magic
tech gf180mcuC
magscale 1 10
timestamp 1694167481
<< nwell >>
rect -3356 -2050 -1223 1494
rect -801 727 1273 1072
rect -801 719 206 727
rect 269 719 1273 727
rect -801 352 1273 719
rect -801 337 -262 352
rect -129 351 1273 352
rect -129 337 596 351
rect -801 333 596 337
rect 734 333 1273 351
rect -3327 -5821 -1192 -2523
rect -801 -3402 1273 333
rect 2328 -2739 4727 1209
rect 2328 -2805 2599 -2739
rect 2677 -2805 4727 -2739
rect 2328 -2977 4727 -2805
rect 5128 -2977 7527 1209
rect 7928 -2977 10327 1209
rect -3327 -5931 -2302 -5821
rect -2291 -5931 -1192 -5821
rect -3327 -6363 -1192 -5931
rect -515 -4375 1318 -4010
rect -515 -4398 -260 -4375
rect -80 -4398 1318 -4375
rect -515 -4553 1318 -4398
rect -515 -4728 -331 -4553
rect -247 -4728 1318 -4553
rect -515 -6334 1318 -4728
rect 1580 -4662 3777 -4275
rect 1580 -4677 2799 -4662
rect 2804 -4677 3777 -4662
rect 1580 -5366 3777 -4677
rect 1580 -5367 2287 -5366
rect 1580 -5443 2071 -5367
rect 2148 -5442 2287 -5367
rect 2364 -5442 3777 -5366
rect 2148 -5443 3777 -5442
rect 1580 -6286 3777 -5443
rect 3985 -6109 6764 -4369
<< pwell >>
rect 8737 -5079 11136 -4680
rect 8737 -5110 9252 -5079
rect 9343 -5080 10204 -5079
rect 9343 -5110 9569 -5080
rect 8737 -5111 9569 -5110
rect 9660 -5111 9886 -5080
rect 9977 -5110 10204 -5080
rect 10295 -5080 11136 -5079
rect 10295 -5110 10536 -5080
rect 9977 -5111 10536 -5110
rect 10627 -5111 11136 -5080
rect -3356 -7177 -1146 -6788
rect -3356 -7348 -2657 -7177
rect -2449 -7348 -1146 -7177
rect -3356 -7994 -1146 -7348
rect -3356 -8131 -1983 -7994
rect -1814 -8131 -1146 -7994
rect -3356 -8780 -1146 -8131
rect -3356 -8919 -1988 -8780
rect -1836 -8919 -1146 -8780
rect -3356 -9589 -1146 -8919
rect -3356 -9741 -2622 -9589
rect -2472 -9741 -1146 -9589
rect -3356 -10473 -1146 -9741
rect -610 -8055 1318 -6466
rect 1570 -7724 4149 -6521
rect 4358 -7533 8117 -6726
rect 4358 -7538 7618 -7533
rect 4358 -7540 7852 -7538
rect 7855 -7540 8117 -7533
rect 4358 -7615 8117 -7540
rect 8737 -7181 11136 -5111
rect 8737 -7183 10209 -7181
rect 8737 -7211 9244 -7183
rect 9343 -7211 9574 -7183
rect 9673 -7211 9887 -7183
rect 9986 -7209 10209 -7183
rect 10308 -7183 11136 -7181
rect 10308 -7209 10522 -7183
rect 9986 -7211 10522 -7209
rect 10621 -7211 11136 -7183
rect 8737 -7573 11136 -7211
rect 4358 -7616 7852 -7615
rect 4358 -7618 7618 -7616
rect 7855 -7618 8117 -7615
rect -610 -8065 389 -8055
rect -610 -8079 287 -8065
rect 292 -8079 389 -8065
rect -610 -8140 389 -8079
rect -610 -8154 284 -8140
rect 292 -8154 389 -8140
rect -610 -8160 389 -8154
rect 395 -8160 1318 -8055
rect -610 -9083 1318 -8160
rect 4358 -8070 8117 -7618
rect 4358 -8079 4610 -8070
rect 4847 -8071 7618 -8070
rect 4844 -8072 7618 -8071
rect 4844 -8074 7852 -8072
rect 7855 -8074 8117 -8070
rect 4844 -8079 8117 -8074
rect 4358 -8149 8117 -8079
rect 4358 -8150 7852 -8149
rect 4358 -8154 7618 -8150
rect 4358 -8155 4610 -8154
rect 4847 -8155 7618 -8154
rect 7855 -8155 8117 -8149
rect -610 -9096 282 -9083
rect 290 -9096 1318 -9083
rect -610 -10718 1318 -9096
rect 1589 -9579 2997 -8253
rect 4358 -9017 8117 -8155
rect 8737 -8079 11136 -7680
rect 8737 -8110 9252 -8079
rect 9343 -8080 10204 -8079
rect 9343 -8110 9569 -8080
rect 8737 -8111 9569 -8110
rect 9660 -8111 9886 -8080
rect 9977 -8110 10204 -8080
rect 10295 -8080 11136 -8079
rect 10295 -8110 10536 -8080
rect 9977 -8111 10536 -8110
rect 10627 -8111 11136 -8080
rect 1589 -9605 1774 -9579
rect 1932 -9605 2997 -9579
rect 1589 -10444 2997 -9605
rect 8737 -10181 11136 -8111
rect 8737 -10183 10209 -10181
rect 8737 -10211 9244 -10183
rect 9343 -10211 9574 -10183
rect 9673 -10211 9887 -10183
rect 9986 -10209 10209 -10183
rect 10308 -10183 11136 -10181
rect 10308 -10209 10522 -10183
rect 9986 -10211 10522 -10209
rect 10621 -10211 11136 -10183
rect 8737 -10573 11136 -10211
<< pdiff >>
rect -2599 -3034 -2531 -2953
rect -2435 -4033 -2373 -3971
<< psubdiff >>
rect 8771 -4734 11101 -4719
rect 8771 -4780 8786 -4734
rect 8832 -4780 8884 -4734
rect 8930 -4780 8982 -4734
rect 9028 -4780 9080 -4734
rect 9126 -4780 9178 -4734
rect 9224 -4780 9276 -4734
rect 9322 -4780 9374 -4734
rect 9420 -4780 9472 -4734
rect 9518 -4780 9570 -4734
rect 9616 -4780 9668 -4734
rect 9714 -4780 9766 -4734
rect 9812 -4780 9864 -4734
rect 9910 -4780 9962 -4734
rect 10008 -4780 10060 -4734
rect 10106 -4780 10158 -4734
rect 10204 -4780 10256 -4734
rect 10302 -4780 10354 -4734
rect 10400 -4780 10452 -4734
rect 10498 -4780 10550 -4734
rect 10596 -4780 10648 -4734
rect 10694 -4780 10746 -4734
rect 10792 -4780 10844 -4734
rect 10890 -4780 10942 -4734
rect 10988 -4780 11040 -4734
rect 11086 -4780 11101 -4734
rect 8771 -4795 11101 -4780
rect 8771 -4832 8847 -4795
rect 8771 -4878 8786 -4832
rect 8832 -4878 8847 -4832
rect 8771 -4930 8847 -4878
rect 8771 -4976 8786 -4930
rect 8832 -4976 8847 -4930
rect 11025 -4832 11101 -4795
rect 11025 -4878 11040 -4832
rect 11086 -4878 11101 -4832
rect 11025 -4930 11101 -4878
rect 8771 -5028 8847 -4976
rect 8771 -5074 8786 -5028
rect 8832 -5074 8847 -5028
rect 8771 -5126 8847 -5074
rect 11025 -4976 11040 -4930
rect 11086 -4976 11101 -4930
rect 11025 -5028 11101 -4976
rect 11025 -5074 11040 -5028
rect 11086 -5074 11101 -5028
rect 8771 -5172 8786 -5126
rect 8832 -5172 8847 -5126
rect 8771 -5224 8847 -5172
rect 8771 -5270 8786 -5224
rect 8832 -5270 8847 -5224
rect 8771 -5322 8847 -5270
rect 8771 -5368 8786 -5322
rect 8832 -5368 8847 -5322
rect 8771 -5420 8847 -5368
rect 8771 -5466 8786 -5420
rect 8832 -5466 8847 -5420
rect 8771 -5518 8847 -5466
rect 8771 -5564 8786 -5518
rect 8832 -5564 8847 -5518
rect 8771 -5616 8847 -5564
rect 8771 -5662 8786 -5616
rect 8832 -5662 8847 -5616
rect 8771 -5714 8847 -5662
rect 8771 -5760 8786 -5714
rect 8832 -5760 8847 -5714
rect 11025 -5126 11101 -5074
rect 11025 -5172 11040 -5126
rect 11086 -5172 11101 -5126
rect 11025 -5224 11101 -5172
rect 11025 -5270 11040 -5224
rect 11086 -5270 11101 -5224
rect 11025 -5322 11101 -5270
rect 11025 -5368 11040 -5322
rect 11086 -5368 11101 -5322
rect 11025 -5420 11101 -5368
rect 11025 -5466 11040 -5420
rect 11086 -5466 11101 -5420
rect 11025 -5518 11101 -5466
rect 11025 -5564 11040 -5518
rect 11086 -5564 11101 -5518
rect 11025 -5616 11101 -5564
rect 11025 -5662 11040 -5616
rect 11086 -5662 11101 -5616
rect 11025 -5714 11101 -5662
rect 8771 -5812 8847 -5760
rect 8771 -5858 8786 -5812
rect 8832 -5858 8847 -5812
rect 11025 -5760 11040 -5714
rect 11086 -5760 11101 -5714
rect 11025 -5812 11101 -5760
rect 8771 -5910 8847 -5858
rect 8771 -5956 8786 -5910
rect 8832 -5956 8847 -5910
rect 8771 -6008 8847 -5956
rect 8771 -6054 8786 -6008
rect 8832 -6054 8847 -6008
rect 8771 -6106 8847 -6054
rect 8771 -6152 8786 -6106
rect 8832 -6152 8847 -6106
rect 8771 -6204 8847 -6152
rect 8771 -6250 8786 -6204
rect 8832 -6250 8847 -6204
rect 8771 -6302 8847 -6250
rect 8771 -6348 8786 -6302
rect 8832 -6348 8847 -6302
rect 8771 -6400 8847 -6348
rect 8771 -6446 8786 -6400
rect 8832 -6446 8847 -6400
rect -564 -6512 1276 -6497
rect -564 -6558 -549 -6512
rect -503 -6558 -451 -6512
rect -405 -6558 -353 -6512
rect -307 -6558 -255 -6512
rect -209 -6558 -157 -6512
rect -111 -6558 -59 -6512
rect -13 -6558 39 -6512
rect 85 -6558 137 -6512
rect 183 -6558 235 -6512
rect 281 -6558 333 -6512
rect 379 -6558 431 -6512
rect 477 -6558 529 -6512
rect 575 -6558 627 -6512
rect 673 -6558 725 -6512
rect 771 -6558 823 -6512
rect 869 -6558 921 -6512
rect 967 -6558 1019 -6512
rect 1065 -6558 1117 -6512
rect 1163 -6558 1215 -6512
rect 1261 -6558 1276 -6512
rect 8771 -6498 8847 -6446
rect 11025 -5858 11040 -5812
rect 11086 -5858 11101 -5812
rect 11025 -5910 11101 -5858
rect 11025 -5956 11040 -5910
rect 11086 -5956 11101 -5910
rect 11025 -6008 11101 -5956
rect 11025 -6054 11040 -6008
rect 11086 -6054 11101 -6008
rect 11025 -6106 11101 -6054
rect 11025 -6152 11040 -6106
rect 11086 -6152 11101 -6106
rect 11025 -6204 11101 -6152
rect 11025 -6250 11040 -6204
rect 11086 -6250 11101 -6204
rect 11025 -6302 11101 -6250
rect 11025 -6348 11040 -6302
rect 11086 -6348 11101 -6302
rect 11025 -6400 11101 -6348
rect 11025 -6446 11040 -6400
rect 11086 -6446 11101 -6400
rect 8771 -6544 8786 -6498
rect 8832 -6544 8847 -6498
rect -564 -6573 1276 -6558
rect -564 -6610 -488 -6573
rect -564 -6656 -549 -6610
rect -503 -6656 -488 -6610
rect -564 -6708 -488 -6656
rect -564 -6754 -549 -6708
rect -503 -6754 -488 -6708
rect -564 -6806 -488 -6754
rect -3310 -6842 -1176 -6827
rect -3310 -6888 -3295 -6842
rect -3249 -6888 -3197 -6842
rect -3151 -6888 -3099 -6842
rect -3053 -6888 -3001 -6842
rect -2955 -6888 -2903 -6842
rect -2857 -6888 -2805 -6842
rect -2759 -6888 -2707 -6842
rect -2661 -6888 -2609 -6842
rect -2563 -6888 -2511 -6842
rect -2465 -6888 -2413 -6842
rect -2367 -6888 -2315 -6842
rect -2269 -6888 -2217 -6842
rect -2171 -6888 -2119 -6842
rect -2073 -6888 -2021 -6842
rect -1975 -6888 -1923 -6842
rect -1877 -6888 -1825 -6842
rect -1779 -6888 -1727 -6842
rect -1681 -6888 -1629 -6842
rect -1583 -6888 -1531 -6842
rect -1485 -6888 -1433 -6842
rect -1387 -6888 -1335 -6842
rect -1289 -6888 -1237 -6842
rect -1191 -6888 -1176 -6842
rect -3310 -6903 -1176 -6888
rect -3310 -6940 -3234 -6903
rect -3310 -6986 -3295 -6940
rect -3249 -6986 -3234 -6940
rect -3310 -7038 -3234 -6986
rect -3310 -7084 -3295 -7038
rect -3249 -7084 -3234 -7038
rect -1252 -6940 -1176 -6903
rect -1252 -6986 -1237 -6940
rect -1191 -6986 -1176 -6940
rect -1252 -7038 -1176 -6986
rect -3310 -7136 -3234 -7084
rect -3310 -7182 -3295 -7136
rect -3249 -7182 -3234 -7136
rect -1252 -7084 -1237 -7038
rect -1191 -7084 -1176 -7038
rect -1252 -7136 -1176 -7084
rect -3310 -7234 -3234 -7182
rect -3310 -7280 -3295 -7234
rect -3249 -7280 -3234 -7234
rect -3310 -7332 -3234 -7280
rect -3310 -7378 -3295 -7332
rect -3249 -7378 -3234 -7332
rect -3310 -7430 -3234 -7378
rect -3310 -7476 -3295 -7430
rect -3249 -7476 -3234 -7430
rect -3310 -7528 -3234 -7476
rect -3310 -7574 -3295 -7528
rect -3249 -7574 -3234 -7528
rect -3310 -7626 -3234 -7574
rect -3310 -7672 -3295 -7626
rect -3249 -7672 -3234 -7626
rect -3310 -7724 -3234 -7672
rect -3310 -7770 -3295 -7724
rect -3249 -7770 -3234 -7724
rect -1252 -7182 -1237 -7136
rect -1191 -7182 -1176 -7136
rect -1252 -7234 -1176 -7182
rect -1252 -7280 -1237 -7234
rect -1191 -7280 -1176 -7234
rect -1252 -7332 -1176 -7280
rect -1252 -7378 -1237 -7332
rect -1191 -7378 -1176 -7332
rect -1252 -7430 -1176 -7378
rect -1252 -7476 -1237 -7430
rect -1191 -7476 -1176 -7430
rect -1252 -7528 -1176 -7476
rect -1252 -7574 -1237 -7528
rect -1191 -7574 -1176 -7528
rect -1252 -7626 -1176 -7574
rect -1252 -7672 -1237 -7626
rect -1191 -7672 -1176 -7626
rect -1252 -7724 -1176 -7672
rect -3310 -7822 -3234 -7770
rect -3310 -7868 -3295 -7822
rect -3249 -7868 -3234 -7822
rect -1252 -7770 -1237 -7724
rect -1191 -7770 -1176 -7724
rect -3310 -7920 -3234 -7868
rect -1252 -7822 -1176 -7770
rect -3310 -7966 -3295 -7920
rect -3249 -7966 -3234 -7920
rect -1252 -7868 -1237 -7822
rect -1191 -7868 -1176 -7822
rect -1252 -7920 -1176 -7868
rect -3310 -8018 -3234 -7966
rect -3310 -8064 -3295 -8018
rect -3249 -8064 -3234 -8018
rect -3310 -8116 -3234 -8064
rect -3310 -8162 -3295 -8116
rect -3249 -8162 -3234 -8116
rect -3310 -8214 -3234 -8162
rect -3310 -8260 -3295 -8214
rect -3249 -8260 -3234 -8214
rect -3310 -8312 -3234 -8260
rect -3310 -8358 -3295 -8312
rect -3249 -8358 -3234 -8312
rect -3310 -8410 -3234 -8358
rect -3310 -8456 -3295 -8410
rect -3249 -8456 -3234 -8410
rect -3310 -8508 -3234 -8456
rect -3310 -8554 -3295 -8508
rect -3249 -8554 -3234 -8508
rect -1252 -7966 -1237 -7920
rect -1191 -7966 -1176 -7920
rect -1252 -8018 -1176 -7966
rect -1252 -8064 -1237 -8018
rect -1191 -8064 -1176 -8018
rect -1252 -8116 -1176 -8064
rect -1252 -8162 -1237 -8116
rect -1191 -8162 -1176 -8116
rect -1252 -8214 -1176 -8162
rect -1252 -8260 -1237 -8214
rect -1191 -8260 -1176 -8214
rect -1252 -8312 -1176 -8260
rect -1252 -8358 -1237 -8312
rect -1191 -8358 -1176 -8312
rect -1252 -8410 -1176 -8358
rect -1252 -8456 -1237 -8410
rect -1191 -8456 -1176 -8410
rect -1252 -8508 -1176 -8456
rect -3310 -8606 -3234 -8554
rect -3310 -8652 -3295 -8606
rect -3249 -8652 -3234 -8606
rect -1252 -8554 -1237 -8508
rect -1191 -8554 -1176 -8508
rect -3310 -8704 -3234 -8652
rect -3310 -8750 -3295 -8704
rect -3249 -8750 -3234 -8704
rect -1252 -8606 -1176 -8554
rect -1252 -8652 -1237 -8606
rect -1191 -8652 -1176 -8606
rect -1252 -8704 -1176 -8652
rect -3310 -8802 -3234 -8750
rect -3310 -8848 -3295 -8802
rect -3249 -8848 -3234 -8802
rect -3310 -8900 -3234 -8848
rect -3310 -8946 -3295 -8900
rect -3249 -8946 -3234 -8900
rect -3310 -8998 -3234 -8946
rect -3310 -9044 -3295 -8998
rect -3249 -9044 -3234 -8998
rect -3310 -9096 -3234 -9044
rect -3310 -9142 -3295 -9096
rect -3249 -9142 -3234 -9096
rect -3310 -9194 -3234 -9142
rect -3310 -9240 -3295 -9194
rect -3249 -9240 -3234 -9194
rect -3310 -9292 -3234 -9240
rect -3310 -9338 -3295 -9292
rect -3249 -9338 -3234 -9292
rect -1252 -8750 -1237 -8704
rect -1191 -8750 -1176 -8704
rect -1252 -8802 -1176 -8750
rect -1252 -8848 -1237 -8802
rect -1191 -8848 -1176 -8802
rect -1252 -8900 -1176 -8848
rect -1252 -8946 -1237 -8900
rect -1191 -8946 -1176 -8900
rect -1252 -8998 -1176 -8946
rect -1252 -9044 -1237 -8998
rect -1191 -9044 -1176 -8998
rect -1252 -9096 -1176 -9044
rect -1252 -9142 -1237 -9096
rect -1191 -9142 -1176 -9096
rect -1252 -9194 -1176 -9142
rect -1252 -9240 -1237 -9194
rect -1191 -9240 -1176 -9194
rect -1252 -9292 -1176 -9240
rect -3310 -9390 -3234 -9338
rect -3310 -9436 -3295 -9390
rect -3249 -9436 -3234 -9390
rect -3310 -9488 -3234 -9436
rect -1252 -9338 -1237 -9292
rect -1191 -9338 -1176 -9292
rect -3310 -9534 -3295 -9488
rect -3249 -9534 -3234 -9488
rect -3310 -9586 -3234 -9534
rect -1252 -9390 -1176 -9338
rect -1252 -9436 -1237 -9390
rect -1191 -9436 -1176 -9390
rect -1252 -9488 -1176 -9436
rect -1252 -9534 -1237 -9488
rect -1191 -9534 -1176 -9488
rect -3310 -9632 -3295 -9586
rect -3249 -9632 -3234 -9586
rect -3310 -9684 -3234 -9632
rect -3310 -9730 -3295 -9684
rect -3249 -9730 -3234 -9684
rect -3310 -9782 -3234 -9730
rect -3310 -9828 -3295 -9782
rect -3249 -9828 -3234 -9782
rect -3310 -9880 -3234 -9828
rect -3310 -9926 -3295 -9880
rect -3249 -9926 -3234 -9880
rect -3310 -9978 -3234 -9926
rect -3310 -10024 -3295 -9978
rect -3249 -10024 -3234 -9978
rect -3310 -10076 -3234 -10024
rect -3310 -10122 -3295 -10076
rect -3249 -10122 -3234 -10076
rect -3310 -10174 -3234 -10122
rect -1252 -9586 -1176 -9534
rect -1252 -9632 -1237 -9586
rect -1191 -9632 -1176 -9586
rect -1252 -9684 -1176 -9632
rect -1252 -9730 -1237 -9684
rect -1191 -9730 -1176 -9684
rect -1252 -9782 -1176 -9730
rect -1252 -9828 -1237 -9782
rect -1191 -9828 -1176 -9782
rect -1252 -9880 -1176 -9828
rect -1252 -9926 -1237 -9880
rect -1191 -9926 -1176 -9880
rect -1252 -9978 -1176 -9926
rect -1252 -10024 -1237 -9978
rect -1191 -10024 -1176 -9978
rect -1252 -10076 -1176 -10024
rect -1252 -10122 -1237 -10076
rect -1191 -10122 -1176 -10076
rect -3310 -10220 -3295 -10174
rect -3249 -10220 -3234 -10174
rect -1252 -10174 -1176 -10122
rect -3310 -10272 -3234 -10220
rect -3310 -10318 -3295 -10272
rect -3249 -10318 -3234 -10272
rect -3310 -10355 -3234 -10318
rect -1252 -10220 -1237 -10174
rect -1191 -10220 -1176 -10174
rect -1252 -10272 -1176 -10220
rect -1252 -10318 -1237 -10272
rect -1191 -10318 -1176 -10272
rect -1252 -10355 -1176 -10318
rect -3310 -10370 -1176 -10355
rect -3310 -10416 -3295 -10370
rect -3249 -10416 -3197 -10370
rect -3151 -10416 -3099 -10370
rect -3053 -10416 -3001 -10370
rect -2955 -10416 -2903 -10370
rect -2857 -10416 -2805 -10370
rect -2759 -10416 -2707 -10370
rect -2661 -10416 -2609 -10370
rect -2563 -10416 -2511 -10370
rect -2465 -10416 -2413 -10370
rect -2367 -10416 -2315 -10370
rect -2269 -10416 -2217 -10370
rect -2171 -10416 -2119 -10370
rect -2073 -10416 -2021 -10370
rect -1975 -10416 -1923 -10370
rect -1877 -10416 -1825 -10370
rect -1779 -10416 -1727 -10370
rect -1681 -10416 -1629 -10370
rect -1583 -10416 -1531 -10370
rect -1485 -10416 -1433 -10370
rect -1387 -10416 -1335 -10370
rect -1289 -10416 -1237 -10370
rect -1191 -10416 -1176 -10370
rect -3310 -10431 -1176 -10416
rect -564 -6852 -549 -6806
rect -503 -6852 -488 -6806
rect 1200 -6610 1276 -6573
rect 1200 -6656 1215 -6610
rect 1261 -6656 1276 -6610
rect 1200 -6708 1276 -6656
rect 1200 -6754 1215 -6708
rect 1261 -6754 1276 -6708
rect 1200 -6806 1276 -6754
rect -564 -6904 -488 -6852
rect -564 -6950 -549 -6904
rect -503 -6950 -488 -6904
rect 1200 -6852 1215 -6806
rect 1261 -6852 1276 -6806
rect 1200 -6904 1276 -6852
rect -564 -7002 -488 -6950
rect -564 -7048 -549 -7002
rect -503 -7048 -488 -7002
rect -564 -7100 -488 -7048
rect -564 -7146 -549 -7100
rect -503 -7146 -488 -7100
rect -564 -7198 -488 -7146
rect -564 -7244 -549 -7198
rect -503 -7244 -488 -7198
rect -564 -7296 -488 -7244
rect -564 -7342 -549 -7296
rect -503 -7342 -488 -7296
rect -564 -7394 -488 -7342
rect -564 -7440 -549 -7394
rect -503 -7440 -488 -7394
rect -564 -7492 -488 -7440
rect -564 -7538 -549 -7492
rect -503 -7538 -488 -7492
rect -564 -7590 -488 -7538
rect -564 -7636 -549 -7590
rect -503 -7636 -488 -7590
rect 1200 -6950 1215 -6904
rect 1261 -6950 1276 -6904
rect 1200 -7002 1276 -6950
rect 1200 -7048 1215 -7002
rect 1261 -7048 1276 -7002
rect 1200 -7100 1276 -7048
rect 1200 -7146 1215 -7100
rect 1261 -7146 1276 -7100
rect 1200 -7198 1276 -7146
rect 1200 -7244 1215 -7198
rect 1261 -7244 1276 -7198
rect 1200 -7296 1276 -7244
rect 1200 -7342 1215 -7296
rect 1261 -7342 1276 -7296
rect 1200 -7394 1276 -7342
rect 1200 -7440 1215 -7394
rect 1261 -7440 1276 -7394
rect 1200 -7492 1276 -7440
rect 1200 -7538 1215 -7492
rect 1261 -7538 1276 -7492
rect 1200 -7590 1276 -7538
rect -564 -7688 -488 -7636
rect -564 -7734 -549 -7688
rect -503 -7734 -488 -7688
rect -564 -7786 -488 -7734
rect -564 -7832 -549 -7786
rect -503 -7832 -488 -7786
rect 1200 -7636 1215 -7590
rect 1261 -7636 1276 -7590
rect 1200 -7688 1276 -7636
rect 1200 -7734 1215 -7688
rect 1261 -7734 1276 -7688
rect 1597 -6562 4123 -6547
rect 1597 -6608 1612 -6562
rect 1658 -6608 1710 -6562
rect 1756 -6608 1808 -6562
rect 1854 -6608 1906 -6562
rect 1952 -6608 2004 -6562
rect 2050 -6608 2102 -6562
rect 2148 -6608 2200 -6562
rect 2246 -6608 2298 -6562
rect 2344 -6608 2396 -6562
rect 2442 -6608 2494 -6562
rect 2540 -6608 2592 -6562
rect 2638 -6608 2690 -6562
rect 2736 -6608 2788 -6562
rect 2834 -6608 2886 -6562
rect 2932 -6608 2984 -6562
rect 3030 -6608 3082 -6562
rect 3128 -6608 3180 -6562
rect 3226 -6608 3278 -6562
rect 3324 -6608 3376 -6562
rect 3422 -6608 3474 -6562
rect 3520 -6608 3572 -6562
rect 3618 -6608 3670 -6562
rect 3716 -6608 3768 -6562
rect 3814 -6608 3866 -6562
rect 3912 -6608 3964 -6562
rect 4010 -6608 4062 -6562
rect 4108 -6608 4123 -6562
rect 1597 -6623 4123 -6608
rect 1597 -6660 1673 -6623
rect 1597 -6706 1612 -6660
rect 1658 -6706 1673 -6660
rect 1597 -6756 1673 -6706
rect 4047 -6660 4123 -6623
rect 4047 -6706 4062 -6660
rect 4108 -6706 4123 -6660
rect 1597 -6802 1612 -6756
rect 1658 -6802 1673 -6756
rect 1597 -6854 1673 -6802
rect 1597 -6900 1612 -6854
rect 1658 -6900 1673 -6854
rect 4047 -6756 4123 -6706
rect 8771 -6596 8847 -6544
rect 11025 -6498 11101 -6446
rect 11025 -6544 11040 -6498
rect 11086 -6544 11101 -6498
rect 8771 -6642 8786 -6596
rect 8832 -6642 8847 -6596
rect 8771 -6694 8847 -6642
rect 8771 -6740 8786 -6694
rect 8832 -6740 8847 -6694
rect 4047 -6802 4062 -6756
rect 4108 -6802 4123 -6756
rect 4047 -6854 4123 -6802
rect 1597 -6952 1673 -6900
rect 4047 -6900 4062 -6854
rect 4108 -6900 4123 -6854
rect 1597 -6998 1612 -6952
rect 1658 -6998 1673 -6952
rect 1597 -7050 1673 -6998
rect 1597 -7096 1612 -7050
rect 1658 -7096 1673 -7050
rect 1597 -7148 1673 -7096
rect 1597 -7194 1612 -7148
rect 1658 -7194 1673 -7148
rect 1597 -7246 1673 -7194
rect 1597 -7292 1612 -7246
rect 1658 -7292 1673 -7246
rect 1597 -7344 1673 -7292
rect 4047 -6952 4123 -6900
rect 4047 -6998 4062 -6952
rect 4108 -6998 4123 -6952
rect 4047 -7050 4123 -6998
rect 4047 -7096 4062 -7050
rect 4108 -7096 4123 -7050
rect 4047 -7148 4123 -7096
rect 4047 -7194 4062 -7148
rect 4108 -7194 4123 -7148
rect 4047 -7246 4123 -7194
rect 4047 -7292 4062 -7246
rect 4108 -7292 4123 -7246
rect 1597 -7390 1612 -7344
rect 1658 -7390 1673 -7344
rect 1597 -7442 1673 -7390
rect 1597 -7488 1612 -7442
rect 1658 -7488 1673 -7442
rect 1597 -7540 1673 -7488
rect 4047 -7344 4123 -7292
rect 4047 -7390 4062 -7344
rect 4108 -7390 4123 -7344
rect 4047 -7442 4123 -7390
rect 4047 -7488 4062 -7442
rect 4108 -7488 4123 -7442
rect 1597 -7586 1612 -7540
rect 1658 -7586 1673 -7540
rect 1597 -7623 1673 -7586
rect 4047 -7540 4123 -7488
rect 4047 -7586 4062 -7540
rect 4108 -7586 4123 -7540
rect 4047 -7623 4123 -7586
rect 1597 -7638 4123 -7623
rect 1597 -7684 1612 -7638
rect 1658 -7684 1710 -7638
rect 1756 -7684 1808 -7638
rect 1854 -7684 1906 -7638
rect 1952 -7684 2004 -7638
rect 2050 -7684 2102 -7638
rect 2148 -7684 2200 -7638
rect 2246 -7684 2298 -7638
rect 2344 -7684 2396 -7638
rect 2442 -7684 2494 -7638
rect 2540 -7684 2592 -7638
rect 2638 -7684 2690 -7638
rect 2736 -7684 2788 -7638
rect 2834 -7684 2886 -7638
rect 2932 -7684 2984 -7638
rect 3030 -7684 3082 -7638
rect 3128 -7684 3180 -7638
rect 3226 -7684 3278 -7638
rect 3324 -7684 3376 -7638
rect 3422 -7684 3474 -7638
rect 3520 -7684 3572 -7638
rect 3618 -7684 3670 -7638
rect 3716 -7684 3768 -7638
rect 3814 -7684 3866 -7638
rect 3912 -7684 3964 -7638
rect 4010 -7684 4062 -7638
rect 4108 -7684 4123 -7638
rect 1597 -7699 4123 -7684
rect 4385 -6765 8087 -6750
rect 4385 -6766 4497 -6765
rect 4385 -6812 4399 -6766
rect 4445 -6811 4497 -6766
rect 4543 -6811 4595 -6765
rect 4641 -6811 4693 -6765
rect 4739 -6811 4791 -6765
rect 4837 -6811 4889 -6765
rect 4935 -6811 4987 -6765
rect 5033 -6811 5085 -6765
rect 5131 -6811 5183 -6765
rect 5229 -6811 5281 -6765
rect 5327 -6811 5379 -6765
rect 5425 -6811 5477 -6765
rect 5523 -6811 5575 -6765
rect 5621 -6811 5673 -6765
rect 5719 -6811 5771 -6765
rect 5817 -6811 5869 -6765
rect 5915 -6811 5967 -6765
rect 6013 -6811 6065 -6765
rect 6111 -6811 6163 -6765
rect 6209 -6811 6261 -6765
rect 6307 -6811 6359 -6765
rect 6405 -6811 6457 -6765
rect 6503 -6811 6555 -6765
rect 6601 -6811 6653 -6765
rect 6699 -6811 6751 -6765
rect 6797 -6811 6849 -6765
rect 6895 -6811 6947 -6765
rect 6993 -6811 7045 -6765
rect 7091 -6811 7143 -6765
rect 7189 -6811 7241 -6765
rect 7287 -6811 7339 -6765
rect 7385 -6811 7437 -6765
rect 7483 -6811 7535 -6765
rect 7581 -6811 7633 -6765
rect 7679 -6811 7731 -6765
rect 7777 -6811 7829 -6765
rect 7875 -6811 7927 -6765
rect 7973 -6811 8025 -6765
rect 8071 -6811 8087 -6765
rect 4445 -6812 8087 -6811
rect 4385 -6826 8087 -6812
rect 4385 -6863 4461 -6826
rect 4385 -6909 4400 -6863
rect 4446 -6909 4461 -6863
rect 8011 -6864 8087 -6826
rect 4385 -6961 4461 -6909
rect 4385 -7007 4400 -6961
rect 4446 -7007 4461 -6961
rect 4385 -7059 4461 -7007
rect 4385 -7105 4400 -7059
rect 4446 -7105 4461 -7059
rect 8011 -6910 8026 -6864
rect 8072 -6910 8087 -6864
rect 8011 -6962 8087 -6910
rect 8011 -7008 8026 -6962
rect 8072 -7008 8087 -6962
rect 8011 -7060 8087 -7008
rect 4385 -7157 4461 -7105
rect 4385 -7203 4400 -7157
rect 4446 -7203 4461 -7157
rect 4385 -7255 4461 -7203
rect 4385 -7301 4400 -7255
rect 4446 -7301 4461 -7255
rect 4385 -7353 4461 -7301
rect 4385 -7399 4400 -7353
rect 4446 -7399 4461 -7353
rect 4385 -7451 4461 -7399
rect 4385 -7497 4400 -7451
rect 4446 -7497 4461 -7451
rect 4385 -7549 4461 -7497
rect 8011 -7106 8026 -7060
rect 8072 -7106 8087 -7060
rect 8011 -7158 8087 -7106
rect 8011 -7204 8026 -7158
rect 8072 -7204 8087 -7158
rect 8011 -7256 8087 -7204
rect 8011 -7302 8026 -7256
rect 8072 -7302 8087 -7256
rect 8011 -7354 8087 -7302
rect 8011 -7400 8026 -7354
rect 8072 -7400 8087 -7354
rect 8011 -7452 8087 -7400
rect 8011 -7498 8026 -7452
rect 8072 -7498 8087 -7452
rect 4385 -7595 4400 -7549
rect 4446 -7595 4461 -7549
rect 4385 -7647 4461 -7595
rect 8011 -7550 8087 -7498
rect 8771 -6792 8847 -6740
rect 8771 -6838 8786 -6792
rect 8832 -6838 8847 -6792
rect 8771 -6890 8847 -6838
rect 8771 -6936 8786 -6890
rect 8832 -6936 8847 -6890
rect 8771 -6988 8847 -6936
rect 8771 -7034 8786 -6988
rect 8832 -7034 8847 -6988
rect 8771 -7086 8847 -7034
rect 8771 -7132 8786 -7086
rect 8832 -7132 8847 -7086
rect 8771 -7184 8847 -7132
rect 8771 -7230 8786 -7184
rect 8832 -7230 8847 -7184
rect 11025 -6596 11101 -6544
rect 11025 -6642 11040 -6596
rect 11086 -6642 11101 -6596
rect 11025 -6694 11101 -6642
rect 11025 -6740 11040 -6694
rect 11086 -6740 11101 -6694
rect 11025 -6792 11101 -6740
rect 11025 -6838 11040 -6792
rect 11086 -6838 11101 -6792
rect 11025 -6890 11101 -6838
rect 11025 -6936 11040 -6890
rect 11086 -6936 11101 -6890
rect 11025 -6988 11101 -6936
rect 11025 -7034 11040 -6988
rect 11086 -7034 11101 -6988
rect 11025 -7086 11101 -7034
rect 11025 -7132 11040 -7086
rect 11086 -7132 11101 -7086
rect 11025 -7184 11101 -7132
rect 8771 -7282 8847 -7230
rect 8771 -7328 8786 -7282
rect 8832 -7328 8847 -7282
rect 8771 -7380 8847 -7328
rect 11025 -7230 11040 -7184
rect 11086 -7230 11101 -7184
rect 11025 -7282 11101 -7230
rect 11025 -7328 11040 -7282
rect 11086 -7328 11101 -7282
rect 8771 -7426 8786 -7380
rect 8832 -7426 8847 -7380
rect 8771 -7463 8847 -7426
rect 11025 -7380 11101 -7328
rect 11025 -7426 11040 -7380
rect 11086 -7426 11101 -7380
rect 11025 -7463 11101 -7426
rect 8771 -7478 11101 -7463
rect 8771 -7524 8786 -7478
rect 8832 -7524 8884 -7478
rect 8930 -7524 8982 -7478
rect 9028 -7524 9080 -7478
rect 9126 -7524 9178 -7478
rect 9224 -7524 9276 -7478
rect 9322 -7524 9374 -7478
rect 9420 -7524 9472 -7478
rect 9518 -7524 9570 -7478
rect 9616 -7524 9668 -7478
rect 9714 -7524 9766 -7478
rect 9812 -7524 9864 -7478
rect 9910 -7524 9962 -7478
rect 10008 -7524 10060 -7478
rect 10106 -7524 10158 -7478
rect 10204 -7524 10256 -7478
rect 10302 -7524 10354 -7478
rect 10400 -7524 10452 -7478
rect 10498 -7524 10550 -7478
rect 10596 -7524 10648 -7478
rect 10694 -7524 10746 -7478
rect 10792 -7524 10844 -7478
rect 10890 -7524 10942 -7478
rect 10988 -7524 11040 -7478
rect 11086 -7524 11101 -7478
rect 8771 -7539 11101 -7524
rect 8011 -7596 8026 -7550
rect 8072 -7596 8087 -7550
rect 4385 -7693 4400 -7647
rect 4446 -7693 4461 -7647
rect 1200 -7786 1276 -7734
rect -564 -7884 -488 -7832
rect -564 -7930 -549 -7884
rect -503 -7930 -488 -7884
rect -564 -7982 -488 -7930
rect -564 -8028 -549 -7982
rect -503 -8028 -488 -7982
rect -564 -8080 -488 -8028
rect -564 -8126 -549 -8080
rect -503 -8126 -488 -8080
rect -564 -8178 -488 -8126
rect -564 -8224 -549 -8178
rect -503 -8224 -488 -8178
rect -564 -8276 -488 -8224
rect -564 -8322 -549 -8276
rect -503 -8322 -488 -8276
rect -564 -8374 -488 -8322
rect -564 -8420 -549 -8374
rect -503 -8420 -488 -8374
rect -564 -8472 -488 -8420
rect -564 -8518 -549 -8472
rect -503 -8518 -488 -8472
rect 1200 -7832 1215 -7786
rect 1261 -7832 1276 -7786
rect 1200 -7884 1276 -7832
rect 1200 -7930 1215 -7884
rect 1261 -7930 1276 -7884
rect 1200 -7982 1276 -7930
rect 1200 -8028 1215 -7982
rect 1261 -8028 1276 -7982
rect 1200 -8080 1276 -8028
rect 1200 -8126 1215 -8080
rect 1261 -8126 1276 -8080
rect 1200 -8178 1276 -8126
rect 1200 -8224 1215 -8178
rect 1261 -8224 1276 -8178
rect 1200 -8276 1276 -8224
rect 1200 -8322 1215 -8276
rect 1261 -8322 1276 -8276
rect 4385 -7745 4461 -7693
rect 4385 -7791 4400 -7745
rect 4446 -7791 4461 -7745
rect 4385 -7843 4461 -7791
rect 4385 -7889 4400 -7843
rect 4446 -7889 4461 -7843
rect 4385 -7941 4461 -7889
rect 4385 -7987 4400 -7941
rect 4446 -7987 4461 -7941
rect 4385 -8039 4461 -7987
rect 4385 -8085 4400 -8039
rect 4446 -8085 4461 -8039
rect 8011 -7648 8087 -7596
rect 8011 -7694 8026 -7648
rect 8072 -7694 8087 -7648
rect 8011 -7746 8087 -7694
rect 8011 -7792 8026 -7746
rect 8072 -7792 8087 -7746
rect 8011 -7844 8087 -7792
rect 8011 -7890 8026 -7844
rect 8072 -7890 8087 -7844
rect 8011 -7942 8087 -7890
rect 8011 -7988 8026 -7942
rect 8072 -7988 8087 -7942
rect 8011 -8040 8087 -7988
rect 4385 -8137 4461 -8085
rect 4385 -8183 4400 -8137
rect 4446 -8183 4461 -8137
rect 8011 -8086 8026 -8040
rect 8072 -8086 8087 -8040
rect 8011 -8138 8087 -8086
rect 4385 -8235 4461 -8183
rect 4385 -8281 4400 -8235
rect 4446 -8281 4461 -8235
rect 2858 -8282 2971 -8281
rect 1200 -8374 1276 -8322
rect 1200 -8420 1215 -8374
rect 1261 -8420 1276 -8374
rect 1200 -8472 1276 -8420
rect -564 -8570 -488 -8518
rect -564 -8616 -549 -8570
rect -503 -8616 -488 -8570
rect -564 -8668 -488 -8616
rect -564 -8714 -549 -8668
rect -503 -8714 -488 -8668
rect -564 -8766 -488 -8714
rect -564 -8812 -549 -8766
rect -503 -8812 -488 -8766
rect 1200 -8518 1215 -8472
rect 1261 -8518 1276 -8472
rect 1200 -8570 1276 -8518
rect 1200 -8616 1215 -8570
rect 1261 -8616 1276 -8570
rect 1200 -8668 1276 -8616
rect 1200 -8714 1215 -8668
rect 1261 -8714 1276 -8668
rect 1200 -8766 1276 -8714
rect -564 -8864 -488 -8812
rect -564 -8910 -549 -8864
rect -503 -8910 -488 -8864
rect -564 -8962 -488 -8910
rect -564 -9008 -549 -8962
rect -503 -9008 -488 -8962
rect -564 -9060 -488 -9008
rect -564 -9106 -549 -9060
rect -503 -9106 -488 -9060
rect -564 -9158 -488 -9106
rect -564 -9204 -549 -9158
rect -503 -9204 -488 -9158
rect -564 -9256 -488 -9204
rect -564 -9302 -549 -9256
rect -503 -9302 -488 -9256
rect -564 -9354 -488 -9302
rect -564 -9400 -549 -9354
rect -503 -9400 -488 -9354
rect -564 -9452 -488 -9400
rect -564 -9498 -549 -9452
rect -503 -9498 -488 -9452
rect 1200 -8812 1215 -8766
rect 1261 -8812 1276 -8766
rect 1200 -8864 1276 -8812
rect 1200 -8910 1215 -8864
rect 1261 -8910 1276 -8864
rect 1200 -8962 1276 -8910
rect 1200 -9008 1215 -8962
rect 1261 -9008 1276 -8962
rect 1200 -9060 1276 -9008
rect 1200 -9106 1215 -9060
rect 1261 -9106 1276 -9060
rect 1200 -9158 1276 -9106
rect 1200 -9204 1215 -9158
rect 1261 -9204 1276 -9158
rect 1200 -9256 1276 -9204
rect 1200 -9302 1215 -9256
rect 1261 -9302 1276 -9256
rect 1200 -9354 1276 -9302
rect 1200 -9400 1215 -9354
rect 1261 -9400 1276 -9354
rect 1200 -9452 1276 -9400
rect -564 -9550 -488 -9498
rect -564 -9596 -549 -9550
rect -503 -9596 -488 -9550
rect -564 -9648 -488 -9596
rect 1200 -9498 1215 -9452
rect 1261 -9498 1276 -9452
rect 1200 -9550 1276 -9498
rect 1200 -9596 1215 -9550
rect 1261 -9596 1276 -9550
rect -564 -9694 -549 -9648
rect -503 -9694 -488 -9648
rect -564 -9746 -488 -9694
rect -564 -9792 -549 -9746
rect -503 -9792 -488 -9746
rect -564 -9844 -488 -9792
rect -564 -9890 -549 -9844
rect -503 -9890 -488 -9844
rect -564 -9942 -488 -9890
rect -564 -9988 -549 -9942
rect -503 -9988 -488 -9942
rect -564 -10040 -488 -9988
rect -564 -10086 -549 -10040
rect -503 -10086 -488 -10040
rect -564 -10138 -488 -10086
rect -564 -10184 -549 -10138
rect -503 -10184 -488 -10138
rect -564 -10236 -488 -10184
rect -564 -10282 -549 -10236
rect -503 -10282 -488 -10236
rect -564 -10334 -488 -10282
rect 1200 -9648 1276 -9596
rect 1200 -9694 1215 -9648
rect 1261 -9694 1276 -9648
rect 1200 -9746 1276 -9694
rect 1200 -9792 1215 -9746
rect 1261 -9792 1276 -9746
rect 1200 -9844 1276 -9792
rect 1200 -9890 1215 -9844
rect 1261 -9890 1276 -9844
rect 1200 -9942 1276 -9890
rect 1200 -9988 1215 -9942
rect 1261 -9988 1276 -9942
rect 1200 -10040 1276 -9988
rect 1200 -10086 1215 -10040
rect 1261 -10086 1276 -10040
rect 1200 -10138 1276 -10086
rect 1200 -10184 1215 -10138
rect 1261 -10184 1276 -10138
rect 1200 -10236 1276 -10184
rect 1200 -10282 1215 -10236
rect 1261 -10282 1276 -10236
rect -564 -10380 -549 -10334
rect -503 -10380 -488 -10334
rect -564 -10432 -488 -10380
rect 1200 -10334 1276 -10282
rect 1200 -10380 1215 -10334
rect 1261 -10380 1276 -10334
rect -564 -10478 -549 -10432
rect -503 -10478 -488 -10432
rect -564 -10530 -488 -10478
rect -564 -10576 -549 -10530
rect -503 -10576 -488 -10530
rect -564 -10613 -488 -10576
rect 1200 -10432 1276 -10380
rect 1621 -8296 2971 -8282
rect 1621 -8342 1636 -8296
rect 1682 -8297 2910 -8296
rect 1682 -8342 1734 -8297
rect 1621 -8343 1734 -8342
rect 1780 -8343 1832 -8297
rect 1878 -8343 1930 -8297
rect 1976 -8343 2028 -8297
rect 2074 -8343 2126 -8297
rect 2172 -8343 2224 -8297
rect 2270 -8343 2322 -8297
rect 2368 -8343 2420 -8297
rect 2466 -8343 2518 -8297
rect 2564 -8343 2616 -8297
rect 2662 -8343 2714 -8297
rect 2760 -8343 2812 -8297
rect 2858 -8342 2910 -8297
rect 2956 -8342 2971 -8296
rect 2858 -8343 2971 -8342
rect 1621 -8358 2971 -8343
rect 1621 -8394 1697 -8358
rect 1621 -8440 1636 -8394
rect 1682 -8440 1697 -8394
rect 1621 -8492 1697 -8440
rect 1621 -8538 1636 -8492
rect 1682 -8538 1697 -8492
rect 1621 -8590 1697 -8538
rect 1621 -8636 1636 -8590
rect 1682 -8636 1697 -8590
rect 1621 -8688 1697 -8636
rect 1621 -8734 1636 -8688
rect 1682 -8734 1697 -8688
rect 1621 -8786 1697 -8734
rect 1621 -8832 1636 -8786
rect 1682 -8832 1697 -8786
rect 1621 -8884 1697 -8832
rect 1621 -8930 1636 -8884
rect 1682 -8930 1697 -8884
rect 1621 -8982 1697 -8930
rect 1621 -9028 1636 -8982
rect 1682 -9028 1697 -8982
rect 1621 -9080 1697 -9028
rect 1621 -9126 1636 -9080
rect 1682 -9126 1697 -9080
rect 1621 -9178 1697 -9126
rect 2895 -8394 2971 -8358
rect 2895 -8440 2910 -8394
rect 2956 -8440 2971 -8394
rect 2895 -8492 2971 -8440
rect 2895 -8538 2910 -8492
rect 2956 -8538 2971 -8492
rect 2895 -8590 2971 -8538
rect 2895 -8636 2910 -8590
rect 2956 -8636 2971 -8590
rect 2895 -8688 2971 -8636
rect 2895 -8734 2910 -8688
rect 2956 -8734 2971 -8688
rect 2895 -8786 2971 -8734
rect 2895 -8832 2910 -8786
rect 2956 -8832 2971 -8786
rect 2895 -8884 2971 -8832
rect 2895 -8930 2910 -8884
rect 2956 -8930 2971 -8884
rect 2895 -8982 2971 -8930
rect 2895 -9028 2910 -8982
rect 2956 -9028 2971 -8982
rect 4385 -8333 4461 -8281
rect 4385 -8379 4400 -8333
rect 4446 -8379 4461 -8333
rect 4385 -8431 4461 -8379
rect 4385 -8477 4400 -8431
rect 4446 -8477 4461 -8431
rect 4385 -8529 4461 -8477
rect 4385 -8575 4400 -8529
rect 4446 -8575 4461 -8529
rect 4385 -8627 4461 -8575
rect 8011 -8184 8026 -8138
rect 8072 -8184 8087 -8138
rect 8011 -8236 8087 -8184
rect 8011 -8282 8026 -8236
rect 8072 -8282 8087 -8236
rect 8011 -8334 8087 -8282
rect 8011 -8380 8026 -8334
rect 8072 -8380 8087 -8334
rect 8011 -8432 8087 -8380
rect 8011 -8478 8026 -8432
rect 8072 -8478 8087 -8432
rect 8011 -8530 8087 -8478
rect 8011 -8576 8026 -8530
rect 8072 -8576 8087 -8530
rect 4385 -8673 4400 -8627
rect 4446 -8673 4461 -8627
rect 4385 -8725 4461 -8673
rect 4385 -8771 4400 -8725
rect 4446 -8771 4461 -8725
rect 4385 -8823 4461 -8771
rect 8011 -8628 8087 -8576
rect 8011 -8674 8026 -8628
rect 8072 -8674 8087 -8628
rect 8011 -8726 8087 -8674
rect 8011 -8772 8026 -8726
rect 8072 -8772 8087 -8726
rect 4385 -8869 4400 -8823
rect 4446 -8869 4461 -8823
rect 4385 -8907 4461 -8869
rect 8011 -8824 8087 -8772
rect 8011 -8870 8026 -8824
rect 8072 -8870 8087 -8824
rect 8011 -8907 8087 -8870
rect 4385 -8921 8087 -8907
rect 4385 -8967 4399 -8921
rect 4445 -8922 8087 -8921
rect 4445 -8967 4497 -8922
rect 4385 -8968 4497 -8967
rect 4543 -8968 4595 -8922
rect 4641 -8968 4693 -8922
rect 4739 -8968 4791 -8922
rect 4837 -8968 4889 -8922
rect 4935 -8968 4987 -8922
rect 5033 -8968 5085 -8922
rect 5131 -8968 5183 -8922
rect 5229 -8968 5281 -8922
rect 5327 -8968 5379 -8922
rect 5425 -8968 5477 -8922
rect 5523 -8968 5575 -8922
rect 5621 -8968 5673 -8922
rect 5719 -8968 5771 -8922
rect 5817 -8968 5869 -8922
rect 5915 -8968 5967 -8922
rect 6013 -8968 6065 -8922
rect 6111 -8968 6163 -8922
rect 6209 -8968 6261 -8922
rect 6307 -8968 6359 -8922
rect 6405 -8968 6457 -8922
rect 6503 -8968 6555 -8922
rect 6601 -8968 6653 -8922
rect 6699 -8968 6751 -8922
rect 6797 -8968 6849 -8922
rect 6895 -8968 6947 -8922
rect 6993 -8968 7045 -8922
rect 7091 -8968 7143 -8922
rect 7189 -8968 7241 -8922
rect 7287 -8968 7339 -8922
rect 7385 -8968 7437 -8922
rect 7483 -8968 7535 -8922
rect 7581 -8968 7633 -8922
rect 7679 -8968 7731 -8922
rect 7777 -8968 7829 -8922
rect 7875 -8968 7927 -8922
rect 7973 -8968 8025 -8922
rect 8071 -8968 8087 -8922
rect 4385 -8983 8087 -8968
rect 8771 -7734 11101 -7719
rect 8771 -7780 8786 -7734
rect 8832 -7780 8884 -7734
rect 8930 -7780 8982 -7734
rect 9028 -7780 9080 -7734
rect 9126 -7780 9178 -7734
rect 9224 -7780 9276 -7734
rect 9322 -7780 9374 -7734
rect 9420 -7780 9472 -7734
rect 9518 -7780 9570 -7734
rect 9616 -7780 9668 -7734
rect 9714 -7780 9766 -7734
rect 9812 -7780 9864 -7734
rect 9910 -7780 9962 -7734
rect 10008 -7780 10060 -7734
rect 10106 -7780 10158 -7734
rect 10204 -7780 10256 -7734
rect 10302 -7780 10354 -7734
rect 10400 -7780 10452 -7734
rect 10498 -7780 10550 -7734
rect 10596 -7780 10648 -7734
rect 10694 -7780 10746 -7734
rect 10792 -7780 10844 -7734
rect 10890 -7780 10942 -7734
rect 10988 -7780 11040 -7734
rect 11086 -7780 11101 -7734
rect 8771 -7795 11101 -7780
rect 8771 -7832 8847 -7795
rect 8771 -7878 8786 -7832
rect 8832 -7878 8847 -7832
rect 8771 -7930 8847 -7878
rect 8771 -7976 8786 -7930
rect 8832 -7976 8847 -7930
rect 11025 -7832 11101 -7795
rect 11025 -7878 11040 -7832
rect 11086 -7878 11101 -7832
rect 11025 -7930 11101 -7878
rect 8771 -8028 8847 -7976
rect 8771 -8074 8786 -8028
rect 8832 -8074 8847 -8028
rect 8771 -8126 8847 -8074
rect 11025 -7976 11040 -7930
rect 11086 -7976 11101 -7930
rect 11025 -8028 11101 -7976
rect 11025 -8074 11040 -8028
rect 11086 -8074 11101 -8028
rect 8771 -8172 8786 -8126
rect 8832 -8172 8847 -8126
rect 8771 -8224 8847 -8172
rect 8771 -8270 8786 -8224
rect 8832 -8270 8847 -8224
rect 8771 -8322 8847 -8270
rect 8771 -8368 8786 -8322
rect 8832 -8368 8847 -8322
rect 8771 -8420 8847 -8368
rect 8771 -8466 8786 -8420
rect 8832 -8466 8847 -8420
rect 8771 -8518 8847 -8466
rect 8771 -8564 8786 -8518
rect 8832 -8564 8847 -8518
rect 8771 -8616 8847 -8564
rect 8771 -8662 8786 -8616
rect 8832 -8662 8847 -8616
rect 8771 -8714 8847 -8662
rect 8771 -8760 8786 -8714
rect 8832 -8760 8847 -8714
rect 11025 -8126 11101 -8074
rect 11025 -8172 11040 -8126
rect 11086 -8172 11101 -8126
rect 11025 -8224 11101 -8172
rect 11025 -8270 11040 -8224
rect 11086 -8270 11101 -8224
rect 11025 -8322 11101 -8270
rect 11025 -8368 11040 -8322
rect 11086 -8368 11101 -8322
rect 11025 -8420 11101 -8368
rect 11025 -8466 11040 -8420
rect 11086 -8466 11101 -8420
rect 11025 -8518 11101 -8466
rect 11025 -8564 11040 -8518
rect 11086 -8564 11101 -8518
rect 11025 -8616 11101 -8564
rect 11025 -8662 11040 -8616
rect 11086 -8662 11101 -8616
rect 11025 -8714 11101 -8662
rect 8771 -8812 8847 -8760
rect 8771 -8858 8786 -8812
rect 8832 -8858 8847 -8812
rect 11025 -8760 11040 -8714
rect 11086 -8760 11101 -8714
rect 11025 -8812 11101 -8760
rect 8771 -8910 8847 -8858
rect 8771 -8956 8786 -8910
rect 8832 -8956 8847 -8910
rect 2895 -9080 2971 -9028
rect 2895 -9126 2910 -9080
rect 2956 -9126 2971 -9080
rect 1621 -9224 1636 -9178
rect 1682 -9224 1697 -9178
rect 2895 -9178 2971 -9126
rect 1621 -9276 1697 -9224
rect 1621 -9322 1636 -9276
rect 1682 -9322 1697 -9276
rect 1621 -9374 1697 -9322
rect 1621 -9420 1636 -9374
rect 1682 -9420 1697 -9374
rect 1621 -9472 1697 -9420
rect 1621 -9518 1636 -9472
rect 1682 -9518 1697 -9472
rect 2895 -9224 2910 -9178
rect 2956 -9224 2971 -9178
rect 2895 -9276 2971 -9224
rect 2895 -9322 2910 -9276
rect 2956 -9322 2971 -9276
rect 2895 -9374 2971 -9322
rect 2895 -9420 2910 -9374
rect 2956 -9420 2971 -9374
rect 2895 -9472 2971 -9420
rect 1621 -9570 1697 -9518
rect 1621 -9616 1636 -9570
rect 1682 -9616 1697 -9570
rect 2895 -9518 2910 -9472
rect 2956 -9518 2971 -9472
rect 2895 -9570 2971 -9518
rect 1621 -9668 1697 -9616
rect 1621 -9714 1636 -9668
rect 1682 -9714 1697 -9668
rect 1621 -9766 1697 -9714
rect 1621 -9812 1636 -9766
rect 1682 -9812 1697 -9766
rect 1621 -9864 1697 -9812
rect 1621 -9910 1636 -9864
rect 1682 -9910 1697 -9864
rect 1621 -9962 1697 -9910
rect 1621 -10008 1636 -9962
rect 1682 -10008 1697 -9962
rect 1621 -10060 1697 -10008
rect 1621 -10106 1636 -10060
rect 1682 -10106 1697 -10060
rect 1621 -10158 1697 -10106
rect 1621 -10204 1636 -10158
rect 1682 -10204 1697 -10158
rect 1621 -10256 1697 -10204
rect 1621 -10302 1636 -10256
rect 1682 -10302 1697 -10256
rect 1621 -10339 1697 -10302
rect 2895 -9616 2910 -9570
rect 2956 -9616 2971 -9570
rect 2895 -9668 2971 -9616
rect 2895 -9714 2910 -9668
rect 2956 -9714 2971 -9668
rect 2895 -9766 2971 -9714
rect 2895 -9812 2910 -9766
rect 2956 -9812 2971 -9766
rect 2895 -9864 2971 -9812
rect 2895 -9910 2910 -9864
rect 2956 -9910 2971 -9864
rect 2895 -9962 2971 -9910
rect 2895 -10008 2910 -9962
rect 2956 -10008 2971 -9962
rect 2895 -10060 2971 -10008
rect 2895 -10106 2910 -10060
rect 2956 -10106 2971 -10060
rect 2895 -10158 2971 -10106
rect 2895 -10204 2910 -10158
rect 2956 -10204 2971 -10158
rect 2895 -10256 2971 -10204
rect 2895 -10302 2910 -10256
rect 2956 -10302 2971 -10256
rect 2895 -10339 2971 -10302
rect 1621 -10354 2971 -10339
rect 1621 -10400 1636 -10354
rect 1682 -10400 1734 -10354
rect 1780 -10400 1832 -10354
rect 1878 -10400 1930 -10354
rect 1976 -10400 2028 -10354
rect 2074 -10400 2126 -10354
rect 2172 -10400 2224 -10354
rect 2270 -10400 2322 -10354
rect 2368 -10400 2420 -10354
rect 2466 -10400 2518 -10354
rect 2564 -10400 2616 -10354
rect 2662 -10400 2714 -10354
rect 2760 -10400 2812 -10354
rect 2858 -10400 2910 -10354
rect 2956 -10400 2971 -10354
rect 1621 -10415 2971 -10400
rect 8771 -9008 8847 -8956
rect 8771 -9054 8786 -9008
rect 8832 -9054 8847 -9008
rect 8771 -9106 8847 -9054
rect 8771 -9152 8786 -9106
rect 8832 -9152 8847 -9106
rect 8771 -9204 8847 -9152
rect 8771 -9250 8786 -9204
rect 8832 -9250 8847 -9204
rect 8771 -9302 8847 -9250
rect 8771 -9348 8786 -9302
rect 8832 -9348 8847 -9302
rect 8771 -9400 8847 -9348
rect 8771 -9446 8786 -9400
rect 8832 -9446 8847 -9400
rect 8771 -9498 8847 -9446
rect 11025 -8858 11040 -8812
rect 11086 -8858 11101 -8812
rect 11025 -8910 11101 -8858
rect 11025 -8956 11040 -8910
rect 11086 -8956 11101 -8910
rect 11025 -9008 11101 -8956
rect 11025 -9054 11040 -9008
rect 11086 -9054 11101 -9008
rect 11025 -9106 11101 -9054
rect 11025 -9152 11040 -9106
rect 11086 -9152 11101 -9106
rect 11025 -9204 11101 -9152
rect 11025 -9250 11040 -9204
rect 11086 -9250 11101 -9204
rect 11025 -9302 11101 -9250
rect 11025 -9348 11040 -9302
rect 11086 -9348 11101 -9302
rect 11025 -9400 11101 -9348
rect 11025 -9446 11040 -9400
rect 11086 -9446 11101 -9400
rect 8771 -9544 8786 -9498
rect 8832 -9544 8847 -9498
rect 8771 -9596 8847 -9544
rect 11025 -9498 11101 -9446
rect 11025 -9544 11040 -9498
rect 11086 -9544 11101 -9498
rect 8771 -9642 8786 -9596
rect 8832 -9642 8847 -9596
rect 8771 -9694 8847 -9642
rect 8771 -9740 8786 -9694
rect 8832 -9740 8847 -9694
rect 8771 -9792 8847 -9740
rect 8771 -9838 8786 -9792
rect 8832 -9838 8847 -9792
rect 8771 -9890 8847 -9838
rect 8771 -9936 8786 -9890
rect 8832 -9936 8847 -9890
rect 8771 -9988 8847 -9936
rect 8771 -10034 8786 -9988
rect 8832 -10034 8847 -9988
rect 8771 -10086 8847 -10034
rect 8771 -10132 8786 -10086
rect 8832 -10132 8847 -10086
rect 8771 -10184 8847 -10132
rect 8771 -10230 8786 -10184
rect 8832 -10230 8847 -10184
rect 11025 -9596 11101 -9544
rect 11025 -9642 11040 -9596
rect 11086 -9642 11101 -9596
rect 11025 -9694 11101 -9642
rect 11025 -9740 11040 -9694
rect 11086 -9740 11101 -9694
rect 11025 -9792 11101 -9740
rect 11025 -9838 11040 -9792
rect 11086 -9838 11101 -9792
rect 11025 -9890 11101 -9838
rect 11025 -9936 11040 -9890
rect 11086 -9936 11101 -9890
rect 11025 -9988 11101 -9936
rect 11025 -10034 11040 -9988
rect 11086 -10034 11101 -9988
rect 11025 -10086 11101 -10034
rect 11025 -10132 11040 -10086
rect 11086 -10132 11101 -10086
rect 11025 -10184 11101 -10132
rect 8771 -10282 8847 -10230
rect 8771 -10328 8786 -10282
rect 8832 -10328 8847 -10282
rect 8771 -10380 8847 -10328
rect 11025 -10230 11040 -10184
rect 11086 -10230 11101 -10184
rect 11025 -10282 11101 -10230
rect 11025 -10328 11040 -10282
rect 11086 -10328 11101 -10282
rect 1200 -10478 1215 -10432
rect 1261 -10478 1276 -10432
rect 1200 -10530 1276 -10478
rect 1200 -10576 1215 -10530
rect 1261 -10576 1276 -10530
rect 8771 -10426 8786 -10380
rect 8832 -10426 8847 -10380
rect 8771 -10463 8847 -10426
rect 11025 -10380 11101 -10328
rect 11025 -10426 11040 -10380
rect 11086 -10426 11101 -10380
rect 11025 -10463 11101 -10426
rect 8771 -10478 11101 -10463
rect 8771 -10524 8786 -10478
rect 8832 -10524 8884 -10478
rect 8930 -10524 8982 -10478
rect 9028 -10524 9080 -10478
rect 9126 -10524 9178 -10478
rect 9224 -10524 9276 -10478
rect 9322 -10524 9374 -10478
rect 9420 -10524 9472 -10478
rect 9518 -10524 9570 -10478
rect 9616 -10524 9668 -10478
rect 9714 -10524 9766 -10478
rect 9812 -10524 9864 -10478
rect 9910 -10524 9962 -10478
rect 10008 -10524 10060 -10478
rect 10106 -10524 10158 -10478
rect 10204 -10524 10256 -10478
rect 10302 -10524 10354 -10478
rect 10400 -10524 10452 -10478
rect 10498 -10524 10550 -10478
rect 10596 -10524 10648 -10478
rect 10694 -10524 10746 -10478
rect 10792 -10524 10844 -10478
rect 10890 -10524 10942 -10478
rect 10988 -10524 11040 -10478
rect 11086 -10524 11101 -10478
rect 8771 -10539 11101 -10524
rect 1200 -10613 1276 -10576
rect -564 -10628 1276 -10613
rect -564 -10674 -549 -10628
rect -503 -10674 -451 -10628
rect -405 -10674 -353 -10628
rect -307 -10674 -255 -10628
rect -209 -10674 -157 -10628
rect -111 -10674 -59 -10628
rect -13 -10674 39 -10628
rect 85 -10674 137 -10628
rect 183 -10674 235 -10628
rect 281 -10674 333 -10628
rect 379 -10674 431 -10628
rect 477 -10674 529 -10628
rect 575 -10674 627 -10628
rect 673 -10674 725 -10628
rect 771 -10674 823 -10628
rect 869 -10674 921 -10628
rect 967 -10674 1019 -10628
rect 1065 -10674 1117 -10628
rect 1163 -10674 1215 -10628
rect 1261 -10674 1276 -10628
rect -564 -10689 1276 -10674
<< nsubdiff >>
rect -3309 1441 -1257 1456
rect -3309 1394 -3294 1441
rect -3247 1395 -3199 1441
rect -3153 1395 -3105 1441
rect -3059 1395 -3011 1441
rect -2965 1395 -2917 1441
rect -2871 1395 -2823 1441
rect -2777 1395 -2729 1441
rect -2683 1395 -2635 1441
rect -2589 1395 -2541 1441
rect -2495 1395 -2447 1441
rect -2401 1395 -2353 1441
rect -2307 1395 -2259 1441
rect -2213 1395 -2165 1441
rect -2119 1395 -2071 1441
rect -2025 1395 -1977 1441
rect -1931 1395 -1883 1441
rect -1837 1395 -1789 1441
rect -1743 1395 -1695 1441
rect -1649 1395 -1601 1441
rect -1555 1395 -1507 1441
rect -1461 1395 -1413 1441
rect -1367 1395 -1319 1441
rect -3247 1394 -1319 1395
rect -1272 1394 -1257 1441
rect -3309 1380 -1257 1394
rect -3309 1346 -3233 1380
rect -3309 1300 -3294 1346
rect -3248 1300 -3233 1346
rect -3309 1252 -3233 1300
rect -1333 1346 -1257 1380
rect -1333 1300 -1318 1346
rect -1272 1300 -1257 1346
rect -3309 1206 -3294 1252
rect -3248 1206 -3233 1252
rect -3309 1158 -3233 1206
rect -1333 1252 -1257 1300
rect -1333 1206 -1318 1252
rect -1272 1206 -1257 1252
rect -3309 1112 -3294 1158
rect -3248 1112 -3233 1158
rect -3309 1064 -3233 1112
rect -3309 1018 -3294 1064
rect -3248 1018 -3233 1064
rect -3309 970 -3233 1018
rect -3309 924 -3294 970
rect -3248 924 -3233 970
rect -3309 876 -3233 924
rect -3309 830 -3294 876
rect -3248 830 -3233 876
rect -3309 782 -3233 830
rect -3309 736 -3294 782
rect -3248 736 -3233 782
rect -3309 688 -3233 736
rect -3309 642 -3294 688
rect -3248 642 -3233 688
rect -3309 594 -3233 642
rect -3309 548 -3294 594
rect -3248 548 -3233 594
rect -3309 500 -3233 548
rect -1333 1158 -1257 1206
rect -1333 1112 -1318 1158
rect -1272 1112 -1257 1158
rect -1333 1064 -1257 1112
rect -1333 1018 -1318 1064
rect -1272 1018 -1257 1064
rect 2361 1155 4695 1170
rect 2361 1109 2377 1155
rect 2423 1109 2471 1155
rect 2517 1109 2565 1155
rect 2611 1109 2659 1155
rect 2705 1109 2753 1155
rect 2799 1109 2847 1155
rect 2893 1109 2941 1155
rect 2987 1109 3035 1155
rect 3081 1109 3129 1155
rect 3175 1109 3223 1155
rect 3269 1109 3317 1155
rect 3363 1109 3411 1155
rect 3457 1109 3505 1155
rect 3551 1109 3599 1155
rect 3645 1109 3693 1155
rect 3739 1109 3787 1155
rect 3833 1109 3881 1155
rect 3927 1109 3975 1155
rect 4021 1109 4069 1155
rect 4115 1109 4163 1155
rect 4209 1109 4257 1155
rect 4303 1109 4351 1155
rect 4397 1109 4445 1155
rect 4491 1109 4539 1155
rect 4585 1109 4633 1155
rect 4679 1109 4695 1155
rect 2361 1094 4695 1109
rect 2361 1061 2437 1094
rect -1333 970 -1257 1018
rect -1333 924 -1318 970
rect -1272 924 -1257 970
rect -1333 876 -1257 924
rect -1333 830 -1318 876
rect -1272 830 -1257 876
rect -1333 782 -1257 830
rect -1333 736 -1318 782
rect -1272 736 -1257 782
rect -1333 688 -1257 736
rect -1333 642 -1318 688
rect -1272 642 -1257 688
rect -1333 594 -1257 642
rect -1333 548 -1318 594
rect -1272 548 -1257 594
rect -3309 454 -3294 500
rect -3248 454 -3233 500
rect -1333 500 -1257 548
rect -3309 406 -3233 454
rect -1333 454 -1318 500
rect -1272 454 -1257 500
rect -3309 360 -3294 406
rect -3248 360 -3233 406
rect -3309 312 -3233 360
rect -3309 266 -3294 312
rect -3248 266 -3233 312
rect -3309 218 -3233 266
rect -3309 172 -3294 218
rect -3248 172 -3233 218
rect -3309 124 -3233 172
rect -3309 78 -3294 124
rect -3248 78 -3233 124
rect -3309 30 -3233 78
rect -3309 -16 -3294 30
rect -3248 -16 -3233 30
rect -3309 -64 -3233 -16
rect -3309 -110 -3294 -64
rect -3248 -110 -3233 -64
rect -3309 -158 -3233 -110
rect -3309 -204 -3294 -158
rect -3248 -204 -3233 -158
rect -3309 -252 -3233 -204
rect -1333 406 -1257 454
rect -1333 360 -1318 406
rect -1272 360 -1257 406
rect -1333 312 -1257 360
rect -1333 266 -1318 312
rect -1272 266 -1257 312
rect -1333 218 -1257 266
rect -1333 172 -1318 218
rect -1272 172 -1257 218
rect -1333 124 -1257 172
rect -1333 78 -1318 124
rect -1272 78 -1257 124
rect -1333 30 -1257 78
rect -1333 -16 -1318 30
rect -1272 -16 -1257 30
rect -1333 -64 -1257 -16
rect -1333 -110 -1318 -64
rect -1272 -110 -1257 -64
rect -1333 -158 -1257 -110
rect -1333 -204 -1318 -158
rect -1272 -204 -1257 -158
rect -3309 -298 -3294 -252
rect -3248 -298 -3233 -252
rect -1333 -252 -1257 -204
rect -3309 -346 -3233 -298
rect -3309 -392 -3294 -346
rect -3248 -392 -3233 -346
rect -3309 -440 -3233 -392
rect -3309 -486 -3294 -440
rect -3248 -486 -3233 -440
rect -3309 -534 -3233 -486
rect -3309 -580 -3294 -534
rect -3248 -580 -3233 -534
rect -3309 -628 -3233 -580
rect -3309 -674 -3294 -628
rect -3248 -674 -3233 -628
rect -3309 -722 -3233 -674
rect -3309 -768 -3294 -722
rect -3248 -768 -3233 -722
rect -3309 -816 -3233 -768
rect -3309 -862 -3294 -816
rect -3248 -862 -3233 -816
rect -3309 -910 -3233 -862
rect -3309 -956 -3294 -910
rect -3248 -956 -3233 -910
rect -1333 -298 -1318 -252
rect -1272 -298 -1257 -252
rect -1333 -346 -1257 -298
rect -1333 -392 -1318 -346
rect -1272 -392 -1257 -346
rect -1333 -440 -1257 -392
rect -1333 -486 -1318 -440
rect -1272 -486 -1257 -440
rect -1333 -534 -1257 -486
rect -1333 -580 -1318 -534
rect -1272 -580 -1257 -534
rect -1333 -628 -1257 -580
rect -1333 -674 -1318 -628
rect -1272 -674 -1257 -628
rect -1333 -722 -1257 -674
rect -1333 -768 -1318 -722
rect -1272 -768 -1257 -722
rect -1333 -816 -1257 -768
rect -1333 -862 -1318 -816
rect -1272 -862 -1257 -816
rect -1333 -910 -1257 -862
rect -3309 -1004 -3233 -956
rect -3309 -1050 -3294 -1004
rect -3248 -1050 -3233 -1004
rect -1333 -956 -1318 -910
rect -1272 -956 -1257 -910
rect -1333 -1004 -1257 -956
rect -3309 -1098 -3233 -1050
rect -3309 -1144 -3294 -1098
rect -3248 -1144 -3233 -1098
rect -3309 -1192 -3233 -1144
rect -3309 -1238 -3294 -1192
rect -3248 -1238 -3233 -1192
rect -3309 -1286 -3233 -1238
rect -3309 -1332 -3294 -1286
rect -3248 -1332 -3233 -1286
rect -3309 -1380 -3233 -1332
rect -3309 -1426 -3294 -1380
rect -3248 -1426 -3233 -1380
rect -3309 -1474 -3233 -1426
rect -3309 -1520 -3294 -1474
rect -3248 -1520 -3233 -1474
rect -3309 -1568 -3233 -1520
rect -3309 -1614 -3294 -1568
rect -3248 -1614 -3233 -1568
rect -3309 -1662 -3233 -1614
rect -3309 -1708 -3294 -1662
rect -3248 -1708 -3233 -1662
rect -3309 -1756 -3233 -1708
rect -3309 -1802 -3294 -1756
rect -3248 -1802 -3233 -1756
rect -3309 -1850 -3233 -1802
rect -3309 -1896 -3294 -1850
rect -3248 -1896 -3233 -1850
rect -3309 -1929 -3233 -1896
rect -1333 -1050 -1318 -1004
rect -1272 -1050 -1257 -1004
rect -1333 -1098 -1257 -1050
rect -1333 -1144 -1318 -1098
rect -1272 -1144 -1257 -1098
rect -1333 -1192 -1257 -1144
rect -1333 -1238 -1318 -1192
rect -1272 -1238 -1257 -1192
rect -1333 -1286 -1257 -1238
rect -1333 -1332 -1318 -1286
rect -1272 -1332 -1257 -1286
rect -1333 -1380 -1257 -1332
rect -1333 -1426 -1318 -1380
rect -1272 -1426 -1257 -1380
rect -1333 -1474 -1257 -1426
rect -1333 -1520 -1318 -1474
rect -1272 -1520 -1257 -1474
rect -1333 -1568 -1257 -1520
rect -1333 -1614 -1318 -1568
rect -1272 -1614 -1257 -1568
rect -1333 -1662 -1257 -1614
rect -1333 -1708 -1318 -1662
rect -1272 -1708 -1257 -1662
rect -1333 -1756 -1257 -1708
rect -1333 -1802 -1318 -1756
rect -1272 -1802 -1257 -1756
rect -1333 -1850 -1257 -1802
rect -1333 -1896 -1318 -1850
rect -1272 -1896 -1257 -1850
rect -1333 -1929 -1257 -1896
rect -3309 -1944 -1257 -1929
rect -3309 -1990 -3293 -1944
rect -3247 -1990 -3199 -1944
rect -3153 -1990 -3105 -1944
rect -3059 -1990 -3011 -1944
rect -2965 -1990 -2917 -1944
rect -2871 -1990 -2823 -1944
rect -2777 -1990 -2729 -1944
rect -2683 -1990 -2635 -1944
rect -2589 -1990 -2541 -1944
rect -2495 -1990 -2447 -1944
rect -2401 -1990 -2353 -1944
rect -2307 -1990 -2259 -1944
rect -2213 -1990 -2165 -1944
rect -2119 -1990 -2071 -1944
rect -2025 -1990 -1977 -1944
rect -1931 -1990 -1883 -1944
rect -1837 -1990 -1789 -1944
rect -1743 -1990 -1695 -1944
rect -1649 -1990 -1601 -1944
rect -1555 -1990 -1507 -1944
rect -1461 -1990 -1413 -1944
rect -1367 -1990 -1319 -1944
rect -1273 -1990 -1257 -1944
rect -3309 -2005 -1257 -1990
rect -762 1013 1233 1028
rect -762 967 -747 1013
rect -701 967 -653 1013
rect -607 967 -552 1013
rect -506 967 -458 1013
rect -412 967 -362 1013
rect -316 967 -268 1013
rect -222 967 -167 1013
rect -121 967 -73 1013
rect -27 967 21 1013
rect 67 967 115 1013
rect 161 967 216 1013
rect 262 967 310 1013
rect 356 967 406 1013
rect 452 967 500 1013
rect 546 967 601 1013
rect 647 967 695 1013
rect 741 967 789 1013
rect 835 967 883 1013
rect 929 967 984 1013
rect 1030 967 1078 1013
rect 1124 967 1172 1013
rect 1218 967 1233 1013
rect -762 952 1233 967
rect -762 917 -686 952
rect -762 871 -747 917
rect -701 871 -686 917
rect -762 823 -686 871
rect 1157 917 1233 952
rect 1157 871 1172 917
rect 1218 871 1233 917
rect -762 777 -747 823
rect -701 777 -686 823
rect -762 727 -686 777
rect 1157 816 1233 871
rect 1157 770 1172 816
rect 1218 770 1233 816
rect -762 681 -747 727
rect -701 681 -686 727
rect -762 633 -686 681
rect -762 587 -747 633
rect -701 587 -686 633
rect -762 539 -686 587
rect -762 493 -747 539
rect -701 493 -686 539
rect -762 438 -686 493
rect -762 392 -747 438
rect -701 392 -686 438
rect -762 344 -686 392
rect -762 298 -747 344
rect -701 298 -686 344
rect -762 248 -686 298
rect -762 202 -747 248
rect -701 202 -686 248
rect -762 154 -686 202
rect -762 108 -747 154
rect -701 108 -686 154
rect -762 53 -686 108
rect 1157 722 1233 770
rect 1157 676 1172 722
rect 1218 676 1233 722
rect 1157 628 1233 676
rect 1157 582 1172 628
rect 1218 582 1233 628
rect 1157 534 1233 582
rect 1157 488 1172 534
rect 1218 488 1233 534
rect 1157 433 1233 488
rect 1157 387 1172 433
rect 1218 387 1233 433
rect 1157 339 1233 387
rect 1157 293 1172 339
rect 1218 293 1233 339
rect 1157 243 1233 293
rect 1157 197 1172 243
rect 1218 197 1233 243
rect 1157 149 1233 197
rect 1157 103 1172 149
rect 1218 103 1233 149
rect -762 7 -747 53
rect -701 7 -686 53
rect -762 -41 -686 7
rect -762 -87 -747 -41
rect -701 -87 -686 -41
rect -762 -135 -686 -87
rect -762 -181 -747 -135
rect -701 -181 -686 -135
rect -762 -229 -686 -181
rect -762 -275 -747 -229
rect -701 -275 -686 -229
rect -762 -330 -686 -275
rect 1157 48 1233 103
rect 1157 2 1172 48
rect 1218 2 1233 48
rect 1157 -46 1233 2
rect 1157 -92 1172 -46
rect 1218 -92 1233 -46
rect 1157 -140 1233 -92
rect 1157 -186 1172 -140
rect 1218 -186 1233 -140
rect 1157 -234 1233 -186
rect 1157 -280 1172 -234
rect 1218 -280 1233 -234
rect -762 -376 -747 -330
rect -701 -376 -686 -330
rect -762 -424 -686 -376
rect -762 -470 -747 -424
rect -701 -470 -686 -424
rect -762 -520 -686 -470
rect -762 -566 -747 -520
rect -701 -566 -686 -520
rect -762 -614 -686 -566
rect -762 -660 -747 -614
rect -701 -660 -686 -614
rect -762 -715 -686 -660
rect -762 -761 -747 -715
rect -701 -761 -686 -715
rect -762 -809 -686 -761
rect -762 -855 -747 -809
rect -701 -855 -686 -809
rect -762 -903 -686 -855
rect -762 -949 -747 -903
rect -701 -949 -686 -903
rect -762 -997 -686 -949
rect 1157 -335 1233 -280
rect 1157 -381 1172 -335
rect 1218 -381 1233 -335
rect 1157 -429 1233 -381
rect 1157 -475 1172 -429
rect 1218 -475 1233 -429
rect 1157 -525 1233 -475
rect 1157 -571 1172 -525
rect 1218 -571 1233 -525
rect 1157 -619 1233 -571
rect 1157 -665 1172 -619
rect 1218 -665 1233 -619
rect 1157 -720 1233 -665
rect 1157 -766 1172 -720
rect 1218 -766 1233 -720
rect 1157 -814 1233 -766
rect 1157 -860 1172 -814
rect 1218 -860 1233 -814
rect 1157 -908 1233 -860
rect 1157 -954 1172 -908
rect 1218 -954 1233 -908
rect -762 -1043 -747 -997
rect -701 -1043 -686 -997
rect -762 -1098 -686 -1043
rect -762 -1144 -747 -1098
rect -701 -1144 -686 -1098
rect -762 -1192 -686 -1144
rect -762 -1238 -747 -1192
rect -701 -1238 -686 -1192
rect -762 -1288 -686 -1238
rect -762 -1334 -747 -1288
rect -701 -1334 -686 -1288
rect 1157 -1004 1233 -954
rect 1157 -1050 1172 -1004
rect 1218 -1050 1233 -1004
rect 1157 -1098 1233 -1050
rect 1157 -1144 1172 -1098
rect 1218 -1144 1233 -1098
rect 1157 -1199 1233 -1144
rect 1157 -1245 1172 -1199
rect 1218 -1245 1233 -1199
rect 1157 -1293 1233 -1245
rect -762 -1382 -686 -1334
rect -762 -1428 -747 -1382
rect -701 -1428 -686 -1382
rect -762 -1476 -686 -1428
rect -762 -1522 -747 -1476
rect -701 -1522 -686 -1476
rect -762 -1577 -686 -1522
rect -762 -1623 -747 -1577
rect -701 -1623 -686 -1577
rect -762 -1671 -686 -1623
rect -762 -1717 -747 -1671
rect -701 -1717 -686 -1671
rect -762 -1767 -686 -1717
rect -762 -1813 -747 -1767
rect -701 -1813 -686 -1767
rect -762 -1861 -686 -1813
rect -762 -1907 -747 -1861
rect -701 -1907 -686 -1861
rect -762 -1962 -686 -1907
rect -762 -2008 -747 -1962
rect -701 -2008 -686 -1962
rect 1157 -1339 1172 -1293
rect 1218 -1339 1233 -1293
rect 1157 -1387 1233 -1339
rect 1157 -1433 1172 -1387
rect 1218 -1433 1233 -1387
rect 1157 -1481 1233 -1433
rect 1157 -1527 1172 -1481
rect 1218 -1527 1233 -1481
rect 1157 -1582 1233 -1527
rect 1157 -1628 1172 -1582
rect 1218 -1628 1233 -1582
rect 1157 -1676 1233 -1628
rect 1157 -1722 1172 -1676
rect 1218 -1722 1233 -1676
rect 1157 -1772 1233 -1722
rect 1157 -1818 1172 -1772
rect 1218 -1818 1233 -1772
rect 1157 -1866 1233 -1818
rect 1157 -1912 1172 -1866
rect 1218 -1912 1233 -1866
rect 1157 -1967 1233 -1912
rect -762 -2056 -686 -2008
rect -762 -2102 -747 -2056
rect -701 -2102 -686 -2056
rect -762 -2150 -686 -2102
rect -762 -2196 -747 -2150
rect -701 -2196 -686 -2150
rect -762 -2244 -686 -2196
rect -762 -2290 -747 -2244
rect -701 -2290 -686 -2244
rect -762 -2345 -686 -2290
rect -762 -2391 -747 -2345
rect -701 -2391 -686 -2345
rect 1157 -2013 1172 -1967
rect 1218 -2013 1233 -1967
rect 1157 -2061 1233 -2013
rect 1157 -2107 1172 -2061
rect 1218 -2107 1233 -2061
rect 1157 -2155 1233 -2107
rect 1157 -2201 1172 -2155
rect 1218 -2201 1233 -2155
rect 1157 -2249 1233 -2201
rect 1157 -2295 1172 -2249
rect 1218 -2295 1233 -2249
rect 1157 -2350 1233 -2295
rect -762 -2439 -686 -2391
rect -762 -2485 -747 -2439
rect -701 -2485 -686 -2439
rect -762 -2535 -686 -2485
rect -3282 -2593 -1230 -2578
rect -3282 -2640 -3267 -2593
rect -3220 -2639 -3172 -2593
rect -3126 -2639 -3078 -2593
rect -3032 -2639 -2984 -2593
rect -2938 -2639 -2890 -2593
rect -2844 -2639 -2796 -2593
rect -2750 -2639 -2702 -2593
rect -2656 -2639 -2608 -2593
rect -2562 -2639 -2514 -2593
rect -2468 -2639 -2420 -2593
rect -2374 -2639 -2326 -2593
rect -2280 -2639 -2232 -2593
rect -2186 -2639 -2138 -2593
rect -2092 -2639 -2044 -2593
rect -1998 -2639 -1950 -2593
rect -1904 -2639 -1856 -2593
rect -1810 -2639 -1762 -2593
rect -1716 -2639 -1668 -2593
rect -1622 -2639 -1574 -2593
rect -1528 -2639 -1480 -2593
rect -1434 -2639 -1386 -2593
rect -1340 -2639 -1292 -2593
rect -3220 -2640 -1292 -2639
rect -1245 -2640 -1230 -2593
rect -3282 -2654 -1230 -2640
rect -3282 -2688 -3206 -2654
rect -3282 -2734 -3267 -2688
rect -3221 -2734 -3206 -2688
rect -1306 -2688 -1230 -2654
rect -3282 -2782 -3206 -2734
rect -3282 -2828 -3267 -2782
rect -3221 -2828 -3206 -2782
rect -3282 -2876 -3206 -2828
rect -1306 -2734 -1291 -2688
rect -1245 -2734 -1230 -2688
rect -1306 -2782 -1230 -2734
rect -1306 -2828 -1291 -2782
rect -1245 -2828 -1230 -2782
rect -3282 -2922 -3267 -2876
rect -3221 -2922 -3206 -2876
rect -3282 -2970 -3206 -2922
rect -1306 -2876 -1230 -2828
rect -1306 -2922 -1291 -2876
rect -1245 -2922 -1230 -2876
rect -3282 -3016 -3267 -2970
rect -3221 -3016 -3206 -2970
rect -3282 -3064 -3206 -3016
rect -1306 -2970 -1230 -2922
rect -1306 -3016 -1291 -2970
rect -1245 -3016 -1230 -2970
rect -3282 -3110 -3267 -3064
rect -3221 -3110 -3206 -3064
rect -3282 -3158 -3206 -3110
rect -3282 -3204 -3267 -3158
rect -3221 -3204 -3206 -3158
rect -3282 -3252 -3206 -3204
rect -3282 -3298 -3267 -3252
rect -3221 -3298 -3206 -3252
rect -3282 -3346 -3206 -3298
rect -3282 -3392 -3267 -3346
rect -3221 -3392 -3206 -3346
rect -3282 -3440 -3206 -3392
rect -3282 -3486 -3267 -3440
rect -3221 -3486 -3206 -3440
rect -3282 -3534 -3206 -3486
rect -1306 -3064 -1230 -3016
rect -1306 -3110 -1291 -3064
rect -1245 -3110 -1230 -3064
rect -1306 -3158 -1230 -3110
rect -1306 -3204 -1291 -3158
rect -1245 -3204 -1230 -3158
rect -1306 -3252 -1230 -3204
rect -1306 -3298 -1291 -3252
rect -1245 -3298 -1230 -3252
rect -1306 -3346 -1230 -3298
rect -1306 -3392 -1291 -3346
rect -1245 -3392 -1230 -3346
rect -762 -2581 -747 -2535
rect -701 -2581 -686 -2535
rect -762 -2629 -686 -2581
rect -762 -2675 -747 -2629
rect -701 -2675 -686 -2629
rect -762 -2730 -686 -2675
rect -762 -2776 -747 -2730
rect -701 -2776 -686 -2730
rect -762 -2824 -686 -2776
rect -762 -2870 -747 -2824
rect -701 -2870 -686 -2824
rect -762 -2918 -686 -2870
rect -762 -2964 -747 -2918
rect -701 -2964 -686 -2918
rect -762 -3012 -686 -2964
rect -762 -3058 -747 -3012
rect -701 -3058 -686 -3012
rect 1157 -2396 1172 -2350
rect 1218 -2396 1233 -2350
rect 1157 -2444 1233 -2396
rect 1157 -2490 1172 -2444
rect 1218 -2490 1233 -2444
rect 1157 -2540 1233 -2490
rect 1157 -2586 1172 -2540
rect 1218 -2586 1233 -2540
rect 1157 -2634 1233 -2586
rect 1157 -2680 1172 -2634
rect 1218 -2680 1233 -2634
rect 1157 -2735 1233 -2680
rect 1157 -2781 1172 -2735
rect 1218 -2781 1233 -2735
rect 1157 -2829 1233 -2781
rect 1157 -2875 1172 -2829
rect 1218 -2875 1233 -2829
rect 1157 -2923 1233 -2875
rect 1157 -2969 1172 -2923
rect 1218 -2969 1233 -2923
rect 2361 1015 2376 1061
rect 2422 1015 2437 1061
rect 2361 967 2437 1015
rect 4619 1061 4695 1094
rect 4619 1015 4634 1061
rect 4680 1015 4695 1061
rect 2361 921 2376 967
rect 2422 921 2437 967
rect 2361 873 2437 921
rect 2361 827 2376 873
rect 2422 827 2437 873
rect 2361 779 2437 827
rect 2361 733 2376 779
rect 2422 733 2437 779
rect 2361 685 2437 733
rect 2361 639 2376 685
rect 2422 639 2437 685
rect 2361 591 2437 639
rect 2361 545 2376 591
rect 2422 545 2437 591
rect 2361 497 2437 545
rect 2361 451 2376 497
rect 2422 451 2437 497
rect 2361 403 2437 451
rect 2361 357 2376 403
rect 2422 357 2437 403
rect 2361 309 2437 357
rect 2361 263 2376 309
rect 2422 263 2437 309
rect 2361 215 2437 263
rect 4619 967 4695 1015
rect 4619 921 4634 967
rect 4680 921 4695 967
rect 4619 873 4695 921
rect 4619 827 4634 873
rect 4680 827 4695 873
rect 4619 779 4695 827
rect 4619 733 4634 779
rect 4680 733 4695 779
rect 4619 685 4695 733
rect 4619 639 4634 685
rect 4680 639 4695 685
rect 4619 591 4695 639
rect 4619 545 4634 591
rect 4680 545 4695 591
rect 4619 497 4695 545
rect 4619 451 4634 497
rect 4680 451 4695 497
rect 4619 403 4695 451
rect 4619 357 4634 403
rect 4680 357 4695 403
rect 4619 309 4695 357
rect 4619 263 4634 309
rect 4680 263 4695 309
rect 2361 169 2376 215
rect 2422 169 2437 215
rect 2361 121 2437 169
rect 4619 215 4695 263
rect 4619 169 4634 215
rect 4680 169 4695 215
rect 2361 75 2376 121
rect 2422 75 2437 121
rect 2361 27 2437 75
rect 2361 -19 2376 27
rect 2422 -19 2437 27
rect 2361 -67 2437 -19
rect 2361 -113 2376 -67
rect 2422 -113 2437 -67
rect 2361 -161 2437 -113
rect 2361 -207 2376 -161
rect 2422 -207 2437 -161
rect 2361 -255 2437 -207
rect 2361 -301 2376 -255
rect 2422 -301 2437 -255
rect 2361 -349 2437 -301
rect 2361 -395 2376 -349
rect 2422 -395 2437 -349
rect 2361 -443 2437 -395
rect 2361 -489 2376 -443
rect 2422 -489 2437 -443
rect 2361 -537 2437 -489
rect 4619 121 4695 169
rect 4619 75 4634 121
rect 4680 75 4695 121
rect 4619 27 4695 75
rect 4619 -19 4634 27
rect 4680 -19 4695 27
rect 4619 -67 4695 -19
rect 4619 -113 4634 -67
rect 4680 -113 4695 -67
rect 4619 -161 4695 -113
rect 4619 -207 4634 -161
rect 4680 -207 4695 -161
rect 4619 -255 4695 -207
rect 4619 -301 4634 -255
rect 4680 -301 4695 -255
rect 4619 -349 4695 -301
rect 4619 -395 4634 -349
rect 4680 -395 4695 -349
rect 4619 -443 4695 -395
rect 4619 -489 4634 -443
rect 4680 -489 4695 -443
rect 2361 -583 2376 -537
rect 2422 -583 2437 -537
rect 2361 -631 2437 -583
rect 4619 -537 4695 -489
rect 4619 -583 4634 -537
rect 4680 -583 4695 -537
rect 2361 -677 2376 -631
rect 2422 -677 2437 -631
rect 2361 -725 2437 -677
rect 2361 -771 2376 -725
rect 2422 -771 2437 -725
rect 2361 -819 2437 -771
rect 2361 -865 2376 -819
rect 2422 -865 2437 -819
rect 2361 -913 2437 -865
rect 2361 -959 2376 -913
rect 2422 -959 2437 -913
rect 2361 -1007 2437 -959
rect 2361 -1053 2376 -1007
rect 2422 -1053 2437 -1007
rect 2361 -1101 2437 -1053
rect 2361 -1147 2376 -1101
rect 2422 -1147 2437 -1101
rect 2361 -1195 2437 -1147
rect 2361 -1241 2376 -1195
rect 2422 -1241 2437 -1195
rect 2361 -1289 2437 -1241
rect 4619 -631 4695 -583
rect 4619 -677 4634 -631
rect 4680 -677 4695 -631
rect 4619 -725 4695 -677
rect 4619 -771 4634 -725
rect 4680 -771 4695 -725
rect 4619 -819 4695 -771
rect 4619 -865 4634 -819
rect 4680 -865 4695 -819
rect 4619 -913 4695 -865
rect 4619 -959 4634 -913
rect 4680 -959 4695 -913
rect 4619 -1007 4695 -959
rect 4619 -1053 4634 -1007
rect 4680 -1053 4695 -1007
rect 4619 -1101 4695 -1053
rect 4619 -1147 4634 -1101
rect 4680 -1147 4695 -1101
rect 4619 -1195 4695 -1147
rect 4619 -1241 4634 -1195
rect 4680 -1241 4695 -1195
rect 2361 -1335 2376 -1289
rect 2422 -1335 2437 -1289
rect 2361 -1383 2437 -1335
rect 4619 -1289 4695 -1241
rect 4619 -1335 4634 -1289
rect 4680 -1335 4695 -1289
rect 2361 -1429 2376 -1383
rect 2422 -1429 2437 -1383
rect 2361 -1477 2437 -1429
rect 2361 -1523 2376 -1477
rect 2422 -1523 2437 -1477
rect 2361 -1571 2437 -1523
rect 2361 -1617 2376 -1571
rect 2422 -1617 2437 -1571
rect 2361 -1665 2437 -1617
rect 2361 -1711 2376 -1665
rect 2422 -1711 2437 -1665
rect 2361 -1759 2437 -1711
rect 2361 -1805 2376 -1759
rect 2422 -1805 2437 -1759
rect 2361 -1853 2437 -1805
rect 2361 -1899 2376 -1853
rect 2422 -1899 2437 -1853
rect 2361 -1947 2437 -1899
rect 2361 -1993 2376 -1947
rect 2422 -1993 2437 -1947
rect 4619 -1383 4695 -1335
rect 4619 -1429 4634 -1383
rect 4680 -1429 4695 -1383
rect 4619 -1477 4695 -1429
rect 4619 -1523 4634 -1477
rect 4680 -1523 4695 -1477
rect 4619 -1571 4695 -1523
rect 4619 -1617 4634 -1571
rect 4680 -1617 4695 -1571
rect 4619 -1665 4695 -1617
rect 4619 -1711 4634 -1665
rect 4680 -1711 4695 -1665
rect 4619 -1759 4695 -1711
rect 4619 -1805 4634 -1759
rect 4680 -1805 4695 -1759
rect 4619 -1853 4695 -1805
rect 4619 -1899 4634 -1853
rect 4680 -1899 4695 -1853
rect 4619 -1947 4695 -1899
rect 2361 -2041 2437 -1993
rect 2361 -2087 2376 -2041
rect 2422 -2087 2437 -2041
rect 4619 -1993 4634 -1947
rect 4680 -1993 4695 -1947
rect 4619 -2041 4695 -1993
rect 2361 -2135 2437 -2087
rect 2361 -2181 2376 -2135
rect 2422 -2181 2437 -2135
rect 2361 -2229 2437 -2181
rect 2361 -2275 2376 -2229
rect 2422 -2275 2437 -2229
rect 2361 -2323 2437 -2275
rect 2361 -2369 2376 -2323
rect 2422 -2369 2437 -2323
rect 2361 -2417 2437 -2369
rect 2361 -2463 2376 -2417
rect 2422 -2463 2437 -2417
rect 2361 -2511 2437 -2463
rect 2361 -2557 2376 -2511
rect 2422 -2557 2437 -2511
rect 2361 -2605 2437 -2557
rect 2361 -2651 2376 -2605
rect 2422 -2651 2437 -2605
rect 2361 -2699 2437 -2651
rect 2361 -2745 2376 -2699
rect 2422 -2745 2437 -2699
rect 2361 -2793 2437 -2745
rect 2361 -2839 2376 -2793
rect 2422 -2839 2437 -2793
rect 4619 -2087 4634 -2041
rect 4680 -2087 4695 -2041
rect 4619 -2135 4695 -2087
rect 4619 -2181 4634 -2135
rect 4680 -2181 4695 -2135
rect 4619 -2229 4695 -2181
rect 4619 -2275 4634 -2229
rect 4680 -2275 4695 -2229
rect 4619 -2323 4695 -2275
rect 4619 -2369 4634 -2323
rect 4680 -2369 4695 -2323
rect 4619 -2417 4695 -2369
rect 4619 -2463 4634 -2417
rect 4680 -2463 4695 -2417
rect 4619 -2511 4695 -2463
rect 4619 -2557 4634 -2511
rect 4680 -2557 4695 -2511
rect 4619 -2605 4695 -2557
rect 4619 -2651 4634 -2605
rect 4680 -2651 4695 -2605
rect 4619 -2699 4695 -2651
rect 4619 -2745 4634 -2699
rect 4680 -2745 4695 -2699
rect 4619 -2793 4695 -2745
rect 2361 -2872 2437 -2839
rect 4619 -2839 4634 -2793
rect 4680 -2839 4695 -2793
rect 4619 -2872 4695 -2839
rect 2361 -2887 4695 -2872
rect 2361 -2933 2377 -2887
rect 2423 -2933 2471 -2887
rect 2517 -2933 2565 -2887
rect 2611 -2933 2659 -2887
rect 2705 -2933 2753 -2887
rect 2799 -2933 2847 -2887
rect 2893 -2933 2941 -2887
rect 2987 -2933 3035 -2887
rect 3081 -2933 3129 -2887
rect 3175 -2933 3223 -2887
rect 3269 -2933 3317 -2887
rect 3363 -2933 3411 -2887
rect 3457 -2933 3505 -2887
rect 3551 -2933 3599 -2887
rect 3645 -2933 3693 -2887
rect 3739 -2933 3787 -2887
rect 3833 -2933 3881 -2887
rect 3927 -2933 3975 -2887
rect 4021 -2933 4069 -2887
rect 4115 -2933 4163 -2887
rect 4209 -2933 4257 -2887
rect 4303 -2933 4351 -2887
rect 4397 -2933 4445 -2887
rect 4491 -2933 4539 -2887
rect 4585 -2933 4633 -2887
rect 4679 -2933 4695 -2887
rect 2361 -2948 4695 -2933
rect 5161 1155 7495 1170
rect 5161 1109 5177 1155
rect 5223 1109 5271 1155
rect 5317 1109 5365 1155
rect 5411 1109 5459 1155
rect 5505 1109 5553 1155
rect 5599 1109 5647 1155
rect 5693 1109 5741 1155
rect 5787 1109 5835 1155
rect 5881 1109 5929 1155
rect 5975 1109 6023 1155
rect 6069 1109 6117 1155
rect 6163 1109 6211 1155
rect 6257 1109 6305 1155
rect 6351 1109 6399 1155
rect 6445 1109 6493 1155
rect 6539 1109 6587 1155
rect 6633 1109 6681 1155
rect 6727 1109 6775 1155
rect 6821 1109 6869 1155
rect 6915 1109 6963 1155
rect 7009 1109 7057 1155
rect 7103 1109 7151 1155
rect 7197 1109 7245 1155
rect 7291 1109 7339 1155
rect 7385 1109 7433 1155
rect 7479 1109 7495 1155
rect 5161 1094 7495 1109
rect 5161 1061 5237 1094
rect 5161 1015 5176 1061
rect 5222 1015 5237 1061
rect 5161 967 5237 1015
rect 7419 1061 7495 1094
rect 7419 1015 7434 1061
rect 7480 1015 7495 1061
rect 5161 921 5176 967
rect 5222 921 5237 967
rect 5161 873 5237 921
rect 5161 827 5176 873
rect 5222 827 5237 873
rect 5161 779 5237 827
rect 5161 733 5176 779
rect 5222 733 5237 779
rect 5161 685 5237 733
rect 5161 639 5176 685
rect 5222 639 5237 685
rect 5161 591 5237 639
rect 5161 545 5176 591
rect 5222 545 5237 591
rect 5161 497 5237 545
rect 5161 451 5176 497
rect 5222 451 5237 497
rect 5161 403 5237 451
rect 5161 357 5176 403
rect 5222 357 5237 403
rect 5161 309 5237 357
rect 5161 263 5176 309
rect 5222 263 5237 309
rect 5161 215 5237 263
rect 7419 967 7495 1015
rect 7419 921 7434 967
rect 7480 921 7495 967
rect 7419 873 7495 921
rect 7419 827 7434 873
rect 7480 827 7495 873
rect 7419 779 7495 827
rect 7419 733 7434 779
rect 7480 733 7495 779
rect 7419 685 7495 733
rect 7419 639 7434 685
rect 7480 639 7495 685
rect 7419 591 7495 639
rect 7419 545 7434 591
rect 7480 545 7495 591
rect 7419 497 7495 545
rect 7419 451 7434 497
rect 7480 451 7495 497
rect 7419 403 7495 451
rect 7419 357 7434 403
rect 7480 357 7495 403
rect 7419 309 7495 357
rect 7419 263 7434 309
rect 7480 263 7495 309
rect 5161 169 5176 215
rect 5222 169 5237 215
rect 5161 121 5237 169
rect 7419 215 7495 263
rect 7419 169 7434 215
rect 7480 169 7495 215
rect 5161 75 5176 121
rect 5222 75 5237 121
rect 5161 27 5237 75
rect 5161 -19 5176 27
rect 5222 -19 5237 27
rect 5161 -67 5237 -19
rect 5161 -113 5176 -67
rect 5222 -113 5237 -67
rect 5161 -161 5237 -113
rect 5161 -207 5176 -161
rect 5222 -207 5237 -161
rect 5161 -255 5237 -207
rect 5161 -301 5176 -255
rect 5222 -301 5237 -255
rect 5161 -349 5237 -301
rect 5161 -395 5176 -349
rect 5222 -395 5237 -349
rect 5161 -443 5237 -395
rect 5161 -489 5176 -443
rect 5222 -489 5237 -443
rect 5161 -537 5237 -489
rect 7419 121 7495 169
rect 7419 75 7434 121
rect 7480 75 7495 121
rect 7419 27 7495 75
rect 7419 -19 7434 27
rect 7480 -19 7495 27
rect 7419 -67 7495 -19
rect 7419 -113 7434 -67
rect 7480 -113 7495 -67
rect 7419 -161 7495 -113
rect 7419 -207 7434 -161
rect 7480 -207 7495 -161
rect 7419 -255 7495 -207
rect 7419 -301 7434 -255
rect 7480 -301 7495 -255
rect 7419 -349 7495 -301
rect 7419 -395 7434 -349
rect 7480 -395 7495 -349
rect 7419 -443 7495 -395
rect 7419 -489 7434 -443
rect 7480 -489 7495 -443
rect 5161 -583 5176 -537
rect 5222 -583 5237 -537
rect 5161 -631 5237 -583
rect 7419 -537 7495 -489
rect 7419 -583 7434 -537
rect 7480 -583 7495 -537
rect 5161 -677 5176 -631
rect 5222 -677 5237 -631
rect 5161 -725 5237 -677
rect 5161 -771 5176 -725
rect 5222 -771 5237 -725
rect 5161 -819 5237 -771
rect 5161 -865 5176 -819
rect 5222 -865 5237 -819
rect 5161 -913 5237 -865
rect 5161 -959 5176 -913
rect 5222 -959 5237 -913
rect 5161 -1007 5237 -959
rect 5161 -1053 5176 -1007
rect 5222 -1053 5237 -1007
rect 5161 -1101 5237 -1053
rect 5161 -1147 5176 -1101
rect 5222 -1147 5237 -1101
rect 5161 -1195 5237 -1147
rect 5161 -1241 5176 -1195
rect 5222 -1241 5237 -1195
rect 5161 -1289 5237 -1241
rect 7419 -631 7495 -583
rect 7419 -677 7434 -631
rect 7480 -677 7495 -631
rect 7419 -725 7495 -677
rect 7419 -771 7434 -725
rect 7480 -771 7495 -725
rect 7419 -819 7495 -771
rect 7419 -865 7434 -819
rect 7480 -865 7495 -819
rect 7419 -913 7495 -865
rect 7419 -959 7434 -913
rect 7480 -959 7495 -913
rect 7419 -1007 7495 -959
rect 7419 -1053 7434 -1007
rect 7480 -1053 7495 -1007
rect 7419 -1101 7495 -1053
rect 7419 -1147 7434 -1101
rect 7480 -1147 7495 -1101
rect 7419 -1195 7495 -1147
rect 7419 -1241 7434 -1195
rect 7480 -1241 7495 -1195
rect 5161 -1335 5176 -1289
rect 5222 -1335 5237 -1289
rect 5161 -1383 5237 -1335
rect 7419 -1289 7495 -1241
rect 7419 -1335 7434 -1289
rect 7480 -1335 7495 -1289
rect 5161 -1429 5176 -1383
rect 5222 -1429 5237 -1383
rect 5161 -1477 5237 -1429
rect 5161 -1523 5176 -1477
rect 5222 -1523 5237 -1477
rect 5161 -1571 5237 -1523
rect 5161 -1617 5176 -1571
rect 5222 -1617 5237 -1571
rect 5161 -1665 5237 -1617
rect 5161 -1711 5176 -1665
rect 5222 -1711 5237 -1665
rect 5161 -1759 5237 -1711
rect 5161 -1805 5176 -1759
rect 5222 -1805 5237 -1759
rect 5161 -1853 5237 -1805
rect 5161 -1899 5176 -1853
rect 5222 -1899 5237 -1853
rect 5161 -1947 5237 -1899
rect 5161 -1993 5176 -1947
rect 5222 -1993 5237 -1947
rect 7419 -1383 7495 -1335
rect 7419 -1429 7434 -1383
rect 7480 -1429 7495 -1383
rect 7419 -1477 7495 -1429
rect 7419 -1523 7434 -1477
rect 7480 -1523 7495 -1477
rect 7419 -1571 7495 -1523
rect 7419 -1617 7434 -1571
rect 7480 -1617 7495 -1571
rect 7419 -1665 7495 -1617
rect 7419 -1711 7434 -1665
rect 7480 -1711 7495 -1665
rect 7419 -1759 7495 -1711
rect 7419 -1805 7434 -1759
rect 7480 -1805 7495 -1759
rect 7419 -1853 7495 -1805
rect 7419 -1899 7434 -1853
rect 7480 -1899 7495 -1853
rect 7419 -1947 7495 -1899
rect 5161 -2041 5237 -1993
rect 5161 -2087 5176 -2041
rect 5222 -2087 5237 -2041
rect 7419 -1993 7434 -1947
rect 7480 -1993 7495 -1947
rect 7419 -2041 7495 -1993
rect 5161 -2135 5237 -2087
rect 5161 -2181 5176 -2135
rect 5222 -2181 5237 -2135
rect 5161 -2229 5237 -2181
rect 5161 -2275 5176 -2229
rect 5222 -2275 5237 -2229
rect 5161 -2323 5237 -2275
rect 5161 -2369 5176 -2323
rect 5222 -2369 5237 -2323
rect 5161 -2417 5237 -2369
rect 5161 -2463 5176 -2417
rect 5222 -2463 5237 -2417
rect 5161 -2511 5237 -2463
rect 5161 -2557 5176 -2511
rect 5222 -2557 5237 -2511
rect 5161 -2605 5237 -2557
rect 5161 -2651 5176 -2605
rect 5222 -2651 5237 -2605
rect 5161 -2699 5237 -2651
rect 5161 -2745 5176 -2699
rect 5222 -2745 5237 -2699
rect 5161 -2793 5237 -2745
rect 5161 -2839 5176 -2793
rect 5222 -2839 5237 -2793
rect 7419 -2087 7434 -2041
rect 7480 -2087 7495 -2041
rect 7419 -2135 7495 -2087
rect 7419 -2181 7434 -2135
rect 7480 -2181 7495 -2135
rect 7419 -2229 7495 -2181
rect 7419 -2275 7434 -2229
rect 7480 -2275 7495 -2229
rect 7419 -2323 7495 -2275
rect 7419 -2369 7434 -2323
rect 7480 -2369 7495 -2323
rect 7419 -2417 7495 -2369
rect 7419 -2463 7434 -2417
rect 7480 -2463 7495 -2417
rect 7419 -2511 7495 -2463
rect 7419 -2557 7434 -2511
rect 7480 -2557 7495 -2511
rect 7419 -2605 7495 -2557
rect 7419 -2651 7434 -2605
rect 7480 -2651 7495 -2605
rect 7419 -2699 7495 -2651
rect 7419 -2745 7434 -2699
rect 7480 -2745 7495 -2699
rect 7419 -2793 7495 -2745
rect 5161 -2872 5237 -2839
rect 7419 -2839 7434 -2793
rect 7480 -2839 7495 -2793
rect 7419 -2872 7495 -2839
rect 5161 -2887 7495 -2872
rect 5161 -2933 5177 -2887
rect 5223 -2933 5271 -2887
rect 5317 -2933 5365 -2887
rect 5411 -2933 5459 -2887
rect 5505 -2933 5553 -2887
rect 5599 -2933 5647 -2887
rect 5693 -2933 5741 -2887
rect 5787 -2933 5835 -2887
rect 5881 -2933 5929 -2887
rect 5975 -2933 6023 -2887
rect 6069 -2933 6117 -2887
rect 6163 -2933 6211 -2887
rect 6257 -2933 6305 -2887
rect 6351 -2933 6399 -2887
rect 6445 -2933 6493 -2887
rect 6539 -2933 6587 -2887
rect 6633 -2933 6681 -2887
rect 6727 -2933 6775 -2887
rect 6821 -2933 6869 -2887
rect 6915 -2933 6963 -2887
rect 7009 -2933 7057 -2887
rect 7103 -2933 7151 -2887
rect 7197 -2933 7245 -2887
rect 7291 -2933 7339 -2887
rect 7385 -2933 7433 -2887
rect 7479 -2933 7495 -2887
rect 5161 -2948 7495 -2933
rect 7961 1155 10295 1170
rect 7961 1109 7977 1155
rect 8023 1109 8071 1155
rect 8117 1109 8165 1155
rect 8211 1109 8259 1155
rect 8305 1109 8353 1155
rect 8399 1109 8447 1155
rect 8493 1109 8541 1155
rect 8587 1109 8635 1155
rect 8681 1109 8729 1155
rect 8775 1109 8823 1155
rect 8869 1109 8917 1155
rect 8963 1109 9011 1155
rect 9057 1109 9105 1155
rect 9151 1109 9199 1155
rect 9245 1109 9293 1155
rect 9339 1109 9387 1155
rect 9433 1109 9481 1155
rect 9527 1109 9575 1155
rect 9621 1109 9669 1155
rect 9715 1109 9763 1155
rect 9809 1109 9857 1155
rect 9903 1109 9951 1155
rect 9997 1109 10045 1155
rect 10091 1109 10139 1155
rect 10185 1109 10233 1155
rect 10279 1109 10295 1155
rect 7961 1094 10295 1109
rect 7961 1061 8037 1094
rect 7961 1015 7976 1061
rect 8022 1015 8037 1061
rect 7961 967 8037 1015
rect 10219 1061 10295 1094
rect 10219 1015 10234 1061
rect 10280 1015 10295 1061
rect 7961 921 7976 967
rect 8022 921 8037 967
rect 7961 873 8037 921
rect 7961 827 7976 873
rect 8022 827 8037 873
rect 7961 779 8037 827
rect 7961 733 7976 779
rect 8022 733 8037 779
rect 7961 685 8037 733
rect 7961 639 7976 685
rect 8022 639 8037 685
rect 7961 591 8037 639
rect 7961 545 7976 591
rect 8022 545 8037 591
rect 7961 497 8037 545
rect 7961 451 7976 497
rect 8022 451 8037 497
rect 7961 403 8037 451
rect 7961 357 7976 403
rect 8022 357 8037 403
rect 7961 309 8037 357
rect 7961 263 7976 309
rect 8022 263 8037 309
rect 7961 215 8037 263
rect 10219 967 10295 1015
rect 10219 921 10234 967
rect 10280 921 10295 967
rect 10219 873 10295 921
rect 10219 827 10234 873
rect 10280 827 10295 873
rect 10219 779 10295 827
rect 10219 733 10234 779
rect 10280 733 10295 779
rect 10219 685 10295 733
rect 10219 639 10234 685
rect 10280 639 10295 685
rect 10219 591 10295 639
rect 10219 545 10234 591
rect 10280 545 10295 591
rect 10219 497 10295 545
rect 10219 451 10234 497
rect 10280 451 10295 497
rect 10219 403 10295 451
rect 10219 357 10234 403
rect 10280 357 10295 403
rect 10219 309 10295 357
rect 10219 263 10234 309
rect 10280 263 10295 309
rect 7961 169 7976 215
rect 8022 169 8037 215
rect 7961 121 8037 169
rect 10219 215 10295 263
rect 10219 169 10234 215
rect 10280 169 10295 215
rect 7961 75 7976 121
rect 8022 75 8037 121
rect 7961 27 8037 75
rect 7961 -19 7976 27
rect 8022 -19 8037 27
rect 7961 -67 8037 -19
rect 7961 -113 7976 -67
rect 8022 -113 8037 -67
rect 7961 -161 8037 -113
rect 7961 -207 7976 -161
rect 8022 -207 8037 -161
rect 7961 -255 8037 -207
rect 7961 -301 7976 -255
rect 8022 -301 8037 -255
rect 7961 -349 8037 -301
rect 7961 -395 7976 -349
rect 8022 -395 8037 -349
rect 7961 -443 8037 -395
rect 7961 -489 7976 -443
rect 8022 -489 8037 -443
rect 7961 -537 8037 -489
rect 10219 121 10295 169
rect 10219 75 10234 121
rect 10280 75 10295 121
rect 10219 27 10295 75
rect 10219 -19 10234 27
rect 10280 -19 10295 27
rect 10219 -67 10295 -19
rect 10219 -113 10234 -67
rect 10280 -113 10295 -67
rect 10219 -161 10295 -113
rect 10219 -207 10234 -161
rect 10280 -207 10295 -161
rect 10219 -255 10295 -207
rect 10219 -301 10234 -255
rect 10280 -301 10295 -255
rect 10219 -349 10295 -301
rect 10219 -395 10234 -349
rect 10280 -395 10295 -349
rect 10219 -443 10295 -395
rect 10219 -489 10234 -443
rect 10280 -489 10295 -443
rect 7961 -583 7976 -537
rect 8022 -583 8037 -537
rect 7961 -631 8037 -583
rect 10219 -537 10295 -489
rect 10219 -583 10234 -537
rect 10280 -583 10295 -537
rect 7961 -677 7976 -631
rect 8022 -677 8037 -631
rect 7961 -725 8037 -677
rect 7961 -771 7976 -725
rect 8022 -771 8037 -725
rect 7961 -819 8037 -771
rect 7961 -865 7976 -819
rect 8022 -865 8037 -819
rect 7961 -913 8037 -865
rect 7961 -959 7976 -913
rect 8022 -959 8037 -913
rect 7961 -1007 8037 -959
rect 7961 -1053 7976 -1007
rect 8022 -1053 8037 -1007
rect 7961 -1101 8037 -1053
rect 7961 -1147 7976 -1101
rect 8022 -1147 8037 -1101
rect 7961 -1195 8037 -1147
rect 7961 -1241 7976 -1195
rect 8022 -1241 8037 -1195
rect 7961 -1289 8037 -1241
rect 10219 -631 10295 -583
rect 10219 -677 10234 -631
rect 10280 -677 10295 -631
rect 10219 -725 10295 -677
rect 10219 -771 10234 -725
rect 10280 -771 10295 -725
rect 10219 -819 10295 -771
rect 10219 -865 10234 -819
rect 10280 -865 10295 -819
rect 10219 -913 10295 -865
rect 10219 -959 10234 -913
rect 10280 -959 10295 -913
rect 10219 -1007 10295 -959
rect 10219 -1053 10234 -1007
rect 10280 -1053 10295 -1007
rect 10219 -1101 10295 -1053
rect 10219 -1147 10234 -1101
rect 10280 -1147 10295 -1101
rect 10219 -1195 10295 -1147
rect 10219 -1241 10234 -1195
rect 10280 -1241 10295 -1195
rect 7961 -1335 7976 -1289
rect 8022 -1335 8037 -1289
rect 7961 -1383 8037 -1335
rect 10219 -1289 10295 -1241
rect 10219 -1335 10234 -1289
rect 10280 -1335 10295 -1289
rect 7961 -1429 7976 -1383
rect 8022 -1429 8037 -1383
rect 7961 -1477 8037 -1429
rect 7961 -1523 7976 -1477
rect 8022 -1523 8037 -1477
rect 7961 -1571 8037 -1523
rect 7961 -1617 7976 -1571
rect 8022 -1617 8037 -1571
rect 7961 -1665 8037 -1617
rect 7961 -1711 7976 -1665
rect 8022 -1711 8037 -1665
rect 7961 -1759 8037 -1711
rect 7961 -1805 7976 -1759
rect 8022 -1805 8037 -1759
rect 7961 -1853 8037 -1805
rect 7961 -1899 7976 -1853
rect 8022 -1899 8037 -1853
rect 7961 -1947 8037 -1899
rect 7961 -1993 7976 -1947
rect 8022 -1993 8037 -1947
rect 10219 -1383 10295 -1335
rect 10219 -1429 10234 -1383
rect 10280 -1429 10295 -1383
rect 10219 -1477 10295 -1429
rect 10219 -1523 10234 -1477
rect 10280 -1523 10295 -1477
rect 10219 -1571 10295 -1523
rect 10219 -1617 10234 -1571
rect 10280 -1617 10295 -1571
rect 10219 -1665 10295 -1617
rect 10219 -1711 10234 -1665
rect 10280 -1711 10295 -1665
rect 10219 -1759 10295 -1711
rect 10219 -1805 10234 -1759
rect 10280 -1805 10295 -1759
rect 10219 -1853 10295 -1805
rect 10219 -1899 10234 -1853
rect 10280 -1899 10295 -1853
rect 10219 -1947 10295 -1899
rect 7961 -2041 8037 -1993
rect 7961 -2087 7976 -2041
rect 8022 -2087 8037 -2041
rect 10219 -1993 10234 -1947
rect 10280 -1993 10295 -1947
rect 10219 -2041 10295 -1993
rect 7961 -2135 8037 -2087
rect 7961 -2181 7976 -2135
rect 8022 -2181 8037 -2135
rect 7961 -2229 8037 -2181
rect 7961 -2275 7976 -2229
rect 8022 -2275 8037 -2229
rect 7961 -2323 8037 -2275
rect 7961 -2369 7976 -2323
rect 8022 -2369 8037 -2323
rect 7961 -2417 8037 -2369
rect 7961 -2463 7976 -2417
rect 8022 -2463 8037 -2417
rect 7961 -2511 8037 -2463
rect 7961 -2557 7976 -2511
rect 8022 -2557 8037 -2511
rect 7961 -2605 8037 -2557
rect 7961 -2651 7976 -2605
rect 8022 -2651 8037 -2605
rect 7961 -2699 8037 -2651
rect 7961 -2745 7976 -2699
rect 8022 -2745 8037 -2699
rect 7961 -2793 8037 -2745
rect 7961 -2839 7976 -2793
rect 8022 -2839 8037 -2793
rect 10219 -2087 10234 -2041
rect 10280 -2087 10295 -2041
rect 10219 -2135 10295 -2087
rect 10219 -2181 10234 -2135
rect 10280 -2181 10295 -2135
rect 10219 -2229 10295 -2181
rect 10219 -2275 10234 -2229
rect 10280 -2275 10295 -2229
rect 10219 -2323 10295 -2275
rect 10219 -2369 10234 -2323
rect 10280 -2369 10295 -2323
rect 10219 -2417 10295 -2369
rect 10219 -2463 10234 -2417
rect 10280 -2463 10295 -2417
rect 10219 -2511 10295 -2463
rect 10219 -2557 10234 -2511
rect 10280 -2557 10295 -2511
rect 10219 -2605 10295 -2557
rect 10219 -2651 10234 -2605
rect 10280 -2651 10295 -2605
rect 10219 -2699 10295 -2651
rect 10219 -2745 10234 -2699
rect 10280 -2745 10295 -2699
rect 10219 -2793 10295 -2745
rect 7961 -2872 8037 -2839
rect 10219 -2839 10234 -2793
rect 10280 -2839 10295 -2793
rect 10219 -2872 10295 -2839
rect 7961 -2887 10295 -2872
rect 7961 -2933 7977 -2887
rect 8023 -2933 8071 -2887
rect 8117 -2933 8165 -2887
rect 8211 -2933 8259 -2887
rect 8305 -2933 8353 -2887
rect 8399 -2933 8447 -2887
rect 8493 -2933 8541 -2887
rect 8587 -2933 8635 -2887
rect 8681 -2933 8729 -2887
rect 8775 -2933 8823 -2887
rect 8869 -2933 8917 -2887
rect 8963 -2933 9011 -2887
rect 9057 -2933 9105 -2887
rect 9151 -2933 9199 -2887
rect 9245 -2933 9293 -2887
rect 9339 -2933 9387 -2887
rect 9433 -2933 9481 -2887
rect 9527 -2933 9575 -2887
rect 9621 -2933 9669 -2887
rect 9715 -2933 9763 -2887
rect 9809 -2933 9857 -2887
rect 9903 -2933 9951 -2887
rect 9997 -2933 10045 -2887
rect 10091 -2933 10139 -2887
rect 10185 -2933 10233 -2887
rect 10279 -2933 10295 -2887
rect 7961 -2948 10295 -2933
rect 1157 -3019 1233 -2969
rect -762 -3113 -686 -3058
rect -762 -3159 -747 -3113
rect -701 -3159 -686 -3113
rect -762 -3207 -686 -3159
rect 1157 -3065 1172 -3019
rect 1218 -3065 1233 -3019
rect 1157 -3113 1233 -3065
rect 1157 -3159 1172 -3113
rect 1218 -3159 1233 -3113
rect -762 -3253 -747 -3207
rect -701 -3253 -686 -3207
rect -762 -3288 -686 -3253
rect 1157 -3207 1233 -3159
rect 1157 -3253 1172 -3207
rect 1218 -3253 1233 -3207
rect 1157 -3288 1233 -3253
rect -762 -3303 1233 -3288
rect -762 -3349 -747 -3303
rect -701 -3349 -653 -3303
rect -607 -3349 -552 -3303
rect -506 -3349 -458 -3303
rect -412 -3349 -362 -3303
rect -316 -3349 -268 -3303
rect -222 -3349 -167 -3303
rect -121 -3349 -73 -3303
rect -27 -3349 21 -3303
rect 67 -3349 115 -3303
rect 161 -3349 216 -3303
rect 262 -3349 310 -3303
rect 356 -3349 406 -3303
rect 452 -3349 500 -3303
rect 546 -3349 601 -3303
rect 647 -3349 695 -3303
rect 741 -3349 789 -3303
rect 835 -3349 883 -3303
rect 929 -3349 984 -3303
rect 1030 -3349 1078 -3303
rect 1124 -3349 1172 -3303
rect 1218 -3349 1233 -3303
rect -762 -3364 1233 -3349
rect -1306 -3440 -1230 -3392
rect -1306 -3486 -1291 -3440
rect -1245 -3486 -1230 -3440
rect -3282 -3580 -3267 -3534
rect -3221 -3580 -3206 -3534
rect -3282 -3628 -3206 -3580
rect -3282 -3674 -3267 -3628
rect -3221 -3674 -3206 -3628
rect -1306 -3534 -1230 -3486
rect -1306 -3580 -1291 -3534
rect -1245 -3580 -1230 -3534
rect -1306 -3628 -1230 -3580
rect -3282 -3722 -3206 -3674
rect -1306 -3674 -1291 -3628
rect -1245 -3674 -1230 -3628
rect -3282 -3768 -3267 -3722
rect -3221 -3768 -3206 -3722
rect -3282 -3816 -3206 -3768
rect -3282 -3862 -3267 -3816
rect -3221 -3862 -3206 -3816
rect -3282 -3910 -3206 -3862
rect -3282 -3956 -3267 -3910
rect -3221 -3956 -3206 -3910
rect -3282 -4004 -3206 -3956
rect -1306 -3722 -1230 -3674
rect -1306 -3768 -1291 -3722
rect -1245 -3768 -1230 -3722
rect -1306 -3816 -1230 -3768
rect -1306 -3862 -1291 -3816
rect -1245 -3862 -1230 -3816
rect -1306 -3910 -1230 -3862
rect -1306 -3956 -1291 -3910
rect -1245 -3956 -1230 -3910
rect -3282 -4050 -3267 -4004
rect -3221 -4050 -3206 -4004
rect -1306 -4004 -1230 -3956
rect -3282 -4098 -3206 -4050
rect -3282 -4144 -3267 -4098
rect -3221 -4144 -3206 -4098
rect -3282 -4192 -3206 -4144
rect -3282 -4238 -3267 -4192
rect -3221 -4238 -3206 -4192
rect -3282 -4286 -3206 -4238
rect -3282 -4332 -3267 -4286
rect -3221 -4332 -3206 -4286
rect -3282 -4380 -3206 -4332
rect -1306 -4050 -1291 -4004
rect -1245 -4050 -1230 -4004
rect -1306 -4098 -1230 -4050
rect -1306 -4144 -1291 -4098
rect -1245 -4144 -1230 -4098
rect -1306 -4192 -1230 -4144
rect -1306 -4238 -1291 -4192
rect -1245 -4238 -1230 -4192
rect -1306 -4286 -1230 -4238
rect -1306 -4332 -1291 -4286
rect -1245 -4332 -1230 -4286
rect -3282 -4426 -3267 -4380
rect -3221 -4426 -3206 -4380
rect -3282 -4474 -3206 -4426
rect -3282 -4520 -3267 -4474
rect -3221 -4520 -3206 -4474
rect -1306 -4380 -1230 -4332
rect -1306 -4426 -1291 -4380
rect -1245 -4426 -1230 -4380
rect -3282 -4568 -3206 -4520
rect -3282 -4614 -3267 -4568
rect -3221 -4614 -3206 -4568
rect -1306 -4474 -1230 -4426
rect -1306 -4520 -1291 -4474
rect -1245 -4520 -1230 -4474
rect -1306 -4568 -1230 -4520
rect -3282 -4662 -3206 -4614
rect -3282 -4708 -3267 -4662
rect -3221 -4708 -3206 -4662
rect -3282 -4756 -3206 -4708
rect -3282 -4802 -3267 -4756
rect -3221 -4802 -3206 -4756
rect -3282 -4850 -3206 -4802
rect -3282 -4896 -3267 -4850
rect -3221 -4896 -3206 -4850
rect -3282 -4944 -3206 -4896
rect -3282 -4990 -3267 -4944
rect -3221 -4990 -3206 -4944
rect -3282 -5038 -3206 -4990
rect -3282 -5084 -3267 -5038
rect -3221 -5084 -3206 -5038
rect -3282 -5132 -3206 -5084
rect -3282 -5178 -3267 -5132
rect -3221 -5178 -3206 -5132
rect -1306 -4614 -1291 -4568
rect -1245 -4614 -1230 -4568
rect -1306 -4662 -1230 -4614
rect -1306 -4708 -1291 -4662
rect -1245 -4708 -1230 -4662
rect -1306 -4756 -1230 -4708
rect -1306 -4802 -1291 -4756
rect -1245 -4802 -1230 -4756
rect -1306 -4850 -1230 -4802
rect -1306 -4896 -1291 -4850
rect -1245 -4896 -1230 -4850
rect -1306 -4944 -1230 -4896
rect -1306 -4990 -1291 -4944
rect -1245 -4990 -1230 -4944
rect -1306 -5038 -1230 -4990
rect -1306 -5084 -1291 -5038
rect -1245 -5084 -1230 -5038
rect -1306 -5132 -1230 -5084
rect -3282 -5226 -3206 -5178
rect -3282 -5272 -3267 -5226
rect -3221 -5272 -3206 -5226
rect -3282 -5320 -3206 -5272
rect -1306 -5178 -1291 -5132
rect -1245 -5178 -1230 -5132
rect -3282 -5366 -3267 -5320
rect -3221 -5366 -3206 -5320
rect -1306 -5226 -1230 -5178
rect -1306 -5272 -1291 -5226
rect -1245 -5272 -1230 -5226
rect -1306 -5320 -1230 -5272
rect -3282 -5414 -3206 -5366
rect -3282 -5460 -3267 -5414
rect -3221 -5460 -3206 -5414
rect -1306 -5366 -1291 -5320
rect -1245 -5366 -1230 -5320
rect -1306 -5414 -1230 -5366
rect -3282 -5508 -3206 -5460
rect -3282 -5554 -3267 -5508
rect -3221 -5554 -3206 -5508
rect -3282 -5602 -3206 -5554
rect -3282 -5648 -3267 -5602
rect -3221 -5648 -3206 -5602
rect -3282 -5696 -3206 -5648
rect -3282 -5742 -3267 -5696
rect -3221 -5742 -3206 -5696
rect -3282 -5790 -3206 -5742
rect -3282 -5836 -3267 -5790
rect -3221 -5836 -3206 -5790
rect -3282 -5884 -3206 -5836
rect -3282 -5930 -3267 -5884
rect -3221 -5930 -3206 -5884
rect -3282 -5978 -3206 -5930
rect -3282 -6024 -3267 -5978
rect -3221 -6024 -3206 -5978
rect -1306 -5460 -1291 -5414
rect -1245 -5460 -1230 -5414
rect -1306 -5508 -1230 -5460
rect -1306 -5554 -1291 -5508
rect -1245 -5554 -1230 -5508
rect -1306 -5602 -1230 -5554
rect -1306 -5648 -1291 -5602
rect -1245 -5648 -1230 -5602
rect -1306 -5696 -1230 -5648
rect -1306 -5742 -1291 -5696
rect -1245 -5742 -1230 -5696
rect -1306 -5790 -1230 -5742
rect -1306 -5836 -1291 -5790
rect -1245 -5836 -1230 -5790
rect -1306 -5884 -1230 -5836
rect -1306 -5930 -1291 -5884
rect -1245 -5930 -1230 -5884
rect -1306 -5978 -1230 -5930
rect -3282 -6072 -3206 -6024
rect -3282 -6118 -3267 -6072
rect -3221 -6118 -3206 -6072
rect -3282 -6166 -3206 -6118
rect -1306 -6024 -1291 -5978
rect -1245 -6024 -1230 -5978
rect -1306 -6072 -1230 -6024
rect -1306 -6118 -1291 -6072
rect -1245 -6118 -1230 -6072
rect -3282 -6212 -3267 -6166
rect -3221 -6212 -3206 -6166
rect -3282 -6245 -3206 -6212
rect -1306 -6166 -1230 -6118
rect -1306 -6212 -1291 -6166
rect -1245 -6212 -1230 -6166
rect -1306 -6245 -1230 -6212
rect -3282 -6260 -1230 -6245
rect -3282 -6306 -3266 -6260
rect -3220 -6306 -3172 -6260
rect -3126 -6306 -3078 -6260
rect -3032 -6306 -2984 -6260
rect -2938 -6306 -2890 -6260
rect -2844 -6306 -2796 -6260
rect -2750 -6306 -2702 -6260
rect -2656 -6306 -2608 -6260
rect -2562 -6306 -2514 -6260
rect -2468 -6306 -2420 -6260
rect -2374 -6306 -2326 -6260
rect -2280 -6306 -2232 -6260
rect -2186 -6306 -2138 -6260
rect -2092 -6306 -2044 -6260
rect -1998 -6306 -1950 -6260
rect -1904 -6306 -1856 -6260
rect -1810 -6306 -1762 -6260
rect -1716 -6306 -1668 -6260
rect -1622 -6306 -1574 -6260
rect -1528 -6306 -1480 -6260
rect -1434 -6306 -1386 -6260
rect -1340 -6306 -1292 -6260
rect -1246 -6306 -1230 -6260
rect -477 -4068 1293 -4053
rect -477 -4115 -462 -4068
rect -415 -4114 -367 -4068
rect -321 -4114 -273 -4068
rect -227 -4114 -179 -4068
rect -133 -4114 -85 -4068
rect -39 -4114 9 -4068
rect 55 -4114 103 -4068
rect 149 -4114 197 -4068
rect 243 -4114 291 -4068
rect 337 -4114 385 -4068
rect 431 -4114 479 -4068
rect 525 -4114 573 -4068
rect 619 -4114 667 -4068
rect 713 -4114 761 -4068
rect 807 -4114 855 -4068
rect 901 -4114 949 -4068
rect 995 -4114 1043 -4068
rect 1089 -4114 1137 -4068
rect 1183 -4114 1231 -4068
rect -415 -4115 1231 -4114
rect 1278 -4115 1293 -4068
rect -477 -4129 1293 -4115
rect -477 -4163 -401 -4129
rect -477 -4213 -462 -4163
rect -416 -4213 -401 -4163
rect -477 -4261 -401 -4213
rect 1217 -4163 1293 -4129
rect 1217 -4213 1232 -4163
rect 1278 -4213 1293 -4163
rect -477 -4307 -462 -4261
rect -416 -4307 -401 -4261
rect -477 -4355 -401 -4307
rect -477 -4401 -462 -4355
rect -416 -4401 -401 -4355
rect -477 -4449 -401 -4401
rect 1217 -4261 1293 -4213
rect 1217 -4307 1232 -4261
rect 1278 -4307 1293 -4261
rect 1217 -4355 1293 -4307
rect 1217 -4401 1232 -4355
rect 1278 -4401 1293 -4355
rect -477 -4495 -462 -4449
rect -416 -4495 -401 -4449
rect -477 -4543 -401 -4495
rect -477 -4589 -462 -4543
rect -416 -4589 -401 -4543
rect -477 -4637 -401 -4589
rect -477 -4683 -462 -4637
rect -416 -4683 -401 -4637
rect -477 -4731 -401 -4683
rect -477 -4777 -462 -4731
rect -416 -4777 -401 -4731
rect -477 -4825 -401 -4777
rect -477 -4871 -462 -4825
rect -416 -4871 -401 -4825
rect -477 -4919 -401 -4871
rect -477 -4965 -462 -4919
rect -416 -4965 -401 -4919
rect -477 -5013 -401 -4965
rect -477 -5059 -462 -5013
rect -416 -5059 -401 -5013
rect -477 -5107 -401 -5059
rect -477 -5153 -462 -5107
rect -416 -5153 -401 -5107
rect 1217 -4449 1293 -4401
rect 1217 -4495 1232 -4449
rect 1278 -4495 1293 -4449
rect 1217 -4543 1293 -4495
rect 1217 -4589 1232 -4543
rect 1278 -4589 1293 -4543
rect 1217 -4637 1293 -4589
rect 1217 -4683 1232 -4637
rect 1278 -4683 1293 -4637
rect 1217 -4731 1293 -4683
rect 1217 -4777 1232 -4731
rect 1278 -4777 1293 -4731
rect 1217 -4825 1293 -4777
rect 1217 -4871 1232 -4825
rect 1278 -4871 1293 -4825
rect 1217 -4919 1293 -4871
rect 1217 -4965 1232 -4919
rect 1278 -4965 1293 -4919
rect 1217 -5013 1293 -4965
rect 1217 -5059 1232 -5013
rect 1278 -5059 1293 -5013
rect 1217 -5107 1293 -5059
rect -477 -5201 -401 -5153
rect -477 -5247 -462 -5201
rect -416 -5247 -401 -5201
rect 1217 -5153 1232 -5107
rect 1278 -5153 1293 -5107
rect 1217 -5201 1293 -5153
rect -477 -5295 -401 -5247
rect -477 -5341 -462 -5295
rect -416 -5341 -401 -5295
rect -477 -5389 -401 -5341
rect -477 -5435 -462 -5389
rect -416 -5435 -401 -5389
rect -477 -5483 -401 -5435
rect -477 -5529 -462 -5483
rect -416 -5529 -401 -5483
rect -477 -5577 -401 -5529
rect -477 -5623 -462 -5577
rect -416 -5623 -401 -5577
rect -477 -5671 -401 -5623
rect -477 -5717 -462 -5671
rect -416 -5717 -401 -5671
rect -477 -5765 -401 -5717
rect -477 -5811 -462 -5765
rect -416 -5811 -401 -5765
rect -477 -5859 -401 -5811
rect -477 -5905 -462 -5859
rect -416 -5905 -401 -5859
rect -477 -5953 -401 -5905
rect -477 -5999 -462 -5953
rect -416 -5999 -401 -5953
rect -477 -6047 -401 -5999
rect -477 -6093 -462 -6047
rect -416 -6093 -401 -6047
rect -477 -6141 -401 -6093
rect -477 -6187 -462 -6141
rect -416 -6187 -401 -6141
rect -477 -6221 -401 -6187
rect 1217 -5247 1232 -5201
rect 1278 -5247 1293 -5201
rect 1217 -5295 1293 -5247
rect 1217 -5341 1232 -5295
rect 1278 -5341 1293 -5295
rect 1217 -5389 1293 -5341
rect 1217 -5435 1232 -5389
rect 1278 -5435 1293 -5389
rect 1217 -5483 1293 -5435
rect 1217 -5529 1232 -5483
rect 1278 -5529 1293 -5483
rect 1217 -5577 1293 -5529
rect 1217 -5623 1232 -5577
rect 1278 -5623 1293 -5577
rect 1217 -5671 1293 -5623
rect 1217 -5717 1232 -5671
rect 1278 -5717 1293 -5671
rect 1217 -5765 1293 -5717
rect 1217 -5811 1232 -5765
rect 1278 -5811 1293 -5765
rect 1217 -5859 1293 -5811
rect 1217 -5905 1232 -5859
rect 1278 -5905 1293 -5859
rect 1217 -5953 1293 -5905
rect 1217 -5999 1232 -5953
rect 1278 -5999 1293 -5953
rect 1217 -6047 1293 -5999
rect 1217 -6093 1232 -6047
rect 1278 -6093 1293 -6047
rect 1217 -6141 1293 -6093
rect 1217 -6187 1232 -6141
rect 1278 -6187 1293 -6141
rect 1217 -6221 1293 -6187
rect -477 -6235 1293 -6221
rect -477 -6282 -462 -6235
rect -415 -6236 1231 -6235
rect -415 -6282 -367 -6236
rect -321 -6282 -273 -6236
rect -227 -6282 -179 -6236
rect -133 -6282 -85 -6236
rect -39 -6282 9 -6236
rect 55 -6282 103 -6236
rect 149 -6282 197 -6236
rect 243 -6282 291 -6236
rect 337 -6282 385 -6236
rect 431 -6282 479 -6236
rect 525 -6282 573 -6236
rect 619 -6282 667 -6236
rect 713 -6282 761 -6236
rect 807 -6282 855 -6236
rect 901 -6282 949 -6236
rect 995 -6282 1043 -6236
rect 1089 -6282 1137 -6236
rect 1183 -6282 1231 -6236
rect 1278 -6282 1293 -6235
rect 1606 -4319 3752 -4304
rect 1606 -4365 1622 -4319
rect 1668 -4365 1716 -4319
rect 1762 -4365 1810 -4319
rect 1856 -4365 1904 -4319
rect 1950 -4365 1998 -4319
rect 2044 -4365 2092 -4319
rect 2138 -4365 2186 -4319
rect 2232 -4365 2280 -4319
rect 2326 -4365 2374 -4319
rect 2420 -4365 2468 -4319
rect 2514 -4365 2562 -4319
rect 2608 -4365 2656 -4319
rect 2702 -4365 2750 -4319
rect 2796 -4365 2844 -4319
rect 2890 -4365 2938 -4319
rect 2984 -4365 3032 -4319
rect 3078 -4365 3126 -4319
rect 3172 -4365 3220 -4319
rect 3266 -4365 3314 -4319
rect 3360 -4365 3408 -4319
rect 3454 -4365 3502 -4319
rect 3548 -4365 3596 -4319
rect 3642 -4365 3690 -4319
rect 3736 -4365 3752 -4319
rect 1606 -4380 3752 -4365
rect 1606 -4413 1682 -4380
rect 1606 -4459 1621 -4413
rect 1667 -4459 1682 -4413
rect 1606 -4507 1682 -4459
rect 1606 -4553 1621 -4507
rect 1667 -4553 1682 -4507
rect 1606 -4601 1682 -4553
rect 3676 -4413 3752 -4380
rect 3676 -4459 3691 -4413
rect 3737 -4459 3752 -4413
rect 3676 -4507 3752 -4459
rect 3676 -4553 3691 -4507
rect 3737 -4553 3752 -4507
rect 1606 -4647 1621 -4601
rect 1667 -4647 1682 -4601
rect 1606 -4695 1682 -4647
rect 3676 -4601 3752 -4553
rect 3676 -4647 3691 -4601
rect 3737 -4647 3752 -4601
rect 1606 -4741 1621 -4695
rect 1667 -4741 1682 -4695
rect 1606 -4789 1682 -4741
rect 1606 -4835 1621 -4789
rect 1667 -4835 1682 -4789
rect 1606 -4883 1682 -4835
rect 1606 -4929 1621 -4883
rect 1667 -4929 1682 -4883
rect 1606 -4977 1682 -4929
rect 1606 -5023 1621 -4977
rect 1667 -5023 1682 -4977
rect 1606 -5071 1682 -5023
rect 1606 -5117 1621 -5071
rect 1667 -5117 1682 -5071
rect 1606 -5165 1682 -5117
rect 3676 -4695 3752 -4647
rect 3676 -4741 3691 -4695
rect 3737 -4741 3752 -4695
rect 3676 -4789 3752 -4741
rect 3676 -4835 3691 -4789
rect 3737 -4835 3752 -4789
rect 3676 -4883 3752 -4835
rect 3676 -4929 3691 -4883
rect 3737 -4929 3752 -4883
rect 3676 -4977 3752 -4929
rect 3676 -5023 3691 -4977
rect 3737 -5023 3752 -4977
rect 3676 -5071 3752 -5023
rect 3676 -5117 3691 -5071
rect 3737 -5117 3752 -5071
rect 1606 -5211 1621 -5165
rect 1667 -5211 1682 -5165
rect 1606 -5259 1682 -5211
rect 1606 -5305 1621 -5259
rect 1667 -5305 1682 -5259
rect 1606 -5353 1682 -5305
rect 3676 -5165 3752 -5117
rect 3676 -5211 3691 -5165
rect 3737 -5211 3752 -5165
rect 3676 -5259 3752 -5211
rect 3676 -5305 3691 -5259
rect 3737 -5305 3752 -5259
rect 1606 -5399 1621 -5353
rect 1667 -5399 1682 -5353
rect 3676 -5353 3752 -5305
rect 1606 -5447 1682 -5399
rect 3676 -5399 3691 -5353
rect 3737 -5399 3752 -5353
rect 1606 -5493 1621 -5447
rect 1667 -5493 1682 -5447
rect 1606 -5541 1682 -5493
rect 1606 -5587 1621 -5541
rect 1667 -5587 1682 -5541
rect 1606 -5635 1682 -5587
rect 1606 -5681 1621 -5635
rect 1667 -5681 1682 -5635
rect 1606 -5729 1682 -5681
rect 1606 -5775 1621 -5729
rect 1667 -5775 1682 -5729
rect 1606 -5823 1682 -5775
rect 1606 -5869 1621 -5823
rect 1667 -5869 1682 -5823
rect 3676 -5447 3752 -5399
rect 3676 -5493 3691 -5447
rect 3737 -5493 3752 -5447
rect 3676 -5541 3752 -5493
rect 3676 -5587 3691 -5541
rect 3737 -5587 3752 -5541
rect 3676 -5635 3752 -5587
rect 3676 -5681 3691 -5635
rect 3737 -5681 3752 -5635
rect 3676 -5729 3752 -5681
rect 3676 -5775 3691 -5729
rect 3737 -5775 3752 -5729
rect 3676 -5823 3752 -5775
rect 1606 -5917 1682 -5869
rect 3676 -5869 3691 -5823
rect 3737 -5869 3752 -5823
rect 1606 -5963 1621 -5917
rect 1667 -5963 1682 -5917
rect 1606 -6011 1682 -5963
rect 1606 -6057 1621 -6011
rect 1667 -6057 1682 -6011
rect 3676 -5917 3752 -5869
rect 3676 -5963 3691 -5917
rect 3737 -5963 3752 -5917
rect 3676 -6011 3752 -5963
rect 1606 -6105 1682 -6057
rect 1606 -6151 1621 -6105
rect 1667 -6151 1682 -6105
rect 1606 -6184 1682 -6151
rect 3676 -6057 3691 -6011
rect 3737 -6057 3752 -6011
rect 3676 -6105 3752 -6057
rect 4013 -4422 6723 -4407
rect 4013 -4468 4029 -4422
rect 4075 -4468 4123 -4422
rect 4169 -4468 4217 -4422
rect 4263 -4468 4311 -4422
rect 4357 -4468 4405 -4422
rect 4451 -4468 4499 -4422
rect 4545 -4468 4593 -4422
rect 4639 -4468 4687 -4422
rect 4733 -4468 4781 -4422
rect 4827 -4468 4875 -4422
rect 4921 -4468 4969 -4422
rect 5015 -4468 5063 -4422
rect 5109 -4468 5157 -4422
rect 5203 -4468 5251 -4422
rect 5297 -4468 5345 -4422
rect 5391 -4468 5439 -4422
rect 5485 -4468 5533 -4422
rect 5579 -4468 5627 -4422
rect 5673 -4468 5721 -4422
rect 5767 -4468 5815 -4422
rect 5861 -4468 5909 -4422
rect 5955 -4468 6003 -4422
rect 6049 -4468 6097 -4422
rect 6143 -4468 6191 -4422
rect 6237 -4468 6285 -4422
rect 6331 -4468 6379 -4422
rect 6425 -4468 6473 -4422
rect 6519 -4468 6567 -4422
rect 6613 -4468 6661 -4422
rect 6707 -4468 6723 -4422
rect 4013 -4483 6723 -4468
rect 4013 -4516 4089 -4483
rect 4013 -4562 4028 -4516
rect 4074 -4562 4089 -4516
rect 4013 -4610 4089 -4562
rect 6647 -4516 6723 -4483
rect 6647 -4562 6662 -4516
rect 6708 -4562 6723 -4516
rect 4013 -4656 4028 -4610
rect 4074 -4656 4089 -4610
rect 4013 -4704 4089 -4656
rect 4013 -4750 4028 -4704
rect 4074 -4750 4089 -4704
rect 6647 -4610 6723 -4562
rect 6647 -4656 6662 -4610
rect 6708 -4656 6723 -4610
rect 6647 -4704 6723 -4656
rect 4013 -4798 4089 -4750
rect 4013 -4844 4028 -4798
rect 4074 -4844 4089 -4798
rect 4013 -4892 4089 -4844
rect 4013 -4938 4028 -4892
rect 4074 -4938 4089 -4892
rect 4013 -4986 4089 -4938
rect 4013 -5032 4028 -4986
rect 4074 -5032 4089 -4986
rect 4013 -5080 4089 -5032
rect 4013 -5126 4028 -5080
rect 4074 -5126 4089 -5080
rect 4013 -5174 4089 -5126
rect 4013 -5220 4028 -5174
rect 4074 -5220 4089 -5174
rect 6647 -4750 6662 -4704
rect 6708 -4750 6723 -4704
rect 6647 -4798 6723 -4750
rect 6647 -4844 6662 -4798
rect 6708 -4844 6723 -4798
rect 6647 -4892 6723 -4844
rect 6647 -4938 6662 -4892
rect 6708 -4938 6723 -4892
rect 6647 -4986 6723 -4938
rect 6647 -5032 6662 -4986
rect 6708 -5032 6723 -4986
rect 6647 -5080 6723 -5032
rect 6647 -5126 6662 -5080
rect 6708 -5126 6723 -5080
rect 6647 -5174 6723 -5126
rect 4013 -5268 4089 -5220
rect 4013 -5314 4028 -5268
rect 4074 -5314 4089 -5268
rect 6647 -5220 6662 -5174
rect 6708 -5220 6723 -5174
rect 6647 -5268 6723 -5220
rect 4013 -5362 4089 -5314
rect 4013 -5408 4028 -5362
rect 4074 -5408 4089 -5362
rect 4013 -5456 4089 -5408
rect 4013 -5502 4028 -5456
rect 4074 -5502 4089 -5456
rect 4013 -5550 4089 -5502
rect 4013 -5596 4028 -5550
rect 4074 -5596 4089 -5550
rect 4013 -5644 4089 -5596
rect 4013 -5690 4028 -5644
rect 4074 -5690 4089 -5644
rect 4013 -5738 4089 -5690
rect 4013 -5784 4028 -5738
rect 4074 -5784 4089 -5738
rect 6647 -5314 6662 -5268
rect 6708 -5314 6723 -5268
rect 6647 -5362 6723 -5314
rect 6647 -5408 6662 -5362
rect 6708 -5408 6723 -5362
rect 6647 -5456 6723 -5408
rect 6647 -5502 6662 -5456
rect 6708 -5502 6723 -5456
rect 6647 -5550 6723 -5502
rect 6647 -5596 6662 -5550
rect 6708 -5596 6723 -5550
rect 6647 -5644 6723 -5596
rect 6647 -5690 6662 -5644
rect 6708 -5690 6723 -5644
rect 6647 -5738 6723 -5690
rect 4013 -5832 4089 -5784
rect 4013 -5878 4028 -5832
rect 4074 -5878 4089 -5832
rect 4013 -5926 4089 -5878
rect 6647 -5784 6662 -5738
rect 6708 -5784 6723 -5738
rect 6647 -5832 6723 -5784
rect 6647 -5878 6662 -5832
rect 6708 -5878 6723 -5832
rect 4013 -5972 4028 -5926
rect 4074 -5972 4089 -5926
rect 4013 -6005 4089 -5972
rect 6647 -5926 6723 -5878
rect 6647 -5972 6662 -5926
rect 6708 -5972 6723 -5926
rect 6647 -6005 6723 -5972
rect 4013 -6020 6723 -6005
rect 4013 -6066 4029 -6020
rect 4075 -6066 4123 -6020
rect 4169 -6066 4217 -6020
rect 4263 -6066 4311 -6020
rect 4357 -6066 4405 -6020
rect 4451 -6066 4499 -6020
rect 4545 -6066 4593 -6020
rect 4639 -6066 4687 -6020
rect 4733 -6066 4781 -6020
rect 4827 -6066 4875 -6020
rect 4921 -6066 4969 -6020
rect 5015 -6066 5063 -6020
rect 5109 -6066 5157 -6020
rect 5203 -6066 5251 -6020
rect 5297 -6066 5345 -6020
rect 5391 -6066 5439 -6020
rect 5485 -6066 5533 -6020
rect 5579 -6066 5627 -6020
rect 5673 -6066 5721 -6020
rect 5767 -6066 5815 -6020
rect 5861 -6066 5909 -6020
rect 5955 -6066 6003 -6020
rect 6049 -6066 6097 -6020
rect 6143 -6066 6191 -6020
rect 6237 -6066 6285 -6020
rect 6331 -6066 6379 -6020
rect 6425 -6066 6473 -6020
rect 6519 -6066 6567 -6020
rect 6613 -6066 6661 -6020
rect 6707 -6066 6723 -6020
rect 4013 -6081 6723 -6066
rect 3676 -6151 3691 -6105
rect 3737 -6151 3752 -6105
rect 3676 -6184 3752 -6151
rect 1606 -6199 3752 -6184
rect 1606 -6245 1622 -6199
rect 1668 -6245 1716 -6199
rect 1762 -6245 1810 -6199
rect 1856 -6245 1904 -6199
rect 1950 -6245 1998 -6199
rect 2044 -6245 2092 -6199
rect 2138 -6245 2186 -6199
rect 2232 -6245 2280 -6199
rect 2326 -6245 2374 -6199
rect 2420 -6245 2468 -6199
rect 2514 -6245 2562 -6199
rect 2608 -6245 2656 -6199
rect 2702 -6245 2750 -6199
rect 2796 -6245 2844 -6199
rect 2890 -6245 2938 -6199
rect 2984 -6245 3032 -6199
rect 3078 -6245 3126 -6199
rect 3172 -6245 3220 -6199
rect 3266 -6245 3314 -6199
rect 3360 -6245 3408 -6199
rect 3454 -6245 3502 -6199
rect 3548 -6245 3596 -6199
rect 3642 -6245 3690 -6199
rect 3736 -6245 3752 -6199
rect 1606 -6260 3752 -6245
rect -477 -6297 1293 -6282
rect -3282 -6321 -1230 -6306
<< psubdiffcont >>
rect 8786 -4780 8832 -4734
rect 8884 -4780 8930 -4734
rect 8982 -4780 9028 -4734
rect 9080 -4780 9126 -4734
rect 9178 -4780 9224 -4734
rect 9276 -4780 9322 -4734
rect 9374 -4780 9420 -4734
rect 9472 -4780 9518 -4734
rect 9570 -4780 9616 -4734
rect 9668 -4780 9714 -4734
rect 9766 -4780 9812 -4734
rect 9864 -4780 9910 -4734
rect 9962 -4780 10008 -4734
rect 10060 -4780 10106 -4734
rect 10158 -4780 10204 -4734
rect 10256 -4780 10302 -4734
rect 10354 -4780 10400 -4734
rect 10452 -4780 10498 -4734
rect 10550 -4780 10596 -4734
rect 10648 -4780 10694 -4734
rect 10746 -4780 10792 -4734
rect 10844 -4780 10890 -4734
rect 10942 -4780 10988 -4734
rect 11040 -4780 11086 -4734
rect 8786 -4878 8832 -4832
rect 8786 -4976 8832 -4930
rect 11040 -4878 11086 -4832
rect 8786 -5074 8832 -5028
rect 11040 -4976 11086 -4930
rect 11040 -5074 11086 -5028
rect 8786 -5172 8832 -5126
rect 8786 -5270 8832 -5224
rect 8786 -5368 8832 -5322
rect 8786 -5466 8832 -5420
rect 8786 -5564 8832 -5518
rect 8786 -5662 8832 -5616
rect 8786 -5760 8832 -5714
rect 11040 -5172 11086 -5126
rect 11040 -5270 11086 -5224
rect 11040 -5368 11086 -5322
rect 11040 -5466 11086 -5420
rect 11040 -5564 11086 -5518
rect 11040 -5662 11086 -5616
rect 8786 -5858 8832 -5812
rect 11040 -5760 11086 -5714
rect 8786 -5956 8832 -5910
rect 8786 -6054 8832 -6008
rect 8786 -6152 8832 -6106
rect 8786 -6250 8832 -6204
rect 8786 -6348 8832 -6302
rect 8786 -6446 8832 -6400
rect -549 -6558 -503 -6512
rect -451 -6558 -405 -6512
rect -353 -6558 -307 -6512
rect -255 -6558 -209 -6512
rect -157 -6558 -111 -6512
rect -59 -6558 -13 -6512
rect 39 -6558 85 -6512
rect 137 -6558 183 -6512
rect 235 -6558 281 -6512
rect 333 -6558 379 -6512
rect 431 -6558 477 -6512
rect 529 -6558 575 -6512
rect 627 -6558 673 -6512
rect 725 -6558 771 -6512
rect 823 -6558 869 -6512
rect 921 -6558 967 -6512
rect 1019 -6558 1065 -6512
rect 1117 -6558 1163 -6512
rect 1215 -6558 1261 -6512
rect 11040 -5858 11086 -5812
rect 11040 -5956 11086 -5910
rect 11040 -6054 11086 -6008
rect 11040 -6152 11086 -6106
rect 11040 -6250 11086 -6204
rect 11040 -6348 11086 -6302
rect 11040 -6446 11086 -6400
rect 8786 -6544 8832 -6498
rect -549 -6656 -503 -6610
rect -549 -6754 -503 -6708
rect -3295 -6888 -3249 -6842
rect -3197 -6888 -3151 -6842
rect -3099 -6888 -3053 -6842
rect -3001 -6888 -2955 -6842
rect -2903 -6888 -2857 -6842
rect -2805 -6888 -2759 -6842
rect -2707 -6888 -2661 -6842
rect -2609 -6888 -2563 -6842
rect -2511 -6888 -2465 -6842
rect -2413 -6888 -2367 -6842
rect -2315 -6888 -2269 -6842
rect -2217 -6888 -2171 -6842
rect -2119 -6888 -2073 -6842
rect -2021 -6888 -1975 -6842
rect -1923 -6888 -1877 -6842
rect -1825 -6888 -1779 -6842
rect -1727 -6888 -1681 -6842
rect -1629 -6888 -1583 -6842
rect -1531 -6888 -1485 -6842
rect -1433 -6888 -1387 -6842
rect -1335 -6888 -1289 -6842
rect -1237 -6888 -1191 -6842
rect -3295 -6986 -3249 -6940
rect -3295 -7084 -3249 -7038
rect -1237 -6986 -1191 -6940
rect -3295 -7182 -3249 -7136
rect -1237 -7084 -1191 -7038
rect -3295 -7280 -3249 -7234
rect -3295 -7378 -3249 -7332
rect -3295 -7476 -3249 -7430
rect -3295 -7574 -3249 -7528
rect -3295 -7672 -3249 -7626
rect -3295 -7770 -3249 -7724
rect -1237 -7182 -1191 -7136
rect -1237 -7280 -1191 -7234
rect -1237 -7378 -1191 -7332
rect -1237 -7476 -1191 -7430
rect -1237 -7574 -1191 -7528
rect -1237 -7672 -1191 -7626
rect -3295 -7868 -3249 -7822
rect -1237 -7770 -1191 -7724
rect -3295 -7966 -3249 -7920
rect -1237 -7868 -1191 -7822
rect -3295 -8064 -3249 -8018
rect -3295 -8162 -3249 -8116
rect -3295 -8260 -3249 -8214
rect -3295 -8358 -3249 -8312
rect -3295 -8456 -3249 -8410
rect -3295 -8554 -3249 -8508
rect -1237 -7966 -1191 -7920
rect -1237 -8064 -1191 -8018
rect -1237 -8162 -1191 -8116
rect -1237 -8260 -1191 -8214
rect -1237 -8358 -1191 -8312
rect -1237 -8456 -1191 -8410
rect -3295 -8652 -3249 -8606
rect -1237 -8554 -1191 -8508
rect -3295 -8750 -3249 -8704
rect -1237 -8652 -1191 -8606
rect -3295 -8848 -3249 -8802
rect -3295 -8946 -3249 -8900
rect -3295 -9044 -3249 -8998
rect -3295 -9142 -3249 -9096
rect -3295 -9240 -3249 -9194
rect -3295 -9338 -3249 -9292
rect -1237 -8750 -1191 -8704
rect -1237 -8848 -1191 -8802
rect -1237 -8946 -1191 -8900
rect -1237 -9044 -1191 -8998
rect -1237 -9142 -1191 -9096
rect -1237 -9240 -1191 -9194
rect -3295 -9436 -3249 -9390
rect -1237 -9338 -1191 -9292
rect -3295 -9534 -3249 -9488
rect -1237 -9436 -1191 -9390
rect -1237 -9534 -1191 -9488
rect -3295 -9632 -3249 -9586
rect -3295 -9730 -3249 -9684
rect -3295 -9828 -3249 -9782
rect -3295 -9926 -3249 -9880
rect -3295 -10024 -3249 -9978
rect -3295 -10122 -3249 -10076
rect -1237 -9632 -1191 -9586
rect -1237 -9730 -1191 -9684
rect -1237 -9828 -1191 -9782
rect -1237 -9926 -1191 -9880
rect -1237 -10024 -1191 -9978
rect -1237 -10122 -1191 -10076
rect -3295 -10220 -3249 -10174
rect -3295 -10318 -3249 -10272
rect -1237 -10220 -1191 -10174
rect -1237 -10318 -1191 -10272
rect -3295 -10416 -3249 -10370
rect -3197 -10416 -3151 -10370
rect -3099 -10416 -3053 -10370
rect -3001 -10416 -2955 -10370
rect -2903 -10416 -2857 -10370
rect -2805 -10416 -2759 -10370
rect -2707 -10416 -2661 -10370
rect -2609 -10416 -2563 -10370
rect -2511 -10416 -2465 -10370
rect -2413 -10416 -2367 -10370
rect -2315 -10416 -2269 -10370
rect -2217 -10416 -2171 -10370
rect -2119 -10416 -2073 -10370
rect -2021 -10416 -1975 -10370
rect -1923 -10416 -1877 -10370
rect -1825 -10416 -1779 -10370
rect -1727 -10416 -1681 -10370
rect -1629 -10416 -1583 -10370
rect -1531 -10416 -1485 -10370
rect -1433 -10416 -1387 -10370
rect -1335 -10416 -1289 -10370
rect -1237 -10416 -1191 -10370
rect -549 -6852 -503 -6806
rect 1215 -6656 1261 -6610
rect 1215 -6754 1261 -6708
rect -549 -6950 -503 -6904
rect 1215 -6852 1261 -6806
rect -549 -7048 -503 -7002
rect -549 -7146 -503 -7100
rect -549 -7244 -503 -7198
rect -549 -7342 -503 -7296
rect -549 -7440 -503 -7394
rect -549 -7538 -503 -7492
rect -549 -7636 -503 -7590
rect 1215 -6950 1261 -6904
rect 1215 -7048 1261 -7002
rect 1215 -7146 1261 -7100
rect 1215 -7244 1261 -7198
rect 1215 -7342 1261 -7296
rect 1215 -7440 1261 -7394
rect 1215 -7538 1261 -7492
rect -549 -7734 -503 -7688
rect -549 -7832 -503 -7786
rect 1215 -7636 1261 -7590
rect 1215 -7734 1261 -7688
rect 1612 -6608 1658 -6562
rect 1710 -6608 1756 -6562
rect 1808 -6608 1854 -6562
rect 1906 -6608 1952 -6562
rect 2004 -6608 2050 -6562
rect 2102 -6608 2148 -6562
rect 2200 -6608 2246 -6562
rect 2298 -6608 2344 -6562
rect 2396 -6608 2442 -6562
rect 2494 -6608 2540 -6562
rect 2592 -6608 2638 -6562
rect 2690 -6608 2736 -6562
rect 2788 -6608 2834 -6562
rect 2886 -6608 2932 -6562
rect 2984 -6608 3030 -6562
rect 3082 -6608 3128 -6562
rect 3180 -6608 3226 -6562
rect 3278 -6608 3324 -6562
rect 3376 -6608 3422 -6562
rect 3474 -6608 3520 -6562
rect 3572 -6608 3618 -6562
rect 3670 -6608 3716 -6562
rect 3768 -6608 3814 -6562
rect 3866 -6608 3912 -6562
rect 3964 -6608 4010 -6562
rect 4062 -6608 4108 -6562
rect 1612 -6706 1658 -6660
rect 4062 -6706 4108 -6660
rect 1612 -6802 1658 -6756
rect 1612 -6900 1658 -6854
rect 11040 -6544 11086 -6498
rect 8786 -6642 8832 -6596
rect 8786 -6740 8832 -6694
rect 4062 -6802 4108 -6756
rect 4062 -6900 4108 -6854
rect 1612 -6998 1658 -6952
rect 1612 -7096 1658 -7050
rect 1612 -7194 1658 -7148
rect 1612 -7292 1658 -7246
rect 4062 -6998 4108 -6952
rect 4062 -7096 4108 -7050
rect 4062 -7194 4108 -7148
rect 4062 -7292 4108 -7246
rect 1612 -7390 1658 -7344
rect 1612 -7488 1658 -7442
rect 4062 -7390 4108 -7344
rect 4062 -7488 4108 -7442
rect 1612 -7586 1658 -7540
rect 4062 -7586 4108 -7540
rect 1612 -7684 1658 -7638
rect 1710 -7684 1756 -7638
rect 1808 -7684 1854 -7638
rect 1906 -7684 1952 -7638
rect 2004 -7684 2050 -7638
rect 2102 -7684 2148 -7638
rect 2200 -7684 2246 -7638
rect 2298 -7684 2344 -7638
rect 2396 -7684 2442 -7638
rect 2494 -7684 2540 -7638
rect 2592 -7684 2638 -7638
rect 2690 -7684 2736 -7638
rect 2788 -7684 2834 -7638
rect 2886 -7684 2932 -7638
rect 2984 -7684 3030 -7638
rect 3082 -7684 3128 -7638
rect 3180 -7684 3226 -7638
rect 3278 -7684 3324 -7638
rect 3376 -7684 3422 -7638
rect 3474 -7684 3520 -7638
rect 3572 -7684 3618 -7638
rect 3670 -7684 3716 -7638
rect 3768 -7684 3814 -7638
rect 3866 -7684 3912 -7638
rect 3964 -7684 4010 -7638
rect 4062 -7684 4108 -7638
rect 4399 -6812 4445 -6766
rect 4497 -6811 4543 -6765
rect 4595 -6811 4641 -6765
rect 4693 -6811 4739 -6765
rect 4791 -6811 4837 -6765
rect 4889 -6811 4935 -6765
rect 4987 -6811 5033 -6765
rect 5085 -6811 5131 -6765
rect 5183 -6811 5229 -6765
rect 5281 -6811 5327 -6765
rect 5379 -6811 5425 -6765
rect 5477 -6811 5523 -6765
rect 5575 -6811 5621 -6765
rect 5673 -6811 5719 -6765
rect 5771 -6811 5817 -6765
rect 5869 -6811 5915 -6765
rect 5967 -6811 6013 -6765
rect 6065 -6811 6111 -6765
rect 6163 -6811 6209 -6765
rect 6261 -6811 6307 -6765
rect 6359 -6811 6405 -6765
rect 6457 -6811 6503 -6765
rect 6555 -6811 6601 -6765
rect 6653 -6811 6699 -6765
rect 6751 -6811 6797 -6765
rect 6849 -6811 6895 -6765
rect 6947 -6811 6993 -6765
rect 7045 -6811 7091 -6765
rect 7143 -6811 7189 -6765
rect 7241 -6811 7287 -6765
rect 7339 -6811 7385 -6765
rect 7437 -6811 7483 -6765
rect 7535 -6811 7581 -6765
rect 7633 -6811 7679 -6765
rect 7731 -6811 7777 -6765
rect 7829 -6811 7875 -6765
rect 7927 -6811 7973 -6765
rect 8025 -6811 8071 -6765
rect 4400 -6909 4446 -6863
rect 4400 -7007 4446 -6961
rect 4400 -7105 4446 -7059
rect 8026 -6910 8072 -6864
rect 8026 -7008 8072 -6962
rect 4400 -7203 4446 -7157
rect 4400 -7301 4446 -7255
rect 4400 -7399 4446 -7353
rect 4400 -7497 4446 -7451
rect 8026 -7106 8072 -7060
rect 8026 -7204 8072 -7158
rect 8026 -7302 8072 -7256
rect 8026 -7400 8072 -7354
rect 8026 -7498 8072 -7452
rect 4400 -7595 4446 -7549
rect 8786 -6838 8832 -6792
rect 8786 -6936 8832 -6890
rect 8786 -7034 8832 -6988
rect 8786 -7132 8832 -7086
rect 8786 -7230 8832 -7184
rect 11040 -6642 11086 -6596
rect 11040 -6740 11086 -6694
rect 11040 -6838 11086 -6792
rect 11040 -6936 11086 -6890
rect 11040 -7034 11086 -6988
rect 11040 -7132 11086 -7086
rect 8786 -7328 8832 -7282
rect 11040 -7230 11086 -7184
rect 11040 -7328 11086 -7282
rect 8786 -7426 8832 -7380
rect 11040 -7426 11086 -7380
rect 8786 -7524 8832 -7478
rect 8884 -7524 8930 -7478
rect 8982 -7524 9028 -7478
rect 9080 -7524 9126 -7478
rect 9178 -7524 9224 -7478
rect 9276 -7524 9322 -7478
rect 9374 -7524 9420 -7478
rect 9472 -7524 9518 -7478
rect 9570 -7524 9616 -7478
rect 9668 -7524 9714 -7478
rect 9766 -7524 9812 -7478
rect 9864 -7524 9910 -7478
rect 9962 -7524 10008 -7478
rect 10060 -7524 10106 -7478
rect 10158 -7524 10204 -7478
rect 10256 -7524 10302 -7478
rect 10354 -7524 10400 -7478
rect 10452 -7524 10498 -7478
rect 10550 -7524 10596 -7478
rect 10648 -7524 10694 -7478
rect 10746 -7524 10792 -7478
rect 10844 -7524 10890 -7478
rect 10942 -7524 10988 -7478
rect 11040 -7524 11086 -7478
rect 8026 -7596 8072 -7550
rect 4400 -7693 4446 -7647
rect -549 -7930 -503 -7884
rect -549 -8028 -503 -7982
rect -549 -8126 -503 -8080
rect -549 -8224 -503 -8178
rect -549 -8322 -503 -8276
rect -549 -8420 -503 -8374
rect -549 -8518 -503 -8472
rect 1215 -7832 1261 -7786
rect 1215 -7930 1261 -7884
rect 1215 -8028 1261 -7982
rect 1215 -8126 1261 -8080
rect 1215 -8224 1261 -8178
rect 1215 -8322 1261 -8276
rect 4400 -7791 4446 -7745
rect 4400 -7889 4446 -7843
rect 4400 -7987 4446 -7941
rect 4400 -8085 4446 -8039
rect 8026 -7694 8072 -7648
rect 8026 -7792 8072 -7746
rect 8026 -7890 8072 -7844
rect 8026 -7988 8072 -7942
rect 4400 -8183 4446 -8137
rect 8026 -8086 8072 -8040
rect 4400 -8281 4446 -8235
rect 1215 -8420 1261 -8374
rect -549 -8616 -503 -8570
rect -549 -8714 -503 -8668
rect -549 -8812 -503 -8766
rect 1215 -8518 1261 -8472
rect 1215 -8616 1261 -8570
rect 1215 -8714 1261 -8668
rect -549 -8910 -503 -8864
rect -549 -9008 -503 -8962
rect -549 -9106 -503 -9060
rect -549 -9204 -503 -9158
rect -549 -9302 -503 -9256
rect -549 -9400 -503 -9354
rect -549 -9498 -503 -9452
rect 1215 -8812 1261 -8766
rect 1215 -8910 1261 -8864
rect 1215 -9008 1261 -8962
rect 1215 -9106 1261 -9060
rect 1215 -9204 1261 -9158
rect 1215 -9302 1261 -9256
rect 1215 -9400 1261 -9354
rect -549 -9596 -503 -9550
rect 1215 -9498 1261 -9452
rect 1215 -9596 1261 -9550
rect -549 -9694 -503 -9648
rect -549 -9792 -503 -9746
rect -549 -9890 -503 -9844
rect -549 -9988 -503 -9942
rect -549 -10086 -503 -10040
rect -549 -10184 -503 -10138
rect -549 -10282 -503 -10236
rect 1215 -9694 1261 -9648
rect 1215 -9792 1261 -9746
rect 1215 -9890 1261 -9844
rect 1215 -9988 1261 -9942
rect 1215 -10086 1261 -10040
rect 1215 -10184 1261 -10138
rect 1215 -10282 1261 -10236
rect -549 -10380 -503 -10334
rect 1215 -10380 1261 -10334
rect -549 -10478 -503 -10432
rect -549 -10576 -503 -10530
rect 1636 -8342 1682 -8296
rect 1734 -8343 1780 -8297
rect 1832 -8343 1878 -8297
rect 1930 -8343 1976 -8297
rect 2028 -8343 2074 -8297
rect 2126 -8343 2172 -8297
rect 2224 -8343 2270 -8297
rect 2322 -8343 2368 -8297
rect 2420 -8343 2466 -8297
rect 2518 -8343 2564 -8297
rect 2616 -8343 2662 -8297
rect 2714 -8343 2760 -8297
rect 2812 -8343 2858 -8297
rect 2910 -8342 2956 -8296
rect 1636 -8440 1682 -8394
rect 1636 -8538 1682 -8492
rect 1636 -8636 1682 -8590
rect 1636 -8734 1682 -8688
rect 1636 -8832 1682 -8786
rect 1636 -8930 1682 -8884
rect 1636 -9028 1682 -8982
rect 1636 -9126 1682 -9080
rect 2910 -8440 2956 -8394
rect 2910 -8538 2956 -8492
rect 2910 -8636 2956 -8590
rect 2910 -8734 2956 -8688
rect 2910 -8832 2956 -8786
rect 2910 -8930 2956 -8884
rect 2910 -9028 2956 -8982
rect 4400 -8379 4446 -8333
rect 4400 -8477 4446 -8431
rect 4400 -8575 4446 -8529
rect 8026 -8184 8072 -8138
rect 8026 -8282 8072 -8236
rect 8026 -8380 8072 -8334
rect 8026 -8478 8072 -8432
rect 8026 -8576 8072 -8530
rect 4400 -8673 4446 -8627
rect 4400 -8771 4446 -8725
rect 8026 -8674 8072 -8628
rect 8026 -8772 8072 -8726
rect 4400 -8869 4446 -8823
rect 8026 -8870 8072 -8824
rect 4399 -8967 4445 -8921
rect 4497 -8968 4543 -8922
rect 4595 -8968 4641 -8922
rect 4693 -8968 4739 -8922
rect 4791 -8968 4837 -8922
rect 4889 -8968 4935 -8922
rect 4987 -8968 5033 -8922
rect 5085 -8968 5131 -8922
rect 5183 -8968 5229 -8922
rect 5281 -8968 5327 -8922
rect 5379 -8968 5425 -8922
rect 5477 -8968 5523 -8922
rect 5575 -8968 5621 -8922
rect 5673 -8968 5719 -8922
rect 5771 -8968 5817 -8922
rect 5869 -8968 5915 -8922
rect 5967 -8968 6013 -8922
rect 6065 -8968 6111 -8922
rect 6163 -8968 6209 -8922
rect 6261 -8968 6307 -8922
rect 6359 -8968 6405 -8922
rect 6457 -8968 6503 -8922
rect 6555 -8968 6601 -8922
rect 6653 -8968 6699 -8922
rect 6751 -8968 6797 -8922
rect 6849 -8968 6895 -8922
rect 6947 -8968 6993 -8922
rect 7045 -8968 7091 -8922
rect 7143 -8968 7189 -8922
rect 7241 -8968 7287 -8922
rect 7339 -8968 7385 -8922
rect 7437 -8968 7483 -8922
rect 7535 -8968 7581 -8922
rect 7633 -8968 7679 -8922
rect 7731 -8968 7777 -8922
rect 7829 -8968 7875 -8922
rect 7927 -8968 7973 -8922
rect 8025 -8968 8071 -8922
rect 8786 -7780 8832 -7734
rect 8884 -7780 8930 -7734
rect 8982 -7780 9028 -7734
rect 9080 -7780 9126 -7734
rect 9178 -7780 9224 -7734
rect 9276 -7780 9322 -7734
rect 9374 -7780 9420 -7734
rect 9472 -7780 9518 -7734
rect 9570 -7780 9616 -7734
rect 9668 -7780 9714 -7734
rect 9766 -7780 9812 -7734
rect 9864 -7780 9910 -7734
rect 9962 -7780 10008 -7734
rect 10060 -7780 10106 -7734
rect 10158 -7780 10204 -7734
rect 10256 -7780 10302 -7734
rect 10354 -7780 10400 -7734
rect 10452 -7780 10498 -7734
rect 10550 -7780 10596 -7734
rect 10648 -7780 10694 -7734
rect 10746 -7780 10792 -7734
rect 10844 -7780 10890 -7734
rect 10942 -7780 10988 -7734
rect 11040 -7780 11086 -7734
rect 8786 -7878 8832 -7832
rect 8786 -7976 8832 -7930
rect 11040 -7878 11086 -7832
rect 8786 -8074 8832 -8028
rect 11040 -7976 11086 -7930
rect 11040 -8074 11086 -8028
rect 8786 -8172 8832 -8126
rect 8786 -8270 8832 -8224
rect 8786 -8368 8832 -8322
rect 8786 -8466 8832 -8420
rect 8786 -8564 8832 -8518
rect 8786 -8662 8832 -8616
rect 8786 -8760 8832 -8714
rect 11040 -8172 11086 -8126
rect 11040 -8270 11086 -8224
rect 11040 -8368 11086 -8322
rect 11040 -8466 11086 -8420
rect 11040 -8564 11086 -8518
rect 11040 -8662 11086 -8616
rect 8786 -8858 8832 -8812
rect 11040 -8760 11086 -8714
rect 8786 -8956 8832 -8910
rect 2910 -9126 2956 -9080
rect 1636 -9224 1682 -9178
rect 1636 -9322 1682 -9276
rect 1636 -9420 1682 -9374
rect 1636 -9518 1682 -9472
rect 2910 -9224 2956 -9178
rect 2910 -9322 2956 -9276
rect 2910 -9420 2956 -9374
rect 1636 -9616 1682 -9570
rect 2910 -9518 2956 -9472
rect 1636 -9714 1682 -9668
rect 1636 -9812 1682 -9766
rect 1636 -9910 1682 -9864
rect 1636 -10008 1682 -9962
rect 1636 -10106 1682 -10060
rect 1636 -10204 1682 -10158
rect 1636 -10302 1682 -10256
rect 2910 -9616 2956 -9570
rect 2910 -9714 2956 -9668
rect 2910 -9812 2956 -9766
rect 2910 -9910 2956 -9864
rect 2910 -10008 2956 -9962
rect 2910 -10106 2956 -10060
rect 2910 -10204 2956 -10158
rect 2910 -10302 2956 -10256
rect 1636 -10400 1682 -10354
rect 1734 -10400 1780 -10354
rect 1832 -10400 1878 -10354
rect 1930 -10400 1976 -10354
rect 2028 -10400 2074 -10354
rect 2126 -10400 2172 -10354
rect 2224 -10400 2270 -10354
rect 2322 -10400 2368 -10354
rect 2420 -10400 2466 -10354
rect 2518 -10400 2564 -10354
rect 2616 -10400 2662 -10354
rect 2714 -10400 2760 -10354
rect 2812 -10400 2858 -10354
rect 2910 -10400 2956 -10354
rect 8786 -9054 8832 -9008
rect 8786 -9152 8832 -9106
rect 8786 -9250 8832 -9204
rect 8786 -9348 8832 -9302
rect 8786 -9446 8832 -9400
rect 11040 -8858 11086 -8812
rect 11040 -8956 11086 -8910
rect 11040 -9054 11086 -9008
rect 11040 -9152 11086 -9106
rect 11040 -9250 11086 -9204
rect 11040 -9348 11086 -9302
rect 11040 -9446 11086 -9400
rect 8786 -9544 8832 -9498
rect 11040 -9544 11086 -9498
rect 8786 -9642 8832 -9596
rect 8786 -9740 8832 -9694
rect 8786 -9838 8832 -9792
rect 8786 -9936 8832 -9890
rect 8786 -10034 8832 -9988
rect 8786 -10132 8832 -10086
rect 8786 -10230 8832 -10184
rect 11040 -9642 11086 -9596
rect 11040 -9740 11086 -9694
rect 11040 -9838 11086 -9792
rect 11040 -9936 11086 -9890
rect 11040 -10034 11086 -9988
rect 11040 -10132 11086 -10086
rect 8786 -10328 8832 -10282
rect 11040 -10230 11086 -10184
rect 11040 -10328 11086 -10282
rect 1215 -10478 1261 -10432
rect 1215 -10576 1261 -10530
rect 8786 -10426 8832 -10380
rect 11040 -10426 11086 -10380
rect 8786 -10524 8832 -10478
rect 8884 -10524 8930 -10478
rect 8982 -10524 9028 -10478
rect 9080 -10524 9126 -10478
rect 9178 -10524 9224 -10478
rect 9276 -10524 9322 -10478
rect 9374 -10524 9420 -10478
rect 9472 -10524 9518 -10478
rect 9570 -10524 9616 -10478
rect 9668 -10524 9714 -10478
rect 9766 -10524 9812 -10478
rect 9864 -10524 9910 -10478
rect 9962 -10524 10008 -10478
rect 10060 -10524 10106 -10478
rect 10158 -10524 10204 -10478
rect 10256 -10524 10302 -10478
rect 10354 -10524 10400 -10478
rect 10452 -10524 10498 -10478
rect 10550 -10524 10596 -10478
rect 10648 -10524 10694 -10478
rect 10746 -10524 10792 -10478
rect 10844 -10524 10890 -10478
rect 10942 -10524 10988 -10478
rect 11040 -10524 11086 -10478
rect -549 -10674 -503 -10628
rect -451 -10674 -405 -10628
rect -353 -10674 -307 -10628
rect -255 -10674 -209 -10628
rect -157 -10674 -111 -10628
rect -59 -10674 -13 -10628
rect 39 -10674 85 -10628
rect 137 -10674 183 -10628
rect 235 -10674 281 -10628
rect 333 -10674 379 -10628
rect 431 -10674 477 -10628
rect 529 -10674 575 -10628
rect 627 -10674 673 -10628
rect 725 -10674 771 -10628
rect 823 -10674 869 -10628
rect 921 -10674 967 -10628
rect 1019 -10674 1065 -10628
rect 1117 -10674 1163 -10628
rect 1215 -10674 1261 -10628
<< nsubdiffcont >>
rect -3294 1394 -3247 1441
rect -3199 1395 -3153 1441
rect -3105 1395 -3059 1441
rect -3011 1395 -2965 1441
rect -2917 1395 -2871 1441
rect -2823 1395 -2777 1441
rect -2729 1395 -2683 1441
rect -2635 1395 -2589 1441
rect -2541 1395 -2495 1441
rect -2447 1395 -2401 1441
rect -2353 1395 -2307 1441
rect -2259 1395 -2213 1441
rect -2165 1395 -2119 1441
rect -2071 1395 -2025 1441
rect -1977 1395 -1931 1441
rect -1883 1395 -1837 1441
rect -1789 1395 -1743 1441
rect -1695 1395 -1649 1441
rect -1601 1395 -1555 1441
rect -1507 1395 -1461 1441
rect -1413 1395 -1367 1441
rect -1319 1394 -1272 1441
rect -3294 1300 -3248 1346
rect -1318 1300 -1272 1346
rect -3294 1206 -3248 1252
rect -1318 1206 -1272 1252
rect -3294 1112 -3248 1158
rect -3294 1018 -3248 1064
rect -3294 924 -3248 970
rect -3294 830 -3248 876
rect -3294 736 -3248 782
rect -3294 642 -3248 688
rect -3294 548 -3248 594
rect -1318 1112 -1272 1158
rect -1318 1018 -1272 1064
rect 2377 1109 2423 1155
rect 2471 1109 2517 1155
rect 2565 1109 2611 1155
rect 2659 1109 2705 1155
rect 2753 1109 2799 1155
rect 2847 1109 2893 1155
rect 2941 1109 2987 1155
rect 3035 1109 3081 1155
rect 3129 1109 3175 1155
rect 3223 1109 3269 1155
rect 3317 1109 3363 1155
rect 3411 1109 3457 1155
rect 3505 1109 3551 1155
rect 3599 1109 3645 1155
rect 3693 1109 3739 1155
rect 3787 1109 3833 1155
rect 3881 1109 3927 1155
rect 3975 1109 4021 1155
rect 4069 1109 4115 1155
rect 4163 1109 4209 1155
rect 4257 1109 4303 1155
rect 4351 1109 4397 1155
rect 4445 1109 4491 1155
rect 4539 1109 4585 1155
rect 4633 1109 4679 1155
rect -1318 924 -1272 970
rect -1318 830 -1272 876
rect -1318 736 -1272 782
rect -1318 642 -1272 688
rect -1318 548 -1272 594
rect -3294 454 -3248 500
rect -1318 454 -1272 500
rect -3294 360 -3248 406
rect -3294 266 -3248 312
rect -3294 172 -3248 218
rect -3294 78 -3248 124
rect -3294 -16 -3248 30
rect -3294 -110 -3248 -64
rect -3294 -204 -3248 -158
rect -1318 360 -1272 406
rect -1318 266 -1272 312
rect -1318 172 -1272 218
rect -1318 78 -1272 124
rect -1318 -16 -1272 30
rect -1318 -110 -1272 -64
rect -1318 -204 -1272 -158
rect -3294 -298 -3248 -252
rect -3294 -392 -3248 -346
rect -3294 -486 -3248 -440
rect -3294 -580 -3248 -534
rect -3294 -674 -3248 -628
rect -3294 -768 -3248 -722
rect -3294 -862 -3248 -816
rect -3294 -956 -3248 -910
rect -1318 -298 -1272 -252
rect -1318 -392 -1272 -346
rect -1318 -486 -1272 -440
rect -1318 -580 -1272 -534
rect -1318 -674 -1272 -628
rect -1318 -768 -1272 -722
rect -1318 -862 -1272 -816
rect -3294 -1050 -3248 -1004
rect -1318 -956 -1272 -910
rect -3294 -1144 -3248 -1098
rect -3294 -1238 -3248 -1192
rect -3294 -1332 -3248 -1286
rect -3294 -1426 -3248 -1380
rect -3294 -1520 -3248 -1474
rect -3294 -1614 -3248 -1568
rect -3294 -1708 -3248 -1662
rect -3294 -1802 -3248 -1756
rect -3294 -1896 -3248 -1850
rect -1318 -1050 -1272 -1004
rect -1318 -1144 -1272 -1098
rect -1318 -1238 -1272 -1192
rect -1318 -1332 -1272 -1286
rect -1318 -1426 -1272 -1380
rect -1318 -1520 -1272 -1474
rect -1318 -1614 -1272 -1568
rect -1318 -1708 -1272 -1662
rect -1318 -1802 -1272 -1756
rect -1318 -1896 -1272 -1850
rect -3293 -1990 -3247 -1944
rect -3199 -1990 -3153 -1944
rect -3105 -1990 -3059 -1944
rect -3011 -1990 -2965 -1944
rect -2917 -1990 -2871 -1944
rect -2823 -1990 -2777 -1944
rect -2729 -1990 -2683 -1944
rect -2635 -1990 -2589 -1944
rect -2541 -1990 -2495 -1944
rect -2447 -1990 -2401 -1944
rect -2353 -1990 -2307 -1944
rect -2259 -1990 -2213 -1944
rect -2165 -1990 -2119 -1944
rect -2071 -1990 -2025 -1944
rect -1977 -1990 -1931 -1944
rect -1883 -1990 -1837 -1944
rect -1789 -1990 -1743 -1944
rect -1695 -1990 -1649 -1944
rect -1601 -1990 -1555 -1944
rect -1507 -1990 -1461 -1944
rect -1413 -1990 -1367 -1944
rect -1319 -1990 -1273 -1944
rect -747 967 -701 1013
rect -653 967 -607 1013
rect -552 967 -506 1013
rect -458 967 -412 1013
rect -362 967 -316 1013
rect -268 967 -222 1013
rect -167 967 -121 1013
rect -73 967 -27 1013
rect 21 967 67 1013
rect 115 967 161 1013
rect 216 967 262 1013
rect 310 967 356 1013
rect 406 967 452 1013
rect 500 967 546 1013
rect 601 967 647 1013
rect 695 967 741 1013
rect 789 967 835 1013
rect 883 967 929 1013
rect 984 967 1030 1013
rect 1078 967 1124 1013
rect 1172 967 1218 1013
rect -747 871 -701 917
rect 1172 871 1218 917
rect -747 777 -701 823
rect 1172 770 1218 816
rect -747 681 -701 727
rect -747 587 -701 633
rect -747 493 -701 539
rect -747 392 -701 438
rect -747 298 -701 344
rect -747 202 -701 248
rect -747 108 -701 154
rect 1172 676 1218 722
rect 1172 582 1218 628
rect 1172 488 1218 534
rect 1172 387 1218 433
rect 1172 293 1218 339
rect 1172 197 1218 243
rect 1172 103 1218 149
rect -747 7 -701 53
rect -747 -87 -701 -41
rect -747 -181 -701 -135
rect -747 -275 -701 -229
rect 1172 2 1218 48
rect 1172 -92 1218 -46
rect 1172 -186 1218 -140
rect 1172 -280 1218 -234
rect -747 -376 -701 -330
rect -747 -470 -701 -424
rect -747 -566 -701 -520
rect -747 -660 -701 -614
rect -747 -761 -701 -715
rect -747 -855 -701 -809
rect -747 -949 -701 -903
rect 1172 -381 1218 -335
rect 1172 -475 1218 -429
rect 1172 -571 1218 -525
rect 1172 -665 1218 -619
rect 1172 -766 1218 -720
rect 1172 -860 1218 -814
rect 1172 -954 1218 -908
rect -747 -1043 -701 -997
rect -747 -1144 -701 -1098
rect -747 -1238 -701 -1192
rect -747 -1334 -701 -1288
rect 1172 -1050 1218 -1004
rect 1172 -1144 1218 -1098
rect 1172 -1245 1218 -1199
rect -747 -1428 -701 -1382
rect -747 -1522 -701 -1476
rect -747 -1623 -701 -1577
rect -747 -1717 -701 -1671
rect -747 -1813 -701 -1767
rect -747 -1907 -701 -1861
rect -747 -2008 -701 -1962
rect 1172 -1339 1218 -1293
rect 1172 -1433 1218 -1387
rect 1172 -1527 1218 -1481
rect 1172 -1628 1218 -1582
rect 1172 -1722 1218 -1676
rect 1172 -1818 1218 -1772
rect 1172 -1912 1218 -1866
rect -747 -2102 -701 -2056
rect -747 -2196 -701 -2150
rect -747 -2290 -701 -2244
rect -747 -2391 -701 -2345
rect 1172 -2013 1218 -1967
rect 1172 -2107 1218 -2061
rect 1172 -2201 1218 -2155
rect 1172 -2295 1218 -2249
rect -747 -2485 -701 -2439
rect -3267 -2640 -3220 -2593
rect -3172 -2639 -3126 -2593
rect -3078 -2639 -3032 -2593
rect -2984 -2639 -2938 -2593
rect -2890 -2639 -2844 -2593
rect -2796 -2639 -2750 -2593
rect -2702 -2639 -2656 -2593
rect -2608 -2639 -2562 -2593
rect -2514 -2639 -2468 -2593
rect -2420 -2639 -2374 -2593
rect -2326 -2639 -2280 -2593
rect -2232 -2639 -2186 -2593
rect -2138 -2639 -2092 -2593
rect -2044 -2639 -1998 -2593
rect -1950 -2639 -1904 -2593
rect -1856 -2639 -1810 -2593
rect -1762 -2639 -1716 -2593
rect -1668 -2639 -1622 -2593
rect -1574 -2639 -1528 -2593
rect -1480 -2639 -1434 -2593
rect -1386 -2639 -1340 -2593
rect -1292 -2640 -1245 -2593
rect -3267 -2734 -3221 -2688
rect -3267 -2828 -3221 -2782
rect -1291 -2734 -1245 -2688
rect -1291 -2828 -1245 -2782
rect -3267 -2922 -3221 -2876
rect -1291 -2922 -1245 -2876
rect -3267 -3016 -3221 -2970
rect -1291 -3016 -1245 -2970
rect -3267 -3110 -3221 -3064
rect -3267 -3204 -3221 -3158
rect -3267 -3298 -3221 -3252
rect -3267 -3392 -3221 -3346
rect -3267 -3486 -3221 -3440
rect -1291 -3110 -1245 -3064
rect -1291 -3204 -1245 -3158
rect -1291 -3298 -1245 -3252
rect -1291 -3392 -1245 -3346
rect -747 -2581 -701 -2535
rect -747 -2675 -701 -2629
rect -747 -2776 -701 -2730
rect -747 -2870 -701 -2824
rect -747 -2964 -701 -2918
rect -747 -3058 -701 -3012
rect 1172 -2396 1218 -2350
rect 1172 -2490 1218 -2444
rect 1172 -2586 1218 -2540
rect 1172 -2680 1218 -2634
rect 1172 -2781 1218 -2735
rect 1172 -2875 1218 -2829
rect 1172 -2969 1218 -2923
rect 2376 1015 2422 1061
rect 4634 1015 4680 1061
rect 2376 921 2422 967
rect 2376 827 2422 873
rect 2376 733 2422 779
rect 2376 639 2422 685
rect 2376 545 2422 591
rect 2376 451 2422 497
rect 2376 357 2422 403
rect 2376 263 2422 309
rect 4634 921 4680 967
rect 4634 827 4680 873
rect 4634 733 4680 779
rect 4634 639 4680 685
rect 4634 545 4680 591
rect 4634 451 4680 497
rect 4634 357 4680 403
rect 4634 263 4680 309
rect 2376 169 2422 215
rect 4634 169 4680 215
rect 2376 75 2422 121
rect 2376 -19 2422 27
rect 2376 -113 2422 -67
rect 2376 -207 2422 -161
rect 2376 -301 2422 -255
rect 2376 -395 2422 -349
rect 2376 -489 2422 -443
rect 4634 75 4680 121
rect 4634 -19 4680 27
rect 4634 -113 4680 -67
rect 4634 -207 4680 -161
rect 4634 -301 4680 -255
rect 4634 -395 4680 -349
rect 4634 -489 4680 -443
rect 2376 -583 2422 -537
rect 4634 -583 4680 -537
rect 2376 -677 2422 -631
rect 2376 -771 2422 -725
rect 2376 -865 2422 -819
rect 2376 -959 2422 -913
rect 2376 -1053 2422 -1007
rect 2376 -1147 2422 -1101
rect 2376 -1241 2422 -1195
rect 4634 -677 4680 -631
rect 4634 -771 4680 -725
rect 4634 -865 4680 -819
rect 4634 -959 4680 -913
rect 4634 -1053 4680 -1007
rect 4634 -1147 4680 -1101
rect 4634 -1241 4680 -1195
rect 2376 -1335 2422 -1289
rect 4634 -1335 4680 -1289
rect 2376 -1429 2422 -1383
rect 2376 -1523 2422 -1477
rect 2376 -1617 2422 -1571
rect 2376 -1711 2422 -1665
rect 2376 -1805 2422 -1759
rect 2376 -1899 2422 -1853
rect 2376 -1993 2422 -1947
rect 4634 -1429 4680 -1383
rect 4634 -1523 4680 -1477
rect 4634 -1617 4680 -1571
rect 4634 -1711 4680 -1665
rect 4634 -1805 4680 -1759
rect 4634 -1899 4680 -1853
rect 2376 -2087 2422 -2041
rect 4634 -1993 4680 -1947
rect 2376 -2181 2422 -2135
rect 2376 -2275 2422 -2229
rect 2376 -2369 2422 -2323
rect 2376 -2463 2422 -2417
rect 2376 -2557 2422 -2511
rect 2376 -2651 2422 -2605
rect 2376 -2745 2422 -2699
rect 2376 -2839 2422 -2793
rect 4634 -2087 4680 -2041
rect 4634 -2181 4680 -2135
rect 4634 -2275 4680 -2229
rect 4634 -2369 4680 -2323
rect 4634 -2463 4680 -2417
rect 4634 -2557 4680 -2511
rect 4634 -2651 4680 -2605
rect 4634 -2745 4680 -2699
rect 4634 -2839 4680 -2793
rect 2377 -2933 2423 -2887
rect 2471 -2933 2517 -2887
rect 2565 -2933 2611 -2887
rect 2659 -2933 2705 -2887
rect 2753 -2933 2799 -2887
rect 2847 -2933 2893 -2887
rect 2941 -2933 2987 -2887
rect 3035 -2933 3081 -2887
rect 3129 -2933 3175 -2887
rect 3223 -2933 3269 -2887
rect 3317 -2933 3363 -2887
rect 3411 -2933 3457 -2887
rect 3505 -2933 3551 -2887
rect 3599 -2933 3645 -2887
rect 3693 -2933 3739 -2887
rect 3787 -2933 3833 -2887
rect 3881 -2933 3927 -2887
rect 3975 -2933 4021 -2887
rect 4069 -2933 4115 -2887
rect 4163 -2933 4209 -2887
rect 4257 -2933 4303 -2887
rect 4351 -2933 4397 -2887
rect 4445 -2933 4491 -2887
rect 4539 -2933 4585 -2887
rect 4633 -2933 4679 -2887
rect 5177 1109 5223 1155
rect 5271 1109 5317 1155
rect 5365 1109 5411 1155
rect 5459 1109 5505 1155
rect 5553 1109 5599 1155
rect 5647 1109 5693 1155
rect 5741 1109 5787 1155
rect 5835 1109 5881 1155
rect 5929 1109 5975 1155
rect 6023 1109 6069 1155
rect 6117 1109 6163 1155
rect 6211 1109 6257 1155
rect 6305 1109 6351 1155
rect 6399 1109 6445 1155
rect 6493 1109 6539 1155
rect 6587 1109 6633 1155
rect 6681 1109 6727 1155
rect 6775 1109 6821 1155
rect 6869 1109 6915 1155
rect 6963 1109 7009 1155
rect 7057 1109 7103 1155
rect 7151 1109 7197 1155
rect 7245 1109 7291 1155
rect 7339 1109 7385 1155
rect 7433 1109 7479 1155
rect 5176 1015 5222 1061
rect 7434 1015 7480 1061
rect 5176 921 5222 967
rect 5176 827 5222 873
rect 5176 733 5222 779
rect 5176 639 5222 685
rect 5176 545 5222 591
rect 5176 451 5222 497
rect 5176 357 5222 403
rect 5176 263 5222 309
rect 7434 921 7480 967
rect 7434 827 7480 873
rect 7434 733 7480 779
rect 7434 639 7480 685
rect 7434 545 7480 591
rect 7434 451 7480 497
rect 7434 357 7480 403
rect 7434 263 7480 309
rect 5176 169 5222 215
rect 7434 169 7480 215
rect 5176 75 5222 121
rect 5176 -19 5222 27
rect 5176 -113 5222 -67
rect 5176 -207 5222 -161
rect 5176 -301 5222 -255
rect 5176 -395 5222 -349
rect 5176 -489 5222 -443
rect 7434 75 7480 121
rect 7434 -19 7480 27
rect 7434 -113 7480 -67
rect 7434 -207 7480 -161
rect 7434 -301 7480 -255
rect 7434 -395 7480 -349
rect 7434 -489 7480 -443
rect 5176 -583 5222 -537
rect 7434 -583 7480 -537
rect 5176 -677 5222 -631
rect 5176 -771 5222 -725
rect 5176 -865 5222 -819
rect 5176 -959 5222 -913
rect 5176 -1053 5222 -1007
rect 5176 -1147 5222 -1101
rect 5176 -1241 5222 -1195
rect 7434 -677 7480 -631
rect 7434 -771 7480 -725
rect 7434 -865 7480 -819
rect 7434 -959 7480 -913
rect 7434 -1053 7480 -1007
rect 7434 -1147 7480 -1101
rect 7434 -1241 7480 -1195
rect 5176 -1335 5222 -1289
rect 7434 -1335 7480 -1289
rect 5176 -1429 5222 -1383
rect 5176 -1523 5222 -1477
rect 5176 -1617 5222 -1571
rect 5176 -1711 5222 -1665
rect 5176 -1805 5222 -1759
rect 5176 -1899 5222 -1853
rect 5176 -1993 5222 -1947
rect 7434 -1429 7480 -1383
rect 7434 -1523 7480 -1477
rect 7434 -1617 7480 -1571
rect 7434 -1711 7480 -1665
rect 7434 -1805 7480 -1759
rect 7434 -1899 7480 -1853
rect 5176 -2087 5222 -2041
rect 7434 -1993 7480 -1947
rect 5176 -2181 5222 -2135
rect 5176 -2275 5222 -2229
rect 5176 -2369 5222 -2323
rect 5176 -2463 5222 -2417
rect 5176 -2557 5222 -2511
rect 5176 -2651 5222 -2605
rect 5176 -2745 5222 -2699
rect 5176 -2839 5222 -2793
rect 7434 -2087 7480 -2041
rect 7434 -2181 7480 -2135
rect 7434 -2275 7480 -2229
rect 7434 -2369 7480 -2323
rect 7434 -2463 7480 -2417
rect 7434 -2557 7480 -2511
rect 7434 -2651 7480 -2605
rect 7434 -2745 7480 -2699
rect 7434 -2839 7480 -2793
rect 5177 -2933 5223 -2887
rect 5271 -2933 5317 -2887
rect 5365 -2933 5411 -2887
rect 5459 -2933 5505 -2887
rect 5553 -2933 5599 -2887
rect 5647 -2933 5693 -2887
rect 5741 -2933 5787 -2887
rect 5835 -2933 5881 -2887
rect 5929 -2933 5975 -2887
rect 6023 -2933 6069 -2887
rect 6117 -2933 6163 -2887
rect 6211 -2933 6257 -2887
rect 6305 -2933 6351 -2887
rect 6399 -2933 6445 -2887
rect 6493 -2933 6539 -2887
rect 6587 -2933 6633 -2887
rect 6681 -2933 6727 -2887
rect 6775 -2933 6821 -2887
rect 6869 -2933 6915 -2887
rect 6963 -2933 7009 -2887
rect 7057 -2933 7103 -2887
rect 7151 -2933 7197 -2887
rect 7245 -2933 7291 -2887
rect 7339 -2933 7385 -2887
rect 7433 -2933 7479 -2887
rect 7977 1109 8023 1155
rect 8071 1109 8117 1155
rect 8165 1109 8211 1155
rect 8259 1109 8305 1155
rect 8353 1109 8399 1155
rect 8447 1109 8493 1155
rect 8541 1109 8587 1155
rect 8635 1109 8681 1155
rect 8729 1109 8775 1155
rect 8823 1109 8869 1155
rect 8917 1109 8963 1155
rect 9011 1109 9057 1155
rect 9105 1109 9151 1155
rect 9199 1109 9245 1155
rect 9293 1109 9339 1155
rect 9387 1109 9433 1155
rect 9481 1109 9527 1155
rect 9575 1109 9621 1155
rect 9669 1109 9715 1155
rect 9763 1109 9809 1155
rect 9857 1109 9903 1155
rect 9951 1109 9997 1155
rect 10045 1109 10091 1155
rect 10139 1109 10185 1155
rect 10233 1109 10279 1155
rect 7976 1015 8022 1061
rect 10234 1015 10280 1061
rect 7976 921 8022 967
rect 7976 827 8022 873
rect 7976 733 8022 779
rect 7976 639 8022 685
rect 7976 545 8022 591
rect 7976 451 8022 497
rect 7976 357 8022 403
rect 7976 263 8022 309
rect 10234 921 10280 967
rect 10234 827 10280 873
rect 10234 733 10280 779
rect 10234 639 10280 685
rect 10234 545 10280 591
rect 10234 451 10280 497
rect 10234 357 10280 403
rect 10234 263 10280 309
rect 7976 169 8022 215
rect 10234 169 10280 215
rect 7976 75 8022 121
rect 7976 -19 8022 27
rect 7976 -113 8022 -67
rect 7976 -207 8022 -161
rect 7976 -301 8022 -255
rect 7976 -395 8022 -349
rect 7976 -489 8022 -443
rect 10234 75 10280 121
rect 10234 -19 10280 27
rect 10234 -113 10280 -67
rect 10234 -207 10280 -161
rect 10234 -301 10280 -255
rect 10234 -395 10280 -349
rect 10234 -489 10280 -443
rect 7976 -583 8022 -537
rect 10234 -583 10280 -537
rect 7976 -677 8022 -631
rect 7976 -771 8022 -725
rect 7976 -865 8022 -819
rect 7976 -959 8022 -913
rect 7976 -1053 8022 -1007
rect 7976 -1147 8022 -1101
rect 7976 -1241 8022 -1195
rect 10234 -677 10280 -631
rect 10234 -771 10280 -725
rect 10234 -865 10280 -819
rect 10234 -959 10280 -913
rect 10234 -1053 10280 -1007
rect 10234 -1147 10280 -1101
rect 10234 -1241 10280 -1195
rect 7976 -1335 8022 -1289
rect 10234 -1335 10280 -1289
rect 7976 -1429 8022 -1383
rect 7976 -1523 8022 -1477
rect 7976 -1617 8022 -1571
rect 7976 -1711 8022 -1665
rect 7976 -1805 8022 -1759
rect 7976 -1899 8022 -1853
rect 7976 -1993 8022 -1947
rect 10234 -1429 10280 -1383
rect 10234 -1523 10280 -1477
rect 10234 -1617 10280 -1571
rect 10234 -1711 10280 -1665
rect 10234 -1805 10280 -1759
rect 10234 -1899 10280 -1853
rect 7976 -2087 8022 -2041
rect 10234 -1993 10280 -1947
rect 7976 -2181 8022 -2135
rect 7976 -2275 8022 -2229
rect 7976 -2369 8022 -2323
rect 7976 -2463 8022 -2417
rect 7976 -2557 8022 -2511
rect 7976 -2651 8022 -2605
rect 7976 -2745 8022 -2699
rect 7976 -2839 8022 -2793
rect 10234 -2087 10280 -2041
rect 10234 -2181 10280 -2135
rect 10234 -2275 10280 -2229
rect 10234 -2369 10280 -2323
rect 10234 -2463 10280 -2417
rect 10234 -2557 10280 -2511
rect 10234 -2651 10280 -2605
rect 10234 -2745 10280 -2699
rect 10234 -2839 10280 -2793
rect 7977 -2933 8023 -2887
rect 8071 -2933 8117 -2887
rect 8165 -2933 8211 -2887
rect 8259 -2933 8305 -2887
rect 8353 -2933 8399 -2887
rect 8447 -2933 8493 -2887
rect 8541 -2933 8587 -2887
rect 8635 -2933 8681 -2887
rect 8729 -2933 8775 -2887
rect 8823 -2933 8869 -2887
rect 8917 -2933 8963 -2887
rect 9011 -2933 9057 -2887
rect 9105 -2933 9151 -2887
rect 9199 -2933 9245 -2887
rect 9293 -2933 9339 -2887
rect 9387 -2933 9433 -2887
rect 9481 -2933 9527 -2887
rect 9575 -2933 9621 -2887
rect 9669 -2933 9715 -2887
rect 9763 -2933 9809 -2887
rect 9857 -2933 9903 -2887
rect 9951 -2933 9997 -2887
rect 10045 -2933 10091 -2887
rect 10139 -2933 10185 -2887
rect 10233 -2933 10279 -2887
rect -747 -3159 -701 -3113
rect 1172 -3065 1218 -3019
rect 1172 -3159 1218 -3113
rect -747 -3253 -701 -3207
rect 1172 -3253 1218 -3207
rect -747 -3349 -701 -3303
rect -653 -3349 -607 -3303
rect -552 -3349 -506 -3303
rect -458 -3349 -412 -3303
rect -362 -3349 -316 -3303
rect -268 -3349 -222 -3303
rect -167 -3349 -121 -3303
rect -73 -3349 -27 -3303
rect 21 -3349 67 -3303
rect 115 -3349 161 -3303
rect 216 -3349 262 -3303
rect 310 -3349 356 -3303
rect 406 -3349 452 -3303
rect 500 -3349 546 -3303
rect 601 -3349 647 -3303
rect 695 -3349 741 -3303
rect 789 -3349 835 -3303
rect 883 -3349 929 -3303
rect 984 -3349 1030 -3303
rect 1078 -3349 1124 -3303
rect 1172 -3349 1218 -3303
rect -1291 -3486 -1245 -3440
rect -3267 -3580 -3221 -3534
rect -3267 -3674 -3221 -3628
rect -1291 -3580 -1245 -3534
rect -1291 -3674 -1245 -3628
rect -3267 -3768 -3221 -3722
rect -3267 -3862 -3221 -3816
rect -3267 -3956 -3221 -3910
rect -1291 -3768 -1245 -3722
rect -1291 -3862 -1245 -3816
rect -1291 -3956 -1245 -3910
rect -3267 -4050 -3221 -4004
rect -3267 -4144 -3221 -4098
rect -3267 -4238 -3221 -4192
rect -3267 -4332 -3221 -4286
rect -1291 -4050 -1245 -4004
rect -1291 -4144 -1245 -4098
rect -1291 -4238 -1245 -4192
rect -1291 -4332 -1245 -4286
rect -3267 -4426 -3221 -4380
rect -3267 -4520 -3221 -4474
rect -1291 -4426 -1245 -4380
rect -3267 -4614 -3221 -4568
rect -1291 -4520 -1245 -4474
rect -3267 -4708 -3221 -4662
rect -3267 -4802 -3221 -4756
rect -3267 -4896 -3221 -4850
rect -3267 -4990 -3221 -4944
rect -3267 -5084 -3221 -5038
rect -3267 -5178 -3221 -5132
rect -1291 -4614 -1245 -4568
rect -1291 -4708 -1245 -4662
rect -1291 -4802 -1245 -4756
rect -1291 -4896 -1245 -4850
rect -1291 -4990 -1245 -4944
rect -1291 -5084 -1245 -5038
rect -3267 -5272 -3221 -5226
rect -1291 -5178 -1245 -5132
rect -3267 -5366 -3221 -5320
rect -1291 -5272 -1245 -5226
rect -3267 -5460 -3221 -5414
rect -1291 -5366 -1245 -5320
rect -3267 -5554 -3221 -5508
rect -3267 -5648 -3221 -5602
rect -3267 -5742 -3221 -5696
rect -3267 -5836 -3221 -5790
rect -3267 -5930 -3221 -5884
rect -3267 -6024 -3221 -5978
rect -1291 -5460 -1245 -5414
rect -1291 -5554 -1245 -5508
rect -1291 -5648 -1245 -5602
rect -1291 -5742 -1245 -5696
rect -1291 -5836 -1245 -5790
rect -1291 -5930 -1245 -5884
rect -3267 -6118 -3221 -6072
rect -1291 -6024 -1245 -5978
rect -1291 -6118 -1245 -6072
rect -3267 -6212 -3221 -6166
rect -1291 -6212 -1245 -6166
rect -3266 -6306 -3220 -6260
rect -3172 -6306 -3126 -6260
rect -3078 -6306 -3032 -6260
rect -2984 -6306 -2938 -6260
rect -2890 -6306 -2844 -6260
rect -2796 -6306 -2750 -6260
rect -2702 -6306 -2656 -6260
rect -2608 -6306 -2562 -6260
rect -2514 -6306 -2468 -6260
rect -2420 -6306 -2374 -6260
rect -2326 -6306 -2280 -6260
rect -2232 -6306 -2186 -6260
rect -2138 -6306 -2092 -6260
rect -2044 -6306 -1998 -6260
rect -1950 -6306 -1904 -6260
rect -1856 -6306 -1810 -6260
rect -1762 -6306 -1716 -6260
rect -1668 -6306 -1622 -6260
rect -1574 -6306 -1528 -6260
rect -1480 -6306 -1434 -6260
rect -1386 -6306 -1340 -6260
rect -1292 -6306 -1246 -6260
rect -462 -4115 -415 -4068
rect -367 -4114 -321 -4068
rect -273 -4114 -227 -4068
rect -179 -4114 -133 -4068
rect -85 -4114 -39 -4068
rect 9 -4114 55 -4068
rect 103 -4114 149 -4068
rect 197 -4114 243 -4068
rect 291 -4114 337 -4068
rect 385 -4114 431 -4068
rect 479 -4114 525 -4068
rect 573 -4114 619 -4068
rect 667 -4114 713 -4068
rect 761 -4114 807 -4068
rect 855 -4114 901 -4068
rect 949 -4114 995 -4068
rect 1043 -4114 1089 -4068
rect 1137 -4114 1183 -4068
rect 1231 -4115 1278 -4068
rect -462 -4213 -416 -4163
rect 1232 -4213 1278 -4163
rect -462 -4307 -416 -4261
rect -462 -4401 -416 -4355
rect 1232 -4307 1278 -4261
rect 1232 -4401 1278 -4355
rect -462 -4495 -416 -4449
rect -462 -4589 -416 -4543
rect -462 -4683 -416 -4637
rect -462 -4777 -416 -4731
rect -462 -4871 -416 -4825
rect -462 -4965 -416 -4919
rect -462 -5059 -416 -5013
rect -462 -5153 -416 -5107
rect 1232 -4495 1278 -4449
rect 1232 -4589 1278 -4543
rect 1232 -4683 1278 -4637
rect 1232 -4777 1278 -4731
rect 1232 -4871 1278 -4825
rect 1232 -4965 1278 -4919
rect 1232 -5059 1278 -5013
rect -462 -5247 -416 -5201
rect 1232 -5153 1278 -5107
rect -462 -5341 -416 -5295
rect -462 -5435 -416 -5389
rect -462 -5529 -416 -5483
rect -462 -5623 -416 -5577
rect -462 -5717 -416 -5671
rect -462 -5811 -416 -5765
rect -462 -5905 -416 -5859
rect -462 -5999 -416 -5953
rect -462 -6093 -416 -6047
rect -462 -6187 -416 -6141
rect 1232 -5247 1278 -5201
rect 1232 -5341 1278 -5295
rect 1232 -5435 1278 -5389
rect 1232 -5529 1278 -5483
rect 1232 -5623 1278 -5577
rect 1232 -5717 1278 -5671
rect 1232 -5811 1278 -5765
rect 1232 -5905 1278 -5859
rect 1232 -5999 1278 -5953
rect 1232 -6093 1278 -6047
rect 1232 -6187 1278 -6141
rect -462 -6282 -415 -6235
rect -367 -6282 -321 -6236
rect -273 -6282 -227 -6236
rect -179 -6282 -133 -6236
rect -85 -6282 -39 -6236
rect 9 -6282 55 -6236
rect 103 -6282 149 -6236
rect 197 -6282 243 -6236
rect 291 -6282 337 -6236
rect 385 -6282 431 -6236
rect 479 -6282 525 -6236
rect 573 -6282 619 -6236
rect 667 -6282 713 -6236
rect 761 -6282 807 -6236
rect 855 -6282 901 -6236
rect 949 -6282 995 -6236
rect 1043 -6282 1089 -6236
rect 1137 -6282 1183 -6236
rect 1231 -6282 1278 -6235
rect 1622 -4365 1668 -4319
rect 1716 -4365 1762 -4319
rect 1810 -4365 1856 -4319
rect 1904 -4365 1950 -4319
rect 1998 -4365 2044 -4319
rect 2092 -4365 2138 -4319
rect 2186 -4365 2232 -4319
rect 2280 -4365 2326 -4319
rect 2374 -4365 2420 -4319
rect 2468 -4365 2514 -4319
rect 2562 -4365 2608 -4319
rect 2656 -4365 2702 -4319
rect 2750 -4365 2796 -4319
rect 2844 -4365 2890 -4319
rect 2938 -4365 2984 -4319
rect 3032 -4365 3078 -4319
rect 3126 -4365 3172 -4319
rect 3220 -4365 3266 -4319
rect 3314 -4365 3360 -4319
rect 3408 -4365 3454 -4319
rect 3502 -4365 3548 -4319
rect 3596 -4365 3642 -4319
rect 3690 -4365 3736 -4319
rect 1621 -4459 1667 -4413
rect 1621 -4553 1667 -4507
rect 3691 -4459 3737 -4413
rect 3691 -4553 3737 -4507
rect 1621 -4647 1667 -4601
rect 3691 -4647 3737 -4601
rect 1621 -4741 1667 -4695
rect 1621 -4835 1667 -4789
rect 1621 -4929 1667 -4883
rect 1621 -5023 1667 -4977
rect 1621 -5117 1667 -5071
rect 3691 -4741 3737 -4695
rect 3691 -4835 3737 -4789
rect 3691 -4929 3737 -4883
rect 3691 -5023 3737 -4977
rect 3691 -5117 3737 -5071
rect 1621 -5211 1667 -5165
rect 1621 -5305 1667 -5259
rect 3691 -5211 3737 -5165
rect 3691 -5305 3737 -5259
rect 1621 -5399 1667 -5353
rect 3691 -5399 3737 -5353
rect 1621 -5493 1667 -5447
rect 1621 -5587 1667 -5541
rect 1621 -5681 1667 -5635
rect 1621 -5775 1667 -5729
rect 1621 -5869 1667 -5823
rect 3691 -5493 3737 -5447
rect 3691 -5587 3737 -5541
rect 3691 -5681 3737 -5635
rect 3691 -5775 3737 -5729
rect 3691 -5869 3737 -5823
rect 1621 -5963 1667 -5917
rect 1621 -6057 1667 -6011
rect 3691 -5963 3737 -5917
rect 1621 -6151 1667 -6105
rect 3691 -6057 3737 -6011
rect 4029 -4468 4075 -4422
rect 4123 -4468 4169 -4422
rect 4217 -4468 4263 -4422
rect 4311 -4468 4357 -4422
rect 4405 -4468 4451 -4422
rect 4499 -4468 4545 -4422
rect 4593 -4468 4639 -4422
rect 4687 -4468 4733 -4422
rect 4781 -4468 4827 -4422
rect 4875 -4468 4921 -4422
rect 4969 -4468 5015 -4422
rect 5063 -4468 5109 -4422
rect 5157 -4468 5203 -4422
rect 5251 -4468 5297 -4422
rect 5345 -4468 5391 -4422
rect 5439 -4468 5485 -4422
rect 5533 -4468 5579 -4422
rect 5627 -4468 5673 -4422
rect 5721 -4468 5767 -4422
rect 5815 -4468 5861 -4422
rect 5909 -4468 5955 -4422
rect 6003 -4468 6049 -4422
rect 6097 -4468 6143 -4422
rect 6191 -4468 6237 -4422
rect 6285 -4468 6331 -4422
rect 6379 -4468 6425 -4422
rect 6473 -4468 6519 -4422
rect 6567 -4468 6613 -4422
rect 6661 -4468 6707 -4422
rect 4028 -4562 4074 -4516
rect 6662 -4562 6708 -4516
rect 4028 -4656 4074 -4610
rect 4028 -4750 4074 -4704
rect 6662 -4656 6708 -4610
rect 4028 -4844 4074 -4798
rect 4028 -4938 4074 -4892
rect 4028 -5032 4074 -4986
rect 4028 -5126 4074 -5080
rect 4028 -5220 4074 -5174
rect 6662 -4750 6708 -4704
rect 6662 -4844 6708 -4798
rect 6662 -4938 6708 -4892
rect 6662 -5032 6708 -4986
rect 6662 -5126 6708 -5080
rect 4028 -5314 4074 -5268
rect 6662 -5220 6708 -5174
rect 4028 -5408 4074 -5362
rect 4028 -5502 4074 -5456
rect 4028 -5596 4074 -5550
rect 4028 -5690 4074 -5644
rect 4028 -5784 4074 -5738
rect 6662 -5314 6708 -5268
rect 6662 -5408 6708 -5362
rect 6662 -5502 6708 -5456
rect 6662 -5596 6708 -5550
rect 6662 -5690 6708 -5644
rect 4028 -5878 4074 -5832
rect 6662 -5784 6708 -5738
rect 6662 -5878 6708 -5832
rect 4028 -5972 4074 -5926
rect 6662 -5972 6708 -5926
rect 4029 -6066 4075 -6020
rect 4123 -6066 4169 -6020
rect 4217 -6066 4263 -6020
rect 4311 -6066 4357 -6020
rect 4405 -6066 4451 -6020
rect 4499 -6066 4545 -6020
rect 4593 -6066 4639 -6020
rect 4687 -6066 4733 -6020
rect 4781 -6066 4827 -6020
rect 4875 -6066 4921 -6020
rect 4969 -6066 5015 -6020
rect 5063 -6066 5109 -6020
rect 5157 -6066 5203 -6020
rect 5251 -6066 5297 -6020
rect 5345 -6066 5391 -6020
rect 5439 -6066 5485 -6020
rect 5533 -6066 5579 -6020
rect 5627 -6066 5673 -6020
rect 5721 -6066 5767 -6020
rect 5815 -6066 5861 -6020
rect 5909 -6066 5955 -6020
rect 6003 -6066 6049 -6020
rect 6097 -6066 6143 -6020
rect 6191 -6066 6237 -6020
rect 6285 -6066 6331 -6020
rect 6379 -6066 6425 -6020
rect 6473 -6066 6519 -6020
rect 6567 -6066 6613 -6020
rect 6661 -6066 6707 -6020
rect 3691 -6151 3737 -6105
rect 1622 -6245 1668 -6199
rect 1716 -6245 1762 -6199
rect 1810 -6245 1856 -6199
rect 1904 -6245 1950 -6199
rect 1998 -6245 2044 -6199
rect 2092 -6245 2138 -6199
rect 2186 -6245 2232 -6199
rect 2280 -6245 2326 -6199
rect 2374 -6245 2420 -6199
rect 2468 -6245 2514 -6199
rect 2562 -6245 2608 -6199
rect 2656 -6245 2702 -6199
rect 2750 -6245 2796 -6199
rect 2844 -6245 2890 -6199
rect 2938 -6245 2984 -6199
rect 3032 -6245 3078 -6199
rect 3126 -6245 3172 -6199
rect 3220 -6245 3266 -6199
rect 3314 -6245 3360 -6199
rect 3408 -6245 3454 -6199
rect 3502 -6245 3548 -6199
rect 3596 -6245 3642 -6199
rect 3690 -6245 3736 -6199
<< polysilicon >>
rect -2679 1263 -1919 1276
rect -2679 1262 -2258 1263
rect -2679 1216 -2413 1262
rect -2367 1217 -2258 1262
rect -2212 1217 -1919 1263
rect -2367 1216 -1919 1217
rect -2679 1192 -1919 1216
rect -2679 507 -1919 517
rect -2895 504 -2783 505
rect -2895 458 -2864 504
rect -2818 458 -2783 504
rect -2895 457 -2783 458
rect -2679 461 -2428 507
rect -2382 504 -1919 507
rect -2382 461 -2215 504
rect -2679 457 -2215 461
rect -2167 457 -1919 504
rect -1815 504 -1703 505
rect -1815 458 -1782 504
rect -1736 458 -1703 504
rect -1815 457 -1703 458
rect -2679 444 -1919 457
rect -2895 -232 -2783 -231
rect -2895 -278 -2864 -232
rect -2818 -278 -2783 -232
rect -2895 -279 -2783 -278
rect -2679 -232 -1919 -219
rect -2679 -278 -2428 -232
rect -2382 -278 -2215 -232
rect -2679 -279 -2215 -278
rect -2167 -279 -1919 -232
rect -1815 -232 -1703 -231
rect -1815 -278 -1781 -232
rect -1735 -278 -1703 -232
rect -1815 -279 -1703 -278
rect -2679 -292 -1919 -279
rect -2895 -968 -2783 -967
rect -2895 -1014 -2863 -968
rect -2817 -1014 -2783 -968
rect -2895 -1015 -2783 -1014
rect -2679 -970 -1919 -955
rect -2679 -971 -2215 -970
rect -2679 -1017 -2428 -971
rect -2382 -1017 -2215 -971
rect -2167 -1017 -1919 -970
rect -1815 -968 -1703 -967
rect -1815 -1014 -1781 -968
rect -1735 -1014 -1703 -968
rect -1815 -1015 -1703 -1014
rect -2679 -1028 -1919 -1017
rect -365 842 -253 863
rect -365 796 -336 842
rect -290 796 -253 842
rect -365 758 -253 796
rect 715 844 827 864
rect 715 798 750 844
rect 796 798 827 844
rect 715 758 827 798
rect -149 -7 -37 70
rect 67 -7 179 70
rect 283 -7 395 70
rect 499 -7 611 70
rect -149 -60 611 -7
rect -149 -106 99 -60
rect 145 -62 611 -60
rect 145 -106 208 -62
rect -149 -108 208 -106
rect 254 -108 611 -62
rect -149 -153 611 -108
rect -149 -280 -37 -153
rect 67 -178 179 -153
rect 67 -224 99 -178
rect 145 -224 179 -178
rect 67 -280 179 -224
rect 283 -280 395 -153
rect 499 -280 611 -153
rect -365 -1122 -253 -968
rect -365 -1170 -330 -1122
rect -283 -1170 -253 -1122
rect -365 -1320 -253 -1170
rect -149 -1080 -37 -968
rect 67 -1028 179 -968
rect 67 -1074 99 -1028
rect 145 -1074 179 -1028
rect 67 -1080 179 -1074
rect 283 -1080 395 -968
rect 499 -1080 611 -968
rect -149 -1135 611 -1080
rect -149 -1181 99 -1135
rect 145 -1181 611 -1135
rect -149 -1226 611 -1181
rect -149 -1320 -37 -1226
rect 67 -1231 179 -1226
rect 67 -1277 99 -1231
rect 145 -1277 179 -1231
rect 67 -1320 179 -1277
rect 283 -1320 395 -1226
rect 499 -1320 611 -1226
rect 715 -1123 827 -968
rect 715 -1169 752 -1123
rect 798 -1169 827 -1123
rect 715 -1320 827 -1169
rect -149 -2117 -37 -2008
rect 67 -2057 179 -2008
rect 67 -2103 99 -2057
rect 145 -2103 179 -2057
rect 67 -2117 179 -2103
rect 283 -2117 395 -2008
rect 499 -2117 611 -2008
rect -149 -2171 611 -2117
rect -149 -2217 130 -2171
rect 176 -2217 611 -2171
rect -149 -2263 611 -2217
rect -149 -2358 -37 -2263
rect 67 -2358 179 -2263
rect 283 -2358 395 -2263
rect 499 -2358 611 -2263
rect -2849 -2747 -2762 -2733
rect -2849 -2793 -2828 -2747
rect -2782 -2793 -2762 -2747
rect -2849 -2813 -2762 -2793
rect -2370 -2747 -2283 -2731
rect -2370 -2793 -2348 -2747
rect -2302 -2793 -2283 -2747
rect -2370 -2811 -2283 -2793
rect -2207 -2747 -2120 -2731
rect -2207 -2793 -2188 -2747
rect -2142 -2793 -2120 -2747
rect -2207 -2811 -2120 -2793
rect -1728 -2747 -1642 -2733
rect -1728 -2793 -1708 -2747
rect -1662 -2793 -1642 -2747
rect -2833 -2865 -2777 -2813
rect -2353 -2821 -2297 -2811
rect -2193 -2821 -2137 -2811
rect -1728 -2813 -1642 -2793
rect -1713 -2865 -1657 -2813
rect 2591 952 2681 973
rect 2591 901 2610 952
rect 2661 901 2681 952
rect 2591 881 2681 901
rect 2767 942 4263 955
rect 2767 892 3488 942
rect 3538 892 4263 942
rect 2607 228 2663 881
rect 2767 877 4263 892
rect 4351 952 4441 973
rect 4351 901 4370 952
rect 4421 901 4441 952
rect 4351 881 4441 901
rect 4367 228 4423 881
rect 2591 207 2681 228
rect 2591 156 2610 207
rect 2661 156 2681 207
rect 2591 136 2681 156
rect 2767 207 4263 220
rect 2767 157 3489 207
rect 3539 157 4263 207
rect 2767 142 4263 157
rect 4351 207 4441 228
rect 4351 156 4370 207
rect 4421 156 4441 207
rect 4351 136 4441 156
rect 2607 -508 2663 136
rect 4367 -508 4423 136
rect 2591 -529 2681 -508
rect 2591 -580 2610 -529
rect 2661 -580 2681 -529
rect 2591 -600 2681 -580
rect 2767 -529 4263 -516
rect 2767 -579 3487 -529
rect 3537 -579 4263 -529
rect 2767 -594 4263 -579
rect 4351 -529 4441 -508
rect 4351 -580 4370 -529
rect 4421 -580 4441 -529
rect 4351 -600 4441 -580
rect 2607 -1245 2663 -600
rect 4367 -1245 4423 -600
rect 2591 -1266 2681 -1245
rect 2591 -1317 2610 -1266
rect 2661 -1317 2681 -1266
rect 2591 -1337 2681 -1317
rect 2767 -1265 4263 -1252
rect 2767 -1315 3487 -1265
rect 3537 -1315 4263 -1265
rect 2767 -1330 4263 -1315
rect 4351 -1266 4441 -1245
rect 4351 -1317 4370 -1266
rect 4421 -1317 4441 -1266
rect 4351 -1337 4441 -1317
rect 2607 -1981 2663 -1337
rect 4367 -1981 4423 -1337
rect 2591 -2002 2681 -1981
rect 2591 -2053 2610 -2002
rect 2661 -2053 2681 -2002
rect 2591 -2073 2681 -2053
rect 2767 -1999 4263 -1986
rect 2767 -2049 3488 -1999
rect 3538 -2049 4263 -1999
rect 2767 -2064 4263 -2049
rect 4351 -2002 4441 -1981
rect 4351 -2053 4370 -2002
rect 4421 -2053 4441 -2002
rect 4351 -2073 4441 -2053
rect 2607 -2739 2663 -2073
rect 2767 -2734 4263 -2721
rect 2767 -2784 3486 -2734
rect 3536 -2784 4263 -2734
rect 4367 -2739 4423 -2073
rect 2767 -2799 4263 -2784
rect 5391 952 5481 973
rect 5391 901 5410 952
rect 5461 901 5481 952
rect 5391 881 5481 901
rect 5567 942 7063 955
rect 5567 892 6288 942
rect 6338 892 7063 942
rect 5407 228 5463 881
rect 5567 877 7063 892
rect 7151 952 7241 973
rect 7151 901 7170 952
rect 7221 901 7241 952
rect 7151 881 7241 901
rect 7167 228 7223 881
rect 5391 207 5481 228
rect 5391 156 5410 207
rect 5461 156 5481 207
rect 5391 136 5481 156
rect 5567 207 7063 220
rect 5567 157 6289 207
rect 6339 157 7063 207
rect 5567 142 7063 157
rect 7151 207 7241 228
rect 7151 156 7170 207
rect 7221 156 7241 207
rect 7151 136 7241 156
rect 5407 -508 5463 136
rect 7167 -508 7223 136
rect 5391 -529 5481 -508
rect 5391 -580 5410 -529
rect 5461 -580 5481 -529
rect 5391 -600 5481 -580
rect 5567 -529 7063 -516
rect 5567 -579 6287 -529
rect 6337 -579 7063 -529
rect 5567 -594 7063 -579
rect 7151 -529 7241 -508
rect 7151 -580 7170 -529
rect 7221 -580 7241 -529
rect 7151 -600 7241 -580
rect 5407 -1245 5463 -600
rect 7167 -1245 7223 -600
rect 5391 -1266 5481 -1245
rect 5391 -1317 5410 -1266
rect 5461 -1317 5481 -1266
rect 5391 -1337 5481 -1317
rect 5567 -1265 7063 -1252
rect 5567 -1315 6287 -1265
rect 6337 -1315 7063 -1265
rect 5567 -1330 7063 -1315
rect 7151 -1266 7241 -1245
rect 7151 -1317 7170 -1266
rect 7221 -1317 7241 -1266
rect 7151 -1337 7241 -1317
rect 5407 -1981 5463 -1337
rect 7167 -1981 7223 -1337
rect 5391 -2002 5481 -1981
rect 5391 -2053 5410 -2002
rect 5461 -2053 5481 -2002
rect 5391 -2073 5481 -2053
rect 5567 -1999 7063 -1986
rect 5567 -2049 6288 -1999
rect 6338 -2049 7063 -1999
rect 5567 -2064 7063 -2049
rect 7151 -2002 7241 -1981
rect 7151 -2053 7170 -2002
rect 7221 -2053 7241 -2002
rect 7151 -2073 7241 -2053
rect 5407 -2739 5463 -2073
rect 5567 -2734 7063 -2721
rect 5567 -2784 6286 -2734
rect 6336 -2784 7063 -2734
rect 7167 -2739 7223 -2073
rect 5567 -2799 7063 -2784
rect 8191 952 8281 973
rect 8191 901 8210 952
rect 8261 901 8281 952
rect 8191 881 8281 901
rect 8367 942 9863 955
rect 8367 892 9088 942
rect 9138 892 9863 942
rect 8207 228 8263 881
rect 8367 877 9863 892
rect 9951 952 10041 973
rect 9951 901 9970 952
rect 10021 901 10041 952
rect 9951 881 10041 901
rect 9967 228 10023 881
rect 8191 207 8281 228
rect 8191 156 8210 207
rect 8261 156 8281 207
rect 8191 136 8281 156
rect 8367 207 9863 220
rect 8367 157 9089 207
rect 9139 157 9863 207
rect 8367 142 9863 157
rect 9951 207 10041 228
rect 9951 156 9970 207
rect 10021 156 10041 207
rect 9951 136 10041 156
rect 8207 -508 8263 136
rect 9967 -508 10023 136
rect 8191 -529 8281 -508
rect 8191 -580 8210 -529
rect 8261 -580 8281 -529
rect 8191 -600 8281 -580
rect 8367 -529 9863 -516
rect 8367 -579 9087 -529
rect 9137 -579 9863 -529
rect 8367 -594 9863 -579
rect 9951 -529 10041 -508
rect 9951 -580 9970 -529
rect 10021 -580 10041 -529
rect 9951 -600 10041 -580
rect 8207 -1245 8263 -600
rect 9967 -1245 10023 -600
rect 8191 -1266 8281 -1245
rect 8191 -1317 8210 -1266
rect 8261 -1317 8281 -1266
rect 8191 -1337 8281 -1317
rect 8367 -1265 9863 -1252
rect 8367 -1315 9087 -1265
rect 9137 -1315 9863 -1265
rect 8367 -1330 9863 -1315
rect 9951 -1266 10041 -1245
rect 9951 -1317 9970 -1266
rect 10021 -1317 10041 -1266
rect 9951 -1337 10041 -1317
rect 8207 -1981 8263 -1337
rect 9967 -1981 10023 -1337
rect 8191 -2002 8281 -1981
rect 8191 -2053 8210 -2002
rect 8261 -2053 8281 -2002
rect 8191 -2073 8281 -2053
rect 8367 -1999 9863 -1986
rect 8367 -2049 9088 -1999
rect 9138 -2049 9863 -1999
rect 8367 -2064 9863 -2049
rect 9951 -2002 10041 -1981
rect 9951 -2053 9970 -2002
rect 10021 -2053 10041 -2002
rect 9951 -2073 10041 -2053
rect 8207 -2739 8263 -2073
rect 8367 -2734 9863 -2721
rect 8367 -2784 9086 -2734
rect 9136 -2784 9863 -2734
rect 9967 -2739 10023 -2073
rect 8367 -2799 9863 -2784
rect -365 -3132 -253 -3045
rect -365 -3184 -333 -3132
rect -276 -3184 -253 -3132
rect -365 -3206 -253 -3184
rect 715 -3128 827 -3046
rect 715 -3182 738 -3128
rect 796 -3182 827 -3128
rect 715 -3202 827 -3182
rect -3077 -3534 -2937 -3509
rect -3077 -3580 -3061 -3534
rect -3015 -3580 -2937 -3534
rect -2673 -3542 -2617 -3497
rect -2513 -3542 -2457 -3497
rect -2033 -3542 -1977 -3497
rect -1873 -3542 -1817 -3497
rect -1553 -3525 -1403 -3509
rect -2684 -3559 -2606 -3542
rect -3077 -3595 -2937 -3580
rect -2845 -3580 -2767 -3563
rect -2845 -3626 -2829 -3580
rect -2783 -3626 -2767 -3580
rect -2684 -3605 -2668 -3559
rect -2622 -3605 -2606 -3559
rect -2684 -3619 -2606 -3605
rect -2524 -3558 -2446 -3542
rect -2524 -3604 -2508 -3558
rect -2462 -3604 -2446 -3558
rect -2044 -3558 -1966 -3542
rect -2524 -3619 -2446 -3604
rect -2363 -3577 -2285 -3563
rect -2845 -3640 -2767 -3626
rect -2363 -3623 -2348 -3577
rect -2302 -3623 -2285 -3577
rect -2363 -3640 -2285 -3623
rect -2205 -3577 -2127 -3563
rect -2205 -3623 -2188 -3577
rect -2142 -3623 -2127 -3577
rect -2044 -3604 -2028 -3558
rect -1982 -3604 -1966 -3558
rect -2044 -3619 -1966 -3604
rect -1884 -3559 -1806 -3542
rect -1884 -3605 -1868 -3559
rect -1822 -3605 -1806 -3559
rect -1884 -3619 -1806 -3605
rect -1723 -3580 -1645 -3563
rect -2205 -3640 -2127 -3623
rect -1723 -3626 -1707 -3580
rect -1661 -3626 -1645 -3580
rect -1553 -3571 -1468 -3525
rect -1422 -3571 -1403 -3525
rect -1553 -3596 -1403 -3571
rect -1723 -3640 -1645 -3626
rect -2833 -3685 -2777 -3640
rect -2353 -3685 -2297 -3640
rect -2193 -3685 -2137 -3640
rect -1713 -3685 -1657 -3640
rect -3086 -4380 -2937 -4361
rect -3086 -4426 -3068 -4380
rect -3022 -4426 -2937 -4380
rect -2673 -4402 -2617 -4361
rect -3086 -4453 -2937 -4426
rect -2688 -4420 -2601 -4402
rect -2513 -4403 -2457 -4361
rect -2033 -4403 -1977 -4361
rect -1873 -4402 -1817 -4361
rect -1553 -4381 -1396 -4361
rect -2688 -4466 -2667 -4420
rect -2621 -4466 -2601 -4420
rect -2688 -4484 -2601 -4466
rect -2529 -4420 -2442 -4403
rect -2529 -4466 -2507 -4420
rect -2461 -4466 -2442 -4420
rect -2529 -4483 -2442 -4466
rect -2048 -4420 -1961 -4403
rect -2048 -4466 -2029 -4420
rect -1983 -4466 -1961 -4420
rect -2048 -4483 -1961 -4466
rect -1889 -4420 -1802 -4402
rect -1889 -4466 -1869 -4420
rect -1823 -4466 -1802 -4420
rect -1553 -4427 -1468 -4381
rect -1422 -4427 -1396 -4381
rect -1553 -4448 -1396 -4427
rect -2993 -4569 -2937 -4525
rect -2833 -4569 -2777 -4525
rect -2673 -4569 -2617 -4484
rect -2513 -4569 -2457 -4483
rect -2353 -4569 -2297 -4525
rect -2193 -4569 -2137 -4525
rect -2033 -4569 -1977 -4483
rect -1889 -4484 -1802 -4466
rect -1873 -4569 -1817 -4484
rect -1713 -4569 -1657 -4525
rect -1553 -4569 -1497 -4525
rect -2993 -5213 -2937 -5169
rect -3083 -5231 -2937 -5213
rect -3083 -5277 -3068 -5231
rect -3022 -5277 -2937 -5231
rect -2833 -5246 -2777 -5169
rect -2673 -5213 -2617 -5169
rect -2513 -5213 -2457 -5169
rect -2353 -5246 -2297 -5169
rect -2193 -5246 -2137 -5169
rect -2033 -5213 -1977 -5169
rect -1873 -5213 -1817 -5169
rect -1713 -5246 -1657 -5169
rect -1553 -5213 -1497 -5169
rect -1553 -5232 -1403 -5213
rect -3083 -5296 -2937 -5277
rect -2845 -5260 -2767 -5246
rect -2845 -5306 -2829 -5260
rect -2783 -5306 -2767 -5260
rect -2363 -5263 -2285 -5246
rect -2845 -5323 -2767 -5306
rect -2684 -5281 -2606 -5267
rect -2684 -5327 -2668 -5281
rect -2622 -5327 -2606 -5281
rect -2684 -5344 -2606 -5327
rect -2524 -5282 -2446 -5267
rect -2524 -5328 -2508 -5282
rect -2462 -5328 -2446 -5282
rect -2363 -5309 -2348 -5263
rect -2302 -5309 -2285 -5263
rect -2363 -5323 -2285 -5309
rect -2205 -5263 -2127 -5246
rect -2205 -5309 -2188 -5263
rect -2142 -5309 -2127 -5263
rect -1723 -5260 -1645 -5246
rect -2205 -5323 -2127 -5309
rect -2044 -5282 -1966 -5267
rect -2524 -5344 -2446 -5328
rect -2044 -5328 -2028 -5282
rect -1982 -5328 -1966 -5282
rect -2044 -5344 -1966 -5328
rect -1884 -5281 -1806 -5267
rect -1884 -5327 -1868 -5281
rect -1822 -5327 -1806 -5281
rect -1723 -5306 -1707 -5260
rect -1661 -5306 -1645 -5260
rect -1553 -5278 -1468 -5232
rect -1422 -5278 -1403 -5232
rect -1553 -5305 -1403 -5278
rect -1723 -5323 -1645 -5306
rect -1884 -5344 -1806 -5327
rect -2993 -5421 -2937 -5377
rect -2833 -5421 -2777 -5377
rect -2673 -5421 -2617 -5344
rect -2513 -5421 -2457 -5344
rect -2353 -5421 -2297 -5377
rect -2193 -5421 -2137 -5377
rect -2033 -5421 -1977 -5344
rect -1873 -5421 -1817 -5344
rect -1713 -5421 -1657 -5377
rect -1553 -5421 -1497 -5377
rect -2993 -6065 -2937 -6021
rect -3086 -6081 -2937 -6065
rect -2833 -6073 -2777 -6021
rect -2673 -6065 -2617 -6021
rect -2513 -6065 -2457 -6021
rect -3086 -6127 -3068 -6081
rect -3022 -6127 -2937 -6081
rect -3086 -6147 -2937 -6127
rect -2849 -6093 -2762 -6073
rect -2353 -6075 -2297 -6021
rect -2193 -6075 -2137 -6021
rect -2033 -6065 -1977 -6021
rect -1873 -6065 -1817 -6021
rect -1713 -6073 -1657 -6021
rect -1553 -6065 -1497 -6021
rect -2849 -6139 -2828 -6093
rect -2782 -6139 -2762 -6093
rect -2849 -6153 -2762 -6139
rect -2370 -6093 -2283 -6075
rect -2370 -6139 -2348 -6093
rect -2302 -6139 -2283 -6093
rect -2370 -6155 -2283 -6139
rect -2207 -6093 -2120 -6075
rect -2207 -6139 -2188 -6093
rect -2142 -6139 -2120 -6093
rect -2207 -6155 -2120 -6139
rect -1728 -6093 -1641 -6073
rect -1728 -6139 -1708 -6093
rect -1662 -6139 -1641 -6093
rect -1728 -6153 -1641 -6139
rect -1553 -6085 -1403 -6065
rect -1553 -6131 -1468 -6085
rect -1422 -6131 -1403 -6085
rect -1553 -6152 -1403 -6131
rect -315 -4246 80 -4226
rect -315 -4304 -295 -4246
rect -230 -4248 80 -4246
rect -230 -4303 -154 -4248
rect -90 -4303 80 -4248
rect -230 -4304 80 -4303
rect -315 -4318 80 -4304
rect -1 -4361 80 -4318
rect -1 -4444 791 -4361
rect -173 -5148 -90 -5132
rect -173 -5194 -156 -5148
rect -110 -5194 -90 -5148
rect -173 -5211 -90 -5194
rect -161 -5224 -105 -5211
rect -1 -5224 791 -5132
rect 895 -5135 951 -5132
rect 884 -5152 967 -5135
rect 884 -5198 901 -5152
rect 947 -5198 967 -5152
rect 884 -5214 967 -5198
rect 895 -5224 951 -5214
rect 2076 -4595 3268 -4562
rect 2076 -4655 2583 -4595
rect 2643 -4655 2713 -4595
rect 2773 -4655 3268 -4595
rect 2076 -4690 3268 -4655
rect 1860 -5180 1972 -5136
rect 1825 -5213 1972 -5180
rect 1825 -5271 1865 -5213
rect 1923 -5271 1972 -5213
rect 1825 -5306 1972 -5271
rect 2076 -5228 2188 -5178
rect 2292 -5228 2404 -5178
rect 2508 -5228 2620 -5178
rect 2724 -5228 2836 -5178
rect 2940 -5228 3052 -5178
rect 3156 -5228 3268 -5173
rect 2076 -5321 3268 -5228
rect 3372 -5180 3484 -5136
rect 3372 -5213 3519 -5180
rect 3372 -5271 3421 -5213
rect 3479 -5271 3519 -5213
rect 3372 -5306 3519 -5271
rect 2076 -5350 2441 -5321
rect 2162 -5398 2274 -5350
rect 2419 -5381 2441 -5350
rect 2501 -5350 3268 -5321
rect 2501 -5381 2620 -5350
rect 2419 -5398 2620 -5381
rect 2724 -5398 2836 -5350
rect 2419 -5404 2550 -5398
rect 1946 -5886 2058 -5842
rect 3070 -5886 3182 -5842
rect 1911 -5919 2058 -5886
rect 1911 -5977 1951 -5919
rect 2009 -5977 2058 -5919
rect 1911 -6012 2058 -5977
rect 3035 -5919 3182 -5886
rect 3035 -5977 3075 -5919
rect 3133 -5977 3182 -5919
rect 3035 -6012 3182 -5977
rect 3286 -5919 3433 -5886
rect 3286 -5977 3335 -5919
rect 3393 -5977 3433 -5919
rect 3286 -6012 3433 -5977
rect 4587 -4629 6141 -4570
rect 4587 -4695 5256 -4629
rect 5322 -4695 5394 -4629
rect 5460 -4695 6141 -4629
rect 4587 -4723 6141 -4695
rect 4283 -5212 4483 -5199
rect 4283 -5262 4302 -5212
rect 4352 -5262 4415 -5212
rect 4465 -5262 4483 -5212
rect 4283 -5274 4483 -5262
rect 4587 -5209 6141 -5198
rect 4587 -5261 5302 -5209
rect 5354 -5261 6141 -5209
rect 4587 -5270 6141 -5261
rect 6245 -5214 6445 -5201
rect 6245 -5264 6264 -5214
rect 6314 -5264 6377 -5214
rect 6427 -5264 6445 -5214
rect 6245 -5276 6445 -5264
rect 4587 -5788 6141 -5747
rect 4587 -5854 5256 -5788
rect 5322 -5854 5394 -5788
rect 5460 -5854 6141 -5788
rect 4587 -5900 6141 -5854
rect 9187 -4966 10683 -4937
rect 9187 -4967 10224 -4966
rect 9187 -4970 9893 -4967
rect 9187 -4971 9576 -4970
rect 9187 -5030 9262 -4971
rect 9321 -5029 9576 -4971
rect 9635 -5026 9893 -4970
rect 9952 -5025 10224 -4967
rect 10283 -4967 10683 -4966
rect 10283 -5025 10543 -4967
rect 9952 -5026 10543 -5025
rect 10602 -5026 10683 -4967
rect 9635 -5029 10683 -5026
rect 9321 -5030 10683 -5029
rect 9187 -5076 10683 -5030
rect 9015 -5754 9095 -5740
rect 9015 -5805 9029 -5754
rect 9080 -5805 9095 -5754
rect 9015 -5819 9095 -5805
rect 9187 -5814 10683 -5743
rect 10774 -5755 10854 -5741
rect 10774 -5806 10788 -5755
rect 10839 -5806 10854 -5755
rect 10774 -5820 10854 -5806
rect -3063 -7053 -2918 -7040
rect -3063 -7099 -3049 -7053
rect -3003 -7099 -2918 -7053
rect -1534 -7053 -1389 -7040
rect -3063 -7112 -2918 -7099
rect -2974 -7139 -2918 -7112
rect -2174 -7139 -2118 -7095
rect -2014 -7139 -1958 -7095
rect -1854 -7139 -1798 -7095
rect -1694 -7139 -1638 -7095
rect -1534 -7099 -1449 -7053
rect -1403 -7099 -1389 -7053
rect -1534 -7112 -1389 -7099
rect -1534 -7139 -1478 -7112
rect -2814 -7789 -2758 -7783
rect -2654 -7789 -2598 -7783
rect -2494 -7789 -2438 -7783
rect -2334 -7789 -2278 -7783
rect -2174 -7789 -2118 -7739
rect -2014 -7789 -1958 -7739
rect -1854 -7789 -1798 -7739
rect -1694 -7789 -1638 -7739
rect -1534 -7783 -1478 -7739
rect -2814 -7815 -1638 -7789
rect -3063 -7853 -2918 -7840
rect -3063 -7899 -3049 -7853
rect -3003 -7899 -2918 -7853
rect -2814 -7864 -2251 -7815
rect -2202 -7864 -1638 -7815
rect -2814 -7887 -1638 -7864
rect -2814 -7895 -2758 -7887
rect -2654 -7895 -2598 -7887
rect -2494 -7895 -2438 -7887
rect -2334 -7895 -2278 -7887
rect -3063 -7912 -2918 -7899
rect -2974 -7939 -2918 -7912
rect -2174 -7939 -2118 -7887
rect -2014 -7939 -1958 -7887
rect -1854 -7939 -1798 -7887
rect -1694 -7939 -1638 -7887
rect -1534 -7853 -1389 -7840
rect -1534 -7899 -1449 -7853
rect -1403 -7899 -1389 -7853
rect -1534 -7912 -1389 -7899
rect -1534 -7939 -1478 -7912
rect -2814 -8589 -2758 -8583
rect -2654 -8589 -2598 -8583
rect -2494 -8589 -2438 -8583
rect -2334 -8589 -2278 -8583
rect -2174 -8589 -2118 -8539
rect -2014 -8589 -1958 -8539
rect -1854 -8589 -1798 -8539
rect -1694 -8589 -1638 -8539
rect -1534 -8583 -1478 -8539
rect -2814 -8616 -1638 -8589
rect -3063 -8651 -2918 -8638
rect -3063 -8697 -3049 -8651
rect -3003 -8697 -2918 -8651
rect -3063 -8710 -2918 -8697
rect -2974 -8737 -2918 -8710
rect -2814 -8665 -2251 -8616
rect -2202 -8665 -1638 -8616
rect -2814 -8687 -1638 -8665
rect -2814 -8737 -2758 -8687
rect -2654 -8737 -2598 -8687
rect -2494 -8737 -2438 -8687
rect -2334 -8737 -2278 -8687
rect -2174 -8737 -2118 -8687
rect -2014 -8737 -1958 -8687
rect -1854 -8737 -1798 -8687
rect -1694 -8737 -1638 -8687
rect -1534 -8651 -1389 -8638
rect -1534 -8697 -1449 -8651
rect -1403 -8697 -1389 -8651
rect -1534 -8710 -1389 -8697
rect -1534 -8737 -1478 -8710
rect -2974 -9381 -2918 -9337
rect -2814 -9389 -2758 -9337
rect -2654 -9389 -2598 -9337
rect -2494 -9389 -2438 -9337
rect -2334 -9389 -2278 -9337
rect -2174 -9389 -2118 -9337
rect -2014 -9389 -1958 -9337
rect -1854 -9389 -1798 -9337
rect -1694 -9389 -1638 -9337
rect -1534 -9381 -1478 -9337
rect -2814 -9416 -1638 -9389
rect -3063 -9451 -2918 -9438
rect -3063 -9497 -3049 -9451
rect -3003 -9497 -2918 -9451
rect -3063 -9510 -2918 -9497
rect -2974 -9537 -2918 -9510
rect -2814 -9465 -2252 -9416
rect -2203 -9465 -1638 -9416
rect -2814 -9487 -1638 -9465
rect -2814 -9537 -2758 -9487
rect -2654 -9537 -2598 -9487
rect -2494 -9537 -2438 -9487
rect -2334 -9537 -2278 -9487
rect -2174 -9537 -2118 -9487
rect -2014 -9537 -1958 -9487
rect -1854 -9537 -1798 -9487
rect -1694 -9537 -1638 -9487
rect -1534 -9451 -1389 -9438
rect -1534 -9497 -1449 -9451
rect -1403 -9497 -1389 -9451
rect -1534 -9510 -1389 -9497
rect -1534 -9537 -1478 -9510
rect -2974 -10181 -2918 -10137
rect -2814 -10181 -2758 -10137
rect -2654 -10181 -2598 -10137
rect -2494 -10181 -2438 -10137
rect -2334 -10181 -2278 -10137
rect -2174 -10181 -2118 -10137
rect -2014 -10181 -1958 -10137
rect -1854 -10181 -1798 -10137
rect -1694 -10181 -1638 -10137
rect -1534 -10181 -1478 -10137
rect -262 -6863 -183 -6842
rect -262 -6909 -245 -6863
rect -199 -6909 -183 -6863
rect -262 -6938 -183 -6909
rect 863 -6885 940 -6871
rect 863 -6931 878 -6885
rect 924 -6931 940 -6885
rect 863 -6946 940 -6931
rect -89 -7645 -33 -7626
rect 232 -7645 288 -7626
rect 392 -7645 448 -7626
rect 713 -7645 769 -7626
rect -89 -7682 769 -7645
rect -260 -7725 -180 -7705
rect -260 -7771 -243 -7725
rect -197 -7771 -180 -7725
rect -260 -7788 -180 -7771
rect -89 -7740 313 -7682
rect 371 -7740 769 -7682
rect -89 -7769 769 -7740
rect -89 -7788 -33 -7769
rect 232 -7788 288 -7769
rect 392 -7788 448 -7769
rect 713 -7788 769 -7769
rect 862 -7743 939 -7729
rect 862 -7789 877 -7743
rect 923 -7789 939 -7743
rect 862 -7803 939 -7789
rect 2046 -6774 2374 -6737
rect 2046 -6835 2113 -6774
rect 2174 -6775 2374 -6774
rect 2174 -6835 2259 -6775
rect 2046 -6836 2259 -6835
rect 2320 -6836 2374 -6775
rect 2046 -6877 2374 -6836
rect 2478 -6772 3498 -6737
rect 2478 -6830 2873 -6772
rect 2931 -6773 3498 -6772
rect 2931 -6830 3010 -6773
rect 2478 -6831 3010 -6830
rect 3068 -6831 3498 -6773
rect 2478 -6877 3498 -6831
rect 9015 -6491 9095 -6477
rect 9015 -6542 9029 -6491
rect 9080 -6542 9095 -6491
rect 9015 -6556 9095 -6542
rect 9187 -6549 10683 -6478
rect 10774 -6491 10854 -6477
rect 10774 -6542 10788 -6491
rect 10839 -6542 10854 -6491
rect 10774 -6556 10854 -6542
rect 2824 -6907 2936 -6877
rect 1830 -7378 1942 -7334
rect 1795 -7411 1942 -7378
rect 1795 -7469 1835 -7411
rect 1893 -7469 1942 -7411
rect 1795 -7504 1942 -7469
rect 3735 -7368 3847 -7324
rect 3735 -7401 3882 -7368
rect 3735 -7459 3784 -7401
rect 3842 -7459 3882 -7401
rect 3735 -7494 3882 -7459
rect 5069 -6952 7397 -6896
rect 5069 -7018 6135 -6952
rect 6201 -7018 6273 -6952
rect 6339 -7018 7397 -6952
rect 5069 -7066 7397 -7018
rect 4627 -7553 4827 -7536
rect 4627 -7603 4646 -7553
rect 4696 -7603 4759 -7553
rect 4809 -7603 4827 -7553
rect 4627 -7616 4827 -7603
rect 5069 -7553 7397 -7538
rect 5069 -7603 6152 -7553
rect 6202 -7603 6265 -7553
rect 6315 -7603 7397 -7553
rect 5069 -7618 7397 -7603
rect 7635 -7553 7835 -7538
rect 7635 -7603 7654 -7553
rect 7704 -7603 7767 -7553
rect 7817 -7603 7835 -7553
rect 7635 -7616 7835 -7603
rect 9187 -7256 10683 -7218
rect 9187 -7259 10540 -7256
rect 9187 -7262 9589 -7259
rect 9187 -7321 9261 -7262
rect 9320 -7318 9589 -7262
rect 9648 -7260 10540 -7259
rect 9648 -7318 9899 -7260
rect 9320 -7319 9899 -7318
rect 9958 -7319 10225 -7260
rect 10284 -7315 10540 -7260
rect 10599 -7315 10683 -7256
rect 10284 -7319 10683 -7315
rect 9320 -7321 10683 -7319
rect 9187 -7354 10683 -7321
rect 9187 -7357 10645 -7354
rect 4627 -8092 4827 -8079
rect 4627 -8142 4646 -8092
rect 4696 -8142 4759 -8092
rect 4809 -8142 4827 -8092
rect 4627 -8155 4827 -8142
rect 5069 -8089 7397 -8074
rect 5069 -8139 6150 -8089
rect 6200 -8139 6263 -8089
rect 6313 -8139 7397 -8089
rect 5069 -8154 7397 -8139
rect 7635 -8087 7835 -8072
rect 7635 -8137 7654 -8087
rect 7704 -8137 7767 -8087
rect 7817 -8137 7835 -8087
rect 7635 -8150 7835 -8137
rect -89 -8562 -33 -8476
rect 232 -8562 288 -8476
rect 392 -8562 448 -8476
rect 713 -8562 769 -8476
rect -89 -8593 984 -8562
rect -89 -8651 908 -8593
rect 966 -8651 984 -8593
rect -89 -8686 984 -8651
rect -89 -8768 -33 -8686
rect 232 -8768 288 -8686
rect 392 -8768 448 -8686
rect 713 -8768 769 -8686
rect -264 -9468 -175 -9453
rect -264 -9514 -243 -9468
rect -197 -9514 -175 -9468
rect -264 -9531 -175 -9514
rect -89 -9475 -33 -9456
rect 232 -9475 288 -9456
rect 392 -9475 448 -9456
rect 713 -9475 769 -9456
rect -89 -9511 769 -9475
rect -89 -9569 304 -9511
rect 362 -9569 769 -9511
rect 858 -9474 948 -9456
rect 858 -9520 880 -9474
rect 926 -9520 948 -9474
rect 858 -9534 948 -9520
rect -89 -9599 769 -9569
rect -89 -9618 -33 -9599
rect 232 -9618 288 -9599
rect 392 -9618 448 -9599
rect 713 -9618 769 -9599
rect -261 -10321 -185 -10306
rect -261 -10367 -246 -10321
rect -200 -10367 -185 -10321
rect -261 -10381 -185 -10367
rect 873 -10329 1019 -10306
rect 873 -10375 957 -10329
rect 1003 -10375 1019 -10329
rect 873 -10396 1019 -10375
rect 5069 -8683 7397 -8626
rect 5069 -8749 6132 -8683
rect 6198 -8749 6270 -8683
rect 6336 -8749 7397 -8683
rect 5069 -8796 7397 -8749
rect 9187 -7966 10683 -7937
rect 9187 -7967 10224 -7966
rect 9187 -7970 9893 -7967
rect 9187 -7971 9576 -7970
rect 9187 -8030 9262 -7971
rect 9321 -8029 9576 -7971
rect 9635 -8026 9893 -7970
rect 9952 -8025 10224 -7967
rect 10283 -7967 10683 -7966
rect 10283 -8025 10543 -7967
rect 9952 -8026 10543 -8025
rect 10602 -8026 10683 -7967
rect 9635 -8029 10683 -8026
rect 9321 -8030 10683 -8029
rect 9187 -8076 10683 -8030
rect 9015 -8754 9095 -8740
rect 9015 -8805 9029 -8754
rect 9080 -8805 9095 -8754
rect 9015 -8819 9095 -8805
rect 9187 -8814 10683 -8743
rect 10774 -8755 10854 -8741
rect 10774 -8806 10788 -8755
rect 10839 -8806 10854 -8755
rect 10774 -8820 10854 -8806
rect 1875 -9150 2731 -9133
rect 1875 -9151 2544 -9150
rect 1875 -9203 1905 -9151
rect 1957 -9152 2544 -9151
rect 1957 -9203 2011 -9152
rect 1875 -9204 2011 -9203
rect 2063 -9204 2223 -9152
rect 2275 -9153 2544 -9152
rect 2275 -9204 2329 -9153
rect 1875 -9205 2329 -9204
rect 2381 -9202 2544 -9153
rect 2596 -9151 2731 -9150
rect 2596 -9202 2650 -9151
rect 2381 -9203 2650 -9202
rect 2702 -9203 2731 -9151
rect 2381 -9205 2731 -9203
rect 1875 -9219 2731 -9205
rect 1868 -9499 2724 -9485
rect 1868 -9500 2322 -9499
rect 1868 -9501 2004 -9500
rect 1868 -9553 1898 -9501
rect 1950 -9552 2004 -9501
rect 2056 -9552 2216 -9500
rect 2268 -9551 2322 -9500
rect 2374 -9501 2724 -9499
rect 2374 -9502 2643 -9501
rect 2374 -9551 2537 -9502
rect 2268 -9552 2537 -9551
rect 1950 -9553 2537 -9552
rect 1868 -9554 2537 -9553
rect 2589 -9553 2643 -9502
rect 2695 -9553 2724 -9501
rect 2589 -9554 2724 -9553
rect 1868 -9571 2724 -9554
rect 9015 -9491 9095 -9477
rect 9015 -9542 9029 -9491
rect 9080 -9542 9095 -9491
rect 9015 -9556 9095 -9542
rect 9187 -9549 10683 -9478
rect 10774 -9491 10854 -9477
rect 10774 -9542 10788 -9491
rect 10839 -9542 10854 -9491
rect 10774 -9556 10854 -9542
rect 9187 -10256 10683 -10218
rect 9187 -10259 10540 -10256
rect 9187 -10262 9589 -10259
rect 9187 -10321 9261 -10262
rect 9320 -10318 9589 -10262
rect 9648 -10260 10540 -10259
rect 9648 -10318 9899 -10260
rect 9320 -10319 9899 -10318
rect 9958 -10319 10225 -10260
rect 10284 -10315 10540 -10260
rect 10599 -10315 10683 -10256
rect 10284 -10319 10683 -10315
rect 9320 -10321 10683 -10319
rect 9187 -10354 10683 -10321
rect 9187 -10357 10645 -10354
<< polycontact >>
rect -2413 1216 -2367 1262
rect -2258 1217 -2212 1263
rect -2864 458 -2818 504
rect -2428 461 -2382 507
rect -2215 457 -2167 504
rect -1782 458 -1736 504
rect -2864 -278 -2818 -232
rect -2428 -278 -2382 -232
rect -2215 -279 -2167 -232
rect -1781 -278 -1735 -232
rect -2863 -1014 -2817 -968
rect -2428 -1017 -2382 -971
rect -2215 -1017 -2167 -970
rect -1781 -1014 -1735 -968
rect -336 796 -290 842
rect 750 798 796 844
rect 99 -106 145 -60
rect 208 -108 254 -62
rect 99 -224 145 -178
rect -330 -1170 -283 -1122
rect 99 -1074 145 -1028
rect 99 -1181 145 -1135
rect 99 -1277 145 -1231
rect 752 -1169 798 -1123
rect 99 -2103 145 -2057
rect 130 -2217 176 -2171
rect -2828 -2793 -2782 -2747
rect -2348 -2793 -2302 -2747
rect -2188 -2793 -2142 -2747
rect -1708 -2793 -1662 -2747
rect 2610 901 2661 952
rect 3488 892 3538 942
rect 4370 901 4421 952
rect 2610 156 2661 207
rect 3489 157 3539 207
rect 4370 156 4421 207
rect 2610 -580 2661 -529
rect 3487 -579 3537 -529
rect 4370 -580 4421 -529
rect 2610 -1317 2661 -1266
rect 3487 -1315 3537 -1265
rect 4370 -1317 4421 -1266
rect 2610 -2053 2661 -2002
rect 3488 -2049 3538 -1999
rect 4370 -2053 4421 -2002
rect 3486 -2784 3536 -2734
rect 5410 901 5461 952
rect 6288 892 6338 942
rect 7170 901 7221 952
rect 5410 156 5461 207
rect 6289 157 6339 207
rect 7170 156 7221 207
rect 5410 -580 5461 -529
rect 6287 -579 6337 -529
rect 7170 -580 7221 -529
rect 5410 -1317 5461 -1266
rect 6287 -1315 6337 -1265
rect 7170 -1317 7221 -1266
rect 5410 -2053 5461 -2002
rect 6288 -2049 6338 -1999
rect 7170 -2053 7221 -2002
rect 6286 -2784 6336 -2734
rect 8210 901 8261 952
rect 9088 892 9138 942
rect 9970 901 10021 952
rect 8210 156 8261 207
rect 9089 157 9139 207
rect 9970 156 10021 207
rect 8210 -580 8261 -529
rect 9087 -579 9137 -529
rect 9970 -580 10021 -529
rect 8210 -1317 8261 -1266
rect 9087 -1315 9137 -1265
rect 9970 -1317 10021 -1266
rect 8210 -2053 8261 -2002
rect 9088 -2049 9138 -1999
rect 9970 -2053 10021 -2002
rect 9086 -2784 9136 -2734
rect -333 -3184 -276 -3132
rect 738 -3182 796 -3128
rect -3061 -3580 -3015 -3534
rect -2829 -3626 -2783 -3580
rect -2668 -3605 -2622 -3559
rect -2508 -3604 -2462 -3558
rect -2348 -3623 -2302 -3577
rect -2188 -3623 -2142 -3577
rect -2028 -3604 -1982 -3558
rect -1868 -3605 -1822 -3559
rect -1707 -3626 -1661 -3580
rect -1468 -3571 -1422 -3525
rect -3068 -4426 -3022 -4380
rect -2667 -4466 -2621 -4420
rect -2507 -4466 -2461 -4420
rect -2029 -4466 -1983 -4420
rect -1869 -4466 -1823 -4420
rect -1468 -4427 -1422 -4381
rect -3068 -5277 -3022 -5231
rect -2829 -5306 -2783 -5260
rect -2668 -5327 -2622 -5281
rect -2508 -5328 -2462 -5282
rect -2348 -5309 -2302 -5263
rect -2188 -5309 -2142 -5263
rect -2028 -5328 -1982 -5282
rect -1868 -5327 -1822 -5281
rect -1707 -5306 -1661 -5260
rect -1468 -5278 -1422 -5232
rect -3068 -6127 -3022 -6081
rect -2828 -6139 -2782 -6093
rect -2348 -6139 -2302 -6093
rect -2188 -6139 -2142 -6093
rect -1708 -6139 -1662 -6093
rect -1468 -6131 -1422 -6085
rect -295 -4304 -230 -4246
rect -154 -4303 -90 -4248
rect -156 -5194 -110 -5148
rect 901 -5198 947 -5152
rect 2583 -4655 2643 -4595
rect 2713 -4655 2773 -4595
rect 1865 -5271 1923 -5213
rect 3421 -5271 3479 -5213
rect 2441 -5381 2501 -5321
rect 1951 -5977 2009 -5919
rect 3075 -5977 3133 -5919
rect 3335 -5977 3393 -5919
rect 5256 -4695 5322 -4629
rect 5394 -4695 5460 -4629
rect 4302 -5262 4352 -5212
rect 4415 -5262 4465 -5212
rect 5302 -5261 5354 -5209
rect 6264 -5264 6314 -5214
rect 6377 -5264 6427 -5214
rect 5256 -5854 5322 -5788
rect 5394 -5854 5460 -5788
rect 9262 -5030 9321 -4971
rect 9576 -5029 9635 -4970
rect 9893 -5026 9952 -4967
rect 10224 -5025 10283 -4966
rect 10543 -5026 10602 -4967
rect 9029 -5805 9080 -5754
rect 10788 -5806 10839 -5755
rect -3049 -7099 -3003 -7053
rect -1449 -7099 -1403 -7053
rect -3049 -7899 -3003 -7853
rect -2251 -7864 -2202 -7815
rect -1449 -7899 -1403 -7853
rect -3049 -8697 -3003 -8651
rect -2251 -8665 -2202 -8616
rect -1449 -8697 -1403 -8651
rect -3049 -9497 -3003 -9451
rect -2252 -9465 -2203 -9416
rect -1449 -9497 -1403 -9451
rect -245 -6909 -199 -6863
rect 878 -6931 924 -6885
rect -243 -7771 -197 -7725
rect 313 -7740 371 -7682
rect 877 -7789 923 -7743
rect 2113 -6835 2174 -6774
rect 2259 -6836 2320 -6775
rect 2873 -6830 2931 -6772
rect 3010 -6831 3068 -6773
rect 9029 -6542 9080 -6491
rect 10788 -6542 10839 -6491
rect 1835 -7469 1893 -7411
rect 3784 -7459 3842 -7401
rect 6135 -7018 6201 -6952
rect 6273 -7018 6339 -6952
rect 4646 -7603 4696 -7553
rect 4759 -7603 4809 -7553
rect 6152 -7603 6202 -7553
rect 6265 -7603 6315 -7553
rect 7654 -7603 7704 -7553
rect 7767 -7603 7817 -7553
rect 9261 -7321 9320 -7262
rect 9589 -7318 9648 -7259
rect 9899 -7319 9958 -7260
rect 10225 -7319 10284 -7260
rect 10540 -7315 10599 -7256
rect 4646 -8142 4696 -8092
rect 4759 -8142 4809 -8092
rect 6150 -8139 6200 -8089
rect 6263 -8139 6313 -8089
rect 7654 -8137 7704 -8087
rect 7767 -8137 7817 -8087
rect 908 -8651 966 -8593
rect -243 -9514 -197 -9468
rect 304 -9569 362 -9511
rect 880 -9520 926 -9474
rect -246 -10367 -200 -10321
rect 957 -10375 1003 -10329
rect 6132 -8749 6198 -8683
rect 6270 -8749 6336 -8683
rect 9262 -8030 9321 -7971
rect 9576 -8029 9635 -7970
rect 9893 -8026 9952 -7967
rect 10224 -8025 10283 -7966
rect 10543 -8026 10602 -7967
rect 9029 -8805 9080 -8754
rect 10788 -8806 10839 -8755
rect 1905 -9203 1957 -9151
rect 2011 -9204 2063 -9152
rect 2223 -9204 2275 -9152
rect 2329 -9205 2381 -9153
rect 2544 -9202 2596 -9150
rect 2650 -9203 2702 -9151
rect 1898 -9553 1950 -9501
rect 2004 -9552 2056 -9500
rect 2216 -9552 2268 -9500
rect 2322 -9551 2374 -9499
rect 2537 -9554 2589 -9502
rect 2643 -9553 2695 -9501
rect 9029 -9542 9080 -9491
rect 10788 -9542 10839 -9491
rect 9261 -10321 9320 -10262
rect 9589 -10318 9648 -10259
rect 9899 -10319 9958 -10260
rect 10225 -10319 10284 -10260
rect 10540 -10315 10599 -10256
<< metal1 >>
rect -2822 1581 -195 1731
rect -3224 1467 12216 1581
rect -3320 1451 12216 1467
rect -3320 1441 -1246 1451
rect -3320 1394 -3294 1441
rect -3247 1395 -3199 1441
rect -3153 1395 -3105 1441
rect -3059 1395 -3011 1441
rect -2965 1395 -2917 1441
rect -2871 1395 -2823 1441
rect -2777 1395 -2729 1441
rect -2683 1395 -2635 1441
rect -2589 1395 -2541 1441
rect -2495 1395 -2447 1441
rect -2401 1395 -2353 1441
rect -2307 1395 -2259 1441
rect -2213 1395 -2165 1441
rect -2119 1395 -2071 1441
rect -2025 1395 -1977 1441
rect -1931 1395 -1883 1441
rect -1837 1395 -1789 1441
rect -1743 1395 -1695 1441
rect -1649 1395 -1601 1441
rect -1555 1395 -1507 1441
rect -1461 1395 -1413 1441
rect -1367 1395 -1319 1441
rect -3247 1394 -1319 1395
rect -1272 1394 -1246 1441
rect -3320 1369 -1246 1394
rect -3320 1346 -3222 1369
rect -3320 1300 -3294 1346
rect -3248 1300 -3222 1346
rect -3320 1252 -3222 1300
rect -3320 1206 -3294 1252
rect -3248 1206 -3222 1252
rect -3320 1158 -3222 1206
rect -3320 1112 -3294 1158
rect -3248 1112 -3222 1158
rect -3320 1064 -3222 1112
rect -3320 1018 -3294 1064
rect -3248 1018 -3222 1064
rect -3320 970 -3222 1018
rect -3320 924 -3294 970
rect -3248 924 -3222 970
rect -3320 876 -3222 924
rect -3320 830 -3294 876
rect -3248 830 -3222 876
rect -3320 782 -3222 830
rect -3320 736 -3294 782
rect -3248 736 -3222 782
rect -3320 688 -3222 736
rect -3320 642 -3294 688
rect -3248 642 -3222 688
rect -3320 594 -3222 642
rect -3320 548 -3294 594
rect -3248 548 -3222 594
rect -3320 500 -3222 548
rect -3320 454 -3294 500
rect -3248 454 -3222 500
rect -3320 406 -3222 454
rect -3320 360 -3294 406
rect -3248 360 -3222 406
rect -3320 312 -3222 360
rect -3320 266 -3294 312
rect -3248 266 -3222 312
rect -3320 218 -3222 266
rect -3320 172 -3294 218
rect -3248 172 -3222 218
rect -3320 124 -3222 172
rect -3320 78 -3294 124
rect -3248 78 -3222 124
rect -3320 30 -3222 78
rect -3320 -16 -3294 30
rect -3248 -16 -3222 30
rect -3320 -64 -3222 -16
rect -3320 -110 -3294 -64
rect -3248 -110 -3222 -64
rect -3320 -158 -3222 -110
rect -3320 -204 -3294 -158
rect -3248 -204 -3222 -158
rect -3320 -252 -3222 -204
rect -3320 -298 -3294 -252
rect -3248 -298 -3222 -252
rect -3320 -346 -3222 -298
rect -3320 -392 -3294 -346
rect -3248 -392 -3222 -346
rect -3320 -440 -3222 -392
rect -3320 -486 -3294 -440
rect -3248 -486 -3222 -440
rect -3320 -534 -3222 -486
rect -3320 -580 -3294 -534
rect -3248 -580 -3222 -534
rect -3320 -628 -3222 -580
rect -3320 -674 -3294 -628
rect -3248 -674 -3222 -628
rect -3320 -722 -3222 -674
rect -3320 -768 -3294 -722
rect -3248 -768 -3222 -722
rect -3320 -816 -3222 -768
rect -3320 -862 -3294 -816
rect -3248 -862 -3222 -816
rect -3320 -910 -3222 -862
rect -3320 -956 -3294 -910
rect -3248 -956 -3222 -910
rect -3320 -1004 -3222 -956
rect -3320 -1050 -3294 -1004
rect -3248 -1050 -3222 -1004
rect -3320 -1098 -3222 -1050
rect -3320 -1144 -3294 -1098
rect -3248 -1144 -3222 -1098
rect -3320 -1192 -3222 -1144
rect -3320 -1238 -3294 -1192
rect -3248 -1238 -3222 -1192
rect -3320 -1286 -3222 -1238
rect -3320 -1332 -3294 -1286
rect -3248 -1332 -3222 -1286
rect -3320 -1380 -3222 -1332
rect -3320 -1426 -3294 -1380
rect -3248 -1426 -3222 -1380
rect -3320 -1474 -3222 -1426
rect -3320 -1520 -3294 -1474
rect -3248 -1520 -3222 -1474
rect -3320 -1568 -3222 -1520
rect -3320 -1614 -3294 -1568
rect -3248 -1614 -3222 -1568
rect -3320 -1662 -3222 -1614
rect -2973 508 -2921 1149
rect -2757 508 -2705 1150
rect -2973 504 -2705 508
rect -2973 458 -2864 504
rect -2818 458 -2705 504
rect -2973 454 -2705 458
rect -2973 -228 -2921 454
rect -2757 -228 -2705 454
rect -2973 -232 -2705 -228
rect -2973 -278 -2864 -232
rect -2818 -278 -2705 -232
rect -2973 -282 -2705 -278
rect -2973 -964 -2921 -282
rect -2757 -964 -2705 -282
rect -2973 -968 -2705 -964
rect -2973 -1014 -2863 -968
rect -2817 -1014 -2705 -968
rect -2973 -1018 -2705 -1014
rect -2973 -1660 -2921 -1018
rect -3320 -1708 -3294 -1662
rect -3248 -1708 -3222 -1662
rect -3320 -1756 -3222 -1708
rect -2757 -1744 -2705 -1018
rect -3320 -1802 -3294 -1756
rect -3248 -1802 -3222 -1756
rect -3320 -1850 -3222 -1802
rect -3320 -1896 -3294 -1850
rect -3248 -1896 -3222 -1850
rect -2791 -1762 -2675 -1744
rect -2791 -1845 -2775 -1762
rect -2691 -1845 -2675 -1762
rect -2791 -1861 -2675 -1845
rect -3320 -1918 -3222 -1896
rect -2541 -1918 -2489 1369
rect -2431 1281 -2312 1320
rect -2431 1266 -2165 1281
rect -2431 1213 -2416 1266
rect -2364 1213 -2304 1266
rect -2252 1263 -2165 1266
rect -2212 1217 -2165 1263
rect -2252 1213 -2165 1217
rect -2431 1201 -2165 1213
rect -2431 507 -2379 1201
rect -2431 461 -2428 507
rect -2382 461 -2379 507
rect -2431 -232 -2379 461
rect -2431 -278 -2428 -232
rect -2382 -278 -2379 -232
rect -2431 -971 -2379 -278
rect -2431 -1017 -2428 -971
rect -2382 -1017 -2379 -971
rect -2431 -1032 -2379 -1017
rect -2325 -1742 -2273 1150
rect -2217 504 -2165 1201
rect -2217 457 -2215 504
rect -2167 457 -2165 504
rect -2217 -232 -2165 457
rect -2217 -279 -2215 -232
rect -2167 -279 -2165 -232
rect -2217 -970 -2165 -279
rect -2217 -1017 -2215 -970
rect -2167 -1017 -2165 -970
rect -2217 -1032 -2165 -1017
rect -2359 -1760 -2243 -1742
rect -2359 -1843 -2343 -1760
rect -2259 -1843 -2243 -1760
rect -2359 -1859 -2243 -1843
rect -2109 -1918 -2057 1369
rect -1344 1346 -1246 1369
rect -1344 1300 -1318 1346
rect -1272 1300 -1246 1346
rect -1344 1252 -1246 1300
rect -1344 1206 -1318 1252
rect -1272 1206 -1246 1252
rect -1344 1158 -1246 1206
rect -1893 507 -1841 1150
rect -1677 507 -1625 1150
rect -1893 504 -1625 507
rect -1893 458 -1782 504
rect -1736 458 -1625 504
rect -1893 453 -1625 458
rect -1893 -228 -1841 453
rect -1677 -228 -1625 453
rect -1893 -232 -1625 -228
rect -1893 -278 -1781 -232
rect -1735 -278 -1625 -232
rect -1893 -282 -1625 -278
rect -1893 -964 -1841 -282
rect -1677 -964 -1625 -282
rect -1893 -968 -1625 -964
rect -1893 -1014 -1781 -968
rect -1735 -1014 -1625 -968
rect -1893 -1018 -1625 -1014
rect -1893 -1742 -1841 -1018
rect -1677 -1659 -1625 -1018
rect -1344 1112 -1318 1158
rect -1272 1112 -1246 1158
rect -1344 1064 -1246 1112
rect -1344 1018 -1318 1064
rect -1272 1018 -1246 1064
rect -1344 970 -1246 1018
rect -1344 924 -1318 970
rect -1272 924 -1246 970
rect -1344 902 -1246 924
rect -1134 1209 -894 1451
rect -485 1209 12216 1451
rect -1134 1173 12216 1209
rect -1134 1039 1063 1173
rect -1134 1013 1244 1039
rect -1134 967 -747 1013
rect -701 967 -653 1013
rect -607 967 -552 1013
rect -506 967 -458 1013
rect -412 967 -362 1013
rect -316 967 -268 1013
rect -222 967 -167 1013
rect -121 967 -73 1013
rect -27 967 21 1013
rect 67 967 115 1013
rect 161 967 216 1013
rect 262 967 310 1013
rect 356 967 406 1013
rect 452 967 500 1013
rect 546 967 601 1013
rect 647 967 695 1013
rect 741 967 789 1013
rect 835 967 883 1013
rect 929 967 984 1013
rect 1030 967 1078 1013
rect 1124 967 1172 1013
rect 1218 970 1244 1013
rect 1858 970 2058 1173
rect 2350 1155 4706 1173
rect 2350 1109 2377 1155
rect 2423 1109 2471 1155
rect 2517 1109 2565 1155
rect 2611 1109 2659 1155
rect 2705 1109 2753 1155
rect 2799 1109 2847 1155
rect 2893 1109 2941 1155
rect 2987 1109 3035 1155
rect 3081 1109 3129 1155
rect 3175 1109 3223 1155
rect 3269 1109 3317 1155
rect 3363 1109 3411 1155
rect 3457 1109 3505 1155
rect 3551 1109 3599 1155
rect 3645 1109 3693 1155
rect 3739 1109 3787 1155
rect 3833 1109 3881 1155
rect 3927 1109 3975 1155
rect 4021 1109 4069 1155
rect 4115 1109 4163 1155
rect 4209 1109 4257 1155
rect 4303 1109 4351 1155
rect 4397 1109 4445 1155
rect 4491 1109 4539 1155
rect 4585 1109 4633 1155
rect 4679 1109 4706 1155
rect 2350 1083 4706 1109
rect 2350 1061 2448 1083
rect 2350 1015 2376 1061
rect 2422 1015 2448 1061
rect 2350 970 2448 1015
rect 1218 967 2448 970
rect -1134 941 2376 967
rect -1134 917 -675 941
rect -1134 902 -747 917
rect -1344 876 -747 902
rect -1344 830 -1318 876
rect -1272 871 -747 876
rect -701 871 -675 917
rect -1272 830 -675 871
rect -255 860 -146 880
rect -1344 823 -675 830
rect -1344 782 -747 823
rect -1344 736 -1318 782
rect -1272 777 -747 782
rect -701 777 -675 823
rect -1272 736 -675 777
rect -1344 727 -675 736
rect -1344 702 -747 727
rect -1344 688 -1246 702
rect -1344 642 -1318 688
rect -1272 642 -1246 688
rect -1344 594 -1246 642
rect -1344 548 -1318 594
rect -1272 548 -1246 594
rect -1344 502 -1246 548
rect -1134 502 -894 702
rect -773 681 -747 702
rect -701 681 -675 727
rect -440 842 -146 860
rect -440 796 -336 842
rect -290 796 -146 842
rect -440 780 -146 796
rect -440 712 -394 780
rect -255 762 -146 780
rect -773 633 -675 681
rect -773 587 -747 633
rect -701 587 -675 633
rect -773 539 -675 587
rect -773 502 -747 539
rect -1344 500 -747 502
rect -1344 454 -1318 500
rect -1272 493 -747 500
rect -701 493 -675 539
rect -1272 454 -675 493
rect -1344 438 -675 454
rect -1344 406 -747 438
rect -1344 360 -1318 406
rect -1272 392 -747 406
rect -701 392 -675 438
rect -1272 360 -675 392
rect -1344 344 -675 360
rect -1344 312 -747 344
rect -1344 266 -1318 312
rect -1272 302 -747 312
rect -1272 266 -1246 302
rect -1344 218 -1246 266
rect -1344 172 -1318 218
rect -1272 172 -1246 218
rect -1344 124 -1246 172
rect -1344 78 -1318 124
rect -1272 102 -1246 124
rect -1134 102 -894 302
rect -773 298 -747 302
rect -701 298 -675 344
rect -235 337 -173 762
rect -8 689 38 941
rect 199 550 261 719
rect 424 712 470 941
rect 1146 921 2376 941
rect 2422 921 2448 967
rect 1146 917 2448 921
rect 608 864 712 876
rect 1146 871 1172 917
rect 1218 873 2448 917
rect 1218 871 2376 873
rect 608 844 902 864
rect 608 798 750 844
rect 796 798 902 844
rect 608 782 902 798
rect 608 773 712 782
rect 175 535 286 550
rect 175 457 191 535
rect 271 457 286 535
rect 175 443 286 457
rect -773 248 -675 298
rect -773 202 -747 248
rect -701 202 -675 248
rect -259 323 -147 337
rect -259 233 -244 323
rect -162 233 -147 323
rect -259 219 -147 233
rect -773 154 -675 202
rect -773 108 -747 154
rect -701 108 -675 154
rect -773 102 -675 108
rect -235 107 -173 219
rect -1272 78 -675 102
rect -1344 53 -675 78
rect -1344 30 -747 53
rect -1344 -16 -1318 30
rect -1272 7 -747 30
rect -701 7 -675 53
rect -1272 -16 -675 7
rect -1344 -41 -675 -16
rect -1344 -64 -747 -41
rect -1344 -110 -1318 -64
rect -1272 -87 -747 -64
rect -701 -87 -675 -41
rect -1272 -98 -675 -87
rect -1272 -110 -1246 -98
rect -1344 -158 -1246 -110
rect -1344 -204 -1318 -158
rect -1272 -204 -1246 -158
rect -1344 -252 -1246 -204
rect -1344 -298 -1318 -252
rect -1272 -298 -1246 -252
rect -1134 -298 -894 -98
rect -773 -135 -675 -98
rect -773 -181 -747 -135
rect -701 -181 -675 -135
rect -260 -66 -144 -44
rect -260 -145 -242 -66
rect -160 -145 -144 -66
rect -260 -160 -144 -145
rect -773 -229 -675 -181
rect -773 -275 -747 -229
rect -701 -275 -675 -229
rect -773 -298 -675 -275
rect -1344 -330 -675 -298
rect -224 -326 -178 -160
rect -8 -326 38 116
rect 199 106 261 443
rect 631 325 693 773
rect 856 712 902 782
rect 1146 827 2376 871
rect 2422 827 2448 873
rect 1146 816 2448 827
rect 1146 770 1172 816
rect 1218 779 2448 816
rect 1218 770 2376 779
rect 1146 722 1244 770
rect 1146 676 1172 722
rect 1218 676 1244 722
rect 1146 628 1244 676
rect 1146 582 1172 628
rect 1218 582 1244 628
rect 1146 570 1244 582
rect 1858 570 2058 770
rect 2350 733 2376 770
rect 2422 733 2448 779
rect 2350 685 2448 733
rect 2350 639 2376 685
rect 2422 639 2448 685
rect 2350 591 2448 639
rect 2350 570 2376 591
rect 1146 545 2376 570
rect 2422 545 2448 591
rect 1146 534 2448 545
rect 1146 488 1172 534
rect 1218 497 2448 534
rect 1218 488 2376 497
rect 1146 451 2376 488
rect 2422 451 2448 497
rect 1146 433 2448 451
rect 1146 387 1172 433
rect 1218 403 2448 433
rect 1218 387 2376 403
rect 1146 370 2376 387
rect 1146 339 1244 370
rect 612 311 713 325
rect 612 237 625 311
rect 700 237 713 311
rect 612 224 713 237
rect 1146 293 1172 339
rect 1218 293 1244 339
rect 1146 243 1244 293
rect 96 -60 276 -36
rect 96 -106 99 -60
rect 145 -62 276 -60
rect 145 -106 208 -62
rect 96 -108 208 -106
rect 254 -108 276 -62
rect 96 -122 276 -108
rect 96 -178 148 -122
rect 96 -224 99 -178
rect 145 -224 148 -178
rect -1344 -346 -747 -330
rect -1344 -392 -1318 -346
rect -1272 -376 -747 -346
rect -701 -376 -675 -330
rect -1272 -392 -675 -376
rect -1344 -424 -675 -392
rect -1344 -440 -747 -424
rect -1344 -486 -1318 -440
rect -1272 -470 -747 -440
rect -701 -470 -675 -424
rect -1272 -486 -675 -470
rect -1344 -498 -675 -486
rect -1344 -534 -1246 -498
rect -1344 -580 -1318 -534
rect -1272 -580 -1246 -534
rect -1344 -628 -1246 -580
rect -1344 -674 -1318 -628
rect -1272 -674 -1246 -628
rect -1344 -698 -1246 -674
rect -1134 -698 -894 -498
rect -773 -520 -675 -498
rect -773 -566 -747 -520
rect -701 -566 -675 -520
rect -257 -456 -146 -437
rect -257 -535 -242 -456
rect -160 -535 -146 -456
rect -257 -550 -146 -535
rect -773 -614 -675 -566
rect -773 -660 -747 -614
rect -701 -660 -675 -614
rect -773 -698 -675 -660
rect -1344 -715 -675 -698
rect -1344 -722 -747 -715
rect -1344 -768 -1318 -722
rect -1272 -761 -747 -722
rect -701 -761 -675 -715
rect -1272 -768 -675 -761
rect -1344 -809 -675 -768
rect -1344 -816 -747 -809
rect -1344 -862 -1318 -816
rect -1272 -855 -747 -816
rect -701 -855 -675 -809
rect -1272 -862 -675 -855
rect -1344 -898 -675 -862
rect -1344 -910 -1246 -898
rect -1344 -956 -1318 -910
rect -1272 -956 -1246 -910
rect -1344 -1004 -1246 -956
rect -1344 -1050 -1318 -1004
rect -1272 -1050 -1246 -1004
rect -1344 -1098 -1246 -1050
rect -1134 -1098 -894 -898
rect -773 -903 -675 -898
rect -773 -949 -747 -903
rect -701 -949 -675 -903
rect -773 -997 -675 -949
rect -773 -1043 -747 -997
rect -701 -1043 -675 -997
rect -773 -1098 -675 -1043
rect -1344 -1144 -1318 -1098
rect -1272 -1144 -747 -1098
rect -701 -1144 -675 -1098
rect -1344 -1192 -675 -1144
rect -1344 -1238 -1318 -1192
rect -1272 -1238 -747 -1192
rect -701 -1238 -675 -1192
rect -1344 -1286 -675 -1238
rect -1344 -1332 -1318 -1286
rect -1272 -1288 -675 -1286
rect -1272 -1298 -747 -1288
rect -1272 -1332 -1246 -1298
rect -1344 -1380 -1246 -1332
rect -1344 -1426 -1318 -1380
rect -1272 -1426 -1246 -1380
rect -1344 -1474 -1246 -1426
rect -1344 -1520 -1318 -1474
rect -1272 -1498 -1246 -1474
rect -1134 -1498 -894 -1298
rect -773 -1334 -747 -1298
rect -701 -1334 -675 -1288
rect -773 -1382 -675 -1334
rect -440 -1121 -394 -922
rect -224 -1121 -178 -922
rect -440 -1122 -178 -1121
rect -440 -1170 -330 -1122
rect -283 -1170 -178 -1122
rect -440 -1172 -178 -1170
rect -440 -1366 -394 -1172
rect -224 -1366 -178 -1172
rect -8 -1366 38 -922
rect 96 -1028 148 -224
rect 96 -1074 99 -1028
rect 145 -1074 148 -1028
rect 96 -1135 148 -1074
rect 96 -1181 99 -1135
rect 145 -1181 148 -1135
rect 96 -1231 148 -1181
rect 96 -1277 99 -1231
rect 145 -1277 148 -1231
rect -773 -1428 -747 -1382
rect -701 -1428 -675 -1382
rect -773 -1476 -675 -1428
rect -773 -1498 -747 -1476
rect -1272 -1520 -747 -1498
rect -1344 -1522 -747 -1520
rect -701 -1522 -675 -1476
rect -1344 -1568 -675 -1522
rect -1344 -1614 -1318 -1568
rect -1272 -1577 -675 -1568
rect -1272 -1614 -747 -1577
rect -1344 -1623 -747 -1614
rect -701 -1623 -675 -1577
rect -1344 -1662 -675 -1623
rect -1344 -1708 -1318 -1662
rect -1272 -1671 -675 -1662
rect -1272 -1698 -747 -1671
rect -1272 -1708 -1246 -1698
rect -1926 -1760 -1810 -1742
rect -1926 -1843 -1910 -1760
rect -1826 -1843 -1810 -1760
rect -1926 -1859 -1810 -1843
rect -1344 -1756 -1246 -1708
rect -1344 -1802 -1318 -1756
rect -1272 -1802 -1246 -1756
rect -1344 -1850 -1246 -1802
rect -1344 -1896 -1318 -1850
rect -1272 -1896 -1246 -1850
rect -1344 -1918 -1246 -1896
rect -3320 -1944 -1246 -1918
rect -3320 -1990 -3293 -1944
rect -3247 -1990 -3199 -1944
rect -3153 -1990 -3105 -1944
rect -3059 -1990 -3011 -1944
rect -2965 -1990 -2917 -1944
rect -2871 -1990 -2823 -1944
rect -2777 -1990 -2729 -1944
rect -2683 -1990 -2635 -1944
rect -2589 -1990 -2541 -1944
rect -2495 -1990 -2447 -1944
rect -2401 -1990 -2353 -1944
rect -2307 -1990 -2259 -1944
rect -2213 -1990 -2165 -1944
rect -2119 -1990 -2071 -1944
rect -2025 -1990 -1977 -1944
rect -1931 -1990 -1883 -1944
rect -1837 -1990 -1789 -1944
rect -1743 -1990 -1695 -1944
rect -1649 -1990 -1601 -1944
rect -1555 -1990 -1507 -1944
rect -1461 -1990 -1413 -1944
rect -1367 -1990 -1319 -1944
rect -1273 -1990 -1246 -1944
rect -3320 -2016 -1246 -1990
rect -3159 -2168 -2959 -2016
rect -2759 -2168 -2559 -2016
rect -2359 -2168 -2159 -2016
rect -1959 -2168 -1759 -2016
rect -1559 -2168 -1359 -2016
rect -1134 -2168 -894 -1698
rect -773 -1717 -747 -1698
rect -701 -1717 -675 -1671
rect -773 -1767 -675 -1717
rect -773 -1813 -747 -1767
rect -701 -1813 -675 -1767
rect -773 -1861 -675 -1813
rect -773 -1907 -747 -1861
rect -701 -1907 -675 -1861
rect -773 -1962 -675 -1907
rect -773 -2008 -747 -1962
rect -701 -2008 -675 -1962
rect -773 -2056 -675 -2008
rect -773 -2102 -747 -2056
rect -701 -2102 -675 -2056
rect -773 -2150 -675 -2102
rect -773 -2168 -747 -2150
rect -3159 -2196 -747 -2168
rect -701 -2196 -675 -2150
rect -3159 -2244 -675 -2196
rect -3159 -2290 -747 -2244
rect -701 -2290 -675 -2244
rect -3159 -2345 -675 -2290
rect -3159 -2391 -747 -2345
rect -701 -2391 -675 -2345
rect -3159 -2408 -675 -2391
rect -4059 -2471 -3700 -2447
rect -4059 -2591 -4042 -2471
rect -3919 -2591 -3842 -2471
rect -3719 -2591 -3700 -2471
rect -3159 -2567 -2959 -2408
rect -2759 -2567 -2559 -2408
rect -2359 -2567 -2159 -2408
rect -1959 -2567 -1759 -2408
rect -1559 -2567 -1359 -2408
rect -4059 -2608 -3700 -2591
rect -3293 -2593 -1219 -2567
rect -3293 -2640 -3267 -2593
rect -3220 -2639 -3172 -2593
rect -3126 -2639 -3078 -2593
rect -3032 -2639 -2984 -2593
rect -2938 -2639 -2890 -2593
rect -2844 -2639 -2796 -2593
rect -2750 -2639 -2702 -2593
rect -2656 -2639 -2608 -2593
rect -2562 -2639 -2514 -2593
rect -2468 -2639 -2420 -2593
rect -2374 -2639 -2326 -2593
rect -2280 -2639 -2232 -2593
rect -2186 -2639 -2138 -2593
rect -2092 -2639 -2044 -2593
rect -1998 -2639 -1950 -2593
rect -1904 -2639 -1856 -2593
rect -1810 -2639 -1762 -2593
rect -1716 -2639 -1668 -2593
rect -1622 -2639 -1574 -2593
rect -1528 -2639 -1480 -2593
rect -1434 -2639 -1386 -2593
rect -1340 -2639 -1292 -2593
rect -3220 -2640 -1292 -2639
rect -1245 -2640 -1219 -2593
rect -3293 -2650 -1219 -2640
rect -1134 -2650 -894 -2408
rect -773 -2439 -675 -2408
rect -773 -2485 -747 -2439
rect -701 -2485 -675 -2439
rect -773 -2535 -675 -2485
rect -773 -2581 -747 -2535
rect -701 -2581 -675 -2535
rect -773 -2629 -675 -2581
rect -773 -2650 -747 -2629
rect -3293 -2665 -747 -2650
rect -3293 -2688 -3195 -2665
rect -4063 -2723 -3687 -2693
rect -4063 -2843 -4039 -2723
rect -3916 -2843 -3839 -2723
rect -3716 -2843 -3687 -2723
rect -4063 -2868 -3687 -2843
rect -3293 -2734 -3267 -2688
rect -3221 -2734 -3195 -2688
rect -1317 -2675 -747 -2665
rect -701 -2675 -675 -2629
rect -1317 -2688 -675 -2675
rect -3293 -2782 -3195 -2734
rect -1750 -2730 -1634 -2712
rect -1750 -2743 -1734 -2730
rect -3293 -2828 -3267 -2782
rect -3221 -2828 -3195 -2782
rect -2849 -2747 -1734 -2743
rect -2849 -2793 -2828 -2747
rect -2782 -2793 -2348 -2747
rect -2302 -2793 -2188 -2747
rect -2142 -2793 -1734 -2747
rect -2849 -2799 -1734 -2793
rect -1750 -2810 -1734 -2799
rect -1654 -2810 -1634 -2730
rect -1750 -2820 -1634 -2810
rect -1317 -2734 -1291 -2688
rect -1245 -2730 -675 -2688
rect -1245 -2734 -747 -2730
rect -1317 -2776 -747 -2734
rect -701 -2776 -675 -2730
rect -1317 -2782 -675 -2776
rect -3293 -2876 -3195 -2828
rect -3293 -2922 -3267 -2876
rect -3221 -2922 -3195 -2876
rect -3293 -2970 -3195 -2922
rect -1317 -2828 -1291 -2782
rect -1245 -2824 -675 -2782
rect -1245 -2828 -747 -2824
rect -1317 -2850 -747 -2828
rect -1317 -2876 -1219 -2850
rect -1317 -2922 -1291 -2876
rect -1245 -2922 -1219 -2876
rect -3293 -3016 -3267 -2970
rect -3221 -3016 -3195 -2970
rect -3293 -3064 -3195 -3016
rect -2614 -2953 -2517 -2940
rect -2614 -3034 -2599 -2953
rect -2531 -3034 -2517 -2953
rect -2614 -3047 -2517 -3034
rect -1978 -2955 -1881 -2942
rect -1978 -3036 -1963 -2955
rect -1895 -3036 -1881 -2955
rect -1978 -3049 -1881 -3036
rect -1317 -2970 -1219 -2922
rect -1317 -3016 -1291 -2970
rect -1245 -3016 -1219 -2970
rect -3293 -3110 -3267 -3064
rect -3221 -3110 -3195 -3064
rect -1317 -3050 -1219 -3016
rect -1134 -3050 -894 -2850
rect -773 -2870 -747 -2850
rect -701 -2870 -675 -2824
rect -773 -2918 -675 -2870
rect -773 -2964 -747 -2918
rect -701 -2964 -675 -2918
rect -773 -3012 -675 -2964
rect -773 -3050 -747 -3012
rect -1317 -3058 -747 -3050
rect -701 -3058 -675 -3012
rect -1317 -3064 -675 -3058
rect -3293 -3158 -3195 -3110
rect -3293 -3204 -3267 -3158
rect -3221 -3204 -3195 -3158
rect -2774 -3109 -2677 -3096
rect -2774 -3190 -2759 -3109
rect -2691 -3190 -2677 -3109
rect -2774 -3203 -2677 -3190
rect -2454 -3101 -2357 -3088
rect -2454 -3182 -2439 -3101
rect -2371 -3182 -2357 -3101
rect -2454 -3195 -2357 -3182
rect -2133 -3109 -2036 -3096
rect -2133 -3190 -2118 -3109
rect -2050 -3190 -2036 -3109
rect -2133 -3203 -2036 -3190
rect -1818 -3105 -1721 -3092
rect -1818 -3186 -1803 -3105
rect -1735 -3186 -1721 -3105
rect -1818 -3199 -1721 -3186
rect -1317 -3110 -1291 -3064
rect -1245 -3110 -675 -3064
rect -1317 -3113 -675 -3110
rect -1317 -3158 -747 -3113
rect -3293 -3252 -3195 -3204
rect -1317 -3204 -1291 -3158
rect -1245 -3159 -747 -3158
rect -701 -3159 -675 -3113
rect -1245 -3204 -675 -3159
rect -440 -3114 -394 -3000
rect -236 -3092 -168 -2402
rect -8 -2404 38 -1962
rect 96 -2057 148 -1277
rect 204 -1088 270 -321
rect 424 -326 470 116
rect 631 110 693 224
rect 1146 197 1172 243
rect 1218 197 1244 243
rect 1146 170 1244 197
rect 1858 170 2058 370
rect 2350 357 2376 370
rect 2422 357 2448 403
rect 2350 309 2448 357
rect 2350 263 2376 309
rect 2422 263 2448 309
rect 2350 215 2448 263
rect 2350 170 2376 215
rect 1146 169 2376 170
rect 2422 169 2448 215
rect 1146 149 2448 169
rect 1146 103 1172 149
rect 1218 121 2448 149
rect 1218 103 2376 121
rect 1146 75 2376 103
rect 2422 75 2448 121
rect 1146 48 2448 75
rect 1146 2 1172 48
rect 1218 27 2448 48
rect 1218 2 2376 27
rect 1146 -19 2376 2
rect 2422 -19 2448 27
rect 1146 -30 2448 -19
rect 1146 -46 1244 -30
rect 605 -71 721 -51
rect 605 -150 621 -71
rect 703 -150 721 -71
rect 605 -167 721 -150
rect 1146 -92 1172 -46
rect 1218 -92 1244 -46
rect 1146 -140 1244 -92
rect 640 -326 686 -167
rect 1146 -186 1172 -140
rect 1218 -186 1244 -140
rect 1146 -230 1244 -186
rect 1858 -230 2058 -30
rect 2350 -67 2448 -30
rect 2350 -113 2376 -67
rect 2422 -113 2448 -67
rect 2350 -161 2448 -113
rect 2350 -207 2376 -161
rect 2422 -207 2448 -161
rect 2350 -230 2448 -207
rect 1146 -234 2448 -230
rect 1146 -280 1172 -234
rect 1218 -255 2448 -234
rect 1218 -280 2376 -255
rect 1146 -301 2376 -280
rect 2422 -301 2448 -255
rect 1146 -335 2448 -301
rect 1146 -381 1172 -335
rect 1218 -349 2448 -335
rect 1218 -381 2376 -349
rect 1146 -395 2376 -381
rect 2422 -395 2448 -349
rect 1146 -429 2448 -395
rect 609 -455 718 -441
rect 609 -534 623 -455
rect 705 -534 718 -455
rect 609 -549 718 -534
rect 1146 -475 1172 -429
rect 1218 -430 2448 -429
rect 1218 -475 1244 -430
rect 1146 -525 1244 -475
rect 1146 -571 1172 -525
rect 1218 -571 1244 -525
rect 1146 -619 1244 -571
rect 1146 -665 1172 -619
rect 1218 -630 1244 -619
rect 1858 -630 2058 -430
rect 2350 -443 2448 -430
rect 2350 -489 2376 -443
rect 2422 -489 2448 -443
rect 2350 -537 2448 -489
rect 2350 -583 2376 -537
rect 2422 -583 2448 -537
rect 2350 -630 2448 -583
rect 1218 -631 2448 -630
rect 1218 -665 2376 -631
rect 1146 -677 2376 -665
rect 2422 -677 2448 -631
rect 1146 -720 2448 -677
rect 1146 -766 1172 -720
rect 1218 -725 2448 -720
rect 1218 -766 2376 -725
rect 1146 -771 2376 -766
rect 2422 -771 2448 -725
rect 1146 -814 2448 -771
rect 1146 -860 1172 -814
rect 1218 -819 2448 -814
rect 1218 -830 2376 -819
rect 1218 -860 1244 -830
rect 1146 -908 1244 -860
rect 204 -1109 366 -1088
rect 204 -1188 270 -1109
rect 353 -1188 366 -1109
rect 204 -1204 366 -1188
rect 204 -1967 270 -1204
rect 424 -1366 470 -922
rect 640 -1121 686 -922
rect 856 -1121 902 -922
rect 640 -1123 902 -1121
rect 640 -1169 752 -1123
rect 798 -1169 902 -1123
rect 640 -1172 902 -1169
rect 640 -1366 686 -1172
rect 856 -1366 902 -1172
rect 1146 -954 1172 -908
rect 1218 -954 1244 -908
rect 1146 -1004 1244 -954
rect 1146 -1050 1172 -1004
rect 1218 -1030 1244 -1004
rect 1858 -1030 2058 -830
rect 2350 -865 2376 -830
rect 2422 -865 2448 -819
rect 2350 -913 2448 -865
rect 2350 -959 2376 -913
rect 2422 -959 2448 -913
rect 2350 -1007 2448 -959
rect 2350 -1030 2376 -1007
rect 1218 -1050 2376 -1030
rect 1146 -1053 2376 -1050
rect 2422 -1053 2448 -1007
rect 1146 -1098 2448 -1053
rect 1146 -1144 1172 -1098
rect 1218 -1101 2448 -1098
rect 1218 -1144 2376 -1101
rect 1146 -1147 2376 -1144
rect 2422 -1147 2448 -1101
rect 1146 -1195 2448 -1147
rect 1146 -1199 2376 -1195
rect 1146 -1245 1172 -1199
rect 1218 -1230 2376 -1199
rect 1218 -1245 1244 -1230
rect 1146 -1293 1244 -1245
rect 1146 -1339 1172 -1293
rect 1218 -1339 1244 -1293
rect 1146 -1387 1244 -1339
rect 1146 -1433 1172 -1387
rect 1218 -1430 1244 -1387
rect 1858 -1430 2058 -1230
rect 2350 -1241 2376 -1230
rect 2422 -1241 2448 -1195
rect 2350 -1289 2448 -1241
rect 2350 -1335 2376 -1289
rect 2422 -1335 2448 -1289
rect 2350 -1383 2448 -1335
rect 2350 -1429 2376 -1383
rect 2422 -1429 2448 -1383
rect 2350 -1430 2448 -1429
rect 1218 -1433 2448 -1430
rect 1146 -1477 2448 -1433
rect 1146 -1481 2376 -1477
rect 1146 -1527 1172 -1481
rect 1218 -1523 2376 -1481
rect 2422 -1523 2448 -1477
rect 1218 -1527 2448 -1523
rect 1146 -1571 2448 -1527
rect 1146 -1582 2376 -1571
rect 1146 -1628 1172 -1582
rect 1218 -1617 2376 -1582
rect 2422 -1617 2448 -1571
rect 1218 -1628 2448 -1617
rect 1146 -1630 2448 -1628
rect 1146 -1676 1244 -1630
rect 1146 -1722 1172 -1676
rect 1218 -1722 1244 -1676
rect 1146 -1772 1244 -1722
rect 1146 -1818 1172 -1772
rect 1218 -1818 1244 -1772
rect 1146 -1830 1244 -1818
rect 1858 -1830 2058 -1630
rect 2350 -1665 2448 -1630
rect 2350 -1711 2376 -1665
rect 2422 -1711 2448 -1665
rect 2350 -1759 2448 -1711
rect 2350 -1805 2376 -1759
rect 2422 -1805 2448 -1759
rect 2350 -1830 2448 -1805
rect 1146 -1853 2448 -1830
rect 1146 -1866 2376 -1853
rect 1146 -1912 1172 -1866
rect 1218 -1899 2376 -1866
rect 2422 -1899 2448 -1853
rect 1218 -1912 2448 -1899
rect 1146 -1947 2448 -1912
rect 96 -2103 99 -2057
rect 145 -2103 148 -2057
rect 96 -2139 148 -2103
rect 96 -2154 281 -2139
rect 96 -2171 185 -2154
rect 96 -2217 130 -2171
rect 176 -2217 185 -2171
rect 96 -2235 185 -2217
rect 266 -2235 281 -2154
rect 96 -2237 281 -2235
rect 171 -2252 281 -2237
rect 424 -2404 470 -1962
rect 1146 -1967 2376 -1947
rect 1146 -2013 1172 -1967
rect 1218 -1993 2376 -1967
rect 2422 -1993 2448 -1947
rect 1218 -2013 2448 -1993
rect 1146 -2030 2448 -2013
rect 1146 -2061 1244 -2030
rect 1146 -2107 1172 -2061
rect 1218 -2107 1244 -2061
rect 1146 -2155 1244 -2107
rect 1146 -2201 1172 -2155
rect 1218 -2201 1244 -2155
rect 1146 -2230 1244 -2201
rect 1858 -2230 2058 -2030
rect 2350 -2041 2448 -2030
rect 2350 -2087 2376 -2041
rect 2422 -2087 2448 -2041
rect 2350 -2135 2448 -2087
rect 2350 -2181 2376 -2135
rect 2422 -2181 2448 -2135
rect 2350 -2229 2448 -2181
rect 2350 -2230 2376 -2229
rect 1146 -2249 2376 -2230
rect 1146 -2295 1172 -2249
rect 1218 -2275 2376 -2249
rect 2422 -2275 2448 -2229
rect 1218 -2295 2448 -2275
rect 1146 -2323 2448 -2295
rect 1146 -2350 2376 -2323
rect 1146 -2396 1172 -2350
rect 1218 -2369 2376 -2350
rect 2422 -2369 2448 -2323
rect 1218 -2396 2448 -2369
rect -264 -3114 -144 -3092
rect -440 -3117 -144 -3114
rect -440 -3132 -243 -3117
rect -440 -3184 -333 -3132
rect -276 -3184 -243 -3132
rect -440 -3197 -243 -3184
rect -163 -3197 -144 -3117
rect -440 -3198 -144 -3197
rect -1317 -3207 -675 -3204
rect -3293 -3298 -3267 -3252
rect -3221 -3298 -3195 -3252
rect -3293 -3346 -3195 -3298
rect -3293 -3392 -3267 -3346
rect -3221 -3392 -3195 -3346
rect -3094 -3260 -2997 -3247
rect -3094 -3341 -3079 -3260
rect -3011 -3341 -2997 -3260
rect -3094 -3354 -2997 -3341
rect -2937 -3262 -2840 -3249
rect -2937 -3343 -2922 -3262
rect -2854 -3343 -2840 -3262
rect -2937 -3356 -2840 -3343
rect -2294 -3261 -2197 -3248
rect -2294 -3342 -2279 -3261
rect -2211 -3342 -2197 -3261
rect -2294 -3355 -2197 -3342
rect -1658 -3264 -1561 -3251
rect -1658 -3345 -1643 -3264
rect -1575 -3345 -1561 -3264
rect -1658 -3358 -1561 -3345
rect -1492 -3260 -1395 -3247
rect -1492 -3341 -1477 -3260
rect -1409 -3341 -1395 -3260
rect -1492 -3354 -1395 -3341
rect -1317 -3250 -747 -3207
rect -1317 -3252 -1219 -3250
rect -1317 -3298 -1291 -3252
rect -1245 -3298 -1219 -3252
rect -1317 -3346 -1219 -3298
rect -3293 -3440 -3195 -3392
rect -3293 -3486 -3267 -3440
rect -3221 -3486 -3195 -3440
rect -1317 -3392 -1291 -3346
rect -1245 -3392 -1219 -3346
rect -1317 -3440 -1219 -3392
rect -3293 -3534 -3195 -3486
rect -3068 -3509 -3022 -3461
rect -3293 -3580 -3267 -3534
rect -3221 -3580 -3195 -3534
rect -3293 -3628 -3195 -3580
rect -3077 -3534 -3003 -3509
rect -1468 -3515 -1422 -3463
rect -1317 -3486 -1291 -3440
rect -1245 -3486 -1219 -3440
rect -3077 -3580 -3061 -3534
rect -3015 -3580 -3003 -3534
rect -1480 -3525 -1410 -3515
rect -3077 -3595 -3003 -3580
rect -2854 -3549 -2750 -3538
rect -3293 -3674 -3267 -3628
rect -3221 -3674 -3195 -3628
rect -2854 -3629 -2844 -3549
rect -2762 -3563 -2750 -3549
rect -2684 -3559 -2606 -3542
rect -2684 -3563 -2668 -3559
rect -2762 -3605 -2668 -3563
rect -2622 -3563 -2606 -3559
rect -2524 -3558 -2446 -3542
rect -2524 -3563 -2508 -3558
rect -2622 -3604 -2508 -3563
rect -2462 -3563 -2446 -3558
rect -2044 -3558 -1966 -3542
rect -2044 -3563 -2028 -3558
rect -2462 -3577 -2028 -3563
rect -2462 -3604 -2348 -3577
rect -2622 -3605 -2348 -3604
rect -2762 -3619 -2348 -3605
rect -2762 -3629 -2750 -3619
rect -2854 -3639 -2750 -3629
rect -2363 -3623 -2348 -3619
rect -2302 -3619 -2188 -3577
rect -2302 -3623 -2285 -3619
rect -2845 -3640 -2767 -3639
rect -2363 -3640 -2285 -3623
rect -2205 -3623 -2188 -3619
rect -2142 -3604 -2028 -3577
rect -1982 -3563 -1966 -3558
rect -1884 -3559 -1806 -3542
rect -1884 -3563 -1868 -3559
rect -1982 -3604 -1868 -3563
rect -2142 -3605 -1868 -3604
rect -1822 -3563 -1806 -3559
rect -1822 -3580 -1645 -3563
rect -1822 -3605 -1707 -3580
rect -2142 -3619 -1707 -3605
rect -2142 -3623 -2127 -3619
rect -2205 -3640 -2127 -3623
rect -1723 -3626 -1707 -3619
rect -1661 -3626 -1645 -3580
rect -1480 -3571 -1468 -3525
rect -1422 -3571 -1410 -3525
rect -1480 -3583 -1410 -3571
rect -1317 -3534 -1219 -3486
rect -1317 -3580 -1291 -3534
rect -1245 -3580 -1219 -3534
rect -1723 -3640 -1645 -3626
rect -1317 -3628 -1219 -3580
rect -3293 -3722 -3195 -3674
rect -3293 -3768 -3267 -3722
rect -3221 -3768 -3195 -3722
rect -3293 -3816 -3195 -3768
rect -1317 -3674 -1291 -3628
rect -1245 -3674 -1219 -3628
rect -1317 -3722 -1219 -3674
rect -1317 -3768 -1291 -3722
rect -1245 -3768 -1219 -3722
rect -3293 -3862 -3267 -3816
rect -3221 -3862 -3195 -3816
rect -3293 -3910 -3195 -3862
rect -2615 -3811 -2518 -3798
rect -2615 -3892 -2600 -3811
rect -2532 -3892 -2518 -3811
rect -2615 -3905 -2518 -3892
rect -1972 -3805 -1875 -3792
rect -1972 -3886 -1957 -3805
rect -1889 -3886 -1875 -3805
rect -1972 -3899 -1875 -3886
rect -1317 -3816 -1219 -3768
rect -1134 -3567 -894 -3250
rect -773 -3253 -747 -3250
rect -701 -3253 -675 -3207
rect -264 -3216 -144 -3198
rect -773 -3277 -675 -3253
rect -8 -3277 38 -2999
rect 208 -3100 254 -3000
rect 174 -3117 285 -3100
rect 174 -3200 189 -3117
rect 271 -3200 285 -3117
rect 174 -3214 285 -3200
rect 424 -3277 470 -2999
rect 628 -3096 696 -2401
rect 1146 -2417 2448 -2396
rect 1146 -2430 2376 -2417
rect 1146 -2444 1244 -2430
rect 1146 -2490 1172 -2444
rect 1218 -2490 1244 -2444
rect 1146 -2540 1244 -2490
rect 1146 -2586 1172 -2540
rect 1218 -2586 1244 -2540
rect 1146 -2630 1244 -2586
rect 1858 -2630 2058 -2430
rect 2350 -2463 2376 -2430
rect 2422 -2463 2448 -2417
rect 2350 -2511 2448 -2463
rect 2350 -2557 2376 -2511
rect 2422 -2557 2448 -2511
rect 2350 -2605 2448 -2557
rect 2350 -2630 2376 -2605
rect 1146 -2634 2376 -2630
rect 1146 -2680 1172 -2634
rect 1218 -2651 2376 -2634
rect 2422 -2651 2448 -2605
rect 1218 -2680 2448 -2651
rect 1146 -2699 2448 -2680
rect 1146 -2735 2376 -2699
rect 1146 -2781 1172 -2735
rect 1218 -2745 2376 -2735
rect 2422 -2745 2448 -2699
rect 1218 -2781 2448 -2745
rect 1146 -2793 2448 -2781
rect 1146 -2829 2376 -2793
rect 1146 -2875 1172 -2829
rect 1218 -2830 2376 -2829
rect 1218 -2875 1244 -2830
rect 1146 -2923 1244 -2875
rect 1146 -2969 1172 -2923
rect 1218 -2969 1244 -2923
rect 607 -3110 718 -3096
rect 607 -3196 620 -3110
rect 704 -3112 718 -3110
rect 856 -3112 902 -3000
rect 704 -3128 902 -3112
rect 704 -3182 738 -3128
rect 796 -3182 902 -3128
rect 704 -3196 902 -3182
rect 607 -3198 902 -3196
rect 1146 -3019 1244 -2969
rect 1146 -3065 1172 -3019
rect 1218 -3065 1244 -3019
rect 1146 -3113 1244 -3065
rect 1146 -3159 1172 -3113
rect 1218 -3159 1244 -3113
rect 607 -3210 718 -3198
rect 1146 -3207 1244 -3159
rect 1146 -3253 1172 -3207
rect 1218 -3253 1244 -3207
rect 1146 -3277 1244 -3253
rect -773 -3303 1244 -3277
rect -773 -3349 -747 -3303
rect -701 -3349 -653 -3303
rect -607 -3349 -552 -3303
rect -506 -3349 -458 -3303
rect -412 -3349 -362 -3303
rect -316 -3349 -268 -3303
rect -222 -3349 -167 -3303
rect -121 -3349 -73 -3303
rect -27 -3349 21 -3303
rect 67 -3349 115 -3303
rect 161 -3349 216 -3303
rect 262 -3349 310 -3303
rect 356 -3349 406 -3303
rect 452 -3349 500 -3303
rect 546 -3349 601 -3303
rect 647 -3349 695 -3303
rect 741 -3349 789 -3303
rect 835 -3349 883 -3303
rect 929 -3349 984 -3303
rect 1030 -3349 1078 -3303
rect 1124 -3349 1172 -3303
rect 1218 -3349 1244 -3303
rect -773 -3375 1244 -3349
rect 1858 -3478 2058 -2830
rect 2350 -2839 2376 -2830
rect 2422 -2839 2448 -2793
rect 2350 -2861 2448 -2839
rect 2524 963 2585 1083
rect 2684 963 2745 1083
rect 2524 952 2745 963
rect 2524 901 2610 952
rect 2661 901 2745 952
rect 2524 889 2745 901
rect 2524 218 2585 889
rect 2684 218 2745 889
rect 2847 661 2903 848
rect 2826 643 2923 661
rect 2826 579 2843 643
rect 2907 579 2923 643
rect 2826 527 2923 579
rect 2826 463 2843 527
rect 2907 463 2923 527
rect 2826 449 2923 463
rect 2524 207 2745 218
rect 2524 156 2610 207
rect 2661 156 2745 207
rect 2524 144 2745 156
rect 2524 -518 2585 144
rect 2684 -518 2745 144
rect 2847 -79 2903 449
rect 2826 -97 2923 -79
rect 2826 -161 2843 -97
rect 2907 -161 2923 -97
rect 2826 -213 2923 -161
rect 2826 -277 2843 -213
rect 2907 -277 2923 -213
rect 2826 -291 2923 -277
rect 2524 -529 2745 -518
rect 2524 -580 2610 -529
rect 2661 -580 2745 -529
rect 2524 -592 2745 -580
rect 2524 -1255 2585 -592
rect 2684 -1255 2745 -592
rect 2847 -842 2903 -291
rect 2826 -860 2923 -842
rect 2826 -924 2843 -860
rect 2907 -924 2923 -860
rect 2826 -976 2923 -924
rect 2826 -1040 2843 -976
rect 2907 -1040 2923 -976
rect 2826 -1054 2923 -1040
rect 2524 -1266 2745 -1255
rect 2524 -1317 2610 -1266
rect 2661 -1317 2745 -1266
rect 2524 -1329 2745 -1317
rect 2524 -1991 2585 -1329
rect 2684 -1991 2745 -1329
rect 2847 -1571 2903 -1054
rect 2826 -1589 2923 -1571
rect 2826 -1653 2843 -1589
rect 2907 -1653 2923 -1589
rect 2826 -1705 2923 -1653
rect 2826 -1769 2843 -1705
rect 2907 -1769 2923 -1705
rect 2826 -1783 2923 -1769
rect 2524 -2002 2745 -1991
rect 2524 -2053 2610 -2002
rect 2661 -2053 2745 -2002
rect 2524 -2065 2745 -2053
rect 2524 -2861 2585 -2065
rect 2684 -2861 2745 -2065
rect 2847 -2289 2903 -1783
rect 2826 -2307 2923 -2289
rect 2826 -2371 2843 -2307
rect 2907 -2371 2923 -2307
rect 2826 -2423 2923 -2371
rect 2826 -2487 2843 -2423
rect 2907 -2487 2923 -2423
rect 2826 -2501 2923 -2487
rect 2847 -2694 2903 -2501
rect 3004 -2861 3065 1083
rect 3167 659 3223 848
rect 3146 641 3243 659
rect 3146 577 3163 641
rect 3227 577 3243 641
rect 3146 525 3243 577
rect 3146 461 3163 525
rect 3227 461 3243 525
rect 3146 447 3243 461
rect 3167 -81 3223 447
rect 3146 -99 3243 -81
rect 3146 -163 3163 -99
rect 3227 -163 3243 -99
rect 3146 -215 3243 -163
rect 3146 -279 3163 -215
rect 3227 -279 3243 -215
rect 3146 -293 3243 -279
rect 3167 -810 3223 -293
rect 3146 -828 3243 -810
rect 3146 -892 3163 -828
rect 3227 -892 3243 -828
rect 3146 -944 3243 -892
rect 3146 -1008 3163 -944
rect 3227 -1008 3243 -944
rect 3146 -1022 3243 -1008
rect 3167 -1550 3223 -1022
rect 3146 -1568 3243 -1550
rect 3146 -1632 3163 -1568
rect 3227 -1632 3243 -1568
rect 3146 -1684 3243 -1632
rect 3146 -1748 3163 -1684
rect 3227 -1748 3243 -1684
rect 3146 -1762 3243 -1748
rect 3167 -2290 3223 -1762
rect 3146 -2308 3243 -2290
rect 3146 -2372 3163 -2308
rect 3227 -2372 3243 -2308
rect 3146 -2424 3243 -2372
rect 3146 -2488 3163 -2424
rect 3227 -2488 3243 -2424
rect 3146 -2502 3243 -2488
rect 3167 -2694 3223 -2502
rect 3324 -2861 3385 1083
rect 3472 942 3557 955
rect 3472 892 3488 942
rect 3538 892 3557 942
rect 3472 877 3557 892
rect 3484 689 3545 877
rect 3466 671 3563 689
rect 3466 607 3483 671
rect 3547 607 3563 671
rect 3466 555 3563 607
rect 3466 491 3483 555
rect 3547 491 3563 555
rect 3466 477 3563 491
rect 3484 220 3545 477
rect 3473 207 3558 220
rect 3473 157 3489 207
rect 3539 157 3558 207
rect 3473 142 3558 157
rect 3484 -62 3545 142
rect 3466 -80 3563 -62
rect 3466 -144 3483 -80
rect 3547 -144 3563 -80
rect 3466 -196 3563 -144
rect 3466 -260 3483 -196
rect 3547 -260 3563 -196
rect 3466 -274 3563 -260
rect 3484 -516 3545 -274
rect 3471 -529 3556 -516
rect 3471 -579 3487 -529
rect 3537 -579 3556 -529
rect 3471 -594 3556 -579
rect 3484 -794 3545 -594
rect 3466 -812 3563 -794
rect 3466 -876 3483 -812
rect 3547 -876 3563 -812
rect 3466 -928 3563 -876
rect 3466 -992 3483 -928
rect 3547 -992 3563 -928
rect 3466 -1006 3563 -992
rect 3484 -1252 3545 -1006
rect 3471 -1265 3556 -1252
rect 3471 -1315 3487 -1265
rect 3537 -1315 3556 -1265
rect 3471 -1330 3556 -1315
rect 3484 -1536 3545 -1330
rect 3466 -1554 3563 -1536
rect 3466 -1618 3483 -1554
rect 3547 -1618 3563 -1554
rect 3466 -1670 3563 -1618
rect 3466 -1734 3483 -1670
rect 3547 -1734 3563 -1670
rect 3466 -1748 3563 -1734
rect 3484 -1986 3545 -1748
rect 3472 -1999 3557 -1986
rect 3472 -2049 3488 -1999
rect 3538 -2049 3557 -1999
rect 3472 -2064 3557 -2049
rect 3484 -2296 3545 -2064
rect 3466 -2314 3563 -2296
rect 3466 -2378 3483 -2314
rect 3547 -2378 3563 -2314
rect 3466 -2430 3563 -2378
rect 3466 -2494 3483 -2430
rect 3547 -2494 3563 -2430
rect 3466 -2508 3563 -2494
rect 3484 -2721 3545 -2508
rect 3470 -2734 3555 -2721
rect 3470 -2784 3486 -2734
rect 3536 -2784 3555 -2734
rect 3470 -2799 3555 -2784
rect 3645 -2861 3706 1083
rect 3807 676 3863 847
rect 3786 658 3883 676
rect 3786 594 3803 658
rect 3867 594 3883 658
rect 3786 542 3883 594
rect 3786 478 3803 542
rect 3867 478 3883 542
rect 3786 464 3883 478
rect 3807 -83 3863 464
rect 3786 -101 3883 -83
rect 3786 -165 3803 -101
rect 3867 -165 3883 -101
rect 3786 -217 3883 -165
rect 3786 -281 3803 -217
rect 3867 -281 3883 -217
rect 3786 -295 3883 -281
rect 3807 -819 3863 -295
rect 3786 -837 3883 -819
rect 3786 -901 3803 -837
rect 3867 -901 3883 -837
rect 3786 -953 3883 -901
rect 3786 -1017 3803 -953
rect 3867 -1017 3883 -953
rect 3786 -1031 3883 -1017
rect 3807 -1544 3863 -1031
rect 3786 -1562 3883 -1544
rect 3786 -1626 3803 -1562
rect 3867 -1626 3883 -1562
rect 3786 -1678 3883 -1626
rect 3786 -1742 3803 -1678
rect 3867 -1742 3883 -1678
rect 3786 -1756 3883 -1742
rect 3807 -2292 3863 -1756
rect 3786 -2310 3883 -2292
rect 3786 -2374 3803 -2310
rect 3867 -2374 3883 -2310
rect 3786 -2426 3883 -2374
rect 3786 -2490 3803 -2426
rect 3867 -2490 3883 -2426
rect 3786 -2504 3883 -2490
rect 3807 -2695 3863 -2504
rect 3965 -2861 4026 1083
rect 4284 963 4345 1083
rect 4443 963 4504 1083
rect 4284 952 4504 963
rect 4284 901 4370 952
rect 4421 901 4504 952
rect 4284 889 4504 901
rect 4127 673 4183 847
rect 4106 655 4203 673
rect 4106 591 4123 655
rect 4187 591 4203 655
rect 4106 539 4203 591
rect 4106 475 4123 539
rect 4187 475 4203 539
rect 4106 461 4203 475
rect 4127 -98 4183 461
rect 4284 218 4345 889
rect 4443 218 4504 889
rect 4284 207 4504 218
rect 4284 156 4370 207
rect 4421 156 4504 207
rect 4284 144 4504 156
rect 4106 -116 4203 -98
rect 4106 -180 4123 -116
rect 4187 -180 4203 -116
rect 4106 -232 4203 -180
rect 4106 -296 4123 -232
rect 4187 -296 4203 -232
rect 4106 -310 4203 -296
rect 4127 -823 4183 -310
rect 4284 -518 4345 144
rect 4443 -518 4504 144
rect 4284 -529 4504 -518
rect 4284 -580 4370 -529
rect 4421 -580 4504 -529
rect 4284 -592 4504 -580
rect 4106 -841 4203 -823
rect 4106 -905 4123 -841
rect 4187 -905 4203 -841
rect 4106 -957 4203 -905
rect 4106 -1021 4123 -957
rect 4187 -1021 4203 -957
rect 4106 -1035 4203 -1021
rect 4127 -1547 4183 -1035
rect 4284 -1255 4345 -592
rect 4443 -1255 4504 -592
rect 4284 -1266 4504 -1255
rect 4284 -1317 4370 -1266
rect 4421 -1317 4504 -1266
rect 4284 -1329 4504 -1317
rect 4106 -1565 4203 -1547
rect 4106 -1629 4123 -1565
rect 4187 -1629 4203 -1565
rect 4106 -1681 4203 -1629
rect 4106 -1745 4123 -1681
rect 4187 -1745 4203 -1681
rect 4106 -1759 4203 -1745
rect 4127 -2295 4183 -1759
rect 4284 -1991 4345 -1329
rect 4443 -1991 4504 -1329
rect 4284 -2002 4504 -1991
rect 4284 -2053 4370 -2002
rect 4421 -2053 4504 -2002
rect 4284 -2065 4504 -2053
rect 4106 -2313 4203 -2295
rect 4106 -2377 4123 -2313
rect 4187 -2377 4203 -2313
rect 4106 -2429 4203 -2377
rect 4106 -2493 4123 -2429
rect 4187 -2493 4203 -2429
rect 4106 -2507 4203 -2493
rect 4127 -2695 4183 -2507
rect 4284 -2861 4345 -2065
rect 4443 -2861 4504 -2065
rect 4608 1061 4706 1083
rect 4608 1015 4634 1061
rect 4680 1015 4706 1061
rect 4608 967 4706 1015
rect 4608 921 4634 967
rect 4680 963 4706 967
rect 4826 963 5022 1173
rect 5150 1155 7506 1173
rect 5150 1109 5177 1155
rect 5223 1109 5271 1155
rect 5317 1109 5365 1155
rect 5411 1109 5459 1155
rect 5505 1109 5553 1155
rect 5599 1109 5647 1155
rect 5693 1109 5741 1155
rect 5787 1109 5835 1155
rect 5881 1109 5929 1155
rect 5975 1109 6023 1155
rect 6069 1109 6117 1155
rect 6163 1109 6211 1155
rect 6257 1109 6305 1155
rect 6351 1109 6399 1155
rect 6445 1109 6493 1155
rect 6539 1109 6587 1155
rect 6633 1109 6681 1155
rect 6727 1109 6775 1155
rect 6821 1109 6869 1155
rect 6915 1109 6963 1155
rect 7009 1109 7057 1155
rect 7103 1109 7151 1155
rect 7197 1109 7245 1155
rect 7291 1109 7339 1155
rect 7385 1109 7433 1155
rect 7479 1109 7506 1155
rect 5150 1083 7506 1109
rect 5150 1061 5248 1083
rect 5150 1015 5176 1061
rect 5222 1015 5248 1061
rect 5150 967 5248 1015
rect 5150 963 5176 967
rect 4680 921 5176 963
rect 5222 921 5248 967
rect 4608 873 5248 921
rect 4608 827 4634 873
rect 4680 827 5176 873
rect 5222 827 5248 873
rect 4608 779 5248 827
rect 4608 733 4634 779
rect 4680 763 5176 779
rect 4680 733 4706 763
rect 4608 685 4706 733
rect 4608 639 4634 685
rect 4680 639 4706 685
rect 4608 591 4706 639
rect 4608 545 4634 591
rect 4680 563 4706 591
rect 4826 563 5022 763
rect 5150 733 5176 763
rect 5222 733 5248 779
rect 5150 685 5248 733
rect 5150 639 5176 685
rect 5222 639 5248 685
rect 5150 591 5248 639
rect 5150 563 5176 591
rect 4680 545 5176 563
rect 5222 545 5248 591
rect 4608 497 5248 545
rect 4608 451 4634 497
rect 4680 451 5176 497
rect 5222 451 5248 497
rect 4608 403 5248 451
rect 4608 357 4634 403
rect 4680 363 5176 403
rect 4680 357 4706 363
rect 4608 309 4706 357
rect 4608 263 4634 309
rect 4680 263 4706 309
rect 4608 215 4706 263
rect 4608 169 4634 215
rect 4680 169 4706 215
rect 4608 163 4706 169
rect 4826 163 5022 363
rect 5150 357 5176 363
rect 5222 357 5248 403
rect 5150 309 5248 357
rect 5150 263 5176 309
rect 5222 263 5248 309
rect 5150 215 5248 263
rect 5150 169 5176 215
rect 5222 169 5248 215
rect 5150 163 5248 169
rect 4608 121 5248 163
rect 4608 75 4634 121
rect 4680 75 5176 121
rect 5222 75 5248 121
rect 4608 27 5248 75
rect 4608 -19 4634 27
rect 4680 -19 5176 27
rect 5222 -19 5248 27
rect 4608 -37 5248 -19
rect 4608 -67 4706 -37
rect 4608 -113 4634 -67
rect 4680 -113 4706 -67
rect 4608 -161 4706 -113
rect 4608 -207 4634 -161
rect 4680 -207 4706 -161
rect 4608 -237 4706 -207
rect 4826 -237 5022 -37
rect 5150 -67 5248 -37
rect 5150 -113 5176 -67
rect 5222 -113 5248 -67
rect 5150 -161 5248 -113
rect 5150 -207 5176 -161
rect 5222 -207 5248 -161
rect 5150 -237 5248 -207
rect 4608 -255 5248 -237
rect 4608 -301 4634 -255
rect 4680 -301 5176 -255
rect 5222 -301 5248 -255
rect 4608 -349 5248 -301
rect 4608 -395 4634 -349
rect 4680 -395 5176 -349
rect 5222 -395 5248 -349
rect 4608 -437 5248 -395
rect 4608 -443 4706 -437
rect 4608 -489 4634 -443
rect 4680 -489 4706 -443
rect 4608 -537 4706 -489
rect 4608 -583 4634 -537
rect 4680 -583 4706 -537
rect 4608 -631 4706 -583
rect 4608 -677 4634 -631
rect 4680 -637 4706 -631
rect 4826 -637 5022 -437
rect 5150 -443 5248 -437
rect 5150 -489 5176 -443
rect 5222 -489 5248 -443
rect 5150 -537 5248 -489
rect 5150 -583 5176 -537
rect 5222 -583 5248 -537
rect 5150 -631 5248 -583
rect 5150 -637 5176 -631
rect 4680 -677 5176 -637
rect 5222 -677 5248 -631
rect 4608 -725 5248 -677
rect 4608 -771 4634 -725
rect 4680 -771 5176 -725
rect 5222 -771 5248 -725
rect 4608 -819 5248 -771
rect 4608 -865 4634 -819
rect 4680 -837 5176 -819
rect 4680 -865 4706 -837
rect 4608 -913 4706 -865
rect 4608 -959 4634 -913
rect 4680 -959 4706 -913
rect 4608 -1007 4706 -959
rect 4608 -1053 4634 -1007
rect 4680 -1037 4706 -1007
rect 4826 -1037 5022 -837
rect 5150 -865 5176 -837
rect 5222 -865 5248 -819
rect 5150 -913 5248 -865
rect 5150 -959 5176 -913
rect 5222 -959 5248 -913
rect 5150 -1007 5248 -959
rect 5150 -1037 5176 -1007
rect 4680 -1053 5176 -1037
rect 5222 -1053 5248 -1007
rect 4608 -1101 5248 -1053
rect 4608 -1147 4634 -1101
rect 4680 -1147 5176 -1101
rect 5222 -1147 5248 -1101
rect 4608 -1195 5248 -1147
rect 4608 -1241 4634 -1195
rect 4680 -1237 5176 -1195
rect 4680 -1241 4706 -1237
rect 4608 -1289 4706 -1241
rect 4608 -1335 4634 -1289
rect 4680 -1335 4706 -1289
rect 4608 -1383 4706 -1335
rect 4608 -1429 4634 -1383
rect 4680 -1429 4706 -1383
rect 4608 -1437 4706 -1429
rect 4826 -1437 5022 -1237
rect 5150 -1241 5176 -1237
rect 5222 -1241 5248 -1195
rect 5150 -1289 5248 -1241
rect 5150 -1335 5176 -1289
rect 5222 -1335 5248 -1289
rect 5150 -1383 5248 -1335
rect 5150 -1429 5176 -1383
rect 5222 -1429 5248 -1383
rect 5150 -1437 5248 -1429
rect 4608 -1477 5248 -1437
rect 4608 -1523 4634 -1477
rect 4680 -1523 5176 -1477
rect 5222 -1523 5248 -1477
rect 4608 -1571 5248 -1523
rect 4608 -1617 4634 -1571
rect 4680 -1617 5176 -1571
rect 5222 -1617 5248 -1571
rect 4608 -1637 5248 -1617
rect 4608 -1665 4706 -1637
rect 4608 -1711 4634 -1665
rect 4680 -1711 4706 -1665
rect 4608 -1759 4706 -1711
rect 4608 -1805 4634 -1759
rect 4680 -1805 4706 -1759
rect 4608 -1837 4706 -1805
rect 4826 -1837 5022 -1637
rect 5150 -1665 5248 -1637
rect 5150 -1711 5176 -1665
rect 5222 -1711 5248 -1665
rect 5150 -1759 5248 -1711
rect 5150 -1805 5176 -1759
rect 5222 -1805 5248 -1759
rect 5150 -1837 5248 -1805
rect 4608 -1853 5248 -1837
rect 4608 -1899 4634 -1853
rect 4680 -1899 5176 -1853
rect 5222 -1899 5248 -1853
rect 4608 -1947 5248 -1899
rect 4608 -1993 4634 -1947
rect 4680 -1993 5176 -1947
rect 5222 -1993 5248 -1947
rect 4608 -2037 5248 -1993
rect 4608 -2041 4706 -2037
rect 4608 -2087 4634 -2041
rect 4680 -2087 4706 -2041
rect 4608 -2135 4706 -2087
rect 4608 -2181 4634 -2135
rect 4680 -2181 4706 -2135
rect 4608 -2229 4706 -2181
rect 4608 -2275 4634 -2229
rect 4680 -2237 4706 -2229
rect 4826 -2237 5022 -2037
rect 5150 -2041 5248 -2037
rect 5150 -2087 5176 -2041
rect 5222 -2087 5248 -2041
rect 5150 -2135 5248 -2087
rect 5150 -2181 5176 -2135
rect 5222 -2181 5248 -2135
rect 5150 -2229 5248 -2181
rect 5150 -2237 5176 -2229
rect 4680 -2275 5176 -2237
rect 5222 -2275 5248 -2229
rect 4608 -2323 5248 -2275
rect 4608 -2369 4634 -2323
rect 4680 -2369 5176 -2323
rect 5222 -2369 5248 -2323
rect 4608 -2417 5248 -2369
rect 4608 -2463 4634 -2417
rect 4680 -2437 5176 -2417
rect 4680 -2463 4706 -2437
rect 4608 -2511 4706 -2463
rect 4608 -2557 4634 -2511
rect 4680 -2557 4706 -2511
rect 4608 -2605 4706 -2557
rect 4608 -2651 4634 -2605
rect 4680 -2637 4706 -2605
rect 4826 -2637 5022 -2437
rect 5150 -2463 5176 -2437
rect 5222 -2463 5248 -2417
rect 5150 -2511 5248 -2463
rect 5150 -2557 5176 -2511
rect 5222 -2557 5248 -2511
rect 5150 -2605 5248 -2557
rect 5150 -2637 5176 -2605
rect 4680 -2651 5176 -2637
rect 5222 -2651 5248 -2605
rect 4608 -2699 5248 -2651
rect 4608 -2745 4634 -2699
rect 4680 -2745 5176 -2699
rect 5222 -2745 5248 -2699
rect 4608 -2793 5248 -2745
rect 4608 -2839 4634 -2793
rect 4680 -2837 5176 -2793
rect 4680 -2839 4706 -2837
rect 4608 -2861 4706 -2839
rect 2350 -2887 4706 -2861
rect 2350 -2933 2377 -2887
rect 2423 -2933 2471 -2887
rect 2517 -2933 2565 -2887
rect 2611 -2933 2659 -2887
rect 2705 -2933 2753 -2887
rect 2799 -2933 2847 -2887
rect 2893 -2933 2941 -2887
rect 2987 -2933 3035 -2887
rect 3081 -2933 3129 -2887
rect 3175 -2933 3223 -2887
rect 3269 -2933 3317 -2887
rect 3363 -2933 3411 -2887
rect 3457 -2933 3505 -2887
rect 3551 -2933 3599 -2887
rect 3645 -2933 3693 -2887
rect 3739 -2933 3787 -2887
rect 3833 -2933 3881 -2887
rect 3927 -2933 3975 -2887
rect 4021 -2933 4069 -2887
rect 4115 -2933 4163 -2887
rect 4209 -2933 4257 -2887
rect 4303 -2933 4351 -2887
rect 4397 -2933 4445 -2887
rect 4491 -2933 4539 -2887
rect 4585 -2933 4633 -2887
rect 4679 -2933 4706 -2887
rect 2350 -2959 4706 -2933
rect 2403 -3478 2603 -2959
rect 2803 -3478 3003 -2959
rect 3203 -3478 3403 -2959
rect 3603 -3478 3803 -2959
rect 4003 -3478 4203 -2959
rect 4403 -3478 4603 -2959
rect 4826 -3478 5022 -2837
rect 5150 -2839 5176 -2837
rect 5222 -2839 5248 -2793
rect 5150 -2861 5248 -2839
rect 5324 963 5385 1083
rect 5484 963 5545 1083
rect 5324 952 5545 963
rect 5324 901 5410 952
rect 5461 901 5545 952
rect 5324 889 5545 901
rect 5324 218 5385 889
rect 5484 218 5545 889
rect 5647 661 5703 848
rect 5626 643 5723 661
rect 5626 579 5643 643
rect 5707 579 5723 643
rect 5626 527 5723 579
rect 5626 463 5643 527
rect 5707 463 5723 527
rect 5626 449 5723 463
rect 5324 207 5545 218
rect 5324 156 5410 207
rect 5461 156 5545 207
rect 5324 144 5545 156
rect 5324 -518 5385 144
rect 5484 -518 5545 144
rect 5647 -79 5703 449
rect 5626 -97 5723 -79
rect 5626 -161 5643 -97
rect 5707 -161 5723 -97
rect 5626 -213 5723 -161
rect 5626 -277 5643 -213
rect 5707 -277 5723 -213
rect 5626 -291 5723 -277
rect 5324 -529 5545 -518
rect 5324 -580 5410 -529
rect 5461 -580 5545 -529
rect 5324 -592 5545 -580
rect 5324 -1255 5385 -592
rect 5484 -1255 5545 -592
rect 5647 -842 5703 -291
rect 5626 -860 5723 -842
rect 5626 -924 5643 -860
rect 5707 -924 5723 -860
rect 5626 -976 5723 -924
rect 5626 -1040 5643 -976
rect 5707 -1040 5723 -976
rect 5626 -1054 5723 -1040
rect 5324 -1266 5545 -1255
rect 5324 -1317 5410 -1266
rect 5461 -1317 5545 -1266
rect 5324 -1329 5545 -1317
rect 5324 -1991 5385 -1329
rect 5484 -1991 5545 -1329
rect 5647 -1571 5703 -1054
rect 5626 -1589 5723 -1571
rect 5626 -1653 5643 -1589
rect 5707 -1653 5723 -1589
rect 5626 -1705 5723 -1653
rect 5626 -1769 5643 -1705
rect 5707 -1769 5723 -1705
rect 5626 -1783 5723 -1769
rect 5324 -2002 5545 -1991
rect 5324 -2053 5410 -2002
rect 5461 -2053 5545 -2002
rect 5324 -2065 5545 -2053
rect 5324 -2861 5385 -2065
rect 5484 -2861 5545 -2065
rect 5647 -2289 5703 -1783
rect 5626 -2307 5723 -2289
rect 5626 -2371 5643 -2307
rect 5707 -2371 5723 -2307
rect 5626 -2423 5723 -2371
rect 5626 -2487 5643 -2423
rect 5707 -2487 5723 -2423
rect 5626 -2501 5723 -2487
rect 5647 -2694 5703 -2501
rect 5804 -2861 5865 1083
rect 5967 659 6023 848
rect 5946 641 6043 659
rect 5946 577 5963 641
rect 6027 577 6043 641
rect 5946 525 6043 577
rect 5946 461 5963 525
rect 6027 461 6043 525
rect 5946 447 6043 461
rect 5967 -81 6023 447
rect 5946 -99 6043 -81
rect 5946 -163 5963 -99
rect 6027 -163 6043 -99
rect 5946 -215 6043 -163
rect 5946 -279 5963 -215
rect 6027 -279 6043 -215
rect 5946 -293 6043 -279
rect 5967 -810 6023 -293
rect 5946 -828 6043 -810
rect 5946 -892 5963 -828
rect 6027 -892 6043 -828
rect 5946 -944 6043 -892
rect 5946 -1008 5963 -944
rect 6027 -1008 6043 -944
rect 5946 -1022 6043 -1008
rect 5967 -1550 6023 -1022
rect 5946 -1568 6043 -1550
rect 5946 -1632 5963 -1568
rect 6027 -1632 6043 -1568
rect 5946 -1684 6043 -1632
rect 5946 -1748 5963 -1684
rect 6027 -1748 6043 -1684
rect 5946 -1762 6043 -1748
rect 5967 -2290 6023 -1762
rect 5946 -2308 6043 -2290
rect 5946 -2372 5963 -2308
rect 6027 -2372 6043 -2308
rect 5946 -2424 6043 -2372
rect 5946 -2488 5963 -2424
rect 6027 -2488 6043 -2424
rect 5946 -2502 6043 -2488
rect 5967 -2694 6023 -2502
rect 6124 -2861 6185 1083
rect 6272 942 6357 955
rect 6272 892 6288 942
rect 6338 892 6357 942
rect 6272 877 6357 892
rect 6284 689 6345 877
rect 6266 671 6363 689
rect 6266 607 6283 671
rect 6347 607 6363 671
rect 6266 555 6363 607
rect 6266 491 6283 555
rect 6347 491 6363 555
rect 6266 477 6363 491
rect 6284 220 6345 477
rect 6273 207 6358 220
rect 6273 157 6289 207
rect 6339 157 6358 207
rect 6273 142 6358 157
rect 6284 -62 6345 142
rect 6266 -80 6363 -62
rect 6266 -144 6283 -80
rect 6347 -144 6363 -80
rect 6266 -196 6363 -144
rect 6266 -260 6283 -196
rect 6347 -260 6363 -196
rect 6266 -274 6363 -260
rect 6284 -516 6345 -274
rect 6271 -529 6356 -516
rect 6271 -579 6287 -529
rect 6337 -579 6356 -529
rect 6271 -594 6356 -579
rect 6284 -794 6345 -594
rect 6266 -812 6363 -794
rect 6266 -876 6283 -812
rect 6347 -876 6363 -812
rect 6266 -928 6363 -876
rect 6266 -992 6283 -928
rect 6347 -992 6363 -928
rect 6266 -1006 6363 -992
rect 6284 -1252 6345 -1006
rect 6271 -1265 6356 -1252
rect 6271 -1315 6287 -1265
rect 6337 -1315 6356 -1265
rect 6271 -1330 6356 -1315
rect 6284 -1536 6345 -1330
rect 6266 -1554 6363 -1536
rect 6266 -1618 6283 -1554
rect 6347 -1618 6363 -1554
rect 6266 -1670 6363 -1618
rect 6266 -1734 6283 -1670
rect 6347 -1734 6363 -1670
rect 6266 -1748 6363 -1734
rect 6284 -1986 6345 -1748
rect 6272 -1999 6357 -1986
rect 6272 -2049 6288 -1999
rect 6338 -2049 6357 -1999
rect 6272 -2064 6357 -2049
rect 6284 -2296 6345 -2064
rect 6266 -2314 6363 -2296
rect 6266 -2378 6283 -2314
rect 6347 -2378 6363 -2314
rect 6266 -2430 6363 -2378
rect 6266 -2494 6283 -2430
rect 6347 -2494 6363 -2430
rect 6266 -2508 6363 -2494
rect 6284 -2721 6345 -2508
rect 6270 -2734 6355 -2721
rect 6270 -2784 6286 -2734
rect 6336 -2784 6355 -2734
rect 6270 -2799 6355 -2784
rect 6445 -2861 6506 1083
rect 6607 676 6663 847
rect 6586 658 6683 676
rect 6586 594 6603 658
rect 6667 594 6683 658
rect 6586 542 6683 594
rect 6586 478 6603 542
rect 6667 478 6683 542
rect 6586 464 6683 478
rect 6607 -83 6663 464
rect 6586 -101 6683 -83
rect 6586 -165 6603 -101
rect 6667 -165 6683 -101
rect 6586 -217 6683 -165
rect 6586 -281 6603 -217
rect 6667 -281 6683 -217
rect 6586 -295 6683 -281
rect 6607 -819 6663 -295
rect 6586 -837 6683 -819
rect 6586 -901 6603 -837
rect 6667 -901 6683 -837
rect 6586 -953 6683 -901
rect 6586 -1017 6603 -953
rect 6667 -1017 6683 -953
rect 6586 -1031 6683 -1017
rect 6607 -1544 6663 -1031
rect 6586 -1562 6683 -1544
rect 6586 -1626 6603 -1562
rect 6667 -1626 6683 -1562
rect 6586 -1678 6683 -1626
rect 6586 -1742 6603 -1678
rect 6667 -1742 6683 -1678
rect 6586 -1756 6683 -1742
rect 6607 -2292 6663 -1756
rect 6586 -2310 6683 -2292
rect 6586 -2374 6603 -2310
rect 6667 -2374 6683 -2310
rect 6586 -2426 6683 -2374
rect 6586 -2490 6603 -2426
rect 6667 -2490 6683 -2426
rect 6586 -2504 6683 -2490
rect 6607 -2695 6663 -2504
rect 6765 -2861 6826 1083
rect 7084 963 7145 1083
rect 7243 963 7304 1083
rect 7084 952 7304 963
rect 7084 901 7170 952
rect 7221 901 7304 952
rect 7084 889 7304 901
rect 6927 673 6983 847
rect 6906 655 7003 673
rect 6906 591 6923 655
rect 6987 591 7003 655
rect 6906 539 7003 591
rect 6906 475 6923 539
rect 6987 475 7003 539
rect 6906 461 7003 475
rect 6927 -98 6983 461
rect 7084 218 7145 889
rect 7243 218 7304 889
rect 7084 207 7304 218
rect 7084 156 7170 207
rect 7221 156 7304 207
rect 7084 144 7304 156
rect 6906 -116 7003 -98
rect 6906 -180 6923 -116
rect 6987 -180 7003 -116
rect 6906 -232 7003 -180
rect 6906 -296 6923 -232
rect 6987 -296 7003 -232
rect 6906 -310 7003 -296
rect 6927 -823 6983 -310
rect 7084 -518 7145 144
rect 7243 -518 7304 144
rect 7084 -529 7304 -518
rect 7084 -580 7170 -529
rect 7221 -580 7304 -529
rect 7084 -592 7304 -580
rect 6906 -841 7003 -823
rect 6906 -905 6923 -841
rect 6987 -905 7003 -841
rect 6906 -957 7003 -905
rect 6906 -1021 6923 -957
rect 6987 -1021 7003 -957
rect 6906 -1035 7003 -1021
rect 6927 -1547 6983 -1035
rect 7084 -1255 7145 -592
rect 7243 -1255 7304 -592
rect 7084 -1266 7304 -1255
rect 7084 -1317 7170 -1266
rect 7221 -1317 7304 -1266
rect 7084 -1329 7304 -1317
rect 6906 -1565 7003 -1547
rect 6906 -1629 6923 -1565
rect 6987 -1629 7003 -1565
rect 6906 -1681 7003 -1629
rect 6906 -1745 6923 -1681
rect 6987 -1745 7003 -1681
rect 6906 -1759 7003 -1745
rect 6927 -2295 6983 -1759
rect 7084 -1991 7145 -1329
rect 7243 -1991 7304 -1329
rect 7084 -2002 7304 -1991
rect 7084 -2053 7170 -2002
rect 7221 -2053 7304 -2002
rect 7084 -2065 7304 -2053
rect 6906 -2313 7003 -2295
rect 6906 -2377 6923 -2313
rect 6987 -2377 7003 -2313
rect 6906 -2429 7003 -2377
rect 6906 -2493 6923 -2429
rect 6987 -2493 7003 -2429
rect 6906 -2507 7003 -2493
rect 6927 -2695 6983 -2507
rect 7084 -2861 7145 -2065
rect 7243 -2861 7304 -2065
rect 7408 1061 7506 1083
rect 7408 1015 7434 1061
rect 7480 1015 7506 1061
rect 7408 967 7506 1015
rect 7408 921 7434 967
rect 7480 966 7506 967
rect 7620 966 7816 1173
rect 7950 1155 12216 1173
rect 7950 1109 7977 1155
rect 8023 1109 8071 1155
rect 8117 1109 8165 1155
rect 8211 1109 8259 1155
rect 8305 1109 8353 1155
rect 8399 1109 8447 1155
rect 8493 1109 8541 1155
rect 8587 1109 8635 1155
rect 8681 1109 8729 1155
rect 8775 1109 8823 1155
rect 8869 1109 8917 1155
rect 8963 1109 9011 1155
rect 9057 1109 9105 1155
rect 9151 1109 9199 1155
rect 9245 1109 9293 1155
rect 9339 1109 9387 1155
rect 9433 1109 9481 1155
rect 9527 1109 9575 1155
rect 9621 1109 9669 1155
rect 9715 1109 9763 1155
rect 9809 1109 9857 1155
rect 9903 1109 9951 1155
rect 9997 1109 10045 1155
rect 10091 1109 10139 1155
rect 10185 1109 10233 1155
rect 10279 1109 10306 1155
rect 7950 1083 10306 1109
rect 7950 1061 8048 1083
rect 7950 1015 7976 1061
rect 8022 1015 8048 1061
rect 7950 967 8048 1015
rect 7950 966 7976 967
rect 7480 921 7976 966
rect 8022 921 8048 967
rect 7408 873 8048 921
rect 7408 827 7434 873
rect 7480 827 7976 873
rect 8022 827 8048 873
rect 7408 779 8048 827
rect 7408 733 7434 779
rect 7480 766 7976 779
rect 7480 733 7506 766
rect 7408 685 7506 733
rect 7408 639 7434 685
rect 7480 639 7506 685
rect 7408 591 7506 639
rect 7408 545 7434 591
rect 7480 566 7506 591
rect 7620 566 7816 766
rect 7950 733 7976 766
rect 8022 733 8048 779
rect 7950 685 8048 733
rect 7950 639 7976 685
rect 8022 639 8048 685
rect 7950 591 8048 639
rect 7950 566 7976 591
rect 7480 545 7976 566
rect 8022 545 8048 591
rect 7408 497 8048 545
rect 7408 451 7434 497
rect 7480 451 7976 497
rect 8022 451 8048 497
rect 7408 403 8048 451
rect 7408 357 7434 403
rect 7480 366 7976 403
rect 7480 357 7506 366
rect 7408 309 7506 357
rect 7408 263 7434 309
rect 7480 263 7506 309
rect 7408 215 7506 263
rect 7408 169 7434 215
rect 7480 169 7506 215
rect 7408 166 7506 169
rect 7620 166 7816 366
rect 7950 357 7976 366
rect 8022 357 8048 403
rect 7950 309 8048 357
rect 7950 263 7976 309
rect 8022 263 8048 309
rect 7950 215 8048 263
rect 7950 169 7976 215
rect 8022 169 8048 215
rect 7950 166 8048 169
rect 7408 121 8048 166
rect 7408 75 7434 121
rect 7480 75 7976 121
rect 8022 75 8048 121
rect 7408 27 8048 75
rect 7408 -19 7434 27
rect 7480 -19 7976 27
rect 8022 -19 8048 27
rect 7408 -34 8048 -19
rect 7408 -67 7506 -34
rect 7408 -113 7434 -67
rect 7480 -113 7506 -67
rect 7408 -161 7506 -113
rect 7408 -207 7434 -161
rect 7480 -207 7506 -161
rect 7408 -234 7506 -207
rect 7620 -234 7816 -34
rect 7950 -67 8048 -34
rect 7950 -113 7976 -67
rect 8022 -113 8048 -67
rect 7950 -161 8048 -113
rect 7950 -207 7976 -161
rect 8022 -207 8048 -161
rect 7950 -234 8048 -207
rect 7408 -255 8048 -234
rect 7408 -301 7434 -255
rect 7480 -301 7976 -255
rect 8022 -301 8048 -255
rect 7408 -349 8048 -301
rect 7408 -395 7434 -349
rect 7480 -395 7976 -349
rect 8022 -395 8048 -349
rect 7408 -434 8048 -395
rect 7408 -443 7506 -434
rect 7408 -489 7434 -443
rect 7480 -489 7506 -443
rect 7408 -537 7506 -489
rect 7408 -583 7434 -537
rect 7480 -583 7506 -537
rect 7408 -631 7506 -583
rect 7408 -677 7434 -631
rect 7480 -634 7506 -631
rect 7620 -634 7816 -434
rect 7950 -443 8048 -434
rect 7950 -489 7976 -443
rect 8022 -489 8048 -443
rect 7950 -537 8048 -489
rect 7950 -583 7976 -537
rect 8022 -583 8048 -537
rect 7950 -631 8048 -583
rect 7950 -634 7976 -631
rect 7480 -677 7976 -634
rect 8022 -677 8048 -631
rect 7408 -725 8048 -677
rect 7408 -771 7434 -725
rect 7480 -771 7976 -725
rect 8022 -771 8048 -725
rect 7408 -819 8048 -771
rect 7408 -865 7434 -819
rect 7480 -834 7976 -819
rect 7480 -865 7506 -834
rect 7408 -913 7506 -865
rect 7408 -959 7434 -913
rect 7480 -959 7506 -913
rect 7408 -1007 7506 -959
rect 7408 -1053 7434 -1007
rect 7480 -1034 7506 -1007
rect 7620 -1034 7816 -834
rect 7950 -865 7976 -834
rect 8022 -865 8048 -819
rect 7950 -913 8048 -865
rect 7950 -959 7976 -913
rect 8022 -959 8048 -913
rect 7950 -1007 8048 -959
rect 7950 -1034 7976 -1007
rect 7480 -1053 7976 -1034
rect 8022 -1053 8048 -1007
rect 7408 -1101 8048 -1053
rect 7408 -1147 7434 -1101
rect 7480 -1147 7976 -1101
rect 8022 -1147 8048 -1101
rect 7408 -1195 8048 -1147
rect 7408 -1241 7434 -1195
rect 7480 -1234 7976 -1195
rect 7480 -1241 7506 -1234
rect 7408 -1289 7506 -1241
rect 7408 -1335 7434 -1289
rect 7480 -1335 7506 -1289
rect 7408 -1383 7506 -1335
rect 7408 -1429 7434 -1383
rect 7480 -1429 7506 -1383
rect 7408 -1434 7506 -1429
rect 7620 -1434 7816 -1234
rect 7950 -1241 7976 -1234
rect 8022 -1241 8048 -1195
rect 7950 -1289 8048 -1241
rect 7950 -1335 7976 -1289
rect 8022 -1335 8048 -1289
rect 7950 -1383 8048 -1335
rect 7950 -1429 7976 -1383
rect 8022 -1429 8048 -1383
rect 7950 -1434 8048 -1429
rect 7408 -1477 8048 -1434
rect 7408 -1523 7434 -1477
rect 7480 -1523 7976 -1477
rect 8022 -1523 8048 -1477
rect 7408 -1571 8048 -1523
rect 7408 -1617 7434 -1571
rect 7480 -1617 7976 -1571
rect 8022 -1617 8048 -1571
rect 7408 -1634 8048 -1617
rect 7408 -1665 7506 -1634
rect 7408 -1711 7434 -1665
rect 7480 -1711 7506 -1665
rect 7408 -1759 7506 -1711
rect 7408 -1805 7434 -1759
rect 7480 -1805 7506 -1759
rect 7408 -1834 7506 -1805
rect 7620 -1834 7816 -1634
rect 7950 -1665 8048 -1634
rect 7950 -1711 7976 -1665
rect 8022 -1711 8048 -1665
rect 7950 -1759 8048 -1711
rect 7950 -1805 7976 -1759
rect 8022 -1805 8048 -1759
rect 7950 -1834 8048 -1805
rect 7408 -1853 8048 -1834
rect 7408 -1899 7434 -1853
rect 7480 -1899 7976 -1853
rect 8022 -1899 8048 -1853
rect 7408 -1947 8048 -1899
rect 7408 -1993 7434 -1947
rect 7480 -1993 7976 -1947
rect 8022 -1993 8048 -1947
rect 7408 -2034 8048 -1993
rect 7408 -2041 7506 -2034
rect 7408 -2087 7434 -2041
rect 7480 -2087 7506 -2041
rect 7408 -2135 7506 -2087
rect 7408 -2181 7434 -2135
rect 7480 -2181 7506 -2135
rect 7408 -2229 7506 -2181
rect 7408 -2275 7434 -2229
rect 7480 -2234 7506 -2229
rect 7620 -2234 7816 -2034
rect 7950 -2041 8048 -2034
rect 7950 -2087 7976 -2041
rect 8022 -2087 8048 -2041
rect 7950 -2135 8048 -2087
rect 7950 -2181 7976 -2135
rect 8022 -2181 8048 -2135
rect 7950 -2229 8048 -2181
rect 7950 -2234 7976 -2229
rect 7480 -2275 7976 -2234
rect 8022 -2275 8048 -2229
rect 7408 -2323 8048 -2275
rect 7408 -2369 7434 -2323
rect 7480 -2369 7976 -2323
rect 8022 -2369 8048 -2323
rect 7408 -2417 8048 -2369
rect 7408 -2463 7434 -2417
rect 7480 -2434 7976 -2417
rect 7480 -2463 7506 -2434
rect 7408 -2511 7506 -2463
rect 7408 -2557 7434 -2511
rect 7480 -2557 7506 -2511
rect 7408 -2605 7506 -2557
rect 7408 -2651 7434 -2605
rect 7480 -2634 7506 -2605
rect 7620 -2634 7816 -2434
rect 7950 -2463 7976 -2434
rect 8022 -2463 8048 -2417
rect 7950 -2511 8048 -2463
rect 7950 -2557 7976 -2511
rect 8022 -2557 8048 -2511
rect 7950 -2605 8048 -2557
rect 7950 -2634 7976 -2605
rect 7480 -2651 7976 -2634
rect 8022 -2651 8048 -2605
rect 7408 -2699 8048 -2651
rect 7408 -2745 7434 -2699
rect 7480 -2745 7976 -2699
rect 8022 -2745 8048 -2699
rect 7408 -2793 8048 -2745
rect 7408 -2839 7434 -2793
rect 7480 -2834 7976 -2793
rect 7480 -2839 7506 -2834
rect 7408 -2861 7506 -2839
rect 5150 -2887 7506 -2861
rect 5150 -2933 5177 -2887
rect 5223 -2933 5271 -2887
rect 5317 -2933 5365 -2887
rect 5411 -2933 5459 -2887
rect 5505 -2933 5553 -2887
rect 5599 -2933 5647 -2887
rect 5693 -2933 5741 -2887
rect 5787 -2933 5835 -2887
rect 5881 -2933 5929 -2887
rect 5975 -2933 6023 -2887
rect 6069 -2933 6117 -2887
rect 6163 -2933 6211 -2887
rect 6257 -2933 6305 -2887
rect 6351 -2933 6399 -2887
rect 6445 -2933 6493 -2887
rect 6539 -2933 6587 -2887
rect 6633 -2933 6681 -2887
rect 6727 -2933 6775 -2887
rect 6821 -2933 6869 -2887
rect 6915 -2933 6963 -2887
rect 7009 -2933 7057 -2887
rect 7103 -2933 7151 -2887
rect 7197 -2933 7245 -2887
rect 7291 -2933 7339 -2887
rect 7385 -2933 7433 -2887
rect 7479 -2933 7506 -2887
rect 5150 -2959 7506 -2933
rect 7950 -2839 7976 -2834
rect 8022 -2839 8048 -2793
rect 7950 -2861 8048 -2839
rect 8124 963 8185 1083
rect 8284 963 8345 1083
rect 8124 952 8345 963
rect 8124 901 8210 952
rect 8261 901 8345 952
rect 8124 889 8345 901
rect 8124 218 8185 889
rect 8284 218 8345 889
rect 8447 661 8503 848
rect 8426 643 8523 661
rect 8426 579 8443 643
rect 8507 579 8523 643
rect 8426 527 8523 579
rect 8426 463 8443 527
rect 8507 463 8523 527
rect 8426 449 8523 463
rect 8124 207 8345 218
rect 8124 156 8210 207
rect 8261 156 8345 207
rect 8124 144 8345 156
rect 8124 -518 8185 144
rect 8284 -518 8345 144
rect 8447 -79 8503 449
rect 8426 -97 8523 -79
rect 8426 -161 8443 -97
rect 8507 -161 8523 -97
rect 8426 -213 8523 -161
rect 8426 -277 8443 -213
rect 8507 -277 8523 -213
rect 8426 -291 8523 -277
rect 8124 -529 8345 -518
rect 8124 -580 8210 -529
rect 8261 -580 8345 -529
rect 8124 -592 8345 -580
rect 8124 -1255 8185 -592
rect 8284 -1255 8345 -592
rect 8447 -842 8503 -291
rect 8426 -860 8523 -842
rect 8426 -924 8443 -860
rect 8507 -924 8523 -860
rect 8426 -976 8523 -924
rect 8426 -1040 8443 -976
rect 8507 -1040 8523 -976
rect 8426 -1054 8523 -1040
rect 8124 -1266 8345 -1255
rect 8124 -1317 8210 -1266
rect 8261 -1317 8345 -1266
rect 8124 -1329 8345 -1317
rect 8124 -1991 8185 -1329
rect 8284 -1991 8345 -1329
rect 8447 -1571 8503 -1054
rect 8426 -1589 8523 -1571
rect 8426 -1653 8443 -1589
rect 8507 -1653 8523 -1589
rect 8426 -1705 8523 -1653
rect 8426 -1769 8443 -1705
rect 8507 -1769 8523 -1705
rect 8426 -1783 8523 -1769
rect 8124 -2002 8345 -1991
rect 8124 -2053 8210 -2002
rect 8261 -2053 8345 -2002
rect 8124 -2065 8345 -2053
rect 8124 -2861 8185 -2065
rect 8284 -2861 8345 -2065
rect 8447 -2289 8503 -1783
rect 8426 -2307 8523 -2289
rect 8426 -2371 8443 -2307
rect 8507 -2371 8523 -2307
rect 8426 -2423 8523 -2371
rect 8426 -2487 8443 -2423
rect 8507 -2487 8523 -2423
rect 8426 -2501 8523 -2487
rect 8447 -2694 8503 -2501
rect 8604 -2861 8665 1083
rect 8767 659 8823 848
rect 8746 641 8843 659
rect 8746 577 8763 641
rect 8827 577 8843 641
rect 8746 525 8843 577
rect 8746 461 8763 525
rect 8827 461 8843 525
rect 8746 447 8843 461
rect 8767 -81 8823 447
rect 8746 -99 8843 -81
rect 8746 -163 8763 -99
rect 8827 -163 8843 -99
rect 8746 -215 8843 -163
rect 8746 -279 8763 -215
rect 8827 -279 8843 -215
rect 8746 -293 8843 -279
rect 8767 -810 8823 -293
rect 8746 -828 8843 -810
rect 8746 -892 8763 -828
rect 8827 -892 8843 -828
rect 8746 -944 8843 -892
rect 8746 -1008 8763 -944
rect 8827 -1008 8843 -944
rect 8746 -1022 8843 -1008
rect 8767 -1550 8823 -1022
rect 8746 -1568 8843 -1550
rect 8746 -1632 8763 -1568
rect 8827 -1632 8843 -1568
rect 8746 -1684 8843 -1632
rect 8746 -1748 8763 -1684
rect 8827 -1748 8843 -1684
rect 8746 -1762 8843 -1748
rect 8767 -2290 8823 -1762
rect 8746 -2308 8843 -2290
rect 8746 -2372 8763 -2308
rect 8827 -2372 8843 -2308
rect 8746 -2424 8843 -2372
rect 8746 -2488 8763 -2424
rect 8827 -2488 8843 -2424
rect 8746 -2502 8843 -2488
rect 8767 -2694 8823 -2502
rect 8924 -2861 8985 1083
rect 9072 942 9157 955
rect 9072 892 9088 942
rect 9138 892 9157 942
rect 9072 877 9157 892
rect 9084 689 9145 877
rect 9066 671 9163 689
rect 9066 607 9083 671
rect 9147 607 9163 671
rect 9066 555 9163 607
rect 9066 491 9083 555
rect 9147 491 9163 555
rect 9066 477 9163 491
rect 9084 220 9145 477
rect 9073 207 9158 220
rect 9073 157 9089 207
rect 9139 157 9158 207
rect 9073 142 9158 157
rect 9084 -62 9145 142
rect 9066 -80 9163 -62
rect 9066 -144 9083 -80
rect 9147 -144 9163 -80
rect 9066 -196 9163 -144
rect 9066 -260 9083 -196
rect 9147 -260 9163 -196
rect 9066 -274 9163 -260
rect 9084 -516 9145 -274
rect 9071 -529 9156 -516
rect 9071 -579 9087 -529
rect 9137 -579 9156 -529
rect 9071 -594 9156 -579
rect 9084 -794 9145 -594
rect 9066 -812 9163 -794
rect 9066 -876 9083 -812
rect 9147 -876 9163 -812
rect 9066 -928 9163 -876
rect 9066 -992 9083 -928
rect 9147 -992 9163 -928
rect 9066 -1006 9163 -992
rect 9084 -1252 9145 -1006
rect 9071 -1265 9156 -1252
rect 9071 -1315 9087 -1265
rect 9137 -1315 9156 -1265
rect 9071 -1330 9156 -1315
rect 9084 -1536 9145 -1330
rect 9066 -1554 9163 -1536
rect 9066 -1618 9083 -1554
rect 9147 -1618 9163 -1554
rect 9066 -1670 9163 -1618
rect 9066 -1734 9083 -1670
rect 9147 -1734 9163 -1670
rect 9066 -1748 9163 -1734
rect 9084 -1986 9145 -1748
rect 9072 -1999 9157 -1986
rect 9072 -2049 9088 -1999
rect 9138 -2049 9157 -1999
rect 9072 -2064 9157 -2049
rect 9084 -2296 9145 -2064
rect 9066 -2314 9163 -2296
rect 9066 -2378 9083 -2314
rect 9147 -2378 9163 -2314
rect 9066 -2430 9163 -2378
rect 9066 -2494 9083 -2430
rect 9147 -2494 9163 -2430
rect 9066 -2508 9163 -2494
rect 9084 -2721 9145 -2508
rect 9070 -2734 9155 -2721
rect 9070 -2784 9086 -2734
rect 9136 -2784 9155 -2734
rect 9070 -2799 9155 -2784
rect 9245 -2861 9306 1083
rect 9407 676 9463 847
rect 9386 658 9483 676
rect 9386 594 9403 658
rect 9467 594 9483 658
rect 9386 542 9483 594
rect 9386 478 9403 542
rect 9467 478 9483 542
rect 9386 464 9483 478
rect 9407 -83 9463 464
rect 9386 -101 9483 -83
rect 9386 -165 9403 -101
rect 9467 -165 9483 -101
rect 9386 -217 9483 -165
rect 9386 -281 9403 -217
rect 9467 -281 9483 -217
rect 9386 -295 9483 -281
rect 9407 -819 9463 -295
rect 9386 -837 9483 -819
rect 9386 -901 9403 -837
rect 9467 -901 9483 -837
rect 9386 -953 9483 -901
rect 9386 -1017 9403 -953
rect 9467 -1017 9483 -953
rect 9386 -1031 9483 -1017
rect 9407 -1544 9463 -1031
rect 9386 -1562 9483 -1544
rect 9386 -1626 9403 -1562
rect 9467 -1626 9483 -1562
rect 9386 -1678 9483 -1626
rect 9386 -1742 9403 -1678
rect 9467 -1742 9483 -1678
rect 9386 -1756 9483 -1742
rect 9407 -2292 9463 -1756
rect 9386 -2310 9483 -2292
rect 9386 -2374 9403 -2310
rect 9467 -2374 9483 -2310
rect 9386 -2426 9483 -2374
rect 9386 -2490 9403 -2426
rect 9467 -2490 9483 -2426
rect 9386 -2504 9483 -2490
rect 9407 -2695 9463 -2504
rect 9565 -2861 9626 1083
rect 9884 963 9945 1083
rect 10043 963 10104 1083
rect 9884 952 10104 963
rect 9884 901 9970 952
rect 10021 901 10104 952
rect 9884 889 10104 901
rect 9727 673 9783 847
rect 9706 655 9803 673
rect 9706 591 9723 655
rect 9787 591 9803 655
rect 9706 539 9803 591
rect 9706 475 9723 539
rect 9787 475 9803 539
rect 9706 461 9803 475
rect 9727 -98 9783 461
rect 9884 218 9945 889
rect 10043 218 10104 889
rect 9884 207 10104 218
rect 9884 156 9970 207
rect 10021 156 10104 207
rect 9884 144 10104 156
rect 9706 -116 9803 -98
rect 9706 -180 9723 -116
rect 9787 -180 9803 -116
rect 9706 -232 9803 -180
rect 9706 -296 9723 -232
rect 9787 -296 9803 -232
rect 9706 -310 9803 -296
rect 9727 -823 9783 -310
rect 9884 -518 9945 144
rect 10043 -518 10104 144
rect 9884 -529 10104 -518
rect 9884 -580 9970 -529
rect 10021 -580 10104 -529
rect 9884 -592 10104 -580
rect 9706 -841 9803 -823
rect 9706 -905 9723 -841
rect 9787 -905 9803 -841
rect 9706 -957 9803 -905
rect 9706 -1021 9723 -957
rect 9787 -1021 9803 -957
rect 9706 -1035 9803 -1021
rect 9727 -1547 9783 -1035
rect 9884 -1255 9945 -592
rect 10043 -1255 10104 -592
rect 9884 -1266 10104 -1255
rect 9884 -1317 9970 -1266
rect 10021 -1317 10104 -1266
rect 9884 -1329 10104 -1317
rect 9706 -1565 9803 -1547
rect 9706 -1629 9723 -1565
rect 9787 -1629 9803 -1565
rect 9706 -1681 9803 -1629
rect 9706 -1745 9723 -1681
rect 9787 -1745 9803 -1681
rect 9706 -1759 9803 -1745
rect 9727 -2295 9783 -1759
rect 9884 -1991 9945 -1329
rect 10043 -1991 10104 -1329
rect 9884 -2002 10104 -1991
rect 9884 -2053 9970 -2002
rect 10021 -2053 10104 -2002
rect 9884 -2065 10104 -2053
rect 9706 -2313 9803 -2295
rect 9706 -2377 9723 -2313
rect 9787 -2377 9803 -2313
rect 9706 -2429 9803 -2377
rect 9706 -2493 9723 -2429
rect 9787 -2493 9803 -2429
rect 9706 -2507 9803 -2493
rect 9727 -2695 9783 -2507
rect 9884 -2861 9945 -2065
rect 10043 -2861 10104 -2065
rect 10208 1061 10306 1083
rect 10208 1015 10234 1061
rect 10280 1015 10306 1061
rect 10208 967 10306 1015
rect 10208 921 10234 967
rect 10280 921 10306 967
rect 10208 873 10306 921
rect 10208 827 10234 873
rect 10280 827 10306 873
rect 10208 779 10306 827
rect 10208 733 10234 779
rect 10280 733 10306 779
rect 10208 685 10306 733
rect 10208 639 10234 685
rect 10280 639 10306 685
rect 10208 591 10306 639
rect 10208 545 10234 591
rect 10280 545 10306 591
rect 10208 520 10306 545
rect 10861 520 11287 1155
rect 11790 520 12216 1155
rect 10208 497 12216 520
rect 10208 451 10234 497
rect 10280 451 12216 497
rect 10208 403 12216 451
rect 10208 357 10234 403
rect 10280 357 12216 403
rect 10208 309 12216 357
rect 10208 263 10234 309
rect 10280 263 12216 309
rect 10208 215 12216 263
rect 10208 169 10234 215
rect 10280 169 12216 215
rect 10208 121 12216 169
rect 10208 75 10234 121
rect 10280 94 12216 121
rect 10280 75 10306 94
rect 10208 27 10306 75
rect 10208 -19 10234 27
rect 10280 -19 10306 27
rect 10208 -67 10306 -19
rect 10208 -113 10234 -67
rect 10280 -113 10306 -67
rect 10208 -161 10306 -113
rect 10208 -207 10234 -161
rect 10280 -207 10306 -161
rect 10208 -255 10306 -207
rect 10208 -301 10234 -255
rect 10280 -273 10306 -255
rect 10861 -273 11287 94
rect 11790 -273 12216 94
rect 10280 -301 12216 -273
rect 10208 -349 12216 -301
rect 10208 -395 10234 -349
rect 10280 -395 12216 -349
rect 10208 -443 12216 -395
rect 10208 -489 10234 -443
rect 10280 -489 12216 -443
rect 10208 -537 12216 -489
rect 10208 -583 10234 -537
rect 10280 -583 12216 -537
rect 10208 -631 12216 -583
rect 10208 -677 10234 -631
rect 10280 -677 12216 -631
rect 10208 -699 12216 -677
rect 10208 -725 10306 -699
rect 10208 -771 10234 -725
rect 10280 -771 10306 -725
rect 10208 -819 10306 -771
rect 10208 -865 10234 -819
rect 10280 -865 10306 -819
rect 10208 -913 10306 -865
rect 10208 -959 10234 -913
rect 10280 -959 10306 -913
rect 10208 -1007 10306 -959
rect 10208 -1053 10234 -1007
rect 10280 -1053 10306 -1007
rect 10208 -1101 10306 -1053
rect 10208 -1147 10234 -1101
rect 10280 -1147 10306 -1101
rect 10861 -1137 11287 -699
rect 11790 -1145 12216 -699
rect 10208 -1195 10306 -1147
rect 10208 -1241 10234 -1195
rect 10280 -1241 10306 -1195
rect 10208 -1289 10306 -1241
rect 10208 -1335 10234 -1289
rect 10280 -1335 10306 -1289
rect 10755 -1328 10922 -1146
rect 11070 -1254 11746 -1239
rect 11070 -1257 11088 -1254
rect 10993 -1329 11088 -1257
rect 10208 -1383 10306 -1335
rect 11070 -1335 11088 -1329
rect 11169 -1335 11228 -1254
rect 11309 -1335 11368 -1254
rect 11449 -1335 11508 -1254
rect 11589 -1335 11648 -1254
rect 11729 -1257 11746 -1254
rect 11729 -1329 11878 -1257
rect 11955 -1327 12122 -1145
rect 11729 -1335 11746 -1329
rect 11070 -1349 11746 -1335
rect 10208 -1429 10234 -1383
rect 10280 -1429 10306 -1383
rect 10208 -1448 10306 -1429
rect 10208 -1477 10643 -1448
rect 10208 -1523 10234 -1477
rect 10280 -1523 10643 -1477
rect 10208 -1571 10643 -1523
rect 10208 -1617 10234 -1571
rect 10280 -1617 10643 -1571
rect 10208 -1648 10643 -1617
rect 10208 -1665 10306 -1648
rect 10208 -1711 10234 -1665
rect 10280 -1711 10306 -1665
rect 10208 -1759 10306 -1711
rect 10208 -1805 10234 -1759
rect 10280 -1805 10306 -1759
rect 10208 -1848 10306 -1805
rect 10208 -1853 10643 -1848
rect 10208 -1899 10234 -1853
rect 10280 -1899 10643 -1853
rect 10208 -1947 10643 -1899
rect 10208 -1993 10234 -1947
rect 10280 -1993 10643 -1947
rect 10208 -2041 10643 -1993
rect 10208 -2087 10234 -2041
rect 10280 -2048 10643 -2041
rect 10280 -2087 10306 -2048
rect 10208 -2135 10306 -2087
rect 10208 -2181 10234 -2135
rect 10280 -2181 10306 -2135
rect 10208 -2229 10306 -2181
rect 10208 -2275 10234 -2229
rect 10280 -2248 10306 -2229
rect 10280 -2275 10643 -2248
rect 10208 -2323 10643 -2275
rect 10208 -2369 10234 -2323
rect 10280 -2369 10643 -2323
rect 10208 -2417 10643 -2369
rect 10208 -2463 10234 -2417
rect 10280 -2448 10643 -2417
rect 10280 -2463 10306 -2448
rect 10208 -2511 10306 -2463
rect 10208 -2557 10234 -2511
rect 10280 -2557 10306 -2511
rect 10208 -2605 10306 -2557
rect 10208 -2651 10234 -2605
rect 10280 -2648 10306 -2605
rect 10280 -2651 10643 -2648
rect 10208 -2699 10643 -2651
rect 11077 -2683 11750 -2666
rect 11077 -2689 11094 -2683
rect 10208 -2745 10234 -2699
rect 10280 -2745 10643 -2699
rect 10208 -2793 10643 -2745
rect 10208 -2839 10234 -2793
rect 10280 -2839 10643 -2793
rect 10208 -2848 10643 -2839
rect 10208 -2861 10306 -2848
rect 7950 -2887 10306 -2861
rect 10753 -2874 10920 -2692
rect 10992 -2761 11094 -2689
rect 11077 -2764 11094 -2761
rect 11175 -2764 11234 -2683
rect 11315 -2764 11374 -2683
rect 11455 -2764 11514 -2683
rect 11595 -2764 11654 -2683
rect 11735 -2689 11750 -2683
rect 11735 -2761 11877 -2689
rect 11735 -2764 11750 -2761
rect 11077 -2778 11750 -2764
rect 11955 -2879 12122 -2697
rect 7950 -2933 7977 -2887
rect 8023 -2933 8071 -2887
rect 8117 -2933 8165 -2887
rect 8211 -2933 8259 -2887
rect 8305 -2933 8353 -2887
rect 8399 -2933 8447 -2887
rect 8493 -2933 8541 -2887
rect 8587 -2933 8635 -2887
rect 8681 -2933 8729 -2887
rect 8775 -2933 8823 -2887
rect 8869 -2933 8917 -2887
rect 8963 -2933 9011 -2887
rect 9057 -2933 9105 -2887
rect 9151 -2933 9199 -2887
rect 9245 -2933 9293 -2887
rect 9339 -2933 9387 -2887
rect 9433 -2933 9481 -2887
rect 9527 -2933 9575 -2887
rect 9621 -2933 9669 -2887
rect 9715 -2933 9763 -2887
rect 9809 -2933 9857 -2887
rect 9903 -2933 9951 -2887
rect 9997 -2933 10045 -2887
rect 10091 -2933 10139 -2887
rect 10185 -2933 10233 -2887
rect 10279 -2933 10306 -2887
rect 7950 -2959 10306 -2933
rect 5203 -3478 5403 -2959
rect 5603 -3478 5803 -2959
rect 6003 -3478 6203 -2959
rect 6403 -3478 6603 -2959
rect 1352 -3557 1486 -3542
rect -308 -3563 1364 -3557
rect -1134 -3807 -716 -3567
rect -308 -3649 -245 -3563
rect -161 -3565 1364 -3563
rect -161 -3649 477 -3565
rect -308 -3651 477 -3649
rect 561 -3651 621 -3565
rect 705 -3651 1364 -3565
rect -308 -3661 1364 -3651
rect 1473 -3661 1486 -3557
rect 1352 -3677 1486 -3661
rect 1858 -3678 6603 -3478
rect 1550 -3753 1688 -3738
rect 1550 -3754 1565 -3753
rect -1317 -3862 -1291 -3816
rect -1245 -3862 -1219 -3816
rect -3293 -3956 -3267 -3910
rect -3221 -3956 -3195 -3910
rect -1317 -3910 -1219 -3862
rect -3293 -4004 -3195 -3956
rect -3293 -4050 -3267 -4004
rect -3221 -4050 -3195 -4004
rect -3293 -4098 -3195 -4050
rect -2772 -3961 -2675 -3948
rect -2772 -4042 -2757 -3961
rect -2689 -4042 -2675 -3961
rect -2772 -4055 -2675 -4042
rect -2455 -3966 -2358 -3953
rect -2455 -4047 -2440 -3966
rect -2372 -4047 -2358 -3966
rect -2455 -4060 -2358 -4047
rect -2135 -3961 -2038 -3948
rect -2135 -4042 -2120 -3961
rect -2052 -4042 -2038 -3961
rect -2135 -4055 -2038 -4042
rect -1815 -3959 -1718 -3946
rect -1815 -4040 -1800 -3959
rect -1732 -4040 -1718 -3959
rect -1815 -4053 -1718 -4040
rect -1317 -3956 -1291 -3910
rect -1245 -3956 -1219 -3910
rect -1317 -4004 -1219 -3956
rect -1317 -4050 -1291 -4004
rect -1245 -4050 -1219 -4004
rect -3293 -4144 -3267 -4098
rect -3221 -4144 -3195 -4098
rect -1317 -4089 -1219 -4050
rect -956 -4089 -716 -3807
rect -308 -3761 1565 -3754
rect -308 -3847 25 -3761
rect 109 -3762 1565 -3761
rect 109 -3847 184 -3762
rect -308 -3848 184 -3847
rect 268 -3848 1565 -3762
rect -308 -3856 1565 -3848
rect 1550 -3858 1565 -3856
rect 1675 -3858 1688 -3753
rect 1550 -3873 1688 -3858
rect -488 -4068 1304 -4042
rect -488 -4089 -462 -4068
rect -1317 -4098 -462 -4089
rect -3293 -4192 -3195 -4144
rect -3293 -4238 -3267 -4192
rect -3221 -4238 -3195 -4192
rect -3095 -4119 -2998 -4106
rect -3095 -4200 -3080 -4119
rect -3012 -4200 -2998 -4119
rect -3095 -4213 -2998 -4200
rect -2938 -4122 -2841 -4109
rect -2938 -4203 -2923 -4122
rect -2855 -4203 -2841 -4122
rect -2938 -4216 -2841 -4203
rect -2295 -4123 -2198 -4110
rect -2295 -4204 -2280 -4123
rect -2212 -4204 -2198 -4123
rect -2295 -4217 -2198 -4204
rect -1658 -4120 -1561 -4107
rect -1658 -4201 -1643 -4120
rect -1575 -4201 -1561 -4120
rect -1658 -4214 -1561 -4201
rect -1493 -4118 -1396 -4105
rect -1493 -4199 -1478 -4118
rect -1410 -4199 -1396 -4118
rect -1493 -4212 -1396 -4199
rect -1317 -4144 -1291 -4098
rect -1245 -4115 -462 -4098
rect -415 -4114 -367 -4068
rect -321 -4114 -273 -4068
rect -227 -4114 -179 -4068
rect -133 -4114 -85 -4068
rect -39 -4114 9 -4068
rect 55 -4114 103 -4068
rect 149 -4114 197 -4068
rect 243 -4114 291 -4068
rect 337 -4114 385 -4068
rect 431 -4114 479 -4068
rect 525 -4114 573 -4068
rect 619 -4114 667 -4068
rect 713 -4114 761 -4068
rect 807 -4114 855 -4068
rect 901 -4114 949 -4068
rect 995 -4114 1043 -4068
rect 1089 -4114 1137 -4068
rect 1183 -4114 1231 -4068
rect -415 -4115 1231 -4114
rect 1278 -4115 1304 -4068
rect -1245 -4140 1304 -4115
rect -1245 -4144 -390 -4140
rect -1317 -4163 -390 -4144
rect -1317 -4192 -462 -4163
rect -3293 -4286 -3195 -4238
rect -3293 -4332 -3267 -4286
rect -3221 -4332 -3195 -4286
rect -1317 -4238 -1291 -4192
rect -1245 -4213 -462 -4192
rect -416 -4213 -390 -4163
rect 1206 -4163 1304 -4140
rect -1245 -4238 -390 -4213
rect 174 -4207 281 -4206
rect 174 -4220 708 -4207
rect -1317 -4261 -390 -4238
rect -1317 -4286 -462 -4261
rect -3293 -4380 -3195 -4332
rect -3068 -4373 -3022 -4315
rect -1468 -4369 -1422 -4315
rect -1317 -4332 -1291 -4286
rect -1245 -4289 -462 -4286
rect -1245 -4332 -1219 -4289
rect -3293 -4426 -3267 -4380
rect -3221 -4426 -3195 -4380
rect -3293 -4474 -3195 -4426
rect -3080 -4380 -3010 -4373
rect -3080 -4426 -3068 -4380
rect -3022 -4426 -3010 -4380
rect -1756 -4393 -1633 -4376
rect -1756 -4415 -1737 -4393
rect -3080 -4439 -3010 -4426
rect -2688 -4420 -1737 -4415
rect -2688 -4466 -2667 -4420
rect -2621 -4466 -2507 -4420
rect -2461 -4466 -2029 -4420
rect -1983 -4466 -1869 -4420
rect -1823 -4466 -1737 -4420
rect -2688 -4471 -1737 -4466
rect -3293 -4520 -3267 -4474
rect -3221 -4520 -3195 -4474
rect -1756 -4478 -1737 -4471
rect -1650 -4478 -1633 -4393
rect -1480 -4381 -1410 -4369
rect -1480 -4427 -1468 -4381
rect -1422 -4427 -1410 -4381
rect -1480 -4439 -1410 -4427
rect -1317 -4380 -1219 -4332
rect -1317 -4426 -1291 -4380
rect -1245 -4426 -1219 -4380
rect -1756 -4491 -1633 -4478
rect -1317 -4474 -1219 -4426
rect -3293 -4568 -3195 -4520
rect -3293 -4614 -3267 -4568
rect -3221 -4614 -3195 -4568
rect -1317 -4520 -1291 -4474
rect -1245 -4489 -1219 -4474
rect -956 -4489 -716 -4289
rect -488 -4307 -462 -4289
rect -416 -4307 -390 -4261
rect -488 -4355 -390 -4307
rect -310 -4245 -53 -4221
rect 174 -4232 189 -4220
rect -310 -4246 -261 -4245
rect -310 -4304 -295 -4246
rect -197 -4248 -145 -4245
rect -197 -4303 -154 -4248
rect -310 -4309 -261 -4304
rect -197 -4309 -145 -4303
rect -81 -4309 -53 -4245
rect -310 -4327 -53 -4309
rect 82 -4292 189 -4232
rect 266 -4272 708 -4220
rect 266 -4292 281 -4272
rect 82 -4306 281 -4292
rect -488 -4401 -462 -4355
rect -416 -4401 -390 -4355
rect -488 -4449 -390 -4401
rect -488 -4489 -462 -4449
rect -1245 -4495 -462 -4489
rect -416 -4495 -390 -4449
rect -1245 -4520 -390 -4495
rect -1317 -4543 -390 -4520
rect -1317 -4568 -462 -4543
rect -3068 -4582 -3022 -4571
rect -2908 -4582 -2862 -4571
rect -2748 -4582 -2702 -4571
rect -2588 -4582 -2542 -4571
rect -2428 -4582 -2382 -4571
rect -2268 -4582 -2222 -4571
rect -2108 -4582 -2062 -4571
rect -1948 -4582 -1902 -4571
rect -1788 -4582 -1742 -4571
rect -1628 -4582 -1582 -4571
rect -1468 -4582 -1422 -4571
rect -3293 -4662 -3195 -4614
rect -1317 -4614 -1291 -4568
rect -1245 -4589 -462 -4568
rect -416 -4589 -390 -4543
rect -1245 -4614 -390 -4589
rect -1317 -4637 -390 -4614
rect -3293 -4708 -3267 -4662
rect -3221 -4708 -3195 -4662
rect -3293 -4756 -3195 -4708
rect -2615 -4661 -2518 -4648
rect -2615 -4742 -2600 -4661
rect -2532 -4742 -2518 -4661
rect -2615 -4755 -2518 -4742
rect -1976 -4665 -1879 -4652
rect -1976 -4746 -1961 -4665
rect -1893 -4746 -1879 -4665
rect -3293 -4802 -3267 -4756
rect -3221 -4802 -3195 -4756
rect -1976 -4759 -1879 -4746
rect -1317 -4662 -462 -4637
rect -1317 -4708 -1291 -4662
rect -1245 -4683 -462 -4662
rect -416 -4683 -390 -4637
rect -1245 -4689 -390 -4683
rect -1245 -4708 -1219 -4689
rect -1317 -4756 -1219 -4708
rect -3293 -4850 -3195 -4802
rect -1317 -4802 -1291 -4756
rect -1245 -4802 -1219 -4756
rect -3293 -4896 -3267 -4850
rect -3221 -4896 -3195 -4850
rect -3293 -4944 -3195 -4896
rect -2775 -4819 -2678 -4806
rect -2775 -4900 -2760 -4819
rect -2692 -4900 -2678 -4819
rect -2775 -4913 -2678 -4900
rect -2457 -4823 -2360 -4810
rect -2457 -4904 -2442 -4823
rect -2374 -4904 -2360 -4823
rect -2457 -4917 -2360 -4904
rect -2131 -4817 -2034 -4804
rect -2131 -4898 -2116 -4817
rect -2048 -4898 -2034 -4817
rect -2131 -4911 -2034 -4898
rect -1817 -4828 -1720 -4815
rect -1817 -4909 -1802 -4828
rect -1734 -4909 -1720 -4828
rect -1817 -4922 -1720 -4909
rect -1317 -4850 -1219 -4802
rect -1317 -4896 -1291 -4850
rect -1245 -4889 -1219 -4850
rect -956 -4889 -716 -4689
rect -488 -4731 -390 -4689
rect -488 -4777 -462 -4731
rect -416 -4777 -390 -4731
rect -488 -4825 -390 -4777
rect -488 -4871 -462 -4825
rect -416 -4871 -390 -4825
rect -488 -4889 -390 -4871
rect -1245 -4896 -390 -4889
rect -1317 -4919 -390 -4896
rect -3293 -4990 -3267 -4944
rect -3221 -4990 -3195 -4944
rect -1317 -4944 -462 -4919
rect -3293 -5038 -3195 -4990
rect -3293 -5084 -3267 -5038
rect -3221 -5084 -3195 -5038
rect -3092 -4969 -2995 -4956
rect -3092 -5050 -3077 -4969
rect -3009 -5050 -2995 -4969
rect -3092 -5063 -2995 -5050
rect -2935 -4972 -2838 -4959
rect -2935 -5053 -2920 -4972
rect -2852 -5053 -2838 -4972
rect -2935 -5066 -2838 -5053
rect -2295 -4974 -2198 -4961
rect -2295 -5055 -2280 -4974
rect -2212 -5055 -2198 -4974
rect -2295 -5068 -2198 -5055
rect -1651 -4975 -1554 -4962
rect -1651 -5056 -1636 -4975
rect -1568 -5056 -1554 -4975
rect -1651 -5069 -1554 -5056
rect -1494 -4971 -1397 -4958
rect -1494 -5052 -1479 -4971
rect -1411 -5052 -1397 -4971
rect -1494 -5065 -1397 -5052
rect -1317 -4990 -1291 -4944
rect -1245 -4965 -462 -4944
rect -416 -4965 -390 -4919
rect -1245 -4990 -390 -4965
rect -1317 -5013 -390 -4990
rect -1317 -5038 -462 -5013
rect -3293 -5132 -3195 -5084
rect -3293 -5178 -3267 -5132
rect -3221 -5178 -3195 -5132
rect -1317 -5084 -1291 -5038
rect -1245 -5059 -462 -5038
rect -416 -5059 -390 -5013
rect -1245 -5084 -390 -5059
rect -1317 -5089 -390 -5084
rect -1317 -5132 -1219 -5089
rect -3293 -5226 -3195 -5178
rect -3068 -5219 -3022 -5156
rect -2908 -5167 -2862 -5156
rect -2748 -5167 -2702 -5156
rect -2588 -5167 -2542 -5156
rect -2428 -5167 -2382 -5156
rect -2268 -5167 -2222 -5156
rect -2108 -5167 -2062 -5156
rect -1948 -5167 -1902 -5156
rect -1788 -5167 -1742 -5156
rect -1628 -5167 -1582 -5156
rect -3293 -5272 -3267 -5226
rect -3221 -5272 -3195 -5226
rect -3293 -5320 -3195 -5272
rect -3081 -5231 -3009 -5219
rect -1468 -5223 -1422 -5156
rect -1317 -5178 -1291 -5132
rect -1245 -5178 -1219 -5132
rect -3081 -5277 -3068 -5231
rect -3022 -5277 -3009 -5231
rect -1480 -5232 -1410 -5223
rect -3081 -5289 -3009 -5277
rect -2861 -5252 -2740 -5234
rect -3293 -5366 -3267 -5320
rect -3221 -5366 -3195 -5320
rect -2861 -5337 -2845 -5252
rect -2759 -5267 -2740 -5252
rect -2363 -5263 -2285 -5246
rect -2363 -5267 -2348 -5263
rect -2759 -5281 -2348 -5267
rect -2759 -5323 -2668 -5281
rect -2759 -5337 -2740 -5323
rect -2861 -5352 -2740 -5337
rect -2684 -5327 -2668 -5323
rect -2622 -5282 -2348 -5281
rect -2622 -5323 -2508 -5282
rect -2622 -5327 -2606 -5323
rect -2684 -5344 -2606 -5327
rect -2524 -5328 -2508 -5323
rect -2462 -5309 -2348 -5282
rect -2302 -5267 -2285 -5263
rect -2205 -5263 -2127 -5246
rect -2205 -5267 -2188 -5263
rect -2302 -5309 -2188 -5267
rect -2142 -5267 -2127 -5263
rect -1723 -5260 -1645 -5246
rect -1723 -5267 -1707 -5260
rect -2142 -5281 -1707 -5267
rect -2142 -5282 -1868 -5281
rect -2142 -5309 -2028 -5282
rect -2462 -5323 -2028 -5309
rect -2462 -5328 -2446 -5323
rect -2524 -5344 -2446 -5328
rect -2044 -5328 -2028 -5323
rect -1982 -5323 -1868 -5282
rect -1982 -5328 -1966 -5323
rect -2044 -5344 -1966 -5328
rect -1884 -5327 -1868 -5323
rect -1822 -5306 -1707 -5281
rect -1661 -5306 -1645 -5260
rect -1480 -5278 -1468 -5232
rect -1422 -5278 -1410 -5232
rect -1480 -5291 -1410 -5278
rect -1317 -5226 -1219 -5178
rect -1317 -5272 -1291 -5226
rect -1245 -5272 -1219 -5226
rect -1317 -5289 -1219 -5272
rect -956 -5289 -716 -5089
rect -488 -5107 -390 -5089
rect -488 -5153 -462 -5107
rect -416 -5153 -390 -5107
rect -488 -5201 -390 -5153
rect -488 -5247 -462 -5201
rect -416 -5247 -390 -5201
rect -488 -5289 -390 -5247
rect -1822 -5323 -1645 -5306
rect -1317 -5295 -390 -5289
rect -1317 -5320 -462 -5295
rect -1822 -5327 -1806 -5323
rect -1884 -5344 -1806 -5327
rect -3293 -5414 -3195 -5366
rect -3293 -5460 -3267 -5414
rect -3221 -5460 -3195 -5414
rect -1317 -5366 -1291 -5320
rect -1245 -5341 -462 -5320
rect -416 -5341 -390 -5295
rect -1245 -5366 -390 -5341
rect -1317 -5389 -390 -5366
rect -1317 -5414 -462 -5389
rect -3068 -5434 -3022 -5423
rect -2908 -5434 -2862 -5423
rect -2748 -5434 -2702 -5423
rect -2588 -5434 -2542 -5423
rect -2428 -5434 -2382 -5423
rect -2268 -5434 -2222 -5423
rect -2108 -5434 -2062 -5423
rect -1948 -5434 -1902 -5423
rect -1788 -5434 -1742 -5423
rect -1628 -5434 -1582 -5423
rect -1468 -5434 -1422 -5423
rect -3293 -5508 -3195 -5460
rect -3293 -5554 -3267 -5508
rect -3221 -5554 -3195 -5508
rect -1317 -5460 -1291 -5414
rect -1245 -5435 -462 -5414
rect -416 -5435 -390 -5389
rect -1245 -5460 -390 -5435
rect -1317 -5483 -390 -5460
rect -1317 -5489 -462 -5483
rect -1317 -5508 -1219 -5489
rect -3293 -5602 -3195 -5554
rect -3293 -5648 -3267 -5602
rect -3221 -5648 -3195 -5602
rect -2613 -5528 -2516 -5515
rect -2613 -5609 -2598 -5528
rect -2530 -5609 -2516 -5528
rect -2613 -5622 -2516 -5609
rect -1970 -5527 -1873 -5514
rect -1970 -5608 -1955 -5527
rect -1887 -5608 -1873 -5527
rect -1970 -5621 -1873 -5608
rect -1317 -5554 -1291 -5508
rect -1245 -5554 -1219 -5508
rect -1317 -5602 -1219 -5554
rect -3293 -5696 -3195 -5648
rect -1317 -5648 -1291 -5602
rect -1245 -5648 -1219 -5602
rect -3293 -5742 -3267 -5696
rect -3221 -5742 -3195 -5696
rect -3293 -5790 -3195 -5742
rect -2778 -5679 -2681 -5666
rect -2778 -5760 -2763 -5679
rect -2695 -5760 -2681 -5679
rect -2778 -5773 -2681 -5760
rect -2456 -5678 -2359 -5665
rect -2456 -5759 -2441 -5678
rect -2373 -5759 -2359 -5678
rect -2456 -5772 -2359 -5759
rect -2141 -5686 -2044 -5673
rect -2141 -5767 -2126 -5686
rect -2058 -5767 -2044 -5686
rect -2141 -5780 -2044 -5767
rect -1812 -5684 -1715 -5671
rect -1812 -5765 -1797 -5684
rect -1729 -5765 -1715 -5684
rect -1812 -5778 -1715 -5765
rect -1317 -5689 -1219 -5648
rect -956 -5689 -716 -5489
rect -488 -5529 -462 -5489
rect -416 -5529 -390 -5483
rect -488 -5577 -390 -5529
rect -488 -5623 -462 -5577
rect -416 -5623 -390 -5577
rect -488 -5671 -390 -5623
rect -488 -5689 -462 -5671
rect -1317 -5696 -462 -5689
rect -1317 -5742 -1291 -5696
rect -1245 -5717 -462 -5696
rect -416 -5717 -390 -5671
rect -1245 -5742 -390 -5717
rect -1317 -5765 -390 -5742
rect -3293 -5836 -3267 -5790
rect -3221 -5836 -3195 -5790
rect -1317 -5790 -462 -5765
rect -3293 -5884 -3195 -5836
rect -3293 -5930 -3267 -5884
rect -3221 -5930 -3195 -5884
rect -3293 -5978 -3195 -5930
rect -3092 -5844 -2995 -5831
rect -3092 -5925 -3077 -5844
rect -3009 -5925 -2995 -5844
rect -3092 -5938 -2995 -5925
rect -2930 -5842 -2833 -5829
rect -2930 -5923 -2915 -5842
rect -2847 -5923 -2833 -5842
rect -2930 -5936 -2833 -5923
rect -2291 -5837 -2197 -5824
rect -2291 -5918 -2279 -5837
rect -2211 -5918 -2197 -5837
rect -2291 -5931 -2197 -5918
rect -1659 -5837 -1562 -5824
rect -1659 -5918 -1644 -5837
rect -1576 -5918 -1562 -5837
rect -1659 -5931 -1562 -5918
rect -1491 -5839 -1394 -5826
rect -1491 -5920 -1476 -5839
rect -1408 -5920 -1394 -5839
rect -1491 -5933 -1394 -5920
rect -1317 -5836 -1291 -5790
rect -1245 -5811 -462 -5790
rect -416 -5811 -390 -5765
rect -1245 -5836 -390 -5811
rect -1317 -5859 -390 -5836
rect -1317 -5884 -462 -5859
rect -1317 -5930 -1291 -5884
rect -1245 -5889 -462 -5884
rect -1245 -5930 -1219 -5889
rect -3293 -6024 -3267 -5978
rect -3221 -6024 -3195 -5978
rect -1317 -5978 -1219 -5930
rect -3293 -6072 -3195 -6024
rect -3068 -6069 -3022 -6008
rect -2908 -6019 -2862 -6008
rect -2748 -6019 -2702 -6008
rect -2588 -6019 -2542 -6008
rect -2428 -6019 -2382 -6008
rect -2268 -6019 -2222 -6008
rect -2108 -6019 -2062 -6008
rect -1948 -6019 -1902 -6008
rect -1788 -6019 -1742 -6008
rect -1628 -6019 -1582 -6008
rect -3293 -6118 -3267 -6072
rect -3221 -6118 -3195 -6072
rect -3293 -6166 -3195 -6118
rect -3080 -6081 -3011 -6069
rect -3080 -6127 -3068 -6081
rect -3022 -6127 -3011 -6081
rect -1744 -6076 -1640 -6065
rect -1468 -6074 -1422 -6008
rect -1317 -6024 -1291 -5978
rect -1245 -6024 -1219 -5978
rect -1317 -6072 -1219 -6024
rect -1744 -6087 -1731 -6076
rect -3080 -6139 -3011 -6127
rect -2849 -6093 -1731 -6087
rect -2849 -6139 -2828 -6093
rect -2782 -6139 -2348 -6093
rect -2302 -6139 -2188 -6093
rect -2142 -6139 -1731 -6093
rect -2849 -6143 -1731 -6139
rect -1744 -6156 -1731 -6143
rect -1651 -6156 -1640 -6076
rect -1481 -6085 -1410 -6074
rect -1481 -6131 -1468 -6085
rect -1422 -6131 -1410 -6085
rect -1481 -6143 -1410 -6131
rect -1317 -6118 -1291 -6072
rect -1245 -6089 -1219 -6072
rect -956 -6089 -716 -5889
rect -488 -5905 -462 -5889
rect -416 -5905 -390 -5859
rect -238 -5142 -188 -4488
rect -97 -5142 -15 -4487
rect -238 -5148 -15 -5142
rect -238 -5194 -156 -5148
rect -110 -5194 -15 -5148
rect -238 -5201 -15 -5194
rect -238 -5868 -188 -5201
rect -488 -5953 -390 -5905
rect -488 -5999 -462 -5953
rect -416 -5999 -390 -5953
rect -488 -6047 -390 -5999
rect -97 -6030 -15 -5201
rect 82 -5868 132 -4306
rect 341 -4336 447 -4319
rect 341 -4415 355 -4336
rect 434 -4415 447 -4336
rect 341 -4430 447 -4415
rect 210 -5950 260 -4488
rect 360 -5871 430 -4430
rect 337 -5939 449 -5922
rect 337 -5950 353 -5939
rect 210 -6000 353 -5950
rect 337 -6024 353 -6000
rect 435 -5950 449 -5939
rect 530 -5950 580 -4488
rect 658 -5868 708 -4272
rect 1206 -4213 1232 -4163
rect 1278 -4213 1304 -4163
rect 1206 -4261 1304 -4213
rect 1206 -4307 1232 -4261
rect 1278 -4307 1304 -4261
rect 1858 -4293 2058 -3678
rect 2403 -4293 2603 -3678
rect 2803 -4293 3003 -3678
rect 3203 -4293 3403 -3678
rect 3603 -4293 3803 -3678
rect 1206 -4320 1304 -4307
rect 1595 -4301 3803 -4293
rect 4003 -3969 4203 -3678
rect 4403 -3969 4603 -3678
rect 4826 -3969 5022 -3678
rect 5203 -3969 5403 -3678
rect 5603 -3969 5803 -3678
rect 6003 -3969 6203 -3678
rect 6403 -3969 6603 -3678
rect 4003 -4169 6603 -3969
rect 1595 -4319 3763 -4301
rect 1595 -4320 1622 -4319
rect 1206 -4355 1622 -4320
rect 1206 -4401 1232 -4355
rect 1278 -4365 1622 -4355
rect 1668 -4365 1716 -4319
rect 1762 -4365 1810 -4319
rect 1856 -4365 1904 -4319
rect 1950 -4365 1998 -4319
rect 2044 -4365 2092 -4319
rect 2138 -4365 2186 -4319
rect 2232 -4365 2280 -4319
rect 2326 -4365 2374 -4319
rect 2420 -4365 2468 -4319
rect 2514 -4365 2562 -4319
rect 2608 -4365 2656 -4319
rect 2702 -4365 2750 -4319
rect 2796 -4365 2844 -4319
rect 2890 -4365 2938 -4319
rect 2984 -4365 3032 -4319
rect 3078 -4365 3126 -4319
rect 3172 -4365 3220 -4319
rect 3266 -4365 3314 -4319
rect 3360 -4365 3408 -4319
rect 3454 -4365 3502 -4319
rect 3548 -4365 3596 -4319
rect 3642 -4365 3690 -4319
rect 3736 -4365 3763 -4319
rect 1278 -4391 3763 -4365
rect 1278 -4401 1693 -4391
rect 1206 -4413 1693 -4401
rect 1206 -4449 1621 -4413
rect 802 -4852 884 -4486
rect 802 -4916 811 -4852
rect 875 -4916 884 -4852
rect 802 -4968 884 -4916
rect 802 -5032 811 -4968
rect 875 -5032 884 -4968
rect 802 -5146 884 -5032
rect 978 -5146 1028 -4488
rect 802 -5152 1028 -5146
rect 802 -5198 901 -5152
rect 947 -5198 1028 -5152
rect 802 -5205 1028 -5198
rect 802 -5533 884 -5205
rect 802 -5597 810 -5533
rect 874 -5597 884 -5533
rect 802 -5649 884 -5597
rect 802 -5713 810 -5649
rect 874 -5713 884 -5649
rect 435 -6000 580 -5950
rect 435 -6024 449 -6000
rect -488 -6089 -462 -6047
rect -1245 -6093 -462 -6089
rect -416 -6093 -390 -6047
rect -1245 -6118 -390 -6093
rect -1317 -6141 -390 -6118
rect -1744 -6166 -1640 -6156
rect -1317 -6166 -462 -6141
rect -3293 -6212 -3267 -6166
rect -3221 -6212 -3195 -6166
rect -3293 -6234 -3195 -6212
rect -1317 -6212 -1291 -6166
rect -1245 -6187 -462 -6166
rect -416 -6187 -390 -6141
rect -146 -6049 148 -6030
rect 337 -6038 449 -6024
rect -146 -6052 50 -6049
rect -146 -6137 -109 -6052
rect -27 -6134 50 -6052
rect 132 -6064 148 -6049
rect 802 -6064 884 -5713
rect 978 -5868 1028 -5205
rect 1206 -4495 1232 -4449
rect 1278 -4459 1621 -4449
rect 1667 -4459 1693 -4413
rect 1278 -4495 1693 -4459
rect 1206 -4507 1693 -4495
rect 1206 -4520 1621 -4507
rect 1206 -4543 1304 -4520
rect 1206 -4589 1232 -4543
rect 1278 -4589 1304 -4543
rect 1206 -4637 1304 -4589
rect 1206 -4683 1232 -4637
rect 1278 -4683 1304 -4637
rect 1206 -4720 1304 -4683
rect 1595 -4553 1621 -4520
rect 1667 -4553 1693 -4507
rect 1595 -4601 1693 -4553
rect 1595 -4647 1621 -4601
rect 1667 -4647 1693 -4601
rect 1595 -4695 1693 -4647
rect 1595 -4720 1621 -4695
rect 1206 -4731 1621 -4720
rect 1206 -4777 1232 -4731
rect 1278 -4741 1621 -4731
rect 1667 -4741 1693 -4695
rect 1278 -4777 1693 -4741
rect 1206 -4789 1693 -4777
rect 1206 -4825 1621 -4789
rect 1206 -4871 1232 -4825
rect 1278 -4835 1621 -4825
rect 1667 -4835 1693 -4789
rect 1278 -4871 1693 -4835
rect 1206 -4883 1693 -4871
rect 1206 -4919 1621 -4883
rect 1206 -4965 1232 -4919
rect 1278 -4920 1621 -4919
rect 1278 -4965 1304 -4920
rect 1206 -5013 1304 -4965
rect 1206 -5059 1232 -5013
rect 1278 -5059 1304 -5013
rect 1206 -5107 1304 -5059
rect 1206 -5153 1232 -5107
rect 1278 -5120 1304 -5107
rect 1595 -4929 1621 -4920
rect 1667 -4929 1693 -4883
rect 1595 -4977 1693 -4929
rect 1595 -5023 1621 -4977
rect 1667 -5023 1693 -4977
rect 1595 -5071 1693 -5023
rect 1595 -5117 1621 -5071
rect 1667 -5117 1693 -5071
rect 1595 -5120 1693 -5117
rect 1278 -5153 1693 -5120
rect 1206 -5165 1693 -5153
rect 1206 -5201 1621 -5165
rect 1206 -5247 1232 -5201
rect 1278 -5211 1621 -5201
rect 1667 -5211 1693 -5165
rect 1278 -5247 1693 -5211
rect 1206 -5259 1693 -5247
rect 1206 -5295 1621 -5259
rect 1206 -5341 1232 -5295
rect 1278 -5305 1621 -5295
rect 1667 -5305 1693 -5259
rect 1779 -5201 1837 -4391
rect 1995 -5135 2053 -4391
rect 2191 -4800 2288 -4782
rect 2191 -4864 2208 -4800
rect 2272 -4864 2288 -4800
rect 2191 -4916 2288 -4864
rect 2191 -4980 2208 -4916
rect 2272 -4980 2288 -4916
rect 2191 -4994 2288 -4980
rect 2427 -5137 2485 -4391
rect 2561 -4479 2799 -4461
rect 2561 -4543 2579 -4479
rect 2643 -4543 2719 -4479
rect 2783 -4543 2799 -4479
rect 2561 -4595 2799 -4543
rect 2561 -4659 2579 -4595
rect 2643 -4655 2713 -4595
rect 2643 -4659 2719 -4655
rect 2783 -4659 2799 -4595
rect 2561 -4677 2799 -4659
rect 1779 -5213 1936 -5201
rect 1779 -5271 1865 -5213
rect 1923 -5271 1936 -5213
rect 1779 -5283 1936 -5271
rect 1278 -5320 1693 -5305
rect 1278 -5341 1304 -5320
rect 1206 -5389 1304 -5341
rect 1206 -5435 1232 -5389
rect 1278 -5435 1304 -5389
rect 1206 -5483 1304 -5435
rect 1206 -5529 1232 -5483
rect 1278 -5520 1304 -5483
rect 1595 -5353 1693 -5320
rect 1595 -5399 1621 -5353
rect 1667 -5399 1693 -5353
rect 1595 -5447 1693 -5399
rect 2427 -5321 2513 -5307
rect 2427 -5381 2441 -5321
rect 2501 -5325 2513 -5321
rect 2644 -5325 2699 -4677
rect 2860 -5136 2918 -4391
rect 3053 -4809 3150 -4791
rect 3053 -4873 3070 -4809
rect 3134 -4873 3150 -4809
rect 3053 -4925 3150 -4873
rect 3053 -4989 3070 -4925
rect 3134 -4989 3150 -4925
rect 3053 -5003 3150 -4989
rect 3291 -5136 3349 -4391
rect 3507 -5201 3565 -4391
rect 3408 -5213 3565 -5201
rect 3408 -5271 3421 -5213
rect 3479 -5271 3565 -5213
rect 3408 -5283 3565 -5271
rect 3665 -4413 3763 -4391
rect 4003 -4396 4203 -4169
rect 4403 -4396 4603 -4169
rect 4826 -4396 5022 -4169
rect 5203 -4396 5403 -4169
rect 5603 -4396 5803 -4169
rect 6003 -4396 6203 -4169
rect 6403 -4396 6603 -4169
rect 3665 -4459 3691 -4413
rect 3737 -4459 3763 -4413
rect 3665 -4507 3763 -4459
rect 3665 -4553 3691 -4507
rect 3737 -4553 3763 -4507
rect 3665 -4601 3763 -4553
rect 3665 -4647 3691 -4601
rect 3737 -4647 3763 -4601
rect 3665 -4665 3763 -4647
rect 4002 -4422 6734 -4396
rect 4002 -4468 4029 -4422
rect 4075 -4468 4123 -4422
rect 4169 -4468 4217 -4422
rect 4263 -4468 4311 -4422
rect 4357 -4468 4405 -4422
rect 4451 -4468 4499 -4422
rect 4545 -4468 4593 -4422
rect 4639 -4468 4687 -4422
rect 4733 -4468 4781 -4422
rect 4827 -4468 4875 -4422
rect 4921 -4468 4969 -4422
rect 5015 -4468 5063 -4422
rect 5109 -4468 5157 -4422
rect 5203 -4468 5251 -4422
rect 5297 -4468 5345 -4422
rect 5391 -4468 5439 -4422
rect 5485 -4468 5533 -4422
rect 5579 -4468 5627 -4422
rect 5673 -4468 5721 -4422
rect 5767 -4468 5815 -4422
rect 5861 -4468 5909 -4422
rect 5955 -4468 6003 -4422
rect 6049 -4468 6097 -4422
rect 6143 -4468 6191 -4422
rect 6237 -4468 6285 -4422
rect 6331 -4468 6379 -4422
rect 6425 -4468 6473 -4422
rect 6519 -4468 6567 -4422
rect 6613 -4468 6661 -4422
rect 6707 -4468 6734 -4422
rect 4002 -4494 6734 -4468
rect 4002 -4516 4100 -4494
rect 4002 -4562 4028 -4516
rect 4074 -4562 4100 -4516
rect 4002 -4610 4100 -4562
rect 4002 -4656 4028 -4610
rect 4074 -4656 4100 -4610
rect 4002 -4665 4100 -4656
rect 3665 -4695 4100 -4665
rect 3665 -4741 3691 -4695
rect 3737 -4704 4100 -4695
rect 3737 -4741 4028 -4704
rect 3665 -4750 4028 -4741
rect 4074 -4750 4100 -4704
rect 3665 -4789 4100 -4750
rect 3665 -4835 3691 -4789
rect 3737 -4798 4100 -4789
rect 3737 -4835 4028 -4798
rect 3665 -4844 4028 -4835
rect 4074 -4844 4100 -4798
rect 3665 -4865 4100 -4844
rect 3665 -4883 3763 -4865
rect 3665 -4929 3691 -4883
rect 3737 -4929 3763 -4883
rect 3665 -4977 3763 -4929
rect 3665 -5023 3691 -4977
rect 3737 -5023 3763 -4977
rect 3665 -5065 3763 -5023
rect 4002 -4892 4100 -4865
rect 4002 -4938 4028 -4892
rect 4074 -4938 4100 -4892
rect 4002 -4986 4100 -4938
rect 4002 -5032 4028 -4986
rect 4074 -5032 4100 -4986
rect 4002 -5065 4100 -5032
rect 3665 -5071 4100 -5065
rect 3665 -5117 3691 -5071
rect 3737 -5080 4100 -5071
rect 3737 -5117 4028 -5080
rect 3665 -5126 4028 -5117
rect 4074 -5126 4100 -5080
rect 3665 -5165 4100 -5126
rect 3665 -5211 3691 -5165
rect 3737 -5174 4100 -5165
rect 3737 -5211 4028 -5174
rect 3665 -5220 4028 -5211
rect 4074 -5220 4100 -5174
rect 3665 -5259 4100 -5220
rect 2501 -5380 2699 -5325
rect 3665 -5305 3691 -5259
rect 3737 -5265 4100 -5259
rect 3737 -5305 3763 -5265
rect 3665 -5353 3763 -5305
rect 2501 -5381 2513 -5380
rect 2427 -5394 2513 -5381
rect 1595 -5493 1621 -5447
rect 1667 -5493 1693 -5447
rect 1595 -5520 1693 -5493
rect 1278 -5529 1693 -5520
rect 1206 -5541 1693 -5529
rect 1206 -5577 1621 -5541
rect 1206 -5623 1232 -5577
rect 1278 -5587 1621 -5577
rect 1667 -5587 1693 -5541
rect 1278 -5623 1693 -5587
rect 1206 -5635 1693 -5623
rect 1206 -5671 1621 -5635
rect 1206 -5717 1232 -5671
rect 1278 -5681 1621 -5671
rect 1667 -5681 1693 -5635
rect 1278 -5717 1693 -5681
rect 1206 -5720 1693 -5717
rect 1206 -5765 1304 -5720
rect 1206 -5811 1232 -5765
rect 1278 -5811 1304 -5765
rect 1206 -5859 1304 -5811
rect 132 -6102 295 -6064
rect 496 -6102 884 -6064
rect 132 -6134 884 -6102
rect -27 -6137 884 -6134
rect -146 -6151 884 -6137
rect 1206 -5905 1232 -5859
rect 1278 -5905 1304 -5859
rect 1206 -5920 1304 -5905
rect 1595 -5729 1693 -5720
rect 1595 -5775 1621 -5729
rect 1667 -5775 1693 -5729
rect 1595 -5823 1693 -5775
rect 1595 -5869 1621 -5823
rect 1667 -5869 1693 -5823
rect 1595 -5917 1693 -5869
rect 1595 -5920 1621 -5917
rect 1206 -5953 1621 -5920
rect 1206 -5999 1232 -5953
rect 1278 -5963 1621 -5953
rect 1667 -5963 1693 -5917
rect 1278 -5999 1693 -5963
rect 1206 -6011 1693 -5999
rect 1206 -6047 1621 -6011
rect 1206 -6093 1232 -6047
rect 1278 -6057 1621 -6047
rect 1667 -6057 1693 -6011
rect 1278 -6093 1693 -6057
rect 1206 -6105 1693 -6093
rect 1206 -6120 1621 -6105
rect 1206 -6141 1304 -6120
rect -146 -6152 547 -6151
rect -146 -6161 148 -6152
rect 275 -6159 547 -6152
rect -1245 -6210 -390 -6187
rect 1206 -6187 1232 -6141
rect 1278 -6187 1304 -6141
rect 1206 -6210 1304 -6187
rect -1245 -6212 1304 -6210
rect -1317 -6234 1304 -6212
rect -3293 -6235 1304 -6234
rect -3293 -6260 -462 -6235
rect -3293 -6306 -3266 -6260
rect -3220 -6306 -3172 -6260
rect -3126 -6306 -3078 -6260
rect -3032 -6306 -2984 -6260
rect -2938 -6306 -2890 -6260
rect -2844 -6306 -2796 -6260
rect -2750 -6306 -2702 -6260
rect -2656 -6306 -2608 -6260
rect -2562 -6306 -2514 -6260
rect -2468 -6306 -2420 -6260
rect -2374 -6306 -2326 -6260
rect -2280 -6306 -2232 -6260
rect -2186 -6306 -2138 -6260
rect -2092 -6306 -2044 -6260
rect -1998 -6306 -1950 -6260
rect -1904 -6306 -1856 -6260
rect -1810 -6306 -1762 -6260
rect -1716 -6306 -1668 -6260
rect -1622 -6306 -1574 -6260
rect -1528 -6306 -1480 -6260
rect -1434 -6306 -1386 -6260
rect -1340 -6306 -1292 -6260
rect -1246 -6282 -462 -6260
rect -415 -6236 1231 -6235
rect -415 -6282 -367 -6236
rect -321 -6282 -273 -6236
rect -227 -6282 -179 -6236
rect -133 -6282 -85 -6236
rect -39 -6282 9 -6236
rect 55 -6282 103 -6236
rect 149 -6282 197 -6236
rect 243 -6282 291 -6236
rect 337 -6282 385 -6236
rect 431 -6282 479 -6236
rect 525 -6282 573 -6236
rect 619 -6282 667 -6236
rect 713 -6282 761 -6236
rect 807 -6282 855 -6236
rect 901 -6282 949 -6236
rect 995 -6282 1043 -6236
rect 1089 -6282 1137 -6236
rect 1183 -6282 1231 -6236
rect 1278 -6282 1304 -6235
rect 1595 -6151 1621 -6120
rect 1667 -6151 1693 -6105
rect 1595 -6173 1693 -6151
rect 1865 -5907 1923 -5440
rect 1865 -5919 2022 -5907
rect 1865 -5977 1951 -5919
rect 2009 -5977 2022 -5919
rect 1865 -5989 2022 -5977
rect 1865 -6173 1923 -5989
rect 2081 -6173 2139 -5443
rect 2294 -5859 2352 -5442
rect 2427 -5842 2485 -5394
rect 3665 -5399 3691 -5353
rect 3737 -5399 3763 -5353
rect 2273 -5877 2370 -5859
rect 2273 -5941 2290 -5877
rect 2354 -5941 2370 -5877
rect 2273 -5993 2370 -5941
rect 2273 -6057 2290 -5993
rect 2354 -6057 2370 -5993
rect 2273 -6071 2370 -6057
rect 2643 -6173 2701 -5444
rect 2829 -5522 2926 -5504
rect 2829 -5586 2846 -5522
rect 2910 -5586 2926 -5522
rect 2829 -5638 2926 -5586
rect 2829 -5702 2846 -5638
rect 2910 -5702 2926 -5638
rect 2829 -5716 2926 -5702
rect 2989 -5872 3047 -5442
rect 2989 -5890 3146 -5872
rect 2989 -5954 3018 -5890
rect 3082 -5919 3146 -5890
rect 2989 -5977 3075 -5954
rect 3133 -5977 3146 -5919
rect 2989 -6006 3146 -5977
rect 2989 -6070 3018 -6006
rect 3082 -6070 3146 -6006
rect 2989 -6091 3146 -6070
rect 3205 -6173 3263 -5441
rect 3421 -5907 3479 -5441
rect 3322 -5919 3479 -5907
rect 3322 -5977 3335 -5919
rect 3393 -5977 3479 -5919
rect 3322 -5989 3479 -5977
rect 3421 -6173 3479 -5989
rect 3665 -5447 3763 -5399
rect 3665 -5493 3691 -5447
rect 3737 -5465 3763 -5447
rect 4002 -5268 4100 -5265
rect 4002 -5314 4028 -5268
rect 4074 -5314 4100 -5268
rect 4002 -5362 4100 -5314
rect 4002 -5408 4028 -5362
rect 4074 -5408 4100 -5362
rect 4002 -5456 4100 -5408
rect 4002 -5465 4028 -5456
rect 3737 -5493 4028 -5465
rect 3665 -5502 4028 -5493
rect 4074 -5502 4100 -5456
rect 3665 -5541 4100 -5502
rect 3665 -5587 3691 -5541
rect 3737 -5550 4100 -5541
rect 3737 -5587 4028 -5550
rect 3665 -5596 4028 -5587
rect 4074 -5596 4100 -5550
rect 3665 -5635 4100 -5596
rect 3665 -5681 3691 -5635
rect 3737 -5644 4100 -5635
rect 3737 -5665 4028 -5644
rect 3737 -5681 3763 -5665
rect 3665 -5729 3763 -5681
rect 3665 -5775 3691 -5729
rect 3737 -5775 3763 -5729
rect 3665 -5823 3763 -5775
rect 3665 -5869 3691 -5823
rect 3737 -5865 3763 -5823
rect 4002 -5690 4028 -5665
rect 4074 -5690 4100 -5644
rect 4002 -5738 4100 -5690
rect 4002 -5784 4028 -5738
rect 4074 -5784 4100 -5738
rect 4002 -5832 4100 -5784
rect 4002 -5865 4028 -5832
rect 3737 -5869 4028 -5865
rect 3665 -5878 4028 -5869
rect 4074 -5878 4100 -5832
rect 3665 -5917 4100 -5878
rect 3665 -5963 3691 -5917
rect 3737 -5926 4100 -5917
rect 3737 -5963 4028 -5926
rect 3665 -5972 4028 -5963
rect 4074 -5972 4100 -5926
rect 3665 -5994 4100 -5972
rect 4199 -5199 4263 -4494
rect 4502 -5199 4566 -4494
rect 4806 -4909 4870 -4755
rect 4790 -4927 4887 -4909
rect 4790 -4991 4807 -4927
rect 4871 -4991 4887 -4927
rect 4790 -5043 4887 -4991
rect 4790 -5107 4807 -5043
rect 4871 -5107 4887 -5043
rect 4790 -5121 4887 -5107
rect 4199 -5212 4566 -5199
rect 4199 -5262 4302 -5212
rect 4352 -5262 4415 -5212
rect 4465 -5262 4566 -5212
rect 4199 -5274 4566 -5262
rect 4199 -5994 4263 -5274
rect 4502 -5994 4566 -5274
rect 4806 -5428 4870 -5121
rect 4790 -5446 4887 -5428
rect 4790 -5510 4807 -5446
rect 4871 -5510 4887 -5446
rect 4790 -5562 4887 -5510
rect 4790 -5626 4807 -5562
rect 4871 -5626 4887 -5562
rect 4790 -5640 4887 -5626
rect 4806 -5743 4870 -5640
rect 5111 -5994 5175 -4494
rect 5241 -4629 5476 -4615
rect 5241 -4695 5256 -4629
rect 5322 -4695 5394 -4629
rect 5460 -4695 5476 -4629
rect 5241 -4708 5476 -4695
rect 5412 -5197 5476 -4708
rect 5289 -5209 5476 -5197
rect 5289 -5261 5302 -5209
rect 5354 -5261 5476 -5209
rect 5289 -5273 5476 -5261
rect 5412 -5390 5476 -5273
rect 5394 -5408 5491 -5390
rect 5394 -5472 5411 -5408
rect 5475 -5472 5491 -5408
rect 5394 -5524 5491 -5472
rect 5394 -5588 5411 -5524
rect 5475 -5588 5491 -5524
rect 5394 -5602 5491 -5588
rect 5412 -5774 5476 -5602
rect 5241 -5788 5476 -5774
rect 5241 -5854 5256 -5788
rect 5322 -5854 5394 -5788
rect 5460 -5854 5476 -5788
rect 5241 -5867 5476 -5854
rect 5555 -5994 5619 -4494
rect 5857 -4906 5921 -4759
rect 5842 -4924 5939 -4906
rect 5842 -4988 5859 -4924
rect 5923 -4988 5939 -4924
rect 5842 -5040 5939 -4988
rect 5842 -5104 5859 -5040
rect 5923 -5104 5939 -5040
rect 5842 -5118 5939 -5104
rect 5857 -5425 5921 -5118
rect 6160 -5201 6224 -4494
rect 6464 -5201 6528 -4494
rect 6160 -5214 6528 -5201
rect 6160 -5264 6264 -5214
rect 6314 -5264 6377 -5214
rect 6427 -5264 6528 -5214
rect 6160 -5276 6528 -5264
rect 5842 -5443 5939 -5425
rect 5842 -5507 5859 -5443
rect 5923 -5507 5939 -5443
rect 5842 -5559 5939 -5507
rect 5842 -5623 5859 -5559
rect 5923 -5623 5939 -5559
rect 5842 -5637 5939 -5623
rect 5857 -5745 5921 -5637
rect 6160 -5994 6224 -5276
rect 6464 -5994 6528 -5276
rect 6636 -4516 6734 -4494
rect 6636 -4562 6662 -4516
rect 6708 -4562 6734 -4516
rect 6636 -4610 6734 -4562
rect 6636 -4656 6662 -4610
rect 6708 -4656 6734 -4610
rect 6636 -4704 6734 -4656
rect 6636 -4750 6662 -4704
rect 6708 -4750 6734 -4704
rect 6636 -4798 6734 -4750
rect 6636 -4844 6662 -4798
rect 6708 -4844 6734 -4798
rect 6636 -4892 6734 -4844
rect 8760 -4734 11112 -4708
rect 8760 -4780 8786 -4734
rect 8832 -4780 8884 -4734
rect 8930 -4780 8982 -4734
rect 9028 -4780 9080 -4734
rect 9126 -4780 9178 -4734
rect 9224 -4780 9276 -4734
rect 9322 -4780 9374 -4734
rect 9420 -4780 9472 -4734
rect 9518 -4780 9570 -4734
rect 9616 -4780 9668 -4734
rect 9714 -4780 9766 -4734
rect 9812 -4780 9864 -4734
rect 9910 -4780 9962 -4734
rect 10008 -4780 10060 -4734
rect 10106 -4780 10158 -4734
rect 10204 -4780 10256 -4734
rect 10302 -4780 10354 -4734
rect 10400 -4780 10452 -4734
rect 10498 -4780 10550 -4734
rect 10596 -4780 10648 -4734
rect 10694 -4780 10746 -4734
rect 10792 -4780 10844 -4734
rect 10890 -4780 10942 -4734
rect 10988 -4780 11040 -4734
rect 11086 -4780 11112 -4734
rect 8760 -4806 11112 -4780
rect 8760 -4832 8858 -4806
rect 8760 -4878 8786 -4832
rect 8832 -4878 8858 -4832
rect 8760 -4889 8858 -4878
rect 6636 -4938 6662 -4892
rect 6708 -4938 6734 -4892
rect 6636 -4986 6734 -4938
rect 6636 -5032 6662 -4986
rect 6708 -5032 6734 -4986
rect 6636 -5080 6734 -5032
rect 6636 -5126 6662 -5080
rect 6708 -5126 6734 -5080
rect 6636 -5174 6734 -5126
rect 6636 -5220 6662 -5174
rect 6708 -5220 6734 -5174
rect 6636 -5268 6734 -5220
rect 6636 -5314 6662 -5268
rect 6708 -5314 6734 -5268
rect 6636 -5362 6734 -5314
rect 6636 -5408 6662 -5362
rect 6708 -5408 6734 -5362
rect 6636 -5456 6734 -5408
rect 6636 -5502 6662 -5456
rect 6708 -5502 6734 -5456
rect 6636 -5550 6734 -5502
rect 6636 -5596 6662 -5550
rect 6708 -5596 6734 -5550
rect 6636 -5644 6734 -5596
rect 6636 -5690 6662 -5644
rect 6708 -5690 6734 -5644
rect 6636 -5738 6734 -5690
rect 6636 -5784 6662 -5738
rect 6708 -5784 6734 -5738
rect 6636 -5832 6734 -5784
rect 6636 -5878 6662 -5832
rect 6708 -5878 6734 -5832
rect 6636 -5926 6734 -5878
rect 6636 -5972 6662 -5926
rect 6708 -5972 6734 -5926
rect 6636 -5994 6734 -5972
rect 3665 -6011 6734 -5994
rect 3665 -6057 3691 -6011
rect 3737 -6020 6734 -6011
rect 3737 -6057 4029 -6020
rect 3665 -6065 4029 -6057
rect 3665 -6105 3763 -6065
rect 4002 -6066 4029 -6065
rect 4075 -6066 4123 -6020
rect 4169 -6066 4217 -6020
rect 4263 -6066 4311 -6020
rect 4357 -6066 4405 -6020
rect 4451 -6066 4499 -6020
rect 4545 -6066 4593 -6020
rect 4639 -6066 4687 -6020
rect 4733 -6066 4781 -6020
rect 4827 -6066 4875 -6020
rect 4921 -6066 4969 -6020
rect 5015 -6066 5063 -6020
rect 5109 -6066 5157 -6020
rect 5203 -6066 5251 -6020
rect 5297 -6066 5345 -6020
rect 5391 -6066 5439 -6020
rect 5485 -6066 5533 -6020
rect 5579 -6066 5627 -6020
rect 5673 -6066 5721 -6020
rect 5767 -6066 5815 -6020
rect 5861 -6066 5909 -6020
rect 5955 -6066 6003 -6020
rect 6049 -6066 6097 -6020
rect 6143 -6066 6191 -6020
rect 6237 -6066 6285 -6020
rect 6331 -6066 6379 -6020
rect 6425 -6066 6473 -6020
rect 6519 -6066 6567 -6020
rect 6613 -6066 6661 -6020
rect 6707 -6066 6734 -6020
rect 4002 -6092 6734 -6066
rect 8298 -4930 8858 -4889
rect 8298 -4976 8786 -4930
rect 8832 -4976 8858 -4930
rect 8298 -5028 8858 -4976
rect 8298 -5074 8786 -5028
rect 8832 -5074 8858 -5028
rect 8298 -5126 8858 -5074
rect 8298 -5153 8786 -5126
rect 8298 -5431 8562 -5153
rect 8760 -5172 8786 -5153
rect 8832 -5172 8858 -5126
rect 8760 -5224 8858 -5172
rect 8760 -5270 8786 -5224
rect 8832 -5270 8858 -5224
rect 8760 -5322 8858 -5270
rect 8760 -5368 8786 -5322
rect 8832 -5368 8858 -5322
rect 8760 -5420 8858 -5368
rect 8760 -5431 8786 -5420
rect 8298 -5466 8786 -5431
rect 8832 -5466 8858 -5420
rect 8298 -5518 8858 -5466
rect 8298 -5564 8786 -5518
rect 8832 -5564 8858 -5518
rect 8298 -5616 8858 -5564
rect 8298 -5662 8786 -5616
rect 8832 -5662 8858 -5616
rect 8298 -5695 8858 -5662
rect 8298 -5889 8562 -5695
rect 8760 -5714 8858 -5695
rect 8760 -5760 8786 -5714
rect 8832 -5760 8858 -5714
rect 8760 -5812 8858 -5760
rect 8760 -5858 8786 -5812
rect 8832 -5858 8858 -5812
rect 8760 -5889 8858 -5858
rect 8298 -5910 8858 -5889
rect 8298 -5956 8786 -5910
rect 8832 -5956 8858 -5910
rect 8298 -6008 8858 -5956
rect 8298 -6054 8786 -6008
rect 8832 -6054 8858 -6008
rect 3665 -6151 3691 -6105
rect 3737 -6151 3763 -6105
rect 3665 -6173 3763 -6151
rect 1595 -6199 3763 -6173
rect 1595 -6245 1622 -6199
rect 1668 -6245 1716 -6199
rect 1762 -6245 1810 -6199
rect 1856 -6245 1904 -6199
rect 1950 -6245 1998 -6199
rect 2044 -6245 2092 -6199
rect 2138 -6245 2186 -6199
rect 2232 -6245 2280 -6199
rect 2326 -6245 2374 -6199
rect 2420 -6245 2468 -6199
rect 2514 -6245 2562 -6199
rect 2608 -6245 2656 -6199
rect 2702 -6245 2750 -6199
rect 2796 -6245 2844 -6199
rect 2890 -6245 2938 -6199
rect 2984 -6245 3032 -6199
rect 3078 -6245 3126 -6199
rect 3172 -6245 3220 -6199
rect 3266 -6245 3314 -6199
rect 3360 -6245 3408 -6199
rect 3454 -6245 3502 -6199
rect 3548 -6245 3596 -6199
rect 3642 -6245 3690 -6199
rect 3736 -6245 3763 -6199
rect 1595 -6271 3763 -6245
rect 8298 -6106 8858 -6054
rect 8298 -6152 8786 -6106
rect 8832 -6152 8858 -6106
rect 8298 -6153 8858 -6152
rect -1246 -6289 1304 -6282
rect -1246 -6306 -1219 -6289
rect -3293 -6332 -1219 -6306
rect -488 -6308 1304 -6289
rect 8298 -6317 8562 -6153
rect 8760 -6204 8858 -6153
rect 8760 -6250 8786 -6204
rect 8832 -6250 8858 -6204
rect 8760 -6302 8858 -6250
rect 8760 -6317 8786 -6302
rect 8298 -6348 8786 -6317
rect 8832 -6348 8858 -6302
rect 8298 -6400 8858 -6348
rect -2030 -6460 -1881 -6426
rect -2030 -6550 -2004 -6460
rect -1908 -6550 -1881 -6460
rect 8298 -6446 8786 -6400
rect 8832 -6446 8858 -6400
rect -2631 -6585 -2482 -6551
rect -2030 -6579 -1881 -6550
rect -574 -6512 1287 -6487
rect -574 -6558 -549 -6512
rect -503 -6558 -451 -6512
rect -405 -6558 -353 -6512
rect -307 -6558 -255 -6512
rect -209 -6558 -157 -6512
rect -111 -6558 -59 -6512
rect -13 -6558 39 -6512
rect 85 -6558 137 -6512
rect 183 -6558 235 -6512
rect 281 -6558 333 -6512
rect 379 -6558 431 -6512
rect 477 -6558 529 -6512
rect 575 -6558 627 -6512
rect 673 -6558 725 -6512
rect 771 -6558 823 -6512
rect 869 -6558 921 -6512
rect 967 -6558 1019 -6512
rect 1065 -6558 1117 -6512
rect 1163 -6558 1215 -6512
rect 1261 -6558 1287 -6512
rect 8298 -6498 8858 -6446
rect -574 -6566 1287 -6558
rect 1587 -6562 4134 -6537
rect 1587 -6566 1612 -6562
rect -2631 -6675 -2605 -6585
rect -2509 -6675 -2482 -6585
rect -2631 -6705 -2482 -6675
rect -574 -6584 1612 -6566
rect -574 -6610 -477 -6584
rect -574 -6656 -549 -6610
rect -503 -6656 -477 -6610
rect -574 -6708 -477 -6656
rect -574 -6754 -549 -6708
rect -503 -6754 -477 -6708
rect 1190 -6608 1612 -6584
rect 1658 -6608 1710 -6562
rect 1756 -6608 1808 -6562
rect 1854 -6608 1906 -6562
rect 1952 -6608 2004 -6562
rect 2050 -6608 2102 -6562
rect 2148 -6608 2200 -6562
rect 2246 -6608 2298 -6562
rect 2344 -6608 2396 -6562
rect 2442 -6608 2494 -6562
rect 2540 -6608 2592 -6562
rect 2638 -6608 2690 -6562
rect 2736 -6608 2788 -6562
rect 2834 -6608 2886 -6562
rect 2932 -6608 2984 -6562
rect 3030 -6608 3082 -6562
rect 3128 -6608 3180 -6562
rect 3226 -6608 3278 -6562
rect 3324 -6608 3376 -6562
rect 3422 -6608 3474 -6562
rect 3520 -6608 3572 -6562
rect 3618 -6608 3670 -6562
rect 3716 -6608 3768 -6562
rect 3814 -6608 3866 -6562
rect 3912 -6608 3964 -6562
rect 4010 -6608 4062 -6562
rect 4108 -6608 4134 -6562
rect 1190 -6610 4134 -6608
rect 1190 -6656 1215 -6610
rect 1261 -6634 4134 -6610
rect 1261 -6656 1684 -6634
rect 1190 -6660 1684 -6656
rect 1190 -6706 1612 -6660
rect 1658 -6706 1684 -6660
rect 1190 -6708 1684 -6706
rect -574 -6806 -477 -6754
rect -3321 -6842 -1166 -6816
rect -3321 -6888 -3295 -6842
rect -3249 -6888 -3197 -6842
rect -3151 -6888 -3099 -6842
rect -3053 -6888 -3001 -6842
rect -2955 -6888 -2903 -6842
rect -2857 -6888 -2805 -6842
rect -2759 -6888 -2707 -6842
rect -2661 -6888 -2609 -6842
rect -2563 -6888 -2511 -6842
rect -2465 -6888 -2413 -6842
rect -2367 -6888 -2315 -6842
rect -2269 -6888 -2217 -6842
rect -2171 -6888 -2119 -6842
rect -2073 -6888 -2021 -6842
rect -1975 -6888 -1923 -6842
rect -1877 -6888 -1825 -6842
rect -1779 -6888 -1727 -6842
rect -1681 -6888 -1629 -6842
rect -1583 -6888 -1531 -6842
rect -1485 -6888 -1433 -6842
rect -1387 -6888 -1335 -6842
rect -1289 -6888 -1237 -6842
rect -1191 -6888 -1166 -6842
rect -3321 -6914 -1166 -6888
rect -3321 -6940 -3223 -6914
rect -3321 -6986 -3295 -6940
rect -3249 -6986 -3223 -6940
rect -3321 -7038 -3223 -6986
rect -3321 -7084 -3295 -7038
rect -3249 -7084 -3223 -7038
rect -3321 -7136 -3223 -7084
rect -3060 -7053 -2992 -7040
rect -3060 -7099 -3049 -7053
rect -3003 -7099 -2992 -7053
rect -3060 -7107 -2992 -7099
rect -3321 -7182 -3295 -7136
rect -3249 -7182 -3223 -7136
rect -3049 -7141 -3003 -7107
rect -3321 -7234 -3223 -7182
rect -3321 -7280 -3295 -7234
rect -3249 -7280 -3223 -7234
rect -3321 -7332 -3223 -7280
rect -3076 -7212 -2979 -7199
rect -3076 -7293 -3061 -7212
rect -2993 -7293 -2979 -7212
rect -3076 -7306 -2979 -7293
rect -2912 -7211 -2815 -7198
rect -2912 -7292 -2897 -7211
rect -2829 -7292 -2815 -7211
rect -2912 -7305 -2815 -7292
rect -3321 -7378 -3295 -7332
rect -3249 -7378 -3223 -7332
rect -3321 -7430 -3223 -7378
rect -3321 -7476 -3295 -7430
rect -3249 -7476 -3223 -7430
rect -3321 -7528 -3223 -7476
rect -3321 -7574 -3295 -7528
rect -3249 -7574 -3223 -7528
rect -3321 -7626 -3223 -7574
rect -3321 -7672 -3295 -7626
rect -3249 -7672 -3223 -7626
rect -3321 -7724 -3223 -7672
rect -3321 -7770 -3295 -7724
rect -3249 -7770 -3223 -7724
rect -3321 -7822 -3223 -7770
rect -3321 -7868 -3295 -7822
rect -3249 -7868 -3223 -7822
rect -3321 -7920 -3223 -7868
rect -3060 -7853 -2992 -7840
rect -3060 -7899 -3049 -7853
rect -3003 -7899 -2992 -7853
rect -3060 -7907 -2992 -7899
rect -3321 -7966 -3295 -7920
rect -3249 -7966 -3223 -7920
rect -3049 -7941 -3003 -7907
rect -3321 -8018 -3223 -7966
rect -3321 -8064 -3295 -8018
rect -3249 -8064 -3223 -8018
rect -3321 -8116 -3223 -8064
rect -3075 -8018 -2978 -8005
rect -3075 -8099 -3060 -8018
rect -2992 -8099 -2978 -8018
rect -3075 -8112 -2978 -8099
rect -2915 -8022 -2818 -8007
rect -2915 -8103 -2901 -8022
rect -2833 -8103 -2818 -8022
rect -2915 -8115 -2818 -8103
rect -3321 -8162 -3295 -8116
rect -3249 -8162 -3223 -8116
rect -3321 -8214 -3223 -8162
rect -3321 -8260 -3295 -8214
rect -3249 -8260 -3223 -8214
rect -3321 -8312 -3223 -8260
rect -3321 -8358 -3295 -8312
rect -3249 -8358 -3223 -8312
rect -3321 -8410 -3223 -8358
rect -3321 -8456 -3295 -8410
rect -3249 -8456 -3223 -8410
rect -3321 -8508 -3223 -8456
rect -3321 -8554 -3295 -8508
rect -3249 -8554 -3223 -8508
rect -3321 -8606 -3223 -8554
rect -3321 -8652 -3295 -8606
rect -3249 -8652 -3223 -8606
rect -3321 -8704 -3223 -8652
rect -3321 -8750 -3295 -8704
rect -3249 -8750 -3223 -8704
rect -3060 -8651 -2992 -8638
rect -3060 -8697 -3049 -8651
rect -3003 -8697 -2992 -8651
rect -3060 -8705 -2992 -8697
rect -3049 -8750 -3003 -8705
rect -2889 -8750 -2843 -8739
rect -3321 -8802 -3223 -8750
rect -3321 -8848 -3295 -8802
rect -3249 -8848 -3223 -8802
rect -3321 -8900 -3223 -8848
rect -3321 -8946 -3295 -8900
rect -3249 -8946 -3223 -8900
rect -3077 -8818 -2980 -8805
rect -3077 -8899 -3062 -8818
rect -2994 -8899 -2980 -8818
rect -3077 -8912 -2980 -8899
rect -2918 -8818 -2821 -8805
rect -2918 -8899 -2903 -8818
rect -2835 -8899 -2821 -8818
rect -2918 -8912 -2821 -8899
rect -3321 -8998 -3223 -8946
rect -3321 -9044 -3295 -8998
rect -3249 -9044 -3223 -8998
rect -3321 -9096 -3223 -9044
rect -3321 -9142 -3295 -9096
rect -3249 -9142 -3223 -9096
rect -3321 -9194 -3223 -9142
rect -3321 -9240 -3295 -9194
rect -3249 -9240 -3223 -9194
rect -3321 -9292 -3223 -9240
rect -3321 -9338 -3295 -9292
rect -3249 -9338 -3223 -9292
rect -3049 -9335 -3003 -9324
rect -2889 -9335 -2843 -9324
rect -3321 -9390 -3223 -9338
rect -3321 -9436 -3295 -9390
rect -3249 -9436 -3223 -9390
rect -3321 -9488 -3223 -9436
rect -3321 -9534 -3295 -9488
rect -3249 -9534 -3223 -9488
rect -3060 -9451 -2992 -9438
rect -3060 -9497 -3049 -9451
rect -3003 -9497 -2992 -9451
rect -3060 -9505 -2992 -9497
rect -3321 -9586 -3223 -9534
rect -3049 -9550 -3003 -9505
rect -2889 -9550 -2843 -9539
rect -3321 -9632 -3295 -9586
rect -3249 -9632 -3223 -9586
rect -3321 -9684 -3223 -9632
rect -3321 -9730 -3295 -9684
rect -3249 -9730 -3223 -9684
rect -3075 -9616 -2978 -9603
rect -3075 -9697 -3060 -9616
rect -2992 -9697 -2978 -9616
rect -3075 -9710 -2978 -9697
rect -2913 -9615 -2816 -9602
rect -2913 -9696 -2898 -9615
rect -2830 -9696 -2816 -9615
rect -2913 -9709 -2816 -9696
rect -3321 -9782 -3223 -9730
rect -3321 -9828 -3295 -9782
rect -3249 -9828 -3223 -9782
rect -3321 -9880 -3223 -9828
rect -3321 -9926 -3295 -9880
rect -3249 -9926 -3223 -9880
rect -3321 -9978 -3223 -9926
rect -3321 -10024 -3295 -9978
rect -3249 -10024 -3223 -9978
rect -3321 -10076 -3223 -10024
rect -3321 -10122 -3295 -10076
rect -3249 -10122 -3223 -10076
rect -3321 -10174 -3223 -10122
rect -3049 -10135 -3003 -10124
rect -2889 -10135 -2843 -10124
rect -3321 -10220 -3295 -10174
rect -3249 -10220 -3223 -10174
rect -3321 -10272 -3223 -10220
rect -3321 -10318 -3295 -10272
rect -3249 -10318 -3223 -10272
rect -3321 -10344 -3223 -10318
rect -2731 -10344 -2681 -6914
rect -2597 -7531 -2500 -7518
rect -2597 -7612 -2582 -7531
rect -2514 -7612 -2500 -7531
rect -2597 -7625 -2500 -7612
rect -2605 -8332 -2491 -8316
rect -2605 -8414 -2589 -8332
rect -2507 -8414 -2491 -8332
rect -2605 -8428 -2491 -8414
rect -2569 -8750 -2523 -8739
rect -2607 -9133 -2493 -9117
rect -2607 -9215 -2591 -9133
rect -2509 -9215 -2493 -9133
rect -2607 -9229 -2493 -9215
rect -2569 -9335 -2523 -9324
rect -2569 -9550 -2523 -9539
rect -2596 -9931 -2499 -9918
rect -2596 -10012 -2581 -9931
rect -2513 -10012 -2499 -9931
rect -2596 -10025 -2499 -10012
rect -2569 -10135 -2523 -10124
rect -2411 -10344 -2361 -6914
rect -2249 -7152 -2203 -7141
rect -2274 -7212 -2177 -7199
rect -2274 -7293 -2259 -7212
rect -2191 -7293 -2177 -7212
rect -2274 -7306 -2177 -7293
rect -2249 -7737 -2203 -7726
rect -2268 -7809 -2184 -7797
rect -2268 -7869 -2256 -7809
rect -2196 -7869 -2184 -7809
rect -2268 -7881 -2184 -7869
rect -2249 -7952 -2203 -7941
rect -2273 -8016 -2176 -8003
rect -2273 -8097 -2258 -8016
rect -2190 -8097 -2176 -8016
rect -2273 -8110 -2176 -8097
rect -2249 -8537 -2203 -8526
rect -2268 -8610 -2184 -8598
rect -2268 -8670 -2256 -8610
rect -2196 -8670 -2184 -8610
rect -2268 -8682 -2184 -8670
rect -2249 -8750 -2203 -8739
rect -2276 -8816 -2179 -8803
rect -2276 -8897 -2261 -8816
rect -2193 -8897 -2179 -8816
rect -2276 -8910 -2179 -8897
rect -2249 -9335 -2203 -9324
rect -2269 -9410 -2185 -9398
rect -2269 -9470 -2257 -9410
rect -2197 -9470 -2185 -9410
rect -2269 -9482 -2185 -9470
rect -2249 -9550 -2203 -9539
rect -2275 -9616 -2178 -9603
rect -2275 -9697 -2260 -9616
rect -2192 -9697 -2178 -9616
rect -2275 -9710 -2178 -9697
rect -2249 -10135 -2203 -10124
rect -2091 -10344 -2041 -6914
rect -1929 -7152 -1883 -7141
rect -1965 -7530 -1851 -7514
rect -1965 -7612 -1949 -7530
rect -1867 -7612 -1851 -7530
rect -1965 -7626 -1851 -7612
rect -1929 -7737 -1883 -7726
rect -1929 -7952 -1883 -7941
rect -1955 -8327 -1858 -8314
rect -1955 -8408 -1940 -8327
rect -1872 -8408 -1858 -8327
rect -1955 -8421 -1858 -8408
rect -1929 -8537 -1883 -8526
rect -1929 -8750 -1883 -8739
rect -1955 -9128 -1858 -9115
rect -1955 -9209 -1940 -9128
rect -1872 -9209 -1858 -9128
rect -1955 -9222 -1858 -9209
rect -1929 -9335 -1883 -9324
rect -1929 -9550 -1883 -9539
rect -1963 -9931 -1849 -9915
rect -1963 -10013 -1947 -9931
rect -1865 -10013 -1849 -9931
rect -1963 -10027 -1849 -10013
rect -1929 -10135 -1883 -10124
rect -1771 -10344 -1721 -6914
rect -1263 -6920 -1166 -6914
rect -574 -6852 -549 -6806
rect -503 -6852 -477 -6806
rect -574 -6904 -477 -6852
rect -164 -6760 844 -6714
rect -164 -6863 -118 -6760
rect 127 -6824 229 -6811
rect 127 -6829 143 -6824
rect -574 -6920 -549 -6904
rect -1263 -6940 -549 -6920
rect -1263 -6986 -1237 -6940
rect -1191 -6950 -549 -6940
rect -503 -6950 -477 -6904
rect -1191 -6986 -477 -6950
rect -1263 -7002 -477 -6986
rect -324 -6909 -245 -6863
rect -199 -6909 -118 -6863
rect -324 -6990 -278 -6909
rect -323 -7001 -278 -6990
rect -164 -6992 -118 -6909
rect -4 -6875 143 -6829
rect -4 -6984 42 -6875
rect 127 -6880 143 -6875
rect 215 -6829 229 -6824
rect 215 -6875 684 -6829
rect 215 -6880 229 -6875
rect 127 -6894 229 -6880
rect 638 -6984 684 -6875
rect 798 -6885 844 -6760
rect 1190 -6754 1215 -6708
rect 1261 -6754 1684 -6708
rect 1190 -6756 1684 -6754
rect 1190 -6766 1612 -6756
rect 1190 -6806 1287 -6766
rect 1190 -6852 1215 -6806
rect 1261 -6852 1287 -6806
rect 798 -6931 878 -6885
rect 924 -6931 1004 -6885
rect 798 -6992 844 -6931
rect 958 -6988 1004 -6931
rect 960 -6997 1004 -6988
rect 1190 -6904 1287 -6852
rect 1190 -6950 1215 -6904
rect 1261 -6950 1287 -6904
rect 1190 -6966 1287 -6950
rect 1381 -6966 1496 -6766
rect 1587 -6802 1612 -6766
rect 1658 -6802 1684 -6756
rect 1587 -6854 1684 -6802
rect 1587 -6900 1612 -6854
rect 1658 -6900 1684 -6854
rect 1587 -6952 1684 -6900
rect 1587 -6966 1612 -6952
rect 1190 -6998 1612 -6966
rect 1658 -6998 1684 -6952
rect -1263 -7038 -549 -7002
rect -1460 -7053 -1392 -7040
rect -1460 -7099 -1449 -7053
rect -1403 -7099 -1392 -7053
rect -1460 -7107 -1392 -7099
rect -1263 -7084 -1237 -7038
rect -1191 -7048 -549 -7038
rect -503 -7048 -477 -7002
rect 1190 -7002 1684 -6998
rect -1191 -7084 -477 -7048
rect -1263 -7100 -477 -7084
rect -1609 -7152 -1563 -7141
rect -1449 -7152 -1403 -7107
rect -1263 -7120 -549 -7100
rect -1263 -7136 -1166 -7120
rect -1263 -7182 -1237 -7136
rect -1191 -7182 -1166 -7136
rect -1638 -7212 -1541 -7199
rect -1638 -7293 -1623 -7212
rect -1555 -7293 -1541 -7212
rect -1638 -7306 -1541 -7293
rect -1475 -7216 -1378 -7203
rect -1475 -7297 -1460 -7216
rect -1392 -7297 -1378 -7216
rect -1475 -7310 -1378 -7297
rect -1263 -7234 -1166 -7182
rect -1263 -7280 -1237 -7234
rect -1191 -7280 -1166 -7234
rect -1263 -7320 -1166 -7280
rect -1011 -7320 -765 -7120
rect -574 -7146 -549 -7120
rect -503 -7146 -477 -7100
rect -184 -7047 -99 -7032
rect -184 -7129 -169 -7047
rect -113 -7129 -99 -7047
rect -184 -7142 -99 -7129
rect 1190 -7048 1215 -7002
rect 1261 -7048 1684 -7002
rect 1190 -7050 1684 -7048
rect 1190 -7096 1612 -7050
rect 1658 -7096 1684 -7050
rect 1190 -7100 1684 -7096
rect -574 -7198 -477 -7146
rect -574 -7244 -549 -7198
rect -503 -7244 -477 -7198
rect 1190 -7146 1215 -7100
rect 1261 -7146 1684 -7100
rect 1190 -7148 1684 -7146
rect 1190 -7166 1612 -7148
rect 1190 -7198 1287 -7166
rect -574 -7296 -477 -7244
rect -574 -7320 -549 -7296
rect -1263 -7332 -549 -7320
rect -1263 -7378 -1237 -7332
rect -1191 -7342 -549 -7332
rect -503 -7342 -477 -7296
rect -185 -7232 -99 -7214
rect -185 -7314 -170 -7232
rect -114 -7314 -99 -7232
rect 298 -7215 381 -7199
rect 298 -7287 312 -7215
rect 368 -7287 381 -7215
rect 298 -7301 381 -7287
rect 1190 -7244 1215 -7198
rect 1261 -7244 1287 -7198
rect 1190 -7296 1287 -7244
rect -185 -7330 -99 -7314
rect -1191 -7378 -477 -7342
rect -1263 -7394 -477 -7378
rect -1263 -7430 -549 -7394
rect -1263 -7476 -1237 -7430
rect -1191 -7440 -549 -7430
rect -503 -7440 -477 -7394
rect -1191 -7476 -477 -7440
rect -1263 -7492 -477 -7476
rect -1263 -7520 -549 -7492
rect -1263 -7528 -1166 -7520
rect -1263 -7574 -1237 -7528
rect -1191 -7574 -1166 -7528
rect -1263 -7626 -1166 -7574
rect -1263 -7672 -1237 -7626
rect -1191 -7672 -1166 -7626
rect -1263 -7720 -1166 -7672
rect -1011 -7720 -765 -7520
rect -574 -7538 -549 -7520
rect -503 -7538 -477 -7492
rect -574 -7590 -477 -7538
rect 1190 -7342 1215 -7296
rect 1261 -7342 1287 -7296
rect 1190 -7366 1287 -7342
rect 1381 -7366 1496 -7166
rect 1587 -7194 1612 -7166
rect 1658 -7194 1684 -7148
rect 1587 -7246 1684 -7194
rect 1587 -7292 1612 -7246
rect 1658 -7292 1684 -7246
rect 1587 -7344 1684 -7292
rect 1587 -7366 1612 -7344
rect 1190 -7390 1612 -7366
rect 1658 -7390 1684 -7344
rect 1190 -7394 1684 -7390
rect 1190 -7440 1215 -7394
rect 1261 -7440 1684 -7394
rect 1190 -7442 1684 -7440
rect 1190 -7488 1612 -7442
rect 1658 -7488 1684 -7442
rect 1190 -7492 1684 -7488
rect 1190 -7538 1215 -7492
rect 1261 -7538 1684 -7492
rect 1190 -7540 1684 -7538
rect 1190 -7566 1612 -7540
rect -574 -7636 -549 -7590
rect -503 -7636 -477 -7590
rect -574 -7688 -477 -7636
rect -574 -7720 -549 -7688
rect -1263 -7724 -549 -7720
rect -1609 -7737 -1563 -7726
rect -1449 -7737 -1403 -7726
rect -1263 -7770 -1237 -7724
rect -1191 -7734 -549 -7724
rect -503 -7734 -477 -7688
rect 157 -7693 203 -7579
rect -1191 -7770 -477 -7734
rect -1263 -7786 -477 -7770
rect -1263 -7822 -549 -7786
rect -1460 -7853 -1392 -7840
rect -1460 -7899 -1449 -7853
rect -1403 -7899 -1392 -7853
rect -1460 -7907 -1392 -7899
rect -1263 -7868 -1237 -7822
rect -1191 -7832 -549 -7822
rect -503 -7832 -477 -7786
rect -1191 -7868 -477 -7832
rect -324 -7771 -243 -7725
rect -197 -7771 -118 -7725
rect -324 -7835 -278 -7771
rect -164 -7839 -118 -7771
rect -4 -7739 203 -7693
rect 297 -7677 387 -7665
rect -1263 -7884 -477 -7868
rect -1609 -7952 -1563 -7941
rect -1449 -7952 -1403 -7907
rect -1263 -7920 -549 -7884
rect -1263 -7966 -1237 -7920
rect -1191 -7966 -1166 -7920
rect -1636 -8015 -1539 -8002
rect -1636 -8096 -1621 -8015
rect -1553 -8096 -1539 -8015
rect -1636 -8109 -1539 -8096
rect -1473 -8015 -1376 -8002
rect -1473 -8096 -1458 -8015
rect -1390 -8096 -1376 -8015
rect -1473 -8109 -1376 -8096
rect -1263 -8018 -1166 -7966
rect -1263 -8064 -1237 -8018
rect -1191 -8064 -1166 -8018
rect -1263 -8116 -1166 -8064
rect -1263 -8162 -1237 -8116
rect -1191 -8120 -1166 -8116
rect -1011 -8120 -765 -7920
rect -574 -7930 -549 -7920
rect -503 -7930 -477 -7884
rect -574 -7982 -477 -7930
rect -574 -8028 -549 -7982
rect -503 -8028 -477 -7982
rect -574 -8080 -477 -8028
rect -574 -8120 -549 -8080
rect -1191 -8126 -549 -8120
rect -503 -8126 -477 -8080
rect -1191 -8162 -477 -8126
rect -1263 -8178 -477 -8162
rect -1263 -8214 -549 -8178
rect -1263 -8260 -1237 -8214
rect -1191 -8224 -549 -8214
rect -503 -8224 -477 -8178
rect -1191 -8260 -477 -8224
rect -1263 -8276 -477 -8260
rect -1263 -8312 -549 -8276
rect -1263 -8358 -1237 -8312
rect -1191 -8320 -549 -8312
rect -1191 -8358 -1166 -8320
rect -1263 -8410 -1166 -8358
rect -1263 -8456 -1237 -8410
rect -1191 -8456 -1166 -8410
rect -1263 -8508 -1166 -8456
rect -1609 -8537 -1563 -8526
rect -1449 -8537 -1403 -8526
rect -1263 -8554 -1237 -8508
rect -1191 -8520 -1166 -8508
rect -1011 -8520 -765 -8320
rect -574 -8322 -549 -8320
rect -503 -8322 -477 -8276
rect -164 -8279 -118 -8188
rect -574 -8374 -477 -8322
rect -574 -8420 -549 -8374
rect -503 -8420 -477 -8374
rect -183 -8295 -100 -8279
rect -183 -8367 -169 -8295
rect -113 -8367 -100 -8295
rect -183 -8381 -100 -8367
rect -574 -8472 -477 -8420
rect -574 -8518 -549 -8472
rect -503 -8518 -477 -8472
rect -574 -8520 -477 -8518
rect -1191 -8554 -477 -8520
rect -1263 -8570 -477 -8554
rect -1263 -8606 -549 -8570
rect -1460 -8651 -1392 -8638
rect -1460 -8697 -1449 -8651
rect -1403 -8697 -1392 -8651
rect -1460 -8705 -1392 -8697
rect -1263 -8652 -1237 -8606
rect -1191 -8616 -549 -8606
rect -503 -8616 -477 -8570
rect -1191 -8652 -477 -8616
rect -1263 -8668 -477 -8652
rect -1263 -8704 -549 -8668
rect -1609 -8750 -1563 -8739
rect -1449 -8750 -1403 -8705
rect -1263 -8750 -1237 -8704
rect -1191 -8714 -549 -8704
rect -503 -8714 -477 -8668
rect -1191 -8720 -477 -8714
rect -1191 -8750 -1166 -8720
rect -1263 -8802 -1166 -8750
rect -1637 -8816 -1540 -8803
rect -1637 -8897 -1622 -8816
rect -1554 -8897 -1540 -8816
rect -1637 -8910 -1540 -8897
rect -1475 -8815 -1378 -8802
rect -1475 -8896 -1460 -8815
rect -1392 -8896 -1378 -8815
rect -1475 -8909 -1378 -8896
rect -1263 -8848 -1237 -8802
rect -1191 -8848 -1166 -8802
rect -1263 -8900 -1166 -8848
rect -1263 -8946 -1237 -8900
rect -1191 -8920 -1166 -8900
rect -1011 -8920 -765 -8720
rect -574 -8766 -477 -8720
rect -574 -8812 -549 -8766
rect -503 -8812 -477 -8766
rect -574 -8864 -477 -8812
rect -574 -8910 -549 -8864
rect -503 -8910 -477 -8864
rect -164 -8879 -118 -8381
rect -4 -8645 42 -7739
rect 297 -7743 309 -7677
rect 375 -7743 387 -7677
rect 477 -7693 523 -7569
rect 1190 -7590 1287 -7566
rect 1190 -7636 1215 -7590
rect 1261 -7636 1287 -7590
rect 1190 -7688 1287 -7636
rect 477 -7739 684 -7693
rect 297 -7755 387 -7743
rect 157 -7897 203 -7834
rect 139 -7913 222 -7897
rect 139 -7985 153 -7913
rect 209 -7985 222 -7913
rect 317 -7977 363 -7834
rect 139 -7999 222 -7985
rect 292 -7995 389 -7977
rect 157 -8489 203 -7999
rect 292 -8059 309 -7995
rect 373 -8059 389 -7995
rect 292 -8079 389 -8059
rect 289 -8111 389 -8079
rect 289 -8140 309 -8111
rect 292 -8175 309 -8140
rect 373 -8175 389 -8111
rect 292 -8189 389 -8175
rect 317 -8410 363 -8189
rect 477 -8488 523 -7834
rect 134 -8505 217 -8489
rect 134 -8577 148 -8505
rect 204 -8577 217 -8505
rect 134 -8591 217 -8577
rect 460 -8504 543 -8488
rect 460 -8576 474 -8504
rect 530 -8576 543 -8504
rect 460 -8590 543 -8576
rect -23 -8661 60 -8645
rect -23 -8733 -9 -8661
rect 47 -8733 60 -8661
rect -23 -8747 60 -8733
rect -574 -8920 -477 -8910
rect -1191 -8946 -477 -8920
rect -1263 -8962 -477 -8946
rect -1263 -8998 -549 -8962
rect -1263 -9044 -1237 -8998
rect -1191 -9008 -549 -8998
rect -503 -9008 -477 -8962
rect -1191 -9044 -477 -9008
rect -1263 -9060 -477 -9044
rect -1263 -9096 -549 -9060
rect -1263 -9142 -1237 -9096
rect -1191 -9106 -549 -9096
rect -503 -9106 -477 -9060
rect -1191 -9120 -477 -9106
rect -1191 -9142 -1166 -9120
rect -1263 -9194 -1166 -9142
rect -1263 -9240 -1237 -9194
rect -1191 -9240 -1166 -9194
rect -1263 -9292 -1166 -9240
rect -1609 -9335 -1563 -9324
rect -1449 -9335 -1403 -9324
rect -1263 -9338 -1237 -9292
rect -1191 -9320 -1166 -9292
rect -1011 -9320 -765 -9120
rect -574 -9158 -477 -9120
rect -574 -9204 -549 -9158
rect -503 -9204 -477 -9158
rect -574 -9256 -477 -9204
rect -574 -9302 -549 -9256
rect -503 -9302 -477 -9256
rect -574 -9320 -477 -9302
rect -1191 -9338 -477 -9320
rect -1263 -9354 -477 -9338
rect -1263 -9390 -549 -9354
rect -1263 -9436 -1237 -9390
rect -1191 -9400 -549 -9390
rect -503 -9400 -477 -9354
rect -1191 -9436 -477 -9400
rect -1460 -9451 -1392 -9438
rect -1460 -9497 -1449 -9451
rect -1403 -9497 -1392 -9451
rect -1460 -9505 -1392 -9497
rect -1263 -9452 -477 -9436
rect -1263 -9488 -549 -9452
rect -1609 -9550 -1563 -9539
rect -1449 -9550 -1403 -9505
rect -1263 -9534 -1237 -9488
rect -1191 -9498 -549 -9488
rect -503 -9498 -477 -9452
rect -1191 -9520 -477 -9498
rect -324 -9468 -278 -9410
rect -164 -9468 -118 -9228
rect -324 -9514 -243 -9468
rect -197 -9514 -118 -9468
rect -4 -9509 42 -8747
rect 157 -9410 203 -8591
rect 317 -8957 363 -8824
rect 290 -8975 390 -8957
rect 290 -9031 304 -8975
rect 376 -9031 390 -8975
rect 290 -9096 390 -9031
rect 288 -9098 390 -9096
rect 288 -9154 304 -9098
rect 376 -9154 390 -9098
rect 288 -9168 390 -9154
rect 317 -9410 363 -9168
rect 477 -9212 523 -8590
rect 638 -8645 684 -7739
rect 1190 -7734 1215 -7688
rect 1261 -7734 1287 -7688
rect 798 -7789 877 -7743
rect 923 -7789 1004 -7743
rect 798 -8141 844 -7789
rect 958 -7843 1004 -7789
rect 1190 -7786 1287 -7734
rect 1190 -7832 1215 -7786
rect 1261 -7832 1287 -7786
rect 1190 -7884 1287 -7832
rect 1190 -7930 1215 -7884
rect 1261 -7913 1287 -7884
rect 1381 -7913 1496 -7566
rect 1587 -7586 1612 -7566
rect 1658 -7586 1684 -7540
rect 1587 -7612 1684 -7586
rect 1749 -7399 1807 -6634
rect 1749 -7411 1906 -7399
rect 1749 -7469 1835 -7411
rect 1893 -7469 1906 -7411
rect 1749 -7481 1906 -7469
rect 1749 -7612 1807 -7481
rect 1965 -7612 2023 -6634
rect 2103 -6768 2330 -6751
rect 2103 -6774 2127 -6768
rect 2103 -6835 2113 -6774
rect 2187 -6828 2241 -6768
rect 2301 -6775 2330 -6768
rect 2174 -6835 2259 -6828
rect 2103 -6836 2259 -6835
rect 2320 -6836 2330 -6775
rect 2103 -6851 2330 -6836
rect 2181 -7325 2239 -6851
rect 2397 -7612 2455 -6634
rect 2611 -7430 2669 -6921
rect 2743 -7329 2801 -6634
rect 2860 -6749 3089 -6734
rect 2860 -6772 2882 -6749
rect 2860 -6830 2873 -6772
rect 2942 -6809 2996 -6749
rect 3056 -6773 3089 -6749
rect 2931 -6830 3010 -6809
rect 2860 -6831 3010 -6830
rect 3068 -6831 3089 -6773
rect 2860 -6842 3089 -6831
rect 2959 -6844 3089 -6842
rect 2959 -7326 3017 -6844
rect 3090 -7413 3148 -6921
rect 3025 -7428 3226 -7413
rect 3025 -7430 3039 -7428
rect 2611 -7488 3039 -7430
rect 3099 -7488 3153 -7428
rect 3213 -7488 3226 -7428
rect 3025 -7502 3226 -7488
rect 3305 -7612 3363 -6634
rect 3499 -7010 3596 -6992
rect 3499 -7074 3516 -7010
rect 3580 -7074 3596 -7010
rect 3499 -7126 3596 -7074
rect 3499 -7190 3516 -7126
rect 3580 -7190 3596 -7126
rect 3499 -7204 3596 -7190
rect 3655 -7612 3713 -6634
rect 3870 -7389 3928 -6634
rect 3771 -7401 3928 -7389
rect 3771 -7459 3784 -7401
rect 3842 -7459 3928 -7401
rect 3771 -7471 3928 -7459
rect 3870 -7612 3928 -7471
rect 4037 -6660 4134 -6634
rect 4037 -6706 4062 -6660
rect 4108 -6706 4134 -6660
rect 4037 -6756 4134 -6706
rect 8298 -6544 8786 -6498
rect 8832 -6544 8858 -6498
rect 8298 -6581 8858 -6544
rect 4037 -6802 4062 -6756
rect 4108 -6802 4134 -6756
rect 4037 -6854 4134 -6802
rect 4037 -6900 4062 -6854
rect 4108 -6900 4134 -6854
rect 4037 -6952 4134 -6900
rect 4037 -6998 4062 -6952
rect 4108 -6989 4134 -6952
rect 4374 -6765 8097 -6740
rect 4374 -6766 4497 -6765
rect 4374 -6812 4399 -6766
rect 4445 -6811 4497 -6766
rect 4543 -6811 4595 -6765
rect 4641 -6811 4693 -6765
rect 4739 -6811 4791 -6765
rect 4837 -6811 4889 -6765
rect 4935 -6811 4987 -6765
rect 5033 -6811 5085 -6765
rect 5131 -6811 5183 -6765
rect 5229 -6811 5281 -6765
rect 5327 -6811 5379 -6765
rect 5425 -6811 5477 -6765
rect 5523 -6811 5575 -6765
rect 5621 -6811 5673 -6765
rect 5719 -6811 5771 -6765
rect 5817 -6811 5869 -6765
rect 5915 -6811 5967 -6765
rect 6013 -6811 6065 -6765
rect 6111 -6811 6163 -6765
rect 6209 -6811 6261 -6765
rect 6307 -6811 6359 -6765
rect 6405 -6811 6457 -6765
rect 6503 -6811 6555 -6765
rect 6601 -6811 6653 -6765
rect 6699 -6811 6751 -6765
rect 6797 -6811 6849 -6765
rect 6895 -6811 6947 -6765
rect 6993 -6811 7045 -6765
rect 7091 -6811 7143 -6765
rect 7189 -6811 7241 -6765
rect 7287 -6811 7339 -6765
rect 7385 -6811 7437 -6765
rect 7483 -6811 7535 -6765
rect 7581 -6811 7633 -6765
rect 7679 -6811 7731 -6765
rect 7777 -6811 7829 -6765
rect 7875 -6811 7927 -6765
rect 7973 -6811 8025 -6765
rect 8071 -6780 8097 -6765
rect 8298 -6780 8562 -6581
rect 8760 -6596 8858 -6581
rect 8760 -6642 8786 -6596
rect 8832 -6642 8858 -6596
rect 8760 -6694 8858 -6642
rect 8760 -6740 8786 -6694
rect 8832 -6740 8858 -6694
rect 8760 -6780 8858 -6740
rect 8071 -6792 8858 -6780
rect 8071 -6811 8786 -6792
rect 4445 -6812 8786 -6811
rect 4374 -6837 8786 -6812
rect 4374 -6863 4471 -6837
rect 4374 -6909 4400 -6863
rect 4446 -6909 4471 -6863
rect 4374 -6961 4471 -6909
rect 4374 -6989 4400 -6961
rect 4108 -6998 4400 -6989
rect 4037 -7007 4400 -6998
rect 4446 -7007 4471 -6961
rect 4037 -7050 4471 -7007
rect 4037 -7096 4062 -7050
rect 4108 -7059 4471 -7050
rect 4108 -7096 4400 -7059
rect 4037 -7105 4400 -7096
rect 4446 -7105 4471 -7059
rect 4037 -7148 4471 -7105
rect 4037 -7194 4062 -7148
rect 4108 -7157 4471 -7148
rect 4108 -7189 4400 -7157
rect 4108 -7194 4134 -7189
rect 4037 -7246 4134 -7194
rect 4037 -7292 4062 -7246
rect 4108 -7292 4134 -7246
rect 4037 -7344 4134 -7292
rect 4037 -7390 4062 -7344
rect 4108 -7389 4134 -7344
rect 4374 -7203 4400 -7189
rect 4446 -7203 4471 -7157
rect 4374 -7255 4471 -7203
rect 4374 -7301 4400 -7255
rect 4446 -7301 4471 -7255
rect 4374 -7353 4471 -7301
rect 4374 -7389 4400 -7353
rect 4108 -7390 4400 -7389
rect 4037 -7399 4400 -7390
rect 4446 -7399 4471 -7353
rect 4037 -7442 4471 -7399
rect 4037 -7488 4062 -7442
rect 4108 -7451 4471 -7442
rect 4108 -7488 4400 -7451
rect 4037 -7497 4400 -7488
rect 4446 -7497 4471 -7451
rect 4037 -7540 4471 -7497
rect 4037 -7586 4062 -7540
rect 4108 -7549 4471 -7540
rect 4108 -7586 4400 -7549
rect 4037 -7589 4400 -7586
rect 4037 -7612 4134 -7589
rect 1587 -7638 4134 -7612
rect 1587 -7684 1612 -7638
rect 1658 -7684 1710 -7638
rect 1756 -7684 1808 -7638
rect 1854 -7684 1906 -7638
rect 1952 -7684 2004 -7638
rect 2050 -7684 2102 -7638
rect 2148 -7684 2200 -7638
rect 2246 -7684 2298 -7638
rect 2344 -7684 2396 -7638
rect 2442 -7684 2494 -7638
rect 2540 -7684 2592 -7638
rect 2638 -7684 2690 -7638
rect 2736 -7684 2788 -7638
rect 2834 -7684 2886 -7638
rect 2932 -7684 2984 -7638
rect 3030 -7684 3082 -7638
rect 3128 -7684 3180 -7638
rect 3226 -7684 3278 -7638
rect 3324 -7684 3376 -7638
rect 3422 -7684 3474 -7638
rect 3520 -7684 3572 -7638
rect 3618 -7684 3670 -7638
rect 3716 -7684 3768 -7638
rect 3814 -7684 3866 -7638
rect 3912 -7684 3964 -7638
rect 4010 -7684 4062 -7638
rect 4108 -7684 4134 -7638
rect 1587 -7709 4134 -7684
rect 4374 -7595 4400 -7589
rect 4446 -7595 4471 -7549
rect 4374 -7647 4471 -7595
rect 4374 -7693 4400 -7647
rect 4446 -7693 4471 -7647
rect 1659 -7913 1859 -7709
rect 2059 -7913 2259 -7709
rect 2459 -7913 2659 -7709
rect 2859 -7913 3059 -7709
rect 3259 -7913 3459 -7709
rect 3659 -7913 3859 -7709
rect 4374 -7745 4471 -7693
rect 4374 -7791 4400 -7745
rect 4446 -7791 4471 -7745
rect 4374 -7843 4471 -7791
rect 4374 -7889 4400 -7843
rect 4446 -7889 4471 -7843
rect 4374 -7913 4471 -7889
rect 1261 -7930 4471 -7913
rect 1190 -7941 4471 -7930
rect 1190 -7982 4400 -7941
rect 1190 -8028 1215 -7982
rect 1261 -7987 4400 -7982
rect 4446 -7987 4471 -7941
rect 1261 -8028 4471 -7987
rect 1190 -8039 4471 -8028
rect 1190 -8080 4400 -8039
rect 1190 -8126 1215 -8080
rect 1261 -8085 4400 -8080
rect 4446 -8085 4471 -8039
rect 1261 -8113 4471 -8085
rect 1261 -8126 1287 -8113
rect 778 -8157 863 -8141
rect 778 -8229 793 -8157
rect 849 -8229 863 -8157
rect 778 -8300 863 -8229
rect 778 -8372 793 -8300
rect 849 -8372 863 -8300
rect 778 -8387 863 -8372
rect 1190 -8178 1287 -8126
rect 1190 -8224 1215 -8178
rect 1261 -8224 1287 -8178
rect 1190 -8276 1287 -8224
rect 1190 -8322 1215 -8276
rect 1261 -8322 1287 -8276
rect 1190 -8374 1287 -8322
rect 620 -8661 703 -8645
rect 620 -8733 634 -8661
rect 690 -8733 703 -8661
rect 620 -8747 703 -8733
rect 457 -9228 540 -9212
rect 457 -9300 471 -9228
rect 527 -9300 540 -9228
rect 457 -9314 540 -9300
rect 477 -9410 523 -9314
rect 288 -9506 378 -9494
rect -1191 -9534 -1166 -9520
rect -1263 -9586 -1166 -9534
rect -1635 -9619 -1538 -9606
rect -1635 -9700 -1620 -9619
rect -1552 -9700 -1538 -9619
rect -1635 -9713 -1538 -9700
rect -1478 -9617 -1381 -9604
rect -1478 -9698 -1463 -9617
rect -1395 -9698 -1381 -9617
rect -1478 -9711 -1381 -9698
rect -1263 -9632 -1237 -9586
rect -1191 -9632 -1166 -9586
rect -1263 -9684 -1166 -9632
rect -1263 -9730 -1237 -9684
rect -1191 -9720 -1166 -9684
rect -1011 -9720 -765 -9520
rect -574 -9550 -477 -9520
rect -574 -9596 -549 -9550
rect -503 -9596 -477 -9550
rect -4 -9555 203 -9509
rect -574 -9648 -477 -9596
rect -574 -9694 -549 -9648
rect -503 -9694 -477 -9648
rect 157 -9681 203 -9555
rect 288 -9572 300 -9506
rect 366 -9572 378 -9506
rect 638 -9509 684 -8747
rect 288 -9584 378 -9572
rect 477 -9555 684 -9509
rect 798 -9473 844 -8387
rect 1190 -8420 1215 -8374
rect 1261 -8420 1287 -8374
rect 1190 -8472 1287 -8420
rect 1190 -8518 1215 -8472
rect 1261 -8518 1287 -8472
rect 1190 -8537 1287 -8518
rect 1381 -8537 1496 -8113
rect 1659 -8271 1859 -8113
rect 2059 -8271 2259 -8113
rect 2459 -8271 2659 -8113
rect 2859 -8271 3059 -8113
rect 3259 -8271 3459 -8113
rect 3659 -8271 3859 -8113
rect 4374 -8137 4471 -8113
rect 4374 -8183 4400 -8137
rect 4446 -8183 4471 -8137
rect 4374 -8235 4471 -8183
rect 4374 -8271 4400 -8235
rect 1611 -8281 4400 -8271
rect 4446 -8281 4471 -8235
rect 1611 -8296 4471 -8281
rect 1611 -8342 1636 -8296
rect 1682 -8297 2910 -8296
rect 1682 -8342 1734 -8297
rect 1611 -8343 1734 -8342
rect 1780 -8343 1832 -8297
rect 1878 -8343 1930 -8297
rect 1976 -8343 2028 -8297
rect 2074 -8343 2126 -8297
rect 2172 -8343 2224 -8297
rect 2270 -8343 2322 -8297
rect 2368 -8343 2420 -8297
rect 2466 -8343 2518 -8297
rect 2564 -8343 2616 -8297
rect 2662 -8343 2714 -8297
rect 2760 -8343 2812 -8297
rect 2858 -8342 2910 -8297
rect 2956 -8333 4471 -8296
rect 2956 -8342 4400 -8333
rect 2858 -8343 4400 -8342
rect 1611 -8368 4400 -8343
rect 1611 -8394 1708 -8368
rect 1611 -8440 1636 -8394
rect 1682 -8440 1708 -8394
rect 1611 -8492 1708 -8440
rect 1611 -8537 1636 -8492
rect 1190 -8538 1636 -8537
rect 1682 -8538 1708 -8492
rect 1190 -8570 1708 -8538
rect 892 -8588 982 -8576
rect 892 -8654 904 -8588
rect 970 -8654 982 -8588
rect 892 -8666 982 -8654
rect 1190 -8616 1215 -8570
rect 1261 -8590 1708 -8570
rect 1261 -8616 1636 -8590
rect 1190 -8636 1636 -8616
rect 1682 -8636 1708 -8590
rect 1190 -8668 1708 -8636
rect 1190 -8714 1215 -8668
rect 1261 -8688 1708 -8668
rect 1261 -8714 1636 -8688
rect 1190 -8734 1636 -8714
rect 1682 -8734 1708 -8688
rect 1190 -8737 1708 -8734
rect 1190 -8766 1287 -8737
rect 1190 -8812 1215 -8766
rect 1261 -8812 1287 -8766
rect 1190 -8864 1287 -8812
rect 1190 -8910 1215 -8864
rect 1261 -8910 1287 -8864
rect 1190 -8937 1287 -8910
rect 1381 -8937 1496 -8737
rect 1611 -8786 1708 -8737
rect 1611 -8832 1636 -8786
rect 1682 -8832 1708 -8786
rect 1611 -8884 1708 -8832
rect 1611 -8930 1636 -8884
rect 1682 -8930 1708 -8884
rect 1611 -8937 1708 -8930
rect 1190 -8962 1708 -8937
rect 1190 -9008 1215 -8962
rect 1261 -8982 1708 -8962
rect 1261 -9008 1636 -8982
rect 1190 -9028 1636 -9008
rect 1682 -9028 1708 -8982
rect 1190 -9060 1708 -9028
rect 1190 -9106 1215 -9060
rect 1261 -9080 1708 -9060
rect 1261 -9106 1636 -9080
rect 1190 -9126 1636 -9106
rect 1682 -9126 1708 -9080
rect 1790 -9089 1856 -8368
rect 1190 -9137 1708 -9126
rect 1190 -9158 1287 -9137
rect 1190 -9204 1215 -9158
rect 1261 -9204 1287 -9158
rect 1190 -9256 1287 -9204
rect 1190 -9302 1215 -9256
rect 1261 -9302 1287 -9256
rect 1190 -9337 1287 -9302
rect 1381 -9337 1496 -9137
rect 1611 -9178 1708 -9137
rect 1950 -9138 2016 -8488
rect 2110 -9089 2176 -8368
rect 2269 -9138 2335 -8489
rect 2430 -9090 2496 -8368
rect 2590 -9138 2656 -8489
rect 2749 -9089 2815 -8368
rect 2884 -8379 4400 -8368
rect 4446 -8379 4471 -8333
rect 2884 -8394 4471 -8379
rect 2884 -8440 2910 -8394
rect 2956 -8431 4471 -8394
rect 2956 -8436 4400 -8431
rect 2956 -8440 2981 -8436
rect 2884 -8492 2981 -8440
rect 2884 -8538 2910 -8492
rect 2956 -8538 2981 -8492
rect 2884 -8590 2981 -8538
rect 2884 -8636 2910 -8590
rect 2956 -8607 2981 -8590
rect 3259 -8607 3459 -8436
rect 3659 -8607 3859 -8436
rect 4374 -8477 4400 -8436
rect 4446 -8477 4471 -8431
rect 4374 -8529 4471 -8477
rect 4374 -8575 4400 -8529
rect 4446 -8575 4471 -8529
rect 4374 -8607 4471 -8575
rect 2956 -8627 4471 -8607
rect 2956 -8636 4400 -8627
rect 2884 -8673 4400 -8636
rect 4446 -8673 4471 -8627
rect 2884 -8688 4471 -8673
rect 2884 -8734 2910 -8688
rect 2956 -8725 4471 -8688
rect 2956 -8734 4400 -8725
rect 2884 -8771 4400 -8734
rect 4446 -8771 4471 -8725
rect 2884 -8786 4471 -8771
rect 2884 -8832 2910 -8786
rect 2956 -8823 4471 -8786
rect 2956 -8832 4400 -8823
rect 2884 -8869 4400 -8832
rect 4446 -8869 4471 -8823
rect 2884 -8884 4471 -8869
rect 2884 -8930 2910 -8884
rect 2956 -8896 4471 -8884
rect 4545 -7540 4609 -6837
rect 4844 -7540 4908 -6837
rect 4988 -7218 5052 -6971
rect 4970 -7232 5067 -7218
rect 4970 -7296 4986 -7232
rect 5050 -7296 5067 -7232
rect 4970 -7348 5067 -7296
rect 4970 -7412 4986 -7348
rect 5050 -7412 5067 -7348
rect 4970 -7430 5067 -7412
rect 4545 -7553 4908 -7540
rect 4545 -7603 4646 -7553
rect 4696 -7603 4759 -7553
rect 4809 -7603 4908 -7553
rect 4545 -7615 4908 -7603
rect 4545 -8079 4609 -7615
rect 4844 -8079 4908 -7615
rect 4988 -7805 5052 -7430
rect 4970 -7819 5067 -7805
rect 4970 -7883 4986 -7819
rect 5050 -7883 5067 -7819
rect 4970 -7935 5067 -7883
rect 4970 -7999 4986 -7935
rect 5050 -7999 5067 -7935
rect 4970 -8017 5067 -7999
rect 4545 -8092 4908 -8079
rect 4545 -8142 4646 -8092
rect 4696 -8142 4759 -8092
rect 4809 -8142 4908 -8092
rect 4545 -8154 4908 -8142
rect 4545 -8896 4609 -8154
rect 4844 -8896 4908 -8154
rect 4988 -8324 5052 -8017
rect 4970 -8338 5067 -8324
rect 4970 -8402 4986 -8338
rect 5050 -8402 5067 -8338
rect 4970 -8454 5067 -8402
rect 4970 -8518 4986 -8454
rect 5050 -8518 5067 -8454
rect 4970 -8536 5067 -8518
rect 4988 -8659 5052 -8536
rect 5289 -8896 5353 -6837
rect 5592 -7219 5656 -6964
rect 5576 -7233 5673 -7219
rect 5576 -7297 5592 -7233
rect 5656 -7297 5673 -7233
rect 5576 -7349 5673 -7297
rect 5576 -7413 5592 -7349
rect 5656 -7413 5673 -7349
rect 5576 -7431 5673 -7413
rect 5592 -7806 5656 -7431
rect 5576 -7820 5673 -7806
rect 5576 -7884 5592 -7820
rect 5656 -7884 5673 -7820
rect 5576 -7936 5673 -7884
rect 5576 -8000 5592 -7936
rect 5656 -8000 5673 -7936
rect 5576 -8018 5673 -8000
rect 5592 -8325 5656 -8018
rect 5576 -8339 5673 -8325
rect 5576 -8403 5592 -8339
rect 5656 -8403 5673 -8339
rect 5576 -8455 5673 -8403
rect 5576 -8519 5592 -8455
rect 5656 -8519 5673 -8455
rect 5576 -8537 5673 -8519
rect 5592 -8652 5656 -8537
rect 5897 -8896 5961 -6837
rect 6120 -6952 6352 -6938
rect 6120 -7018 6135 -6952
rect 6201 -7018 6273 -6952
rect 6339 -7018 6352 -6952
rect 6120 -7031 6352 -7018
rect 6201 -7217 6265 -7031
rect 6185 -7231 6282 -7217
rect 6185 -7295 6201 -7231
rect 6265 -7295 6282 -7231
rect 6185 -7347 6282 -7295
rect 6185 -7411 6201 -7347
rect 6265 -7411 6282 -7347
rect 6185 -7429 6282 -7411
rect 6201 -7541 6265 -7429
rect 6140 -7553 6327 -7541
rect 6140 -7603 6152 -7553
rect 6202 -7603 6265 -7553
rect 6315 -7603 6327 -7553
rect 6140 -7614 6327 -7603
rect 6201 -7804 6265 -7614
rect 6185 -7818 6282 -7804
rect 6185 -7882 6201 -7818
rect 6265 -7882 6282 -7818
rect 6185 -7934 6282 -7882
rect 6185 -7998 6201 -7934
rect 6265 -7998 6282 -7934
rect 6185 -8016 6282 -7998
rect 6201 -8077 6265 -8016
rect 6138 -8089 6325 -8077
rect 6138 -8139 6150 -8089
rect 6200 -8139 6263 -8089
rect 6313 -8139 6325 -8089
rect 6138 -8150 6325 -8139
rect 6201 -8323 6265 -8150
rect 6185 -8337 6282 -8323
rect 6185 -8401 6201 -8337
rect 6265 -8401 6282 -8337
rect 6185 -8453 6282 -8401
rect 6185 -8517 6201 -8453
rect 6265 -8517 6282 -8453
rect 6185 -8535 6282 -8517
rect 6201 -8669 6265 -8535
rect 6117 -8683 6349 -8669
rect 6117 -8749 6132 -8683
rect 6198 -8749 6270 -8683
rect 6336 -8749 6349 -8683
rect 6117 -8762 6349 -8749
rect 6505 -8896 6569 -6837
rect 6809 -7220 6873 -6980
rect 6794 -7234 6891 -7220
rect 6794 -7298 6810 -7234
rect 6874 -7298 6891 -7234
rect 6794 -7350 6891 -7298
rect 6794 -7414 6810 -7350
rect 6874 -7414 6891 -7350
rect 6794 -7432 6891 -7414
rect 6809 -7807 6873 -7432
rect 6794 -7821 6891 -7807
rect 6794 -7885 6810 -7821
rect 6874 -7885 6891 -7821
rect 6794 -7937 6891 -7885
rect 6794 -8001 6810 -7937
rect 6874 -8001 6891 -7937
rect 6794 -8019 6891 -8001
rect 6809 -8326 6873 -8019
rect 6794 -8340 6891 -8326
rect 6794 -8404 6810 -8340
rect 6874 -8404 6891 -8340
rect 6794 -8456 6891 -8404
rect 6794 -8520 6810 -8456
rect 6874 -8520 6891 -8456
rect 6794 -8538 6891 -8520
rect 6809 -8668 6873 -8538
rect 7113 -8896 7177 -6837
rect 7417 -7228 7481 -6976
rect 7397 -7242 7494 -7228
rect 7397 -7306 7413 -7242
rect 7477 -7306 7494 -7242
rect 7397 -7358 7494 -7306
rect 7397 -7422 7413 -7358
rect 7477 -7422 7494 -7358
rect 7397 -7440 7494 -7422
rect 7417 -7815 7481 -7440
rect 7554 -7540 7618 -6837
rect 7855 -7540 7919 -6837
rect 7554 -7553 7919 -7540
rect 7554 -7603 7654 -7553
rect 7704 -7603 7767 -7553
rect 7817 -7603 7919 -7553
rect 7554 -7615 7919 -7603
rect 7397 -7829 7494 -7815
rect 7397 -7893 7413 -7829
rect 7477 -7893 7494 -7829
rect 7397 -7945 7494 -7893
rect 7397 -8009 7413 -7945
rect 7477 -8009 7494 -7945
rect 7397 -8027 7494 -8009
rect 7417 -8334 7481 -8027
rect 7554 -8074 7618 -7615
rect 7855 -8074 7919 -7615
rect 7554 -8087 7919 -8074
rect 7554 -8137 7654 -8087
rect 7704 -8137 7767 -8087
rect 7817 -8137 7919 -8087
rect 7554 -8149 7919 -8137
rect 7397 -8348 7494 -8334
rect 7397 -8412 7413 -8348
rect 7477 -8412 7494 -8348
rect 7397 -8464 7494 -8412
rect 7397 -8528 7413 -8464
rect 7477 -8528 7494 -8464
rect 7397 -8546 7494 -8528
rect 7417 -8664 7481 -8546
rect 7554 -8896 7618 -8149
rect 7855 -8896 7919 -8149
rect 8000 -6838 8786 -6837
rect 8832 -6838 8858 -6792
rect 8000 -6864 8858 -6838
rect 8000 -6910 8026 -6864
rect 8072 -6890 8858 -6864
rect 8072 -6910 8786 -6890
rect 8000 -6936 8786 -6910
rect 8832 -6936 8858 -6890
rect 8000 -6962 8858 -6936
rect 8000 -7008 8026 -6962
rect 8072 -6988 8858 -6962
rect 8072 -7008 8786 -6988
rect 8000 -7034 8786 -7008
rect 8832 -7034 8858 -6988
rect 8000 -7039 8858 -7034
rect 8000 -7060 8097 -7039
rect 8000 -7106 8026 -7060
rect 8072 -7106 8097 -7060
rect 8000 -7158 8097 -7106
rect 8000 -7204 8026 -7158
rect 8072 -7204 8097 -7158
rect 8000 -7219 8097 -7204
rect 8298 -7219 8562 -7039
rect 8760 -7086 8858 -7039
rect 8760 -7132 8786 -7086
rect 8832 -7132 8858 -7086
rect 8760 -7184 8858 -7132
rect 8760 -7219 8786 -7184
rect 8000 -7230 8786 -7219
rect 8832 -7230 8858 -7184
rect 8000 -7256 8858 -7230
rect 8000 -7302 8026 -7256
rect 8072 -7282 8858 -7256
rect 8072 -7302 8786 -7282
rect 8000 -7328 8786 -7302
rect 8832 -7328 8858 -7282
rect 8000 -7354 8858 -7328
rect 8000 -7400 8026 -7354
rect 8072 -7380 8858 -7354
rect 8072 -7400 8786 -7380
rect 8000 -7426 8786 -7400
rect 8832 -7426 8858 -7380
rect 8000 -7452 8858 -7426
rect 8945 -5742 9006 -4806
rect 9104 -5742 9165 -4806
rect 9246 -4967 9336 -4955
rect 9246 -5034 9259 -4967
rect 9324 -5034 9336 -4967
rect 9246 -5046 9336 -5034
rect 9264 -5319 9325 -5110
rect 9246 -5333 9343 -5319
rect 9246 -5397 9262 -5333
rect 9326 -5397 9343 -5333
rect 9246 -5449 9343 -5397
rect 9246 -5513 9262 -5449
rect 9326 -5513 9343 -5449
rect 9246 -5531 9343 -5513
rect 8945 -5754 9165 -5742
rect 8945 -5805 9029 -5754
rect 9080 -5805 9165 -5754
rect 8945 -5817 9165 -5805
rect 8945 -6479 9006 -5817
rect 9104 -6479 9165 -5817
rect 9264 -6045 9325 -5531
rect 9248 -6059 9345 -6045
rect 9248 -6123 9264 -6059
rect 9328 -6123 9345 -6059
rect 9248 -6175 9345 -6123
rect 9248 -6239 9264 -6175
rect 9328 -6239 9345 -6175
rect 9248 -6257 9345 -6239
rect 8945 -6491 9165 -6479
rect 8945 -6542 9029 -6491
rect 9080 -6542 9165 -6491
rect 8945 -6554 9165 -6542
rect 8945 -7452 9006 -6554
rect 9104 -7452 9165 -6554
rect 9264 -6776 9325 -6257
rect 9246 -6790 9343 -6776
rect 9246 -6854 9262 -6790
rect 9326 -6854 9343 -6790
rect 9246 -6906 9343 -6854
rect 9246 -6970 9262 -6906
rect 9326 -6970 9343 -6906
rect 9246 -6988 9343 -6970
rect 9264 -7183 9325 -6988
rect 9245 -7258 9335 -7246
rect 9245 -7325 9258 -7258
rect 9323 -7325 9335 -7258
rect 9245 -7337 9335 -7325
rect 9424 -7452 9485 -4806
rect 9560 -4966 9650 -4954
rect 9560 -5033 9573 -4966
rect 9638 -5033 9650 -4966
rect 9560 -5045 9650 -5033
rect 9585 -5319 9646 -5111
rect 9566 -5333 9663 -5319
rect 9566 -5397 9582 -5333
rect 9646 -5397 9663 -5333
rect 9566 -5449 9663 -5397
rect 9566 -5513 9582 -5449
rect 9646 -5513 9663 -5449
rect 9566 -5531 9663 -5513
rect 9585 -6047 9646 -5531
rect 9568 -6061 9665 -6047
rect 9568 -6125 9584 -6061
rect 9648 -6125 9665 -6061
rect 9568 -6177 9665 -6125
rect 9568 -6241 9584 -6177
rect 9648 -6241 9665 -6177
rect 9568 -6259 9665 -6241
rect 9585 -6776 9646 -6259
rect 9568 -6790 9665 -6776
rect 9568 -6854 9584 -6790
rect 9648 -6854 9665 -6790
rect 9568 -6906 9665 -6854
rect 9568 -6970 9584 -6906
rect 9648 -6970 9665 -6906
rect 9568 -6988 9665 -6970
rect 9585 -7183 9646 -6988
rect 9573 -7255 9663 -7243
rect 9573 -7322 9586 -7255
rect 9651 -7322 9663 -7255
rect 9573 -7334 9663 -7322
rect 9745 -7452 9806 -4806
rect 9877 -4963 9967 -4951
rect 9877 -5030 9890 -4963
rect 9955 -5030 9967 -4963
rect 9877 -5042 9967 -5030
rect 9904 -5319 9965 -5111
rect 9887 -5333 9984 -5319
rect 9887 -5397 9903 -5333
rect 9967 -5397 9984 -5333
rect 9887 -5449 9984 -5397
rect 9887 -5513 9903 -5449
rect 9967 -5513 9984 -5449
rect 9887 -5531 9984 -5513
rect 9904 -6049 9965 -5531
rect 9888 -6063 9985 -6049
rect 9888 -6127 9904 -6063
rect 9968 -6127 9985 -6063
rect 9888 -6179 9985 -6127
rect 9888 -6243 9904 -6179
rect 9968 -6243 9985 -6179
rect 9888 -6261 9985 -6243
rect 9904 -6776 9965 -6261
rect 9887 -6790 9984 -6776
rect 9887 -6854 9903 -6790
rect 9967 -6854 9984 -6790
rect 9887 -6906 9984 -6854
rect 9887 -6970 9903 -6906
rect 9967 -6970 9984 -6906
rect 9887 -6988 9984 -6970
rect 9904 -7183 9965 -6988
rect 9883 -7256 9973 -7244
rect 9883 -7323 9896 -7256
rect 9961 -7323 9973 -7256
rect 9883 -7335 9973 -7323
rect 10064 -7452 10125 -4806
rect 10208 -4962 10298 -4950
rect 10208 -5029 10221 -4962
rect 10286 -5029 10298 -4962
rect 10208 -5041 10298 -5029
rect 10224 -5322 10285 -5110
rect 10207 -5336 10304 -5322
rect 10207 -5400 10223 -5336
rect 10287 -5400 10304 -5336
rect 10207 -5452 10304 -5400
rect 10207 -5516 10223 -5452
rect 10287 -5516 10304 -5452
rect 10207 -5534 10304 -5516
rect 10224 -6049 10285 -5534
rect 10208 -6063 10305 -6049
rect 10208 -6127 10224 -6063
rect 10288 -6127 10305 -6063
rect 10208 -6179 10305 -6127
rect 10208 -6243 10224 -6179
rect 10288 -6243 10305 -6179
rect 10208 -6261 10305 -6243
rect 10224 -6778 10285 -6261
rect 10207 -6792 10304 -6778
rect 10207 -6856 10223 -6792
rect 10287 -6856 10304 -6792
rect 10207 -6908 10304 -6856
rect 10207 -6972 10223 -6908
rect 10287 -6972 10304 -6908
rect 10207 -6990 10304 -6972
rect 10224 -7181 10285 -6990
rect 10209 -7256 10299 -7244
rect 10209 -7323 10222 -7256
rect 10287 -7323 10299 -7256
rect 10209 -7335 10299 -7323
rect 10384 -7452 10445 -4806
rect 10527 -4963 10617 -4951
rect 10527 -5030 10540 -4963
rect 10605 -5030 10617 -4963
rect 10527 -5042 10617 -5030
rect 10544 -5320 10605 -5111
rect 10527 -5334 10624 -5320
rect 10527 -5398 10543 -5334
rect 10607 -5398 10624 -5334
rect 10527 -5450 10624 -5398
rect 10527 -5514 10543 -5450
rect 10607 -5514 10624 -5450
rect 10527 -5532 10624 -5514
rect 10544 -6049 10605 -5532
rect 10704 -5743 10765 -4806
rect 10864 -5743 10925 -4806
rect 10704 -5755 10925 -5743
rect 10704 -5806 10788 -5755
rect 10839 -5806 10925 -5755
rect 10704 -5818 10925 -5806
rect 10525 -6063 10622 -6049
rect 10525 -6127 10541 -6063
rect 10605 -6127 10622 -6063
rect 10525 -6179 10622 -6127
rect 10525 -6243 10541 -6179
rect 10605 -6243 10622 -6179
rect 10525 -6261 10622 -6243
rect 10544 -6778 10605 -6261
rect 10704 -6479 10765 -5818
rect 10864 -6479 10925 -5818
rect 10704 -6491 10925 -6479
rect 10704 -6542 10788 -6491
rect 10839 -6542 10925 -6491
rect 10704 -6554 10925 -6542
rect 10527 -6792 10624 -6778
rect 10527 -6856 10543 -6792
rect 10607 -6856 10624 -6792
rect 10527 -6908 10624 -6856
rect 10527 -6972 10543 -6908
rect 10607 -6972 10624 -6908
rect 10527 -6990 10624 -6972
rect 10544 -7183 10605 -6990
rect 10524 -7252 10614 -7240
rect 10524 -7319 10537 -7252
rect 10602 -7319 10614 -7252
rect 10524 -7331 10614 -7319
rect 10704 -7452 10765 -6554
rect 10864 -7452 10925 -6554
rect 11014 -4832 11112 -4806
rect 11014 -4878 11040 -4832
rect 11086 -4878 11112 -4832
rect 11014 -4930 11112 -4878
rect 11014 -4976 11040 -4930
rect 11086 -4976 11112 -4930
rect 11014 -5028 11112 -4976
rect 11014 -5074 11040 -5028
rect 11086 -5074 11112 -5028
rect 11014 -5126 11112 -5074
rect 11014 -5172 11040 -5126
rect 11086 -5172 11112 -5126
rect 11014 -5224 11112 -5172
rect 11014 -5270 11040 -5224
rect 11086 -5270 11112 -5224
rect 11014 -5322 11112 -5270
rect 11014 -5368 11040 -5322
rect 11086 -5368 11112 -5322
rect 11014 -5420 11112 -5368
rect 11014 -5466 11040 -5420
rect 11086 -5466 11112 -5420
rect 11014 -5518 11112 -5466
rect 11014 -5564 11040 -5518
rect 11086 -5564 11112 -5518
rect 11014 -5616 11112 -5564
rect 11014 -5662 11040 -5616
rect 11086 -5662 11112 -5616
rect 11014 -5714 11112 -5662
rect 11014 -5760 11040 -5714
rect 11086 -5760 11112 -5714
rect 11014 -5812 11112 -5760
rect 11014 -5858 11040 -5812
rect 11086 -5858 11112 -5812
rect 11014 -5910 11112 -5858
rect 11014 -5956 11040 -5910
rect 11086 -5956 11112 -5910
rect 11014 -6008 11112 -5956
rect 11014 -6054 11040 -6008
rect 11086 -6054 11112 -6008
rect 11014 -6106 11112 -6054
rect 11014 -6152 11040 -6106
rect 11086 -6152 11112 -6106
rect 11014 -6204 11112 -6152
rect 11014 -6250 11040 -6204
rect 11086 -6250 11112 -6204
rect 11014 -6302 11112 -6250
rect 11014 -6348 11040 -6302
rect 11086 -6348 11112 -6302
rect 11014 -6400 11112 -6348
rect 11014 -6446 11040 -6400
rect 11086 -6446 11112 -6400
rect 11014 -6498 11112 -6446
rect 11014 -6544 11040 -6498
rect 11086 -6544 11112 -6498
rect 11014 -6596 11112 -6544
rect 11014 -6642 11040 -6596
rect 11086 -6642 11112 -6596
rect 11014 -6694 11112 -6642
rect 11014 -6740 11040 -6694
rect 11086 -6740 11112 -6694
rect 11014 -6792 11112 -6740
rect 11014 -6838 11040 -6792
rect 11086 -6838 11112 -6792
rect 11014 -6890 11112 -6838
rect 11014 -6936 11040 -6890
rect 11086 -6936 11112 -6890
rect 11014 -6988 11112 -6936
rect 11014 -7034 11040 -6988
rect 11086 -7034 11112 -6988
rect 11014 -7086 11112 -7034
rect 11014 -7132 11040 -7086
rect 11086 -7132 11112 -7086
rect 11014 -7184 11112 -7132
rect 11014 -7230 11040 -7184
rect 11086 -7230 11112 -7184
rect 11014 -7282 11112 -7230
rect 11014 -7328 11040 -7282
rect 11086 -7328 11112 -7282
rect 11014 -7380 11112 -7328
rect 11014 -7426 11040 -7380
rect 11086 -7426 11112 -7380
rect 11014 -7452 11112 -7426
rect 8000 -7498 8026 -7452
rect 8072 -7478 11112 -7452
rect 8072 -7498 8786 -7478
rect 8000 -7499 8786 -7498
rect 8000 -7550 8097 -7499
rect 8000 -7596 8026 -7550
rect 8072 -7596 8097 -7550
rect 8000 -7648 8097 -7596
rect 8000 -7694 8026 -7648
rect 8072 -7694 8097 -7648
rect 8000 -7746 8097 -7694
rect 8000 -7792 8026 -7746
rect 8072 -7792 8097 -7746
rect 8000 -7826 8097 -7792
rect 8298 -7826 8562 -7499
rect 8760 -7524 8786 -7499
rect 8832 -7524 8884 -7478
rect 8930 -7524 8982 -7478
rect 9028 -7524 9080 -7478
rect 9126 -7524 9178 -7478
rect 9224 -7524 9276 -7478
rect 9322 -7524 9374 -7478
rect 9420 -7524 9472 -7478
rect 9518 -7524 9570 -7478
rect 9616 -7524 9668 -7478
rect 9714 -7524 9766 -7478
rect 9812 -7524 9864 -7478
rect 9910 -7524 9962 -7478
rect 10008 -7524 10060 -7478
rect 10106 -7524 10158 -7478
rect 10204 -7524 10256 -7478
rect 10302 -7524 10354 -7478
rect 10400 -7524 10452 -7478
rect 10498 -7524 10550 -7478
rect 10596 -7524 10648 -7478
rect 10694 -7524 10746 -7478
rect 10792 -7524 10844 -7478
rect 10890 -7524 10942 -7478
rect 10988 -7524 11040 -7478
rect 11086 -7524 11112 -7478
rect 8760 -7550 11112 -7524
rect 8846 -7708 9046 -7550
rect 9246 -7708 9446 -7550
rect 9646 -7708 9846 -7550
rect 10046 -7708 10246 -7550
rect 10446 -7708 10646 -7550
rect 10846 -7708 11046 -7550
rect 8760 -7734 11112 -7708
rect 8760 -7780 8786 -7734
rect 8832 -7780 8884 -7734
rect 8930 -7780 8982 -7734
rect 9028 -7780 9080 -7734
rect 9126 -7780 9178 -7734
rect 9224 -7780 9276 -7734
rect 9322 -7780 9374 -7734
rect 9420 -7780 9472 -7734
rect 9518 -7780 9570 -7734
rect 9616 -7780 9668 -7734
rect 9714 -7780 9766 -7734
rect 9812 -7780 9864 -7734
rect 9910 -7780 9962 -7734
rect 10008 -7780 10060 -7734
rect 10106 -7780 10158 -7734
rect 10204 -7780 10256 -7734
rect 10302 -7780 10354 -7734
rect 10400 -7780 10452 -7734
rect 10498 -7780 10550 -7734
rect 10596 -7780 10648 -7734
rect 10694 -7780 10746 -7734
rect 10792 -7780 10844 -7734
rect 10890 -7780 10942 -7734
rect 10988 -7780 11040 -7734
rect 11086 -7780 11112 -7734
rect 8760 -7806 11112 -7780
rect 8760 -7826 8858 -7806
rect 8000 -7832 8858 -7826
rect 8000 -7844 8786 -7832
rect 8000 -7890 8026 -7844
rect 8072 -7878 8786 -7844
rect 8832 -7878 8858 -7832
rect 8072 -7890 8858 -7878
rect 8000 -7930 8858 -7890
rect 8000 -7942 8786 -7930
rect 8000 -7988 8026 -7942
rect 8072 -7976 8786 -7942
rect 8832 -7976 8858 -7930
rect 8072 -7988 8858 -7976
rect 8000 -8028 8858 -7988
rect 8000 -8040 8786 -8028
rect 8000 -8086 8026 -8040
rect 8072 -8074 8786 -8040
rect 8832 -8074 8858 -8028
rect 8072 -8086 8858 -8074
rect 8000 -8106 8858 -8086
rect 8000 -8138 8097 -8106
rect 8000 -8184 8026 -8138
rect 8072 -8184 8097 -8138
rect 8000 -8236 8097 -8184
rect 8000 -8282 8026 -8236
rect 8072 -8282 8097 -8236
rect 8000 -8334 8097 -8282
rect 8000 -8380 8026 -8334
rect 8072 -8380 8097 -8334
rect 8000 -8409 8097 -8380
rect 8298 -8409 8562 -8106
rect 8760 -8126 8858 -8106
rect 8760 -8172 8786 -8126
rect 8832 -8172 8858 -8126
rect 8760 -8224 8858 -8172
rect 8760 -8270 8786 -8224
rect 8832 -8270 8858 -8224
rect 8760 -8322 8858 -8270
rect 8760 -8368 8786 -8322
rect 8832 -8368 8858 -8322
rect 8760 -8409 8858 -8368
rect 8000 -8420 8858 -8409
rect 8000 -8432 8786 -8420
rect 8000 -8478 8026 -8432
rect 8072 -8466 8786 -8432
rect 8832 -8466 8858 -8420
rect 8072 -8478 8858 -8466
rect 8000 -8518 8858 -8478
rect 8000 -8530 8786 -8518
rect 8000 -8576 8026 -8530
rect 8072 -8564 8786 -8530
rect 8832 -8564 8858 -8518
rect 8072 -8576 8858 -8564
rect 8000 -8616 8858 -8576
rect 8000 -8628 8786 -8616
rect 8000 -8674 8026 -8628
rect 8072 -8662 8786 -8628
rect 8832 -8662 8858 -8616
rect 8072 -8674 8858 -8662
rect 8000 -8689 8858 -8674
rect 8000 -8726 8097 -8689
rect 8000 -8772 8026 -8726
rect 8072 -8772 8097 -8726
rect 8000 -8824 8097 -8772
rect 8000 -8870 8026 -8824
rect 8072 -8870 8097 -8824
rect 8000 -8896 8097 -8870
rect 2956 -8898 8097 -8896
rect 2956 -8930 2981 -8898
rect 2884 -8982 2981 -8930
rect 2884 -9028 2910 -8982
rect 2956 -9028 2981 -8982
rect 2884 -9080 2981 -9028
rect 2884 -9126 2910 -9080
rect 2956 -9126 2981 -9080
rect 1611 -9224 1636 -9178
rect 1682 -9224 1708 -9178
rect 1611 -9276 1708 -9224
rect 1892 -9150 2715 -9138
rect 1892 -9151 2544 -9150
rect 1892 -9203 1905 -9151
rect 1957 -9152 2544 -9151
rect 1957 -9177 2011 -9152
rect 1892 -9241 1928 -9203
rect 1992 -9204 2011 -9177
rect 2063 -9179 2223 -9152
rect 2275 -9153 2544 -9152
rect 2063 -9204 2073 -9179
rect 1992 -9241 2073 -9204
rect 1892 -9243 2073 -9241
rect 2137 -9243 2207 -9179
rect 2275 -9204 2329 -9153
rect 2271 -9205 2329 -9204
rect 2381 -9202 2544 -9153
rect 2596 -9151 2715 -9150
rect 2596 -9202 2650 -9151
rect 2381 -9203 2650 -9202
rect 2702 -9203 2715 -9151
rect 2381 -9205 2715 -9203
rect 2271 -9243 2715 -9205
rect 1892 -9264 2715 -9243
rect 2884 -9178 2981 -9126
rect 2884 -9224 2910 -9178
rect 2956 -9224 2981 -9178
rect 1611 -9322 1636 -9276
rect 1682 -9322 1708 -9276
rect 1611 -9337 1708 -9322
rect 1190 -9354 1708 -9337
rect 1190 -9400 1215 -9354
rect 1261 -9374 1708 -9354
rect 1261 -9400 1636 -9374
rect 958 -9473 1004 -9410
rect 798 -9474 1004 -9473
rect 798 -9520 880 -9474
rect 926 -9520 1004 -9474
rect 1190 -9420 1636 -9400
rect 1682 -9420 1708 -9374
rect 1190 -9452 1708 -9420
rect 2884 -9276 2981 -9224
rect 2884 -9322 2910 -9276
rect 2956 -9309 2981 -9276
rect 3259 -9309 3459 -8898
rect 3659 -9309 3859 -8898
rect 4374 -8921 8097 -8898
rect 4374 -8967 4399 -8921
rect 4445 -8922 8097 -8921
rect 4445 -8967 4497 -8922
rect 4374 -8968 4497 -8967
rect 4543 -8968 4595 -8922
rect 4641 -8968 4693 -8922
rect 4739 -8968 4791 -8922
rect 4837 -8968 4889 -8922
rect 4935 -8968 4987 -8922
rect 5033 -8968 5085 -8922
rect 5131 -8968 5183 -8922
rect 5229 -8968 5281 -8922
rect 5327 -8968 5379 -8922
rect 5425 -8968 5477 -8922
rect 5523 -8968 5575 -8922
rect 5621 -8968 5673 -8922
rect 5719 -8968 5771 -8922
rect 5817 -8968 5869 -8922
rect 5915 -8968 5967 -8922
rect 6013 -8968 6065 -8922
rect 6111 -8968 6163 -8922
rect 6209 -8968 6261 -8922
rect 6307 -8968 6359 -8922
rect 6405 -8968 6457 -8922
rect 6503 -8968 6555 -8922
rect 6601 -8968 6653 -8922
rect 6699 -8968 6751 -8922
rect 6797 -8968 6849 -8922
rect 6895 -8968 6947 -8922
rect 6993 -8968 7045 -8922
rect 7091 -8968 7143 -8922
rect 7189 -8968 7241 -8922
rect 7287 -8968 7339 -8922
rect 7385 -8968 7437 -8922
rect 7483 -8968 7535 -8922
rect 7581 -8968 7633 -8922
rect 7679 -8968 7731 -8922
rect 7777 -8968 7829 -8922
rect 7875 -8968 7927 -8922
rect 7973 -8968 8025 -8922
rect 8071 -8968 8097 -8922
rect 8298 -8968 8562 -8689
rect 8760 -8714 8858 -8689
rect 8760 -8760 8786 -8714
rect 8832 -8760 8858 -8714
rect 8760 -8812 8858 -8760
rect 8760 -8858 8786 -8812
rect 8832 -8858 8858 -8812
rect 8760 -8910 8858 -8858
rect 8760 -8956 8786 -8910
rect 8832 -8956 8858 -8910
rect 8760 -8968 8858 -8956
rect 4374 -8993 8858 -8968
rect 4437 -9008 8858 -8993
rect 4437 -9054 8786 -9008
rect 8832 -9054 8858 -9008
rect 4437 -9106 8858 -9054
rect 4437 -9152 8786 -9106
rect 8832 -9152 8858 -9106
rect 4437 -9204 8858 -9152
rect 4437 -9244 8786 -9204
rect 4437 -9309 4696 -9244
rect 2956 -9322 4696 -9309
rect 2884 -9374 4696 -9322
rect 2884 -9420 2910 -9374
rect 2956 -9404 4696 -9374
rect 6080 -9404 6620 -9244
rect 8298 -9404 8562 -9244
rect 8760 -9250 8786 -9244
rect 8832 -9250 8858 -9204
rect 8760 -9302 8858 -9250
rect 8760 -9348 8786 -9302
rect 8832 -9348 8858 -9302
rect 8760 -9400 8858 -9348
rect 8760 -9404 8786 -9400
rect 2956 -9420 8786 -9404
rect 1190 -9498 1215 -9452
rect 1261 -9472 1708 -9452
rect 1261 -9498 1636 -9472
rect 1190 -9518 1636 -9498
rect 1682 -9518 1708 -9472
rect 1190 -9537 1708 -9518
rect 1190 -9550 1287 -9537
rect 477 -9681 523 -9555
rect 1190 -9596 1215 -9550
rect 1261 -9596 1287 -9550
rect 1190 -9648 1287 -9596
rect -574 -9720 -477 -9694
rect -1191 -9730 -477 -9720
rect -1263 -9746 -477 -9730
rect -1263 -9782 -549 -9746
rect -1263 -9828 -1237 -9782
rect -1191 -9792 -549 -9782
rect -503 -9792 -477 -9746
rect -1191 -9828 -477 -9792
rect 1190 -9694 1215 -9648
rect 1261 -9694 1287 -9648
rect 1190 -9737 1287 -9694
rect 1381 -9737 1496 -9537
rect 1611 -9570 1708 -9537
rect 1885 -9461 2708 -9440
rect 1885 -9463 2066 -9461
rect 1885 -9501 1921 -9463
rect 1985 -9500 2066 -9463
rect 1885 -9553 1898 -9501
rect 1985 -9527 2004 -9500
rect 1950 -9552 2004 -9527
rect 2056 -9525 2066 -9500
rect 2130 -9525 2200 -9461
rect 2264 -9499 2708 -9461
rect 2264 -9500 2322 -9499
rect 2056 -9552 2216 -9525
rect 2268 -9551 2322 -9500
rect 2374 -9501 2708 -9499
rect 2374 -9502 2643 -9501
rect 2374 -9551 2537 -9502
rect 2268 -9552 2537 -9551
rect 1950 -9553 2537 -9552
rect 1885 -9554 2537 -9553
rect 2589 -9553 2643 -9502
rect 2695 -9553 2708 -9501
rect 2589 -9554 2708 -9553
rect 1885 -9566 2708 -9554
rect 2884 -9446 8786 -9420
rect 8832 -9446 8858 -9400
rect 2884 -9472 8858 -9446
rect 2884 -9518 2910 -9472
rect 2956 -9498 8858 -9472
rect 2956 -9518 8786 -9498
rect 2884 -9544 8786 -9518
rect 8832 -9544 8858 -9498
rect 1611 -9616 1636 -9570
rect 1682 -9616 1708 -9570
rect 1611 -9668 1708 -9616
rect 1611 -9714 1636 -9668
rect 1682 -9714 1708 -9668
rect 1611 -9737 1708 -9714
rect 1190 -9746 1708 -9737
rect 1190 -9792 1215 -9746
rect 1261 -9766 1708 -9746
rect 1261 -9792 1636 -9766
rect 1190 -9812 1636 -9792
rect 1682 -9812 1708 -9766
rect -1263 -9844 -477 -9828
rect -1263 -9880 -549 -9844
rect -1263 -9926 -1237 -9880
rect -1191 -9890 -549 -9880
rect -503 -9890 -477 -9844
rect -1191 -9920 -477 -9890
rect -1191 -9926 -1166 -9920
rect -1263 -9978 -1166 -9926
rect -1263 -10024 -1237 -9978
rect -1191 -10024 -1166 -9978
rect -1263 -10076 -1166 -10024
rect -1263 -10122 -1237 -10076
rect -1191 -10120 -1166 -10076
rect -1011 -10120 -765 -9920
rect -574 -9942 -477 -9920
rect -574 -9988 -549 -9942
rect -503 -9988 -477 -9942
rect 299 -9835 382 -9819
rect 299 -9907 313 -9835
rect 369 -9907 382 -9835
rect 299 -9970 382 -9907
rect -574 -10040 -477 -9988
rect -574 -10086 -549 -10040
rect -503 -10086 -477 -10040
rect -574 -10120 -477 -10086
rect -1191 -10122 -477 -10120
rect -1609 -10135 -1563 -10124
rect -1449 -10135 -1403 -10124
rect -1263 -10138 -477 -10122
rect -1263 -10174 -549 -10138
rect -1263 -10220 -1237 -10174
rect -1191 -10184 -549 -10174
rect -503 -10184 -477 -10138
rect -184 -9998 -99 -9980
rect -184 -10054 -169 -9998
rect -113 -10054 -99 -9998
rect -184 -10112 -99 -10054
rect 299 -10042 313 -9970
rect 369 -10042 382 -9970
rect 299 -10055 382 -10042
rect 1190 -9844 1708 -9812
rect 1190 -9890 1215 -9844
rect 1261 -9864 1708 -9844
rect 1261 -9890 1636 -9864
rect 1190 -9910 1636 -9890
rect 1682 -9910 1708 -9864
rect 1190 -9937 1708 -9910
rect 1190 -9942 1287 -9937
rect 1190 -9988 1215 -9942
rect 1261 -9988 1287 -9942
rect 1190 -10040 1287 -9988
rect -184 -10168 -169 -10112
rect -113 -10168 -99 -10112
rect -184 -10184 -99 -10168
rect 1190 -10086 1215 -10040
rect 1261 -10086 1287 -10040
rect 1190 -10137 1287 -10086
rect 1381 -10137 1496 -9937
rect 1611 -9962 1708 -9937
rect 1611 -10008 1636 -9962
rect 1682 -10008 1708 -9962
rect 1611 -10060 1708 -10008
rect 1611 -10106 1636 -10060
rect 1682 -10106 1708 -10060
rect 1611 -10137 1708 -10106
rect 1190 -10138 1708 -10137
rect 1190 -10184 1215 -10138
rect 1261 -10158 1708 -10138
rect 1261 -10184 1636 -10158
rect -1191 -10220 -477 -10184
rect -1263 -10236 -477 -10220
rect -1263 -10272 -549 -10236
rect -1263 -10318 -1237 -10272
rect -1191 -10282 -549 -10272
rect -503 -10282 -477 -10236
rect 1190 -10204 1636 -10184
rect 1682 -10204 1708 -10158
rect 1190 -10236 1708 -10204
rect -1191 -10318 -477 -10282
rect -1263 -10320 -477 -10318
rect -1263 -10344 -1166 -10320
rect -3321 -10370 -1166 -10344
rect -3321 -10416 -3295 -10370
rect -3249 -10416 -3197 -10370
rect -3151 -10416 -3099 -10370
rect -3053 -10416 -3001 -10370
rect -2955 -10416 -2903 -10370
rect -2857 -10416 -2805 -10370
rect -2759 -10416 -2707 -10370
rect -2661 -10416 -2609 -10370
rect -2563 -10416 -2511 -10370
rect -2465 -10416 -2413 -10370
rect -2367 -10416 -2315 -10370
rect -2269 -10416 -2217 -10370
rect -2171 -10416 -2119 -10370
rect -2073 -10416 -2021 -10370
rect -1975 -10416 -1923 -10370
rect -1877 -10416 -1825 -10370
rect -1779 -10416 -1727 -10370
rect -1681 -10416 -1629 -10370
rect -1583 -10416 -1531 -10370
rect -1485 -10416 -1433 -10370
rect -1387 -10416 -1335 -10370
rect -1289 -10416 -1237 -10370
rect -1191 -10416 -1166 -10370
rect -3321 -10441 -1166 -10416
rect -3321 -10694 -1321 -10441
rect -1011 -10694 -765 -10320
rect -574 -10334 -477 -10320
rect -574 -10380 -549 -10334
rect -503 -10380 -477 -10334
rect -324 -10321 -278 -10237
rect -164 -10321 -118 -10254
rect -324 -10367 -246 -10321
rect -200 -10367 -118 -10321
rect -574 -10432 -477 -10380
rect -574 -10478 -549 -10432
rect -503 -10478 -477 -10432
rect -574 -10530 -477 -10478
rect -164 -10481 -118 -10367
rect -4 -10369 42 -10260
rect 444 -10364 546 -10351
rect 444 -10369 460 -10364
rect -4 -10415 460 -10369
rect 444 -10420 460 -10415
rect 532 -10369 546 -10364
rect 638 -10369 684 -10260
rect 532 -10415 684 -10369
rect 798 -10328 844 -10260
rect 958 -10318 1004 -10259
rect 1190 -10282 1215 -10236
rect 1261 -10256 1708 -10236
rect 1261 -10282 1636 -10256
rect 1190 -10302 1636 -10282
rect 1682 -10302 1708 -10256
rect 944 -10328 1011 -10318
rect 798 -10329 1011 -10328
rect 798 -10375 957 -10329
rect 1003 -10375 1011 -10329
rect 798 -10376 1011 -10375
rect 532 -10420 546 -10415
rect 444 -10434 546 -10420
rect 798 -10481 844 -10376
rect 944 -10388 1011 -10376
rect 1190 -10328 1708 -10302
rect 1783 -10328 1849 -9615
rect 1943 -10216 2009 -9566
rect 2103 -10328 2169 -9615
rect 2262 -10215 2328 -9566
rect 2423 -10328 2489 -9614
rect 2583 -10215 2649 -9566
rect 2884 -9568 8858 -9544
rect 2884 -9570 2981 -9568
rect 2742 -10328 2808 -9615
rect 2884 -9616 2910 -9570
rect 2956 -9616 2981 -9570
rect 2884 -9668 2981 -9616
rect 2884 -9714 2910 -9668
rect 2956 -9714 2981 -9668
rect 2884 -9766 2981 -9714
rect 2884 -9812 2910 -9766
rect 2956 -9812 2981 -9766
rect 2884 -9864 2981 -9812
rect 2884 -9910 2910 -9864
rect 2956 -9879 2981 -9864
rect 3259 -9879 3459 -9568
rect 3659 -9879 3859 -9568
rect 4437 -9596 8858 -9568
rect 4437 -9642 8786 -9596
rect 8832 -9642 8858 -9596
rect 4437 -9663 8858 -9642
rect 4437 -9879 4696 -9663
rect 6080 -9879 6620 -9663
rect 8298 -9879 8562 -9663
rect 8760 -9694 8858 -9663
rect 8760 -9740 8786 -9694
rect 8832 -9740 8858 -9694
rect 8760 -9792 8858 -9740
rect 8760 -9838 8786 -9792
rect 8832 -9838 8858 -9792
rect 8760 -9879 8858 -9838
rect 2956 -9890 8858 -9879
rect 2956 -9910 8786 -9890
rect 2884 -9936 8786 -9910
rect 8832 -9936 8858 -9890
rect 2884 -9962 8858 -9936
rect 2884 -10008 2910 -9962
rect 2956 -9988 8858 -9962
rect 2956 -10008 8786 -9988
rect 2884 -10034 8786 -10008
rect 8832 -10034 8858 -9988
rect 2884 -10060 8858 -10034
rect 2884 -10106 2910 -10060
rect 2956 -10086 8858 -10060
rect 2956 -10106 8786 -10086
rect 2884 -10132 8786 -10106
rect 8832 -10132 8858 -10086
rect 2884 -10138 8858 -10132
rect 2884 -10158 2981 -10138
rect 2884 -10204 2910 -10158
rect 2956 -10204 2981 -10158
rect 2884 -10256 2981 -10204
rect 2884 -10302 2910 -10256
rect 2956 -10302 2981 -10256
rect 2884 -10328 2981 -10302
rect 1190 -10334 2981 -10328
rect 1190 -10380 1215 -10334
rect 1261 -10337 2981 -10334
rect 1261 -10380 1287 -10337
rect -164 -10527 844 -10481
rect 1190 -10432 1287 -10380
rect 1611 -10354 2981 -10337
rect 1611 -10400 1636 -10354
rect 1682 -10400 1734 -10354
rect 1780 -10400 1832 -10354
rect 1878 -10400 1930 -10354
rect 1976 -10400 2028 -10354
rect 2074 -10400 2126 -10354
rect 2172 -10400 2224 -10354
rect 2270 -10400 2322 -10354
rect 2368 -10400 2420 -10354
rect 2466 -10400 2518 -10354
rect 2564 -10400 2616 -10354
rect 2662 -10400 2714 -10354
rect 2760 -10400 2812 -10354
rect 2858 -10400 2910 -10354
rect 2956 -10400 2981 -10354
rect 3259 -10400 3459 -10138
rect 3659 -10400 3859 -10138
rect 4437 -10400 4696 -10138
rect 6080 -10400 6620 -10138
rect 8298 -10400 8562 -10138
rect 8760 -10184 8858 -10138
rect 8760 -10230 8786 -10184
rect 8832 -10230 8858 -10184
rect 8760 -10282 8858 -10230
rect 8760 -10328 8786 -10282
rect 8832 -10328 8858 -10282
rect 8760 -10380 8858 -10328
rect 8760 -10400 8786 -10380
rect 1611 -10425 8786 -10400
rect 1190 -10478 1215 -10432
rect 1261 -10478 1287 -10432
rect -574 -10576 -549 -10530
rect -503 -10576 -477 -10530
rect -574 -10602 -477 -10576
rect 1190 -10530 1287 -10478
rect 1190 -10576 1215 -10530
rect 1261 -10576 1287 -10530
rect 1190 -10602 1287 -10576
rect -574 -10628 1287 -10602
rect -574 -10674 -549 -10628
rect -503 -10674 -451 -10628
rect -405 -10674 -353 -10628
rect -307 -10674 -255 -10628
rect -209 -10674 -157 -10628
rect -111 -10674 -59 -10628
rect -13 -10674 39 -10628
rect 85 -10674 137 -10628
rect 183 -10674 235 -10628
rect 281 -10674 333 -10628
rect 379 -10674 431 -10628
rect 477 -10674 529 -10628
rect 575 -10674 627 -10628
rect 673 -10674 725 -10628
rect 771 -10674 823 -10628
rect 869 -10674 921 -10628
rect 967 -10674 1019 -10628
rect 1065 -10674 1117 -10628
rect 1163 -10674 1215 -10628
rect 1261 -10674 1287 -10628
rect -574 -10694 1287 -10674
rect 1739 -10426 8786 -10425
rect 8832 -10426 8858 -10380
rect 1739 -10452 8858 -10426
rect 8945 -8742 9006 -7806
rect 9104 -8742 9165 -7806
rect 9246 -7967 9336 -7955
rect 9246 -8034 9259 -7967
rect 9324 -8034 9336 -7967
rect 9246 -8046 9336 -8034
rect 9264 -8319 9325 -8110
rect 9246 -8333 9343 -8319
rect 9246 -8397 9262 -8333
rect 9326 -8397 9343 -8333
rect 9246 -8449 9343 -8397
rect 9246 -8513 9262 -8449
rect 9326 -8513 9343 -8449
rect 9246 -8531 9343 -8513
rect 8945 -8754 9165 -8742
rect 8945 -8805 9029 -8754
rect 9080 -8805 9165 -8754
rect 8945 -8817 9165 -8805
rect 8945 -9479 9006 -8817
rect 9104 -9479 9165 -8817
rect 9264 -9045 9325 -8531
rect 9248 -9059 9345 -9045
rect 9248 -9123 9264 -9059
rect 9328 -9123 9345 -9059
rect 9248 -9175 9345 -9123
rect 9248 -9239 9264 -9175
rect 9328 -9239 9345 -9175
rect 9248 -9257 9345 -9239
rect 8945 -9491 9165 -9479
rect 8945 -9542 9029 -9491
rect 9080 -9542 9165 -9491
rect 8945 -9554 9165 -9542
rect 8945 -10452 9006 -9554
rect 9104 -10452 9165 -9554
rect 9264 -9776 9325 -9257
rect 9246 -9790 9343 -9776
rect 9246 -9854 9262 -9790
rect 9326 -9854 9343 -9790
rect 9246 -9906 9343 -9854
rect 9246 -9970 9262 -9906
rect 9326 -9970 9343 -9906
rect 9246 -9988 9343 -9970
rect 9264 -10183 9325 -9988
rect 9245 -10258 9335 -10246
rect 9245 -10325 9258 -10258
rect 9323 -10325 9335 -10258
rect 9245 -10337 9335 -10325
rect 9424 -10452 9485 -7806
rect 9560 -7966 9650 -7954
rect 9560 -8033 9573 -7966
rect 9638 -8033 9650 -7966
rect 9560 -8045 9650 -8033
rect 9585 -8319 9646 -8111
rect 9566 -8333 9663 -8319
rect 9566 -8397 9582 -8333
rect 9646 -8397 9663 -8333
rect 9566 -8449 9663 -8397
rect 9566 -8513 9582 -8449
rect 9646 -8513 9663 -8449
rect 9566 -8531 9663 -8513
rect 9585 -9047 9646 -8531
rect 9568 -9061 9665 -9047
rect 9568 -9125 9584 -9061
rect 9648 -9125 9665 -9061
rect 9568 -9177 9665 -9125
rect 9568 -9241 9584 -9177
rect 9648 -9241 9665 -9177
rect 9568 -9259 9665 -9241
rect 9585 -9776 9646 -9259
rect 9568 -9790 9665 -9776
rect 9568 -9854 9584 -9790
rect 9648 -9854 9665 -9790
rect 9568 -9906 9665 -9854
rect 9568 -9970 9584 -9906
rect 9648 -9970 9665 -9906
rect 9568 -9988 9665 -9970
rect 9585 -10183 9646 -9988
rect 9573 -10255 9663 -10243
rect 9573 -10322 9586 -10255
rect 9651 -10322 9663 -10255
rect 9573 -10334 9663 -10322
rect 9745 -10452 9806 -7806
rect 9877 -7963 9967 -7951
rect 9877 -8030 9890 -7963
rect 9955 -8030 9967 -7963
rect 9877 -8042 9967 -8030
rect 9904 -8319 9965 -8111
rect 9887 -8333 9984 -8319
rect 9887 -8397 9903 -8333
rect 9967 -8397 9984 -8333
rect 9887 -8449 9984 -8397
rect 9887 -8513 9903 -8449
rect 9967 -8513 9984 -8449
rect 9887 -8531 9984 -8513
rect 9904 -9049 9965 -8531
rect 9888 -9063 9985 -9049
rect 9888 -9127 9904 -9063
rect 9968 -9127 9985 -9063
rect 9888 -9179 9985 -9127
rect 9888 -9243 9904 -9179
rect 9968 -9243 9985 -9179
rect 9888 -9261 9985 -9243
rect 9904 -9776 9965 -9261
rect 9887 -9790 9984 -9776
rect 9887 -9854 9903 -9790
rect 9967 -9854 9984 -9790
rect 9887 -9906 9984 -9854
rect 9887 -9970 9903 -9906
rect 9967 -9970 9984 -9906
rect 9887 -9988 9984 -9970
rect 9904 -10183 9965 -9988
rect 9883 -10256 9973 -10244
rect 9883 -10323 9896 -10256
rect 9961 -10323 9973 -10256
rect 9883 -10335 9973 -10323
rect 10064 -10452 10125 -7806
rect 10208 -7962 10298 -7950
rect 10208 -8029 10221 -7962
rect 10286 -8029 10298 -7962
rect 10208 -8041 10298 -8029
rect 10224 -8322 10285 -8110
rect 10207 -8336 10304 -8322
rect 10207 -8400 10223 -8336
rect 10287 -8400 10304 -8336
rect 10207 -8452 10304 -8400
rect 10207 -8516 10223 -8452
rect 10287 -8516 10304 -8452
rect 10207 -8534 10304 -8516
rect 10224 -9049 10285 -8534
rect 10208 -9063 10305 -9049
rect 10208 -9127 10224 -9063
rect 10288 -9127 10305 -9063
rect 10208 -9179 10305 -9127
rect 10208 -9243 10224 -9179
rect 10288 -9243 10305 -9179
rect 10208 -9261 10305 -9243
rect 10224 -9778 10285 -9261
rect 10207 -9792 10304 -9778
rect 10207 -9856 10223 -9792
rect 10287 -9856 10304 -9792
rect 10207 -9908 10304 -9856
rect 10207 -9972 10223 -9908
rect 10287 -9972 10304 -9908
rect 10207 -9990 10304 -9972
rect 10224 -10181 10285 -9990
rect 10209 -10256 10299 -10244
rect 10209 -10323 10222 -10256
rect 10287 -10323 10299 -10256
rect 10209 -10335 10299 -10323
rect 10384 -10452 10445 -7806
rect 10527 -7963 10617 -7951
rect 10527 -8030 10540 -7963
rect 10605 -8030 10617 -7963
rect 10527 -8042 10617 -8030
rect 10544 -8320 10605 -8111
rect 10527 -8334 10624 -8320
rect 10527 -8398 10543 -8334
rect 10607 -8398 10624 -8334
rect 10527 -8450 10624 -8398
rect 10527 -8514 10543 -8450
rect 10607 -8514 10624 -8450
rect 10527 -8532 10624 -8514
rect 10544 -9049 10605 -8532
rect 10704 -8743 10765 -7806
rect 10864 -8743 10925 -7806
rect 10704 -8755 10925 -8743
rect 10704 -8806 10788 -8755
rect 10839 -8806 10925 -8755
rect 10704 -8818 10925 -8806
rect 10525 -9063 10622 -9049
rect 10525 -9127 10541 -9063
rect 10605 -9127 10622 -9063
rect 10525 -9179 10622 -9127
rect 10525 -9243 10541 -9179
rect 10605 -9243 10622 -9179
rect 10525 -9261 10622 -9243
rect 10544 -9778 10605 -9261
rect 10704 -9479 10765 -8818
rect 10864 -9479 10925 -8818
rect 10704 -9491 10925 -9479
rect 10704 -9542 10788 -9491
rect 10839 -9542 10925 -9491
rect 10704 -9554 10925 -9542
rect 10527 -9792 10624 -9778
rect 10527 -9856 10543 -9792
rect 10607 -9856 10624 -9792
rect 10527 -9908 10624 -9856
rect 10527 -9972 10543 -9908
rect 10607 -9972 10624 -9908
rect 10527 -9990 10624 -9972
rect 10544 -10183 10605 -9990
rect 10524 -10252 10614 -10240
rect 10524 -10319 10537 -10252
rect 10602 -10319 10614 -10252
rect 10524 -10331 10614 -10319
rect 10704 -10452 10765 -9554
rect 10864 -10452 10925 -9554
rect 11014 -7832 11112 -7806
rect 11014 -7878 11040 -7832
rect 11086 -7878 11112 -7832
rect 11014 -7930 11112 -7878
rect 11014 -7976 11040 -7930
rect 11086 -7976 11112 -7930
rect 11014 -8028 11112 -7976
rect 11014 -8074 11040 -8028
rect 11086 -8074 11112 -8028
rect 11014 -8126 11112 -8074
rect 11014 -8172 11040 -8126
rect 11086 -8172 11112 -8126
rect 11014 -8224 11112 -8172
rect 11014 -8270 11040 -8224
rect 11086 -8270 11112 -8224
rect 11014 -8322 11112 -8270
rect 11014 -8368 11040 -8322
rect 11086 -8368 11112 -8322
rect 11014 -8420 11112 -8368
rect 11014 -8466 11040 -8420
rect 11086 -8466 11112 -8420
rect 11014 -8518 11112 -8466
rect 11014 -8564 11040 -8518
rect 11086 -8564 11112 -8518
rect 11014 -8616 11112 -8564
rect 11014 -8662 11040 -8616
rect 11086 -8662 11112 -8616
rect 11014 -8714 11112 -8662
rect 11014 -8760 11040 -8714
rect 11086 -8760 11112 -8714
rect 11014 -8812 11112 -8760
rect 11014 -8858 11040 -8812
rect 11086 -8858 11112 -8812
rect 11014 -8910 11112 -8858
rect 11014 -8956 11040 -8910
rect 11086 -8956 11112 -8910
rect 11014 -9008 11112 -8956
rect 11014 -9054 11040 -9008
rect 11086 -9054 11112 -9008
rect 11014 -9106 11112 -9054
rect 11014 -9152 11040 -9106
rect 11086 -9152 11112 -9106
rect 11014 -9204 11112 -9152
rect 11014 -9250 11040 -9204
rect 11086 -9250 11112 -9204
rect 11014 -9302 11112 -9250
rect 11014 -9348 11040 -9302
rect 11086 -9348 11112 -9302
rect 11014 -9400 11112 -9348
rect 11014 -9446 11040 -9400
rect 11086 -9446 11112 -9400
rect 11014 -9498 11112 -9446
rect 11014 -9544 11040 -9498
rect 11086 -9544 11112 -9498
rect 11014 -9596 11112 -9544
rect 11014 -9642 11040 -9596
rect 11086 -9642 11112 -9596
rect 11014 -9694 11112 -9642
rect 11014 -9740 11040 -9694
rect 11086 -9740 11112 -9694
rect 11014 -9792 11112 -9740
rect 11014 -9838 11040 -9792
rect 11086 -9838 11112 -9792
rect 11014 -9890 11112 -9838
rect 11014 -9936 11040 -9890
rect 11086 -9936 11112 -9890
rect 11014 -9988 11112 -9936
rect 11014 -10034 11040 -9988
rect 11086 -10034 11112 -9988
rect 11014 -10086 11112 -10034
rect 11014 -10132 11040 -10086
rect 11086 -10132 11112 -10086
rect 11014 -10184 11112 -10132
rect 11014 -10230 11040 -10184
rect 11086 -10230 11112 -10184
rect 11014 -10282 11112 -10230
rect 11014 -10328 11040 -10282
rect 11086 -10328 11112 -10282
rect 11014 -10380 11112 -10328
rect 11014 -10426 11040 -10380
rect 11086 -10426 11112 -10380
rect 11014 -10452 11112 -10426
rect 1739 -10478 11112 -10452
rect 1739 -10524 8786 -10478
rect 8832 -10524 8884 -10478
rect 8930 -10524 8982 -10478
rect 9028 -10524 9080 -10478
rect 9126 -10524 9178 -10478
rect 9224 -10524 9276 -10478
rect 9322 -10524 9374 -10478
rect 9420 -10524 9472 -10478
rect 9518 -10524 9570 -10478
rect 9616 -10524 9668 -10478
rect 9714 -10524 9766 -10478
rect 9812 -10524 9864 -10478
rect 9910 -10524 9962 -10478
rect 10008 -10524 10060 -10478
rect 10106 -10524 10158 -10478
rect 10204 -10524 10256 -10478
rect 10302 -10524 10354 -10478
rect 10400 -10524 10452 -10478
rect 10498 -10524 10550 -10478
rect 10596 -10524 10648 -10478
rect 10694 -10524 10746 -10478
rect 10792 -10524 10844 -10478
rect 10890 -10524 10942 -10478
rect 10988 -10524 11040 -10478
rect 11086 -10524 11112 -10478
rect 1739 -10550 11112 -10524
rect 1739 -10694 11084 -10550
rect -3321 -10940 11084 -10694
<< via1 >>
rect -2775 -1845 -2691 -1762
rect -2416 1262 -2364 1266
rect -2416 1216 -2413 1262
rect -2413 1216 -2367 1262
rect -2367 1216 -2364 1262
rect -2416 1213 -2364 1216
rect -2304 1263 -2252 1266
rect -2304 1217 -2258 1263
rect -2258 1217 -2252 1263
rect -2304 1213 -2252 1217
rect -2343 -1843 -2259 -1760
rect 191 457 271 535
rect -244 233 -162 323
rect -242 -145 -160 -66
rect 625 237 700 311
rect -242 -535 -160 -456
rect -1910 -1843 -1826 -1760
rect -4042 -2591 -3919 -2471
rect -3842 -2591 -3719 -2471
rect -4039 -2843 -3916 -2723
rect -3839 -2843 -3716 -2723
rect -1734 -2747 -1654 -2730
rect -1734 -2793 -1708 -2747
rect -1708 -2793 -1662 -2747
rect -1662 -2793 -1654 -2747
rect -1734 -2810 -1654 -2793
rect -2599 -3034 -2531 -2953
rect -1963 -3036 -1895 -2955
rect -2759 -3190 -2691 -3109
rect -2439 -3182 -2371 -3101
rect -2118 -3190 -2050 -3109
rect -1803 -3186 -1735 -3105
rect 621 -150 703 -71
rect 623 -534 705 -455
rect 270 -1188 353 -1109
rect 185 -2235 266 -2154
rect -243 -3197 -163 -3117
rect -3079 -3341 -3011 -3260
rect -2922 -3343 -2854 -3262
rect -2279 -3342 -2211 -3261
rect -1643 -3345 -1575 -3264
rect -1477 -3341 -1409 -3260
rect -2844 -3580 -2762 -3549
rect -2844 -3626 -2829 -3580
rect -2829 -3626 -2783 -3580
rect -2783 -3626 -2762 -3580
rect -2844 -3629 -2762 -3626
rect -2600 -3892 -2532 -3811
rect -1957 -3886 -1889 -3805
rect 189 -3200 271 -3117
rect 620 -3196 704 -3110
rect 2843 579 2907 643
rect 2843 463 2907 527
rect 2843 -161 2907 -97
rect 2843 -277 2907 -213
rect 2843 -924 2907 -860
rect 2843 -1040 2907 -976
rect 2843 -1653 2907 -1589
rect 2843 -1769 2907 -1705
rect 2843 -2371 2907 -2307
rect 2843 -2487 2907 -2423
rect 3163 577 3227 641
rect 3163 461 3227 525
rect 3163 -163 3227 -99
rect 3163 -279 3227 -215
rect 3163 -892 3227 -828
rect 3163 -1008 3227 -944
rect 3163 -1632 3227 -1568
rect 3163 -1748 3227 -1684
rect 3163 -2372 3227 -2308
rect 3163 -2488 3227 -2424
rect 3483 607 3547 671
rect 3483 491 3547 555
rect 3483 -144 3547 -80
rect 3483 -260 3547 -196
rect 3483 -876 3547 -812
rect 3483 -992 3547 -928
rect 3483 -1618 3547 -1554
rect 3483 -1734 3547 -1670
rect 3483 -2378 3547 -2314
rect 3483 -2494 3547 -2430
rect 3803 594 3867 658
rect 3803 478 3867 542
rect 3803 -165 3867 -101
rect 3803 -281 3867 -217
rect 3803 -901 3867 -837
rect 3803 -1017 3867 -953
rect 3803 -1626 3867 -1562
rect 3803 -1742 3867 -1678
rect 3803 -2374 3867 -2310
rect 3803 -2490 3867 -2426
rect 4123 591 4187 655
rect 4123 475 4187 539
rect 4123 -180 4187 -116
rect 4123 -296 4187 -232
rect 4123 -905 4187 -841
rect 4123 -1021 4187 -957
rect 4123 -1629 4187 -1565
rect 4123 -1745 4187 -1681
rect 4123 -2377 4187 -2313
rect 4123 -2493 4187 -2429
rect 5643 579 5707 643
rect 5643 463 5707 527
rect 5643 -161 5707 -97
rect 5643 -277 5707 -213
rect 5643 -924 5707 -860
rect 5643 -1040 5707 -976
rect 5643 -1653 5707 -1589
rect 5643 -1769 5707 -1705
rect 5643 -2371 5707 -2307
rect 5643 -2487 5707 -2423
rect 5963 577 6027 641
rect 5963 461 6027 525
rect 5963 -163 6027 -99
rect 5963 -279 6027 -215
rect 5963 -892 6027 -828
rect 5963 -1008 6027 -944
rect 5963 -1632 6027 -1568
rect 5963 -1748 6027 -1684
rect 5963 -2372 6027 -2308
rect 5963 -2488 6027 -2424
rect 6283 607 6347 671
rect 6283 491 6347 555
rect 6283 -144 6347 -80
rect 6283 -260 6347 -196
rect 6283 -876 6347 -812
rect 6283 -992 6347 -928
rect 6283 -1618 6347 -1554
rect 6283 -1734 6347 -1670
rect 6283 -2378 6347 -2314
rect 6283 -2494 6347 -2430
rect 6603 594 6667 658
rect 6603 478 6667 542
rect 6603 -165 6667 -101
rect 6603 -281 6667 -217
rect 6603 -901 6667 -837
rect 6603 -1017 6667 -953
rect 6603 -1626 6667 -1562
rect 6603 -1742 6667 -1678
rect 6603 -2374 6667 -2310
rect 6603 -2490 6667 -2426
rect 6923 591 6987 655
rect 6923 475 6987 539
rect 6923 -180 6987 -116
rect 6923 -296 6987 -232
rect 6923 -905 6987 -841
rect 6923 -1021 6987 -957
rect 6923 -1629 6987 -1565
rect 6923 -1745 6987 -1681
rect 6923 -2377 6987 -2313
rect 6923 -2493 6987 -2429
rect 8443 579 8507 643
rect 8443 463 8507 527
rect 8443 -161 8507 -97
rect 8443 -277 8507 -213
rect 8443 -924 8507 -860
rect 8443 -1040 8507 -976
rect 8443 -1653 8507 -1589
rect 8443 -1769 8507 -1705
rect 8443 -2371 8507 -2307
rect 8443 -2487 8507 -2423
rect 8763 577 8827 641
rect 8763 461 8827 525
rect 8763 -163 8827 -99
rect 8763 -279 8827 -215
rect 8763 -892 8827 -828
rect 8763 -1008 8827 -944
rect 8763 -1632 8827 -1568
rect 8763 -1748 8827 -1684
rect 8763 -2372 8827 -2308
rect 8763 -2488 8827 -2424
rect 9083 607 9147 671
rect 9083 491 9147 555
rect 9083 -144 9147 -80
rect 9083 -260 9147 -196
rect 9083 -876 9147 -812
rect 9083 -992 9147 -928
rect 9083 -1618 9147 -1554
rect 9083 -1734 9147 -1670
rect 9083 -2378 9147 -2314
rect 9083 -2494 9147 -2430
rect 9403 594 9467 658
rect 9403 478 9467 542
rect 9403 -165 9467 -101
rect 9403 -281 9467 -217
rect 9403 -901 9467 -837
rect 9403 -1017 9467 -953
rect 9403 -1626 9467 -1562
rect 9403 -1742 9467 -1678
rect 9403 -2374 9467 -2310
rect 9403 -2490 9467 -2426
rect 9723 591 9787 655
rect 9723 475 9787 539
rect 9723 -180 9787 -116
rect 9723 -296 9787 -232
rect 9723 -905 9787 -841
rect 9723 -1021 9787 -957
rect 9723 -1629 9787 -1565
rect 9723 -1745 9787 -1681
rect 9723 -2377 9787 -2313
rect 9723 -2493 9787 -2429
rect 11088 -1335 11169 -1254
rect 11228 -1335 11309 -1254
rect 11368 -1335 11449 -1254
rect 11508 -1335 11589 -1254
rect 11648 -1335 11729 -1254
rect 11094 -2764 11175 -2683
rect 11234 -2764 11315 -2683
rect 11374 -2764 11455 -2683
rect 11514 -2764 11595 -2683
rect 11654 -2764 11735 -2683
rect -245 -3649 -161 -3563
rect 477 -3651 561 -3565
rect 621 -3651 705 -3565
rect 1364 -3661 1473 -3557
rect -2757 -4042 -2689 -3961
rect -2440 -4047 -2372 -3966
rect -2120 -4042 -2052 -3961
rect -1800 -4040 -1732 -3959
rect 25 -3847 109 -3761
rect 184 -3848 268 -3762
rect 1565 -3858 1675 -3753
rect -3080 -4200 -3012 -4119
rect -2923 -4203 -2855 -4122
rect -2280 -4204 -2212 -4123
rect -1643 -4201 -1575 -4120
rect -1478 -4199 -1410 -4118
rect -1737 -4478 -1650 -4393
rect -261 -4246 -197 -4245
rect -261 -4304 -230 -4246
rect -230 -4304 -197 -4246
rect -145 -4248 -81 -4245
rect -145 -4303 -90 -4248
rect -90 -4303 -81 -4248
rect -261 -4309 -197 -4304
rect -145 -4309 -81 -4303
rect 189 -4292 266 -4220
rect -2600 -4742 -2532 -4661
rect -1961 -4746 -1893 -4665
rect -2760 -4900 -2692 -4819
rect -2442 -4904 -2374 -4823
rect -2116 -4898 -2048 -4817
rect -1802 -4909 -1734 -4828
rect -3077 -5050 -3009 -4969
rect -2920 -5053 -2852 -4972
rect -2280 -5055 -2212 -4974
rect -1636 -5056 -1568 -4975
rect -1479 -5052 -1411 -4971
rect -2845 -5260 -2759 -5252
rect -2845 -5306 -2829 -5260
rect -2829 -5306 -2783 -5260
rect -2783 -5306 -2759 -5260
rect -2845 -5337 -2759 -5306
rect -2598 -5609 -2530 -5528
rect -1955 -5608 -1887 -5527
rect -2763 -5760 -2695 -5679
rect -2441 -5759 -2373 -5678
rect -2126 -5767 -2058 -5686
rect -1797 -5765 -1729 -5684
rect -3077 -5925 -3009 -5844
rect -2915 -5923 -2847 -5842
rect -2279 -5918 -2211 -5837
rect -1644 -5918 -1576 -5837
rect -1476 -5920 -1408 -5839
rect -1731 -6093 -1651 -6076
rect -1731 -6139 -1708 -6093
rect -1708 -6139 -1662 -6093
rect -1662 -6139 -1651 -6093
rect -1731 -6156 -1651 -6139
rect 355 -4415 434 -4336
rect 353 -6024 435 -5939
rect 811 -4916 875 -4852
rect 811 -5032 875 -4968
rect 810 -5597 874 -5533
rect 810 -5713 874 -5649
rect -109 -6137 -27 -6052
rect 50 -6134 132 -6049
rect 2208 -4864 2272 -4800
rect 2208 -4980 2272 -4916
rect 2579 -4543 2643 -4479
rect 2719 -4543 2783 -4479
rect 2579 -4655 2583 -4595
rect 2583 -4655 2643 -4595
rect 2719 -4655 2773 -4595
rect 2773 -4655 2783 -4595
rect 2579 -4659 2643 -4655
rect 2719 -4659 2783 -4655
rect 3070 -4873 3134 -4809
rect 3070 -4989 3134 -4925
rect 2290 -5941 2354 -5877
rect 2290 -6057 2354 -5993
rect 2846 -5586 2910 -5522
rect 2846 -5702 2910 -5638
rect 3018 -5919 3082 -5890
rect 3018 -5954 3075 -5919
rect 3075 -5954 3082 -5919
rect 3018 -6070 3082 -6006
rect 4807 -4991 4871 -4927
rect 4807 -5107 4871 -5043
rect 4807 -5510 4871 -5446
rect 4807 -5626 4871 -5562
rect 5411 -5472 5475 -5408
rect 5411 -5588 5475 -5524
rect 5859 -4988 5923 -4924
rect 5859 -5104 5923 -5040
rect 5859 -5507 5923 -5443
rect 5859 -5623 5923 -5559
rect -2004 -6550 -1908 -6460
rect -2605 -6675 -2509 -6585
rect -3061 -7293 -2993 -7212
rect -2897 -7292 -2829 -7211
rect -3060 -8099 -2992 -8018
rect -2901 -8103 -2833 -8022
rect -3062 -8899 -2994 -8818
rect -2903 -8899 -2835 -8818
rect -3060 -9697 -2992 -9616
rect -2898 -9696 -2830 -9615
rect -2582 -7612 -2514 -7531
rect -2589 -8414 -2507 -8332
rect -2591 -9215 -2509 -9133
rect -2581 -10012 -2513 -9931
rect -2259 -7293 -2191 -7212
rect -2256 -7815 -2196 -7809
rect -2256 -7864 -2251 -7815
rect -2251 -7864 -2202 -7815
rect -2202 -7864 -2196 -7815
rect -2256 -7869 -2196 -7864
rect -2258 -8097 -2190 -8016
rect -2256 -8616 -2196 -8610
rect -2256 -8665 -2251 -8616
rect -2251 -8665 -2202 -8616
rect -2202 -8665 -2196 -8616
rect -2256 -8670 -2196 -8665
rect -2261 -8897 -2193 -8816
rect -2257 -9416 -2197 -9410
rect -2257 -9465 -2252 -9416
rect -2252 -9465 -2203 -9416
rect -2203 -9465 -2197 -9416
rect -2257 -9470 -2197 -9465
rect -2260 -9697 -2192 -9616
rect -1949 -7612 -1867 -7530
rect -1940 -8408 -1872 -8327
rect -1940 -9209 -1872 -9128
rect -1947 -10013 -1865 -9931
rect 143 -6880 215 -6824
rect -1623 -7293 -1555 -7212
rect -1460 -7297 -1392 -7216
rect -169 -7129 -113 -7047
rect -170 -7314 -114 -7232
rect 312 -7287 368 -7215
rect -1621 -8096 -1553 -8015
rect -1458 -8096 -1390 -8015
rect -169 -8367 -113 -8295
rect -1622 -8897 -1554 -8816
rect -1460 -8896 -1392 -8815
rect 309 -7682 375 -7677
rect 309 -7740 313 -7682
rect 313 -7740 371 -7682
rect 371 -7740 375 -7682
rect 309 -7743 375 -7740
rect 153 -7985 209 -7913
rect 309 -8059 373 -7995
rect 309 -8175 373 -8111
rect 148 -8577 204 -8505
rect 474 -8576 530 -8504
rect -9 -8733 47 -8661
rect 304 -9031 376 -8975
rect 304 -9154 376 -9098
rect 2127 -6774 2187 -6768
rect 2127 -6828 2174 -6774
rect 2174 -6828 2187 -6774
rect 2241 -6775 2301 -6768
rect 2241 -6828 2259 -6775
rect 2259 -6828 2301 -6775
rect 2882 -6772 2942 -6749
rect 2882 -6809 2931 -6772
rect 2931 -6809 2942 -6772
rect 2996 -6773 3056 -6749
rect 2996 -6809 3010 -6773
rect 3010 -6809 3056 -6773
rect 3039 -7488 3099 -7428
rect 3153 -7488 3213 -7428
rect 3516 -7074 3580 -7010
rect 3516 -7190 3580 -7126
rect 793 -8229 849 -8157
rect 793 -8372 849 -8300
rect 634 -8733 690 -8661
rect 471 -9300 527 -9228
rect -1620 -9700 -1552 -9619
rect -1463 -9698 -1395 -9617
rect 300 -9511 366 -9506
rect 300 -9569 304 -9511
rect 304 -9569 362 -9511
rect 362 -9569 366 -9511
rect 300 -9572 366 -9569
rect 904 -8593 970 -8588
rect 904 -8651 908 -8593
rect 908 -8651 966 -8593
rect 966 -8651 970 -8593
rect 904 -8654 970 -8651
rect 4986 -7296 5050 -7232
rect 4986 -7412 5050 -7348
rect 4986 -7883 5050 -7819
rect 4986 -7999 5050 -7935
rect 4986 -8402 5050 -8338
rect 4986 -8518 5050 -8454
rect 5592 -7297 5656 -7233
rect 5592 -7413 5656 -7349
rect 5592 -7884 5656 -7820
rect 5592 -8000 5656 -7936
rect 5592 -8403 5656 -8339
rect 5592 -8519 5656 -8455
rect 6201 -7295 6265 -7231
rect 6201 -7411 6265 -7347
rect 6201 -7882 6265 -7818
rect 6201 -7998 6265 -7934
rect 6201 -8401 6265 -8337
rect 6201 -8517 6265 -8453
rect 6810 -7298 6874 -7234
rect 6810 -7414 6874 -7350
rect 6810 -7885 6874 -7821
rect 6810 -8001 6874 -7937
rect 6810 -8404 6874 -8340
rect 6810 -8520 6874 -8456
rect 7413 -7306 7477 -7242
rect 7413 -7422 7477 -7358
rect 7413 -7893 7477 -7829
rect 7413 -8009 7477 -7945
rect 7413 -8412 7477 -8348
rect 7413 -8528 7477 -8464
rect 9259 -4971 9324 -4967
rect 9259 -5030 9262 -4971
rect 9262 -5030 9321 -4971
rect 9321 -5030 9324 -4971
rect 9259 -5034 9324 -5030
rect 9262 -5397 9326 -5333
rect 9262 -5513 9326 -5449
rect 9264 -6123 9328 -6059
rect 9264 -6239 9328 -6175
rect 9262 -6854 9326 -6790
rect 9262 -6970 9326 -6906
rect 9258 -7262 9323 -7258
rect 9258 -7321 9261 -7262
rect 9261 -7321 9320 -7262
rect 9320 -7321 9323 -7262
rect 9258 -7325 9323 -7321
rect 9573 -4970 9638 -4966
rect 9573 -5029 9576 -4970
rect 9576 -5029 9635 -4970
rect 9635 -5029 9638 -4970
rect 9573 -5033 9638 -5029
rect 9582 -5397 9646 -5333
rect 9582 -5513 9646 -5449
rect 9584 -6125 9648 -6061
rect 9584 -6241 9648 -6177
rect 9584 -6854 9648 -6790
rect 9584 -6970 9648 -6906
rect 9586 -7259 9651 -7255
rect 9586 -7318 9589 -7259
rect 9589 -7318 9648 -7259
rect 9648 -7318 9651 -7259
rect 9586 -7322 9651 -7318
rect 9890 -4967 9955 -4963
rect 9890 -5026 9893 -4967
rect 9893 -5026 9952 -4967
rect 9952 -5026 9955 -4967
rect 9890 -5030 9955 -5026
rect 9903 -5397 9967 -5333
rect 9903 -5513 9967 -5449
rect 9904 -6127 9968 -6063
rect 9904 -6243 9968 -6179
rect 9903 -6854 9967 -6790
rect 9903 -6970 9967 -6906
rect 9896 -7260 9961 -7256
rect 9896 -7319 9899 -7260
rect 9899 -7319 9958 -7260
rect 9958 -7319 9961 -7260
rect 9896 -7323 9961 -7319
rect 10221 -4966 10286 -4962
rect 10221 -5025 10224 -4966
rect 10224 -5025 10283 -4966
rect 10283 -5025 10286 -4966
rect 10221 -5029 10286 -5025
rect 10223 -5400 10287 -5336
rect 10223 -5516 10287 -5452
rect 10224 -6127 10288 -6063
rect 10224 -6243 10288 -6179
rect 10223 -6856 10287 -6792
rect 10223 -6972 10287 -6908
rect 10222 -7260 10287 -7256
rect 10222 -7319 10225 -7260
rect 10225 -7319 10284 -7260
rect 10284 -7319 10287 -7260
rect 10222 -7323 10287 -7319
rect 10540 -4967 10605 -4963
rect 10540 -5026 10543 -4967
rect 10543 -5026 10602 -4967
rect 10602 -5026 10605 -4967
rect 10540 -5030 10605 -5026
rect 10543 -5398 10607 -5334
rect 10543 -5514 10607 -5450
rect 10541 -6127 10605 -6063
rect 10541 -6243 10605 -6179
rect 10543 -6856 10607 -6792
rect 10543 -6972 10607 -6908
rect 10537 -7256 10602 -7252
rect 10537 -7315 10540 -7256
rect 10540 -7315 10599 -7256
rect 10599 -7315 10602 -7256
rect 10537 -7319 10602 -7315
rect 1928 -9203 1957 -9177
rect 1957 -9203 1992 -9177
rect 1928 -9241 1992 -9203
rect 2073 -9243 2137 -9179
rect 2207 -9204 2223 -9179
rect 2223 -9204 2271 -9179
rect 2207 -9243 2271 -9204
rect 1921 -9501 1985 -9463
rect 1921 -9527 1950 -9501
rect 1950 -9527 1985 -9501
rect 2066 -9525 2130 -9461
rect 2200 -9500 2264 -9461
rect 2200 -9525 2216 -9500
rect 2216 -9525 2264 -9500
rect 313 -9907 369 -9835
rect -169 -10054 -113 -9998
rect 313 -10042 369 -9970
rect -169 -10168 -113 -10112
rect 460 -10420 532 -10364
rect 9259 -7971 9324 -7967
rect 9259 -8030 9262 -7971
rect 9262 -8030 9321 -7971
rect 9321 -8030 9324 -7971
rect 9259 -8034 9324 -8030
rect 9262 -8397 9326 -8333
rect 9262 -8513 9326 -8449
rect 9264 -9123 9328 -9059
rect 9264 -9239 9328 -9175
rect 9262 -9854 9326 -9790
rect 9262 -9970 9326 -9906
rect 9258 -10262 9323 -10258
rect 9258 -10321 9261 -10262
rect 9261 -10321 9320 -10262
rect 9320 -10321 9323 -10262
rect 9258 -10325 9323 -10321
rect 9573 -7970 9638 -7966
rect 9573 -8029 9576 -7970
rect 9576 -8029 9635 -7970
rect 9635 -8029 9638 -7970
rect 9573 -8033 9638 -8029
rect 9582 -8397 9646 -8333
rect 9582 -8513 9646 -8449
rect 9584 -9125 9648 -9061
rect 9584 -9241 9648 -9177
rect 9584 -9854 9648 -9790
rect 9584 -9970 9648 -9906
rect 9586 -10259 9651 -10255
rect 9586 -10318 9589 -10259
rect 9589 -10318 9648 -10259
rect 9648 -10318 9651 -10259
rect 9586 -10322 9651 -10318
rect 9890 -7967 9955 -7963
rect 9890 -8026 9893 -7967
rect 9893 -8026 9952 -7967
rect 9952 -8026 9955 -7967
rect 9890 -8030 9955 -8026
rect 9903 -8397 9967 -8333
rect 9903 -8513 9967 -8449
rect 9904 -9127 9968 -9063
rect 9904 -9243 9968 -9179
rect 9903 -9854 9967 -9790
rect 9903 -9970 9967 -9906
rect 9896 -10260 9961 -10256
rect 9896 -10319 9899 -10260
rect 9899 -10319 9958 -10260
rect 9958 -10319 9961 -10260
rect 9896 -10323 9961 -10319
rect 10221 -7966 10286 -7962
rect 10221 -8025 10224 -7966
rect 10224 -8025 10283 -7966
rect 10283 -8025 10286 -7966
rect 10221 -8029 10286 -8025
rect 10223 -8400 10287 -8336
rect 10223 -8516 10287 -8452
rect 10224 -9127 10288 -9063
rect 10224 -9243 10288 -9179
rect 10223 -9856 10287 -9792
rect 10223 -9972 10287 -9908
rect 10222 -10260 10287 -10256
rect 10222 -10319 10225 -10260
rect 10225 -10319 10284 -10260
rect 10284 -10319 10287 -10260
rect 10222 -10323 10287 -10319
rect 10540 -7967 10605 -7963
rect 10540 -8026 10543 -7967
rect 10543 -8026 10602 -7967
rect 10602 -8026 10605 -7967
rect 10540 -8030 10605 -8026
rect 10543 -8398 10607 -8334
rect 10543 -8514 10607 -8450
rect 10541 -9127 10605 -9063
rect 10541 -9243 10605 -9179
rect 10543 -9856 10607 -9792
rect 10543 -9972 10607 -9908
rect 10537 -10256 10602 -10252
rect 10537 -10315 10540 -10256
rect 10540 -10315 10599 -10256
rect 10599 -10315 10602 -10256
rect 10537 -10319 10602 -10315
<< metal2 >>
rect -2441 1297 -522 1496
rect -2441 1266 -2242 1297
rect -2441 1213 -2416 1266
rect -2364 1213 -2304 1266
rect -2252 1213 -2242 1266
rect -2441 1180 -2242 1213
rect -2791 -1762 -2675 -1744
rect -2791 -1845 -2775 -1762
rect -2691 -1845 -2675 -1762
rect -2791 -1861 -2675 -1845
rect -2359 -1760 -2243 -1742
rect -2359 -1843 -2343 -1760
rect -2259 -1843 -2243 -1760
rect -2359 -1859 -2243 -1843
rect -1926 -1760 -1810 -1742
rect -1926 -1843 -1910 -1760
rect -1826 -1843 -1810 -1760
rect -1926 -1859 -1810 -1843
rect -3492 -2170 -3232 -2168
rect -2774 -2170 -2691 -1861
rect -2342 -2170 -2259 -1859
rect -1911 -2170 -1828 -1859
rect -721 -2121 -522 1297
rect 2806 643 2940 712
rect 2806 579 2843 643
rect 2907 579 2940 643
rect 169 535 1681 553
rect 169 457 191 535
rect 271 457 1681 535
rect 169 439 1681 457
rect -259 333 -146 337
rect -259 323 1474 333
rect -259 233 -244 323
rect -162 311 1474 323
rect -162 237 625 311
rect 700 237 1474 311
rect -162 233 1474 237
rect -259 222 1474 233
rect -259 219 -147 222
rect -260 -66 -144 -44
rect -260 -145 -242 -66
rect -160 -145 -144 -66
rect -260 -160 -144 -145
rect 605 -71 721 -51
rect 605 -150 621 -71
rect 703 -150 721 -71
rect -236 -437 -164 -160
rect 605 -167 721 -150
rect -257 -456 -146 -437
rect 628 -441 699 -167
rect -257 -535 -242 -456
rect -160 -535 -146 -456
rect -257 -550 -146 -535
rect 609 -455 718 -441
rect 609 -534 623 -455
rect 705 -534 718 -455
rect 609 -549 718 -534
rect 243 -1109 366 -1088
rect 243 -1188 270 -1109
rect 353 -1188 366 -1109
rect 243 -1204 366 -1188
rect 1363 -1108 1474 222
rect 1363 -1186 1377 -1108
rect 1461 -1186 1474 -1108
rect -721 -2154 1135 -2121
rect -3492 -2373 -1760 -2170
rect -721 -2235 185 -2154
rect 266 -2235 1135 -2154
rect -721 -2320 1135 -2235
rect -3492 -2420 -3232 -2373
rect -4059 -2471 -3700 -2447
rect -4059 -2591 -4042 -2471
rect -3919 -2591 -3842 -2471
rect -3719 -2591 -3700 -2471
rect -4059 -2608 -3700 -2591
rect -4063 -2723 -3687 -2693
rect -4063 -2843 -4039 -2723
rect -3916 -2843 -3839 -2723
rect -3716 -2843 -3687 -2723
rect -4063 -2868 -3687 -2843
rect -3472 -3116 -3269 -2420
rect -1750 -2730 -1634 -2712
rect -1750 -2810 -1734 -2730
rect -1654 -2810 -1634 -2730
rect -1750 -2825 -1634 -2810
rect -2614 -2953 -2517 -2940
rect -1978 -2952 -1881 -2942
rect -2614 -3034 -2599 -2953
rect -2531 -2965 -2517 -2953
rect -2156 -2955 -1881 -2952
rect -2156 -2965 -1963 -2955
rect -2531 -3021 -2142 -2965
rect -2086 -3021 -2032 -2965
rect -1976 -3021 -1963 -2965
rect -2531 -3025 -1963 -3021
rect -2531 -3034 -2517 -3025
rect -2614 -3047 -2517 -3034
rect -2156 -3036 -1963 -3025
rect -1895 -3036 -1881 -2955
rect -1978 -3049 -1881 -3036
rect -2774 -3109 -2677 -3096
rect -2774 -3116 -2759 -3109
rect -3472 -3177 -2759 -3116
rect -3472 -3973 -3269 -3177
rect -2774 -3190 -2759 -3177
rect -2691 -3116 -2677 -3109
rect -2454 -3101 -2357 -3088
rect -2454 -3116 -2439 -3101
rect -2691 -3177 -2439 -3116
rect -2691 -3190 -2677 -3177
rect -2774 -3203 -2677 -3190
rect -2454 -3182 -2439 -3177
rect -2371 -3116 -2357 -3101
rect -2133 -3109 -2036 -3096
rect -2133 -3116 -2118 -3109
rect -2371 -3177 -2118 -3116
rect -2371 -3182 -2357 -3177
rect -2454 -3195 -2357 -3182
rect -2133 -3190 -2118 -3177
rect -2050 -3116 -2036 -3109
rect -1818 -3105 -1721 -3092
rect -1818 -3116 -1803 -3105
rect -2050 -3177 -1803 -3116
rect -2050 -3190 -2036 -3177
rect -2133 -3203 -2036 -3190
rect -1818 -3186 -1803 -3177
rect -1735 -3186 -1721 -3105
rect -1818 -3199 -1721 -3186
rect -264 -3117 -144 -3092
rect -264 -3197 -243 -3117
rect -163 -3197 -144 -3117
rect -264 -3216 -144 -3197
rect 174 -3117 285 -3100
rect 174 -3200 189 -3117
rect 271 -3200 285 -3117
rect 174 -3214 285 -3200
rect 607 -3110 718 -3096
rect 607 -3196 620 -3110
rect 704 -3196 718 -3110
rect 607 -3210 718 -3196
rect -3094 -3260 -2997 -3247
rect -3094 -3341 -3079 -3260
rect -3011 -3272 -2997 -3260
rect -2937 -3262 -2840 -3249
rect -2937 -3272 -2922 -3262
rect -3011 -3332 -2922 -3272
rect -3011 -3341 -2997 -3332
rect -3094 -3354 -2997 -3341
rect -2937 -3343 -2922 -3332
rect -2854 -3272 -2840 -3262
rect -2547 -3272 -2355 -3260
rect -2294 -3261 -2197 -3248
rect -2294 -3272 -2279 -3261
rect -2854 -3273 -2279 -3272
rect -2854 -3329 -2533 -3273
rect -2477 -3329 -2423 -3273
rect -2367 -3329 -2279 -3273
rect -2854 -3332 -2279 -3329
rect -2854 -3343 -2840 -3332
rect -2937 -3356 -2840 -3343
rect -2547 -3344 -2355 -3332
rect -2294 -3342 -2279 -3332
rect -2211 -3272 -2197 -3261
rect -1658 -3264 -1561 -3251
rect -1658 -3272 -1643 -3264
rect -2211 -3332 -1643 -3272
rect -2211 -3342 -2197 -3332
rect -2294 -3355 -2197 -3342
rect -1658 -3345 -1643 -3332
rect -1575 -3272 -1561 -3264
rect -1492 -3260 -1395 -3247
rect -1492 -3272 -1477 -3260
rect -1575 -3332 -1477 -3272
rect -1575 -3345 -1561 -3332
rect -1658 -3358 -1561 -3345
rect -1492 -3341 -1477 -3332
rect -1409 -3341 -1395 -3260
rect -1492 -3354 -1395 -3341
rect -2854 -3549 -2750 -3538
rect -238 -3544 -168 -3216
rect -2854 -3629 -2844 -3549
rect -2762 -3629 -2750 -3549
rect -2854 -3639 -2750 -3629
rect -265 -3563 -143 -3544
rect -265 -3649 -245 -3563
rect -161 -3649 -143 -3563
rect -265 -3662 -143 -3649
rect 194 -3730 264 -3214
rect 634 -3513 693 -3210
rect 633 -3546 694 -3513
rect 465 -3565 723 -3546
rect 465 -3651 477 -3565
rect 561 -3651 621 -3565
rect 705 -3651 723 -3565
rect 465 -3667 723 -3651
rect 8 -3761 316 -3730
rect -2615 -3806 -2518 -3798
rect -1972 -3805 -1875 -3792
rect -2615 -3811 -2332 -3806
rect -2615 -3892 -2600 -3811
rect -2532 -3819 -2332 -3811
rect -2532 -3875 -2510 -3819
rect -2454 -3875 -2400 -3819
rect -2344 -3820 -2332 -3819
rect -1972 -3820 -1957 -3805
rect -2344 -3875 -1957 -3820
rect -2532 -3880 -1957 -3875
rect -2532 -3890 -2332 -3880
rect -1972 -3886 -1957 -3880
rect -1889 -3886 -1875 -3805
rect 8 -3847 25 -3761
rect 109 -3762 316 -3761
rect 109 -3847 184 -3762
rect 8 -3848 184 -3847
rect 268 -3848 316 -3762
rect 8 -3860 316 -3848
rect -2532 -3892 -2518 -3890
rect -2615 -3905 -2518 -3892
rect -1972 -3899 -1875 -3886
rect 149 -3863 285 -3860
rect -2772 -3961 -2675 -3948
rect -2772 -3973 -2757 -3961
rect -3472 -4034 -2757 -3973
rect -3472 -4837 -3269 -4034
rect -2772 -4042 -2757 -4034
rect -2689 -3973 -2675 -3961
rect -2455 -3966 -2358 -3953
rect -2455 -3973 -2440 -3966
rect -2689 -4034 -2440 -3973
rect -2689 -4042 -2675 -4034
rect -2772 -4055 -2675 -4042
rect -2455 -4047 -2440 -4034
rect -2372 -3973 -2358 -3966
rect -2135 -3961 -2038 -3948
rect -2135 -3973 -2120 -3961
rect -2372 -4034 -2120 -3973
rect -2372 -4047 -2358 -4034
rect -2455 -4060 -2358 -4047
rect -2135 -4042 -2120 -4034
rect -2052 -3973 -2038 -3961
rect -1815 -3959 -1718 -3946
rect -1815 -3973 -1800 -3959
rect -2052 -4034 -1800 -3973
rect -2052 -4042 -2038 -4034
rect -2135 -4055 -2038 -4042
rect -1815 -4040 -1800 -4034
rect -1732 -4040 -1718 -3959
rect -1815 -4053 -1718 -4040
rect -3095 -4119 -2998 -4106
rect -3095 -4200 -3080 -4119
rect -3012 -4132 -2998 -4119
rect -2938 -4122 -2841 -4109
rect -2938 -4132 -2923 -4122
rect -3012 -4192 -2923 -4132
rect -3012 -4200 -2998 -4192
rect -3095 -4213 -2998 -4200
rect -2938 -4203 -2923 -4192
rect -2855 -4132 -2841 -4122
rect -2295 -4123 -2198 -4110
rect -2295 -4132 -2280 -4123
rect -2855 -4192 -2280 -4132
rect -2855 -4203 -2841 -4192
rect -2938 -4216 -2841 -4203
rect -2295 -4204 -2280 -4192
rect -2212 -4132 -2198 -4123
rect -2121 -4131 -1929 -4118
rect -2121 -4132 -2107 -4131
rect -2212 -4187 -2107 -4132
rect -2051 -4187 -1997 -4131
rect -1941 -4132 -1929 -4131
rect -1658 -4120 -1561 -4107
rect -1658 -4132 -1643 -4120
rect -1941 -4187 -1643 -4132
rect -2212 -4192 -1643 -4187
rect -2212 -4204 -2198 -4192
rect -2121 -4202 -1929 -4192
rect -1658 -4201 -1643 -4192
rect -1575 -4132 -1561 -4120
rect -1493 -4118 -1396 -4105
rect -1493 -4132 -1478 -4118
rect -1575 -4192 -1478 -4132
rect -1575 -4201 -1561 -4192
rect -2295 -4217 -2198 -4204
rect -1658 -4214 -1561 -4201
rect -1493 -4199 -1478 -4192
rect -1410 -4199 -1396 -4118
rect -1493 -4212 -1396 -4199
rect 149 -4220 283 -3863
rect -281 -4245 -53 -4221
rect -281 -4309 -261 -4245
rect -197 -4309 -145 -4245
rect -81 -4309 -53 -4245
rect 149 -4292 189 -4220
rect 266 -4292 283 -4220
rect 149 -4309 283 -4292
rect -281 -4327 -53 -4309
rect 584 -4318 705 -3667
rect 936 -4062 1135 -2320
rect 1363 -3542 1474 -1186
rect 1567 -71 1681 439
rect 1567 -149 1583 -71
rect 1666 -149 1681 -71
rect 1352 -3557 1486 -3542
rect 1352 -3661 1364 -3557
rect 1473 -3661 1486 -3557
rect 1352 -3676 1486 -3661
rect 1567 -3739 1681 -149
rect 2806 527 2940 579
rect 2806 463 2843 527
rect 2907 463 2940 527
rect 2806 -97 2940 463
rect 2806 -161 2843 -97
rect 2907 -161 2940 -97
rect 2806 -213 2940 -161
rect 2806 -277 2843 -213
rect 2907 -277 2940 -213
rect 2806 -860 2940 -277
rect 2806 -924 2843 -860
rect 2907 -924 2940 -860
rect 2806 -976 2940 -924
rect 2806 -1040 2843 -976
rect 2907 -1040 2940 -976
rect 2806 -1589 2940 -1040
rect 2806 -1653 2843 -1589
rect 2907 -1653 2940 -1589
rect 2806 -1705 2940 -1653
rect 2806 -1769 2843 -1705
rect 2907 -1769 2940 -1705
rect 2806 -2307 2940 -1769
rect 2806 -2371 2843 -2307
rect 2907 -2371 2940 -2307
rect 2806 -2423 2940 -2371
rect 2806 -2487 2843 -2423
rect 2907 -2487 2940 -2423
rect 2806 -3446 2940 -2487
rect 3127 641 3261 707
rect 3127 577 3163 641
rect 3227 577 3261 641
rect 3127 525 3261 577
rect 3127 461 3163 525
rect 3227 461 3261 525
rect 3127 -99 3261 461
rect 3127 -163 3163 -99
rect 3227 -163 3261 -99
rect 3127 -215 3261 -163
rect 3127 -279 3163 -215
rect 3227 -279 3261 -215
rect 3127 -828 3261 -279
rect 3127 -892 3163 -828
rect 3227 -892 3261 -828
rect 3127 -944 3261 -892
rect 3127 -1008 3163 -944
rect 3227 -1008 3261 -944
rect 3127 -1568 3261 -1008
rect 3127 -1632 3163 -1568
rect 3227 -1632 3261 -1568
rect 3127 -1684 3261 -1632
rect 3127 -1748 3163 -1684
rect 3227 -1748 3261 -1684
rect 3127 -2308 3261 -1748
rect 3127 -2372 3163 -2308
rect 3227 -2372 3261 -2308
rect 3127 -2424 3261 -2372
rect 3127 -2488 3163 -2424
rect 3227 -2488 3261 -2424
rect 3127 -3446 3261 -2488
rect 3444 671 3578 704
rect 3444 607 3483 671
rect 3547 607 3578 671
rect 3444 555 3578 607
rect 3444 491 3483 555
rect 3547 491 3578 555
rect 3444 -80 3578 491
rect 3444 -144 3483 -80
rect 3547 -144 3578 -80
rect 3444 -196 3578 -144
rect 3444 -260 3483 -196
rect 3547 -260 3578 -196
rect 3444 -812 3578 -260
rect 3444 -876 3483 -812
rect 3547 -876 3578 -812
rect 3444 -928 3578 -876
rect 3444 -992 3483 -928
rect 3547 -992 3578 -928
rect 3444 -1554 3578 -992
rect 3444 -1618 3483 -1554
rect 3547 -1618 3578 -1554
rect 3444 -1670 3578 -1618
rect 3444 -1734 3483 -1670
rect 3547 -1734 3578 -1670
rect 3444 -2314 3578 -1734
rect 3444 -2378 3483 -2314
rect 3547 -2378 3578 -2314
rect 3444 -2430 3578 -2378
rect 3444 -2494 3483 -2430
rect 3547 -2494 3578 -2430
rect 3444 -3105 3578 -2494
rect 3765 658 3899 709
rect 3765 594 3803 658
rect 3867 594 3899 658
rect 3765 542 3899 594
rect 3765 478 3803 542
rect 3867 478 3899 542
rect 3765 -101 3899 478
rect 3765 -165 3803 -101
rect 3867 -165 3899 -101
rect 3765 -217 3899 -165
rect 3765 -281 3803 -217
rect 3867 -281 3899 -217
rect 3765 -837 3899 -281
rect 3765 -901 3803 -837
rect 3867 -901 3899 -837
rect 3765 -953 3899 -901
rect 3765 -1017 3803 -953
rect 3867 -1017 3899 -953
rect 3765 -1562 3899 -1017
rect 3765 -1626 3803 -1562
rect 3867 -1626 3899 -1562
rect 3765 -1678 3899 -1626
rect 3765 -1742 3803 -1678
rect 3867 -1742 3899 -1678
rect 3765 -2310 3899 -1742
rect 3765 -2374 3803 -2310
rect 3867 -2374 3899 -2310
rect 3765 -2426 3899 -2374
rect 3765 -2490 3803 -2426
rect 3867 -2490 3899 -2426
rect 3400 -3119 3615 -3105
rect 3400 -3183 3417 -3119
rect 3481 -3183 3537 -3119
rect 3601 -3183 3615 -3119
rect 3400 -3239 3615 -3183
rect 3400 -3303 3417 -3239
rect 3481 -3303 3537 -3239
rect 3601 -3303 3615 -3239
rect 3400 -3317 3615 -3303
rect 2761 -3460 2976 -3446
rect 2761 -3524 2778 -3460
rect 2842 -3524 2898 -3460
rect 2962 -3524 2976 -3460
rect 2761 -3580 2976 -3524
rect 2761 -3644 2778 -3580
rect 2842 -3644 2898 -3580
rect 2962 -3644 2976 -3580
rect 2761 -3658 2976 -3644
rect 3089 -3460 3304 -3446
rect 3765 -3447 3899 -2490
rect 4086 655 4220 712
rect 4086 591 4123 655
rect 4187 591 4220 655
rect 4086 539 4220 591
rect 4086 475 4123 539
rect 4187 475 4220 539
rect 4086 -116 4220 475
rect 4086 -180 4123 -116
rect 4187 -180 4220 -116
rect 4086 -232 4220 -180
rect 4086 -296 4123 -232
rect 4187 -296 4220 -232
rect 4086 -841 4220 -296
rect 4086 -905 4123 -841
rect 4187 -905 4220 -841
rect 4086 -957 4220 -905
rect 4086 -1021 4123 -957
rect 4187 -1021 4220 -957
rect 4086 -1565 4220 -1021
rect 4086 -1629 4123 -1565
rect 4187 -1629 4220 -1565
rect 4086 -1681 4220 -1629
rect 4086 -1745 4123 -1681
rect 4187 -1745 4220 -1681
rect 4086 -2313 4220 -1745
rect 4086 -2377 4123 -2313
rect 4187 -2377 4220 -2313
rect 4086 -2429 4220 -2377
rect 4086 -2493 4123 -2429
rect 4187 -2493 4220 -2429
rect 4086 -3446 4220 -2493
rect 5606 643 5740 712
rect 5606 579 5643 643
rect 5707 579 5740 643
rect 5606 527 5740 579
rect 5606 463 5643 527
rect 5707 463 5740 527
rect 5606 -97 5740 463
rect 5606 -161 5643 -97
rect 5707 -161 5740 -97
rect 5606 -213 5740 -161
rect 5606 -277 5643 -213
rect 5707 -277 5740 -213
rect 5606 -860 5740 -277
rect 5606 -924 5643 -860
rect 5707 -924 5740 -860
rect 5606 -976 5740 -924
rect 5606 -1040 5643 -976
rect 5707 -1040 5740 -976
rect 5606 -1589 5740 -1040
rect 5606 -1653 5643 -1589
rect 5707 -1653 5740 -1589
rect 5606 -1705 5740 -1653
rect 5606 -1769 5643 -1705
rect 5707 -1769 5740 -1705
rect 5606 -2307 5740 -1769
rect 5606 -2371 5643 -2307
rect 5707 -2371 5740 -2307
rect 5606 -2423 5740 -2371
rect 5606 -2487 5643 -2423
rect 5707 -2487 5740 -2423
rect 5606 -3446 5740 -2487
rect 5927 641 6061 707
rect 5927 577 5963 641
rect 6027 577 6061 641
rect 5927 525 6061 577
rect 5927 461 5963 525
rect 6027 461 6061 525
rect 5927 -99 6061 461
rect 5927 -163 5963 -99
rect 6027 -163 6061 -99
rect 5927 -215 6061 -163
rect 5927 -279 5963 -215
rect 6027 -279 6061 -215
rect 5927 -828 6061 -279
rect 5927 -892 5963 -828
rect 6027 -892 6061 -828
rect 5927 -944 6061 -892
rect 5927 -1008 5963 -944
rect 6027 -1008 6061 -944
rect 5927 -1568 6061 -1008
rect 5927 -1632 5963 -1568
rect 6027 -1632 6061 -1568
rect 5927 -1684 6061 -1632
rect 5927 -1748 5963 -1684
rect 6027 -1748 6061 -1684
rect 5927 -2308 6061 -1748
rect 5927 -2372 5963 -2308
rect 6027 -2372 6061 -2308
rect 5927 -2424 6061 -2372
rect 5927 -2488 5963 -2424
rect 6027 -2488 6061 -2424
rect 5927 -3446 6061 -2488
rect 6244 671 6378 704
rect 6244 607 6283 671
rect 6347 607 6378 671
rect 6244 555 6378 607
rect 6244 491 6283 555
rect 6347 491 6378 555
rect 6244 -80 6378 491
rect 6244 -144 6283 -80
rect 6347 -144 6378 -80
rect 6244 -196 6378 -144
rect 6244 -260 6283 -196
rect 6347 -260 6378 -196
rect 6244 -812 6378 -260
rect 6244 -876 6283 -812
rect 6347 -876 6378 -812
rect 6244 -928 6378 -876
rect 6244 -992 6283 -928
rect 6347 -992 6378 -928
rect 6244 -1554 6378 -992
rect 6244 -1618 6283 -1554
rect 6347 -1618 6378 -1554
rect 6244 -1670 6378 -1618
rect 6244 -1734 6283 -1670
rect 6347 -1734 6378 -1670
rect 6244 -2314 6378 -1734
rect 6244 -2378 6283 -2314
rect 6347 -2378 6378 -2314
rect 6244 -2430 6378 -2378
rect 6244 -2494 6283 -2430
rect 6347 -2494 6378 -2430
rect 6244 -3105 6378 -2494
rect 6565 658 6699 709
rect 6565 594 6603 658
rect 6667 594 6699 658
rect 6565 542 6699 594
rect 6565 478 6603 542
rect 6667 478 6699 542
rect 6565 -101 6699 478
rect 6565 -165 6603 -101
rect 6667 -165 6699 -101
rect 6565 -217 6699 -165
rect 6565 -281 6603 -217
rect 6667 -281 6699 -217
rect 6565 -837 6699 -281
rect 6565 -901 6603 -837
rect 6667 -901 6699 -837
rect 6565 -953 6699 -901
rect 6565 -1017 6603 -953
rect 6667 -1017 6699 -953
rect 6565 -1562 6699 -1017
rect 6565 -1626 6603 -1562
rect 6667 -1626 6699 -1562
rect 6565 -1678 6699 -1626
rect 6565 -1742 6603 -1678
rect 6667 -1742 6699 -1678
rect 6565 -2310 6699 -1742
rect 6565 -2374 6603 -2310
rect 6667 -2374 6699 -2310
rect 6565 -2426 6699 -2374
rect 6565 -2490 6603 -2426
rect 6667 -2490 6699 -2426
rect 6200 -3119 6415 -3105
rect 6200 -3183 6217 -3119
rect 6281 -3183 6337 -3119
rect 6401 -3183 6415 -3119
rect 6200 -3239 6415 -3183
rect 6200 -3303 6217 -3239
rect 6281 -3303 6337 -3239
rect 6401 -3303 6415 -3239
rect 6200 -3317 6415 -3303
rect 3089 -3524 3106 -3460
rect 3170 -3524 3226 -3460
rect 3290 -3524 3304 -3460
rect 3089 -3580 3304 -3524
rect 3089 -3644 3106 -3580
rect 3170 -3644 3226 -3580
rect 3290 -3644 3304 -3580
rect 3089 -3658 3304 -3644
rect 3717 -3461 3932 -3447
rect 3717 -3525 3734 -3461
rect 3798 -3525 3854 -3461
rect 3918 -3525 3932 -3461
rect 3717 -3581 3932 -3525
rect 3717 -3645 3734 -3581
rect 3798 -3645 3854 -3581
rect 3918 -3645 3932 -3581
rect 3717 -3659 3932 -3645
rect 4043 -3460 4258 -3446
rect 4043 -3524 4060 -3460
rect 4124 -3524 4180 -3460
rect 4244 -3524 4258 -3460
rect 4043 -3580 4258 -3524
rect 4043 -3644 4060 -3580
rect 4124 -3644 4180 -3580
rect 4244 -3644 4258 -3580
rect 4043 -3658 4258 -3644
rect 5561 -3460 5776 -3446
rect 5561 -3524 5578 -3460
rect 5642 -3524 5698 -3460
rect 5762 -3524 5776 -3460
rect 5561 -3580 5776 -3524
rect 5561 -3644 5578 -3580
rect 5642 -3644 5698 -3580
rect 5762 -3644 5776 -3580
rect 5561 -3658 5776 -3644
rect 5889 -3460 6104 -3446
rect 6565 -3447 6699 -2490
rect 6886 655 7020 712
rect 6886 591 6923 655
rect 6987 591 7020 655
rect 6886 539 7020 591
rect 6886 475 6923 539
rect 6987 475 7020 539
rect 6886 -116 7020 475
rect 6886 -180 6923 -116
rect 6987 -180 7020 -116
rect 6886 -232 7020 -180
rect 6886 -296 6923 -232
rect 6987 -296 7020 -232
rect 6886 -841 7020 -296
rect 6886 -905 6923 -841
rect 6987 -905 7020 -841
rect 6886 -957 7020 -905
rect 6886 -1021 6923 -957
rect 6987 -1021 7020 -957
rect 6886 -1565 7020 -1021
rect 6886 -1629 6923 -1565
rect 6987 -1629 7020 -1565
rect 6886 -1681 7020 -1629
rect 6886 -1745 6923 -1681
rect 6987 -1745 7020 -1681
rect 6886 -2313 7020 -1745
rect 6886 -2377 6923 -2313
rect 6987 -2377 7020 -2313
rect 6886 -2429 7020 -2377
rect 6886 -2493 6923 -2429
rect 6987 -2493 7020 -2429
rect 6886 -3446 7020 -2493
rect 8406 643 8540 712
rect 8406 579 8443 643
rect 8507 579 8540 643
rect 8406 527 8540 579
rect 8406 463 8443 527
rect 8507 463 8540 527
rect 8406 -97 8540 463
rect 8406 -161 8443 -97
rect 8507 -161 8540 -97
rect 8406 -213 8540 -161
rect 8406 -277 8443 -213
rect 8507 -277 8540 -213
rect 8406 -860 8540 -277
rect 8406 -924 8443 -860
rect 8507 -924 8540 -860
rect 8406 -976 8540 -924
rect 8406 -1040 8443 -976
rect 8507 -1040 8540 -976
rect 8406 -1589 8540 -1040
rect 8406 -1653 8443 -1589
rect 8507 -1653 8540 -1589
rect 8406 -1705 8540 -1653
rect 8406 -1769 8443 -1705
rect 8507 -1769 8540 -1705
rect 8406 -2307 8540 -1769
rect 8406 -2371 8443 -2307
rect 8507 -2371 8540 -2307
rect 8406 -2423 8540 -2371
rect 8406 -2487 8443 -2423
rect 8507 -2487 8540 -2423
rect 7330 -3098 7784 -3082
rect 7330 -3162 7347 -3098
rect 7411 -3162 7467 -3098
rect 7531 -3162 7587 -3098
rect 7651 -3162 7707 -3098
rect 7771 -3162 7784 -3098
rect 7330 -3218 7784 -3162
rect 7330 -3282 7347 -3218
rect 7411 -3282 7467 -3218
rect 7531 -3282 7587 -3218
rect 7651 -3282 7707 -3218
rect 7771 -3282 7784 -3218
rect 7330 -3296 7784 -3282
rect 5889 -3524 5906 -3460
rect 5970 -3524 6026 -3460
rect 6090 -3524 6104 -3460
rect 5889 -3580 6104 -3524
rect 5889 -3644 5906 -3580
rect 5970 -3644 6026 -3580
rect 6090 -3644 6104 -3580
rect 5889 -3658 6104 -3644
rect 6517 -3461 6732 -3447
rect 6517 -3525 6534 -3461
rect 6598 -3525 6654 -3461
rect 6718 -3525 6732 -3461
rect 6517 -3581 6732 -3525
rect 6517 -3645 6534 -3581
rect 6598 -3645 6654 -3581
rect 6718 -3645 6732 -3581
rect 6517 -3659 6732 -3645
rect 6843 -3460 7058 -3446
rect 6843 -3524 6860 -3460
rect 6924 -3524 6980 -3460
rect 7044 -3524 7058 -3460
rect 6843 -3580 7058 -3524
rect 6843 -3644 6860 -3580
rect 6924 -3644 6980 -3580
rect 7044 -3644 7058 -3580
rect 6843 -3658 7058 -3644
rect 1552 -3753 1687 -3739
rect 1552 -3858 1565 -3753
rect 1675 -3858 1687 -3753
rect 1552 -3874 1687 -3858
rect 936 -4261 2779 -4062
rect -1756 -4393 -1633 -4376
rect -1756 -4478 -1737 -4393
rect -1650 -4478 -1633 -4393
rect -1756 -4491 -1633 -4478
rect -247 -4565 -97 -4327
rect 340 -4336 705 -4318
rect 340 -4415 355 -4336
rect 434 -4415 705 -4336
rect 340 -4439 705 -4415
rect 2580 -4461 2779 -4261
rect 2561 -4479 2799 -4461
rect 2561 -4543 2579 -4479
rect 2643 -4543 2719 -4479
rect 2783 -4543 2799 -4479
rect -2615 -4661 -2518 -4648
rect -2615 -4742 -2600 -4661
rect -2532 -4666 -2518 -4661
rect -1976 -4665 -1879 -4652
rect -2532 -4679 -2332 -4666
rect -2532 -4735 -2510 -4679
rect -2454 -4735 -2400 -4679
rect -2344 -4680 -2332 -4679
rect -1976 -4680 -1961 -4665
rect -2344 -4735 -1961 -4680
rect -2532 -4740 -1961 -4735
rect -2532 -4742 -2332 -4740
rect -2615 -4750 -2332 -4742
rect -1976 -4746 -1961 -4740
rect -1893 -4746 -1879 -4665
rect -247 -4715 1509 -4565
rect 2561 -4595 2799 -4543
rect 2561 -4659 2579 -4595
rect 2643 -4659 2719 -4595
rect 2783 -4659 2799 -4595
rect 2561 -4677 2799 -4659
rect -2615 -4755 -2518 -4750
rect -1976 -4759 -1879 -4746
rect -2775 -4819 -2678 -4806
rect -2775 -4837 -2760 -4819
rect -3472 -4898 -2760 -4837
rect -3472 -5691 -3269 -4898
rect -2775 -4900 -2760 -4898
rect -2692 -4837 -2678 -4819
rect -2457 -4823 -2360 -4810
rect -2457 -4837 -2442 -4823
rect -2692 -4898 -2442 -4837
rect -2692 -4900 -2678 -4898
rect -2775 -4913 -2678 -4900
rect -2457 -4904 -2442 -4898
rect -2374 -4837 -2360 -4823
rect -2131 -4817 -2034 -4804
rect -2131 -4837 -2116 -4817
rect -2374 -4898 -2116 -4837
rect -2048 -4837 -2034 -4817
rect -1817 -4828 -1720 -4815
rect -1817 -4837 -1802 -4828
rect -2048 -4898 -1802 -4837
rect -2374 -4904 -2360 -4898
rect -2457 -4917 -2360 -4904
rect -2131 -4911 -2034 -4898
rect -1817 -4909 -1802 -4898
rect -1734 -4909 -1720 -4828
rect -1817 -4922 -1720 -4909
rect 793 -4852 891 -4830
rect 793 -4916 811 -4852
rect 875 -4916 891 -4852
rect -3092 -4969 -2995 -4956
rect -3092 -5050 -3077 -4969
rect -3009 -4987 -2995 -4969
rect -2935 -4972 -2838 -4959
rect -2935 -4987 -2920 -4972
rect -3009 -5047 -2920 -4987
rect -3009 -5050 -2995 -5047
rect -3092 -5063 -2995 -5050
rect -2935 -5053 -2920 -5047
rect -2852 -4987 -2838 -4972
rect -2295 -4974 -2198 -4961
rect -2295 -4987 -2280 -4974
rect -2852 -5047 -2280 -4987
rect -2852 -5053 -2838 -5047
rect -2935 -5066 -2838 -5053
rect -2295 -5055 -2280 -5047
rect -2212 -4987 -2198 -4974
rect -1651 -4975 -1554 -4962
rect -2120 -4987 -1928 -4976
rect -1651 -4987 -1636 -4975
rect -2212 -4989 -1636 -4987
rect -2212 -5045 -2106 -4989
rect -2050 -5045 -1996 -4989
rect -1940 -5045 -1636 -4989
rect -2212 -5047 -1636 -5045
rect -2212 -5055 -2198 -5047
rect -2295 -5068 -2198 -5055
rect -2120 -5060 -1928 -5047
rect -1651 -5056 -1636 -5047
rect -1568 -4987 -1554 -4975
rect -1494 -4971 -1397 -4958
rect -1494 -4987 -1479 -4971
rect -1568 -5047 -1479 -4987
rect -1568 -5056 -1554 -5047
rect -1651 -5069 -1554 -5056
rect -1494 -5052 -1479 -5047
rect -1411 -5052 -1397 -4971
rect -1494 -5065 -1397 -5052
rect 793 -4968 891 -4916
rect 793 -5032 811 -4968
rect 875 -4978 891 -4968
rect 875 -5032 890 -4978
rect -2861 -5252 -2740 -5234
rect -2861 -5337 -2845 -5252
rect -2759 -5337 -2740 -5252
rect -2861 -5352 -2740 -5337
rect -2613 -5528 -2516 -5515
rect -1970 -5527 -1873 -5514
rect -2613 -5609 -2598 -5528
rect -2530 -5540 -2516 -5528
rect -2155 -5540 -1955 -5527
rect -2530 -5596 -2141 -5540
rect -2085 -5596 -2031 -5540
rect -1975 -5596 -1955 -5540
rect -2530 -5600 -1955 -5596
rect -2530 -5609 -2516 -5600
rect -2613 -5622 -2516 -5609
rect -2155 -5608 -1955 -5600
rect -1887 -5608 -1873 -5527
rect -2155 -5611 -1873 -5608
rect -1970 -5621 -1873 -5611
rect 793 -5533 890 -5032
rect 793 -5597 810 -5533
rect 874 -5567 890 -5533
rect 874 -5597 891 -5567
rect 793 -5649 891 -5597
rect -2778 -5679 -2681 -5666
rect -2778 -5691 -2763 -5679
rect -3472 -5752 -2763 -5691
rect -3472 -5826 -3269 -5752
rect -2778 -5760 -2763 -5752
rect -2695 -5691 -2681 -5679
rect -2456 -5678 -2359 -5665
rect -2456 -5691 -2441 -5678
rect -2695 -5752 -2441 -5691
rect -2695 -5760 -2681 -5752
rect -2778 -5773 -2681 -5760
rect -2456 -5759 -2441 -5752
rect -2373 -5691 -2359 -5678
rect -2141 -5686 -2044 -5673
rect -2141 -5691 -2126 -5686
rect -2373 -5752 -2126 -5691
rect -2373 -5759 -2359 -5752
rect -2456 -5772 -2359 -5759
rect -2141 -5767 -2126 -5752
rect -2058 -5691 -2044 -5686
rect -1812 -5684 -1715 -5671
rect -1812 -5691 -1797 -5684
rect -2058 -5752 -1797 -5691
rect -2058 -5767 -2044 -5752
rect -2141 -5780 -2044 -5767
rect -1812 -5765 -1797 -5752
rect -1729 -5765 -1715 -5684
rect -1812 -5778 -1715 -5765
rect 793 -5713 810 -5649
rect 874 -5700 891 -5649
rect 874 -5713 890 -5700
rect -3092 -5844 -2995 -5831
rect -3092 -5925 -3077 -5844
rect -3009 -5847 -2995 -5844
rect -2930 -5842 -2833 -5829
rect -2930 -5847 -2915 -5842
rect -3009 -5907 -2915 -5847
rect -3009 -5925 -2995 -5907
rect -3092 -5938 -2995 -5925
rect -2930 -5923 -2915 -5907
rect -2847 -5847 -2833 -5842
rect -2540 -5847 -2348 -5835
rect -2291 -5837 -2197 -5824
rect -2291 -5847 -2279 -5837
rect -2847 -5848 -2279 -5847
rect -2847 -5904 -2526 -5848
rect -2470 -5904 -2416 -5848
rect -2360 -5904 -2279 -5848
rect -2847 -5907 -2279 -5904
rect -2847 -5923 -2833 -5907
rect -2540 -5919 -2348 -5907
rect -2291 -5918 -2279 -5907
rect -2211 -5847 -2197 -5837
rect -1659 -5837 -1562 -5824
rect -1659 -5847 -1644 -5837
rect -2211 -5907 -1644 -5847
rect -2211 -5918 -2197 -5907
rect -2930 -5936 -2833 -5923
rect -2291 -5931 -2197 -5918
rect -1659 -5918 -1644 -5907
rect -1576 -5847 -1562 -5837
rect -1491 -5839 -1394 -5826
rect -1491 -5847 -1476 -5839
rect -1576 -5907 -1476 -5847
rect -1576 -5918 -1562 -5907
rect -1659 -5931 -1562 -5918
rect -1491 -5920 -1476 -5907
rect -1408 -5920 -1394 -5839
rect -1491 -5933 -1394 -5920
rect 337 -5939 449 -5922
rect 337 -6024 353 -5939
rect 435 -6024 449 -5939
rect -146 -6049 148 -6030
rect 337 -6038 449 -6024
rect -146 -6052 50 -6049
rect -1744 -6076 -1640 -6065
rect -1744 -6156 -1731 -6076
rect -1651 -6156 -1640 -6076
rect -1744 -6166 -1640 -6156
rect -146 -6137 -109 -6052
rect -27 -6134 50 -6052
rect 132 -6134 148 -6049
rect -27 -6137 148 -6134
rect -146 -6164 148 -6137
rect 793 -6164 890 -5713
rect -146 -6261 890 -6164
rect -2030 -6460 -1881 -6426
rect -2030 -6550 -2004 -6460
rect -1908 -6550 -1881 -6460
rect -2631 -6585 -2482 -6551
rect -2030 -6579 -1881 -6550
rect -2631 -6675 -2605 -6585
rect -2509 -6675 -2482 -6585
rect -2631 -6705 -2482 -6675
rect -2286 -6657 -2167 -6644
rect -2286 -6738 -2267 -6657
rect -2186 -6670 -2167 -6657
rect -424 -6663 -329 -6651
rect -424 -6670 -411 -6663
rect -2186 -6733 -411 -6670
rect -341 -6670 -329 -6663
rect -341 -6733 372 -6670
rect -2186 -6734 372 -6733
rect -2186 -6738 -2167 -6734
rect -2286 -6749 -2167 -6738
rect -424 -6745 -329 -6734
rect 127 -6824 229 -6811
rect 127 -6880 143 -6824
rect 215 -6880 229 -6824
rect 127 -6894 229 -6880
rect -184 -7047 -99 -7032
rect -184 -7129 -169 -7047
rect -113 -7129 -99 -7047
rect -184 -7142 -99 -7129
rect -3076 -7212 -2979 -7199
rect -3076 -7293 -3061 -7212
rect -2993 -7225 -2979 -7212
rect -2912 -7211 -2815 -7198
rect -2912 -7225 -2897 -7211
rect -2993 -7289 -2897 -7225
rect -2993 -7293 -2979 -7289
rect -3076 -7306 -2979 -7293
rect -2912 -7292 -2897 -7289
rect -2829 -7225 -2815 -7211
rect -2612 -7212 -2486 -7163
rect -2612 -7225 -2589 -7212
rect -2829 -7289 -2589 -7225
rect -2829 -7292 -2815 -7289
rect -2912 -7305 -2815 -7292
rect -2612 -7298 -2589 -7289
rect -2503 -7225 -2486 -7212
rect -2274 -7212 -2177 -7199
rect -2274 -7225 -2259 -7212
rect -2503 -7289 -2259 -7225
rect -2503 -7298 -2486 -7289
rect -2612 -7314 -2486 -7298
rect -2274 -7293 -2259 -7289
rect -2191 -7225 -2177 -7212
rect -1638 -7212 -1541 -7199
rect -1638 -7225 -1623 -7212
rect -2191 -7289 -1623 -7225
rect -2191 -7293 -2177 -7289
rect -2274 -7306 -2177 -7293
rect -1638 -7293 -1623 -7289
rect -1555 -7225 -1541 -7212
rect -1475 -7216 -1378 -7203
rect -1475 -7225 -1460 -7216
rect -1555 -7289 -1460 -7225
rect -1555 -7293 -1541 -7289
rect -1638 -7306 -1541 -7293
rect -1475 -7297 -1460 -7289
rect -1392 -7297 -1378 -7216
rect -1475 -7310 -1378 -7297
rect -185 -7232 -99 -7214
rect -185 -7314 -170 -7232
rect -114 -7314 -99 -7232
rect -185 -7330 -99 -7314
rect -2597 -7531 -2500 -7518
rect -2597 -7612 -2582 -7531
rect -2514 -7538 -2500 -7531
rect -1965 -7530 -1851 -7514
rect -1965 -7538 -1949 -7530
rect -2514 -7612 -1949 -7538
rect -1867 -7538 -1851 -7530
rect -1867 -7612 -732 -7538
rect -2597 -7659 -732 -7612
rect -2268 -7809 -2184 -7797
rect -2268 -7869 -2256 -7809
rect -2196 -7869 -2184 -7809
rect -2268 -7881 -2184 -7869
rect -3075 -8018 -2978 -8005
rect -3075 -8099 -3060 -8018
rect -2992 -8026 -2978 -8018
rect -2915 -8022 -2818 -8007
rect -2915 -8026 -2901 -8022
rect -2992 -8090 -2901 -8026
rect -2992 -8099 -2978 -8090
rect -3075 -8112 -2978 -8099
rect -2915 -8103 -2901 -8090
rect -2833 -8026 -2818 -8022
rect -2273 -8016 -2176 -8003
rect -2273 -8026 -2258 -8016
rect -2833 -8090 -2258 -8026
rect -2833 -8103 -2818 -8090
rect -2915 -8115 -2818 -8103
rect -2273 -8097 -2258 -8090
rect -2190 -8026 -2176 -8016
rect -1968 -8014 -1853 -7997
rect -1968 -8026 -1952 -8014
rect -2190 -8090 -1952 -8026
rect -2190 -8097 -2176 -8090
rect -2273 -8110 -2176 -8097
rect -1968 -8098 -1952 -8090
rect -1868 -8026 -1853 -8014
rect -1636 -8015 -1539 -8002
rect -1636 -8026 -1621 -8015
rect -1868 -8090 -1621 -8026
rect -1868 -8098 -1853 -8090
rect -1968 -8113 -1853 -8098
rect -1636 -8096 -1621 -8090
rect -1553 -8026 -1539 -8015
rect -1473 -8015 -1376 -8002
rect -1473 -8026 -1458 -8015
rect -1553 -8090 -1458 -8026
rect -1553 -8096 -1539 -8090
rect -1636 -8109 -1539 -8096
rect -1473 -8096 -1458 -8090
rect -1390 -8096 -1376 -8015
rect -1473 -8109 -1376 -8096
rect -2605 -8332 -2491 -8316
rect -2605 -8414 -2589 -8332
rect -2507 -8339 -2491 -8332
rect -1955 -8327 -1858 -8314
rect -1955 -8339 -1940 -8327
rect -2507 -8403 -1940 -8339
rect -2507 -8414 -2491 -8403
rect -2605 -8428 -2491 -8414
rect -1955 -8408 -1940 -8403
rect -1872 -8339 -1858 -8327
rect -1872 -8402 -962 -8339
rect -1872 -8408 -1858 -8402
rect -1955 -8421 -1858 -8408
rect -2268 -8610 -2184 -8598
rect -2268 -8670 -2256 -8610
rect -2196 -8670 -2184 -8610
rect -2268 -8682 -2184 -8670
rect -1025 -8664 -962 -8402
rect -796 -8346 -732 -7659
rect 148 -7897 211 -6894
rect 308 -7199 372 -6734
rect 1359 -7179 1509 -4715
rect 2191 -4800 2288 -4782
rect 2191 -4830 2208 -4800
rect 1920 -4864 2208 -4830
rect 2272 -4835 2288 -4800
rect 3053 -4809 3150 -4791
rect 3053 -4835 3070 -4809
rect 2272 -4864 3070 -4835
rect 1920 -4873 3070 -4864
rect 3134 -4873 3150 -4809
rect 1920 -4916 3150 -4873
rect 1920 -4957 2208 -4916
rect 1920 -6389 2047 -4957
rect 2191 -4980 2208 -4957
rect 2272 -4925 3150 -4916
rect 2272 -4943 3070 -4925
rect 2272 -4980 2288 -4943
rect 2191 -5121 2288 -4980
rect 3053 -4989 3070 -4943
rect 3134 -4989 3150 -4925
rect 3053 -5003 3150 -4989
rect 4781 -4927 4895 -4862
rect 4781 -4991 4807 -4927
rect 4871 -4975 4895 -4927
rect 5817 -4924 5959 -4854
rect 5817 -4975 5859 -4924
rect 4871 -4988 5859 -4975
rect 5923 -4988 5959 -4924
rect 4871 -4991 5959 -4988
rect 4781 -5040 5959 -4991
rect 4781 -5043 5859 -5040
rect 4781 -5107 4807 -5043
rect 4871 -5104 5859 -5043
rect 5923 -5104 5959 -5040
rect 4871 -5107 5959 -5104
rect 4781 -5144 5959 -5107
rect 4781 -5446 4895 -5144
rect 2829 -5522 2926 -5504
rect 2829 -5550 2846 -5522
rect 2273 -5586 2846 -5550
rect 2910 -5586 2926 -5522
rect 2273 -5638 2926 -5586
rect 2273 -5647 2846 -5638
rect 2273 -5877 2370 -5647
rect 2829 -5702 2846 -5647
rect 2910 -5702 2926 -5638
rect 2829 -5716 2926 -5702
rect 4781 -5510 4807 -5446
rect 4871 -5510 4895 -5446
rect 4781 -5562 4895 -5510
rect 4781 -5626 4807 -5562
rect 4871 -5626 4895 -5562
rect 4781 -5730 4895 -5626
rect 5372 -5408 5495 -5381
rect 5372 -5472 5411 -5408
rect 5475 -5472 5495 -5408
rect 5372 -5524 5495 -5472
rect 5372 -5588 5411 -5524
rect 5475 -5588 5495 -5524
rect 5372 -5857 5495 -5588
rect 2273 -5941 2290 -5877
rect 2354 -5911 2370 -5877
rect 2989 -5890 3146 -5872
rect 2354 -5941 2671 -5911
rect 2273 -5993 2671 -5941
rect 2273 -6057 2290 -5993
rect 2354 -6044 2671 -5993
rect 2354 -6057 2370 -6044
rect 2273 -6071 2370 -6057
rect 2538 -6317 2671 -6044
rect 2989 -5954 3018 -5890
rect 3082 -5926 3146 -5890
rect 3082 -5954 3382 -5926
rect 2989 -6006 3382 -5954
rect 2989 -6070 3018 -6006
rect 3082 -6054 3382 -6006
rect 3082 -6070 3146 -6054
rect 2989 -6091 3146 -6070
rect 1920 -6516 2263 -6389
rect 2538 -6450 3035 -6317
rect 2136 -6723 2263 -6516
rect 2076 -6755 2332 -6723
rect 2902 -6734 3035 -6450
rect 2076 -6826 2103 -6755
rect 2174 -6757 2332 -6755
rect 2174 -6768 2239 -6757
rect 2076 -6828 2127 -6826
rect 2187 -6828 2239 -6768
rect 2310 -6828 2332 -6757
rect 2868 -6749 3069 -6734
rect 2868 -6809 2882 -6749
rect 2942 -6809 2996 -6749
rect 3056 -6809 3069 -6749
rect 2868 -6823 3069 -6809
rect 2076 -6841 2332 -6828
rect 2113 -6842 2314 -6841
rect 3254 -7061 3382 -6054
rect 3905 -5980 5495 -5857
rect 5817 -5443 5959 -5144
rect 5817 -5507 5859 -5443
rect 5923 -5507 5959 -5443
rect 5817 -5559 5959 -5507
rect 5817 -5623 5859 -5559
rect 5923 -5623 5959 -5559
rect 5817 -5759 5959 -5623
rect 5817 -5901 6306 -5759
rect 3060 -7179 3382 -7061
rect 1359 -7189 3382 -7179
rect 3499 -7010 3596 -6992
rect 3499 -7074 3516 -7010
rect 3580 -7038 3596 -7010
rect 3905 -7038 4028 -5980
rect 4941 -6430 5155 -6414
rect 4941 -6494 4958 -6430
rect 5022 -6494 5078 -6430
rect 5142 -6494 5155 -6430
rect 4941 -6550 5155 -6494
rect 4941 -6614 4958 -6550
rect 5022 -6614 5078 -6550
rect 5142 -6614 5155 -6550
rect 4941 -6628 5155 -6614
rect 5514 -6433 5728 -6417
rect 5514 -6497 5531 -6433
rect 5595 -6497 5651 -6433
rect 5715 -6497 5728 -6433
rect 5514 -6553 5728 -6497
rect 5514 -6617 5531 -6553
rect 5595 -6617 5651 -6553
rect 5715 -6617 5728 -6553
rect 3580 -7074 4028 -7038
rect 3499 -7126 4028 -7074
rect 298 -7215 381 -7199
rect 298 -7287 312 -7215
rect 368 -7287 381 -7215
rect 298 -7301 381 -7287
rect 1359 -7329 3188 -7189
rect 3499 -7190 3516 -7126
rect 3580 -7161 4028 -7126
rect 3580 -7190 3596 -7161
rect 3499 -7204 3596 -7190
rect 3060 -7413 3188 -7329
rect 4962 -7232 5076 -6628
rect 5514 -6631 5728 -6617
rect 4962 -7296 4986 -7232
rect 5050 -7296 5076 -7232
rect 4962 -7348 5076 -7296
rect 4962 -7412 4986 -7348
rect 5050 -7412 5076 -7348
rect 3025 -7428 3226 -7413
rect 3025 -7488 3039 -7428
rect 3099 -7488 3153 -7428
rect 3213 -7488 3226 -7428
rect 3025 -7502 3226 -7488
rect 297 -7677 387 -7665
rect 297 -7743 309 -7677
rect 375 -7743 387 -7677
rect 297 -7755 387 -7743
rect 4962 -7819 5076 -7412
rect 4962 -7883 4986 -7819
rect 5050 -7883 5076 -7819
rect -190 -7934 -93 -7912
rect -190 -8004 -177 -7934
rect -107 -8004 -93 -7934
rect 139 -7913 222 -7897
rect 139 -7985 153 -7913
rect 209 -7985 222 -7913
rect 4962 -7935 5076 -7883
rect 139 -7999 222 -7985
rect 292 -7995 389 -7977
rect -190 -8074 -93 -8004
rect -190 -8144 -175 -8074
rect -105 -8079 -93 -8074
rect 292 -8059 309 -7995
rect 373 -8059 389 -7995
rect 292 -8079 389 -8059
rect -105 -8111 389 -8079
rect -105 -8140 309 -8111
rect -105 -8144 -93 -8140
rect -190 -8162 -93 -8144
rect 292 -8175 309 -8140
rect 373 -8175 389 -8111
rect 4962 -7999 4986 -7935
rect 5050 -7999 5076 -7935
rect 292 -8189 389 -8175
rect 778 -8157 863 -8141
rect 778 -8229 793 -8157
rect 849 -8229 863 -8157
rect -422 -8293 -327 -8283
rect -183 -8293 -100 -8279
rect -422 -8295 -100 -8293
rect -796 -8506 -730 -8346
rect -422 -8365 -409 -8295
rect -339 -8365 -169 -8295
rect -422 -8367 -169 -8365
rect -113 -8299 -100 -8295
rect 778 -8299 863 -8229
rect -113 -8300 863 -8299
rect -113 -8367 793 -8300
rect -422 -8368 793 -8367
rect -422 -8377 -327 -8368
rect -183 -8370 793 -8368
rect -183 -8381 -100 -8370
rect 778 -8372 793 -8370
rect 849 -8372 863 -8300
rect 778 -8387 863 -8372
rect 4962 -8338 5076 -7999
rect 4962 -8402 4986 -8338
rect 5050 -8402 5076 -8338
rect 4962 -8454 5076 -8402
rect 134 -8505 217 -8489
rect 134 -8506 148 -8505
rect -796 -8572 148 -8506
rect 134 -8577 148 -8572
rect 204 -8506 217 -8505
rect 460 -8504 543 -8488
rect 460 -8506 474 -8504
rect 204 -8572 474 -8506
rect 204 -8577 217 -8572
rect 134 -8591 217 -8577
rect 460 -8576 474 -8572
rect 530 -8576 543 -8504
rect 4962 -8518 4986 -8454
rect 5050 -8518 5076 -8454
rect 460 -8590 543 -8576
rect 892 -8588 982 -8576
rect 4962 -8583 5076 -8518
rect 5568 -7233 5682 -6631
rect 5568 -7297 5592 -7233
rect 5656 -7297 5682 -7233
rect 5568 -7349 5682 -7297
rect 5568 -7413 5592 -7349
rect 5656 -7413 5682 -7349
rect 5568 -7820 5682 -7413
rect 5568 -7884 5592 -7820
rect 5656 -7884 5682 -7820
rect 5568 -7936 5682 -7884
rect 5568 -8000 5592 -7936
rect 5656 -8000 5682 -7936
rect 5568 -8339 5682 -8000
rect 5568 -8403 5592 -8339
rect 5656 -8403 5682 -8339
rect 5568 -8455 5682 -8403
rect 5568 -8519 5592 -8455
rect 5656 -8519 5682 -8455
rect 5568 -8584 5682 -8519
rect 6164 -7231 6306 -5901
rect 6729 -6394 6943 -6378
rect 7368 -6381 7742 -3296
rect 8406 -3445 8540 -2487
rect 8727 641 8861 707
rect 8727 577 8763 641
rect 8827 577 8861 641
rect 8727 525 8861 577
rect 8727 461 8763 525
rect 8827 461 8861 525
rect 8727 -99 8861 461
rect 8727 -163 8763 -99
rect 8827 -163 8861 -99
rect 8727 -215 8861 -163
rect 8727 -279 8763 -215
rect 8827 -279 8861 -215
rect 8727 -828 8861 -279
rect 8727 -892 8763 -828
rect 8827 -892 8861 -828
rect 8727 -944 8861 -892
rect 8727 -1008 8763 -944
rect 8827 -1008 8861 -944
rect 8727 -1568 8861 -1008
rect 8727 -1632 8763 -1568
rect 8827 -1632 8861 -1568
rect 8727 -1684 8861 -1632
rect 8727 -1748 8763 -1684
rect 8827 -1748 8861 -1684
rect 8727 -2308 8861 -1748
rect 8727 -2372 8763 -2308
rect 8827 -2372 8861 -2308
rect 8727 -2424 8861 -2372
rect 8727 -2488 8763 -2424
rect 8827 -2488 8861 -2424
rect 8727 -3445 8861 -2488
rect 9044 671 9178 704
rect 9044 607 9083 671
rect 9147 607 9178 671
rect 9044 555 9178 607
rect 9044 491 9083 555
rect 9147 491 9178 555
rect 9044 -80 9178 491
rect 9044 -144 9083 -80
rect 9147 -144 9178 -80
rect 9044 -196 9178 -144
rect 9044 -260 9083 -196
rect 9147 -260 9178 -196
rect 9044 -812 9178 -260
rect 9044 -876 9083 -812
rect 9147 -876 9178 -812
rect 9044 -928 9178 -876
rect 9044 -992 9083 -928
rect 9147 -992 9178 -928
rect 9044 -1554 9178 -992
rect 9044 -1618 9083 -1554
rect 9147 -1618 9178 -1554
rect 9044 -1670 9178 -1618
rect 9044 -1734 9083 -1670
rect 9147 -1734 9178 -1670
rect 9044 -2314 9178 -1734
rect 9044 -2378 9083 -2314
rect 9147 -2378 9178 -2314
rect 9044 -2430 9178 -2378
rect 9044 -2494 9083 -2430
rect 9147 -2494 9178 -2430
rect 9044 -3105 9178 -2494
rect 9365 658 9499 709
rect 9365 594 9403 658
rect 9467 594 9499 658
rect 9365 542 9499 594
rect 9365 478 9403 542
rect 9467 478 9499 542
rect 9365 -101 9499 478
rect 9365 -165 9403 -101
rect 9467 -165 9499 -101
rect 9365 -217 9499 -165
rect 9365 -281 9403 -217
rect 9467 -281 9499 -217
rect 9365 -837 9499 -281
rect 9365 -901 9403 -837
rect 9467 -901 9499 -837
rect 9365 -953 9499 -901
rect 9365 -1017 9403 -953
rect 9467 -1017 9499 -953
rect 9365 -1562 9499 -1017
rect 9365 -1626 9403 -1562
rect 9467 -1626 9499 -1562
rect 9365 -1678 9499 -1626
rect 9365 -1742 9403 -1678
rect 9467 -1742 9499 -1678
rect 9365 -2310 9499 -1742
rect 9365 -2374 9403 -2310
rect 9467 -2374 9499 -2310
rect 9365 -2426 9499 -2374
rect 9365 -2490 9403 -2426
rect 9467 -2490 9499 -2426
rect 9000 -3119 9215 -3105
rect 9000 -3183 9017 -3119
rect 9081 -3183 9137 -3119
rect 9201 -3183 9215 -3119
rect 9000 -3239 9215 -3183
rect 9000 -3303 9017 -3239
rect 9081 -3303 9137 -3239
rect 9201 -3303 9215 -3239
rect 9000 -3317 9215 -3303
rect 9365 -3445 9499 -2490
rect 9686 655 9820 712
rect 9686 591 9723 655
rect 9787 591 9820 655
rect 9686 539 9820 591
rect 9686 475 9723 539
rect 9787 475 9820 539
rect 9686 -116 9820 475
rect 9686 -180 9723 -116
rect 9787 -180 9820 -116
rect 9686 -232 9820 -180
rect 9686 -296 9723 -232
rect 9787 -296 9820 -232
rect 9686 -841 9820 -296
rect 9686 -905 9723 -841
rect 9787 -905 9820 -841
rect 9686 -957 9820 -905
rect 9686 -1021 9723 -957
rect 9787 -1021 9820 -957
rect 9686 -1565 9820 -1021
rect 11070 -1254 11746 -1239
rect 11070 -1335 11088 -1254
rect 11169 -1335 11228 -1254
rect 11309 -1335 11368 -1254
rect 11449 -1335 11508 -1254
rect 11589 -1335 11648 -1254
rect 11729 -1335 11746 -1254
rect 11070 -1349 11746 -1335
rect 9686 -1629 9723 -1565
rect 9787 -1629 9820 -1565
rect 9686 -1681 9820 -1629
rect 9686 -1745 9723 -1681
rect 9787 -1745 9820 -1681
rect 9686 -2313 9820 -1745
rect 9686 -2377 9723 -2313
rect 9787 -2377 9820 -2313
rect 9686 -2429 9820 -2377
rect 9686 -2493 9723 -2429
rect 9787 -2493 9820 -2429
rect 9686 -3445 9820 -2493
rect 11077 -2683 11750 -2666
rect 11077 -2764 11094 -2683
rect 11175 -2764 11234 -2683
rect 11315 -2764 11374 -2683
rect 11455 -2764 11514 -2683
rect 11595 -2764 11654 -2683
rect 11735 -2764 11750 -2683
rect 11077 -2778 11750 -2764
rect 8200 -3460 10133 -3445
rect 8200 -3524 8378 -3460
rect 8442 -3524 8498 -3460
rect 8562 -3524 8706 -3460
rect 8770 -3524 8826 -3460
rect 8890 -3461 9660 -3460
rect 8890 -3524 9334 -3461
rect 8200 -3525 9334 -3524
rect 9398 -3525 9454 -3461
rect 9518 -3524 9660 -3461
rect 9724 -3524 9780 -3460
rect 9844 -3524 10133 -3460
rect 9518 -3525 10133 -3524
rect 8200 -3580 10133 -3525
rect 8200 -3644 8378 -3580
rect 8442 -3644 8498 -3580
rect 8562 -3644 8706 -3580
rect 8770 -3644 8826 -3580
rect 8890 -3581 9660 -3580
rect 8890 -3644 9334 -3581
rect 8200 -3645 9334 -3644
rect 9398 -3645 9454 -3581
rect 9518 -3644 9660 -3581
rect 9724 -3644 9780 -3580
rect 9844 -3644 10133 -3580
rect 9518 -3645 10133 -3644
rect 8200 -3782 10133 -3645
rect 8200 -5340 8537 -3782
rect 11255 -4942 11469 -4932
rect 9195 -4948 11469 -4942
rect 9195 -4962 11272 -4948
rect 9195 -4963 10221 -4962
rect 9195 -4966 9890 -4963
rect 9195 -4967 9573 -4966
rect 9195 -5034 9259 -4967
rect 9324 -5033 9573 -4967
rect 9638 -5030 9890 -4966
rect 9955 -5029 10221 -4963
rect 10286 -4963 11272 -4962
rect 10286 -5029 10540 -4963
rect 9955 -5030 10540 -5029
rect 10605 -5012 11272 -4963
rect 11336 -5012 11392 -4948
rect 11456 -5012 11469 -4948
rect 10605 -5030 11469 -5012
rect 9638 -5033 11469 -5030
rect 9324 -5034 11469 -5033
rect 9195 -5064 11469 -5034
rect 11255 -5068 11469 -5064
rect 11255 -5132 11272 -5068
rect 11336 -5132 11392 -5068
rect 11456 -5132 11469 -5068
rect 11255 -5146 11469 -5132
rect 9246 -5333 9343 -5319
rect 9246 -5340 9262 -5333
rect 8200 -5397 9262 -5340
rect 9326 -5340 9343 -5333
rect 9566 -5333 9663 -5319
rect 9566 -5340 9582 -5333
rect 9326 -5397 9582 -5340
rect 9646 -5340 9663 -5333
rect 9887 -5333 9984 -5319
rect 9887 -5340 9903 -5333
rect 9646 -5397 9903 -5340
rect 9967 -5340 9984 -5333
rect 10207 -5336 10304 -5322
rect 10207 -5340 10223 -5336
rect 9967 -5397 10223 -5340
rect 8200 -5400 10223 -5397
rect 10287 -5340 10304 -5336
rect 10527 -5334 10624 -5320
rect 10527 -5340 10543 -5334
rect 10287 -5398 10543 -5340
rect 10607 -5398 10624 -5334
rect 10287 -5400 10624 -5398
rect 8200 -5449 10624 -5400
rect 8200 -5504 9262 -5449
rect 8200 -6070 8537 -5504
rect 9246 -5513 9262 -5504
rect 9326 -5504 9582 -5449
rect 9326 -5513 9343 -5504
rect 9246 -5531 9343 -5513
rect 9566 -5513 9582 -5504
rect 9646 -5504 9903 -5449
rect 9646 -5513 9663 -5504
rect 9566 -5531 9663 -5513
rect 9887 -5513 9903 -5504
rect 9967 -5450 10624 -5449
rect 9967 -5452 10543 -5450
rect 9967 -5504 10223 -5452
rect 9967 -5513 9984 -5504
rect 9887 -5531 9984 -5513
rect 10207 -5516 10223 -5504
rect 10287 -5504 10543 -5452
rect 10287 -5516 10304 -5504
rect 10207 -5534 10304 -5516
rect 10527 -5514 10543 -5504
rect 10607 -5514 10624 -5450
rect 10527 -5532 10624 -5514
rect 9248 -6059 9345 -6045
rect 9248 -6070 9264 -6059
rect 8200 -6123 9264 -6070
rect 9328 -6070 9345 -6059
rect 9568 -6061 9665 -6047
rect 9568 -6070 9584 -6061
rect 9328 -6123 9584 -6070
rect 8200 -6125 9584 -6123
rect 9648 -6070 9665 -6061
rect 9888 -6063 9985 -6049
rect 9888 -6070 9904 -6063
rect 9648 -6125 9904 -6070
rect 8200 -6127 9904 -6125
rect 9968 -6070 9985 -6063
rect 10208 -6063 10305 -6049
rect 10208 -6070 10224 -6063
rect 9968 -6127 10224 -6070
rect 10288 -6070 10305 -6063
rect 10525 -6063 10622 -6049
rect 10525 -6070 10541 -6063
rect 10288 -6127 10541 -6070
rect 10605 -6127 10622 -6063
rect 8200 -6175 10622 -6127
rect 8200 -6234 9264 -6175
rect 6729 -6458 6746 -6394
rect 6810 -6458 6866 -6394
rect 6930 -6458 6943 -6394
rect 6729 -6514 6943 -6458
rect 6729 -6578 6746 -6514
rect 6810 -6578 6866 -6514
rect 6930 -6578 6943 -6514
rect 6729 -6592 6943 -6578
rect 7330 -6397 7784 -6381
rect 7330 -6461 7347 -6397
rect 7411 -6461 7467 -6397
rect 7531 -6461 7587 -6397
rect 7651 -6461 7707 -6397
rect 7771 -6461 7784 -6397
rect 7330 -6517 7784 -6461
rect 7330 -6581 7347 -6517
rect 7411 -6581 7467 -6517
rect 7531 -6581 7587 -6517
rect 7651 -6581 7707 -6517
rect 7771 -6581 7784 -6517
rect 6164 -7295 6201 -7231
rect 6265 -7295 6306 -7231
rect 6164 -7347 6306 -7295
rect 6164 -7411 6201 -7347
rect 6265 -7411 6306 -7347
rect 6164 -7818 6306 -7411
rect 6164 -7882 6201 -7818
rect 6265 -7882 6306 -7818
rect 6164 -7934 6306 -7882
rect 6164 -7998 6201 -7934
rect 6265 -7998 6306 -7934
rect 6164 -8337 6306 -7998
rect 6164 -8401 6201 -8337
rect 6265 -8401 6306 -8337
rect 6164 -8453 6306 -8401
rect 6164 -8517 6201 -8453
rect 6265 -8517 6306 -8453
rect -23 -8661 60 -8645
rect -23 -8664 -9 -8661
rect -1025 -8729 -9 -8664
rect -23 -8733 -9 -8729
rect 47 -8664 60 -8661
rect 620 -8661 703 -8645
rect 620 -8664 634 -8661
rect 47 -8729 634 -8664
rect 47 -8733 60 -8729
rect -23 -8747 60 -8733
rect 620 -8733 634 -8729
rect 690 -8733 703 -8661
rect 892 -8654 904 -8588
rect 970 -8654 982 -8588
rect 6164 -8595 6306 -8517
rect 6786 -7234 6900 -6592
rect 7330 -6595 7784 -6581
rect 6786 -7298 6810 -7234
rect 6874 -7298 6900 -7234
rect 6786 -7350 6900 -7298
rect 6786 -7414 6810 -7350
rect 6874 -7414 6900 -7350
rect 6786 -7821 6900 -7414
rect 6786 -7885 6810 -7821
rect 6874 -7885 6900 -7821
rect 6786 -7937 6900 -7885
rect 6786 -8001 6810 -7937
rect 6874 -8001 6900 -7937
rect 6786 -8340 6900 -8001
rect 6786 -8404 6810 -8340
rect 6874 -8404 6900 -8340
rect 6786 -8456 6900 -8404
rect 6786 -8520 6810 -8456
rect 6874 -8520 6900 -8456
rect 6786 -8585 6900 -8520
rect 7389 -7242 7503 -6595
rect 7389 -7306 7413 -7242
rect 7477 -7306 7503 -7242
rect 7389 -7358 7503 -7306
rect 7389 -7422 7413 -7358
rect 7477 -7422 7503 -7358
rect 7389 -7829 7503 -7422
rect 7389 -7893 7413 -7829
rect 7477 -7893 7503 -7829
rect 7389 -7945 7503 -7893
rect 7389 -8009 7413 -7945
rect 7477 -8009 7503 -7945
rect 7389 -8348 7503 -8009
rect 7389 -8412 7413 -8348
rect 7477 -8412 7503 -8348
rect 7389 -8464 7503 -8412
rect 7389 -8528 7413 -8464
rect 7477 -8528 7503 -8464
rect 7389 -8593 7503 -8528
rect 8200 -6801 8537 -6234
rect 9248 -6239 9264 -6234
rect 9328 -6177 10622 -6175
rect 9328 -6234 9584 -6177
rect 9328 -6239 9345 -6234
rect 9248 -6257 9345 -6239
rect 9568 -6241 9584 -6234
rect 9648 -6179 10622 -6177
rect 9648 -6234 9904 -6179
rect 9648 -6241 9665 -6234
rect 9568 -6259 9665 -6241
rect 9888 -6243 9904 -6234
rect 9968 -6234 10224 -6179
rect 9968 -6243 9985 -6234
rect 9888 -6261 9985 -6243
rect 10208 -6243 10224 -6234
rect 10288 -6234 10541 -6179
rect 10288 -6243 10305 -6234
rect 10208 -6261 10305 -6243
rect 10525 -6243 10541 -6234
rect 10605 -6243 10622 -6179
rect 10525 -6261 10622 -6243
rect 9246 -6790 9343 -6776
rect 9246 -6801 9262 -6790
rect 8200 -6854 9262 -6801
rect 9326 -6801 9343 -6790
rect 9568 -6790 9665 -6776
rect 9568 -6801 9584 -6790
rect 9326 -6854 9584 -6801
rect 9648 -6801 9665 -6790
rect 9887 -6790 9984 -6776
rect 9887 -6801 9903 -6790
rect 9648 -6854 9903 -6801
rect 9967 -6801 9984 -6790
rect 10207 -6792 10304 -6778
rect 10207 -6801 10223 -6792
rect 9967 -6854 10223 -6801
rect 8200 -6856 10223 -6854
rect 10287 -6801 10304 -6792
rect 10527 -6792 10624 -6778
rect 10527 -6801 10543 -6792
rect 10287 -6856 10543 -6801
rect 10607 -6856 10624 -6792
rect 8200 -6906 10624 -6856
rect 8200 -6965 9262 -6906
rect 8200 -8340 8537 -6965
rect 9246 -6970 9262 -6965
rect 9326 -6965 9584 -6906
rect 9326 -6970 9343 -6965
rect 9246 -6988 9343 -6970
rect 9568 -6970 9584 -6965
rect 9648 -6965 9903 -6906
rect 9648 -6970 9665 -6965
rect 9568 -6988 9665 -6970
rect 9887 -6970 9903 -6965
rect 9967 -6908 10624 -6906
rect 9967 -6965 10223 -6908
rect 9967 -6970 9984 -6965
rect 9887 -6988 9984 -6970
rect 10207 -6972 10223 -6965
rect 10287 -6965 10543 -6908
rect 10287 -6972 10304 -6965
rect 10207 -6990 10304 -6972
rect 10527 -6972 10543 -6965
rect 10607 -6972 10624 -6908
rect 10527 -6990 10624 -6972
rect 11274 -7226 11431 -5146
rect 9193 -7252 11431 -7226
rect 9193 -7255 10537 -7252
rect 9193 -7258 9586 -7255
rect 9193 -7325 9258 -7258
rect 9323 -7322 9586 -7258
rect 9651 -7256 10537 -7255
rect 9651 -7322 9896 -7256
rect 9323 -7323 9896 -7322
rect 9961 -7323 10222 -7256
rect 10287 -7319 10537 -7256
rect 10602 -7319 11431 -7252
rect 10287 -7323 11431 -7319
rect 9323 -7325 11431 -7323
rect 9193 -7348 11431 -7325
rect 11274 -7538 11431 -7348
rect 11245 -7554 11459 -7538
rect 11245 -7618 11262 -7554
rect 11326 -7618 11382 -7554
rect 11446 -7618 11459 -7554
rect 11245 -7674 11459 -7618
rect 11245 -7738 11262 -7674
rect 11326 -7738 11382 -7674
rect 11446 -7738 11459 -7674
rect 11245 -7752 11459 -7738
rect 11274 -7942 11431 -7752
rect 9195 -7962 11433 -7942
rect 9195 -7963 10221 -7962
rect 9195 -7966 9890 -7963
rect 9195 -7967 9573 -7966
rect 9195 -8034 9259 -7967
rect 9324 -8033 9573 -7967
rect 9638 -8030 9890 -7966
rect 9955 -8029 10221 -7963
rect 10286 -7963 11433 -7962
rect 10286 -8029 10540 -7963
rect 9955 -8030 10540 -8029
rect 10605 -8030 11433 -7963
rect 9638 -8033 11433 -8030
rect 9324 -8034 11433 -8033
rect 9195 -8064 11433 -8034
rect 9246 -8333 9343 -8319
rect 9246 -8340 9262 -8333
rect 8200 -8397 9262 -8340
rect 9326 -8340 9343 -8333
rect 9566 -8333 9663 -8319
rect 9566 -8340 9582 -8333
rect 9326 -8397 9582 -8340
rect 9646 -8340 9663 -8333
rect 9887 -8333 9984 -8319
rect 9887 -8340 9903 -8333
rect 9646 -8397 9903 -8340
rect 9967 -8340 9984 -8333
rect 10207 -8336 10304 -8322
rect 10207 -8340 10223 -8336
rect 9967 -8397 10223 -8340
rect 8200 -8400 10223 -8397
rect 10287 -8340 10304 -8336
rect 10527 -8334 10624 -8320
rect 10527 -8340 10543 -8334
rect 10287 -8398 10543 -8340
rect 10607 -8398 10624 -8334
rect 10287 -8400 10624 -8398
rect 8200 -8449 10624 -8400
rect 8200 -8504 9262 -8449
rect 892 -8666 982 -8654
rect 620 -8747 703 -8733
rect -3077 -8818 -2980 -8805
rect -3077 -8899 -3062 -8818
rect -2994 -8827 -2980 -8818
rect -2918 -8818 -2821 -8805
rect -2918 -8827 -2903 -8818
rect -2994 -8891 -2903 -8827
rect -2994 -8899 -2980 -8891
rect -3077 -8912 -2980 -8899
rect -2918 -8899 -2903 -8891
rect -2835 -8827 -2821 -8818
rect -2276 -8816 -2179 -8803
rect -2276 -8827 -2261 -8816
rect -2835 -8891 -2261 -8827
rect -2835 -8899 -2821 -8891
rect -2918 -8912 -2821 -8899
rect -2276 -8897 -2261 -8891
rect -2193 -8827 -2179 -8816
rect -1965 -8816 -1853 -8802
rect -1965 -8827 -1952 -8816
rect -2193 -8891 -1952 -8827
rect -2193 -8897 -2179 -8891
rect -2276 -8910 -2179 -8897
rect -1965 -8902 -1952 -8891
rect -1866 -8827 -1853 -8816
rect -1637 -8816 -1540 -8803
rect -1637 -8827 -1622 -8816
rect -1866 -8891 -1622 -8827
rect -1866 -8902 -1853 -8891
rect -1965 -8915 -1853 -8902
rect -1637 -8897 -1622 -8891
rect -1554 -8827 -1540 -8816
rect -1475 -8815 -1378 -8802
rect -1475 -8827 -1460 -8815
rect -1554 -8891 -1460 -8827
rect -1554 -8897 -1540 -8891
rect -1637 -8910 -1540 -8897
rect -1475 -8896 -1460 -8891
rect -1392 -8896 -1378 -8815
rect -1475 -8909 -1378 -8896
rect -189 -8941 -92 -8921
rect -189 -9011 -175 -8941
rect -105 -9011 -92 -8941
rect -189 -9081 -92 -9011
rect 290 -8975 390 -8957
rect 290 -9031 304 -8975
rect 376 -9031 390 -8975
rect -189 -9093 -91 -9081
rect -2607 -9133 -2493 -9117
rect -2607 -9215 -2591 -9133
rect -2509 -9140 -2493 -9133
rect -1955 -9128 -1858 -9115
rect -1955 -9140 -1940 -9128
rect -2509 -9204 -1940 -9140
rect -2509 -9215 -2493 -9204
rect -2607 -9229 -2493 -9215
rect -1955 -9209 -1940 -9204
rect -1872 -9209 -1858 -9128
rect -189 -9163 -173 -9093
rect -103 -9096 -91 -9093
rect 290 -9096 390 -9031
rect -103 -9098 390 -9096
rect -103 -9154 304 -9098
rect 376 -9154 390 -9098
rect 8200 -9070 8537 -8504
rect 9246 -8513 9262 -8504
rect 9326 -8504 9582 -8449
rect 9326 -8513 9343 -8504
rect 9246 -8531 9343 -8513
rect 9566 -8513 9582 -8504
rect 9646 -8504 9903 -8449
rect 9646 -8513 9663 -8504
rect 9566 -8531 9663 -8513
rect 9887 -8513 9903 -8504
rect 9967 -8450 10624 -8449
rect 9967 -8452 10543 -8450
rect 9967 -8504 10223 -8452
rect 9967 -8513 9984 -8504
rect 9887 -8531 9984 -8513
rect 10207 -8516 10223 -8504
rect 10287 -8504 10543 -8452
rect 10287 -8516 10304 -8504
rect 10207 -8534 10304 -8516
rect 10527 -8514 10543 -8504
rect 10607 -8514 10624 -8450
rect 10527 -8532 10624 -8514
rect 9248 -9059 9345 -9045
rect 9248 -9070 9264 -9059
rect 8200 -9123 9264 -9070
rect 9328 -9070 9345 -9059
rect 9568 -9061 9665 -9047
rect 9568 -9070 9584 -9061
rect 9328 -9123 9584 -9070
rect 8200 -9125 9584 -9123
rect 9648 -9070 9665 -9061
rect 9888 -9063 9985 -9049
rect 9888 -9070 9904 -9063
rect 9648 -9125 9904 -9070
rect 8200 -9127 9904 -9125
rect 9968 -9070 9985 -9063
rect 10208 -9063 10305 -9049
rect 10208 -9070 10224 -9063
rect 9968 -9127 10224 -9070
rect 10288 -9070 10305 -9063
rect 10525 -9063 10622 -9049
rect 10525 -9070 10541 -9063
rect 10288 -9127 10541 -9070
rect 10605 -9127 10622 -9063
rect -103 -9157 390 -9154
rect -103 -9163 -91 -9157
rect -189 -9175 -91 -9163
rect 288 -9168 390 -9157
rect -189 -9178 -92 -9175
rect 1893 -9177 2701 -9143
rect -1955 -9222 -1858 -9209
rect 457 -9228 540 -9212
rect 457 -9300 471 -9228
rect 527 -9300 540 -9228
rect 457 -9314 540 -9300
rect 1893 -9241 1928 -9177
rect 1992 -9179 2701 -9177
rect 1992 -9241 2073 -9179
rect 1893 -9243 2073 -9241
rect 2137 -9243 2207 -9179
rect 2271 -9243 2701 -9179
rect 1893 -9303 2701 -9243
rect -2269 -9410 -2185 -9398
rect -2269 -9470 -2257 -9410
rect -2197 -9470 -2185 -9410
rect -2269 -9482 -2185 -9470
rect 288 -9506 378 -9494
rect 288 -9572 300 -9506
rect 366 -9572 378 -9506
rect 288 -9584 378 -9572
rect -3075 -9616 -2978 -9603
rect -3075 -9697 -3060 -9616
rect -2992 -9628 -2978 -9616
rect -2913 -9615 -2816 -9602
rect -2913 -9628 -2898 -9615
rect -2992 -9692 -2898 -9628
rect -2992 -9697 -2978 -9692
rect -3075 -9710 -2978 -9697
rect -2913 -9696 -2898 -9692
rect -2830 -9628 -2816 -9615
rect -2604 -9616 -2491 -9600
rect -2604 -9628 -2591 -9616
rect -2830 -9692 -2591 -9628
rect -2830 -9696 -2816 -9692
rect -2913 -9709 -2816 -9696
rect -2604 -9702 -2591 -9692
rect -2505 -9628 -2491 -9616
rect -2275 -9616 -2178 -9603
rect -2275 -9628 -2260 -9616
rect -2505 -9692 -2260 -9628
rect -2505 -9702 -2491 -9692
rect -2604 -9719 -2491 -9702
rect -2275 -9697 -2260 -9692
rect -2192 -9628 -2178 -9616
rect -1635 -9619 -1538 -9606
rect -1635 -9628 -1620 -9619
rect -2192 -9692 -1620 -9628
rect -2192 -9697 -2178 -9692
rect -2275 -9710 -2178 -9697
rect -1635 -9700 -1620 -9692
rect -1552 -9628 -1538 -9619
rect -1478 -9617 -1381 -9604
rect -1478 -9628 -1463 -9617
rect -1552 -9692 -1463 -9628
rect -1552 -9700 -1538 -9692
rect -1635 -9713 -1538 -9700
rect -1478 -9698 -1463 -9692
rect -1395 -9698 -1381 -9617
rect -1478 -9711 -1381 -9698
rect -425 -9834 -330 -9822
rect 299 -9834 382 -9819
rect -425 -9904 -412 -9834
rect -342 -9835 382 -9834
rect -342 -9904 313 -9835
rect -425 -9907 313 -9904
rect 369 -9907 382 -9835
rect -425 -9908 382 -9907
rect -2596 -9931 -2499 -9918
rect -2596 -10012 -2581 -9931
rect -2513 -9941 -2499 -9931
rect -1963 -9931 -1849 -9915
rect -425 -9916 -330 -9908
rect -1963 -9941 -1947 -9931
rect -2513 -10005 -1947 -9941
rect -2513 -10012 -2499 -10005
rect -2596 -10025 -2499 -10012
rect -1963 -10013 -1947 -10005
rect -1865 -10013 -1849 -9931
rect 299 -9970 382 -9908
rect -1963 -10027 -1849 -10013
rect -184 -9998 -99 -9980
rect -184 -10054 -169 -9998
rect -113 -10054 -99 -9998
rect -184 -10112 -99 -10054
rect 299 -10042 313 -9970
rect 369 -10042 382 -9970
rect 299 -10055 382 -10042
rect -184 -10168 -169 -10112
rect -113 -10168 -99 -10112
rect -184 -10184 -99 -10168
rect 469 -10351 529 -9314
rect 1861 -9461 2302 -9412
rect 1861 -9463 2066 -9461
rect 1861 -9527 1921 -9463
rect 1985 -9525 2066 -9463
rect 2130 -9525 2200 -9461
rect 2264 -9525 2302 -9461
rect 1985 -9527 2302 -9525
rect 1861 -9548 2302 -9527
rect 444 -10364 546 -10351
rect 444 -10420 460 -10364
rect 532 -10420 546 -10364
rect 444 -10434 546 -10420
rect 2023 -10530 2183 -9548
rect 2541 -10264 2701 -9303
rect 8200 -9175 10622 -9127
rect 8200 -9234 9264 -9175
rect 8200 -9801 8537 -9234
rect 9248 -9239 9264 -9234
rect 9328 -9177 10622 -9175
rect 9328 -9234 9584 -9177
rect 9328 -9239 9345 -9234
rect 9248 -9257 9345 -9239
rect 9568 -9241 9584 -9234
rect 9648 -9179 10622 -9177
rect 9648 -9234 9904 -9179
rect 9648 -9241 9665 -9234
rect 9568 -9259 9665 -9241
rect 9888 -9243 9904 -9234
rect 9968 -9234 10224 -9179
rect 9968 -9243 9985 -9234
rect 9888 -9261 9985 -9243
rect 10208 -9243 10224 -9234
rect 10288 -9234 10541 -9179
rect 10288 -9243 10305 -9234
rect 10208 -9261 10305 -9243
rect 10525 -9243 10541 -9234
rect 10605 -9243 10622 -9179
rect 10525 -9261 10622 -9243
rect 9246 -9790 9343 -9776
rect 9246 -9801 9262 -9790
rect 8200 -9854 9262 -9801
rect 9326 -9801 9343 -9790
rect 9568 -9790 9665 -9776
rect 9568 -9801 9584 -9790
rect 9326 -9854 9584 -9801
rect 9648 -9801 9665 -9790
rect 9887 -9790 9984 -9776
rect 9887 -9801 9903 -9790
rect 9648 -9854 9903 -9801
rect 9967 -9801 9984 -9790
rect 10207 -9792 10304 -9778
rect 10207 -9801 10223 -9792
rect 9967 -9854 10223 -9801
rect 8200 -9856 10223 -9854
rect 10287 -9801 10304 -9792
rect 10527 -9792 10624 -9778
rect 10527 -9801 10543 -9792
rect 10287 -9856 10543 -9801
rect 10607 -9856 10624 -9792
rect 11274 -9836 11431 -8064
rect 8200 -9906 10624 -9856
rect 8200 -9965 9262 -9906
rect 9246 -9970 9262 -9965
rect 9326 -9965 9584 -9906
rect 9326 -9970 9343 -9965
rect 9246 -9988 9343 -9970
rect 9568 -9970 9584 -9965
rect 9648 -9965 9903 -9906
rect 9648 -9970 9665 -9965
rect 9568 -9988 9665 -9970
rect 9887 -9970 9903 -9965
rect 9967 -9908 10624 -9906
rect 9967 -9965 10223 -9908
rect 9967 -9970 9984 -9965
rect 9887 -9988 9984 -9970
rect 10207 -9972 10223 -9965
rect 10287 -9965 10543 -9908
rect 10287 -9972 10304 -9965
rect 10207 -9990 10304 -9972
rect 10527 -9972 10543 -9965
rect 10607 -9972 10624 -9908
rect 10527 -9990 10624 -9972
rect 11240 -9852 11454 -9836
rect 11240 -9916 11257 -9852
rect 11321 -9916 11377 -9852
rect 11441 -9916 11454 -9852
rect 11240 -9972 11454 -9916
rect 11240 -10036 11257 -9972
rect 11321 -10036 11377 -9972
rect 11441 -10036 11454 -9972
rect 11240 -10050 11454 -10036
rect 11274 -10226 11431 -10050
rect 9193 -10252 11431 -10226
rect 9193 -10255 10537 -10252
rect 9193 -10258 9586 -10255
rect 2514 -10280 2728 -10264
rect 2514 -10344 2531 -10280
rect 2595 -10344 2651 -10280
rect 2715 -10344 2728 -10280
rect 2514 -10400 2728 -10344
rect 9193 -10325 9258 -10258
rect 9323 -10322 9586 -10258
rect 9651 -10256 10537 -10255
rect 9651 -10322 9896 -10256
rect 9323 -10323 9896 -10322
rect 9961 -10323 10222 -10256
rect 10287 -10319 10537 -10256
rect 10602 -10319 11431 -10252
rect 10287 -10323 11431 -10319
rect 9323 -10325 11431 -10323
rect 9193 -10348 11431 -10325
rect 2514 -10464 2531 -10400
rect 2595 -10464 2651 -10400
rect 2715 -10464 2728 -10400
rect 2514 -10478 2728 -10464
rect 1994 -10546 2208 -10530
rect 1994 -10610 2011 -10546
rect 2075 -10610 2131 -10546
rect 2195 -10610 2208 -10546
rect 1994 -10666 2208 -10610
rect 1994 -10730 2011 -10666
rect 2075 -10730 2131 -10666
rect 2195 -10730 2208 -10666
rect 1994 -10744 2208 -10730
<< via2 >>
rect -242 -145 -160 -66
rect 621 -150 703 -71
rect 270 -1188 353 -1109
rect 1377 -1186 1461 -1108
rect -4042 -2591 -3919 -2471
rect -3842 -2591 -3719 -2471
rect -4039 -2843 -3916 -2723
rect -3839 -2843 -3716 -2723
rect -1734 -2810 -1654 -2730
rect -2142 -3021 -2086 -2965
rect -2032 -3021 -1976 -2965
rect -2533 -3329 -2477 -3273
rect -2423 -3329 -2367 -3273
rect -2844 -3629 -2762 -3549
rect -2510 -3875 -2454 -3819
rect -2400 -3875 -2344 -3819
rect -2107 -4187 -2051 -4131
rect -1997 -4187 -1941 -4131
rect 1583 -149 1666 -71
rect 3417 -3183 3481 -3119
rect 3537 -3183 3601 -3119
rect 3417 -3303 3481 -3239
rect 3537 -3303 3601 -3239
rect 2778 -3524 2842 -3460
rect 2898 -3524 2962 -3460
rect 2778 -3644 2842 -3580
rect 2898 -3644 2962 -3580
rect 6217 -3183 6281 -3119
rect 6337 -3183 6401 -3119
rect 6217 -3303 6281 -3239
rect 6337 -3303 6401 -3239
rect 3106 -3524 3170 -3460
rect 3226 -3524 3290 -3460
rect 3106 -3644 3170 -3580
rect 3226 -3644 3290 -3580
rect 3734 -3525 3798 -3461
rect 3854 -3525 3918 -3461
rect 3734 -3645 3798 -3581
rect 3854 -3645 3918 -3581
rect 4060 -3524 4124 -3460
rect 4180 -3524 4244 -3460
rect 4060 -3644 4124 -3580
rect 4180 -3644 4244 -3580
rect 5578 -3524 5642 -3460
rect 5698 -3524 5762 -3460
rect 5578 -3644 5642 -3580
rect 5698 -3644 5762 -3580
rect 7347 -3162 7411 -3098
rect 7467 -3162 7531 -3098
rect 7587 -3162 7651 -3098
rect 7707 -3162 7771 -3098
rect 7347 -3282 7411 -3218
rect 7467 -3282 7531 -3218
rect 7587 -3282 7651 -3218
rect 7707 -3282 7771 -3218
rect 5906 -3524 5970 -3460
rect 6026 -3524 6090 -3460
rect 5906 -3644 5970 -3580
rect 6026 -3644 6090 -3580
rect 6534 -3525 6598 -3461
rect 6654 -3525 6718 -3461
rect 6534 -3645 6598 -3581
rect 6654 -3645 6718 -3581
rect 6860 -3524 6924 -3460
rect 6980 -3524 7044 -3460
rect 6860 -3644 6924 -3580
rect 6980 -3644 7044 -3580
rect -1737 -4478 -1650 -4393
rect -2510 -4735 -2454 -4679
rect -2400 -4735 -2344 -4679
rect -2106 -5045 -2050 -4989
rect -1996 -5045 -1940 -4989
rect -2845 -5337 -2759 -5252
rect -2141 -5596 -2085 -5540
rect -2031 -5596 -1975 -5540
rect -2526 -5904 -2470 -5848
rect -2416 -5904 -2360 -5848
rect 353 -6024 435 -5939
rect -1731 -6156 -1651 -6076
rect -109 -6137 -27 -6052
rect 50 -6134 132 -6049
rect -2004 -6550 -1908 -6460
rect -2605 -6675 -2509 -6585
rect -2267 -6738 -2186 -6657
rect -411 -6733 -341 -6663
rect -169 -7129 -113 -7047
rect -2589 -7298 -2503 -7212
rect -170 -7314 -114 -7232
rect -1949 -7612 -1867 -7530
rect -2256 -7869 -2196 -7809
rect -1952 -8098 -1868 -8014
rect -2589 -8414 -2507 -8332
rect -2256 -8670 -2196 -8610
rect 2103 -6768 2174 -6755
rect 2239 -6768 2310 -6757
rect 2103 -6826 2127 -6768
rect 2127 -6826 2174 -6768
rect 2239 -6828 2241 -6768
rect 2241 -6828 2301 -6768
rect 2301 -6828 2310 -6768
rect 4958 -6494 5022 -6430
rect 5078 -6494 5142 -6430
rect 4958 -6614 5022 -6550
rect 5078 -6614 5142 -6550
rect 5531 -6497 5595 -6433
rect 5651 -6497 5715 -6433
rect 5531 -6617 5595 -6553
rect 5651 -6617 5715 -6553
rect 309 -7743 375 -7677
rect -177 -8004 -107 -7934
rect -175 -8144 -105 -8074
rect -409 -8365 -339 -8295
rect 9017 -3183 9081 -3119
rect 9137 -3183 9201 -3119
rect 9017 -3303 9081 -3239
rect 9137 -3303 9201 -3239
rect 11088 -1335 11169 -1254
rect 11228 -1335 11309 -1254
rect 11368 -1335 11449 -1254
rect 11508 -1335 11589 -1254
rect 11648 -1335 11729 -1254
rect 11094 -2764 11175 -2683
rect 11234 -2764 11315 -2683
rect 11374 -2764 11455 -2683
rect 11514 -2764 11595 -2683
rect 11654 -2764 11735 -2683
rect 8378 -3524 8442 -3460
rect 8498 -3524 8562 -3460
rect 8706 -3524 8770 -3460
rect 8826 -3524 8890 -3460
rect 9334 -3525 9398 -3461
rect 9454 -3525 9518 -3461
rect 9660 -3524 9724 -3460
rect 9780 -3524 9844 -3460
rect 8378 -3644 8442 -3580
rect 8498 -3644 8562 -3580
rect 8706 -3644 8770 -3580
rect 8826 -3644 8890 -3580
rect 9334 -3645 9398 -3581
rect 9454 -3645 9518 -3581
rect 9660 -3644 9724 -3580
rect 9780 -3644 9844 -3580
rect 11272 -5012 11336 -4948
rect 11392 -5012 11456 -4948
rect 11272 -5132 11336 -5068
rect 11392 -5132 11456 -5068
rect 6746 -6458 6810 -6394
rect 6866 -6458 6930 -6394
rect 6746 -6578 6810 -6514
rect 6866 -6578 6930 -6514
rect 7347 -6461 7411 -6397
rect 7467 -6461 7531 -6397
rect 7587 -6461 7651 -6397
rect 7707 -6461 7771 -6397
rect 7347 -6581 7411 -6517
rect 7467 -6581 7531 -6517
rect 7587 -6581 7651 -6517
rect 7707 -6581 7771 -6517
rect 904 -8654 970 -8588
rect 11262 -7618 11326 -7554
rect 11382 -7618 11446 -7554
rect 11262 -7738 11326 -7674
rect 11382 -7738 11446 -7674
rect -1952 -8902 -1866 -8816
rect -175 -9011 -105 -8941
rect -2591 -9215 -2509 -9133
rect -173 -9163 -103 -9093
rect -2257 -9470 -2197 -9410
rect 300 -9572 366 -9506
rect -2591 -9702 -2505 -9616
rect -412 -9904 -342 -9834
rect -1947 -10013 -1865 -9931
rect -169 -10054 -113 -9998
rect -169 -10168 -113 -10112
rect 11257 -9916 11321 -9852
rect 11377 -9916 11441 -9852
rect 11257 -10036 11321 -9972
rect 11377 -10036 11441 -9972
rect 2531 -10344 2595 -10280
rect 2651 -10344 2715 -10280
rect 2531 -10464 2595 -10400
rect 2651 -10464 2715 -10400
rect 2011 -10610 2075 -10546
rect 2131 -10610 2195 -10546
rect 2011 -10730 2075 -10666
rect 2131 -10730 2195 -10666
<< metal3 >>
rect -300 -66 1710 -20
rect -300 -145 -242 -66
rect -160 -71 1710 -66
rect -160 -145 621 -71
rect -300 -150 621 -145
rect 703 -149 1583 -71
rect 1666 -149 1710 -71
rect 703 -150 1710 -149
rect -300 -200 1710 -150
rect 240 -1108 1500 -1050
rect 240 -1109 1377 -1108
rect 240 -1188 270 -1109
rect 353 -1186 1377 -1109
rect 1461 -1186 1500 -1108
rect 353 -1188 1500 -1186
rect 240 -1230 1500 -1188
rect 11070 -1254 11746 -1239
rect 11070 -1335 11088 -1254
rect 11169 -1335 11228 -1254
rect 11309 -1335 11368 -1254
rect 11449 -1335 11508 -1254
rect 11589 -1335 11648 -1254
rect 11729 -1335 11746 -1254
rect 11070 -1349 11746 -1335
rect -4059 -2464 -3700 -2447
rect -4059 -2471 -1621 -2464
rect -4059 -2591 -4042 -2471
rect -3919 -2591 -3842 -2471
rect -3719 -2591 -1621 -2471
rect -4059 -2593 -1621 -2591
rect -4059 -2608 -3700 -2593
rect -4063 -2710 -3687 -2693
rect -4063 -2723 -2730 -2710
rect -4063 -2843 -4039 -2723
rect -3916 -2843 -3839 -2723
rect -3716 -2840 -2730 -2723
rect -3716 -2843 -3687 -2840
rect -4063 -2868 -3687 -2843
rect -2860 -3549 -2730 -2840
rect -1750 -2730 -1621 -2593
rect -1750 -2810 -1734 -2730
rect -1654 -2810 -1621 -2730
rect -2156 -2965 -1964 -2952
rect -2156 -3021 -2142 -2965
rect -2086 -3021 -2032 -2965
rect -1976 -3021 -1964 -2965
rect -2156 -3036 -1964 -3021
rect -2547 -3273 -2355 -3260
rect -2547 -3329 -2533 -3273
rect -2477 -3329 -2423 -3273
rect -2367 -3329 -2355 -3273
rect -2547 -3344 -2355 -3329
rect -2860 -3629 -2844 -3549
rect -2762 -3629 -2730 -3549
rect -2860 -5234 -2730 -3629
rect -2505 -3806 -2375 -3344
rect -2524 -3819 -2332 -3806
rect -2524 -3875 -2510 -3819
rect -2454 -3875 -2400 -3819
rect -2344 -3875 -2332 -3819
rect -2524 -3890 -2332 -3875
rect -2505 -4666 -2375 -3890
rect -2123 -4118 -1993 -3036
rect -2123 -4131 -1929 -4118
rect -2123 -4187 -2107 -4131
rect -2051 -4187 -1997 -4131
rect -1941 -4187 -1929 -4131
rect -2123 -4202 -1929 -4187
rect -2524 -4679 -2332 -4666
rect -2524 -4735 -2510 -4679
rect -2454 -4735 -2400 -4679
rect -2344 -4735 -2332 -4679
rect -2524 -4750 -2332 -4735
rect -2861 -5252 -2730 -5234
rect -2861 -5337 -2845 -5252
rect -2759 -5337 -2730 -5252
rect -2861 -5352 -2730 -5337
rect -2860 -6191 -2730 -5352
rect -2505 -5835 -2375 -4750
rect -2123 -4976 -1993 -4202
rect -1750 -4376 -1621 -2810
rect 10928 -2683 11892 -2628
rect 10928 -2764 11094 -2683
rect 11175 -2764 11234 -2683
rect 11315 -2764 11374 -2683
rect 11455 -2764 11514 -2683
rect 11595 -2764 11654 -2683
rect 11735 -2764 11892 -2683
rect 10928 -2953 11892 -2764
rect 3357 -3098 9263 -3036
rect 3357 -3119 7347 -3098
rect 3357 -3183 3417 -3119
rect 3481 -3183 3537 -3119
rect 3601 -3183 6217 -3119
rect 6281 -3183 6337 -3119
rect 6401 -3162 7347 -3119
rect 7411 -3162 7467 -3098
rect 7531 -3162 7587 -3098
rect 7651 -3162 7707 -3098
rect 7771 -3119 9263 -3098
rect 7771 -3162 9017 -3119
rect 6401 -3183 9017 -3162
rect 9081 -3183 9137 -3119
rect 9201 -3183 9263 -3119
rect 3357 -3218 9263 -3183
rect 3357 -3239 7347 -3218
rect 3357 -3303 3417 -3239
rect 3481 -3303 3537 -3239
rect 3601 -3303 6217 -3239
rect 6281 -3303 6337 -3239
rect 6401 -3282 7347 -3239
rect 7411 -3282 7467 -3218
rect 7531 -3282 7587 -3218
rect 7651 -3282 7707 -3218
rect 7771 -3239 9263 -3218
rect 7771 -3282 9017 -3239
rect 6401 -3303 9017 -3282
rect 9081 -3303 9137 -3239
rect 9201 -3303 9263 -3239
rect 3357 -3324 9263 -3303
rect 11157 -3443 11482 -2953
rect 2602 -3460 11482 -3443
rect 2602 -3524 2778 -3460
rect 2842 -3524 2898 -3460
rect 2962 -3524 3106 -3460
rect 3170 -3524 3226 -3460
rect 3290 -3461 4060 -3460
rect 3290 -3524 3734 -3461
rect 2602 -3525 3734 -3524
rect 3798 -3525 3854 -3461
rect 3918 -3524 4060 -3461
rect 4124 -3524 4180 -3460
rect 4244 -3524 5578 -3460
rect 5642 -3524 5698 -3460
rect 5762 -3524 5906 -3460
rect 5970 -3524 6026 -3460
rect 6090 -3461 6860 -3460
rect 6090 -3524 6534 -3461
rect 3918 -3525 6534 -3524
rect 6598 -3525 6654 -3461
rect 6718 -3524 6860 -3461
rect 6924 -3524 6980 -3460
rect 7044 -3524 8378 -3460
rect 8442 -3524 8498 -3460
rect 8562 -3524 8706 -3460
rect 8770 -3524 8826 -3460
rect 8890 -3461 9660 -3460
rect 8890 -3524 9334 -3461
rect 6718 -3525 9334 -3524
rect 9398 -3525 9454 -3461
rect 9518 -3524 9660 -3461
rect 9724 -3524 9780 -3460
rect 9844 -3524 11482 -3460
rect 9518 -3525 11482 -3524
rect 2602 -3580 11482 -3525
rect 2602 -3644 2778 -3580
rect 2842 -3644 2898 -3580
rect 2962 -3644 3106 -3580
rect 3170 -3644 3226 -3580
rect 3290 -3581 4060 -3580
rect 3290 -3644 3734 -3581
rect 2602 -3645 3734 -3644
rect 3798 -3645 3854 -3581
rect 3918 -3644 4060 -3581
rect 4124 -3644 4180 -3580
rect 4244 -3644 5578 -3580
rect 5642 -3644 5698 -3580
rect 5762 -3644 5906 -3580
rect 5970 -3644 6026 -3580
rect 6090 -3581 6860 -3580
rect 6090 -3644 6534 -3581
rect 3918 -3645 6534 -3644
rect 6598 -3645 6654 -3581
rect 6718 -3644 6860 -3581
rect 6924 -3644 6980 -3580
rect 7044 -3644 8378 -3580
rect 8442 -3644 8498 -3580
rect 8562 -3644 8706 -3580
rect 8770 -3644 8826 -3580
rect 8890 -3581 9660 -3580
rect 8890 -3644 9334 -3581
rect 6718 -3645 9334 -3644
rect 9398 -3645 9454 -3581
rect 9518 -3644 9660 -3581
rect 9724 -3644 9780 -3580
rect 9844 -3644 11482 -3580
rect 9518 -3645 11482 -3644
rect 2602 -3768 11482 -3645
rect -1756 -4393 -1621 -4376
rect -1756 -4478 -1737 -4393
rect -1650 -4478 -1621 -4393
rect -1756 -4491 -1621 -4478
rect -2123 -4989 -1928 -4976
rect -2123 -5045 -2106 -4989
rect -2050 -5045 -1996 -4989
rect -1940 -5045 -1928 -4989
rect -2123 -5060 -1928 -5045
rect -2123 -5527 -1993 -5060
rect -2155 -5540 -1963 -5527
rect -2155 -5596 -2141 -5540
rect -2085 -5596 -2031 -5540
rect -1975 -5596 -1963 -5540
rect -2155 -5611 -1963 -5596
rect -2540 -5848 -2348 -5835
rect -2540 -5904 -2526 -5848
rect -2470 -5904 -2416 -5848
rect -2360 -5904 -2348 -5848
rect -2540 -5919 -2348 -5904
rect -2505 -6444 -2375 -5919
rect -2631 -6566 -2375 -6444
rect -2123 -6423 -1993 -5611
rect -1750 -6076 -1621 -4491
rect 11241 -4948 11481 -4917
rect 9246 -5046 9336 -4955
rect 9560 -5045 9650 -4954
rect 9877 -5042 9967 -4951
rect 10208 -5041 10298 -4950
rect 10527 -5042 10617 -4951
rect 11241 -5012 11272 -4948
rect 11336 -5012 11392 -4948
rect 11456 -5012 11481 -4948
rect 11241 -5068 11481 -5012
rect 11241 -5132 11272 -5068
rect 11336 -5132 11392 -5068
rect 11456 -5132 11481 -5068
rect -1750 -6156 -1731 -6076
rect -1651 -6156 -1621 -6076
rect -1750 -6179 -1621 -6156
rect -449 -5939 460 -5809
rect -2123 -6456 -1880 -6423
rect -2123 -6460 -1840 -6456
rect -2123 -6550 -2004 -6460
rect -1908 -6550 -1840 -6460
rect -2123 -6553 -1840 -6550
rect -2631 -6585 -2481 -6566
rect -2030 -6579 -1840 -6553
rect -2631 -6675 -2605 -6585
rect -2509 -6675 -2481 -6585
rect -2631 -7212 -2481 -6675
rect -2631 -7298 -2589 -7212
rect -2503 -7298 -2481 -7212
rect -2631 -8332 -2481 -7298
rect -2631 -8414 -2589 -8332
rect -2507 -8414 -2481 -8332
rect -2631 -9133 -2481 -8414
rect -2631 -9215 -2591 -9133
rect -2509 -9215 -2481 -9133
rect -2631 -9505 -2481 -9215
rect -2635 -9616 -2481 -9505
rect -2298 -6657 -2136 -6635
rect -2298 -6738 -2267 -6657
rect -2186 -6738 -2136 -6657
rect -2298 -7809 -2136 -6738
rect -2298 -7869 -2256 -7809
rect -2196 -7869 -2136 -7809
rect -2298 -8610 -2136 -7869
rect -2298 -8670 -2256 -8610
rect -2196 -8670 -2136 -8610
rect -2298 -9410 -2136 -8670
rect -2298 -9470 -2257 -9410
rect -2197 -9470 -2136 -9410
rect -2298 -9507 -2136 -9470
rect -1977 -7530 -1840 -6579
rect -1977 -7612 -1949 -7530
rect -1867 -7612 -1840 -7530
rect -1977 -8014 -1840 -7612
rect -1977 -8098 -1952 -8014
rect -1868 -8098 -1840 -8014
rect -1977 -8816 -1840 -8098
rect -1977 -8902 -1952 -8816
rect -1866 -8902 -1840 -8816
rect -2635 -9702 -2591 -9616
rect -2505 -9702 -2481 -9616
rect -2635 -10535 -2481 -9702
rect -1977 -9931 -1840 -8902
rect -449 -6663 -319 -5939
rect 327 -6024 353 -5939
rect 435 -6024 460 -5939
rect -146 -6033 148 -6030
rect -449 -6733 -411 -6663
rect -341 -6733 -319 -6663
rect -449 -8295 -319 -6733
rect -449 -8365 -409 -8295
rect -339 -8365 -319 -8295
rect -449 -9834 -319 -8365
rect -449 -9904 -412 -9834
rect -342 -9904 -319 -9834
rect -449 -9924 -319 -9904
rect -195 -6049 148 -6033
rect 327 -6040 460 -6024
rect -195 -6052 50 -6049
rect -195 -6137 -109 -6052
rect -27 -6134 50 -6052
rect 132 -6134 148 -6049
rect 11241 -6087 11481 -5132
rect -27 -6137 148 -6134
rect -195 -6161 148 -6137
rect 11228 -6123 11519 -6087
rect -195 -7047 -67 -6161
rect 11228 -6204 11263 -6123
rect 11344 -6204 11413 -6123
rect 11494 -6204 11519 -6123
rect 11228 -6273 11519 -6204
rect 4914 -6394 7982 -6277
rect 4914 -6430 6746 -6394
rect 4914 -6494 4958 -6430
rect 5022 -6494 5078 -6430
rect 5142 -6433 6746 -6430
rect 5142 -6494 5531 -6433
rect 4914 -6497 5531 -6494
rect 5595 -6497 5651 -6433
rect 5715 -6458 6746 -6433
rect 6810 -6458 6866 -6394
rect 6930 -6397 7982 -6394
rect 6930 -6458 7347 -6397
rect 5715 -6461 7347 -6458
rect 7411 -6461 7467 -6397
rect 7531 -6461 7587 -6397
rect 7651 -6461 7707 -6397
rect 7771 -6461 7982 -6397
rect 5715 -6497 7982 -6461
rect 4914 -6514 7982 -6497
rect 4914 -6550 6746 -6514
rect 4914 -6614 4958 -6550
rect 5022 -6614 5078 -6550
rect 5142 -6553 6746 -6550
rect 5142 -6614 5531 -6553
rect 4914 -6617 5531 -6614
rect 5595 -6617 5651 -6553
rect 5715 -6578 6746 -6553
rect 6810 -6578 6866 -6514
rect 6930 -6517 7982 -6514
rect 6930 -6578 7347 -6517
rect 5715 -6581 7347 -6578
rect 7411 -6581 7467 -6517
rect 7531 -6581 7587 -6517
rect 7651 -6581 7707 -6517
rect 7771 -6581 7982 -6517
rect 5715 -6617 7982 -6581
rect 4914 -6696 7982 -6617
rect 11228 -6354 11263 -6273
rect 11344 -6354 11413 -6273
rect 11494 -6354 11519 -6273
rect 11228 -6418 11519 -6354
rect 11228 -6499 11267 -6418
rect 11348 -6499 11417 -6418
rect 11498 -6499 11519 -6418
rect 11228 -6568 11519 -6499
rect 11228 -6649 11267 -6568
rect 11348 -6649 11417 -6568
rect 11498 -6649 11519 -6568
rect 11228 -6685 11519 -6649
rect 2076 -6755 2332 -6723
rect 2076 -6826 2103 -6755
rect 2174 -6757 2332 -6755
rect 2174 -6826 2239 -6757
rect 2076 -6828 2239 -6826
rect 2310 -6828 2332 -6757
rect 2076 -6841 2332 -6828
rect -195 -7129 -169 -7047
rect -113 -7129 -67 -7047
rect -195 -7232 -67 -7129
rect -195 -7314 -170 -7232
rect -114 -7314 -67 -7232
rect -195 -7934 -67 -7314
rect 2087 -7571 2301 -6841
rect 9245 -7337 9335 -7246
rect 9573 -7334 9663 -7243
rect 9883 -7335 9973 -7244
rect 10209 -7335 10299 -7244
rect 10524 -7331 10614 -7240
rect 286 -7677 2301 -7571
rect 286 -7743 309 -7677
rect 375 -7743 2301 -7677
rect 286 -7785 2301 -7743
rect 11241 -7554 11481 -6685
rect 11241 -7618 11262 -7554
rect 11326 -7618 11382 -7554
rect 11446 -7618 11481 -7554
rect 11241 -7674 11481 -7618
rect 11241 -7738 11262 -7674
rect 11326 -7738 11382 -7674
rect 11446 -7738 11481 -7674
rect -195 -8004 -177 -7934
rect -107 -8004 -67 -7934
rect -195 -8074 -67 -8004
rect -195 -8144 -175 -8074
rect -105 -8144 -67 -8074
rect -195 -8941 -67 -8144
rect -195 -9011 -175 -8941
rect -105 -9011 -67 -8941
rect -195 -9093 -67 -9011
rect -195 -9163 -173 -9093
rect -103 -9163 -67 -9093
rect -195 -9816 -67 -9163
rect 855 -8588 1035 -7785
rect 9246 -8046 9336 -7955
rect 9560 -8045 9650 -7954
rect 9877 -8042 9967 -7951
rect 10208 -8041 10298 -7950
rect 10527 -8042 10617 -7951
rect 855 -8654 904 -8588
rect 970 -8654 1035 -8588
rect 855 -9468 1035 -8654
rect 11241 -8770 11481 -7738
rect 11222 -8806 11513 -8770
rect 11222 -8887 11257 -8806
rect 11338 -8887 11407 -8806
rect 11488 -8887 11513 -8806
rect 11222 -8956 11513 -8887
rect 11222 -9037 11257 -8956
rect 11338 -9037 11407 -8956
rect 11488 -9037 11513 -8956
rect 11222 -9101 11513 -9037
rect 11222 -9182 11261 -9101
rect 11342 -9182 11411 -9101
rect 11492 -9182 11513 -9101
rect 11222 -9251 11513 -9182
rect 11222 -9332 11261 -9251
rect 11342 -9332 11411 -9251
rect 11492 -9332 11513 -9251
rect 11222 -9368 11513 -9332
rect 251 -9506 1035 -9468
rect 251 -9572 300 -9506
rect 366 -9572 1035 -9506
rect 251 -9614 1035 -9572
rect 11241 -9816 11481 -9368
rect -195 -9852 11481 -9816
rect -195 -9916 11257 -9852
rect 11321 -9916 11377 -9852
rect 11441 -9916 11481 -9852
rect -1977 -10013 -1947 -9931
rect -1865 -10013 -1840 -9931
rect -1977 -10289 -1840 -10013
rect -195 -9972 11481 -9916
rect -195 -9998 11257 -9972
rect -195 -10054 -169 -9998
rect -113 -10036 11257 -9998
rect 11321 -10036 11377 -9972
rect 11441 -10036 11481 -9972
rect -113 -10054 11481 -10036
rect -195 -10056 11481 -10054
rect -195 -10112 -67 -10056
rect -195 -10136 -169 -10112
rect -184 -10168 -169 -10136
rect -113 -10136 -67 -10112
rect -113 -10168 -99 -10136
rect -184 -10184 -99 -10168
rect 2514 -10280 2728 -10264
rect 2514 -10289 2531 -10280
rect -1977 -10344 2531 -10289
rect 2595 -10344 2651 -10280
rect 2715 -10344 2728 -10280
rect 9245 -10337 9335 -10246
rect 9573 -10334 9663 -10243
rect 9883 -10335 9973 -10244
rect 10209 -10335 10299 -10244
rect 10524 -10331 10614 -10240
rect -1977 -10400 2728 -10344
rect -1977 -10448 2531 -10400
rect 2514 -10464 2531 -10448
rect 2595 -10464 2651 -10400
rect 2715 -10464 2728 -10400
rect 2514 -10478 2728 -10464
rect 1994 -10535 2208 -10530
rect -2635 -10546 2208 -10535
rect -2635 -10610 2011 -10546
rect 2075 -10610 2131 -10546
rect 2195 -10610 2208 -10546
rect -2635 -10666 2208 -10610
rect -2635 -10691 2011 -10666
rect 1994 -10730 2011 -10691
rect 2075 -10730 2131 -10666
rect 2195 -10730 2208 -10666
rect 1994 -10744 2208 -10730
<< via3 >>
rect 11088 -1335 11169 -1254
rect 11228 -1335 11309 -1254
rect 11368 -1335 11449 -1254
rect 11508 -1335 11589 -1254
rect 11648 -1335 11729 -1254
rect 11263 -6204 11344 -6123
rect 11413 -6204 11494 -6123
rect 11263 -6354 11344 -6273
rect 11413 -6354 11494 -6273
rect 11267 -6499 11348 -6418
rect 11417 -6499 11498 -6418
rect 11267 -6649 11348 -6568
rect 11417 -6649 11498 -6568
rect 11257 -8887 11338 -8806
rect 11407 -8887 11488 -8806
rect 11257 -9037 11338 -8956
rect 11407 -9037 11488 -8956
rect 11261 -9182 11342 -9101
rect 11411 -9182 11492 -9101
rect 11261 -9332 11342 -9251
rect 11411 -9332 11492 -9251
<< metal4 >>
rect 11070 -1254 11746 -1239
rect 11070 -1335 11088 -1254
rect 11169 -1335 11228 -1254
rect 11309 -1335 11368 -1254
rect 11449 -1335 11508 -1254
rect 11589 -1335 11648 -1254
rect 11729 -1335 11746 -1254
rect 11070 -1349 11746 -1335
rect 11228 -6123 11519 -6087
rect 11228 -6204 11263 -6123
rect 11344 -6204 11413 -6123
rect 11494 -6204 11519 -6123
rect 11228 -6273 11519 -6204
rect 11228 -6354 11263 -6273
rect 11344 -6354 11413 -6273
rect 11494 -6354 11519 -6273
rect 11228 -6418 11519 -6354
rect 11228 -6499 11267 -6418
rect 11348 -6499 11417 -6418
rect 11498 -6499 11519 -6418
rect 11228 -6568 11519 -6499
rect 11228 -6649 11267 -6568
rect 11348 -6649 11417 -6568
rect 11498 -6649 11519 -6568
rect 11228 -6685 11519 -6649
rect 11222 -8806 11513 -8770
rect 11222 -8887 11257 -8806
rect 11338 -8887 11407 -8806
rect 11488 -8887 11513 -8806
rect 11222 -8956 11513 -8887
rect 11222 -9037 11257 -8956
rect 11338 -9037 11407 -8956
rect 11488 -9037 11513 -8956
rect 11222 -9101 11513 -9037
rect 11222 -9182 11261 -9101
rect 11342 -9182 11411 -9101
rect 11492 -9182 11513 -9101
rect 11222 -9251 11513 -9182
rect 11222 -9332 11261 -9251
rect 11342 -9332 11411 -9251
rect 11492 -9332 11513 -9251
rect 11222 -9368 11513 -9332
<< via4 >>
rect 11088 -1335 11169 -1254
rect 11228 -1335 11309 -1254
rect 11368 -1335 11449 -1254
rect 11508 -1335 11589 -1254
rect 11648 -1335 11729 -1254
rect 11263 -6204 11344 -6123
rect 11413 -6204 11494 -6123
rect 11263 -6354 11344 -6273
rect 11413 -6354 11494 -6273
rect 11267 -6499 11348 -6418
rect 11417 -6499 11498 -6418
rect 11267 -6649 11348 -6568
rect 11417 -6649 11498 -6568
rect 11257 -8887 11338 -8806
rect 11407 -8887 11488 -8806
rect 11257 -9037 11338 -8956
rect 11407 -9037 11488 -8956
rect 11261 -9182 11342 -9101
rect 11411 -9182 11492 -9101
rect 11261 -9332 11342 -9251
rect 11411 -9332 11492 -9251
<< metal5 >>
rect 10970 -1254 12660 -1183
rect 10970 -1335 11088 -1254
rect 11169 -1335 11228 -1254
rect 11309 -1335 11368 -1254
rect 11449 -1335 11508 -1254
rect 11589 -1335 11648 -1254
rect 11729 -1335 12660 -1254
rect 10970 -1456 12660 -1335
rect 12387 -4068 12660 -1456
rect 12387 -4341 14684 -4068
rect 11228 -6123 11519 -6087
rect 11228 -6204 11263 -6123
rect 11344 -6204 11413 -6123
rect 11494 -6156 11519 -6123
rect 11494 -6204 12002 -6156
rect 11228 -6273 12002 -6204
rect 11228 -6354 11263 -6273
rect 11344 -6354 11413 -6273
rect 11494 -6354 12002 -6273
rect 11228 -6418 12002 -6354
rect 11228 -6499 11267 -6418
rect 11348 -6499 11417 -6418
rect 11498 -6499 12002 -6418
rect 11228 -6568 12002 -6499
rect 11228 -6649 11267 -6568
rect 11348 -6649 11417 -6568
rect 11498 -6640 12002 -6568
rect 11498 -6649 11519 -6640
rect 11228 -6685 11519 -6649
rect 11222 -8806 11513 -8770
rect 11222 -8887 11257 -8806
rect 11338 -8887 11407 -8806
rect 11488 -8873 11513 -8806
rect 11488 -8887 11989 -8873
rect 11222 -8956 11989 -8887
rect 11222 -9037 11257 -8956
rect 11338 -9037 11407 -8956
rect 11488 -9037 11989 -8956
rect 11222 -9101 11989 -9037
rect 11222 -9182 11261 -9101
rect 11342 -9182 11411 -9101
rect 11492 -9182 11989 -9101
rect 11222 -9251 11989 -9182
rect 11222 -9332 11261 -9251
rect 11342 -9332 11411 -9251
rect 11492 -9332 11989 -9251
rect 11222 -9357 11989 -9332
rect 11222 -9368 11513 -9357
use cap_mim_2p0fF_XHV85N  cap_mim_2p0fF_XHV85N_0
timestamp 1694159936
transform -1 0 14432 0 -1 -7788
box -2640 -3460 2640 3460
use nmos_3p3_4F3WC4  nmos_3p3_4F3WC4_0
timestamp 1693997255
transform 1 0 5473 0 1 -7846
box -516 -804 516 804
use nmos_3p3_4F3WC4  nmos_3p3_4F3WC4_1
timestamp 1693997255
transform 1 0 6993 0 1 -7846
box -516 -804 516 804
use nmos_3p3_5F3WC4  nmos_3p3_5F3WC4_0
timestamp 1693997255
transform 1 0 6233 0 1 -7846
box -364 -804 364 804
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_0
timestamp 1692712407
transform 1 0 -2546 0 -1 -9037
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_1
timestamp 1692712407
transform 1 0 -2546 0 -1 -9837
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_2
timestamp 1692712407
transform -1 0 -1906 0 -1 -9037
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_3
timestamp 1692712407
transform -1 0 -1906 0 -1 -9837
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_4
timestamp 1692712407
transform 1 0 -2546 0 1 -8239
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_5
timestamp 1692712407
transform -1 0 -1906 0 1 -8239
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_6
timestamp 1692712407
transform 1 0 -2546 0 1 -7439
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_7
timestamp 1692712407
transform -1 0 -1906 0 1 -7439
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_8
timestamp 1692712407
transform 1 0 340 0 1 -9962
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_9
timestamp 1692712407
transform 1 0 340 0 1 -9112
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_10
timestamp 1692712407
transform 1 0 340 0 1 -8132
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_11
timestamp 1692712407
transform 1 0 340 0 1 -7282
box -220 -368 220 368
use nmos_3p3_676RTJ  nmos_3p3_676RTJ_0
timestamp 1693916241
transform 1 0 2303 0 1 -8789
box -540 -368 540 368
use nmos_3p3_676RTJ  nmos_3p3_676RTJ_1
timestamp 1693916241
transform 1 0 2296 0 -1 -9915
box -540 -368 540 368
use nmos_3p3_M56RTJ  nmos_3p3_M56RTJ_0
timestamp 1694074718
transform 1 0 10815 0 1 -9146
box -140 -1104 140 1104
use nmos_3p3_M56RTJ  nmos_3p3_M56RTJ_1
timestamp 1694074718
transform 1 0 9055 0 1 -6146
box -140 -1104 140 1104
use nmos_3p3_M56RTJ  nmos_3p3_M56RTJ_2
timestamp 1694074718
transform 1 0 10815 0 1 -6146
box -140 -1104 140 1104
use nmos_3p3_M56RTJ  nmos_3p3_M56RTJ_3
timestamp 1694074718
transform 1 0 9055 0 1 -9146
box -140 -1104 140 1104
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_0
timestamp 1692712407
transform 1 0 -2946 0 -1 -9037
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_1
timestamp 1692712407
transform 1 0 -2306 0 -1 -9037
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_2
timestamp 1692712407
transform 1 0 -2786 0 -1 -9037
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_3
timestamp 1692712407
transform 1 0 -2306 0 -1 -9837
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_4
timestamp 1692712407
transform 1 0 -2946 0 -1 -9837
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_5
timestamp 1692712407
transform 1 0 -2786 0 -1 -9837
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_6
timestamp 1692712407
transform -1 0 -2146 0 -1 -9037
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_7
timestamp 1692712407
transform -1 0 -1666 0 -1 -9037
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_8
timestamp 1692712407
transform -1 0 -1506 0 -1 -9037
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_9
timestamp 1692712407
transform -1 0 -2146 0 -1 -9837
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_10
timestamp 1692712407
transform -1 0 -1506 0 -1 -9837
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_11
timestamp 1692712407
transform -1 0 -1666 0 -1 -9837
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_12
timestamp 1692712407
transform 1 0 -2306 0 1 -8239
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_13
timestamp 1692712407
transform 1 0 -2786 0 1 -8239
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_14
timestamp 1692712407
transform 1 0 -2946 0 1 -8239
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_15
timestamp 1692712407
transform -1 0 -1506 0 1 -8239
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_16
timestamp 1692712407
transform -1 0 -1666 0 1 -8239
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_17
timestamp 1692712407
transform -1 0 -2146 0 1 -8239
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_18
timestamp 1692712407
transform 1 0 -2306 0 1 -7439
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_19
timestamp 1692712407
transform 1 0 -2946 0 1 -7439
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_20
timestamp 1692712407
transform 1 0 -2786 0 1 -7439
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_21
timestamp 1692712407
transform -1 0 -2146 0 1 -7439
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_22
timestamp 1692712407
transform -1 0 -1666 0 1 -7439
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_23
timestamp 1692712407
transform -1 0 -1506 0 1 -7439
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_24
timestamp 1692712407
transform -1 0 741 0 1 -9962
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_25
timestamp 1692712407
transform -1 0 901 0 1 -9962
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_26
timestamp 1692712407
transform -1 0 -221 0 1 -9962
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_27
timestamp 1692712407
transform -1 0 -61 0 1 -9962
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_28
timestamp 1692712407
transform -1 0 901 0 1 -9112
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_29
timestamp 1692712407
transform -1 0 741 0 1 -9112
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_30
timestamp 1692712407
transform -1 0 -221 0 1 -9112
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_31
timestamp 1692712407
transform -1 0 -61 0 1 -9112
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_32
timestamp 1692712407
transform -1 0 -61 0 1 -8132
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_33
timestamp 1692712407
transform -1 0 -221 0 1 -8132
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_34
timestamp 1692712407
transform -1 0 901 0 1 -8132
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_35
timestamp 1692712407
transform -1 0 741 0 1 -8132
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_36
timestamp 1692712407
transform -1 0 -221 0 1 -7282
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_37
timestamp 1692712407
transform -1 0 -61 0 1 -7282
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_38
timestamp 1692712407
transform -1 0 901 0 1 -7282
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_39
timestamp 1692712407
transform -1 0 741 0 1 -7282
box -140 -368 140 368
use nmos_3p3_N3WVC4  nmos_3p3_N3WVC4_0
timestamp 1693997255
transform 1 0 4727 0 1 -7846
box -212 -804 212 804
use nmos_3p3_N3WVC4  nmos_3p3_N3WVC4_1
timestamp 1693997255
transform 1 0 7735 0 1 -7846
box -212 -804 212 804
use nmos_3p3_NQ5EG7  nmos_3p3_NQ5EG7_0
timestamp 1694074718
transform 1 0 9935 0 1 -6146
box -860 -1104 860 1104
use nmos_3p3_NQ5EG7  nmos_3p3_NQ5EG7_1
timestamp 1694074718
transform 1 0 9935 0 1 -9146
box -860 -1104 860 1104
use nmos_3p3_QNHHV5  nmos_3p3_QNHHV5_0
timestamp 1693997255
transform 1 0 2318 0 1 -7121
box -168 -268 168 268
use nmos_3p3_QNHHV5  nmos_3p3_QNHHV5_1
timestamp 1693997255
transform 1 0 1886 0 1 -7121
box -168 -268 168 268
use nmos_3p3_QNHHV5  nmos_3p3_QNHHV5_2
timestamp 1693997255
transform 1 0 2102 0 1 -7121
box -168 -268 168 268
use nmos_3p3_QNHHV5  nmos_3p3_QNHHV5_3
timestamp 1693997255
transform 1 0 3442 0 1 -7121
box -168 -268 168 268
use nmos_3p3_QNHHV5  nmos_3p3_QNHHV5_4
timestamp 1693997255
transform 1 0 2534 0 1 -7121
box -168 -268 168 268
use nmos_3p3_QNHHV5  nmos_3p3_QNHHV5_5
timestamp 1693997255
transform 1 0 2880 0 1 -7121
box -168 -268 168 268
use nmos_3p3_QNHHV5  nmos_3p3_QNHHV5_6
timestamp 1693997255
transform 1 0 3226 0 1 -7121
box -168 -268 168 268
use nmos_3p3_QNHHV5  nmos_3p3_QNHHV5_8
timestamp 1693997255
transform 1 0 3791 0 1 -7121
box -168 -268 168 268
use pmos_3p3_9BLZD7  pmos_3p3_9BLZD7_0
timestamp 1692615943
transform 1 0 -2299 0 1 -255
box -554 -1534 554 1534
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_0
timestamp 1692615943
transform 1 0 771 0 1 -1664
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_1
timestamp 1692615943
transform 1 0 -309 0 1 -2702
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_2
timestamp 1692615943
transform 1 0 -93 0 1 -2702
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_3
timestamp 1692615943
transform 1 0 555 0 1 -1664
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_4
timestamp 1692615943
transform 1 0 771 0 1 -2702
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_5
timestamp 1692615943
transform 1 0 555 0 1 -2702
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_6
timestamp 1692615943
transform 1 0 -309 0 1 -1664
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_7
timestamp 1692615943
transform 1 0 -93 0 1 -1664
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_8
timestamp 1692615943
transform 1 0 771 0 1 -624
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_9
timestamp 1692615943
transform 1 0 555 0 1 -624
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_10
timestamp 1692615943
transform 1 0 555 0 1 414
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_11
timestamp 1692615943
transform 1 0 771 0 1 414
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_12
timestamp 1692615943
transform 1 0 -93 0 1 -624
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_13
timestamp 1692615943
transform 1 0 -309 0 1 -624
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_14
timestamp 1692615943
transform 1 0 -309 0 1 414
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_15
timestamp 1692615943
transform 1 0 -93 0 1 414
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_16
timestamp 1692615943
transform 1 0 -2839 0 1 -1359
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_17
timestamp 1692615943
transform 1 0 -1759 0 1 -1359
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_18
timestamp 1692615943
transform 1 0 -2839 0 1 113
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_19
timestamp 1692615943
transform 1 0 -2839 0 1 -623
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_20
timestamp 1692615943
transform 1 0 -2839 0 1 849
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_21
timestamp 1692615943
transform 1 0 -1759 0 1 849
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_22
timestamp 1692615943
transform 1 0 -1759 0 1 113
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_23
timestamp 1692615943
transform 1 0 -1759 0 1 -623
box -230 -430 230 430
use pmos_3p3_H6V2RY  pmos_3p3_H6V2RY_0
timestamp 1694004920
transform 1 0 4839 0 1 -5235
box -426 -598 426 598
use pmos_3p3_H6V2RY  pmos_3p3_H6V2RY_1
timestamp 1694004920
transform 1 0 5889 0 1 -5235
box -426 -598 426 598
use pmos_3p3_HWZ2RY  pmos_3p3_HWZ2RY_0
timestamp 1694004920
transform 1 0 4383 0 1 -5235
box -274 -598 274 598
use pmos_3p3_HWZ2RY  pmos_3p3_HWZ2RY_1
timestamp 1694004920
transform 1 0 6345 0 1 -5235
box -274 -598 274 598
use pmos_3p3_HWZ2RY  pmos_3p3_HWZ2RY_2
timestamp 1694004920
transform 1 0 5295 0 1 -5235
box -274 -598 274 598
use pmos_3p3_M2JNAR  pmos_3p3_M2JNAR_0
timestamp 1693911244
transform 1 0 6315 0 1 -923
box -282 -1902 282 1902
use pmos_3p3_M2JNAR  pmos_3p3_M2JNAR_1
timestamp 1693911244
transform 1 0 9115 0 1 -923
box -282 -1902 282 1902
use pmos_3p3_M2JNAR  pmos_3p3_M2JNAR_2
timestamp 1693911244
transform 1 0 3515 0 1 -923
box -282 -1902 282 1902
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_0
timestamp 1692683681
transform 1 0 395 0 1 -5568
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_1
timestamp 1692683681
transform 1 0 395 0 1 -4788
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_2
timestamp 1692683681
transform -1 0 -1925 0 -1 -4869
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_3
timestamp 1692683681
transform -1 0 -1925 0 -1 -5721
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_4
timestamp 1692683681
transform 1 0 -2565 0 -1 -4869
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_5
timestamp 1692683681
transform 1 0 -2565 0 -1 -5721
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_6
timestamp 1692683681
transform 1 0 -2565 0 1 -4017
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_7
timestamp 1692683681
transform -1 0 -1925 0 1 -4017
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_8
timestamp 1692683681
transform 1 0 -2565 0 1 -3165
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_9
timestamp 1692683681
transform -1 0 -1925 0 1 -3165
box -282 -430 282 430
use pmos_3p3_M22VUP  pmos_3p3_M22VUP_0
timestamp 1691491496
transform 1 0 231 0 1 -1664
box -338 -430 338 430
use pmos_3p3_M22VUP  pmos_3p3_M22VUP_1
timestamp 1691491496
transform 1 0 231 0 1 -2702
box -338 -430 338 430
use pmos_3p3_M22VUP  pmos_3p3_M22VUP_2
timestamp 1691491496
transform 1 0 231 0 1 -624
box -338 -430 338 430
use pmos_3p3_M22VUP  pmos_3p3_M22VUP_3
timestamp 1691491496
transform 1 0 231 0 1 414
box -338 -430 338 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_0
timestamp 1692683681
transform 1 0 27 0 1 -5568
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_1
timestamp 1692683681
transform 1 0 -133 0 1 -5568
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_2
timestamp 1692683681
transform 1 0 923 0 1 -5568
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_3
timestamp 1692683681
transform 1 0 763 0 1 -5568
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_4
timestamp 1692683681
transform 1 0 -133 0 1 -4788
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_5
timestamp 1692683681
transform 1 0 27 0 1 -4788
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_6
timestamp 1692683681
transform 1 0 923 0 1 -4788
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_7
timestamp 1692683681
transform 1 0 763 0 1 -4788
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_8
timestamp 1692683681
transform -1 0 -1525 0 -1 -4869
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_9
timestamp 1692683681
transform -1 0 -1685 0 -1 -4869
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_10
timestamp 1692683681
transform -1 0 -2165 0 -1 -4869
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_11
timestamp 1692683681
transform -1 0 -1685 0 -1 -5721
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_12
timestamp 1692683681
transform -1 0 -1525 0 -1 -5721
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_13
timestamp 1692683681
transform -1 0 -2165 0 -1 -5721
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_14
timestamp 1692683681
transform 1 0 -2805 0 1 -4017
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_15
timestamp 1692683681
transform 1 0 -2965 0 1 -4017
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_16
timestamp 1692683681
transform 1 0 -2805 0 -1 -4869
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_17
timestamp 1692683681
transform 1 0 -2965 0 -1 -4869
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_18
timestamp 1692683681
transform 1 0 -2325 0 -1 -4869
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_19
timestamp 1692683681
transform -1 0 -2165 0 1 -4017
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_20
timestamp 1692683681
transform 1 0 -2805 0 -1 -5721
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_21
timestamp 1692683681
transform 1 0 -2965 0 -1 -5721
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_22
timestamp 1692683681
transform 1 0 -2325 0 -1 -5721
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_23
timestamp 1692683681
transform 1 0 -2325 0 1 -4017
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_24
timestamp 1692683681
transform 1 0 -2805 0 1 -3165
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_25
timestamp 1692683681
transform 1 0 -2965 0 1 -3165
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_26
timestamp 1692683681
transform -1 0 -2165 0 1 -3165
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_27
timestamp 1692683681
transform -1 0 -1685 0 1 -4017
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_28
timestamp 1692683681
transform -1 0 -1525 0 1 -4017
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_29
timestamp 1692683681
transform -1 0 -1525 0 1 -3165
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_30
timestamp 1692683681
transform -1 0 -1685 0 1 -3165
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_31
timestamp 1692683681
transform 1 0 -2325 0 1 -3165
box -202 -430 202 430
use pmos_3p3_MAJNAR  pmos_3p3_MAJNAR_0
timestamp 1693911244
transform 1 0 5435 0 1 -923
box -202 -1902 202 1902
use pmos_3p3_MAJNAR  pmos_3p3_MAJNAR_1
timestamp 1693911244
transform 1 0 7195 0 1 -923
box -202 -1902 202 1902
use pmos_3p3_MAJNAR  pmos_3p3_MAJNAR_2
timestamp 1693911244
transform 1 0 8235 0 1 -923
box -202 -1902 202 1902
use pmos_3p3_MAJNAR  pmos_3p3_MAJNAR_3
timestamp 1693911244
transform 1 0 9995 0 1 -923
box -202 -1902 202 1902
use pmos_3p3_MAJNAR  pmos_3p3_MAJNAR_4
timestamp 1693911244
transform 1 0 4395 0 1 -923
box -202 -1902 202 1902
use pmos_3p3_MAJNAR  pmos_3p3_MAJNAR_5
timestamp 1693911244
transform 1 0 2635 0 1 -923
box -202 -1902 202 1902
use pmos_3p3_MJGNAR  pmos_3p3_MJGNAR_0
timestamp 1693911244
transform 1 0 5835 0 1 -923
box -442 -1902 442 1902
use pmos_3p3_MJGNAR  pmos_3p3_MJGNAR_1
timestamp 1693911244
transform 1 0 6795 0 1 -923
box -442 -1902 442 1902
use pmos_3p3_MJGNAR  pmos_3p3_MJGNAR_2
timestamp 1693911244
transform 1 0 8635 0 1 -923
box -442 -1902 442 1902
use pmos_3p3_MJGNAR  pmos_3p3_MJGNAR_3
timestamp 1693911244
transform 1 0 9595 0 1 -923
box -442 -1902 442 1902
use pmos_3p3_MJGNAR  pmos_3p3_MJGNAR_4
timestamp 1693911244
transform 1 0 3995 0 1 -923
box -442 -1902 442 1902
use pmos_3p3_MJGNAR  pmos_3p3_MJGNAR_5
timestamp 1693911244
transform 1 0 3035 0 1 -923
box -442 -1902 442 1902
use pmos_3p3_VK6RD7  pmos_3p3_VK6RD7_0
timestamp 1693470477
transform 1 0 1916 0 1 -4934
box -230 -330 230 330
use pmos_3p3_VK6RD7  pmos_3p3_VK6RD7_1
timestamp 1693470477
transform 1 0 3342 0 1 -5642
box -230 -330 230 330
use pmos_3p3_VK6RD7  pmos_3p3_VK6RD7_2
timestamp 1693470477
transform 1 0 2564 0 1 -5642
box -230 -330 230 330
use pmos_3p3_VK6RD7  pmos_3p3_VK6RD7_3
timestamp 1693470477
transform 1 0 2780 0 1 -5642
box -230 -330 230 330
use pmos_3p3_VK6RD7  pmos_3p3_VK6RD7_4
timestamp 1693470477
transform 1 0 3126 0 1 -5642
box -230 -330 230 330
use pmos_3p3_VK6RD7  pmos_3p3_VK6RD7_5
timestamp 1693470477
transform 1 0 2218 0 1 -5642
box -230 -330 230 330
use pmos_3p3_VK6RD7  pmos_3p3_VK6RD7_6
timestamp 1693470477
transform 1 0 2002 0 1 -5642
box -230 -330 230 330
use pmos_3p3_VK6RD7  pmos_3p3_VK6RD7_7
timestamp 1693470477
transform 1 0 3428 0 1 -4934
box -230 -330 230 330
use pmos_3p3_VTYQD7  pmos_3p3_VTYQD7_0
timestamp 1693470477
transform 1 0 2240 0 1 -4934
box -338 -330 338 330
use pmos_3p3_VTYQD7  pmos_3p3_VTYQD7_1
timestamp 1693470477
transform 1 0 3104 0 1 -4934
box -338 -330 338 330
use pmos_3p3_VTYQD7  pmos_3p3_VTYQD7_2
timestamp 1693470477
transform 1 0 2672 0 1 -4934
box -338 -330 338 330
use ppolyf_u_WRMTN3  ppolyf_u_WRMTN3_0
timestamp 1694159936
transform 1 0 11437 0 1 -2013
box -864 -932 864 932
<< labels >>
flabel metal1 672 -6091 672 -6091 0 FreeSans 640 0 0 0 OUT
port 7 nsew
flabel via2 -3767 -2533 -3767 -2533 0 FreeSans 480 0 0 0 VINN
port 3 nsew
flabel metal3 -2619 -6615 -2619 -6615 0 FreeSans 1600 0 0 0 VC
port 11 nsew
flabel metal3 -2024 -6512 -2024 -6512 0 FreeSans 1600 0 0 0 VD
port 13 nsew
flabel metal1 276 -5980 276 -5980 0 FreeSans 960 0 0 0 VX
port 15 nsew
flabel metal2 -74 -4260 -74 -4260 0 FreeSans 960 0 0 0 VBS2
port 20 nsew
flabel via2 -3963 -2776 -3963 -2776 0 FreeSans 480 0 0 0 VINP
port 2 nsew
flabel metal3 2214 -6861 2214 -6861 0 FreeSans 960 0 0 0 VBS3
port 22 nsew
flabel metal1 2990 -6842 2990 -6842 0 FreeSans 960 0 0 0 VBIASN
port 24 nsew
flabel metal1 21 -3616 21 -3616 0 FreeSans 960 0 0 0 VA
port 16 nsew
flabel metal1 991 -3795 991 -3795 0 FreeSans 960 0 0 0 VB
port 18 nsew
flabel metal1 3371 -10582 3371 -10582 0 FreeSans 1600 0 0 0 VSS
port 1 nsew
flabel metal1 5365 -4651 5365 -4651 0 FreeSans 960 0 0 0 IBIAS2
port 26 nsew
flabel metal1 6234 -8706 6234 -8706 0 FreeSans 960 0 0 0 VBIASN2
port 28 nsew
flabel metal2 5019 -7015 5019 -7015 0 FreeSans 960 0 0 0 IBIAS3
port 30 nsew
flabel metal1 -2185 1254 -2185 1254 0 FreeSans 960 0 0 0 IBIAS
port 32 nsew
flabel metal3 9104 -3600 9104 -3600 0 FreeSans 960 0 0 0 OUTo
port 34 nsew
flabel metal2 -3378 -2243 -3378 -2241 0 FreeSans 960 0 0 0 VP
port 36 nsew
flabel metal1 221 1353 221 1353 0 FreeSans 1600 0 0 0 VDD
port 0 nsew
flabel metal5 11203 -1294 11203 -1294 0 FreeSans 800 0 0 0 c_mid
port 38 nsew
<< end >>
