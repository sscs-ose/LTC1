magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1880 -1319 1880 1319
<< metal4 >>
rect -877 311 877 316
rect -877 283 -872 311
rect -844 283 -806 311
rect -778 283 -740 311
rect -712 283 -674 311
rect -646 283 -608 311
rect -580 283 -542 311
rect -514 283 -476 311
rect -448 283 -410 311
rect -382 283 -344 311
rect -316 283 -278 311
rect -250 283 -212 311
rect -184 283 -146 311
rect -118 283 -80 311
rect -52 283 -14 311
rect 14 283 52 311
rect 80 283 118 311
rect 146 283 184 311
rect 212 283 250 311
rect 278 283 316 311
rect 344 283 382 311
rect 410 283 448 311
rect 476 283 514 311
rect 542 283 580 311
rect 608 283 646 311
rect 674 283 712 311
rect 740 283 778 311
rect 806 283 844 311
rect 872 283 877 311
rect -877 245 877 283
rect -877 217 -872 245
rect -844 217 -806 245
rect -778 217 -740 245
rect -712 217 -674 245
rect -646 217 -608 245
rect -580 217 -542 245
rect -514 217 -476 245
rect -448 217 -410 245
rect -382 217 -344 245
rect -316 217 -278 245
rect -250 217 -212 245
rect -184 217 -146 245
rect -118 217 -80 245
rect -52 217 -14 245
rect 14 217 52 245
rect 80 217 118 245
rect 146 217 184 245
rect 212 217 250 245
rect 278 217 316 245
rect 344 217 382 245
rect 410 217 448 245
rect 476 217 514 245
rect 542 217 580 245
rect 608 217 646 245
rect 674 217 712 245
rect 740 217 778 245
rect 806 217 844 245
rect 872 217 877 245
rect -877 179 877 217
rect -877 151 -872 179
rect -844 151 -806 179
rect -778 151 -740 179
rect -712 151 -674 179
rect -646 151 -608 179
rect -580 151 -542 179
rect -514 151 -476 179
rect -448 151 -410 179
rect -382 151 -344 179
rect -316 151 -278 179
rect -250 151 -212 179
rect -184 151 -146 179
rect -118 151 -80 179
rect -52 151 -14 179
rect 14 151 52 179
rect 80 151 118 179
rect 146 151 184 179
rect 212 151 250 179
rect 278 151 316 179
rect 344 151 382 179
rect 410 151 448 179
rect 476 151 514 179
rect 542 151 580 179
rect 608 151 646 179
rect 674 151 712 179
rect 740 151 778 179
rect 806 151 844 179
rect 872 151 877 179
rect -877 113 877 151
rect -877 85 -872 113
rect -844 85 -806 113
rect -778 85 -740 113
rect -712 85 -674 113
rect -646 85 -608 113
rect -580 85 -542 113
rect -514 85 -476 113
rect -448 85 -410 113
rect -382 85 -344 113
rect -316 85 -278 113
rect -250 85 -212 113
rect -184 85 -146 113
rect -118 85 -80 113
rect -52 85 -14 113
rect 14 85 52 113
rect 80 85 118 113
rect 146 85 184 113
rect 212 85 250 113
rect 278 85 316 113
rect 344 85 382 113
rect 410 85 448 113
rect 476 85 514 113
rect 542 85 580 113
rect 608 85 646 113
rect 674 85 712 113
rect 740 85 778 113
rect 806 85 844 113
rect 872 85 877 113
rect -877 47 877 85
rect -877 19 -872 47
rect -844 19 -806 47
rect -778 19 -740 47
rect -712 19 -674 47
rect -646 19 -608 47
rect -580 19 -542 47
rect -514 19 -476 47
rect -448 19 -410 47
rect -382 19 -344 47
rect -316 19 -278 47
rect -250 19 -212 47
rect -184 19 -146 47
rect -118 19 -80 47
rect -52 19 -14 47
rect 14 19 52 47
rect 80 19 118 47
rect 146 19 184 47
rect 212 19 250 47
rect 278 19 316 47
rect 344 19 382 47
rect 410 19 448 47
rect 476 19 514 47
rect 542 19 580 47
rect 608 19 646 47
rect 674 19 712 47
rect 740 19 778 47
rect 806 19 844 47
rect 872 19 877 47
rect -877 -19 877 19
rect -877 -47 -872 -19
rect -844 -47 -806 -19
rect -778 -47 -740 -19
rect -712 -47 -674 -19
rect -646 -47 -608 -19
rect -580 -47 -542 -19
rect -514 -47 -476 -19
rect -448 -47 -410 -19
rect -382 -47 -344 -19
rect -316 -47 -278 -19
rect -250 -47 -212 -19
rect -184 -47 -146 -19
rect -118 -47 -80 -19
rect -52 -47 -14 -19
rect 14 -47 52 -19
rect 80 -47 118 -19
rect 146 -47 184 -19
rect 212 -47 250 -19
rect 278 -47 316 -19
rect 344 -47 382 -19
rect 410 -47 448 -19
rect 476 -47 514 -19
rect 542 -47 580 -19
rect 608 -47 646 -19
rect 674 -47 712 -19
rect 740 -47 778 -19
rect 806 -47 844 -19
rect 872 -47 877 -19
rect -877 -85 877 -47
rect -877 -113 -872 -85
rect -844 -113 -806 -85
rect -778 -113 -740 -85
rect -712 -113 -674 -85
rect -646 -113 -608 -85
rect -580 -113 -542 -85
rect -514 -113 -476 -85
rect -448 -113 -410 -85
rect -382 -113 -344 -85
rect -316 -113 -278 -85
rect -250 -113 -212 -85
rect -184 -113 -146 -85
rect -118 -113 -80 -85
rect -52 -113 -14 -85
rect 14 -113 52 -85
rect 80 -113 118 -85
rect 146 -113 184 -85
rect 212 -113 250 -85
rect 278 -113 316 -85
rect 344 -113 382 -85
rect 410 -113 448 -85
rect 476 -113 514 -85
rect 542 -113 580 -85
rect 608 -113 646 -85
rect 674 -113 712 -85
rect 740 -113 778 -85
rect 806 -113 844 -85
rect 872 -113 877 -85
rect -877 -151 877 -113
rect -877 -179 -872 -151
rect -844 -179 -806 -151
rect -778 -179 -740 -151
rect -712 -179 -674 -151
rect -646 -179 -608 -151
rect -580 -179 -542 -151
rect -514 -179 -476 -151
rect -448 -179 -410 -151
rect -382 -179 -344 -151
rect -316 -179 -278 -151
rect -250 -179 -212 -151
rect -184 -179 -146 -151
rect -118 -179 -80 -151
rect -52 -179 -14 -151
rect 14 -179 52 -151
rect 80 -179 118 -151
rect 146 -179 184 -151
rect 212 -179 250 -151
rect 278 -179 316 -151
rect 344 -179 382 -151
rect 410 -179 448 -151
rect 476 -179 514 -151
rect 542 -179 580 -151
rect 608 -179 646 -151
rect 674 -179 712 -151
rect 740 -179 778 -151
rect 806 -179 844 -151
rect 872 -179 877 -151
rect -877 -217 877 -179
rect -877 -245 -872 -217
rect -844 -245 -806 -217
rect -778 -245 -740 -217
rect -712 -245 -674 -217
rect -646 -245 -608 -217
rect -580 -245 -542 -217
rect -514 -245 -476 -217
rect -448 -245 -410 -217
rect -382 -245 -344 -217
rect -316 -245 -278 -217
rect -250 -245 -212 -217
rect -184 -245 -146 -217
rect -118 -245 -80 -217
rect -52 -245 -14 -217
rect 14 -245 52 -217
rect 80 -245 118 -217
rect 146 -245 184 -217
rect 212 -245 250 -217
rect 278 -245 316 -217
rect 344 -245 382 -217
rect 410 -245 448 -217
rect 476 -245 514 -217
rect 542 -245 580 -217
rect 608 -245 646 -217
rect 674 -245 712 -217
rect 740 -245 778 -217
rect 806 -245 844 -217
rect 872 -245 877 -217
rect -877 -283 877 -245
rect -877 -311 -872 -283
rect -844 -311 -806 -283
rect -778 -311 -740 -283
rect -712 -311 -674 -283
rect -646 -311 -608 -283
rect -580 -311 -542 -283
rect -514 -311 -476 -283
rect -448 -311 -410 -283
rect -382 -311 -344 -283
rect -316 -311 -278 -283
rect -250 -311 -212 -283
rect -184 -311 -146 -283
rect -118 -311 -80 -283
rect -52 -311 -14 -283
rect 14 -311 52 -283
rect 80 -311 118 -283
rect 146 -311 184 -283
rect 212 -311 250 -283
rect 278 -311 316 -283
rect 344 -311 382 -283
rect 410 -311 448 -283
rect 476 -311 514 -283
rect 542 -311 580 -283
rect 608 -311 646 -283
rect 674 -311 712 -283
rect 740 -311 778 -283
rect 806 -311 844 -283
rect 872 -311 877 -283
rect -877 -316 877 -311
<< via4 >>
rect -872 283 -844 311
rect -806 283 -778 311
rect -740 283 -712 311
rect -674 283 -646 311
rect -608 283 -580 311
rect -542 283 -514 311
rect -476 283 -448 311
rect -410 283 -382 311
rect -344 283 -316 311
rect -278 283 -250 311
rect -212 283 -184 311
rect -146 283 -118 311
rect -80 283 -52 311
rect -14 283 14 311
rect 52 283 80 311
rect 118 283 146 311
rect 184 283 212 311
rect 250 283 278 311
rect 316 283 344 311
rect 382 283 410 311
rect 448 283 476 311
rect 514 283 542 311
rect 580 283 608 311
rect 646 283 674 311
rect 712 283 740 311
rect 778 283 806 311
rect 844 283 872 311
rect -872 217 -844 245
rect -806 217 -778 245
rect -740 217 -712 245
rect -674 217 -646 245
rect -608 217 -580 245
rect -542 217 -514 245
rect -476 217 -448 245
rect -410 217 -382 245
rect -344 217 -316 245
rect -278 217 -250 245
rect -212 217 -184 245
rect -146 217 -118 245
rect -80 217 -52 245
rect -14 217 14 245
rect 52 217 80 245
rect 118 217 146 245
rect 184 217 212 245
rect 250 217 278 245
rect 316 217 344 245
rect 382 217 410 245
rect 448 217 476 245
rect 514 217 542 245
rect 580 217 608 245
rect 646 217 674 245
rect 712 217 740 245
rect 778 217 806 245
rect 844 217 872 245
rect -872 151 -844 179
rect -806 151 -778 179
rect -740 151 -712 179
rect -674 151 -646 179
rect -608 151 -580 179
rect -542 151 -514 179
rect -476 151 -448 179
rect -410 151 -382 179
rect -344 151 -316 179
rect -278 151 -250 179
rect -212 151 -184 179
rect -146 151 -118 179
rect -80 151 -52 179
rect -14 151 14 179
rect 52 151 80 179
rect 118 151 146 179
rect 184 151 212 179
rect 250 151 278 179
rect 316 151 344 179
rect 382 151 410 179
rect 448 151 476 179
rect 514 151 542 179
rect 580 151 608 179
rect 646 151 674 179
rect 712 151 740 179
rect 778 151 806 179
rect 844 151 872 179
rect -872 85 -844 113
rect -806 85 -778 113
rect -740 85 -712 113
rect -674 85 -646 113
rect -608 85 -580 113
rect -542 85 -514 113
rect -476 85 -448 113
rect -410 85 -382 113
rect -344 85 -316 113
rect -278 85 -250 113
rect -212 85 -184 113
rect -146 85 -118 113
rect -80 85 -52 113
rect -14 85 14 113
rect 52 85 80 113
rect 118 85 146 113
rect 184 85 212 113
rect 250 85 278 113
rect 316 85 344 113
rect 382 85 410 113
rect 448 85 476 113
rect 514 85 542 113
rect 580 85 608 113
rect 646 85 674 113
rect 712 85 740 113
rect 778 85 806 113
rect 844 85 872 113
rect -872 19 -844 47
rect -806 19 -778 47
rect -740 19 -712 47
rect -674 19 -646 47
rect -608 19 -580 47
rect -542 19 -514 47
rect -476 19 -448 47
rect -410 19 -382 47
rect -344 19 -316 47
rect -278 19 -250 47
rect -212 19 -184 47
rect -146 19 -118 47
rect -80 19 -52 47
rect -14 19 14 47
rect 52 19 80 47
rect 118 19 146 47
rect 184 19 212 47
rect 250 19 278 47
rect 316 19 344 47
rect 382 19 410 47
rect 448 19 476 47
rect 514 19 542 47
rect 580 19 608 47
rect 646 19 674 47
rect 712 19 740 47
rect 778 19 806 47
rect 844 19 872 47
rect -872 -47 -844 -19
rect -806 -47 -778 -19
rect -740 -47 -712 -19
rect -674 -47 -646 -19
rect -608 -47 -580 -19
rect -542 -47 -514 -19
rect -476 -47 -448 -19
rect -410 -47 -382 -19
rect -344 -47 -316 -19
rect -278 -47 -250 -19
rect -212 -47 -184 -19
rect -146 -47 -118 -19
rect -80 -47 -52 -19
rect -14 -47 14 -19
rect 52 -47 80 -19
rect 118 -47 146 -19
rect 184 -47 212 -19
rect 250 -47 278 -19
rect 316 -47 344 -19
rect 382 -47 410 -19
rect 448 -47 476 -19
rect 514 -47 542 -19
rect 580 -47 608 -19
rect 646 -47 674 -19
rect 712 -47 740 -19
rect 778 -47 806 -19
rect 844 -47 872 -19
rect -872 -113 -844 -85
rect -806 -113 -778 -85
rect -740 -113 -712 -85
rect -674 -113 -646 -85
rect -608 -113 -580 -85
rect -542 -113 -514 -85
rect -476 -113 -448 -85
rect -410 -113 -382 -85
rect -344 -113 -316 -85
rect -278 -113 -250 -85
rect -212 -113 -184 -85
rect -146 -113 -118 -85
rect -80 -113 -52 -85
rect -14 -113 14 -85
rect 52 -113 80 -85
rect 118 -113 146 -85
rect 184 -113 212 -85
rect 250 -113 278 -85
rect 316 -113 344 -85
rect 382 -113 410 -85
rect 448 -113 476 -85
rect 514 -113 542 -85
rect 580 -113 608 -85
rect 646 -113 674 -85
rect 712 -113 740 -85
rect 778 -113 806 -85
rect 844 -113 872 -85
rect -872 -179 -844 -151
rect -806 -179 -778 -151
rect -740 -179 -712 -151
rect -674 -179 -646 -151
rect -608 -179 -580 -151
rect -542 -179 -514 -151
rect -476 -179 -448 -151
rect -410 -179 -382 -151
rect -344 -179 -316 -151
rect -278 -179 -250 -151
rect -212 -179 -184 -151
rect -146 -179 -118 -151
rect -80 -179 -52 -151
rect -14 -179 14 -151
rect 52 -179 80 -151
rect 118 -179 146 -151
rect 184 -179 212 -151
rect 250 -179 278 -151
rect 316 -179 344 -151
rect 382 -179 410 -151
rect 448 -179 476 -151
rect 514 -179 542 -151
rect 580 -179 608 -151
rect 646 -179 674 -151
rect 712 -179 740 -151
rect 778 -179 806 -151
rect 844 -179 872 -151
rect -872 -245 -844 -217
rect -806 -245 -778 -217
rect -740 -245 -712 -217
rect -674 -245 -646 -217
rect -608 -245 -580 -217
rect -542 -245 -514 -217
rect -476 -245 -448 -217
rect -410 -245 -382 -217
rect -344 -245 -316 -217
rect -278 -245 -250 -217
rect -212 -245 -184 -217
rect -146 -245 -118 -217
rect -80 -245 -52 -217
rect -14 -245 14 -217
rect 52 -245 80 -217
rect 118 -245 146 -217
rect 184 -245 212 -217
rect 250 -245 278 -217
rect 316 -245 344 -217
rect 382 -245 410 -217
rect 448 -245 476 -217
rect 514 -245 542 -217
rect 580 -245 608 -217
rect 646 -245 674 -217
rect 712 -245 740 -217
rect 778 -245 806 -217
rect 844 -245 872 -217
rect -872 -311 -844 -283
rect -806 -311 -778 -283
rect -740 -311 -712 -283
rect -674 -311 -646 -283
rect -608 -311 -580 -283
rect -542 -311 -514 -283
rect -476 -311 -448 -283
rect -410 -311 -382 -283
rect -344 -311 -316 -283
rect -278 -311 -250 -283
rect -212 -311 -184 -283
rect -146 -311 -118 -283
rect -80 -311 -52 -283
rect -14 -311 14 -283
rect 52 -311 80 -283
rect 118 -311 146 -283
rect 184 -311 212 -283
rect 250 -311 278 -283
rect 316 -311 344 -283
rect 382 -311 410 -283
rect 448 -311 476 -283
rect 514 -311 542 -283
rect 580 -311 608 -283
rect 646 -311 674 -283
rect 712 -311 740 -283
rect 778 -311 806 -283
rect 844 -311 872 -283
<< metal5 >>
rect -880 311 880 319
rect -880 283 -872 311
rect -844 283 -806 311
rect -778 283 -740 311
rect -712 283 -674 311
rect -646 283 -608 311
rect -580 283 -542 311
rect -514 283 -476 311
rect -448 283 -410 311
rect -382 283 -344 311
rect -316 283 -278 311
rect -250 283 -212 311
rect -184 283 -146 311
rect -118 283 -80 311
rect -52 283 -14 311
rect 14 283 52 311
rect 80 283 118 311
rect 146 283 184 311
rect 212 283 250 311
rect 278 283 316 311
rect 344 283 382 311
rect 410 283 448 311
rect 476 283 514 311
rect 542 283 580 311
rect 608 283 646 311
rect 674 283 712 311
rect 740 283 778 311
rect 806 283 844 311
rect 872 283 880 311
rect -880 245 880 283
rect -880 217 -872 245
rect -844 217 -806 245
rect -778 217 -740 245
rect -712 217 -674 245
rect -646 217 -608 245
rect -580 217 -542 245
rect -514 217 -476 245
rect -448 217 -410 245
rect -382 217 -344 245
rect -316 217 -278 245
rect -250 217 -212 245
rect -184 217 -146 245
rect -118 217 -80 245
rect -52 217 -14 245
rect 14 217 52 245
rect 80 217 118 245
rect 146 217 184 245
rect 212 217 250 245
rect 278 217 316 245
rect 344 217 382 245
rect 410 217 448 245
rect 476 217 514 245
rect 542 217 580 245
rect 608 217 646 245
rect 674 217 712 245
rect 740 217 778 245
rect 806 217 844 245
rect 872 217 880 245
rect -880 179 880 217
rect -880 151 -872 179
rect -844 151 -806 179
rect -778 151 -740 179
rect -712 151 -674 179
rect -646 151 -608 179
rect -580 151 -542 179
rect -514 151 -476 179
rect -448 151 -410 179
rect -382 151 -344 179
rect -316 151 -278 179
rect -250 151 -212 179
rect -184 151 -146 179
rect -118 151 -80 179
rect -52 151 -14 179
rect 14 151 52 179
rect 80 151 118 179
rect 146 151 184 179
rect 212 151 250 179
rect 278 151 316 179
rect 344 151 382 179
rect 410 151 448 179
rect 476 151 514 179
rect 542 151 580 179
rect 608 151 646 179
rect 674 151 712 179
rect 740 151 778 179
rect 806 151 844 179
rect 872 151 880 179
rect -880 113 880 151
rect -880 85 -872 113
rect -844 85 -806 113
rect -778 85 -740 113
rect -712 85 -674 113
rect -646 85 -608 113
rect -580 85 -542 113
rect -514 85 -476 113
rect -448 85 -410 113
rect -382 85 -344 113
rect -316 85 -278 113
rect -250 85 -212 113
rect -184 85 -146 113
rect -118 85 -80 113
rect -52 85 -14 113
rect 14 85 52 113
rect 80 85 118 113
rect 146 85 184 113
rect 212 85 250 113
rect 278 85 316 113
rect 344 85 382 113
rect 410 85 448 113
rect 476 85 514 113
rect 542 85 580 113
rect 608 85 646 113
rect 674 85 712 113
rect 740 85 778 113
rect 806 85 844 113
rect 872 85 880 113
rect -880 47 880 85
rect -880 19 -872 47
rect -844 19 -806 47
rect -778 19 -740 47
rect -712 19 -674 47
rect -646 19 -608 47
rect -580 19 -542 47
rect -514 19 -476 47
rect -448 19 -410 47
rect -382 19 -344 47
rect -316 19 -278 47
rect -250 19 -212 47
rect -184 19 -146 47
rect -118 19 -80 47
rect -52 19 -14 47
rect 14 19 52 47
rect 80 19 118 47
rect 146 19 184 47
rect 212 19 250 47
rect 278 19 316 47
rect 344 19 382 47
rect 410 19 448 47
rect 476 19 514 47
rect 542 19 580 47
rect 608 19 646 47
rect 674 19 712 47
rect 740 19 778 47
rect 806 19 844 47
rect 872 19 880 47
rect -880 -19 880 19
rect -880 -47 -872 -19
rect -844 -47 -806 -19
rect -778 -47 -740 -19
rect -712 -47 -674 -19
rect -646 -47 -608 -19
rect -580 -47 -542 -19
rect -514 -47 -476 -19
rect -448 -47 -410 -19
rect -382 -47 -344 -19
rect -316 -47 -278 -19
rect -250 -47 -212 -19
rect -184 -47 -146 -19
rect -118 -47 -80 -19
rect -52 -47 -14 -19
rect 14 -47 52 -19
rect 80 -47 118 -19
rect 146 -47 184 -19
rect 212 -47 250 -19
rect 278 -47 316 -19
rect 344 -47 382 -19
rect 410 -47 448 -19
rect 476 -47 514 -19
rect 542 -47 580 -19
rect 608 -47 646 -19
rect 674 -47 712 -19
rect 740 -47 778 -19
rect 806 -47 844 -19
rect 872 -47 880 -19
rect -880 -85 880 -47
rect -880 -113 -872 -85
rect -844 -113 -806 -85
rect -778 -113 -740 -85
rect -712 -113 -674 -85
rect -646 -113 -608 -85
rect -580 -113 -542 -85
rect -514 -113 -476 -85
rect -448 -113 -410 -85
rect -382 -113 -344 -85
rect -316 -113 -278 -85
rect -250 -113 -212 -85
rect -184 -113 -146 -85
rect -118 -113 -80 -85
rect -52 -113 -14 -85
rect 14 -113 52 -85
rect 80 -113 118 -85
rect 146 -113 184 -85
rect 212 -113 250 -85
rect 278 -113 316 -85
rect 344 -113 382 -85
rect 410 -113 448 -85
rect 476 -113 514 -85
rect 542 -113 580 -85
rect 608 -113 646 -85
rect 674 -113 712 -85
rect 740 -113 778 -85
rect 806 -113 844 -85
rect 872 -113 880 -85
rect -880 -151 880 -113
rect -880 -179 -872 -151
rect -844 -179 -806 -151
rect -778 -179 -740 -151
rect -712 -179 -674 -151
rect -646 -179 -608 -151
rect -580 -179 -542 -151
rect -514 -179 -476 -151
rect -448 -179 -410 -151
rect -382 -179 -344 -151
rect -316 -179 -278 -151
rect -250 -179 -212 -151
rect -184 -179 -146 -151
rect -118 -179 -80 -151
rect -52 -179 -14 -151
rect 14 -179 52 -151
rect 80 -179 118 -151
rect 146 -179 184 -151
rect 212 -179 250 -151
rect 278 -179 316 -151
rect 344 -179 382 -151
rect 410 -179 448 -151
rect 476 -179 514 -151
rect 542 -179 580 -151
rect 608 -179 646 -151
rect 674 -179 712 -151
rect 740 -179 778 -151
rect 806 -179 844 -151
rect 872 -179 880 -151
rect -880 -217 880 -179
rect -880 -245 -872 -217
rect -844 -245 -806 -217
rect -778 -245 -740 -217
rect -712 -245 -674 -217
rect -646 -245 -608 -217
rect -580 -245 -542 -217
rect -514 -245 -476 -217
rect -448 -245 -410 -217
rect -382 -245 -344 -217
rect -316 -245 -278 -217
rect -250 -245 -212 -217
rect -184 -245 -146 -217
rect -118 -245 -80 -217
rect -52 -245 -14 -217
rect 14 -245 52 -217
rect 80 -245 118 -217
rect 146 -245 184 -217
rect 212 -245 250 -217
rect 278 -245 316 -217
rect 344 -245 382 -217
rect 410 -245 448 -217
rect 476 -245 514 -217
rect 542 -245 580 -217
rect 608 -245 646 -217
rect 674 -245 712 -217
rect 740 -245 778 -217
rect 806 -245 844 -217
rect 872 -245 880 -217
rect -880 -283 880 -245
rect -880 -311 -872 -283
rect -844 -311 -806 -283
rect -778 -311 -740 -283
rect -712 -311 -674 -283
rect -646 -311 -608 -283
rect -580 -311 -542 -283
rect -514 -311 -476 -283
rect -448 -311 -410 -283
rect -382 -311 -344 -283
rect -316 -311 -278 -283
rect -250 -311 -212 -283
rect -184 -311 -146 -283
rect -118 -311 -80 -283
rect -52 -311 -14 -283
rect 14 -311 52 -283
rect 80 -311 118 -283
rect 146 -311 184 -283
rect 212 -311 250 -283
rect 278 -311 316 -283
rect 344 -311 382 -283
rect 410 -311 448 -283
rect 476 -311 514 -283
rect 542 -311 580 -283
rect 608 -311 646 -283
rect 674 -311 712 -283
rect 740 -311 778 -283
rect 806 -311 844 -283
rect 872 -311 880 -283
rect -880 -319 880 -311
<< end >>
