magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -7445 -2195 7445 2195
<< psubdiff >>
rect -5445 173 5445 195
rect -5445 -173 -5423 173
rect 5423 -173 5445 173
rect -5445 -195 5445 -173
<< psubdiffcont >>
rect -5423 -173 5423 173
<< metal1 >>
rect -5434 173 5434 184
rect -5434 -173 -5423 173
rect 5423 -173 5434 173
rect -5434 -184 5434 -173
<< end >>
