* NGSPICE file created from TG_flat.ext - technology: gf180mcuC

.subckt TG_flat VSS SD0_1 G0_2 G0_1 VDD G1_2 G1_1 SD2_0 G3_2 G3_1
X0 G3_2 G3_2.t36 G3_1.t31 VSS.t106 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X1 G3_2 G3_2.t44 G3_1.t30 VSS.t105 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X2 G1_2 G1_2.t12 VDD.t127 VDD.t89 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X3 G3_2 G3_2.t32 G3_1.t29 VSS.t104 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X4 VDD G1_2.t97 SD2_0.t37 VDD.t6 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X5 SD2_0 G1_2.t98 VDD.t124 VDD.t59 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X6 SD0_1 G0_2.t0 G1_1.t95 VSS.t11 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X7 G1_2 G1_2.t14 VDD.t123 VDD.t87 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X8 SD2_0 G1_2.t100 VDD.t122 VDD.t73 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X9 G1_1 G0_2.t1 SD0_1.t30 VSS.t71 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X10 SD0_1 G0_2.t2 G1_1.t94 VSS.t14 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X11 VDD G1_2.t50 G1_2.t51 VDD.t66 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X12 SD2_0 G1_2.t101 VDD.t119 VDD.t52 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X13 G3_2 G3_2.t46 G3_1.t28 VSS.t103 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X14 G1_2 G1_1.t62 G1_1.t63 VDD.t0 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X15 G3_1 G3_2.t90 G3_2.t91 VSS.t102 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X16 VDD G1_2.t48 G1_2.t49 VDD.t61 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X17 VSS G0_1.t0 SD0_1.t42 VSS.t0 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X18 G1_2 G1_2.t8 VDD.t116 VDD.t10 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X19 VDD G1_2.t46 G1_2.t47 VDD.t9 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X20 VSS G3_1.t84 G3_1.t85 VSS.t105 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X21 G3_1 G3_1.t40 VSS.t152 VSS.t100 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X22 SD0_1 G0_1.t1 VSS.t39 VSS.t38 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X23 G1_1 G0_2.t3 SD0_1.t28 VSS.t25 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X24 G1_1 G1_1.t60 G1_2.t92 VDD.t1 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X25 SD2_0 G1_1.t97 G3_2.t6 VDD.t36 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X26 SD2_0 G1_1.t98 G3_2.t7 VDD.t43 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X27 VDD G1_2.t103 SD2_0.t33 VDD.t50 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X28 G1_1 G1_1.t58 G1_2.t91 VDD.t2 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X29 SD0_1 G0_1.t2 VSS.t41 VSS.t40 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X30 VSS G0_1.t3 SD0_1.t61 VSS.t3 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X31 G3_1 G3_1.t38 VSS.t151 VSS.t102 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X32 G3_2 G3_2.t40 G3_1.t26 VSS.t101 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X33 G1_2 G1_1.t56 G1_1.t57 VDD.t89 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X34 VSS G0_1.t4 SD0_1.t62 VSS.t74 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X35 SD0_1 G0_2.t4 G1_1.t93 VSS.t2 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X36 VDD G1_2.t44 G1_2.t45 VDD.t5 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X37 G3_1 G3_2.t88 G3_2.t89 VSS.t100 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X38 G3_2 G3_2.t58 G3_1.t24 VSS.t99 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X39 G1_2 G1_1.t54 G1_1.t55 VDD.t87 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X40 G1_1 G0_2.t5 SD0_1.t26 VSS.t22 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X41 G1_1 G0_2.t6 SD0_1.t25 VSS.t28 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X42 G3_2 G1_1.t100 SD2_0.t40 VDD.t25 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X43 SD0_1 G0_2.t7 G1_1.t92 VSS.t31 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X44 G3_2 G1_1.t101 SD2_0.t50 VDD.t15 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X45 VDD G1_2.t104 SD2_0.t32 VDD.t45 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X46 SD0_1 G0_1.t5 VSS.t159 VSS.t19 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X47 G3_2 G3_2.t48 G3_1.t23 VSS.t98 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X48 G3_2 G1_1.t102 SD2_0.t51 VDD.t29 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X49 VSS G0_1.t6 SD0_1.t32 VSS.t6 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X50 G3_2 G1_1.t103 SD2_0.t52 VDD.t17 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X51 G1_2 G1_2.t10 VDD.t107 VDD.t0 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X52 G1_2 G1_1.t52 G1_1.t53 VDD.t10 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X53 G3_1 G3_1.t36 VSS.t150 VSS.t97 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X54 G1_1 G1_1.t50 G1_2.t4 VDD.t9 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X55 SD0_1 G0_2.t8 G1_1.t91 VSS.t9 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X56 SD0_1 G0_1.t7 VSS.t10 VSS.t9 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X57 G1_2 G1_1.t48 G1_1.t49 VDD.t38 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X58 VSS G3_1.t82 G3_1.t83 VSS.t101 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X59 VDD G1_2.t42 G1_2.t43 VDD.t1 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X60 G1_1 G0_2.t9 SD0_1.t22 VSS.t0 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X61 VSS G3_1.t80 G3_1.t81 VSS.t99 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X62 SD2_0 G1_1.t105 G3_2.t24 VDD.t59 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X63 SD0_1 G0_1.t8 VSS.t32 VSS.t31 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X64 G1_2 G1_1.t46 G1_1.t47 VDD.t8 pfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X65 SD2_0 G1_2.t106 VDD.t104 VDD.t41 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X66 SD2_0 G1_1.t106 G3_2.t25 VDD.t13 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X67 G1_2 G1_1.t44 G1_1.t45 VDD.t7 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X68 VSS G3_1.t78 G3_1.t79 VSS.t98 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X69 G3_1 G3_1.t34 VSS.t143 VSS.t96 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X70 SD2_0 G1_2.t107 VDD.t103 VDD.t3 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X71 VSS G0_1.t9 SD0_1.t41 VSS.t33 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X72 G1_2 G1_1.t42 G1_1.t43 VDD.t32 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X73 SD2_0 G1_1.t107 G3_2.t26 VDD.t52 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X74 G1_1 G1_1.t40 G1_2.t89 VDD.t5 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X75 SD0_1 G0_1.t10 VSS.t66 VSS.t4 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X76 SD0_1 G0_1.t11 VSS.t67 VSS.t2 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X77 SD0_1 G0_2.t10 G1_1.t90 VSS.t5 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X78 G3_1 G3_2.t86 G3_2.t87 VSS.t97 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X79 VSS G0_1.t12 SD0_1.t47 VSS.t43 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X80 G1_1 G0_2.t11 SD0_1.t20 VSS.t1 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X81 SD0_1 G0_2.t12 G1_1.t89 VSS.t12 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X82 G1_1 G1_1.t38 G1_2.t95 VDD.t20 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X83 G3_2 G1_1.t110 SD2_0.t41 VDD.t66 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X84 SD0_1 G0_2.t13 G1_1.t88 VSS.t13 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X85 G1_1 G0_2.t14 SD0_1.t17 VSS.t16 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X86 G1_1 G1_1.t36 G1_2.t94 VDD.t4 pfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X87 VDD G1_2.t40 G1_2.t41 VDD.t48 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X88 G3_1 G3_2.t84 G3_2.t85 VSS.t96 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X89 SD2_0 G1_2.t108 VDD.t100 VDD.t43 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X90 G1_1 G0_2.t15 SD0_1.t16 VSS.t3 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X91 SD0_1 G0_2.t16 G1_1.t87 VSS.t59 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X92 SD0_1 G0_1.t13 VSS.t51 VSS.t50 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X93 G3_2 G1_1.t112 SD2_0.t42 VDD.t50 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X94 G1_2 G1_2.t58 VDD.t99 VDD.t38 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X95 VSS G0_1.t14 SD0_1.t38 VSS.t25 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X96 G3_2 G3_2.t34 G3_1.t20 VSS.t95 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X97 G3_2 G1_1.t113 SD2_0.t43 VDD.t61 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X98 VSS G3_1.t76 G3_1.t77 VSS.t94 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X99 G1_2 G1_2.t64 VDD.t98 VDD.t8 pfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X100 VSS G0_1.t15 SD0_1.t39 VSS.t28 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X101 G1_1 G1_1.t34 G1_2.t93 VDD.t6 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X102 VSS G3_1.t74 G3_1.t75 VSS.t90 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X103 G1_2 G1_2.t56 VDD.t97 VDD.t7 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X104 G3_1 G3_1.t32 VSS.t138 VSS.t89 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X105 G3_2 G1_1.t115 SD2_0.t44 VDD.t45 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X106 G1_2 G1_2.t60 VDD.t96 VDD.t32 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X107 SD0_1 G0_1.t16 VSS.t63 VSS.t20 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X108 G1_2 G1_1.t32 G1_1.t33 VDD.t73 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X109 VDD G1_2.t113 SD2_0.t28 VDD.t29 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X110 VSS G0_1.t17 SD0_1.t56 VSS.t1 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X111 VDD G1_2.t114 SD2_0.t27 VDD.t17 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X112 G3_1 G3_1.t52 VSS.t137 VSS.t88 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X113 VDD G1_2.t115 SD2_0.t26 VDD.t2 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X114 SD0_1 G0_1.t18 VSS.t60 VSS.t59 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X115 VSS G3_1.t72 G3_1.t73 VSS.t95 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X116 SD2_0 G1_2.t116 VDD.t90 VDD.t89 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X117 G3_2 G3_2.t42 G3_1.t19 VSS.t94 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X118 G3_1 G3_2.t82 G3_2.t83 VSS.t93 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X119 G3_1 G3_2.t80 G3_2.t81 VSS.t92 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X120 SD2_0 G1_2.t117 VDD.t88 VDD.t87 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X121 VDD G1_2.t38 G1_2.t39 VDD.t20 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X122 G1_1 G1_1.t30 G1_2.t87 VDD.t48 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X123 G1_1 G0_2.t17 SD0_1.t14 VSS.t42 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X124 G1_2 G1_2.t62 VDD.t84 VDD.t36 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X125 G3_1 G3_2.t78 G3_2.t79 VSS.t91 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X126 VDD G1_2.t36 G1_2.t37 VDD.t4 pfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X127 SD0_1 G0_2.t18 G1_1.t86 VSS.t40 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X128 G3_2 G3_2.t94 G3_1.t15 VSS.t90 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X129 G3_1 G3_2.t76 G3_2.t77 VSS.t89 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X130 SD2_0 G1_1.t117 G3_2.t13 VDD.t41 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X131 SD2_0 G1_2.t119 VDD.t80 VDD.t13 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X132 SD2_0 G1_1.t118 G3_2.t14 VDD.t3 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X133 G1_1 G0_2.t19 SD0_1.t12 VSS.t68 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X134 SD0_1 G0_2.t20 G1_1.t85 VSS.t50 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X135 G3_1 G3_2.t74 G3_2.t75 VSS.t88 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X136 SD2_0 G1_1.t119 G3_2.t0 VDD.t0 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X137 SD2_0 G1_2.t120 VDD.t79 VDD.t10 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X138 SD0_1 G0_2.t21 G1_1.t84 VSS.t38 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X139 G3_1 G3_2.t72 G3_2.t73 VSS.t87 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X140 VDD G1_2.t121 SD2_0.t21 VDD.t9 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X141 G3_2 G1_1.t120 SD2_0.t1 VDD.t1 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X142 VDD G1_2.t34 G1_2.t35 VDD.t6 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X143 G3_1 G3_1.t50 VSS.t134 VSS.t93 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X144 G3_1 G3_1.t48 VSS.t133 VSS.t92 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X145 G1_2 G1_2.t54 VDD.t74 VDD.t73 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X146 SD0_1 G0_1.t19 VSS.t62 VSS.t61 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X147 VDD G1_2.t32 G1_2.t33 VDD.t25 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X148 VDD G1_2.t30 G1_2.t31 VDD.t15 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X149 G3_1 G3_1.t46 VSS.t132 VSS.t91 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X150 VDD G1_2.t123 SD2_0.t20 VDD.t66 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X151 SD0_1 G0_1.t20 VSS.t15 VSS.t14 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X152 VSS G3_1.t70 G3_1.t71 VSS.t84 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X153 VSS G0_1.t21 SD0_1.t35 VSS.t16 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X154 VDD G1_2.t124 SD2_0.t19 VDD.t5 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X155 SD0_1 G0_2.t22 G1_1.t83 VSS.t19 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X156 G3_1 G3_1.t44 VSS.t129 VSS.t87 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X157 G3_2 G3_2.t92 G3_1.t11 VSS.t86 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X158 VSS G0_1.t22 SD0_1.t59 VSS.t68 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X159 VDD G1_2.t125 SD2_0.t18 VDD.t61 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X160 G1_2 G1_1.t28 G1_1.t29 VDD.t36 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X161 G1_1 G0_2.t23 SD0_1.t8 VSS.t43 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X162 G1_2 G1_2.t68 VDD.t60 VDD.t59 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X163 G1_1 G0_2.t24 SD0_1.t7 VSS.t33 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X164 G3_1 G3_2.t70 G3_2.t71 VSS.t85 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X165 G1_2 G1_2.t18 VDD.t53 VDD.t52 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X166 G3_2 G3_2.t50 G3_1.t9 VSS.t84 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X167 G3_1 G3_2.t68 G3_2.t69 VSS.t83 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X168 G3_2 G1_1.t121 SD2_0.t2 VDD.t2 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X169 SD2_0 G1_1.t122 G3_2.t29 VDD.t38 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X170 G1_1 G0_2.t25 SD0_1.t6 VSS.t45 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X171 VSS G3_1.t68 G3_1.t69 VSS.t86 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X172 SD2_0 G1_1.t123 G3_2.t30 VDD.t89 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X173 G1_1 G1_1.t26 G1_2.t82 VDD.t25 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X174 SD0_1 G0_2.t26 G1_1.t82 VSS.t61 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X175 SD2_0 G1_1.t125 G3_2.t31 VDD.t87 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X176 G1_1 G1_1.t24 G1_2.t86 VDD.t15 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X177 VSS G0_1.t23 SD0_1.t60 VSS.t71 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X178 SD2_0 G1_1.t127 G3_2.t21 VDD.t8 pfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X179 SD2_0 G1_1.t128 G3_2.t22 VDD.t7 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X180 G3_1 G3_2.t66 G3_2.t67 VSS.t82 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X181 SD2_0 G1_1.t129 G3_2.t23 VDD.t32 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X182 G1_2 G1_1.t22 G1_1.t23 VDD.t43 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X183 G3_2 G3_2.t52 G3_1.t6 VSS.t81 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X184 G3_1 G3_1.t42 VSS.t126 VSS.t79 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X185 G3_2 G3_2.t56 G3_1.t5 VSS.t80 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X186 VDD G1_2.t28 G1_2.t29 VDD.t50 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X187 G3_1 G3_1.t94 VSS.t125 VSS.t85 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X188 SD2_0 G1_2.t128 VDD.t57 VDD.t0 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X189 SD2_0 G1_1.t130 G3_2.t15 VDD.t10 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X190 G3_1 G3_1.t92 VSS.t124 VSS.t83 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X191 G3_2 G1_1.t131 SD2_0.t48 VDD.t9 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X192 VDD G1_2.t129 SD2_0.t16 VDD.t1 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X193 G1_2 G1_1.t20 G1_1.t21 VDD.t59 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X194 SD0_1 G0_1.t24 VSS.t55 VSS.t5 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X195 VSS G0_1.t25 SD0_1.t52 VSS.t56 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X196 G3_2 G1_1.t132 SD2_0.t49 VDD.t20 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X197 VDD G1_2.t130 SD2_0.t15 VDD.t48 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X198 G3_2 G1_1.t133 SD2_0.t3 VDD.t4 pfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X199 G3_1 G3_1.t90 VSS.t123 VSS.t82 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X200 G1_2 G1_1.t18 G1_1.t19 VDD.t52 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X201 G1_1 G1_1.t16 G1_2.t74 VDD.t29 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X202 VDD G1_2.t26 G1_2.t27 VDD.t45 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X203 VSS G3_1.t66 G3_1.t67 VSS.t81 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X204 G3_1 G3_2.t64 G3_2.t65 VSS.t79 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X205 VSS G3_1.t64 G3_1.t65 VSS.t80 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X206 VSS G3_1.t62 G3_1.t63 VSS.t78 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X207 G1_1 G1_1.t14 G1_2.t73 VDD.t17 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X208 G3_2 G1_1.t136 SD2_0.t4 VDD.t5 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X209 G3_2 G1_1.t137 SD2_0.t5 VDD.t6 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X210 SD2_0 G1_1.t138 G3_2.t27 VDD.t73 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X211 G1_2 G1_2.t52 VDD.t44 VDD.t43 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X212 G1_2 G1_2.t6 VDD.t42 VDD.t41 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X213 G1_1 G1_1.t12 G1_2.t80 VDD.t50 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X214 G1_2 G1_2.t16 VDD.t40 VDD.t3 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X215 G1_2 G1_1.t10 G1_1.t11 VDD.t13 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X216 G3_2 G3_2.t54 G3_1.t3 VSS.t78 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X217 VSS G0_1.t26 SD0_1.t49 VSS.t42 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X218 SD0_1 G0_1.t27 VSS.t54 VSS.t12 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X219 SD2_0 G1_2.t134 VDD.t39 VDD.t38 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X220 G3_1 G3_1.t88 VSS.t116 VSS.t77 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X221 G3_1 G3_1.t86 VSS.t115 VSS.t76 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X222 SD2_0 G1_2.t135 VDD.t37 VDD.t36 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X223 G1_1 G0_2.t27 SD0_1.t4 VSS.t74 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X224 SD2_0 G1_2.t136 VDD.t35 VDD.t8 pfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X225 SD2_0 G1_2.t137 VDD.t34 VDD.t7 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X226 SD0_1 G0_2.t28 G1_1.t81 VSS.t4 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X227 SD2_0 G1_2.t138 VDD.t33 VDD.t32 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X228 G1_1 G1_1.t8 G1_2.t78 VDD.t45 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X229 VDD G1_2.t24 G1_2.t25 VDD.t29 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X230 VDD G1_2.t22 G1_2.t23 VDD.t17 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X231 G1_1 G1_1.t6 G1_2.t77 VDD.t66 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X232 SD0_1 G0_1.t28 VSS.t21 VSS.t13 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X233 G1_1 G0_2.t29 SD0_1.t2 VSS.t6 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X234 VSS G3_1.t60 G3_1.t61 VSS.t75 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X235 SD0_1 G0_2.t30 G1_1.t80 VSS.t20 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X236 G3_1 G3_2.t62 G3_2.t63 VSS.t77 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X237 VSS G3_1.t58 G3_1.t59 VSS.t106 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X238 G1_1 G1_1.t4 G1_2.t76 VDD.t61 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X239 G3_1 G3_2.t60 G3_2.t61 VSS.t76 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X240 VSS G3_1.t56 G3_1.t57 VSS.t104 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X241 VDD G1_2.t139 SD2_0.t9 VDD.t25 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X242 VDD G1_2.t140 SD2_0.t8 VDD.t20 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X243 G3_2 G1_1.t143 SD2_0.t60 VDD.t48 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X244 VDD G1_2.t141 SD2_0.t7 VDD.t4 pfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X245 VDD G1_2.t142 SD2_0.t6 VDD.t15 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X246 G1_2 G1_1.t2 G1_1.t3 VDD.t41 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X247 G1_2 G1_2.t66 VDD.t14 VDD.t13 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X248 G1_2 G1_1.t0 G1_1.t1 VDD.t3 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X249 G1_1 G0_2.t31 SD0_1.t0 VSS.t56 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X250 VSS G0_1.t29 SD0_1.t37 VSS.t22 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X251 SD0_1 G0_1.t30 VSS.t44 VSS.t11 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X252 VSS G3_1.t54 G3_1.t55 VSS.t103 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X253 VSS G0_1.t31 SD0_1.t46 VSS.t45 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X254 G3_2 G3_2.t38 G3_1.t0 VSS.t75 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X255 VDD G1_2.t20 G1_2.t21 VDD.t2 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
R0 G3_2.n117 G3_2.n116 107.18
R1 G3_2.n96 G3_2.n95 107.18
R2 G3_2.n125 G3_2.n124 103.823
R3 G3_2.n123 G3_2.n122 103.823
R4 G3_2.n121 G3_2.n120 103.823
R5 G3_2.n119 G3_2.n118 103.823
R6 G3_2.n136 G3_2.n47 103.823
R7 G3_2.n135 G3_2.n134 103.823
R8 G3_2.n24 G3_2.n23 103.823
R9 G3_2.n29 G3_2.n28 103.823
R10 G3_2.n34 G3_2.n33 103.823
R11 G3_2.n39 G3_2.n38 103.823
R12 G3_2.n40 G3_2.n2 103.823
R13 G3_2.n149 G3_2.n148 103.823
R14 G3_2.n154 G3_2.n153 103.823
R15 G3_2.n23 G3_2.n22 23.4254
R16 G3_2.n155 G3_2.n154 23.2794
R17 G3_2.n124 G3_2.n123 21.0894
R18 G3_2.n122 G3_2.n121 21.0894
R19 G3_2.n120 G3_2.n119 21.0894
R20 G3_2.n118 G3_2.n117 21.0894
R21 G3_2.n95 G3_2.n47 21.0894
R22 G3_2.n136 G3_2.n135 21.0894
R23 G3_2.n134 G3_2.n125 21.0894
R24 G3_2.n28 G3_2.n24 21.0894
R25 G3_2.n33 G3_2.n29 21.0894
R26 G3_2.n38 G3_2.n34 21.0894
R27 G3_2.n148 G3_2.n2 21.0894
R28 G3_2.n40 G3_2.n39 21.0894
R29 G3_2.n153 G3_2.n149 21.0894
R30 G3_2.n125 G3_2.t64 14.0895
R31 G3_2.n123 G3_2.t84 14.0895
R32 G3_2.n121 G3_2.t88 14.0895
R33 G3_2.n119 G3_2.t76 14.0895
R34 G3_2.n117 G3_2.t62 14.0895
R35 G3_2.n47 G3_2.t74 14.0895
R36 G3_2.n135 G3_2.t60 14.0895
R37 G3_2.n23 G3_2.t56 12.7025
R38 G3_2.n24 G3_2.t70 12.7025
R39 G3_2.n29 G3_2.t90 12.7025
R40 G3_2.n34 G3_2.t72 12.7025
R41 G3_2.n39 G3_2.t66 12.7025
R42 G3_2.n2 G3_2.t78 12.7025
R43 G3_2.n149 G3_2.t68 12.7025
R44 G3_2.n154 G3_2.t82 12.7025
R45 G3_2.n50 G3_2.t54 10.7315
R46 G3_2.n53 G3_2.t46 10.7315
R47 G3_2.n56 G3_2.t50 10.7315
R48 G3_2.n59 G3_2.t42 10.7315
R49 G3_2.n116 G3_2.t36 10.7315
R50 G3_2.n96 G3_2.t86 10.7315
R51 G3_2.n94 G3_2.t38 10.7315
R52 G3_2.n22 G3_2.t80 10.3665
R53 G3_2.n27 G3_2.t40 10.3665
R54 G3_2.n32 G3_2.t92 10.3665
R55 G3_2.n37 G3_2.t44 10.3665
R56 G3_2.n152 G3_2.t58 10.3665
R57 G3_2.n156 G3_2.t52 10.3665
R58 G3_2.n142 G3_2.t94 9.7761
R59 G3_2.n130 G3_2.t32 8.1765
R60 G3_2.n8 G3_2.t34 8.1765
R61 G3_2.n148 G3_2.n147 8.17038
R62 G3_2.n42 G3_2.n41 8.02202
R63 G3_2.n8 G3_2.n7 8.01152
R64 G3_2.n6 G3_2.n3 8.008
R65 G3_2.n141 G3_2.n140 8.0005
R66 G3_2.n130 G3_2.n126 8.0005
R67 G3_2.n132 G3_2.n129 8.0005
R68 G3_2.n12 G3_2.n11 8.0005
R69 G3_2.n17 G3_2.n13 8.0005
R70 G3_2.n19 G3_2.n18 8.0005
R71 G3_2.n10 G3_2.n9 8.0005
R72 G3_2.n12 G3_2.t48 7.8845
R73 G3_2.n53 G3_2.n52 7.59736
R74 G3_2.n50 G3_2.n49 7.58813
R75 G3_2.n59 G3_2.n58 7.50659
R76 G3_2.n94 G3_2.n93 7.50659
R77 G3_2.n56 G3_2.n55 7.50213
R78 G3_2.n32 G3_2.n31 7.49478
R79 G3_2.n22 G3_2.n21 7.49191
R80 G3_2.n152 G3_2.n151 7.49008
R81 G3_2.n27 G3_2.n26 7.48719
R82 G3_2.n37 G3_2.n36 7.47354
R83 G3_2.n114 G3_2.n61 6.0756
R84 G3_2.n98 G3_2.t21 6.0756
R85 G3_2.n115 G3_2.n60 6.03311
R86 G3_2.n97 G3_2.t87 6.01354
R87 G3_2.n97 G3_2.n96 4.09218
R88 G3_2.n116 G3_2.n115 4.07208
R89 G3_2.n157 G3_2.n156 4.0005
R90 G3_2.n140 G3_2.n139 3.56662
R91 G3_2.n133 G3_2.n126 3.54789
R92 G3_2.n137 G3_2.n46 3.51501
R93 G3_2.n157 G3_2.n1 3.49193
R94 G3_2.n6 G3_2.n5 3.48507
R95 G3_2.n16 G3_2.n15 3.48115
R96 G3_2.n129 G3_2.n128 3.47959
R97 G3_2.n124 G3_2.n50 3.3585
R98 G3_2.n122 G3_2.n53 3.3585
R99 G3_2.n120 G3_2.n56 3.3585
R100 G3_2.n118 G3_2.n59 3.3585
R101 G3_2.n95 G3_2.n94 3.3585
R102 G3_2.n63 G3_2.t14 3.03383
R103 G3_2.n63 G3_2.n62 3.03383
R104 G3_2.n67 G3_2.t30 3.03383
R105 G3_2.n67 G3_2.n66 3.03383
R106 G3_2.n71 G3_2.t6 3.03383
R107 G3_2.n71 G3_2.n70 3.03383
R108 G3_2.n75 G3_2.t26 3.03383
R109 G3_2.n75 G3_2.n74 3.03383
R110 G3_2.n79 G3_2.t15 3.03383
R111 G3_2.n79 G3_2.n78 3.03383
R112 G3_2.n83 G3_2.t24 3.03383
R113 G3_2.n83 G3_2.n82 3.03383
R114 G3_2.n87 G3_2.t31 3.03383
R115 G3_2.n87 G3_2.n86 3.03383
R116 G3_2.n91 G3_2.t13 3.03383
R117 G3_2.n91 G3_2.n90 3.03383
R118 G3_2.n89 G3_2.t0 3.03383
R119 G3_2.n89 G3_2.n88 3.03383
R120 G3_2.n85 G3_2.t23 3.03383
R121 G3_2.n85 G3_2.n84 3.03383
R122 G3_2.n81 G3_2.t25 3.03383
R123 G3_2.n81 G3_2.n80 3.03383
R124 G3_2.n77 G3_2.t27 3.03383
R125 G3_2.n77 G3_2.n76 3.03383
R126 G3_2.n73 G3_2.t29 3.03383
R127 G3_2.n73 G3_2.n72 3.03383
R128 G3_2.n69 G3_2.t7 3.03383
R129 G3_2.n69 G3_2.n68 3.03383
R130 G3_2.n65 G3_2.t22 3.03383
R131 G3_2.n65 G3_2.n64 3.03383
R132 G3_2.n113 G3_2.n63 3.00941
R133 G3_2.n111 G3_2.n67 3.00941
R134 G3_2.n109 G3_2.n71 3.00941
R135 G3_2.n107 G3_2.n75 3.00941
R136 G3_2.n105 G3_2.n79 3.00941
R137 G3_2.n103 G3_2.n83 3.00941
R138 G3_2.n101 G3_2.n87 3.00941
R139 G3_2.n99 G3_2.n91 3.00941
R140 G3_2.n100 G3_2.n89 2.99767
R141 G3_2.n102 G3_2.n85 2.99767
R142 G3_2.n104 G3_2.n81 2.99767
R143 G3_2.n106 G3_2.n77 2.99767
R144 G3_2.n108 G3_2.n73 2.99767
R145 G3_2.n110 G3_2.n69 2.99767
R146 G3_2.n112 G3_2.n65 2.99767
R147 G3_2.n132 G3_2.n131 2.88412
R148 G3_2.n144 G3_2.n143 2.88107
R149 G3_2.n43 G3_2.n13 2.8805
R150 G3_2.n146 G3_2.n3 2.8805
R151 G3_2.n1 G3_2.t83 2.7305
R152 G3_2.n1 G3_2.n0 2.7305
R153 G3_2.n49 G3_2.t85 2.7305
R154 G3_2.n49 G3_2.n48 2.7305
R155 G3_2.n52 G3_2.t89 2.7305
R156 G3_2.n52 G3_2.n51 2.7305
R157 G3_2.n55 G3_2.t77 2.7305
R158 G3_2.n55 G3_2.n54 2.7305
R159 G3_2.n58 G3_2.t63 2.7305
R160 G3_2.n58 G3_2.n57 2.7305
R161 G3_2.n93 G3_2.t75 2.7305
R162 G3_2.n93 G3_2.n92 2.7305
R163 G3_2.n139 G3_2.t61 2.7305
R164 G3_2.n139 G3_2.n138 2.7305
R165 G3_2.n128 G3_2.t65 2.7305
R166 G3_2.n128 G3_2.n127 2.7305
R167 G3_2.n21 G3_2.t81 2.7305
R168 G3_2.n21 G3_2.n20 2.7305
R169 G3_2.n26 G3_2.t71 2.7305
R170 G3_2.n26 G3_2.n25 2.7305
R171 G3_2.n31 G3_2.t91 2.7305
R172 G3_2.n31 G3_2.n30 2.7305
R173 G3_2.n36 G3_2.t73 2.7305
R174 G3_2.n36 G3_2.n35 2.7305
R175 G3_2.n15 G3_2.t67 2.7305
R176 G3_2.n15 G3_2.n14 2.7305
R177 G3_2.n5 G3_2.t79 2.7305
R178 G3_2.n5 G3_2.n4 2.7305
R179 G3_2.n151 G3_2.t69 2.7305
R180 G3_2.n151 G3_2.n150 2.7305
R181 G3_2.n28 G3_2.n27 2.3365
R182 G3_2.n33 G3_2.n32 2.3365
R183 G3_2.n38 G3_2.n37 2.3365
R184 G3_2.n153 G3_2.n152 2.3365
R185 G3_2.n44 G3_2.n43 2.2505
R186 G3_2.n131 G3_2.n45 2.2505
R187 G3_2.n146 G3_2.n145 2.2505
R188 G3_2.n134 G3_2.n133 2.22123
R189 G3_2.n13 G3_2.n12 2.1905
R190 G3_2.n41 G3_2.n19 2.1905
R191 G3_2.n9 G3_2.n8 2.1905
R192 G3_2.n137 G3_2.n136 2.09002
R193 G3_2.n132 G3_2.n130 2.0445
R194 G3_2.n148 G3_2.n3 2.0445
R195 G3_2.n143 G3_2.n142 1.75738
R196 G3_2.n115 G3_2.n114 1.74861
R197 G3_2.n98 G3_2.n97 1.7405
R198 G3_2.n45 G3_2.n44 1.6125
R199 G3_2.n133 G3_2.n132 1.41823
R200 G3_2.n145 G3_2.n44 1.27751
R201 G3_2.n141 G3_2.n137 1.06317
R202 G3_2.n145 G3_2.n144 0.952132
R203 G3_2.n144 G3_2.n45 0.640509
R204 G3_2.n142 G3_2.n141 0.495409
R205 G3_2.n113 G3_2.n112 0.331311
R206 G3_2.n112 G3_2.n111 0.331311
R207 G3_2.n111 G3_2.n110 0.331311
R208 G3_2.n110 G3_2.n109 0.331311
R209 G3_2.n109 G3_2.n108 0.331311
R210 G3_2.n108 G3_2.n107 0.331311
R211 G3_2.n107 G3_2.n106 0.331311
R212 G3_2.n106 G3_2.n105 0.331311
R213 G3_2.n105 G3_2.n104 0.331311
R214 G3_2.n104 G3_2.n103 0.331311
R215 G3_2.n103 G3_2.n102 0.331311
R216 G3_2.n102 G3_2.n101 0.331311
R217 G3_2.n101 G3_2.n100 0.331311
R218 G3_2.n100 G3_2.n99 0.331311
R219 G3_2.n19 G3_2.n13 0.2925
R220 G3_2.n9 G3_2.n3 0.2925
R221 G3_2.n114 G3_2.n113 0.259959
R222 G3_2.n99 G3_2.n98 0.259959
R223 G3_2.n41 G3_2.n40 0.1465
R224 G3_2.n156 G3_2.n155 0.1465
R225 G3_2.n43 G3_2.n42 0.0475455
R226 G3_2.n43 G3_2.n11 0.0474565
R227 G3_2.n10 G3_2.n7 0.0445816
R228 G3_2.n16 G3_2.n11 0.0435435
R229 G3_2.n7 G3_2.n6 0.0396304
R230 G3_2.n147 G3_2.n6 0.038
R231 G3_2.n42 G3_2.n18 0.0376739
R232 G3_2.n147 G3_2.n146 0.0317245
R233 G3_2.n129 G3_2.n126 0.0275
R234 G3_2.n131 G3_2.n126 0.0085
R235 G3_2.n18 G3_2.n17 0.00832609
R236 G3_2.n146 G3_2.n10 0.00784694
R237 G3_2 G3_2.n157 0.0075
R238 G3_2.n17 G3_2.n16 0.00636957
R239 G3_2.n140 G3_2.n46 0.00523684
R240 G3_2.n143 G3_2.n46 0.00176761
R241 G3_1.n179 G3_1.t36 34.1564
R242 G3_1.n135 G3_1.t72 12.0455
R243 G3_1.n132 G3_1.t46 12.0455
R244 G3_1.n113 G3_1.t78 12.0455
R245 G3_1.n110 G3_1.t90 12.0455
R246 G3_1.n91 G3_1.t84 12.0455
R247 G3_1.n88 G3_1.t44 12.0455
R248 G3_1.n69 G3_1.t68 12.0455
R249 G3_1.n66 G3_1.t38 12.0455
R250 G3_1.n47 G3_1.t82 12.0455
R251 G3_1.n44 G3_1.t94 12.0455
R252 G3_1.n25 G3_1.t64 12.0455
R253 G3_1.n22 G3_1.t48 12.0455
R254 G3_1.n176 G3_1.t50 12.0455
R255 G3_1.n178 G3_1.t66 11.9725
R256 G3_1.n157 G3_1.t80 11.5345
R257 G3_1.n154 G3_1.t92 10.8775
R258 G3_1.n169 G3_1.t60 10.7315
R259 G3_1.n166 G3_1.t52 10.7315
R260 G3_1.n144 G3_1.t86 10.7315
R261 G3_1.n125 G3_1.t56 10.7315
R262 G3_1.n122 G3_1.t42 10.7315
R263 G3_1.n103 G3_1.t62 10.7315
R264 G3_1.n100 G3_1.t34 10.7315
R265 G3_1.n81 G3_1.t54 10.7315
R266 G3_1.n78 G3_1.t40 10.7315
R267 G3_1.n59 G3_1.t70 10.7315
R268 G3_1.n56 G3_1.t32 10.7315
R269 G3_1.n37 G3_1.t76 10.7315
R270 G3_1.n34 G3_1.t88 10.7315
R271 G3_1.n16 G3_1.t58 10.7315
R272 G3_1.n147 G3_1.t74 10.5125
R273 G3_1.n19 G3_1.n16 4.05396
R274 G3_1.n23 G3_1.n22 4.0005
R275 G3_1.n26 G3_1.n25 4.0005
R276 G3_1.n35 G3_1.n34 4.0005
R277 G3_1.n38 G3_1.n37 4.0005
R278 G3_1.n45 G3_1.n44 4.0005
R279 G3_1.n48 G3_1.n47 4.0005
R280 G3_1.n57 G3_1.n56 4.0005
R281 G3_1.n60 G3_1.n59 4.0005
R282 G3_1.n67 G3_1.n66 4.0005
R283 G3_1.n70 G3_1.n69 4.0005
R284 G3_1.n79 G3_1.n78 4.0005
R285 G3_1.n82 G3_1.n81 4.0005
R286 G3_1.n89 G3_1.n88 4.0005
R287 G3_1.n92 G3_1.n91 4.0005
R288 G3_1.n101 G3_1.n100 4.0005
R289 G3_1.n104 G3_1.n103 4.0005
R290 G3_1.n111 G3_1.n110 4.0005
R291 G3_1.n114 G3_1.n113 4.0005
R292 G3_1.n123 G3_1.n122 4.0005
R293 G3_1.n126 G3_1.n125 4.0005
R294 G3_1.n133 G3_1.n132 4.0005
R295 G3_1.n136 G3_1.n135 4.0005
R296 G3_1.n145 G3_1.n144 4.0005
R297 G3_1.n148 G3_1.n147 4.0005
R298 G3_1.n155 G3_1.n154 4.0005
R299 G3_1.n158 G3_1.n157 4.0005
R300 G3_1.n167 G3_1.n166 4.0005
R301 G3_1.n170 G3_1.n169 4.0005
R302 G3_1.n177 G3_1.n176 4.0005
R303 G3_1.n181 G3_1.n180 4.0005
R304 G3_1.n154 G3_1.n153 3.5045
R305 G3_1.n19 G3_1.n18 3.4792
R306 G3_1.n32 G3_1.n31 3.4792
R307 G3_1.n41 G3_1.n40 3.4792
R308 G3_1.n54 G3_1.n53 3.4792
R309 G3_1.n63 G3_1.n62 3.4792
R310 G3_1.n76 G3_1.n75 3.4792
R311 G3_1.n85 G3_1.n84 3.4792
R312 G3_1.n98 G3_1.n97 3.4792
R313 G3_1.n107 G3_1.n106 3.4792
R314 G3_1.n120 G3_1.n119 3.4792
R315 G3_1.n129 G3_1.n128 3.4792
R316 G3_1.n142 G3_1.n141 3.4792
R317 G3_1.n164 G3_1.n163 3.4792
R318 G3_1.n173 G3_1.n172 3.4792
R319 G3_1.n151 G3_1.n150 3.47724
R320 G3_1.n186 G3_1.n185 3.47528
R321 G3_1.n20 G3_1.n15 3.47333
R322 G3_1.n29 G3_1.n28 3.47333
R323 G3_1.n42 G3_1.n13 3.47333
R324 G3_1.n51 G3_1.n50 3.47333
R325 G3_1.n64 G3_1.n11 3.47333
R326 G3_1.n73 G3_1.n72 3.47333
R327 G3_1.n86 G3_1.n9 3.47333
R328 G3_1.n95 G3_1.n94 3.47333
R329 G3_1.n108 G3_1.n7 3.47333
R330 G3_1.n117 G3_1.n116 3.47333
R331 G3_1.n130 G3_1.n5 3.47333
R332 G3_1.n139 G3_1.n138 3.47333
R333 G3_1.n174 G3_1.n1 3.47333
R334 G3_1.n161 G3_1.n160 3.45963
R335 G3_1.n152 G3_1.n3 3.44202
R336 G3_1.n186 G3_1.n183 3.38528
R337 G3_1.n157 G3_1.n156 2.8475
R338 G3_1.n185 G3_1.t6 2.7305
R339 G3_1.n185 G3_1.n184 2.7305
R340 G3_1.n183 G3_1.t67 2.7305
R341 G3_1.n183 G3_1.n182 2.7305
R342 G3_1.n172 G3_1.t61 2.7305
R343 G3_1.n172 G3_1.n171 2.7305
R344 G3_1.n1 G3_1.t0 2.7305
R345 G3_1.n1 G3_1.n0 2.7305
R346 G3_1.n160 G3_1.t81 2.7305
R347 G3_1.n160 G3_1.n159 2.7305
R348 G3_1.n163 G3_1.t24 2.7305
R349 G3_1.n163 G3_1.n162 2.7305
R350 G3_1.n3 G3_1.t15 2.7305
R351 G3_1.n3 G3_1.n2 2.7305
R352 G3_1.n150 G3_1.t75 2.7305
R353 G3_1.n150 G3_1.n149 2.7305
R354 G3_1.n138 G3_1.t73 2.7305
R355 G3_1.n138 G3_1.n137 2.7305
R356 G3_1.n141 G3_1.t20 2.7305
R357 G3_1.n141 G3_1.n140 2.7305
R358 G3_1.n128 G3_1.t57 2.7305
R359 G3_1.n128 G3_1.n127 2.7305
R360 G3_1.n5 G3_1.t29 2.7305
R361 G3_1.n5 G3_1.n4 2.7305
R362 G3_1.n116 G3_1.t79 2.7305
R363 G3_1.n116 G3_1.n115 2.7305
R364 G3_1.n119 G3_1.t23 2.7305
R365 G3_1.n119 G3_1.n118 2.7305
R366 G3_1.n106 G3_1.t63 2.7305
R367 G3_1.n106 G3_1.n105 2.7305
R368 G3_1.n7 G3_1.t3 2.7305
R369 G3_1.n7 G3_1.n6 2.7305
R370 G3_1.n94 G3_1.t85 2.7305
R371 G3_1.n94 G3_1.n93 2.7305
R372 G3_1.n97 G3_1.t30 2.7305
R373 G3_1.n97 G3_1.n96 2.7305
R374 G3_1.n84 G3_1.t55 2.7305
R375 G3_1.n84 G3_1.n83 2.7305
R376 G3_1.n9 G3_1.t28 2.7305
R377 G3_1.n9 G3_1.n8 2.7305
R378 G3_1.n72 G3_1.t69 2.7305
R379 G3_1.n72 G3_1.n71 2.7305
R380 G3_1.n75 G3_1.t11 2.7305
R381 G3_1.n75 G3_1.n74 2.7305
R382 G3_1.n62 G3_1.t71 2.7305
R383 G3_1.n62 G3_1.n61 2.7305
R384 G3_1.n11 G3_1.t9 2.7305
R385 G3_1.n11 G3_1.n10 2.7305
R386 G3_1.n50 G3_1.t83 2.7305
R387 G3_1.n50 G3_1.n49 2.7305
R388 G3_1.n53 G3_1.t26 2.7305
R389 G3_1.n53 G3_1.n52 2.7305
R390 G3_1.n40 G3_1.t77 2.7305
R391 G3_1.n40 G3_1.n39 2.7305
R392 G3_1.n13 G3_1.t19 2.7305
R393 G3_1.n13 G3_1.n12 2.7305
R394 G3_1.n28 G3_1.t65 2.7305
R395 G3_1.n28 G3_1.n27 2.7305
R396 G3_1.n31 G3_1.t5 2.7305
R397 G3_1.n31 G3_1.n30 2.7305
R398 G3_1.n18 G3_1.t59 2.7305
R399 G3_1.n18 G3_1.n17 2.7305
R400 G3_1.n15 G3_1.t31 2.7305
R401 G3_1.n15 G3_1.n14 2.7305
R402 G3_1.n147 G3_1.n146 2.5555
R403 G3_1.n169 G3_1.n168 2.3365
R404 G3_1.n166 G3_1.n165 2.3365
R405 G3_1.n144 G3_1.n143 2.3365
R406 G3_1.n135 G3_1.n134 2.3365
R407 G3_1.n132 G3_1.n131 2.3365
R408 G3_1.n125 G3_1.n124 2.3365
R409 G3_1.n122 G3_1.n121 2.3365
R410 G3_1.n113 G3_1.n112 2.3365
R411 G3_1.n110 G3_1.n109 2.3365
R412 G3_1.n103 G3_1.n102 2.3365
R413 G3_1.n100 G3_1.n99 2.3365
R414 G3_1.n91 G3_1.n90 2.3365
R415 G3_1.n88 G3_1.n87 2.3365
R416 G3_1.n81 G3_1.n80 2.3365
R417 G3_1.n78 G3_1.n77 2.3365
R418 G3_1.n69 G3_1.n68 2.3365
R419 G3_1.n66 G3_1.n65 2.3365
R420 G3_1.n59 G3_1.n58 2.3365
R421 G3_1.n56 G3_1.n55 2.3365
R422 G3_1.n47 G3_1.n46 2.3365
R423 G3_1.n44 G3_1.n43 2.3365
R424 G3_1.n37 G3_1.n36 2.3365
R425 G3_1.n34 G3_1.n33 2.3365
R426 G3_1.n25 G3_1.n24 2.3365
R427 G3_1.n22 G3_1.n21 2.3365
R428 G3_1.n176 G3_1.n175 2.3365
R429 G3_1.n180 G3_1.n179 2.3365
R430 G3_1.n181 G3_1.n177 0.313543
R431 G3_1.n26 G3_1.n23 0.313543
R432 G3_1.n48 G3_1.n45 0.313543
R433 G3_1.n70 G3_1.n67 0.313543
R434 G3_1.n92 G3_1.n89 0.313543
R435 G3_1.n114 G3_1.n111 0.313543
R436 G3_1.n136 G3_1.n133 0.313543
R437 G3_1.n158 G3_1.n155 0.313543
R438 G3_1.n38 G3_1.n35 0.284446
R439 G3_1.n60 G3_1.n57 0.284446
R440 G3_1.n82 G3_1.n79 0.284446
R441 G3_1.n104 G3_1.n101 0.284446
R442 G3_1.n126 G3_1.n123 0.284446
R443 G3_1.n170 G3_1.n167 0.284446
R444 G3_1.n148 G3_1.n145 0.283774
R445 G3_1.n152 G3_1.n151 0.117891
R446 G3_1 G3_1.n186 0.1015
R447 G3_1.n164 G3_1.n161 0.0983261
R448 G3_1.n20 G3_1.n19 0.0846304
R449 G3_1.n32 G3_1.n29 0.0846304
R450 G3_1.n42 G3_1.n41 0.0846304
R451 G3_1.n54 G3_1.n51 0.0846304
R452 G3_1.n64 G3_1.n63 0.0846304
R453 G3_1.n76 G3_1.n73 0.0846304
R454 G3_1.n86 G3_1.n85 0.0846304
R455 G3_1.n98 G3_1.n95 0.0846304
R456 G3_1.n108 G3_1.n107 0.0846304
R457 G3_1.n120 G3_1.n117 0.0846304
R458 G3_1.n130 G3_1.n129 0.0846304
R459 G3_1.n142 G3_1.n139 0.0846304
R460 G3_1.n174 G3_1.n173 0.0846304
R461 G3_1.n23 G3_1.n20 0.0795
R462 G3_1.n29 G3_1.n26 0.0795
R463 G3_1.n45 G3_1.n42 0.0795
R464 G3_1.n51 G3_1.n48 0.0795
R465 G3_1.n67 G3_1.n64 0.0795
R466 G3_1.n73 G3_1.n70 0.0795
R467 G3_1.n89 G3_1.n86 0.0795
R468 G3_1.n95 G3_1.n92 0.0795
R469 G3_1.n111 G3_1.n108 0.0795
R470 G3_1.n117 G3_1.n114 0.0795
R471 G3_1.n133 G3_1.n130 0.0795
R472 G3_1.n139 G3_1.n136 0.0795
R473 G3_1.n155 G3_1.n152 0.0795
R474 G3_1.n161 G3_1.n158 0.0795
R475 G3_1.n177 G3_1.n174 0.0795
R476 G3_1.n180 G3_1.n178 0.0735
R477 G3_1.n35 G3_1.n32 0.0539586
R478 G3_1.n41 G3_1.n38 0.0539586
R479 G3_1.n57 G3_1.n54 0.0539586
R480 G3_1.n63 G3_1.n60 0.0539586
R481 G3_1.n79 G3_1.n76 0.0539586
R482 G3_1.n85 G3_1.n82 0.0539586
R483 G3_1.n101 G3_1.n98 0.0539586
R484 G3_1.n107 G3_1.n104 0.0539586
R485 G3_1.n123 G3_1.n120 0.0539586
R486 G3_1.n129 G3_1.n126 0.0539586
R487 G3_1.n145 G3_1.n142 0.0539586
R488 G3_1.n167 G3_1.n164 0.0539586
R489 G3_1.n173 G3_1.n170 0.0539586
R490 G3_1.n151 G3_1.n148 0.0527794
R491 G3_1 G3_1.n181 0.0015
R492 VSS.n174 VSS.t76 284.212
R493 VSS.n23 VSS.t22 278.649
R494 VSS.n149 VSS.t101 273.685
R495 VSS.n160 VSS.t105 273.685
R496 VSS.n304 VSS.t59 267.932
R497 VSS.n283 VSS.t14 267.932
R498 VSS.n149 VSS.t85 263.159
R499 VSS.n160 VSS.t96 263.159
R500 VSS.n264 VSS.t1 257.214
R501 VSS.n322 VSS.t6 257.214
R502 VSS.n174 VSS.t90 252.632
R503 VSS.n246 VSS.t38 246.496
R504 VSS.n171 VSS.t95 215.79
R505 VSS.n26 VSS.t4 208.987
R506 VSS.n150 VSS.t89 205.263
R507 VSS.n159 VSS.t87 205.263
R508 VSS.n306 VSS.t0 198.269
R509 VSS.n280 VSS.t74 198.269
R510 VSS.n148 VSS.t94 194.738
R511 VSS.n163 VSS.t78 194.738
R512 VSS.n262 VSS.t61 187.553
R513 VSS.n324 VSS.t12 187.553
R514 VSS.n175 VSS.t83 184.212
R515 VSS.n244 VSS.t28 176.834
R516 VSS.n182 VSS.t81 157.895
R517 VSS.n170 VSS.t91 147.369
R518 VSS.n27 VSS.t71 139.325
R519 VSS.n293 VSS.t33 139.325
R520 VSS.n153 VSS.t84 136.843
R521 VSS.n158 VSS.t103 136.843
R522 VSS.n308 VSS.t20 128.607
R523 VSS.n278 VSS.t11 128.607
R524 VSS.n145 VSS.t77 126.317
R525 VSS.n164 VSS.t82 126.317
R526 VSS.n260 VSS.t45 117.891
R527 VSS.n327 VSS.t56 117.891
R528 VSS.n176 VSS.t99 115.79
R529 VSS.n351 VSS.t2 112.531
R530 VSS.n241 VSS.t5 107.172
R531 VSS.n188 VSS.t97 97.3689
R532 VSS.n181 VSS.t93 89.4742
R533 VSS.n169 VSS.t104 78.9479
R534 VSS.n28 VSS.t13 69.6625
R535 VSS.n292 VSS.t50 69.6625
R536 VSS.n154 VSS.t102 68.4216
R537 VSS.n155 VSS.t100 68.4216
R538 VSS.n311 VSS.t43 58.9453
R539 VSS.n276 VSS.t25 58.9453
R540 VSS.n144 VSS.t80 57.8952
R541 VSS.n165 VSS.t98 57.8952
R542 VSS.n257 VSS.t40 48.228
R543 VSS.n329 VSS.t19 48.228
R544 VSS.n177 VSS.t88 47.3689
R545 VSS.n239 VSS.t3 37.5108
R546 VSS.n66 VSS.t106 34.211
R547 VSS.n180 VSS.t75 21.0531
R548 VSS.n17 VSS.t9 10.7177
R549 VSS.n273 VSS.t31 10.7177
R550 VSS.n143 VSS.t92 10.5268
R551 VSS.n166 VSS.t79 10.5268
R552 VSS.n133 VSS.n132 6.37382
R553 VSS.n16 VSS.n15 6.36926
R554 VSS.n183 VSS.t150 6.35593
R555 VSS.n354 VSS.t67 6.35232
R556 VSS.n85 VSS.n84 6.04912
R557 VSS.n88 VSS.n87 5.2005
R558 VSS.n67 VSS.n66 5.2005
R559 VSS.n67 VSS.n65 5.2005
R560 VSS.n192 VSS.n190 5.2005
R561 VSS.n142 VSS.n140 5.2005
R562 VSS.n142 VSS.n138 5.2005
R563 VSS.n227 VSS.n143 5.2005
R564 VSS.n226 VSS.n144 5.2005
R565 VSS.n225 VSS.n145 5.2005
R566 VSS.n223 VSS.n148 5.2005
R567 VSS.n222 VSS.n149 5.2005
R568 VSS.n221 VSS.n150 5.2005
R569 VSS.n219 VSS.n153 5.2005
R570 VSS.n218 VSS.n154 5.2005
R571 VSS.n217 VSS.t86 5.2005
R572 VSS.n216 VSS.n155 5.2005
R573 VSS.n214 VSS.n158 5.2005
R574 VSS.n213 VSS.n159 5.2005
R575 VSS.n212 VSS.n160 5.2005
R576 VSS.n210 VSS.n163 5.2005
R577 VSS.n209 VSS.n164 5.2005
R578 VSS.n208 VSS.n165 5.2005
R579 VSS.n207 VSS.n166 5.2005
R580 VSS.n205 VSS.n169 5.2005
R581 VSS.n204 VSS.n170 5.2005
R582 VSS.n203 VSS.n171 5.2005
R583 VSS.n201 VSS.n174 5.2005
R584 VSS.n200 VSS.n175 5.2005
R585 VSS.n199 VSS.n176 5.2005
R586 VSS.n198 VSS.n177 5.2005
R587 VSS.n196 VSS.n180 5.2005
R588 VSS.n195 VSS.n181 5.2005
R589 VSS.n194 VSS.n182 5.2005
R590 VSS.n192 VSS.n188 5.2005
R591 VSS.n346 VSS.n344 5.2005
R592 VSS.n60 VSS.n58 5.2005
R593 VSS.n60 VSS.n56 5.2005
R594 VSS.n51 VSS.n17 5.2005
R595 VSS.n49 VSS.n20 5.2005
R596 VSS.n48 VSS.n21 5.2005
R597 VSS.n47 VSS.n22 5.2005
R598 VSS.n46 VSS.n23 5.2005
R599 VSS.n44 VSS.n26 5.2005
R600 VSS.n43 VSS.n27 5.2005
R601 VSS.n42 VSS.n28 5.2005
R602 VSS.n40 VSS.t68 5.2005
R603 VSS.n39 VSS.n31 5.2005
R604 VSS.n38 VSS.n32 5.2005
R605 VSS.n37 VSS.n33 5.2005
R606 VSS.n305 VSS.n304 5.2005
R607 VSS.n307 VSS.n306 5.2005
R608 VSS.n309 VSS.n308 5.2005
R609 VSS.n312 VSS.n311 5.2005
R610 VSS.n314 VSS.n313 5.2005
R611 VSS.n316 VSS.n315 5.2005
R612 VSS.n318 VSS.n317 5.2005
R613 VSS.n321 VSS.n320 5.2005
R614 VSS.n323 VSS.n322 5.2005
R615 VSS.n325 VSS.n324 5.2005
R616 VSS.n328 VSS.n327 5.2005
R617 VSS.n330 VSS.n329 5.2005
R618 VSS.n332 VSS.n331 5.2005
R619 VSS.n334 VSS.n333 5.2005
R620 VSS.n337 VSS.n336 5.2005
R621 VSS.n346 VSS.n342 5.2005
R622 VSS.n14 VSS.n12 5.2005
R623 VSS.n238 VSS.n237 5.2005
R624 VSS.n240 VSS.n239 5.2005
R625 VSS.n242 VSS.n241 5.2005
R626 VSS.n245 VSS.n244 5.2005
R627 VSS.n247 VSS.n246 5.2005
R628 VSS.n249 VSS.n248 5.2005
R629 VSS.n252 VSS.n251 5.2005
R630 VSS.n254 VSS.n253 5.2005
R631 VSS.n256 VSS.n255 5.2005
R632 VSS.n258 VSS.n257 5.2005
R633 VSS.n261 VSS.n260 5.2005
R634 VSS.n263 VSS.n262 5.2005
R635 VSS.n265 VSS.n264 5.2005
R636 VSS.n268 VSS.n267 5.2005
R637 VSS.n270 VSS.n269 5.2005
R638 VSS.n272 VSS.n271 5.2005
R639 VSS.n274 VSS.n273 5.2005
R640 VSS.n277 VSS.n276 5.2005
R641 VSS.n279 VSS.n278 5.2005
R642 VSS.n281 VSS.n280 5.2005
R643 VSS.n364 VSS.n287 5.2005
R644 VSS.n363 VSS.n288 5.2005
R645 VSS.n362 VSS.n289 5.2005
R646 VSS.n360 VSS.t42 5.2005
R647 VSS.n359 VSS.n292 5.2005
R648 VSS.n358 VSS.n293 5.2005
R649 VSS.n353 VSS.n351 5.2005
R650 VSS.n353 VSS.n352 5.2005
R651 VSS.n14 VSS.n10 5.2005
R652 VSS.n355 VSS.n348 5.00675
R653 VSS.n90 VSS.n89 4.5005
R654 VSS.n142 VSS.n141 4.5005
R655 VSS.n192 VSS.n191 4.5005
R656 VSS.n60 VSS.n59 4.5005
R657 VSS.n346 VSS.n345 4.5005
R658 VSS.n353 VSS.n349 4.5005
R659 VSS.n14 VSS.n13 4.5005
R660 VSS.n230 VSS.n131 3.76894
R661 VSS.n232 VSS.n231 3.72662
R662 VSS.n335 VSS.n297 3.65528
R663 VSS.n326 VSS.n299 3.65528
R664 VSS.n319 VSS.n301 3.65528
R665 VSS.n310 VSS.n303 3.65528
R666 VSS.n36 VSS.n35 3.65528
R667 VSS.n41 VSS.n30 3.65528
R668 VSS.n45 VSS.n25 3.65528
R669 VSS.n50 VSS.n19 3.65528
R670 VSS.n96 VSS.n83 3.6318
R671 VSS.n101 VSS.n81 3.6318
R672 VSS.n105 VSS.n79 3.6318
R673 VSS.n110 VSS.n77 3.6318
R674 VSS.n114 VSS.n75 3.6318
R675 VSS.n119 VSS.n73 3.6318
R676 VSS.n123 VSS.n71 3.6318
R677 VSS.n128 VSS.n69 3.6318
R678 VSS.n224 VSS.n147 3.62593
R679 VSS.n220 VSS.n152 3.62593
R680 VSS.n215 VSS.n157 3.62593
R681 VSS.n211 VSS.n162 3.62593
R682 VSS.n206 VSS.n168 3.62593
R683 VSS.n202 VSS.n173 3.62593
R684 VSS.n197 VSS.n179 3.62593
R685 VSS.n243 VSS.n9 3.61811
R686 VSS.n250 VSS.n7 3.61811
R687 VSS.n259 VSS.n5 3.61811
R688 VSS.n266 VSS.n3 3.61811
R689 VSS.n275 VSS.n1 3.61811
R690 VSS.n365 VSS.n286 3.61811
R691 VSS.n361 VSS.n291 3.61811
R692 VSS.n231 VSS.n230 3.26287
R693 VSS.n147 VSS.t116 2.7305
R694 VSS.n147 VSS.n146 2.7305
R695 VSS.n152 VSS.t138 2.7305
R696 VSS.n152 VSS.n151 2.7305
R697 VSS.n157 VSS.t152 2.7305
R698 VSS.n157 VSS.n156 2.7305
R699 VSS.n162 VSS.t143 2.7305
R700 VSS.n162 VSS.n161 2.7305
R701 VSS.n168 VSS.t126 2.7305
R702 VSS.n168 VSS.n167 2.7305
R703 VSS.n173 VSS.t115 2.7305
R704 VSS.n173 VSS.n172 2.7305
R705 VSS.n179 VSS.t137 2.7305
R706 VSS.n179 VSS.n178 2.7305
R707 VSS.n297 VSS.t51 2.7305
R708 VSS.n297 VSS.n296 2.7305
R709 VSS.n299 VSS.t54 2.7305
R710 VSS.n299 VSS.n298 2.7305
R711 VSS.n301 VSS.t44 2.7305
R712 VSS.n301 VSS.n300 2.7305
R713 VSS.n303 VSS.t63 2.7305
R714 VSS.n303 VSS.n302 2.7305
R715 VSS.n35 VSS.t62 2.7305
R716 VSS.n35 VSS.n34 2.7305
R717 VSS.n30 VSS.t21 2.7305
R718 VSS.n30 VSS.n29 2.7305
R719 VSS.n25 VSS.t39 2.7305
R720 VSS.n25 VSS.n24 2.7305
R721 VSS.n19 VSS.t10 2.7305
R722 VSS.n19 VSS.n18 2.7305
R723 VSS.n83 VSS.t134 2.7305
R724 VSS.n83 VSS.n82 2.7305
R725 VSS.n81 VSS.t124 2.7305
R726 VSS.n81 VSS.n80 2.7305
R727 VSS.n79 VSS.t132 2.7305
R728 VSS.n79 VSS.n78 2.7305
R729 VSS.n77 VSS.t123 2.7305
R730 VSS.n77 VSS.n76 2.7305
R731 VSS.n75 VSS.t129 2.7305
R732 VSS.n75 VSS.n74 2.7305
R733 VSS.n73 VSS.t151 2.7305
R734 VSS.n73 VSS.n72 2.7305
R735 VSS.n71 VSS.t125 2.7305
R736 VSS.n71 VSS.n70 2.7305
R737 VSS.n69 VSS.t133 2.7305
R738 VSS.n69 VSS.n68 2.7305
R739 VSS.n9 VSS.t55 2.7305
R740 VSS.n9 VSS.n8 2.7305
R741 VSS.n7 VSS.t66 2.7305
R742 VSS.n7 VSS.n6 2.7305
R743 VSS.n5 VSS.t41 2.7305
R744 VSS.n5 VSS.n4 2.7305
R745 VSS.n3 VSS.t60 2.7305
R746 VSS.n3 VSS.n2 2.7305
R747 VSS.n1 VSS.t32 2.7305
R748 VSS.n1 VSS.n0 2.7305
R749 VSS.n286 VSS.t15 2.7305
R750 VSS.n286 VSS.n285 2.7305
R751 VSS.n291 VSS.t159 2.7305
R752 VSS.n291 VSS.n290 2.7305
R753 VSS.n12 VSS.t16 2.67981
R754 VSS.n135 VSS.n134 2.63208
R755 VSS.n341 VSS.n340 2.60175
R756 VSS.n137 VSS.n136 2.60175
R757 VSS.n185 VSS.n184 2.60175
R758 VSS.n64 VSS.n62 2.60175
R759 VSS.n235 VSS.n234 2.60175
R760 VSS.n356 VSS.n295 2.60175
R761 VSS.n55 VSS.n54 2.60175
R762 VSS.n295 VSS.n294 2.601
R763 VSS.n54 VSS.n53 2.601
R764 VSS.n340 VSS.n339 2.601
R765 VSS.n136 VSS.n135 2.601
R766 VSS.n234 VSS.n233 2.601
R767 VSS VSS.n284 2.6005
R768 VSS.n284 VSS.n283 2.6005
R769 VSS.n348 VSS.n347 2.55463
R770 VSS.n61 VSS.n60 2.41795
R771 VSS.n347 VSS.n346 2.41733
R772 VSS.n354 VSS.n353 2.41463
R773 VSS.n193 VSS.n192 2.40822
R774 VSS.n16 VSS.n14 2.40807
R775 VSS.n228 VSS.n142 2.4075
R776 VSS.n130 VSS.n67 2.40736
R777 VSS.n231 VSS.n61 2.26028
R778 VSS.n187 VSS.n186 2.25438
R779 VSS.n230 VSS.n229 2.25101
R780 VSS.n64 VSS.n63 2.21822
R781 VSS.n86 VSS.n85 2.0261
R782 VSS.n92 VSS.n88 1.88512
R783 VSS.n192 VSS.n189 1.87311
R784 VSS.n142 VSS.n139 1.82853
R785 VSS.n60 VSS.n57 1.78394
R786 VSS.n346 VSS.n343 1.78394
R787 VSS.n92 VSS.n91 1.73383
R788 VSS.n93 VSS.n92 1.73383
R789 VSS.n353 VSS.n350 1.6056
R790 VSS.n14 VSS.n11 1.6056
R791 VSS.n284 VSS.n282 0.312602
R792 VSS.n227 VSS.n226 0.133192
R793 VSS.n226 VSS.n225 0.133192
R794 VSS.n223 VSS.n222 0.133192
R795 VSS.n222 VSS.n221 0.133192
R796 VSS.n219 VSS.n218 0.133192
R797 VSS.n218 VSS.n217 0.133192
R798 VSS.n217 VSS.n216 0.133192
R799 VSS.n214 VSS.n213 0.133192
R800 VSS.n213 VSS.n212 0.133192
R801 VSS.n210 VSS.n209 0.133192
R802 VSS.n209 VSS.n208 0.133192
R803 VSS.n208 VSS.n207 0.133192
R804 VSS.n205 VSS.n204 0.133192
R805 VSS.n204 VSS.n203 0.133192
R806 VSS.n201 VSS.n200 0.133192
R807 VSS.n200 VSS.n199 0.133192
R808 VSS.n199 VSS.n198 0.133192
R809 VSS.n196 VSS.n195 0.133192
R810 VSS.n195 VSS.n194 0.133192
R811 VSS.n49 VSS.n48 0.133192
R812 VSS.n48 VSS.n47 0.133192
R813 VSS.n47 VSS.n46 0.133192
R814 VSS.n44 VSS.n43 0.133192
R815 VSS.n43 VSS.n42 0.133192
R816 VSS.n40 VSS.n39 0.133192
R817 VSS.n39 VSS.n38 0.133192
R818 VSS.n38 VSS.n37 0.133192
R819 VSS.n307 VSS.n305 0.133192
R820 VSS.n309 VSS.n307 0.133192
R821 VSS.n314 VSS.n312 0.133192
R822 VSS.n316 VSS.n314 0.133192
R823 VSS.n318 VSS.n316 0.133192
R824 VSS.n323 VSS.n321 0.133192
R825 VSS.n325 VSS.n323 0.133192
R826 VSS.n330 VSS.n328 0.133192
R827 VSS.n332 VSS.n330 0.133192
R828 VSS.n334 VSS.n332 0.133192
R829 VSS.n127 VSS.n126 0.133192
R830 VSS.n126 VSS.n125 0.133192
R831 VSS.n125 VSS.n124 0.133192
R832 VSS.n122 VSS.n121 0.133192
R833 VSS.n121 VSS.n120 0.133192
R834 VSS.n118 VSS.n117 0.133192
R835 VSS.n117 VSS.n116 0.133192
R836 VSS.n116 VSS.n115 0.133192
R837 VSS.n113 VSS.n112 0.133192
R838 VSS.n112 VSS.n111 0.133192
R839 VSS.n109 VSS.n108 0.133192
R840 VSS.n108 VSS.n107 0.133192
R841 VSS.n107 VSS.n106 0.133192
R842 VSS.n104 VSS.n103 0.133192
R843 VSS.n103 VSS.n102 0.133192
R844 VSS.n100 VSS.n99 0.133192
R845 VSS.n99 VSS.n98 0.133192
R846 VSS.n98 VSS.n97 0.133192
R847 VSS.n240 VSS.n238 0.133192
R848 VSS.n242 VSS.n240 0.133192
R849 VSS.n247 VSS.n245 0.133192
R850 VSS.n249 VSS.n247 0.133192
R851 VSS.n254 VSS.n252 0.133192
R852 VSS.n256 VSS.n254 0.133192
R853 VSS.n258 VSS.n256 0.133192
R854 VSS.n263 VSS.n261 0.133192
R855 VSS.n265 VSS.n263 0.133192
R856 VSS.n270 VSS.n268 0.133192
R857 VSS.n272 VSS.n270 0.133192
R858 VSS.n274 VSS.n272 0.133192
R859 VSS.n279 VSS.n277 0.133192
R860 VSS.n281 VSS.n279 0.133192
R861 VSS VSS.n281 0.133192
R862 VSS.n364 VSS.n363 0.133192
R863 VSS.n363 VSS.n362 0.133192
R864 VSS.n360 VSS.n359 0.133192
R865 VSS.n359 VSS.n358 0.133192
R866 VSS.n45 VSS.n44 0.132038
R867 VSS.n123 VSS.n122 0.132038
R868 VSS.n365 VSS.n364 0.132038
R869 VSS.n203 VSS.n202 0.129731
R870 VSS.n130 VSS.n129 0.121842
R871 VSS.n266 VSS.n265 0.121654
R872 VSS.n228 VSS.n227 0.120957
R873 VSS.n114 VSS.n113 0.119346
R874 VSS.n212 VSS.n211 0.117038
R875 VSS.n194 VSS.n193 0.116533
R876 VSS.n338 VSS.n337 0.112423
R877 VSS.n358 VSS.n357 0.112423
R878 VSS.n238 VSS.n236 0.111846
R879 VSS.n52 VSS.n51 0.109538
R880 VSS.n95 VSS.n94 0.108962
R881 VSS.n250 VSS.n249 0.108962
R882 VSS.n321 VSS.n319 0.106654
R883 VSS.n105 VSS.n104 0.106654
R884 VSS.n221 VSS.n220 0.104346
R885 VSS.n224 VSS.n223 0.102038
R886 VSS.n326 VSS.n325 0.0997308
R887 VSS.n102 VSS.n101 0.0997308
R888 VSS.n245 VSS.n243 0.0974231
R889 VSS.n337 VSS.n335 0.0939615
R890 VSS.n96 VSS.n95 0.0939615
R891 VSS.n92 VSS.n90 0.0902436
R892 VSS.n215 VSS.n214 0.0893462
R893 VSS.n310 VSS.n309 0.0870385
R894 VSS.n111 VSS.n110 0.0870385
R895 VSS.n261 VSS.n259 0.0847308
R896 VSS.n206 VSS.n205 0.0766538
R897 VSS.n42 VSS.n41 0.0743462
R898 VSS.n120 VSS.n119 0.0743462
R899 VSS.n362 VSS.n361 0.0743462
R900 VSS.n50 VSS.n49 0.0720385
R901 VSS.n128 VSS.n127 0.0720385
R902 VSS.n277 VSS.n275 0.0720385
R903 VSS.n198 VSS.n197 0.0697308
R904 VSS.n197 VSS.n196 0.0639615
R905 VSS.n51 VSS.n50 0.0616538
R906 VSS.n129 VSS.n128 0.0616538
R907 VSS.n275 VSS.n274 0.0616538
R908 VSS.n41 VSS.n40 0.0593462
R909 VSS.n119 VSS.n118 0.0593462
R910 VSS.n361 VSS.n360 0.0593462
R911 VSS.n207 VSS.n206 0.0570385
R912 VSS.n259 VSS.n258 0.0489615
R913 VSS.n312 VSS.n310 0.0466538
R914 VSS.n110 VSS.n109 0.0466538
R915 VSS.n216 VSS.n215 0.0443462
R916 VSS.n335 VSS.n334 0.0397308
R917 VSS.n97 VSS.n96 0.0397308
R918 VSS.n243 VSS.n242 0.0362692
R919 VSS.n328 VSS.n326 0.0339615
R920 VSS.n101 VSS.n100 0.0339615
R921 VSS.n225 VSS.n224 0.0316538
R922 VSS.n220 VSS.n219 0.0293462
R923 VSS.n319 VSS.n318 0.0270385
R924 VSS.n106 VSS.n105 0.0270385
R925 VSS.n94 VSS.n93 0.0247308
R926 VSS.n252 VSS.n250 0.0247308
R927 VSS.n137 VSS.n133 0.0241538
R928 VSS.n55 VSS.n52 0.0241538
R929 VSS.n236 VSS.n235 0.0218462
R930 VSS.n341 VSS.n338 0.0212692
R931 VSS.n357 VSS.n356 0.0212692
R932 VSS.n211 VSS.n210 0.0166538
R933 VSS.n37 VSS.n36 0.0143462
R934 VSS.n115 VSS.n114 0.0143462
R935 VSS.n131 VSS.n130 0.0122131
R936 VSS.n268 VSS.n266 0.0120385
R937 VSS.n229 VSS.n228 0.0119467
R938 VSS.n232 VSS.n16 0.0108811
R939 VSS.n193 VSS.n187 0.0106146
R940 VSS.n185 VSS.n183 0.00973077
R941 VSS.n187 VSS.n185 0.008
R942 VSS.n347 VSS.n341 0.008
R943 VSS.n356 VSS.n355 0.00742308
R944 VSS.n235 VSS.n232 0.00684615
R945 VSS.n355 VSS.n354 0.00420487
R946 VSS.n202 VSS.n201 0.00396154
R947 VSS.n229 VSS.n137 0.00223077
R948 VSS.n61 VSS.n55 0.00165385
R949 VSS.n46 VSS.n45 0.00165385
R950 VSS.n124 VSS.n123 0.00165385
R951 VSS.n93 VSS.n86 0.00165385
R952 VSS VSS.n365 0.00165385
R953 VSS.n131 VSS.n64 0.00107692
R954 G1_2.n9 G1_2.t141 110.841
R955 G1_2.n137 G1_2.t36 104.368
R956 G1_2.n11 G1_2.n10 98.3584
R957 G1_2.n13 G1_2.n12 98.3584
R958 G1_2.n15 G1_2.n14 98.3584
R959 G1_2.n17 G1_2.n16 98.3584
R960 G1_2.n19 G1_2.n18 98.3584
R961 G1_2.n21 G1_2.n20 98.3584
R962 G1_2.n30 G1_2.n29 98.3584
R963 G1_2.n28 G1_2.n27 98.3584
R964 G1_2.n26 G1_2.n25 98.3584
R965 G1_2.n144 G1_2.n143 98.3584
R966 G1_2.n146 G1_2.n145 98.3584
R967 G1_2.n148 G1_2.n147 98.3584
R968 G1_2.n23 G1_2.n22 91.8697
R969 G1_2.n163 G1_2.n162 89.3295
R970 G1_2.n195 G1_2.t46 50.286
R971 G1_2.n166 G1_2.n165 39.19
R972 G1_2.n120 G1_2.n119 39.19
R973 G1_2.n102 G1_2.n101 39.19
R974 G1_2.n84 G1_2.n83 39.19
R975 G1_2.n66 G1_2.n65 39.19
R976 G1_2.n48 G1_2.n47 39.19
R977 G1_2.n162 G1_2.t16 32.4624
R978 G1_2.n108 G1_2.n107 21.3797
R979 G1_2.n54 G1_2.n53 21.3765
R980 G1_2.n90 G1_2.n89 21.3729
R981 G1_2.n126 G1_2.n125 21.3689
R982 G1_2.n72 G1_2.n71 21.2844
R983 G1_2.n149 G1_2.n148 21.2613
R984 G1_2.n31 G1_2.n30 20.7384
R985 G1_2.n10 G1_2.n9 19.9794
R986 G1_2.n12 G1_2.n11 19.9794
R987 G1_2.n14 G1_2.n13 19.9794
R988 G1_2.n16 G1_2.n15 19.9794
R989 G1_2.n18 G1_2.n17 19.9794
R990 G1_2.n20 G1_2.n19 19.9794
R991 G1_2.n22 G1_2.n21 19.9794
R992 G1_2.n29 G1_2.n28 19.9794
R993 G1_2.n27 G1_2.n26 19.9794
R994 G1_2.n25 G1_2.n24 19.9794
R995 G1_2.n143 G1_2.n142 19.9794
R996 G1_2.n145 G1_2.n144 19.9794
R997 G1_2.n147 G1_2.n146 19.9794
R998 G1_2.n136 G1_2.n135 19.9794
R999 G1_2.n5 G1_2.n4 19.9794
R1000 G1_2.n9 G1_2.t137 12.4835
R1001 G1_2.n10 G1_2.t113 12.4835
R1002 G1_2.n11 G1_2.t108 12.4835
R1003 G1_2.n12 G1_2.t125 12.4835
R1004 G1_2.n13 G1_2.t134 12.4835
R1005 G1_2.n14 G1_2.t97 12.4835
R1006 G1_2.n15 G1_2.t100 12.4835
R1007 G1_2.n16 G1_2.t123 12.4835
R1008 G1_2.n17 G1_2.t119 12.4835
R1009 G1_2.n18 G1_2.t129 12.4835
R1010 G1_2.n19 G1_2.t138 12.4835
R1011 G1_2.n20 G1_2.t114 12.4835
R1012 G1_2.n21 G1_2.t128 12.4835
R1013 G1_2.n22 G1_2.t140 12.4835
R1014 G1_2.n30 G1_2.t106 12.4835
R1015 G1_2.n29 G1_2.t142 12.4835
R1016 G1_2.n28 G1_2.t117 12.4835
R1017 G1_2.n27 G1_2.t104 12.4835
R1018 G1_2.n26 G1_2.t98 12.4835
R1019 G1_2.n25 G1_2.t130 12.4835
R1020 G1_2.n24 G1_2.t120 12.4835
R1021 G1_2.n142 G1_2.t124 12.4835
R1022 G1_2.n143 G1_2.t101 12.4835
R1023 G1_2.n144 G1_2.t103 12.4835
R1024 G1_2.n145 G1_2.t135 12.4835
R1025 G1_2.n146 G1_2.t139 12.4835
R1026 G1_2.n147 G1_2.t116 12.4835
R1027 G1_2.n148 G1_2.t115 12.4835
R1028 G1_2.n135 G1_2.t24 12.4835
R1029 G1_2.n125 G1_2.t48 12.4835
R1030 G1_2.n107 G1_2.t34 12.4835
R1031 G1_2.n89 G1_2.t50 12.4835
R1032 G1_2.n71 G1_2.t42 12.4835
R1033 G1_2.n53 G1_2.t22 12.4835
R1034 G1_2.n4 G1_2.t38 12.4835
R1035 G1_2.n162 G1_2.t20 12.4835
R1036 G1_2.n23 G1_2.t136 12.0283
R1037 G1_2.n181 G1_2.t64 11.7766
R1038 G1_2.n31 G1_2.t121 11.6536
R1039 G1_2.n7 G1_2.t10 11.2425
R1040 G1_2.n72 G1_2.t66 11.0965
R1041 G1_2.n165 G1_2.t32 11.0965
R1042 G1_2.n119 G1_2.t28 11.0965
R1043 G1_2.n101 G1_2.t44 11.0965
R1044 G1_2.n83 G1_2.t40 11.0965
R1045 G1_2.n65 G1_2.t26 11.0965
R1046 G1_2.n47 G1_2.t30 11.0965
R1047 G1_2.n149 G1_2.t107 11.0781
R1048 G1_2.n126 G1_2.t52 11.0235
R1049 G1_2.n108 G1_2.t58 11.0235
R1050 G1_2.n90 G1_2.t54 11.0235
R1051 G1_2.n54 G1_2.t60 11.0235
R1052 G1_2.n195 G1_2.n194 10.5803
R1053 G1_2.n138 G1_2.t56 9.7825
R1054 G1_2.n193 G1_2.t6 9.4175
R1055 G1_2.n46 G1_2.t14 9.4175
R1056 G1_2.n64 G1_2.t68 9.3445
R1057 G1_2.n100 G1_2.t18 9.2715
R1058 G1_2.n82 G1_2.t8 9.2715
R1059 G1_2.n164 G1_2.t12 9.1985
R1060 G1_2.n118 G1_2.t62 9.1985
R1061 G1_2.n164 G1_2.n163 6.91629
R1062 G1_2.n64 G1_2.n63 6.67631
R1063 G1_2.n150 G1_2.n149 6.39681
R1064 G1_2.n32 G1_2.n31 6.38115
R1065 G1_2.n194 G1_2.n193 6.29484
R1066 G1_2.n100 G1_2.n99 5.98304
R1067 G1_2.n118 G1_2.n117 5.73461
R1068 G1_2.n82 G1_2.n81 5.57314
R1069 G1_2.n32 G1_2.n23 5.25845
R1070 G1_2.n68 G1_2.n67 5.13202
R1071 G1_2.n104 G1_2.n103 4.86134
R1072 G1_2.n122 G1_2.n121 4.85769
R1073 G1_2.n50 G1_2.n49 4.77802
R1074 G1_2.n86 G1_2.n85 4.77215
R1075 G1_2.n168 G1_2.n167 4.67852
R1076 G1_2.n46 G1_2.n45 4.53834
R1077 G1_2.n112 G1_2.n109 4.52266
R1078 G1_2.n76 G1_2.n73 4.43719
R1079 G1_2.n58 G1_2.n55 4.43328
R1080 G1_2.n130 G1_2.n127 4.36026
R1081 G1_2.n184 G1_2.n181 4.28703
R1082 G1_2.n94 G1_2.n91 4.27334
R1083 G1_2.n197 G1_2.n196 4.0005
R1084 G1_2.n139 G1_2.n137 3.53989
R1085 G1_2.n158 G1_2.n157 3.1855
R1086 G1_2.n159 G1_2.n134 3.1855
R1087 G1_2.n170 G1_2.n124 3.1855
R1088 G1_2.n172 G1_2.n106 3.1855
R1089 G1_2.n174 G1_2.n88 3.1855
R1090 G1_2.n176 G1_2.n70 3.1855
R1091 G1_2.n178 G1_2.n52 3.1855
R1092 G1_2.n180 G1_2.n3 3.1855
R1093 G1_2.n187 G1_2.n186 3.1855
R1094 G1_2.n7 G1_2.n6 3.15726
R1095 G1_2.n161 G1_2.t74 3.03383
R1096 G1_2.n161 G1_2.n160 3.03383
R1097 G1_2.n132 G1_2.t25 3.03383
R1098 G1_2.n132 G1_2.n131 3.03383
R1099 G1_2.n157 G1_2.t94 3.03383
R1100 G1_2.n157 G1_2.n156 3.03383
R1101 G1_2.n155 G1_2.t37 3.03383
R1102 G1_2.n155 G1_2.n154 3.03383
R1103 G1_2.n134 G1_2.t21 3.03383
R1104 G1_2.n134 G1_2.n133 3.03383
R1105 G1_2.n124 G1_2.t33 3.03383
R1106 G1_2.n124 G1_2.n123 3.03383
R1107 G1_2.n116 G1_2.t76 3.03383
R1108 G1_2.n116 G1_2.n115 3.03383
R1109 G1_2.n114 G1_2.t49 3.03383
R1110 G1_2.n114 G1_2.n113 3.03383
R1111 G1_2.n106 G1_2.t29 3.03383
R1112 G1_2.n106 G1_2.n105 3.03383
R1113 G1_2.n98 G1_2.t93 3.03383
R1114 G1_2.n98 G1_2.n97 3.03383
R1115 G1_2.n96 G1_2.t35 3.03383
R1116 G1_2.n96 G1_2.n95 3.03383
R1117 G1_2.n88 G1_2.t45 3.03383
R1118 G1_2.n88 G1_2.n87 3.03383
R1119 G1_2.n80 G1_2.t77 3.03383
R1120 G1_2.n80 G1_2.n79 3.03383
R1121 G1_2.n78 G1_2.t51 3.03383
R1122 G1_2.n78 G1_2.n77 3.03383
R1123 G1_2.n70 G1_2.t41 3.03383
R1124 G1_2.n70 G1_2.n69 3.03383
R1125 G1_2.n62 G1_2.t92 3.03383
R1126 G1_2.n62 G1_2.n61 3.03383
R1127 G1_2.n60 G1_2.t43 3.03383
R1128 G1_2.n60 G1_2.n59 3.03383
R1129 G1_2.n52 G1_2.t27 3.03383
R1130 G1_2.n52 G1_2.n51 3.03383
R1131 G1_2.n44 G1_2.t73 3.03383
R1132 G1_2.n44 G1_2.n43 3.03383
R1133 G1_2.n42 G1_2.t23 3.03383
R1134 G1_2.n42 G1_2.n41 3.03383
R1135 G1_2.n3 G1_2.t31 3.03383
R1136 G1_2.n3 G1_2.n2 3.03383
R1137 G1_2.n190 G1_2.t95 3.03383
R1138 G1_2.n190 G1_2.n189 3.03383
R1139 G1_2.n1 G1_2.t39 3.03383
R1140 G1_2.n1 G1_2.n0 3.03383
R1141 G1_2.n186 G1_2.t47 3.03383
R1142 G1_2.n186 G1_2.n185 3.03383
R1143 G1_2.n183 G1_2.t4 3.03383
R1144 G1_2.n183 G1_2.n182 3.03383
R1145 G1_2.n57 G1_2.t78 3.03383
R1146 G1_2.n57 G1_2.n56 3.03383
R1147 G1_2.n75 G1_2.t87 3.03383
R1148 G1_2.n75 G1_2.n74 3.03383
R1149 G1_2.n93 G1_2.t89 3.03383
R1150 G1_2.n93 G1_2.n92 3.03383
R1151 G1_2.n111 G1_2.t80 3.03383
R1152 G1_2.n111 G1_2.n110 3.03383
R1153 G1_2.n129 G1_2.t82 3.03383
R1154 G1_2.n129 G1_2.n128 3.03383
R1155 G1_2.n39 G1_2.t86 3.03383
R1156 G1_2.n39 G1_2.n38 3.03383
R1157 G1_2.n152 G1_2.t91 3.03383
R1158 G1_2.n152 G1_2.n151 3.03383
R1159 G1_2.n35 G1_2.n8 2.88206
R1160 G1_2.n141 G1_2.n140 2.84775
R1161 G1_2.n169 G1_2.n132 2.84507
R1162 G1_2.n158 G1_2.n155 2.84507
R1163 G1_2.n171 G1_2.n114 2.84507
R1164 G1_2.n173 G1_2.n96 2.84507
R1165 G1_2.n175 G1_2.n78 2.84507
R1166 G1_2.n177 G1_2.n60 2.84507
R1167 G1_2.n179 G1_2.n42 2.84507
R1168 G1_2.n188 G1_2.n1 2.84507
R1169 G1_2.n122 G1_2.n116 2.6005
R1170 G1_2.n104 G1_2.n98 2.6005
R1171 G1_2.n86 G1_2.n80 2.6005
R1172 G1_2.n68 G1_2.n62 2.6005
R1173 G1_2.n50 G1_2.n44 2.6005
R1174 G1_2.n191 G1_2.n190 2.6005
R1175 G1_2.n58 G1_2.n57 2.6005
R1176 G1_2.n76 G1_2.n75 2.6005
R1177 G1_2.n94 G1_2.n93 2.6005
R1178 G1_2.n112 G1_2.n111 2.6005
R1179 G1_2.n130 G1_2.n129 2.6005
R1180 G1_2.n40 G1_2.n39 2.6005
R1181 G1_2.n153 G1_2.n152 2.6005
R1182 G1_2.n184 G1_2.n183 2.6005
R1183 G1_2.n168 G1_2.n161 2.6005
R1184 G1_2.n33 G1_2.n32 1.65279
R1185 G1_2.n139 G1_2.n138 1.4605
R1186 G1_2.n49 G1_2.n46 1.3145
R1187 G1_2.n103 G1_2.n100 1.2415
R1188 G1_2.n85 G1_2.n82 1.2415
R1189 G1_2.n67 G1_2.n64 1.2415
R1190 G1_2.n167 G1_2.n164 1.1685
R1191 G1_2.n121 G1_2.n118 1.1685
R1192 G1_2.n193 G1_2.n192 1.1685
R1193 G1_2.n35 G1_2.n34 1.13001
R1194 G1_2.n153 G1_2.n150 1.01243
R1195 G1_2.n197 G1_2.n191 1.00561
R1196 G1_2.n8 G1_2.n5 0.8765
R1197 G1_2.n40 G1_2.n37 0.804097
R1198 G1_2.n140 G1_2.n136 0.782953
R1199 G1_2.n167 G1_2.n166 0.7305
R1200 G1_2.n121 G1_2.n120 0.7305
R1201 G1_2.n127 G1_2.n126 0.712695
R1202 G1_2.n171 G1_2.n122 0.5855
R1203 G1_2.n173 G1_2.n104 0.5855
R1204 G1_2.n175 G1_2.n86 0.5855
R1205 G1_2.n177 G1_2.n68 0.5855
R1206 G1_2.n179 G1_2.n50 0.5855
R1207 G1_2.n191 G1_2.n188 0.5855
R1208 G1_2.n169 G1_2.n168 0.5855
R1209 G1_2.n103 G1_2.n102 0.5845
R1210 G1_2.n85 G1_2.n84 0.5845
R1211 G1_2.n91 G1_2.n90 0.534646
R1212 G1_2.n67 G1_2.n66 0.5115
R1213 G1_2.n140 G1_2.n139 0.458361
R1214 G1_2.n159 G1_2.n158 0.44291
R1215 G1_2.n169 G1_2.n159 0.44291
R1216 G1_2.n170 G1_2.n169 0.44291
R1217 G1_2.n171 G1_2.n170 0.44291
R1218 G1_2.n172 G1_2.n171 0.44291
R1219 G1_2.n173 G1_2.n172 0.44291
R1220 G1_2.n174 G1_2.n173 0.44291
R1221 G1_2.n175 G1_2.n174 0.44291
R1222 G1_2.n176 G1_2.n175 0.44291
R1223 G1_2.n177 G1_2.n176 0.44291
R1224 G1_2.n178 G1_2.n177 0.44291
R1225 G1_2.n179 G1_2.n178 0.44291
R1226 G1_2.n180 G1_2.n179 0.44291
R1227 G1_2.n188 G1_2.n180 0.44291
R1228 G1_2.n188 G1_2.n187 0.44291
R1229 G1_2.n8 G1_2.n7 0.3655
R1230 G1_2.n49 G1_2.n48 0.3655
R1231 G1_2.n196 G1_2.n195 0.3655
R1232 G1_2.n73 G1_2.n72 0.267573
R1233 G1_2.n55 G1_2.n54 0.267573
R1234 G1_2.n178 G1_2.n58 0.245065
R1235 G1_2.n176 G1_2.n76 0.245065
R1236 G1_2.n174 G1_2.n94 0.245065
R1237 G1_2.n172 G1_2.n112 0.245065
R1238 G1_2.n170 G1_2.n130 0.245065
R1239 G1_2.n180 G1_2.n40 0.245065
R1240 G1_2.n159 G1_2.n153 0.245065
R1241 G1_2.n187 G1_2.n184 0.245065
R1242 G1_2.n196 G1_2.n192 0.1465
R1243 G1_2.n109 G1_2.n108 0.0895244
R1244 G1_2.n34 G1_2.n33 0.0332273
R1245 G1_2.n36 G1_2.n35 0.0241243
R1246 G1_2.n37 G1_2.n36 0.0141364
R1247 G1_2.n150 G1_2.n141 0.0133843
R1248 G1_2 G1_2.n197 0.0123033
R1249 VDD.n255 VDD.t32 42.5052
R1250 VDD.n91 VDD.t5 40.9872
R1251 VDD.n73 VDD.t89 39.4692
R1252 VDD.n73 VDD.t25 37.9512
R1253 VDD.n91 VDD.t73 36.4331
R1254 VDD.n255 VDD.t17 34.9151
R1255 VDD.n107 VDD.t45 32.6381
R1256 VDD.n88 VDD.t52 31.12
R1257 VDD.n70 VDD.t29 29.602
R1258 VDD.n75 VDD.t43 28.084
R1259 VDD.n93 VDD.t66 26.566
R1260 VDD.n109 VDD.t87 25.0479
R1261 VDD.n104 VDD.t59 22.7709
R1262 VDD.n86 VDD.t6 21.2529
R1263 VDD.n68 VDD.t7 19.7348
R1264 VDD.n77 VDD.t61 18.2168
R1265 VDD.n95 VDD.t10 16.6988
R1266 VDD.n118 VDD.t9 15.9398
R1267 VDD.n112 VDD.t15 15.1808
R1268 VDD.n115 VDD.t41 14.4218
R1269 VDD.n102 VDD.t1 12.9037
R1270 VDD.n84 VDD.t38 11.3857
R1271 VDD.n129 VDD.t8 10.6267
R1272 VDD.n66 VDD.t2 9.86767
R1273 VDD.n18 VDD.n14 9.71606
R1274 VDD.n79 VDD.t36 8.34965
R1275 VDD.n98 VDD.t48 6.83162
R1276 VDD.n243 VDD.n135 6.37537
R1277 VDD.n130 VDD.n129 6.3005
R1278 VDD.n18 VDD.n16 6.3005
R1279 VDD.n64 VDD.t3 6.3005
R1280 VDD.n67 VDD.n66 6.3005
R1281 VDD.n69 VDD.n68 6.3005
R1282 VDD.n71 VDD.n70 6.3005
R1283 VDD.n74 VDD.n73 6.3005
R1284 VDD.n76 VDD.n75 6.3005
R1285 VDD.n78 VDD.n77 6.3005
R1286 VDD.n80 VDD.n79 6.3005
R1287 VDD.n83 VDD.n82 6.3005
R1288 VDD.n85 VDD.n84 6.3005
R1289 VDD.n87 VDD.n86 6.3005
R1290 VDD.n89 VDD.n88 6.3005
R1291 VDD.n92 VDD.n91 6.3005
R1292 VDD.n94 VDD.n93 6.3005
R1293 VDD.n96 VDD.n95 6.3005
R1294 VDD.n99 VDD.n98 6.3005
R1295 VDD.n101 VDD.n100 6.3005
R1296 VDD.n103 VDD.n102 6.3005
R1297 VDD.n105 VDD.n104 6.3005
R1298 VDD.n108 VDD.n107 6.3005
R1299 VDD.n253 VDD.n109 6.3005
R1300 VDD.n251 VDD.n112 6.3005
R1301 VDD.n250 VDD.n113 6.3005
R1302 VDD.n249 VDD.n114 6.3005
R1303 VDD.n248 VDD.n115 6.3005
R1304 VDD.n123 VDD.n119 6.3005
R1305 VDD.n51 VDD.n38 6.13519
R1306 VDD.n37 VDD.n36 6.1324
R1307 VDD.n200 VDD.t98 6.12266
R1308 VDD.n238 VDD.t35 6.11709
R1309 VDD.n16 VDD.n15 6.07261
R1310 VDD.n113 VDD.t0 5.31359
R1311 VDD.n241 VDD.n240 4.85382
R1312 VDD.n53 VDD.n52 4.68801
R1313 VDD.n114 VDD.t20 4.55458
R1314 VDD.n132 VDD.n131 4.5005
R1315 VDD.n123 VDD.n122 4.5005
R1316 VDD.n18 VDD.n17 4.5005
R1317 VDD.n243 VDD.n242 4.2252
R1318 VDD.n52 VDD.n37 4.08027
R1319 VDD.n47 VDD.n40 3.15224
R1320 VDD.n162 VDD.n161 3.15224
R1321 VDD.n168 VDD.n157 3.15224
R1322 VDD.n174 VDD.n153 3.15224
R1323 VDD.n179 VDD.n149 3.15224
R1324 VDD.n185 VDD.n145 3.15224
R1325 VDD.n190 VDD.n141 3.15224
R1326 VDD.n196 VDD.n137 3.15224
R1327 VDD.n61 VDD.n60 3.15175
R1328 VDD.n245 VDD.n128 3.15175
R1329 VDD.n62 VDD.n61 3.151
R1330 VDD.n60 VDD.n59 3.151
R1331 VDD.n60 VDD.n56 3.151
R1332 VDD.n128 VDD.n127 3.151
R1333 VDD.n127 VDD.n126 3.151
R1334 VDD.n257 VDD.n256 3.1505
R1335 VDD.n256 VDD.n255 3.1505
R1336 VDD.n193 VDD.n139 3.08376
R1337 VDD.n187 VDD.n143 3.08376
R1338 VDD.n182 VDD.n147 3.08376
R1339 VDD.n176 VDD.n151 3.08376
R1340 VDD.n171 VDD.n155 3.08376
R1341 VDD.n165 VDD.n159 3.08376
R1342 VDD.n44 VDD.n42 3.08376
R1343 VDD.n233 VDD.n204 3.08376
R1344 VDD.n228 VDD.n206 3.08376
R1345 VDD.n224 VDD.n208 3.08376
R1346 VDD.n219 VDD.n210 3.08376
R1347 VDD.n215 VDD.n212 3.08376
R1348 VDD.n25 VDD.n22 3.08376
R1349 VDD.n29 VDD.n20 3.08376
R1350 VDD.n65 VDD.n11 3.05441
R1351 VDD.n72 VDD.n9 3.05441
R1352 VDD.n81 VDD.n7 3.05441
R1353 VDD.n90 VDD.n5 3.05441
R1354 VDD.n97 VDD.n3 3.05441
R1355 VDD.n106 VDD.n1 3.05441
R1356 VDD.n252 VDD.n111 3.05441
R1357 VDD.n247 VDD.n117 3.05441
R1358 VDD.n100 VDD.t13 3.03655
R1359 VDD.n40 VDD.t103 3.03383
R1360 VDD.n40 VDD.n39 3.03383
R1361 VDD.n161 VDD.t90 3.03383
R1362 VDD.n161 VDD.n160 3.03383
R1363 VDD.n157 VDD.t37 3.03383
R1364 VDD.n157 VDD.n156 3.03383
R1365 VDD.n153 VDD.t119 3.03383
R1366 VDD.n153 VDD.n152 3.03383
R1367 VDD.n149 VDD.t79 3.03383
R1368 VDD.n149 VDD.n148 3.03383
R1369 VDD.n145 VDD.t124 3.03383
R1370 VDD.n145 VDD.n144 3.03383
R1371 VDD.n141 VDD.t88 3.03383
R1372 VDD.n141 VDD.n140 3.03383
R1373 VDD.n137 VDD.t104 3.03383
R1374 VDD.n137 VDD.n136 3.03383
R1375 VDD.n139 VDD.t107 3.03383
R1376 VDD.n139 VDD.n138 3.03383
R1377 VDD.n143 VDD.t96 3.03383
R1378 VDD.n143 VDD.n142 3.03383
R1379 VDD.n147 VDD.t14 3.03383
R1380 VDD.n147 VDD.n146 3.03383
R1381 VDD.n151 VDD.t74 3.03383
R1382 VDD.n151 VDD.n150 3.03383
R1383 VDD.n155 VDD.t99 3.03383
R1384 VDD.n155 VDD.n154 3.03383
R1385 VDD.n159 VDD.t44 3.03383
R1386 VDD.n159 VDD.n158 3.03383
R1387 VDD.n42 VDD.t97 3.03383
R1388 VDD.n42 VDD.n41 3.03383
R1389 VDD.n204 VDD.t57 3.03383
R1390 VDD.n204 VDD.n203 3.03383
R1391 VDD.n206 VDD.t33 3.03383
R1392 VDD.n206 VDD.n205 3.03383
R1393 VDD.n208 VDD.t80 3.03383
R1394 VDD.n208 VDD.n207 3.03383
R1395 VDD.n210 VDD.t122 3.03383
R1396 VDD.n210 VDD.n209 3.03383
R1397 VDD.n212 VDD.t39 3.03383
R1398 VDD.n212 VDD.n211 3.03383
R1399 VDD.n22 VDD.t100 3.03383
R1400 VDD.n22 VDD.n21 3.03383
R1401 VDD.n20 VDD.t34 3.03383
R1402 VDD.n20 VDD.n19 3.03383
R1403 VDD.n11 VDD.t40 3.03383
R1404 VDD.n11 VDD.n10 3.03383
R1405 VDD.n9 VDD.t127 3.03383
R1406 VDD.n9 VDD.n8 3.03383
R1407 VDD.n7 VDD.t84 3.03383
R1408 VDD.n7 VDD.n6 3.03383
R1409 VDD.n5 VDD.t53 3.03383
R1410 VDD.n5 VDD.n4 3.03383
R1411 VDD.n3 VDD.t116 3.03383
R1412 VDD.n3 VDD.n2 3.03383
R1413 VDD.n1 VDD.t60 3.03383
R1414 VDD.n1 VDD.n0 3.03383
R1415 VDD.n111 VDD.t123 3.03383
R1416 VDD.n111 VDD.n110 3.03383
R1417 VDD.n117 VDD.t42 3.03383
R1418 VDD.n117 VDD.n116 3.03383
R1419 VDD.n53 VDD.n18 2.62871
R1420 VDD.n119 VDD.n118 2.27754
R1421 VDD.n122 VDD.n121 2.27754
R1422 VDD.n242 VDD.n202 2.25504
R1423 VDD.n52 VDD.n51 2.2505
R1424 VDD.n135 VDD.n134 1.7738
R1425 VDD.n18 VDD.n12 1.5755
R1426 VDD.n82 VDD.t50 1.51853
R1427 VDD.n58 VDD.n57 1.4255
R1428 VDD.n125 VDD.n124 1.3505
R1429 VDD.n55 VDD.n54 1.313
R1430 VDD.n133 VDD.n132 1.24541
R1431 VDD.n123 VDD.n120 1.238
R1432 VDD.n128 VDD.n123 1.15979
R1433 VDD.n132 VDD.n130 1.09451
R1434 VDD.n56 VDD.n55 1.02276
R1435 VDD.n126 VDD.n125 0.954149
R1436 VDD.n59 VDD.n58 0.77924
R1437 VDD.n14 VDD.n13 0.759513
R1438 VDD.n256 VDD.n254 0.679542
R1439 VDD.n15 VDD.t4 0.380007
R1440 VDD.n134 VDD.n133 0.113071
R1441 VDD.n46 VDD.n45 0.107201
R1442 VDD.n164 VDD.n163 0.107201
R1443 VDD.n167 VDD.n166 0.107201
R1444 VDD.n170 VDD.n169 0.107201
R1445 VDD.n173 VDD.n172 0.107201
R1446 VDD.n178 VDD.n177 0.107201
R1447 VDD.n181 VDD.n180 0.107201
R1448 VDD.n184 VDD.n183 0.107201
R1449 VDD.n189 VDD.n188 0.107201
R1450 VDD.n192 VDD.n191 0.107201
R1451 VDD.n195 VDD.n194 0.107201
R1452 VDD.n32 VDD.n31 0.107201
R1453 VDD.n31 VDD.n30 0.107201
R1454 VDD.n28 VDD.n27 0.107201
R1455 VDD.n27 VDD.n26 0.107201
R1456 VDD.n24 VDD.n23 0.107201
R1457 VDD.n214 VDD.n213 0.107201
R1458 VDD.n217 VDD.n216 0.107201
R1459 VDD.n218 VDD.n217 0.107201
R1460 VDD.n221 VDD.n220 0.107201
R1461 VDD.n222 VDD.n221 0.107201
R1462 VDD.n223 VDD.n222 0.107201
R1463 VDD.n226 VDD.n225 0.107201
R1464 VDD.n227 VDD.n226 0.107201
R1465 VDD.n230 VDD.n229 0.107201
R1466 VDD.n231 VDD.n230 0.107201
R1467 VDD.n232 VDD.n231 0.107201
R1468 VDD.n235 VDD.n234 0.107201
R1469 VDD.n236 VDD.n235 0.107201
R1470 VDD.n187 VDD.n186 0.102562
R1471 VDD.n228 VDD.n227 0.102562
R1472 VDD.n69 VDD.n67 0.0995431
R1473 VDD.n71 VDD.n69 0.0995431
R1474 VDD.n76 VDD.n74 0.0995431
R1475 VDD.n78 VDD.n76 0.0995431
R1476 VDD.n80 VDD.n78 0.0995431
R1477 VDD.n85 VDD.n83 0.0995431
R1478 VDD.n87 VDD.n85 0.0995431
R1479 VDD.n89 VDD.n87 0.0995431
R1480 VDD.n94 VDD.n92 0.0995431
R1481 VDD.n96 VDD.n94 0.0995431
R1482 VDD.n101 VDD.n99 0.0995431
R1483 VDD.n103 VDD.n101 0.0995431
R1484 VDD.n105 VDD.n103 0.0995431
R1485 VDD.n257 VDD.n253 0.0995431
R1486 VDD.n251 VDD.n250 0.0995431
R1487 VDD.n250 VDD.n249 0.0995431
R1488 VDD.n249 VDD.n248 0.0995431
R1489 VDD.n72 VDD.n71 0.0986818
R1490 VDD.n175 VDD.n174 0.0979227
R1491 VDD.n49 VDD.n48 0.0951392
R1492 VDD.n33 VDD.n32 0.0946753
R1493 VDD.n176 VDD.n175 0.0923557
R1494 VDD.n219 VDD.n218 0.0923557
R1495 VDD VDD.n108 0.0917919
R1496 VDD.n92 VDD.n90 0.0909306
R1497 VDD.n186 VDD.n185 0.0877165
R1498 VDD.n44 VDD.n43 0.0840052
R1499 VDD.n29 VDD.n28 0.0840052
R1500 VDD.n165 VDD.n164 0.0821495
R1501 VDD.n26 VDD.n25 0.0821495
R1502 VDD.n108 VDD.n106 0.0814569
R1503 VDD.n64 VDD.n63 0.0810263
R1504 VDD.n190 VDD.n189 0.0784381
R1505 VDD.n237 VDD.n236 0.0784381
R1506 VDD.n201 VDD.n200 0.0765825
R1507 VDD.n172 VDD.n171 0.073799
R1508 VDD.n216 VDD.n215 0.073799
R1509 VDD.n253 VDD.n252 0.0728445
R1510 VDD.n179 VDD.n178 0.068232
R1511 VDD.n197 VDD.n196 0.0673041
R1512 VDD.n247 VDD.n246 0.0650933
R1513 VDD.n183 VDD.n182 0.0635928
R1514 VDD.n225 VDD.n224 0.0635928
R1515 VDD.n97 VDD.n96 0.0633708
R1516 VDD.n47 VDD.n46 0.0598814
R1517 VDD.n168 VDD.n167 0.0580258
R1518 VDD.n67 VDD.n65 0.0556196
R1519 VDD.n193 VDD.n192 0.0543144
R1520 VDD.n233 VDD.n232 0.0543144
R1521 VDD.n81 VDD.n80 0.0538971
R1522 VDD.n194 VDD.n193 0.0533866
R1523 VDD.n234 VDD.n233 0.0533866
R1524 VDD.n169 VDD.n168 0.0496753
R1525 VDD.n48 VDD.n47 0.0478196
R1526 VDD.n83 VDD.n81 0.0461459
R1527 VDD.n65 VDD.n64 0.0444234
R1528 VDD.n182 VDD.n181 0.0441082
R1529 VDD.n224 VDD.n223 0.0441082
R1530 VDD.n180 VDD.n179 0.0394691
R1531 VDD.n99 VDD.n97 0.0366722
R1532 VDD.n171 VDD.n170 0.0339021
R1533 VDD.n215 VDD.n214 0.0339021
R1534 VDD.n196 VDD.n195 0.0301907
R1535 VDD.n191 VDD.n190 0.0292629
R1536 VDD.n248 VDD.n247 0.0280598
R1537 VDD.n252 VDD.n251 0.0271986
R1538 VDD.n166 VDD.n165 0.0255515
R1539 VDD.n25 VDD.n24 0.0255515
R1540 VDD.n45 VDD.n44 0.0236959
R1541 VDD.n30 VDD.n29 0.0236959
R1542 VDD.n242 VDD.n241 0.021875
R1543 VDD.n245 VDD.n244 0.0203086
R1544 VDD.n185 VDD.n184 0.0199845
R1545 VDD.n199 VDD.n198 0.0190567
R1546 VDD.n63 VDD.n62 0.0190167
R1547 VDD.n106 VDD.n105 0.0185861
R1548 VDD.n51 VDD.n50 0.0176649
R1549 VDD.n35 VDD.n34 0.0167371
R1550 VDD.n240 VDD.n239 0.0158093
R1551 VDD.n177 VDD.n176 0.0153454
R1552 VDD.n220 VDD.n219 0.0153454
R1553 VDD.n240 VDD.n237 0.0139536
R1554 VDD.n34 VDD.n33 0.0130258
R1555 VDD.n50 VDD.n49 0.0125619
R1556 VDD.n202 VDD.n201 0.0121334
R1557 VDD.n198 VDD.n197 0.0107062
R1558 VDD.n174 VDD.n173 0.00977835
R1559 VDD.n90 VDD.n89 0.00911244
R1560 VDD VDD.n257 0.0082512
R1561 VDD.n246 VDD.n245 0.00738995
R1562 VDD.n244 VDD.n243 0.00684906
R1563 VDD.n37 VDD.n35 0.00618398
R1564 VDD.n239 VDD.n238 0.00606701
R1565 VDD.n188 VDD.n187 0.00513918
R1566 VDD.n229 VDD.n228 0.00513918
R1567 VDD.n202 VDD.n199 0.00192811
R1568 VDD.n62 VDD.n53 0.00179187
R1569 VDD.n163 VDD.n162 0.00142783
R1570 VDD.n74 VDD.n72 0.00136124
R1571 SD2_0.n56 SD2_0.n55 3.51036
R1572 SD2_0.n72 SD2_0.n35 3.49563
R1573 SD2_0.n100 SD2_0.n3 3.49081
R1574 SD2_0.n115 SD2_0.n114 3.09757
R1575 SD2_0 SD2_0.n1 3.08774
R1576 SD2_0.n66 SD2_0.n37 3.08345
R1577 SD2_0.n63 SD2_0.n42 3.08151
R1578 SD2_0.n84 SD2_0.n23 3.07949
R1579 SD2_0.n78 SD2_0.n33 3.07685
R1580 SD2_0.n57 SD2_0.n51 3.0768
R1581 SD2_0.n91 SD2_0.n17 3.07536
R1582 SD2_0.n89 SD2_0.n21 3.07535
R1583 SD2_0.n60 SD2_0.n47 3.07497
R1584 SD2_0.n81 SD2_0.n28 3.07433
R1585 SD2_0.n97 SD2_0.n8 3.07386
R1586 SD2_0.n94 SD2_0.n13 3.07165
R1587 SD2_0.n112 SD2_0.t21 3.03383
R1588 SD2_0.n112 SD2_0.n111 3.03383
R1589 SD2_0.n114 SD2_0.t48 3.03383
R1590 SD2_0.n114 SD2_0.n113 3.03383
R1591 SD2_0.n102 SD2_0.t6 3.03383
R1592 SD2_0.n102 SD2_0.n101 3.03383
R1593 SD2_0.n5 SD2_0.t52 3.03383
R1594 SD2_0.n5 SD2_0.n4 3.03383
R1595 SD2_0.n10 SD2_0.t32 3.03383
R1596 SD2_0.n10 SD2_0.n9 3.03383
R1597 SD2_0.n15 SD2_0.t1 3.03383
R1598 SD2_0.n15 SD2_0.n14 3.03383
R1599 SD2_0.n19 SD2_0.t15 3.03383
R1600 SD2_0.n19 SD2_0.n18 3.03383
R1601 SD2_0.n86 SD2_0.t41 3.03383
R1602 SD2_0.n86 SD2_0.n85 3.03383
R1603 SD2_0.n25 SD2_0.t19 3.03383
R1604 SD2_0.n25 SD2_0.n24 3.03383
R1605 SD2_0.n30 SD2_0.t5 3.03383
R1606 SD2_0.n30 SD2_0.n29 3.03383
R1607 SD2_0.n35 SD2_0.t42 3.03383
R1608 SD2_0.n35 SD2_0.n34 3.03383
R1609 SD2_0.n74 SD2_0.t33 3.03383
R1610 SD2_0.n74 SD2_0.n73 3.03383
R1611 SD2_0.n37 SD2_0.t18 3.03383
R1612 SD2_0.n37 SD2_0.n36 3.03383
R1613 SD2_0.n68 SD2_0.t43 3.03383
R1614 SD2_0.n68 SD2_0.n67 3.03383
R1615 SD2_0.n39 SD2_0.t9 3.03383
R1616 SD2_0.n39 SD2_0.n38 3.03383
R1617 SD2_0.n44 SD2_0.t51 3.03383
R1618 SD2_0.n44 SD2_0.n43 3.03383
R1619 SD2_0.n49 SD2_0.t26 3.03383
R1620 SD2_0.n49 SD2_0.n48 3.03383
R1621 SD2_0.n53 SD2_0.t3 3.03383
R1622 SD2_0.n53 SD2_0.n52 3.03383
R1623 SD2_0.n55 SD2_0.t7 3.03383
R1624 SD2_0.n55 SD2_0.n54 3.03383
R1625 SD2_0.n51 SD2_0.t2 3.03383
R1626 SD2_0.n51 SD2_0.n50 3.03383
R1627 SD2_0.n47 SD2_0.t28 3.03383
R1628 SD2_0.n47 SD2_0.n46 3.03383
R1629 SD2_0.n42 SD2_0.t40 3.03383
R1630 SD2_0.n42 SD2_0.n41 3.03383
R1631 SD2_0.n33 SD2_0.t37 3.03383
R1632 SD2_0.n33 SD2_0.n32 3.03383
R1633 SD2_0.n28 SD2_0.t4 3.03383
R1634 SD2_0.n28 SD2_0.n27 3.03383
R1635 SD2_0.n23 SD2_0.t20 3.03383
R1636 SD2_0.n23 SD2_0.n22 3.03383
R1637 SD2_0.n21 SD2_0.t60 3.03383
R1638 SD2_0.n21 SD2_0.n20 3.03383
R1639 SD2_0.n17 SD2_0.t16 3.03383
R1640 SD2_0.n17 SD2_0.n16 3.03383
R1641 SD2_0.n13 SD2_0.t44 3.03383
R1642 SD2_0.n13 SD2_0.n12 3.03383
R1643 SD2_0.n8 SD2_0.t27 3.03383
R1644 SD2_0.n8 SD2_0.n7 3.03383
R1645 SD2_0.n3 SD2_0.t50 3.03383
R1646 SD2_0.n3 SD2_0.n2 3.03383
R1647 SD2_0.n1 SD2_0.t8 3.03383
R1648 SD2_0.n1 SD2_0.n0 3.03383
R1649 SD2_0.n106 SD2_0.t49 3.03383
R1650 SD2_0.n106 SD2_0.n105 3.03383
R1651 SD2_0.n92 SD2_0.n15 2.75441
R1652 SD2_0.n58 SD2_0.n49 2.75441
R1653 SD2_0.n90 SD2_0.n19 2.75396
R1654 SD2_0.n115 SD2_0.n112 2.38302
R1655 SD2_0.n56 SD2_0.n53 2.38112
R1656 SD2_0.n104 SD2_0.n103 2.24447
R1657 SD2_0.n70 SD2_0.n69 2.24419
R1658 SD2_0.n76 SD2_0.n75 2.24419
R1659 SD2_0.n110 SD2_0.n109 1.49481
R1660 SD2_0.n88 SD2_0.n87 1.4947
R1661 SD2_0.n79 SD2_0.n31 1.49456
R1662 SD2_0.n98 SD2_0.n6 1.49456
R1663 SD2_0.n61 SD2_0.n45 1.49431
R1664 SD2_0.n64 SD2_0.n40 1.49431
R1665 SD2_0.n82 SD2_0.n26 1.49431
R1666 SD2_0.n95 SD2_0.n11 1.49431
R1667 SD2_0.n6 SD2_0.n5 1.26105
R1668 SD2_0.n11 SD2_0.n10 1.26092
R1669 SD2_0.n45 SD2_0.n44 1.2606
R1670 SD2_0.n103 SD2_0.n102 1.26047
R1671 SD2_0.n26 SD2_0.n25 1.26047
R1672 SD2_0.n31 SD2_0.n30 1.26016
R1673 SD2_0.n87 SD2_0.n86 1.25971
R1674 SD2_0.n75 SD2_0.n74 1.25971
R1675 SD2_0.n69 SD2_0.n68 1.25971
R1676 SD2_0.n40 SD2_0.n39 1.25957
R1677 SD2_0.n108 SD2_0.n106 1.25796
R1678 SD2_0.n57 SD2_0.n56 0.612813
R1679 SD2_0.n99 SD2_0.n98 0.611577
R1680 SD2_0.n89 SD2_0.n88 0.610706
R1681 SD2_0.n91 SD2_0.n90 0.608363
R1682 SD2_0.n65 SD2_0.n64 0.596198
R1683 SD2_0.n110 SD2_0.n104 0.591867
R1684 SD2_0.n71 SD2_0.n70 0.591483
R1685 SD2_0.n116 SD2_0.n115 0.585815
R1686 SD2_0.n80 SD2_0.n79 0.584906
R1687 SD2_0.n62 SD2_0.n61 0.583676
R1688 SD2_0.n59 SD2_0.n58 0.582832
R1689 SD2_0.n93 SD2_0.n92 0.582832
R1690 SD2_0.n96 SD2_0.n95 0.582069
R1691 SD2_0.n83 SD2_0.n82 0.579994
R1692 SD2_0.n77 SD2_0.n76 0.577353
R1693 SD2_0 SD2_0.n116 0.0278418
R1694 SD2_0.n63 SD2_0.n62 0.0244241
R1695 SD2_0.n84 SD2_0.n83 0.0244241
R1696 SD2_0.n94 SD2_0.n93 0.0244241
R1697 SD2_0.n97 SD2_0.n96 0.0232848
R1698 SD2_0.n78 SD2_0.n77 0.0221456
R1699 SD2_0.n81 SD2_0.n80 0.0221456
R1700 SD2_0.n60 SD2_0.n59 0.0210063
R1701 SD2_0.n61 SD2_0.n60 0.0183749
R1702 SD2_0.n79 SD2_0.n78 0.0176185
R1703 SD2_0.n82 SD2_0.n81 0.0172357
R1704 SD2_0.n66 SD2_0.n65 0.016908
R1705 SD2_0.n76 SD2_0.n72 0.016908
R1706 SD2_0.n98 SD2_0.n97 0.0164793
R1707 SD2_0.n104 SD2_0.n100 0.0163417
R1708 SD2_0.n58 SD2_0.n57 0.015337
R1709 SD2_0.n90 SD2_0.n89 0.015337
R1710 SD2_0.n88 SD2_0.n84 0.0150107
R1711 SD2_0.n64 SD2_0.n63 0.0149572
R1712 SD2_0.n95 SD2_0.n94 0.0149572
R1713 SD2_0.n70 SD2_0.n66 0.0146295
R1714 SD2_0.n72 SD2_0.n71 0.0146295
R1715 SD2_0.n92 SD2_0.n91 0.0141978
R1716 SD2_0 SD2_0.n110 0.0123049
R1717 SD2_0.n108 SD2_0.n107 0.00342725
R1718 SD2_0.n109 SD2_0.n108 0.00324374
R1719 SD2_0.n100 SD2_0.n99 0.00277848
R1720 G0_2.n20 G0_2.t14 117.912
R1721 G0_2.n34 G0_2.n33 105.725
R1722 G0_2.n22 G0_2.n21 103.823
R1723 G0_2.n24 G0_2.n23 103.823
R1724 G0_2.n26 G0_2.n25 103.823
R1725 G0_2.n28 G0_2.n27 103.823
R1726 G0_2.n30 G0_2.n29 103.823
R1727 G0_2.n32 G0_2.n31 103.823
R1728 G0_2.n3 G0_2.n2 103.823
R1729 G0_2.n5 G0_2.n4 103.823
R1730 G0_2.n7 G0_2.n6 103.823
R1731 G0_2.n9 G0_2.n8 103.823
R1732 G0_2.n11 G0_2.n10 103.823
R1733 G0_2.n13 G0_2.n12 103.823
R1734 G0_2.n15 G0_2.n14 103.823
R1735 G0_2.n2 G0_2.t8 33.7914
R1736 G0_2.n16 G0_2.n15 22.1091
R1737 G0_2.n21 G0_2.n20 21.0894
R1738 G0_2.n23 G0_2.n22 21.0894
R1739 G0_2.n25 G0_2.n24 21.0894
R1740 G0_2.n27 G0_2.n26 21.0894
R1741 G0_2.n29 G0_2.n28 21.0894
R1742 G0_2.n31 G0_2.n30 21.0894
R1743 G0_2.n33 G0_2.n32 21.0894
R1744 G0_2.n4 G0_2.n3 21.0894
R1745 G0_2.n6 G0_2.n5 21.0894
R1746 G0_2.n8 G0_2.n7 21.0894
R1747 G0_2.n10 G0_2.n9 21.0894
R1748 G0_2.n12 G0_2.n11 21.0894
R1749 G0_2.n14 G0_2.n13 21.0894
R1750 G0_2.n20 G0_2.t10 14.0895
R1751 G0_2.n21 G0_2.t6 14.0895
R1752 G0_2.n22 G0_2.t28 14.0895
R1753 G0_2.n23 G0_2.t1 14.0895
R1754 G0_2.n24 G0_2.t18 14.0895
R1755 G0_2.n25 G0_2.t25 14.0895
R1756 G0_2.n26 G0_2.t16 14.0895
R1757 G0_2.n27 G0_2.t9 14.0895
R1758 G0_2.n28 G0_2.t7 14.0895
R1759 G0_2.n29 G0_2.t3 14.0895
R1760 G0_2.n30 G0_2.t2 14.0895
R1761 G0_2.n31 G0_2.t29 14.0895
R1762 G0_2.n32 G0_2.t22 14.0895
R1763 G0_2.n33 G0_2.t17 14.0895
R1764 G0_2.n2 G0_2.t15 12.7025
R1765 G0_2.n3 G0_2.t21 12.7025
R1766 G0_2.n4 G0_2.t5 12.7025
R1767 G0_2.n5 G0_2.t13 12.7025
R1768 G0_2.n6 G0_2.t19 12.7025
R1769 G0_2.n7 G0_2.t26 12.7025
R1770 G0_2.n8 G0_2.t11 12.7025
R1771 G0_2.n9 G0_2.t30 12.7025
R1772 G0_2.n10 G0_2.t23 12.7025
R1773 G0_2.n11 G0_2.t0 12.7025
R1774 G0_2.n12 G0_2.t27 12.7025
R1775 G0_2.n13 G0_2.t12 12.7025
R1776 G0_2.n14 G0_2.t31 12.7025
R1777 G0_2.n15 G0_2.t20 12.7025
R1778 G0_2.n34 G0_2.t4 11.1355
R1779 G0_2.n17 G0_2.n1 8.0195
R1780 G0_2.n0 G0_2.t24 7.9575
R1781 G0_2 G0_2.n34 4.35404
R1782 G0_2.n18 G0_2.n16 3.4914
R1783 G0_2.n19 G0_2.n1 2.88425
R1784 G0_2.n1 G0_2.n0 2.3365
R1785 G0_2 G0_2.n19 2.2655
R1786 G0_2.n18 G0_2.n17 0.0105
R1787 G0_2.n19 G0_2.n18 0.0045
R1788 G1_1.n103 G1_1.n100 31.7026
R1789 G1_1.n65 G1_1.n64 28.879
R1790 G1_1.n63 G1_1.t131 24.5285
R1791 G1_1.n62 G1_1.t117 24.5285
R1792 G1_1.n59 G1_1.t101 24.5285
R1793 G1_1.n58 G1_1.t125 24.5285
R1794 G1_1.n55 G1_1.t115 24.5285
R1795 G1_1.n54 G1_1.t105 24.5285
R1796 G1_1.n51 G1_1.t143 24.5285
R1797 G1_1.n50 G1_1.t130 24.5285
R1798 G1_1.n86 G1_1.t136 24.5285
R1799 G1_1.n87 G1_1.t107 24.5285
R1800 G1_1.n90 G1_1.t112 24.5285
R1801 G1_1.n91 G1_1.t97 24.5285
R1802 G1_1.n94 G1_1.t100 24.5285
R1803 G1_1.n95 G1_1.t123 24.5285
R1804 G1_1.n98 G1_1.t121 24.5285
R1805 G1_1.n99 G1_1.t118 24.5285
R1806 G1_1.n186 G1_1.t46 23.86
R1807 G1_1.n110 G1_1.t36 23.86
R1808 G1_1.n186 G1_1.t50 23.1415
R1809 G1_1.n187 G1_1.t2 23.1415
R1810 G1_1.n184 G1_1.t24 23.1415
R1811 G1_1.n177 G1_1.t54 23.1415
R1812 G1_1.n175 G1_1.t8 23.1415
R1813 G1_1.n165 G1_1.t20 23.1415
R1814 G1_1.n163 G1_1.t30 23.1415
R1815 G1_1.n152 G1_1.t52 23.1415
R1816 G1_1.n150 G1_1.t40 23.1415
R1817 G1_1.n139 G1_1.t18 23.1415
R1818 G1_1.n137 G1_1.t12 23.1415
R1819 G1_1.n126 G1_1.t28 23.1415
R1820 G1_1.n124 G1_1.t26 23.1415
R1821 G1_1.n113 G1_1.t56 23.1415
R1822 G1_1.n110 G1_1.t0 23.1415
R1823 G1_1.n111 G1_1.t58 23.1415
R1824 G1_1.n188 G1_1.t38 13.8705
R1825 G1_1.n185 G1_1.t62 13.8705
R1826 G1_1.n178 G1_1.t14 13.8705
R1827 G1_1.n176 G1_1.t42 13.8705
R1828 G1_1.n166 G1_1.t60 13.8705
R1829 G1_1.n164 G1_1.t10 13.8705
R1830 G1_1.n153 G1_1.t6 13.8705
R1831 G1_1.n151 G1_1.t32 13.8705
R1832 G1_1.n140 G1_1.t34 13.8705
R1833 G1_1.n138 G1_1.t48 13.8705
R1834 G1_1.n127 G1_1.t4 13.8705
R1835 G1_1.n125 G1_1.t22 13.8705
R1836 G1_1.n114 G1_1.t16 13.8705
R1837 G1_1.n112 G1_1.t44 13.8705
R1838 G1_1.n64 G1_1.t127 13.6515
R1839 G1_1.n61 G1_1.t132 13.6515
R1840 G1_1.n60 G1_1.t119 13.6515
R1841 G1_1.n57 G1_1.t103 13.6515
R1842 G1_1.n56 G1_1.t129 13.6515
R1843 G1_1.n53 G1_1.t120 13.6515
R1844 G1_1.n52 G1_1.t106 13.6515
R1845 G1_1.n49 G1_1.t110 13.6515
R1846 G1_1.n85 G1_1.t138 13.6515
R1847 G1_1.n88 G1_1.t137 13.6515
R1848 G1_1.n89 G1_1.t122 13.6515
R1849 G1_1.n92 G1_1.t113 13.6515
R1850 G1_1.n93 G1_1.t98 13.6515
R1851 G1_1.n96 G1_1.t102 13.6515
R1852 G1_1.n97 G1_1.t128 13.6515
R1853 G1_1.n100 G1_1.t133 13.6515
R1854 G1_1.n64 G1_1.n63 10.6935
R1855 G1_1.n63 G1_1.n62 10.6935
R1856 G1_1.n62 G1_1.n61 10.6935
R1857 G1_1.n61 G1_1.n60 10.6935
R1858 G1_1.n60 G1_1.n59 10.6935
R1859 G1_1.n59 G1_1.n58 10.6935
R1860 G1_1.n58 G1_1.n57 10.6935
R1861 G1_1.n57 G1_1.n56 10.6935
R1862 G1_1.n56 G1_1.n55 10.6935
R1863 G1_1.n55 G1_1.n54 10.6935
R1864 G1_1.n54 G1_1.n53 10.6935
R1865 G1_1.n53 G1_1.n52 10.6935
R1866 G1_1.n52 G1_1.n51 10.6935
R1867 G1_1.n51 G1_1.n50 10.6935
R1868 G1_1.n50 G1_1.n49 10.6935
R1869 G1_1.n86 G1_1.n85 10.6935
R1870 G1_1.n87 G1_1.n86 10.6935
R1871 G1_1.n88 G1_1.n87 10.6935
R1872 G1_1.n89 G1_1.n88 10.6935
R1873 G1_1.n90 G1_1.n89 10.6935
R1874 G1_1.n91 G1_1.n90 10.6935
R1875 G1_1.n92 G1_1.n91 10.6935
R1876 G1_1.n93 G1_1.n92 10.6935
R1877 G1_1.n94 G1_1.n93 10.6935
R1878 G1_1.n95 G1_1.n94 10.6935
R1879 G1_1.n96 G1_1.n95 10.6935
R1880 G1_1.n97 G1_1.n96 10.6935
R1881 G1_1.n98 G1_1.n97 10.6935
R1882 G1_1.n99 G1_1.n98 10.6935
R1883 G1_1.n100 G1_1.n99 10.6935
R1884 G1_1.n187 G1_1.n186 9.98997
R1885 G1_1.n188 G1_1.n187 9.98997
R1886 G1_1.n185 G1_1.n184 9.98997
R1887 G1_1.n178 G1_1.n177 9.98997
R1888 G1_1.n176 G1_1.n175 9.98997
R1889 G1_1.n166 G1_1.n165 9.98997
R1890 G1_1.n164 G1_1.n163 9.98997
R1891 G1_1.n153 G1_1.n152 9.98997
R1892 G1_1.n151 G1_1.n150 9.98997
R1893 G1_1.n140 G1_1.n139 9.98997
R1894 G1_1.n138 G1_1.n137 9.98997
R1895 G1_1.n127 G1_1.n126 9.98997
R1896 G1_1.n125 G1_1.n124 9.98997
R1897 G1_1.n114 G1_1.n113 9.98997
R1898 G1_1.n111 G1_1.n110 9.98997
R1899 G1_1.n112 G1_1.n111 9.98997
R1900 G1_1.n115 G1_1.n112 6.72418
R1901 G1_1.n102 G1_1.n101 6.14854
R1902 G1_1.n48 G1_1.t93 6.14854
R1903 G1_1.n179 G1_1.n176 5.85971
R1904 G1_1.n128 G1_1.n125 5.85971
R1905 G1_1.n154 G1_1.n151 5.37945
R1906 G1_1.n2 G1_1.n1 5.24336
R1907 G1_1.n189 G1_1.n188 5.18734
R1908 G1_1.n167 G1_1.n164 5.18734
R1909 G1_1.n141 G1_1.n140 5.18734
R1910 G1_1.n189 G1_1.n185 4.80313
R1911 G1_1.n167 G1_1.n166 4.80313
R1912 G1_1.n141 G1_1.n138 4.80313
R1913 G1_1.n154 G1_1.n153 4.61103
R1914 G1_1.n104 G1_1.n84 4.29029
R1915 G1_1.n179 G1_1.n178 4.13076
R1916 G1_1.n128 G1_1.n127 4.13076
R1917 G1_1.n47 G1_1.n4 3.44202
R1918 G1_1.n45 G1_1.n8 3.44202
R1919 G1_1.n43 G1_1.n12 3.44202
R1920 G1_1.n41 G1_1.n16 3.44202
R1921 G1_1.n39 G1_1.n20 3.44202
R1922 G1_1.n37 G1_1.n24 3.44202
R1923 G1_1.n35 G1_1.n28 3.44202
R1924 G1_1.n33 G1_1.n32 3.44202
R1925 G1_1.n34 G1_1.n30 3.41854
R1926 G1_1.n36 G1_1.n26 3.41854
R1927 G1_1.n38 G1_1.n22 3.41854
R1928 G1_1.n40 G1_1.n18 3.41854
R1929 G1_1.n42 G1_1.n14 3.41854
R1930 G1_1.n44 G1_1.n10 3.41854
R1931 G1_1.n46 G1_1.n6 3.41854
R1932 G1_1.n115 G1_1.n114 3.26629
R1933 G1_1.n2 G1_1.t47 3.03383
R1934 G1_1.n122 G1_1.t23 3.03383
R1935 G1_1.n122 G1_1.n121 3.03383
R1936 G1_1.n135 G1_1.t49 3.03383
R1937 G1_1.n135 G1_1.n134 3.03383
R1938 G1_1.n148 G1_1.t33 3.03383
R1939 G1_1.n148 G1_1.n147 3.03383
R1940 G1_1.n161 G1_1.t11 3.03383
R1941 G1_1.n161 G1_1.n160 3.03383
R1942 G1_1.n173 G1_1.t43 3.03383
R1943 G1_1.n173 G1_1.n172 3.03383
R1944 G1_1.n192 G1_1.t63 3.03383
R1945 G1_1.n192 G1_1.n191 3.03383
R1946 G1_1.n108 G1_1.t45 3.03383
R1947 G1_1.n108 G1_1.n107 3.03383
R1948 G1_1.n83 G1_1.t1 3.03383
R1949 G1_1.n83 G1_1.n82 3.03383
R1950 G1_1.n81 G1_1.t57 3.03383
R1951 G1_1.n81 G1_1.n80 3.03383
R1952 G1_1.n79 G1_1.t29 3.03383
R1953 G1_1.n79 G1_1.n78 3.03383
R1954 G1_1.n77 G1_1.t19 3.03383
R1955 G1_1.n77 G1_1.n76 3.03383
R1956 G1_1.n75 G1_1.t53 3.03383
R1957 G1_1.n75 G1_1.n74 3.03383
R1958 G1_1.n73 G1_1.t21 3.03383
R1959 G1_1.n73 G1_1.n72 3.03383
R1960 G1_1.n71 G1_1.t55 3.03383
R1961 G1_1.n71 G1_1.n70 3.03383
R1962 G1_1.n69 G1_1.t3 3.03383
R1963 G1_1.n69 G1_1.n68 3.03383
R1964 G1_1.n193 G1_1.n192 2.91531
R1965 G1_1.n136 G1_1.n135 2.89977
R1966 G1_1.n123 G1_1.n122 2.89762
R1967 G1_1.n162 G1_1.n161 2.89762
R1968 G1_1.n149 G1_1.n148 2.89547
R1969 G1_1.n174 G1_1.n173 2.88224
R1970 G1_1.n190 G1_1.n189 2.8805
R1971 G1_1.n180 G1_1.n179 2.8805
R1972 G1_1.n168 G1_1.n167 2.8805
R1973 G1_1.n155 G1_1.n154 2.8805
R1974 G1_1.n142 G1_1.n141 2.8805
R1975 G1_1.n129 G1_1.n128 2.8805
R1976 G1_1.n116 G1_1.n115 2.8805
R1977 G1_1.n109 G1_1.n108 2.87637
R1978 G1_1.n182 G1_1.n71 2.79692
R1979 G1_1.n157 G1_1.n75 2.7913
R1980 G1_1.n105 G1_1.n83 2.7872
R1981 G1_1.n131 G1_1.n79 2.78609
R1982 G1_1.n196 G1_1.n69 2.78592
R1983 G1_1.n118 G1_1.n81 2.78535
R1984 G1_1.n170 G1_1.n73 2.78042
R1985 G1_1.n144 G1_1.n77 2.78024
R1986 G1_1.n30 G1_1.t90 2.7305
R1987 G1_1.n30 G1_1.n29 2.7305
R1988 G1_1.n26 G1_1.t81 2.7305
R1989 G1_1.n26 G1_1.n25 2.7305
R1990 G1_1.n22 G1_1.t86 2.7305
R1991 G1_1.n22 G1_1.n21 2.7305
R1992 G1_1.n18 G1_1.t87 2.7305
R1993 G1_1.n18 G1_1.n17 2.7305
R1994 G1_1.n14 G1_1.t92 2.7305
R1995 G1_1.n14 G1_1.n13 2.7305
R1996 G1_1.n10 G1_1.t94 2.7305
R1997 G1_1.n10 G1_1.n9 2.7305
R1998 G1_1.n6 G1_1.t83 2.7305
R1999 G1_1.n6 G1_1.n5 2.7305
R2000 G1_1.n4 G1_1.t85 2.7305
R2001 G1_1.n4 G1_1.n3 2.7305
R2002 G1_1.n8 G1_1.t89 2.7305
R2003 G1_1.n8 G1_1.n7 2.7305
R2004 G1_1.n12 G1_1.t95 2.7305
R2005 G1_1.n12 G1_1.n11 2.7305
R2006 G1_1.n16 G1_1.t80 2.7305
R2007 G1_1.n16 G1_1.n15 2.7305
R2008 G1_1.n20 G1_1.t82 2.7305
R2009 G1_1.n20 G1_1.n19 2.7305
R2010 G1_1.n24 G1_1.t88 2.7305
R2011 G1_1.n24 G1_1.n23 2.7305
R2012 G1_1.n28 G1_1.t84 2.7305
R2013 G1_1.n28 G1_1.n27 2.7305
R2014 G1_1.n32 G1_1.t91 2.7305
R2015 G1_1.n32 G1_1.n31 2.7305
R2016 G1_1.n199 G1_1.n67 2.25044
R2017 G1_1.n105 G1_1.n104 1.80349
R2018 G1_1.n65 G1_1.n48 1.70664
R2019 G1_1.n66 G1_1.n2 1.65036
R2020 G1_1.n103 G1_1.n102 1.58193
R2021 G1_1.n194 G1_1.n193 1.1231
R2022 G1_1.n130 G1_1.n129 1.12283
R2023 G1_1.n143 G1_1.n142 1.12283
R2024 G1_1.n156 G1_1.n155 1.12283
R2025 G1_1.n169 G1_1.n168 1.12283
R2026 G1_1.n117 G1_1.n116 0.897749
R2027 G1_1.n181 G1_1.n180 0.897685
R2028 G1_1.n106 G1_1.n105 0.815399
R2029 G1_1.n171 G1_1.n170 0.807847
R2030 G1_1.n197 G1_1.n196 0.567009
R2031 G1_1.n34 G1_1.n33 0.525071
R2032 G1_1.n35 G1_1.n34 0.525071
R2033 G1_1.n36 G1_1.n35 0.525071
R2034 G1_1.n37 G1_1.n36 0.525071
R2035 G1_1.n38 G1_1.n37 0.525071
R2036 G1_1.n39 G1_1.n38 0.525071
R2037 G1_1.n40 G1_1.n39 0.525071
R2038 G1_1.n41 G1_1.n40 0.525071
R2039 G1_1.n42 G1_1.n41 0.525071
R2040 G1_1.n43 G1_1.n42 0.525071
R2041 G1_1.n44 G1_1.n43 0.525071
R2042 G1_1.n45 G1_1.n44 0.525071
R2043 G1_1.n46 G1_1.n45 0.525071
R2044 G1_1.n47 G1_1.n46 0.525071
R2045 G1_1.n48 G1_1.n47 0.525071
R2046 G1_1.n144 G1_1.n143 0.472321
R2047 G1_1.n157 G1_1.n156 0.470978
R2048 G1_1.n170 G1_1.n169 0.463775
R2049 G1_1.n182 G1_1.n181 0.463101
R2050 G1_1.n131 G1_1.n130 0.459551
R2051 G1_1.n196 G1_1.n195 0.454175
R2052 G1_1.n118 G1_1.n117 0.450213
R2053 G1_1.n119 G1_1.n118 0.444603
R2054 G1_1.n145 G1_1.n144 0.440282
R2055 G1_1.n158 G1_1.n157 0.434458
R2056 G1_1.n132 G1_1.n131 0.434202
R2057 G1_1.n183 G1_1.n182 0.430393
R2058 G1_1.n66 G1_1.n65 0.320822
R2059 G1_1.n104 G1_1.n103 0.306943
R2060 G1_1.n198 G1_1.n197 0.103625
R2061 G1_1.n181 G1_1.n171 0.0335252
R2062 G1_1.n117 G1_1.n106 0.0328885
R2063 G1_1.n195 G1_1.n194 0.0292629
R2064 G1_1.n120 G1_1.n119 0.0283351
R2065 G1_1.n133 G1_1.n132 0.0283351
R2066 G1_1.n146 G1_1.n145 0.0283351
R2067 G1_1.n159 G1_1.n158 0.0283351
R2068 G1_1.n194 G1_1.n183 0.0283351
R2069 G1_1.n129 G1_1.n123 0.0278529
R2070 G1_1.n142 G1_1.n136 0.0278529
R2071 G1_1.n155 G1_1.n149 0.0278529
R2072 G1_1.n168 G1_1.n162 0.0278529
R2073 G1_1 G1_1.n200 0.017375
R2074 G1_1.n116 G1_1.n109 0.0163824
R2075 G1_1.n1 G1_1.n0 0.00907143
R2076 G1_1 G1_1.n199 0.00887472
R2077 G1_1.n180 G1_1.n174 0.0086
R2078 G1_1.n130 G1_1.n120 0.00817049
R2079 G1_1.n143 G1_1.n133 0.00817049
R2080 G1_1.n156 G1_1.n146 0.00817049
R2081 G1_1.n169 G1_1.n159 0.00817049
R2082 G1_1.n193 G1_1.n190 0.00782059
R2083 G1_1.n67 G1_1.n66 0.00615724
R2084 G1_1.n199 G1_1.n198 0.00324972
R2085 G1_1.n67 G1_1.n0 0.00192857
R2086 SD0_1.n103 SD0_1.n101 6.33762
R2087 SD0_1.n107 SD0_1.n106 4.5005
R2088 SD0_1.n88 SD0_1.n5 3.43055
R2089 SD0_1.n73 SD0_1.n13 3.42597
R2090 SD0_1.n37 SD0_1.n36 3.01986
R2091 SD0_1.n41 SD0_1.n28 3.00577
R2092 SD0_1.n94 SD0_1.n3 3.00356
R2093 SD0_1.n38 SD0_1.n32 3.00189
R2094 SD0_1.n47 SD0_1.n26 3.00189
R2095 SD0_1.n62 SD0_1.n17 3.00176
R2096 SD0_1.n71 SD0_1.n15 2.99921
R2097 SD0_1.n59 SD0_1.n19 2.99854
R2098 SD0_1.n100 SD0_1.n1 2.99694
R2099 SD0_1.n79 SD0_1.n9 2.99611
R2100 SD0_1.n114 SD0_1.n113 2.9953
R2101 SD0_1.n85 SD0_1.n7 2.99257
R2102 SD0_1.n119 SD0_1.n109 2.98849
R2103 SD0_1.n50 SD0_1.n21 2.98849
R2104 SD0_1.n39 SD0_1.n30 2.93125
R2105 SD0_1.n34 SD0_1.n33 2.90218
R2106 SD0_1.n7 SD0_1.n6 2.90217
R2107 SD0_1.n113 SD0_1.n112 2.90217
R2108 SD0_1.n17 SD0_1.n16 2.90217
R2109 SD0_1.n19 SD0_1.n18 2.90217
R2110 SD0_1.n1 SD0_1.n0 2.90217
R2111 SD0_1.n68 SD0_1.n67 2.90215
R2112 SD0_1.n76 SD0_1.n75 2.90213
R2113 SD0_1.n3 SD0_1.n2 2.90213
R2114 SD0_1.n32 SD0_1.n31 2.90211
R2115 SD0_1.n26 SD0_1.n25 2.90211
R2116 SD0_1.n116 SD0_1.n115 2.90211
R2117 SD0_1.n82 SD0_1.n81 2.90211
R2118 SD0_1.n11 SD0_1.n10 2.90211
R2119 SD0_1.n36 SD0_1.n35 2.90209
R2120 SD0_1.n111 SD0_1.n110 2.90198
R2121 SD0_1.n106 SD0_1.n102 2.89755
R2122 SD0_1.n109 SD0_1.n108 2.87832
R2123 SD0_1.n43 SD0_1.n42 2.87832
R2124 SD0_1.n21 SD0_1.n20 2.87832
R2125 SD0_1.n15 SD0_1.n14 2.87832
R2126 SD0_1.n28 SD0_1.n27 2.87826
R2127 SD0_1.n96 SD0_1.n95 2.87826
R2128 SD0_1.n90 SD0_1.n89 2.87826
R2129 SD0_1.n9 SD0_1.n8 2.87826
R2130 SD0_1.n64 SD0_1.t6 2.7305
R2131 SD0_1.n64 SD0_1.n63 2.7305
R2132 SD0_1.n56 SD0_1.t59 2.7305
R2133 SD0_1.n56 SD0_1.n55 2.7305
R2134 SD0_1.n52 SD0_1.t30 2.7305
R2135 SD0_1.n52 SD0_1.n51 2.7305
R2136 SD0_1.n23 SD0_1.t37 2.7305
R2137 SD0_1.n23 SD0_1.n22 2.7305
R2138 SD0_1.n30 SD0_1.t61 2.7305
R2139 SD0_1.n30 SD0_1.n29 2.7305
R2140 SD0_1.n13 SD0_1.t42 2.7305
R2141 SD0_1.n13 SD0_1.n12 2.7305
R2142 SD0_1.n5 SD0_1.t4 2.7305
R2143 SD0_1.n5 SD0_1.n4 2.7305
R2144 SD0_1.n105 SD0_1.n104 2.66916
R2145 SD0_1.n106 SD0_1.n105 2.60815
R2146 SD0_1.n114 SD0_1.n111 2.51423
R2147 SD0_1.n37 SD0_1.n34 2.50503
R2148 SD0_1.n74 SD0_1.n11 2.50485
R2149 SD0_1.n96 SD0_1.t2 2.43825
R2150 SD0_1.n90 SD0_1.t62 2.43825
R2151 SD0_1.n9 SD0_1.t8 2.43825
R2152 SD0_1.n28 SD0_1.t39 2.43825
R2153 SD0_1.n15 SD0_1.t20 2.43821
R2154 SD0_1.n109 SD0_1.t49 2.4382
R2155 SD0_1.n43 SD0_1.t25 2.4382
R2156 SD0_1.n21 SD0_1.t60 2.4382
R2157 SD0_1.n36 SD0_1.t35 2.40706
R2158 SD0_1.n116 SD0_1.t14 2.40704
R2159 SD0_1.n82 SD0_1.t28 2.40704
R2160 SD0_1.n11 SD0_1.t22 2.40704
R2161 SD0_1.n32 SD0_1.t16 2.40704
R2162 SD0_1.n26 SD0_1.t26 2.40704
R2163 SD0_1.n3 SD0_1.t32 2.40703
R2164 SD0_1.n76 SD0_1.t47 2.40702
R2165 SD0_1.n68 SD0_1.t56 2.40701
R2166 SD0_1.n113 SD0_1.t7 2.407
R2167 SD0_1.n17 SD0_1.t46 2.407
R2168 SD0_1.n19 SD0_1.t12 2.407
R2169 SD0_1.n1 SD0_1.t0 2.407
R2170 SD0_1.n7 SD0_1.t38 2.40699
R2171 SD0_1.n34 SD0_1.t17 2.40698
R2172 SD0_1.n111 SD0_1.t41 2.40627
R2173 SD0_1.n58 SD0_1.n57 2.24993
R2174 SD0_1.n70 SD0_1.n69 2.24993
R2175 SD0_1.n84 SD0_1.n83 2.24993
R2176 SD0_1.n78 SD0_1.n77 2.24966
R2177 SD0_1.n45 SD0_1.n44 2.24539
R2178 SD0_1.n92 SD0_1.n91 2.24539
R2179 SD0_1.n98 SD0_1.n97 2.24539
R2180 SD0_1.n118 SD0_1.n117 2.24512
R2181 SD0_1.n54 SD0_1.n53 2.24486
R2182 SD0_1.n66 SD0_1.n65 2.24459
R2183 SD0_1.n102 SD0_1.t52 2.1354
R2184 SD0_1.n48 SD0_1.n24 1.49518
R2185 SD0_1.n65 SD0_1.n64 1.43739
R2186 SD0_1.n57 SD0_1.n56 1.43704
R2187 SD0_1.n53 SD0_1.n52 1.43704
R2188 SD0_1.n24 SD0_1.n23 1.43704
R2189 SD0_1.n69 SD0_1.n68 1.01061
R2190 SD0_1.n77 SD0_1.n76 1.01054
R2191 SD0_1.n117 SD0_1.n116 1.01041
R2192 SD0_1.n83 SD0_1.n82 1.01041
R2193 SD0_1.n44 SD0_1.n43 1.00827
R2194 SD0_1.n97 SD0_1.n96 1.00786
R2195 SD0_1.n91 SD0_1.n90 1.00786
R2196 SD0_1.n40 SD0_1.n39 0.607669
R2197 SD0_1.n78 SD0_1.n74 0.607459
R2198 SD0_1.n70 SD0_1.n66 0.604141
R2199 SD0_1.n58 SD0_1.n54 0.601465
R2200 SD0_1.n118 SD0_1.n114 0.60093
R2201 SD0_1.n38 SD0_1.n37 0.598744
R2202 SD0_1.n99 SD0_1.n98 0.597758
R2203 SD0_1.n93 SD0_1.n92 0.595615
R2204 SD0_1.n49 SD0_1.n48 0.594387
R2205 SD0_1.n87 SD0_1.n86 0.588179
R2206 SD0_1.n84 SD0_1.n80 0.586535
R2207 SD0_1.n121 SD0_1.n120 0.58175
R2208 SD0_1.n73 SD0_1.n72 0.580143
R2209 SD0_1.n61 SD0_1.n60 0.570963
R2210 SD0_1.n46 SD0_1.n45 0.564543
R2211 SD0_1.n105 SD0_1.n103 0.0618334
R2212 SD0_1.n47 SD0_1.n46 0.0251429
R2213 SD0_1.n60 SD0_1.n59 0.0240714
R2214 SD0_1.n72 SD0_1.n71 0.023
R2215 SD0_1.n80 SD0_1.n79 0.023
R2216 SD0_1.n86 SD0_1.n85 0.023
R2217 SD0_1 SD0_1.n121 0.0219286
R2218 SD0_1.n74 SD0_1.n73 0.017366
R2219 SD0_1.n62 SD0_1.n61 0.0159634
R2220 SD0_1.n50 SD0_1.n49 0.0154306
R2221 SD0_1.n119 SD0_1.n118 0.0148978
R2222 SD0_1.n39 SD0_1.n38 0.0145059
R2223 SD0_1.n45 SD0_1.n41 0.0143648
R2224 SD0_1.n92 SD0_1.n88 0.0143648
R2225 SD0_1.n54 SD0_1.n50 0.0143592
R2226 SD0_1.n66 SD0_1.n62 0.0138205
R2227 SD0_1.n98 SD0_1.n94 0.0132934
R2228 SD0_1.n48 SD0_1.n47 0.011654
R2229 SD0_1.n106 SD0_1.n101 0.006125
R2230 SD0_1.n100 SD0_1.n99 0.00585714
R2231 SD0_1.n41 SD0_1.n40 0.00478571
R2232 SD0_1.n88 SD0_1.n87 0.00478571
R2233 SD0_1.n94 SD0_1.n93 0.00478571
R2234 SD0_1.n79 SD0_1.n78 0.00474841
R2235 SD0_1.n59 SD0_1.n58 0.00421327
R2236 SD0_1.n71 SD0_1.n70 0.00421327
R2237 SD0_1.n85 SD0_1.n84 0.00421327
R2238 SD0_1.n120 SD0_1.n119 0.00264286
R2239 SD0_1.n107 SD0_1.n100 0.00157143
R2240 SD0_1 SD0_1.n107 0.00157143
R2241 G0_1.n31 G0_1.n30 53.6251
R2242 G0_1.n0 G0_1.t21 33.7184
R2243 G0_1.n1 G0_1.n0 21.0894
R2244 G0_1.n2 G0_1.n1 21.0894
R2245 G0_1.n3 G0_1.n2 21.0894
R2246 G0_1.n4 G0_1.n3 21.0894
R2247 G0_1.n5 G0_1.n4 21.0894
R2248 G0_1.n6 G0_1.n5 21.0894
R2249 G0_1.n7 G0_1.n6 21.0894
R2250 G0_1.n8 G0_1.n7 21.0894
R2251 G0_1.n9 G0_1.n8 21.0894
R2252 G0_1.n10 G0_1.n9 21.0894
R2253 G0_1.n11 G0_1.n10 21.0894
R2254 G0_1.n12 G0_1.n11 21.0894
R2255 G0_1.n13 G0_1.n12 21.0894
R2256 G0_1.n14 G0_1.n13 21.0894
R2257 G0_1.n15 G0_1.n14 21.0894
R2258 G0_1.n16 G0_1.n15 21.0894
R2259 G0_1.n17 G0_1.n16 21.0894
R2260 G0_1.n18 G0_1.n17 21.0894
R2261 G0_1.n19 G0_1.n18 21.0894
R2262 G0_1.n20 G0_1.n19 21.0894
R2263 G0_1.n21 G0_1.n20 21.0894
R2264 G0_1.n22 G0_1.n21 21.0894
R2265 G0_1.n23 G0_1.n22 21.0894
R2266 G0_1.n24 G0_1.n23 21.0894
R2267 G0_1.n25 G0_1.n24 21.0894
R2268 G0_1.n26 G0_1.n25 21.0894
R2269 G0_1.n27 G0_1.n26 21.0894
R2270 G0_1.n28 G0_1.n27 21.0894
R2271 G0_1.n29 G0_1.n28 21.0894
R2272 G0_1.n30 G0_1.n29 21.0894
R2273 G0_1.n0 G0_1.t7 13.3595
R2274 G0_1.n1 G0_1.t3 13.3595
R2275 G0_1.n4 G0_1.t1 13.3595
R2276 G0_1.n5 G0_1.t29 13.3595
R2277 G0_1.n8 G0_1.t28 13.3595
R2278 G0_1.n9 G0_1.t22 13.3595
R2279 G0_1.n12 G0_1.t19 13.3595
R2280 G0_1.n13 G0_1.t17 13.3595
R2281 G0_1.n16 G0_1.t16 13.3595
R2282 G0_1.n17 G0_1.t12 13.3595
R2283 G0_1.n20 G0_1.t30 13.3595
R2284 G0_1.n21 G0_1.t4 13.3595
R2285 G0_1.n24 G0_1.t27 13.3595
R2286 G0_1.n25 G0_1.t25 13.3595
R2287 G0_1.n28 G0_1.t13 13.3595
R2288 G0_1.n29 G0_1.t9 13.3595
R2289 G0_1.n2 G0_1.t24 12.6295
R2290 G0_1.n3 G0_1.t15 12.6295
R2291 G0_1.n6 G0_1.t10 12.6295
R2292 G0_1.n7 G0_1.t23 12.6295
R2293 G0_1.n10 G0_1.t2 12.6295
R2294 G0_1.n11 G0_1.t31 12.6295
R2295 G0_1.n14 G0_1.t18 12.6295
R2296 G0_1.n15 G0_1.t0 12.6295
R2297 G0_1.n18 G0_1.t8 12.6295
R2298 G0_1.n19 G0_1.t14 12.6295
R2299 G0_1.n22 G0_1.t20 12.6295
R2300 G0_1.n23 G0_1.t6 12.6295
R2301 G0_1.n26 G0_1.t5 12.6295
R2302 G0_1.n27 G0_1.t26 12.6295
R2303 G0_1.n30 G0_1.t11 12.6295
R2304 G0_1 G0_1.n31 4.09609
C0 G1_1 SD0_1 3.89f
C1 G1_1 VDD 18.4f
C2 VDD G3_1 0.00847f
C3 G1_1 G3_1 4.91e-19
C4 G3_2 G1_2 0.714f
C5 G0_2 G0_1 2.02f
C6 SD2_0 VDD 3.06f
C7 G0_1 SD0_1 0.653f
C8 G1_1 SD2_0 1.14f
C9 G0_1 VDD 0.00465f
C10 SD2_0 G3_1 0.0258f
C11 G1_1 G0_1 1.13f
C12 G0_2 G1_2 0.136f
C13 VDD G3_2 3.44f
C14 SD0_1 G1_2 0.0537f
C15 G1_1 G3_2 2.33f
C16 VDD G1_2 28.1f
C17 G3_2 G3_1 4.76f
C18 G1_1 G1_2 10.9f
C19 G3_1 G1_2 0.00788f
C20 G0_2 SD0_1 0.908f
C21 SD2_0 G3_2 3.46f
C22 G0_2 VDD 0.291f
C23 G1_1 G0_2 0.8f
C24 SD0_1 VDD 0.173f
C25 SD2_0 G1_2 1.43f
.ends

