* NGSPICE file created from GF_INV4_flat.ext - technology: gf180mcuC

.subckt GF_INV_4_PEX VSS VDD OUT IN
X0 VDD IN.t0 OUT.t2 VDD.t2 pfet_03v3 ad=0.616p pd=3.68u as=0.364p ps=1.92u w=1.4u l=0.35u
X1 VSS IN.t1 OUT.t3 VSS.t2 nfet_03v3 ad=0.308p pd=2.28u as=0.182p ps=1.22u w=0.7u l=0.35u
X2 OUT IN.t2 VDD.t1 VDD.t0 pfet_03v3 ad=0.364p pd=1.92u as=0.616p ps=3.68u w=1.4u l=0.35u
X3 OUT IN.t3 VSS.t1 VSS.t0 nfet_03v3 ad=0.182p pd=1.22u as=0.308p ps=2.28u w=0.7u l=0.35u
R0 IN.n0 IN.t0 21.9005
R1 IN.n1 IN.t2 20.5448
R2 IN.n1 IN.n0 16.59
R3 IN.n0 IN.t1 14.9134
R4 IN.n1 IN.t3 13.9748
R5 IN IN.n1 9.21196
R6 OUT.n4 OUT.n3 3.44007
R7 OUT.n4 OUT.n1 3.05441
R8 OUT.n3 OUT.t3 2.3405
R9 OUT.n3 OUT.n2 2.3405
R10 OUT.n1 OUT.t2 1.3005
R11 OUT.n1 OUT.n0 1.3005
R12 OUT OUT.n4 0.335065
R13 VDD.n8 VDD.t0 39.8225
R14 VDD.n2 VDD.t2 9.67173
R15 VDD.n11 VDD.t1 4.3192
R16 VDD.n1 VDD.n0 4.3192
R17 VDD.n4 VDD.n3 3.1505
R18 VDD.n7 VDD.n6 3.1505
R19 VDD.n6 VDD.n5 3.1505
R20 VDD.n10 VDD.n9 3.1505
R21 VDD.n3 VDD.n2 0.125861
R22 VDD.n9 VDD.n8 0.125617
R23 VDD.n7 VDD.n4 0.102773
R24 VDD.n10 VDD.n7 0.102773
R25 VDD.n4 VDD.n1 0.0853864
R26 VDD VDD.n10 0.0526591
R27 VDD VDD.n11 0.0148182
R28 VSS.n46 VSS.n45 548.402
R29 VSS.n86 VSS.t0 342.526
R30 VSS.n8 VSS.n7 337.918
R31 VSS.n38 VSS.t2 262.868
R32 VSS.n75 VSS.n74 135.417
R33 VSS.n28 VSS.n27 95.5887
R34 VSS.n85 VSS.t1 5.80213
R35 VSS.n37 VSS.n0 5.80209
R36 VSS.n56 VSS.n46 2.60441
R37 VSS.n81 VSS.n80 2.60148
R38 VSS.n62 VSS.n61 2.6005
R39 VSS.n61 VSS.n60 2.6005
R40 VSS.n65 VSS.n64 2.6005
R41 VSS.n64 VSS.n63 2.6005
R42 VSS.n68 VSS.n67 2.6005
R43 VSS.n67 VSS.n66 2.6005
R44 VSS.n71 VSS.n70 2.6005
R45 VSS.n70 VSS.n69 2.6005
R46 VSS.n73 VSS.n72 2.6005
R47 VSS.n78 VSS.n77 2.6005
R48 VSS.n59 VSS.n58 2.6005
R49 VSS.n58 VSS.n57 2.6005
R50 VSS.n9 VSS.n8 2.6005
R51 VSS.n6 VSS.n5 2.6005
R52 VSS.n5 VSS.n4 2.6005
R53 VSS.n3 VSS.n2 2.6005
R54 VSS.n2 VSS.n1 2.6005
R55 VSS.n49 VSS.n48 2.6005
R56 VSS.n48 VSS.n47 2.6005
R57 VSS.n52 VSS.n51 2.6005
R58 VSS.n51 VSS.n50 2.6005
R59 VSS.n55 VSS.n54 2.6005
R60 VSS.n54 VSS.n53 2.6005
R61 VSS.n31 VSS.n30 2.6005
R62 VSS.n26 VSS.n25 2.6005
R63 VSS.n24 VSS.n23 2.6005
R64 VSS.n23 VSS.n22 2.6005
R65 VSS.n21 VSS.n20 2.6005
R66 VSS.n20 VSS.n19 2.6005
R67 VSS.n18 VSS.n17 2.6005
R68 VSS.n17 VSS.n16 2.6005
R69 VSS.n15 VSS.n14 2.6005
R70 VSS.n14 VSS.n13 2.6005
R71 VSS.n12 VSS.n11 2.6005
R72 VSS.n11 VSS.n10 2.6005
R73 VSS.n36 VSS.n35 2.6005
R74 VSS.n35 VSS.n34 2.6005
R75 VSS.n40 VSS.n39 2.6005
R76 VSS.n39 VSS.n38 2.6005
R77 VSS.n43 VSS.n42 2.6005
R78 VSS.n42 VSS.n41 2.6005
R79 VSS.n88 VSS.n87 2.6005
R80 VSS.n87 VSS.n86 2.6005
R81 VSS.n84 VSS.n83 2.6005
R82 VSS.n83 VSS.n82 2.6005
R83 VSS.n33 VSS.n32 2.6005
R84 VSS.n30 VSS.n29 1.74053
R85 VSS.n77 VSS.n76 1.72725
R86 VSS.n76 VSS.n75 0.438169
R87 VSS.n29 VSS.n28 0.431816
R88 VSS.n46 VSS.n44 0.304848
R89 VSS.n15 VSS.n12 0.1355
R90 VSS.n18 VSS.n15 0.1355
R91 VSS.n21 VSS.n18 0.1355
R92 VSS.n24 VSS.n21 0.1355
R93 VSS.n26 VSS.n24 0.1355
R94 VSS.n31 VSS.n26 0.1355
R95 VSS.n62 VSS.n59 0.132565
R96 VSS.n65 VSS.n62 0.132565
R97 VSS.n68 VSS.n65 0.132565
R98 VSS.n71 VSS.n68 0.132565
R99 VSS.n73 VSS.n71 0.132565
R100 VSS.n78 VSS.n73 0.132565
R101 VSS.n59 VSS.n56 0.128652
R102 VSS.n9 VSS.n6 0.1255
R103 VSS.n6 VSS.n3 0.1255
R104 VSS.n52 VSS.n49 0.1255
R105 VSS.n55 VSS.n52 0.1255
R106 VSS.n36 VSS.n33 0.1255
R107 VSS.n43 VSS.n40 0.1255
R108 VSS.n81 VSS.n78 0.0983261
R109 VSS.n33 VSS.n31 0.0945
R110 VSS.n56 VSS.n55 0.0815
R111 VSS.n85 VSS.n84 0.0815
R112 VSS.n84 VSS.n81 0.0805
R113 VSS.n80 VSS.n79 0.076587
R114 VSS.n37 VSS.n36 0.0725
R115 VSS VSS.n88 0.0655
R116 VSS VSS.n43 0.0605
R117 VSS.n12 VSS.n9 0.0565
R118 VSS.n40 VSS.n37 0.0535
R119 VSS.n88 VSS.n85 0.0445
C0 VDD OUT 0.286f
C1 IN VDD 0.358f
C2 IN OUT 0.118f
.ends

