* NGSPICE file created from CLK_DIV_11_mag_new_flat.ext - technology: gf180mcuC

.subckt CLK_DIV_11_mag_new_flat VSS RST CLK Vdiv11 Q2 Q1 Q0 Q3 VDD
X0 VDD CLK.t0 JK_FF_mag_1.nand3_mag_2.OUT VDD.t37 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1 a_6046_4917# CLK.t1 a_5886_4917# VSS.t22 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2 JK_FF_mag_3.nand3_mag_2.OUT JK_FF_mag_3.K.t2 VDD.t214 VDD.t213 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X3 JK_FF_mag_3.QB JK_FF_mag_3.nand2_mag_4.IN2 VDD.t77 VDD.t76 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X4 and2_mag_3.OUT and2_mag_3.GF_INV_MAG_0.IN VDD.t1 VDD.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X5 JK_FF_mag_1.nand3_mag_2.OUT JK_FF_mag_1.K.t2 VDD.t216 VDD.t215 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X6 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.K VDD.t224 VDD.t223 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X7 JK_FF_mag_1.QB JK_FF_mag_1.nand2_mag_4.IN2 VDD.t128 VDD.t127 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X8 a_2751_4915# JK_FF_mag_0.K VSS.t153 VSS.t152 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X9 a_5886_4917# JK_FF_mag_1.K.t3 VSS.t1 VSS.t0 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X10 a_7898_4917# JK_FF_mag_1.nand2_mag_4.IN2 VSS.t90 VSS.t89 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X11 JK_FF_mag_1.nand3_mag_2.OUT Q2.t3 VDD.t240 VDD.t239 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X12 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand3_mag_2.OUT VDD.t156 VDD.t155 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X13 and2_mag_3.GF_INV_MAG_0.IN Q1.t3 VDD.t193 VDD.t192 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X14 JK_FF_mag_1.nand3_mag_2.OUT Q2.t4 a_6046_4917# VSS.t107 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X15 a_8344_1618# Q1.t4 VSS.t47 VSS.t46 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X16 a_6610_4917# JK_FF_mag_1.nand3_mag_2.OUT VSS.t111 VSS.t110 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X17 JK_FF_mag_1.nand2_mag_4.IN2 JK_FF_mag_1.nand3_mag_1.OUT VDD.t238 VDD.t237 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X18 VDD Q1.t5 and2_mag_1.GF_INV_MAG_0.IN VDD.t208 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X19 Q0 JK_FF_mag_3.nand2_mag_1.IN2 VDD.t233 VDD.t232 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X20 a_14017_3822# JK_FF_mag_3.nand2_mag_1.IN2 VSS.t157 VSS.t156 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X21 a_7334_4917# JK_FF_mag_1.nand3_mag_1.OUT VSS.t159 VSS.t158 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X22 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand3_mag_1.OUT VDD.t122 VDD.t121 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X23 JK_FF_mag_2.K or_2_mag_1.GF_INV_MAG_1.IN VDD.t167 VDD.t166 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X24 a_4199_4915# JK_FF_mag_0.nand3_mag_1.OUT VSS.t85 VSS.t84 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X25 VDD Q2.t5 JK_FF_mag_1.QB VDD.t110 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X26 JK_FF_mag_3.nand2_mag_1.IN2 JK_FF_mag_3.nand3_mag_1.IN1 VDD.t146 VDD.t145 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X27 a_13453_3822# JK_FF_mag_3.nand3_mag_1.IN1 VSS.t102 VSS.t101 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X28 JK_FF_mag_1.QB Q2.t6 a_7898_4917# VSS.t57 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X29 and2_mag_1.GF_INV_MAG_0.IN Q0.t3 VDD.t5 VDD.t4 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X30 or_2_mag_0.IN1 and2_mag_0.GF_INV_MAG_0.IN VDD.t53 VDD.t52 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X31 VDD JK_FF_mag_3.QB Q0.t1 VDD.t102 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X32 VDD CLK.t2 JK_FF_mag_1.nand3_mag_0.OUT VDD.t34 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X33 Q0 JK_FF_mag_3.QB a_14017_3822# VSS.t77 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X34 Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN Q2.t7 VDD.t197 VDD.t196 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X35 a_6052_3820# CLK.t3 a_5892_3820# VSS.t21 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X36 JK_FF_mag_0.K or_2_mag_0.GF_INV_MAG_1.IN VDD.t49 VDD.t48 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X37 VDD JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand3_mag_1.IN1 VDD.t234 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X38 a_2849_1480# or_2_mag_3.IN2 VDD.t165 VDD.t164 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X39 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand3_mag_1.OUT a_6616_3820# VSS.t87 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X40 JK_FF_mag_1.nand2_mag_3.IN1 CLK.t4 VDD.t33 VDD.t32 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X41 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_1.K.t4 VDD.t88 VDD.t87 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X42 a_11241_1205# and2_mag_3.OUT a_11081_1205# VDD.t40 pfet_03v3 ad=0.624p pd=2.92u as=0.624p ps=2.92u w=2.4u l=0.28u
X43 VDD JK_FF_mag_1.QB Q2.t1 VDD.t227 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X44 a_5892_3820# JK_FF_mag_1.K.t5 VSS.t104 VSS.t21 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X45 Q2 JK_FF_mag_1.QB a_7744_3820# VSS.t87 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X46 Q3 JK_FF_mag_0.nand2_mag_1.IN2 VDD.t264 VDD.t263 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X47 Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN Q2.t8 VSS.t49 VSS.t48 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X48 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_1.QB VDD.t226 VDD.t225 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X49 a_4609_3818# JK_FF_mag_0.nand2_mag_1.IN2 VSS.t170 VSS.t169 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X50 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_1.QB a_6052_3820# VSS.t21 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X51 a_11081_1205# nor_3_mag_0.IN3 VDD.t195 VDD.t194 pfet_03v3 ad=0.624p pd=2.92u as=1.06p ps=5.68u w=2.4u l=0.28u
X52 VSS or_2_mag_3.IN1.t3 or_2_mag_3.GF_INV_MAG_1.IN VSS.t52 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X53 JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_2.nand3_mag_1.IN1 VDD.t247 VDD.t246 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X54 JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_2.nand3_mag_1.IN1 a_9884_4915# VSS.t163 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X55 VDD Q0.t4 nand3_mag_0.OUT VDD.t68 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X56 JK_FF_mag_0.nand2_mag_3.IN1 CLK.t5 VSS.t20 VSS.t19 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X57 JK_FF_mag_1.nand2_mag_3.IN1 CLK.t6 VSS.t18 VSS.t17 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X58 or_2_mag_0.IN1 and2_mag_0.GF_INV_MAG_0.IN VSS.t36 VSS.t35 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X59 VDD RST.t0 JK_FF_mag_2.nand3_mag_1.OUT VDD.t78 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X60 a_9884_4915# RST.t1 a_9724_4915# VSS.t125 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X61 JK_FF_mag_0.K or_2_mag_0.GF_INV_MAG_1.IN VSS.t32 VSS.t31 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X62 nand3_mag_0.OUT Q2.t9 VDD.t45 VDD.t44 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X63 or_2_mag_3.GF_INV_MAG_1.IN or_2_mag_3.IN2 VSS.t116 VSS.t52 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X64 or_2_mag_0.GF_INV_MAG_1.IN or_2_mag_0.IN1 a_939_3715# VDD.t172 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X65 Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN GF_INV_MAG_1.OUT VDD.t169 VDD.t168 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X66 or_2_mag_1.IN1 and2_mag_2.GF_INV_MAG_0.IN VDD.t43 VDD.t42 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X67 or_2_mag_0.IN2 nand3_mag_0.OUT VDD.t152 VDD.t151 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X68 nand3_mag_0.OUT Q1.t6 VDD.t242 VDD.t241 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X69 VDD JK_FF_mag_2.nand2_mag_3.IN1 JK_FF_mag_2.nand2_mag_4.IN2 VDD.t254 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X70 JK_FF_mag_1.K and2_mag_1.GF_INV_MAG_0.IN VDD.t218 VDD.t217 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X71 VDD JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_2.nand3_mag_1.IN1 VDD.t115 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X72 JK_FF_mag_2.nand2_mag_4.IN2 JK_FF_mag_2.nand2_mag_3.IN1 a_10448_4915# VSS.t165 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X73 or_2_mag_3.IN1 JK_FF_mag_2.nand2_mag_4.IN2 VDD.t51 VDD.t50 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X74 JK_FF_mag_2.nand3_mag_1.IN1 JK_FF_mag_2.nand3_mag_1.OUT a_9730_3818# VSS.t82 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X75 JK_FF_mag_2.nand2_mag_3.IN1 CLK.t7 VDD.t31 VDD.t30 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X76 a_11012_4915# JK_FF_mag_2.nand2_mag_4.IN2 VSS.t34 VSS.t33 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X77 Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN GF_INV_MAG_1.OUT VSS.t120 VSS.t119 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X78 a_13043_4919# RST.t2 a_12883_4919# VSS.t75 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X79 VDD Q1.t7 or_2_mag_3.IN1.t1 VDD.t173 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X80 nand3_mag_1.OUT CLK.t8 VDD.t29 VDD.t28 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X81 and2_mag_3.OUT and2_mag_3.GF_INV_MAG_0.IN VSS.t3 VSS.t2 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X82 or_2_mag_3.IN1 Q1.t8 a_11012_4915# VSS.t166 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X83 JK_FF_mag_3.nand2_mag_4.IN2 JK_FF_mag_3.nand2_mag_3.IN1 a_13607_4919# VSS.t43 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X84 nand3_mag_1.OUT CLK.t9 a_7639_1615# VSS.t16 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X85 JK_FF_mag_3.nand3_mag_2.OUT Q0.t5 a_12319_4919# VSS.t136 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X86 a_12883_4919# JK_FF_mag_3.nand3_mag_2.OUT VSS.t5 VSS.t4 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X87 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand3_mag_1.IN1 a_13043_4919# VSS.t100 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X88 VDD or_2_mag_3.IN1.t4 Q1.t2 VDD.t198 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X89 Q1 or_2_mag_3.IN1.t5 a_10858_3818# VSS.t63 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X90 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand3_mag_0.OUT VDD.t205 VDD.t204 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X91 a_6616_3820# JK_FF_mag_1.nand3_mag_0.OUT VSS.t142 VSS.t87 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X92 VDD JK_FF_mag_2.nand2_mag_3.IN1 JK_FF_mag_2.nand2_mag_1.IN2 VDD.t251 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X93 JK_FF_mag_2.nand2_mag_1.IN2 JK_FF_mag_2.nand2_mag_3.IN1 a_10294_3818# VSS.t164 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X94 Q2 JK_FF_mag_1.nand2_mag_1.IN2 VDD.t148 VDD.t147 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X95 VDD JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.nand2_mag_1.IN2 VDD.t132 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X96 JK_FF_mag_1.nand2_mag_1.IN2 JK_FF_mag_1.nand2_mag_3.IN1 a_7180_3820# VSS.t87 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X97 a_7744_3820# JK_FF_mag_1.nand2_mag_1.IN2 VSS.t103 VSS.t87 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X98 or_2_mag_1.GF_INV_MAG_1.IN or_2_mag_1.IN1 a_1377_1477# VDD.t86 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X99 Q1 JK_FF_mag_2.nand2_mag_1.IN2 VDD.t158 VDD.t157 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X100 a_10858_3818# JK_FF_mag_2.nand2_mag_1.IN2 VSS.t113 VSS.t112 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X101 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.IN1 VDD.t187 VDD.t186 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X102 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.IN1 a_3635_4915# VSS.t131 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X103 JK_FF_mag_2.nand2_mag_1.IN2 JK_FF_mag_2.nand3_mag_1.IN1 VDD.t245 VDD.t244 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X104 JK_FF_mag_1.nand2_mag_1.IN2 JK_FF_mag_1.nand3_mag_1.IN1 VDD.t126 VDD.t125 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X105 a_10294_3818# JK_FF_mag_2.nand3_mag_1.IN1 VSS.t162 VSS.t161 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X106 JK_FF_mag_2.K or_2_mag_1.GF_INV_MAG_1.IN VSS.t118 VSS.t117 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X107 a_140_2787# Q0.t6 a_n20_2787# VSS.t28 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X108 a_7180_3820# JK_FF_mag_1.nand3_mag_1.IN1 VSS.t88 VSS.t87 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X109 a_1377_1477# Q0.t7 VDD.t90 VDD.t89 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X110 JK_FF_mag_3.nand2_mag_3.IN1 CLK.t10 VDD.t27 VDD.t26 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X111 JK_FF_mag_2.nand3_mag_2.OUT JK_FF_mag_2.K VDD.t142 VDD.t141 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X112 JK_FF_mag_3.nand3_mag_0.OUT JK_FF_mag_3.QB VDD.t101 VDD.t100 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X113 a_9000_4915# JK_FF_mag_2.K VSS.t99 VSS.t98 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X114 JK_FF_mag_2.nand3_mag_2.OUT Q1.t9 VDD.t94 VDD.t93 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X115 JK_FF_mag_3.nand3_mag_0.OUT JK_FF_mag_3.QB a_12325_3822# VSS.t76 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X116 JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_2.nand3_mag_2.OUT VDD.t207 VDD.t206 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X117 Vdiv11 nor_3_mag_0.OUT VDD.t171 VDD.t170 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X118 JK_FF_mag_2.nand3_mag_2.OUT Q1.t10 a_9160_4915# VSS.t72 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X119 a_9724_4915# JK_FF_mag_2.nand3_mag_2.OUT VSS.t144 VSS.t143 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X120 VSS or_2_mag_1.IN1 or_2_mag_1.GF_INV_MAG_1.IN VSS.t68 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X121 nand3_mag_0.OUT Q2.t10 a_140_2787# VSS.t28 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X122 VDD CLK.t11 JK_FF_mag_2.nand3_mag_2.OUT VDD.t23 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X123 JK_FF_mag_3.nand2_mag_3.IN1 CLK.t12 VSS.t15 VSS.t14 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X124 a_9160_4915# CLK.t13 a_9000_4915# VSS.t13 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X125 and2_mag_1.GF_INV_MAG_0.IN Q1.t11 a_1385_2540# VSS.t78 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X126 a_939_3715# or_2_mag_0.IN2 VDD.t67 VDD.t66 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X127 a_n20_2787# Q1.t12 VSS.t60 VSS.t28 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X128 JK_FF_mag_2.nand3_mag_0.OUT JK_FF_mag_2.K VDD.t140 VDD.t139 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X129 a_9006_3818# JK_FF_mag_2.K VSS.t97 VSS.t96 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X130 JK_FF_mag_2.nand2_mag_4.IN2 JK_FF_mag_2.nand3_mag_1.OUT VDD.t114 VDD.t113 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X131 JK_FF_mag_2.nand3_mag_1.IN1 JK_FF_mag_2.nand3_mag_0.OUT VDD.t220 VDD.t219 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X132 JK_FF_mag_2.nand3_mag_0.OUT or_2_mag_3.IN1.t6 VDD.t99 VDD.t98 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X133 a_10448_4915# JK_FF_mag_2.nand3_mag_1.OUT VSS.t81 VSS.t80 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X134 JK_FF_mag_2.nand3_mag_0.OUT or_2_mag_3.IN1.t7 a_9166_3818# VSS.t37 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X135 a_9730_3818# JK_FF_mag_2.nand3_mag_0.OUT VSS.t149 VSS.t148 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X136 or_2_mag_1.GF_INV_MAG_1.IN Q0.t8 VSS.t160 VSS.t68 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X137 a_1385_2540# Q0.t9 VSS.t145 VSS.t78 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X138 VDD CLK.t14 JK_FF_mag_2.nand3_mag_0.OUT VDD.t20 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X139 VDD RST.t3 JK_FF_mag_3.nand3_mag_1.OUT VDD.t248 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X140 a_9166_3818# CLK.t15 a_9006_3818# VSS.t12 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X141 VDD Q0.t10 nand3_mag_1.OUT VDD.t181 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X142 a_13607_4919# JK_FF_mag_3.nand3_mag_1.OUT VSS.t128 VSS.t127 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X143 VDD JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_3.nand2_mag_4.IN2 VDD.t60 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X144 and2_mag_3.IN1 Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VDD.t136 VDD.t135 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X145 a_7639_1615# Q0.t11 a_7479_1615# VSS.t79 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X146 a_12319_4919# CLK.t16 a_12159_4919# VSS.t11 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X147 JK_FF_mag_3.nand3_mag_2.OUT Q0.t12 VDD.t106 VDD.t105 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X148 GF_INV_MAG_1.OUT nand3_mag_1.OUT VDD.t138 VDD.t137 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X149 JK_FF_mag_3.QB Q0.t13 a_14171_4919# VSS.t71 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X150 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand3_mag_2.OUT VDD.t3 VDD.t2 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X151 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand3_mag_1.IN1 VDD.t144 VDD.t143 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X152 JK_FF_mag_2.nand2_mag_3.IN1 CLK.t17 VSS.t10 VSS.t9 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X153 VDD Q3.t3 and2_mag_2.GF_INV_MAG_0.IN VDD.t71 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X154 nand3_mag_1.OUT and2_mag_3.IN1 VDD.t85 VDD.t84 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X155 or_2_mag_1.IN1 and2_mag_2.GF_INV_MAG_0.IN VSS.t27 VSS.t26 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X156 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand3_mag_1.IN1 VDD.t124 VDD.t123 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X157 a_7479_1615# and2_mag_3.IN1 VSS.t66 VSS.t65 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X158 a_12159_4919# JK_FF_mag_3.K.t3 VSS.t51 VSS.t50 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X159 and2_mag_3.IN1 Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS.t93 VSS.t92 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X160 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand3_mag_1.IN1 a_6770_4917# VSS.t86 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X161 a_14171_4919# JK_FF_mag_3.nand2_mag_4.IN2 VSS.t59 VSS.t58 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X162 nor_3_mag_0.IN3 Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN VDD.t47 VDD.t46 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X163 VDD JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand3_mag_1.IN1 VDD.t178 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X164 VDD CLK.t18 JK_FF_mag_0.nand3_mag_2.OUT VDD.t17 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X165 GF_INV_MAG_1.OUT nand3_mag_1.OUT VSS.t95 VSS.t94 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X166 and2_mag_2.GF_INV_MAG_0.IN Q1.t13 VDD.t150 VDD.t149 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X167 JK_FF_mag_3.nand3_mag_1.IN1 JK_FF_mag_3.nand3_mag_1.OUT a_12889_3822# VSS.t126 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X168 a_2911_4915# CLK.t19 a_2751_4915# VSS.t8 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X169 VDD Q3.t4 or_2_mag_3.IN2 VDD.t63 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X170 VDD RST.t4 JK_FF_mag_1.nand3_mag_1.OUT VDD.t54 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X171 VDD and2_mag_3.IN1 and2_mag_3.GF_INV_MAG_0.IN VDD.t81 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X172 or_2_mag_3.IN2 Q3.t5 a_4763_4915# VSS.t62 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X173 VDD RST.t5 JK_FF_mag_0.nand3_mag_1.OUT VDD.t201 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X174 and2_mag_3.GF_INV_MAG_0.IN and2_mag_3.IN1 a_8344_1618# VSS.t64 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X175 and2_mag_2.GF_INV_MAG_0.IN Q3.t6 a_n27_2146# VSS.t134 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X176 a_3635_4915# RST.t6 a_3475_4915# VSS.t61 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X177 a_6770_4917# RST.t7 a_6610_4917# VSS.t137 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X178 VDD JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.nand2_mag_4.IN2 VDD.t129 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X179 VDD Q3.t7 and2_mag_0.GF_INV_MAG_0.IN VDD.t68 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X180 nor_3_mag_0.IN3 Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN VSS.t30 VSS.t29 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X181 nor_3_mag_0.OUT nor_3_mag_0.IN3 VSS.t139 VSS.t138 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X182 JK_FF_mag_3.nand3_mag_1.IN1 JK_FF_mag_3.nand3_mag_0.OUT VDD.t75 VDD.t74 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X183 JK_FF_mag_1.nand2_mag_4.IN2 JK_FF_mag_1.nand2_mag_3.IN1 a_7334_4917# VSS.t91 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X184 VDD JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand2_mag_4.IN2 VDD.t260 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X185 a_12889_3822# JK_FF_mag_3.nand3_mag_0.OUT VSS.t56 VSS.t55 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X186 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand2_mag_3.IN1 a_4199_4915# VSS.t168 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X187 JK_FF_mag_0.nand3_mag_2.OUT Q3.t8 VDD.t109 VDD.t108 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X188 or_2_mag_3.IN2 JK_FF_mag_0.nand2_mag_4.IN2 VDD.t191 VDD.t190 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X189 VDD JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_3.nand2_mag_1.IN2 VDD.t57 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X190 a_4763_4915# JK_FF_mag_0.nand2_mag_4.IN2 VSS.t133 VSS.t132 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X191 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_2.OUT VDD.t231 VDD.t230 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X192 VDD CLK.t20 JK_FF_mag_3.nand3_mag_0.OUT VDD.t14 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X193 JK_FF_mag_3.nand2_mag_1.IN2 JK_FF_mag_3.nand2_mag_3.IN1 a_13453_3822# VSS.t42 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X194 JK_FF_mag_0.nand3_mag_2.OUT Q3.t9 a_2911_4915# VSS.t67 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X195 a_3475_4915# JK_FF_mag_0.nand3_mag_2.OUT VSS.t155 VSS.t154 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X196 JK_FF_mag_3.K or_2_mag_3.GF_INV_MAG_1.IN VDD.t154 VDD.t153 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X197 a_n27_2146# Q1.t14 VSS.t135 VSS.t134 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X198 a_12325_3822# CLK.t21 a_12165_3822# VSS.t7 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X199 and2_mag_0.GF_INV_MAG_0.IN Q3.t10 a_n20_4333# VSS.t40 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X200 VDD CLK.t22 JK_FF_mag_0.nand3_mag_0.OUT VDD.t11 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X201 a_2917_3818# CLK.t23 a_2757_3818# VSS.t6 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X202 JK_FF_mag_3.nand3_mag_0.OUT JK_FF_mag_3.K.t4 VDD.t189 VDD.t188 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X203 VDD JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.IN1 VDD.t118 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X204 a_12165_3822# JK_FF_mag_3.K.t5 VSS.t39 VSS.t38 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X205 VSS or_2_mag_0.IN1 or_2_mag_0.GF_INV_MAG_1.IN VSS.t44 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X206 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand3_mag_1.OUT a_3481_3818# VSS.t83 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X207 JK_FF_mag_0.nand2_mag_3.IN1 CLK.t24 VDD.t10 VDD.t9 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X208 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_0.nand3_mag_1.IN1 VDD.t185 VDD.t184 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X209 or_2_mag_3.GF_INV_MAG_1.IN or_2_mag_3.IN1.t8 a_2849_1480# VDD.t107 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X210 or_2_mag_0.IN2 nand3_mag_0.OUT VSS.t106 VSS.t105 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X211 a_4045_3818# JK_FF_mag_0.nand3_mag_1.IN1 VSS.t130 VSS.t129 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X212 nor_3_mag_0.OUT Q3.t11 a_11241_1205# VDD.t41 pfet_03v3 ad=1.06p pd=5.68u as=0.624p ps=2.92u w=2.4u l=0.28u
X213 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.K VDD.t222 VDD.t221 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X214 nor_3_mag_0.OUT Q3.t12 VSS.t141 VSS.t140 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X215 and2_mag_0.GF_INV_MAG_0.IN Q1.t15 VDD.t243 VDD.t241 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X216 a_2757_3818# JK_FF_mag_0.K VSS.t151 VSS.t150 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X217 JK_FF_mag_0.nand3_mag_0.OUT or_2_mag_3.IN2 VDD.t163 VDD.t162 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X218 VDD or_2_mag_3.IN2 Q3.t1 VDD.t159 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X219 Q3 or_2_mag_3.IN2 a_4609_3818# VSS.t115 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X220 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand3_mag_0.OUT VDD.t92 VDD.t91 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X221 Vdiv11 nor_3_mag_0.OUT VSS.t122 VSS.t121 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X222 JK_FF_mag_0.nand3_mag_0.OUT or_2_mag_3.IN2 a_2917_3818# VSS.t114 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X223 a_3481_3818# JK_FF_mag_0.nand3_mag_0.OUT VSS.t74 VSS.t73 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X224 VDD JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand2_mag_1.IN2 VDD.t257 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X225 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_0.nand2_mag_3.IN1 a_4045_3818# VSS.t167 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X226 JK_FF_mag_3.K or_2_mag_3.GF_INV_MAG_1.IN VSS.t109 VSS.t108 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X227 JK_FF_mag_1.K and2_mag_1.GF_INV_MAG_0.IN VSS.t147 VSS.t146 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X228 a_n20_4333# Q1.t16 VSS.t41 VSS.t40 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X229 VSS and2_mag_3.OUT nor_3_mag_0.OUT VSS.t23 nfet_03v3 ad=86.8f pd=0.92u as=86.8f ps=0.92u w=0.22u l=0.28u
X230 JK_FF_mag_3.nand2_mag_4.IN2 JK_FF_mag_3.nand3_mag_1.OUT VDD.t177 VDD.t176 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X231 or_2_mag_0.GF_INV_MAG_1.IN or_2_mag_0.IN2 VSS.t45 VSS.t44 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X232 VDD CLK.t25 JK_FF_mag_3.nand3_mag_2.OUT VDD.t6 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X233 VDD Q0.t14 JK_FF_mag_3.QB VDD.t95 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
R0 CLK.n12 CLK.t3 36.935
R1 CLK.n6 CLK.t1 36.935
R2 CLK.n48 CLK.t15 36.935
R3 CLK.n42 CLK.t13 36.935
R4 CLK.n57 CLK.t9 36.935
R5 CLK.n30 CLK.t21 36.935
R6 CLK.n24 CLK.t16 36.935
R7 CLK.n72 CLK.t23 36.935
R8 CLK.n66 CLK.t19 36.935
R9 CLK.n77 CLK.t24 25.4742
R10 CLK.n38 CLK.t7 25.4742
R11 CLK.n2 CLK.t4 25.4739
R12 CLK.n20 CLK.t10 25.4739
R13 CLK.n12 CLK.t2 18.1962
R14 CLK.n6 CLK.t0 18.1962
R15 CLK.n48 CLK.t14 18.1962
R16 CLK.n42 CLK.t11 18.1962
R17 CLK.n57 CLK.t8 18.1962
R18 CLK.n30 CLK.t20 18.1962
R19 CLK.n24 CLK.t25 18.1962
R20 CLK.n72 CLK.t22 18.1962
R21 CLK.n66 CLK.t18 18.1962
R22 CLK.n77 CLK.t5 14.142
R23 CLK.n38 CLK.t17 14.142
R24 CLK.n2 CLK.t6 14.1414
R25 CLK.n20 CLK.t12 14.1414
R26 CLK.n62 CLK 5.77975
R27 CLK.n79 CLK.n63 5.11742
R28 CLK.n7 CLK.n4 4.5005
R29 CLK.n9 CLK.n8 4.5005
R30 CLK.n11 CLK.n10 4.5005
R31 CLK.n13 CLK.n10 4.5005
R32 CLK.n17 CLK.n3 4.5005
R33 CLK.n18 CLK.n17 4.5005
R34 CLK.n43 CLK.n40 4.5005
R35 CLK.n45 CLK.n44 4.5005
R36 CLK.n47 CLK.n46 4.5005
R37 CLK.n49 CLK.n46 4.5005
R38 CLK.n54 CLK.n53 4.5005
R39 CLK.n53 CLK.n39 4.5005
R40 CLK.n58 CLK.n55 4.5005
R41 CLK.n25 CLK.n22 4.5005
R42 CLK.n27 CLK.n26 4.5005
R43 CLK.n29 CLK.n28 4.5005
R44 CLK.n31 CLK.n28 4.5005
R45 CLK.n35 CLK.n21 4.5005
R46 CLK.n36 CLK.n35 4.5005
R47 CLK.n69 CLK.n68 4.5005
R48 CLK.n67 CLK.n64 4.5005
R49 CLK.n71 CLK.n70 4.5005
R50 CLK.n73 CLK.n70 4.5005
R51 CLK.n79 CLK.n78 4.5005
R52 CLK.n80 CLK.n79 4.5005
R53 CLK.n63 CLK 4.43115
R54 CLK.n82 CLK 4.16645
R55 CLK.n61 CLK.n60 4.05271
R56 CLK.n62 CLK.n61 3.52625
R57 CLK.n61 CLK 2.3355
R58 CLK.n82 CLK.n81 2.25561
R59 CLK.n51 CLK.n50 2.25147
R60 CLK.n75 CLK.n74 2.25147
R61 CLK.n15 CLK.n14 2.25107
R62 CLK.n33 CLK.n32 2.25107
R63 CLK.n56 CLK.n55 2.24785
R64 CLK.n60 CLK.n59 2.24572
R65 CLK.n16 CLK.n1 2.24196
R66 CLK.n52 CLK.n37 2.24196
R67 CLK.n34 CLK.n19 2.24196
R68 CLK.n76 CLK.n0 2.24196
R69 CLK.n58 CLK.n57 2.12226
R70 CLK.n13 CLK.n12 2.12175
R71 CLK.n7 CLK.n6 2.12175
R72 CLK.n49 CLK.n48 2.12175
R73 CLK.n43 CLK.n42 2.12175
R74 CLK.n31 CLK.n30 2.12175
R75 CLK.n25 CLK.n24 2.12175
R76 CLK.n73 CLK.n72 2.12175
R77 CLK.n67 CLK.n66 2.12075
R78 CLK.n10 CLK.n9 1.71671
R79 CLK.n28 CLK.n27 1.71671
R80 CLK.n46 CLK.n45 1.71071
R81 CLK.n70 CLK.n69 1.71071
R82 CLK.n63 CLK.n62 1.62531
R83 CLK.n5 CLK.n4 1.49782
R84 CLK.n41 CLK.n40 1.49782
R85 CLK.n23 CLK.n22 1.49782
R86 CLK.n65 CLK.n64 1.49782
R87 CLK.n3 CLK.n2 1.4219
R88 CLK.n21 CLK.n20 1.4219
R89 CLK.n39 CLK.n38 1.42126
R90 CLK.n78 CLK.n77 1.42126
R91 CLK.n16 CLK.n15 0.970654
R92 CLK.n34 CLK.n33 0.970654
R93 CLK.n52 CLK.n51 0.968731
R94 CLK.n76 CLK.n75 0.968731
R95 CLK CLK.n18 0.1605
R96 CLK CLK.n54 0.1605
R97 CLK CLK.n36 0.1605
R98 CLK CLK.n80 0.1605
R99 CLK.n5 CLK 0.0714821
R100 CLK.n41 CLK 0.0714821
R101 CLK.n23 CLK 0.0714821
R102 CLK.n65 CLK 0.0714821
R103 CLK.n56 CLK 0.0529963
R104 CLK.n11 CLK 0.0473512
R105 CLK.n47 CLK 0.0473512
R106 CLK.n29 CLK 0.0473512
R107 CLK.n71 CLK 0.0473512
R108 CLK.n9 CLK.n4 0.0386356
R109 CLK.n45 CLK.n40 0.0386356
R110 CLK.n27 CLK.n22 0.0386356
R111 CLK.n69 CLK.n64 0.0386356
R112 CLK.n14 CLK.n11 0.0361897
R113 CLK.n50 CLK.n47 0.0361897
R114 CLK.n32 CLK.n29 0.0361897
R115 CLK.n74 CLK.n71 0.0361897
R116 CLK.n18 CLK.n1 0.03175
R117 CLK.n54 CLK.n37 0.03175
R118 CLK.n36 CLK.n19 0.03175
R119 CLK.n80 CLK.n0 0.03175
R120 CLK.n17 CLK.n16 0.0238218
R121 CLK.n53 CLK.n52 0.0238218
R122 CLK.n35 CLK.n34 0.0238218
R123 CLK.n79 CLK.n76 0.0238218
R124 CLK.n59 CLK.n58 0.0210263
R125 CLK.n59 CLK.n56 0.0183441
R126 CLK.n8 CLK.n5 0.0128713
R127 CLK.n44 CLK.n41 0.0128713
R128 CLK.n26 CLK.n23 0.0128713
R129 CLK.n68 CLK.n65 0.0128713
R130 CLK.n60 CLK.n55 0.0124457
R131 CLK.n15 CLK.n10 0.0122182
R132 CLK.n33 CLK.n28 0.0122182
R133 CLK.n51 CLK.n46 0.00986143
R134 CLK.n75 CLK.n70 0.00986143
R135 CLK CLK.n82 0.00567241
R136 CLK.n14 CLK.n13 0.00515517
R137 CLK.n8 CLK.n7 0.00515517
R138 CLK.n50 CLK.n49 0.00515517
R139 CLK.n44 CLK.n43 0.00515517
R140 CLK.n32 CLK.n31 0.00515517
R141 CLK.n26 CLK.n25 0.00515517
R142 CLK.n74 CLK.n73 0.00515517
R143 CLK.n68 CLK.n67 0.00515517
R144 CLK.n3 CLK.n1 0.00175
R145 CLK.n39 CLK.n37 0.00175
R146 CLK.n21 CLK.n19 0.00175
R147 CLK.n78 CLK.n0 0.00175
R148 VDD.t223 VDD.n175 57397.6
R149 VDD.t141 VDD.n78 57397.6
R150 VDD.n19 VDD.t194 3502.08
R151 VDD.n31 VDD.t135 1105.93
R152 VDD.n22 VDD.t46 1105.93
R153 VDD.t41 VDD.n13 1011.51
R154 VDD.t260 VDD.t190 961.905
R155 VDD.t108 VDD.t230 961.905
R156 VDD.t254 VDD.t50 961.905
R157 VDD.t93 VDD.t206 961.905
R158 VDD.n175 VDD.t121 864.287
R159 VDD.n78 VDD.t113 864.287
R160 VDD.n25 VDD.t81 857.144
R161 VDD.t132 VDD.t147 765.152
R162 VDD.t125 VDD.t234 765.152
R163 VDD.t225 VDD.t204 765.152
R164 VDD.t257 VDD.t263 765.152
R165 VDD.t118 VDD.t184 765.152
R166 VDD.t162 VDD.t91 765.152
R167 VDD.t157 VDD.t251 765.152
R168 VDD.t115 VDD.t244 765.152
R169 VDD.t219 VDD.t98 765.152
R170 VDD.t232 VDD.t57 765.152
R171 VDD.t178 VDD.t145 765.152
R172 VDD.t74 VDD.t100 765.152
R173 VDD.t60 VDD.t76 765.152
R174 VDD.t143 VDD.t176 765.152
R175 VDD.t105 VDD.t2 765.152
R176 VDD.t129 VDD.t127 765.152
R177 VDD.t123 VDD.t237 765.152
R178 VDD.t239 VDD.t155 765.152
R179 VDD.n23 VDD.t168 581.375
R180 VDD VDD.n23 569.634
R181 VDD.n220 VDD.t151 480.199
R182 VDD VDD.n165 426.699
R183 VDD VDD.n150 426.699
R184 VDD VDD.n133 426.699
R185 VDD.n253 VDD 424.618
R186 VDD.n213 VDD 424.618
R187 VDD.n249 VDD 424.618
R188 VDD.n258 VDD 422.557
R189 VDD.n13 VDD.t170 420.793
R190 VDD.n165 VDD.t87 386.365
R191 VDD.n197 VDD.t221 386.365
R192 VDD.n150 VDD.t139 386.365
R193 VDD.n133 VDD.t188 386.365
R194 VDD.t186 VDD.t201 380.952
R195 VDD.t17 VDD.t108 380.952
R196 VDD.t246 VDD.t78 380.952
R197 VDD.t23 VDD.t93 380.952
R198 VDD.t71 VDD.n258 378.788
R199 VDD.t208 VDD.n201 375
R200 VDD.n198 VDD.n197 365.673
R201 VDD.n201 VDD.n199 343.137
R202 VDD.t86 VDD.n253 309.341
R203 VDD.t107 VDD.n249 309.341
R204 VDD.t172 VDD.n213 306.118
R205 VDD.t34 VDD.t225 303.031
R206 VDD.t11 VDD.t162 303.031
R207 VDD.t98 VDD.t20 303.031
R208 VDD.t100 VDD.t14 303.031
R209 VDD.t248 VDD.t143 303.031
R210 VDD.t6 VDD.t105 303.031
R211 VDD.t54 VDD.t123 303.031
R212 VDD.t37 VDD.t239 303.031
R213 VDD.t181 VDD.t28 303.031
R214 VDD.n216 VDD.n204 298.536
R215 VDD.n220 VDD.n204 288
R216 VDD.n167 VDD.t63 242.857
R217 VDD.n169 VDD.t260 242.857
R218 VDD.t201 VDD.n172 242.857
R219 VDD.n176 VDD.t17 242.857
R220 VDD.n70 VDD.t173 242.857
R221 VDD.n72 VDD.t254 242.857
R222 VDD.t78 VDD.n75 242.857
R223 VDD.n79 VDD.t23 242.857
R224 VDD.t81 VDD.n24 217.337
R225 VDD.n259 VDD.t71 193.183
R226 VDD.n156 VDD.t227 193.183
R227 VDD.n157 VDD.t132 193.183
R228 VDD.n163 VDD.t234 193.183
R229 VDD.n164 VDD.t34 193.183
R230 VDD.n189 VDD.t159 193.183
R231 VDD.n191 VDD.t257 193.183
R232 VDD.n193 VDD.t118 193.183
R233 VDD.n196 VDD.t11 193.183
R234 VDD.n202 VDD.t208 193.183
R235 VDD.n137 VDD.t198 193.183
R236 VDD.n143 VDD.t251 193.183
R237 VDD.n144 VDD.t115 193.183
R238 VDD.n149 VDD.t20 193.183
R239 VDD.n120 VDD.t102 193.183
R240 VDD.n126 VDD.t57 193.183
R241 VDD.n127 VDD.t178 193.183
R242 VDD.n132 VDD.t14 193.183
R243 VDD.n99 VDD.t95 193.183
R244 VDD.n101 VDD.t60 193.183
R245 VDD.n104 VDD.t248 193.183
R246 VDD.n107 VDD.t6 193.183
R247 VDD.n42 VDD.t110 193.183
R248 VDD.n44 VDD.t129 193.183
R249 VDD.n47 VDD.t54 193.183
R250 VDD.n50 VDD.t37 193.183
R251 VDD.n3 VDD.t181 193.183
R252 VDD.n215 VDD.t44 191.288
R253 VDD.t40 VDD.t41 175.631
R254 VDD.t194 VDD.n18 153.678
R255 VDD.t44 VDD.t68 151.516
R256 VDD.t190 VDD.n167 138.095
R257 VDD.t121 VDD.n169 138.095
R258 VDD.t230 VDD.n172 138.095
R259 VDD.n176 VDD.t223 138.095
R260 VDD.t50 VDD.n70 138.095
R261 VDD.t113 VDD.n72 138.095
R262 VDD.t206 VDD.n75 138.095
R263 VDD.n79 VDD.t141 138.095
R264 VDD.n254 VDD.t86 137.826
R265 VDD.n250 VDD.t107 137.826
R266 VDD.n201 VDD.t217 132.353
R267 VDD.n212 VDD.t52 124.511
R268 VDD.n24 VDD.t192 123.258
R269 VDD.n216 VDD.n215 115.385
R270 VDD.n199 VDD.n198 112.746
R271 VDD.n259 VDD.t149 109.849
R272 VDD.t147 VDD.n156 109.849
R273 VDD.n157 VDD.t125 109.849
R274 VDD.t204 VDD.n163 109.849
R275 VDD.t87 VDD.n164 109.849
R276 VDD.t263 VDD.n189 109.849
R277 VDD.t184 VDD.n191 109.849
R278 VDD.t91 VDD.n193 109.849
R279 VDD.t221 VDD.n196 109.849
R280 VDD.n202 VDD.t4 109.849
R281 VDD.n137 VDD.t157 109.849
R282 VDD.t244 VDD.n143 109.849
R283 VDD.n144 VDD.t219 109.849
R284 VDD.t139 VDD.n149 109.849
R285 VDD.n120 VDD.t232 109.849
R286 VDD.t145 VDD.n126 109.849
R287 VDD.n127 VDD.t74 109.849
R288 VDD.t188 VDD.n132 109.849
R289 VDD.t76 VDD.n99 109.849
R290 VDD.t176 VDD.n101 109.849
R291 VDD.t2 VDD.n104 109.849
R292 VDD.n107 VDD.t213 109.849
R293 VDD.t127 VDD.n42 109.849
R294 VDD.t237 VDD.n44 109.849
R295 VDD.t155 VDD.n47 109.849
R296 VDD.n50 VDD.t215 109.849
R297 VDD.n3 VDD.t84 109.849
R298 VDD.n254 VDD.t89 107.198
R299 VDD.n250 VDD.t164 107.198
R300 VDD.n175 VDD.t186 97.6195
R301 VDD.n78 VDD.t246 97.6195
R302 VDD.t68 VDD.n211 96.5914
R303 VDD.n214 VDD.n212 90.2261
R304 VDD.n23 VDD.t137 83.3338
R305 VDD.n214 VDD.t172 76.2337
R306 VDD.n13 VDD 65.7064
R307 VDD.n165 VDD.t32 62.1896
R308 VDD.n197 VDD.t9 62.1896
R309 VDD.n150 VDD.t30 62.1896
R310 VDD.n133 VDD.t26 62.1896
R311 VDD.n253 VDD.t166 61.8817
R312 VDD.n213 VDD.t48 61.8817
R313 VDD.n249 VDD.t153 61.8817
R314 VDD.n258 VDD.t42 61.5769
R315 VDD.t135 VDD 61.3852
R316 VDD VDD.n198 61.0269
R317 VDD.n31 VDD.t196 55.0852
R318 VDD.n19 VDD.t46 55.0852
R319 VDD.t168 VDD.n22 55.0852
R320 VDD.n211 VDD.t241 54.9247
R321 VDD.n215 VDD.n214 21.9785
R322 VDD.n18 VDD.t40 21.9544
R323 VDD.n9 VDD.t169 14.0055
R324 VDD.n0 VDD.t136 12.3869
R325 VDD.n10 VDD.t47 12.3869
R326 VDD.n9 VDD.t138 10.1341
R327 VDD.n218 VDD.n217 9.64171
R328 VDD.n16 VDD.n15 7.9205
R329 VDD.n219 VDD.n218 6.69176
R330 VDD.n24 VDD.n7 6.40987
R331 VDD.n260 VDD.n259 6.3005
R332 VDD.n263 VDD.n254 6.3005
R333 VDD VDD.n220 6.3005
R334 VDD.n222 VDD.n204 6.3005
R335 VDD VDD.n216 6.3005
R336 VDD.n225 VDD.n202 6.3005
R337 VDD VDD.n199 6.3005
R338 VDD.n177 VDD.n176 6.3005
R339 VDD.n180 VDD.n172 6.3005
R340 VDD.n183 VDD.n169 6.3005
R341 VDD.n186 VDD.n167 6.3005
R342 VDD.n230 VDD.n196 6.3005
R343 VDD.n233 VDD.n193 6.3005
R344 VDD.n236 VDD.n191 6.3005
R345 VDD.n239 VDD.n189 6.3005
R346 VDD.n117 VDD.n99 6.3005
R347 VDD.n114 VDD.n101 6.3005
R348 VDD.n111 VDD.n104 6.3005
R349 VDD.n108 VDD.n107 6.3005
R350 VDD.n121 VDD.n120 6.3005
R351 VDD.n126 VDD.n125 6.3005
R352 VDD.n128 VDD.n127 6.3005
R353 VDD.n132 VDD.n131 6.3005
R354 VDD.n89 VDD.n70 6.3005
R355 VDD.n86 VDD.n72 6.3005
R356 VDD.n83 VDD.n75 6.3005
R357 VDD.n80 VDD.n79 6.3005
R358 VDD.n138 VDD.n137 6.3005
R359 VDD.n143 VDD.n142 6.3005
R360 VDD.n145 VDD.n144 6.3005
R361 VDD.n149 VDD.n148 6.3005
R362 VDD.n60 VDD.n42 6.3005
R363 VDD.n57 VDD.n44 6.3005
R364 VDD.n54 VDD.n47 6.3005
R365 VDD.n51 VDD.n50 6.3005
R366 VDD.n156 VDD.n155 6.3005
R367 VDD.n158 VDD.n157 6.3005
R368 VDD.n163 VDD.n162 6.3005
R369 VDD.n244 VDD.n164 6.3005
R370 VDD.n18 VDD.n17 6.3005
R371 VDD VDD.n19 6.3005
R372 VDD.n22 VDD.n21 6.3005
R373 VDD VDD.n25 6.3005
R374 VDD.n4 VDD.n3 6.3005
R375 VDD.n32 VDD.n31 6.3005
R376 VDD.n251 VDD.n250 6.3005
R377 VDD.n227 VDD.t218 5.85907
R378 VDD.n246 VDD.n245 5.69603
R379 VDD VDD.t193 5.26433
R380 VDD.n177 VDD.t224 5.213
R381 VDD.n108 VDD.t214 5.213
R382 VDD.n80 VDD.t142 5.213
R383 VDD.n51 VDD.t216 5.213
R384 VDD.n30 VDD.t85 5.16519
R385 VDD.n224 VDD.t5 5.15377
R386 VDD.n256 VDD.n255 5.13287
R387 VDD.n261 VDD.t150 5.13287
R388 VDD.n208 VDD.n205 5.13287
R389 VDD.n209 VDD.t243 5.13287
R390 VDD.n209 VDD.t242 5.13287
R391 VDD.n226 VDD.n200 5.13287
R392 VDD.n187 VDD.n166 5.13287
R393 VDD.n185 VDD.t191 5.13287
R394 VDD.n184 VDD.n168 5.13287
R395 VDD.n182 VDD.t122 5.13287
R396 VDD.n179 VDD.t231 5.13287
R397 VDD.n240 VDD.n188 5.13287
R398 VDD.n238 VDD.t264 5.13287
R399 VDD.n237 VDD.n190 5.13287
R400 VDD.n235 VDD.t185 5.13287
R401 VDD.n234 VDD.n192 5.13287
R402 VDD.n232 VDD.t92 5.13287
R403 VDD.n229 VDD.t222 5.13287
R404 VDD.n118 VDD.n98 5.13287
R405 VDD.n116 VDD.t77 5.13287
R406 VDD.n115 VDD.n100 5.13287
R407 VDD.n113 VDD.t177 5.13287
R408 VDD.n110 VDD.t3 5.13287
R409 VDD.n119 VDD.n97 5.13287
R410 VDD.n122 VDD.t233 5.13287
R411 VDD.n123 VDD.n96 5.13287
R412 VDD.n124 VDD.t146 5.13287
R413 VDD.n95 VDD.n94 5.13287
R414 VDD.n129 VDD.t75 5.13287
R415 VDD.n91 VDD.t189 5.13287
R416 VDD.n90 VDD.n69 5.13287
R417 VDD.n88 VDD.t51 5.13287
R418 VDD.n87 VDD.n71 5.13287
R419 VDD.n85 VDD.t114 5.13287
R420 VDD.n82 VDD.t207 5.13287
R421 VDD.n136 VDD.n68 5.13287
R422 VDD.n139 VDD.t158 5.13287
R423 VDD.n140 VDD.n67 5.13287
R424 VDD.n141 VDD.t245 5.13287
R425 VDD.n66 VDD.n65 5.13287
R426 VDD.n146 VDD.t220 5.13287
R427 VDD.n62 VDD.t140 5.13287
R428 VDD.n61 VDD.n41 5.13287
R429 VDD.n59 VDD.t128 5.13287
R430 VDD.n58 VDD.n43 5.13287
R431 VDD.n56 VDD.t238 5.13287
R432 VDD.n53 VDD.t156 5.13287
R433 VDD.n153 VDD.n40 5.13287
R434 VDD.n154 VDD.t148 5.13287
R435 VDD.n39 VDD.n38 5.13287
R436 VDD.n159 VDD.t126 5.13287
R437 VDD.n160 VDD.n37 5.13287
R438 VDD.n161 VDD.t205 5.13287
R439 VDD.n243 VDD.t88 5.13287
R440 VDD.n6 VDD.n5 5.13287
R441 VDD.n257 VDD.t43 5.09407
R442 VDD.n252 VDD.t167 5.09407
R443 VDD.n217 VDD.t53 5.09407
R444 VDD.n219 VDD.t152 5.09407
R445 VDD.n203 VDD.t49 5.09407
R446 VDD.n228 VDD.t10 5.09407
R447 VDD.n242 VDD.t33 5.09407
R448 VDD.n134 VDD.t27 5.09407
R449 VDD.n151 VDD.t31 5.09407
R450 VDD.n26 VDD.t1 5.09407
R451 VDD.n12 VDD.t171 5.09407
R452 VDD.n248 VDD.t154 5.09407
R453 VDD.n33 VDD.t197 4.9655
R454 VDD.n25 VDD.t0 4.26489
R455 VDD.n262 VDD.t90 4.12326
R456 VDD.n265 VDD.t165 4.12326
R457 VDD.n221 VDD.t67 4.11379
R458 VDD.n16 VDD.t195 4.09193
R459 VDD.n16 VDD.n8 4.0205
R460 VDD.n135 VDD.n90 3.90405
R461 VDD.n211 VDD.n210 3.1505
R462 VDD.n14 VDD.n11 3.0905
R463 VDD VDD.n2 3.04833
R464 VDD.n208 VDD.n207 2.85787
R465 VDD.n181 VDD.n171 2.85787
R466 VDD.n178 VDD.n174 2.85787
R467 VDD.n231 VDD.n195 2.85787
R468 VDD.n112 VDD.n103 2.85787
R469 VDD.n109 VDD.n106 2.85787
R470 VDD.n130 VDD.n93 2.85787
R471 VDD.n84 VDD.n74 2.85787
R472 VDD.n81 VDD.n77 2.85787
R473 VDD.n147 VDD.n64 2.85787
R474 VDD.n55 VDD.n46 2.85787
R475 VDD.n52 VDD.n49 2.85787
R476 VDD.n36 VDD.n35 2.85787
R477 VDD.n229 VDD 2.30404
R478 VDD.n207 VDD.t45 2.2755
R479 VDD.n207 VDD.n206 2.2755
R480 VDD.n171 VDD.t187 2.2755
R481 VDD.n171 VDD.n170 2.2755
R482 VDD.n174 VDD.t109 2.2755
R483 VDD.n174 VDD.n173 2.2755
R484 VDD.n195 VDD.t163 2.2755
R485 VDD.n195 VDD.n194 2.2755
R486 VDD.n103 VDD.t144 2.2755
R487 VDD.n103 VDD.n102 2.2755
R488 VDD.n106 VDD.t106 2.2755
R489 VDD.n106 VDD.n105 2.2755
R490 VDD.n93 VDD.t101 2.2755
R491 VDD.n93 VDD.n92 2.2755
R492 VDD.n74 VDD.t247 2.2755
R493 VDD.n74 VDD.n73 2.2755
R494 VDD.n77 VDD.t94 2.2755
R495 VDD.n77 VDD.n76 2.2755
R496 VDD.n64 VDD.t99 2.2755
R497 VDD.n64 VDD.n63 2.2755
R498 VDD.n46 VDD.t124 2.2755
R499 VDD.n46 VDD.n45 2.2755
R500 VDD.n49 VDD.t240 2.2755
R501 VDD.n49 VDD.n48 2.2755
R502 VDD.n35 VDD.t226 2.2755
R503 VDD.n35 VDD.n34 2.2755
R504 VDD.n2 VDD.t29 2.2755
R505 VDD.n2 VDD.n1 2.2755
R506 VDD.n17 VDD.n15 2.09907
R507 VDD.n20 VDD.n8 1.81414
R508 VDD.n10 VDD.n9 1.81414
R509 VDD.n14 VDD.n8 1.08595
R510 VDD.n241 VDD.n187 1.02928
R511 VDD.n152 VDD.n61 1.02928
R512 VDD VDD.n11 1.01181
R513 VDD.n119 VDD.n118 0.881662
R514 VDD.n212 VDD.t66 0.783764
R515 VDD.n15 VDD.n14 0.5405
R516 VDD.n247 VDD.n246 0.493148
R517 VDD VDD.n30 0.469361
R518 VDD.n20 VDD.n10 0.461409
R519 VDD.n29 VDD.n28 0.402136
R520 VDD.n262 VDD.n261 0.38985
R521 VDD.n27 VDD 0.268397
R522 VDD.n182 VDD.n181 0.233919
R523 VDD.n179 VDD.n178 0.233919
R524 VDD.n113 VDD.n112 0.233919
R525 VDD.n110 VDD.n109 0.233919
R526 VDD.n85 VDD.n84 0.233919
R527 VDD.n82 VDD.n81 0.233919
R528 VDD.n56 VDD.n55 0.233919
R529 VDD.n53 VDD.n52 0.233919
R530 VDD.n26 VDD.n6 0.228212
R531 VDD.n223 VDD.n222 0.224447
R532 VDD.n28 VDD.n27 0.204472
R533 VDD.n228 VDD.n227 0.204322
R534 VDD.n224 VDD.n223 0.202146
R535 VDD.n21 VDD.n20 0.19522
R536 VDD VDD.n226 0.179806
R537 VDD.n265 VDD.n264 0.173131
R538 VDD.n257 VDD.n256 0.170231
R539 VDD.n242 VDD.n241 0.167533
R540 VDD.n28 VDD.n6 0.165331
R541 VDD VDD.n62 0.160716
R542 VDD.n243 VDD 0.158984
R543 VDD VDD.n91 0.157289
R544 VDD.n152 VDD.n151 0.155496
R545 VDD.n135 VDD.n134 0.154581
R546 VDD.n185 VDD.n184 0.141016
R547 VDD.n116 VDD.n115 0.141016
R548 VDD.n88 VDD.n87 0.141016
R549 VDD.n59 VDD.n58 0.141016
R550 VDD.n223 VDD.n203 0.137126
R551 VDD.n12 VDD.n11 0.136815
R552 VDD.n264 VDD.n252 0.13637
R553 VDD.n248 VDD.n247 0.13637
R554 VDD.n136 VDD.n135 0.131861
R555 VDD.n238 VDD.n237 0.123551
R556 VDD.n235 VDD.n234 0.123551
R557 VDD.n140 VDD.n139 0.123551
R558 VDD.n141 VDD.n66 0.123551
R559 VDD.n154 VDD.n39 0.122176
R560 VDD.n160 VDD.n159 0.122176
R561 VDD.n123 VDD.n122 0.120831
R562 VDD.n124 VDD.n95 0.120831
R563 VDD.n241 VDD.n240 0.116432
R564 VDD.n153 VDD.n152 0.115137
R565 VDD.n260 VDD.n256 0.107339
R566 VDD.n226 VDD.n225 0.107339
R567 VDD.n187 VDD.n186 0.107339
R568 VDD.n184 VDD.n183 0.107339
R569 VDD.n118 VDD.n117 0.107339
R570 VDD.n115 VDD.n114 0.107339
R571 VDD.n90 VDD.n89 0.107339
R572 VDD.n87 VDD.n86 0.107339
R573 VDD.n61 VDD.n60 0.107339
R574 VDD.n58 VDD.n57 0.107339
R575 VDD.n232 VDD 0.10728
R576 VDD VDD.n146 0.10728
R577 VDD.n181 VDD 0.106177
R578 VDD.n178 VDD 0.106177
R579 VDD.n112 VDD 0.106177
R580 VDD.n109 VDD 0.106177
R581 VDD.n84 VDD 0.106177
R582 VDD.n81 VDD 0.106177
R583 VDD.n55 VDD 0.106177
R584 VDD.n52 VDD 0.106177
R585 VDD.n161 VDD 0.106087
R586 VDD VDD.n129 0.10492
R587 VDD VDD.n231 0.0981271
R588 VDD.n147 VDD 0.0981271
R589 VDD VDD.n36 0.0970363
R590 VDD.n130 VDD 0.0959696
R591 VDD.n240 VDD.n239 0.0940593
R592 VDD.n237 VDD.n236 0.0940593
R593 VDD.n234 VDD.n233 0.0940593
R594 VDD.n138 VDD.n136 0.0940593
R595 VDD.n142 VDD.n140 0.0940593
R596 VDD.n145 VDD.n66 0.0940593
R597 VDD.n231 VDD 0.0930424
R598 VDD VDD.n147 0.0930424
R599 VDD.n155 VDD.n153 0.093014
R600 VDD.n158 VDD.n39 0.093014
R601 VDD.n162 VDD.n160 0.093014
R602 VDD.n121 VDD.n119 0.0919917
R603 VDD.n125 VDD.n123 0.0919917
R604 VDD.n128 VDD.n95 0.0919917
R605 VDD VDD.n130 0.0909972
R606 VDD.n180 VDD.n179 0.080629
R607 VDD.n111 VDD.n110 0.080629
R608 VDD.n83 VDD.n82 0.080629
R609 VDD.n54 VDD.n53 0.080629
R610 VDD VDD.n185 0.0794677
R611 VDD VDD.n182 0.0794677
R612 VDD VDD.n116 0.0794677
R613 VDD VDD.n113 0.0794677
R614 VDD VDD.n88 0.0794677
R615 VDD VDD.n85 0.0794677
R616 VDD VDD.n59 0.0794677
R617 VDD VDD.n56 0.0794677
R618 VDD.n261 VDD 0.0759839
R619 VDD VDD.n26 0.0759545
R620 VDD.n29 VDD.n4 0.0727093
R621 VDD VDD.n257 0.0709717
R622 VDD VDD.n252 0.0709717
R623 VDD.n217 VDD 0.0709717
R624 VDD VDD.n203 0.0709717
R625 VDD VDD.n228 0.0709717
R626 VDD VDD.n248 0.0709717
R627 VDD.n230 VDD.n229 0.0706695
R628 VDD.n148 VDD.n62 0.0706695
R629 VDD.n244 VDD.n243 0.0698855
R630 VDD VDD.n238 0.0696525
R631 VDD VDD.n235 0.0696525
R632 VDD VDD.n232 0.0696525
R633 VDD.n139 VDD 0.0696525
R634 VDD VDD.n141 0.0696525
R635 VDD.n146 VDD 0.0696525
R636 VDD.n131 VDD.n91 0.0691188
R637 VDD VDD.n154 0.0688799
R638 VDD.n159 VDD 0.0688799
R639 VDD VDD.n161 0.0688799
R640 VDD.n122 VDD 0.0681243
R641 VDD VDD.n124 0.0681243
R642 VDD.n129 VDD 0.0681243
R643 VDD.n32 VDD.n0 0.064413
R644 VDD VDD.n0 0.0557174
R645 VDD VDD.n221 0.0555633
R646 VDD VDD.n224 0.0550806
R647 VDD.n264 VDD.n263 0.0545
R648 VDD VDD.n208 0.0533387
R649 VDD.n245 VDD.n36 0.0532933
R650 VDD.n151 VDD 0.0404465
R651 VDD VDD.n242 0.0400238
R652 VDD.n134 VDD 0.0396099
R653 VDD.n245 VDD 0.0392151
R654 VDD.n30 VDD.n29 0.0386026
R655 VDD VDD.n209 0.0382419
R656 VDD.n33 VDD 0.0363979
R657 VDD.n20 VDD 0.0362477
R658 VDD.n218 VDD.n208 0.0344677
R659 VDD.n251 VDD 0.0325968
R660 VDD VDD.n219 0.032019
R661 VDD VDD.n12 0.030261
R662 VDD.n246 VDD.n33 0.024997
R663 VDD VDD.n262 0.0240135
R664 VDD VDD.n265 0.0238871
R665 VDD.n247 VDD 0.0221129
R666 VDD.n28 VDD.n7 0.021736
R667 VDD VDD.n16 0.00978571
R668 VDD.n7 VDD 0.00858989
R669 VDD.n221 VDD 0.00543671
R670 VDD VDD.n260 0.00514516
R671 VDD.n225 VDD 0.00514516
R672 VDD.n222 VDD 0.00315823
R673 VDD.n210 VDD 0.00282258
R674 VDD.n4 VDD 0.00259302
R675 VDD.n27 VDD 0.00231818
R676 VDD.n186 VDD 0.00166129
R677 VDD.n183 VDD 0.00166129
R678 VDD VDD.n180 0.00166129
R679 VDD VDD.n177 0.00166129
R680 VDD.n117 VDD 0.00166129
R681 VDD.n114 VDD 0.00166129
R682 VDD VDD.n111 0.00166129
R683 VDD VDD.n108 0.00166129
R684 VDD.n89 VDD 0.00166129
R685 VDD.n86 VDD 0.00166129
R686 VDD VDD.n83 0.00166129
R687 VDD VDD.n80 0.00166129
R688 VDD.n60 VDD 0.00166129
R689 VDD.n57 VDD 0.00166129
R690 VDD VDD.n54 0.00166129
R691 VDD VDD.n51 0.00166129
R692 VDD.n263 VDD 0.00163514
R693 VDD VDD.n251 0.00162903
R694 VDD.n227 VDD 0.00159756
R695 VDD.n239 VDD 0.00151695
R696 VDD.n236 VDD 0.00151695
R697 VDD.n233 VDD 0.00151695
R698 VDD VDD.n230 0.00151695
R699 VDD VDD.n138 0.00151695
R700 VDD.n142 VDD 0.00151695
R701 VDD VDD.n145 0.00151695
R702 VDD.n148 VDD 0.00151695
R703 VDD.n155 VDD 0.00150559
R704 VDD VDD.n158 0.00150559
R705 VDD.n162 VDD 0.00150559
R706 VDD VDD.n244 0.00150559
R707 VDD VDD.n121 0.00149448
R708 VDD.n125 VDD 0.00149448
R709 VDD VDD.n128 0.00149448
R710 VDD.n131 VDD 0.00149448
R711 VDD.n21 VDD 0.00134112
R712 VDD.n17 VDD 0.00121429
R713 VDD.n210 VDD 0.00108064
R714 VDD VDD.n32 0.000934783
R715 VSS.n177 VSS.n176 19658.7
R716 VSS.t9 VSS.n37 17230
R717 VSS.n179 VSS.n177 16363.2
R718 VSS.n175 VSS.n35 14313.1
R719 VSS.n180 VSS.n179 12992.6
R720 VSS.n143 VSS.t23 10467.5
R721 VSS.n181 VSS.n22 8017.2
R722 VSS.n41 VSS.t140 7006.49
R723 VSS.n179 VSS.n178 6922.48
R724 VSS.t71 VSS.n48 6724.15
R725 VSS.n218 VSS.n184 6418.54
R726 VSS.n96 VSS.n95 4521.5
R727 VSS.n218 VSS.n183 4422.88
R728 VSS.n227 VSS.n10 3462.29
R729 VSS.n110 VSS.n109 3119.27
R730 VSS.n170 VSS.n169 2659.14
R731 VSS.n143 VSS.n142 2588.5
R732 VSS.t169 VSS.t167 2307.56
R733 VSS.t129 VSS.t83 2307.56
R734 VSS.t73 VSS.t114 2307.56
R735 VSS.t112 VSS.t164 2307.56
R736 VSS.t82 VSS.t161 2307.56
R737 VSS.t148 VSS.t37 2307.56
R738 VSS.t156 VSS.t42 2307.56
R739 VSS.t126 VSS.t101 2307.56
R740 VSS.t55 VSS.t76 2307.56
R741 VSS.n142 VSS.t138 2166.67
R742 VSS.n95 VSS.t98 2068.58
R743 VSS.t43 VSS.t58 1783.97
R744 VSS.t136 VSS.t4 1783.97
R745 VSS.t91 VSS.t89 1779.13
R746 VSS.t107 VSS.t110 1779.13
R747 VSS.t168 VSS.t132 1774.32
R748 VSS.t67 VSS.t154 1774.32
R749 VSS.t165 VSS.t33 1774.32
R750 VSS.t72 VSS.t143 1774.32
R751 VSS.t63 VSS.n79 1732.15
R752 VSS.n35 VSS.t115 1719.81
R753 VSS.n160 VSS.t2 1635.55
R754 VSS.t166 VSS.n54 1448.32
R755 VSS.n182 VSS.n181 1399.37
R756 VSS.n110 VSS.t62 1388.52
R757 VSS.n41 VSS.n40 1310.77
R758 VSS.n64 VSS.t14 1272.1
R759 VSS.n79 VSS.n78 1249.13
R760 VSS.t150 VSS.n10 1199.47
R761 VSS.n94 VSS.t96 1199.47
R762 VSS.n77 VSS.t38 1199.47
R763 VSS.n228 VSS.n227 1161.67
R764 VSS.n174 VSS.t92 1143.48
R765 VSS.n54 VSS.t50 1138.43
R766 VSS.n15 VSS.t105 1134.57
R767 VSS.n175 VSS.t48 1103.42
R768 VSS.t0 VSS.n110 1088.19
R769 VSS.t16 VSS.t46 1058.09
R770 VSS.n218 VSS.n182 1002.52
R771 VSS.n219 VSS.n218 988.177
R772 VSS.n154 VSS.t29 985.303
R773 VSS.n180 VSS.n175 947.745
R774 VSS.n198 VSS.n182 943.441
R775 VSS.n45 VSS.t121 927.716
R776 VSS.t114 VSS.t6 913.885
R777 VSS.t37 VSS.t12 913.885
R778 VSS.t76 VSS.t7 913.885
R779 VSS.n143 VSS.n42 766.241
R780 VSS.n93 VSS.t9 730.073
R781 VSS.t75 VSS.t100 706.523
R782 VSS.t11 VSS.t136 706.523
R783 VSS.t137 VSS.t86 704.607
R784 VSS.t22 VSS.t107 704.607
R785 VSS.t61 VSS.t131 702.703
R786 VSS.t8 VSS.t67 702.703
R787 VSS.t125 VSS.t163 702.703
R788 VSS.t13 VSS.t72 702.703
R789 VSS.t94 VSS.t119 696.831
R790 VSS.n9 VSS.t19 598.279
R791 VSS.n155 VSS.t64 578.554
R792 VSS.t115 VSS.n34 548.331
R793 VSS.t167 VSS.n33 548.331
R794 VSS.t83 VSS.n32 548.331
R795 VSS.t6 VSS.n31 548.331
R796 VSS.n80 VSS.t63 548.331
R797 VSS.n85 VSS.t164 548.331
R798 VSS.n86 VSS.t82 548.331
R799 VSS.n91 VSS.t12 548.331
R800 VSS.n65 VSS.t77 548.331
R801 VSS.n70 VSS.t42 548.331
R802 VSS.n71 VSS.t126 548.331
R803 VSS.n76 VSS.t7 548.331
R804 VSS.n156 VSS.n155 500.144
R805 VSS.n18 VSS.t28 490.991
R806 VSS.n144 VSS.n143 468.3
R807 VSS.n227 VSS.n226 429.526
R808 VSS.n78 VSS.n77 426.769
R809 VSS.n6 VSS.t44 426.396
R810 VSS.n194 VSS.t52 426.396
R811 VSS.n201 VSS.t68 426.396
R812 VSS.n49 VSS.t71 423.913
R813 VSS.n50 VSS.t43 423.913
R814 VSS.n51 VSS.t75 423.913
R815 VSS.n52 VSS.t11 423.913
R816 VSS.n60 VSS.t57 422.764
R817 VSS.n61 VSS.t91 422.764
R818 VSS.n62 VSS.t137 422.764
R819 VSS.n111 VSS.t22 422.764
R820 VSS.t62 VSS.n1 421.623
R821 VSS.n2 VSS.t168 421.623
R822 VSS.n3 VSS.t61 421.623
R823 VSS.n4 VSS.t8 421.623
R824 VSS.n55 VSS.t166 421.623
R825 VSS.n56 VSS.t165 421.623
R826 VSS.n57 VSS.t125 421.623
R827 VSS.n58 VSS.t13 421.623
R828 VSS.n34 VSS.t169 365.555
R829 VSS.n33 VSS.t129 365.555
R830 VSS.n32 VSS.t73 365.555
R831 VSS.n31 VSS.t150 365.555
R832 VSS.n80 VSS.t112 365.555
R833 VSS.t161 VSS.n85 365.555
R834 VSS.n86 VSS.t148 365.555
R835 VSS.t96 VSS.n91 365.555
R836 VSS.n65 VSS.t156 365.555
R837 VSS.t101 VSS.n70 365.555
R838 VSS.n71 VSS.t55 365.555
R839 VSS.t38 VSS.n76 365.555
R840 VSS.n96 VSS.n35 329.288
R841 VSS.t78 VSS.t146 329.029
R842 VSS.n157 VSS.n156 307.205
R843 VSS.n220 VSS.n219 288.551
R844 VSS.n42 VSS.n41 287.635
R845 VSS.t58 VSS.n49 282.61
R846 VSS.n50 VSS.t127 282.61
R847 VSS.t4 VSS.n51 282.61
R848 VSS.t50 VSS.n52 282.61
R849 VSS.t89 VSS.n60 281.844
R850 VSS.n61 VSS.t158 281.844
R851 VSS.t110 VSS.n62 281.844
R852 VSS.n111 VSS.t0 281.844
R853 VSS.t132 VSS.n1 281.082
R854 VSS.n2 VSS.t84 281.082
R855 VSS.t154 VSS.n3 281.082
R856 VSS.n4 VSS.t152 281.082
R857 VSS.t33 VSS.n55 281.082
R858 VSS.n56 VSS.t80 281.082
R859 VSS.t143 VSS.n57 281.082
R860 VSS.t98 VSS.n58 281.082
R861 VSS.t134 VSS.t26 220.721
R862 VSS.t40 VSS.t35 207.357
R863 VSS.n190 VSS.t78 191.375
R864 VSS.n109 VSS.n96 186.862
R865 VSS.n166 VSS.t79 186.381
R866 VSS.n165 VSS.t16 176.673
R867 VSS.n221 VSS.n220 162.162
R868 VSS.t79 VSS.n165 133.962
R869 VSS.n207 VSS.t134 128.379
R870 VSS.t46 VSS.n164 124.254
R871 VSS.n166 VSS.t65 124.254
R872 VSS.n12 VSS.t40 120.606
R873 VSS.t87 VSS.t17 112.944
R874 VSS.t64 VSS.n37 99.0148
R875 VSS.t44 VSS.t31 94.0088
R876 VSS.t52 VSS.t108 94.0088
R877 VSS.t68 VSS.t117 94.0088
R878 VSS.n164 VSS.n37 87.3661
R879 VSS.n218 VSS.n217 77.2216
R880 VSS.n170 VSS.t92 47.8266
R881 VSS.t48 VSS.n174 47.8266
R882 VSS.t119 VSS.n154 41.2109
R883 VSS.n103 VSS.t21 40.3374
R884 VSS.n77 VSS.n64 32.8288
R885 VSS.n148 VSS.t29 31.8449
R886 VSS.t21 VSS.t87 25.3551
R887 VSS.n181 VSS.n180 21.1044
R888 VSS.n94 VSS.n93 18.8411
R889 VSS.n10 VSS.n9 15.4399
R890 VSS.n109 VSS.n108 14.8335
R891 VSS.n146 VSS.n145 13.6116
R892 VSS.n157 VSS.t94 11.2397
R893 VSS.n96 VSS.n94 9.42079
R894 VSS.n173 VSS.t49 9.40866
R895 VSS.n104 VSS.t18 9.3736
R896 VSS.n8 VSS.t20 9.3736
R897 VSS.n63 VSS.t15 9.3736
R898 VSS.n92 VSS.t10 9.3736
R899 VSS.n148 VSS.n147 9.36649
R900 VSS.n203 VSS.t118 9.36362
R901 VSS.n212 VSS.t160 9.3221
R902 VSS.n205 VSS.n189 9.3221
R903 VSS.n200 VSS.t116 9.3221
R904 VSS.n197 VSS.n193 9.3221
R905 VSS.n14 VSS.t36 9.30652
R906 VSS.n17 VSS.t106 9.30652
R907 VSS.n192 VSS.t147 9.30652
R908 VSS.n196 VSS.t109 9.30652
R909 VSS.n162 VSS.t3 9.30652
R910 VSS.n152 VSS.t120 9.30652
R911 VSS.n47 VSS.t122 9.30652
R912 VSS.n208 VSS.t27 9.30607
R913 VSS.n159 VSS.t95 9.30518
R914 VSS.n151 VSS.t30 9.30518
R915 VSS.n140 VSS.t139 9.30323
R916 VSS.n231 VSS.t32 9.3025
R917 VSS.n11 VSS.t45 9.30189
R918 VSS.n230 VSS.n7 9.30189
R919 VSS.n172 VSS.t93 9.29981
R920 VSS.n210 VSS.n188 7.39136
R921 VSS.n213 VSS.t145 7.19156
R922 VSS.n238 VSS.t85 7.17323
R923 VSS.n240 VSS.t133 7.17323
R924 VSS.n125 VSS.t81 7.17323
R925 VSS.n127 VSS.t34 7.17323
R926 VSS.n36 VSS.t47 7.17156
R927 VSS.n116 VSS.t159 7.16989
R928 VSS.n118 VSS.t90 7.16989
R929 VSS.n134 VSS.t128 7.16656
R930 VSS.n136 VSS.t59 7.16656
R931 VSS.n224 VSS.t41 7.15156
R932 VSS.n88 VSS.t149 7.13489
R933 VSS.n83 VSS.t162 7.13489
R934 VSS.n82 VSS.t113 7.13489
R935 VSS.n28 VSS.t74 7.13323
R936 VSS.n26 VSS.t130 7.13323
R937 VSS.n24 VSS.t170 7.13323
R938 VSS.n102 VSS.t142 7.13156
R939 VSS.n100 VSS.t88 7.13156
R940 VSS.n98 VSS.t103 7.13156
R941 VSS.n73 VSS.t56 7.12823
R942 VSS.n68 VSS.t102 7.12823
R943 VSS.n67 VSS.t157 7.12823
R944 VSS.n223 VSS.t135 7.11732
R945 VSS.n224 VSS.n223 6.35063
R946 VSS VSS.t60 6.02876
R947 VSS.n44 VSS.n43 6.01414
R948 VSS.n44 VSS.t141 6.01414
R949 VSS.n168 VSS.t66 5.89898
R950 VSS.n121 VSS.t99 5.89565
R951 VSS.n123 VSS.t144 5.89565
R952 VSS.n234 VSS.t153 5.89565
R953 VSS.n236 VSS.t155 5.89565
R954 VSS.n112 VSS.t1 5.89232
R955 VSS.n114 VSS.t111 5.89232
R956 VSS.n130 VSS.t51 5.88898
R957 VSS.n132 VSS.t5 5.88898
R958 VSS.n89 VSS.t97 5.85732
R959 VSS.n29 VSS.t151 5.85565
R960 VSS.n106 VSS.t104 5.85398
R961 VSS.n74 VSS.t39 5.85065
R962 VSS VSS.n103 5.20137
R963 VSS.n108 VSS.n107 5.2005
R964 VSS.n108 VSS.n101 5.2005
R965 VSS.n108 VSS.n99 5.2005
R966 VSS.n108 VSS.n97 5.2005
R967 VSS.n237 VSS.n3 5.2005
R968 VSS.n235 VSS.n4 5.2005
R969 VSS.n229 VSS.n228 5.2005
R970 VSS.n232 VSS.n6 5.2005
R971 VSS.n226 VSS.n225 5.2005
R972 VSS.n13 VSS.n12 5.2005
R973 VSS.n19 VSS.n18 5.2005
R974 VSS.n222 VSS.n221 5.2005
R975 VSS.n209 VSS.n207 5.2005
R976 VSS.n199 VSS.n198 5.2005
R977 VSS.n195 VSS.n194 5.2005
R978 VSS.n186 VSS.n185 5.2005
R979 VSS.n191 VSS.n190 5.2005
R980 VSS.n202 VSS.n201 5.2005
R981 VSS.n16 VSS.n15 5.2005
R982 VSS.n9 VSS.n8 5.2005
R983 VSS.n31 VSS.n30 5.2005
R984 VSS.n32 VSS.n27 5.2005
R985 VSS.n33 VSS.n25 5.2005
R986 VSS.n34 VSS.n23 5.2005
R987 VSS.n64 VSS.n63 5.2005
R988 VSS.n91 VSS.n90 5.2005
R989 VSS.n87 VSS.n86 5.2005
R990 VSS.n85 VSS.n84 5.2005
R991 VSS.n81 VSS.n80 5.2005
R992 VSS.n93 VSS.n92 5.2005
R993 VSS.n171 VSS.n170 5.2005
R994 VSS.n174 VSS.n173 5.2005
R995 VSS.n164 VSS.n163 5.2005
R996 VSS.n167 VSS.n166 5.2005
R997 VSS.n161 VSS.n160 5.2005
R998 VSS.n142 VSS.n141 5.2005
R999 VSS.n150 VSS.n149 5.2005
R1000 VSS.n149 VSS.n148 5.2005
R1001 VSS.n154 VSS.n153 5.2005
R1002 VSS.n158 VSS.n157 5.2005
R1003 VSS.n46 VSS.n45 5.2005
R1004 VSS.n76 VSS.n75 5.2005
R1005 VSS.n72 VSS.n71 5.2005
R1006 VSS.n70 VSS.n69 5.2005
R1007 VSS.n66 VSS.n65 5.2005
R1008 VSS.n119 VSS.n60 5.2005
R1009 VSS.n117 VSS.n61 5.2005
R1010 VSS.n115 VSS.n62 5.2005
R1011 VSS.n113 VSS.n111 5.2005
R1012 VSS.n137 VSS.n49 5.2005
R1013 VSS.n135 VSS.n50 5.2005
R1014 VSS.n133 VSS.n51 5.2005
R1015 VSS.n131 VSS.n52 5.2005
R1016 VSS.n128 VSS.n55 5.2005
R1017 VSS.n126 VSS.n56 5.2005
R1018 VSS.n124 VSS.n57 5.2005
R1019 VSS.n122 VSS.n58 5.2005
R1020 VSS.n241 VSS.n1 5.2005
R1021 VSS.n239 VSS.n2 5.2005
R1022 VSS.n103 VSS.n96 4.61043
R1023 VSS.n211 VSS.n210 4.5005
R1024 VSS.n145 VSS.n39 4.5005
R1025 VSS.n145 VSS.n144 4.5005
R1026 VSS.n211 VSS 4.12355
R1027 VSS.n139 VSS.n44 3.28959
R1028 VSS.n216 VSS.n215 2.6005
R1029 VSS.n217 VSS.n216 2.6005
R1030 VSS.n140 VSS.n39 2.1373
R1031 VSS.n138 VSS 2.03738
R1032 VSS VSS.n200 1.00141
R1033 VSS.n233 VSS 0.930989
R1034 VSS.n225 VSS.n14 0.930556
R1035 VSS.n129 VSS.n53 0.844504
R1036 VSS.n120 VSS.n59 0.73994
R1037 VSS VSS.n159 0.676801
R1038 VSS.n233 VSS.n5 0.645242
R1039 VSS.n138 VSS.n47 0.616742
R1040 VSS.n105 VSS.n0 0.605616
R1041 VSS.n149 VSS.n146 0.486611
R1042 VSS.n167 VSS.n36 0.439554
R1043 VSS.n188 VSS.n187 0.349684
R1044 VSS.n20 VSS.n17 0.338437
R1045 VSS.n163 VSS.n162 0.316175
R1046 VSS VSS.n168 0.311851
R1047 VSS.n238 VSS.n237 0.286539
R1048 VSS.n222 VSS.n21 0.277931
R1049 VSS.n20 VSS.n19 0.272151
R1050 VSS.n234 VSS.n233 0.262771
R1051 VSS VSS.n82 0.261689
R1052 VSS.n83 VSS 0.261689
R1053 VSS VSS.n24 0.259875
R1054 VSS VSS.n26 0.259875
R1055 VSS VSS.n98 0.258086
R1056 VSS VSS.n100 0.258086
R1057 VSS VSS.n67 0.254582
R1058 VSS.n68 VSS 0.254582
R1059 VSS VSS.n172 0.223676
R1060 VSS.n90 VSS 0.22078
R1061 VSS.n30 VSS 0.21925
R1062 VSS.n107 VSS 0.217741
R1063 VSS.n75 VSS 0.214786
R1064 VSS.n129 VSS 0.206405
R1065 VSS VSS.n0 0.19412
R1066 VSS.n120 VSS 0.192251
R1067 VSS.n204 VSS.n192 0.188412
R1068 VSS.n197 VSS.n196 0.184546
R1069 VSS VSS.n151 0.182492
R1070 VSS.n139 VSS.n138 0.180913
R1071 VSS.n236 VSS.n235 0.156125
R1072 VSS.n134 VSS.n133 0.155663
R1073 VSS.n132 VSS.n131 0.155663
R1074 VSS.n125 VSS.n124 0.155663
R1075 VSS.n123 VSS.n122 0.155663
R1076 VSS.n116 VSS.n115 0.155663
R1077 VSS.n114 VSS.n113 0.155663
R1078 VSS VSS.n88 0.145885
R1079 VSS VSS.n28 0.144875
R1080 VSS VSS.n102 0.143879
R1081 VSS VSS.n73 0.141929
R1082 VSS.n199 VSS.n197 0.136634
R1083 VSS.n223 VSS 0.128863
R1084 VSS VSS.n5 0.127807
R1085 VSS VSS.n53 0.126709
R1086 VSS.n208 VSS.n21 0.12579
R1087 VSS.n200 VSS 0.115458
R1088 VSS.n136 VSS 0.111331
R1089 VSS.n127 VSS 0.111331
R1090 VSS.n118 VSS 0.111331
R1091 VSS.n152 VSS 0.109909
R1092 VSS.n172 VSS.n171 0.109351
R1093 VSS VSS.n59 0.106075
R1094 VSS VSS.n11 0.0924934
R1095 VSS.n82 VSS.n81 0.0905
R1096 VSS.n84 VSS.n83 0.0905
R1097 VSS.n88 VSS.n87 0.0905
R1098 VSS.n24 VSS.n23 0.089875
R1099 VSS.n26 VSS.n25 0.089875
R1100 VSS.n28 VSS.n27 0.089875
R1101 VSS.n153 VSS.n152 0.0895055
R1102 VSS.n98 VSS.n97 0.0892586
R1103 VSS.n100 VSS.n99 0.0892586
R1104 VSS.n102 VSS.n101 0.0892586
R1105 VSS.n67 VSS.n66 0.088051
R1106 VSS.n69 VSS.n68 0.088051
R1107 VSS.n73 VSS.n72 0.088051
R1108 VSS VSS.n224 0.0879825
R1109 VSS VSS.n89 0.0879825
R1110 VSS VSS.n29 0.087375
R1111 VSS.n151 VSS.n150 0.0869264
R1112 VSS VSS.n106 0.0867759
R1113 VSS VSS.n74 0.085602
R1114 VSS VSS.n36 0.085027
R1115 VSS.n168 VSS 0.085027
R1116 VSS.n89 VSS.n59 0.0779126
R1117 VSS.n21 VSS.n20 0.0777727
R1118 VSS.n29 VSS.n5 0.077375
R1119 VSS.n106 VSS.n105 0.0768448
R1120 VSS.n141 VSS.n139 0.0760505
R1121 VSS.n74 VSS.n53 0.0758061
R1122 VSS.n105 VSS.n104 0.0723269
R1123 VSS.n216 VSS.n188 0.071566
R1124 VSS.n206 VSS.n205 0.0706762
R1125 VSS.n39 VSS 0.0691188
R1126 VSS.n231 VSS.n230 0.0689718
R1127 VSS.n17 VSS.n16 0.0675755
R1128 VSS.n209 VSS.n208 0.0675755
R1129 VSS.n192 VSS.n191 0.0675755
R1130 VSS.n196 VSS.n195 0.0675755
R1131 VSS.n162 VSS.n161 0.0675755
R1132 VSS.n47 VSS.n46 0.0675755
R1133 VSS.n112 VSS.n0 0.0669985
R1134 VSS VSS.n236 0.0666607
R1135 VSS.n121 VSS.n120 0.0632596
R1136 VSS VSS.n140 0.0624266
R1137 VSS.n130 VSS.n129 0.0611231
R1138 VSS VSS.n213 0.0548172
R1139 VSS.n230 VSS.n229 0.0543206
R1140 VSS.n11 VSS 0.0459485
R1141 VSS.n205 VSS.n204 0.0449053
R1142 VSS.n159 VSS.n158 0.04
R1143 VSS.n137 VSS.n136 0.0386899
R1144 VSS.n135 VSS.n134 0.0386899
R1145 VSS.n128 VSS.n127 0.0386899
R1146 VSS.n126 VSS.n125 0.0386899
R1147 VSS.n119 VSS.n118 0.0386899
R1148 VSS.n117 VSS.n116 0.0386899
R1149 VSS.n241 VSS.n240 0.0386899
R1150 VSS.n239 VSS.n238 0.0386899
R1151 VSS VSS.n234 0.0377321
R1152 VSS VSS.n132 0.0376217
R1153 VSS VSS.n130 0.0376217
R1154 VSS VSS.n123 0.0376217
R1155 VSS VSS.n121 0.0376217
R1156 VSS VSS.n114 0.0376217
R1157 VSS VSS.n112 0.0376217
R1158 VSS.n216 VSS.n186 0.036033
R1159 VSS.n203 VSS.n202 0.0263217
R1160 VSS.n232 VSS.n231 0.0241213
R1161 VSS.n14 VSS.n13 0.0235097
R1162 VSS.n212 VSS.n211 0.0211167
R1163 VSS.n240 VSS 0.0154555
R1164 VSS.n204 VSS.n203 0.00960656
R1165 VSS.n213 VSS.n212 0.00644714
R1166 VSS.n81 VSS 0.00427622
R1167 VSS.n84 VSS 0.00427622
R1168 VSS.n87 VSS 0.00427622
R1169 VSS.n23 VSS 0.00425
R1170 VSS.n25 VSS 0.00425
R1171 VSS.n27 VSS 0.00425
R1172 VSS.n97 VSS 0.00422414
R1173 VSS.n99 VSS 0.00422414
R1174 VSS.n101 VSS 0.00422414
R1175 VSS.n66 VSS 0.00417347
R1176 VSS.n69 VSS 0.00417347
R1177 VSS.n72 VSS 0.00417347
R1178 VSS.n19 VSS 0.00380275
R1179 VSS VSS.n222 0.00380275
R1180 VSS VSS.n199 0.00352521
R1181 VSS.n237 VSS 0.0035
R1182 VSS.n225 VSS 0.00301748
R1183 VSS.n90 VSS 0.00301748
R1184 VSS.n30 VSS 0.003
R1185 VSS.n150 VSS.n38 0.00298619
R1186 VSS.n107 VSS 0.00298276
R1187 VSS.n75 VSS 0.00294898
R1188 VSS.n163 VSS 0.00293243
R1189 VSS VSS.n167 0.00293243
R1190 VSS.n8 VSS 0.00219811
R1191 VSS.n16 VSS 0.00219811
R1192 VSS VSS.n209 0.00219811
R1193 VSS.n191 VSS 0.00219811
R1194 VSS.n195 VSS 0.00219811
R1195 VSS.n63 VSS 0.00219811
R1196 VSS.n92 VSS 0.00219811
R1197 VSS.n161 VSS 0.00219811
R1198 VSS.n46 VSS 0.00219811
R1199 VSS.n141 VSS 0.00215138
R1200 VSS VSS.n137 0.00210237
R1201 VSS VSS.n135 0.00210237
R1202 VSS VSS.n128 0.00210237
R1203 VSS VSS.n126 0.00210237
R1204 VSS VSS.n119 0.00210237
R1205 VSS VSS.n117 0.00210237
R1206 VSS VSS.n241 0.00210237
R1207 VSS VSS.n239 0.00210237
R1208 VSS.n171 VSS 0.00171622
R1209 VSS.n173 VSS 0.00171622
R1210 VSS.n229 VSS 0.00169601
R1211 VSS.n235 VSS 0.00157143
R1212 VSS.n133 VSS 0.00156825
R1213 VSS.n131 VSS 0.00156825
R1214 VSS.n124 VSS 0.00156825
R1215 VSS.n122 VSS 0.00156825
R1216 VSS.n115 VSS 0.00156825
R1217 VSS.n113 VSS 0.00156825
R1218 VSS.n158 VSS 0.0015
R1219 VSS.n153 VSS 0.00149448
R1220 VSS VSS.n38 0.00149448
R1221 VSS.n104 VSS 0.00136539
R1222 VSS.n202 VSS 0.0013
R1223 VSS.n215 VSS.n214 0.00129295
R1224 VSS.n214 VSS 0.00129295
R1225 VSS VSS.n232 0.00109801
R1226 VSS.n13 VSS 0.00108252
R1227 VSS.n215 VSS.n206 0.000896476
R1228 JK_FF_mag_3.K.n0 JK_FF_mag_3.K.t2 30.9379
R1229 JK_FF_mag_3.K.n1 JK_FF_mag_3.K.t4 30.664
R1230 JK_FF_mag_3.K.n1 JK_FF_mag_3.K.t5 24.5385
R1231 JK_FF_mag_3.K.n0 JK_FF_mag_3.K.t3 24.5101
R1232 JK_FF_mag_3.K JK_FF_mag_3.K.n2 21.2236
R1233 JK_FF_mag_3.K JK_FF_mag_3.K.n3 5.29319
R1234 JK_FF_mag_3.K JK_FF_mag_3.K.n0 4.09208
R1235 JK_FF_mag_3.K.n2 JK_FF_mag_3.K 3.35432
R1236 JK_FF_mag_3.K.n2 JK_FF_mag_3.K 1.6274
R1237 JK_FF_mag_3.K JK_FF_mag_3.K.n1 1.4252
R1238 JK_FF_mag_1.K.n0 JK_FF_mag_1.K.t2 30.9379
R1239 JK_FF_mag_1.K.n1 JK_FF_mag_1.K.t4 30.664
R1240 JK_FF_mag_1.K.n1 JK_FF_mag_1.K.t5 24.5385
R1241 JK_FF_mag_1.K.n0 JK_FF_mag_1.K.t3 24.5101
R1242 JK_FF_mag_1.K JK_FF_mag_1.K.n2 7.46763
R1243 JK_FF_mag_1.K JK_FF_mag_1.K.n0 4.09208
R1244 JK_FF_mag_1.K.n2 JK_FF_mag_1.K 3.12156
R1245 JK_FF_mag_1.K.n2 JK_FF_mag_1.K 1.86016
R1246 JK_FF_mag_1.K JK_FF_mag_1.K.n1 1.4252
R1247 Q2.n0 Q2.t4 36.935
R1248 Q2.n7 Q2.t10 36.935
R1249 Q2.n2 Q2.t6 31.528
R1250 Q2.n0 Q2.t3 18.1962
R1251 Q2.n7 Q2.t9 18.1962
R1252 Q2.n12 Q2.n11 18.1259
R1253 Q2.n2 Q2.t5 15.3826
R1254 Q2.n13 Q2.n12 7.78566
R1255 Q2.n5 Q2.t7 7.483
R1256 Q2.n17 Q2.n14 7.09905
R1257 Q2.n3 Q2.n2 6.86029
R1258 Q2.n12 Q2 6.27254
R1259 Q2.n4 Q2.n1 5.01233
R1260 Q2.n5 Q2.t8 4.636
R1261 Q2.n10 Q2.n8 4.5005
R1262 Q2 Q2.n5 4.17425
R1263 Q2.n17 Q2.n16 3.24912
R1264 Q2.n18 Q2.n13 2.32428
R1265 Q2.n16 Q2.t1 2.2755
R1266 Q2.n16 Q2.n15 2.2755
R1267 Q2.n11 Q2.n6 2.251
R1268 Q2.n10 Q2.n9 2.24392
R1269 Q2.n1 Q2.n0 2.13398
R1270 Q2.n8 Q2.n7 2.12359
R1271 Q2.n13 Q2.n4 1.36395
R1272 Q2.n4 Q2.n3 1.12067
R1273 Q2.n18 Q2.n17 0.0919062
R1274 Q2.n3 Q2 0.0857632
R1275 Q2.n1 Q2 0.0810725
R1276 Q2 Q2.n18 0.073625
R1277 Q2.n9 Q2 0.0483237
R1278 Q2.n8 Q2.n6 0.0226053
R1279 Q2.n9 Q2.n6 0.0151658
R1280 Q2.n11 Q2.n10 0.0150625
R1281 Q1.n12 Q1.t10 36.935
R1282 Q1.n14 Q1.t8 31.528
R1283 Q1.n7 Q1.t11 31.528
R1284 Q1.n2 Q1.t15 30.9379
R1285 Q1.n1 Q1.t6 30.9379
R1286 Q1.n0 Q1.t13 30.9379
R1287 Q1.n23 Q1.t3 30.2877
R1288 Q1.n1 Q1.t12 24.5101
R1289 Q1.n23 Q1.t4 22.0463
R1290 Q1.n2 Q1.t16 21.6422
R1291 Q1.n0 Q1.t14 21.6422
R1292 Q1.n12 Q1.t9 18.1962
R1293 Q1.n26 Q1.n25 17.4222
R1294 Q1.n14 Q1.t7 15.3826
R1295 Q1.n7 Q1.t5 15.3826
R1296 Q1.n8 Q1.n7 7.62076
R1297 Q1.n20 Q1.n17 7.09905
R1298 Q1.n15 Q1.n14 6.86029
R1299 Q1.n25 Q1.n22 6.54023
R1300 Q1.n16 Q1.n13 5.01233
R1301 Q1.n11 Q1.n10 4.68036
R1302 Q1.n4 Q1.n3 4.64138
R1303 Q1.n25 Q1.n24 4.57443
R1304 Q1 Q1.n1 4.11094
R1305 Q1 Q1.n0 4.11094
R1306 Q1.n20 Q1.n19 3.24912
R1307 Q1.n3 Q1.n2 2.88363
R1308 Q1.n19 Q1.t2 2.2755
R1309 Q1.n19 Q1.n18 2.2755
R1310 Q1.n10 Q1.n9 2.251
R1311 Q1.n22 Q1.n21 2.2505
R1312 Q1.n6 Q1.n5 2.24218
R1313 Q1.n13 Q1.n12 2.13398
R1314 Q1.n24 Q1.n23 1.82835
R1315 Q1 Q1.n16 1.46982
R1316 Q1.n16 Q1.n15 1.12067
R1317 Q1.n26 Q1.n11 0.551624
R1318 Q1.n11 Q1.n4 0.525331
R1319 Q1.n4 Q1 0.299223
R1320 Q1 Q1.n26 0.285819
R1321 Q1.n24 Q1 0.10558
R1322 Q1.n21 Q1.n20 0.0919062
R1323 Q1.n15 Q1 0.0857632
R1324 Q1.n13 Q1 0.0810725
R1325 Q1.n21 Q1 0.073625
R1326 Q1.n3 Q1 0.0725473
R1327 Q1.n5 Q1 0.0496191
R1328 Q1.n9 Q1.n8 0.0226311
R1329 Q1.n10 Q1.n6 0.0148889
R1330 Q1.n22 Q1 0.0128158
R1331 Q0.n21 Q0.t7 40.1505
R1332 Q0.n7 Q0.t5 36.935
R1333 Q0.n16 Q0.t6 36.935
R1334 Q0.n0 Q0.t11 36.935
R1335 Q0.n9 Q0.t13 31.528
R1336 Q0.n13 Q0.t3 30.9379
R1337 Q0.n13 Q0.t9 21.6422
R1338 Q0.n23 Q0.n22 19.2517
R1339 Q0.n7 Q0.t12 18.1962
R1340 Q0.n16 Q0.t4 18.1962
R1341 Q0.n0 Q0.t10 18.1962
R1342 Q0.n21 Q0.t8 15.484
R1343 Q0.n9 Q0.t14 15.3826
R1344 Q0.n23 Q0 8.45416
R1345 Q0.n5 Q0.n2 7.09905
R1346 Q0.n10 Q0.n9 6.86029
R1347 Q0.n11 Q0.n8 5.01233
R1348 Q0.n15 Q0.n14 4.50508
R1349 Q0.n19 Q0.n18 4.5005
R1350 Q0.n20 Q0.n19 4.10652
R1351 Q0 Q0.n21 4.07224
R1352 Q0.n20 Q0.n13 4.06648
R1353 Q0.n25 Q0.n23 3.89052
R1354 Q0.n5 Q0.n4 3.24912
R1355 Q0.n12 Q0.n6 2.28145
R1356 Q0.n4 Q0.t1 2.2755
R1357 Q0.n4 Q0.n3 2.2755
R1358 Q0.n17 Q0.n16 2.14002
R1359 Q0.n8 Q0.n7 2.13398
R1360 Q0.n1 Q0.n0 2.12188
R1361 Q0.n22 Q0 1.75611
R1362 Q0.n12 Q0.n11 1.65779
R1363 Q0.n17 Q0.n14 1.5013
R1364 Q0.n26 Q0.n25 1.49857
R1365 Q0.n11 Q0.n10 1.12067
R1366 Q0.n22 Q0 0.487022
R1367 Q0.n6 Q0.n5 0.0919062
R1368 Q0.n10 Q0 0.0857632
R1369 Q0.n8 Q0 0.0810725
R1370 Q0.n6 Q0 0.073625
R1371 Q0 Q0.n12 0.0448919
R1372 Q0 Q0.n27 0.0442477
R1373 Q0.n27 Q0.n26 0.0361897
R1374 Q0.n19 Q0.n14 0.0309225
R1375 Q0.n15 Q0 0.0270574
R1376 Q0 Q0.n20 0.0200181
R1377 Q0.n18 Q0.n15 0.0182049
R1378 Q0.n25 Q0.n24 0.0102158
R1379 Q0.n18 Q0.n17 0.0082131
R1380 Q0.n26 Q0.n1 0.0067069
R1381 Q3.n0 Q3.t11 40.3485
R1382 Q3.n3 Q3.t9 36.935
R1383 Q3.n14 Q3.t5 31.528
R1384 Q3.n10 Q3.t10 31.528
R1385 Q3.n6 Q3.t6 31.528
R1386 Q3.n0 Q3.t12 30.0906
R1387 Q3.n3 Q3.t8 18.1962
R1388 Q3.n14 Q3.t4 15.3826
R1389 Q3.n10 Q3.t7 15.3826
R1390 Q3.n6 Q3.t3 15.3826
R1391 Q3.n8 Q3.n7 9.56316
R1392 Q3.n13 Q3.n12 9.38651
R1393 Q3.n23 Q3.n22 8.68206
R1394 Q3.n20 Q3.n17 7.09905
R1395 Q3.n15 Q3.n14 6.86029
R1396 Q3.n7 Q3.n6 6.15125
R1397 Q3.n11 Q3.n10 5.68213
R1398 Q3.n12 Q3.n5 4.5005
R1399 Q3.n12 Q3.n11 4.5005
R1400 Q3.n16 Q3.n13 3.42123
R1401 Q3.n20 Q3.n19 3.24912
R1402 Q3.n19 Q3.t1 2.2755
R1403 Q3.n19 Q3.n18 2.2755
R1404 Q3.n22 Q3.n21 2.2505
R1405 Q3.n24 Q3.n23 2.2441
R1406 Q3.n9 Q3.n8 2.24309
R1407 Q3.n4 Q3.n3 2.13398
R1408 Q3.n1 Q3.n0 2.1259
R1409 Q3.n13 Q3.n4 1.5916
R1410 Q3 Q3.n16 1.46621
R1411 Q3.n16 Q3.n15 1.12067
R1412 Q3.n21 Q3.n20 0.0919062
R1413 Q3.n15 Q3 0.0857632
R1414 Q3.n4 Q3 0.0810725
R1415 Q3.n21 Q3 0.073625
R1416 Q3.n5 Q3 0.0522241
R1417 Q3.n7 Q3 0.0515305
R1418 Q3.n9 Q3.n5 0.0361897
R1419 Q3.n25 Q3.n24 0.0251575
R1420 Q3 Q3.n25 0.0239247
R1421 Q3.n12 Q3.n8 0.0194736
R1422 Q3.n23 Q3.n2 0.0159575
R1423 Q3.n22 Q3 0.0141047
R1424 Q3.n11 Q3.n9 0.00515517
R1425 Q3.n24 Q3.n1 0.00470694
R1426 or_2_mag_3.IN1.n1 or_2_mag_3.IN1.t7 37.1981
R1427 or_2_mag_3.IN1.n2 or_2_mag_3.IN1.t5 31.528
R1428 or_2_mag_3.IN1.n0 or_2_mag_3.IN1.t8 30.5358
R1429 or_2_mag_3.IN1.n0 or_2_mag_3.IN1.t3 27.4841
R1430 or_2_mag_3.IN1.n1 or_2_mag_3.IN1.t6 17.6611
R1431 or_2_mag_3.IN1.n2 or_2_mag_3.IN1.t4 15.3826
R1432 or_2_mag_3.IN1 or_2_mag_3.IN1.n2 7.62758
R1433 or_2_mag_3.IN1.n3 or_2_mag_3.IN1 6.09789
R1434 or_2_mag_3.IN1 or_2_mag_3.IN1.n0 2.8878
R1435 or_2_mag_3.IN1.n3 or_2_mag_3.IN1 2.66613
R1436 or_2_mag_3.IN1.t1 or_2_mag_3.IN1.n3 2.2505
R1437 or_2_mag_3.IN1 or_2_mag_3.IN1.n1 1.43706
R1438 or_2_mag_3.IN1.t1 or_2_mag_3.IN1 0.4325
R1439 RST.n1 RST.t7 36.935
R1440 RST.n20 RST.t1 36.935
R1441 RST.n8 RST.t2 36.935
R1442 RST.n32 RST.t6 36.935
R1443 RST.n1 RST.t4 18.1962
R1444 RST.n20 RST.t0 18.1962
R1445 RST.n8 RST.t3 18.1962
R1446 RST.n32 RST.t5 18.1962
R1447 RST RST.n0 4.56717
R1448 RST RST.n0 4.5005
R1449 RST.n11 RST.n10 2.2505
R1450 RST.n22 RST.n17 2.24984
R1451 RST.n22 RST.n21 2.24984
R1452 RST.n24 RST.n23 2.24707
R1453 RST.n21 RST.n20 2.12601
R1454 RST.n2 RST.n1 2.12318
R1455 RST.n33 RST.n32 2.1224
R1456 RST.n9 RST.n8 2.12207
R1457 RST.n16 RST.n15 1.90023
R1458 RST.n28 RST.n27 1.87776
R1459 RST.n26 RST.n25 1.87165
R1460 RST.n35 RST.n34 1.5005
R1461 RST.n37 RST.n36 1.5005
R1462 RST.n14 RST.n13 1.5005
R1463 RST.n27 RST.n5 1.13106
R1464 RST.n40 RST.n0 1.12313
R1465 RST.n4 RST.n3 0.89746
R1466 RST.n40 RST.n39 0.63397
R1467 RST.n3 RST 0.0499589
R1468 RST.n31 RST 0.0363802
R1469 RST.n10 RST.n7 0.0361897
R1470 RST.n34 RST.n31 0.0346379
R1471 RST.n7 RST 0.031725
R1472 RST.n17 RST 0.0298963
R1473 RST.n3 RST.n2 0.0268355
R1474 RST.n22 RST.n18 0.0236959
R1475 RST.n15 RST.n14 0.0205676
R1476 RST.n37 RST.n28 0.0193514
R1477 RST.n36 RST.n29 0.0181289
R1478 RST.n25 RST.n24 0.0144865
R1479 RST.n23 RST.n22 0.0130264
R1480 RST.n10 RST.n9 0.0129138
R1481 RST.n27 RST.n26 0.0117737
R1482 RST.n11 RST.n6 0.0116103
R1483 RST.n21 RST.n19 0.011085
R1484 RST RST.n40 0.0100811
R1485 RST.n34 RST.n33 0.00825862
R1486 RST.n24 RST.n16 0.0077973
R1487 RST.n13 RST.n12 0.00513918
R1488 RST.n35 RST.n30 0.00513918
R1489 RST.n5 RST.n4 0.00504545
R1490 RST.n13 RST.n11 0.00328351
R1491 RST.n36 RST.n35 0.00328351
R1492 RST.n38 RST.n37 0.00232432
R1493 RST.n39 RST.n38 0.00232432
R1494 Vdiv11.n2 Vdiv11.n0 9.33985
R1495 Vdiv11.n2 Vdiv11.n1 5.17836
R1496 Vdiv11 Vdiv11.n2 0.115328
C0 a_939_3715# or_2_mag_0.IN1 0.0178f
C1 Q1 and2_mag_3.IN1 0.106f
C2 JK_FF_mag_3.nand2_mag_4.IN2 a_13607_4919# 0.069f
C3 a_12889_3822# JK_FF_mag_3.QB 3.33e-19
C4 JK_FF_mag_2.K JK_FF_mag_0.K 2.21e-19
C5 or_2_mag_0.GF_INV_MAG_1.IN VDD 0.411f
C6 and2_mag_0.GF_INV_MAG_0.IN CLK 1.93e-20
C7 a_2757_3818# a_2917_3818# 0.0504f
C8 a_9000_4915# VDD 2.21e-19
C9 nand3_mag_1.OUT and2_mag_3.OUT 0.109f
C10 Q0 and2_mag_1.GF_INV_MAG_0.IN 0.107f
C11 JK_FF_mag_3.nand3_mag_0.OUT VDD 0.647f
C12 a_4199_4915# or_2_mag_3.IN2 0.00964f
C13 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C14 JK_FF_mag_2.nand3_mag_2.OUT JK_FF_mag_2.K 0.105f
C15 JK_FF_mag_3.nand2_mag_3.IN1 a_12325_3822# 0.00119f
C16 JK_FF_mag_2.nand3_mag_1.IN1 a_9730_3818# 0.0697f
C17 JK_FF_mag_2.nand2_mag_4.IN2 CLK 0.01f
C18 JK_FF_mag_2.nand3_mag_0.OUT Q0 3.4e-19
C19 JK_FF_mag_0.nand3_mag_1.IN1 or_2_mag_3.IN1 6.57e-19
C20 a_939_3715# and2_mag_0.GF_INV_MAG_0.IN 1.14e-19
C21 or_2_mag_0.GF_INV_MAG_1.IN or_2_mag_0.IN1 0.226f
C22 or_2_mag_0.GF_INV_MAG_1.IN Q3 1.51e-19
C23 or_2_mag_0.IN1 VDD 0.378f
C24 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_3.K 0.00544f
C25 Q3 VDD 4.24f
C26 Q0 a_14017_3822# 0.069f
C27 a_3635_4915# JK_FF_mag_0.nand3_mag_1.IN1 8.64e-19
C28 a_13607_4919# JK_FF_mag_3.QB 0.00964f
C29 JK_FF_mag_0.nand3_mag_0.OUT a_2917_3818# 0.0732f
C30 JK_FF_mag_2.K Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 4.04e-19
C31 JK_FF_mag_2.nand3_mag_2.OUT JK_FF_mag_2.nand3_mag_1.IN1 0.00158f
C32 JK_FF_mag_0.nand2_mag_1.IN2 CLK 0.00637f
C33 or_2_mag_3.IN2 JK_FF_mag_0.K 2.8e-19
C34 JK_FF_mag_3.K JK_FF_mag_2.nand3_mag_0.OUT 1.83e-19
C35 or_2_mag_0.GF_INV_MAG_1.IN and2_mag_0.GF_INV_MAG_0.IN 9.6e-19
C36 or_2_mag_0.IN1 Q3 0.00935f
C37 and2_mag_0.GF_INV_MAG_0.IN VDD 0.433f
C38 Q1 JK_FF_mag_2.nand2_mag_3.IN1 0.0309f
C39 JK_FF_mag_3.nand3_mag_2.OUT JK_FF_mag_3.nand3_mag_1.IN1 0.00156f
C40 JK_FF_mag_3.QB JK_FF_mag_3.nand3_mag_1.IN1 0.0404f
C41 a_7639_1615# CLK 0.00487f
C42 JK_FF_mag_0.nand3_mag_0.OUT a_2757_3818# 0.0203f
C43 JK_FF_mag_2.nand2_mag_4.IN2 VDD 0.391f
C44 Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN Vdiv11 1.71e-21
C45 Q1 or_2_mag_1.IN1 0.203f
C46 and2_mag_0.GF_INV_MAG_0.IN or_2_mag_0.IN1 0.126f
C47 or_2_mag_3.IN1 GF_INV_MAG_1.OUT 1.2e-19
C48 or_2_mag_0.IN2 CLK 6.61e-20
C49 and2_mag_0.GF_INV_MAG_0.IN Q3 0.329f
C50 Q1 a_n20_2787# 0.00369f
C51 JK_FF_mag_3.nand2_mag_3.IN1 CLK 0.416f
C52 JK_FF_mag_1.nand2_mag_3.IN1 a_7334_4917# 0.0036f
C53 JK_FF_mag_1.nand2_mag_1.IN2 or_2_mag_3.IN1 6.18e-19
C54 JK_FF_mag_0.nand2_mag_1.IN2 VDD 0.397f
C55 JK_FF_mag_1.nand2_mag_4.IN2 Q0 1.65e-21
C56 a_939_3715# or_2_mag_0.IN2 0.0177f
C57 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_2.K 2.01e-19
C58 a_12319_4919# JK_FF_mag_3.nand2_mag_3.IN1 1.46e-19
C59 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_1.K 2.39e-21
C60 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.nand2_mag_1.IN2 0.36f
C61 Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN a_11241_1205# 2.31e-19
C62 a_2751_4915# JK_FF_mag_0.K 8.64e-19
C63 Q1 and2_mag_2.GF_INV_MAG_0.IN 0.146f
C64 JK_FF_mag_1.QB or_2_mag_3.IN1 0.00209f
C65 or_2_mag_3.IN1 and2_mag_3.GF_INV_MAG_0.IN 5.73e-20
C66 Q2 and2_mag_3.IN1 0.00392f
C67 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_1.K 3.98e-19
C68 or_2_mag_3.IN2 a_2849_1480# 8.64e-19
C69 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.QB 0.28f
C70 Q1 RST 0.16f
C71 JK_FF_mag_0.nand2_mag_1.IN2 Q3 0.11f
C72 a_7744_3820# Q2 0.069f
C73 Q1 a_10448_4915# 0.00859f
C74 JK_FF_mag_1.K or_2_mag_3.IN1 2.19f
C75 or_2_mag_0.GF_INV_MAG_1.IN or_2_mag_0.IN2 0.0512f
C76 or_2_mag_3.GF_INV_MAG_1.IN CLK 5.45e-20
C77 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_2.OUT 0.121f
C78 Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN and2_mag_3.IN1 2.29e-19
C79 or_2_mag_0.IN2 VDD 0.657f
C80 Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN a_11081_1205# 3.59e-19
C81 JK_FF_mag_3.K a_12165_3822# 0.00472f
C82 CLK and2_mag_3.OUT 0.00104f
C83 Q0 a_13607_4919# 0.00859f
C84 JK_FF_mag_1.K JK_FF_mag_1.nand2_mag_3.IN1 0.0702f
C85 JK_FF_mag_1.K nand3_mag_0.OUT 7.98e-20
C86 JK_FF_mag_3.nand2_mag_3.IN1 VDD 1.16f
C87 RST JK_FF_mag_2.nand2_mag_3.IN1 0.0695f
C88 and2_mag_2.GF_INV_MAG_0.IN or_2_mag_1.IN1 0.124f
C89 JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_3.nand3_mag_0.OUT 0.0894f
C90 a_140_2787# Q3 6.63e-20
C91 or_2_mag_3.IN2 a_1377_1477# 2.69e-22
C92 JK_FF_mag_0.nand3_mag_1.IN1 or_2_mag_3.IN2 0.0379f
C93 JK_FF_mag_2.nand2_mag_3.IN1 a_10448_4915# 0.0036f
C94 Q0 Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00776f
C95 a_7479_1615# VDD 5.08e-19
C96 Q1 a_n27_2146# 0.00544f
C97 or_2_mag_0.IN1 or_2_mag_0.IN2 0.209f
C98 Q1 Q2 2.34f
C99 nor_3_mag_0.IN3 VDD 0.514f
C100 or_2_mag_0.IN2 Q3 8e-19
C101 Q0 JK_FF_mag_3.nand3_mag_1.IN1 0.00425f
C102 RST JK_FF_mag_1.nand3_mag_2.OUT 0.0903f
C103 a_3635_4915# JK_FF_mag_0.nand3_mag_2.OUT 2.88e-20
C104 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C105 JK_FF_mag_2.K JK_FF_mag_1.nand2_mag_1.IN2 0.0052f
C106 JK_FF_mag_3.K Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 9.58e-19
C107 JK_FF_mag_0.nand2_mag_3.IN1 CLK 0.519f
C108 Q1 Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 3.09e-19
C109 Q0 a_2849_1480# 0.00589f
C110 and2_mag_1.GF_INV_MAG_0.IN CLK 0.00323f
C111 nor_3_mag_0.IN3 Q3 0.0224f
C112 and2_mag_0.GF_INV_MAG_0.IN or_2_mag_0.IN2 0.0108f
C113 or_2_mag_3.GF_INV_MAG_1.IN VDD 0.409f
C114 Q1 a_1385_2540# 0.0205f
C115 JK_FF_mag_3.K JK_FF_mag_3.nand3_mag_1.IN1 2.51e-19
C116 Q1 or_2_mag_1.GF_INV_MAG_1.IN 0.0364f
C117 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.QB 0.0377f
C118 JK_FF_mag_2.K JK_FF_mag_1.QB 0.00917f
C119 JK_FF_mag_0.nand3_mag_0.OUT a_3481_3818# 0.00378f
C120 JK_FF_mag_2.K and2_mag_3.GF_INV_MAG_0.IN 0.00118f
C121 and2_mag_3.OUT VDD 0.303f
C122 JK_FF_mag_2.nand3_mag_0.OUT CLK 0.276f
C123 nand3_mag_1.OUT Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 2.25e-19
C124 a_3475_4915# JK_FF_mag_0.nand3_mag_2.OUT 9.1e-19
C125 JK_FF_mag_0.nand3_mag_0.OUT Q2 8.93e-19
C126 or_2_mag_1.IN1 Q2 0.026f
C127 Q2 JK_FF_mag_1.nand3_mag_2.OUT 0.338f
C128 a_5892_3820# a_6052_3820# 0.0504f
C129 JK_FF_mag_1.K JK_FF_mag_1.nand3_mag_1.IN1 2.56e-19
C130 JK_FF_mag_1.K JK_FF_mag_2.K 1.57f
C131 Q0 a_1377_1477# 0.00718f
C132 or_2_mag_3.GF_INV_MAG_1.IN Q3 1.34e-19
C133 RST a_10448_4915# 0.00107f
C134 a_9166_3818# or_2_mag_3.IN1 0.00392f
C135 a_12165_3822# a_12325_3822# 0.0504f
C136 Q3 and2_mag_3.OUT 0.161f
C137 JK_FF_mag_2.K a_8344_1618# 2.5e-19
C138 and2_mag_2.GF_INV_MAG_0.IN a_n27_2146# 0.069f
C139 or_2_mag_1.IN1 or_2_mag_1.GF_INV_MAG_1.IN 0.205f
C140 or_2_mag_1.IN1 a_1385_2540# 1.78e-20
C141 and2_mag_2.GF_INV_MAG_0.IN Q2 9.25e-19
C142 Q2 a_6052_3820# 2.79e-20
C143 a_11241_1205# or_2_mag_3.IN1 1.9e-19
C144 or_2_mag_0.GF_INV_MAG_1.IN and2_mag_1.GF_INV_MAG_0.IN 1.84e-19
C145 JK_FF_mag_1.nand2_mag_4.IN2 JK_FF_mag_1.nand3_mag_1.OUT 0.122f
C146 JK_FF_mag_0.nand2_mag_3.IN1 VDD 1.15f
C147 JK_FF_mag_3.K JK_FF_mag_0.nand3_mag_1.IN1 8.28e-20
C148 JK_FF_mag_1.QB or_2_mag_3.IN2 2.25e-21
C149 and2_mag_1.GF_INV_MAG_0.IN VDD 0.423f
C150 RST Q2 0.163f
C151 JK_FF_mag_2.nand3_mag_0.OUT VDD 0.647f
C152 and2_mag_2.GF_INV_MAG_0.IN or_2_mag_1.GF_INV_MAG_1.IN 4.7e-20
C153 JK_FF_mag_1.K or_2_mag_3.IN2 0.412f
C154 or_2_mag_3.IN1 and2_mag_3.IN1 2.11e-19
C155 JK_FF_mag_0.nand2_mag_3.IN1 Q3 0.0281f
C156 Q1 JK_FF_mag_2.nand3_mag_1.OUT 0.0346f
C157 a_14017_3822# VDD 3.56e-19
C158 a_12889_3822# CLK 6.43e-21
C159 Q0 GF_INV_MAG_1.OUT 1.61e-19
C160 a_7479_1615# a_7639_1615# 0.0504f
C161 JK_FF_mag_0.nand3_mag_2.OUT or_2_mag_3.IN2 0.103f
C162 a_9730_3818# CLK 3.8e-19
C163 JK_FF_mag_1.nand2_mag_4.IN2 CLK 0.00995f
C164 JK_FF_mag_0.K CLK 0.779f
C165 JK_FF_mag_1.nand3_mag_1.OUT Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 2.98e-19
C166 JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_2.nand2_mag_3.IN1 0.16f
C167 Q0 JK_FF_mag_1.nand2_mag_1.IN2 6.35e-19
C168 a_7744_3820# JK_FF_mag_1.nand2_mag_3.IN1 0.00118f
C169 JK_FF_mag_1.K a_4763_4915# 1.44e-21
C170 a_12165_3822# CLK 0.0101f
C171 Q1 a_9884_4915# 0.0101f
C172 JK_FF_mag_1.QB JK_FF_mag_1.nand3_mag_0.OUT 0.342f
C173 a_9166_3818# JK_FF_mag_2.K 8.21e-19
C174 JK_FF_mag_3.K GF_INV_MAG_1.OUT 1.89e-19
C175 a_13453_3822# VDD 3.14e-19
C176 JK_FF_mag_1.QB Q0 0.00121f
C177 JK_FF_mag_2.nand3_mag_2.OUT CLK 0.26f
C178 Q0 and2_mag_3.GF_INV_MAG_0.IN 8.33e-20
C179 a_4199_4915# VDD 3.14e-19
C180 or_2_mag_1.GF_INV_MAG_1.IN Q2 0.0766f
C181 Q1 or_2_mag_3.IN1 2.57f
C182 a_2911_4915# JK_FF_mag_0.nand3_mag_2.OUT 0.0731f
C183 Q1 JK_FF_mag_2.nand2_mag_1.IN2 0.11f
C184 JK_FF_mag_3.K JK_FF_mag_1.nand2_mag_1.IN2 8.26e-20
C185 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand2_mag_1.IN2 0.00975f
C186 JK_FF_mag_1.K JK_FF_mag_1.nand3_mag_0.OUT 0.0951f
C187 nand3_mag_1.OUT GF_INV_MAG_1.OUT 0.131f
C188 a_7180_3820# JK_FF_mag_1.nand2_mag_3.IN1 0.011f
C189 JK_FF_mag_1.nand2_mag_3.IN1 Q1 0.00917f
C190 Q1 nand3_mag_0.OUT 0.117f
C191 JK_FF_mag_1.K Q0 0.0709f
C192 Q1 a_9724_4915# 0.0102f
C193 JK_FF_mag_3.K JK_FF_mag_1.QB 3.18e-19
C194 JK_FF_mag_2.nand3_mag_2.OUT a_9160_4915# 0.0731f
C195 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_0.nand2_mag_3.IN1 0.36f
C196 CLK Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 6.86e-20
C197 or_2_mag_3.IN1 JK_FF_mag_2.nand2_mag_3.IN1 0.306f
C198 a_9006_3818# JK_FF_mag_2.K 0.00598f
C199 a_12889_3822# VDD 3.14e-19
C200 JK_FF_mag_3.K and2_mag_3.GF_INV_MAG_0.IN 4.11e-19
C201 JK_FF_mag_2.nand2_mag_1.IN2 JK_FF_mag_2.nand2_mag_3.IN1 0.36f
C202 a_12889_3822# JK_FF_mag_3.nand3_mag_0.OUT 0.00378f
C203 a_4199_4915# Q3 0.00859f
C204 a_9730_3818# VDD 3.14e-19
C205 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.nand3_mag_1.OUT 0.0622f
C206 JK_FF_mag_1.nand2_mag_4.IN2 VDD 0.391f
C207 or_2_mag_0.GF_INV_MAG_1.IN JK_FF_mag_0.K 0.129f
C208 JK_FF_mag_1.QB a_6610_4917# 0.00695f
C209 Q1 a_11012_4915# 0.0157f
C210 JK_FF_mag_3.nand3_mag_1.IN1 CLK 9.85e-20
C211 a_2751_4915# JK_FF_mag_0.nand3_mag_2.OUT 0.0202f
C212 JK_FF_mag_0.K VDD 0.592f
C213 JK_FF_mag_2.K and2_mag_3.IN1 0.00441f
C214 JK_FF_mag_1.QB nand3_mag_1.OUT 9.75e-21
C215 JK_FF_mag_0.nand3_mag_0.OUT or_2_mag_3.IN1 6.36e-19
C216 a_12165_3822# VDD 2.21e-19
C217 JK_FF_mag_3.K JK_FF_mag_1.K 0.00238f
C218 nor_3_mag_0.IN3 and2_mag_3.OUT 0.191f
C219 a_12165_3822# JK_FF_mag_3.nand3_mag_0.OUT 0.0203f
C220 nand3_mag_1.OUT and2_mag_3.GF_INV_MAG_0.IN 0.048f
C221 JK_FF_mag_2.nand3_mag_1.OUT RST 0.284f
C222 Q1 a_10858_3818# 0.069f
C223 JK_FF_mag_2.nand3_mag_1.OUT a_10448_4915# 0.00378f
C224 JK_FF_mag_2.nand3_mag_2.OUT a_9000_4915# 0.0202f
C225 JK_FF_mag_2.nand3_mag_2.OUT VDD 0.642f
C226 a_7744_3820# JK_FF_mag_2.K 8.11e-19
C227 CLK a_2849_1480# 1.64e-20
C228 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.nand3_mag_2.OUT 0.00118f
C229 or_2_mag_0.IN1 JK_FF_mag_0.K 0.00265f
C230 or_2_mag_1.IN1 nand3_mag_0.OUT 1.74e-19
C231 Q3 JK_FF_mag_0.K 0.133f
C232 JK_FF_mag_0.nand2_mag_4.IN2 RST 0.0306f
C233 and2_mag_1.GF_INV_MAG_0.IN or_2_mag_0.IN2 0.00574f
C234 a_n20_2787# nand3_mag_0.OUT 0.0202f
C235 a_10858_3818# JK_FF_mag_2.nand2_mag_3.IN1 0.00118f
C236 a_13607_4919# VDD 3.14e-19
C237 JK_FF_mag_3.nand2_mag_4.IN2 JK_FF_mag_3.nand2_mag_1.IN2 8.16e-20
C238 JK_FF_mag_3.nand3_mag_1.OUT RST 0.265f
C239 JK_FF_mag_1.QB a_6616_3820# 3.12e-19
C240 nand3_mag_1.OUT a_8344_1618# 2.05e-19
C241 a_9884_4915# RST 0.00193f
C242 JK_FF_mag_0.nand3_mag_1.OUT RST 0.278f
C243 Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VDD 0.52f
C244 Q1 JK_FF_mag_1.nand3_mag_1.IN1 1.17e-19
C245 JK_FF_mag_2.K Q1 1.93f
C246 JK_FF_mag_0.nand3_mag_1.IN1 CLK 0.0844f
C247 a_7180_3820# JK_FF_mag_1.nand3_mag_1.IN1 0.0059f
C248 a_7180_3820# JK_FF_mag_2.K 3.47e-19
C249 JK_FF_mag_1.nand2_mag_3.IN1 a_6052_3820# 0.00119f
C250 and2_mag_0.GF_INV_MAG_0.IN JK_FF_mag_0.K 1.5e-20
C251 and2_mag_2.GF_INV_MAG_0.IN nand3_mag_0.OUT 1.01e-19
C252 RST or_2_mag_3.IN1 0.376f
C253 JK_FF_mag_2.nand2_mag_1.IN2 RST 1.36e-19
C254 JK_FF_mag_3.nand3_mag_1.IN1 VDD 0.66f
C255 JK_FF_mag_3.nand3_mag_1.IN1 JK_FF_mag_3.nand3_mag_0.OUT 0.122f
C256 Q1 JK_FF_mag_3.QB 1.76e-21
C257 or_2_mag_3.IN1 a_10448_4915# 0.00964f
C258 Q1 JK_FF_mag_3.nand3_mag_2.OUT 3.39e-20
C259 a_2917_3818# or_2_mag_3.IN2 0.00392f
C260 a_10294_3818# JK_FF_mag_2.nand2_mag_3.IN1 0.011f
C261 a_13043_4919# RST 0.00162f
C262 JK_FF_mag_1.nand2_mag_3.IN1 RST 0.0703f
C263 a_7334_4917# JK_FF_mag_1.nand3_mag_1.OUT 0.00378f
C264 a_14017_3822# JK_FF_mag_3.nand2_mag_3.IN1 0.00118f
C265 a_9724_4915# RST 0.00176f
C266 JK_FF_mag_2.K JK_FF_mag_2.nand2_mag_3.IN1 0.0707f
C267 Q3 Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.013f
C268 JK_FF_mag_0.nand2_mag_4.IN2 a_4609_3818# 4.52e-20
C269 a_3635_4915# RST 0.00327f
C270 a_3481_3818# JK_FF_mag_0.nand3_mag_1.OUT 0.0195f
C271 JK_FF_mag_0.nand3_mag_1.OUT Q2 1.05e-19
C272 a_2849_1480# VDD 0.165f
C273 JK_FF_mag_2.nand3_mag_1.IN1 Q1 0.00403f
C274 JK_FF_mag_0.nand2_mag_3.IN1 or_2_mag_3.GF_INV_MAG_1.IN 7.97e-19
C275 JK_FF_mag_1.nand2_mag_1.IN2 JK_FF_mag_1.nand3_mag_1.OUT 0.00975f
C276 nor_3_mag_0.OUT Vdiv11 0.119f
C277 JK_FF_mag_3.QB JK_FF_mag_3.nand2_mag_1.IN2 0.0592f
C278 RST a_11012_4915# 0.00106f
C279 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_2.K 2.01e-19
C280 Q2 or_2_mag_3.IN1 0.109f
C281 JK_FF_mag_2.K or_2_mag_1.IN1 2.75e-19
C282 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand3_mag_2.OUT 0.00156f
C283 JK_FF_mag_1.QB JK_FF_mag_1.nand3_mag_1.OUT 0.25f
C284 Q1 or_2_mag_3.IN2 0.0161f
C285 RST JK_FF_mag_3.nand2_mag_4.IN2 0.00146f
C286 a_12883_4919# RST 0.00176f
C287 JK_FF_mag_2.nand3_mag_1.IN1 JK_FF_mag_2.nand2_mag_3.IN1 0.233f
C288 a_13453_3822# JK_FF_mag_3.nand2_mag_3.IN1 0.011f
C289 JK_FF_mag_1.nand2_mag_3.IN1 Q2 0.0274f
C290 Q2 nand3_mag_0.OUT 0.306f
C291 JK_FF_mag_2.nand3_mag_0.OUT and2_mag_3.OUT 1.39e-19
C292 a_3475_4915# RST 0.00183f
C293 JK_FF_mag_1.nand3_mag_2.OUT a_6046_4917# 0.0731f
C294 a_1377_1477# VDD 0.165f
C295 JK_FF_mag_0.nand3_mag_1.IN1 VDD 0.651f
C296 nor_3_mag_0.OUT a_11241_1205# 0.198f
C297 Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN or_2_mag_3.IN1 1.2e-19
C298 Q0 and2_mag_3.IN1 0.104f
C299 JK_FF_mag_1.K JK_FF_mag_1.nand3_mag_1.OUT 2.51e-19
C300 or_2_mag_1.GF_INV_MAG_1.IN or_2_mag_3.IN1 9.22e-20
C301 JK_FF_mag_0.nand3_mag_1.OUT a_4045_3818# 4.52e-20
C302 JK_FF_mag_2.K and2_mag_2.GF_INV_MAG_0.IN 1.64e-20
C303 JK_FF_mag_1.nand2_mag_1.IN2 CLK 0.00639f
C304 JK_FF_mag_1.QB a_6770_4917# 0.00696f
C305 a_12889_3822# JK_FF_mag_3.nand2_mag_3.IN1 1.43e-19
C306 or_2_mag_0.IN2 JK_FF_mag_0.K 0.00121f
C307 JK_FF_mag_0.nand3_mag_1.IN1 Q3 0.00397f
C308 JK_FF_mag_0.nand3_mag_0.OUT or_2_mag_3.IN2 0.342f
C309 JK_FF_mag_1.nand3_mag_2.OUT or_2_mag_3.IN2 7.36e-21
C310 a_7898_4917# VDD 3.14e-19
C311 or_2_mag_1.IN1 or_2_mag_3.IN2 9.21e-19
C312 JK_FF_mag_1.nand3_mag_1.IN1 RST 0.186f
C313 JK_FF_mag_2.K RST 0.0781f
C314 JK_FF_mag_3.K and2_mag_3.IN1 0.00243f
C315 JK_FF_mag_1.QB CLK 0.484f
C316 nor_3_mag_0.OUT a_11081_1205# 0.0135f
C317 and2_mag_3.GF_INV_MAG_0.IN CLK 5.73e-19
C318 JK_FF_mag_3.nand3_mag_2.OUT RST 0.0957f
C319 RST JK_FF_mag_3.QB 0.141f
C320 RST a_6046_4917# 0.00201f
C321 Q1 JK_FF_mag_1.nand3_mag_0.OUT 1.17e-19
C322 and2_mag_3.IN1 nand3_mag_1.OUT 0.407f
C323 a_11081_1205# nand3_mag_1.OUT 8.09e-22
C324 JK_FF_mag_1.K CLK 0.631f
C325 Q1 Q0 3.23f
C326 JK_FF_mag_2.nand3_mag_1.IN1 RST 0.185f
C327 a_7639_1615# Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 8.5e-20
C328 a_7334_4917# VDD 3.14e-19
C329 GF_INV_MAG_1.OUT VDD 0.569f
C330 a_6052_3820# or_2_mag_3.IN2 1.24e-20
C331 JK_FF_mag_1.K a_5886_4917# 8.64e-19
C332 JK_FF_mag_1.nand3_mag_1.IN1 Q2 0.00391f
C333 JK_FF_mag_2.K Q2 0.291f
C334 JK_FF_mag_3.nand2_mag_3.IN1 a_13607_4919# 0.0036f
C335 JK_FF_mag_0.nand3_mag_2.OUT CLK 0.271f
C336 JK_FF_mag_1.nand2_mag_1.IN2 VDD 0.397f
C337 a_9884_4915# JK_FF_mag_2.nand3_mag_1.OUT 0.0733f
C338 Q0 JK_FF_mag_2.nand2_mag_3.IN1 0.0143f
C339 RST or_2_mag_3.IN2 0.299f
C340 Q2 a_6046_4917# 0.00789f
C341 JK_FF_mag_3.K Q1 3.7f
C342 Q0 JK_FF_mag_3.nand2_mag_1.IN2 0.11f
C343 nor_3_mag_0.OUT Q1 3.11e-19
C344 JK_FF_mag_0.nand2_mag_3.IN1 a_4199_4915# 0.0036f
C345 JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_3.nand3_mag_1.IN1 0.24f
C346 JK_FF_mag_2.nand3_mag_1.OUT or_2_mag_3.IN1 0.25f
C347 Q3 GF_INV_MAG_1.OUT 0.0238f
C348 a_7479_1615# Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 1.32e-19
C349 JK_FF_mag_2.nand2_mag_1.IN2 JK_FF_mag_2.nand3_mag_1.OUT 0.00975f
C350 JK_FF_mag_1.QB VDD 0.904f
C351 JK_FF_mag_1.nand3_mag_2.OUT JK_FF_mag_1.nand3_mag_0.OUT 0.00183f
C352 and2_mag_3.GF_INV_MAG_0.IN VDD 0.423f
C353 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand2_mag_4.IN2 0.122f
C354 a_5892_3820# or_2_mag_3.IN2 1.59e-20
C355 or_2_mag_1.IN1 Q0 0.205f
C356 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_0.nand3_mag_1.IN1 0.109f
C357 JK_FF_mag_2.K or_2_mag_1.GF_INV_MAG_1.IN 0.133f
C358 Q1 nand3_mag_1.OUT 0.0409f
C359 JK_FF_mag_3.K JK_FF_mag_2.nand2_mag_3.IN1 0.0129f
C360 JK_FF_mag_0.nand2_mag_4.IN2 or_2_mag_3.IN1 3.61e-21
C361 Q0 a_n20_2787# 0.00765f
C362 RST a_4763_4915# 0.00131f
C363 a_9724_4915# JK_FF_mag_2.nand3_mag_1.OUT 0.0203f
C364 a_3481_3818# or_2_mag_3.IN2 3.33e-19
C365 a_2911_4915# RST 6.39e-19
C366 JK_FF_mag_1.K VDD 0.881f
C367 Q2 or_2_mag_3.IN2 0.0661f
C368 Q1 a_12159_4919# 5.5e-19
C369 JK_FF_mag_1.QB Q3 9.05e-22
C370 a_n20_4333# VDD 3.14e-19
C371 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_3.K 8.64e-20
C372 a_9884_4915# or_2_mag_3.IN1 0.00696f
C373 JK_FF_mag_0.nand3_mag_1.OUT or_2_mag_3.IN1 7.17e-19
C374 a_8344_1618# VDD 3.14e-19
C375 a_6052_3820# JK_FF_mag_1.nand3_mag_0.OUT 0.0732f
C376 a_4609_3818# or_2_mag_3.IN2 0.0114f
C377 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.K 0.0502f
C378 and2_mag_2.GF_INV_MAG_0.IN Q0 0.00525f
C379 a_13043_4919# JK_FF_mag_3.nand3_mag_1.OUT 0.0733f
C380 JK_FF_mag_1.nand3_mag_2.OUT a_6610_4917# 9.1e-19
C381 JK_FF_mag_0.nand3_mag_2.OUT VDD 0.642f
C382 and2_mag_1.GF_INV_MAG_0.IN JK_FF_mag_0.K 4.68e-20
C383 JK_FF_mag_2.nand2_mag_1.IN2 or_2_mag_3.IN1 0.0598f
C384 JK_FF_mag_2.nand3_mag_0.OUT a_9730_3818# 0.00378f
C385 a_9724_4915# a_9884_4915# 0.0504f
C386 RST JK_FF_mag_1.nand3_mag_0.OUT 5.45e-20
C387 JK_FF_mag_1.K Q3 0.0703f
C388 a_3635_4915# JK_FF_mag_0.nand3_mag_1.OUT 0.0733f
C389 a_2751_4915# RST 5.07e-19
C390 or_2_mag_1.GF_INV_MAG_1.IN or_2_mag_3.IN2 0.00397f
C391 Q0 RST 0.0664f
C392 a_9166_3818# CLK 0.0105f
C393 Q3 a_n20_4333# 0.0111f
C394 JK_FF_mag_1.nand2_mag_3.IN1 or_2_mag_3.IN1 0.0231f
C395 a_9724_4915# or_2_mag_3.IN1 0.00695f
C396 a_5892_3820# JK_FF_mag_1.nand3_mag_0.OUT 0.0203f
C397 a_4045_3818# or_2_mag_3.IN2 2.96e-19
C398 Q3 JK_FF_mag_0.nand3_mag_2.OUT 0.349f
C399 or_2_mag_3.GF_INV_MAG_1.IN a_2849_1480# 0.132f
C400 a_12883_4919# JK_FF_mag_3.nand3_mag_1.OUT 0.0203f
C401 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand2_mag_4.IN2 0.122f
C402 a_11012_4915# or_2_mag_3.IN1 0.0811f
C403 JK_FF_mag_2.nand3_mag_2.OUT JK_FF_mag_2.nand3_mag_0.OUT 0.00183f
C404 JK_FF_mag_2.nand3_mag_1.OUT a_10294_3818# 4.52e-20
C405 JK_FF_mag_3.K RST 0.0864f
C406 and2_mag_0.GF_INV_MAG_0.IN a_n20_4333# 0.069f
C407 a_3475_4915# JK_FF_mag_0.nand3_mag_1.OUT 0.0203f
C408 JK_FF_mag_2.K JK_FF_mag_2.nand3_mag_1.OUT 0.00188f
C409 Q2 JK_FF_mag_1.nand3_mag_0.OUT 9.75e-19
C410 a_9006_3818# CLK 0.0114f
C411 JK_FF_mag_3.K a_10448_4915# 5.58e-22
C412 Q0 Q2 0.888f
C413 RST a_6610_4917# 0.00176f
C414 a_10858_3818# or_2_mag_3.IN1 0.0114f
C415 JK_FF_mag_2.nand2_mag_1.IN2 a_10858_3818# 0.00372f
C416 Vdiv11 VDD 0.153f
C417 and2_mag_3.IN1 CLK 0.0765f
C418 a_7180_3820# JK_FF_mag_1.nand3_mag_1.OUT 4.52e-20
C419 a_12883_4919# a_13043_4919# 0.0504f
C420 Q1 JK_FF_mag_1.nand3_mag_1.OUT 1.36e-19
C421 JK_FF_mag_1.nand2_mag_1.IN2 a_7639_1615# 4.33e-21
C422 JK_FF_mag_2.nand3_mag_1.IN1 JK_FF_mag_2.nand3_mag_1.OUT 0.768f
C423 RST a_12159_4919# 0.00201f
C424 a_2917_3818# CLK 0.0105f
C425 a_3475_4915# a_3635_4915# 0.0504f
C426 Q0 Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 1.61e-19
C427 a_7744_3820# CLK 9.33e-19
C428 JK_FF_mag_3.K Q2 4.54f
C429 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_2.K 2.33e-19
C430 Q0 a_1385_2540# 0.00379f
C431 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_1.K 3.43e-19
C432 or_2_mag_1.GF_INV_MAG_1.IN Q0 0.0582f
C433 a_10294_3818# or_2_mag_3.IN1 2.96e-19
C434 JK_FF_mag_3.nand3_mag_2.OUT JK_FF_mag_3.nand3_mag_1.OUT 0.121f
C435 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.QB 0.249f
C436 Q2 a_6610_4917# 0.0102f
C437 Vdiv11 Q3 0.00291f
C438 JK_FF_mag_2.nand2_mag_1.IN2 a_10294_3818# 0.069f
C439 a_11241_1205# VDD 0.0418f
C440 a_7639_1615# and2_mag_3.GF_INV_MAG_0.IN 4.43e-21
C441 JK_FF_mag_1.nand3_mag_1.IN1 or_2_mag_3.IN1 6.51e-19
C442 JK_FF_mag_2.K or_2_mag_3.IN1 0.161f
C443 nor_3_mag_0.IN3 GF_INV_MAG_1.OUT 1.5e-20
C444 RST a_6616_3820# 3.08e-20
C445 JK_FF_mag_3.nand3_mag_2.OUT or_2_mag_3.IN1 1.47e-20
C446 JK_FF_mag_3.K Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 1.89e-19
C447 nor_3_mag_0.OUT Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 0.00307f
C448 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.nand3_mag_1.IN1 0.233f
C449 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_2.K 0.0106f
C450 JK_FF_mag_2.nand3_mag_1.IN1 a_9884_4915# 8.64e-19
C451 JK_FF_mag_1.nand3_mag_2.OUT JK_FF_mag_1.nand3_mag_1.OUT 0.121f
C452 a_9006_3818# VDD 2.21e-19
C453 a_2757_3818# CLK 0.0114f
C454 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand3_mag_1.IN1 0.233f
C455 JK_FF_mag_3.K or_2_mag_1.GF_INV_MAG_1.IN 1.84e-21
C456 a_7180_3820# CLK 9.25e-19
C457 Q1 CLK 0.554f
C458 JK_FF_mag_0.nand2_mag_4.IN2 or_2_mag_3.IN2 0.198f
C459 JK_FF_mag_3.nand3_mag_2.OUT a_13043_4919# 2.88e-20
C460 a_13043_4919# JK_FF_mag_3.QB 0.00696f
C461 a_11241_1205# Q3 0.0504f
C462 JK_FF_mag_2.nand3_mag_1.IN1 or_2_mag_3.IN1 0.0385f
C463 JK_FF_mag_1.nand2_mag_3.IN1 a_6046_4917# 1.46e-19
C464 and2_mag_3.IN1 VDD 0.795f
C465 a_7479_1615# and2_mag_3.GF_INV_MAG_0.IN 3.44e-21
C466 JK_FF_mag_2.nand3_mag_1.IN1 JK_FF_mag_2.nand2_mag_1.IN2 0.109f
C467 a_11081_1205# VDD 0.235f
C468 Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN nand3_mag_1.OUT 9.5e-19
C469 a_13453_3822# JK_FF_mag_3.nand3_mag_1.IN1 0.00605f
C470 Q1 a_12319_4919# 4.28e-19
C471 RST a_12325_3822# 7.84e-19
C472 JK_FF_mag_0.nand3_mag_1.OUT or_2_mag_3.IN2 0.25f
C473 or_2_mag_0.GF_INV_MAG_1.IN a_2917_3818# 1.03e-20
C474 or_2_mag_0.IN2 a_n20_4333# 3.93e-20
C475 GF_INV_MAG_1.OUT and2_mag_3.OUT 0.00982f
C476 JK_FF_mag_2.nand2_mag_3.IN1 CLK 0.527f
C477 Q1 a_9160_4915# 0.00789f
C478 a_7744_3820# VDD 3.56e-19
C479 JK_FF_mag_3.nand2_mag_1.IN2 CLK 1.48e-20
C480 JK_FF_mag_1.nand3_mag_2.OUT a_6770_4917# 2.88e-20
C481 or_2_mag_3.IN1 or_2_mag_3.IN2 0.211f
C482 JK_FF_mag_0.nand2_mag_4.IN2 a_4763_4915# 0.00372f
C483 JK_FF_mag_3.nand3_mag_2.OUT a_12883_4919# 9.1e-19
C484 a_12883_4919# JK_FF_mag_3.QB 0.00695f
C485 Q3 and2_mag_3.IN1 0.119f
C486 a_11081_1205# Q3 0.0186f
C487 JK_FF_mag_3.nand2_mag_4.IN2 JK_FF_mag_3.QB 0.198f
C488 JK_FF_mag_0.nand3_mag_0.OUT CLK 0.275f
C489 JK_FF_mag_1.nand3_mag_2.OUT CLK 0.26f
C490 JK_FF_mag_1.nand2_mag_3.IN1 or_2_mag_3.IN2 5.42e-20
C491 a_12889_3822# JK_FF_mag_3.nand3_mag_1.IN1 0.0697f
C492 RST JK_FF_mag_1.nand3_mag_1.OUT 0.284f
C493 a_9160_4915# JK_FF_mag_2.nand2_mag_3.IN1 1.46e-19
C494 or_2_mag_0.GF_INV_MAG_1.IN a_2757_3818# 1.29e-20
C495 a_3635_4915# or_2_mag_3.IN2 0.00696f
C496 JK_FF_mag_1.nand3_mag_2.OUT a_5886_4917# 0.0202f
C497 and2_mag_3.GF_INV_MAG_0.IN and2_mag_3.OUT 0.129f
C498 Q1 or_2_mag_0.GF_INV_MAG_1.IN 8.19e-19
C499 JK_FF_mag_0.nand3_mag_1.OUT a_2911_4915# 1.5e-20
C500 a_2917_3818# Q3 3.43e-19
C501 Q0 JK_FF_mag_2.nand3_mag_1.OUT 3.94e-19
C502 a_2757_3818# VDD 2.21e-19
C503 Q1 a_9000_4915# 0.00335f
C504 Q1 VDD 3.43f
C505 a_7180_3820# VDD 3.14e-19
C506 or_2_mag_3.GF_INV_MAG_1.IN JK_FF_mag_1.K 2.04e-19
C507 JK_FF_mag_2.K JK_FF_mag_1.nand3_mag_1.IN1 0.00254f
C508 JK_FF_mag_3.nand2_mag_4.IN2 a_14171_4919# 0.00372f
C509 a_6052_3820# CLK 0.0105f
C510 RST a_6770_4917# 0.00192f
C511 Q0 JK_FF_mag_3.nand3_mag_1.OUT 0.0349f
C512 JK_FF_mag_3.K JK_FF_mag_2.nand3_mag_1.OUT 2.12e-19
C513 Q2 JK_FF_mag_1.nand3_mag_1.OUT 0.0345f
C514 JK_FF_mag_2.nand2_mag_3.IN1 VDD 1.17f
C515 a_3475_4915# or_2_mag_3.IN2 0.00695f
C516 Q1 or_2_mag_0.IN1 3.8e-20
C517 a_8344_1618# and2_mag_3.OUT 6.43e-19
C518 a_2757_3818# Q3 4.47e-19
C519 JK_FF_mag_0.nand3_mag_1.OUT a_2751_4915# 1.17e-20
C520 JK_FF_mag_3.nand2_mag_1.IN2 VDD 0.397f
C521 JK_FF_mag_2.nand3_mag_1.IN1 a_10294_3818# 0.0059f
C522 Q1 Q3 1.83f
C523 JK_FF_mag_3.nand3_mag_2.OUT JK_FF_mag_3.QB 0.103f
C524 RST CLK 3.44f
C525 JK_FF_mag_1.nand3_mag_0.OUT or_2_mag_3.IN1 6.18e-19
C526 JK_FF_mag_2.nand3_mag_1.IN1 JK_FF_mag_2.K 0.00154f
C527 Q0 or_2_mag_3.IN1 4.75f
C528 JK_FF_mag_0.nand3_mag_0.OUT VDD 0.647f
C529 JK_FF_mag_2.nand2_mag_1.IN2 Q0 3.4e-19
C530 JK_FF_mag_1.nand3_mag_2.OUT VDD 0.642f
C531 or_2_mag_1.IN1 VDD 0.338f
C532 RST a_5886_4917# 0.00201f
C533 a_12319_4919# RST 0.00201f
C534 JK_FF_mag_3.K JK_FF_mag_3.nand3_mag_1.OUT 2.47e-19
C535 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.nand3_mag_0.OUT 0.0894f
C536 a_5892_3820# CLK 0.0114f
C537 Q0 a_13043_4919# 0.0101f
C538 JK_FF_mag_1.QB JK_FF_mag_2.nand3_mag_0.OUT 2.46e-20
C539 a_n20_2787# VDD 2.21e-19
C540 JK_FF_mag_1.nand2_mag_3.IN1 Q0 0.0187f
C541 Q2 a_6770_4917# 0.0101f
C542 Q0 nand3_mag_0.OUT 0.305f
C543 Q1 and2_mag_0.GF_INV_MAG_0.IN 0.116f
C544 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_1.K 0.0135f
C545 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_3.K 5.2e-20
C546 a_9160_4915# RST 0.00202f
C547 JK_FF_mag_1.K and2_mag_1.GF_INV_MAG_0.IN 0.121f
C548 JK_FF_mag_2.K or_2_mag_3.IN2 1.93f
C549 a_14171_4919# JK_FF_mag_3.QB 0.0811f
C550 a_3481_3818# CLK 3.8e-19
C551 nor_3_mag_0.OUT or_2_mag_3.IN1 1.2e-19
C552 JK_FF_mag_3.K or_2_mag_3.IN1 0.507f
C553 JK_FF_mag_3.K JK_FF_mag_2.nand2_mag_1.IN2 1.83e-19
C554 JK_FF_mag_0.nand3_mag_0.OUT Q3 0.00107f
C555 Q2 CLK 1.48f
C556 JK_FF_mag_1.nand3_mag_2.OUT Q3 3.26e-20
C557 or_2_mag_1.IN1 Q3 0.0145f
C558 Q1 JK_FF_mag_2.nand2_mag_4.IN2 0.0635f
C559 and2_mag_2.GF_INV_MAG_0.IN VDD 0.423f
C560 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand3_mag_2.OUT 0.00118f
C561 JK_FF_mag_1.nand2_mag_4.IN2 a_7898_4917# 0.00372f
C562 and2_mag_3.IN1 a_7639_1615# 0.00107f
C563 Q2 a_5886_4917# 0.00335f
C564 JK_FF_mag_3.K JK_FF_mag_1.nand2_mag_3.IN1 0.00301f
C565 a_4609_3818# CLK 9.34e-19
C566 a_n20_2787# Q3 4.15e-19
C567 nor_3_mag_0.IN3 a_11241_1205# 2.84e-20
C568 JK_FF_mag_3.nand3_mag_1.OUT a_12159_4919# 1.17e-20
C569 Q0 JK_FF_mag_3.nand2_mag_4.IN2 0.0635f
C570 Q0 a_12883_4919# 0.0102f
C571 or_2_mag_3.IN1 nand3_mag_1.OUT 4.78e-20
C572 a_939_3715# Q2 0.00208f
C573 a_9000_4915# RST 0.00202f
C574 RST VDD 0.972f
C575 RST JK_FF_mag_3.nand3_mag_0.OUT 0.00543f
C576 a_9160_4915# Q2 4.66e-19
C577 JK_FF_mag_2.nand2_mag_3.IN1 JK_FF_mag_2.nand2_mag_4.IN2 0.321f
C578 a_10448_4915# VDD 3.14e-19
C579 JK_FF_mag_3.K a_11012_4915# 2.75e-21
C580 or_2_mag_1.GF_INV_MAG_1.IN CLK 1.48e-19
C581 JK_FF_mag_0.nand2_mag_1.IN2 Q1 1.32e-19
C582 and2_mag_2.GF_INV_MAG_0.IN Q3 0.299f
C583 JK_FF_mag_1.nand2_mag_4.IN2 a_7334_4917# 0.069f
C584 a_5892_3820# VDD 2.21e-19
C585 and2_mag_3.IN1 a_7479_1615# 0.00271f
C586 a_4045_3818# CLK 9.23e-19
C587 nor_3_mag_0.IN3 a_11081_1205# 9.09e-19
C588 a_11241_1205# and2_mag_3.OUT 8.64e-19
C589 RST Q3 0.144f
C590 or_2_mag_0.GF_INV_MAG_1.IN Q2 0.0131f
C591 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand3_mag_0.OUT 0.122f
C592 JK_FF_mag_2.K JK_FF_mag_1.nand3_mag_0.OUT 2e-19
C593 JK_FF_mag_1.nand2_mag_4.IN2 JK_FF_mag_1.nand2_mag_1.IN2 8.16e-20
C594 Q1 a_140_2787# 1.75e-19
C595 a_3481_3818# VDD 3.14e-19
C596 a_9000_4915# Q2 6.02e-19
C597 a_n27_2146# VDD 3.14e-19
C598 Q1 a_7639_1615# 5.19e-20
C599 JK_FF_mag_1.nand3_mag_1.IN1 Q0 3.53e-19
C600 JK_FF_mag_2.K Q0 1.76f
C601 a_4199_4915# JK_FF_mag_1.K 4.96e-22
C602 Q2 VDD 2.58f
C603 JK_FF_mag_1.nand2_mag_3.IN1 a_6616_3820# 1.43e-19
C604 Q0 JK_FF_mag_3.nand3_mag_2.OUT 0.338f
C605 Q0 JK_FF_mag_3.QB 1.99f
C606 JK_FF_mag_1.nand2_mag_4.IN2 JK_FF_mag_1.QB 0.198f
C607 Q1 or_2_mag_0.IN2 0.00103f
C608 a_4763_4915# or_2_mag_3.IN2 0.0811f
C609 a_4609_3818# VDD 3.56e-19
C610 or_2_mag_0.IN1 Q2 0.0814f
C611 or_2_mag_3.IN1 a_12325_3822# 1.19e-20
C612 and2_mag_3.IN1 and2_mag_3.OUT 0.012f
C613 a_11081_1205# and2_mag_3.OUT 0.0105f
C614 or_2_mag_0.GF_INV_MAG_1.IN a_1385_2540# 3.01e-20
C615 Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN VDD 0.512f
C616 JK_FF_mag_3.K JK_FF_mag_1.nand3_mag_1.IN1 8.26e-20
C617 JK_FF_mag_3.K JK_FF_mag_2.K 0.195f
C618 a_n27_2146# Q3 0.00572f
C619 JK_FF_mag_2.nand3_mag_1.IN1 Q0 3.56e-19
C620 Q2 Q3 1.19f
C621 Q1 a_7479_1615# 3.35e-20
C622 a_1385_2540# VDD 3.14e-19
C623 or_2_mag_1.GF_INV_MAG_1.IN VDD 0.408f
C624 RST JK_FF_mag_2.nand2_mag_4.IN2 0.0287f
C625 JK_FF_mag_3.K JK_FF_mag_3.nand3_mag_2.OUT 0.105f
C626 JK_FF_mag_3.K JK_FF_mag_3.QB 6.93e-19
C627 nor_3_mag_0.IN3 Q1 4.07e-19
C628 a_9166_3818# JK_FF_mag_2.nand3_mag_0.OUT 0.0732f
C629 a_4609_3818# Q3 0.069f
C630 JK_FF_mag_1.K JK_FF_mag_0.K 3.43e-19
C631 Q0 a_14171_4919# 0.0157f
C632 JK_FF_mag_2.nand2_mag_4.IN2 a_10448_4915# 0.069f
C633 JK_FF_mag_1.nand3_mag_0.OUT or_2_mag_3.IN2 2.62e-20
C634 a_4045_3818# VDD 3.14e-19
C635 JK_FF_mag_2.K nand3_mag_1.OUT 1.32e-19
C636 a_n20_2787# a_140_2787# 0.0504f
C637 JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_3.nand2_mag_1.IN2 0.36f
C638 Q0 or_2_mag_3.IN2 0.0485f
C639 JK_FF_mag_2.nand3_mag_1.IN1 JK_FF_mag_3.K 1.83e-19
C640 JK_FF_mag_2.nand3_mag_1.OUT CLK 0.0833f
C641 Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN Q3 0.029f
C642 or_2_mag_3.IN1 JK_FF_mag_1.nand3_mag_1.OUT 7.11e-19
C643 and2_mag_0.GF_INV_MAG_0.IN Q2 0.0609f
C644 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.K 0.105f
C645 or_2_mag_1.GF_INV_MAG_1.IN Q3 1.4e-20
C646 JK_FF_mag_0.nand2_mag_1.IN2 RST 1.36e-19
C647 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.nand3_mag_1.OUT 0.16f
C648 or_2_mag_3.GF_INV_MAG_1.IN Q1 0.0248f
C649 and2_mag_3.GF_INV_MAG_0.IN Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 1.05e-20
C650 JK_FF_mag_0.nand2_mag_4.IN2 CLK 0.01f
C651 a_9006_3818# JK_FF_mag_2.nand3_mag_0.OUT 0.0203f
C652 JK_FF_mag_3.nand3_mag_2.OUT a_12159_4919# 0.0202f
C653 Q1 and2_mag_3.OUT 0.209f
C654 JK_FF_mag_3.K or_2_mag_3.IN2 1.08f
C655 JK_FF_mag_1.nand3_mag_1.IN1 a_6616_3820# 0.0697f
C656 a_9160_4915# JK_FF_mag_2.nand3_mag_1.OUT 1.5e-20
C657 JK_FF_mag_0.nand2_mag_3.IN1 a_2917_3818# 0.00119f
C658 JK_FF_mag_3.nand3_mag_1.OUT CLK 9.66e-19
C659 a_2751_4915# a_2911_4915# 0.0504f
C660 JK_FF_mag_0.nand3_mag_1.OUT CLK 0.0854f
C661 JK_FF_mag_2.nand2_mag_3.IN1 and2_mag_3.OUT 0.00359f
C662 a_12319_4919# JK_FF_mag_3.nand3_mag_1.OUT 1.5e-20
C663 JK_FF_mag_0.nand2_mag_1.IN2 Q2 6.62e-20
C664 a_8344_1618# Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 3.04e-20
C665 or_2_mag_3.IN1 CLK 0.748f
C666 JK_FF_mag_2.nand2_mag_1.IN2 CLK 0.00637f
C667 JK_FF_mag_0.nand3_mag_0.OUT or_2_mag_3.GF_INV_MAG_1.IN 2.76e-19
C668 a_9000_4915# JK_FF_mag_2.nand3_mag_1.OUT 1.17e-20
C669 Q0 JK_FF_mag_1.nand3_mag_0.OUT 3.38e-19
C670 RST JK_FF_mag_3.nand2_mag_3.IN1 0.00535f
C671 JK_FF_mag_1.nand2_mag_3.IN1 CLK 0.519f
C672 JK_FF_mag_2.nand3_mag_1.OUT VDD 0.994f
C673 JK_FF_mag_0.nand2_mag_1.IN2 a_4609_3818# 0.00372f
C674 nand3_mag_0.OUT CLK 1.69e-19
C675 JK_FF_mag_0.nand2_mag_3.IN1 Q1 0.00367f
C676 JK_FF_mag_3.QB a_12325_3822# 0.00392f
C677 Q1 and2_mag_1.GF_INV_MAG_0.IN 0.316f
C678 Q2 a_140_2787# 8.95e-19
C679 JK_FF_mag_0.nand2_mag_4.IN2 VDD 0.391f
C680 Q1 JK_FF_mag_2.nand3_mag_0.OUT 0.00101f
C681 JK_FF_mag_3.K JK_FF_mag_1.nand3_mag_0.OUT 8.26e-20
C682 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand3_mag_1.OUT 0.768f
C683 or_2_mag_0.IN2 Q2 0.149f
C684 JK_FF_mag_2.K JK_FF_mag_1.nand3_mag_1.OUT 3.72e-19
C685 JK_FF_mag_3.nand3_mag_1.OUT VDD 0.994f
C686 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand3_mag_0.OUT 0.0622f
C687 JK_FF_mag_3.K Q0 2.42f
C688 JK_FF_mag_0.nand2_mag_1.IN2 a_4045_3818# 0.069f
C689 nor_3_mag_0.OUT Q0 6.99e-20
C690 a_10858_3818# CLK 9.36e-19
C691 JK_FF_mag_0.nand3_mag_1.OUT VDD 0.994f
C692 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_1.K 3.6e-19
C693 a_3475_4915# CLK 6.8e-19
C694 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.nand2_mag_3.IN1 0.0894f
C695 a_6046_4917# JK_FF_mag_1.nand3_mag_1.OUT 1.5e-20
C696 or_2_mag_3.IN1 VDD 9.71f
C697 JK_FF_mag_2.nand3_mag_0.OUT JK_FF_mag_2.nand2_mag_3.IN1 0.0899f
C698 JK_FF_mag_0.nand2_mag_4.IN2 Q3 0.0635f
C699 JK_FF_mag_2.nand2_mag_1.IN2 VDD 0.397f
C700 or_2_mag_3.IN1 JK_FF_mag_3.nand3_mag_0.OUT 2.67e-20
C701 JK_FF_mag_1.QB a_7898_4917# 0.0811f
C702 Q0 nand3_mag_1.OUT 0.242f
C703 or_2_mag_1.IN1 and2_mag_1.GF_INV_MAG_0.IN 2.39e-20
C704 JK_FF_mag_3.K nor_3_mag_0.OUT 0.00134f
C705 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand3_mag_2.OUT 0.00158f
C706 JK_FF_mag_1.nand3_mag_1.IN1 a_6770_4917# 8.64e-19
C707 JK_FF_mag_1.nand2_mag_3.IN1 VDD 1.18f
C708 nand3_mag_0.OUT VDD 0.664f
C709 JK_FF_mag_0.nand3_mag_1.OUT Q3 0.0346f
C710 a_9724_4915# VDD 2.21e-19
C711 Q0 a_12159_4919# 0.00335f
C712 a_10294_3818# CLK 9.24e-19
C713 a_14017_3822# JK_FF_mag_3.nand2_mag_1.IN2 0.00372f
C714 JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_2.nand2_mag_4.IN2 0.122f
C715 JK_FF_mag_1.nand3_mag_1.IN1 CLK 0.0843f
C716 JK_FF_mag_2.K CLK 0.925f
C717 or_2_mag_3.IN1 Q3 0.0631f
C718 nor_3_mag_0.IN3 Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 0.104f
C719 a_7744_3820# JK_FF_mag_1.nand2_mag_4.IN2 4.52e-20
C720 JK_FF_mag_3.K nand3_mag_1.OUT 0.00452f
C721 JK_FF_mag_1.nand3_mag_0.OUT a_6616_3820# 0.00378f
C722 a_11012_4915# VDD 3.14e-19
C723 JK_FF_mag_1.QB a_7334_4917# 0.00964f
C724 or_2_mag_3.GF_INV_MAG_1.IN Q2 0.0515f
C725 and2_mag_3.GF_INV_MAG_0.IN GF_INV_MAG_1.OUT 1.48e-19
C726 or_2_mag_0.IN1 nand3_mag_0.OUT 0.00125f
C727 JK_FF_mag_3.nand3_mag_2.OUT CLK 0.237f
C728 JK_FF_mag_3.QB CLK 0.307f
C729 CLK a_6046_4917# 0.00164f
C730 nand3_mag_0.OUT Q3 0.00154f
C731 a_12883_4919# VDD 2.21e-19
C732 JK_FF_mag_3.K a_12159_4919# 8.64e-19
C733 JK_FF_mag_3.nand2_mag_4.IN2 VDD 0.391f
C734 JK_FF_mag_0.nand2_mag_3.IN1 RST 0.0694f
C735 a_3635_4915# Q3 0.0101f
C736 a_10858_3818# VDD 3.56e-19
C737 JK_FF_mag_1.QB JK_FF_mag_1.nand2_mag_1.IN2 0.0592f
C738 a_3475_4915# VDD 2.21e-19
C739 a_13453_3822# JK_FF_mag_3.nand2_mag_1.IN2 0.069f
C740 a_5886_4917# a_6046_4917# 0.0504f
C741 JK_FF_mag_3.nand3_mag_2.OUT a_12319_4919# 0.0731f
C742 JK_FF_mag_2.nand3_mag_1.IN1 CLK 0.0846f
C743 a_2757_3818# JK_FF_mag_0.K 0.00472f
C744 or_2_mag_3.GF_INV_MAG_1.IN or_2_mag_1.GF_INV_MAG_1.IN 5.88e-19
C745 JK_FF_mag_2.nand3_mag_0.OUT RST 5.36e-20
C746 Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN and2_mag_3.OUT 0.0022f
C747 and2_mag_3.IN1 Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.111f
C748 Q0 a_12325_3822# 2.79e-20
C749 Q1 JK_FF_mag_0.K 9.69e-19
C750 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_0.nand2_mag_4.IN2 8.16e-20
C751 and2_mag_0.GF_INV_MAG_0.IN nand3_mag_0.OUT 9.87e-20
C752 or_2_mag_3.IN1 JK_FF_mag_2.nand2_mag_4.IN2 0.198f
C753 JK_FF_mag_2.nand2_mag_1.IN2 JK_FF_mag_2.nand2_mag_4.IN2 8.16e-20
C754 or_2_mag_3.IN2 CLK 0.64f
C755 a_10294_3818# VDD 3.14e-19
C756 a_3475_4915# Q3 0.0102f
C757 a_3481_3818# JK_FF_mag_0.nand2_mag_3.IN1 1.43e-19
C758 a_9730_3818# JK_FF_mag_2.nand2_mag_3.IN1 1.43e-19
C759 JK_FF_mag_2.K a_9000_4915# 8.64e-19
C760 JK_FF_mag_0.nand2_mag_3.IN1 Q2 0.00952f
C761 JK_FF_mag_1.nand3_mag_1.IN1 VDD 0.651f
C762 JK_FF_mag_2.K VDD 0.866f
C763 JK_FF_mag_1.K JK_FF_mag_1.QB 7.07e-19
C764 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_0.nand3_mag_1.OUT 0.00975f
C765 JK_FF_mag_2.nand3_mag_2.OUT Q1 0.338f
C766 and2_mag_1.GF_INV_MAG_0.IN Q2 0.0549f
C767 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_1.nand3_mag_1.OUT 0.0622f
C768 JK_FF_mag_0.nand2_mag_3.IN1 a_4609_3818# 0.00118f
C769 Q0 JK_FF_mag_1.nand3_mag_1.OUT 3.92e-19
C770 JK_FF_mag_3.nand3_mag_2.OUT VDD 0.642f
C771 JK_FF_mag_3.QB VDD 0.904f
C772 JK_FF_mag_3.nand3_mag_2.OUT JK_FF_mag_3.nand3_mag_0.OUT 0.00183f
C773 JK_FF_mag_3.QB JK_FF_mag_3.nand3_mag_0.OUT 0.342f
C774 JK_FF_mag_0.nand2_mag_1.IN2 or_2_mag_3.IN1 6.23e-19
C775 a_8344_1618# and2_mag_3.GF_INV_MAG_0.IN 0.069f
C776 a_11012_4915# JK_FF_mag_2.nand2_mag_4.IN2 0.00372f
C777 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.K 0.0934f
C778 a_2911_4915# CLK 0.00253f
C779 JK_FF_mag_2.nand3_mag_2.OUT JK_FF_mag_2.nand2_mag_3.IN1 0.00118f
C780 JK_FF_mag_2.nand3_mag_1.IN1 VDD 0.651f
C781 JK_FF_mag_2.K Q3 0.0683f
C782 Q1 Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 7.38e-19
C783 a_10858_3818# JK_FF_mag_2.nand2_mag_4.IN2 4.52e-20
C784 and2_mag_1.GF_INV_MAG_0.IN a_1385_2540# 0.069f
C785 or_2_mag_1.GF_INV_MAG_1.IN and2_mag_1.GF_INV_MAG_0.IN 0.00165f
C786 a_4199_4915# RST 0.00162f
C787 JK_FF_mag_3.K JK_FF_mag_1.nand3_mag_1.OUT 9.58e-20
C788 a_14171_4919# VDD 3.14e-19
C789 JK_FF_mag_0.nand2_mag_3.IN1 a_4045_3818# 0.011f
C790 Q3 a_6046_4917# 4.52e-19
C791 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand2_mag_3.IN1 0.16f
C792 a_6610_4917# JK_FF_mag_1.nand3_mag_1.OUT 0.0203f
C793 or_2_mag_3.IN2 VDD 1.32f
C794 a_140_2787# nand3_mag_0.OUT 0.0732f
C795 JK_FF_mag_1.nand3_mag_0.OUT CLK 0.275f
C796 a_2751_4915# CLK 0.00224f
C797 Q0 CLK 0.538f
C798 or_2_mag_3.IN1 JK_FF_mag_3.nand2_mag_3.IN1 1.1e-19
C799 a_12889_3822# RST 2.67e-19
C800 Q1 a_2849_1480# 0.015f
C801 JK_FF_mag_1.nand2_mag_4.IN2 RST 0.0287f
C802 a_9730_3818# RST 3.68e-20
C803 JK_FF_mag_3.nand3_mag_1.IN1 JK_FF_mag_3.nand2_mag_1.IN2 0.109f
C804 or_2_mag_0.IN2 nand3_mag_0.OUT 0.139f
C805 JK_FF_mag_2.nand3_mag_1.OUT and2_mag_3.OUT 2.6e-20
C806 RST JK_FF_mag_0.K 0.00254f
C807 Q0 a_12319_4919# 0.00789f
C808 nor_3_mag_0.IN3 or_2_mag_3.IN1 6.71e-19
C809 Q3 or_2_mag_3.IN2 2.92f
C810 nor_3_mag_0.IN3 JK_FF_mag_2.nand2_mag_1.IN2 1.89e-20
C811 a_939_3715# Q0 3.17e-19
C812 a_6610_4917# a_6770_4917# 0.0504f
C813 RST a_12165_3822# 9.41e-19
C814 a_4763_4915# VDD 3.14e-19
C815 JK_FF_mag_3.K CLK 0.579f
C816 a_6616_3820# JK_FF_mag_1.nand3_mag_1.OUT 0.0195f
C817 a_9166_3818# JK_FF_mag_1.QB 1.16e-20
C818 Q1 a_1377_1477# 0.0186f
C819 JK_FF_mag_0.nand3_mag_1.IN1 Q1 1.86e-19
C820 JK_FF_mag_2.nand3_mag_2.OUT RST 0.0901f
C821 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_2.K 2.01e-19
C822 JK_FF_mag_1.nand2_mag_4.IN2 Q2 0.0635f
C823 nand3_mag_1.OUT CLK 0.32f
C824 JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_3.nand2_mag_4.IN2 0.321f
C825 or_2_mag_3.GF_INV_MAG_1.IN or_2_mag_3.IN1 0.211f
C826 and2_mag_3.IN1 GF_INV_MAG_1.OUT 0.00147f
C827 Q2 JK_FF_mag_0.K 0.0579f
C828 Q3 a_4763_4915# 0.0157f
C829 or_2_mag_0.GF_INV_MAG_1.IN Q0 0.00129f
C830 JK_FF_mag_1.nand3_mag_0.OUT VDD 0.648f
C831 a_2911_4915# Q3 0.0152f
C832 or_2_mag_3.IN1 and2_mag_3.OUT 0.00165f
C833 a_2751_4915# VDD 2.21e-19
C834 JK_FF_mag_2.nand2_mag_1.IN2 and2_mag_3.OUT 3.83e-19
C835 Q0 VDD 3.8f
C836 a_12159_4919# CLK 0.00117f
C837 Q0 JK_FF_mag_3.nand3_mag_0.OUT 0.00123f
C838 a_9006_3818# JK_FF_mag_1.QB 1.49e-20
C839 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand2_mag_4.IN2 0.321f
C840 JK_FF_mag_2.nand3_mag_0.OUT JK_FF_mag_2.nand3_mag_1.OUT 0.0622f
C841 JK_FF_mag_2.nand3_mag_2.OUT Q2 4.01e-20
C842 RST JK_FF_mag_3.nand3_mag_1.IN1 0.16f
C843 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.nand3_mag_1.IN1 0.122f
C844 a_12319_4919# a_12159_4919# 0.0504f
C845 or_2_mag_1.IN1 a_1377_1477# 0.0202f
C846 a_6616_3820# CLK 3.81e-19
C847 a_7744_3820# JK_FF_mag_1.nand2_mag_1.IN2 0.00372f
C848 and2_mag_3.IN1 and2_mag_3.GF_INV_MAG_0.IN 0.294f
C849 Q0 or_2_mag_0.IN1 0.0128f
C850 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C851 JK_FF_mag_3.K VDD 0.827f
C852 nor_3_mag_0.OUT VDD 0.343f
C853 Q0 Q3 0.128f
C854 a_2751_4915# Q3 0.0124f
C855 JK_FF_mag_3.K JK_FF_mag_3.nand3_mag_0.OUT 0.0951f
C856 JK_FF_mag_0.nand2_mag_1.IN2 or_2_mag_3.IN2 0.0593f
C857 a_6610_4917# VDD 2.21e-19
C858 a_7744_3820# JK_FF_mag_1.QB 0.0114f
C859 JK_FF_mag_0.nand2_mag_3.IN1 or_2_mag_3.IN1 0.0306f
C860 Q2 Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.101f
C861 JK_FF_mag_3.nand3_mag_2.OUT JK_FF_mag_3.nand2_mag_3.IN1 0.00118f
C862 JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_3.QB 0.28f
C863 Q1 GF_INV_MAG_1.OUT 3.09e-19
C864 and2_mag_1.GF_INV_MAG_0.IN or_2_mag_3.IN1 0.00126f
C865 nand3_mag_1.OUT VDD 1.19f
C866 and2_mag_2.GF_INV_MAG_0.IN a_1377_1477# 2.7e-20
C867 a_12325_3822# CLK 0.00939f
C868 Q0 and2_mag_0.GF_INV_MAG_0.IN 0.00115f
C869 a_7180_3820# JK_FF_mag_1.nand2_mag_1.IN2 0.069f
C870 nor_3_mag_0.OUT Q3 0.257f
C871 Q1 JK_FF_mag_1.nand2_mag_1.IN2 1.17e-19
C872 JK_FF_mag_0.nand2_mag_3.IN1 nand3_mag_0.OUT 5.63e-21
C873 JK_FF_mag_3.K Q3 0.076f
C874 and2_mag_3.IN1 a_8344_1618# 0.00476f
C875 JK_FF_mag_2.nand3_mag_0.OUT or_2_mag_3.IN1 0.343f
C876 and2_mag_1.GF_INV_MAG_0.IN nand3_mag_0.OUT 4.36e-19
C877 a_12159_4919# VDD 2.21e-19
C878 JK_FF_mag_0.nand3_mag_1.IN1 RST 0.188f
C879 a_6770_4917# JK_FF_mag_1.nand3_mag_1.OUT 0.0733f
C880 a_7180_3820# JK_FF_mag_1.QB 2.96e-19
C881 Q1 JK_FF_mag_1.QB 6.01e-19
C882 Q2 a_2849_1480# 0.0115f
C883 Q0 JK_FF_mag_2.nand2_mag_4.IN2 1.71e-21
C884 Q3 nand3_mag_1.OUT 0.299f
C885 Q1 and2_mag_3.GF_INV_MAG_0.IN 0.111f
C886 or_2_mag_3.GF_INV_MAG_1.IN JK_FF_mag_2.K 0.00584f
C887 a_6616_3820# VDD 3.14e-19
C888 CLK JK_FF_mag_1.nand3_mag_1.OUT 0.0834f
C889 JK_FF_mag_0.nand2_mag_4.IN2 a_4199_4915# 0.069f
C890 JK_FF_mag_3.nand3_mag_1.OUT a_13453_3822# 4.52e-20
C891 a_5886_4917# JK_FF_mag_1.nand3_mag_1.OUT 1.17e-20
C892 JK_FF_mag_1.K Q1 0.00825f
C893 JK_FF_mag_1.QB JK_FF_mag_2.nand2_mag_3.IN1 5.48e-20
C894 a_9730_3818# JK_FF_mag_2.nand3_mag_1.OUT 0.0195f
C895 JK_FF_mag_3.K JK_FF_mag_2.nand2_mag_4.IN2 1.32e-21
C896 RST a_7898_4917# 0.00106f
C897 JK_FF_mag_0.nand3_mag_1.OUT a_4199_4915# 0.00378f
C898 JK_FF_mag_0.nand2_mag_1.IN2 Q0 2.13e-20
C899 a_3481_3818# JK_FF_mag_0.nand3_mag_1.IN1 0.0697f
C900 Q1 a_n20_4333# 0.00347f
C901 or_2_mag_1.GF_INV_MAG_1.IN a_2849_1480# 2.4e-20
C902 Q2 a_1377_1477# 0.00186f
C903 JK_FF_mag_0.nand3_mag_1.IN1 Q2 1.12e-19
C904 Q1 a_8344_1618# 0.015f
C905 JK_FF_mag_2.nand3_mag_1.IN1 and2_mag_3.OUT 2.22e-20
C906 a_12325_3822# JK_FF_mag_3.nand3_mag_0.OUT 0.0732f
C907 JK_FF_mag_1.QB JK_FF_mag_1.nand3_mag_2.OUT 0.103f
C908 JK_FF_mag_3.nand3_mag_1.OUT a_12889_3822# 0.0195f
C909 a_9006_3818# a_9166_3818# 0.0504f
C910 a_14017_3822# JK_FF_mag_3.nand2_mag_4.IN2 4.52e-20
C911 Q0 a_140_2787# 0.0177f
C912 JK_FF_mag_2.nand3_mag_2.OUT JK_FF_mag_2.nand3_mag_1.OUT 0.121f
C913 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_2.K 0.00808f
C914 or_2_mag_3.GF_INV_MAG_1.IN or_2_mag_3.IN2 0.0432f
C915 Q0 a_7639_1615# 0.0121f
C916 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_3.K 8.28e-20
C917 JK_FF_mag_2.K and2_mag_1.GF_INV_MAG_0.IN 0.00253f
C918 RST a_7334_4917# 0.00106f
C919 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_1.K 3.43e-19
C920 JK_FF_mag_1.K JK_FF_mag_1.nand3_mag_2.OUT 0.105f
C921 or_2_mag_1.GF_INV_MAG_1.IN a_1377_1477# 0.132f
C922 Q2 a_7898_4917# 0.0157f
C923 a_5886_4917# CLK 0.00117f
C924 Q0 or_2_mag_0.IN2 0.0444f
C925 JK_FF_mag_1.nand3_mag_1.OUT VDD 0.994f
C926 JK_FF_mag_1.nand2_mag_4.IN2 or_2_mag_3.IN1 3.6e-21
C927 a_12319_4919# CLK 0.00164f
C928 a_9730_3818# or_2_mag_3.IN1 3.08e-19
C929 RST JK_FF_mag_1.nand2_mag_1.IN2 1.38e-19
C930 JK_FF_mag_2.K JK_FF_mag_2.nand3_mag_0.OUT 0.0998f
C931 Q0 JK_FF_mag_3.nand2_mag_3.IN1 0.0399f
C932 JK_FF_mag_1.QB a_6052_3820# 0.00392f
C933 JK_FF_mag_0.nand3_mag_1.IN1 a_4045_3818# 0.0059f
C934 a_939_3715# CLK 2.02e-20
C935 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.nand3_mag_2.OUT 0.00183f
C936 a_11081_1205# a_11241_1205# 0.186f
C937 a_9160_4915# CLK 0.00164f
C938 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.nand2_mag_4.IN2 0.321f
C939 a_12165_3822# or_2_mag_3.IN1 1.52e-20
C940 JK_FF_mag_2.nand3_mag_2.OUT a_9884_4915# 2.88e-20
C941 Q0 a_7479_1615# 0.00747f
C942 JK_FF_mag_1.QB RST 0.293f
C943 nor_3_mag_0.IN3 Q0 1.32e-19
C944 JK_FF_mag_3.nand3_mag_1.OUT a_13607_4919# 0.00378f
C945 Q2 a_7334_4917# 0.00859f
C946 JK_FF_mag_2.nand3_mag_2.OUT or_2_mag_3.IN1 0.103f
C947 JK_FF_mag_2.nand3_mag_1.IN1 JK_FF_mag_2.nand3_mag_0.OUT 0.122f
C948 a_14017_3822# JK_FF_mag_3.QB 0.0114f
C949 a_7639_1615# nand3_mag_1.OUT 0.0731f
C950 JK_FF_mag_3.K JK_FF_mag_3.nand2_mag_3.IN1 0.0715f
C951 JK_FF_mag_0.nand2_mag_3.IN1 or_2_mag_3.IN2 0.289f
C952 or_2_mag_0.GF_INV_MAG_1.IN CLK 0.0011f
C953 Q2 JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C954 JK_FF_mag_1.K RST 0.0767f
C955 a_9000_4915# CLK 0.00117f
C956 a_9166_3818# Q1 2.79e-20
C957 CLK VDD 5.61f
C958 JK_FF_mag_3.K nor_3_mag_0.IN3 1.82e-19
C959 JK_FF_mag_3.nand3_mag_0.OUT CLK 0.267f
C960 nor_3_mag_0.IN3 nor_3_mag_0.OUT 0.0121f
C961 JK_FF_mag_2.nand3_mag_2.OUT a_9724_4915# 9.1e-19
C962 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand3_mag_1.IN1 0.777f
C963 or_2_mag_3.GF_INV_MAG_1.IN Q0 0.0072f
C964 Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN GF_INV_MAG_1.OUT 0.116f
C965 a_5886_4917# VDD 2.21e-19
C966 or_2_mag_3.IN1 Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 1.74e-19
C967 JK_FF_mag_1.QB Q2 1.97f
C968 Q0 and2_mag_3.OUT 0.00187f
C969 JK_FF_mag_1.K a_5892_3820# 0.00472f
C970 or_2_mag_0.GF_INV_MAG_1.IN a_939_3715# 0.132f
C971 RST JK_FF_mag_0.nand3_mag_2.OUT 0.0571f
C972 a_13453_3822# JK_FF_mag_3.QB 2.96e-19
C973 a_7479_1615# nand3_mag_1.OUT 0.0202f
C974 nor_3_mag_0.IN3 nand3_mag_1.OUT 1.03e-19
C975 a_9166_3818# JK_FF_mag_2.nand2_mag_3.IN1 0.00119f
C976 a_939_3715# VDD 0.167f
C977 JK_FF_mag_0.nand2_mag_3.IN1 a_2911_4915# 8.66e-20
C978 or_2_mag_0.IN1 CLK 5.92e-19
C979 a_9000_4915# a_9160_4915# 0.0504f
C980 Q3 CLK 0.389f
C981 JK_FF_mag_3.K or_2_mag_3.GF_INV_MAG_1.IN 0.132f
C982 JK_FF_mag_1.K Q2 0.0398f
C983 a_13043_4919# JK_FF_mag_3.nand3_mag_1.IN1 8.64e-19
C984 Q3 a_5886_4917# 5.83e-19
C985 nor_3_mag_0.OUT and2_mag_3.OUT 0.163f
C986 Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN and2_mag_3.GF_INV_MAG_0.IN 4.69e-20
C987 JK_FF_mag_3.K and2_mag_3.OUT 0.00252f
C988 JK_FF_mag_2.K a_9730_3818# 1.39e-19
C989 JK_FF_mag_1.nand2_mag_4.IN2 JK_FF_mag_2.K 4.67e-22
C990 or_2_mag_3.IN1 a_2849_1480# 0.0131f
C991 Vdiv11 VSS 0.226f
C992 a_11241_1205# VSS 0.0376f
C993 a_11081_1205# VSS 0.0391f
C994 Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN VSS 0.676f
C995 GF_INV_MAG_1.OUT VSS 0.678f
C996 and2_mag_3.GF_INV_MAG_0.IN VSS 0.457f
C997 a_8344_1618# VSS 0.0693f
C998 nand3_mag_1.OUT VSS 0.741f
C999 a_7639_1615# VSS 0.0362f
C1000 a_7479_1615# VSS 0.0901f
C1001 and2_mag_3.IN1 VSS 0.834f
C1002 and2_mag_3.OUT VSS 1.93f
C1003 Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS 0.701f
C1004 a_2849_1480# VSS 0.0247f
C1005 a_1377_1477# VSS 0.0247f
C1006 nor_3_mag_0.OUT VSS 1.03f
C1007 nor_3_mag_0.IN3 VSS 0.555f
C1008 or_2_mag_3.GF_INV_MAG_1.IN VSS 0.597f
C1009 or_2_mag_1.GF_INV_MAG_1.IN VSS 0.589f
C1010 or_2_mag_1.IN1 VSS 0.532f
C1011 and2_mag_2.GF_INV_MAG_0.IN VSS 0.453f
C1012 a_n27_2146# VSS 0.0678f
C1013 a_1385_2540# VSS 0.0676f
C1014 a_140_2787# VSS 0.0343f
C1015 a_n20_2787# VSS 0.0881f
C1016 and2_mag_1.GF_INV_MAG_0.IN VSS 0.464f
C1017 a_14017_3822# VSS 0.0744f
C1018 a_13453_3822# VSS 0.0745f
C1019 a_12889_3822# VSS 0.0744f
C1020 JK_FF_mag_3.nand2_mag_1.IN2 VSS 0.425f
C1021 JK_FF_mag_3.nand3_mag_0.OUT VSS 0.549f
C1022 a_12325_3822# VSS 0.047f
C1023 a_12165_3822# VSS 0.101f
C1024 nand3_mag_0.OUT VSS 0.585f
C1025 a_10858_3818# VSS 0.0734f
C1026 a_10294_3818# VSS 0.0735f
C1027 a_9730_3818# VSS 0.0735f
C1028 JK_FF_mag_2.nand2_mag_1.IN2 VSS 0.424f
C1029 JK_FF_mag_2.nand3_mag_0.OUT VSS 0.543f
C1030 a_9166_3818# VSS 0.0449f
C1031 a_9006_3818# VSS 0.0987f
C1032 a_7744_3820# VSS 0.0739f
C1033 a_7180_3820# VSS 0.074f
C1034 a_6616_3820# VSS 0.0739f
C1035 JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.424f
C1036 JK_FF_mag_1.nand3_mag_0.OUT VSS 0.546f
C1037 a_6052_3820# VSS 0.0459f
C1038 a_5892_3820# VSS 0.0997f
C1039 a_4609_3818# VSS 0.0737f
C1040 a_4045_3818# VSS 0.0737f
C1041 a_3481_3818# VSS 0.0737f
C1042 JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.424f
C1043 JK_FF_mag_0.nand3_mag_0.OUT VSS 0.544f
C1044 a_2917_3818# VSS 0.0454f
C1045 a_2757_3818# VSS 0.0992f
C1046 a_939_3715# VSS 0.0247f
C1047 or_2_mag_0.GF_INV_MAG_1.IN VSS 0.612f
C1048 or_2_mag_0.IN2 VSS 0.402f
C1049 or_2_mag_0.IN1 VSS 0.511f
C1050 and2_mag_0.GF_INV_MAG_0.IN VSS 0.449f
C1051 a_n20_4333# VSS 0.0716f
C1052 JK_FF_mag_3.QB VSS 0.954f
C1053 a_14171_4919# VSS 0.0696f
C1054 a_13607_4919# VSS 0.0698f
C1055 JK_FF_mag_3.nand2_mag_4.IN2 VSS 0.42f
C1056 JK_FF_mag_3.nand2_mag_3.IN1 VSS 0.907f
C1057 JK_FF_mag_3.nand3_mag_1.OUT VSS 0.831f
C1058 a_13043_4919# VSS 0.0378f
C1059 a_12883_4919# VSS 0.0916f
C1060 a_12319_4919# VSS 0.0378f
C1061 a_12159_4919# VSS 0.0917f
C1062 or_2_mag_3.IN1 VSS 18.7f
C1063 a_11012_4915# VSS 0.069f
C1064 a_10448_4915# VSS 0.0691f
C1065 JK_FF_mag_2.nand2_mag_4.IN2 VSS 0.419f
C1066 JK_FF_mag_2.nand2_mag_3.IN1 VSS 0.86f
C1067 JK_FF_mag_2.nand3_mag_1.OUT VSS 0.827f
C1068 a_9884_4915# VSS 0.0367f
C1069 a_9724_4915# VSS 0.0905f
C1070 a_9160_4915# VSS 0.0368f
C1071 a_9000_4915# VSS 0.0906f
C1072 JK_FF_mag_1.QB VSS 0.912f
C1073 a_7898_4917# VSS 0.0693f
C1074 a_7334_4917# VSS 0.0694f
C1075 JK_FF_mag_3.nand3_mag_1.IN1 VSS 0.756f
C1076 JK_FF_mag_3.nand3_mag_2.OUT VSS 0.552f
C1077 Q0 VSS 8.73f
C1078 JK_FF_mag_3.K VSS 7.6f
C1079 JK_FF_mag_2.nand3_mag_1.IN1 VSS 0.743f
C1080 JK_FF_mag_2.nand3_mag_2.OUT VSS 0.549f
C1081 Q1 VSS 7.36f
C1082 JK_FF_mag_2.K VSS 2.89f
C1083 JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.42f
C1084 JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.832f
C1085 JK_FF_mag_1.nand3_mag_1.OUT VSS 0.829f
C1086 a_6770_4917# VSS 0.0372f
C1087 a_6610_4917# VSS 0.0911f
C1088 a_6046_4917# VSS 0.0373f
C1089 a_5886_4917# VSS 0.0911f
C1090 or_2_mag_3.IN2 VSS 2.53f
C1091 a_4763_4915# VSS 0.069f
C1092 a_4199_4915# VSS 0.0691f
C1093 JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.419f
C1094 JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.844f
C1095 JK_FF_mag_0.nand3_mag_1.OUT VSS 0.828f
C1096 a_3635_4915# VSS 0.0367f
C1097 a_3475_4915# VSS 0.0905f
C1098 a_2911_4915# VSS 0.0368f
C1099 a_2751_4915# VSS 0.0906f
C1100 JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.744f
C1101 JK_FF_mag_1.nand3_mag_2.OUT VSS 0.551f
C1102 Q2 VSS 7.49f
C1103 JK_FF_mag_1.K VSS 3.16f
C1104 JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.742f
C1105 RST VSS 2.97f
C1106 JK_FF_mag_0.nand3_mag_2.OUT VSS 0.548f
C1107 Q3 VSS 7.55f
C1108 CLK VSS 7.56f
C1109 JK_FF_mag_0.K VSS 1.92f
C1110 VDD VSS 77.3f
C1111 RST.n0 VSS 0.0309f
C1112 RST.t7 VSS 0.019f
C1113 RST.t4 VSS 0.0125f
C1114 RST.n1 VSS 0.0335f
C1115 RST.n2 VSS 0.00617f
C1116 RST.n3 VSS 0.00211f
C1117 RST.n4 VSS 0.00774f
C1118 RST.n5 VSS 0.0118f
C1119 RST.n6 VSS 0.0069f
C1120 RST.n7 VSS 0.00257f
C1121 RST.t2 VSS 0.019f
C1122 RST.t3 VSS 0.0125f
C1123 RST.n8 VSS 0.0335f
C1124 RST.n9 VSS 0.00474f
C1125 RST.n10 VSS 0.00184f
C1126 RST.n11 VSS 0.00258f
C1127 RST.n12 VSS 0.009f
C1128 RST.n13 VSS 7.93e-19
C1129 RST.n14 VSS 0.0237f
C1130 RST.n15 VSS 0.478f
C1131 RST.n16 VSS 0.475f
C1132 RST.n17 VSS 0.00227f
C1133 RST.n18 VSS 0.00685f
C1134 RST.n19 VSS 0.00169f
C1135 RST.t1 VSS 0.019f
C1136 RST.t0 VSS 0.0125f
C1137 RST.n20 VSS 0.0335f
C1138 RST.n21 VSS 0.00525f
C1139 RST.n22 VSS 0.00488f
C1140 RST.n23 VSS 0.00751f
C1141 RST.n24 VSS 0.00532f
C1142 RST.n25 VSS 0.47f
C1143 RST.n26 VSS 0.47f
C1144 RST.n27 VSS 0.469f
C1145 RST.n28 VSS 0.473f
C1146 RST.n29 VSS 0.00704f
C1147 RST.n30 VSS 0.00805f
C1148 RST.n31 VSS 0.00268f
C1149 RST.t6 VSS 0.019f
C1150 RST.t5 VSS 0.0125f
C1151 RST.n32 VSS 0.0335f
C1152 RST.n33 VSS 0.00468f
C1153 RST.n34 VSS 0.0016f
C1154 RST.n35 VSS 7.93e-19
C1155 RST.n36 VSS 0.00218f
C1156 RST.n37 VSS 0.00515f
C1157 RST.n38 VSS 9.09e-19
C1158 RST.n39 VSS 0.0599f
C1159 RST.n40 VSS 0.0464f
C1160 or_2_mag_3.IN1.t3 VSS 0.0462f
C1161 or_2_mag_3.IN1.t8 VSS 0.154f
C1162 or_2_mag_3.IN1.n0 VSS 0.159f
C1163 or_2_mag_3.IN1.t6 VSS 0.0699f
C1164 or_2_mag_3.IN1.t7 VSS 0.11f
C1165 or_2_mag_3.IN1.n1 VSS 0.194f
C1166 or_2_mag_3.IN1.t4 VSS 0.0624f
C1167 or_2_mag_3.IN1.t5 VSS 0.0782f
C1168 or_2_mag_3.IN1.n2 VSS 0.185f
C1169 or_2_mag_3.IN1.n3 VSS 1.79f
C1170 or_2_mag_3.IN1.t1 VSS 0.507f
C1171 Q3.t12 VSS 0.012f
C1172 Q3.t11 VSS 0.0631f
C1173 Q3.n0 VSS 0.0501f
C1174 Q3.n1 VSS 0.00745f
C1175 Q3.n2 VSS 0.0122f
C1176 Q3.t9 VSS 0.0297f
C1177 Q3.t8 VSS 0.0196f
C1178 Q3.n3 VSS 0.0527f
C1179 Q3.n4 VSS 0.0246f
C1180 Q3.n5 VSS 0.0052f
C1181 Q3.t3 VSS 0.017f
C1182 Q3.t6 VSS 0.0214f
C1183 Q3.n6 VSS 0.049f
C1184 Q3.n7 VSS 0.468f
C1185 Q3.n8 VSS 0.507f
C1186 Q3.n9 VSS 0.00242f
C1187 Q3.t7 VSS 0.017f
C1188 Q3.t10 VSS 0.0214f
C1189 Q3.n10 VSS 0.0489f
C1190 Q3.n11 VSS 0.0191f
C1191 Q3.n12 VSS 0.518f
C1192 Q3.n13 VSS 0.742f
C1193 Q3.t4 VSS 0.017f
C1194 Q3.t5 VSS 0.0214f
C1195 Q3.n14 VSS 0.0494f
C1196 Q3.n15 VSS 0.0307f
C1197 Q3.n16 VSS 0.306f
C1198 Q3.n17 VSS 0.0162f
C1199 Q3.t1 VSS 0.0133f
C1200 Q3.n18 VSS 0.0133f
C1201 Q3.n19 VSS 0.032f
C1202 Q3.n20 VSS 0.0997f
C1203 Q3.n21 VSS 0.012f
C1204 Q3.n22 VSS 1.94f
C1205 Q3.n23 VSS 1.69f
C1206 Q3.n24 VSS 0.00308f
C1207 Q3.n25 VSS 0.00456f
C1208 Q0.t11 VSS 0.0536f
C1209 Q0.t10 VSS 0.0353f
C1210 Q0.n0 VSS 0.0948f
C1211 Q0.n1 VSS 0.0127f
C1212 Q0.n2 VSS 0.0292f
C1213 Q0.t1 VSS 0.0241f
C1214 Q0.n3 VSS 0.0241f
C1215 Q0.n4 VSS 0.0578f
C1216 Q0.n5 VSS 0.18f
C1217 Q0.n6 VSS 0.0219f
C1218 Q0.t5 VSS 0.0536f
C1219 Q0.t12 VSS 0.0353f
C1220 Q0.n7 VSS 0.0952f
C1221 Q0.n8 VSS 0.373f
C1222 Q0.t14 VSS 0.0308f
C1223 Q0.t13 VSS 0.0386f
C1224 Q0.n9 VSS 0.0892f
C1225 Q0.n10 VSS 0.0554f
C1226 Q0.n11 VSS 0.679f
C1227 Q0.n12 VSS 0.377f
C1228 Q0.t3 VSS 0.0502f
C1229 Q0.t9 VSS 0.0274f
C1230 Q0.n13 VSS 0.0949f
C1231 Q0.n14 VSS 0.0274f
C1232 Q0.n15 VSS 0.0053f
C1233 Q0.t4 VSS 0.0353f
C1234 Q0.t6 VSS 0.0536f
C1235 Q0.n16 VSS 0.0949f
C1236 Q0.n17 VSS 0.0188f
C1237 Q0.n18 VSS 0.00464f
C1238 Q0.n19 VSS 0.502f
C1239 Q0.n20 VSS 0.204f
C1240 Q0.t8 VSS 0.0129f
C1241 Q0.t7 VSS 0.0878f
C1242 Q0.n21 VSS 0.0733f
C1243 Q0.n22 VSS 1.82f
C1244 Q0.n23 VSS 6.05f
C1245 Q0.n24 VSS 0.0192f
C1246 Q0.n25 VSS 0.517f
C1247 Q0.n26 VSS 0.0046f
C1248 Q0.n27 VSS 0.00856f
C1249 Q1.t14 VSS 0.0299f
C1250 Q1.t13 VSS 0.0547f
C1251 Q1.n0 VSS 0.104f
C1252 Q1.t6 VSS 0.0547f
C1253 Q1.t12 VSS 0.0415f
C1254 Q1.n1 VSS 0.108f
C1255 Q1.t16 VSS 0.0299f
C1256 Q1.t15 VSS 0.0547f
C1257 Q1.n2 VSS 0.103f
C1258 Q1.n3 VSS 0.234f
C1259 Q1.n4 VSS 0.769f
C1260 Q1.n5 VSS 0.00545f
C1261 Q1.n6 VSS 0.00467f
C1262 Q1.t5 VSS 0.0335f
C1263 Q1.t11 VSS 0.042f
C1264 Q1.n7 VSS 0.0993f
C1265 Q1.n8 VSS 0.0372f
C1266 Q1.n9 VSS 0.00755f
C1267 Q1.n10 VSS 0.853f
C1268 Q1.n11 VSS 0.597f
C1269 Q1.t10 VSS 0.0584f
C1270 Q1.t9 VSS 0.0385f
C1271 Q1.n12 VSS 0.104f
C1272 Q1.n13 VSS 0.407f
C1273 Q1.t7 VSS 0.0335f
C1274 Q1.t8 VSS 0.042f
C1275 Q1.n14 VSS 0.0972f
C1276 Q1.n15 VSS 0.0604f
C1277 Q1.n16 VSS 0.768f
C1278 Q1.n17 VSS 0.0318f
C1279 Q1.t2 VSS 0.0262f
C1280 Q1.n18 VSS 0.0262f
C1281 Q1.n19 VSS 0.0629f
C1282 Q1.n20 VSS 0.196f
C1283 Q1.n21 VSS 0.0236f
C1284 Q1.n22 VSS 0.75f
C1285 Q1.t4 VSS 0.0309f
C1286 Q1.t3 VSS 0.0536f
C1287 Q1.n23 VSS 0.103f
C1288 Q1.n24 VSS 0.4f
C1289 Q1.n25 VSS 4.87f
C1290 Q1.n26 VSS 3.32f
C1291 Q2.t4 VSS 0.0473f
C1292 Q2.t3 VSS 0.0312f
C1293 Q2.n0 VSS 0.084f
C1294 Q2.n1 VSS 0.329f
C1295 Q2.t5 VSS 0.0272f
C1296 Q2.t6 VSS 0.034f
C1297 Q2.n2 VSS 0.0787f
C1298 Q2.n3 VSS 0.0489f
C1299 Q2.n4 VSS 0.612f
C1300 Q2.t8 VSS 0.0424f
C1301 Q2.t7 VSS 0.141f
C1302 Q2.n5 VSS 0.171f
C1303 Q2.n6 VSS 0.00472f
C1304 Q2.t9 VSS 0.0312f
C1305 Q2.t10 VSS 0.0473f
C1306 Q2.n7 VSS 0.0808f
C1307 Q2.n8 VSS 0.0139f
C1308 Q2.n9 VSS 0.00393f
C1309 Q2.n10 VSS 0.0097f
C1310 Q2.n11 VSS 1.89f
C1311 Q2.n12 VSS 3.87f
C1312 Q2.n13 VSS 0.891f
C1313 Q2.n14 VSS 0.0258f
C1314 Q2.t1 VSS 0.0212f
C1315 Q2.n15 VSS 0.0212f
C1316 Q2.n16 VSS 0.051f
C1317 Q2.n17 VSS 0.159f
C1318 Q2.n18 VSS 0.0199f
C1319 JK_FF_mag_1.K.t3 VSS 0.0207f
C1320 JK_FF_mag_1.K.t2 VSS 0.0273f
C1321 JK_FF_mag_1.K.n0 VSS 0.0537f
C1322 JK_FF_mag_1.K.t5 VSS 0.0207f
C1323 JK_FF_mag_1.K.t4 VSS 0.0271f
C1324 JK_FF_mag_1.K.n1 VSS 0.0537f
C1325 JK_FF_mag_1.K.n2 VSS 0.675f
C1326 JK_FF_mag_3.K.t3 VSS 0.0552f
C1327 JK_FF_mag_3.K.t2 VSS 0.0727f
C1328 JK_FF_mag_3.K.n0 VSS 0.143f
C1329 JK_FF_mag_3.K.t5 VSS 0.0553f
C1330 JK_FF_mag_3.K.t4 VSS 0.0722f
C1331 JK_FF_mag_3.K.n1 VSS 0.143f
C1332 JK_FF_mag_3.K.n2 VSS 5.28f
C1333 JK_FF_mag_3.K.n3 VSS 0.0872f
C1334 VDD.t153 VSS 0.0793f
C1335 VDD.t154 VSS 0.00889f
C1336 VDD.t197 VSS 0.00853f
C1337 VDD.t136 VSS 0.0186f
C1338 VDD.n0 VSS 0.107f
C1339 VDD.t29 VSS 0.00367f
C1340 VDD.n1 VSS 0.00367f
C1341 VDD.n2 VSS 0.00969f
C1342 VDD.t28 VSS -0.00413f
C1343 VDD.t181 VSS 0.0611f
C1344 VDD.t84 VSS 0.107f
C1345 VDD.n3 VSS 0.0554f
C1346 VDD.n4 VSS 0.0208f
C1347 VDD.n5 VSS 0.00892f
C1348 VDD.n6 VSS 0.0308f
C1349 VDD.t193 VSS 0.00968f
C1350 VDD.n7 VSS 0.0199f
C1351 VDD.t137 VSS 0.0589f
C1352 VDD.t46 VSS 0.114f
C1353 VDD.n8 VSS 0.0167f
C1354 VDD.t47 VSS 0.0186f
C1355 VDD.t169 VSS 0.0194f
C1356 VDD.t138 VSS 0.0172f
C1357 VDD.n9 VSS 0.0311f
C1358 VDD.n10 VSS 0.0191f
C1359 VDD.n11 VSS 0.0813f
C1360 VDD.t170 VSS 0.105f
C1361 VDD.t171 VSS 0.00889f
C1362 VDD.n12 VSS 0.0687f
C1363 VDD.n13 VSS 0.0693f
C1364 VDD.t41 VSS 0.217f
C1365 VDD.t40 VSS 0.0724f
C1366 VDD.n14 VSS 0.00596f
C1367 VDD.n15 VSS 0.00166f
C1368 VDD.t195 VSS 0.0362f
C1369 VDD.n16 VSS 0.0542f
C1370 VDD.n17 VSS 0.0465f
C1371 VDD.n18 VSS 0.0839f
C1372 VDD.t194 VSS 0.227f
C1373 VDD.n19 VSS 0.133f
C1374 VDD.n20 VSS 0.0639f
C1375 VDD.n21 VSS 0.0556f
C1376 VDD.n22 VSS 0.126f
C1377 VDD.t168 VSS 0.0625f
C1378 VDD.n23 VSS 0.0831f
C1379 VDD.t0 VSS 0.084f
C1380 VDD.t192 VSS 0.0962f
C1381 VDD.n24 VSS 0.0738f
C1382 VDD.t81 VSS 0.11f
C1383 VDD.n25 VSS 0.0953f
C1384 VDD.t1 VSS 0.00889f
C1385 VDD.n26 VSS 0.0305f
C1386 VDD.n27 VSS 0.124f
C1387 VDD.n28 VSS 0.143f
C1388 VDD.n29 VSS 0.16f
C1389 VDD.t85 VSS 0.00916f
C1390 VDD.n30 VSS 0.0413f
C1391 VDD.t135 VSS 0.123f
C1392 VDD.t196 VSS 0.044f
C1393 VDD.n31 VSS 0.126f
C1394 VDD.n32 VSS 0.0658f
C1395 VDD.n33 VSS 0.0771f
C1396 VDD.t226 VSS 0.00367f
C1397 VDD.n34 VSS 0.00367f
C1398 VDD.n35 VSS 0.00802f
C1399 VDD.n36 VSS 0.0344f
C1400 VDD.t234 VSS 0.118f
C1401 VDD.n37 VSS 0.00892f
C1402 VDD.t126 VSS 0.00893f
C1403 VDD.n38 VSS 0.00892f
C1404 VDD.n39 VSS 0.0487f
C1405 VDD.t227 VSS 0.116f
C1406 VDD.n40 VSS 0.00892f
C1407 VDD.n41 VSS 0.00892f
C1408 VDD.t110 VSS 0.116f
C1409 VDD.n42 VSS 0.0554f
C1410 VDD.t128 VSS 0.00893f
C1411 VDD.n43 VSS 0.00892f
C1412 VDD.t127 VSS 0.108f
C1413 VDD.t129 VSS 0.118f
C1414 VDD.n44 VSS 0.0554f
C1415 VDD.t238 VSS 0.00893f
C1416 VDD.t124 VSS 0.00367f
C1417 VDD.n45 VSS 0.00367f
C1418 VDD.n46 VSS 0.00802f
C1419 VDD.t237 VSS 0.108f
C1420 VDD.t123 VSS 0.131f
C1421 VDD.t54 VSS 0.0611f
C1422 VDD.n47 VSS 0.0554f
C1423 VDD.t156 VSS 0.00893f
C1424 VDD.t240 VSS 0.00367f
C1425 VDD.n48 VSS 0.00367f
C1426 VDD.n49 VSS 0.00802f
C1427 VDD.t155 VSS 0.108f
C1428 VDD.t239 VSS 0.131f
C1429 VDD.t37 VSS 0.0611f
C1430 VDD.t215 VSS 0.107f
C1431 VDD.n50 VSS 0.0554f
C1432 VDD.t216 VSS 0.00957f
C1433 VDD.n51 VSS 0.0687f
C1434 VDD.n52 VSS 0.0509f
C1435 VDD.n53 VSS 0.0522f
C1436 VDD.n54 VSS 0.0277f
C1437 VDD.n55 VSS 0.0509f
C1438 VDD.n56 VSS 0.0521f
C1439 VDD.n57 VSS 0.0308f
C1440 VDD.n58 VSS 0.0442f
C1441 VDD.n59 VSS 0.0411f
C1442 VDD.n60 VSS 0.0308f
C1443 VDD.n61 VSS 0.0774f
C1444 VDD.t31 VSS 0.00889f
C1445 VDD.t140 VSS 0.00893f
C1446 VDD.n62 VSS 0.0517f
C1447 VDD.t30 VSS 0.079f
C1448 VDD.t20 VSS 0.0611f
C1449 VDD.t99 VSS 0.00367f
C1450 VDD.n63 VSS 0.00367f
C1451 VDD.n64 VSS 0.00802f
C1452 VDD.t220 VSS 0.00893f
C1453 VDD.n65 VSS 0.00892f
C1454 VDD.n66 VSS 0.0484f
C1455 VDD.t251 VSS 0.118f
C1456 VDD.n67 VSS 0.00892f
C1457 VDD.t158 VSS 0.00893f
C1458 VDD.n68 VSS 0.00892f
C1459 VDD.n69 VSS 0.00892f
C1460 VDD.t173 VSS 0.0938f
C1461 VDD.n70 VSS 0.0478f
C1462 VDD.t51 VSS 0.00893f
C1463 VDD.n71 VSS 0.00892f
C1464 VDD.t50 VSS 0.0856f
C1465 VDD.t254 VSS 0.0938f
C1466 VDD.n72 VSS 0.0478f
C1467 VDD.t114 VSS 0.00893f
C1468 VDD.t247 VSS 0.00367f
C1469 VDD.n73 VSS 0.00367f
C1470 VDD.n74 VSS 0.00802f
C1471 VDD.n75 VSS 0.0478f
C1472 VDD.t207 VSS 0.00893f
C1473 VDD.t94 VSS 0.00367f
C1474 VDD.n76 VSS 0.00367f
C1475 VDD.n77 VSS 0.00802f
C1476 VDD.t206 VSS 0.0856f
C1477 VDD.t93 VSS 0.105f
C1478 VDD.t23 VSS 0.0486f
C1479 VDD.t113 VSS 0.078f
C1480 VDD.t78 VSS 0.0486f
C1481 VDD.t246 VSS 0.0373f
C1482 VDD.n78 VSS 0.308f
C1483 VDD.t141 VSS 0.0982f
C1484 VDD.n79 VSS 0.0478f
C1485 VDD.t142 VSS 0.00957f
C1486 VDD.n80 VSS 0.0687f
C1487 VDD.n81 VSS 0.0509f
C1488 VDD.n82 VSS 0.0522f
C1489 VDD.n83 VSS 0.0277f
C1490 VDD.n84 VSS 0.0509f
C1491 VDD.n85 VSS 0.0521f
C1492 VDD.n86 VSS 0.0308f
C1493 VDD.n87 VSS 0.0442f
C1494 VDD.n88 VSS 0.0411f
C1495 VDD.n89 VSS 0.0308f
C1496 VDD.n90 VSS 0.105f
C1497 VDD.t27 VSS 0.00889f
C1498 VDD.t189 VSS 0.00893f
C1499 VDD.n91 VSS 0.0525f
C1500 VDD.t26 VSS 0.079f
C1501 VDD.t14 VSS 0.0611f
C1502 VDD.t101 VSS 0.00367f
C1503 VDD.n92 VSS 0.00367f
C1504 VDD.n93 VSS 0.00802f
C1505 VDD.t75 VSS 0.00893f
C1506 VDD.n94 VSS 0.00892f
C1507 VDD.n95 VSS 0.0491f
C1508 VDD.t57 VSS 0.118f
C1509 VDD.n96 VSS 0.00892f
C1510 VDD.t233 VSS 0.00893f
C1511 VDD.n97 VSS 0.00892f
C1512 VDD.n98 VSS 0.00892f
C1513 VDD.t95 VSS 0.116f
C1514 VDD.n99 VSS 0.0554f
C1515 VDD.t77 VSS 0.00893f
C1516 VDD.n100 VSS 0.00892f
C1517 VDD.t76 VSS 0.108f
C1518 VDD.t60 VSS 0.118f
C1519 VDD.n101 VSS 0.0554f
C1520 VDD.t177 VSS 0.00893f
C1521 VDD.t144 VSS 0.00367f
C1522 VDD.n102 VSS 0.00367f
C1523 VDD.n103 VSS 0.00802f
C1524 VDD.t176 VSS 0.108f
C1525 VDD.t143 VSS 0.131f
C1526 VDD.t248 VSS 0.0611f
C1527 VDD.n104 VSS 0.0554f
C1528 VDD.t3 VSS 0.00893f
C1529 VDD.t106 VSS 0.00367f
C1530 VDD.n105 VSS 0.00367f
C1531 VDD.n106 VSS 0.00802f
C1532 VDD.t2 VSS 0.108f
C1533 VDD.t105 VSS 0.131f
C1534 VDD.t6 VSS 0.0611f
C1535 VDD.t213 VSS 0.107f
C1536 VDD.n107 VSS 0.0554f
C1537 VDD.t214 VSS 0.00957f
C1538 VDD.n108 VSS 0.0687f
C1539 VDD.n109 VSS 0.0509f
C1540 VDD.n110 VSS 0.0522f
C1541 VDD.n111 VSS 0.0277f
C1542 VDD.n112 VSS 0.0509f
C1543 VDD.n113 VSS 0.0521f
C1544 VDD.n114 VSS 0.0308f
C1545 VDD.n115 VSS 0.0442f
C1546 VDD.n116 VSS 0.0411f
C1547 VDD.n117 VSS 0.0308f
C1548 VDD.n118 VSS 0.105f
C1549 VDD.n119 VSS 0.121f
C1550 VDD.t102 VSS 0.116f
C1551 VDD.t232 VSS 0.108f
C1552 VDD.n120 VSS 0.0554f
C1553 VDD.n121 VSS 0.033f
C1554 VDD.n122 VSS 0.0455f
C1555 VDD.n123 VSS 0.0491f
C1556 VDD.t146 VSS 0.00893f
C1557 VDD.n124 VSS 0.0455f
C1558 VDD.n125 VSS 0.033f
C1559 VDD.n126 VSS 0.0554f
C1560 VDD.t145 VSS 0.108f
C1561 VDD.t178 VSS 0.118f
C1562 VDD.t100 VSS 0.131f
C1563 VDD.t74 VSS 0.108f
C1564 VDD.n127 VSS 0.0554f
C1565 VDD.n128 VSS 0.033f
C1566 VDD.n129 VSS 0.0429f
C1567 VDD.n130 VSS 0.0408f
C1568 VDD.n131 VSS 0.0293f
C1569 VDD.n132 VSS 0.0554f
C1570 VDD.t188 VSS 0.0611f
C1571 VDD.n133 VSS 0.0829f
C1572 VDD.n134 VSS 0.0499f
C1573 VDD.n135 VSS 0.0557f
C1574 VDD.n136 VSS 0.0497f
C1575 VDD.t198 VSS 0.116f
C1576 VDD.t157 VSS 0.108f
C1577 VDD.n137 VSS 0.0554f
C1578 VDD.n138 VSS 0.0327f
C1579 VDD.n139 VSS 0.0448f
C1580 VDD.n140 VSS 0.0484f
C1581 VDD.t245 VSS 0.00893f
C1582 VDD.n141 VSS 0.0448f
C1583 VDD.n142 VSS 0.0327f
C1584 VDD.n143 VSS 0.0554f
C1585 VDD.t244 VSS 0.108f
C1586 VDD.t115 VSS 0.118f
C1587 VDD.t98 VSS 0.131f
C1588 VDD.t219 VSS 0.108f
C1589 VDD.n144 VSS 0.0554f
C1590 VDD.n145 VSS 0.0327f
C1591 VDD.n146 VSS 0.0423f
C1592 VDD.n147 VSS 0.0401f
C1593 VDD.n148 VSS 0.0291f
C1594 VDD.n149 VSS 0.0554f
C1595 VDD.t139 VSS 0.0611f
C1596 VDD.n150 VSS 0.0829f
C1597 VDD.n151 VSS 0.0478f
C1598 VDD.n152 VSS 0.0784f
C1599 VDD.n153 VSS 0.0476f
C1600 VDD.t148 VSS 0.00893f
C1601 VDD.n154 VSS 0.0451f
C1602 VDD.n155 VSS 0.0328f
C1603 VDD.n156 VSS 0.0554f
C1604 VDD.t147 VSS 0.108f
C1605 VDD.t132 VSS 0.118f
C1606 VDD.t125 VSS 0.108f
C1607 VDD.n157 VSS 0.0554f
C1608 VDD.n158 VSS 0.0328f
C1609 VDD.n159 VSS 0.0451f
C1610 VDD.n160 VSS 0.0487f
C1611 VDD.t205 VSS 0.00893f
C1612 VDD.n161 VSS 0.0426f
C1613 VDD.n162 VSS 0.0328f
C1614 VDD.n163 VSS 0.0554f
C1615 VDD.t204 VSS 0.108f
C1616 VDD.t225 VSS 0.131f
C1617 VDD.t34 VSS 0.0611f
C1618 VDD.n164 VSS 0.0554f
C1619 VDD.t88 VSS 0.00893f
C1620 VDD.t87 VSS 0.0611f
C1621 VDD.t32 VSS 0.079f
C1622 VDD.n165 VSS 0.0829f
C1623 VDD.t33 VSS 0.00889f
C1624 VDD.n166 VSS 0.00892f
C1625 VDD.t63 VSS 0.0938f
C1626 VDD.n167 VSS 0.0478f
C1627 VDD.t191 VSS 0.00893f
C1628 VDD.n168 VSS 0.00892f
C1629 VDD.t190 VSS 0.0856f
C1630 VDD.t260 VSS 0.0938f
C1631 VDD.n169 VSS 0.0478f
C1632 VDD.t122 VSS 0.00893f
C1633 VDD.t187 VSS 0.00367f
C1634 VDD.n170 VSS 0.00367f
C1635 VDD.n171 VSS 0.00802f
C1636 VDD.n172 VSS 0.0478f
C1637 VDD.t231 VSS 0.00893f
C1638 VDD.t109 VSS 0.00367f
C1639 VDD.n173 VSS 0.00367f
C1640 VDD.n174 VSS 0.00802f
C1641 VDD.t230 VSS 0.0856f
C1642 VDD.t108 VSS 0.105f
C1643 VDD.t17 VSS 0.0486f
C1644 VDD.t121 VSS 0.078f
C1645 VDD.t201 VSS 0.0486f
C1646 VDD.t186 VSS 0.0373f
C1647 VDD.n175 VSS 0.308f
C1648 VDD.t223 VSS 0.0982f
C1649 VDD.n176 VSS 0.0478f
C1650 VDD.t224 VSS 0.00957f
C1651 VDD.n177 VSS 0.0687f
C1652 VDD.n178 VSS 0.0509f
C1653 VDD.n179 VSS 0.0522f
C1654 VDD.n180 VSS 0.0277f
C1655 VDD.n181 VSS 0.0509f
C1656 VDD.n182 VSS 0.0521f
C1657 VDD.n183 VSS 0.0308f
C1658 VDD.n184 VSS 0.0442f
C1659 VDD.n185 VSS 0.0411f
C1660 VDD.n186 VSS 0.0308f
C1661 VDD.n187 VSS 0.0774f
C1662 VDD.n188 VSS 0.00892f
C1663 VDD.t159 VSS 0.116f
C1664 VDD.n189 VSS 0.0554f
C1665 VDD.t264 VSS 0.00893f
C1666 VDD.n190 VSS 0.00892f
C1667 VDD.t263 VSS 0.108f
C1668 VDD.t257 VSS 0.118f
C1669 VDD.n191 VSS 0.0554f
C1670 VDD.t185 VSS 0.00893f
C1671 VDD.n192 VSS 0.00892f
C1672 VDD.t184 VSS 0.108f
C1673 VDD.t118 VSS 0.118f
C1674 VDD.n193 VSS 0.0554f
C1675 VDD.t92 VSS 0.00893f
C1676 VDD.t163 VSS 0.00367f
C1677 VDD.n194 VSS 0.00367f
C1678 VDD.n195 VSS 0.00802f
C1679 VDD.t91 VSS 0.108f
C1680 VDD.t162 VSS 0.131f
C1681 VDD.t11 VSS 0.0611f
C1682 VDD.n196 VSS 0.0554f
C1683 VDD.t222 VSS 0.00893f
C1684 VDD.t221 VSS 0.0611f
C1685 VDD.t9 VSS 0.079f
C1686 VDD.n197 VSS 0.0781f
C1687 VDD.n198 VSS 0.0736f
C1688 VDD.t10 VSS 0.00889f
C1689 VDD.t218 VSS 0.0112f
C1690 VDD.n199 VSS 0.0452f
C1691 VDD.n200 VSS 0.00892f
C1692 VDD.t217 VSS 0.0854f
C1693 VDD.n201 VSS 0.0811f
C1694 VDD.t208 VSS 0.0699f
C1695 VDD.t4 VSS 0.107f
C1696 VDD.n202 VSS 0.0554f
C1697 VDD.t49 VSS 0.00889f
C1698 VDD.n203 VSS 0.0291f
C1699 VDD.n204 VSS 0.0955f
C1700 VDD.t67 VSS 0.0213f
C1701 VDD.t152 VSS 0.00889f
C1702 VDD.n205 VSS 0.00892f
C1703 VDD.t45 VSS 0.00367f
C1704 VDD.n206 VSS 0.00367f
C1705 VDD.n207 VSS 0.00802f
C1706 VDD.n208 VSS 0.0669f
C1707 VDD.t53 VSS 0.00889f
C1708 VDD.t241 VSS 0.215f
C1709 VDD.t243 VSS 0.00893f
C1710 VDD.t242 VSS 0.00893f
C1711 VDD.n209 VSS 0.0822f
C1712 VDD.n210 VSS 0.0376f
C1713 VDD.n211 VSS 0.111f
C1714 VDD.t68 VSS 0.122f
C1715 VDD.t44 VSS 0.169f
C1716 VDD.t52 VSS 0.119f
C1717 VDD.t66 VSS 0.0287f
C1718 VDD.t48 VSS 0.0793f
C1719 VDD.n213 VSS 0.0937f
C1720 VDD.t172 VSS 0.0746f
C1721 VDD.n214 VSS 0.0322f
C1722 VDD.n215 VSS 0.112f
C1723 VDD.n216 VSS 0.0662f
C1724 VDD.n217 VSS 0.0315f
C1725 VDD.n218 VSS 0.0171f
C1726 VDD.n219 VSS 0.0928f
C1727 VDD.t151 VSS 0.109f
C1728 VDD.n220 VSS 0.076f
C1729 VDD.n221 VSS 0.0401f
C1730 VDD.n222 VSS 0.0444f
C1731 VDD.n223 VSS 0.0343f
C1732 VDD.t5 VSS 0.00907f
C1733 VDD.n224 VSS 0.0496f
C1734 VDD.n225 VSS 0.0313f
C1735 VDD.n226 VSS 0.0498f
C1736 VDD.n227 VSS 0.0418f
C1737 VDD.n228 VSS 0.0366f
C1738 VDD.n229 VSS 0.0457f
C1739 VDD.n230 VSS 0.0291f
C1740 VDD.n231 VSS 0.0401f
C1741 VDD.n232 VSS 0.0423f
C1742 VDD.n233 VSS 0.0327f
C1743 VDD.n234 VSS 0.0484f
C1744 VDD.n235 VSS 0.0448f
C1745 VDD.n236 VSS 0.0327f
C1746 VDD.n237 VSS 0.0484f
C1747 VDD.n238 VSS 0.0448f
C1748 VDD.n239 VSS 0.0327f
C1749 VDD.n240 VSS 0.0473f
C1750 VDD.n241 VSS 0.0794f
C1751 VDD.n242 VSS 0.0496f
C1752 VDD.n243 VSS 0.0521f
C1753 VDD.n244 VSS 0.0292f
C1754 VDD.n245 VSS 0.137f
C1755 VDD.n246 VSS 0.774f
C1756 VDD.n247 VSS 0.665f
C1757 VDD.n248 VSS 0.029f
C1758 VDD.n249 VSS 0.0938f
C1759 VDD.t107 VSS 0.0842f
C1760 VDD.t164 VSS 0.137f
C1761 VDD.n250 VSS 0.0657f
C1762 VDD.n251 VSS 0.0703f
C1763 VDD.t165 VSS 0.0214f
C1764 VDD.t167 VSS 0.00889f
C1765 VDD.n252 VSS 0.029f
C1766 VDD.t166 VSS 0.0793f
C1767 VDD.n253 VSS 0.0938f
C1768 VDD.t86 VSS 0.0842f
C1769 VDD.t89 VSS 0.137f
C1770 VDD.n254 VSS 0.0657f
C1771 VDD.t90 VSS 0.0214f
C1772 VDD.t150 VSS 0.00893f
C1773 VDD.n255 VSS 0.00892f
C1774 VDD.n256 VSS 0.0439f
C1775 VDD.t42 VSS 0.0797f
C1776 VDD.t43 VSS 0.00889f
C1777 VDD.n257 VSS 0.0314f
C1778 VDD.n258 VSS 0.0823f
C1779 VDD.t71 VSS 0.0704f
C1780 VDD.t149 VSS 0.107f
C1781 VDD.n259 VSS 0.0554f
C1782 VDD.n260 VSS 0.0313f
C1783 VDD.n261 VSS 0.279f
C1784 VDD.n262 VSS 0.515f
C1785 VDD.n263 VSS 0.103f
C1786 VDD.n264 VSS 0.31f
C1787 VDD.n265 VSS 0.287f
C1788 CLK.n0 VSS 0.0027f
C1789 CLK.n1 VSS 0.0027f
C1790 CLK.t6 VSS 0.0057f
C1791 CLK.t4 VSS 0.022f
C1792 CLK.n2 VSS 0.0365f
C1793 CLK.n3 VSS 0.00774f
C1794 CLK.n4 VSS 0.00871f
C1795 CLK.n5 VSS 0.00292f
C1796 CLK.t1 VSS 0.0267f
C1797 CLK.t0 VSS 0.0176f
C1798 CLK.n6 VSS 0.0472f
C1799 CLK.n7 VSS 0.00608f
C1800 CLK.n8 VSS 0.00221f
C1801 CLK.n9 VSS 0.0885f
C1802 CLK.n10 VSS 0.0872f
C1803 CLK.n11 VSS 0.00443f
C1804 CLK.t3 VSS 0.0267f
C1805 CLK.t2 VSS 0.0176f
C1806 CLK.n12 VSS 0.0472f
C1807 CLK.n13 VSS 0.00608f
C1808 CLK.n14 VSS 0.00219f
C1809 CLK.n15 VSS 0.0559f
C1810 CLK.n16 VSS 0.0552f
C1811 CLK.n17 VSS 0.00785f
C1812 CLK.n18 VSS 0.0159f
C1813 CLK.n19 VSS 0.0027f
C1814 CLK.t12 VSS 0.0057f
C1815 CLK.t10 VSS 0.022f
C1816 CLK.n20 VSS 0.0365f
C1817 CLK.n21 VSS 0.00774f
C1818 CLK.n22 VSS 0.00871f
C1819 CLK.n23 VSS 0.00292f
C1820 CLK.t16 VSS 0.0267f
C1821 CLK.t25 VSS 0.0176f
C1822 CLK.n24 VSS 0.0472f
C1823 CLK.n25 VSS 0.00608f
C1824 CLK.n26 VSS 0.00221f
C1825 CLK.n27 VSS 0.0885f
C1826 CLK.n28 VSS 0.0872f
C1827 CLK.n29 VSS 0.00443f
C1828 CLK.t21 VSS 0.0267f
C1829 CLK.t20 VSS 0.0176f
C1830 CLK.n30 VSS 0.0472f
C1831 CLK.n31 VSS 0.00608f
C1832 CLK.n32 VSS 0.00219f
C1833 CLK.n33 VSS 0.0559f
C1834 CLK.n34 VSS 0.0552f
C1835 CLK.n35 VSS 0.00785f
C1836 CLK.n36 VSS 0.0159f
C1837 CLK.n37 VSS 0.0027f
C1838 CLK.t7 VSS 0.022f
C1839 CLK.t17 VSS 0.0057f
C1840 CLK.n38 VSS 0.0365f
C1841 CLK.n39 VSS 0.00775f
C1842 CLK.n40 VSS 0.00871f
C1843 CLK.n41 VSS 0.00292f
C1844 CLK.t13 VSS 0.0267f
C1845 CLK.t11 VSS 0.0176f
C1846 CLK.n42 VSS 0.0472f
C1847 CLK.n43 VSS 0.00608f
C1848 CLK.n44 VSS 0.00221f
C1849 CLK.n45 VSS 0.0882f
C1850 CLK.n46 VSS 0.0898f
C1851 CLK.n47 VSS 0.00443f
C1852 CLK.t15 VSS 0.0267f
C1853 CLK.t14 VSS 0.0176f
C1854 CLK.n48 VSS 0.0472f
C1855 CLK.n49 VSS 0.00608f
C1856 CLK.n50 VSS 0.00219f
C1857 CLK.n51 VSS 0.0581f
C1858 CLK.n52 VSS 0.0551f
C1859 CLK.n53 VSS 0.00785f
C1860 CLK.n54 VSS 0.0159f
C1861 CLK.n55 VSS 0.0141f
C1862 CLK.n56 VSS 0.00239f
C1863 CLK.t9 VSS 0.0267f
C1864 CLK.t8 VSS 0.0176f
C1865 CLK.n57 VSS 0.0473f
C1866 CLK.n58 VSS 0.00712f
C1867 CLK.n59 VSS 0.0029f
C1868 CLK.n60 VSS 0.238f
C1869 CLK.n61 VSS 0.372f
C1870 CLK.n62 VSS 2.2f
C1871 CLK.n63 VSS 2.1f
C1872 CLK.n64 VSS 0.00871f
C1873 CLK.n65 VSS 0.00292f
C1874 CLK.t19 VSS 0.0267f
C1875 CLK.t18 VSS 0.0176f
C1876 CLK.n66 VSS 0.0472f
C1877 CLK.n67 VSS 0.00608f
C1878 CLK.n68 VSS 0.00221f
C1879 CLK.n69 VSS 0.0882f
C1880 CLK.n70 VSS 0.0898f
C1881 CLK.n71 VSS 0.00443f
C1882 CLK.t23 VSS 0.0267f
C1883 CLK.t22 VSS 0.0176f
C1884 CLK.n72 VSS 0.0472f
C1885 CLK.n73 VSS 0.00608f
C1886 CLK.n74 VSS 0.00219f
C1887 CLK.n75 VSS 0.0581f
C1888 CLK.n76 VSS 0.0551f
C1889 CLK.t24 VSS 0.022f
C1890 CLK.t5 VSS 0.0057f
C1891 CLK.n77 VSS 0.0365f
C1892 CLK.n78 VSS 0.00775f
C1893 CLK.n79 VSS 0.365f
C1894 CLK.n80 VSS 0.0159f
C1895 CLK.n81 VSS 0.0215f
C1896 CLK.n82 VSS 0.326f
.ends

