magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2088 -2044 2472 2844
<< mvnmos >>
rect 0 0 140 800
rect 244 0 384 800
<< mvndiff >>
rect -88 787 0 800
rect -88 741 -75 787
rect -29 741 0 787
rect -88 683 0 741
rect -88 637 -75 683
rect -29 637 0 683
rect -88 579 0 637
rect -88 533 -75 579
rect -29 533 0 579
rect -88 475 0 533
rect -88 429 -75 475
rect -29 429 0 475
rect -88 371 0 429
rect -88 325 -75 371
rect -29 325 0 371
rect -88 267 0 325
rect -88 221 -75 267
rect -29 221 0 267
rect -88 163 0 221
rect -88 117 -75 163
rect -29 117 0 163
rect -88 59 0 117
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 140 787 244 800
rect 140 741 169 787
rect 215 741 244 787
rect 140 683 244 741
rect 140 637 169 683
rect 215 637 244 683
rect 140 579 244 637
rect 140 533 169 579
rect 215 533 244 579
rect 140 475 244 533
rect 140 429 169 475
rect 215 429 244 475
rect 140 371 244 429
rect 140 325 169 371
rect 215 325 244 371
rect 140 267 244 325
rect 140 221 169 267
rect 215 221 244 267
rect 140 163 244 221
rect 140 117 169 163
rect 215 117 244 163
rect 140 59 244 117
rect 140 13 169 59
rect 215 13 244 59
rect 140 0 244 13
rect 384 787 472 800
rect 384 741 413 787
rect 459 741 472 787
rect 384 683 472 741
rect 384 637 413 683
rect 459 637 472 683
rect 384 579 472 637
rect 384 533 413 579
rect 459 533 472 579
rect 384 475 472 533
rect 384 429 413 475
rect 459 429 472 475
rect 384 371 472 429
rect 384 325 413 371
rect 459 325 472 371
rect 384 267 472 325
rect 384 221 413 267
rect 459 221 472 267
rect 384 163 472 221
rect 384 117 413 163
rect 459 117 472 163
rect 384 59 472 117
rect 384 13 413 59
rect 459 13 472 59
rect 384 0 472 13
<< mvndiffc >>
rect -75 741 -29 787
rect -75 637 -29 683
rect -75 533 -29 579
rect -75 429 -29 475
rect -75 325 -29 371
rect -75 221 -29 267
rect -75 117 -29 163
rect -75 13 -29 59
rect 169 741 215 787
rect 169 637 215 683
rect 169 533 215 579
rect 169 429 215 475
rect 169 325 215 371
rect 169 221 215 267
rect 169 117 215 163
rect 169 13 215 59
rect 413 741 459 787
rect 413 637 459 683
rect 413 533 459 579
rect 413 429 459 475
rect 413 325 459 371
rect 413 221 459 267
rect 413 117 459 163
rect 413 13 459 59
<< polysilicon >>
rect 0 800 140 844
rect 244 800 384 844
rect 0 -44 140 0
rect 244 -44 384 0
<< metal1 >>
rect -75 787 -29 800
rect -75 683 -29 741
rect -75 579 -29 637
rect -75 475 -29 533
rect -75 371 -29 429
rect -75 267 -29 325
rect -75 163 -29 221
rect -75 59 -29 117
rect -75 0 -29 13
rect 169 787 215 800
rect 169 683 215 741
rect 169 579 215 637
rect 169 475 215 533
rect 169 371 215 429
rect 169 267 215 325
rect 169 163 215 221
rect 169 59 215 117
rect 169 0 215 13
rect 413 787 459 800
rect 413 683 459 741
rect 413 579 459 637
rect 413 475 459 533
rect 413 371 459 429
rect 413 267 459 325
rect 413 163 459 221
rect 413 59 459 117
rect 413 0 459 13
<< labels >>
rlabel metal1 192 400 192 400 4 D
rlabel metal1 436 400 436 400 4 S
rlabel metal1 -52 400 -52 400 4 S
<< end >>
