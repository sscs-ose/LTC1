* NGSPICE file created from nand3_mag_flat.ext - technology: gf180mcuC

.subckt pex_nand3_mag_ibr IN3 IN2 IN1 VDD VSS OUT
X0 a_168_24# IN3.t0 VSS.t2 VSS.t1 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1 OUT IN3.t1 VDD.t4 VDD.t3 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2 VDD IN2.t0 OUT.t0 VDD.t0 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X3 OUT IN1.t0 a_328_24# VSS.t3 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X4 OUT IN1.t1 VDD.t6 VDD.t5 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X5 a_328_24# IN2.t1 a_168_24# VSS.t0 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
R0 IN3.n0 IN3.t1 30.9379
R1 IN3.n0 IN3.t0 24.5101
R2 IN3 IN3.n0 4.11094
R3 VSS.t0 VSS.t3 994.264
R4 VSS.n0 VSS.t0 596.558
R5 VSS.n0 VSS.t1 397.707
R6 VSS VSS.t2 6.02876
R7 VSS VSS.n2 2.6038
R8 VSS.n2 VSS.n0 2.6005
R9 VSS.n2 VSS.n1 0.368921
R10 VDD.t0 VDD.t5 303.031
R11 VDD.n3 VDD.t0 193.183
R12 VDD.n3 VDD.t3 109.849
R13 VDD.n5 VDD.t4 5.213
R14 VDD.n5 VDD.n4 3.1505
R15 VDD.n4 VDD.n3 3.1505
R16 VDD VDD.n1 2.96355
R17 VDD.n1 VDD.t6 2.2755
R18 VDD.n1 VDD.n0 2.2755
R19 VDD.n4 VDD.n2 0.109121
R20 VDD VDD.n5 0.00166129
R21 OUT.n4 OUT.n3 5.89611
R22 OUT OUT.n0 5.22702
R23 OUT.n4 OUT.n2 3.63901
R24 OUT.n2 OUT.t0 2.2755
R25 OUT.n2 OUT.n1 2.2755
R26 OUT OUT.n4 0.00152273
R27 IN2.n0 IN2.t1 36.935
R28 IN2.n0 IN2.t0 18.1962
R29 IN2 IN2.n0 4.0877
R30 IN1.n0 IN1.t0 36.935
R31 IN1.n0 IN1.t1 18.1962
R32 IN1 IN1.n0 4.09366
C0 IN3 IN2 0.0466f
C1 VDD IN2 0.171f
C2 IN1 IN3 1.3e-19
C3 VDD IN1 0.137f
C4 a_328_24# OUT 0.0731f
C5 a_328_24# a_168_24# 0.0504f
C6 OUT IN2 0.209f
C7 VDD IN3 0.158f
C8 OUT IN1 0.246f
C9 a_168_24# IN2 8.64e-19
C10 OUT IN3 0.0904f
C11 OUT VDD 0.318f
C12 a_168_24# IN3 8.64e-19
C13 VDD a_168_24# 2.21e-19
C14 a_328_24# IN2 0.00103f
C15 a_328_24# IN1 8.64e-19
C16 IN1 IN2 0.115f
C17 OUT a_168_24# 0.0202f
.ends

