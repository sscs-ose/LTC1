* NGSPICE file created from PLL_TOP_MUX_flat.ext - technology: gf180mcuC

.subckt pex_PLL_TOP_MUX UP_INPUT VDD DN_INPUT VSS PRE_SCALAR UP F_IN DN ITAIL DIV_OUT S1 ITAIL1 VCTRL_IN S6 VCTRL2 S2 OUT
X0 a_42928_8770.t0 a_43228_8148.t0 VDD.t98 ppolyf_u r_width=1.1u r_length=2.6u
X1 RES_74k_1.M.t1 VSS.t131 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X2 PFD_T2_0.INV_mag_1.OUT PFD_T2_0.INV_mag_1.IN.t17 VSS.t579 VSS.t578 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.5u
X3 PFD_T2_0.Buffer_V_2_0.IN PFD_T2_0.INV_mag_1.IN.t18 VDD.t466 VDD.t244 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X4 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t31 VSS.t265 VSS.t264 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X5 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t32 VDD.t161 VDD.t160 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X6 RES_74k_1.M.t1 VSS.t130 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X7 VSS VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t31 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t3 VSS.t764 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X8 VSS VCTRL2.t1 a_25706_n567.t38 VSS.t276 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X9 VSS mux_magic_3.OR_magic_0.A.t3 a_21443_9476.t0 VSS.t250 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X10 a_43528_12082.t0 a_43828_11460.t0 VDD.t4 ppolyf_u r_width=1.1u r_length=2.6u
X11 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t31 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t3 VDD.t162 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X12 VSS PFD_T2_0.Buffer_V_2_0.IN.t11 a_25557_8739.t0 VSS.t436 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X13 VSS.t241 VSS.t239 VSS.t241 VSS.t240 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X14 RES_74k_1.M.t1 VSS.t129 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X15 RES_74k_1.M.t1 VSS.t128 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X16 RES_74k_1.P.t12 RES_74k_1.P.t13 VDD.t79 ppolyf_u r_width=1.1u r_length=2.6u
X17 RES_74k_1.P A_MUX_0.Tr_Gate_1.CLK.t12 VCO_DFF_C_0.VCTRL.t3 VSS.t449 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X18 VDD a_22967_8787.t4 PFD_T2_0.INV_mag_1.IN.t13 VDD.t731 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X19 RES_74k_1.P.t10 RES_74k_1.P.t11 VDD.t98 ppolyf_u r_width=1.1u r_length=2.6u
X20 VSS VCTRL2.t3 a_34443_2598.t38 VSS.t281 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X21 RES_74k_1.M.t1 VSS.t127 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X22 VSS VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t12 VCO_DFF_C_0.VCO_C_0.OUTB.t3 VSS.t699 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X23 VSS S6.t0 mux_magic_3.AND2_magic_0.A.t2 VSS.t253 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X24 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN OUT.t12 VSS.t533 VSS.t519 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X25 VDD a_22967_8787.t5 PFD_T2_0.INV_mag_1.IN.t14 VDD.t734 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X26 a_43828_11254.t0 a_43528_10632.t0 VDD.t4 ppolyf_u r_width=1.1u r_length=2.6u
X27 VSS VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t16 OUT.t0 VSS.t511 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X28 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCTRL.t16 VDD.t776 VDD.t47 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X29 VSS PFD_T2_0.INV_mag_1.OUT.t3 a_22879_10704.t1 VSS.t569 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X30 PFD_T2_0.INV_mag_1.OUT PFD_T2_0.INV_mag_1.IN.t19 VDD.t467 VDD.t462 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X31 VDD.t77 VDD.t75 VDD.t77 VDD.t76 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X32 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t31 VDD.t365 VDD.t364 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X33 VDD.t74 VDD.t73 VDD.t74 VDD.t13 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X34 RES_74k_1.M.t1 VSS.t126 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X35 VSS.t238 VSS.t237 VSS.t238 VSS.t176 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X36 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t12 a_34443_2598.t59 VSS.t439 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X37 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t32 VDD.t611 VDD.t160 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X38 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCTRL.t17 VDD.t784 VDD.t66 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X39 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t33 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t16 VDD.t162 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X40 VDD.t72 VDD.t70 VDD.t72 VDD.t71 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X41 RES_74k_1.M.t1 VSS.t125 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X42 mux_magic_2.OR_magic_0.B a_19897_10547.t6 VDD.t320 VDD.t319 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X43 RES_74k_1.M.t1 VSS.t124 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X44 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t12 a_34443_2598.t40 VSS.t478 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X45 RES_74k_1.M.t1 VSS.t123 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X46 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t34 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t15 VDD.t165 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X47 VSS VCTRL2.t6 a_34443_2598.t36 VSS.t288 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X48 VSS VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t12 a_44716_n517.t1 VSS.t665 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X49 VSS.t236 VSS.t235 VSS.t236 VSS.t228 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X50 VDD mux_magic_1.AND2_magic_0.A.t10 a_27875_8520.t0 VDD.t116 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X51 VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t12 VSS.t592 VSS.t591 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X52 VDD VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t13 VCO_DFF_C_0.VCO_C_0.OUT.t11 VDD.t479 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X53 VSS ITAIL1.t6 ITAIL1.t7 VSS.t618 nfet_03v3 ad=92.8f pd=0.92u as=0.158p ps=1.64u w=0.28u l=0.56u
X54 RES_74k_1.P.t18 RES_74k_1.P.t19 VDD.t106 ppolyf_u r_width=1.1u r_length=2.6u
X55 RES_74k_1.M.t1 VSS.t122 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X56 VSS.t234 VSS.t232 VSS.t234 VSS.t233 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X57 mux_magic_3.AND2_magic_0.A S6.t1 VDD.t133 VDD.t132 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X58 VDD S3.t1 a_27875_9714.t4 VDD.t561 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X59 VSS.t231 VSS.t230 VSS.t231 VSS.t187 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X60 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t32 VDD.t788 VDD.t396 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X61 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCTRL.t18 VDD.t93 VDD.t88 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X62 a_44728_10426.t1 a_44428_9804.t0 VDD.t106 ppolyf_u r_width=1.1u r_length=2.6u
X63 VDD S4.t0 A_MUX_0.Tr_Gate_1.CLK.t0 VDD.t698 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X64 RES_74k_1.M.t1 VSS.t121 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X65 a_42628_9598.t0 a_42928_8976.t1 VDD.t101 ppolyf_u r_width=1.1u r_length=2.6u
X66 VSS.t229 VSS.t227 VSS.t229 VSS.t228 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X67 a_44728_12082.t0 a_44428_11460.t0 VDD.t106 ppolyf_u r_width=1.1u r_length=2.6u
X68 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t33 VSS.t688 VSS.t266 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X69 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.VCO_C_0.OUTB.t12 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t2 VSS.t736 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X70 PFD_T2_0.FIN a_21437_10708.t6 VSS.t259 VSS.t258 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X71 PFD_T2_0.INV_mag_0.OUT PFD_T2_0.INV_mag_0.IN.t18 VDD.t463 VDD.t462 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X72 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.OUT.t13 a_25706_n567.t41 VSS.t658 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X73 VSS S1.t0 mux_magic_2.AND2_magic_0.A.t0 VSS.t457 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X74 a_44428_11254.t1 a_44728_10632.t1 VDD.t106 ppolyf_u r_width=1.1u r_length=2.6u
X75 VSS OUT.t13 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t2 VSS.t511 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X76 VSS VCTRL2.t8 a_25706_n567.t35 VSS.t292 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X77 ITAIL ITAIL.t14 VDD.t144 VDD.t143 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X78 VSS PFD_T2_0.INV_mag_0.IN.t19 a_23836_10693.t2 VSS.t564 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X79 VSS S3.t2 mux_magic_1.AND2_magic_0.A.t4 VSS.t654 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X80 a_45928_10426.t1 a_46228_9804.t0 VDD.t107 ppolyf_u r_width=1.1u r_length=2.6u
X81 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t33 VDD.t790 VDD.t789 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X82 a_44428_9598.t0 a_44128_8976.t0 VDD.t105 ppolyf_u r_width=1.1u r_length=2.6u
X83 VDD S4.t1 a_42763_5679.t5 VDD.t255 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X84 RES_74k_1.M.t1 VSS.t120 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X85 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.VCO_C_0.OUTB.t13 VSS.t738 VSS.t737 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X86 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t13 VDD.t662 VDD.t660 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X87 RES_74k_1.M.t1 VSS.t119 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X88 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t35 VDD.t169 VDD.t168 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X89 a_45928_8770.t0 a_45628_8148.t0 VDD.t100 ppolyf_u r_width=1.1u r_length=2.6u
X90 OUTB a_41879_1284.t6 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t8 VDD.t146 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X91 a_42628_8770.t0 a_42628_8148.t0 VDD.t78 ppolyf_u r_width=1.1u r_length=2.6u
X92 RES_74k_1.M.t1 VSS.t118 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X93 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.OUT.t14 a_25706_n567.t42 VSS.t659 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X94 VSS DIV_OUT.t1 a_20103_8443.t2 VSS.t711 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X95 RES_74k_1.P.t0 RES_74k_1.P.t1 VDD.t3 ppolyf_u r_width=1.1u r_length=2.6u
X96 VSS VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t14 VCO_DFF_C_0.VCO_C_0.OUT.t2 VSS.t593 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X97 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t34 VDD.t791 VDD.t364 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X98 VDD.t69 VDD.t68 VDD.t69 VDD.t37 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X99 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t20 VDD.t447 VDD.t446 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X100 VSS VCTRL2.t9 a_25706_n567.t34 VSS.t292 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X101 RES_74k_1.P.t85 RES_74k_1.P.t86 VDD.t100 ppolyf_u r_width=1.1u r_length=2.6u
X102 VSS OUT.t14 OUTB.t3 VSS.t536 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X103 PFD_T2_0.FDIV a_21443_9476.t6 VDD.t82 VDD.t81 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X104 RES_74k_1.P.t14 RES_74k_1.P.t15 VDD.t78 ppolyf_u r_width=1.1u r_length=2.6u
X105 VDD.t67 VDD.t65 VDD.t67 VDD.t66 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X106 PFD_T2_0.INV_mag_1.IN a_22967_8787.t6 VDD.t737 VDD.t720 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X107 VDD ITAIL.t12 ITAIL.t13 VDD.t136 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X108 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t35 VDD.t792 VDD.t382 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X109 RES_74k_1.M.t1 VSS.t117 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X110 VSS VSS.t220 a_20103_9637.t0 VSS.t221 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X111 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t36 VDD.t794 VDD.t793 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X112 VDD A_MUX_0.Tr_Gate_1.CLK.t13 a_45158_5339.t5 VDD.t252 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X113 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t34 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t5 VDD.t175 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X114 mux_magic_0.OR_magic_0.B a_27722_10564.t6 VSS.t451 VSS.t450 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X115 a_45328_12082.t0 a_45628_11460.t0 VDD.t3 ppolyf_u r_width=1.1u r_length=2.6u
X116 a_44128_8770.t0 a_43828_8148.t0 VDD.t5 ppolyf_u r_width=1.1u r_length=2.6u
X117 mux_magic_1.AND2_magic_0.A S3.t3 VDD.t488 VDD.t487 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X118 VDD.t64 VDD.t62 VDD.t64 VDD.t63 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X119 VDD S2.t2 a_27722_10564.t1 VDD.t329 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X120 RES_74k_1.P ITAIL.t18 a_31732_10267.t6 VDD.t139 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X121 VSS VCTRL2.t10 a_25706_n567.t33 VSS.t297 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X122 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t32 VSS.t522 VSS.t521 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X123 RES_74k_1.M.t1 VSS.t116 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X124 mux_magic_0.OR_magic_0.A a_27722_11758.t6 VSS.t550 VSS.t549 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X125 RES_74k_1.M.t1 VSS.t115 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X126 VDD a_31468_10271.t6 a_31732_10267.t8 VDD.t599 pfet_03v3 ad=0.308p pd=2.28u as=0.308p ps=2.28u w=0.7u l=0.56u
X127 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t36 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t11 VDD.t170 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X128 RES_74k_1.M.t1 VSS.t114 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X129 a_45628_11254.t0 a_45328_10632.t0 VDD.t3 ppolyf_u r_width=1.1u r_length=2.6u
X130 VDD A_MUX_0.Tr_Gate_1.CLK.t14 a_45158_5339.t4 VDD.t722 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X131 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t13 a_34443_2598.t58 VSS.t480 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X132 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.VCO_C_0.OUTB.t15 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t1 VSS.t739 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X133 VDD VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t16 a_41879_1284.t3 VDD.t146 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X134 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t33 VDD.t367 VDD.t366 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X135 VDD OUT.t15 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t11 VDD.t418 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X136 VDD.t61 VDD.t60 VDD.t61 VDD.t13 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X137 VDD a_22966_11778.t4 PFD_T2_0.INV_mag_0.IN.t4 VDD.t305 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X138 RES_74k_1.P.t16 RES_74k_1.P.t17 VDD.t5 ppolyf_u r_width=1.1u r_length=2.6u
X139 VSS VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t34 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t2 VSS.t523 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X140 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t37 VDD.t174 VDD.t173 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X141 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t35 VDD.t615 VDD.t614 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X142 RES_74k_1.M.t2 VSS.t113 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X143 VSS UP.t5 a_31940_9626.t6 VSS.t600 nfet_03v3 ad=92.8f pd=0.92u as=92.8f ps=0.92u w=0.28u l=0.56u
X144 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t37 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t9 VDD.t795 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X145 mux_magic_3.OR_magic_0.A a_19903_8443.t6 VDD.t557 VDD.t556 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X146 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t38 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t13 VDD.t175 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X147 RES_74k_1.M.t1 VSS.t112 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X148 RES_74k_1.M.t1 VSS.t111 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X149 VDD VCO_DFF_C_0.VCO_C_0.OUTB.t16 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t11 VDD.t688 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X150 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t38 VSS.t768 VSS.t767 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X151 VDD a_31468_10271.t7 a_31732_10267.t9 VDD.t599 pfet_03v3 ad=0.308p pd=2.28u as=0.308p ps=2.28u w=0.7u l=0.56u
X152 VDD VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t21 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t5 VDD.t448 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X153 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t14 VSS.t426 VSS.t425 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X154 RES_74k_1.M.t3 VSS.t110 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X155 VDD mux_magic_2.OR_magic_0.A.t3 a_21437_12116.t7 VDD.t549 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X156 RES_74k_1.M.t1 VSS.t109 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X157 VDD VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t17 OUT.t1 VDD.t347 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X158 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.VCO_C_0.OUTB.t17 VDD.t745 VDD.t679 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X159 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t15 VCO_DFF_C_0.VCO_C_0.OUTB.t10 VDD.t216 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X160 RES_74k_1.M.t1 VSS.t108 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X161 VSS VCTRL2.t12 a_25706_n567.t32 VSS.t276 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X162 VDD.t59 VDD.t57 VDD.t59 VDD.t58 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X163 RES_74k_1.P.t2 RES_74k_1.P.t3 VDD.t78 ppolyf_u r_width=1.1u r_length=2.6u
X164 VSS VCTRL2.t13 a_25706_n567.t31 VSS.t276 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X165 RES_74k_1.P.t99 RES_74k_1.P.t100 VDD.t79 ppolyf_u r_width=1.1u r_length=2.6u
X166 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t35 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t1 VDD.t368 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X167 UP a_29262_10725.t6 VDD.t214 VDD.t213 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X168 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t36 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t6 VDD.t187 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X169 mux_magic_2.OR_magic_0.A a_19897_11741.t6 VSS.t695 VSS.t694 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X170 VSS a_22967_8787.t7 a_22881_9554.t1 VSS.t733 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X171 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t39 VDD.t798 VDD.t396 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X172 RES_74k_1.M.t1 VSS.t107 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X173 VDD a_25557_8739.t3 PFD_T2_0.DOWN.t2 VDD.t667 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X174 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t37 VDD.t619 VDD.t618 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X175 RES_74k_1.M.t0 a_42628_11460.t1 VDD.t78 ppolyf_u r_width=1.1u r_length=2.6u
X176 VDD OUT.t16 OUTB.t11 VDD.t350 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X177 mux_magic_0.AND2_magic_0.A S2.t3 VDD.t333 VDD.t332 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X178 a_46528_12082.t1 a_46228_11460.t1 VDD.t79 ppolyf_u r_width=1.1u r_length=2.6u
X179 VSS.t219 VSS.t218 VSS.t219 VSS.t139 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X180 PFD_T2_0.INV_mag_0.IN a_22966_11778.t6 VDD.t309 VDD.t308 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X181 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t16 VDD.t678 VDD.t677 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X182 a_45328_10426.t1 a_45628_9804.t1 VDD.t3 ppolyf_u r_width=1.1u r_length=2.6u
X183 VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t15 VDD.t486 VDD.t482 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X184 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t36 VDD.t371 VDD.t364 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X185 RES_74k_1.P.t97 RES_74k_1.P.t98 VDD.t108 ppolyf_u r_width=1.1u r_length=2.6u
X186 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.INV_mag_0.IN.t20 VDD.t786 VDD.t308 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X187 VDD a_22967_8787.t8 PFD_T2_0.INV_mag_1.IN.t16 VDD.t724 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X188 DN a_29415_9553.t6 VDD.t8 VDD.t7 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X189 a_43828_9598.t0 a_43528_8976.t1 VDD.t4 ppolyf_u r_width=1.1u r_length=2.6u
X190 VCO_DFF_C_0.VCTRL S4.t3 VCTRL_IN.t3 VSS.t714 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X191 VCTRL_IN a_42763_5679.t6 VCO_DFF_C_0.VCTRL.t4 VDD.t255 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X192 VSS VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t37 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t1 VSS.t526 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X193 RES_74k_1.M.t1 VSS.t106 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X194 mux_magic_2.AND2_magic_0.A S1.t2 VDD.t270 VDD.t269 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X195 a_42628_11254.t0 a_42628_10426.t1 VDD.t78 ppolyf_u r_width=1.1u r_length=2.6u
X196 a_46228_11254.t0 a_46528_10632.t0 VDD.t79 ppolyf_u r_width=1.1u r_length=2.6u
X197 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t38 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t3 VDD.t372 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X198 RES_74k_1.M.t1 VSS.t105 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X199 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t14 a_34443_2598.t42 VSS.t480 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X200 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t39 VDD.t376 VDD.t375 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X201 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t18 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t8 VSS.t670 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X202 PFD_T2_0.Buffer_V_2_0.IN PFD_T2_0.INV_mag_0.OUT.t6 VSS.t488 VSS.t487 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X203 VDD DIV_OUT.t2 a_19903_8443.t5 VDD.t693 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X204 VDD mux_magic_1.OR_magic_0.A.t3 a_29415_8145.t4 VDD.t285 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X205 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t39 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t12 VDD.t165 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X206 VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t16 VDD.t490 VDD.t489 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X207 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t40 VSS.t267 VSS.t266 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X208 RES_74k_1.M.t1 VSS.t104 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X209 RES_74k_1.M.t1 VSS.t103 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X210 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.OUTB.t18 a_25706_n567.t51 VSS.t659 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X211 mux_magic_0.OR_magic_0.A a_27722_11758.t7 VDD.t535 VDD.t534 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X212 RES_74k_1.P.t44 RES_74k_1.P.t45 VDD.t80 ppolyf_u r_width=1.1u r_length=2.6u
X213 VSS.t217 VSS.t215 VSS.t217 VSS.t216 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X214 RES_74k_1.M.t1 VSS.t102 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X215 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t40 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t10 VDD.t377 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X216 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT a_44716_n517.t6 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t12 VDD.t564 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X217 VSS ITAIL1.t4 ITAIL1.t5 VSS.t615 nfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X218 a_45028_9598.t0 a_45328_8976.t1 VDD.t103 ppolyf_u r_width=1.1u r_length=2.6u
X219 VSS VCTRL2.t16 a_34443_2598.t33 VSS.t309 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X220 RES_74k_1.P.t79 RES_74k_1.P.t80 VDD.t104 ppolyf_u r_width=1.1u r_length=2.6u
X221 RES_74k_1.P a_45158_5339.t6 VCO_DFF_C_0.VCTRL.t12 VDD.t252 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X222 VSS VCTRL2.t18 a_34443_2598.t32 VSS.t281 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X223 VDD F_IN.t1 a_19897_10547.t4 VDD.t589 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X224 RES_74k_1.P ITAIL.t19 a_31732_10267.t5 VDD.t143 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X225 VDD PFD_T2_0.FDIV.t4 a_22967_8787.t3 VDD.t724 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X226 a_46528_8770.t1 RES_74k_1.P.t72 VDD.t102 ppolyf_u r_width=1.1u r_length=2.6u
X227 mux_magic_0.AND2_magic_0.A S2.t4 VDD.t335 VDD.t334 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X228 a_43528_8770.t0 a_43228_8148.t1 VDD.t104 ppolyf_u r_width=1.1u r_length=2.6u
X229 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t38 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t7 VDD.t165 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X230 VDD S4.t4 A_MUX_0.Tr_Gate_1.CLK.t1 VDD.t698 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X231 VDD VCO_DFF_C_0.VCO_C_0.OUTB.t19 a_44716_1837.t5 VDD.t566 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X232 VDD.t56 VDD.t55 VDD.t56 VDD.t28 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X233 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.INV_mag_1.OUT.t5 VSS.t573 VSS.t572 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X234 a_43528_12082.t1 a_43228_11460.t1 VDD.t104 ppolyf_u r_width=1.1u r_length=2.6u
X235 RES_74k_1.P a_45158_5339.t7 VCO_DFF_C_0.VCTRL.t13 VDD.t722 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X236 VSS.t214 VSS.t212 VSS.t214 VSS.t213 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X237 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t15 a_34443_2598.t43 VSS.t481 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X238 RES_74k_1.P.t60 RES_74k_1.P.t61 VDD.t102 ppolyf_u r_width=1.1u r_length=2.6u
X239 VSS VCTRL2.t21 a_34443_2598.t30 VSS.t281 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X240 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t40 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t11 VDD.t368 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X241 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.INV_mag_0.IN.t21 a_23836_10693.t4 VSS.t561 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X242 ITAIL1 ITAIL1.t2 VSS.t614 VSS.t613 nfet_03v3 ad=0.158p pd=1.64u as=92.8f ps=0.92u w=0.28u l=0.56u
X243 mux_magic_1.AND2_magic_0.A S3.t4 VDD.t497 VDD.t303 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X244 RES_74k_1.P.t62 RES_74k_1.P.t63 VDD.t104 ppolyf_u r_width=1.1u r_length=2.6u
X245 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN a_41879_n196.t6 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t16 VDD.t148 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X246 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t41 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t10 VDD.t398 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X247 VDD mux_magic_3.OR_magic_0.A.t5 a_21443_8068.t2 VDD.t9 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X248 RES_74k_1.P A_MUX_0.Tr_Gate_1.CLK.t16 VCO_DFF_C_0.VCTRL.t2 VSS.t249 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X249 RES_74k_1.M.t1 VSS.t101 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X250 VSS.t211 VSS.t210 VSS.t211 VSS.t133 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X251 VSS S4.t5 A_MUX_0.Tr_Gate_1.CLK.t2 VSS.t715 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X252 mux_magic_2.AND2_magic_0.A S1.t3 VDD.t272 VDD.t271 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X253 a_43228_11254.t0 a_43528_10632.t1 VDD.t104 ppolyf_u r_width=1.1u r_length=2.6u
X254 RES_74k_1.M.t1 VSS.t100 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X255 VSS PFD_T2_0.INV_mag_1.IN.t22 a_23837_9553.t2 VSS.t260 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X256 a_44728_8770.t0 a_45028_8148.t0 VDD.t99 ppolyf_u r_width=1.1u r_length=2.6u
X257 VDD VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t20 a_44716_n517.t3 VDD.t565 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X258 RES_74k_1.M.t1 VSS.t99 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X259 VSS.t209 VSS.t208 VSS.t209 VSS.t136 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X260 VDD S4.t6 A_MUX_0.Tr_Gate_1.CLK.t3 VDD.t706 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X261 RES_74k_1.M.t1 VSS.t98 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X262 VDD mux_magic_2.AND2_magic_0.A.t11 a_19897_11741.t0 VDD.t670 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X263 VCO_DFF_C_0.VCTRL a_42763_5679.t7 VCTRL_IN.t6 VDD.t256 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X264 VDD.t54 VDD.t52 VDD.t54 VDD.t53 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X265 VDD VCO_DFF_C_0.VCTRL.t19 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t29 VDD.t66 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X266 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t42 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t9 VDD.t368 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X267 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VCO_DFF_C_0.VCO_C_0.OUTB.t20 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t3 VSS.t740 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X268 VDD mux_magic_0.OR_magic_0.A.t5 a_29262_12133.t1 VDD.t264 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X269 RES_74k_1.P.t73 RES_74k_1.P.t74 VDD.t99 ppolyf_u r_width=1.1u r_length=2.6u
X270 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t41 VDD.t381 VDD.t380 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X271 RES_74k_1.M.t1 VSS.t97 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X272 VSS PFD_T2_0.DOWN.t4 a_28075_8520.t0 VSS.t420 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X273 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN a_44716_n517.t7 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t5 VDD.t565 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X274 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t16 a_34443_2598.t44 VSS.t482 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X275 VSS VCTRL2.t22 a_25706_n567.t27 VSS.t320 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X276 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t42 VDD.t383 VDD.t382 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X277 VDD.t51 VDD.t49 VDD.t51 VDD.t50 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X278 RES_74k_1.M.t1 VSS.t96 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X279 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.OUTB.t21 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t5 VSS.t741 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X280 RES_74k_1.P.t56 RES_74k_1.P.t57 VDD.t105 ppolyf_u r_width=1.1u r_length=2.6u
X281 VSS VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t39 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t2 VSS.t268 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X282 mux_magic_3.AND2_magic_0.A S6.t3 VSS.t257 VSS.t256 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X283 RES_74k_1.M.t1 VSS.t95 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X284 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.OUT.t15 a_25706_n567.t43 VSS.t659 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X285 ITAIL ITAIL.t10 VDD.t140 VDD.t139 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X286 VSS DN_INPUT.t2 a_28075_9714.t2 VSS.t644 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X287 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t43 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t8 VDD.t377 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X288 VSS VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t21 a_41879_1284.t0 VSS.t671 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X289 PFD_T2_0.INV_mag_0.IN a_22966_11778.t7 VDD.t310 VDD.t223 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X290 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t40 VDD.t622 VDD.t193 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X291 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t43 VDD.t805 VDD.t793 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X292 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t44 VSS.t530 VSS.t529 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X293 PFD_T2_0.INV_mag_0.IN a_22966_11778.t8 VDD.t311 VDD.t225 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X294 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.INV_mag_0.IN.t22 VDD.t224 VDD.t223 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X295 RES_74k_1.M.t1 VSS.t94 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X296 RES_74k_1.M.t1 VSS.t93 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X297 RES_74k_1.M.t1 VSS.t92 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X298 ITAIL1 ITAIL1.t0 VSS.t612 VSS.t611 nfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X299 VSS VCTRL2.t24 a_34443_2598.t28 VSS.t325 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X300 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t16 VDD.t220 VDD.t219 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X301 a_44128_12082.t0 a_44428_11460.t1 VDD.t105 ppolyf_u r_width=1.1u r_length=2.6u
X302 RES_74k_1.P.t109 VSS.t431 cap_mim_2f0_m4m5_noshield c_width=30u c_length=30u
X303 VDD VCO_DFF_C_0.VCTRL.t20 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t27 VDD.t47 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X304 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.INV_mag_0.IN.t23 VDD.t226 VDD.t225 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X305 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.OUTB.t23 a_25706_n567.t52 VSS.t659 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X306 VSS.t207 VSS.t206 VSS.t207 VSS.t195 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X307 RES_74k_1.M.t1 VSS.t91 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X308 VSS VCO_DFF_C_0.VCO_C_0.OUTB.t24 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t2 VSS.t743 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X309 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t44 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t8 VDD.t372 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X310 VSS S2.t5 mux_magic_0.AND2_magic_0.A.t2 VSS.t502 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X311 mux_magic_1.OR_magic_0.A a_27875_8520.t6 VDD.t325 VDD.t324 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X312 RES_74k_1.M.t1 VSS.t90 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X313 RES_74k_1.M.t1 VSS.t89 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X314 VSS mux_magic_2.OR_magic_0.A.t4 a_21437_10708.t5 VSS.t647 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X315 VSS.t205 VSS.t203 VSS.t205 VSS.t204 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X316 RES_74k_1.M.t1 VSS.t88 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X317 VDD VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t22 a_44716_n517.t2 VDD.t566 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X318 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN a_41879_1284.t7 OUTB.t18 VDD.t147 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X319 PFD_T2_0.UP a_25556_11637.t3 VDD.t514 VDD.t513 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X320 a_44428_11254.t0 a_44128_10632.t1 VDD.t105 ppolyf_u r_width=1.1u r_length=2.6u
X321 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCTRL.t21 VDD.t767 VDD.t85 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.84u
X322 mux_magic_1.OR_magic_0.B a_27875_9714.t6 VDD.t666 VDD.t665 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X323 a_46528_10426.t0 a_46228_9804.t1 VDD.t79 ppolyf_u r_width=1.1u r_length=2.6u
X324 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t45 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t7 VDD.t389 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X325 a_42928_10426.t0 a_43228_9804.t0 VDD.t98 ppolyf_u r_width=1.1u r_length=2.6u
X326 VSS OUT.t17 OUTB.t2 VSS.t539 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X327 VDD.t48 VDD.t46 VDD.t48 VDD.t47 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X328 a_44428_9598.t1 a_44728_8976.t0 VDD.t106 ppolyf_u r_width=1.1u r_length=2.6u
X329 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT a_41879_n196.t7 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t13 VDD.t149 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X330 PFD_T2_0.DOWN a_25557_8739.t4 VDD.t664 VDD.t663 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X331 RES_74k_1.M.t1 VSS.t87 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X332 RES_74k_1.M.t1 VSS.t86 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X333 VDD VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t22 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t6 VDD.t451 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X334 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t41 VDD.t623 VDD.t168 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X335 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t46 VDD.t810 VDD.t375 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X336 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t17 VSS.t703 VSS.t551 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X337 VSS VCTRL2.t27 a_25706_n567.t25 VSS.t297 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X338 a_42928_8770.t1 a_42628_8148.t1 VDD.t101 ppolyf_u r_width=1.1u r_length=2.6u
X339 RES_74k_1.M.t1 VSS.t85 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X340 VSS F_IN.t2 a_20097_10547.t2 VSS.t680 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X341 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t47 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t7 VDD.t811 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X342 VDD VCO_DFF_C_0.VCTRL.t22 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t28 VDD.t88 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X343 VDD ITAIL.t8 ITAIL.t9 VDD.t136 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X344 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t45 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t7 VDD.t386 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X345 RES_74k_1.P.t48 RES_74k_1.P.t49 VDD.t103 ppolyf_u r_width=1.1u r_length=2.6u
X346 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t15 a_34443_2598.t56 VSS.t482 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X347 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t41 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t9 VDD.t180 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X348 RES_74k_1.M.t1 VSS.t84 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X349 mux_magic_2.OR_magic_0.A a_19897_11741.t7 VDD.t653 VDD.t652 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X350 RES_74k_1.M.t4 VSS.t83 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X351 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT a_44716_1837.t6 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t12 VDD.t566 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X352 VDD mux_magic_0.AND2_magic_0.A.t11 a_27722_11758.t3 VDD.t259 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X353 RES_74k_1.P.t28 RES_74k_1.P.t29 VDD.t101 ppolyf_u r_width=1.1u r_length=2.6u
X354 RES_74k_1.P.t110 VSS.t432 cap_mim_2f0_m4m5_noshield c_width=30u c_length=30u
X355 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.INV_mag_0.IN.t24 a_23836_10693.t3 VSS.t564 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X356 a_46228_9598.t1 a_45928_8976.t1 VDD.t107 ppolyf_u r_width=1.1u r_length=2.6u
X357 RES_74k_1.M.t1 VSS.t82 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X358 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t42 VDD.t184 VDD.t183 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X359 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t42 VDD.t624 VDD.t618 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X360 VSS.t202 VSS.t201 VSS.t202 VSS.t139 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X361 VSS.t200 VSS.t199 VSS.t200 VSS.t133 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X362 RES_74k_1.M.t1 VSS.t81 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X363 VDD OUT.t18 OUTB.t10 VDD.t347 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X364 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t17 VCO_DFF_C_0.VCO_C_0.OUTB.t8 VDD.t657 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X365 PFD_T2_0.Buffer_V_2_0.IN PFD_T2_0.INV_mag_1.IN.t23 a_23837_9553.t4 VSS.t263 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X366 VSS.t198 VSS.t197 VSS.t198 VSS.t179 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X367 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN OUT.t19 VDD.t426 VDD.t425 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X368 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t48 VDD.t814 VDD.t382 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X369 VDD S1.t4 mux_magic_2.AND2_magic_0.A.t3 VDD.t273 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X370 a_45328_12082.t1 a_45028_11460.t0 VDD.t103 ppolyf_u r_width=1.1u r_length=2.6u
X371 a_44128_8770.t1 a_44428_8148.t0 VDD.t105 ppolyf_u r_width=1.1u r_length=2.6u
X372 mux_magic_1.AND2_magic_0.A S3.t6 VSS.t475 VSS.t474 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X373 RES_74k_1.M.t1 VSS.t80 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X374 VSS.t196 VSS.t194 VSS.t196 VSS.t195 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X375 RES_74k_1.M.t5 VSS.t79 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X376 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN OUT.t20 VDD.t428 VDD.t427 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X377 VDD OUT.t21 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t8 VDD.t429 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X378 VDD VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t18 OUT.t2 VDD.t350 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X379 VSS VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t49 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t1 VSS.t769 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X380 mux_magic_3.OR_magic_0.B a_19903_9637.t6 VDD.t499 VDD.t498 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X381 OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t19 VDD.t354 VDD.t353 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X382 PFD_T2_0.FIN a_21437_10708.t7 VDD.t151 VDD.t150 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X383 VDD.t45 VDD.t43 VDD.t45 VDD.t44 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X384 VDD VCO_DFF_C_0.VCTRL.t23 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t26 VDD.t85 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X385 a_45028_11254.t0 a_45328_10632.t1 VDD.t103 ppolyf_u r_width=1.1u r_length=2.6u
X386 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t43 VDD.t186 VDD.t185 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X387 VDD VCO_DFF_C_0.VCO_C_0.OUTB.t27 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t9 VDD.t682 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X388 RES_74k_1.M.t1 VSS.t78 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X389 VSS.t193 VSS.t191 VSS.t193 VSS.t192 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X390 RES_74k_1.P.t30 RES_74k_1.P.t31 VDD.t105 ppolyf_u r_width=1.1u r_length=2.6u
X391 VSS.t190 VSS.t189 VSS.t190 VSS.t133 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X392 RES_74k_1.P.t111 VSS.t433 cap_mim_2f0_m4m5_noshield c_width=30u c_length=30u
X393 RES_74k_1.M.t1 VSS.t77 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X394 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t23 OUTB.t15 VSS.t674 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X395 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t46 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t6 VDD.t389 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X396 VSS A_MUX_0.Tr_Gate_1.CLK.t18 a_45158_5339.t0 VSS.t449 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X397 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t16 a_34443_2598.t55 VSS.t439 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X398 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.VCO_C_0.OUTB.t28 VDD.t751 VDD.t677 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X399 VDD a_22967_8787.t9 PFD_T2_0.INV_mag_1.IN.t4 VDD.t120 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X400 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t23 VDD.t455 VDD.t454 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X401 DN a_29415_9553.t7 VDD.t417 VDD.t7 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X402 RES_74k_1.M.t1 VSS.t76 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X403 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t47 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t7 VDD.t372 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X404 VSS VCTRL2.t32 a_34443_2598.t24 VSS.t309 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X405 VDD a_19903_8443.t7 mux_magic_3.OR_magic_0.A.t1 VDD.t558 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X406 mux_magic_3.AND2_magic_0.A S6.t4 VDD.t229 VDD.t228 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X407 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t43 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t8 VDD.t625 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X408 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t18 VDD.t680 VDD.t679 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X409 VDD a_19897_10547.t7 mux_magic_2.OR_magic_0.B.t1 VDD.t321 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X410 OUTB OUT.t22 VDD.t432 VDD.t355 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X411 VDD UP_INPUT.t1 a_27722_10564.t4 VDD.t508 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X412 RES_74k_1.M.t1 VSS.t75 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X413 RES_74k_1.M.t1 VSS.t74 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X414 VDD a_22967_8787.t10 PFD_T2_0.INV_mag_1.IN.t5 VDD.t123 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X415 PFD_T2_0.INV_mag_0.IN a_22966_11778.t9 VDD.t313 VDD.t312 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X416 RES_74k_1.P.t40 RES_74k_1.P.t41 VDD.t108 ppolyf_u r_width=1.1u r_length=2.6u
X417 RES_74k_1.P.t42 RES_74k_1.P.t43 VDD.t107 ppolyf_u r_width=1.1u r_length=2.6u
X418 OUTB OUT.t23 VDD.t433 VDD.t353 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X419 VSS.t188 VSS.t186 VSS.t188 VSS.t187 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X420 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t48 VDD.t394 VDD.t375 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X421 VSS VCTRL2.t33 a_25706_n567.t22 VSS.t320 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X422 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t44 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t10 VDD.t187 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X423 VSS VCTRL2.t34 a_34443_2598.t23 VSS.t342 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X424 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCTRL.t24 VDD.t783 VDD.t88 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X425 VSS.t185 VSS.t183 VSS.t185 VSS.t184 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X426 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t24 VSS.t552 VSS.t551 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X427 RES_74k_1.P.t24 RES_74k_1.P.t25 VDD.t108 ppolyf_u r_width=1.1u r_length=2.6u
X428 VCTRL_IN S4.t8 VCO_DFF_C_0.VCTRL.t9 VSS.t720 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X429 VDD.t42 VDD.t41 VDD.t42 VDD.t37 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X430 VSS.t182 VSS.t181 VSS.t182 VSS.t136 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X431 VSS PFD_T2_0.INV_mag_0.OUT.t8 PFD_T2_0.Buffer_V_2_0.IN.t9 VSS.t490 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X432 a_45928_12082.t0 a_46228_11460.t0 VDD.t107 ppolyf_u r_width=1.1u r_length=2.6u
X433 VSS.t180 VSS.t178 VSS.t180 VSS.t179 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X434 VSS VCTRL2.t35 a_34443_2598.t22 VSS.t345 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X435 VDD VSS.t775 a_19903_9637.t1 VDD.t109 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X436 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.VCO_C_0.OUTB.t29 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t3 VSS.t746 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X437 VSS VCTRL2.t36 a_25706_n567.t21 VSS.t297 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X438 VDD PFD_T2_0.INV_mag_1.IN.t24 PFD_T2_0.Buffer_V_2_0.IN.t3 VDD.t120 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X439 a_45928_10426.t0 a_45628_9804.t0 VDD.t100 ppolyf_u r_width=1.1u r_length=2.6u
X440 RES_74k_1.M.t1 VSS.t73 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X441 VSS.t177 VSS.t175 VSS.t177 VSS.t176 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X442 a_42628_10426.t0 a_42628_9804.t0 VDD.t78 ppolyf_u r_width=1.1u r_length=2.6u
X443 VSS VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t45 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t1 VSS.t268 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X444 RES_74k_1.M.t1 VSS.t72 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X445 RES_74k_1.M.t1 VSS.t71 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X446 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT a_44716_1837.t7 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t17 VDD.t567 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X447 mux_magic_0.AND2_magic_0.A S2.t7 VDD.t338 VDD.t332 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X448 VSS VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t19 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t6 VSS.t553 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X449 VSS mux_magic_0.OR_magic_0.A.t6 a_29262_10725.t0 VSS.t454 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X450 OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t20 VSS.t515 VSS.t514 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X451 PFD_T2_0.DOWN a_25557_8739.t5 VSS.t430 VSS.t429 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X452 RES_74k_1.P.t46 RES_74k_1.P.t47 VDD.t108 ppolyf_u r_width=1.1u r_length=2.6u
X453 a_46228_11254.t1 a_45928_10632.t0 VDD.t107 ppolyf_u r_width=1.1u r_length=2.6u
X454 RES_74k_1.M.t1 VSS.t70 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X455 RES_74k_1.M.t1 VSS.t69 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X456 VSS.t174 VSS.t173 VSS.t174 VSS.t136 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X457 VSS.t172 VSS.t171 VSS.t172 VSS.t167 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X458 VDD a_31468_10271.t8 a_31732_10267.t10 VDD.t599 pfet_03v3 ad=0.308p pd=2.28u as=0.308p ps=2.28u w=0.7u l=0.56u
X459 VDD PFD_T2_0.INV_mag_1.IN.t25 PFD_T2_0.Buffer_V_2_0.IN.t2 VDD.t123 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X460 VSS.t170 VSS.t169 VSS.t170 VSS.t142 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X461 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.OUTB.t30 a_25706_n567.t54 VSS.t658 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X462 VDD PFD_T2_0.INV_mag_0.IN.t25 a_24437_9224.t2 VDD.t740 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X463 VSS.t168 VSS.t166 VSS.t168 VSS.t167 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X464 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t49 VDD.t395 VDD.t366 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X465 VDD S4.t9 A_MUX_0.Tr_Gate_1.CLK.t4 VDD.t706 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X466 VDD S6.t6 mux_magic_3.AND2_magic_0.A.t6 VDD.t230 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X467 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t50 VDD.t397 VDD.t396 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X468 VDD PFD_T2_0.INV_mag_1.IN.t26 PFD_T2_0.INV_mag_1.OUT.t1 VDD.t157 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X469 RES_74k_1.M.t1 VSS.t68 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X470 RES_74k_1.M.t6 VSS.t67 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X471 mux_magic_1.AND2_magic_0.A S3.t7 VDD.t304 VDD.t303 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X472 RES_74k_1.M.t1 VSS.t66 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X473 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCTRL.t25 VDD.t119 VDD.t85 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X474 VDD a_27722_10564.t7 mux_magic_0.OR_magic_0.B.t2 VDD.t0 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X475 RES_74k_1.P ITAIL.t22 a_31732_10267.t3 VDD.t143 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X476 RES_74k_1.M.t1 VSS.t65 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X477 PFD_T2_0.INV_mag_1.IN a_22967_8787.t11 VDD.t127 VDD.t126 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X478 a_44128_10426.t0 a_43828_9804.t0 VDD.t5 ppolyf_u r_width=1.1u r_length=2.6u
X479 a_45628_9598.t0 a_45328_8976.t0 VDD.t3 ppolyf_u r_width=1.1u r_length=2.6u
X480 RES_74k_1.P.t64 RES_74k_1.P.t65 VDD.t108 ppolyf_u r_width=1.1u r_length=2.6u
X481 RES_74k_1.M.t1 VSS.t64 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X482 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.OUT.t18 a_25706_n567.t46 VSS.t658 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X483 VCO_DFF_C_0.VCTRL a_45158_5339.t8 RES_74k_1.P.t105 VDD.t248 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X484 RES_74k_1.M.t1 VSS.t63 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X485 PFD_T2_0.UP a_25556_11637.t4 VSS.t631 VSS.t623 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X486 PFD_T2_0.INV_mag_1.IN a_22967_8787.t12 VDD.t129 VDD.t128 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X487 RES_74k_1.P.t66 RES_74k_1.P.t67 VDD.t98 ppolyf_u r_width=1.1u r_length=2.6u
X488 RES_74k_1.P.t68 RES_74k_1.P.t69 VDD.t80 ppolyf_u r_width=1.1u r_length=2.6u
X489 VSS S4.t10 A_MUX_0.Tr_Gate_1.CLK.t5 VSS.t715 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X490 a_43528_8770.t1 a_43828_8148.t1 VDD.t4 ppolyf_u r_width=1.1u r_length=2.6u
X491 VSS VCTRL2.t39 a_34443_2598.t20 VSS.t325 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X492 RES_74k_1.M.t1 VSS.t62 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X493 VDD a_31468_10271.t9 a_31732_10267.t11 VDD.t599 pfet_03v3 ad=0.308p pd=2.28u as=0.308p ps=2.28u w=0.7u l=0.56u
X494 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t44 VDD.t628 VDD.t160 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X495 PFD_T2_0.INV_mag_0.IN a_22966_11778.t10 VDD.t315 VDD.t314 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X496 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t51 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t10 VDD.t398 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X497 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t46 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t9 VDD.t162 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X498 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t20 VDD.t681 VDD.t677 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X499 mux_magic_0.AND2_magic_0.A S2.t8 VDD.t339 VDD.t334 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X500 a_42928_12082.t1 a_43228_11460.t0 VDD.t98 ppolyf_u r_width=1.1u r_length=2.6u
X501 VDD VCO_DFF_C_0.VCTRL.t26 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t2 VDD.t66 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.84u
X502 RES_74k_1.M.t1 VSS.t61 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X503 VSS UP.t6 a_31940_9626.t5 VSS.t600 nfet_03v3 ad=0.158p pd=1.64u as=92.8f ps=0.92u w=0.28u l=0.56u
X504 RES_74k_1.P.t4 RES_74k_1.P.t5 VDD.t80 ppolyf_u r_width=1.1u r_length=2.6u
X505 RES_74k_1.P.t6 RES_74k_1.P.t7 VDD.t4 ppolyf_u r_width=1.1u r_length=2.6u
X506 RES_74k_1.M.t1 VSS.t60 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X507 RES_74k_1.P.t8 RES_74k_1.P.t9 VDD.t80 ppolyf_u r_width=1.1u r_length=2.6u
X508 A_MUX_0.Tr_Gate_1.CLK S4.t11 VDD.t712 VDD.t711 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X509 RES_74k_1.M.t1 VSS.t59 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X510 RES_74k_1.M.t2 VSS.t58 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X511 RES_74k_1.M.t1 VSS.t57 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X512 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t45 VDD.t629 VDD.t168 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X513 VSS VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t46 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t1 VSS.t271 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X514 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN OUT.t24 VSS.t542 VSS.t514 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X515 a_43228_11254.t1 a_42928_10632.t0 VDD.t98 ppolyf_u r_width=1.1u r_length=2.6u
X516 RES_74k_1.P.t101 RES_74k_1.P.t102 VDD.t80 ppolyf_u r_width=1.1u r_length=2.6u
X517 a_45328_8770.t1 a_45028_8148.t1 VDD.t103 ppolyf_u r_width=1.1u r_length=2.6u
X518 VSS VCTRL2.t43 a_34443_2598.t18 VSS.t358 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X519 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t21 VSS.t706 VSS.t556 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X520 VSS VCTRL2.t44 a_25706_n567.t17 VSS.t297 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X521 PFD_T2_0.Buffer_V_2_0.IN PFD_T2_0.INV_mag_1.IN.t28 VDD.t474 VDD.t128 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X522 A_MUX_0.Tr_Gate_1.CLK S4.t12 VDD.t714 VDD.t713 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X523 RES_74k_1.M.t3 VSS.t56 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X524 mux_magic_2.AND2_magic_0.A S1.t5 VDD.t276 VDD.t271 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X525 UP a_29262_10725.t7 VSS.t424 VSS.t423 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X526 RES_74k_1.P.t20 RES_74k_1.P.t21 VDD.t103 ppolyf_u r_width=1.1u r_length=2.6u
X527 RES_74k_1.M.t1 VSS.t55 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X528 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t50 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t6 VDD.t811 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X529 RES_74k_1.M.t5 VSS.t54 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X530 VSS VCO_DFF_C_0.VCO_C_0.OUTB.t33 a_41879_n196.t0 VSS.t741 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X531 VSS VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t25 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t9 VSS.t553 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X532 VSS VCO_DFF_C_0.VCO_C_0.OUTB.t34 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t1 VSS.t750 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X533 VDD S3.t8 mux_magic_1.AND2_magic_0.A.t5 VDD.t570 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X534 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t47 VDD.t192 VDD.t168 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X535 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCTRL.t27 VDD.t778 VDD.t85 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X536 RES_74k_1.P.t22 RES_74k_1.P.t23 VDD.t5 ppolyf_u r_width=1.1u r_length=2.6u
X537 VSS.t165 VSS.t164 VSS.t165 VSS.t139 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X538 VSS.t163 VSS.t162 VSS.t163 VSS.t133 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X539 RES_74k_1.M.t1 VSS.t53 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X540 RES_74k_1.M.t1 VSS.t52 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X541 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t24 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t17 VSS.t675 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X542 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t48 VDD.t194 VDD.t193 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X543 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT a_41879_n196.t8 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t14 VDD.t146 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X544 VDD mux_magic_3.AND2_magic_0.A.t10 a_19903_8443.t1 VDD.t412 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X545 mux_magic_2.AND2_magic_0.A S1.t6 VSS.t462 VSS.t461 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X546 a_44128_12082.t1 a_43828_11460.t1 VDD.t5 ppolyf_u r_width=1.1u r_length=2.6u
X547 VSS VCTRL2.t46 a_25706_n567.t16 VSS.t292 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X548 RES_74k_1.M.t1 VSS.t51 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X549 VDD VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t26 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t10 VDD.t448 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X550 OUTB OUT.t25 VSS.t544 VSS.t543 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X551 VDD PRE_SCALAR.t2 a_19897_11741.t5 VDD.t527 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X552 PFD_T2_0.INV_mag_1.IN PFD_T2_0.FDIV.t5 a_22881_9554.t3 VSS.t728 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X553 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t25 OUTB.t14 VSS.t668 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X554 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCTRL.t28 VDD.t94 VDD.t66 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X555 UP a_29262_10725.t8 VDD.t215 VDD.t213 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X556 PFD_T2_0.INV_mag_0.IN PFD_T2_0.INV_mag_0.IN.t14 a_24436_11277.t2 VDD.t227 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X557 RES_74k_1.M.t1 VSS.t50 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X558 OUTB OUT.t26 VSS.t546 VSS.t545 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X559 VDD a_27875_8520.t7 mux_magic_1.OR_magic_0.A.t1 VDD.t326 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X560 RES_74k_1.M.t1 VSS.t49 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X561 VSS.t161 VSS.t159 VSS.t161 VSS.t160 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X562 RES_74k_1.M.t1 VSS.t48 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X563 VDD PFD_T2_0.INV_mag_1.IN.t29 a_24436_11277.t0 VDD.t475 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X564 a_43828_11254.t1 a_44128_10632.t0 VDD.t5 ppolyf_u r_width=1.1u r_length=2.6u
X565 a_46528_10426.t1 a_46828_9598.t1 VDD.t102 ppolyf_u r_width=1.1u r_length=2.6u
X566 PFD_T2_0.FDIV a_21443_9476.t7 VSS.t759 VSS.t758 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X567 a_43528_10426.t0 a_43228_9804.t1 VDD.t104 ppolyf_u r_width=1.1u r_length=2.6u
X568 VDD a_27875_9714.t7 mux_magic_1.OR_magic_0.B.t1 VDD.t828 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X569 PFD_T2_0.FDIV a_21443_9476.t8 VDD.t787 VDD.t81 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X570 VDD OUT.t27 OUTB.t7 VDD.t350 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X571 VSS PFD_T2_0.INV_mag_1.OUT.t7 a_22880_9797.t2 VSS.t493 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X572 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t49 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t7 VDD.t170 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X573 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t47 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t7 VDD.t625 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X574 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t50 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t6 VDD.t187 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X575 VDD.t40 VDD.t39 VDD.t40 VDD.t19 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X576 RES_74k_1.M.t1 VSS.t47 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X577 VSS VCTRL2.t49 a_25706_n567.t15 VSS.t320 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X578 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t18 VDD.t661 VDD.t660 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X579 VDD OUT.t28 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t7 VDD.t418 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X580 VDD VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t22 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t12 VDD.t682 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X581 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t51 VDD.t199 VDD.t173 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X582 VSS VCTRL2.t51 a_34443_2598.t13 VSS.t342 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X583 RES_74k_1.P ITAIL1.t11 a_31940_9626.t2 VSS.t613 nfet_03v3 ad=0.158p pd=1.64u as=92.8f ps=0.92u w=0.28u l=0.56u
X584 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t51 VDD.t817 VDD.t364 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X585 RES_74k_1.P.t87 RES_74k_1.P.t88 VDD.t99 ppolyf_u r_width=1.1u r_length=2.6u
X586 VDD.t38 VDD.t36 VDD.t38 VDD.t37 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X587 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.VCO_C_0.OUTB.t35 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t2 VSS.t753 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X588 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t52 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t5 VDD.t386 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X589 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t27 VSS.t557 VSS.t556 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X590 OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t21 VDD.t356 VDD.t355 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X591 VDD VCO_DFF_C_0.VCO_C_0.OUTB.t36 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t7 VDD.t688 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X592 PFD_T2_0.INV_mag_0.IN a_22966_11778.t11 VDD.t317 VDD.t316 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X593 a_44728_10426.t0 a_45028_9804.t0 VDD.t99 ppolyf_u r_width=1.1u r_length=2.6u
X594 VSS VCTRL2.t53 a_25706_n567.t13 VSS.t276 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X595 RES_74k_1.M.t1 VSS.t46 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X596 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.OUT.t20 a_25706_n567.t48 VSS.t658 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X597 VDD PFD_T2_0.DOWN.t5 a_27875_8520.t4 VDD.t208 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X598 a_46228_9598.t0 a_46528_8976.t0 VDD.t79 ppolyf_u r_width=1.1u r_length=2.6u
X599 RES_74k_1.M.t1 VSS.t45 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X600 a_43228_9598.t0 a_42928_8976.t0 VDD.t98 ppolyf_u r_width=1.1u r_length=2.6u
X601 VDD ITAIL.t6 ITAIL.t7 VDD.t145 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X602 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t52 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t5 VDD.t175 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X603 RES_74k_1.M.t1 VSS.t44 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X604 VDD S2.t9 mux_magic_0.AND2_magic_0.A.t4 VDD.t340 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X605 OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t22 VDD.t357 VDD.t353 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X606 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.VCO_C_0.OUTB.t37 VDD.t754 VDD.t679 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X607 mux_magic_3.AND2_magic_0.A S6.t7 VDD.t233 VDD.t228 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X608 VDD S4.t14 a_42763_5679.t2 VDD.t258 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X609 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t28 VDD.t458 VDD.t446 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X610 a_44728_12082.t1 a_45028_11460.t1 VDD.t99 ppolyf_u r_width=1.1u r_length=2.6u
X611 VSS.t158 VSS.t156 VSS.t158 VSS.t157 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X612 VSS VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t23 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t4 VSS.t558 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X613 VSS VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t19 VCO_DFF_C_0.VCO_C_0.OUTB.t1 VSS.t696 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X614 VDD DN_INPUT.t3 a_27875_9714.t0 VDD.t546 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X615 a_44728_8770.t1 a_44428_8148.t1 VDD.t106 ppolyf_u r_width=1.1u r_length=2.6u
X616 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t48 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t12 VDD.t187 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X617 RES_74k_1.M.t1 VSS.t43 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X618 RES_74k_1.M.t1 VSS.t42 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X619 VSS.t155 VSS.t153 VSS.t155 VSS.t154 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X620 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t49 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t6 VDD.t634 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X621 VSS VCTRL2.t54 a_34443_2598.t12 VSS.t309 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X622 VDD S1.t8 mux_magic_2.AND2_magic_0.A.t6 VDD.t273 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X623 VSS PRE_SCALAR.t3 a_20097_11741.t3 VSS.t639 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X624 PFD_T2_0.FIN a_21437_10708.t8 VDD.t152 VDD.t150 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X625 ITAIL ITAIL.t4 VDD.t541 VDD.t143 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X626 VSS VCTRL2.t55 a_34443_2598.t11 VSS.t379 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X627 VDD.t35 VDD.t33 VDD.t35 VDD.t34 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X628 VDD a_19903_9637.t7 mux_magic_3.OR_magic_0.B.t1 VDD.t500 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X629 RES_74k_1.M.t1 VSS.t41 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X630 VDD VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t24 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t11 VDD.t682 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X631 a_45028_11254.t1 a_44728_10632.t0 VDD.t99 ppolyf_u r_width=1.1u r_length=2.6u
X632 RES_74k_1.P.t54 RES_74k_1.P.t55 VDD.t106 ppolyf_u r_width=1.1u r_length=2.6u
X633 VDD.t32 VDD.t30 VDD.t32 VDD.t31 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X634 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t50 VDD.t637 VDD.t185 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X635 RES_74k_1.M.t1 VSS.t40 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X636 VSS VCO_DFF_C_0.VCO_C_0.OUTB.t39 a_44716_1837.t0 VSS.t746 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X637 VDD PFD_T2_0.INV_mag_0.IN.t28 PFD_T2_0.INV_mag_0.OUT.t1 VDD.t157 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X638 VSS.t152 VSS.t150 VSS.t152 VSS.t151 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X639 VSS.t149 VSS.t147 VSS.t149 VSS.t148 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X640 VDD PFD_T2_0.UP.t4 a_27722_11758.t4 VDD.t518 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X641 PFD_T2_0.INV_mag_0.OUT PFD_T2_0.INV_mag_0.IN.t29 VSS.t582 VSS.t581 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.5u
X642 PFD_T2_0.INV_mag_1.IN a_22967_8787.t13 VDD.t131 VDD.t130 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X643 VDD a_22966_11778.t12 PFD_T2_0.INV_mag_0.IN.t0 VDD.t291 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X644 VSS VCTRL2.t56 a_34443_2598.t10 VSS.t309 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X645 VDD PFD_T2_0.INV_mag_0.IN.t30 PFD_T2_0.Buffer_V_2_1.IN.t4 VDD.t291 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X646 VSS PFD_T2_0.INV_mag_1.IN.t30 a_23837_9553.t0 VSS.t263 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X647 RES_74k_1.M.t1 VSS.t39 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X648 VDD a_22966_11778.t13 PFD_T2_0.INV_mag_0.IN.t1 VDD.t294 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X649 a_45928_8770.t1 a_46228_8148.t1 VDD.t107 ppolyf_u r_width=1.1u r_length=2.6u
X650 RES_74k_1.M.t1 VSS.t38 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X651 VSS PFD_T2_0.INV_mag_0.OUT.t9 PFD_T2_0.Buffer_V_2_0.IN.t10 VSS.t493 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X652 VDD VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t17 VCO_DFF_C_0.VCO_C_0.OUT.t8 VDD.t491 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X653 VDD PFD_T2_0.FIN.t5 a_22966_11778.t2 VDD.t294 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X654 ITAIL ITAIL.t2 VDD.t540 VDD.t139 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X655 VSS VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t53 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t0 VSS.t271 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X656 DN a_29415_9553.t8 VSS.t243 VSS.t242 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X657 VCO_DFF_C_0.VCTRL a_42763_5679.t8 VCTRL_IN.t5 VDD.t257 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X658 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t53 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t11 VDD.t368 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X659 RES_74k_1.M.t1 VSS.t37 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X660 RES_74k_1.P.t70 RES_74k_1.P.t71 VDD.t107 ppolyf_u r_width=1.1u r_length=2.6u
X661 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t25 VDD.t687 VDD.t679 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X662 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t20 VCO_DFF_C_0.VCO_C_0.OUTB.t6 VDD.t216 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X663 VDD PFD_T2_0.Buffer_V_2_1.IN.t12 a_25556_11637.t1 VDD.t505 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X664 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN a_44716_n517.t8 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t6 VDD.t566 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X665 VDD VCO_DFF_C_0.VCO_C_0.OUTB.t40 a_41879_n196.t5 VDD.t149 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X666 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t52 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t3 VDD.t398 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X667 PFD_T2_0.INV_mag_1.IN PFD_T2_0.INV_mag_1.IN.t0 a_24437_9224.t0 VDD.t464 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X668 VDD S6.t8 mux_magic_3.AND2_magic_0.A.t4 VDD.t230 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X669 VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t18 VDD.t494 VDD.t489 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X670 RES_74k_1.M.t1 VSS.t36 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X671 VDD VCO_DFF_C_0.VCTRL.t29 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t29 VDD.t88 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X672 RES_74k_1.M.t1 VSS.t35 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X673 RES_74k_1.M.t1 VSS.t34 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X674 PFD_T2_0.Buffer_V_2_0.IN PFD_T2_0.INV_mag_1.IN.t32 VDD.t478 VDD.t130 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X675 RES_74k_1.M.t1 VSS.t33 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X676 RES_74k_1.M.t1 VSS.t32 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X677 VDD VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t23 OUT.t7 VDD.t347 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X678 a_42928_10426.t1 a_42628_9804.t1 VDD.t101 ppolyf_u r_width=1.1u r_length=2.6u
X679 A_MUX_0.Tr_Gate_1.CLK S4.t15 VDD.t718 VDD.t711 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X680 VCO_DFF_C_0.VCTRL A_MUX_0.Tr_Gate_1.CLK.t20 RES_74k_1.P.t26 VSS.t248 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X681 VDD.t29 VDD.t27 VDD.t29 VDD.t28 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X682 VCO_DFF_C_0.VCTRL a_45158_5339.t9 RES_74k_1.P.t106 VDD.t723 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X683 VDD a_27722_11758.t8 mux_magic_0.OR_magic_0.A.t1 VDD.t531 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X684 VDD.t26 VDD.t24 VDD.t26 VDD.t25 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X685 VSS UP_INPUT.t3 a_27922_10564.t3 VSS.t628 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X686 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t51 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t14 VDD.t165 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X687 RES_74k_1.M.t1 VSS.t31 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X688 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t26 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t10 VSS.t665 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X689 A_MUX_0.Tr_Gate_1.CLK S4.t16 VDD.t719 VDD.t713 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X690 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN a_41879_1284.t8 OUTB.t17 VDD.t148 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X691 A_MUX_0.Tr_Gate_1.CLK S4.t17 VSS.t723 VSS.t715 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X692 VSS VCTRL2.t61 a_34443_2598.t8 VSS.t325 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X693 VSS VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t29 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t13 VSS.t558 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X694 VSS PFD_T2_0.UP.t5 a_27922_11758.t3 VSS.t634 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X695 mux_magic_1.AND2_magic_0.A S3.t9 VSS.t664 VSS.t663 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X696 VCO_DFF_C_0.VCTRL S4.t18 VCTRL_IN.t1 VSS.t724 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X697 RES_74k_1.M.t1 VSS.t30 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X698 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCTRL.t30 VDD.t785 VDD.t47 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.84u
X699 a_44128_10426.t1 a_44428_9804.t1 VDD.t105 ppolyf_u r_width=1.1u r_length=2.6u
X700 VSS VCTRL2.t62 a_25706_n567.t9 VSS.t292 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X701 RES_74k_1.M.t1 VSS.t29 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X702 a_45628_9598.t1 a_45928_8976.t0 VDD.t100 ppolyf_u r_width=1.1u r_length=2.6u
X703 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t54 VDD.t202 VDD.t193 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X704 VSS a_22966_11778.t14 a_22880_10947.t0 VSS.t470 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X705 a_42628_9598.t1 a_42628_8770.t1 VDD.t78 ppolyf_u r_width=1.1u r_length=2.6u
X706 RES_74k_1.M.t4 VSS.t28 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X707 A_MUX_0.Tr_Gate_1.CLK S4.t19 VSS.t725 VSS.t715 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X708 VDD.t23 VDD.t21 VDD.t23 VDD.t22 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X709 VCTRL_IN a_42763_5679.t9 VCO_DFF_C_0.VCTRL.t7 VDD.t258 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X710 VSS VCTRL2.t64 a_34443_2598.t6 VSS.t325 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X711 RES_74k_1.M.t1 VSS.t27 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X712 RES_74k_1.M.t1 VSS.t26 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X713 VSS VCTRL2.t65 a_25706_n567.t8 VSS.t320 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X714 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t55 VDD.t203 VDD.t160 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X715 VSS.t146 VSS.t144 VSS.t146 VSS.t145 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X716 VDD a_19897_11741.t8 mux_magic_2.OR_magic_0.A.t1 VDD.t654 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X717 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t52 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t15 VDD.t162 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X718 VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t19 VSS.t607 VSS.t606 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X719 VSS VCTRL2.t67 a_34443_2598.t4 VSS.t281 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X720 mux_magic_3.AND2_magic_0.A S6.t10 VDD.t236 VDD.t132 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X721 RES_74k_1.M.t1 VSS.t25 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X722 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t53 VDD.t642 VDD.t193 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X723 VDD S3.t10 mux_magic_1.AND2_magic_0.A.t7 VDD.t570 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X724 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.OUTB.t42 a_25706_n567.t57 VSS.t659 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X725 a_43828_9598.t1 a_44128_8976.t1 VDD.t5 ppolyf_u r_width=1.1u r_length=2.6u
X726 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT a_44716_n517.t9 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t15 VDD.t567 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X727 VSS VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t24 OUT.t8 VSS.t516 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X728 VDD a_22966_11778.t15 PFD_T2_0.INV_mag_0.IN.t2 VDD.t297 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X729 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t54 VSS.t693 VSS.t264 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X730 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t54 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t12 VDD.t398 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X731 RES_74k_1.M.t1 VSS.t24 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X732 VSS.t143 VSS.t141 VSS.t143 VSS.t142 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X733 a_45328_8770.t0 a_45628_8148.t1 VDD.t3 ppolyf_u r_width=1.1u r_length=2.6u
X734 PFD_T2_0.INV_mag_1.IN a_22967_8787.t14 VDD.t243 VDD.t242 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X735 RES_74k_1.P.t89 RES_74k_1.P.t90 VDD.t108 ppolyf_u r_width=1.1u r_length=2.6u
X736 VSS.t140 VSS.t138 VSS.t140 VSS.t139 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X737 RES_74k_1.M.t1 VSS.t23 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X738 RES_74k_1.P.t91 RES_74k_1.P.t92 VDD.t100 ppolyf_u r_width=1.1u r_length=2.6u
X739 VSS VCTRL2.t69 a_25706_n567.t6 VSS.t276 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X740 VDD VCO_DFF_C_0.VCO_C_0.OUTB.t43 a_44716_1837.t2 VDD.t565 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X741 RES_74k_1.M.t1 VSS.t22 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X742 RES_74k_1.P A_MUX_0.Tr_Gate_1.CLK.t21 VCO_DFF_C_0.VCTRL.t0 VSS.t249 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X743 VDD VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t26 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t9 VDD.t688 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X744 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t21 VCO_DFF_C_0.VCO_C_0.OUTB.t5 VDD.t657 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X745 RES_74k_1.M.t7 VSS.t21 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X746 RES_74k_1.P.t93 RES_74k_1.P.t94 VDD.t3 ppolyf_u r_width=1.1u r_length=2.6u
X747 RES_74k_1.P.t95 RES_74k_1.P.t96 VDD.t108 ppolyf_u r_width=1.1u r_length=2.6u
X748 RES_74k_1.M.t1 VSS.t20 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X749 RES_74k_1.P.t112 VSS.t435 cap_mim_2f0_m4m5_noshield c_width=30u c_length=30u
X750 VDD VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t20 VCO_DFF_C_0.VCO_C_0.OUT.t6 VDD.t491 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X751 RES_74k_1.M.t1 VSS.t19 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X752 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN a_41879_n196.t9 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t19 VDD.t147 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X753 VDD.t20 VDD.t18 VDD.t20 VDD.t19 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X754 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.VCO_C_0.OUTB.t45 VSS.t757 VSS.t756 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X755 VDD VCO_DFF_C_0.VCTRL.t31 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t17 VDD.t47 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X756 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t55 VDD.t407 VDD.t382 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X757 VDD S6.t11 a_19903_9637.t2 VDD.t237 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X758 RES_74k_1.M.t1 VSS.t18 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X759 a_45928_12082.t1 a_45628_11460.t1 VDD.t100 ppolyf_u r_width=1.1u r_length=2.6u
X760 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t19 a_34443_2598.t47 VSS.t481 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X761 RES_74k_1.M.t1 VSS.t17 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X762 VDD a_25556_11637.t5 PFD_T2_0.UP.t2 VDD.t515 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X763 OUTB a_41879_1284.t9 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t11 VDD.t149 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X764 RES_74k_1.P.t81 RES_74k_1.P.t82 VDD.t80 ppolyf_u r_width=1.1u r_length=2.6u
X765 RES_74k_1.M.t1 VSS.t16 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X766 OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t25 VDD.t361 VDD.t355 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X767 OUTB VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t27 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t0 VSS.t671 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X768 RES_74k_1.M.t1 VSS.t15 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X769 RES_74k_1.M.t1 VSS.t14 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X770 RES_74k_1.P.t113 VSS.t434 cap_mim_2f0_m4m5_noshield c_width=30u c_length=30u
X771 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t21 a_34443_2598.t50 VSS.t245 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X772 mux_magic_0.AND2_magic_0.A S2.t10 VSS.t506 VSS.t505 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X773 VDD PFD_T2_0.Buffer_V_2_0.IN.t13 a_25557_8739.t1 VDD.t95 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X774 a_45628_11254.t1 a_45928_10632.t1 VDD.t100 ppolyf_u r_width=1.1u r_length=2.6u
X775 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t30 VDD.t459 VDD.t454 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X776 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.VCO_C_0.OUTB.t46 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t1 VSS.t753 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X777 mux_magic_2.OR_magic_0.B a_19897_10547.t8 VSS.t497 VSS.t496 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X778 RES_74k_1.P.t83 RES_74k_1.P.t84 VDD.t80 ppolyf_u r_width=1.1u r_length=2.6u
X779 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t55 VDD.t643 VDD.t185 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X780 RES_74k_1.M.t1 VSS.t13 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X781 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.VCO_C_0.OUTB.t47 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t0 VSS.t739 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X782 RES_74k_1.P ITAIL.t26 a_31732_10267.t1 VDD.t139 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X783 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t53 VDD.t820 VDD.t789 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X784 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t54 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t2 VDD.t372 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X785 VSS PFD_T2_0.INV_mag_1.OUT.t8 PFD_T2_0.Buffer_V_2_1.IN.t1 VSS.t569 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X786 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t56 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t5 VDD.t180 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X787 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t56 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t5 VDD.t634 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X788 VSS.t137 VSS.t135 VSS.t137 VSS.t136 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X789 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t56 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t14 VDD.t389 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X790 OUTB OUT.t29 VDD.t438 VDD.t355 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X791 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t29 OUTB.t12 VSS.t677 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X792 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t22 VDD.t221 VDD.t219 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X793 VDD.t17 VDD.t15 VDD.t17 VDD.t16 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X794 VSS OUT.t30 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t0 VSS.t516 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X795 VSS VCTRL2.t73 a_25706_n567.t4 VSS.t292 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X796 VSS PFD_T2_0.INV_mag_1.OUT.t9 PFD_T2_0.Buffer_V_2_1.IN.t0 VSS.t575 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X797 mux_magic_1.OR_magic_0.A a_27875_8520.t8 VSS.t499 VSS.t498 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X798 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t57 VDD.t206 VDD.t183 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X799 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT a_44716_1837.t8 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t18 VDD.t564 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X800 VSS PFD_T2_0.Buffer_V_2_1.IN.t13 a_25556_11637.t0 VSS.t623 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X801 RES_74k_1.M.t6 VSS.t12 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X802 OUTB OUT.t31 VDD.t439 VDD.t353 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X803 a_43528_10426.t1 a_43828_9804.t1 VDD.t4 ppolyf_u r_width=1.1u r_length=2.6u
X804 VSS S4.t20 a_42763_5679.t0 VSS.t720 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X805 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN OUT.t32 VDD.t440 VDD.t425 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X806 VSS VCTRL2.t74 a_34443_2598.t1 VSS.t342 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X807 mux_magic_1.OR_magic_0.B a_27875_9714.t8 VSS.t761 VSS.t760 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X808 mux_magic_1.AND2_magic_0.A S3.t11 VDD.t575 VDD.t487 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X809 RES_74k_1.P.t50 RES_74k_1.P.t51 VDD.t101 ppolyf_u r_width=1.1u r_length=2.6u
X810 PFD_T2_0.INV_mag_0.IN PFD_T2_0.FIN.t6 a_22880_10947.t2 VSS.t485 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X811 RES_74k_1.P.t52 RES_74k_1.P.t53 VDD.t102 ppolyf_u r_width=1.1u r_length=2.6u
X812 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t55 VDD.t823 VDD.t375 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X813 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t57 VDD.t410 VDD.t380 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X814 RES_74k_1.M.t1 VSS.t11 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X815 VDD OUT.t33 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t5 VDD.t429 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X816 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN OUT.t34 VDD.t443 VDD.t427 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X817 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t58 VDD.t207 VDD.t185 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X818 VDD VCO_DFF_C_0.VCTRL.t32 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t16 VDD.t85 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X819 RES_74k_1.M.t1 VSS.t10 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X820 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t56 VSS.t773 VSS.t772 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X821 VDD VCO_DFF_C_0.VCO_C_0.OUTB.t49 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t5 VDD.t682 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X822 VDD.t14 VDD.t12 VDD.t14 VDD.t13 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X823 VSS VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t21 VCO_DFF_C_0.VCO_C_0.OUT.t0 VSS.t608 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X824 RES_74k_1.M.t1 VSS.t9 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X825 VDD VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t31 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t15 VDD.t451 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X826 VDD VCO_DFF_C_0.VCO_C_0.OUTB.t51 a_41879_n196.t2 VDD.t146 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X827 VDD ITAIL.t0 ITAIL.t1 VDD.t145 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X828 a_42928_12082.t0 a_42628_11460.t0 VDD.t101 ppolyf_u r_width=1.1u r_length=2.6u
X829 a_46528_12082.t0 a_46828_11254.t0 VDD.t102 ppolyf_u r_width=1.1u r_length=2.6u
X830 VSS VCTRL2.t77 a_34443_2598.t0 VSS.t342 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X831 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t23 VSS.t428 VSS.t427 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X832 RES_74k_1.M.t1 VSS.t8 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X833 mux_magic_0.AND2_magic_0.A S2.t11 VSS.t508 VSS.t507 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X834 RES_74k_1.M.t1 VSS.t7 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X835 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.VCO_C_0.OUTB.t52 VDD.t766 VDD.t677 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X836 mux_magic_2.AND2_magic_0.A S1.t10 VDD.t281 VDD.t269 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X837 a_45328_10426.t0 a_45028_9804.t1 VDD.t103 ppolyf_u r_width=1.1u r_length=2.6u
X838 OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t26 VSS.t520 VSS.t519 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X839 VDD VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t27 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t8 VDD.t688 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X840 a_46828_9598.t0 a_46528_8976.t1 VDD.t102 ppolyf_u r_width=1.1u r_length=2.6u
X841 RES_74k_1.M.t1 VSS.t6 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X842 VSS mux_magic_1.OR_magic_0.A.t7 a_29415_9553.t5 VSS.t466 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X843 a_43228_9598.t1 a_43528_8976.t0 VDD.t104 ppolyf_u r_width=1.1u r_length=2.6u
X844 VDD VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t27 OUT.t11 VDD.t350 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X845 VDD VCO_DFF_C_0.VCTRL.t33 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t0 VDD.t66 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X846 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t57 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t18 VDD.t175 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X847 VDD S1.t11 a_19897_10547.t3 VDD.t282 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X848 PFD_T2_0.INV_mag_1.IN a_22967_8787.t16 VDD.t245 VDD.t244 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X849 a_42628_11254.t1 a_42928_10632.t1 VDD.t101 ppolyf_u r_width=1.1u r_length=2.6u
X850 VSS.t134 VSS.t132 VSS.t134 VSS.t133 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X851 VDD a_22966_11778.t16 PFD_T2_0.INV_mag_0.IN.t3 VDD.t300 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X852 mux_magic_3.AND2_magic_0.A S6.t12 VSS.t444 VSS.t443 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X853 a_46828_11254.t1 a_46528_10632.t1 VDD.t102 ppolyf_u r_width=1.1u r_length=2.6u
X854 mux_magic_3.OR_magic_0.A a_19903_8443.t8 VSS.t653 VSS.t652 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X855 RES_74k_1.M.t1 VSS.t5 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X856 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t30 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t11 VSS.t670 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X857 RES_74k_1.P ITAIL1.t13 a_31940_9626.t0 VSS.t611 nfet_03v3 ad=0.158p pd=1.64u as=92.8f ps=0.92u w=0.28u l=0.56u
X858 VDD PFD_T2_0.INV_mag_0.IN.t32 PFD_T2_0.Buffer_V_2_1.IN.t3 VDD.t300 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X859 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t58 VDD.t648 VDD.t614 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X860 VDD S2.t12 mux_magic_0.AND2_magic_0.A.t3 VDD.t340 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X861 VDD VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t22 VCO_DFF_C_0.VCO_C_0.OUT.t5 VDD.t479 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X862 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.OUTB.t53 a_25706_n567.t59 VSS.t658 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X863 RES_74k_1.M.t1 VSS.t4 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X864 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t57 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t4 VDD.t795 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X865 VDD OUT.t35 OUTB.t4 VDD.t347 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X866 mux_magic_2.AND2_magic_0.A S1.t12 VSS.t465 VSS.t464 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X867 VDD VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t31 a_41879_1284.t2 VDD.t149 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X868 mux_magic_3.OR_magic_0.B a_19903_9637.t8 VSS.t622 VSS.t621 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X869 VCO_DFF_C_0.VCTRL S4.t21 VCTRL_IN.t0 VSS.t718 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X870 RES_74k_1.P.t114 VSS.t762 cap_mim_2f0_m4m5_noshield c_width=30u c_length=30u
X871 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t58 VDD.t411 VDD.t396 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X872 VSS VCTRL2.t78 a_25706_n567.t1 VSS.t297 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X873 VSS PFD_T2_0.INV_mag_0.IN.t33 a_23836_10693.t0 VSS.t561 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X874 VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t23 VDD.t483 VDD.t482 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X875 RES_74k_1.M.t1 VSS.t3 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X876 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT a_44716_1837.t9 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t15 VDD.t565 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X877 a_45028_9598.t1 a_44728_8976.t1 VDD.t99 ppolyf_u r_width=1.1u r_length=2.6u
X878 RES_74k_1.M.t1 VSS.t2 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X879 VDD VCO_DFF_C_0.VCTRL.t34 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t0 VDD.t88 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.84u
X880 RES_74k_1.P.t107 RES_74k_1.P.t108 VDD.t4 ppolyf_u r_width=1.1u r_length=2.6u
X881 RES_74k_1.M.t1 VSS.t1 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X882 mux_magic_0.OR_magic_0.B a_27722_10564.t8 VDD.t537 VDD.t536 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X883 VSS VCTRL2.t79 a_25706_n567.t0 VSS.t320 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X884 RES_74k_1.M.t5 VSS.t0 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X885 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t58 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t0 VDD.t389 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X886 PFD_T2_0.Buffer_V_2_0.IN PFD_T2_0.INV_mag_1.IN.t33 a_23837_9553.t3 VSS.t260 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X887 a_46528_8770.t0 a_46228_8148.t0 VDD.t79 ppolyf_u r_width=1.1u r_length=2.6u
X888 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCTRL.t35 VDD.t777 VDD.t47 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
R0 a_42928_8770.t0 a_42928_8770.t1 12.9675
R1 a_43228_8148.t0 a_43228_8148.t1 12.9675
R2 VDD.n1619 VDD.n421 130000
R3 VDD.n1400 VDD.n570 129000
R4 VDD.n1620 VDD.n1619 65000
R5 VDD.n1355 VDD.n570 64500
R6 VDD.n1809 VDD.n1808 6501.29
R7 VDD.n1567 VDD.n1566 947.995
R8 VDD.n1621 VDD.n413 947.995
R9 VDD.n1372 VDD.n1348 947.995
R10 VDD.n1363 VDD.n1356 947.995
R11 VDD.n1566 VDD.n1557 944.883
R12 VDD.n1557 VDD.n420 944.883
R13 VDD.n1365 VDD.n1364 944.883
R14 VDD.n1364 VDD.n1363 944.883
R15 VDD.n1621 VDD.n1620 842.52
R16 VDD.n1355 VDD.n1348 842.52
R17 VDD.t523 VDD.t332 669.359
R18 VDD.t269 VDD.t774 669.359
R19 VDD.t228 VDD.t415 669.359
R20 VDD.t303 VDD.t114 669.359
R21 VDD.n1809 VDD.n1748 447.029
R22 VDD.t465 VDD.t240 432.243
R23 VDD.t531 VDD.n84 421.245
R24 VDD.n84 VDD.t0 421.245
R25 VDD.n141 VDD.t654 421.245
R26 VDD.t321 VDD.n141 421.245
R27 VDD.n240 VDD.t558 421.245
R28 VDD.t500 VDD.n240 421.245
R29 VDD.n1898 VDD.t326 421.245
R30 VDD.t828 VDD.n1898 421.245
R31 VDD.t534 VDD.t531 395.604
R32 VDD.t518 VDD.t534 395.604
R33 VDD.t521 VDD.t259 395.604
R34 VDD.t259 VDD.t523 395.604
R35 VDD.t0 VDD.t536 395.604
R36 VDD.t536 VDD.t508 395.604
R37 VDD.t511 VDD.t329 395.604
R38 VDD.t329 VDD.t336 395.604
R39 VDD.t654 VDD.t652 395.604
R40 VDD.t652 VDD.t527 395.604
R41 VDD.t670 VDD.t525 395.604
R42 VDD.t774 VDD.t670 395.604
R43 VDD.t319 VDD.t321 395.604
R44 VDD.t589 VDD.t319 395.604
R45 VDD.t592 VDD.t282 395.604
R46 VDD.t282 VDD.t279 395.604
R47 VDD.t558 VDD.t556 395.604
R48 VDD.t556 VDD.t693 395.604
R49 VDD.t412 VDD.t696 395.604
R50 VDD.t415 VDD.t412 395.604
R51 VDD.t498 VDD.t500 395.604
R52 VDD.t109 VDD.t498 395.604
R53 VDD.t112 VDD.t237 395.604
R54 VDD.t237 VDD.t134 395.604
R55 VDD.t326 VDD.t324 395.604
R56 VDD.t324 VDD.t208 395.604
R57 VDD.t116 VDD.t211 395.604
R58 VDD.t114 VDD.t116 395.604
R59 VDD.t665 VDD.t828 395.604
R60 VDD.t546 VDD.t665 395.604
R61 VDD.t544 VDD.t561 395.604
R62 VDD.t561 VDD.t568 395.604
R63 VDD.n1618 VDD.n379 371.986
R64 VDD.n1388 VDD.n577 371.986
R65 VDD.n1606 VDD.n1605 353.928
R66 VDD.n1403 VDD.n567 353.928
R67 VDD.n1607 VDD.n1606 350.877
R68 VDD.n1611 VDD.n422 350.877
R69 VDD.n1399 VDD.n572 350.877
R70 VDD.n1403 VDD.n1402 350.877
R71 VDD.t503 VDD.t222 339.613
R72 VDD.t663 VDD.t667 316.279
R73 VDD.t240 VDD.t95 316.279
R74 VDD.n1611 VDD.n421 312.866
R75 VDD.n1400 VDD.n1399 312.866
R76 VDD.n1773 VDD.n1772 310.428
R77 VDD.n1774 VDD.n1773 307.495
R78 VDD.n1774 VDD.n1757 307.495
R79 VDD.n1759 VDD.n1758 307.495
R80 VDD.n1783 VDD.n1759 307.495
R81 VDD.n1806 VDD.n1750 307.495
R82 VDD.n1799 VDD.n1750 307.495
R83 VDD.n1797 VDD.n1796 307.495
R84 VDD.n1796 VDD.n1784 307.495
R85 VDD.n1789 VDD.n1748 307.495
R86 VDD.n1807 VDD.n1749 304.911
R87 VDD.t53 VDD.n1618 283.627
R88 VDD.n1388 VDD.t58 283.627
R89 VDD.t513 VDD.t515 282.159
R90 VDD.t505 VDD.t503 282.159
R91 VDD.n1609 VDD.t66 279.885
R92 VDD.t47 VDD.n1401 279.885
R93 VDD.t37 VDD.n1797 263.567
R94 VDD.t37 VDD.n1758 235.143
R95 VDD.t332 VDD.t340 233.011
R96 VDD.t273 VDD.t269 233.011
R97 VDD.t230 VDD.t228 233.011
R98 VDD.t570 VDD.t303 233.011
R99 VDD.n1922 VDD.t334 226.537
R100 VDD.n151 VDD.t271 226.537
R101 VDD.n250 VDD.t132 226.537
R102 VDD.n1908 VDD.t487 226.537
R103 VDD.t37 VDD.n1783 209.303
R104 VDD.n1923 VDD.t518 197.803
R105 VDD.n1923 VDD.t521 197.803
R106 VDD.t508 VDD.n83 197.803
R107 VDD.n83 VDD.t511 197.803
R108 VDD.t527 VDD.n132 197.803
R109 VDD.t525 VDD.n132 197.803
R110 VDD.n142 VDD.t589 197.803
R111 VDD.n142 VDD.t592 197.803
R112 VDD.t693 VDD.n231 197.803
R113 VDD.t696 VDD.n231 197.803
R114 VDD.n241 VDD.t109 197.803
R115 VDD.n241 VDD.t112 197.803
R116 VDD.n1907 VDD.t208 197.803
R117 VDD.t211 VDD.n1907 197.803
R118 VDD.n1899 VDD.t546 197.803
R119 VDD.n1899 VDD.t544 197.803
R120 VDD.t297 VDD.t308 188.018
R121 VDD.t308 VDD.t300 188.018
R122 VDD.t300 VDD.t223 188.018
R123 VDD.t223 VDD.t291 188.018
R124 VDD.t291 VDD.t225 188.018
R125 VDD.t225 VDD.t294 188.018
R126 VDD.t294 VDD.t312 188.018
R127 VDD.t95 VDD.n204 184.496
R128 VDD.n1784 VDD.t25 180.88
R129 VDD.t128 VDD.t734 180.213
R130 VDD.t120 VDD.t128 180.213
R131 VDD.t244 VDD.t123 180.213
R132 VDD.t123 VDD.t130 180.213
R133 VDD.t130 VDD.t724 180.213
R134 VDD.t724 VDD.t720 180.213
R135 VDD.n96 VDD.t505 164.593
R136 VDD.n205 VDD.t244 161.661
R137 VDD.n1436 VDD.t22 160.7
R138 VDD.n1595 VDD.t50 160.284
R139 VDD.n84 VDD.t264 145.662
R140 VDD.n141 VDD.t549 145.662
R141 VDD.n240 VDD.t9 145.662
R142 VDD.n1898 VDD.t285 145.662
R143 VDD.t608 VDD.t213 136.796
R144 VDD.t264 VDD.t262 136.796
R145 VDD.t576 VDD.t150 136.796
R146 VDD.t549 VDD.t318 136.796
R147 VDD.t555 VDD.t81 136.796
R148 VDD.t9 VDD.t250 136.796
R149 VDD.t358 VDD.t7 136.796
R150 VDD.t285 VDD.t6 136.796
R151 VDD.n1536 VDD.n1535 132.696
R152 VDD.n1527 VDD.n1526 132.696
R153 VDD.n1461 VDD.n1460 132.696
R154 VDD.n545 VDD.n502 132.696
R155 VDD.n527 VDD.n526 132.696
R156 VDD.n966 VDD.n965 132.696
R157 VDD.n1056 VDD.n1055 132.696
R158 VDD.n1475 VDD.n1472 132.696
R159 VDD.n204 VDD.t663 131.784
R160 VDD.n1537 VDD.n1536 128.591
R161 VDD.t618 VDD.n446 128.591
R162 VDD.n1543 VDD.n446 128.591
R163 VDD.n1545 VDD.n1544 128.591
R164 VDD.n1526 VDD.n1499 128.591
R165 VDD.n1509 VDD.t183 128.591
R166 VDD.n1519 VDD.n1509 128.591
R167 VDD.n1518 VDD.n1517 128.591
R168 VDD.n1453 VDD.n473 128.591
R169 VDD.n1455 VDD.n1454 128.591
R170 VDD.n1455 VDD.t386 128.591
R171 VDD.n1460 VDD.n464 128.591
R172 VDD.n559 VDD.n493 128.591
R173 VDD.n553 VDD.n552 128.591
R174 VDD.n552 VDD.t811 128.591
R175 VDD.n551 VDD.n502 128.591
R176 VDD.n536 VDD.n535 128.591
R177 VDD.n534 VDD.n511 128.591
R178 VDD.t657 VDD.n511 128.591
R179 VDD.n527 VDD.n522 128.591
R180 VDD.n957 VDD.n956 128.591
R181 VDD.n963 VDD.n940 128.591
R182 VDD.t429 VDD.n963 128.591
R183 VDD.n966 VDD.n964 128.591
R184 VDD.n1063 VDD.n1041 128.591
R185 VDD.t451 VDD.n1041 128.591
R186 VDD.n1056 VDD.n1049 128.591
R187 VDD.n1471 VDD.n1470 128.591
R188 VDD.n1484 VDD.n1483 128.591
R189 VDD.n1483 VDD.t491 128.591
R190 VDD.n1482 VDD.n1472 128.591
R191 VDD.n1789 VDD.t25 126.615
R192 VDD.n73 VDD.t608 122.23
R193 VDD.n124 VDD.t576 122.23
R194 VDD.n223 VDD.t555 122.23
R195 VDD.n1897 VDD.t358 122.23
R196 VDD.n1942 VDD.t255 122.1
R197 VDD.t723 VDD.n2004 121.091
R198 VDD.n1914 VDD.t157 120.213
R199 VDD.t222 VDD.t316 118.191
R200 VDD.t227 VDD.t305 118.191
R201 VDD.t468 VDD.t314 118.191
R202 VDD.n1490 VDD.t634 118.061
R203 VDD.n1528 VDD.t180 118.061
R204 VDD.n1462 VDD.t380 118.061
R205 VDD.t789 VDD.n544 118.061
R206 VDD.t660 VDD.n525 118.061
R207 VDD.t454 VDD.n1054 118.061
R208 VDD.n1476 VDD.t489 118.061
R209 VDD.n96 VDD.t513 117.567
R210 VDD.t256 VDD.n1940 116.044
R211 VDD.t242 VDD.t465 113.275
R212 VDD.t731 VDD.t464 113.275
R213 VDD.t126 VDD.t649 113.275
R214 VDD.n1544 VDD.t625 110.808
R215 VDD.t170 VDD.n1518 110.808
R216 VDD.t366 VDD.n1453 110.808
R217 VDD.t793 VDD.n493 110.808
R218 VDD.n535 VDD.t219 110.808
R219 VDD.n957 VDD.t425 110.808
R220 VDD.t482 VDD.n1471 110.808
R221 VDD.n1064 VDD.t446 109.439
R222 VDD.t475 VDD.t297 108.948
R223 VDD.n1941 VDD.t256 105.954
R224 VDD.n2005 VDD.t722 104.945
R225 VDD.t734 VDD.t740 104.418
R226 VDD.n1620 VDD.n420 102.362
R227 VDD.n1365 VDD.n1355 102.362
R228 VDD.n2005 VDD.t723 100.909
R229 VDD.t255 VDD.n1941 99.8996
R230 VDD.n1619 VDD.t66 99.5009
R231 VDD.t47 VDD.n570 99.0846
R232 VDD.n972 VDD.t427 98.4957
R233 VDD.t37 VDD.n1749 98.1917
R234 VDD.n1547 VDD.t614 97.5562
R235 VDD.n1914 VDD.t462 96.809
R236 VDD.t418 VDD.n955 95.9239
R237 VDD.n1512 VDD.t173 95.9239
R238 VDD.n1446 VDD.t377 95.9239
R239 VDD.n560 VDD.t795 95.9239
R240 VDD.n539 VDD.t216 95.9239
R241 VDD.n1467 VDD.t479 95.9239
R242 VDD.t44 VDD.n381 92.4235
R243 VDD.t34 VDD.n1387 92.4235
R244 VDD.n1940 VDD.t258 89.8088
R245 VDD.n2007 VDD.t248 88.7997
R246 VDD.n663 VDD.n662 86.1787
R247 VDD.t448 VDD.n1030 84.8158
R248 VDD.n2004 VDD.t252 84.7634
R249 VDD.n1942 VDD.t257 83.7543
R250 VDD.n1075 VDD.n1031 73.8719
R251 VDD.t37 VDD.n1757 72.3519
R252 VDD.t316 VDD.t227 70.1759
R253 VDD.t305 VDD.t468 70.1759
R254 VDD.t314 VDD.t475 70.1759
R255 VDD.n1607 VDD.t66 70.1759
R256 VDD.n1402 VDD.t47 70.1759
R257 VDD.t464 VDD.t242 67.2571
R258 VDD.t649 VDD.t731 67.2571
R259 VDD.t740 VDD.t126 67.2571
R260 VDD.t53 VDD.n422 67.252
R261 VDD.t58 VDD.n572 67.252
R262 VDD.n894 VDD.n878 66.348
R263 VDD.n895 VDD.n894 64.296
R264 VDD.t355 VDD.n874 64.296
R265 VDD.n911 VDD.n874 64.296
R266 VDD.n915 VDD.n914 64.296
R267 VDD.n921 VDD.n920 64.296
R268 VDD.n782 VDD.t148 61.8854
R269 VDD.n994 VDD.t565 60.8721
R270 VDD.n781 VDD.t149 60.7435
R271 VDD.t567 VDD.n996 59.702
R272 VDD.t147 VDD.n778 59.0509
R273 VDD.t564 VDD.n998 58.9084
R274 VDD.t566 VDD.n999 57.7119
R275 VDD.n888 VDD.t350 57.456
R276 VDD.n701 VDD.n700 56.5021
R277 VDD.n763 VDD.n762 56.5021
R278 VDD.n914 VDD.t347 55.4041
R279 VDD.n1816 VDD.n1742 54.5384
R280 VDD.n1133 VDD.n1132 54.5384
R281 VDD.n833 VDD.n692 53.3521
R282 VDD.n819 VDD.n740 53.3521
R283 VDD.n816 VDD.n815 53.3521
R284 VDD.n761 VDD.n757 53.3521
R285 VDD.n779 VDD.t147 52.7113
R286 VDD.n1672 VDD.n1671 52.4568
R287 VDD.n1287 VDD.n592 52.0405
R288 VDD.n1000 VDD.t566 51.7418
R289 VDD.n15 VDD.t143 51.2378
R290 VDD.t58 VDD.n570 50.3542
R291 VDD.n1619 VDD.t53 49.9381
R292 VDD.n1000 VDD.t567 49.7517
R293 VDD.n779 VDD.t149 49.6993
R294 VDD.t80 VDD.t102 49.5054
R295 VDD.t102 VDD.t79 49.5054
R296 VDD.t79 VDD.t107 49.5054
R297 VDD.t3 VDD.t100 49.5054
R298 VDD.t103 VDD.t3 49.5054
R299 VDD.t99 VDD.t103 49.5054
R300 VDD.t106 VDD.t99 49.5054
R301 VDD.t106 VDD.t105 49.5054
R302 VDD.t105 VDD.t5 49.5054
R303 VDD.t5 VDD.t4 49.5054
R304 VDD.t4 VDD.t104 49.5054
R305 VDD.t101 VDD.t98 49.5054
R306 VDD.t78 VDD.t101 49.5054
R307 VDD.t108 VDD.t78 49.5054
R308 VDD.n24 VDD.t145 47.9334
R309 VDD.t677 VDD.n807 46.5121
R310 VDD.n920 VDD.t353 46.5121
R311 VDD.n1679 VDD.n369 45.7957
R312 VDD.n1678 VDD.n370 45.7957
R313 VDD.n1685 VDD.n365 45.7957
R314 VDD.t168 VDD.n1686 45.7957
R315 VDD.n1705 VDD.n341 45.7957
R316 VDD.n1696 VDD.n1693 45.7957
R317 VDD.n1861 VDD.n275 45.7957
R318 VDD.n283 VDD.n282 45.7957
R319 VDD.n1854 VDD.n1853 45.7957
R320 VDD.n290 VDD.n284 45.7957
R321 VDD.n1847 VDD.n291 45.7957
R322 VDD.n302 VDD.n301 45.7957
R323 VDD.n310 VDD.n303 45.7957
R324 VDD.n1831 VDD.n309 45.7957
R325 VDD.n1732 VDD.n1731 45.7957
R326 VDD.n1740 VDD.n1733 45.7957
R327 VDD.n1817 VDD.n1741 45.7957
R328 VDD.n1140 VDD.n653 45.7957
R329 VDD.n1139 VDD.n655 45.7957
R330 VDD.n1148 VDD.n1147 45.7957
R331 VDD.n1157 VDD.n641 45.7957
R332 VDD.n646 VDD.n645 45.7957
R333 VDD.n1221 VDD.n632 45.7957
R334 VDD.n1231 VDD.n1230 45.7957
R335 VDD.n1238 VDD.n620 45.7957
R336 VDD.n1237 VDD.n621 45.7957
R337 VDD.n1245 VDD.n616 45.7957
R338 VDD.n1255 VDD.n610 45.7957
R339 VDD.n1262 VDD.n606 45.7957
R340 VDD.n1272 VDD.n600 45.7957
R341 VDD.n1278 VDD.n596 45.7957
R342 VDD.n1280 VDD.n1279 45.7957
R343 VDD.n1288 VDD.n591 45.7957
R344 VDD.n1271 VDD.t398 45.3794
R345 VDD.n820 VDD.n739 45.1441
R346 VDD.n1799 VDD.t37 43.9281
R347 VDD.n999 VDD.t564 43.7816
R348 VDD.t165 VDD.n1823 43.2978
R349 VDD.n654 VDD.t382 42.8814
R350 VDD.t364 VDD.n1246 42.8814
R351 VDD.n1860 VDD.t162 42.4651
R352 VDD.n996 VDD.t565 41.7915
R353 VDD.n0 VDD.t80 41.7644
R354 VDD.n1930 VDD.t108 41.7644
R355 VDD.t148 VDD.n781 41.6672
R356 VDD.n1545 VDD.t614 39.6722
R357 VDD.n1517 VDD.t173 39.6722
R358 VDD.t377 VDD.n473 39.6722
R359 VDD.t795 VDD.n559 39.6722
R360 VDD.n536 VDD.t216 39.6722
R361 VDD.n746 VDD.n745 39.6722
R362 VDD.n956 VDD.t418 39.6722
R363 VDD.n1470 VDD.t479 39.6722
R364 VDD.n1966 VDD.t713 39.6722
R365 VDD.n1670 VDD.n374 39.5509
R366 VDD.n1378 VDD.n586 39.5509
R367 VDD.n1658 VDD.n381 38.3019
R368 VDD.n643 VDD.t372 38.3019
R369 VDD.n1387 VDD.n578 38.3019
R370 VDD.n1609 VDD.n421 37.9019
R371 VDD.n1401 VDD.n1400 37.9019
R372 VDD.n311 VDD.t185 37.8856
R373 VDD.n300 VDD.t193 36.2203
R374 VDD.n1597 VDD.n429 35.8675
R375 VDD.n1409 VDD.n1408 35.8675
R376 VDD.n631 VDD.t368 35.804
R377 VDD.n718 VDD.t688 35.5682
R378 VDD.n28 VDD.t136 33.5535
R379 VDD.n1077 VDD.t448 32.8322
R380 VDD.n1569 VDD.n1568 32.7175
R381 VDD.n1438 VDD.n477 32.7175
R382 VDD.n1658 VDD.n382 32.0571
R383 VDD.n1379 VDD.n578 32.0571
R384 VDD.n661 VDD.t63 31.6415
R385 VDD.n1692 VDD.t187 31.6408
R386 VDD.n1264 VDD.t396 31.2245
R387 VDD.n5 VDD.t594 31.1569
R388 VDD.n382 VDD.n374 30.8082
R389 VDD.n1379 VDD.n1378 30.8082
R390 VDD.n1065 VDD.n1031 30.0963
R391 VDD.n1029 VDD.n1020 28.8809
R392 VDD.t389 VDD.n611 28.7266
R393 VDD.n1698 VDD.t160 28.3102
R394 VDD.n1628 VDD.n1627 28.1746
R395 VDD.n1373 VDD.n588 28.1746
R396 VDD.n175 VDD.n93 26.1348
R397 VDD.n778 VDD.t146 24.6667
R398 VDD.n1076 VDD.n1075 24.6243
R399 VDD.n1222 VDD.t375 24.147
R400 VDD.n1839 VDD.t175 23.7307
R401 VDD.n1553 VDD.n1552 23.2342
R402 VDD.n1969 VDD.n1964 23.2342
R403 VDD.t175 VDD.n1838 22.0654
R404 VDD.t625 VDD.n1543 21.8883
R405 VDD.n1519 VDD.t170 21.8883
R406 VDD.n1454 VDD.t366 21.8883
R407 VDD.n553 VDD.t793 21.8883
R408 VDD.t219 VDD.n534 21.8883
R409 VDD.t425 VDD.n940 21.8883
R410 VDD.t446 VDD.n1063 21.8883
R411 VDD.n1484 VDD.t482 21.8883
R412 VDD.n1982 VDD.t698 21.8883
R413 VDD.n644 VDD.t375 21.6491
R414 VDD.n1131 VDD.t13 21.2328
R415 VDD.t37 VDD.n1798 20.8165
R416 VDD.n1554 VDD.n1553 20.395
R417 VDD.n1969 VDD.n1965 20.3898
R418 VDD.n915 VDD.t353 19.8363
R419 VDD.t76 VDD.n1670 19.5675
R420 VDD.t16 VDD.n586 19.5675
R421 VDD.n973 VDD.n972 19.0194
R422 VDD.n205 VDD.t120 18.5517
R423 VDD.n1094 VDD.n658 17.5593
R424 VDD.t160 VDD.n1697 17.4859
R425 VDD.n1254 VDD.t389 17.0696
R426 VDD.n1772 VDD.n1765 16.2393
R427 VDD.t396 VDD.n1263 14.5717
R428 VDD.t262 VDD.n73 14.5667
R429 VDD.t318 VDD.n124 14.5667
R430 VDD.t250 VDD.n223 14.5667
R431 VDD.t6 VDD.n1897 14.5667
R432 VDD.n1704 VDD.t187 14.1554
R433 VDD.n1535 VDD.t634 13.6804
R434 VDD.t180 VDD.n1527 13.6804
R435 VDD.t380 VDD.n1461 13.6804
R436 VDD.n545 VDD.t789 13.6804
R437 VDD.n526 VDD.t660 13.6804
R438 VDD.n745 VDD.n693 13.6804
R439 VDD.n965 VDD.t427 13.6804
R440 VDD.n1055 VDD.t454 13.6804
R441 VDD.t489 VDD.n1475 13.6804
R442 VDD.n1993 VDD.t706 13.6804
R443 VDD.n1669 VDD.n368 13.33
R444 VDD.n1286 VDD.n585 13.2637
R445 VDD.n717 VDD.n692 12.9964
R446 VDD.n808 VDD.n761 12.9964
R447 VDD.n1673 VDD.n373 11.6418
R448 VDD.n1377 VDD.n587 11.6418
R449 VDD.n1617 VDD.n424 11.2373
R450 VDD.n1669 VDD.n375 11.2079
R451 VDD.n1380 VDD.n585 11.2079
R452 VDD.n1389 VDD.n576 11.1709
R453 VDD.n1126 VDD.n659 11.094
R454 VDD.n718 VDD.n716 10.9444
R455 VDD.n820 VDD.n819 10.9444
R456 VDD.t682 VDD.n740 10.9444
R457 VDD.n815 VDD.n757 10.9444
R458 VDD.n807 VDD.n762 10.9444
R459 VDD.n911 VDD.t347 10.9444
R460 VDD.n955 VDD.n954 10.723
R461 VDD.n1513 VDD.n1512 10.7223
R462 VDD.n1446 VDD.n1445 10.7223
R463 VDD.n561 VDD.n560 10.7223
R464 VDD.n540 VDD.n539 10.7223
R465 VDD.n1467 VDD.n1466 10.7223
R466 VDD.n1765 VDD.n1739 10.4784
R467 VDD.n1134 VDD.n658 10.4784
R468 VDD.n1815 VDD.n1744 10.3407
R469 VDD.n1130 VDD.n652 10.3407
R470 VDD.n1638 VDD.n1637 10.2548
R471 VDD.n1338 VDD.n1337 10.2548
R472 VDD.n1126 VDD.n663 10.2279
R473 VDD.n1788 VDD.n1747 10.1865
R474 VDD.n1126 VDD.n1125 10.1865
R475 VDD.n1672 VDD.t19 9.99217
R476 VDD.n1229 VDD.t368 9.99217
R477 VDD.n592 VDD.t28 9.99217
R478 VDD.n1811 VDD.n1744 9.86137
R479 VDD.n1130 VDD.n659 9.86137
R480 VDD.n1628 VDD.n373 9.78981
R481 VDD.n1377 VDD.n588 9.78981
R482 VDD.n1932 VDD.n1931 9.6468
R483 VDD.n1846 VDD.t193 9.57585
R484 VDD.n677 VDD.t12 9.55982
R485 VDD.n673 VDD.t73 9.55982
R486 VDD.n669 VDD.t60 9.55982
R487 VDD.n665 VDD.t62 9.55982
R488 VDD.n1767 VDD.t68 9.51591
R489 VDD.n1761 VDD.t36 9.51591
R490 VDD.n1754 VDD.t41 9.51591
R491 VDD.n1786 VDD.t24 9.51591
R492 VDD.n43 VDD.n42 9.4133
R493 VDD.n1818 VDD.n1739 9.28471
R494 VDD.n1134 VDD.n656 9.28471
R495 VDD.n1673 VDD.n371 9.24507
R496 VDD.n1289 VDD.n587 9.17659
R497 VDD.n1023 VDD.n1020 9.16567
R498 VDD.n2 VDD.n1 9.09976
R499 VDD.n580 VDD.n579 9.08576
R500 VDD.n6 VDD.t598 9.02932
R501 VDD.n1663 VDD.n1662 9.01945
R502 VDD.n833 VDD.n832 8.89243
R503 VDD.n45 VDD.n44 8.82188
R504 VDD.n1571 VDD.n433 8.80618
R505 VDD.n43 VDD.t540 8.79795
R506 VDD.n1656 VDD.n389 8.78029
R507 VDD.n1651 VDD.n1650 8.78029
R508 VDD.n1325 VDD.n1324 8.78029
R509 VDD.n1322 VDD.n1311 8.78029
R510 VDD.n1646 VDD.n1645 8.71327
R511 VDD.n1633 VDD.n1632 8.71327
R512 VDD.n1343 VDD.n1342 8.71327
R513 VDD.n1330 VDD.n1329 8.71327
R514 VDD.n6 VDD.t597 8.6005
R515 VDD.n7 VDD.t595 8.6005
R516 VDD.n8 VDD.t596 8.6005
R517 VDD.n1604 VDD.n427 8.59141
R518 VDD.n1608 VDD.n427 8.59141
R519 VDD.n1610 VDD.n1608 8.59141
R520 VDD.n1612 VDD.n1610 8.59141
R521 VDD.n1612 VDD.n423 8.59141
R522 VDD.n1617 VDD.n423 8.59141
R523 VDD.n1565 VDD.n1556 8.59141
R524 VDD.n1565 VDD.n1558 8.59141
R525 VDD.n1558 VDD.n418 8.59141
R526 VDD.n1622 VDD.n418 8.59141
R527 VDD.n1623 VDD.n1622 8.59141
R528 VDD.n1371 VDD.n1349 8.59141
R529 VDD.n1366 VDD.n1349 8.59141
R530 VDD.n1366 VDD.n1354 8.59141
R531 VDD.n1362 VDD.n1354 8.59141
R532 VDD.n1362 VDD.n1357 8.59141
R533 VDD.n1389 VDD.n573 8.59141
R534 VDD.n1398 VDD.n573 8.59141
R535 VDD.n1398 VDD.n571 8.59141
R536 VDD.n571 VDD.n569 8.59141
R537 VDD.n1404 VDD.n569 8.59141
R538 VDD.n1405 VDD.n1404 8.59141
R539 VDD.n1534 VDD.n1489 8.488
R540 VDD.n1538 VDD.n447 8.488
R541 VDD.n1542 VDD.n445 8.488
R542 VDD.n1525 VDD.n1498 8.488
R543 VDD.n1501 VDD.n1500 8.488
R544 VDD.n1520 VDD.n1508 8.488
R545 VDD.n1516 VDD.n1510 8.488
R546 VDD.n1447 VDD.n474 8.488
R547 VDD.n1452 VDD.n472 8.488
R548 VDD.n1456 VDD.n465 8.488
R549 VDD.n1459 VDD.n463 8.488
R550 VDD.n558 VDD.n492 8.488
R551 VDD.n554 VDD.n494 8.488
R552 VDD.n550 VDD.n501 8.488
R553 VDD.n546 VDD.n503 8.488
R554 VDD.n538 VDD.n537 8.488
R555 VDD.n533 VDD.n509 8.488
R556 VDD.n519 VDD.n512 8.488
R557 VDD.n528 VDD.n521 8.488
R558 VDD.n818 VDD.n817 8.488
R559 VDD.n809 VDD.n755 8.488
R560 VDD.n834 VDD.n690 8.488
R561 VDD.n821 VDD.n691 8.488
R562 VDD.n814 VDD.n738 8.488
R563 VDD.n806 VDD.n758 8.488
R564 VDD.n949 VDD.n948 8.488
R565 VDD.n958 VDD.n941 8.488
R566 VDD.n962 VDD.n939 8.488
R567 VDD.n967 VDD.n937 8.488
R568 VDD.n893 VDD.n892 8.488
R569 VDD.n909 VDD.n875 8.488
R570 VDD.n910 VDD.n871 8.488
R571 VDD.n916 VDD.n868 8.488
R572 VDD.n890 VDD.n877 8.488
R573 VDD.n896 VDD.n872 8.488
R574 VDD.n913 VDD.n912 8.488
R575 VDD.n919 VDD.n869 8.488
R576 VDD.n1058 VDD.n1042 8.488
R577 VDD.n1057 VDD.n1050 8.488
R578 VDD.n1469 VDD.n1468 8.488
R579 VDD.n1481 VDD.n456 8.488
R580 VDD.n1480 VDD.n1473 8.488
R581 VDD.n1568 VDD.n1567 8.48682
R582 VDD.n1627 VDD.n413 8.48682
R583 VDD.n1373 VDD.n1372 8.48682
R584 VDD.n1356 VDD.n477 8.48682
R585 VDD.n1062 VDD.n1040 8.4005
R586 VDD.n1574 VDD.n433 8.37664
R587 VDD.n1798 VDD.n1742 8.32689
R588 VDD.n1133 VDD.n1131 8.32689
R589 VDD.n1605 VDD.n429 8.31689
R590 VDD.n1408 VDD.n567 8.31615
R591 VDD.n1534 VDD.n1490 8.2255
R592 VDD.n1538 VDD.n1489 8.2255
R593 VDD.n1542 VDD.n447 8.2255
R594 VDD.n1546 VDD.n445 8.2255
R595 VDD.n1528 VDD.n1498 8.2255
R596 VDD.n1525 VDD.n1500 8.2255
R597 VDD.n1520 VDD.n1501 8.2255
R598 VDD.n1516 VDD.n1508 8.2255
R599 VDD.n1452 VDD.n474 8.2255
R600 VDD.n1456 VDD.n472 8.2255
R601 VDD.n1459 VDD.n465 8.2255
R602 VDD.n1462 VDD.n463 8.2255
R603 VDD.n558 VDD.n494 8.2255
R604 VDD.n554 VDD.n501 8.2255
R605 VDD.n550 VDD.n503 8.2255
R606 VDD.n546 VDD.n544 8.2255
R607 VDD.n537 VDD.n509 8.2255
R608 VDD.n533 VDD.n512 8.2255
R609 VDD.n528 VDD.n519 8.2255
R610 VDD.n525 VDD.n521 8.2255
R611 VDD.n817 VDD.n755 8.2255
R612 VDD.n809 VDD.n760 8.2255
R613 VDD.n710 VDD.n690 8.2255
R614 VDD.n834 VDD.n691 8.2255
R615 VDD.n821 VDD.n738 8.2255
R616 VDD.n814 VDD.n758 8.2255
R617 VDD.n806 VDD.n763 8.2255
R618 VDD.n958 VDD.n948 8.2255
R619 VDD.n962 VDD.n941 8.2255
R620 VDD.n967 VDD.n939 8.2255
R621 VDD.n892 VDD.n879 8.2255
R622 VDD.n893 VDD.n875 8.2255
R623 VDD.n910 VDD.n909 8.2255
R624 VDD.n916 VDD.n871 8.2255
R625 VDD.n922 VDD.n868 8.2255
R626 VDD.n890 VDD.n889 8.2255
R627 VDD.n896 VDD.n877 8.2255
R628 VDD.n912 VDD.n872 8.2255
R629 VDD.n913 VDD.n869 8.2255
R630 VDD.n919 VDD.n867 8.2255
R631 VDD.n1062 VDD.n1042 8.2255
R632 VDD.n1058 VDD.n1057 8.2255
R633 VDD.n1054 VDD.n1050 8.2255
R634 VDD.n1469 VDD.n455 8.2255
R635 VDD.n1485 VDD.n456 8.2255
R636 VDD.n1481 VDD.n1480 8.2255
R637 VDD.n1476 VDD.n1473 8.2255
R638 VDD.n1985 VDD.n1983 8.2255
R639 VDD.n747 VDD.n739 8.20843
R640 VDD.n1030 VDD.n1029 8.20843
R641 VDD.n1677 VDD.n371 8.14941
R642 VDD.n1677 VDD.n364 8.14941
R643 VDD.n1687 VDD.n364 8.14941
R644 VDD.n1687 VDD.n342 8.14941
R645 VDD.n1703 VDD.n342 8.14941
R646 VDD.n1703 VDD.n343 8.14941
R647 VDD.n1699 VDD.n343 8.14941
R648 VDD.n1699 VDD.n276 8.14941
R649 VDD.n1859 VDD.n276 8.14941
R650 VDD.n1859 VDD.n277 8.14941
R651 VDD.n1855 VDD.n277 8.14941
R652 VDD.n1855 VDD.n280 8.14941
R653 VDD.n292 VDD.n280 8.14941
R654 VDD.n1845 VDD.n292 8.14941
R655 VDD.n1845 VDD.n293 8.14941
R656 VDD.n1840 VDD.n293 8.14941
R657 VDD.n1840 VDD.n299 8.14941
R658 VDD.n312 VDD.n299 8.14941
R659 VDD.n1830 VDD.n312 8.14941
R660 VDD.n1830 VDD.n313 8.14941
R661 VDD.n1825 VDD.n313 8.14941
R662 VDD.n1825 VDD.n1730 8.14941
R663 VDD.n1743 VDD.n1730 8.14941
R664 VDD.n1815 VDD.n1743 8.14941
R665 VDD.n1141 VDD.n652 8.14941
R666 VDD.n1141 VDD.n650 8.14941
R667 VDD.n1145 VDD.n650 8.14941
R668 VDD.n1145 VDD.n639 8.14941
R669 VDD.n1158 VDD.n639 8.14941
R670 VDD.n1158 VDD.n640 8.14941
R671 VDD.n640 VDD.n630 8.14941
R672 VDD.n1223 VDD.n630 8.14941
R673 VDD.n1223 VDD.n625 8.14941
R674 VDD.n1228 VDD.n625 8.14941
R675 VDD.n1228 VDD.n619 8.14941
R676 VDD.n1239 VDD.n619 8.14941
R677 VDD.n1239 VDD.n617 8.14941
R678 VDD.n1244 VDD.n617 8.14941
R679 VDD.n1244 VDD.n609 8.14941
R680 VDD.n1256 VDD.n609 8.14941
R681 VDD.n1256 VDD.n607 8.14941
R682 VDD.n1261 VDD.n607 8.14941
R683 VDD.n1261 VDD.n599 8.14941
R684 VDD.n1273 VDD.n599 8.14941
R685 VDD.n1273 VDD.n597 8.14941
R686 VDD.n1277 VDD.n597 8.14941
R687 VDD.n1277 VDD.n590 8.14941
R688 VDD.n1289 VDD.n590 8.14941
R689 VDD.n831 VDD.n720 7.963
R690 VDD.n1832 VDD.t185 7.91057
R691 VDD.n1680 VDD.n368 7.89208
R692 VDD.n1680 VDD.n366 7.89208
R693 VDD.n1684 VDD.n366 7.89208
R694 VDD.n1684 VDD.n339 7.89208
R695 VDD.n1706 VDD.n339 7.89208
R696 VDD.n1706 VDD.n340 7.89208
R697 VDD.n1695 VDD.n340 7.89208
R698 VDD.n1695 VDD.n273 7.89208
R699 VDD.n1862 VDD.n273 7.89208
R700 VDD.n1862 VDD.n274 7.89208
R701 VDD.n285 VDD.n274 7.89208
R702 VDD.n1852 VDD.n285 7.89208
R703 VDD.n1852 VDD.n286 7.89208
R704 VDD.n1848 VDD.n286 7.89208
R705 VDD.n1848 VDD.n289 7.89208
R706 VDD.n304 VDD.n289 7.89208
R707 VDD.n1837 VDD.n304 7.89208
R708 VDD.n1837 VDD.n305 7.89208
R709 VDD.n1833 VDD.n305 7.89208
R710 VDD.n1833 VDD.n308 7.89208
R711 VDD.n1734 VDD.n308 7.89208
R712 VDD.n1822 VDD.n1734 7.89208
R713 VDD.n1822 VDD.n1735 7.89208
R714 VDD.n1818 VDD.n1735 7.89208
R715 VDD.n1138 VDD.n656 7.89208
R716 VDD.n1138 VDD.n649 7.89208
R717 VDD.n1149 VDD.n649 7.89208
R718 VDD.n1149 VDD.n642 7.89208
R719 VDD.n1155 VDD.n642 7.89208
R720 VDD.n1155 VDD.n647 7.89208
R721 VDD.n647 VDD.n633 7.89208
R722 VDD.n1220 VDD.n633 7.89208
R723 VDD.n1220 VDD.n624 7.89208
R724 VDD.n1232 VDD.n624 7.89208
R725 VDD.n1232 VDD.n622 7.89208
R726 VDD.n1236 VDD.n622 7.89208
R727 VDD.n1236 VDD.n615 7.89208
R728 VDD.n1248 VDD.n615 7.89208
R729 VDD.n1248 VDD.n612 7.89208
R730 VDD.n1253 VDD.n612 7.89208
R731 VDD.n1253 VDD.n605 7.89208
R732 VDD.n1265 VDD.n605 7.89208
R733 VDD.n1265 VDD.n602 7.89208
R734 VDD.n1270 VDD.n602 7.89208
R735 VDD.n1270 VDD.n595 7.89208
R736 VDD.n1281 VDD.n595 7.89208
R737 VDD.n1281 VDD.n593 7.89208
R738 VDD.n1286 VDD.n593 7.89208
R739 VDD.n714 VDD.n701 7.613
R740 VDD.n55 VDD.t541 7.58462
R741 VDD.n56 VDD.t144 7.58462
R742 VDD.n37 VDD.n23 7.58109
R743 VDD.n1078 VDD.n1018 7.5255
R744 VDD.n748 VDD.n747 7.52444
R745 VDD.n1156 VDD.t372 7.49426
R746 VDD.n1642 VDD.n1641 7.30582
R747 VDD.n1334 VDD.n1333 7.30582
R748 VDD.n1382 VDD.n584 7.30582
R749 VDD.n26 VDD.t139 7.19043
R750 VDD.n3 VDD.t599 7.19043
R751 VDD.n818 VDD.n754 7.1755
R752 VDD.n971 VDD.n937 7.1755
R753 VDD.n720 VDD.n719 7.088
R754 VDD.n1771 VDD.n1763 7.00704
R755 VDD.n1775 VDD.n1763 7.00704
R756 VDD.n1776 VDD.n1775 7.00704
R757 VDD.n1777 VDD.n1776 7.00704
R758 VDD.n1777 VDD.n1760 7.00704
R759 VDD.n1782 VDD.n1760 7.00704
R760 VDD.n1782 VDD.n1751 7.00704
R761 VDD.n1805 VDD.n1751 7.00704
R762 VDD.n1805 VDD.n1752 7.00704
R763 VDD.n1800 VDD.n1752 7.00704
R764 VDD.n1800 VDD.n1756 7.00704
R765 VDD.n1795 VDD.n1756 7.00704
R766 VDD.n1795 VDD.n1785 7.00704
R767 VDD.n1790 VDD.n1785 7.00704
R768 VDD.n1790 VDD.n1788 7.00704
R769 VDD.n1123 VDD.n664 7.00704
R770 VDD.n1118 VDD.n1117 7.00704
R771 VDD.n1115 VDD.n668 7.00704
R772 VDD.n1110 VDD.n1109 7.00704
R773 VDD.n1107 VDD.n672 7.00704
R774 VDD.n1102 VDD.n1101 7.00704
R775 VDD.n1099 VDD.n676 7.00704
R776 VDD.n122 VDD.t530 6.94485
R777 VDD.n220 VDD.t721 6.94485
R778 VDD.n409 VDD.n407 6.94485
R779 VDD.n1295 VDD.t785 6.94485
R780 VDD.t688 VDD.n717 6.84045
R781 VDD.n808 VDD.t677 6.84045
R782 VDD.t350 VDD.n878 6.84045
R783 VDD.n1077 VDD.n1076 6.84045
R784 VDD.n1496 VDD.n1495 6.70224
R785 VDD.n1493 VDD.n1491 6.70224
R786 VDD.n523 VDD.t662 6.70224
R787 VDD.n504 VDD.t790 6.70224
R788 VDD.n765 VDD.t766 6.70224
R789 VDD.n704 VDD.n703 6.70224
R790 VDD.n934 VDD.t443 6.70224
R791 VDD.n882 VDD.n880 6.70224
R792 VDD.n885 VDD.n884 6.70224
R793 VDD.n1052 VDD.t459 6.70224
R794 VDD.n461 VDD.t381 6.70224
R795 VDD.n1474 VDD.t494 6.70224
R796 VDD.n1990 VDD.n1989 6.70224
R797 VDD.n443 VDD.t648 6.68489
R798 VDD.n564 VDD.n562 6.68371
R799 VDD.n173 VDD.t504 6.68267
R800 VDD.n1511 VDD.t174 6.65503
R801 VDD.n507 VDD.n505 6.65503
R802 VDD.n793 VDD.t681 6.65503
R803 VDD.n707 VDD.n705 6.65503
R804 VDD.n952 VDD.n950 6.65503
R805 VDD.n849 VDD.t433 6.65503
R806 VDD.n1026 VDD.n1024 6.65503
R807 VDD.n1444 VDD.n1443 6.65503
R808 VDD.n460 VDD.n459 6.65503
R809 VDD.n1965 VDD.t719 6.65503
R810 VDD.n927 VDD.t354 6.64521
R811 VDD.n1661 VDD.n1660 6.63561
R812 VDD.n1917 VDD.n1916 6.61305
R813 VDD.n178 VDD.n177 6.58706
R814 VDD.n1382 VDD.n1381 6.56859
R815 VDD.n1915 VDD.t463 6.54616
R816 VDD.n1915 VDD.t467 6.54616
R817 VDD.n201 VDD.t241 6.52811
R818 VDD.n181 VDD.n180 6.52199
R819 VDD.n1918 VDD.n1913 6.51831
R820 VDD.t35 VDD.n1350 6.50716
R821 VDD.n415 VDD.t45 6.50716
R822 VDD.t340 VDD.n1922 6.47299
R823 VDD.n151 VDD.t273 6.47299
R824 VDD.n250 VDD.t230 6.47299
R825 VDD.n1908 VDD.t570 6.47299
R826 VDD.n51 VDD.n50 6.44895
R827 VDD.n1308 VDD.t15 6.43191
R828 VDD.n1294 VDD.t55 6.43124
R829 VDD.n1317 VDD.t27 6.4298
R830 VDD.n390 VDD.t18 6.42961
R831 VDD.n398 VDD.t75 6.37351
R832 VDD.n1298 VDD.t70 6.37275
R833 VDD.n405 VDD.t30 6.37256
R834 VDD.n411 VDD.t39 6.37217
R835 VDD.n425 VDD.t52 6.36486
R836 VDD.n1600 VDD.t65 6.36262
R837 VDD.n1560 VDD.t49 6.36128
R838 VDD.n1393 VDD.t46 6.30795
R839 VDD.n574 VDD.t57 6.30193
R840 VDD.n83 VDD.n82 6.3005
R841 VDD.n143 VDD.n142 6.3005
R842 VDD VDD.n151 6.3005
R843 VDD.n157 VDD.n132 6.3005
R844 VDD.n161 VDD.n124 6.3005
R845 VDD.n97 VDD.n96 6.3005
R846 VDD.n242 VDD.n241 6.3005
R847 VDD.n204 VDD.n203 6.3005
R848 VDD VDD.n205 6.3005
R849 VDD.n260 VDD.n223 6.3005
R850 VDD.n256 VDD.n231 6.3005
R851 VDD VDD.n250 6.3005
R852 VDD.n1900 VDD.n1899 6.3005
R853 VDD.n744 VDD.n743 6.3005
R854 VDD.n745 VDD.n744 6.3005
R855 VDD.n750 VDD.n749 6.3005
R856 VDD.n749 VDD.n748 6.3005
R857 VDD.n714 VDD.n713 6.3005
R858 VDD.n715 VDD.n714 6.3005
R859 VDD.n971 VDD.n970 6.3005
R860 VDD.n972 VDD.n971 6.3005
R861 VDD.n1022 VDD.n1021 6.3005
R862 VDD.n1040 VDD.n1039 6.3005
R863 VDD.n1064 VDD.n1040 6.3005
R864 VDD.n1079 VDD.n1078 6.3005
R865 VDD.n1078 VDD.n1077 6.3005
R866 VDD.n1019 VDD.n1017 6.3005
R867 VDD.n1076 VDD.n1019 6.3005
R868 VDD.n1067 VDD.n1066 6.3005
R869 VDD.n1066 VDD.n1065 6.3005
R870 VDD VDD.n1908 6.3005
R871 VDD.n1897 VDD.n1896 6.3005
R872 VDD.n1907 VDD.n1906 6.3005
R873 VDD.n1922 VDD 6.3005
R874 VDD.n73 VDD.n72 6.3005
R875 VDD.n1926 VDD.n1923 6.3005
R876 VDD.n10 VDD.n5 6.3005
R877 VDD.n11 VDD.n4 6.3005
R878 VDD.n12 VDD.n3 6.3005
R879 VDD.n14 VDD.n13 6.3005
R880 VDD.n30 VDD.n29 6.3005
R881 VDD.n31 VDD.n28 6.3005
R882 VDD.n32 VDD.n27 6.3005
R883 VDD.n33 VDD.n26 6.3005
R884 VDD.n34 VDD.n25 6.3005
R885 VDD.n35 VDD.n24 6.3005
R886 VDD.n1950 VDD.n1940 6.3005
R887 VDD VDD.n1941 6.3005
R888 VDD.n1949 VDD.n1942 6.3005
R889 VDD.n2004 VDD.n2003 6.3005
R890 VDD.n2006 VDD.n2005 6.3005
R891 VDD.n2008 VDD.n2007 6.3005
R892 VDD.n1358 VDD.t21 6.29942
R893 VDD.n415 VDD.t43 6.29685
R894 VDD.n46 VDD.t140 6.27989
R895 VDD.n927 VDD.t357 6.26273
R896 VDD.n564 VDD.n563 6.24167
R897 VDD.n122 VDD.t313 6.2405
R898 VDD.n220 VDD.t737 6.2405
R899 VDD.n409 VDD.n408 6.2405
R900 VDD.n443 VDD.t615 6.2405
R901 VDD.n1511 VDD.t199 6.2405
R902 VDD.n1496 VDD.n1494 6.2405
R903 VDD.n1493 VDD.n1492 6.2405
R904 VDD.n1351 VDD.t35 6.2405
R905 VDD.n1295 VDD.t767 6.2405
R906 VDD.n523 VDD.t661 6.2405
R907 VDD.n507 VDD.n506 6.2405
R908 VDD.n504 VDD.t820 6.2405
R909 VDD.n765 VDD.t751 6.2405
R910 VDD.n793 VDD.t678 6.2405
R911 VDD.n707 VDD.n706 6.2405
R912 VDD.n704 VDD.n702 6.2405
R913 VDD.n952 VDD.n951 6.2405
R914 VDD.n934 VDD.t428 6.2405
R915 VDD.n885 VDD.n883 6.2405
R916 VDD.n882 VDD.n881 6.2405
R917 VDD.n849 VDD.t439 6.2405
R918 VDD.n1052 VDD.t455 6.2405
R919 VDD.n1026 VDD.n1025 6.2405
R920 VDD.n1444 VDD.n1442 6.2405
R921 VDD.n461 VDD.t410 6.2405
R922 VDD.n460 VDD.n458 6.2405
R923 VDD.n1474 VDD.t490 6.2405
R924 VDD.t45 VDD.n414 6.2405
R925 VDD.n1965 VDD.t714 6.2405
R926 VDD.n1990 VDD.n1988 6.2405
R927 VDD.n1350 VDD.t33 6.23498
R928 VDD.n715 VDD.n700 6.15645
R929 VDD.n1381 VDD.n579 6.03524
R930 VDD.n254 VDD.n244 6.01865
R931 VDD.n1904 VDD.n1902 6.01865
R932 VDD.n80 VDD.n60 6.01863
R933 VDD.n155 VDD.n145 6.01863
R934 VDD.n1662 VDD.n1661 5.96892
R935 VDD.n786 VDD.n785 5.77744
R936 VDD.n775 VDD.n774 5.77744
R937 VDD.n991 VDD.t582 5.77744
R938 VDD.n986 VDD.t757 5.77744
R939 VDD.n1946 VDD.n1945 5.77744
R940 VDD.n1999 VDD.t249 5.77744
R941 VDD.n749 VDD.n744 5.7755
R942 VDD.n20 VDD.n19 5.7405
R943 VDD.n974 VDD.n973 5.2962
R944 VDD.n226 VDD.t651 5.20342
R945 VDD.n1891 VDD.t288 5.20342
R946 VDD.n67 VDD.t265 5.20242
R947 VDD.n127 VDD.t554 5.20242
R948 VDD.n22 VDD.n16 5.2005
R949 VDD.n21 VDD.n17 5.2005
R950 VDD.n20 VDD.n18 5.2005
R951 VDD.n64 VDD.t214 5.17246
R952 VDD.n123 VDD.t152 5.17246
R953 VDD.n222 VDD.t82 5.17246
R954 VDD.n1888 VDD.t8 5.17246
R955 VDD.n77 VDD.n76 5.107
R956 VDD.n140 VDD.n139 5.107
R957 VDD.n239 VDD.n238 5.107
R958 VDD.n1887 VDD.n1886 5.107
R959 VDD.n1661 VDD.n375 5.10682
R960 VDD.n1381 VDD.n1380 5.10682
R961 VDD.n776 VDD.t761 5.07264
R962 VDD.n993 VDD.n992 5.07264
R963 VDD.n988 VDD.n987 5.07264
R964 VDD.n1947 VDD.t715 5.07264
R965 VDD.n2001 VDD.n2000 5.07264
R966 VDD.n179 VDD.n93 5.0405
R967 VDD.n1808 VDD.t25 4.99634
R968 VDD.n152 VDD.t272 4.92985
R969 VDD.n251 VDD.t133 4.92985
R970 VDD.n267 VDD.t488 4.92985
R971 VDD.n92 VDD.t335 4.92985
R972 VDD.n790 VDD.t578 4.79075
R973 VDD.n716 VDD.n715 4.78846
R974 VDD.n1074 VDD.n1032 4.7255
R975 VDD.n80 VDD.t337 4.64447
R976 VDD.n145 VDD.t280 4.64447
R977 VDD.n244 VDD.t135 4.64447
R978 VDD.n1902 VDD.t569 4.64447
R979 VDD.n70 VDD.n69 4.60311
R980 VDD.n154 VDD.t775 4.60311
R981 VDD.n159 VDD.n129 4.60311
R982 VDD.n258 VDD.n228 4.60311
R983 VDD.n253 VDD.t416 4.60311
R984 VDD.n1894 VDD.n1893 4.60311
R985 VDD.n1903 VDD.t115 4.60311
R986 VDD.n90 VDD.t524 4.60311
R987 VDD.n801 VDD.n768 4.52789
R988 VDD.n1070 VDD.n1069 4.52785
R989 VDD.n699 VDD.n684 4.51855
R990 VDD.n974 VDD.n933 4.5152
R991 VDD.n825 VDD.n824 4.5084
R992 VDD.n863 VDD.n862 4.50489
R993 VDD.n800 VDD.n799 4.5005
R994 VDD.n798 VDD.n769 4.5005
R995 VDD.n794 VDD.n767 4.5005
R996 VDD.n768 VDD.n759 4.5005
R997 VDD.n804 VDD.n764 4.5005
R998 VDD.n753 VDD.n752 4.5005
R999 VDD.n754 VDD.n753 4.5005
R1000 VDD.n754 VDD.n739 4.5005
R1001 VDD.n837 VDD.n836 4.5005
R1002 VDD.n830 VDD.n829 4.5005
R1003 VDD.n831 VDD.n830 4.5005
R1004 VDD.n832 VDD.n831 4.5005
R1005 VDD.n719 VDD.n699 4.5005
R1006 VDD.n719 VDD.n718 4.5005
R1007 VDD.n696 VDD.n686 4.5005
R1008 VDD.n840 VDD.n839 4.5005
R1009 VDD.n826 VDD.n723 4.5005
R1010 VDD.n828 VDD.n827 4.5005
R1011 VDD.n838 VDD.n685 4.5005
R1012 VDD.n978 VDD.n932 4.5005
R1013 VDD.n979 VDD.n931 4.5005
R1014 VDD.n863 VDD.n852 4.5005
R1015 VDD.n866 VDD.n853 4.5005
R1016 VDD.n924 VDD.n923 4.5005
R1017 VDD.n925 VDD.n924 4.5005
R1018 VDD.n866 VDD.n865 4.5005
R1019 VDD.n859 VDD.n854 4.5005
R1020 VDD.n856 VDD.n855 4.5005
R1021 VDD.n847 VDD.n846 4.5005
R1022 VDD.n861 VDD.n860 4.5005
R1023 VDD.n1011 VDD.n1010 4.5005
R1024 VDD.n1005 VDD.n1004 4.5005
R1025 VDD.n1006 VDD.n844 4.5005
R1026 VDD.n1009 VDD.n843 4.5005
R1027 VDD.n1069 VDD.n1068 4.5005
R1028 VDD.n1068 VDD.n1032 4.5005
R1029 VDD.n1032 VDD.n1031 4.5005
R1030 VDD.n1038 VDD.n1035 4.5005
R1031 VDD.n1073 VDD.n1072 4.5005
R1032 VDD.n1074 VDD.n1073 4.5005
R1033 VDD.n1075 VDD.n1074 4.5005
R1034 VDD.n1037 VDD.n1034 4.5005
R1035 VDD.n1036 VDD.n1015 4.5005
R1036 VDD.n1081 VDD.n1080 4.5005
R1037 VDD.n1085 VDD.n1084 4.5005
R1038 VDD.n1022 VDD.n682 4.5005
R1039 VDD.n1022 VDD.n1018 4.5005
R1040 VDD.n1030 VDD.n1018 4.5005
R1041 VDD.n683 VDD.n681 4.5005
R1042 VDD.n1869 VDD.n1868 4.5005
R1043 VDD.n54 VDD.n53 4.5005
R1044 VDD.n64 VDD.t215 4.2255
R1045 VDD.n152 VDD.t276 4.2255
R1046 VDD.n123 VDD.t151 4.2255
R1047 VDD.n222 VDD.t787 4.2255
R1048 VDD.n251 VDD.t236 4.2255
R1049 VDD.n1888 VDD.t417 4.2255
R1050 VDD.n267 VDD.t575 4.2255
R1051 VDD.n92 VDD.t339 4.2255
R1052 VDD.n1537 VDD.t618 4.10447
R1053 VDD.t183 VDD.n1499 4.10447
R1054 VDD.t386 VDD.n464 4.10447
R1055 VDD.t811 VDD.n551 4.10447
R1056 VDD.n522 VDD.t657 4.10447
R1057 VDD.n964 VDD.t429 4.10447
R1058 VDD.n1049 VDD.t451 4.10447
R1059 VDD.t491 VDD.n1482 4.10447
R1060 VDD.n1975 VDD.t711 4.10447
R1061 VDD.n190 VDD.n189 3.99669
R1062 VDD.n102 VDD.n101 3.99665
R1063 VDD.n189 VDD.t650 3.80383
R1064 VDD.n101 VDD.t469 3.80304
R1065 VDD.n1671 VDD.n369 3.74738
R1066 VDD.n1679 VDD.n1678 3.74738
R1067 VDD.n370 VDD.n365 3.74738
R1068 VDD.t168 VDD.n1685 3.74738
R1069 VDD.n1686 VDD.n341 3.74738
R1070 VDD.n1705 VDD.n1704 3.74738
R1071 VDD.n1693 VDD.n1692 3.74738
R1072 VDD.n1698 VDD.n1696 3.74738
R1073 VDD.n1697 VDD.n275 3.74738
R1074 VDD.n1861 VDD.n1860 3.74738
R1075 VDD.n282 VDD.n281 3.74738
R1076 VDD.n1854 VDD.n283 3.74738
R1077 VDD.n1853 VDD.n284 3.74738
R1078 VDD.n291 VDD.n290 3.74738
R1079 VDD.n1847 VDD.n1846 3.74738
R1080 VDD.n301 VDD.n300 3.74738
R1081 VDD.n1839 VDD.n302 3.74738
R1082 VDD.n1838 VDD.n303 3.74738
R1083 VDD.n311 VDD.n310 3.74738
R1084 VDD.n1832 VDD.n1831 3.74738
R1085 VDD.n1731 VDD.n309 3.74738
R1086 VDD.n1824 VDD.n1732 3.74738
R1087 VDD.n1823 VDD.n1733 3.74738
R1088 VDD.n1741 VDD.n1740 3.74738
R1089 VDD.n1817 VDD.n1816 3.74738
R1090 VDD.n1132 VDD.n653 3.74738
R1091 VDD.n1140 VDD.n1139 3.74738
R1092 VDD.n655 VDD.n654 3.74738
R1093 VDD.n1148 VDD.n1146 3.74738
R1094 VDD.n1147 VDD.n641 3.74738
R1095 VDD.n1157 VDD.n1156 3.74738
R1096 VDD.n646 VDD.n643 3.74738
R1097 VDD.n645 VDD.n644 3.74738
R1098 VDD.n1222 VDD.n1221 3.74738
R1099 VDD.n632 VDD.n631 3.74738
R1100 VDD.n1231 VDD.n1229 3.74738
R1101 VDD.n1230 VDD.n620 3.74738
R1102 VDD.n1238 VDD.n1237 3.74738
R1103 VDD.n621 VDD.n616 3.74738
R1104 VDD.n1247 VDD.n1245 3.74738
R1105 VDD.n1246 VDD.n610 3.74738
R1106 VDD.n1255 VDD.n1254 3.74738
R1107 VDD.n611 VDD.n606 3.74738
R1108 VDD.n1264 VDD.n1262 3.74738
R1109 VDD.n1263 VDD.n600 3.74738
R1110 VDD.n1272 VDD.n1271 3.74738
R1111 VDD.n601 VDD.n596 3.74738
R1112 VDD.n1280 VDD.n1278 3.74738
R1113 VDD.n1279 VDD.n591 3.74738
R1114 VDD.n1288 VDD.n1287 3.74738
R1115 VDD.n111 VDD.t311 3.6405
R1116 VDD.n111 VDD.n110 3.6405
R1117 VDD.n113 VDD.t226 3.6405
R1118 VDD.n113 VDD.n112 3.6405
R1119 VDD.n115 VDD.t224 3.6405
R1120 VDD.n115 VDD.n114 3.6405
R1121 VDD.n117 VDD.t786 3.6405
R1122 VDD.n117 VDD.n116 3.6405
R1123 VDD.n109 VDD.t310 3.6405
R1124 VDD.n109 VDD.n108 3.6405
R1125 VDD.n106 VDD.t309 3.6405
R1126 VDD.n106 VDD.n105 3.6405
R1127 VDD.n104 VDD.t315 3.6405
R1128 VDD.n104 VDD.n103 3.6405
R1129 VDD.n99 VDD.t317 3.6405
R1130 VDD.n99 VDD.n98 3.6405
R1131 VDD.n95 VDD.t514 3.6405
R1132 VDD.n95 VDD.n94 3.6405
R1133 VDD.n200 VDD.t664 3.6405
R1134 VDD.n200 VDD.n199 3.6405
R1135 VDD.n187 VDD.t243 3.6405
R1136 VDD.n187 VDD.n186 3.6405
R1137 VDD.n185 VDD.t127 3.6405
R1138 VDD.n185 VDD.n184 3.6405
R1139 VDD.n197 VDD.t129 3.6405
R1140 VDD.n197 VDD.n196 3.6405
R1141 VDD.n195 VDD.t245 3.6405
R1142 VDD.n195 VDD.n194 3.6405
R1143 VDD.n217 VDD.t131 3.6405
R1144 VDD.n217 VDD.n216 3.6405
R1145 VDD.n209 VDD.t478 3.6405
R1146 VDD.n209 VDD.n208 3.6405
R1147 VDD.n213 VDD.t474 3.6405
R1148 VDD.n213 VDD.n212 3.6405
R1149 VDD.n211 VDD.t466 3.6405
R1150 VDD.n211 VDD.n210 3.6405
R1151 VDD.n1711 VDD.t629 3.6405
R1152 VDD.n1711 VDD.n1710 3.6405
R1153 VDD.n348 VDD.t611 3.6405
R1154 VDD.n348 VDD.n347 3.6405
R1155 VDD.n332 VDD.t628 3.6405
R1156 VDD.n332 VDD.n331 3.6405
R1157 VDD.n329 VDD.t161 3.6405
R1158 VDD.n329 VDD.n328 3.6405
R1159 VDD.n326 VDD.t622 3.6405
R1160 VDD.n326 VDD.n325 3.6405
R1161 VDD.n354 VDD.t642 3.6405
R1162 VDD.n354 VDD.n353 3.6405
R1163 VDD.n1723 VDD.t207 3.6405
R1164 VDD.n1723 VDD.n1722 3.6405
R1165 VDD.n1720 VDD.t186 3.6405
R1166 VDD.n1720 VDD.n1719 3.6405
R1167 VDD.n317 VDD.t643 3.6405
R1168 VDD.n317 VDD.n316 3.6405
R1169 VDD.n396 VDD.t93 3.6405
R1170 VDD.n396 VDD.n395 3.6405
R1171 VDD.n394 VDD.t94 3.6405
R1172 VDD.n394 VDD.n393 3.6405
R1173 VDD.n402 VDD.t783 3.6405
R1174 VDD.n402 VDD.n401 3.6405
R1175 VDD.n400 VDD.t784 3.6405
R1176 VDD.n400 VDD.n399 3.6405
R1177 VDD.n1551 VDD.t624 3.6405
R1178 VDD.n1551 VDD.n1550 3.6405
R1179 VDD.n1549 VDD.t619 3.6405
R1180 VDD.n1549 VDD.n1548 3.6405
R1181 VDD.n1503 VDD.t206 3.6405
R1182 VDD.n1503 VDD.n1502 3.6405
R1183 VDD.n1505 VDD.t184 3.6405
R1184 VDD.n1505 VDD.n1504 3.6405
R1185 VDD.n1313 VDD.t119 3.6405
R1186 VDD.n1313 VDD.n1312 3.6405
R1187 VDD.n1315 VDD.t777 3.6405
R1188 VDD.n1315 VDD.n1314 3.6405
R1189 VDD.n1302 VDD.t778 3.6405
R1190 VDD.n1302 VDD.n1301 3.6405
R1191 VDD.n1304 VDD.t776 3.6405
R1192 VDD.n1304 VDD.n1303 3.6405
R1193 VDD.n1192 VDD.t788 3.6405
R1194 VDD.n1192 VDD.n1191 3.6405
R1195 VDD.n1178 VDD.t791 3.6405
R1196 VDD.n1178 VDD.n1177 3.6405
R1197 VDD.n1180 VDD.t817 3.6405
R1198 VDD.n1180 VDD.n1179 3.6405
R1199 VDD.n1186 VDD.t411 3.6405
R1200 VDD.n1186 VDD.n1185 3.6405
R1201 VDD.n1189 VDD.t397 3.6405
R1202 VDD.n1189 VDD.n1188 3.6405
R1203 VDD.n1174 VDD.t798 3.6405
R1204 VDD.n1174 VDD.n1173 3.6405
R1205 VDD.n517 VDD.t221 3.6405
R1206 VDD.n517 VDD.n516 3.6405
R1207 VDD.n515 VDD.t220 3.6405
R1208 VDD.n515 VDD.n514 3.6405
R1209 VDD.n498 VDD.t794 3.6405
R1210 VDD.n498 VDD.n497 3.6405
R1211 VDD.n496 VDD.t805 3.6405
R1212 VDD.n496 VDD.n495 3.6405
R1213 VDD.n1182 VDD.t371 3.6405
R1214 VDD.n1182 VDD.n1181 3.6405
R1215 VDD.n1215 VDD.t394 3.6405
R1216 VDD.n1215 VDD.n1214 3.6405
R1217 VDD.n1210 VDD.t814 3.6405
R1218 VDD.n1210 VDD.n1209 3.6405
R1219 VDD.n1204 VDD.t383 3.6405
R1220 VDD.n1204 VDD.n1203 3.6405
R1221 VDD.n1207 VDD.t407 3.6405
R1222 VDD.n1207 VDD.n1206 3.6405
R1223 VDD.n1162 VDD.t792 3.6405
R1224 VDD.n1162 VDD.n1161 3.6405
R1225 VDD.n1167 VDD.t823 3.6405
R1226 VDD.n1167 VDD.n1166 3.6405
R1227 VDD.n1165 VDD.t810 3.6405
R1228 VDD.n1165 VDD.n1164 3.6405
R1229 VDD.n1171 VDD.t365 3.6405
R1230 VDD.n1171 VDD.n1170 3.6405
R1231 VDD.n627 VDD.t376 3.6405
R1232 VDD.n627 VDD.n626 3.6405
R1233 VDD.n730 VDD.t754 3.6405
R1234 VDD.n730 VDD.n729 3.6405
R1235 VDD.n728 VDD.t745 3.6405
R1236 VDD.n728 VDD.n727 3.6405
R1237 VDD.n734 VDD.t680 3.6405
R1238 VDD.n734 VDD.n733 3.6405
R1239 VDD.n736 VDD.t687 3.6405
R1240 VDD.n736 VDD.n735 3.6405
R1241 VDD.n945 VDD.t426 3.6405
R1242 VDD.n945 VDD.n944 3.6405
R1243 VDD.n943 VDD.t440 3.6405
R1244 VDD.n943 VDD.n942 3.6405
R1245 VDD.n904 VDD.t356 3.6405
R1246 VDD.n904 VDD.n903 3.6405
R1247 VDD.n906 VDD.t361 3.6405
R1248 VDD.n906 VDD.n905 3.6405
R1249 VDD.n901 VDD.t438 3.6405
R1250 VDD.n901 VDD.n900 3.6405
R1251 VDD.n899 VDD.t432 3.6405
R1252 VDD.n899 VDD.n898 3.6405
R1253 VDD.n1046 VDD.t458 3.6405
R1254 VDD.n1046 VDD.n1045 3.6405
R1255 VDD.n1044 VDD.t447 3.6405
R1256 VDD.n1044 VDD.n1043 3.6405
R1257 VDD.n467 VDD.t367 3.6405
R1258 VDD.n467 VDD.n466 3.6405
R1259 VDD.n469 VDD.t395 3.6405
R1260 VDD.n469 VDD.n468 3.6405
R1261 VDD.n450 VDD.t486 3.6405
R1262 VDD.n450 VDD.n449 3.6405
R1263 VDD.n452 VDD.t483 3.6405
R1264 VDD.n452 VDD.n451 3.6405
R1265 VDD.n1727 VDD.t637 3.6405
R1266 VDD.n1727 VDD.n1726 3.6405
R1267 VDD.n296 VDD.t194 3.6405
R1268 VDD.n296 VDD.n295 3.6405
R1269 VDD.n351 VDD.t203 3.6405
R1270 VDD.n351 VDD.n350 3.6405
R1271 VDD.n361 VDD.t623 3.6405
R1272 VDD.n361 VDD.n360 3.6405
R1273 VDD.n335 VDD.t169 3.6405
R1274 VDD.n335 VDD.n334 3.6405
R1275 VDD.n345 VDD.t192 3.6405
R1276 VDD.n345 VDD.n344 3.6405
R1277 VDD.n323 VDD.t202 3.6405
R1278 VDD.n323 VDD.n322 3.6405
R1279 VDD.n1961 VDD.t712 3.6405
R1280 VDD.n1961 VDD.n1960 3.6405
R1281 VDD.n1963 VDD.t718 3.6405
R1282 VDD.n1963 VDD.n1962 3.6405
R1283 VDD.n227 VDD.n226 3.60762
R1284 VDD.n1892 VDD.n1891 3.60762
R1285 VDD.n68 VDD.n67 3.60724
R1286 VDD.n128 VDD.n127 3.60724
R1287 VDD.n118 VDD.n117 3.54622
R1288 VDD.n214 VDD.n213 3.54622
R1289 VDD.n748 VDD.t679 3.42047
R1290 VDD.n281 VDD.t162 3.33106
R1291 VDD.n1090 VDD.n1088 3.32815
R1292 VDD.n150 VDD.n149 3.30485
R1293 VDD.n249 VDD.n246 3.30485
R1294 VDD.n1875 VDD.n1872 3.30485
R1295 VDD.n397 VDD.n394 3.30485
R1296 VDD.n403 VDD.n400 3.30485
R1297 VDD.n1316 VDD.n1315 3.30485
R1298 VDD.n1305 VDD.n1304 3.30485
R1299 VDD.n89 VDD.n88 3.30485
R1300 VDD.n1345 VDD.n588 3.28454
R1301 VDD.n1610 VDD.n1609 3.2486
R1302 VDD.n1401 VDD.n571 3.2486
R1303 VDD.n1767 VDD.t69 3.22394
R1304 VDD.n1761 VDD.t38 3.22394
R1305 VDD.n1754 VDD.t42 3.22394
R1306 VDD.n1786 VDD.t26 3.22394
R1307 VDD.n677 VDD.t14 3.22347
R1308 VDD.n673 VDD.t74 3.22347
R1309 VDD.n669 VDD.t61 3.22347
R1310 VDD.n665 VDD.t64 3.22347
R1311 VDD.n1298 VDD.t72 3.21802
R1312 VDD.n405 VDD.t32 3.21788
R1313 VDD.n390 VDD.t20 3.21785
R1314 VDD.n1294 VDD.t56 3.21781
R1315 VDD.n411 VDD.t40 3.21767
R1316 VDD.n1317 VDD.t29 3.21766
R1317 VDD.n1629 VDD.n1628 3.21752
R1318 VDD.n1308 VDD.t17 3.21671
R1319 VDD.n398 VDD.t77 3.21657
R1320 VDD.n55 VDD.n54 3.21512
R1321 VDD.n189 VDD.n188 3.20353
R1322 VDD.n101 VDD.n100 3.20342
R1323 VDD.n1393 VDD.t48 3.19864
R1324 VDD.n1358 VDD.t23 3.19113
R1325 VDD.n1560 VDD.t51 3.19113
R1326 VDD.n1600 VDD.t67 3.18927
R1327 VDD.n425 VDD.t54 3.1878
R1328 VDD.n574 VDD.t59 3.1878
R1329 VDD.n1127 VDD.n1126 3.16769
R1330 VDD.n1747 VDD.n1746 3.16769
R1331 VDD.n57 VDD.n56 3.16326
R1332 VDD.n47 VDD.n46 3.15744
R1333 VDD.n781 VDD.n780 3.15287
R1334 VDD VDD.n779 3.15287
R1335 VDD.n999 VDD.n997 3.15287
R1336 VDD.n1001 VDD.n1000 3.15287
R1337 VDD.n996 VDD.n995 3.15287
R1338 VDD VDD.n1914 3.15269
R1339 VDD.n1665 VDD.n377 3.15151
R1340 VDD.n1599 VDD.n429 3.1505
R1341 VDD.n1604 VDD.n1603 3.1505
R1342 VDD.n1602 VDD.n427 3.1505
R1343 VDD.n1606 VDD.n427 3.1505
R1344 VDD.n1608 VDD.n428 3.1505
R1345 VDD.n1608 VDD.n1607 3.1505
R1346 VDD.n1610 VDD.n426 3.1505
R1347 VDD.n1613 VDD.n1612 3.1505
R1348 VDD.n1612 VDD.n1611 3.1505
R1349 VDD.n1615 VDD.n423 3.1505
R1350 VDD.n423 VDD.n422 3.1505
R1351 VDD.n1617 VDD.n1616 3.1505
R1352 VDD.n1618 VDD.n1617 3.1505
R1353 VDD.n424 VDD.n378 3.1505
R1354 VDD.n1664 VDD.n1663 3.1505
R1355 VDD.n381 VDD.n377 3.1505
R1356 VDD.n1667 VDD.n375 3.1505
R1357 VDD.n382 VDD.n375 3.1505
R1358 VDD.n1669 VDD.n1668 3.1505
R1359 VDD.n1670 VDD.n1669 3.1505
R1360 VDD.n368 VDD.n367 3.1505
R1361 VDD.n1671 VDD.n368 3.1505
R1362 VDD.n1681 VDD.n1680 3.1505
R1363 VDD.n1680 VDD.n1679 3.1505
R1364 VDD.n1682 VDD.n366 3.1505
R1365 VDD.n370 VDD.n366 3.1505
R1366 VDD.n1684 VDD.n1683 3.1505
R1367 VDD.n1685 VDD.n1684 3.1505
R1368 VDD.n339 VDD.n337 3.1505
R1369 VDD.n1686 VDD.n339 3.1505
R1370 VDD.n1707 VDD.n1706 3.1505
R1371 VDD.n1706 VDD.n1705 3.1505
R1372 VDD.n340 VDD.n338 3.1505
R1373 VDD.n1692 VDD.n340 3.1505
R1374 VDD.n1695 VDD.n1694 3.1505
R1375 VDD.n1696 VDD.n1695 3.1505
R1376 VDD.n273 VDD.n270 3.1505
R1377 VDD.n1697 VDD.n273 3.1505
R1378 VDD.n1660 VDD.n376 3.1505
R1379 VDD.n391 VDD.n380 3.1505
R1380 VDD.n1656 VDD.n1655 3.1505
R1381 VDD.n1653 VDD.n389 3.1505
R1382 VDD.n1652 VDD.n1651 3.1505
R1383 VDD.n1650 VDD.n1649 3.1505
R1384 VDD.n1647 VDD.n1646 3.1505
R1385 VDD.n1645 VDD.n1644 3.1505
R1386 VDD.n1643 VDD.n1642 3.1505
R1387 VDD.n1641 VDD.n1640 3.1505
R1388 VDD.n1639 VDD.n1638 3.1505
R1389 VDD.n1637 VDD.n1636 3.1505
R1390 VDD.n1634 VDD.n1633 3.1505
R1391 VDD.n1632 VDD.n1631 3.1505
R1392 VDD.n1630 VDD.n1629 3.1505
R1393 VDD.n1575 VDD.n1574 3.1505
R1394 VDD.n1577 VDD.n1576 3.1505
R1395 VDD.n1579 VDD.n1578 3.1505
R1396 VDD.n1581 VDD.n1580 3.1505
R1397 VDD.n1583 VDD.n1582 3.1505
R1398 VDD.n1585 VDD.n1584 3.1505
R1399 VDD.n1587 VDD.n1586 3.1505
R1400 VDD.n1589 VDD.n1588 3.1505
R1401 VDD.n1591 VDD.n1590 3.1505
R1402 VDD.n1593 VDD.n1592 3.1505
R1403 VDD.n431 VDD.n430 3.1505
R1404 VDD.n1598 VDD.n1597 3.1505
R1405 VDD VDD.n1501 3.1505
R1406 VDD.n1509 VDD.n1501 3.1505
R1407 VDD.n1521 VDD.n1520 3.1505
R1408 VDD.n1520 VDD.n1519 3.1505
R1409 VDD.n1508 VDD.n1507 3.1505
R1410 VDD.n1518 VDD.n1508 3.1505
R1411 VDD.n1516 VDD.n1515 3.1505
R1412 VDD.n1517 VDD.n1516 3.1505
R1413 VDD.n1514 VDD.n1510 3.1505
R1414 VDD.n1529 VDD.n1528 3.1505
R1415 VDD.n1498 VDD.n1497 3.1505
R1416 VDD.n1527 VDD.n1498 3.1505
R1417 VDD.n1525 VDD.n1524 3.1505
R1418 VDD.n1526 VDD.n1525 3.1505
R1419 VDD.n1523 VDD.n1500 3.1505
R1420 VDD.n1500 VDD.n1499 3.1505
R1421 VDD.n1489 VDD.n1488 3.1505
R1422 VDD.n1536 VDD.n1489 3.1505
R1423 VDD.n1534 VDD.n1533 3.1505
R1424 VDD.n1535 VDD.n1534 3.1505
R1425 VDD.n1532 VDD.n1490 3.1505
R1426 VDD.n530 VDD.n519 3.1505
R1427 VDD.n522 VDD.n519 3.1505
R1428 VDD.n529 VDD.n528 3.1505
R1429 VDD.n528 VDD.n527 3.1505
R1430 VDD.n521 VDD.n520 3.1505
R1431 VDD.n526 VDD.n521 3.1505
R1432 VDD.n525 VDD.n524 3.1505
R1433 VDD.n538 VDD.n508 3.1505
R1434 VDD.n537 VDD.n510 3.1505
R1435 VDD.n537 VDD.n536 3.1505
R1436 VDD.n513 VDD.n509 3.1505
R1437 VDD.n535 VDD.n509 3.1505
R1438 VDD.n533 VDD.n532 3.1505
R1439 VDD.n534 VDD.n533 3.1505
R1440 VDD VDD.n512 3.1505
R1441 VDD.n512 VDD.n511 3.1505
R1442 VDD.n544 VDD.n543 3.1505
R1443 VDD.n550 VDD.n549 3.1505
R1444 VDD.n551 VDD.n550 3.1505
R1445 VDD.n548 VDD.n503 3.1505
R1446 VDD.n503 VDD.n502 3.1505
R1447 VDD.n547 VDD.n546 3.1505
R1448 VDD.n546 VDD.n545 3.1505
R1449 VDD.n492 VDD.n491 3.1505
R1450 VDD.n558 VDD.n557 3.1505
R1451 VDD.n559 VDD.n558 3.1505
R1452 VDD.n556 VDD.n494 3.1505
R1453 VDD.n494 VDD.n493 3.1505
R1454 VDD.n555 VDD.n554 3.1505
R1455 VDD.n554 VDD.n553 3.1505
R1456 VDD VDD.n501 3.1505
R1457 VDD.n552 VDD.n501 3.1505
R1458 VDD.n1408 VDD.n1407 3.1505
R1459 VDD.n1391 VDD.n573 3.1505
R1460 VDD.n573 VDD.n572 3.1505
R1461 VDD.n1398 VDD.n1397 3.1505
R1462 VDD.n1399 VDD.n1398 3.1505
R1463 VDD.n1396 VDD.n571 3.1505
R1464 VDD.n1395 VDD.n569 3.1505
R1465 VDD.n1402 VDD.n569 3.1505
R1466 VDD.n1404 VDD.n568 3.1505
R1467 VDD.n1404 VDD.n1403 3.1505
R1468 VDD.n1406 VDD.n1405 3.1505
R1469 VDD.n1390 VDD.n1389 3.1505
R1470 VDD.n1389 VDD.n1388 3.1505
R1471 VDD.n581 VDD.n580 3.1505
R1472 VDD.n576 VDD.n575 3.1505
R1473 VDD.n1135 VDD.n1134 3.1505
R1474 VDD.n1134 VDD.n1133 3.1505
R1475 VDD.n1136 VDD.n656 3.1505
R1476 VDD.n656 VDD.n653 3.1505
R1477 VDD.n1138 VDD.n1137 3.1505
R1478 VDD.n1139 VDD.n1138 3.1505
R1479 VDD.n649 VDD.n648 3.1505
R1480 VDD.n654 VDD.n649 3.1505
R1481 VDD.n1150 VDD.n1149 3.1505
R1482 VDD.n1149 VDD.n1148 3.1505
R1483 VDD.n1151 VDD.n642 3.1505
R1484 VDD.n642 VDD.n641 3.1505
R1485 VDD.n1155 VDD.n1154 3.1505
R1486 VDD.n1156 VDD.n1155 3.1505
R1487 VDD.n1153 VDD.n647 3.1505
R1488 VDD.n647 VDD.n646 3.1505
R1489 VDD.n634 VDD.n633 3.1505
R1490 VDD.n644 VDD.n633 3.1505
R1491 VDD.n1220 VDD.n1219 3.1505
R1492 VDD.n1221 VDD.n1220 3.1505
R1493 VDD.n624 VDD.n623 3.1505
R1494 VDD.n631 VDD.n624 3.1505
R1495 VDD.n1233 VDD.n1232 3.1505
R1496 VDD.n1232 VDD.n1231 3.1505
R1497 VDD.n1234 VDD.n622 3.1505
R1498 VDD.n622 VDD.n620 3.1505
R1499 VDD.n1236 VDD.n1235 3.1505
R1500 VDD.n1237 VDD.n1236 3.1505
R1501 VDD.n615 VDD.n614 3.1505
R1502 VDD.n616 VDD.n615 3.1505
R1503 VDD.n1249 VDD.n1248 3.1505
R1504 VDD.n1248 VDD.n1247 3.1505
R1505 VDD.n1250 VDD.n612 3.1505
R1506 VDD.n612 VDD.n610 3.1505
R1507 VDD.n1253 VDD.n1252 3.1505
R1508 VDD.n1254 VDD.n1253 3.1505
R1509 VDD.n605 VDD.n604 3.1505
R1510 VDD.n606 VDD.n605 3.1505
R1511 VDD.n1266 VDD.n1265 3.1505
R1512 VDD.n1265 VDD.n1264 3.1505
R1513 VDD.n1267 VDD.n602 3.1505
R1514 VDD.n602 VDD.n600 3.1505
R1515 VDD.n658 VDD.n657 3.1505
R1516 VDD.n661 VDD.n658 3.1505
R1517 VDD.n795 VDD.n763 3.1505
R1518 VDD.n738 VDD.n732 3.1505
R1519 VDD.n740 VDD.n738 3.1505
R1520 VDD.n814 VDD.n813 3.1505
R1521 VDD.n815 VDD.n814 3.1505
R1522 VDD.n811 VDD.n758 3.1505
R1523 VDD.n761 VDD.n758 3.1505
R1524 VDD.n806 VDD.n805 3.1505
R1525 VDD.n807 VDD.n806 3.1505
R1526 VDD.n817 VDD.n756 3.1505
R1527 VDD.n817 VDD.n816 3.1505
R1528 VDD.n812 VDD.n755 3.1505
R1529 VDD.n757 VDD.n755 3.1505
R1530 VDD.n810 VDD.n809 3.1505
R1531 VDD.n809 VDD.n808 3.1505
R1532 VDD VDD.n821 3.1505
R1533 VDD.n821 VDD.n820 3.1505
R1534 VDD.n818 VDD 3.1505
R1535 VDD.n819 VDD.n818 3.1505
R1536 VDD.n695 VDD.n690 3.1505
R1537 VDD.n717 VDD.n690 3.1505
R1538 VDD.n835 VDD.n834 3.1505
R1539 VDD.n834 VDD.n833 3.1505
R1540 VDD.n742 VDD.n691 3.1505
R1541 VDD.n746 VDD.n691 3.1505
R1542 VDD.n711 VDD.n710 3.1505
R1543 VDD.n710 VDD.n700 3.1505
R1544 VDD.n721 VDD.n693 3.1505
R1545 VDD.n722 VDD.n721 3.1505
R1546 VDD.n751 VDD.n741 3.1505
R1547 VDD.n747 VDD.n741 3.1505
R1548 VDD.n716 VDD.n694 3.1505
R1549 VDD.n708 VDD.n701 3.1505
R1550 VDD.n712 VDD.n694 3.1505
R1551 VDD.n720 VDD.n688 3.1505
R1552 VDD.n720 VDD.n692 3.1505
R1553 VDD.n953 VDD.n949 3.1505
R1554 VDD.n948 VDD.n947 3.1505
R1555 VDD.n956 VDD.n948 3.1505
R1556 VDD.n959 VDD.n958 3.1505
R1557 VDD.n958 VDD.n957 3.1505
R1558 VDD.n960 VDD.n941 3.1505
R1559 VDD.n941 VDD.n940 3.1505
R1560 VDD.n962 VDD 3.1505
R1561 VDD.n963 VDD.n962 3.1505
R1562 VDD.n939 VDD.n938 3.1505
R1563 VDD.n964 VDD.n939 3.1505
R1564 VDD.n968 VDD.n967 3.1505
R1565 VDD.n967 VDD.n966 3.1505
R1566 VDD.n969 VDD.n937 3.1505
R1567 VDD.n965 VDD.n937 3.1505
R1568 VDD.n936 VDD.n935 3.1505
R1569 VDD.n889 VDD.n887 3.1505
R1570 VDD.n889 VDD.n888 3.1505
R1571 VDD.n891 VDD.n890 3.1505
R1572 VDD.n890 VDD.n878 3.1505
R1573 VDD.n877 VDD.n876 3.1505
R1574 VDD.n894 VDD.n877 3.1505
R1575 VDD.n897 VDD.n896 3.1505
R1576 VDD.n896 VDD.n895 3.1505
R1577 VDD.n887 VDD.n879 3.1505
R1578 VDD.n888 VDD.n879 3.1505
R1579 VDD.n892 VDD.n891 3.1505
R1580 VDD.n892 VDD.n878 3.1505
R1581 VDD.n893 VDD.n876 3.1505
R1582 VDD.n894 VDD.n893 3.1505
R1583 VDD.n897 VDD.n875 3.1505
R1584 VDD.n895 VDD.n875 3.1505
R1585 VDD VDD.n872 3.1505
R1586 VDD.n874 VDD.n872 3.1505
R1587 VDD.n912 VDD.n873 3.1505
R1588 VDD.n912 VDD.n911 3.1505
R1589 VDD.n913 VDD.n870 3.1505
R1590 VDD.n914 VDD.n913 3.1505
R1591 VDD.n917 VDD.n869 3.1505
R1592 VDD.n915 VDD.n869 3.1505
R1593 VDD.n919 VDD.n918 3.1505
R1594 VDD.n920 VDD.n919 3.1505
R1595 VDD.n923 VDD.n867 3.1505
R1596 VDD.n921 VDD.n867 3.1505
R1597 VDD.n909 VDD 3.1505
R1598 VDD.n909 VDD.n874 3.1505
R1599 VDD.n910 VDD.n873 3.1505
R1600 VDD.n911 VDD.n910 3.1505
R1601 VDD.n871 VDD.n870 3.1505
R1602 VDD.n914 VDD.n871 3.1505
R1603 VDD.n917 VDD.n916 3.1505
R1604 VDD.n916 VDD.n915 3.1505
R1605 VDD.n918 VDD.n868 3.1505
R1606 VDD.n920 VDD.n868 3.1505
R1607 VDD.n1059 VDD.n1058 3.1505
R1608 VDD.n1058 VDD.n1049 3.1505
R1609 VDD.n1057 VDD.n1048 3.1505
R1610 VDD.n1057 VDD.n1056 3.1505
R1611 VDD.n1051 VDD.n1050 3.1505
R1612 VDD.n1055 VDD.n1050 3.1505
R1613 VDD.n1054 VDD.n1053 3.1505
R1614 VDD.n1029 VDD.n1028 3.1505
R1615 VDD.n1062 VDD.n1061 3.1505
R1616 VDD.n1063 VDD.n1062 3.1505
R1617 VDD VDD.n1042 3.1505
R1618 VDD.n1042 VDD.n1041 3.1505
R1619 VDD.n1125 VDD.n660 3.1505
R1620 VDD.n1123 VDD.n1122 3.1505
R1621 VDD.n1121 VDD.n664 3.1505
R1622 VDD.n1119 VDD.n1118 3.1505
R1623 VDD.n1117 VDD.n666 3.1505
R1624 VDD.n1115 VDD.n1114 3.1505
R1625 VDD.n1113 VDD.n668 3.1505
R1626 VDD.n1111 VDD.n1110 3.1505
R1627 VDD.n1109 VDD.n670 3.1505
R1628 VDD.n1107 VDD.n1106 3.1505
R1629 VDD.n1104 VDD.n672 3.1505
R1630 VDD.n1103 VDD.n1102 3.1505
R1631 VDD.n1101 VDD.n674 3.1505
R1632 VDD.n1099 VDD.n1098 3.1505
R1633 VDD.n1096 VDD.n676 3.1505
R1634 VDD.n1095 VDD.n1094 3.1505
R1635 VDD.n1128 VDD.n659 3.1505
R1636 VDD.n662 VDD.n659 3.1505
R1637 VDD.n1130 VDD.n1129 3.1505
R1638 VDD.n1131 VDD.n1130 3.1505
R1639 VDD.n652 VDD.n651 3.1505
R1640 VDD.n1132 VDD.n652 3.1505
R1641 VDD.n1142 VDD.n1141 3.1505
R1642 VDD.n1141 VDD.n1140 3.1505
R1643 VDD.n1143 VDD.n650 3.1505
R1644 VDD.n655 VDD.n650 3.1505
R1645 VDD.n1145 VDD.n1144 3.1505
R1646 VDD.n1146 VDD.n1145 3.1505
R1647 VDD.n639 VDD.n637 3.1505
R1648 VDD.n1147 VDD.n639 3.1505
R1649 VDD.n1159 VDD.n1158 3.1505
R1650 VDD.n1158 VDD.n1157 3.1505
R1651 VDD.n640 VDD.n638 3.1505
R1652 VDD.n643 VDD.n640 3.1505
R1653 VDD.n630 VDD.n629 3.1505
R1654 VDD.n645 VDD.n630 3.1505
R1655 VDD.n1224 VDD.n1223 3.1505
R1656 VDD.n1223 VDD.n1222 3.1505
R1657 VDD.n1226 VDD.n625 3.1505
R1658 VDD.n632 VDD.n625 3.1505
R1659 VDD.n1228 VDD.n1227 3.1505
R1660 VDD.n1229 VDD.n1228 3.1505
R1661 VDD.n619 VDD.n618 3.1505
R1662 VDD.n1230 VDD.n619 3.1505
R1663 VDD.n1240 VDD.n1239 3.1505
R1664 VDD.n1239 VDD.n1238 3.1505
R1665 VDD.n1241 VDD.n617 3.1505
R1666 VDD.n621 VDD.n617 3.1505
R1667 VDD.n1244 VDD.n1243 3.1505
R1668 VDD.n1245 VDD.n1244 3.1505
R1669 VDD.n1242 VDD.n609 3.1505
R1670 VDD.n1246 VDD.n609 3.1505
R1671 VDD.n1257 VDD.n1256 3.1505
R1672 VDD.n1256 VDD.n1255 3.1505
R1673 VDD.n1258 VDD.n607 3.1505
R1674 VDD.n611 VDD.n607 3.1505
R1675 VDD.n1261 VDD.n1260 3.1505
R1676 VDD.n1262 VDD.n1261 3.1505
R1677 VDD.n1259 VDD.n599 3.1505
R1678 VDD.n1263 VDD.n599 3.1505
R1679 VDD.n1274 VDD.n1273 3.1505
R1680 VDD.n1273 VDD.n1272 3.1505
R1681 VDD.n1275 VDD.n597 3.1505
R1682 VDD.n601 VDD.n597 3.1505
R1683 VDD.n1277 VDD.n1276 3.1505
R1684 VDD.n1278 VDD.n1277 3.1505
R1685 VDD.n590 VDD.n589 3.1505
R1686 VDD.n1279 VDD.n590 3.1505
R1687 VDD.n1290 VDD.n1289 3.1505
R1688 VDD.n1289 VDD.n1288 3.1505
R1689 VDD.n1291 VDD.n587 3.1505
R1690 VDD.n592 VDD.n587 3.1505
R1691 VDD.n1377 VDD.n1376 3.1505
R1692 VDD.n1378 VDD.n1377 3.1505
R1693 VDD.n1270 VDD.n1269 3.1505
R1694 VDD.n1271 VDD.n1270 3.1505
R1695 VDD.n595 VDD.n594 3.1505
R1696 VDD.n596 VDD.n595 3.1505
R1697 VDD.n1282 VDD.n1281 3.1505
R1698 VDD.n1281 VDD.n1280 3.1505
R1699 VDD.n1283 VDD.n593 3.1505
R1700 VDD.n593 VDD.n591 3.1505
R1701 VDD.n1286 VDD.n1285 3.1505
R1702 VDD.n1287 VDD.n1286 3.1505
R1703 VDD.n1284 VDD.n585 3.1505
R1704 VDD.n586 VDD.n585 3.1505
R1705 VDD.n1380 VDD.n582 3.1505
R1706 VDD.n1380 VDD.n1379 3.1505
R1707 VDD.n1386 VDD.n1385 3.1505
R1708 VDD.n1387 VDD.n1386 3.1505
R1709 VDD.n1343 VDD.n1292 3.1505
R1710 VDD.n1342 VDD.n1341 3.1505
R1711 VDD.n1339 VDD.n1338 3.1505
R1712 VDD.n1337 VDD.n1336 3.1505
R1713 VDD.n1335 VDD.n1334 3.1505
R1714 VDD.n1333 VDD.n1332 3.1505
R1715 VDD.n1331 VDD.n1330 3.1505
R1716 VDD.n1329 VDD.n1328 3.1505
R1717 VDD.n1326 VDD.n1325 3.1505
R1718 VDD.n1324 VDD.n1309 3.1505
R1719 VDD.n1322 VDD.n1321 3.1505
R1720 VDD.n1319 VDD.n1311 3.1505
R1721 VDD.n584 VDD.n583 3.1505
R1722 VDD.n1383 VDD.n1382 3.1505
R1723 VDD.n1382 VDD.n578 3.1505
R1724 VDD.n1346 VDD.n1345 3.1505
R1725 VDD.n1374 VDD.n1373 3.1505
R1726 VDD.n1371 VDD.n1370 3.1505
R1727 VDD.n1368 VDD.n1349 3.1505
R1728 VDD.n1349 VDD.n1348 3.1505
R1729 VDD.n1367 VDD.n1366 3.1505
R1730 VDD.n1366 VDD.n1365 3.1505
R1731 VDD.n1354 VDD.n1353 3.1505
R1732 VDD.n1364 VDD.n1354 3.1505
R1733 VDD.n1362 VDD.n1361 3.1505
R1734 VDD.n1363 VDD.n1362 3.1505
R1735 VDD.n1360 VDD.n1357 3.1505
R1736 VDD.n477 VDD.n475 3.1505
R1737 VDD.n1410 VDD.n1409 3.1505
R1738 VDD.n1412 VDD.n1411 3.1505
R1739 VDD.n1414 VDD.n1413 3.1505
R1740 VDD.n1416 VDD.n1415 3.1505
R1741 VDD.n1418 VDD.n1417 3.1505
R1742 VDD.n1420 VDD.n1419 3.1505
R1743 VDD.n1422 VDD.n1421 3.1505
R1744 VDD.n1424 VDD.n1423 3.1505
R1745 VDD.n1426 VDD.n1425 3.1505
R1746 VDD.n1428 VDD.n1427 3.1505
R1747 VDD.n1430 VDD.n1429 3.1505
R1748 VDD.n1432 VDD.n1431 3.1505
R1749 VDD.n1434 VDD.n1433 3.1505
R1750 VDD.n478 VDD.n476 3.1505
R1751 VDD.n1439 VDD.n1438 3.1505
R1752 VDD VDD.n1456 3.1505
R1753 VDD.n1456 VDD.n1455 3.1505
R1754 VDD.n1448 VDD.n1447 3.1505
R1755 VDD.n1449 VDD.n474 3.1505
R1756 VDD.n474 VDD.n473 3.1505
R1757 VDD.n1452 VDD.n1451 3.1505
R1758 VDD.n1453 VDD.n1452 3.1505
R1759 VDD.n1450 VDD.n472 3.1505
R1760 VDD.n1454 VDD.n472 3.1505
R1761 VDD.n1457 VDD.n465 3.1505
R1762 VDD.n465 VDD.n464 3.1505
R1763 VDD.n1459 VDD.n1458 3.1505
R1764 VDD.n1460 VDD.n1459 3.1505
R1765 VDD.n463 VDD.n462 3.1505
R1766 VDD.n1461 VDD.n463 3.1505
R1767 VDD.n1463 VDD.n1462 3.1505
R1768 VDD.n1477 VDD.n1476 3.1505
R1769 VDD.n1481 VDD.n448 3.1505
R1770 VDD.n1482 VDD.n1481 3.1505
R1771 VDD.n1480 VDD.n1479 3.1505
R1772 VDD.n1480 VDD.n1472 3.1505
R1773 VDD.n1478 VDD.n1473 3.1505
R1774 VDD.n1475 VDD.n1473 3.1505
R1775 VDD.n456 VDD 3.1505
R1776 VDD.n1483 VDD.n456 3.1505
R1777 VDD.n1468 VDD.n457 3.1505
R1778 VDD.n1469 VDD.n454 3.1505
R1779 VDD.n1470 VDD.n1469 3.1505
R1780 VDD.n1471 VDD.n455 3.1505
R1781 VDD.n1485 VDD.n1484 3.1505
R1782 VDD.n1539 VDD.n1538 3.1505
R1783 VDD.n1538 VDD.n1537 3.1505
R1784 VDD VDD.n447 3.1505
R1785 VDD.n447 VDD.n446 3.1505
R1786 VDD.n1542 VDD.n1541 3.1505
R1787 VDD.n1543 VDD.n1542 3.1505
R1788 VDD.n445 VDD.n444 3.1505
R1789 VDD.n1544 VDD.n445 3.1505
R1790 VDD.n1546 VDD.n1545 3.1505
R1791 VDD.n1573 VDD.n433 3.1505
R1792 VDD.n1595 VDD.n433 3.1505
R1793 VDD.n1572 VDD.n1571 3.1505
R1794 VDD.n1570 VDD.n1569 3.1505
R1795 VDD.n1559 VDD.n1556 3.1505
R1796 VDD.n1565 VDD.n1564 3.1505
R1797 VDD.n1566 VDD.n1565 3.1505
R1798 VDD.n1562 VDD.n1558 3.1505
R1799 VDD.n1558 VDD.n1557 3.1505
R1800 VDD.n1561 VDD.n418 3.1505
R1801 VDD.n420 VDD.n418 3.1505
R1802 VDD.n1622 VDD.n419 3.1505
R1803 VDD.n1622 VDD.n1621 3.1505
R1804 VDD.n1624 VDD.n1623 3.1505
R1805 VDD.n1627 VDD.n1626 3.1505
R1806 VDD.n1568 VDD.n1555 3.1505
R1807 VDD.n373 VDD.n372 3.1505
R1808 VDD.n374 VDD.n373 3.1505
R1809 VDD.n1674 VDD.n1673 3.1505
R1810 VDD.n1673 VDD.n1672 3.1505
R1811 VDD.n1675 VDD.n371 3.1505
R1812 VDD.n371 VDD.n369 3.1505
R1813 VDD.n1677 VDD.n1676 3.1505
R1814 VDD.n1678 VDD.n1677 3.1505
R1815 VDD.n364 VDD.n363 3.1505
R1816 VDD.n365 VDD.n364 3.1505
R1817 VDD.n1688 VDD.n1687 3.1505
R1818 VDD.n1687 VDD.t168 3.1505
R1819 VDD.n1689 VDD.n342 3.1505
R1820 VDD.n342 VDD.n341 3.1505
R1821 VDD.n1703 VDD.n1702 3.1505
R1822 VDD.n1704 VDD.n1703 3.1505
R1823 VDD.n1701 VDD.n343 3.1505
R1824 VDD.n1693 VDD.n343 3.1505
R1825 VDD.n1700 VDD.n1699 3.1505
R1826 VDD.n1699 VDD.n1698 3.1505
R1827 VDD.n1691 VDD.n276 3.1505
R1828 VDD.n276 VDD.n275 3.1505
R1829 VDD.n1859 VDD.n1858 3.1505
R1830 VDD.n1860 VDD.n1859 3.1505
R1831 VDD.n1857 VDD.n277 3.1505
R1832 VDD.n282 VDD.n277 3.1505
R1833 VDD.n1856 VDD.n1855 3.1505
R1834 VDD.n1855 VDD.n1854 3.1505
R1835 VDD.n280 VDD.n279 3.1505
R1836 VDD.n284 VDD.n280 3.1505
R1837 VDD.n294 VDD.n292 3.1505
R1838 VDD.n292 VDD.n291 3.1505
R1839 VDD.n1845 VDD.n1844 3.1505
R1840 VDD.n1846 VDD.n1845 3.1505
R1841 VDD.n1843 VDD.n293 3.1505
R1842 VDD.n301 VDD.n293 3.1505
R1843 VDD.n1841 VDD.n1840 3.1505
R1844 VDD.n1840 VDD.n1839 3.1505
R1845 VDD.n299 VDD.n298 3.1505
R1846 VDD.n303 VDD.n299 3.1505
R1847 VDD.n314 VDD.n312 3.1505
R1848 VDD.n312 VDD.n311 3.1505
R1849 VDD.n1830 VDD.n1829 3.1505
R1850 VDD.n1831 VDD.n1830 3.1505
R1851 VDD.n1827 VDD.n313 3.1505
R1852 VDD.n1731 VDD.n313 3.1505
R1853 VDD.n1826 VDD.n1825 3.1505
R1854 VDD.n1825 VDD.n1824 3.1505
R1855 VDD.n1730 VDD.n1729 3.1505
R1856 VDD.n1733 VDD.n1730 3.1505
R1857 VDD.n1745 VDD.n1743 3.1505
R1858 VDD.n1743 VDD.n1741 3.1505
R1859 VDD.n1815 VDD.n1814 3.1505
R1860 VDD.n1816 VDD.n1815 3.1505
R1861 VDD.n1813 VDD.n1744 3.1505
R1862 VDD.n1798 VDD.n1744 3.1505
R1863 VDD.n1812 VDD.n1811 3.1505
R1864 VDD.n1769 VDD.n1763 3.1505
R1865 VDD.n1773 VDD.n1763 3.1505
R1866 VDD.n1775 VDD.n1764 3.1505
R1867 VDD.n1775 VDD.n1774 3.1505
R1868 VDD.n1776 VDD.n1762 3.1505
R1869 VDD.n1776 VDD.n1757 3.1505
R1870 VDD.n1778 VDD.n1777 3.1505
R1871 VDD.n1777 VDD.n1758 3.1505
R1872 VDD.n1779 VDD.n1760 3.1505
R1873 VDD.n1760 VDD.n1759 3.1505
R1874 VDD.n1782 VDD.n1781 3.1505
R1875 VDD.n1783 VDD.n1782 3.1505
R1876 VDD.n1753 VDD.n1751 3.1505
R1877 VDD.n1751 VDD.n1749 3.1505
R1878 VDD.n1805 VDD.n1804 3.1505
R1879 VDD.n1806 VDD.n1805 3.1505
R1880 VDD.n1802 VDD.n1752 3.1505
R1881 VDD.n1752 VDD.n1750 3.1505
R1882 VDD.n1801 VDD.n1800 3.1505
R1883 VDD.n1800 VDD.n1799 3.1505
R1884 VDD.n1756 VDD.n1755 3.1505
R1885 VDD.n1797 VDD.n1756 3.1505
R1886 VDD.n1795 VDD.n1794 3.1505
R1887 VDD.n1796 VDD.n1795 3.1505
R1888 VDD.n1792 VDD.n1785 3.1505
R1889 VDD.n1785 VDD.n1784 3.1505
R1890 VDD.n1791 VDD.n1790 3.1505
R1891 VDD.n1790 VDD.n1789 3.1505
R1892 VDD.n1788 VDD.n1787 3.1505
R1893 VDD.n1788 VDD.n1748 3.1505
R1894 VDD.n1771 VDD.n1770 3.1505
R1895 VDD.n1766 VDD.n1765 3.1505
R1896 VDD.n1739 VDD.n1738 3.1505
R1897 VDD.n1742 VDD.n1739 3.1505
R1898 VDD.n274 VDD.n271 3.1505
R1899 VDD.n281 VDD.n274 3.1505
R1900 VDD.n287 VDD.n285 3.1505
R1901 VDD.n285 VDD.n283 3.1505
R1902 VDD.n1852 VDD.n1851 3.1505
R1903 VDD.n1853 VDD.n1852 3.1505
R1904 VDD.n1850 VDD.n286 3.1505
R1905 VDD.n290 VDD.n286 3.1505
R1906 VDD.n1849 VDD.n1848 3.1505
R1907 VDD.n1848 VDD.n1847 3.1505
R1908 VDD.n289 VDD.n288 3.1505
R1909 VDD.n300 VDD.n289 3.1505
R1910 VDD.n306 VDD.n304 3.1505
R1911 VDD.n304 VDD.n302 3.1505
R1912 VDD.n1837 VDD.n1836 3.1505
R1913 VDD.n1838 VDD.n1837 3.1505
R1914 VDD.n1835 VDD.n305 3.1505
R1915 VDD.n310 VDD.n305 3.1505
R1916 VDD.n1834 VDD.n1833 3.1505
R1917 VDD.n1833 VDD.n1832 3.1505
R1918 VDD.n1736 VDD.n308 3.1505
R1919 VDD.n309 VDD.n308 3.1505
R1920 VDD.n1737 VDD.n1734 3.1505
R1921 VDD.n1734 VDD.n1732 3.1505
R1922 VDD.n1822 VDD.n1821 3.1505
R1923 VDD.n1823 VDD.n1822 3.1505
R1924 VDD.n1820 VDD.n1735 3.1505
R1925 VDD.n1740 VDD.n1735 3.1505
R1926 VDD.n1819 VDD.n1818 3.1505
R1927 VDD.n1818 VDD.n1817 3.1505
R1928 VDD.n1863 VDD.n1862 3.1505
R1929 VDD.n1862 VDD.n1861 3.1505
R1930 VDD.n1995 VDD.n1994 3.1505
R1931 VDD.n1994 VDD.n1993 3.1505
R1932 VDD.n1974 VDD.n1973 3.1505
R1933 VDD.n1973 VDD.n1972 3.1505
R1934 VDD.n1977 VDD.n1976 3.1505
R1935 VDD.n1976 VDD.n1975 3.1505
R1936 VDD VDD.n1985 3.1505
R1937 VDD.n1985 VDD.n1984 3.1505
R1938 VDD.n1983 VDD.n1981 3.1505
R1939 VDD.n1983 VDD.n1982 3.1505
R1940 VDD.n1980 VDD.n1979 3.1505
R1941 VDD.n1979 VDD.n1978 3.1505
R1942 VDD.n1968 VDD.n1967 3.1505
R1943 VDD.n1967 VDD.n1966 3.1505
R1944 VDD.n1955 VDD.n1954 3.1505
R1945 VDD.n1992 VDD.n1991 3.1505
R1946 VDD.n2028 VDD.n2027 3.1505
R1947 VDD.n2027 VDD.t106 3.1505
R1948 VDD.n1931 VDD.n1930 3.1505
R1949 VDD.n2026 VDD.n2025 3.1505
R1950 VDD.t106 VDD.n2026 3.1505
R1951 VDD.n1 VDD.n0 3.1505
R1952 VDD.n1028 VDD.n1027 3.14819
R1953 VDD.n168 VDD.n109 3.13854
R1954 VDD.n170 VDD.n106 3.13854
R1955 VDD.n171 VDD.n104 3.13854
R1956 VDD.n192 VDD.n185 3.13659
R1957 VDD.n198 VDD.n197 3.13659
R1958 VDD.n206 VDD.n195 3.13659
R1959 VDD.n1437 VDD.n478 3.09085
R1960 VDD.n1552 VDD.n1549 3.06224
R1961 VDD.n1506 VDD.n1505 3.06224
R1962 VDD.n518 VDD.n515 3.06224
R1963 VDD.n499 VDD.n496 3.06224
R1964 VDD.n737 VDD.n736 3.06224
R1965 VDD.n731 VDD.n728 3.06224
R1966 VDD.n946 VDD.n943 3.06224
R1967 VDD.n902 VDD.n899 3.06224
R1968 VDD.n907 VDD.n906 3.06224
R1969 VDD.n1047 VDD.n1044 3.06224
R1970 VDD.n470 VDD.n469 3.06224
R1971 VDD.n453 VDD.n452 3.06224
R1972 VDD.n1964 VDD.n1963 3.06224
R1973 VDD.n1596 VDD.n431 3.04049
R1974 VDD.n1576 VDD.n434 3.03982
R1975 VDD.n1411 VDD.n479 3.03982
R1976 VDD.n81 VDD.n79 2.98985
R1977 VDD.n77 VDD.n75 2.98985
R1978 VDD.n144 VDD.n136 2.98985
R1979 VDD.n140 VDD.n138 2.98985
R1980 VDD.n239 VDD.n237 2.98985
R1981 VDD.n243 VDD.n235 2.98985
R1982 VDD.n1887 VDD.n1885 2.98985
R1983 VDD.n1901 VDD.n1883 2.98985
R1984 VDD.n1926 VDD.n1925 2.98721
R1985 VDD.n63 VDD.n62 2.97811
R1986 VDD.n156 VDD.n134 2.97811
R1987 VDD.n158 VDD.n131 2.97811
R1988 VDD.n257 VDD.n230 2.97811
R1989 VDD.n255 VDD.n233 2.97811
R1990 VDD.n1879 VDD.n1878 2.97811
R1991 VDD.n1905 VDD.n1881 2.97811
R1992 VDD.n1146 VDD.t382 2.91474
R1993 VDD.n1247 VDD.t364 2.91474
R1994 VDD.n202 VDD.n200 2.88811
R1995 VDD.n786 VDD.n784 2.87637
R1996 VDD.n775 VDD.n773 2.87637
R1997 VDD.n991 VDD.n990 2.87637
R1998 VDD.n986 VDD.n985 2.87637
R1999 VDD.n1946 VDD.n1944 2.87637
R2000 VDD.n1999 VDD.n1998 2.87637
R2001 VDD.n67 VDD.t268 2.84673
R2002 VDD.n127 VDD.t552 2.84673
R2003 VDD.n226 VDD.t730 2.84631
R2004 VDD.n1891 VDD.t289 2.84631
R2005 VDD.n37 VDD.n36 2.82741
R2006 VDD.n119 VDD.n113 2.78441
R2007 VDD.n118 VDD.n115 2.78441
R2008 VDD.n215 VDD.n209 2.78441
R2009 VDD.n214 VDD.n211 2.78441
R2010 VDD.n1659 VDD.n380 2.7478
R2011 VDD.n1657 VDD.n380 2.7478
R2012 VDD.n176 VDD.n95 2.74538
R2013 VDD.n2025 VDD.n2024 2.60854
R2014 VDD.n150 VDD.n147 2.6005
R2015 VDD.n120 VDD.n111 2.6005
R2016 VDD.n218 VDD.n217 2.6005
R2017 VDD.n249 VDD.n248 2.6005
R2018 VDD.n1875 VDD.n1874 2.6005
R2019 VDD.n330 VDD.n329 2.6005
R2020 VDD.n397 VDD.n396 2.6005
R2021 VDD.n403 VDD.n402 2.6005
R2022 VDD.n1552 VDD.n1551 2.6005
R2023 VDD.n1506 VDD.n1503 2.6005
R2024 VDD.n1316 VDD.n1313 2.6005
R2025 VDD.n1305 VDD.n1302 2.6005
R2026 VDD.n518 VDD.n517 2.6005
R2027 VDD.n499 VDD.n498 2.6005
R2028 VDD.n1183 VDD.n1182 2.6005
R2029 VDD.n1163 VDD.n1162 2.6005
R2030 VDD.n1169 VDD.n1165 2.6005
R2031 VDD.n1168 VDD.n1167 2.6005
R2032 VDD.n1172 VDD.n1171 2.6005
R2033 VDD.n628 VDD.n627 2.6005
R2034 VDD.n1208 VDD.n1207 2.6005
R2035 VDD.n1205 VDD.n1204 2.6005
R2036 VDD.n1211 VDD.n1210 2.6005
R2037 VDD.n1216 VDD.n1215 2.6005
R2038 VDD.n737 VDD.n734 2.6005
R2039 VDD.n731 VDD.n730 2.6005
R2040 VDD.n946 VDD.n945 2.6005
R2041 VDD.n902 VDD.n901 2.6005
R2042 VDD.n907 VDD.n904 2.6005
R2043 VDD.n1047 VDD.n1046 2.6005
R2044 VDD.n1175 VDD.n1174 2.6005
R2045 VDD.n1190 VDD.n1189 2.6005
R2046 VDD.n1187 VDD.n1186 2.6005
R2047 VDD.n1196 VDD.n1180 2.6005
R2048 VDD.n1197 VDD.n1178 2.6005
R2049 VDD.n1193 VDD.n1192 2.6005
R2050 VDD.n470 VDD.n467 2.6005
R2051 VDD.n453 VDD.n450 2.6005
R2052 VDD.n346 VDD.n345 2.6005
R2053 VDD.n336 VDD.n335 2.6005
R2054 VDD.n362 VDD.n361 2.6005
R2055 VDD.n352 VDD.n351 2.6005
R2056 VDD.n297 VDD.n296 2.6005
R2057 VDD.n1728 VDD.n1727 2.6005
R2058 VDD.n324 VDD.n323 2.6005
R2059 VDD.n318 VDD.n317 2.6005
R2060 VDD.n1721 VDD.n1720 2.6005
R2061 VDD.n1724 VDD.n1723 2.6005
R2062 VDD.n355 VDD.n354 2.6005
R2063 VDD.n327 VDD.n326 2.6005
R2064 VDD.n333 VDD.n332 2.6005
R2065 VDD.n349 VDD.n348 2.6005
R2066 VDD.n1712 VDD.n1711 2.6005
R2067 VDD.n89 VDD.n86 2.6005
R2068 VDD.n1964 VDD.n1961 2.6005
R2069 VDD.n1590 VDD.n442 2.59264
R2070 VDD.n1586 VDD.n440 2.59264
R2071 VDD.n1582 VDD.n438 2.59264
R2072 VDD.n1578 VDD.n436 2.59264
R2073 VDD.n1593 VDD.n442 2.59264
R2074 VDD.n1588 VDD.n440 2.59264
R2075 VDD.n1584 VDD.n438 2.59264
R2076 VDD.n1580 VDD.n436 2.59264
R2077 VDD.n1435 VDD.n1434 2.59264
R2078 VDD.n1429 VDD.n489 2.59264
R2079 VDD.n1425 VDD.n487 2.59264
R2080 VDD.n1421 VDD.n485 2.59264
R2081 VDD.n1417 VDD.n483 2.59264
R2082 VDD.n1413 VDD.n481 2.59264
R2083 VDD.n1435 VDD.n478 2.59264
R2084 VDD.n1431 VDD.n489 2.59264
R2085 VDD.n1427 VDD.n487 2.59264
R2086 VDD.n1423 VDD.n485 2.59264
R2087 VDD.n1419 VDD.n483 2.59264
R2088 VDD.n1415 VDD.n481 2.59264
R2089 VDD.n178 VDD.n176 2.588
R2090 VDD.n1807 VDD.n1806 2.58448
R2091 VDD.n1588 VDD.n441 2.5167
R2092 VDD.n1584 VDD.n439 2.5167
R2093 VDD.n1580 VDD.n437 2.5167
R2094 VDD.n1576 VDD.n435 2.5167
R2095 VDD.n1590 VDD.n441 2.5167
R2096 VDD.n1586 VDD.n439 2.5167
R2097 VDD.n1582 VDD.n437 2.5167
R2098 VDD.n1578 VDD.n435 2.5167
R2099 VDD.n1431 VDD.n490 2.5167
R2100 VDD.n1427 VDD.n488 2.5167
R2101 VDD.n1423 VDD.n486 2.5167
R2102 VDD.n1419 VDD.n484 2.5167
R2103 VDD.n1415 VDD.n482 2.5167
R2104 VDD.n1434 VDD.n490 2.5167
R2105 VDD.n1429 VDD.n488 2.5167
R2106 VDD.n1425 VDD.n486 2.5167
R2107 VDD.n1421 VDD.n484 2.5167
R2108 VDD.n1417 VDD.n482 2.5167
R2109 VDD.n1824 VDD.t165 2.49842
R2110 VDD.n1808 VDD.n1807 2.49842
R2111 VDD.n662 VDD.n661 2.49842
R2112 VDD.n1594 VDD.n1593 2.47755
R2113 VDD.n1594 VDD.n431 2.47755
R2114 VDD.n1411 VDD.n480 2.47755
R2115 VDD.n1413 VDD.n480 2.47755
R2116 VDD.n1091 VDD.n1090 2.37611
R2117 VDD.n1929 VDD.n1928 2.36122
R2118 VDD.n2018 VDD.n1957 2.35567
R2119 VDD.n1088 VDD.n1087 2.34319
R2120 VDD.n1087 VDD.n679 2.33916
R2121 VDD.n2023 VDD.n2022 2.32106
R2122 VDD.n929 VDD.n928 2.31932
R2123 VDD.n791 VDD.n790 2.29638
R2124 VDD.n791 VDD.n770 2.29115
R2125 VDD.n1087 VDD.n1086 2.28732
R2126 VDD.n797 VDD.n796 2.2804
R2127 VDD.n1867 VDD.n1866 2.27396
R2128 VDD.n1531 VDD.n1530 2.25904
R2129 VDD.n1936 VDD.n1935 2.25144
R2130 VDD.n1865 VDD.n269 2.25144
R2131 VDD.n803 VDD.n802 2.2505
R2132 VDD.n689 VDD.n687 2.2505
R2133 VDD.n698 VDD.n697 2.2505
R2134 VDD.n726 VDD.n725 2.2505
R2135 VDD.n1008 VDD.n845 2.2505
R2136 VDD.n977 VDD.n976 2.2505
R2137 VDD.n858 VDD.n848 2.2505
R2138 VDD.n998 VDD.n842 2.2505
R2139 VDD.n1003 VDD.n1002 2.2505
R2140 VDD.n48 VDD.n47 2.2505
R2141 VDD.n2017 VDD.n2016 2.2505
R2142 VDD.n1082 VDD.n680 2.24806
R2143 VDD.n784 VDD.t577 2.16717
R2144 VDD.n784 VDD.n783 2.16717
R2145 VDD.n773 VDD.t760 2.16717
R2146 VDD.n773 VDD.n772 2.16717
R2147 VDD.n990 VDD.t581 2.16717
R2148 VDD.n990 VDD.n989 2.16717
R2149 VDD.n985 VDD.t748 2.16717
R2150 VDD.n985 VDD.n984 2.16717
R2151 VDD.n1944 VDD.t703 2.16717
R2152 VDD.n1944 VDD.n1943 2.16717
R2153 VDD.n1998 VDD.t727 2.16717
R2154 VDD.n1998 VDD.n1997 2.16717
R2155 VDD.n1909 VDD.n1870 2.06447
R2156 VDD VDD.n1888 2.06161
R2157 VDD.n832 VDD.n693 2.05248
R2158 VDD.t679 VDD.n746 2.05248
R2159 VDD.n816 VDD.t682 2.05248
R2160 VDD.n895 VDD.t355 2.05248
R2161 VDD.n1342 VDD.n1293 2.04683
R2162 VDD.n1338 VDD.n1293 2.04625
R2163 VDD.n1633 VDD.n384 2.04615
R2164 VDD.n1637 VDD.n384 2.04615
R2165 VDD VDD.n64 2.01923
R2166 VDD.n1811 VDD.n1810 2.00622
R2167 VDD.n1810 VDD.n1747 2.00565
R2168 VDD.n1337 VDD.n1297 1.94801
R2169 VDD.n1334 VDD.n1297 1.94746
R2170 VDD.n1638 VDD.n385 1.94734
R2171 VDD.n1641 VDD.n385 1.94734
R2172 VDD.n792 VDD.n791 1.94241
R2173 VDD.n1066 VDD.n1032 1.9255
R2174 VDD.n1595 VDD.n1594 1.91272
R2175 VDD.n1436 VDD.n480 1.91272
R2176 VDD.n1547 VDD.n1546 1.8985
R2177 VDD.n1595 VDD.n435 1.89315
R2178 VDD.n1595 VDD.n437 1.89315
R2179 VDD.n1595 VDD.n439 1.89315
R2180 VDD.n1595 VDD.n441 1.89315
R2181 VDD.n1436 VDD.n482 1.89315
R2182 VDD.n1436 VDD.n484 1.89315
R2183 VDD.n1436 VDD.n486 1.89315
R2184 VDD.n1436 VDD.n488 1.89315
R2185 VDD.n1436 VDD.n490 1.89315
R2186 VDD.n162 VDD.n123 1.87485
R2187 VDD.n261 VDD.n222 1.87485
R2188 VDD.n424 VDD.n379 1.87282
R2189 VDD.n580 VDD.n577 1.87282
R2190 VDD.n1663 VDD.n379 1.87228
R2191 VDD.n577 VDD.n576 1.87228
R2192 VDD.n1569 VDD.n432 1.8617
R2193 VDD.n1571 VDD.n432 1.8617
R2194 VDD.n1595 VDD.n436 1.85518
R2195 VDD.n1595 VDD.n438 1.85518
R2196 VDD.n1595 VDD.n440 1.85518
R2197 VDD.n1595 VDD.n442 1.85518
R2198 VDD.n1436 VDD.n481 1.85518
R2199 VDD.n1436 VDD.n483 1.85518
R2200 VDD.n1436 VDD.n485 1.85518
R2201 VDD.n1436 VDD.n487 1.85518
R2202 VDD.n1436 VDD.n489 1.85518
R2203 VDD.n1436 VDD.n1435 1.85518
R2204 VDD.n762 VDD.n760 1.85344
R2205 VDD.n804 VDD.n760 1.85344
R2206 VDD.n922 VDD.n921 1.85344
R2207 VDD.n923 VDD.n922 1.85344
R2208 VDD.n1329 VDD.n1307 1.83567
R2209 VDD.n1325 VDD.n1307 1.83513
R2210 VDD.n1646 VDD.n387 1.835
R2211 VDD.n1650 VDD.n387 1.835
R2212 VDD.n1324 VDD.n1323 1.82979
R2213 VDD.n1323 VDD.n1322 1.82925
R2214 VDD.n1651 VDD.n388 1.82912
R2215 VDD.n389 VDD.n388 1.82912
R2216 VDD VDD.n778 1.82452
R2217 VDD.n1486 VDD.n455 1.80965
R2218 VDD.n1486 VDD.n1485 1.80912
R2219 VDD.n744 VDD.n721 1.7505
R2220 VDD.n2021 VDD.n2020 1.71333
R2221 VDD.n1344 VDD.n1343 1.69304
R2222 VDD.n1333 VDD.n1300 1.69304
R2223 VDD.n1311 VDD.n1310 1.69304
R2224 VDD.n1310 VDD.n584 1.69252
R2225 VDD.n1330 VDD.n1300 1.69252
R2226 VDD.n1345 VDD.n1344 1.69252
R2227 VDD.n1642 VDD.n386 1.69238
R2228 VDD.n1629 VDD.n383 1.69238
R2229 VDD.n1645 VDD.n386 1.69238
R2230 VDD.n1632 VDD.n383 1.69238
R2231 VDD.n1125 VDD.n1124 1.66029
R2232 VDD.n1124 VDD.n1123 1.65977
R2233 VDD.n1118 VDD.n667 1.65963
R2234 VDD.n1116 VDD.n1115 1.65963
R2235 VDD.n1110 VDD.n671 1.65963
R2236 VDD.n1108 VDD.n1107 1.65963
R2237 VDD.n1102 VDD.n675 1.65963
R2238 VDD.n1100 VDD.n1099 1.65963
R2239 VDD.n1094 VDD.n1093 1.65963
R2240 VDD.n667 VDD.n664 1.65963
R2241 VDD.n1117 VDD.n1116 1.65963
R2242 VDD.n671 VDD.n668 1.65963
R2243 VDD.n1109 VDD.n1108 1.65963
R2244 VDD.n675 VDD.n672 1.65963
R2245 VDD.n1101 VDD.n1100 1.65963
R2246 VDD.n1093 VDD.n676 1.65963
R2247 VDD.n102 VDD.n99 1.64018
R2248 VDD.n190 VDD.n187 1.64018
R2249 VDD.n62 VDD.t535 1.6255
R2250 VDD.n62 VDD.n61 1.6255
R2251 VDD.n66 VDD.t263 1.6255
R2252 VDD.n66 VDD.n65 1.6255
R2253 VDD.n79 VDD.t512 1.6255
R2254 VDD.n79 VDD.n78 1.6255
R2255 VDD.n75 VDD.t537 1.6255
R2256 VDD.n75 VDD.n74 1.6255
R2257 VDD.n136 VDD.t593 1.6255
R2258 VDD.n136 VDD.n135 1.6255
R2259 VDD.n138 VDD.t320 1.6255
R2260 VDD.n138 VDD.n137 1.6255
R2261 VDD.n147 VDD.t270 1.6255
R2262 VDD.n147 VDD.n146 1.6255
R2263 VDD.n149 VDD.t281 1.6255
R2264 VDD.n149 VDD.n148 1.6255
R2265 VDD.n134 VDD.t526 1.6255
R2266 VDD.n134 VDD.n133 1.6255
R2267 VDD.n131 VDD.t653 1.6255
R2268 VDD.n131 VDD.n130 1.6255
R2269 VDD.n126 VDD.t553 1.6255
R2270 VDD.n126 VDD.n125 1.6255
R2271 VDD.n237 VDD.t499 1.6255
R2272 VDD.n237 VDD.n236 1.6255
R2273 VDD.n235 VDD.t113 1.6255
R2274 VDD.n235 VDD.n234 1.6255
R2275 VDD.n225 VDD.t251 1.6255
R2276 VDD.n225 VDD.n224 1.6255
R2277 VDD.n230 VDD.t557 1.6255
R2278 VDD.n230 VDD.n229 1.6255
R2279 VDD.n233 VDD.t697 1.6255
R2280 VDD.n233 VDD.n232 1.6255
R2281 VDD.n248 VDD.t229 1.6255
R2282 VDD.n248 VDD.n247 1.6255
R2283 VDD.n246 VDD.t233 1.6255
R2284 VDD.n246 VDD.n245 1.6255
R2285 VDD.n1885 VDD.t666 1.6255
R2286 VDD.n1885 VDD.n1884 1.6255
R2287 VDD.n1883 VDD.t545 1.6255
R2288 VDD.n1883 VDD.n1882 1.6255
R2289 VDD.n1890 VDD.t290 1.6255
R2290 VDD.n1890 VDD.n1889 1.6255
R2291 VDD.n1878 VDD.t325 1.6255
R2292 VDD.n1878 VDD.n1877 1.6255
R2293 VDD.n1881 VDD.t212 1.6255
R2294 VDD.n1881 VDD.n1880 1.6255
R2295 VDD.n1874 VDD.t497 1.6255
R2296 VDD.n1874 VDD.n1873 1.6255
R2297 VDD.n1872 VDD.t304 1.6255
R2298 VDD.n1872 VDD.n1871 1.6255
R2299 VDD.n86 VDD.t338 1.6255
R2300 VDD.n86 VDD.n85 1.6255
R2301 VDD.n88 VDD.t333 1.6255
R2302 VDD.n88 VDD.n87 1.6255
R2303 VDD.n1925 VDD.t522 1.6255
R2304 VDD.n1925 VDD.n1924 1.6255
R2305 VDD.n1184 VDD.n636 1.5755
R2306 VDD.n1074 VDD.n1019 1.5755
R2307 VDD.n1716 VDD.n1715 1.5755
R2308 VDD.n1200 VDD.n1199 1.57159
R2309 VDD.n357 VDD.n356 1.57159
R2310 VDD.n1438 VDD.n1437 1.54574
R2311 VDD.n1597 VDD.n1596 1.52056
R2312 VDD.n1574 VDD.n434 1.52041
R2313 VDD.n1409 VDD.n479 1.52041
R2314 VDD.n1071 VDD.n1033 1.5005
R2315 VDD.n1217 VDD.n613 1.49724
R2316 VDD.n321 VDD.n272 1.49724
R2317 VDD.n1028 VDD.n1021 1.488
R2318 VDD.n1014 VDD.n1013 1.42211
R2319 VDD.n982 VDD.n981 1.42018
R2320 VDD.n719 VDD.n694 1.4005
R2321 VDD.n1660 VDD.n1659 1.3744
R2322 VDD.n1657 VDD.n1656 1.3744
R2323 VDD.n1065 VDD.n1064 1.36849
R2324 VDD.n1573 VDD.n1554 1.35142
R2325 VDD.n2019 VDD.n2018 1.25782
R2326 VDD.t50 VDD.t66 1.24946
R2327 VDD.t47 VDD.t22 1.24946
R2328 VDD.n980 VDD.n932 1.2474
R2329 VDD.n68 VDD.n66 1.23637
R2330 VDD.n128 VDD.n126 1.23637
R2331 VDD.n227 VDD.n225 1.23591
R2332 VDD.n1892 VDD.n1890 1.23591
R2333 VDD.n2022 VDD.n2021 1.19777
R2334 VDD.n1659 VDD.n1658 1.1854
R2335 VDD.n1658 VDD.n1657 1.1854
R2336 VDD.n1920 VDD.n1919 1.17953
R2337 VDD.n1090 VDD.n1089 1.14837
R2338 VDD.n802 VDD.n801 1.1255
R2339 VDD.n724 VDD.n687 1.1255
R2340 VDD.n858 VDD.n857 1.1255
R2341 VDD.n1008 VDD.n1007 1.1255
R2342 VDD.n1071 VDD.n1070 1.1255
R2343 VDD.n1083 VDD.n1082 1.1255
R2344 VDD.n862 VDD.n851 1.12549
R2345 VDD.n1866 VDD.n268 1.11762
R2346 VDD.n1596 VDD.n1595 1.08825
R2347 VDD.n1595 VDD.n434 1.08806
R2348 VDD.n1436 VDD.n479 1.08806
R2349 VDD.n1437 VDD.n1436 1.07146
R2350 VDD.n1919 VDD.n1912 1.06955
R2351 VDD.n1202 VDD.n1201 1.06485
R2352 VDD.n1213 VDD.n1212 1.06485
R2353 VDD.n1198 VDD.n1176 1.06485
R2354 VDD.n1195 VDD.n1194 1.06485
R2355 VDD.n359 VDD.n358 1.06485
R2356 VDD.n1725 VDD.n315 1.06485
R2357 VDD.n1718 VDD.n1717 1.06485
R2358 VDD.n1714 VDD.n1713 1.06485
R2359 VDD.n754 VDD.n741 1.0505
R2360 VDD.n971 VDD.n936 1.0505
R2361 VDD.n1217 VDD.n635 1.01789
R2362 VDD.n613 VDD.n603 1.01789
R2363 VDD.n321 VDD.n320 1.01789
R2364 VDD.n1709 VDD.n272 1.01789
R2365 VDD.n1441 VDD.n1440 0.984049
R2366 VDD.n749 VDD.n741 0.963
R2367 VDD.n983 VDD.n982 0.950899
R2368 VDD.n38 VDD.n37 0.93487
R2369 VDD.n1092 VDD.n1091 0.931466
R2370 VDD.n826 VDD.n825 0.927241
R2371 VDD.n683 VDD.n678 0.92659
R2372 VDD.n933 VDD.n931 0.925561
R2373 VDD.n841 VDD.n684 0.904541
R2374 VDD.n930 VDD.n929 0.899617
R2375 VDD.n797 VDD.n792 0.898206
R2376 VDD.n1003 VDD.n983 0.897926
R2377 VDD.n1012 VDD.n842 0.897926
R2378 VDD.n57 VDD.n22 0.873239
R2379 VDD.n56 VDD.n55 0.847535
R2380 VDD.t31 VDD.t76 0.833139
R2381 VDD.t19 VDD.t31 0.833139
R2382 VDD.t37 VDD.t25 0.833139
R2383 VDD.t28 VDD.t71 0.833139
R2384 VDD.t71 VDD.t16 0.833139
R2385 VDD.n1089 VDD 0.830218
R2386 VDD.n1169 VDD.n1168 0.802674
R2387 VDD.n1208 VDD.n1205 0.802674
R2388 VDD.n1190 VDD.n1187 0.802674
R2389 VDD.n1197 VDD.n1196 0.802674
R2390 VDD.n346 VDD.n336 0.802674
R2391 VDD.n1724 VDD.n1721 0.802674
R2392 VDD.n355 VDD.n327 0.802674
R2393 VDD.n349 VDD.n333 0.802674
R2394 VDD.n119 VDD.n118 0.798761
R2395 VDD.n215 VDD.n214 0.798761
R2396 VDD.n264 VDD.n263 0.795258
R2397 VDD.n566 VDD.n565 0.795217
R2398 VDD.n1013 VDD.n1012 0.792748
R2399 VDD.n1124 VDD.n663 0.746922
R2400 VDD.n667 VDD.n663 0.746686
R2401 VDD.n1116 VDD.n663 0.746686
R2402 VDD.n671 VDD.n663 0.746686
R2403 VDD.n1108 VDD.n663 0.746686
R2404 VDD.n675 VDD.n663 0.746686
R2405 VDD.n1100 VDD.n663 0.746686
R2406 VDD.n1093 VDD.n663 0.746686
R2407 VDD.n46 VDD.n45 0.735716
R2408 VDD.n1300 VDD.n578 0.730547
R2409 VDD.n1310 VDD.n578 0.730547
R2410 VDD.n1344 VDD.n578 0.730547
R2411 VDD.n1658 VDD.n386 0.73031
R2412 VDD.n1658 VDD.n383 0.73031
R2413 VDD.n787 VDD.n786 0.7187
R2414 VDD.n1487 VDD.n1486 0.674731
R2415 VDD.n1323 VDD.n578 0.662176
R2416 VDD.n1658 VDD.n388 0.661938
R2417 VDD.n1869 VDD.n269 0.660673
R2418 VDD.n1307 VDD.n578 0.659239
R2419 VDD.n1658 VDD.n387 0.659
R2420 VDD VDD.n251 0.650002
R2421 VDD.n1595 VDD.n432 0.645651
R2422 VDD VDD.n2 0.642616
R2423 VDD VDD.n152 0.641056
R2424 VDD.n776 VDD.n775 0.6395
R2425 VDD.n993 VDD.n991 0.6395
R2426 VDD.n988 VDD.n986 0.6395
R2427 VDD.n1947 VDD.n1946 0.6395
R2428 VDD.n2001 VDD.n1999 0.6395
R2429 VDD.n265 VDD.n264 0.626871
R2430 VDD.n714 VDD.n694 0.613
R2431 VDD.n1297 VDD.n578 0.60307
R2432 VDD.n1658 VDD.n385 0.602829
R2433 VDD.n2010 VDD.n2009 0.597767
R2434 VDD.n1599 VDD.n1598 0.593699
R2435 VDD.n1870 VDD.n268 0.587674
R2436 VDD VDD.n1927 0.582694
R2437 VDD.n1163 VDD.n1160 0.581587
R2438 VDD.n1172 VDD.n608 0.581587
R2439 VDD.n1225 VDD.n628 0.581587
R2440 VDD.n1175 VDD.n598 0.581587
R2441 VDD.n1690 VDD.n362 0.581587
R2442 VDD.n352 VDD.n278 0.581587
R2443 VDD.n1842 VDD.n297 0.581587
R2444 VDD.n1828 VDD.n1728 0.581587
R2445 VDD.n45 VDD.n43 0.576883
R2446 VDD.n1810 VDD.n1809 0.573969
R2447 VDD.n1553 VDD.n1547 0.569476
R2448 VDD.n1293 VDD.n578 0.553668
R2449 VDD.n1658 VDD.n384 0.553425
R2450 VDD.n22 VDD.n21 0.5405
R2451 VDD.n21 VDD.n20 0.5405
R2452 VDD.n1013 VDD.n841 0.539532
R2453 VDD.n221 VDD.n220 0.539417
R2454 VDD.n164 VDD.n122 0.538543
R2455 VDD.n166 VDD.n120 0.538543
R2456 VDD.n219 VDD.n218 0.536587
R2457 VDD.n1654 VDD.n397 0.536587
R2458 VDD.n404 VDD.n403 0.536587
R2459 VDD.n410 VDD.n409 0.536587
R2460 VDD.n1320 VDD.n1316 0.536587
R2461 VDD.n1306 VDD.n1305 0.536587
R2462 VDD.n1296 VDD.n1295 0.536587
R2463 VDD.n1028 VDD.n1018 0.5255
R2464 VDD.n266 VDD.n265 0.50421
R2465 VDD.n172 VDD.n102 0.502171
R2466 VDD.n191 VDD.n190 0.500214
R2467 VDD.n1570 VDD.n1555 0.495796
R2468 VDD.n2028 VDD.n1932 0.489544
R2469 VDD VDD.n731 0.485717
R2470 VDD VDD.n737 0.485717
R2471 VDD.n71 VDD.n68 0.476034
R2472 VDD.n160 VDD.n128 0.476034
R2473 VDD.n259 VDD.n227 0.475523
R2474 VDD.n1895 VDD.n1892 0.475523
R2475 VDD VDD.n453 0.474784
R2476 VDD.n1217 VDD.n1216 0.467817
R2477 VDD.n324 VDD.n321 0.467817
R2478 VDD.n1193 VDD.n603 0.466777
R2479 VDD.n1712 VDD.n1709 0.466777
R2480 VDD.n81 VDD.n80 0.463032
R2481 VDD.n145 VDD.n144 0.463032
R2482 VDD.n244 VDD.n243 0.463032
R2483 VDD.n1902 VDD.n1901 0.463032
R2484 VDD.n981 VDD.n980 0.462817
R2485 VDD.n9 VDD.n8 0.446529
R2486 VDD.n261 VDD 0.44179
R2487 VDD.n1205 VDD.n1202 0.440717
R2488 VDD.n1725 VDD.n1724 0.440717
R2489 VDD.n1078 VDD.n1019 0.438
R2490 VDD.n120 VDD.n119 0.430935
R2491 VDD.n218 VDD.n215 0.430935
R2492 VDD.n330 VDD.n272 0.430935
R2493 VDD.n1183 VDD.n613 0.430935
R2494 VDD.n1211 VDD.n635 0.430935
R2495 VDD.n320 VDD.n318 0.430935
R2496 VDD.n8 VDD.n7 0.429324
R2497 VDD.n7 VDD.n6 0.429324
R2498 VDD.n1928 VDD.n59 0.428242
R2499 VDD.n162 VDD 0.424686
R2500 VDD.n1212 VDD.n1208 0.421152
R2501 VDD.n1194 VDD.n1193 0.421152
R2502 VDD.n1721 VDD.n1718 0.421152
R2503 VDD.n1713 VDD.n1712 0.421152
R2504 VDD.n2015 VDD.n1971 0.419346
R2505 VDD.n2013 VDD.n1987 0.419346
R2506 VDD.n2011 VDD.n2010 0.419346
R2507 VDD.n1957 VDD.n1952 0.419346
R2508 VDD.n153 VDD.n150 0.419196
R2509 VDD.n252 VDD.n249 0.419196
R2510 VDD.n1876 VDD.n1875 0.419196
R2511 VDD.n1910 VDD.n267 0.419196
R2512 VDD.n1921 VDD.n92 0.419196
R2513 VDD.n91 VDD.n89 0.419196
R2514 VDD.t53 VDD.t88 0.41682
R2515 VDD.t88 VDD.t44 0.41682
R2516 VDD.t63 VDD.t13 0.41682
R2517 VDD.t398 VDD.n601 0.41682
R2518 VDD.t85 VDD.t34 0.41682
R2519 VDD.t58 VDD.t85 0.41682
R2520 VDD.n1375 VDD.n1374 0.405977
R2521 VDD.n1626 VDD.n412 0.405977
R2522 VDD.n1928 VDD 0.40579
R2523 VDD.n1218 VDD.n1217 0.394968
R2524 VDD.n1268 VDD.n603 0.394968
R2525 VDD.n321 VDD.n319 0.394968
R2526 VDD.n1709 VDD.n1708 0.394968
R2527 VDD.n1863 VDD.n272 0.39039
R2528 VDD.n1176 VDD.n1175 0.389848
R2529 VDD.n362 VDD.n359 0.389848
R2530 VDD.n524 VDD.n523 0.389323
R2531 VDD.n1053 VDD.n1052 0.389323
R2532 VDD.n1477 VDD.n1474 0.389323
R2533 VDD.n1992 VDD.n1990 0.389323
R2534 VDD.n1952 VDD.n1951 0.388557
R2535 VDD.n1530 VDD.n1496 0.376152
R2536 VDD.n1531 VDD.n1493 0.376152
R2537 VDD.n542 VDD.n504 0.376152
R2538 VDD.n766 VDD.n765 0.376152
R2539 VDD.n709 VDD.n704 0.376152
R2540 VDD.n975 VDD.n934 0.376152
R2541 VDD.n886 VDD.n882 0.376152
R2542 VDD.n886 VDD.n885 0.376152
R2543 VDD.n1464 VDD.n461 0.376152
R2544 VDD.n1522 VDD.n1506 0.374196
R2545 VDD.n531 VDD.n518 0.374196
R2546 VDD.n500 VDD.n499 0.374196
R2547 VDD.n961 VDD.n946 0.374196
R2548 VDD.n908 VDD.n902 0.374196
R2549 VDD.n908 VDD.n907 0.374196
R2550 VDD.n1060 VDD.n1047 0.374196
R2551 VDD.n471 VDD.n470 0.374196
R2552 VDD.n1540 VDD.n1487 0.372931
R2553 VDD.n1410 VDD.n566 0.359918
R2554 VDD.n1152 VDD.n635 0.358543
R2555 VDD.n1251 VDD.n613 0.358543
R2556 VDD.n320 VDD.n307 0.358543
R2557 VDD.n262 VDD.n261 0.357597
R2558 VDD.n1021 VDD.n1020 0.350287
R2559 VDD.n259 VDD.n258 0.334371
R2560 VDD.n253 VDD.n252 0.334371
R2561 VDD.n263 VDD.n262 0.332919
R2562 VDD.n1200 VDD.n1169 0.327239
R2563 VDD.n356 VDD.n355 0.327239
R2564 VDD.n1187 VDD.n1176 0.323326
R2565 VDD.n1198 VDD.n1197 0.323326
R2566 VDD.n359 VDD.n346 0.323326
R2567 VDD.n358 VDD.n349 0.323326
R2568 VDD.n160 VDD.n159 0.32143
R2569 VDD.n154 VDD.n153 0.32143
R2570 VDD.n163 VDD.n162 0.31864
R2571 VDD.n258 VDD.n257 0.314048
R2572 VDD.n542 VDD.n541 0.312794
R2573 VDD.n1715 VDD.n330 0.311587
R2574 VDD.n1184 VDD.n1183 0.311587
R2575 VDD.n1465 VDD.n1464 0.306039
R2576 VDD.n159 VDD.n158 0.301895
R2577 VDD.n58 VDD.n15 0.3007
R2578 VDD.n255 VDD.n254 0.295177
R2579 VDD.n263 VDD.n207 0.292274
R2580 VDD.n264 VDD.n193 0.292274
R2581 VDD.n265 VDD.n183 0.292274
R2582 VDD.n266 VDD.n182 0.292274
R2583 VDD.n262 VDD.n221 0.292274
R2584 VDD.n1097 VDD.n677 0.292144
R2585 VDD.n1105 VDD.n673 0.292144
R2586 VDD.n1112 VDD.n669 0.292144
R2587 VDD.n1212 VDD.n1211 0.292022
R2588 VDD.n1216 VDD.n1213 0.292022
R2589 VDD.n1194 VDD.n1190 0.292022
R2590 VDD.n1196 VDD.n1195 0.292022
R2591 VDD.n1713 VDD.n336 0.292022
R2592 VDD.n1717 VDD.n324 0.292022
R2593 VDD.n1718 VDD.n318 0.292022
R2594 VDD.n1714 VDD.n333 0.292022
R2595 VDD.n1768 VDD.n1767 0.291683
R2596 VDD.n1780 VDD.n1761 0.291683
R2597 VDD.n1803 VDD.n1754 0.291683
R2598 VDD.n1120 VDD.n665 0.288544
R2599 VDD.n1793 VDD.n1786 0.288083
R2600 VDD.n1770 VDD.n1766 0.284207
R2601 VDD.n156 VDD.n155 0.283756
R2602 VDD.n1168 VDD.n636 0.278326
R2603 VDD.n1716 VDD.n327 0.278326
R2604 VDD.n1202 VDD.n1163 0.272457
R2605 VDD.n1201 VDD.n628 0.272457
R2606 VDD.n315 VDD.n297 0.272457
R2607 VDD.n1728 VDD.n1725 0.272457
R2608 VDD.n1199 VDD.n1172 0.266587
R2609 VDD.n357 VDD.n352 0.266587
R2610 VDD.n1635 VDD.n411 0.266523
R2611 VDD.n1340 VDD.n1294 0.26536
R2612 VDD.n392 VDD.n390 0.264528
R2613 VDD.n1318 VDD.n1317 0.263373
R2614 VDD.n831 VDD.n721 0.263
R2615 VDD.n406 VDD.n405 0.262011
R2616 VDD.n1299 VDD.n1298 0.260887
R2617 VDD.n1648 VDD.n398 0.257984
R2618 VDD.n1327 VDD.n1308 0.257526
R2619 VDD.n1601 VDD.n1600 0.25389
R2620 VDD.n1027 VDD.n1026 0.253803
R2621 VDD.n1092 VDD.n657 0.252505
R2622 VDD.n789 VDD.n788 0.252091
R2623 VDD.n1912 VDD.n1911 0.251788
R2624 VDD.n1440 VDD.n475 0.248505
R2625 VDD.n82 VDD.n77 0.246576
R2626 VDD.n143 VDD.n140 0.246576
R2627 VDD.n242 VDD.n239 0.246576
R2628 VDD.n1900 VDD.n1887 0.246576
R2629 VDD VDD.n81 0.245437
R2630 VDD.n144 VDD 0.245437
R2631 VDD.n243 VDD 0.245437
R2632 VDD.n1901 VDD 0.245437
R2633 VDD.n1614 VDD.n425 0.238241
R2634 VDD.n1394 VDD.n1393 0.238069
R2635 VDD.n1392 VDD.n574 0.237294
R2636 VDD.n1513 VDD.n1511 0.237044
R2637 VDD.n954 VDD.n952 0.237044
R2638 VDD.n1445 VDD.n1444 0.237044
R2639 VDD.n708 VDD.n707 0.233429
R2640 VDD.n541 VDD.n507 0.229786
R2641 VDD.n796 VDD.n793 0.229786
R2642 VDD.n850 VDD.n849 0.229786
R2643 VDD.n1465 VDD.n460 0.229786
R2644 VDD.n169 VDD.n107 0.228829
R2645 VDD.n1911 VDD.n266 0.228403
R2646 VDD.n1359 VDD.n1358 0.221442
R2647 VDD.n1563 VDD.n1560 0.220495
R2648 VDD VDD.n2028 0.218882
R2649 VDD.n982 VDD.n930 0.217222
R2650 VDD.n1987 VDD 0.215115
R2651 VDD.n1128 VDD.n1127 0.209826
R2652 VDD.n1812 VDD.n1746 0.209826
R2653 VDD.n163 VDD.n121 0.209105
R2654 VDD.n176 VDD.n175 0.208053
R2655 VDD.n1911 VDD.n1910 0.202732
R2656 VDD.n121 VDD.n107 0.19985
R2657 VDD.n1772 VDD.n1771 0.183919
R2658 VDD.n955 VDD.n949 0.182274
R2659 VDD.n1954 VDD.n1953 0.182274
R2660 VDD.n1512 VDD.n1510 0.182033
R2661 VDD.n539 VDD.n538 0.182033
R2662 VDD.n560 VDD.n492 0.182033
R2663 VDD.n1447 VDD.n1446 0.182033
R2664 VDD.n1468 VDD.n1467 0.182033
R2665 VDD.n1625 VDD.n414 0.178585
R2666 VDD.n1351 VDD.n1347 0.17667
R2667 VDD.n1616 VDD.n378 0.176655
R2668 VDD.n1390 VDD.n575 0.176655
R2669 VDD.n1950 VDD 0.174184
R2670 VDD VDD.n1949 0.174184
R2671 VDD.n2008 VDD.n2006 0.174184
R2672 VDD.n565 VDD.n561 0.174122
R2673 VDD.n2003 VDD 0.173395
R2674 VDD.n1376 VDD.n1291 0.17241
R2675 VDD.n1674 VDD.n372 0.17241
R2676 VDD.n1668 VDD.n1667 0.171399
R2677 VDD.n1284 VDD.n582 0.171399
R2678 VDD.n1640 VDD.n1639 0.163357
R2679 VDD.n1336 VDD.n1335 0.163357
R2680 VDD.n1951 VDD.n1950 0.158395
R2681 VDD.n2009 VDD.n2008 0.158395
R2682 VDD.n1668 VDD.n367 0.157434
R2683 VDD.n257 VDD.n256 0.157274
R2684 VDD.n1285 VDD.n1284 0.15672
R2685 VDD VDD.n255 0.156548
R2686 VDD.n1921 VDD.n1920 0.153813
R2687 VDD.n1129 VDD.n651 0.153197
R2688 VDD.n1814 VDD.n1813 0.153197
R2689 VDD.n158 VDD.n157 0.151198
R2690 VDD VDD.n156 0.1505
R2691 VDD.n1766 VDD.n1738 0.146319
R2692 VDD.n1635 VDD.n1634 0.146214
R2693 VDD.n1341 VDD.n1340 0.146214
R2694 VDD.n1129 VDD.n1128 0.146118
R2695 VDD.n1813 VDD.n1812 0.146118
R2696 VDD.n1135 VDD.n657 0.146022
R2697 VDD.n928 VDD.n926 0.143441
R2698 VDD.n1385 VDD.n581 0.143084
R2699 VDD.n1636 VDD.n410 0.143
R2700 VDD.n1376 VDD.n1375 0.142944
R2701 VDD.n412 VDD.n372 0.142944
R2702 VDD.n1352 VDD.n1351 0.142202
R2703 VDD.n416 VDD.n414 0.142202
R2704 VDD.n1665 VDD.n1664 0.142073
R2705 VDD.n1339 VDD.n1296 0.141929
R2706 VDD.n1895 VDD.n1894 0.141797
R2707 VDD.n1903 VDD.n1876 0.141797
R2708 VDD.n1664 VDD.n378 0.141062
R2709 VDD.n581 VDD.n575 0.141062
R2710 VDD.n1652 VDD.n1649 0.140857
R2711 VDD.n1326 VDD.n1309 0.140857
R2712 VDD.n2023 VDD.n1938 0.140627
R2713 VDD.n1127 VDD.n660 0.14038
R2714 VDD.n1787 VDD.n1746 0.14038
R2715 VDD.n1653 VDD.n1652 0.139786
R2716 VDD.n1634 VDD.n1631 0.139786
R2717 VDD.n1341 VDD.n1292 0.139786
R2718 VDD.n1321 VDD.n1309 0.139786
R2719 VDD VDD.n787 0.139763
R2720 VDD.n1440 VDD.n1439 0.139295
R2721 VDD.n1919 VDD.n1918 0.1385
R2722 VDD.n1439 VDD.n476 0.138211
R2723 VDD.n1572 VDD.n1570 0.138211
R2724 VDD.n1648 VDD.n1647 0.137643
R2725 VDD.n1328 VDD.n1327 0.137643
R2726 VDD.n1675 VDD.n1674 0.137017
R2727 VDD.n1291 VDD.n1290 0.136006
R2728 VDD.n2003 VDD.n2002 0.1355
R2729 VDD.n2017 VDD.n1959 0.1355
R2730 VDD.n1949 VDD.n1948 0.134711
R2731 VDD.n1598 VDD.n430 0.133873
R2732 VDD.n1592 VDD.n1591 0.133873
R2733 VDD.n1589 VDD.n1587 0.133873
R2734 VDD.n1585 VDD.n1583 0.133873
R2735 VDD.n1581 VDD.n1579 0.133873
R2736 VDD.n1577 VDD.n1575 0.133873
R2737 VDD.n1433 VDD.n476 0.133873
R2738 VDD.n1432 VDD.n1430 0.133873
R2739 VDD.n1428 VDD.n1426 0.133873
R2740 VDD.n1424 VDD.n1422 0.133873
R2741 VDD.n1420 VDD.n1418 0.133873
R2742 VDD.n1416 VDD.n1414 0.133873
R2743 VDD.n1412 VDD.n1410 0.133873
R2744 VDD.n1603 VDD.n1602 0.133833
R2745 VDD.n428 VDD.n426 0.133833
R2746 VDD.n1613 VDD.n426 0.133833
R2747 VDD.n1616 VDD.n1615 0.133833
R2748 VDD.n1391 VDD.n1390 0.133833
R2749 VDD.n1397 VDD.n1396 0.133833
R2750 VDD.n1396 VDD.n1395 0.133833
R2751 VDD.n1406 VDD.n568 0.133833
R2752 VDD.n1894 VDD.n1879 0.133196
R2753 VDD.n1662 VDD.n377 0.133132
R2754 VDD.n823 VDD 0.131587
R2755 VDD.n1369 VDD.n1352 0.131498
R2756 VDD.n417 VDD.n416 0.13055
R2757 VDD.n1328 VDD.n1306 0.130143
R2758 VDD.n822 VDD 0.12963
R2759 VDD.n1122 VDD.n660 0.129536
R2760 VDD.n1122 VDD.n1121 0.129536
R2761 VDD.n1119 VDD.n666 0.129536
R2762 VDD.n1114 VDD.n666 0.129536
R2763 VDD.n1114 VDD.n1113 0.129536
R2764 VDD.n1111 VDD.n670 0.129536
R2765 VDD.n1106 VDD.n670 0.129536
R2766 VDD.n1104 VDD.n1103 0.129536
R2767 VDD.n1103 VDD.n674 0.129536
R2768 VDD.n1098 VDD.n674 0.129536
R2769 VDD.n1096 VDD.n1095 0.129536
R2770 VDD.n1770 VDD.n1769 0.129536
R2771 VDD.n1764 VDD.n1762 0.129536
R2772 VDD.n1778 VDD.n1762 0.129536
R2773 VDD.n1779 VDD.n1778 0.129536
R2774 VDD.n1781 VDD.n1753 0.129536
R2775 VDD.n1804 VDD.n1753 0.129536
R2776 VDD.n1802 VDD.n1801 0.129536
R2777 VDD.n1801 VDD.n1755 0.129536
R2778 VDD.n1794 VDD.n1755 0.129536
R2779 VDD.n1792 VDD.n1791 0.129536
R2780 VDD.n1791 VDD.n1787 0.129536
R2781 VDD.n973 VDD.n936 0.129141
R2782 VDD.n1647 VDD.n404 0.129071
R2783 VDD.n1959 VDD.n1958 0.128577
R2784 VDD.n1352 VDD.n1350 0.128395
R2785 VDD.n416 VDD.n415 0.128395
R2786 VDD.n1591 VDD.n1589 0.127367
R2787 VDD.n1587 VDD.n1585 0.127367
R2788 VDD.n1583 VDD.n1581 0.127367
R2789 VDD.n1579 VDD.n1577 0.127367
R2790 VDD.n1097 VDD.n1096 0.127367
R2791 VDD.n1433 VDD.n1432 0.127367
R2792 VDD.n1430 VDD.n1428 0.127367
R2793 VDD.n1426 VDD.n1424 0.127367
R2794 VDD.n1422 VDD.n1420 0.127367
R2795 VDD.n1418 VDD.n1416 0.127367
R2796 VDD.n1769 VDD.n1768 0.127367
R2797 VDD.n2020 VDD.n2019 0.12616
R2798 VDD.n925 VDD.n848 0.126143
R2799 VDD.n1905 VDD.n1904 0.12521
R2800 VDD.n1592 VDD.n430 0.124114
R2801 VDD.n1414 VDD.n1412 0.124114
R2802 VDD.n1368 VDD.n1367 0.123227
R2803 VDD.n1367 VDD.n1353 0.123227
R2804 VDD.n1361 VDD.n1360 0.123227
R2805 VDD.n1360 VDD.n475 0.123227
R2806 VDD.n1559 VDD.n1555 0.123227
R2807 VDD.n1564 VDD.n1559 0.123227
R2808 VDD.n1562 VDD.n1561 0.123227
R2809 VDD.n1561 VDD.n419 0.123227
R2810 VDD.n1112 VDD.n1111 0.12303
R2811 VDD.n1804 VDD.n1803 0.12303
R2812 VDD.n1359 VDD.n1353 0.122205
R2813 VDD.n1563 VDD.n1562 0.122205
R2814 VDD.n1142 VDD.n651 0.120837
R2815 VDD.n1143 VDD.n1142 0.120837
R2816 VDD.n1144 VDD.n1143 0.120837
R2817 VDD.n1144 VDD.n637 0.120837
R2818 VDD.n1159 VDD.n638 0.120837
R2819 VDD.n638 VDD.n629 0.120837
R2820 VDD.n1224 VDD.n629 0.120837
R2821 VDD.n1227 VDD.n1226 0.120837
R2822 VDD.n1227 VDD.n618 0.120837
R2823 VDD.n1240 VDD.n618 0.120837
R2824 VDD.n1241 VDD.n1240 0.120837
R2825 VDD.n1243 VDD.n1241 0.120837
R2826 VDD.n1243 VDD.n1242 0.120837
R2827 VDD.n1258 VDD.n1257 0.120837
R2828 VDD.n1260 VDD.n1258 0.120837
R2829 VDD.n1260 VDD.n1259 0.120837
R2830 VDD.n1275 VDD.n1274 0.120837
R2831 VDD.n1276 VDD.n1275 0.120837
R2832 VDD.n1276 VDD.n589 0.120837
R2833 VDD.n1290 VDD.n589 0.120837
R2834 VDD.n1676 VDD.n1675 0.120837
R2835 VDD.n1676 VDD.n363 0.120837
R2836 VDD.n1688 VDD.n363 0.120837
R2837 VDD.n1689 VDD.n1688 0.120837
R2838 VDD.n1702 VDD.n1701 0.120837
R2839 VDD.n1701 VDD.n1700 0.120837
R2840 VDD.n1700 VDD.n1691 0.120837
R2841 VDD.n1858 VDD.n1857 0.120837
R2842 VDD.n1857 VDD.n1856 0.120837
R2843 VDD.n1856 VDD.n279 0.120837
R2844 VDD.n294 VDD.n279 0.120837
R2845 VDD.n1844 VDD.n294 0.120837
R2846 VDD.n1844 VDD.n1843 0.120837
R2847 VDD.n1841 VDD.n298 0.120837
R2848 VDD.n314 VDD.n298 0.120837
R2849 VDD.n1829 VDD.n314 0.120837
R2850 VDD.n1827 VDD.n1826 0.120837
R2851 VDD.n1826 VDD.n1729 0.120837
R2852 VDD.n1745 VDD.n1729 0.120837
R2853 VDD.n1814 VDD.n1745 0.120837
R2854 VDD.n1407 VDD.n566 0.119037
R2855 VDD.n391 VDD.n376 0.117286
R2856 VDD.n1644 VDD.n1643 0.117286
R2857 VDD.n1631 VDD.n1630 0.117286
R2858 VDD.n1346 VDD.n1292 0.117286
R2859 VDD.n1332 VDD.n1331 0.117286
R2860 VDD.n1383 VDD.n583 0.117286
R2861 VDD.n202 VDD.n201 0.115972
R2862 VDD.n192 VDD.n191 0.115972
R2863 VDD.n1937 VDD.n1936 0.115087
R2864 VDD.n221 VDD.n219 0.113142
R2865 VDD.n1370 VDD.n1369 0.113
R2866 VDD.n1624 VDD.n417 0.111977
R2867 VDD.n1160 VDD.n1159 0.110725
R2868 VDD.n191 VDD.n183 0.109745
R2869 VDD.n91 VDD.n90 0.109735
R2870 VDD.n71 VDD.n70 0.109735
R2871 VDD.n1829 VDD.n1828 0.109713
R2872 VDD.n1666 VDD.n376 0.108714
R2873 VDD.n2015 VDD.n2014 0.108385
R2874 VDD.n2024 VDD.n2023 0.108044
R2875 VDD.n1320 VDD.n1319 0.107643
R2876 VDD.n1384 VDD.n1383 0.107643
R2877 VDD.n980 VDD.n979 0.106797
R2878 VDD.n1655 VDD.n1654 0.106571
R2879 VDD.n1702 VDD.n1690 0.103646
R2880 VDD.n70 VDD.n63 0.103086
R2881 VDD.n1259 VDD.n598 0.102635
R2882 VDD.n1865 VDD.n1864 0.101533
R2883 VDD.n1084 VDD.n683 0.101088
R2884 VDD.n1136 VDD.n1135 0.1005
R2885 VDD.n1819 VDD.n1738 0.1005
R2886 VDD.n207 VDD.n206 0.0989906
R2887 VDD.n2013 VDD.n2012 0.0985769
R2888 VDD.n1615 VDD.n1614 0.0971667
R2889 VDD.n1392 VDD.n1391 0.0971667
R2890 VDD.n198 VDD.n193 0.0964434
R2891 VDD.n260 VDD.n259 0.0955806
R2892 VDD.n392 VDD.n391 0.0947857
R2893 VDD.n1318 VDD.n583 0.0947857
R2894 VDD.n1385 VDD.n1384 0.0945449
R2895 VDD.n1603 VDD.n1599 0.0938198
R2896 VDD.n1407 VDD.n1406 0.0938198
R2897 VDD.n1666 VDD.n1665 0.0935337
R2898 VDD.n1910 VDD.n1909 0.0920358
R2899 VDD.n161 VDD.n160 0.0918953
R2900 VDD.n12 VDD.n11 0.0914091
R2901 VDD.n11 VDD.n10 0.0914091
R2902 VDD.n36 VDD.n35 0.0914091
R2903 VDD.n35 VDD.n34 0.0914091
R2904 VDD.n34 VDD.n33 0.0914091
R2905 VDD.n33 VDD.n32 0.0914091
R2906 VDD.n32 VDD.n31 0.0914091
R2907 VDD.n31 VDD.n30 0.0914091
R2908 VDD VDD.n14 0.0900455
R2909 VDD.n777 VDD.n776 0.0893158
R2910 VDD.n994 VDD.n988 0.0893158
R2911 VDD.n994 VDD.n993 0.0893158
R2912 VDD.n1948 VDD.n1947 0.0893158
R2913 VDD.n2002 VDD.n2001 0.0893158
R2914 VDD.n1374 VDD.n1347 0.0884545
R2915 VDD.n1066 VDD.n1040 0.088
R2916 VDD.n1257 VDD.n608 0.0874663
R2917 VDD.n1626 VDD.n1625 0.0874318
R2918 VDD.n1936 VDD.n1933 0.0865195
R2919 VDD.n1691 VDD.n278 0.0864551
R2920 VDD.n1601 VDD.n428 0.0860556
R2921 VDD.n1395 VDD.n1394 0.0860556
R2922 VDD.n1681 VDD.n367 0.0855
R2923 VDD.n1682 VDD.n1681 0.0855
R2924 VDD.n1683 VDD.n1682 0.0855
R2925 VDD.n1683 VDD.n337 0.0855
R2926 VDD.n1707 VDD.n338 0.0855
R2927 VDD.n1694 VDD.n338 0.0855
R2928 VDD.n1694 VDD.n270 0.0855
R2929 VDD.n1137 VDD.n1136 0.0855
R2930 VDD.n1137 VDD.n648 0.0855
R2931 VDD.n1150 VDD.n648 0.0855
R2932 VDD.n1151 VDD.n1150 0.0855
R2933 VDD.n1154 VDD.n1153 0.0855
R2934 VDD.n1153 VDD.n634 0.0855
R2935 VDD.n1219 VDD.n634 0.0855
R2936 VDD.n1233 VDD.n623 0.0855
R2937 VDD.n1234 VDD.n1233 0.0855
R2938 VDD.n1235 VDD.n614 0.0855
R2939 VDD.n1249 VDD.n614 0.0855
R2940 VDD.n1250 VDD.n1249 0.0855
R2941 VDD.n1252 VDD.n604 0.0855
R2942 VDD.n1266 VDD.n604 0.0855
R2943 VDD.n1267 VDD.n1266 0.0855
R2944 VDD.n1269 VDD.n594 0.0855
R2945 VDD.n1282 VDD.n594 0.0855
R2946 VDD.n1283 VDD.n1282 0.0855
R2947 VDD.n1285 VDD.n1283 0.0855
R2948 VDD.n287 VDD.n271 0.0855
R2949 VDD.n1851 VDD.n287 0.0855
R2950 VDD.n1850 VDD.n1849 0.0855
R2951 VDD.n1849 VDD.n288 0.0855
R2952 VDD.n1836 VDD.n306 0.0855
R2953 VDD.n1836 VDD.n1835 0.0855
R2954 VDD.n1835 VDD.n1834 0.0855
R2955 VDD.n1737 VDD.n1736 0.0855
R2956 VDD.n1821 VDD.n1737 0.0855
R2957 VDD.n1821 VDD.n1820 0.0855
R2958 VDD.n1820 VDD.n1819 0.0855
R2959 VDD.n173 VDD.n172 0.0853962
R2960 VDD.n1121 VDD.n1120 0.0850783
R2961 VDD.n1793 VDD.n1792 0.0850783
R2962 VDD.n1154 VDD.n1152 0.0847857
R2963 VDD.n1834 VDD.n307 0.0840714
R2964 VDD.n780 VDD 0.0836933
R2965 VDD.n252 VDD 0.0832419
R2966 VDD.n1575 VDD.n1573 0.0818253
R2967 VDD.n172 VDD.n171 0.0817389
R2968 VDD.n171 VDD.n170 0.0817389
R2969 VDD.n206 VDD 0.0811604
R2970 VDD.n1842 VDD.n1841 0.0803876
R2971 VDD.n153 VDD 0.0800349
R2972 VDD VDD.n1915 0.0798636
R2973 VDD.n1225 VDD.n1224 0.0793764
R2974 VDD.n1004 VDD.n844 0.0790106
R2975 VDD.n1917 VDD 0.0778182
R2976 VDD.n995 VDD 0.0774922
R2977 VDD.n1667 VDD.n1666 0.0773539
R2978 VDD.n1384 VDD.n582 0.0773539
R2979 VDD.n1640 VDD.n406 0.0765714
R2980 VDD.n1335 VDD.n1299 0.0765714
R2981 VDD VDD.n1921 0.0760145
R2982 VDD.n1605 VDD.n1604 0.0752312
R2983 VDD.n10 VDD.n9 0.0750455
R2984 VDD.n1405 VDD.n567 0.074985
R2985 VDD.n1106 VDD.n1105 0.0742349
R2986 VDD.n1781 VDD.n1780 0.0742349
R2987 VDD.n928 VDD.n927 0.07388
R2988 VDD.n1573 VDD.n1572 0.0731506
R2989 VDD.n800 VDD.n769 0.0717174
R2990 VDD.n799 VDD.n798 0.0717174
R2991 VDD.n1524 VDD.n1497 0.0714756
R2992 VDD.n1533 VDD.n1488 0.0714756
R2993 VDD.n529 VDD.n520 0.0714756
R2994 VDD.n548 VDD.n547 0.0714756
R2995 VDD.n969 VDD.n968 0.0714756
R2996 VDD.n1051 VDD.n1048 0.0714756
R2997 VDD.n1458 VDD.n462 0.0714756
R2998 VDD.n1479 VDD.n1478 0.0714756
R2999 VDD.n1541 VDD.n444 0.0714756
R3000 VDD.n1981 VDD.n1980 0.0714756
R3001 VDD.n1006 VDD.n1005 0.0714615
R3002 VDD.n1523 VDD 0.0713871
R3003 VDD VDD.n530 0.0713871
R3004 VDD.n549 VDD 0.0713871
R3005 VDD VDD.n938 0.0713871
R3006 VDD VDD.n1059 0.0713871
R3007 VDD.n1457 VDD 0.0713871
R3008 VDD.n1521 VDD.n1507 0.0709032
R3009 VDD.n1515 VDD.n1514 0.0709032
R3010 VDD.n510 VDD.n508 0.0709032
R3011 VDD.n532 VDD.n513 0.0709032
R3012 VDD.n557 VDD.n491 0.0709032
R3013 VDD.n556 VDD.n555 0.0709032
R3014 VDD.n953 VDD.n947 0.0709032
R3015 VDD.n960 VDD.n959 0.0709032
R3016 VDD.n1449 VDD.n1448 0.0709032
R3017 VDD.n1451 VDD.n1450 0.0709032
R3018 VDD.n457 VDD.n454 0.0709032
R3019 VDD.n1061 VDD.n1039 0.0701774
R3020 VDD.n1529 VDD.n1497 0.0692805
R3021 VDD.n1524 VDD.n1523 0.0692805
R3022 VDD.n1533 VDD.n1532 0.0692805
R3023 VDD.n1539 VDD.n1488 0.0692805
R3024 VDD.n530 VDD.n529 0.0692805
R3025 VDD.n524 VDD.n520 0.0692805
R3026 VDD.n549 VDD.n548 0.0692805
R3027 VDD.n547 VDD.n543 0.0692805
R3028 VDD.n968 VDD.n938 0.0692805
R3029 VDD.n1059 VDD.n1048 0.0692805
R3030 VDD.n1053 VDD.n1051 0.0692805
R3031 VDD.n1458 VDD.n1457 0.0692805
R3032 VDD.n1463 VDD.n462 0.0692805
R3033 VDD.n1479 VDD.n448 0.0692805
R3034 VDD.n1478 VDD.n1477 0.0692805
R3035 VDD.n1541 VDD 0.0692805
R3036 VDD.n1995 VDD.n1992 0.0692805
R3037 VDD.n1977 VDD.n1974 0.0692805
R3038 VDD VDD.n1981 0.0692805
R3039 VDD.n1932 VDD.n1929 0.0692083
R3040 VDD.n1515 VDD.n1507 0.0687258
R3041 VDD.n1514 VDD.n1513 0.0687258
R3042 VDD.n540 VDD.n508 0.0687258
R3043 VDD.n513 VDD.n510 0.0687258
R3044 VDD.n561 VDD.n491 0.0687258
R3045 VDD.n557 VDD.n556 0.0687258
R3046 VDD.n954 VDD.n953 0.0687258
R3047 VDD.n959 VDD.n947 0.0687258
R3048 VDD.n1451 VDD.n1449 0.0687258
R3049 VDD.n1466 VDD.n457 0.0687258
R3050 VDD.n2018 VDD.n2017 0.0685545
R3051 VDD.n1252 VDD.n1251 0.0683571
R3052 VDD.n174 VDD.n173 0.0676691
R3053 VDD.n2022 VDD.n1939 0.0669557
R3054 VDD.n828 VDD.n723 0.0669486
R3055 VDD.n827 VDD.n826 0.0669486
R3056 VDD.n1906 VDD.n1879 0.0668481
R3057 VDD.n1386 VDD.n579 0.0668158
R3058 VDD VDD.n1905 0.066541
R3059 VDD.n1708 VDD.n1707 0.0662143
R3060 VDD.n1268 VDD.n1267 0.0662143
R3061 VDD.n839 VDD.n838 0.0661075
R3062 VDD.n840 VDD.n685 0.0661075
R3063 VDD.n780 VDD.n777 0.0647857
R3064 VDD.n1010 VDD.n1009 0.0646489
R3065 VDD.n170 VDD.n169 0.0643765
R3066 VDD.n2011 VDD.n1996 0.0639615
R3067 VDD.n2013 VDD.n1986 0.0639615
R3068 VDD.n2015 VDD.n1970 0.0639615
R3069 VDD.n1957 VDD.n1956 0.0639615
R3070 VDD.n1522 VDD.n1521 0.0629194
R3071 VDD.n532 VDD.n531 0.0629194
R3072 VDD.n555 VDD.n500 0.0629194
R3073 VDD.n961 VDD.n960 0.0629194
R3074 VDD.n1061 VDD.n1060 0.0629194
R3075 VDD.n1450 VDD.n471 0.0629194
R3076 VDD VDD.n1971 0.0616538
R3077 VDD.n995 VDD.n994 0.0606172
R3078 VDD.n970 VDD.n969 0.0605
R3079 VDD.n1487 VDD.n448 0.0605
R3080 VDD.n164 VDD.n163 0.0603822
R3081 VDD.n1935 VDD.n1934 0.0593952
R3082 VDD.n1011 VDD.n843 0.0584808
R3083 VDD VDD.n182 0.0582358
R3084 VDD.n1986 VDD.n1977 0.0561098
R3085 VDD.n1105 VDD.n1104 0.0558012
R3086 VDD.n1780 VDD.n1779 0.0558012
R3087 VDD VDD.n1540 0.055378
R3088 VDD.n1956 VDD.n1955 0.055378
R3089 VDD.n167 VDD.n107 0.0549355
R3090 VDD.n165 VDD.n121 0.0542097
R3091 VDD.n1927 VDD.n60 0.0539301
R3092 VDD.n165 VDD.n164 0.0538628
R3093 VDD.n1037 VDD.n1036 0.0534412
R3094 VDD.n1034 VDD.n1015 0.0534412
R3095 VDD.n1213 VDD.n636 0.0533261
R3096 VDD.n1717 VDD.n1716 0.0533261
R3097 VDD.n168 VDD.n167 0.0530664
R3098 VDD.n1375 VDD.n1346 0.053
R3099 VDD.n1553 VDD.n444 0.0524512
R3100 VDD.n182 VDD.n181 0.0522925
R3101 VDD.n1630 VDD.n412 0.0519286
R3102 VDD.n59 VDD.n14 0.0518636
R3103 VDD.n771 VDD.n770 0.0509
R3104 VDD.n1002 VDD.n845 0.0504219
R3105 VDD.n1487 VDD.n454 0.0498548
R3106 VDD.n1219 VDD.n1218 0.0497857
R3107 VDD.n319 VDD.n306 0.0497857
R3108 VDD.n1851 VDD 0.0483571
R3109 VDD.n1602 VDD.n1601 0.0482778
R3110 VDD.n1394 VDD.n568 0.0482778
R3111 VDD.n1235 VDD 0.0462143
R3112 VDD.n789 VDD.n771 0.0458103
R3113 VDD.n1120 VDD.n1119 0.0449578
R3114 VDD.n1794 VDD.n1793 0.0449578
R3115 VDD.n179 VDD 0.0440029
R3116 VDD.n1226 VDD.n1225 0.0419607
R3117 VDD.n1868 VDD.n268 0.0414381
R3118 VDD.n1864 VDD.n270 0.0412143
R3119 VDD.n1643 VDD.n406 0.0412143
R3120 VDD.n1636 VDD.n1635 0.0412143
R3121 VDD.n1340 VDD.n1339 0.0412143
R3122 VDD.n1332 VDD.n1299 0.0412143
R3123 VDD.n1080 VDD.n1079 0.0411452
R3124 VDD.n1843 VDD.n1842 0.0409494
R3125 VDD.n1086 VDD.n681 0.0408043
R3126 VDD.n1896 VDD.n1895 0.0407389
R3127 VDD.n1920 VDD.n179 0.0401282
R3128 VDD VDD.n1234 0.0397857
R3129 VDD.n1095 VDD.n1092 0.0395361
R3130 VDD.n1091 VDD 0.0393983
R3131 VDD.n175 VDD.n174 0.0391413
R3132 VDD VDD.n1850 0.0376429
R3133 VDD.n928 VDD.n848 0.0375588
R3134 VDD.n1445 VDD.n1441 0.0375161
R3135 VDD.n1614 VDD.n1613 0.0371667
R3136 VDD.n1397 VDD.n1392 0.0371667
R3137 VDD.n1864 VDD.n271 0.0369286
R3138 VDD.n565 VDD.n564 0.0369005
R3139 VDD.n998 VDD.n997 0.0367109
R3140 VDD.n1918 VDD.n1917 0.0363784
R3141 VDD.n1625 VDD.n1624 0.0362955
R3142 VDD.n1218 VDD.n623 0.0362143
R3143 VDD.n319 VDD.n288 0.0362143
R3144 VDD.n891 VDD.n876 0.0359878
R3145 VDD VDD.n897 0.0359436
R3146 VDD.n873 VDD.n870 0.0357016
R3147 VDD.n918 VDD.n917 0.0357016
R3148 VDD.n1927 VDD.n63 0.0356451
R3149 VDD VDD.n1876 0.0355171
R3150 VDD.n1912 VDD.n181 0.0353113
R3151 VDD VDD.n198 0.0353113
R3152 VDD.n1370 VDD.n1347 0.0352727
R3153 VDD.n891 VDD.n887 0.0348902
R3154 VDD.n897 VDD.n876 0.0348902
R3155 VDD.n1858 VDD.n278 0.034882
R3156 VDD.n1654 VDD.n1653 0.0347857
R3157 VDD.n917 VDD.n870 0.0346129
R3158 VDD.n860 VDD.n859 0.0340503
R3159 VDD.n1242 VDD.n608 0.0338708
R3160 VDD.n1199 VDD.n1198 0.0337609
R3161 VDD.n358 VDD.n357 0.0337609
R3162 VDD.n1321 VDD.n1320 0.0337143
R3163 VDD.n855 VDD.n847 0.0335178
R3164 VDD.n1012 VDD.n1011 0.0331389
R3165 VDD.n2012 VDD.n2011 0.0328077
R3166 VDD.n1970 VDD.n1969 0.0326951
R3167 VDD.n1005 VDD.n983 0.0322736
R3168 VDD.n908 VDD.n873 0.0317097
R3169 VDD.n1448 VDD.n1441 0.0317097
R3170 VDD.n72 VDD.n71 0.0316082
R3171 VDD.n1996 VDD.n1995 0.0305
R3172 VDD.n2014 VDD.n2013 0.0305
R3173 VDD.n1010 VDD.n842 0.0301809
R3174 VDD.n792 VDD.n769 0.0299176
R3175 VDD.n1004 VDD.n1003 0.0292234
R3176 VDD.n1008 VDD.n844 0.0292234
R3177 VDD.n1009 VDD.n1008 0.0292234
R3178 VDD.n1372 VDD.n1371 0.0291956
R3179 VDD.n1357 VDD.n1356 0.0291956
R3180 VDD.n1567 VDD.n1556 0.0291956
R3181 VDD.n1623 VDD.n413 0.0291956
R3182 VDD.n167 VDD.n166 0.0291726
R3183 VDD.n813 VDD.n756 0.0289211
R3184 VDD.n812 VDD.n811 0.0289211
R3185 VDD.n39 VDD.n38 0.028625
R3186 VDD.n166 VDD.n165 0.0283761
R3187 VDD.n1084 VDD.n1083 0.0278529
R3188 VDD.n1070 VDD.n1037 0.0278529
R3189 VDD.n1927 VDD 0.0277903
R3190 VDD.n861 VDD.n854 0.0277596
R3191 VDD.n2016 VDD.n2015 0.0276154
R3192 VDD VDD.n91 0.0275712
R3193 VDD.n856 VDD.n846 0.0273269
R3194 VDD.n1554 VDD.n443 0.0270909
R3195 VDD.n724 VDD.n685 0.0265748
R3196 VDD.n1007 VDD.n1006 0.0264615
R3197 VDD.n1007 VDD.n843 0.0264615
R3198 VDD.n54 VDD.n48 0.026375
R3199 VDD.n827 VDD.n724 0.0257336
R3200 VDD.n810 VDD.n759 0.0256417
R3201 VDD.n918 VDD.n852 0.0251774
R3202 VDD.n1087 VDD.n680 0.0247707
R3203 VDD.n798 VDD.n797 0.0247609
R3204 VDD.n1201 VDD.n1200 0.0239783
R3205 VDD.n801 VDD.n800 0.0239783
R3206 VDD.n356 VDD.n315 0.0239783
R3207 VDD.n1866 VDD.n1865 0.0237036
R3208 VDD.n864 VDD.n863 0.0235488
R3209 VDD.n822 VDD.n732 0.0234555
R3210 VDD.n1083 VDD.n1014 0.0234412
R3211 VDD.n1655 VDD.n392 0.023
R3212 VDD.n1336 VDD.n1296 0.023
R3213 VDD.n1319 VDD.n1318 0.023
R3214 VDD.n836 VDD.n688 0.0227267
R3215 VDD.n1072 VDD.n1071 0.0225588
R3216 VDD.n1069 VDD.n1035 0.0225588
R3217 VDD.n709 VDD.n708 0.0223623
R3218 VDD.n1639 VDD.n410 0.0219286
R3219 VDD.n743 VDD.n742 0.0216336
R3220 VDD.n841 VDD.n840 0.0206869
R3221 VDD.n1980 VDD.n1970 0.0202561
R3222 VDD.n768 VDD.n764 0.0200652
R3223 VDD.n802 VDD.n767 0.0200652
R3224 VDD.n1195 VDD.n1184 0.0200652
R3225 VDD.n1715 VDD.n1714 0.0200652
R3226 VDD.n193 VDD.n192 0.0200283
R3227 VDD.n839 VDD.n686 0.0198458
R3228 VDD.n1708 VDD.n337 0.0197857
R3229 VDD.n1269 VDD.n1268 0.0197857
R3230 VDD.n254 VDD.n253 0.019371
R3231 VDD.n1002 VDD.n1001 0.0191328
R3232 VDD.n790 VDD.n789 0.0191207
R3233 VDD.n795 VDD.n794 0.019083
R3234 VDD.n981 VDD.n931 0.0190047
R3235 VDD.n1274 VDD.n598 0.0187022
R3236 VDD.n1073 VDD.n1033 0.0186452
R3237 VDD.n1068 VDD.n1038 0.0186452
R3238 VDD.n155 VDD.n154 0.0186395
R3239 VDD.n201 VDD.n183 0.0180472
R3240 VDD.n1690 VDD.n1689 0.017691
R3241 VDD.n1251 VDD.n1250 0.0176429
R3242 VDD.n219 VDD.n207 0.0174811
R3243 VDD.n1969 VDD.n1968 0.0173293
R3244 VDD.n837 VDD.n687 0.0173224
R3245 VDD.n829 VDD.n828 0.0173224
R3246 VDD.n1868 VDD.n1867 0.0167254
R3247 VDD.n1540 VDD.n1539 0.0165976
R3248 VDD.n1068 VDD.n1067 0.0164677
R3249 VDD.n930 VDD.n846 0.0160453
R3250 VDD.n859 VDD.n858 0.0159438
R3251 VDD.n858 VDD.n855 0.0159438
R3252 VDD.n929 VDD.n847 0.0159438
R3253 VDD.n1986 VDD 0.0158659
R3254 VDD.n1088 VDD.n678 0.0157992
R3255 VDD.n752 VDD.n725 0.0156402
R3256 VDD.n979 VDD.n978 0.0156402
R3257 VDD.n1082 VDD.n1081 0.015009
R3258 VDD.n788 VDD.n770 0.0149
R3259 VDD VDD.n178 0.0147661
R3260 VDD.n787 VDD.n771 0.014
R3261 VDD.n1870 VDD.n1869 0.0136831
R3262 VDD.n1530 VDD.n1529 0.0136707
R3263 VDD.n1532 VDD.n1531 0.0136707
R3264 VDD.n543 VDD.n542 0.0136707
R3265 VDD.n1464 VDD.n1463 0.0136707
R3266 VDD.n1073 VDD.n1017 0.0135645
R3267 VDD.n58 VDD.n57 0.0134677
R3268 VDD.n862 VDD.n861 0.0130481
R3269 VDD.n857 VDD.n854 0.0130481
R3270 VDD.n857 VDD.n856 0.0130481
R3271 VDD.n1864 VDD.n1863 0.0122692
R3272 VDD.n681 VDD.n679 0.0122391
R3273 VDD.n696 VDD.n695 0.0121599
R3274 VDD.n1080 VDD.n1016 0.0121129
R3275 VDD.n1081 VDD.n1015 0.0119706
R3276 VDD.n782 VDD.n777 0.0118445
R3277 VDD.n419 VDD.n417 0.01175
R3278 VDD.n1828 VDD.n1827 0.0116236
R3279 VDD.n752 VDD.n723 0.0114346
R3280 VDD.n1644 VDD.n404 0.0112143
R3281 VDD.n1369 VDD.n1368 0.0107273
R3282 VDD.n1160 VDD.n637 0.0106124
R3283 VDD.n978 VDD.n977 0.0105935
R3284 VDD.n59 VDD.n12 0.0105
R3285 VDD.n169 VDD.n168 0.0104739
R3286 VDD.n52 VDD.n51 0.0103544
R3287 VDD.n1331 VDD.n1306 0.0101429
R3288 VDD.n860 VDD.n853 0.0100858
R3289 VDD.n923 VDD.n852 0.00993548
R3290 VDD.n838 VDD.n837 0.00975234
R3291 VDD.n1487 VDD 0.00932353
R3292 VDD.n997 VDD.n845 0.00928906
R3293 VDD.n970 VDD.n935 0.00928049
R3294 VDD.n976 VDD.n932 0.00928049
R3295 VDD.n829 VDD.n687 0.00891121
R3296 VDD.n699 VDD.n698 0.00888057
R3297 VDD.n974 VDD.n935 0.00854878
R3298 VDD.n976 VDD.n975 0.00854878
R3299 VDD.n924 VDD.n851 0.00853674
R3300 VDD.n824 VDD.n823 0.00851619
R3301 VDD.n1904 VDD.n1903 0.00848635
R3302 VDD.n787 VDD.n782 0.00806303
R3303 VDD.n743 VDD.n722 0.00778745
R3304 VDD.n541 VDD.n540 0.00775806
R3305 VDD.n1466 VDD.n1465 0.00775806
R3306 VDD.n1085 VDD.n682 0.00754348
R3307 VDD.n756 VDD.n732 0.00742308
R3308 VDD.n811 VDD.n810 0.00742308
R3309 VDD.n695 VDD.n688 0.00742308
R3310 VDD.n1016 VDD.n680 0.00738437
R3311 VDD.n53 VDD.n49 0.00725
R3312 VDD.n53 VDD.n52 0.00725
R3313 VDD.n887 VDD.n886 0.00708537
R3314 VDD.n711 VDD.n709 0.0070587
R3315 VDD.n753 VDD.n726 0.0070587
R3316 VDD.n1113 VDD.n1112 0.00700602
R3317 VDD.n1803 VDD.n1802 0.00700602
R3318 VDD.n836 VDD.n835 0.00669433
R3319 VDD.n90 VDD.n60 0.00667414
R3320 VDD.n1909 VDD 0.00664335
R3321 VDD.n1027 VDD.n1023 0.00661998
R3322 VDD.n697 VDD.n686 0.00638785
R3323 VDD.n813 VDD.n812 0.00632996
R3324 VDD.n805 VDD.n804 0.00632996
R3325 VDD.n803 VDD.n766 0.00632996
R3326 VDD.n712 VDD.n699 0.00632996
R3327 VDD VDD.n1522 0.00630645
R3328 VDD.n531 VDD 0.00630645
R3329 VDD VDD.n500 0.00630645
R3330 VDD VDD.n961 0.00630645
R3331 VDD.n1060 VDD 0.00630645
R3332 VDD VDD.n471 0.00630645
R3333 VDD.n864 VDD.n853 0.00582544
R3334 VDD.n1072 VDD.n1034 0.00579412
R3335 VDD.n697 VDD.n684 0.00572908
R3336 VDD.n1938 VDD.n1937 0.00562658
R3337 VDD.n975 VDD.n974 0.00562195
R3338 VDD.n1082 VDD.n682 0.00558696
R3339 VDD.n203 VDD.n202 0.00531132
R3340 VDD.n977 VDD.n933 0.00489628
R3341 VDD.n753 VDD.n751 0.00487247
R3342 VDD.n1086 VDD.n1085 0.00480435
R3343 VDD.n751 VDD.n750 0.0045081
R3344 VDD.n824 VDD.n726 0.0045081
R3345 VDD.n799 VDD.n767 0.00441304
R3346 VDD.n796 VDD.n795 0.00414372
R3347 VDD.n830 VDD.n689 0.00414372
R3348 VDD.n926 VDD.n850 0.00412903
R3349 VDD.n1079 VDD.n1017 0.00412903
R3350 VDD.n1036 VDD.n1014 0.00402941
R3351 VDD.n1071 VDD.n1035 0.00402941
R3352 VDD.n40 VDD.n39 0.003875
R3353 VDD.n174 VDD.n97 0.00380882
R3354 VDD.n805 VDD.n759 0.00377935
R3355 VDD.n794 VDD.n766 0.00377935
R3356 VDD.n713 VDD.n711 0.00377935
R3357 VDD.n866 VDD.n850 0.00376613
R3358 VDD.n1649 VDD.n1648 0.00371429
R3359 VDD.n1327 VDD.n1326 0.00371429
R3360 VDD.n679 VDD.n678 0.00360796
R3361 VDD.n865 VDD.n851 0.00350186
R3362 VDD.n750 VDD.n742 0.00341498
R3363 VDD VDD.n908 0.00340323
R3364 VDD.n1038 VDD.n1033 0.00340323
R3365 VDD.n713 VDD.n712 0.00305061
R3366 VDD.n698 VDD.n696 0.00305061
R3367 VDD.n926 VDD.n925 0.00304032
R3368 VDD.n47 VDD.n41 0.00283766
R3369 VDD.n825 VDD.n725 0.00283401
R3370 VDD.n48 VDD.n40 0.00275
R3371 VDD.n1098 VDD.n1097 0.00266867
R3372 VDD.n1768 VDD.n1764 0.00266867
R3373 VDD.n788 VDD 0.00254545
R3374 VDD.n1022 VDD.n1016 0.00254545
R3375 VDD.n823 VDD.n822 0.00245652
R3376 VDD.n802 VDD.n764 0.00206522
R3377 VDD.n1736 VDD.n307 0.00192857
R3378 VDD.n30 VDD 0.00186364
R3379 VDD.n82 VDD 0.00163924
R3380 VDD VDD.n143 0.00163924
R3381 VDD VDD.n242 0.00163924
R3382 VDD VDD.n1900 0.00163924
R3383 VDD.n835 VDD.n689 0.00159312
R3384 VDD.n830 VDD.n722 0.00159312
R3385 VDD.n1361 VDD.n1359 0.00152273
R3386 VDD.n1564 VDD.n1563 0.00152273
R3387 VDD.n1089 VDD 0.00151695
R3388 VDD.n203 VDD 0.00134906
R3389 VDD.n1867 VDD.n269 0.00132534
R3390 VDD.n2006 VDD 0.00128947
R3391 VDD.n804 VDD.n803 0.00122874
R3392 VDD VDD.n260 0.00122581
R3393 VDD.n256 VDD 0.00122581
R3394 VDD.n1067 VDD.n1039 0.00122581
R3395 VDD.n1152 VDD.n1151 0.00121429
R3396 VDD VDD.n161 0.00119767
R3397 VDD.n157 VDD 0.00119767
R3398 VDD.n865 VDD.n864 0.00103254
R3399 VDD.n1023 VDD.n1022 0.00101136
R3400 VDD.n923 VDD.n866 0.000862903
R3401 VDD.n1001 VDD 0.000851563
R3402 VDD.n1896 VDD 0.000807167
R3403 VDD.n1906 VDD 0.000807167
R3404 VDD.n72 VDD 0.000737467
R3405 VDD VDD.n1926 0.000693548
R3406 VDD.n59 VDD.n58 0.000693548
R3407 VDD.n97 VDD.n93 0.000665441
R3408 RES_74k_1.M.t1 RES_74k_1.M.t7 3.92959
R3409 RES_74k_1.M.t1 RES_74k_1.M.n0 3.19141
R3410 RES_74k_1.M.t1 RES_74k_1.M 6.92211
R3411 RES_74k_1.M RES_74k_1.M.t0 6.14618
R3412 RES_74k_1.M.t1 RES_74k_1.M.t6 5.18834
R3413 RES_74k_1.M.t1 RES_74k_1.M.t4 5.18264
R3414 RES_74k_1.M.t1 RES_74k_1.M.t2 3.07204
R3415 RES_74k_1.M.t1 RES_74k_1.M.t3 3.0618
R3416 RES_74k_1.M.t1 RES_74k_1.M.t5 3.0279
R3417 VSS.n4304 VSS.n4303 5.941e+06
R3418 VSS.n5667 VSS.n5664 5.941e+06
R3419 VSS.n5667 VSS.n5666 3.75375e+06
R3420 VSS.n5718 VSS.n5717 3.75375e+06
R3421 VSS.n5724 VSS.n5723 548485
R3422 VSS.t621 VSS.t647 44337.9
R3423 VSS.n5723 VSS.n5722 42998.3
R3424 VSS.n5722 VSS.n5720 37872
R3425 VSS.n5725 VSS.n5724 28016
R3426 VSS.n5720 VSS.n5719 26587
R3427 VSS.n4305 VSS.n4304 15212.8
R3428 VSS.n5889 VSS.n5887 10655.7
R3429 VSS.n4997 VSS.n4996 10552.3
R3430 VSS.n5868 VSS.n5867 9445.69
R3431 VSS.n5768 VSS.t466 8953.91
R3432 VSS.n5820 VSS.n5758 8778.74
R3433 VSS.n5768 VSS.t454 7394.69
R3434 VSS.n5722 VSS.n5721 7304.73
R3435 VSS.t501 VSS.n5811 7210.65
R3436 VSS.n5719 VSS.t683 6204.1
R3437 VSS.n4996 VSS.n4995 6119.25
R3438 VSS.t578 VSS.n5750 4486.13
R3439 VSS.t532 VSS.t652 3685.04
R3440 VSS.n5810 VSS.t246 3621.08
R3441 VSS.n4303 VSS.n4302 3301.18
R3442 VSS.n5338 VSS.n5337 2891.56
R3443 VSS.n5891 VSS.n5890 2413.12
R3444 VSS.t763 VSS.t694 2166.67
R3445 VSS.t452 VSS.t549 2166.67
R3446 VSS.t247 VSS.t498 2166.67
R3447 VSS.n4735 VSS.n4734 1890.45
R3448 VSS.t709 VSS.t711 1842.52
R3449 VSS.t711 VSS.t531 1842.52
R3450 VSS.t724 VSS.t714 1822.88
R3451 VSS.t179 VSS.t445 1805.06
R3452 VSS.t195 VSS.t482 1778.39
R3453 VSS.n5821 VSS.n5820 1752.01
R3454 VSS.n959 VSS.t724 1720.94
R3455 VSS.t611 VSS.t618 1717.16
R3456 VSS.t613 VSS.t615 1707.46
R3457 VSS.t683 VSS.t596 1707.46
R3458 VSS.t204 VSS.t446 1657.99
R3459 VSS.t187 VSS.t439 1649.75
R3460 VSS.n4248 VSS.t677 1557.29
R3461 VSS.n6034 VSS.n6033 1536.82
R3462 VSS.n4841 VSS.n4840 1514.17
R3463 VSS.t464 VSS.n5891 1469.82
R3464 VSS.n4571 VSS.t195 1404.92
R3465 VSS.n48 VSS.t179 1316.01
R3466 VSS.n4590 VSS.t187 1303.3
R3467 VSS.n4392 VSS.t216 1229.06
R3468 VSS.n4669 VSS.t213 1229.06
R3469 VSS.n4590 VSS.t139 1224.94
R3470 VSS.t482 VSS.t244 1209.3
R3471 VSS.t445 VSS.t480 1209.3
R3472 VSS.t702 VSS.n5868 1153.55
R3473 VSS.n5811 VSS.t453 1153.55
R3474 VSS.t439 VSS.t483 1121.83
R3475 VSS.t446 VSS.t481 1121.83
R3476 VSS.t618 VSS.t613 1086.57
R3477 VSS.t598 VSS.t611 1086.57
R3478 VSS.t600 VSS.t598 1086.57
R3479 VSS.t596 VSS.t600 1086.57
R3480 VSS.t637 VSS.t639 1083.33
R3481 VSS.t639 VSS.t702 1083.33
R3482 VSS.t632 VSS.t634 1083.33
R3483 VSS.t634 VSS.t453 1083.33
R3484 VSS.t420 VSS.t418 1083.33
R3485 VSS.t246 VSS.t420 1083.33
R3486 VSS.n5825 VSS.t436 1074.31
R3487 VSS.n5757 VSS.t623 1061.73
R3488 VSS.t442 VSS.t496 1060.11
R3489 VSS.t466 VSS.t509 1047.76
R3490 VSS.n5890 VSS.n5718 1046.74
R3491 VSS.n5751 VSS.t581 967.024
R3492 VSS.n860 VSS.n859 953.981
R3493 VSS.n424 VSS.n423 944.048
R3494 VSS.n1479 VSS.n1478 929.726
R3495 VSS.n5867 VSS.t532 921.26
R3496 VSS.n5867 VSS.t709 921.26
R3497 VSS.n5889 VSS.n5888 914.569
R3498 VSS.t154 VSS.t342 855.827
R3499 VSS.n5750 VSS.t493 797.606
R3500 VSS.t454 VSS.t686 781.737
R3501 VSS.n5869 VSS.t637 767.361
R3502 VSS.n5798 VSS.t632 767.361
R3503 VSS.t418 VSS.n5809 767.361
R3504 VSS.t758 VSS.n5725 756.434
R3505 VSS.n5887 VSS.t484 750.444
R3506 VSS.t469 VSS.t450 727.73
R3507 VSS.n5719 VSS.t423 720.212
R3508 VSS.n5840 VSS.t258 658.784
R3509 VSS.t447 VSS.n5886 650.385
R3510 VSS.n114 VSS.t184 617.99
R3511 VSS.t281 VSS.t279 581.962
R3512 VSS.t300 VSS.t281 581.962
R3513 VSS.t309 VSS.t300 581.962
R3514 VSS.t323 VSS.t325 581.962
R3515 VSS.t325 VSS.t335 581.962
R3516 VSS.n4954 VSS.n4953 572.302
R3517 VSS.n939 VSS.t715 561.086
R3518 VSS.n5867 VSS 552.953
R3519 VSS.t678 VSS.t221 522.588
R3520 VSS.t680 VSS.t441 522.588
R3521 VSS.n5819 VSS.t507 515.361
R3522 VSS.n5822 VSS.t578 481.087
R3523 VSS.n5319 VSS.n5318 477.231
R3524 VSS.n4468 VSS.t309 421.495
R3525 VSS.t250 VSS.t661 419.226
R3526 VSS.n591 VSS.n590 407.524
R3527 VSS.t450 VSS.t760 399.077
R3528 VSS.t642 VSS.t626 399.077
R3529 VSS.t644 VSS.t628 399.077
R3530 VSS.t473 VSS.t501 399.077
R3531 VSS.t561 VSS.t580 390.616
R3532 VSS.t583 VSS.t263 390.616
R3533 VSS.t733 VSS.t476 390.616
R3534 VSS.t729 VSS.t470 390.616
R3535 VSS.t575 VSS.t260 390.344
R3536 VSS.t572 VSS.t490 390.154
R3537 VSS.t728 VSS.t489 388.692
R3538 VSS.n5852 VSS.t225 365.812
R3539 VSS.n5823 VSS.n5822 352.084
R3540 VSS.n5869 VSS.t763 315.973
R3541 VSS.n5798 VSS.t452 315.973
R3542 VSS.n5809 VSS.t247 315.973
R3543 VSS.n162 VSS.t370 297.88
R3544 VSS.n199 VSS.t286 288.988
R3545 VSS.n5749 VSS.t487 282.526
R3546 VSS.n4998 VSS.n4997 281.462
R3547 VSS.n5758 VSS.n5757 279.142
R3548 VSS.n4611 VSS.t145 266.759
R3549 VSS.n202 VSS.t288 253.421
R3550 VSS.n5868 VSS.t443 248.296
R3551 VSS.n165 VSS.t358 244.529
R3552 VSS.n5820 VSS.n5819 240.343
R3553 VSS.t457 VSS.t256 232.776
R3554 VSS.t461 VSS.n5866 231.668
R3555 VSS.n5719 VSS.t242 223.135
R3556 VSS.t760 VSS.n5768 200.844
R3557 VSS.n4635 VSS.t479 191.177
R3558 VSS.n149 VSS.t160 186.731
R3559 VSS.t663 VSS.t505 182.947
R3560 VSS.n4617 VSS.t478 182.286
R3561 VSS.n5817 VSS.t654 181.751
R3562 VSS.t650 VSS.n5841 179.668
R3563 VSS.n121 VSS.t379 164.501
R3564 VSS.n5769 VSS.t469 164.327
R3565 VSS.t642 VSS.t500 164.327
R3566 VSS.t626 VSS.t644 164.327
R3567 VSS.t628 VSS.t473 164.327
R3568 VSS.n4468 VSS.t323 160.468
R3569 VSS.n5822 VSS.n5821 160.02
R3570 VSS.n5818 VSS.t474 156.163
R3571 VSS.n410 VSS.t675 154.649
R3572 VSS.n1526 VSS.n1525 145.089
R3573 VSS.n5851 VSS.t463 141.845
R3574 VSS.n465 VSS.t736 137.732
R3575 VSS.t746 VSS.t750 134.906
R3576 VSS.n456 VSS.n455 132.9
R3577 VSS.n5717 VSS.n5716 130.788
R3578 VSS.n206 VSS.t332 128.934
R3579 VSS.n1201 VSS.n1200 127.87
R3580 VSS.n4697 VSS.t271 127.856
R3581 VSS.n4984 VSS.n4983 127.537
R3582 VSS.n5890 VSS.n5889 126.573
R3583 VSS.n189 VSS.t355 120.041
R3584 VSS.n568 VSS.n567 116.502
R3585 VSS.n4210 VSS.t674 115.596
R3586 VSS.n391 VSS.n390 109.445
R3587 VSS.t569 VSS.n5749 107.629
R3588 VSS.n5821 VSS.t429 92.842
R3589 VSS.t772 VSS.t521 88.6679
R3590 VSS.n5668 VSS.n5667 82.9732
R3591 VSS.n4940 VSS.t606 81.8473
R3592 VSS.n5693 VSS.n5692 81.5669
R3593 VSS.n5811 VSS.n5810 80.7206
R3594 VSS.t474 VSS.t502 75.3316
R3595 VSS.t505 VSS.n5771 74.1359
R3596 VSS.n569 VSS.n568 71.3171
R3597 VSS.n4724 VSS.t264 70.1147
R3598 VSS.n804 VSS.t558 68.7194
R3599 VSS.n854 VSS.t551 68.7194
R3600 VSS.n1432 VSS.t511 68.7194
R3601 VSS.n1489 VSS.t514 68.7194
R3602 VSS.n4629 VSS.t245 66.69
R3603 VSS.n325 VSS.t670 64.2392
R3604 VSS.n4711 VSS.t266 61.866
R3605 VSS.n474 VSS.t741 60.4094
R3606 VSS.n4847 VSS.t764 57.9753
R3607 VSS.n4922 VSS.t699 57.9753
R3608 VSS.n4881 VSS.t593 57.9753
R3609 VSS.n4623 VSS.t440 57.798
R3610 VSS.n4644 VSS.t148 57.798
R3611 VSS.n6017 VSS.n6016 57.7657
R3612 VSS.n6027 VSS.n6026 55.1928
R3613 VSS.n5503 VSS.t136 51.6521
R3614 VSS.n4818 VSS.t526 51.1548
R3615 VSS.n4931 VSS.t696 51.1548
R3616 VSS.n4890 VSS.t608 51.1548
R3617 VSS.n5417 VSS.t233 49.6265
R3618 VSS.n4249 VSS.n4248 49.1159
R3619 VSS.n4897 VSS.n4896 44.3342
R3620 VSS.t776 VSS.t775 44.058
R3621 VSS.n5339 VSS.n5338 43.5499
R3622 VSS.n1226 VSS.n1225 42.6234
R3623 VSS.n5035 VSS.t660 41.5243
R3624 VSS.n5133 VSS.t133 41.5243
R3625 VSS.n5857 VSS.t224 38.8649
R3626 VSS.n4818 VSS.t769 37.5136
R3627 VSS.n5666 VSS.n5665 36.2122
R3628 VSS.n5479 VSS.t659 35.4477
R3629 VSS.n4103 VSS.n4102 32.9568
R3630 VSS.n4494 VSS.n4493 31.0858
R3631 VSS.n4847 VSS.t523 30.6931
R3632 VSS.n1295 VSS.n1294 29.9489
R3633 VSS.n5971 VSS.n5970 29.3566
R3634 VSS.n3932 VSS.n3931 29.0184
R3635 VSS.n1285 VSS.t671 28.751
R3636 VSS.n1389 VSS.n1388 28.7316
R3637 VSS.t224 VSS.t776 28.6791
R3638 VSS.n5575 VSS.t274 28.3582
R3639 VSS.n4898 VSS.t427 27.2828
R3640 VSS.n5182 VSS.t320 26.3327
R3641 VSS.n4113 VSS.n4112 26.1965
R3642 VSS.n414 VSS.t665 26.1718
R3643 VSS.n495 VSS.n494 26.0884
R3644 VSS.n5952 VSS.n5951 25.5687
R3645 VSS.n4102 VSS.t746 25.3911
R3646 VSS.n953 VSS.t756 25.3179
R3647 VSS.n480 VSS.t739 24.1641
R3648 VSS.n4898 VSS.n4897 23.8725
R3649 VSS.n4077 VSS.t248 21.9714
R3650 VSS.n5812 VSS.n5770 21.6
R3651 VSS.n4306 VSS.n4305 20.5962
R3652 VSS.n913 VSS.t449 19.4363
R3653 VSS.n425 VSS.n424 19.0342
R3654 VSS.n5396 VSS.t297 18.2305
R3655 VSS.t507 VSS.n5818 17.9365
R3656 VSS.n5575 VSS.n5574 17.2177
R3657 VSS.n4824 VSS.t772 17.0519
R3658 VSS.n4086 VSS.n4085 15.2111
R3659 VSS.n4109 VSS.t740 15.2111
R3660 VSS.n5440 VSS.t292 15.1921
R3661 VSS.t496 VSS.t621 14.9316
R3662 VSS.t463 VSS.t442 14.9316
R3663 VSS.n5852 VSS.n5851 14.9316
R3664 VSS.t225 VSS.t678 14.9316
R3665 VSS.t221 VSS.t680 14.9316
R3666 VSS.t441 VSS.t460 14.9316
R3667 VSS.n5008 VSS.t176 13.1666
R3668 VSS.n5029 VSS.t658 13.1666
R3669 VSS.n5434 VSS.t306 13.1666
R3670 VSS.n5829 VSS.n5746 12.9101
R3671 VSS.t258 VSS.t758 11.9784
R3672 VSS.n5841 VSS.n5840 11.9784
R3673 VSS.t661 VSS.t650 11.9784
R3674 VSS.t647 VSS.t250 11.9784
R3675 VSS.n1010 VSS.t612 11.3982
R3676 VSS.n3991 VSS.t545 11.0483
R3677 VSS.n5810 VSS.t663 10.9931
R3678 VSS.n1015 VSS.n1014 10.7852
R3679 VSS.n4051 VSS.t539 10.3984
R3680 VSS.n4188 VSS.t718 10.315
R3681 VSS.n5540 VSS.t312 10.1283
R3682 VSS.n4017 VSS.t543 9.74855
R3683 VSS.n5886 VSS.t564 9.62158
R3684 VSS.n508 VSS.n507 9.61182
R3685 VSS.n5060 VSS.t173 9.55913
R3686 VSS.n4510 VSS.t194 9.55885
R3687 VSS.n76 VSS.t230 9.54136
R3688 VSS.n5047 VSS.t208 9.54089
R3689 VSS.n5048 VSS.t135 9.51568
R3690 VSS.n87 VSS.t186 9.5154
R3691 VSS.n5046 VSS.t239 9.5085
R3692 VSS.n63 VSS.t144 9.50824
R3693 VSS.n4509 VSS.t206 9.49457
R3694 VSS.n33 VSS.t178 9.49428
R3695 VSS.n32 VSS.t197 9.49428
R3696 VSS.n31 VSS.t212 9.49428
R3697 VSS.n58 VSS.t203 9.49428
R3698 VSS.n4948 VSS.t227 9.49403
R3699 VSS.n4947 VSS.t235 9.49403
R3700 VSS.n4908 VSS.t191 9.49403
R3701 VSS.n4790 VSS.t175 9.49403
R3702 VSS.n5049 VSS.t181 9.49372
R3703 VSS.n59 VSS.t147 9.45083
R3704 VSS.n4789 VSS.t237 9.45057
R3705 VSS.n85 VSS.t201 9.43205
R3706 VSS.n4507 VSS.t138 9.43205
R3707 VSS.n93 VSS.t164 9.43205
R3708 VSS.n74 VSS.t218 9.43205
R3709 VSS.n65 VSS.t159 9.43205
R3710 VSS.n5058 VSS.t162 9.43205
R3711 VSS.n5093 VSS.t210 9.43205
R3712 VSS.n5114 VSS.t189 9.43205
R3713 VSS.n5086 VSS.t199 9.43205
R3714 VSS.n5105 VSS.t132 9.43205
R3715 VSS.n4378 VSS.t156 9.3886
R3716 VSS.n5281 VSS.t171 9.3886
R3717 VSS.n5305 VSS.t232 9.3886
R3718 VSS.n4409 VSS.t153 9.3886
R3719 VSS.n243 VSS.t183 9.34514
R3720 VSS.n4382 VSS.t215 9.34514
R3721 VSS.n108 VSS.t150 9.34514
R3722 VSS.n5236 VSS.t169 9.34514
R3723 VSS.n5257 VSS.t141 9.34514
R3724 VSS.n5241 VSS.t166 9.34514
R3725 VSS.n1460 VSS.n1458 9.13939
R3726 VSS.n4716 VSS.n4714 9.13939
R3727 VSS.n4718 VSS.n4716 9.13939
R3728 VSS.n4712 VSS.n4710 9.13939
R3729 VSS.n4710 VSS.n4709 9.13939
R3730 VSS.n839 VSS.n837 9.13939
R3731 VSS.n4930 VSS.n4913 9.13939
R3732 VSS.n4932 VSS.n4930 9.13939
R3733 VSS.n4817 VSS.n4801 9.13939
R3734 VSS.n4819 VSS.n4817 9.13939
R3735 VSS.n4855 VSS.n4838 9.13939
R3736 VSS.n4857 VSS.n4855 9.13939
R3737 VSS.n4889 VSS.n4795 9.13939
R3738 VSS.n4891 VSS.n4889 9.13939
R3739 VSS.n5008 VSS.n5007 9.11549
R3740 VSS.n6058 VSS.t685 8.89703
R3741 VSS.n26 VSS.n25 8.78137
R3742 VSS.n27 VSS.t597 8.5505
R3743 VSS.n28 VSS.t605 8.5505
R3744 VSS.n6058 VSS.t684 8.5505
R3745 VSS.n1010 VSS.n1009 8.5505
R3746 VSS.t213 VSS.t204 8.24923
R3747 VSS.n4157 VSS.n4155 8.16717
R3748 VSS.n1078 VSS.n1077 7.61323
R3749 VSS.n1468 VSS.n1466 7.58383
R3750 VSS.n5829 VSS.n5828 7.54047
R3751 VSS.n957 VSS.n956 7.50194
R3752 VSS.n830 VSS.n828 7.48661
R3753 VSS.n5857 VSS.t220 7.3005
R3754 VSS.n5485 VSS.t657 7.08994
R3755 VSS.n5832 VSS.n5731 6.8902
R3756 VSS.n5833 VSS.n5730 6.87063
R3757 VSS.n1382 VSS.n1381 6.76077
R3758 VSS.n5746 VSS.t582 6.68867
R3759 VSS.n5828 VSS.t579 6.68867
R3760 VSS.n924 VSS.n923 6.65541
R3761 VSS.n948 VSS.t725 6.65541
R3762 VSS.n1425 VSS.n1418 6.65541
R3763 VSS.n1425 VSS.n1419 6.65541
R3764 VSS.n1482 VSS.t515 6.65541
R3765 VSS.n1482 VSS.t542 6.65541
R3766 VSS.n1405 VSS.t546 6.65541
R3767 VSS.n3981 VSS.n1524 6.65541
R3768 VSS.n797 VSS.n790 6.65541
R3769 VSS.n797 VSS.n791 6.65541
R3770 VSS.n863 VSS.t703 6.65541
R3771 VSS.n863 VSS.t552 6.65541
R3772 VSS.n4868 VSS.t773 6.65541
R3773 VSS.n4843 VSS.n4839 6.65541
R3774 VSS.n4805 VSS.n4802 6.65541
R3775 VSS.n4830 VSS.t522 6.65541
R3776 VSS.n4877 VSS.n4796 6.65541
R3777 VSS.n4904 VSS.t607 6.65541
R3778 VSS.n4943 VSS.t428 6.65541
R3779 VSS.n4918 VSS.n4914 6.65541
R3780 VSS.n4198 VSS.t757 6.65541
R3781 VSS.n4138 VSS.n890 6.65541
R3782 VSS.n4691 VSS.n29 6.65541
R3783 VSS.n4691 VSS.n30 6.65541
R3784 VSS.n4732 VSS.t265 6.65541
R3785 VSS.n4732 VSS.t693 6.65541
R3786 VSS.t443 VSS.t461 6.65125
R3787 VSS.t256 VSS.t464 6.65125
R3788 VSS.n4508 VSS.t140 6.63905
R3789 VSS.n5059 VSS.t163 6.63905
R3790 VSS.n4379 VSS.t158 6.63522
R3791 VSS.n5306 VSS.t234 6.63522
R3792 VSS.n5282 VSS.t172 6.63522
R3793 VSS.n4410 VSS.t155 6.63522
R3794 VSS.n4383 VSS.t217 6.63331
R3795 VSS.n5258 VSS.t143 6.63331
R3796 VSS.n5735 VSS.t574 6.62607
R3797 VSS.n5743 VSS.t590 6.62607
R3798 VSS.n5736 VSS.n5732 6.6202
R3799 VSS.n5744 VSS.n5740 6.6202
R3800 VSS.n244 VSS.t185 6.5165
R3801 VSS.n5237 VSS.t170 6.5165
R3802 VSS.n109 VSS.t152 6.50525
R3803 VSS.n5242 VSS.t168 6.50525
R3804 VSS.n148 VSS.t371 6.4265
R3805 VSS.n146 VSS.t404 6.4265
R3806 VSS.n141 VSS.t367 6.4265
R3807 VSS.n77 VSS.t202 6.4265
R3808 VSS.n88 VSS.t165 6.4265
R3809 VSS.n64 VSS.t219 6.4265
R3810 VSS.n66 VSS.t161 6.4265
R3811 VSS.n4357 VSS.n4356 6.4265
R3812 VSS.n105 VSS.n104 6.4265
R3813 VSS.n103 VSS.n102 6.4265
R3814 VSS.n5104 VSS.t190 6.4265
R3815 VSS.n5151 VSS.n5146 6.4265
R3816 VSS.n5081 VSS.n5080 6.4265
R3817 VSS.n5302 VSS.t291 6.4265
R3818 VSS.n5233 VSS.t374 6.4265
R3819 VSS.n5238 VSS.t350 6.4265
R3820 VSS.n5079 VSS.t200 6.4265
R3821 VSS.n5088 VSS.t211 6.4265
R3822 VSS.n5153 VSS.n5145 6.4265
R3823 VSS.n5106 VSS.t134 6.4265
R3824 VSS.n5738 VSS.n5737 6.4265
R3825 VSS.n5745 VSS.n5739 6.4265
R3826 VSS.n3738 VSS.n3737 6.39416
R3827 VSS.n5862 VSS.n5846 6.23171
R3828 VSS.n5877 VSS.n5876 6.23168
R3829 VSS.n5794 VSS.n5772 6.23168
R3830 VSS.n5873 VSS.n5872 6.02724
R3831 VSS.n5875 VSS.n5874 6.02724
R3832 VSS.n5802 VSS.n5801 6.02724
R3833 VSS.n4123 VSS.n4122 5.91574
R3834 VSS.n1176 VSS.n1175 5.84933
R3835 VSS.n259 VSS.n258 5.80511
R3836 VSS.n528 VSS.n527 5.60395
R3837 VSS.n5892 VSS.t253 5.54279
R3838 VSS.n1028 VSS.n1027 5.4005
R3839 VSS.n1028 VSS.t614 5.4005
R3840 VSS.n24 VSS.n23 5.4005
R3841 VSS.n24 VSS.t599 5.4005
R3842 VSS VSS.t508 5.34447
R3843 VSS VSS.t257 5.34447
R3844 VSS VSS.t465 5.34447
R3845 VSS VSS.t475 5.34447
R3846 VSS VSS.n5857 5.27587
R3847 VSS.n270 VSS.n269 5.26318
R3848 VSS.n6060 VSS.n6059 5.24323
R3849 VSS.n5862 VSS.t695 5.23126
R3850 VSS.n5876 VSS.t653 5.23126
R3851 VSS.n5850 VSS.t497 5.23126
R3852 VSS.n5849 VSS.t622 5.23126
R3853 VSS.n5797 VSS.t550 5.23126
R3854 VSS.n5772 VSS.t499 5.23126
R3855 VSS.n5803 VSS.t451 5.23126
R3856 VSS.n5796 VSS.t761 5.23126
R3857 VSS.n1012 VSS.n1011 5.20095
R3858 VSS.n952 VSS.n951 5.2005
R3859 VSS.n954 VSS.n953 5.2005
R3860 VSS.n3998 VSS.n3997 5.2005
R3861 VSS.n4022 VSS.n4021 5.2005
R3862 VSS.n4016 VSS.n4015 5.2005
R3863 VSS.n4015 VSS.n4014 5.2005
R3864 VSS.n1516 VSS.n1515 5.2005
R3865 VSS.n286 VSS.n285 5.2005
R3866 VSS.n285 VSS.n284 5.2005
R3867 VSS.n289 VSS.n288 5.2005
R3868 VSS.n288 VSS.n287 5.2005
R3869 VSS.n293 VSS.n291 5.2005
R3870 VSS.n293 VSS.n292 5.2005
R3871 VSS.n278 VSS.n277 5.2005
R3872 VSS.n466 VSS.n465 5.2005
R3873 VSS.n830 VSS.n820 5.2005
R3874 VSS.n830 VSS.n829 5.2005
R3875 VSS.n359 VSS.n338 5.2005
R3876 VSS.n330 VSS.n329 5.2005
R3877 VSS.n329 VSS.n328 5.2005
R3878 VSS.n333 VSS.n332 5.2005
R3879 VSS.n332 VSS.n331 5.2005
R3880 VSS.n341 VSS.n340 5.2005
R3881 VSS.n4134 VSS.n4133 5.2005
R3882 VSS.n4192 VSS.n4191 5.2005
R3883 VSS.n4157 VSS.n4156 5.2005
R3884 VSS.n4178 VSS.n4177 5.2005
R3885 VSS.n4218 VSS.n4217 5.2005
R3886 VSS.n4217 VSS.n4216 5.2005
R3887 VSS.n4215 VSS.n4214 5.2005
R3888 VSS.n4214 VSS.n4213 5.2005
R3889 VSS.n4687 VSS.n4686 5.2005
R3890 VSS VSS.n5869 5.2005
R3891 VSS VSS.n5892 5.2005
R3892 VSS.n5866 VSS 5.2005
R3893 VSS VSS.n5852 5.2005
R3894 VSS VSS.n5851 5.2005
R3895 VSS.n5881 VSS.n5840 5.2005
R3896 VSS.n5880 VSS.n5841 5.2005
R3897 VSS.n5886 VSS 5.2005
R3898 VSS VSS.n5798 5.2005
R3899 VSS.n5809 VSS 5.2005
R3900 VSS.n1466 VSS.n1465 5.2005
R3901 VSS.n1395 VSS.n1394 5.2005
R3902 VSS.n4122 VSS.n4121 5.2005
R3903 VSS.n4120 VSS.n917 5.2005
R3904 VSS.n1397 VSS.n1396 5.2005
R3905 VSS.n914 VSS.n913 5.2005
R3906 VSS.n4129 VSS.n4128 5.2005
R3907 VSS.n4132 VSS.n4131 5.2005
R3908 VSS.n916 VSS.n915 5.2005
R3909 VSS.n960 VSS.n959 5.2005
R3910 VSS.n964 VSS.n963 5.2005
R3911 VSS.n4203 VSS.n4202 5.2005
R3912 VSS.n4205 VSS.n4204 5.2005
R3913 VSS.n4207 VSS.n4206 5.2005
R3914 VSS.n5817 VSS 5.2005
R3915 VSS.n5771 VSS 5.2005
R3916 VSS.n5791 VSS.n5790 5.2005
R3917 VSS.n5785 VSS.n5784 5.2005
R3918 VSS.n1030 VSS.n1026 5.2005
R3919 VSS.n999 VSS.n0 5.2005
R3920 VSS VSS.n1 5.2005
R3921 VSS.n6068 VSS.n2 5.2005
R3922 VSS.n6067 VSS.n18 5.2005
R3923 VSS.n6066 VSS.n19 5.2005
R3924 VSS.n6064 VSS.n22 5.2005
R3925 VSS.n6062 VSS.n6056 5.2005
R3926 VSS.n6061 VSS.n6057 5.2005
R3927 VSS.n1024 VSS.n1023 5.2005
R3928 VSS.n1031 VSS.n1025 5.2005
R3929 VSS.n144 VSS.t336 5.1234
R3930 VSS.n4502 VSS.t403 5.12337
R3931 VSS.n5528 VSS.n5527 5.12337
R3932 VSS.n4406 VSS.n4395 5.12334
R3933 VSS.n5301 VSS.t275 5.12332
R3934 VSS.n5149 VSS.n5147 5.12328
R3935 VSS.n5265 VSS.t316 5.12118
R3936 VSS.n4360 VSS.n4359 5.12105
R3937 VSS.n5787 VSS.t243 5.06622
R3938 VSS.n5882 VSS.t259 5.06496
R3939 VSS.n5883 VSS.t759 5.06496
R3940 VSS.n5786 VSS.t424 5.06496
R3941 VSS.n4088 VSS.n1393 4.88533
R3942 VSS.n327 VSS.n324 4.88449
R3943 VSS.n283 VSS.n280 4.88277
R3944 VSS.n4212 VSS.n4209 4.88215
R3945 VSS.n4177 VSS.t743 4.6889
R3946 VSS.n5895 VSS.n5894 4.63868
R3947 VSS.n2795 VSS.n2794 4.50764
R3948 VSS.n2662 VSS.n2661 4.50764
R3949 VSS.n2791 VSS.n2790 4.50622
R3950 VSS.n2724 VSS.n2723 4.50622
R3951 VSS.n2562 VSS.n2561 4.50565
R3952 VSS.n2658 VSS.n2657 4.50564
R3953 VSS.n2197 VSS.n2195 4.50554
R3954 VSS.n2881 VSS.n2880 4.50542
R3955 VSS.n2582 VSS.n2581 4.50495
R3956 VSS.n2493 VSS.n2492 4.5026
R3957 VSS.n2492 VSS.n2491 4.50224
R3958 VSS.n2882 VSS.n2881 4.50095
R3959 VSS.n2794 VSS.n2793 4.50095
R3960 VSS.n2792 VSS.n2791 4.50095
R3961 VSS.n2726 VSS.n2197 4.50095
R3962 VSS.n2725 VSS.n2724 4.50095
R3963 VSS.n2661 VSS.n2660 4.50095
R3964 VSS.n2563 VSS.n2562 4.50089
R3965 VSS.n2659 VSS.n2658 4.50089
R3966 VSS.n2582 VSS.n2564 4.50089
R3967 VSS.n4011 VSS.n4008 4.5005
R3968 VSS.n4011 VSS.n4010 4.5005
R3969 VSS.n4001 VSS.n4000 4.5005
R3970 VSS.n1519 VSS.n1518 4.5005
R3971 VSS.n296 VSS.n295 4.5005
R3972 VSS.n295 VSS.n294 4.5005
R3973 VSS.n468 VSS.n467 4.5005
R3974 VSS.n283 VSS.n282 4.5005
R3975 VSS.n282 VSS.n281 4.5005
R3976 VSS.n833 VSS.n826 4.5005
R3977 VSS.n833 VSS.n832 4.5005
R3978 VSS.n262 VSS.n261 4.5005
R3979 VSS.n261 VSS.n260 4.5005
R3980 VSS.n327 VSS.n326 4.5005
R3981 VSS.n326 VSS.n325 4.5005
R3982 VSS.n346 VSS.n345 4.5005
R3983 VSS.n345 VSS.n344 4.5005
R3984 VSS.n2001 VSS.n1996 4.5005
R3985 VSS.n2018 VSS.n2004 4.5005
R3986 VSS.n2015 VSS.n2014 4.5005
R3987 VSS.n2019 VSS.n2005 4.5005
R3988 VSS.n2070 VSS.n2069 4.5005
R3989 VSS.n2083 VSS.n2082 4.5005
R3990 VSS.n2842 VSS.n2841 4.5005
R3991 VSS.n2025 VSS.n2023 4.5005
R3992 VSS.n2804 VSS.n2803 4.5005
R3993 VSS.n2817 VSS.n2816 4.5005
R3994 VSS.n2829 VSS.n2828 4.5005
R3995 VSS.n2878 VSS.n2877 4.5005
R3996 VSS.n2815 VSS.n2814 4.5005
R3997 VSS.n2827 VSS.n2826 4.5005
R3998 VSS.n2068 VSS.n2067 4.5005
R3999 VSS.n2031 VSS.n2016 4.5005
R4000 VSS.n2858 VSS.n2857 4.5005
R4001 VSS.n2039 VSS.n2038 4.5005
R4002 VSS.n2876 VSS.n2875 4.5005
R4003 VSS.n2867 VSS.n2866 4.5005
R4004 VSS.n2037 VSS.n2027 4.5005
R4005 VSS.n2840 VSS.n2839 4.5005
R4006 VSS.n2831 VSS.n2830 4.5005
R4007 VSS.n2081 VSS.n2078 4.5005
R4008 VSS.n2046 VSS.n2045 4.5005
R4009 VSS.n2041 VSS.n2040 4.5005
R4010 VSS.n2000 VSS.n1997 4.5005
R4011 VSS.n2088 VSS.n2085 4.5005
R4012 VSS.n2806 VSS.n2805 4.5005
R4013 VSS.n2825 VSS.n2824 4.5005
R4014 VSS.n2012 VSS.n2008 4.5005
R4015 VSS.n2813 VSS.n2812 4.5005
R4016 VSS.n2846 VSS.n2845 4.5005
R4017 VSS.n2036 VSS.n2035 4.5005
R4018 VSS.n2860 VSS.n2859 4.5005
R4019 VSS.n2065 VSS.n2063 4.5005
R4020 VSS.n2071 VSS.n2066 4.5005
R4021 VSS.n2869 VSS.n2868 4.5005
R4022 VSS.n2187 VSS.n2178 4.5005
R4023 VSS.n2732 VSS.n2175 4.5005
R4024 VSS.n2133 VSS.n2132 4.5005
R4025 VSS.n2138 VSS.n2117 4.5005
R4026 VSS.n2106 VSS.n2103 4.5005
R4027 VSS.n2136 VSS.n2135 4.5005
R4028 VSS.n2107 VSS.n2105 4.5005
R4029 VSS.n2139 VSS.n2118 4.5005
R4030 VSS.n2176 VSS.n2174 4.5005
R4031 VSS.n2184 VSS.n2165 4.5005
R4032 VSS.n2186 VSS.n2185 4.5005
R4033 VSS.n2731 VSS.n2730 4.5005
R4034 VSS.n2101 VSS.n2095 4.5005
R4035 VSS.n2788 VSS.n2787 4.5005
R4036 VSS.n2734 VSS.n2733 4.5005
R4037 VSS.n2164 VSS.n2129 4.5005
R4038 VSS.n2099 VSS.n2096 4.5005
R4039 VSS.n2776 VSS.n2775 4.5005
R4040 VSS.n2745 VSS.n2744 4.5005
R4041 VSS.n2145 VSS.n2128 4.5005
R4042 VSS.n2196 VSS.n2194 4.5005
R4043 VSS.n2778 VSS.n2777 4.5005
R4044 VSS.n2113 VSS.n2109 4.5005
R4045 VSS.n2758 VSS.n2757 4.5005
R4046 VSS.n2183 VSS.n2182 4.5005
R4047 VSS.n2200 VSS.n2199 4.5005
R4048 VSS.n2147 VSS.n2144 4.5005
R4049 VSS.n2124 VSS.n2120 4.5005
R4050 VSS.n2736 VSS.n2735 4.5005
R4051 VSS.n2786 VSS.n2785 4.5005
R4052 VSS.n2134 VSS.n2114 4.5005
R4053 VSS.n2181 VSS.n2180 4.5005
R4054 VSS.n2767 VSS.n2766 4.5005
R4055 VSS.n2747 VSS.n2746 4.5005
R4056 VSS.n2202 VSS.n2201 4.5005
R4057 VSS.n2765 VSS.n2764 4.5005
R4058 VSS.n2721 VSS.n2720 4.5005
R4059 VSS.n2702 VSS.n2701 4.5005
R4060 VSS.n2282 VSS.n2278 4.5005
R4061 VSS.n2218 VSS.n2213 4.5005
R4062 VSS.n2246 VSS.n2237 4.5005
R4063 VSS.n2233 VSS.n2229 4.5005
R4064 VSS.n2291 VSS.n2290 4.5005
R4065 VSS.n2305 VSS.n2304 4.5005
R4066 VSS.n2302 VSS.n2270 4.5005
R4067 VSS.n2283 VSS.n2280 4.5005
R4068 VSS.n2700 VSS.n2699 4.5005
R4069 VSS.n2301 VSS.n2269 4.5005
R4070 VSS.n2300 VSS.n2299 4.5005
R4071 VSS.n2285 VSS.n2248 4.5005
R4072 VSS.n2231 VSS.n2221 4.5005
R4073 VSS.n2287 VSS.n2286 4.5005
R4074 VSS.n2665 VSS.n2664 4.5005
R4075 VSS.n2232 VSS.n2222 4.5005
R4076 VSS.n2710 VSS.n2709 4.5005
R4077 VSS.n2239 VSS.n2236 4.5005
R4078 VSS.n2313 VSS.n2281 4.5005
R4079 VSS.n2303 VSS.n2272 4.5005
R4080 VSS.n2217 VSS.n2214 4.5005
R4081 VSS.n2712 VSS.n2711 4.5005
R4082 VSS.n2677 VSS.n2676 4.5005
R4083 VSS.n2289 VSS.n2251 4.5005
R4084 VSS.n2298 VSS.n2254 4.5005
R4085 VSS.n2669 VSS.n2668 4.5005
R4086 VSS.n2690 VSS.n2689 4.5005
R4087 VSS.n2667 VSS.n2666 4.5005
R4088 VSS.n2228 VSS.n2224 4.5005
R4089 VSS.n2698 VSS.n2697 4.5005
R4090 VSS.n2288 VSS.n2249 4.5005
R4091 VSS.n2679 VSS.n2678 4.5005
R4092 VSS.n2244 VSS.n2238 4.5005
R4093 VSS.n2719 VSS.n2718 4.5005
R4094 VSS.n2655 VSS.n2654 4.5005
R4095 VSS.n2345 VSS.n2344 4.5005
R4096 VSS.n2631 VSS.n2630 4.5005
R4097 VSS.n2343 VSS.n2333 4.5005
R4098 VSS.n2391 VSS.n2390 4.5005
R4099 VSS.n2591 VSS.n2590 4.5005
R4100 VSS.n2566 VSS.n2404 4.5005
R4101 VSS.n2328 VSS.n2321 4.5005
R4102 VSS.n2643 VSS.n2642 4.5005
R4103 VSS.n2629 VSS.n2628 4.5005
R4104 VSS.n2403 VSS.n2401 4.5005
R4105 VSS.n2606 VSS.n2605 4.5005
R4106 VSS.n2622 VSS.n2621 4.5005
R4107 VSS.n2350 VSS.n2348 4.5005
R4108 VSS.n2604 VSS.n2603 4.5005
R4109 VSS.n2593 VSS.n2592 4.5005
R4110 VSS.n2618 VSS.n2363 4.5005
R4111 VSS.n2389 VSS.n2388 4.5005
R4112 VSS.n2620 VSS.n2619 4.5005
R4113 VSS.n2641 VSS.n2330 4.5005
R4114 VSS.n2645 VSS.n2644 4.5005
R4115 VSS.n2342 VSS.n2340 4.5005
R4116 VSS.n2347 VSS.n2341 4.5005
R4117 VSS.n2339 VSS.n2335 4.5005
R4118 VSS.n2386 VSS.n2384 4.5005
R4119 VSS.n2589 VSS.n2588 4.5005
R4120 VSS.n2565 VSS.n2405 4.5005
R4121 VSS.n2355 VSS.n2349 4.5005
R4122 VSS.n2608 VSS.n2607 4.5005
R4123 VSS.n2595 VSS.n2594 4.5005
R4124 VSS.n2334 VSS.n2327 4.5005
R4125 VSS.n2324 VSS.n2322 4.5005
R4126 VSS.n2406 VSS.n2402 4.5005
R4127 VSS.n2392 VSS.n2387 4.5005
R4128 VSS.n2617 VSS.n2616 4.5005
R4129 VSS.n2627 VSS.n2626 4.5005
R4130 VSS.n2602 VSS.n2601 4.5005
R4131 VSS.n2653 VSS.n2652 4.5005
R4132 VSS.n2529 VSS.n2528 4.5005
R4133 VSS.n2518 VSS.n2517 4.5005
R4134 VSS.n2428 VSS.n2427 4.5005
R4135 VSS.n2532 VSS.n2531 4.5005
R4136 VSS.n2520 VSS.n2519 4.5005
R4137 VSS.n2472 VSS.n2453 4.5005
R4138 VSS.n2489 VSS.n2481 4.5005
R4139 VSS.n2437 VSS.n2430 4.5005
R4140 VSS.n2557 VSS.n2414 4.5005
R4141 VSS.n2450 VSS.n2442 4.5005
R4142 VSS.n2506 VSS.n2505 4.5005
R4143 VSS.n2494 VSS.n2493 4.5005
R4144 VSS.n2559 VSS.n2558 4.5005
R4145 VSS.n2504 VSS.n2503 4.5005
R4146 VSS.n2417 VSS.n2415 4.5005
R4147 VSS.n2424 VSS.n2422 4.5005
R4148 VSS.n2508 VSS.n2507 4.5005
R4149 VSS.n2534 VSS.n2533 4.5005
R4150 VSS.n2476 VSS.n2473 4.5005
R4151 VSS.n2443 VSS.n2441 4.5005
R4152 VSS.n2452 VSS.n2448 4.5005
R4153 VSS.n2556 VSS.n2555 4.5005
R4154 VSS.n2470 VSS.n2454 4.5005
R4155 VSS.n2496 VSS.n2495 4.5005
R4156 VSS.n2449 VSS.n2444 4.5005
R4157 VSS.n2435 VSS.n2431 4.5005
R4158 VSS.n2490 VSS.n2482 4.5005
R4159 VSS.n2516 VSS.n2515 4.5005
R4160 VSS.n2420 VSS.n2419 4.5005
R4161 VSS.n2457 VSS.n2455 4.5005
R4162 VSS.n2536 VSS.n2535 4.5005
R4163 VSS.n2524 VSS.n2523 4.5005
R4164 VSS.n2537 VSS.n2432 4.5005
R4165 VSS.n2511 VSS.n2456 4.5005
R4166 VSS.n2480 VSS.n2478 4.5005
R4167 VSS.n2554 VSS.n2553 4.5005
R4168 VSS.n2510 VSS.n2509 4.5005
R4169 VSS.n2514 VSS.n2513 4.5005
R4170 VSS.n2446 VSS.n2445 4.5005
R4171 VSS.n2471 VSS.n2469 4.5005
R4172 VSS.n2551 VSS.n2550 4.5005
R4173 VSS.n2358 VSS.n2351 4.5005
R4174 VSS.n2615 VSS.n2614 4.5005
R4175 VSS.n2585 VSS.n2408 4.5005
R4176 VSS.n2409 VSS.n2407 4.5005
R4177 VSS.n2396 VSS.n2385 4.5005
R4178 VSS.n2647 VSS.n2646 4.5005
R4179 VSS.n2354 VSS.n2353 4.5005
R4180 VSS.n2636 VSS.n2337 4.5005
R4181 VSS.n2397 VSS.n2393 4.5005
R4182 VSS.n2587 VSS.n2586 4.5005
R4183 VSS.n2611 VSS.n2610 4.5005
R4184 VSS.n2370 VSS.n2369 4.5005
R4185 VSS.n2371 VSS.n2365 4.5005
R4186 VSS.n2336 VSS.n2326 4.5005
R4187 VSS.n2649 VSS.n2323 4.5005
R4188 VSS.n2400 VSS.n2398 4.5005
R4189 VSS.n2609 VSS.n2383 4.5005
R4190 VSS.n2357 VSS.n2356 4.5005
R4191 VSS.n2635 VSS.n2634 4.5005
R4192 VSS.n2651 VSS.n2650 4.5005
R4193 VSS.n2311 VSS.n2276 4.5005
R4194 VSS.n2245 VSS.n2243 4.5005
R4195 VSS.n2681 VSS.n2680 4.5005
R4196 VSS.n2717 VSS.n2716 4.5005
R4197 VSS.n2242 VSS.n2240 4.5005
R4198 VSS.n2315 VSS.n2314 4.5005
R4199 VSS.n2675 VSS.n2674 4.5005
R4200 VSS.n2688 VSS.n2687 4.5005
R4201 VSS.n2268 VSS.n2267 4.5005
R4202 VSS.n2708 VSS.n2707 4.5005
R4203 VSS.n2696 VSS.n2695 4.5005
R4204 VSS.n2273 VSS.n2271 4.5005
R4205 VSS.n2312 VSS.n2279 4.5005
R4206 VSS.n2686 VSS.n2685 4.5005
R4207 VSS.n2694 VSS.n2241 4.5005
R4208 VSS.n2715 VSS.n2215 4.5005
R4209 VSS.n2220 VSS.n2216 4.5005
R4210 VSS.n2225 VSS.n2223 4.5005
R4211 VSS.n2741 VSS.n2167 4.5005
R4212 VSS.n2206 VSS.n2198 4.5005
R4213 VSS.n2163 VSS.n2162 4.5005
R4214 VSS.n2759 VSS.n2123 4.5005
R4215 VSS.n2771 VSS.n2110 4.5005
R4216 VSS.n2121 VSS.n2116 4.5005
R4217 VSS.n2100 VSS.n2098 4.5005
R4218 VSS.n2770 VSS.n2769 4.5005
R4219 VSS.n2122 VSS.n2119 4.5005
R4220 VSS.n2160 VSS.n2146 4.5005
R4221 VSS.n2782 VSS.n2097 4.5005
R4222 VSS.n2203 VSS.n2173 4.5005
R4223 VSS.n2168 VSS.n2166 4.5005
R4224 VSS.n2749 VSS.n2748 4.5005
R4225 VSS.n2208 VSS.n2207 4.5005
R4226 VSS.n2743 VSS.n2742 4.5005
R4227 VSS.n2763 VSS.n2762 4.5005
R4228 VSS.n2111 VSS.n2104 4.5005
R4229 VSS.n2784 VSS.n2783 4.5005
R4230 VSS.n2205 VSS.n2204 4.5005
R4231 VSS.n2009 VSS.n2006 4.5005
R4232 VSS.n2863 VSS.n2862 4.5005
R4233 VSS.n2838 VSS.n2837 4.5005
R4234 VSS.n2043 VSS.n2042 4.5005
R4235 VSS.n2030 VSS.n2029 4.5005
R4236 VSS.n2049 VSS.n2044 4.5005
R4237 VSS.n2003 VSS.n1999 4.5005
R4238 VSS.n2872 VSS.n1998 4.5005
R4239 VSS.n2861 VSS.n2010 4.5005
R4240 VSS.n2075 VSS.n2064 4.5005
R4241 VSS.n2807 VSS.n2086 4.5005
R4242 VSS.n2832 VSS.n2062 4.5005
R4243 VSS.n2809 VSS.n2808 4.5005
R4244 VSS.n2076 VSS.n2072 4.5005
R4245 VSS.n2034 VSS.n2033 4.5005
R4246 VSS.n2834 VSS.n2833 4.5005
R4247 VSS.n2848 VSS.n2847 4.5005
R4248 VSS.n2084 VSS.n2077 4.5005
R4249 VSS.n2811 VSS.n2810 4.5005
R4250 VSS.n2874 VSS.n2873 4.5005
R4251 VSS.n4189 VSS.n4188 4.5005
R4252 VSS.n4149 VSS.n4148 4.5005
R4253 VSS.n4212 VSS.n4211 4.5005
R4254 VSS.n4211 VSS.n4210 4.5005
R4255 VSS.n4685 VSS.n4684 4.5005
R4256 VSS.n1416 VSS.n1415 4.5005
R4257 VSS.n4088 VSS.n4087 4.5005
R4258 VSS.n4087 VSS.n4086 4.5005
R4259 VSS.n4125 VSS.n4124 4.5005
R4260 VSS.n4124 VSS.n4123 4.5005
R4261 VSS.n966 VSS.n965 4.5005
R4262 VSS.n212 VSS.t345 4.44646
R4263 VSS.t154 VSS.t157 4.44646
R4264 VSS.n4137 VSS.n4136 4.25879
R4265 VSS.n919 VSS.n918 4.25822
R4266 VSS.t216 VSS.t151 4.12487
R4267 VSS.t151 VSS.t154 4.12487
R4268 VSS.n4717 VSS.t268 4.12487
R4269 VSS.n5885 VSS.n5837 4.11115
R4270 VSS.n5884 VSS.n5839 4.09159
R4271 VSS VSS.n5871 4.0484
R4272 VSS VSS.n5848 4.0484
R4273 VSS VSS.n5800 4.0484
R4274 VSS VSS.n5808 4.0484
R4275 VSS.n816 VSS.t556 4.04279
R4276 VSS.n841 VSS.t553 4.04279
R4277 VSS.n1457 VSS.t519 4.04279
R4278 VSS.n1473 VSS.t516 4.04279
R4279 VSS.n5797 VSS.n5773 3.98171
R4280 VSS.n911 VSS.n910 3.95365
R4281 VSS.n971 VSS.n970 3.95358
R4282 VSS.n5860 VSS.n5856 3.76876
R4283 VSS.n5861 VSS.n5854 3.76876
R4284 VSS.n5814 VSS.n5765 3.76876
R4285 VSS.n5813 VSS.n5767 3.76876
R4286 VSS.n5806 VSS.n5805 3.75997
R4287 VSS.n4199 VSS.t720 3.75122
R4288 VSS.n26 VSS.n24 3.68267
R4289 VSS.n5816 VSS.n5760 3.66898
R4290 VSS.n5865 VSS.n5864 3.66898
R4291 VSS.n5893 VSS.n4747 3.66898
R4292 VSS.n5763 VSS.n5762 3.66898
R4293 VSS.n5834 VSS.n5729 3.60687
R4294 VSS.n5878 VSS.n5845 3.60246
R4295 VSS.n5879 VSS.n5843 3.60246
R4296 VSS.n5793 VSS.n5775 3.60246
R4297 VSS.n5792 VSS.n5777 3.60246
R4298 VSS.n4274 VSS.n4273 3.59971
R4299 VSS.n5835 VSS.n5727 3.5873
R4300 VSS.n1029 VSS.n1028 3.48846
R4301 VSS.n1719 VSS.t762 3.45416
R4302 VSS.n1728 VSS.t433 3.45416
R4303 VSS.n1720 VSS.t434 3.45416
R4304 VSS.n1754 VSS.t49 3.41655
R4305 VSS.n2458 VSS.t103 3.41655
R4306 VSS.n2372 VSS.t25 3.41655
R4307 VSS.n2255 VSS.t55 3.41655
R4308 VSS.n2148 VSS.t8 3.41655
R4309 VSS.n2051 VSS.t85 3.41655
R4310 VSS.n1981 VSS.t84 3.41655
R4311 VSS.n1826 VSS.t81 3.41655
R4312 VSS.n1792 VSS.t36 3.41655
R4313 VSS.n1771 VSS.t32 3.41655
R4314 VSS.n1743 VSS.t59 3.41655
R4315 VSS.n4837 VSS.t767 3.41078
R4316 VSS.n4800 VSS.t529 3.41078
R4317 VSS.n4912 VSS.t425 3.41078
R4318 VSS.n4794 VSS.t591 3.41078
R4319 VSS.n5755 VSS.n5754 3.40289
R4320 VSS.n5827 VSS.n5748 3.40289
R4321 VSS.n1382 VSS.t249 3.38064
R4322 VSS.n4094 VSS.t753 3.38064
R4323 VSS.n922 VSS.n921 3.37941
R4324 VSS.n1414 VSS.n1411 3.37941
R4325 VSS.n1414 VSS.n1413 3.37941
R4326 VSS.n4013 VSS.n3986 3.37941
R4327 VSS.n835 VSS.n822 3.37941
R4328 VSS.n835 VSS.n824 3.37941
R4329 VSS.n4836 VSS.n4835 3.37941
R4330 VSS.n4799 VSS.n4798 3.37941
R4331 VSS.n4793 VSS.n4792 3.37941
R4332 VSS.n4911 VSS.n4910 3.37941
R4333 VSS.n4153 VSS.n4152 3.37941
R4334 VSS.n4708 VSS.n4705 3.37941
R4335 VSS.n4708 VSS.n4707 3.37941
R4336 VSS.n4116 VSS.n4115 3.3685
R4337 VSS.n4108 VSS.n4107 3.35882
R4338 VSS.n5735 VSS.n5734 3.3442
R4339 VSS.n5743 VSS.n5742 3.3442
R4340 VSS.n4509 VSS.t207 3.333
R4341 VSS.n5049 VSS.t182 3.33271
R4342 VSS.n76 VSS.t231 3.33057
R4343 VSS.n5047 VSS.t209 3.33036
R4344 VSS.n4948 VSS.t229 3.32608
R4345 VSS.n4947 VSS.t236 3.32608
R4346 VSS.n4908 VSS.t193 3.32608
R4347 VSS.n4790 VSS.t177 3.32608
R4348 VSS.n33 VSS.t180 3.32582
R4349 VSS.n32 VSS.t198 3.32582
R4350 VSS.n31 VSS.t214 3.32582
R4351 VSS.n58 VSS.t205 3.32582
R4352 VSS.n4789 VSS.t238 3.32512
R4353 VSS.n59 VSS.t149 3.32486
R4354 VSS.n4510 VSS.t196 3.31238
R4355 VSS.n5060 VSS.t174 3.31209
R4356 VSS.n63 VSS.t146 3.31186
R4357 VSS.n5046 VSS.t241 3.3116
R4358 VSS.n87 VSS.t188 3.31143
R4359 VSS.n5048 VSS.t137 3.31114
R4360 VSS.n231 VSS.t397 3.2765
R4361 VSS.n231 VSS.n230 3.2765
R4362 VSS.n234 VSS.t317 3.2765
R4363 VSS.n234 VSS.n233 3.2765
R4364 VSS.n237 VSS.t287 3.2765
R4365 VSS.n237 VSS.n236 3.2765
R4366 VSS.n179 VSS.t392 3.2765
R4367 VSS.n179 VSS.n178 3.2765
R4368 VSS.n182 VSS.t356 3.2765
R4369 VSS.n182 VSS.n181 3.2765
R4370 VSS.n176 VSS.t324 3.2765
R4371 VSS.n176 VSS.n175 3.2765
R4372 VSS.n172 VSS.t351 3.2765
R4373 VSS.n172 VSS.n171 3.2765
R4374 VSS.n169 VSS.t387 3.2765
R4375 VSS.n169 VSS.n168 3.2765
R4376 VSS.n125 VSS.t363 3.2765
R4377 VSS.n125 VSS.n124 3.2765
R4378 VSS.n129 VSS.t328 3.2765
R4379 VSS.n129 VSS.n128 3.2765
R4380 VSS.n133 VSS.t301 3.2765
R4381 VSS.n133 VSS.n132 3.2765
R4382 VSS.n136 VSS.t366 3.2765
R4383 VSS.n136 VSS.n135 3.2765
R4384 VSS.n139 VSS.t333 3.2765
R4385 VSS.n139 VSS.n138 3.2765
R4386 VSS.n223 VSS.t308 3.2765
R4387 VSS.n223 VSS.n222 3.2765
R4388 VSS.n227 VSS.t280 3.2765
R4389 VSS.n227 VSS.n226 3.2765
R4390 VSS.n921 VSS.t723 3.2765
R4391 VSS.n921 VSS.n920 3.2765
R4392 VSS.n1413 VSS.t533 3.2765
R4393 VSS.n1413 VSS.n1412 3.2765
R4394 VSS.n1411 VSS.t520 3.2765
R4395 VSS.n1411 VSS.n1410 3.2765
R4396 VSS.n3986 VSS.t544 3.2765
R4397 VSS.n3986 VSS.n3985 3.2765
R4398 VSS.n824 VSS.t557 3.2765
R4399 VSS.n824 VSS.n823 3.2765
R4400 VSS.n822 VSS.t706 3.2765
R4401 VSS.n822 VSS.n821 3.2765
R4402 VSS.n5166 VSS.t313 3.2765
R4403 VSS.n5166 VSS.n5165 3.2765
R4404 VSS.n5168 VSS.t384 3.2765
R4405 VSS.n5168 VSS.n5167 3.2765
R4406 VSS.n5170 VSS.t410 3.2765
R4407 VSS.n5170 VSS.n5169 3.2765
R4408 VSS.n5195 VSS.t386 3.2765
R4409 VSS.n5195 VSS.n5194 3.2765
R4410 VSS.n5193 VSS.t354 3.2765
R4411 VSS.n5193 VSS.n5192 3.2765
R4412 VSS.n5191 VSS.t329 3.2765
R4413 VSS.n5191 VSS.n5190 3.2765
R4414 VSS.n5187 VSS.t285 3.2765
R4415 VSS.n5187 VSS.n5186 3.2765
R4416 VSS.n5189 VSS.t400 3.2765
R4417 VSS.n5189 VSS.n5188 3.2765
R4418 VSS.n5162 VSS.t411 3.2765
R4419 VSS.n5162 VSS.n5161 3.2765
R4420 VSS.n5164 VSS.t385 3.2765
R4421 VSS.n5164 VSS.n5163 3.2765
R4422 VSS.n4775 VSS.t337 3.2765
R4423 VSS.n4775 VSS.n4774 3.2765
R4424 VSS.n4773 VSS.t307 3.2765
R4425 VSS.n4773 VSS.n4772 3.2765
R4426 VSS.n4771 VSS.t405 3.2765
R4427 VSS.n4771 VSS.n4770 3.2765
R4428 VSS.n4769 VSS.t334 3.2765
R4429 VSS.n4769 VSS.n4768 3.2765
R4430 VSS.n4767 VSS.t357 3.2765
R4431 VSS.n4767 VSS.n4766 3.2765
R4432 VSS.n4835 VSS.t768 3.2765
R4433 VSS.n4835 VSS.n4834 3.2765
R4434 VSS.n4798 VSS.t530 3.2765
R4435 VSS.n4798 VSS.n4797 3.2765
R4436 VSS.n4792 VSS.t592 3.2765
R4437 VSS.n4792 VSS.n4791 3.2765
R4438 VSS.n4910 VSS.t426 3.2765
R4439 VSS.n4910 VSS.n4909 3.2765
R4440 VSS.n4152 VSS.t738 3.2765
R4441 VSS.n4152 VSS.n4151 3.2765
R4442 VSS.n4707 VSS.t688 3.2765
R4443 VSS.n4707 VSS.n4706 3.2765
R4444 VSS.n4705 VSS.t267 3.2765
R4445 VSS.n4705 VSS.n4704 3.2765
R4446 VSS.n5754 VSS.t631 3.2765
R4447 VSS.n5754 VSS.n5753 3.2765
R4448 VSS.n5748 VSS.t430 3.2765
R4449 VSS.n5748 VSS.n5747 3.2765
R4450 VSS.n5734 VSS.t573 3.2765
R4451 VSS.n5734 VSS.n5733 3.2765
R4452 VSS.n5727 VSS.t584 3.2765
R4453 VSS.n5727 VSS.n5726 3.2765
R4454 VSS.n5839 VSS.t477 3.2765
R4455 VSS.n5839 VSS.n5838 3.2765
R4456 VSS.n5837 VSS.t448 3.2765
R4457 VSS.n5837 VSS.n5836 3.2765
R4458 VSS.n5729 VSS.t585 3.2765
R4459 VSS.n5729 VSS.n5728 3.2765
R4460 VSS.n5742 VSS.t488 3.2765
R4461 VSS.n5742 VSS.n5741 3.2765
R4462 VSS.n4744 VSS.n4742 3.17523
R4463 VSS.n140 VSS.n139 3.1505
R4464 VSS.n137 VSS.n136 3.1505
R4465 VSS.n130 VSS.n129 3.1505
R4466 VSS.n228 VSS.n227 3.1505
R4467 VSS.n173 VSS.n172 3.1505
R4468 VSS.n183 VSS.n182 3.1505
R4469 VSS.n180 VSS.n179 3.1505
R4470 VSS.n238 VSS.n237 3.1505
R4471 VSS.n235 VSS.n234 3.1505
R4472 VSS.n5175 VSS.n5164 3.1505
R4473 VSS.n5176 VSS.n5162 3.1505
R4474 VSS.n5201 VSS.n5189 3.1505
R4475 VSS.n5202 VSS.n5187 3.1505
R4476 VSS.n5198 VSS.n5193 3.1505
R4477 VSS.n4782 VSS.n4767 3.1505
R4478 VSS.n4781 VSS.n4769 3.1505
R4479 VSS.n4778 VSS.n4773 3.1505
R4480 VSS.n5172 VSS.n5168 3.1505
R4481 VSS.n5945 VSS.n5944 3.08765
R4482 VSS.n4681 VSS.n4680 3.07743
R4483 VSS.n4124 VSS.n916 2.9883
R4484 VSS.n4087 VSS.n1397 2.9883
R4485 VSS.n4744 VSS.n4743 2.91648
R4486 VSS.n4976 VSS.n4975 2.83943
R4487 VSS.n4972 VSS.n4971 2.83943
R4488 VSS.n4968 VSS.n4967 2.83943
R4489 VSS.n4678 VSS.n4677 2.83943
R4490 VSS.n4675 VSS.n4674 2.83943
R4491 VSS.n4661 VSS.n4660 2.83943
R4492 VSS.n4583 VSS.n4582 2.83943
R4493 VSS.n4587 VSS.n4586 2.83943
R4494 VSS.n1311 VSS.n1310 2.81354
R4495 VSS.n3914 VSS.n3908 2.7874
R4496 VSS.n4236 VSS.n4235 2.75024
R4497 VSS.n1021 VSS.n1017 2.65705
R4498 VSS.n1021 VSS.n1020 2.65638
R4499 VSS.n4843 VSS.n4842 2.64393
R4500 VSS.n4805 VSS.n4804 2.64393
R4501 VSS.n134 VSS.n133 2.6255
R4502 VSS.n170 VSS.n169 2.6255
R4503 VSS.n177 VSS.n176 2.6255
R4504 VSS.n232 VSS.n231 2.6255
R4505 VSS.n5200 VSS.n5191 2.6255
R4506 VSS.n4780 VSS.n4771 2.6255
R4507 VSS.n5171 VSS.n5170 2.6255
R4508 VSS.n5174 VSS.n5166 2.6255
R4509 VSS.n5443 VSS.n5403 2.61042
R4510 VSS.n5427 VSS.n5405 2.61042
R4511 VSS.n5538 VSS.n5457 2.61042
R4512 VSS.n5602 VSS.n5601 2.60873
R4513 VSS.n4064 VSS.n1399 2.60616
R4514 VSS.n4040 VSS.n4039 2.60562
R4515 VSS.n1424 VSS.n1421 2.60491
R4516 VSS.n1481 VSS.n1480 2.60491
R4517 VSS.n796 VSS.n793 2.60491
R4518 VSS.n862 VSS.n861 2.60491
R4519 VSS.n4761 VSS.n4760 2.60246
R4520 VSS.n5308 VSS.n5307 2.60244
R4521 VSS.n5287 VSS.n5283 2.60244
R4522 VSS.n117 VSS.n110 2.60148
R4523 VSS.n4411 VSS.n4394 2.60147
R4524 VSS.n1308 VSS.n958 2.6005
R4525 VSS.n958 VSS.n957 2.6005
R4526 VSS.n1324 VSS.n1323 2.6005
R4527 VSS.n1323 VSS.n1322 2.6005
R4528 VSS.n1320 VSS.n1319 2.6005
R4529 VSS.n1319 VSS.n1318 2.6005
R4530 VSS.n1316 VSS.n1315 2.6005
R4531 VSS.n1315 VSS.n1314 2.6005
R4532 VSS.n1313 VSS.n1312 2.6005
R4533 VSS.n1312 VSS.n1311 2.6005
R4534 VSS.n1326 VSS.n1325 2.6005
R4535 VSS.n926 VSS.n925 2.6005
R4536 VSS.n929 VSS.n928 2.6005
R4537 VSS.n931 VSS.n930 2.6005
R4538 VSS.n933 VSS.n932 2.6005
R4539 VSS VSS.n935 2.6005
R4540 VSS.n937 VSS.n936 2.6005
R4541 VSS.n942 VSS.n941 2.6005
R4542 VSS.n945 VSS.n944 2.6005
R4543 VSS.n947 VSS.n946 2.6005
R4544 VSS.n950 VSS.n949 2.6005
R4545 VSS.n1340 VSS.n1339 2.6005
R4546 VSS.n1338 VSS.n1337 2.6005
R4547 VSS.n1336 VSS.n1335 2.6005
R4548 VSS.n1332 VSS.n1331 2.6005
R4549 VSS.n1330 VSS.n1329 2.6005
R4550 VSS.n1403 VSS.n1400 2.6005
R4551 VSS.n1520 VSS.n1517 2.6005
R4552 VSS.n4002 VSS.n3999 2.6005
R4553 VSS.n4012 VSS.n4009 2.6005
R4554 VSS.n4025 VSS.n4023 2.6005
R4555 VSS.n3984 VSS.n3983 2.6005
R4556 VSS.n3983 VSS.n3982 2.6005
R4557 VSS.n4030 VSS.n4029 2.6005
R4558 VSS.n4029 VSS.n4028 2.6005
R4559 VSS.n4026 VSS.n4025 2.6005
R4560 VSS.n4019 VSS.n4018 2.6005
R4561 VSS.n4018 VSS.n4017 2.6005
R4562 VSS VSS.n4012 2.6005
R4563 VSS.n4007 VSS.n4006 2.6005
R4564 VSS.n4006 VSS.n4005 2.6005
R4565 VSS.n4003 VSS.n4002 2.6005
R4566 VSS.n3993 VSS.n3992 2.6005
R4567 VSS.n3992 VSS.n3991 2.6005
R4568 VSS.n1521 VSS.n1520 2.6005
R4569 VSS.n3980 VSS.n3979 2.6005
R4570 VSS.n3979 VSS.n3978 2.6005
R4571 VSS.n4994 VSS.n4788 2.6005
R4572 VSS.n4788 VSS.n4787 2.6005
R4573 VSS.n4986 VSS.n4985 2.6005
R4574 VSS.n4985 VSS.n4984 2.6005
R4575 VSS.n4989 VSS.n4988 2.6005
R4576 VSS.n4988 VSS.n4987 2.6005
R4577 VSS.n4993 VSS.n4992 2.6005
R4578 VSS.n4992 VSS.n4991 2.6005
R4579 VSS.n5000 VSS.n4999 2.6005
R4580 VSS.n4999 VSS.n4998 2.6005
R4581 VSS.n4956 VSS.n4955 2.6005
R4582 VSS.n5469 VSS.n5468 2.6005
R4583 VSS.n5468 VSS.n5467 2.6005
R4584 VSS.n5466 VSS.n5465 2.6005
R4585 VSS.n5465 VSS.n5464 2.6005
R4586 VSS.n4952 VSS.n4951 2.6005
R4587 VSS.n4951 VSS.n4950 2.6005
R4588 VSS.n4955 VSS.n4954 2.6005
R4589 VSS.n5472 VSS.n5471 2.6005
R4590 VSS.n5471 VSS.n5470 2.6005
R4591 VSS.n4959 VSS.n4958 2.6005
R4592 VSS.n4958 VSS.n4957 2.6005
R4593 VSS.n4963 VSS.n4962 2.6005
R4594 VSS.n4965 VSS.n4964 2.6005
R4595 VSS.n4969 VSS.n4968 2.6005
R4596 VSS.n4973 VSS.n4972 2.6005
R4597 VSS.n4876 VSS.n4875 2.6005
R4598 VSS.n4875 VSS.n4874 2.6005
R4599 VSS.n4880 VSS.n4879 2.6005
R4600 VSS.n4879 VSS.n4878 2.6005
R4601 VSS.n4883 VSS.n4882 2.6005
R4602 VSS.n4882 VSS.n4881 2.6005
R4603 VSS.n4886 VSS.n4885 2.6005
R4604 VSS.n4885 VSS.n4884 2.6005
R4605 VSS.n4887 VSS.n4795 2.6005
R4606 VSS.n4795 VSS.n4794 2.6005
R4607 VSS.n4889 VSS 2.6005
R4608 VSS.n4889 VSS.n4888 2.6005
R4609 VSS.n4892 VSS.n4891 2.6005
R4610 VSS.n4891 VSS.n4890 2.6005
R4611 VSS.n4895 VSS.n4894 2.6005
R4612 VSS.n4894 VSS.n4893 2.6005
R4613 VSS.n4900 VSS.n4899 2.6005
R4614 VSS.n4899 VSS.n4898 2.6005
R4615 VSS.n4903 VSS.n4902 2.6005
R4616 VSS.n4902 VSS.n4901 2.6005
R4617 VSS.n4907 VSS.n4906 2.6005
R4618 VSS.n4906 VSS.n4905 2.6005
R4619 VSS.n4977 VSS.n4976 2.6005
R4620 VSS.n4982 VSS.n4981 2.6005
R4621 VSS.n4871 VSS.n4870 2.6005
R4622 VSS.n4870 VSS.n4869 2.6005
R4623 VSS.n4846 VSS.n4845 2.6005
R4624 VSS.n4845 VSS.n4844 2.6005
R4625 VSS.n4849 VSS.n4848 2.6005
R4626 VSS.n4848 VSS.n4847 2.6005
R4627 VSS.n4852 VSS.n4851 2.6005
R4628 VSS.n4851 VSS.n4850 2.6005
R4629 VSS.n4853 VSS.n4838 2.6005
R4630 VSS.n4838 VSS.n4837 2.6005
R4631 VSS.n4855 VSS 2.6005
R4632 VSS.n4855 VSS.n4854 2.6005
R4633 VSS.n4858 VSS.n4857 2.6005
R4634 VSS.n4857 VSS.n4856 2.6005
R4635 VSS.n4861 VSS.n4860 2.6005
R4636 VSS.n4860 VSS.n4859 2.6005
R4637 VSS.n4864 VSS.n4863 2.6005
R4638 VSS.n4863 VSS.n4862 2.6005
R4639 VSS.n4867 VSS.n4866 2.6005
R4640 VSS.n4866 VSS.n4865 2.6005
R4641 VSS.n4842 VSS.n4841 2.6005
R4642 VSS.n4804 VSS.n4803 2.6005
R4643 VSS.n4808 VSS.n4807 2.6005
R4644 VSS.n4807 VSS.n4806 2.6005
R4645 VSS.n4811 VSS.n4810 2.6005
R4646 VSS.n4810 VSS.n4809 2.6005
R4647 VSS.n4814 VSS.n4813 2.6005
R4648 VSS.n4813 VSS.n4812 2.6005
R4649 VSS.n4815 VSS.n4801 2.6005
R4650 VSS.n4801 VSS.n4800 2.6005
R4651 VSS.n4817 VSS 2.6005
R4652 VSS.n4817 VSS.n4816 2.6005
R4653 VSS.n4820 VSS.n4819 2.6005
R4654 VSS.n4819 VSS.n4818 2.6005
R4655 VSS.n4823 VSS.n4822 2.6005
R4656 VSS.n4822 VSS.n4821 2.6005
R4657 VSS.n4826 VSS.n4825 2.6005
R4658 VSS.n4825 VSS.n4824 2.6005
R4659 VSS.n4829 VSS.n4828 2.6005
R4660 VSS.n4828 VSS.n4827 2.6005
R4661 VSS.n4833 VSS.n4832 2.6005
R4662 VSS.n4832 VSS.n4831 2.6005
R4663 VSS.n4917 VSS.n4916 2.6005
R4664 VSS.n4916 VSS.n4915 2.6005
R4665 VSS.n4921 VSS.n4920 2.6005
R4666 VSS.n4920 VSS.n4919 2.6005
R4667 VSS.n4924 VSS.n4923 2.6005
R4668 VSS.n4923 VSS.n4922 2.6005
R4669 VSS.n4927 VSS.n4926 2.6005
R4670 VSS.n4926 VSS.n4925 2.6005
R4671 VSS.n4928 VSS.n4913 2.6005
R4672 VSS.n4913 VSS.n4912 2.6005
R4673 VSS.n4930 VSS 2.6005
R4674 VSS.n4930 VSS.n4929 2.6005
R4675 VSS.n4933 VSS.n4932 2.6005
R4676 VSS.n4932 VSS.n4931 2.6005
R4677 VSS.n4936 VSS.n4935 2.6005
R4678 VSS.n4935 VSS.n4934 2.6005
R4679 VSS.n4939 VSS.n4938 2.6005
R4680 VSS.n4938 VSS.n4937 2.6005
R4681 VSS.n4942 VSS.n4941 2.6005
R4682 VSS.n4941 VSS.n4940 2.6005
R4683 VSS.n4946 VSS.n4945 2.6005
R4684 VSS.n4945 VSS.n4944 2.6005
R4685 VSS.n470 VSS.n469 2.6005
R4686 VSS.n862 VSS.n858 2.6005
R4687 VSS.n858 VSS.n857 2.6005
R4688 VSS.n800 VSS.n799 2.6005
R4689 VSS.n799 VSS.n798 2.6005
R4690 VSS.n806 VSS.n805 2.6005
R4691 VSS.n805 VSS.n804 2.6005
R4692 VSS.n812 VSS.n811 2.6005
R4693 VSS.n811 VSS.n810 2.6005
R4694 VSS.n818 VSS.n817 2.6005
R4695 VSS.n817 VSS.n816 2.6005
R4696 VSS.n837 VSS 2.6005
R4697 VSS.n837 VSS.n836 2.6005
R4698 VSS.n840 VSS.n839 2.6005
R4699 VSS.n839 VSS.n838 2.6005
R4700 VSS.n846 VSS.n845 2.6005
R4701 VSS.n845 VSS.n844 2.6005
R4702 VSS.n853 VSS.n852 2.6005
R4703 VSS.n852 VSS.n851 2.6005
R4704 VSS.n869 VSS.n868 2.6005
R4705 VSS.n868 VSS.n867 2.6005
R4706 VSS.n793 VSS.n792 2.6005
R4707 VSS.n834 VSS.n831 2.6005
R4708 VSS.n803 VSS.n802 2.6005
R4709 VSS.n802 VSS.n801 2.6005
R4710 VSS.n809 VSS.n808 2.6005
R4711 VSS.n808 VSS.n807 2.6005
R4712 VSS.n815 VSS.n814 2.6005
R4713 VSS.n814 VSS.n813 2.6005
R4714 VSS.n828 VSS.n827 2.6005
R4715 VSS VSS.n834 2.6005
R4716 VSS.n843 VSS.n842 2.6005
R4717 VSS.n842 VSS.n841 2.6005
R4718 VSS.n850 VSS.n849 2.6005
R4719 VSS.n849 VSS.n848 2.6005
R4720 VSS.n856 VSS.n855 2.6005
R4721 VSS.n855 VSS.n854 2.6005
R4722 VSS.n866 VSS.n865 2.6005
R4723 VSS.n865 VSS.n864 2.6005
R4724 VSS.n861 VSS.n860 2.6005
R4725 VSS.n796 VSS.n795 2.6005
R4726 VSS.n795 VSS.n794 2.6005
R4727 VSS.n257 VSS.n256 2.6005
R4728 VSS.n342 VSS.n339 2.6005
R4729 VSS.n343 VSS.n342 2.6005
R4730 VSS.n4049 VSS.n4048 2.6005
R4731 VSS.n4067 VSS.n4066 2.6005
R4732 VSS.n4066 VSS.n4065 2.6005
R4733 VSS.n1399 VSS.n1398 2.6005
R4734 VSS.n4063 VSS.n4062 2.6005
R4735 VSS.n4062 VSS.n4061 2.6005
R4736 VSS.n4060 VSS.n4059 2.6005
R4737 VSS.n4059 VSS.n4058 2.6005
R4738 VSS.n4057 VSS.n4056 2.6005
R4739 VSS.n4056 VSS.n4055 2.6005
R4740 VSS.n4053 VSS.n4052 2.6005
R4741 VSS.n4052 VSS.n4051 2.6005
R4742 VSS.n4048 VSS.n4047 2.6005
R4743 VSS.n371 VSS.n370 2.6005
R4744 VSS.n370 VSS.n369 2.6005
R4745 VSS.n374 VSS.n373 2.6005
R4746 VSS.n373 VSS.n372 2.6005
R4747 VSS.n377 VSS.n376 2.6005
R4748 VSS.n376 VSS.n375 2.6005
R4749 VSS.n380 VSS.n379 2.6005
R4750 VSS.n379 VSS.n378 2.6005
R4751 VSS.n383 VSS.n382 2.6005
R4752 VSS.n382 VSS.n381 2.6005
R4753 VSS.n386 VSS.n385 2.6005
R4754 VSS.n385 VSS.n384 2.6005
R4755 VSS.n389 VSS.n388 2.6005
R4756 VSS.n388 VSS.n387 2.6005
R4757 VSS.n393 VSS.n392 2.6005
R4758 VSS.n392 VSS.n391 2.6005
R4759 VSS.n396 VSS.n395 2.6005
R4760 VSS.n395 VSS.n394 2.6005
R4761 VSS.n399 VSS.n398 2.6005
R4762 VSS.n398 VSS.n397 2.6005
R4763 VSS.n402 VSS.n401 2.6005
R4764 VSS.n401 VSS.n400 2.6005
R4765 VSS.n405 VSS.n404 2.6005
R4766 VSS.n404 VSS.n403 2.6005
R4767 VSS.n409 VSS.n408 2.6005
R4768 VSS.n408 VSS.n407 2.6005
R4769 VSS.n412 VSS.n411 2.6005
R4770 VSS.n411 VSS.n410 2.6005
R4771 VSS.n416 VSS.n415 2.6005
R4772 VSS.n415 VSS.n414 2.6005
R4773 VSS.n419 VSS.n418 2.6005
R4774 VSS.n418 VSS.n417 2.6005
R4775 VSS.n422 VSS.n421 2.6005
R4776 VSS.n421 VSS.n420 2.6005
R4777 VSS.n427 VSS.n426 2.6005
R4778 VSS.n426 VSS.n425 2.6005
R4779 VSS.n430 VSS.n429 2.6005
R4780 VSS.n429 VSS.n428 2.6005
R4781 VSS.n433 VSS.n432 2.6005
R4782 VSS.n432 VSS.n431 2.6005
R4783 VSS.n436 VSS.n435 2.6005
R4784 VSS.n435 VSS.n434 2.6005
R4785 VSS.n439 VSS.n438 2.6005
R4786 VSS.n438 VSS.n437 2.6005
R4787 VSS.n442 VSS.n441 2.6005
R4788 VSS.n441 VSS.n440 2.6005
R4789 VSS.n445 VSS.n444 2.6005
R4790 VSS.n444 VSS.n443 2.6005
R4791 VSS.n448 VSS.n447 2.6005
R4792 VSS.n447 VSS.n446 2.6005
R4793 VSS.n451 VSS.n450 2.6005
R4794 VSS.n450 VSS.n449 2.6005
R4795 VSS.n454 VSS.n453 2.6005
R4796 VSS.n453 VSS.n452 2.6005
R4797 VSS.n458 VSS.n457 2.6005
R4798 VSS.n457 VSS.n456 2.6005
R4799 VSS.n461 VSS.n460 2.6005
R4800 VSS.n460 VSS.n459 2.6005
R4801 VSS.n464 VSS.n463 2.6005
R4802 VSS.n463 VSS.n462 2.6005
R4803 VSS.n473 VSS.n472 2.6005
R4804 VSS.n472 VSS.n471 2.6005
R4805 VSS.n476 VSS.n475 2.6005
R4806 VSS.n475 VSS.n474 2.6005
R4807 VSS.n479 VSS.n478 2.6005
R4808 VSS.n478 VSS.n477 2.6005
R4809 VSS.n482 VSS.n481 2.6005
R4810 VSS.n481 VSS.n480 2.6005
R4811 VSS.n485 VSS.n484 2.6005
R4812 VSS.n484 VSS.n483 2.6005
R4813 VSS.n487 VSS.n486 2.6005
R4814 VSS.n491 VSS.n490 2.6005
R4815 VSS.n493 VSS.n492 2.6005
R4816 VSS.n763 VSS.n762 2.6005
R4817 VSS.n716 VSS.n715 2.6005
R4818 VSS.n715 VSS.n714 2.6005
R4819 VSS.n762 VSS.n761 2.6005
R4820 VSS.n760 VSS.n759 2.6005
R4821 VSS.n759 VSS.n758 2.6005
R4822 VSS.n757 VSS.n756 2.6005
R4823 VSS.n756 VSS.n755 2.6005
R4824 VSS.n754 VSS.n753 2.6005
R4825 VSS.n753 VSS.n752 2.6005
R4826 VSS.n732 VSS.n731 2.6005
R4827 VSS.n731 VSS.n730 2.6005
R4828 VSS.n728 VSS.n727 2.6005
R4829 VSS.n727 VSS.n726 2.6005
R4830 VSS.n725 VSS.n724 2.6005
R4831 VSS.n724 VSS.n723 2.6005
R4832 VSS.n722 VSS.n721 2.6005
R4833 VSS.n721 VSS.n720 2.6005
R4834 VSS.n719 VSS.n718 2.6005
R4835 VSS.n718 VSS.n717 2.6005
R4836 VSS.n497 VSS.n496 2.6005
R4837 VSS.n496 VSS.n495 2.6005
R4838 VSS.n500 VSS.n499 2.6005
R4839 VSS.n502 VSS.n501 2.6005
R4840 VSS.n5336 VSS.n5335 2.6005
R4841 VSS.n5332 VSS.n5331 2.6005
R4842 VSS.n5329 VSS.n5328 2.6005
R4843 VSS.n5326 VSS.n5325 2.6005
R4844 VSS.n5324 VSS.n5323 2.6005
R4845 VSS.n5321 VSS.n5320 2.6005
R4846 VSS.n5320 VSS.n5319 2.6005
R4847 VSS.n5317 VSS.n5316 2.6005
R4848 VSS.n5316 VSS.n5315 2.6005
R4849 VSS.n514 VSS.n513 2.6005
R4850 VSS.n513 VSS.n512 2.6005
R4851 VSS.n517 VSS.n516 2.6005
R4852 VSS.n516 VSS.n515 2.6005
R4853 VSS.n520 VSS.n519 2.6005
R4854 VSS.n519 VSS.n518 2.6005
R4855 VSS.n523 VSS.n522 2.6005
R4856 VSS.n522 VSS.n521 2.6005
R4857 VSS.n526 VSS.n525 2.6005
R4858 VSS.n525 VSS.n524 2.6005
R4859 VSS.n530 VSS.n529 2.6005
R4860 VSS.n529 VSS.n528 2.6005
R4861 VSS.n533 VSS.n532 2.6005
R4862 VSS.n532 VSS.n531 2.6005
R4863 VSS.n536 VSS.n535 2.6005
R4864 VSS.n535 VSS.n534 2.6005
R4865 VSS.n539 VSS.n538 2.6005
R4866 VSS.n538 VSS.n537 2.6005
R4867 VSS.n542 VSS.n541 2.6005
R4868 VSS.n541 VSS.n540 2.6005
R4869 VSS.n545 VSS.n544 2.6005
R4870 VSS.n544 VSS.n543 2.6005
R4871 VSS.n548 VSS.n547 2.6005
R4872 VSS.n547 VSS.n546 2.6005
R4873 VSS.n551 VSS.n550 2.6005
R4874 VSS.n550 VSS.n549 2.6005
R4875 VSS.n554 VSS.n553 2.6005
R4876 VSS.n556 VSS.n555 2.6005
R4877 VSS.n559 VSS.n558 2.6005
R4878 VSS.n562 VSS.n561 2.6005
R4879 VSS.n566 VSS.n565 2.6005
R4880 VSS.n571 VSS.n570 2.6005
R4881 VSS.n570 VSS.n569 2.6005
R4882 VSS.n574 VSS.n573 2.6005
R4883 VSS.n573 VSS.n572 2.6005
R4884 VSS.n577 VSS.n576 2.6005
R4885 VSS.n576 VSS.n575 2.6005
R4886 VSS.n580 VSS.n579 2.6005
R4887 VSS.n579 VSS.n578 2.6005
R4888 VSS.n583 VSS.n582 2.6005
R4889 VSS.n582 VSS.n581 2.6005
R4890 VSS.n586 VSS.n585 2.6005
R4891 VSS.n585 VSS.n584 2.6005
R4892 VSS.n589 VSS.n588 2.6005
R4893 VSS.n588 VSS.n587 2.6005
R4894 VSS.n593 VSS.n592 2.6005
R4895 VSS.n592 VSS.n591 2.6005
R4896 VSS.n595 VSS.n594 2.6005
R4897 VSS.n598 VSS.n597 2.6005
R4898 VSS.n601 VSS.n600 2.6005
R4899 VSS.n600 VSS.n599 2.6005
R4900 VSS.n604 VSS.n603 2.6005
R4901 VSS.n603 VSS.n602 2.6005
R4902 VSS.n607 VSS.n606 2.6005
R4903 VSS.n606 VSS.n605 2.6005
R4904 VSS.n610 VSS.n609 2.6005
R4905 VSS.n609 VSS.n608 2.6005
R4906 VSS.n613 VSS.n612 2.6005
R4907 VSS.n612 VSS.n611 2.6005
R4908 VSS.n616 VSS.n615 2.6005
R4909 VSS.n615 VSS.n614 2.6005
R4910 VSS.n619 VSS.n618 2.6005
R4911 VSS.n618 VSS.n617 2.6005
R4912 VSS.n622 VSS.n621 2.6005
R4913 VSS.n621 VSS.n620 2.6005
R4914 VSS.n625 VSS.n624 2.6005
R4915 VSS.n624 VSS.n623 2.6005
R4916 VSS.n628 VSS.n627 2.6005
R4917 VSS.n627 VSS.n626 2.6005
R4918 VSS.n631 VSS.n630 2.6005
R4919 VSS.n630 VSS.n629 2.6005
R4920 VSS.n634 VSS.n633 2.6005
R4921 VSS.n633 VSS.n632 2.6005
R4922 VSS.n637 VSS.n636 2.6005
R4923 VSS.n636 VSS.n635 2.6005
R4924 VSS.n640 VSS.n639 2.6005
R4925 VSS.n639 VSS.n638 2.6005
R4926 VSS.n643 VSS.n642 2.6005
R4927 VSS.n642 VSS.n641 2.6005
R4928 VSS.n646 VSS.n645 2.6005
R4929 VSS.n645 VSS.n644 2.6005
R4930 VSS.n649 VSS.n648 2.6005
R4931 VSS.n648 VSS.n647 2.6005
R4932 VSS.n652 VSS.n651 2.6005
R4933 VSS.n651 VSS.n650 2.6005
R4934 VSS.n655 VSS.n654 2.6005
R4935 VSS.n654 VSS.n653 2.6005
R4936 VSS.n658 VSS.n657 2.6005
R4937 VSS.n657 VSS.n656 2.6005
R4938 VSS.n661 VSS.n660 2.6005
R4939 VSS.n660 VSS.n659 2.6005
R4940 VSS.n664 VSS.n663 2.6005
R4941 VSS.n663 VSS.n662 2.6005
R4942 VSS.n667 VSS.n666 2.6005
R4943 VSS.n666 VSS.n665 2.6005
R4944 VSS.n670 VSS.n669 2.6005
R4945 VSS.n669 VSS.n668 2.6005
R4946 VSS.n673 VSS.n672 2.6005
R4947 VSS.n675 VSS.n674 2.6005
R4948 VSS.n678 VSS.n677 2.6005
R4949 VSS.n681 VSS.n680 2.6005
R4950 VSS.n685 VSS.n684 2.6005
R4951 VSS.n691 VSS.n690 2.6005
R4952 VSS.n687 VSS.n686 2.6005
R4953 VSS.n735 VSS.n734 2.6005
R4954 VSS.n734 VSS.n733 2.6005
R4955 VSS.n713 VSS.n712 2.6005
R4956 VSS.n712 VSS.n711 2.6005
R4957 VSS.n710 VSS.n709 2.6005
R4958 VSS.n709 VSS.n708 2.6005
R4959 VSS.n707 VSS.n706 2.6005
R4960 VSS.n706 VSS.n705 2.6005
R4961 VSS.n704 VSS.n703 2.6005
R4962 VSS.n703 VSS.n702 2.6005
R4963 VSS.n506 VSS.n505 2.6005
R4964 VSS.n509 VSS.n508 2.6005
R4965 VSS.n700 VSS.n699 2.6005
R4966 VSS.n699 VSS.n698 2.6005
R4967 VSS.n697 VSS.n696 2.6005
R4968 VSS.n696 VSS.n695 2.6005
R4969 VSS.n694 VSS.n693 2.6005
R4970 VSS.n693 VSS.n692 2.6005
R4971 VSS.n775 VSS.n255 2.6005
R4972 VSS.n255 VSS.n254 2.6005
R4973 VSS.n787 VSS.n786 2.6005
R4974 VSS.n786 VSS.n785 2.6005
R4975 VSS.n784 VSS.n783 2.6005
R4976 VSS.n783 VSS.n782 2.6005
R4977 VSS.n781 VSS.n780 2.6005
R4978 VSS.n780 VSS.n779 2.6005
R4979 VSS.n778 VSS.n777 2.6005
R4980 VSS.n777 VSS.n776 2.6005
R4981 VSS.n751 VSS.n750 2.6005
R4982 VSS.n750 VSS.n749 2.6005
R4983 VSS.n748 VSS.n747 2.6005
R4984 VSS.n747 VSS.n746 2.6005
R4985 VSS.n745 VSS.n744 2.6005
R4986 VSS.n744 VSS.n743 2.6005
R4987 VSS.n742 VSS.n741 2.6005
R4988 VSS.n741 VSS.n740 2.6005
R4989 VSS.n739 VSS.n738 2.6005
R4990 VSS.n738 VSS.n737 2.6005
R4991 VSS.n770 VSS.n769 2.6005
R4992 VSS.n769 VSS.n768 2.6005
R4993 VSS.n773 VSS.n772 2.6005
R4994 VSS.n772 VSS.n771 2.6005
R4995 VSS.n766 VSS.n765 2.6005
R4996 VSS.n765 VSS.n764 2.6005
R4997 VSS.n4298 VSS.n4297 2.6005
R4998 VSS.n4297 VSS.n4296 2.6005
R4999 VSS.n4295 VSS.n4294 2.6005
R5000 VSS.n4294 VSS.n4293 2.6005
R5001 VSS.n4292 VSS.n4291 2.6005
R5002 VSS.n4291 VSS.n4290 2.6005
R5003 VSS.n4289 VSS.n4288 2.6005
R5004 VSS.n4288 VSS.n4287 2.6005
R5005 VSS.n4301 VSS.n4300 2.6005
R5006 VSS.n4312 VSS.n4311 2.6005
R5007 VSS.n4307 VSS.n4306 2.6005
R5008 VSS.n1174 VSS.n1173 2.6005
R5009 VSS.n1173 VSS.n1172 2.6005
R5010 VSS.n1178 VSS.n1177 2.6005
R5011 VSS.n1177 VSS.n1176 2.6005
R5012 VSS.n1181 VSS.n1180 2.6005
R5013 VSS.n1180 VSS.n1179 2.6005
R5014 VSS.n1184 VSS.n1183 2.6005
R5015 VSS.n1183 VSS.n1182 2.6005
R5016 VSS.n1187 VSS.n1186 2.6005
R5017 VSS.n1186 VSS.n1185 2.6005
R5018 VSS.n1190 VSS.n1189 2.6005
R5019 VSS.n1189 VSS.n1188 2.6005
R5020 VSS.n1193 VSS.n1192 2.6005
R5021 VSS.n1192 VSS.n1191 2.6005
R5022 VSS.n1196 VSS.n1195 2.6005
R5023 VSS.n1195 VSS.n1194 2.6005
R5024 VSS.n1199 VSS.n1198 2.6005
R5025 VSS.n1198 VSS.n1197 2.6005
R5026 VSS.n1171 VSS.n1170 2.6005
R5027 VSS.n1342 VSS.n1341 2.6005
R5028 VSS.n1345 VSS.n1344 2.6005
R5029 VSS.n1347 VSS.n1346 2.6005
R5030 VSS.n1350 VSS.n1349 2.6005
R5031 VSS.n1352 VSS.n1351 2.6005
R5032 VSS.n1355 VSS.n1354 2.6005
R5033 VSS.n1357 VSS.n1356 2.6005
R5034 VSS.n1360 VSS.n1359 2.6005
R5035 VSS.n1362 VSS.n1361 2.6005
R5036 VSS.n1365 VSS.n1364 2.6005
R5037 VSS.n1367 VSS.n1366 2.6005
R5038 VSS.n1371 VSS.n1370 2.6005
R5039 VSS.n1377 VSS.n1376 2.6005
R5040 VSS.n1376 VSS.n1375 2.6005
R5041 VSS.n1374 VSS.n1373 2.6005
R5042 VSS.n1373 VSS.n1372 2.6005
R5043 VSS.n4193 VSS.n4190 2.6005
R5044 VSS.n4158 VSS.n4150 2.6005
R5045 VSS.n4140 VSS.n4139 2.6005
R5046 VSS.n4143 VSS.n4142 2.6005
R5047 VSS.n4145 VSS.n4144 2.6005
R5048 VSS.n4159 VSS.n4158 2.6005
R5049 VSS.n4155 VSS 2.6005
R5050 VSS.n4155 VSS.n4154 2.6005
R5051 VSS.n4180 VSS.n4179 2.6005
R5052 VSS.n4184 VSS.n4183 2.6005
R5053 VSS.n4183 VSS.n4182 2.6005
R5054 VSS.n4194 VSS.n4193 2.6005
R5055 VSS.n4197 VSS.n4196 2.6005
R5056 VSS.n4201 VSS.n4200 2.6005
R5057 VSS.n4200 VSS.n4199 2.6005
R5058 VSS.n4229 VSS.n4228 2.6005
R5059 VSS.n4228 VSS.n4227 2.6005
R5060 VSS.n4226 VSS.n4225 2.6005
R5061 VSS.n4225 VSS.n4224 2.6005
R5062 VSS.n4223 VSS.n4222 2.6005
R5063 VSS.n4222 VSS.n4221 2.6005
R5064 VSS.n893 VSS.n892 2.6005
R5065 VSS.n892 VSS.n891 2.6005
R5066 VSS.n895 VSS.n894 2.6005
R5067 VSS.n897 VSS.n896 2.6005
R5068 VSS.n899 VSS.n898 2.6005
R5069 VSS.n902 VSS.n901 2.6005
R5070 VSS.n905 VSS.n904 2.6005
R5071 VSS.n907 VSS.n906 2.6005
R5072 VSS.n4255 VSS.n4254 2.6005
R5073 VSS.n4349 VSS.n4348 2.6005
R5074 VSS.n4345 VSS.n4344 2.6005
R5075 VSS.n4343 VSS.n4342 2.6005
R5076 VSS.n4340 VSS.n4339 2.6005
R5077 VSS.n4337 VSS.n4336 2.6005
R5078 VSS.n4270 VSS.n4269 2.6005
R5079 VSS.n4269 VSS.n4268 2.6005
R5080 VSS.n4267 VSS.n4266 2.6005
R5081 VSS.n4266 VSS.n4265 2.6005
R5082 VSS.n4264 VSS.n4263 2.6005
R5083 VSS.n4263 VSS.n4262 2.6005
R5084 VSS.n4261 VSS.n4260 2.6005
R5085 VSS.n4260 VSS.n4259 2.6005
R5086 VSS.n4258 VSS.n4257 2.6005
R5087 VSS.n4257 VSS.n4256 2.6005
R5088 VSS.n4254 VSS.n4253 2.6005
R5089 VSS.n4319 VSS.n4318 2.6005
R5090 VSS.n4315 VSS.n4314 2.6005
R5091 VSS.n4286 VSS.n4285 2.6005
R5092 VSS.n4285 VSS.n4284 2.6005
R5093 VSS.n4334 VSS.n4333 2.6005
R5094 VSS.n4330 VSS.n4329 2.6005
R5095 VSS.n4327 VSS.n4326 2.6005
R5096 VSS.n4324 VSS.n4323 2.6005
R5097 VSS.n4321 VSS.n4320 2.6005
R5098 VSS.n4278 VSS.n4277 2.6005
R5099 VSS.n4280 VSS.n4279 2.6005
R5100 VSS.n4283 VSS.n4282 2.6005
R5101 VSS.n4613 VSS.n4612 2.6005
R5102 VSS.n4612 VSS.n4611 2.6005
R5103 VSS.n4616 VSS.n4615 2.6005
R5104 VSS.n4615 VSS.n4614 2.6005
R5105 VSS.n4619 VSS.n4618 2.6005
R5106 VSS.n4618 VSS.n4617 2.6005
R5107 VSS.n4622 VSS.n4621 2.6005
R5108 VSS.n4621 VSS.n4620 2.6005
R5109 VSS.n4625 VSS.n4624 2.6005
R5110 VSS.n4624 VSS.n4623 2.6005
R5111 VSS.n4628 VSS.n4627 2.6005
R5112 VSS.n4627 VSS.n4626 2.6005
R5113 VSS.n4631 VSS.n4630 2.6005
R5114 VSS.n4630 VSS.n4629 2.6005
R5115 VSS.n4634 VSS.n4633 2.6005
R5116 VSS.n4633 VSS.n4632 2.6005
R5117 VSS.n4637 VSS.n4636 2.6005
R5118 VSS.n4636 VSS.n4635 2.6005
R5119 VSS.n4640 VSS.n4639 2.6005
R5120 VSS.n4639 VSS.n4638 2.6005
R5121 VSS.n4643 VSS.n4642 2.6005
R5122 VSS.n4642 VSS.n4641 2.6005
R5123 VSS.n4646 VSS.n4645 2.6005
R5124 VSS.n4645 VSS.n4644 2.6005
R5125 VSS.n4649 VSS.n4648 2.6005
R5126 VSS.n4648 VSS.n4647 2.6005
R5127 VSS.n4652 VSS.n4651 2.6005
R5128 VSS.n4651 VSS.n4650 2.6005
R5129 VSS.n116 VSS.n115 2.6005
R5130 VSS.n115 VSS.n114 2.6005
R5131 VSS.n113 VSS.n112 2.6005
R5132 VSS.n112 VSS.n111 2.6005
R5133 VSS.n123 VSS.n122 2.6005
R5134 VSS.n122 VSS.n121 2.6005
R5135 VSS.n198 VSS.n197 2.6005
R5136 VSS.n197 VSS.n196 2.6005
R5137 VSS.n201 VSS.n200 2.6005
R5138 VSS.n200 VSS.n199 2.6005
R5139 VSS.n204 VSS.n203 2.6005
R5140 VSS.n203 VSS.n202 2.6005
R5141 VSS.n194 VSS.n193 2.6005
R5142 VSS.n193 VSS.n192 2.6005
R5143 VSS.n208 VSS.n207 2.6005
R5144 VSS.n207 VSS.n206 2.6005
R5145 VSS.n211 VSS.n210 2.6005
R5146 VSS.n210 VSS.n209 2.6005
R5147 VSS.n214 VSS.n213 2.6005
R5148 VSS.n213 VSS.n212 2.6005
R5149 VSS.n218 VSS.n217 2.6005
R5150 VSS.n217 VSS.n216 2.6005
R5151 VSS.n191 VSS.n190 2.6005
R5152 VSS.n190 VSS.n189 2.6005
R5153 VSS.n187 VSS.n186 2.6005
R5154 VSS.n186 VSS.n185 2.6005
R5155 VSS.n167 VSS.n166 2.6005
R5156 VSS.n166 VSS.n165 2.6005
R5157 VSS.n164 VSS.n163 2.6005
R5158 VSS.n163 VSS.n162 2.6005
R5159 VSS.n251 VSS.n250 2.6005
R5160 VSS.n247 VSS.n246 2.6005
R5161 VSS.n120 VSS.n119 2.6005
R5162 VSS.n4391 VSS.n4390 2.6005
R5163 VSS.n4389 VSS.n4388 2.6005
R5164 VSS.n4385 VSS.n4384 2.6005
R5165 VSS.n101 VSS.n100 2.6005
R5166 VSS.n160 VSS.n159 2.6005
R5167 VSS.n159 VSS.n158 2.6005
R5168 VSS.n157 VSS.n156 2.6005
R5169 VSS.n156 VSS.n155 2.6005
R5170 VSS.n154 VSS.n153 2.6005
R5171 VSS.n153 VSS.n152 2.6005
R5172 VSS.n151 VSS.n150 2.6005
R5173 VSS.n150 VSS.n149 2.6005
R5174 VSS.n62 VSS.n61 2.6005
R5175 VSS.n61 VSS.n60 2.6005
R5176 VSS.n4610 VSS.n4609 2.6005
R5177 VSS.n4604 VSS.n4603 2.6005
R5178 VSS.n4599 VSS.n4598 2.6005
R5179 VSS.n4607 VSS.n4606 2.6005
R5180 VSS.n4596 VSS.n4595 2.6005
R5181 VSS.n4593 VSS.n4592 2.6005
R5182 VSS.n4588 VSS.n4587 2.6005
R5183 VSS.n4584 VSS.n4583 2.6005
R5184 VSS.n4580 VSS.n4579 2.6005
R5185 VSS.n4577 VSS.n4576 2.6005
R5186 VSS.n4655 VSS.n4654 2.6005
R5187 VSS.n4654 VSS.n4653 2.6005
R5188 VSS.n4659 VSS.n4658 2.6005
R5189 VSS.n4662 VSS.n4661 2.6005
R5190 VSS.n4665 VSS.n4664 2.6005
R5191 VSS.n4668 VSS.n4667 2.6005
R5192 VSS.n4672 VSS.n4671 2.6005
R5193 VSS.n4676 VSS.n4675 2.6005
R5194 VSS.n4679 VSS.n4678 2.6005
R5195 VSS.n54 VSS.n53 2.6005
R5196 VSS.n56 VSS.n55 2.6005
R5197 VSS.n4737 VSS.n4733 2.6005
R5198 VSS.n4695 VSS.n4693 2.6005
R5199 VSS.n4693 VSS.n4692 2.6005
R5200 VSS.n4699 VSS.n4696 2.6005
R5201 VSS.n4703 VSS.n4700 2.6005
R5202 VSS.n4714 VSS.n4713 2.6005
R5203 VSS.n4716 VSS 2.6005
R5204 VSS.n4716 VSS.n4715 2.6005
R5205 VSS.n4719 VSS.n4718 2.6005
R5206 VSS.n4718 VSS.n4717 2.6005
R5207 VSS.n4723 VSS.n4720 2.6005
R5208 VSS.n4727 VSS.n4725 2.6005
R5209 VSS.n4725 VSS.n4724 2.6005
R5210 VSS.n4731 VSS.n4728 2.6005
R5211 VSS.n4689 VSS.n4683 2.6005
R5212 VSS.n4683 VSS.n4682 2.6005
R5213 VSS.n4695 VSS.n4694 2.6005
R5214 VSS.n4699 VSS.n4698 2.6005
R5215 VSS.n4698 VSS.n4697 2.6005
R5216 VSS.n4703 VSS.n4702 2.6005
R5217 VSS.n4702 VSS.n4701 2.6005
R5218 VSS.n4713 VSS.n4712 2.6005
R5219 VSS.n4712 VSS.n4711 2.6005
R5220 VSS.n4710 VSS 2.6005
R5221 VSS.n4723 VSS.n4722 2.6005
R5222 VSS.n4722 VSS.n4721 2.6005
R5223 VSS.n4727 VSS.n4726 2.6005
R5224 VSS.n4731 VSS.n4730 2.6005
R5225 VSS.n4730 VSS.n4729 2.6005
R5226 VSS.n4737 VSS.n4736 2.6005
R5227 VSS.n4736 VSS.n4735 2.6005
R5228 VSS.n4689 VSS.n4688 2.6005
R5229 VSS.n5756 VSS 2.6005
R5230 VSS.n5757 VSS.n5756 2.6005
R5231 VSS VSS.n5752 2.6005
R5232 VSS.n5752 VSS.n5751 2.6005
R5233 VSS.n5824 VSS 2.6005
R5234 VSS.n5824 VSS.n5823 2.6005
R5235 VSS VSS.n5826 2.6005
R5236 VSS.n5826 VSS.n5825 2.6005
R5237 VSS.n1531 VSS.n1530 2.6005
R5238 VSS.n1530 VSS.n1529 2.6005
R5239 VSS.n1534 VSS.n1533 2.6005
R5240 VSS.n1533 VSS.n1532 2.6005
R5241 VSS.n3910 VSS.n3909 2.6005
R5242 VSS.n3912 VSS.n3911 2.6005
R5243 VSS.n3918 VSS.n3917 2.6005
R5244 VSS.n3917 VSS.n3916 2.6005
R5245 VSS.n3921 VSS.n3920 2.6005
R5246 VSS.n3920 VSS.n3919 2.6005
R5247 VSS.n3924 VSS.n3923 2.6005
R5248 VSS.n3923 VSS.n3922 2.6005
R5249 VSS.n3927 VSS.n3926 2.6005
R5250 VSS.n3926 VSS.n3925 2.6005
R5251 VSS.n3930 VSS.n3929 2.6005
R5252 VSS.n3929 VSS.n3928 2.6005
R5253 VSS.n3934 VSS.n3933 2.6005
R5254 VSS.n3933 VSS.n3932 2.6005
R5255 VSS.n3937 VSS.n3936 2.6005
R5256 VSS.n3936 VSS.n3935 2.6005
R5257 VSS.n3940 VSS.n3939 2.6005
R5258 VSS.n3939 VSS.n3938 2.6005
R5259 VSS.n3943 VSS.n3942 2.6005
R5260 VSS.n3942 VSS.n3941 2.6005
R5261 VSS.n3946 VSS.n3945 2.6005
R5262 VSS.n3945 VSS.n3944 2.6005
R5263 VSS.n3949 VSS.n3948 2.6005
R5264 VSS.n3948 VSS.n3947 2.6005
R5265 VSS.n3952 VSS.n3951 2.6005
R5266 VSS.n3951 VSS.n3950 2.6005
R5267 VSS.n3955 VSS.n3954 2.6005
R5268 VSS.n3954 VSS.n3953 2.6005
R5269 VSS.n3958 VSS.n3957 2.6005
R5270 VSS.n3957 VSS.n3956 2.6005
R5271 VSS.n3961 VSS.n3960 2.6005
R5272 VSS.n3960 VSS.n3959 2.6005
R5273 VSS.n3964 VSS.n3963 2.6005
R5274 VSS.n3963 VSS.n3962 2.6005
R5275 VSS.n3967 VSS.n3966 2.6005
R5276 VSS.n3966 VSS.n3965 2.6005
R5277 VSS.n3970 VSS.n3969 2.6005
R5278 VSS.n3969 VSS.n3968 2.6005
R5279 VSS.n3973 VSS.n3972 2.6005
R5280 VSS.n3972 VSS.n3971 2.6005
R5281 VSS.n3976 VSS.n3975 2.6005
R5282 VSS.n3975 VSS.n3974 2.6005
R5283 VSS.n4039 VSS.n4038 2.6005
R5284 VSS.n4046 VSS.n4045 2.6005
R5285 VSS.n4042 VSS.n4041 2.6005
R5286 VSS.n4037 VSS.n4036 2.6005
R5287 VSS.n4036 VSS.n4035 2.6005
R5288 VSS.n4034 VSS.n4033 2.6005
R5289 VSS.n4033 VSS.n4032 2.6005
R5290 VSS.n1528 VSS.n1527 2.6005
R5291 VSS.n1527 VSS.n1526 2.6005
R5292 VSS.n366 VSS.n365 2.6005
R5293 VSS.n368 VSS.n367 2.6005
R5294 VSS.n362 VSS.n361 2.6005
R5295 VSS.n1481 VSS.n1477 2.6005
R5296 VSS.n1477 VSS.n1476 2.6005
R5297 VSS.n1428 VSS.n1427 2.6005
R5298 VSS.n1427 VSS.n1426 2.6005
R5299 VSS.n1434 VSS.n1433 2.6005
R5300 VSS.n1433 VSS.n1432 2.6005
R5301 VSS.n1440 VSS.n1439 2.6005
R5302 VSS.n1439 VSS.n1438 2.6005
R5303 VSS.n1458 VSS.n1456 2.6005
R5304 VSS.n1458 VSS.n1457 2.6005
R5305 VSS VSS.n1460 2.6005
R5306 VSS.n1460 VSS.n1459 2.6005
R5307 VSS.n1472 VSS.n1471 2.6005
R5308 VSS.n1471 VSS.n1470 2.6005
R5309 VSS.n1500 VSS.n1499 2.6005
R5310 VSS.n1499 VSS.n1498 2.6005
R5311 VSS.n1494 VSS.n1493 2.6005
R5312 VSS.n1493 VSS.n1492 2.6005
R5313 VSS.n1488 VSS.n1487 2.6005
R5314 VSS.n1487 VSS.n1486 2.6005
R5315 VSS.n1421 VSS.n1420 2.6005
R5316 VSS VSS.n1468 2.6005
R5317 VSS.n1468 VSS.n1467 2.6005
R5318 VSS.n1475 VSS.n1474 2.6005
R5319 VSS.n1474 VSS.n1473 2.6005
R5320 VSS.n1497 VSS.n1496 2.6005
R5321 VSS.n1496 VSS.n1495 2.6005
R5322 VSS.n1491 VSS.n1490 2.6005
R5323 VSS.n1490 VSS.n1489 2.6005
R5324 VSS.n1485 VSS.n1484 2.6005
R5325 VSS.n1484 VSS.n1483 2.6005
R5326 VSS.n1480 VSS.n1479 2.6005
R5327 VSS.n1424 VSS.n1423 2.6005
R5328 VSS.n1423 VSS.n1422 2.6005
R5329 VSS.n1431 VSS.n1430 2.6005
R5330 VSS.n1430 VSS.n1429 2.6005
R5331 VSS.n1437 VSS.n1436 2.6005
R5332 VSS.n1436 VSS.n1435 2.6005
R5333 VSS.n1443 VSS.n1442 2.6005
R5334 VSS.n1442 VSS.n1441 2.6005
R5335 VSS.n1464 VSS.n1462 2.6005
R5336 VSS.n1464 VSS.n1463 2.6005
R5337 VSS.n1380 VSS.n1379 2.6005
R5338 VSS.n1379 VSS.n1378 2.6005
R5339 VSS.n1384 VSS.n1383 2.6005
R5340 VSS.n1383 VSS.n1382 2.6005
R5341 VSS.n1387 VSS.n1386 2.6005
R5342 VSS.n1386 VSS.n1385 2.6005
R5343 VSS.n1391 VSS.n1390 2.6005
R5344 VSS.n1390 VSS.n1389 2.6005
R5345 VSS.n4096 VSS.n4095 2.6005
R5346 VSS.n4095 VSS.n4094 2.6005
R5347 VSS.n4099 VSS.n4098 2.6005
R5348 VSS.n4098 VSS.n4097 2.6005
R5349 VSS.n4117 VSS.n4101 2.6005
R5350 VSS.n4101 VSS.n4100 2.6005
R5351 VSS.n4114 VSS.n4113 2.6005
R5352 VSS.n4104 VSS.n4103 2.6005
R5353 VSS.n4111 VSS.n4110 2.6005
R5354 VSS.n4110 VSS.n4109 2.6005
R5355 VSS.n4073 VSS.n4072 2.6005
R5356 VSS.n4072 VSS.n4071 2.6005
R5357 VSS.n4076 VSS.n4075 2.6005
R5358 VSS.n4075 VSS.n4074 2.6005
R5359 VSS.n4079 VSS.n4078 2.6005
R5360 VSS.n4078 VSS.n4077 2.6005
R5361 VSS.n4082 VSS.n4081 2.6005
R5362 VSS.n4081 VSS.n4080 2.6005
R5363 VSS.n4084 VSS.n4083 2.6005
R5364 VSS.n4085 VSS.n4084 2.6005
R5365 VSS.n4070 VSS.n4069 2.6005
R5366 VSS.n4069 VSS.n4068 2.6005
R5367 VSS.n1203 VSS.n1202 2.6005
R5368 VSS.n1202 VSS.n1201 2.6005
R5369 VSS.n1206 VSS.n1205 2.6005
R5370 VSS.n1205 VSS.n1204 2.6005
R5371 VSS.n1209 VSS.n1208 2.6005
R5372 VSS.n1208 VSS.n1207 2.6005
R5373 VSS.n1212 VSS.n1211 2.6005
R5374 VSS.n1211 VSS.n1210 2.6005
R5375 VSS.n1215 VSS.n1214 2.6005
R5376 VSS.n1214 VSS.n1213 2.6005
R5377 VSS.n1218 VSS.n1217 2.6005
R5378 VSS.n1217 VSS.n1216 2.6005
R5379 VSS.n1221 VSS.n1220 2.6005
R5380 VSS.n1220 VSS.n1219 2.6005
R5381 VSS.n1224 VSS.n1223 2.6005
R5382 VSS.n1223 VSS.n1222 2.6005
R5383 VSS.n1228 VSS.n1227 2.6005
R5384 VSS.n1227 VSS.n1226 2.6005
R5385 VSS.n1231 VSS.n1230 2.6005
R5386 VSS.n1230 VSS.n1229 2.6005
R5387 VSS.n1234 VSS.n1233 2.6005
R5388 VSS.n1233 VSS.n1232 2.6005
R5389 VSS.n1237 VSS.n1236 2.6005
R5390 VSS.n1236 VSS.n1235 2.6005
R5391 VSS.n1240 VSS.n1239 2.6005
R5392 VSS.n1239 VSS.n1238 2.6005
R5393 VSS.n1243 VSS.n1242 2.6005
R5394 VSS.n1242 VSS.n1241 2.6005
R5395 VSS.n1246 VSS.n1245 2.6005
R5396 VSS.n1245 VSS.n1244 2.6005
R5397 VSS.n1249 VSS.n1248 2.6005
R5398 VSS.n1248 VSS.n1247 2.6005
R5399 VSS.n1307 VSS.n1306 2.6005
R5400 VSS.n1304 VSS.n1303 2.6005
R5401 VSS.n1301 VSS.n1300 2.6005
R5402 VSS.n4241 VSS.n4240 2.6005
R5403 VSS.n4237 VSS.n4236 2.6005
R5404 VSS.n4234 VSS.n4233 2.6005
R5405 VSS.n4232 VSS.n4231 2.6005
R5406 VSS.n1283 VSS.n1282 2.6005
R5407 VSS.n1280 VSS.n1279 2.6005
R5408 VSS.n1277 VSS.n1276 2.6005
R5409 VSS.n1274 VSS.n1273 2.6005
R5410 VSS.n1271 VSS.n1270 2.6005
R5411 VSS.n1268 VSS.n1267 2.6005
R5412 VSS.n1265 VSS.n1264 2.6005
R5413 VSS.n1262 VSS.n1261 2.6005
R5414 VSS.n1259 VSS.n1258 2.6005
R5415 VSS.n1257 VSS.n1256 2.6005
R5416 VSS.n1251 VSS.n1250 2.6005
R5417 VSS.n1250 VSS.t668 2.6005
R5418 VSS.n1254 VSS.n1253 2.6005
R5419 VSS.n1253 VSS.n1252 2.6005
R5420 VSS.n1284 VSS.n974 2.6005
R5421 VSS.n1290 VSS.n1289 2.6005
R5422 VSS.n1297 VSS.n1296 2.6005
R5423 VSS.n1296 VSS.n1295 2.6005
R5424 VSS.n1293 VSS.n1292 2.6005
R5425 VSS.n1292 VSS.n1291 2.6005
R5426 VSS.n4251 VSS.n4250 2.6005
R5427 VSS.n4250 VSS.n4249 2.6005
R5428 VSS.n4247 VSS.n4246 2.6005
R5429 VSS.n4246 VSS.n4245 2.6005
R5430 VSS.n4244 VSS.n4243 2.6005
R5431 VSS.n4243 VSS.n4242 2.6005
R5432 VSS.n1288 VSS.n1287 2.6005
R5433 VSS.n38 VSS.n37 2.6005
R5434 VSS.n41 VSS.n40 2.6005
R5435 VSS.n44 VSS.n43 2.6005
R5436 VSS.n46 VSS.n45 2.6005
R5437 VSS.n51 VSS.n50 2.6005
R5438 VSS.n4574 VSS.n4573 2.6005
R5439 VSS.n4568 VSS.n4567 2.6005
R5440 VSS.n4563 VSS.n4562 2.6005
R5441 VSS.n4566 VSS.n4565 2.6005
R5442 VSS.n4559 VSS.n4558 2.6005
R5443 VSS.n4427 VSS.n4426 2.6005
R5444 VSS.n4424 VSS.n4423 2.6005
R5445 VSS.n4422 VSS.n4421 2.6005
R5446 VSS.n99 VSS.n98 2.6005
R5447 VSS.n976 VSS.n975 2.6005
R5448 VSS.n980 VSS.n979 2.6005
R5449 VSS.n4354 VSS.n4353 2.6005
R5450 VSS.n4418 VSS.n4417 2.6005
R5451 VSS.n4413 VSS.n4412 2.6005
R5452 VSS.n4351 VSS.n4350 2.6005
R5453 VSS.n4430 VSS.n4429 2.6005
R5454 VSS.n4429 VSS.n4428 2.6005
R5455 VSS.n4439 VSS.n4438 2.6005
R5456 VSS.n4438 VSS.n4437 2.6005
R5457 VSS.n4443 VSS.n4442 2.6005
R5458 VSS.n4442 VSS.n4441 2.6005
R5459 VSS.n4446 VSS.n4445 2.6005
R5460 VSS.n4445 VSS.n4444 2.6005
R5461 VSS.n4449 VSS.n4448 2.6005
R5462 VSS.n4448 VSS.n4447 2.6005
R5463 VSS.n4452 VSS.n4451 2.6005
R5464 VSS.n4451 VSS.n4450 2.6005
R5465 VSS.n4455 VSS.n4454 2.6005
R5466 VSS.n4454 VSS.n4453 2.6005
R5467 VSS.n4458 VSS.n4457 2.6005
R5468 VSS.n4457 VSS.n4456 2.6005
R5469 VSS.n4461 VSS.n4460 2.6005
R5470 VSS.n4460 VSS.n4459 2.6005
R5471 VSS.n4464 VSS.n4463 2.6005
R5472 VSS.n4463 VSS.n4462 2.6005
R5473 VSS.n4467 VSS.n4466 2.6005
R5474 VSS.n4466 VSS.n4465 2.6005
R5475 VSS.n4471 VSS.n4470 2.6005
R5476 VSS.n4470 VSS.n4469 2.6005
R5477 VSS.n4474 VSS.n4473 2.6005
R5478 VSS.n4473 VSS.n4472 2.6005
R5479 VSS.n4477 VSS.n4476 2.6005
R5480 VSS.n4476 VSS.n4475 2.6005
R5481 VSS.n4480 VSS.n4479 2.6005
R5482 VSS.n4479 VSS.n4478 2.6005
R5483 VSS.n4483 VSS.n4482 2.6005
R5484 VSS.n4482 VSS.n4481 2.6005
R5485 VSS.n4486 VSS.n4485 2.6005
R5486 VSS.n4485 VSS.n4484 2.6005
R5487 VSS.n4499 VSS.n4498 2.6005
R5488 VSS.n4498 VSS.n4497 2.6005
R5489 VSS.n4496 VSS.n4495 2.6005
R5490 VSS.n4495 VSS.n4494 2.6005
R5491 VSS.n4492 VSS.n4491 2.6005
R5492 VSS.n4491 VSS.n4490 2.6005
R5493 VSS.n4489 VSS.n4488 2.6005
R5494 VSS.n4488 VSS.n4487 2.6005
R5495 VSS.n4557 VSS.n4556 2.6005
R5496 VSS.n4554 VSS.n4553 2.6005
R5497 VSS.n4553 VSS.n4552 2.6005
R5498 VSS.n4551 VSS.n4550 2.6005
R5499 VSS.n4550 VSS.n4549 2.6005
R5500 VSS.n4548 VSS.n4547 2.6005
R5501 VSS.n4547 VSS.n4546 2.6005
R5502 VSS.n4545 VSS.n4544 2.6005
R5503 VSS.n4544 VSS.n4543 2.6005
R5504 VSS.n4542 VSS.n4541 2.6005
R5505 VSS.n4541 VSS.n4540 2.6005
R5506 VSS.n4539 VSS.n4538 2.6005
R5507 VSS.n4538 VSS.n4537 2.6005
R5508 VSS.n4536 VSS.n4535 2.6005
R5509 VSS.n4535 VSS.n4534 2.6005
R5510 VSS.n4533 VSS.n4532 2.6005
R5511 VSS.n4532 VSS.n4531 2.6005
R5512 VSS.n4530 VSS.n4529 2.6005
R5513 VSS.n4529 VSS.n4528 2.6005
R5514 VSS.n4527 VSS.n4526 2.6005
R5515 VSS.n4526 VSS.n4525 2.6005
R5516 VSS.n4524 VSS.n4523 2.6005
R5517 VSS.n4523 VSS.n4522 2.6005
R5518 VSS.n4521 VSS.n4520 2.6005
R5519 VSS.n4520 VSS.n4519 2.6005
R5520 VSS.n4518 VSS.n4517 2.6005
R5521 VSS.n4517 VSS.n4516 2.6005
R5522 VSS.n4515 VSS.n4514 2.6005
R5523 VSS.n4514 VSS.n4513 2.6005
R5524 VSS.n4512 VSS.n4511 2.6005
R5525 VSS.n35 VSS.n34 2.6005
R5526 VSS.n4433 VSS.n4432 2.6005
R5527 VSS.n4432 VSS.n4431 2.6005
R5528 VSS.n4436 VSS.n4435 2.6005
R5529 VSS.n4435 VSS.n4434 2.6005
R5530 VSS.n983 VSS.n982 2.6005
R5531 VSS.n985 VSS.n984 2.6005
R5532 VSS.n988 VSS.n987 2.6005
R5533 VSS.n992 VSS.n991 2.6005
R5534 VSS.n6029 VSS.n6028 2.6005
R5535 VSS.n6028 VSS.n6027 2.6005
R5536 VSS.n6032 VSS.n6031 2.6005
R5537 VSS.n6031 VSS.n6030 2.6005
R5538 VSS.n6036 VSS.n6035 2.6005
R5539 VSS.n6035 VSS.n6034 2.6005
R5540 VSS.n6040 VSS.n6039 2.6005
R5541 VSS.n6039 VSS.n6038 2.6005
R5542 VSS.n6043 VSS.n6042 2.6005
R5543 VSS.n6042 VSS.n6041 2.6005
R5544 VSS.n6046 VSS.n6045 2.6005
R5545 VSS.n6045 VSS.n6044 2.6005
R5546 VSS.n6049 VSS.n6048 2.6005
R5547 VSS.n6048 VSS.n6047 2.6005
R5548 VSS.n6052 VSS.n6051 2.6005
R5549 VSS.n6051 VSS.n6050 2.6005
R5550 VSS.n6054 VSS.n6053 2.6005
R5551 VSS.n6055 VSS.n6054 2.6005
R5552 VSS.n8 VSS.n7 2.6005
R5553 VSS.n7 VSS.n6 2.6005
R5554 VSS.n11 VSS.n10 2.6005
R5555 VSS.n10 VSS.n9 2.6005
R5556 VSS.n14 VSS.n13 2.6005
R5557 VSS.n13 VSS.n12 2.6005
R5558 VSS.n16 VSS.n15 2.6005
R5559 VSS.n17 VSS.n16 2.6005
R5560 VSS.n5 VSS.n4 2.6005
R5561 VSS.n4 VSS.n3 2.6005
R5562 VSS.n995 VSS.n994 2.6005
R5563 VSS.n994 VSS.n993 2.6005
R5564 VSS.n998 VSS.n997 2.6005
R5565 VSS.n997 VSS.n996 2.6005
R5566 VSS.n1002 VSS.n1001 2.6005
R5567 VSS.n1001 VSS.n1000 2.6005
R5568 VSS.n1005 VSS.n1004 2.6005
R5569 VSS.n1004 VSS.n1003 2.6005
R5570 VSS.n1008 VSS.n1007 2.6005
R5571 VSS.n1007 VSS.n1006 2.6005
R5572 VSS.n1037 VSS.n1036 2.6005
R5573 VSS.n1036 VSS.n1035 2.6005
R5574 VSS.n1040 VSS.n1039 2.6005
R5575 VSS.n1039 VSS.n1038 2.6005
R5576 VSS.n1043 VSS.n1042 2.6005
R5577 VSS.n1042 VSS.n1041 2.6005
R5578 VSS.n1046 VSS.n1045 2.6005
R5579 VSS.n1045 VSS.n1044 2.6005
R5580 VSS.n1049 VSS.n1048 2.6005
R5581 VSS.n1048 VSS.n1047 2.6005
R5582 VSS.n1052 VSS.n1051 2.6005
R5583 VSS.n1051 VSS.n1050 2.6005
R5584 VSS.n1055 VSS.n1054 2.6005
R5585 VSS.n1054 VSS.n1053 2.6005
R5586 VSS.n1058 VSS.n1057 2.6005
R5587 VSS.n1057 VSS.n1056 2.6005
R5588 VSS.n1061 VSS.n1060 2.6005
R5589 VSS.n1060 VSS.n1059 2.6005
R5590 VSS.n1064 VSS.n1063 2.6005
R5591 VSS.n1063 VSS.n1062 2.6005
R5592 VSS.n1067 VSS.n1066 2.6005
R5593 VSS.n1066 VSS.n1065 2.6005
R5594 VSS.n1070 VSS.n1069 2.6005
R5595 VSS.n1069 VSS.n1068 2.6005
R5596 VSS.n1073 VSS.n1072 2.6005
R5597 VSS.n1072 VSS.n1071 2.6005
R5598 VSS.n1076 VSS.n1075 2.6005
R5599 VSS.n1075 VSS.n1074 2.6005
R5600 VSS.n1080 VSS.n1079 2.6005
R5601 VSS.n1079 VSS.n1078 2.6005
R5602 VSS.n1083 VSS.n1082 2.6005
R5603 VSS.n1082 VSS.n1081 2.6005
R5604 VSS.n1086 VSS.n1085 2.6005
R5605 VSS.n1085 VSS.n1084 2.6005
R5606 VSS.n1089 VSS.n1088 2.6005
R5607 VSS.n1088 VSS.n1087 2.6005
R5608 VSS.n1092 VSS.n1091 2.6005
R5609 VSS.n1091 VSS.n1090 2.6005
R5610 VSS.n1095 VSS.n1094 2.6005
R5611 VSS.n1094 VSS.n1093 2.6005
R5612 VSS.n1098 VSS.n1097 2.6005
R5613 VSS.n1097 VSS.n1096 2.6005
R5614 VSS.n1101 VSS.n1100 2.6005
R5615 VSS.n1100 VSS.n1099 2.6005
R5616 VSS.n1104 VSS.n1103 2.6005
R5617 VSS.n1103 VSS.n1102 2.6005
R5618 VSS.n1107 VSS.n1106 2.6005
R5619 VSS.n1106 VSS.n1105 2.6005
R5620 VSS.n1110 VSS.n1109 2.6005
R5621 VSS.n1109 VSS.n1108 2.6005
R5622 VSS.n1113 VSS.n1112 2.6005
R5623 VSS.n1112 VSS.n1111 2.6005
R5624 VSS.n1116 VSS.n1115 2.6005
R5625 VSS.n1115 VSS.n1114 2.6005
R5626 VSS.n1119 VSS.n1118 2.6005
R5627 VSS.n1118 VSS.n1117 2.6005
R5628 VSS.n1122 VSS.n1121 2.6005
R5629 VSS.n1121 VSS.n1120 2.6005
R5630 VSS.n1125 VSS.n1124 2.6005
R5631 VSS.n1124 VSS.n1123 2.6005
R5632 VSS.n1128 VSS.n1127 2.6005
R5633 VSS.n1127 VSS.n1126 2.6005
R5634 VSS.n1131 VSS.n1130 2.6005
R5635 VSS.n1130 VSS.n1129 2.6005
R5636 VSS.n1134 VSS.n1133 2.6005
R5637 VSS.n1133 VSS.n1132 2.6005
R5638 VSS.n1137 VSS.n1136 2.6005
R5639 VSS.n1136 VSS.n1135 2.6005
R5640 VSS.n1140 VSS.n1139 2.6005
R5641 VSS.n1139 VSS.n1138 2.6005
R5642 VSS.n1143 VSS.n1142 2.6005
R5643 VSS.n1142 VSS.n1141 2.6005
R5644 VSS.n1146 VSS.n1145 2.6005
R5645 VSS.n1145 VSS.n1144 2.6005
R5646 VSS.n1149 VSS.n1148 2.6005
R5647 VSS.n1148 VSS.n1147 2.6005
R5648 VSS.n1152 VSS.n1151 2.6005
R5649 VSS.n1151 VSS.n1150 2.6005
R5650 VSS.n1155 VSS.n1154 2.6005
R5651 VSS.n1154 VSS.n1153 2.6005
R5652 VSS.n1158 VSS.n1157 2.6005
R5653 VSS.n1157 VSS.n1156 2.6005
R5654 VSS.n1161 VSS.n1160 2.6005
R5655 VSS.n1160 VSS.n1159 2.6005
R5656 VSS.n1168 VSS.n1167 2.6005
R5657 VSS.n1164 VSS.n1163 2.6005
R5658 VSS.n1163 VSS.n1162 2.6005
R5659 VSS.n5954 VSS.n5953 2.6005
R5660 VSS.n5953 VSS.n5952 2.6005
R5661 VSS.n5957 VSS.n5956 2.6005
R5662 VSS.n5956 VSS.n5955 2.6005
R5663 VSS.n5960 VSS.n5959 2.6005
R5664 VSS.n5959 VSS.n5958 2.6005
R5665 VSS.n5963 VSS.n5962 2.6005
R5666 VSS.n5962 VSS.n5961 2.6005
R5667 VSS.n5966 VSS.n5965 2.6005
R5668 VSS.n5965 VSS.n5964 2.6005
R5669 VSS.n5969 VSS.n5968 2.6005
R5670 VSS.n5968 VSS.n5967 2.6005
R5671 VSS.n5973 VSS.n5972 2.6005
R5672 VSS.n5972 VSS.n5971 2.6005
R5673 VSS.n5976 VSS.n5975 2.6005
R5674 VSS.n5975 VSS.n5974 2.6005
R5675 VSS.n5979 VSS.n5978 2.6005
R5676 VSS.n5978 VSS.n5977 2.6005
R5677 VSS.n5982 VSS.n5981 2.6005
R5678 VSS.n5981 VSS.n5980 2.6005
R5679 VSS.n5985 VSS.n5984 2.6005
R5680 VSS.n5984 VSS.n5983 2.6005
R5681 VSS.n5988 VSS.n5987 2.6005
R5682 VSS.n5987 VSS.n5986 2.6005
R5683 VSS.n5991 VSS.n5990 2.6005
R5684 VSS.n5990 VSS.n5989 2.6005
R5685 VSS.n5994 VSS.n5993 2.6005
R5686 VSS.n5993 VSS.n5992 2.6005
R5687 VSS.n5997 VSS.n5996 2.6005
R5688 VSS.n5996 VSS.n5995 2.6005
R5689 VSS.n6000 VSS.n5999 2.6005
R5690 VSS.n5999 VSS.n5998 2.6005
R5691 VSS.n6003 VSS.n6002 2.6005
R5692 VSS.n6002 VSS.n6001 2.6005
R5693 VSS.n6006 VSS.n6005 2.6005
R5694 VSS.n6005 VSS.n6004 2.6005
R5695 VSS.n6009 VSS.n6008 2.6005
R5696 VSS.n6008 VSS.n6007 2.6005
R5697 VSS.n6012 VSS.n6011 2.6005
R5698 VSS.n6011 VSS.n6010 2.6005
R5699 VSS.n6015 VSS.n6014 2.6005
R5700 VSS.n6014 VSS.n6013 2.6005
R5701 VSS.n6019 VSS.n6018 2.6005
R5702 VSS.n6018 VSS.n6017 2.6005
R5703 VSS.n6022 VSS.n6021 2.6005
R5704 VSS.n6021 VSS.n6020 2.6005
R5705 VSS.n6025 VSS.n6024 2.6005
R5706 VSS.n6024 VSS.n6023 2.6005
R5707 VSS.n5605 VSS.n5604 2.6005
R5708 VSS.n5607 VSS.n5606 2.6005
R5709 VSS.n5609 VSS.n5608 2.6005
R5710 VSS.n5612 VSS.n5611 2.6005
R5711 VSS.n5615 VSS.n5614 2.6005
R5712 VSS.n5513 VSS.n5512 2.6005
R5713 VSS.n5419 VSS.n5418 2.6005
R5714 VSS.n5418 VSS.n5417 2.6005
R5715 VSS.n5416 VSS.n5415 2.6005
R5716 VSS.n5415 VSS.n5414 2.6005
R5717 VSS.n5413 VSS.n5412 2.6005
R5718 VSS.n5412 VSS.n5411 2.6005
R5719 VSS.n5409 VSS.n5408 2.6005
R5720 VSS.n5314 VSS.n5313 2.6005
R5721 VSS.n5045 VSS.n5044 2.6005
R5722 VSS.n5003 VSS.n5002 2.6005
R5723 VSS.n5002 VSS.n5001 2.6005
R5724 VSS.n5006 VSS.n5005 2.6005
R5725 VSS.n5005 VSS.n5004 2.6005
R5726 VSS.n5010 VSS.n5009 2.6005
R5727 VSS.n5009 VSS.n5008 2.6005
R5728 VSS.n5013 VSS.n5012 2.6005
R5729 VSS.n5012 VSS.n5011 2.6005
R5730 VSS.n5016 VSS.n5015 2.6005
R5731 VSS.n5015 VSS.n5014 2.6005
R5732 VSS.n5019 VSS.n5018 2.6005
R5733 VSS.n5018 VSS.n5017 2.6005
R5734 VSS.n5022 VSS.n5021 2.6005
R5735 VSS.n5021 VSS.n5020 2.6005
R5736 VSS.n5025 VSS.n5024 2.6005
R5737 VSS.n5024 VSS.n5023 2.6005
R5738 VSS.n5028 VSS.n5027 2.6005
R5739 VSS.n5027 VSS.n5026 2.6005
R5740 VSS.n5031 VSS.n5030 2.6005
R5741 VSS.n5030 VSS.n5029 2.6005
R5742 VSS.n5034 VSS.n5033 2.6005
R5743 VSS.n5033 VSS.n5032 2.6005
R5744 VSS.n5037 VSS.n5036 2.6005
R5745 VSS.n5036 VSS.n5035 2.6005
R5746 VSS.n5040 VSS.n5039 2.6005
R5747 VSS.n5039 VSS.n5038 2.6005
R5748 VSS.n5043 VSS.n5042 2.6005
R5749 VSS.n5042 VSS.n5041 2.6005
R5750 VSS.n5262 VSS.n5261 2.6005
R5751 VSS.n5632 VSS.n5631 2.6005
R5752 VSS.n5312 VSS.n5311 2.6005
R5753 VSS.n5290 VSS.n5289 2.6005
R5754 VSS.n5286 VSS.n5285 2.6005
R5755 VSS.n5622 VSS.n5621 2.6005
R5756 VSS.n5624 VSS.n5623 2.6005
R5757 VSS.n5627 VSS.n5626 2.6005
R5758 VSS.n5630 VSS.n5629 2.6005
R5759 VSS.n5619 VSS.n5618 2.6005
R5760 VSS.n4765 VSS.n4764 2.6005
R5761 VSS.n5650 VSS.n5649 2.6005
R5762 VSS.n5652 VSS.n5651 2.6005
R5763 VSS.n5655 VSS.n5654 2.6005
R5764 VSS.n5660 VSS.n5659 2.6005
R5765 VSS.n5646 VSS.n5645 2.6005
R5766 VSS.n5643 VSS.n5642 2.6005
R5767 VSS.n5641 VSS.n5640 2.6005
R5768 VSS.n5638 VSS.n5637 2.6005
R5769 VSS.n5636 VSS.n5635 2.6005
R5770 VSS.n5250 VSS.n5249 2.6005
R5771 VSS.n5252 VSS.n5251 2.6005
R5772 VSS.n5246 VSS.n5245 2.6005
R5773 VSS.n5244 VSS.n5243 2.6005
R5774 VSS.n5063 VSS.n5062 2.6005
R5775 VSS.n5065 VSS.n5064 2.6005
R5776 VSS.n5052 VSS.n5051 2.6005
R5777 VSS.n5068 VSS.n5067 2.6005
R5778 VSS.n5071 VSS.n5070 2.6005
R5779 VSS.n5074 VSS.n5073 2.6005
R5780 VSS.n5078 VSS.n5077 2.6005
R5781 VSS.n5097 VSS.n5096 2.6005
R5782 VSS.n5101 VSS.n5100 2.6005
R5783 VSS.n5103 VSS.n5102 2.6005
R5784 VSS.n5122 VSS.n5121 2.6005
R5785 VSS.n5125 VSS.n5124 2.6005
R5786 VSS.n5459 VSS.n5458 2.6005
R5787 VSS.n5128 VSS.n5127 2.6005
R5788 VSS.n5132 VSS.n5131 2.6005
R5789 VSS.n5131 VSS.n5130 2.6005
R5790 VSS.n5135 VSS.n5134 2.6005
R5791 VSS.n5134 VSS.n5133 2.6005
R5792 VSS.n5138 VSS.n5137 2.6005
R5793 VSS.n5137 VSS.n5136 2.6005
R5794 VSS.n5141 VSS.n5140 2.6005
R5795 VSS.n5140 VSS.n5139 2.6005
R5796 VSS.n5144 VSS.n5143 2.6005
R5797 VSS.n5143 VSS.n5142 2.6005
R5798 VSS.n5157 VSS.n5156 2.6005
R5799 VSS.n5156 VSS.n5155 2.6005
R5800 VSS.n5160 VSS.n5159 2.6005
R5801 VSS.n5159 VSS.n5158 2.6005
R5802 VSS.n5180 VSS.n5179 2.6005
R5803 VSS.n5179 VSS.n5178 2.6005
R5804 VSS.n5184 VSS.n5183 2.6005
R5805 VSS.n5183 VSS.n5182 2.6005
R5806 VSS.n5207 VSS.n5206 2.6005
R5807 VSS.n5206 VSS.n5205 2.6005
R5808 VSS.n5211 VSS.n5210 2.6005
R5809 VSS.n5210 VSS.n5209 2.6005
R5810 VSS.n5214 VSS.n5213 2.6005
R5811 VSS.n5213 VSS.n5212 2.6005
R5812 VSS.n5217 VSS.n5216 2.6005
R5813 VSS.n5216 VSS.n5215 2.6005
R5814 VSS.n4786 VSS.n4785 2.6005
R5815 VSS.n4785 VSS.n4784 2.6005
R5816 VSS.n5221 VSS.n5220 2.6005
R5817 VSS.n5220 VSS.n5219 2.6005
R5818 VSS.n5224 VSS.n5223 2.6005
R5819 VSS.n5223 VSS.n5222 2.6005
R5820 VSS.n5227 VSS.n5226 2.6005
R5821 VSS.n5226 VSS.n5225 2.6005
R5822 VSS.n5231 VSS.n5230 2.6005
R5823 VSS.n5230 VSS.n5229 2.6005
R5824 VSS.n4755 VSS.n4754 2.6005
R5825 VSS.n4754 VSS.n4753 2.6005
R5826 VSS.n4758 VSS.n4757 2.6005
R5827 VSS.n4757 VSS.n4756 2.6005
R5828 VSS.n5422 VSS.n5421 2.6005
R5829 VSS.n5421 VSS.n5420 2.6005
R5830 VSS.n5426 VSS.n5425 2.6005
R5831 VSS.n5425 VSS.n5424 2.6005
R5832 VSS.n5405 VSS.n5404 2.6005
R5833 VSS.n5430 VSS.n5429 2.6005
R5834 VSS.n5429 VSS.n5428 2.6005
R5835 VSS.n5433 VSS.n5432 2.6005
R5836 VSS.n5432 VSS.n5431 2.6005
R5837 VSS.n5436 VSS.n5435 2.6005
R5838 VSS.n5435 VSS.n5434 2.6005
R5839 VSS.n5439 VSS.n5438 2.6005
R5840 VSS.n5438 VSS.n5437 2.6005
R5841 VSS.n5442 VSS.n5441 2.6005
R5842 VSS.n5441 VSS.n5440 2.6005
R5843 VSS.n5403 VSS.n5402 2.6005
R5844 VSS.n5446 VSS.n5445 2.6005
R5845 VSS.n5445 VSS.n5444 2.6005
R5846 VSS.n5449 VSS.n5448 2.6005
R5847 VSS.n5448 VSS.n5447 2.6005
R5848 VSS.n5452 VSS.n5451 2.6005
R5849 VSS.n5451 VSS.n5450 2.6005
R5850 VSS.n5455 VSS.n5454 2.6005
R5851 VSS.n5454 VSS.n5453 2.6005
R5852 VSS.n5457 VSS.n5456 2.6005
R5853 VSS.n5537 VSS.n5536 2.6005
R5854 VSS.n5536 VSS.n5535 2.6005
R5855 VSS.n5534 VSS.n5533 2.6005
R5856 VSS.n5533 VSS.n5532 2.6005
R5857 VSS.n5526 VSS.n5525 2.6005
R5858 VSS.n5525 VSS.n5524 2.6005
R5859 VSS.n5523 VSS.n5522 2.6005
R5860 VSS.n5522 VSS.n5521 2.6005
R5861 VSS.n5520 VSS.n5519 2.6005
R5862 VSS.n5519 VSS.n5518 2.6005
R5863 VSS.n5517 VSS.n5516 2.6005
R5864 VSS.n5516 VSS.n5515 2.6005
R5865 VSS.n5463 VSS.n5462 2.6005
R5866 VSS.n5462 VSS.n5461 2.6005
R5867 VSS.n5478 VSS.n5477 2.6005
R5868 VSS.n5477 VSS.n5476 2.6005
R5869 VSS.n5481 VSS.n5480 2.6005
R5870 VSS.n5480 VSS.n5479 2.6005
R5871 VSS.n5484 VSS.n5483 2.6005
R5872 VSS.n5483 VSS.n5482 2.6005
R5873 VSS.n5487 VSS.n5486 2.6005
R5874 VSS.n5486 VSS.n5485 2.6005
R5875 VSS.n5490 VSS.n5489 2.6005
R5876 VSS.n5489 VSS.n5488 2.6005
R5877 VSS.n5493 VSS.n5492 2.6005
R5878 VSS.n5492 VSS.n5491 2.6005
R5879 VSS.n5496 VSS.n5495 2.6005
R5880 VSS.n5495 VSS.n5494 2.6005
R5881 VSS.n5499 VSS.n5498 2.6005
R5882 VSS.n5498 VSS.n5497 2.6005
R5883 VSS.n5502 VSS.n5501 2.6005
R5884 VSS.n5501 VSS.n5500 2.6005
R5885 VSS.n5505 VSS.n5504 2.6005
R5886 VSS.n5504 VSS.n5503 2.6005
R5887 VSS.n5508 VSS.n5507 2.6005
R5888 VSS.n5507 VSS.n5506 2.6005
R5889 VSS.n5511 VSS.n5510 2.6005
R5890 VSS.n5510 VSS.n5509 2.6005
R5891 VSS.n5475 VSS.n5474 2.6005
R5892 VSS.n5474 VSS.n5473 2.6005
R5893 VSS.n5599 VSS.n5598 2.6005
R5894 VSS.n5598 VSS.n5597 2.6005
R5895 VSS.n5596 VSS.n5595 2.6005
R5896 VSS.n5595 VSS.n5594 2.6005
R5897 VSS.n5593 VSS.n5592 2.6005
R5898 VSS.n5592 VSS.n5591 2.6005
R5899 VSS.n5589 VSS.n5588 2.6005
R5900 VSS.n5588 VSS.n5587 2.6005
R5901 VSS.n5586 VSS.n5585 2.6005
R5902 VSS.n5585 VSS.n5584 2.6005
R5903 VSS.n5583 VSS.n5582 2.6005
R5904 VSS.n5582 VSS.n5581 2.6005
R5905 VSS.n5580 VSS.n5579 2.6005
R5906 VSS.n5579 VSS.n5578 2.6005
R5907 VSS.n5577 VSS.n5576 2.6005
R5908 VSS.n5576 VSS.n5575 2.6005
R5909 VSS.n5573 VSS.n5572 2.6005
R5910 VSS.n5572 VSS.n5571 2.6005
R5911 VSS.n5569 VSS.n5568 2.6005
R5912 VSS.n5568 VSS.t276 2.6005
R5913 VSS.n5567 VSS.n5566 2.6005
R5914 VSS.n5566 VSS.n5565 2.6005
R5915 VSS.n5564 VSS.n5563 2.6005
R5916 VSS.n5563 VSS.n5562 2.6005
R5917 VSS.n5561 VSS.n5560 2.6005
R5918 VSS.n5560 VSS.n5559 2.6005
R5919 VSS.n5558 VSS.n5557 2.6005
R5920 VSS.n5557 VSS.n5556 2.6005
R5921 VSS.n5554 VSS.n5553 2.6005
R5922 VSS.n5553 VSS.n5552 2.6005
R5923 VSS.n5551 VSS.n5550 2.6005
R5924 VSS.n5550 VSS.n5549 2.6005
R5925 VSS.n5548 VSS.n5547 2.6005
R5926 VSS.n5547 VSS.n5546 2.6005
R5927 VSS.n5545 VSS.n5544 2.6005
R5928 VSS.n5544 VSS.n5543 2.6005
R5929 VSS.n5542 VSS.n5541 2.6005
R5930 VSS.n5541 VSS.n5540 2.6005
R5931 VSS.n5401 VSS.n5400 2.6005
R5932 VSS.n5400 VSS.n5399 2.6005
R5933 VSS.n5398 VSS.n5397 2.6005
R5934 VSS.n5397 VSS.n5396 2.6005
R5935 VSS.n5395 VSS.n5394 2.6005
R5936 VSS.n5394 VSS.n5393 2.6005
R5937 VSS.n5392 VSS.n5391 2.6005
R5938 VSS.n5391 VSS.n5390 2.6005
R5939 VSS.n5389 VSS.n5388 2.6005
R5940 VSS.n5388 VSS.n5387 2.6005
R5941 VSS.n5386 VSS.n5385 2.6005
R5942 VSS.n5385 VSS.n5384 2.6005
R5943 VSS.n5383 VSS.n5382 2.6005
R5944 VSS.n5382 VSS.n5381 2.6005
R5945 VSS.n5380 VSS.n5379 2.6005
R5946 VSS.n5379 VSS.n5378 2.6005
R5947 VSS.n5377 VSS.n5376 2.6005
R5948 VSS.n5376 VSS.n5375 2.6005
R5949 VSS.n5374 VSS.n5373 2.6005
R5950 VSS.n5373 VSS.n5372 2.6005
R5951 VSS.n5371 VSS.n5370 2.6005
R5952 VSS.n5370 VSS.n5369 2.6005
R5953 VSS.n5368 VSS.n5367 2.6005
R5954 VSS.n5367 VSS.n5366 2.6005
R5955 VSS.n5365 VSS.n5364 2.6005
R5956 VSS.n5364 VSS.n5363 2.6005
R5957 VSS.n5362 VSS.n5361 2.6005
R5958 VSS.n5361 VSS.n5360 2.6005
R5959 VSS.n5359 VSS.n5358 2.6005
R5960 VSS.n5358 VSS.n5357 2.6005
R5961 VSS.n5356 VSS.n5355 2.6005
R5962 VSS.n5355 VSS.n5354 2.6005
R5963 VSS.n5353 VSS.n5352 2.6005
R5964 VSS.n5352 VSS.n5351 2.6005
R5965 VSS.n5350 VSS.n5349 2.6005
R5966 VSS.n5349 VSS.n5348 2.6005
R5967 VSS.n5347 VSS.n5346 2.6005
R5968 VSS.n5346 VSS.n5345 2.6005
R5969 VSS.n5344 VSS.n5343 2.6005
R5970 VSS.n5343 VSS.n5342 2.6005
R5971 VSS.n5341 VSS.n5340 2.6005
R5972 VSS.n5340 VSS.n5339 2.6005
R5973 VSS.n5663 VSS.n5662 2.6005
R5974 VSS.n5662 VSS.n5661 2.6005
R5975 VSS.n5670 VSS.n5669 2.6005
R5976 VSS.n5669 VSS.n5668 2.6005
R5977 VSS.n5673 VSS.n5672 2.6005
R5978 VSS.n5672 VSS.n5671 2.6005
R5979 VSS.n5676 VSS.n5675 2.6005
R5980 VSS.n5675 VSS.n5674 2.6005
R5981 VSS.n5679 VSS.n5678 2.6005
R5982 VSS.n5678 VSS.n5677 2.6005
R5983 VSS.n5682 VSS.n5681 2.6005
R5984 VSS.n5681 VSS.n5680 2.6005
R5985 VSS.n5685 VSS.n5684 2.6005
R5986 VSS.n5684 VSS.n5683 2.6005
R5987 VSS.n5688 VSS.n5687 2.6005
R5988 VSS.n5687 VSS.n5686 2.6005
R5989 VSS.n5691 VSS.n5690 2.6005
R5990 VSS.n5690 VSS.n5689 2.6005
R5991 VSS.n5695 VSS.n5694 2.6005
R5992 VSS.n5694 VSS.n5693 2.6005
R5993 VSS.n5698 VSS.n5697 2.6005
R5994 VSS.n5697 VSS.n5696 2.6005
R5995 VSS.n5701 VSS.n5700 2.6005
R5996 VSS.n5700 VSS.n5699 2.6005
R5997 VSS.n5704 VSS.n5703 2.6005
R5998 VSS.n5703 VSS.n5702 2.6005
R5999 VSS.n5707 VSS.n5706 2.6005
R6000 VSS.n5706 VSS.n5705 2.6005
R6001 VSS.n5710 VSS.n5709 2.6005
R6002 VSS.n5709 VSS.n5708 2.6005
R6003 VSS.n5713 VSS.n5712 2.6005
R6004 VSS.n5712 VSS.n5711 2.6005
R6005 VSS.n5715 VSS.n5714 2.6005
R6006 VSS.n5716 VSS.n5715 2.6005
R6007 VSS.n5901 VSS.n5900 2.6005
R6008 VSS.n5900 VSS.n5899 2.6005
R6009 VSS.n5904 VSS.n5903 2.6005
R6010 VSS.n5903 VSS.n5902 2.6005
R6011 VSS.n5907 VSS.n5906 2.6005
R6012 VSS.n5906 VSS.n5905 2.6005
R6013 VSS.n5910 VSS.n5909 2.6005
R6014 VSS.n5909 VSS.n5908 2.6005
R6015 VSS.n5913 VSS.n5912 2.6005
R6016 VSS.n5912 VSS.n5911 2.6005
R6017 VSS.n5916 VSS.n5915 2.6005
R6018 VSS.n5915 VSS.n5914 2.6005
R6019 VSS.n5919 VSS.n5918 2.6005
R6020 VSS.n5918 VSS.n5917 2.6005
R6021 VSS.n5922 VSS.n5921 2.6005
R6022 VSS.n5921 VSS.n5920 2.6005
R6023 VSS.n5925 VSS.n5924 2.6005
R6024 VSS.n5924 VSS.n5923 2.6005
R6025 VSS.n5928 VSS.n5927 2.6005
R6026 VSS.n5927 VSS.n5926 2.6005
R6027 VSS.n5931 VSS.n5930 2.6005
R6028 VSS.n5930 VSS.n5929 2.6005
R6029 VSS.n5934 VSS.n5933 2.6005
R6030 VSS.n5933 VSS.n5932 2.6005
R6031 VSS.n5937 VSS.n5936 2.6005
R6032 VSS.n5936 VSS.n5935 2.6005
R6033 VSS.n5940 VSS.n5939 2.6005
R6034 VSS.n5939 VSS.n5938 2.6005
R6035 VSS.n5943 VSS.n5942 2.6005
R6036 VSS.n5942 VSS.n5941 2.6005
R6037 VSS.n5947 VSS.n5946 2.6005
R6038 VSS.n5946 VSS.n5945 2.6005
R6039 VSS.n5950 VSS.n5949 2.6005
R6040 VSS.n5949 VSS.n5948 2.6005
R6041 VSS.n4752 VSS.n4751 2.6005
R6042 VSS.n4749 VSS.n4748 2.6005
R6043 VSS.n4740 VSS.n4739 2.6005
R6044 VSS.n5898 VSS.n5897 2.6005
R6045 VSS VSS.n5812 2.6005
R6046 VSS.n5812 VSS.t642 2.6005
R6047 VSS.n5770 VSS 2.6005
R6048 VSS.n5770 VSS.n5769 2.6005
R6049 VSS.n1019 VSS.n1018 2.6005
R6050 VSS.n1022 VSS.n1021 2.6005
R6051 VSS.n1016 VSS.n1015 2.6005
R6052 VSS.n4055 VSS.n4054 2.59998
R6053 VSS.n1566 VSS.n1565 2.53192
R6054 VSS.n1261 VSS.n1260 2.48961
R6055 VSS.n1264 VSS.n1263 2.48961
R6056 VSS.n1267 VSS.n1266 2.48961
R6057 VSS.n1270 VSS.n1269 2.48961
R6058 VSS.n1273 VSS.n1272 2.48961
R6059 VSS.n1276 VSS.n1275 2.48961
R6060 VSS.n1279 VSS.n1278 2.48961
R6061 VSS.n471 VSS.n470 2.41686
R6062 VSS.n5789 VSS.n5788 2.36862
R6063 VSS.n5884 VSS.n5883 2.34081
R6064 VSS.n1646 VSS.n1554 2.3405
R6065 VSS.n1647 VSS.n1544 2.33208
R6066 VSS.n1566 VSS.n1561 2.33079
R6067 VSS.n5781 VSS.n21 2.30179
R6068 VSS.n987 VSS.n986 2.29396
R6069 VSS.n5788 VSS.n5787 2.29248
R6070 VSS.n2802 VSS.n2801 2.28632
R6071 VSS.n5328 VSS.n5327 2.28399
R6072 VSS.n5331 VSS.n5330 2.28399
R6073 VSS.n558 VSS.n557 2.28399
R6074 VSS.n561 VSS.n560 2.28399
R6075 VSS.n677 VSS.n676 2.28399
R6076 VSS.n680 VSS.n679 2.28399
R6077 VSS.n5654 VSS.n5653 2.28399
R6078 VSS.n5626 VSS.n5625 2.28399
R6079 VSS.n5614 VSS.n5613 2.28399
R6080 VSS.n5611 VSS.n5610 2.28399
R6081 VSS.n4739 VSS.n4738 2.28399
R6082 VSS.n5858 VSS 2.28174
R6083 VSS.n2722 VSS.n2212 2.2791
R6084 VSS.n2580 VSS.n2579 2.27836
R6085 VSS.n2193 VSS.n2192 2.27834
R6086 VSS.n2879 VSS.n1995 2.27413
R6087 VSS.n2789 VSS.n2094 2.27187
R6088 VSS.n2656 VSS.n2320 2.26934
R6089 VSS.n2663 VSS.n2308 2.25712
R6090 VSS.n4371 VSS.n4370 2.25676
R6091 VSS.n5275 VSS.n5274 2.25635
R6092 VSS.n2560 VSS.n2413 2.25613
R6093 VSS.n874 VSS.n870 2.25575
R6094 VSS.n1754 VSS.t57 2.25428
R6095 VSS.n1755 VSS.t37 2.25428
R6096 VSS.n1756 VSS.t109 2.25428
R6097 VSS.n1757 VSS.t118 2.25428
R6098 VSS.n1758 VSS.t35 2.25428
R6099 VSS.n1759 VSS.t44 2.25428
R6100 VSS.n1760 VSS.t22 2.25428
R6101 VSS.n1761 VSS.t102 2.25428
R6102 VSS.n1762 VSS.t105 2.25428
R6103 VSS.n1763 VSS.t83 2.25428
R6104 VSS.n1764 VSS.t28 2.25428
R6105 VSS.n2458 VSS.t112 2.25428
R6106 VSS.n2459 VSS.t94 2.25428
R6107 VSS.n2460 VSS.t30 2.25428
R6108 VSS.n2461 VSS.t39 2.25428
R6109 VSS.n2462 VSS.t90 2.25428
R6110 VSS.n2463 VSS.t101 2.25428
R6111 VSS.n2464 VSS.t75 2.25428
R6112 VSS.n2465 VSS.t21 2.25428
R6113 VSS.n2466 VSS.t24 2.25428
R6114 VSS.n2467 VSS.t128 2.25428
R6115 VSS.n2468 VSS.t82 2.25428
R6116 VSS.n2372 VSS.t33 2.25428
R6117 VSS.n2373 VSS.t10 2.25428
R6118 VSS.n2374 VSS.t87 2.25428
R6119 VSS.n2375 VSS.t99 2.25428
R6120 VSS.n2376 VSS.t7 2.25428
R6121 VSS.n2377 VSS.t16 2.25428
R6122 VSS.n2378 VSS.t123 2.25428
R6123 VSS.n2379 VSS.t77 2.25428
R6124 VSS.n2380 VSS.t79 2.25428
R6125 VSS.n2381 VSS.t54 2.25428
R6126 VSS.n2382 VSS.t0 2.25428
R6127 VSS.n2255 VSS.t65 2.25428
R6128 VSS.n2256 VSS.t43 2.25428
R6129 VSS.n2257 VSS.t117 2.25428
R6130 VSS.n2258 VSS.t121 2.25428
R6131 VSS.n2259 VSS.t41 2.25428
R6132 VSS.n2260 VSS.t48 2.25428
R6133 VSS.n2261 VSS.t27 2.25428
R6134 VSS.n2262 VSS.t107 2.25428
R6135 VSS.n2263 VSS.t108 2.25428
R6136 VSS.n2264 VSS.t91 2.25428
R6137 VSS.n2265 VSS.t34 2.25428
R6138 VSS.n2148 VSS.t17 2.25428
R6139 VSS.n2149 VSS.t124 2.25428
R6140 VSS.n2150 VSS.t73 2.25428
R6141 VSS.n2151 VSS.t80 2.25428
R6142 VSS.n2152 VSS.t122 2.25428
R6143 VSS.n2153 VSS.t1 2.25428
R6144 VSS.n2154 VSS.t114 2.25428
R6145 VSS.n2155 VSS.t60 2.25428
R6146 VSS.n2156 VSS.t62 2.25428
R6147 VSS.n2157 VSS.t40 2.25428
R6148 VSS.n2158 VSS.t120 2.25428
R6149 VSS.n2051 VSS.t97 2.25428
R6150 VSS.n2052 VSS.t72 2.25428
R6151 VSS.n2053 VSS.t9 2.25428
R6152 VSS.n2054 VSS.t18 2.25428
R6153 VSS.n2055 VSS.t69 2.25428
R6154 VSS.n2056 VSS.t78 2.25428
R6155 VSS.n2057 VSS.t53 2.25428
R6156 VSS.n2058 VSS.t130 2.25428
R6157 VSS.n2059 VSS.t2 2.25428
R6158 VSS.n2060 VSS.t116 2.25428
R6159 VSS.n2061 VSS.t61 2.25428
R6160 VSS.n1981 VSS.t95 2.25428
R6161 VSS.n1982 VSS.t70 2.25428
R6162 VSS.n1983 VSS.t6 2.25428
R6163 VSS.n1984 VSS.t14 2.25428
R6164 VSS.n1985 VSS.t66 2.25428
R6165 VSS.n1986 VSS.t76 2.25428
R6166 VSS.n1987 VSS.t51 2.25428
R6167 VSS.n1988 VSS.t127 2.25428
R6168 VSS.n1989 VSS.t131 2.25428
R6169 VSS.n1990 VSS.t113 2.25428
R6170 VSS.n1991 VSS.t58 2.25428
R6171 VSS.n1826 VSS.t93 2.25428
R6172 VSS.n1827 VSS.t68 2.25428
R6173 VSS.n1828 VSS.t5 2.25428
R6174 VSS.n1829 VSS.t13 2.25428
R6175 VSS.n1830 VSS.t63 2.25428
R6176 VSS.n1831 VSS.t74 2.25428
R6177 VSS.n1832 VSS.t50 2.25428
R6178 VSS.n1833 VSS.t126 2.25428
R6179 VSS.n1834 VSS.t129 2.25428
R6180 VSS.n1835 VSS.t110 2.25428
R6181 VSS.n1836 VSS.t56 2.25428
R6182 VSS.n1792 VSS.t45 2.25428
R6183 VSS.n1793 VSS.t23 2.25428
R6184 VSS.n1794 VSS.t100 2.25428
R6185 VSS.n1795 VSS.t106 2.25428
R6186 VSS.n1796 VSS.t19 2.25428
R6187 VSS.n1797 VSS.t29 2.25428
R6188 VSS.n1798 VSS.t4 2.25428
R6189 VSS.n1799 VSS.t88 2.25428
R6190 VSS.n1800 VSS.t92 2.25428
R6191 VSS.n1801 VSS.t67 2.25428
R6192 VSS.n1802 VSS.t12 2.25428
R6193 VSS.n1771 VSS.t42 2.25428
R6194 VSS.n1772 VSS.t20 2.25428
R6195 VSS.n1773 VSS.t98 2.25428
R6196 VSS.n1774 VSS.t104 2.25428
R6197 VSS.n1775 VSS.t15 2.25428
R6198 VSS.n1776 VSS.t26 2.25428
R6199 VSS.n1777 VSS.t3 2.25428
R6200 VSS.n1778 VSS.t86 2.25428
R6201 VSS.n1779 VSS.t89 2.25428
R6202 VSS.n1780 VSS.t64 2.25428
R6203 VSS.n1781 VSS.t11 2.25428
R6204 VSS.n1743 VSS.t71 2.25428
R6205 VSS.n1744 VSS.t47 2.25428
R6206 VSS.n1745 VSS.t119 2.25428
R6207 VSS.n1746 VSS.t125 2.25428
R6208 VSS.n1747 VSS.t46 2.25428
R6209 VSS.n1748 VSS.t52 2.25428
R6210 VSS.n1749 VSS.t31 2.25428
R6211 VSS.n1750 VSS.t111 2.25428
R6212 VSS.n1751 VSS.t115 2.25428
R6213 VSS.n1752 VSS.t96 2.25428
R6214 VSS.n1753 VSS.t38 2.25428
R6215 VSS.n1719 VSS.t431 2.25416
R6216 VSS.n1728 VSS.t432 2.25416
R6217 VSS.n1720 VSS.t435 2.25416
R6218 VSS.n1662 VSS.n1661 2.2531
R6219 VSS.n1669 VSS.n1665 2.2531
R6220 VSS.n3907 VSS.n3906 2.25293
R6221 VSS.n1402 VSS.n1401 2.25285
R6222 VSS.n1656 VSS.n1654 2.25253
R6223 VSS.n2491 VSS.n2478 2.25113
R6224 VSS.n1686 VSS.n1685 2.25077
R6225 VSS.n319 VSS.n318 2.2505
R6226 VSS.n1455 VSS.n1454 2.2505
R6227 VSS.n1513 VSS.n1512 2.2505
R6228 VSS.n3995 VSS.n3990 2.2505
R6229 VSS.n1502 VSS.n1501 2.2505
R6230 VSS.n337 VSS.n336 2.2505
R6231 VSS.n357 VSS.n356 2.2505
R6232 VSS.n1645 VSS.n1644 2.2505
R6233 VSS.n1579 VSS.n1578 2.2505
R6234 VSS.n1571 VSS.n1570 2.2505
R6235 VSS.n1569 VSS.n1568 2.2505
R6236 VSS.n1577 VSS.n1576 2.2505
R6237 VSS.n3397 VSS.n3369 2.2505
R6238 VSS.n3388 VSS.n3372 2.2505
R6239 VSS.n3403 VSS.n3367 2.2505
R6240 VSS.n3396 VSS.n3370 2.2505
R6241 VSS.n3386 VSS.n3373 2.2505
R6242 VSS.n3398 VSS.n3368 2.2505
R6243 VSS.n3379 VSS.n3375 2.2505
R6244 VSS.n3382 VSS.n3374 2.2505
R6245 VSS.n3390 VSS.n3371 2.2505
R6246 VSS.n3078 VSS.n3077 2.2505
R6247 VSS.n3229 VSS.n3206 2.2505
R6248 VSS.n3074 VSS.n3073 2.2505
R6249 VSS.n3082 VSS.n3081 2.2505
R6250 VSS.n3213 VSS.n3212 2.2505
R6251 VSS.n3224 VSS.n3223 2.2505
R6252 VSS.n3219 VSS.n3208 2.2505
R6253 VSS.n3225 VSS.n3207 2.2505
R6254 VSS.n3216 VSS.n3209 2.2505
R6255 VSS.n2923 VSS.n2922 2.2505
R6256 VSS.n2952 VSS.n2951 2.2505
R6257 VSS.n2938 VSS.n2937 2.2505
R6258 VSS.n2927 VSS.n2926 2.2505
R6259 VSS.n2948 VSS.n2947 2.2505
R6260 VSS.n2942 VSS.n2941 2.2505
R6261 VSS.n2931 VSS.n2930 2.2505
R6262 VSS.n2950 VSS.n2949 2.2505
R6263 VSS.n2936 VSS.n2935 2.2505
R6264 VSS.n1858 VSS.n1857 2.2505
R6265 VSS.n1847 VSS.n1843 2.2505
R6266 VSS.n1854 VSS.n1840 2.2505
R6267 VSS.n1870 VSS.n1837 2.2505
R6268 VSS.n1859 VSS.n1839 2.2505
R6269 VSS.n1849 VSS.n1841 2.2505
R6270 VSS.n1864 VSS.n1863 2.2505
R6271 VSS.n1848 VSS.n1842 2.2505
R6272 VSS.n1867 VSS.n1838 2.2505
R6273 VSS.n2798 VSS.n2797 2.2505
R6274 VSS.n2017 VSS.n1995 2.2505
R6275 VSS.n2801 VSS.n2080 2.2505
R6276 VSS.n2024 VSS.n2022 2.2505
R6277 VSS.n2021 VSS.n2020 2.2505
R6278 VSS.n2844 VSS.n2843 2.2505
R6279 VSS.n2796 VSS.n2047 2.2505
R6280 VSS.n2856 VSS.n2855 2.2505
R6281 VSS.n2800 VSS.n2799 2.2505
R6282 VSS.n2854 VSS.n2853 2.2505
R6283 VSS.n2130 VSS.n2108 2.2505
R6284 VSS.n2192 VSS.n2191 2.2505
R6285 VSS.n2753 VSS.n2143 2.2505
R6286 VSS.n2137 VSS.n2131 2.2505
R6287 VSS.n2190 VSS.n2177 2.2505
R6288 VSS.n2189 VSS.n2179 2.2505
R6289 VSS.n2141 VSS.n2140 2.2505
R6290 VSS.n2755 VSS.n2754 2.2505
R6291 VSS.n2142 VSS.n2127 2.2505
R6292 VSS.n2102 VSS.n2094 2.2505
R6293 VSS.n2293 VSS.n2235 2.2505
R6294 VSS.n2292 VSS.n2234 2.2505
R6295 VSS.n2308 VSS.n2277 2.2505
R6296 VSS.n2307 VSS.n2306 2.2505
R6297 VSS.n2297 VSS.n2284 2.2505
R6298 VSS.n2296 VSS.n2295 2.2505
R6299 VSS.n2230 VSS.n2212 2.2505
R6300 VSS.n2294 VSS.n2247 2.2505
R6301 VSS.n2571 VSS.n2361 2.2505
R6302 VSS.n2579 VSS.n2578 2.2505
R6303 VSS.n2570 VSS.n2360 2.2505
R6304 VSS.n2331 VSS.n2320 2.2505
R6305 VSS.n2575 VSS.n2574 2.2505
R6306 VSS.n2577 VSS.n2568 2.2505
R6307 VSS.n2573 VSS.n2572 2.2505
R6308 VSS.n2569 VSS.n2346 2.2505
R6309 VSS.n2640 VSS.n2332 2.2505
R6310 VSS.n2368 VSS.n2362 2.2505
R6311 VSS.n2485 VSS.n2451 2.2505
R6312 VSS.n2484 VSS.n2440 2.2505
R6313 VSS.n2486 VSS.n2474 2.2505
R6314 VSS.n2546 VSS.n2545 2.2505
R6315 VSS.n2530 VSS.n2439 2.2505
R6316 VSS.n2543 VSS.n2542 2.2505
R6317 VSS.n2426 VSS.n2413 2.2505
R6318 VSS.n2541 VSS.n2540 2.2505
R6319 VSS.n2548 VSS.n2547 2.2505
R6320 VSS.n2549 VSS.n2421 2.2505
R6321 VSS.n2539 VSS.n2538 2.2505
R6322 VSS.n3908 VSS.n3907 2.2505
R6323 VSS.n1673 VSS.n1672 2.2505
R6324 VSS.n1687 VSS.n1686 2.2505
R6325 VSS.n4162 VSS.n4161 2.2505
R6326 VSS.n4174 VSS.n4173 2.2505
R6327 VSS.n5795 VSS.n5773 2.2505
R6328 VSS.n5805 VSS.n5804 2.2505
R6329 VSS.n3845 VSS.n1727 2.24994
R6330 VSS.n1678 VSS.n1677 2.24918
R6331 VSS.n972 VSS.n971 2.24654
R6332 VSS.n912 VSS.n911 2.24654
R6333 VSS.n3844 VSS.n3843 2.24495
R6334 VSS.n1662 VSS.n1660 2.24449
R6335 VSS.n1656 VSS.n1655 2.24449
R6336 VSS.n1669 VSS.n1668 2.24449
R6337 VSS.n3907 VSS.n1690 2.24449
R6338 VSS.n469 VSS.n468 2.22001
R6339 VSS.n295 VSS.n293 2.04928
R6340 VSS.n5878 VSS.n5877 2.03445
R6341 VSS.n910 VSS.t747 2.02838
R6342 VSS.n1393 VSS.t732 2.02837
R6343 VSS.n324 VSS.t676 2.02837
R6344 VSS.t192 VSS.t228 2.02605
R6345 VSS.t176 VSS.t192 2.02605
R6346 VSS.n5209 VSS.t284 2.02605
R6347 VSS.n4209 VSS.n4208 2.0097
R6348 VSS.n970 VSS.n969 2.00969
R6349 VSS.n280 VSS.n279 2.00969
R6350 VSS.n293 VSS.n278 1.96391
R6351 VSS VSS.n4737 1.9362
R6352 VSS.t260 VSS.t561 1.92472
R6353 VSS.t580 VSS.t583 1.92472
R6354 VSS.t263 VSS.t564 1.92472
R6355 VSS.t476 VSS.t447 1.92472
R6356 VSS.t470 VSS.t733 1.92472
R6357 VSS.t486 VSS.t729 1.92472
R6358 VSS.t489 VSS.t486 1.92472
R6359 VSS.t485 VSS.t728 1.92472
R6360 VSS.t484 VSS.t485 1.92472
R6361 VSS.t493 VSS.t569 1.92244
R6362 VSS.t487 VSS.t572 1.92244
R6363 VSS.t490 VSS.t575 1.92244
R6364 VSS.n4469 VSS.n4468 1.90368
R6365 VSS.n1318 VSS.n1317 1.87586
R6366 VSS.n4221 VSS.n4220 1.87586
R6367 VSS.n224 VSS.n223 1.85787
R6368 VSS.n126 VSS.n125 1.85767
R6369 VSS.n5196 VSS.n5195 1.85765
R6370 VSS.n4776 VSS.n4775 1.85765
R6371 VSS.n5887 VSS.n5725 1.85285
R6372 VSS.n250 VSS.n249 1.83785
R6373 VSS.n4388 VSS.n4387 1.83785
R6374 VSS.n4562 VSS.n4561 1.83785
R6375 VSS.n4394 VSS.n4393 1.83724
R6376 VSS.n5261 VSS.n5260 1.83716
R6377 VSS.n50 VSS.n49 1.83716
R6378 VSS.n4417 VSS.n4416 1.83716
R6379 VSS.n5311 VSS.n5310 1.83716
R6380 VSS.n5289 VSS.n5288 1.83716
R6381 VSS.n4764 VSS.n4763 1.83716
R6382 VSS.n5249 VSS.n5248 1.83716
R6383 VSS.n5051 VSS.n5050 1.83716
R6384 VSS.n5070 VSS.n5069 1.83716
R6385 VSS.n5077 VSS.n5076 1.83716
R6386 VSS.n5100 VSS.n5099 1.83716
R6387 VSS.n5121 VSS.n5120 1.83716
R6388 VSS.n884 VSS.n883 1.82536
R6389 VSS.n970 VSS.t719 1.82525
R6390 VSS.n280 VSS.t742 1.82525
R6391 VSS.n4209 VSS.t669 1.82525
R6392 VSS.n1507 VSS.n1506 1.82479
R6393 VSS.n5788 VSS.n5783 1.80764
R6394 VSS.n1393 VSS.n1392 1.80405
R6395 VSS.n324 VSS.n323 1.80405
R6396 VSS.n910 VSS.n909 1.80404
R6397 VSS.n503 VSS.n500 1.8001
R6398 VSS.n4308 VSS.n4301 1.8001
R6399 VSS.n3913 VSS.n3910 1.8001
R6400 VSS.n4045 VSS.n4044 1.8001
R6401 VSS.n365 VSS.n364 1.8001
R6402 VSS.n490 VSS.n489 1.79951
R6403 VSS.n503 VSS.n502 1.79951
R6404 VSS.n4308 VSS.n4307 1.79951
R6405 VSS.n4274 VSS.n4271 1.79951
R6406 VSS.n3913 VSS.n3912 1.79951
R6407 VSS.n4108 VSS.n4104 1.79951
R6408 VSS.n4282 VSS.n4281 1.79942
R6409 VSS.n901 VSS.n900 1.79942
R6410 VSS.n469 VSS.n466 1.79318
R6411 VSS.n4025 VSS.n4022 1.7505
R6412 VSS.n119 VSS.n118 1.7445
R6413 VSS.n1329 VSS.n1328 1.68421
R6414 VSS.n1335 VSS.n1334 1.68421
R6415 VSS.n4116 VSS.n4114 1.68421
R6416 VSS.n1349 VSS.n1348 1.68411
R6417 VSS.n1354 VSS.n1353 1.68411
R6418 VSS.n1359 VSS.n1358 1.68411
R6419 VSS.n1364 VSS.n1363 1.68411
R6420 VSS.n1370 VSS.n1369 1.68411
R6421 VSS.n1287 VSS.n1286 1.68411
R6422 VSS.n928 VSS.n927 1.65879
R6423 VSS.n934 VSS.n933 1.65879
R6424 VSS.n944 VSS.n943 1.65879
R6425 VSS.n935 VSS.n934 1.65822
R6426 VSS.n941 VSS.n940 1.65822
R6427 VSS.n4142 VSS.n4141 1.65811
R6428 VSS.n834 VSS.n830 1.65328
R6429 VSS.n342 VSS.n341 1.62245
R6430 VSS.n4981 VSS.n4980 1.60209
R6431 VSS.n4595 VSS.n4594 1.60209
R6432 VSS.n4576 VSS.n4575 1.60209
R6433 VSS.n4667 VSS.n4666 1.60209
R6434 VSS.n4565 VSS.n4564 1.60209
R6435 VSS.n5285 VSS.n5284 1.60209
R6436 VSS.n5408 VSS.n5407 1.60199
R6437 VSS.n4962 VSS.n4961 1.60199
R6438 VSS.n37 VSS.n36 1.60199
R6439 VSS.n43 VSS.n42 1.60199
R6440 VSS.n53 VSS.n52 1.60199
R6441 VSS.n4671 VSS.n4670 1.60199
R6442 VSS.n4658 VSS.n4657 1.60199
R6443 VSS.n4573 VSS.n4572 1.60199
R6444 VSS.n4592 VSS.n4591 1.60199
R6445 VSS.n4603 VSS.n4602 1.60199
R6446 VSS.n4426 VSS.n4425 1.60199
R6447 VSS.n4421 VSS.n4420 1.60199
R6448 VSS.n510 VSS.n506 1.59295
R6449 VSS.n4318 VSS.n4317 1.59295
R6450 VSS.n510 VSS.n509 1.5924
R6451 VSS.n4339 VSS.n4338 1.59228
R6452 VSS.n4323 VSS.n4322 1.59228
R6453 VSS.n4353 VSS.n4352 1.59228
R6454 VSS.n690 VSS.n689 1.58814
R6455 VSS.n597 VSS.n596 1.58759
R6456 VSS.n5635 VSS.n5634 1.58759
R6457 VSS.n5645 VSS.n5644 1.58747
R6458 VSS.n5640 VSS.n5639 1.58747
R6459 VSS.n262 VSS.n259 1.56241
R6460 VSS.n4231 VSS.n4230 1.55933
R6461 VSS.n904 VSS.n903 1.55922
R6462 VSS.n4240 VSS.n4239 1.55922
R6463 VSS.n1466 VSS.n1464 1.55606
R6464 VSS.n1648 VSS.n1647 1.50717
R6465 VSS.n1647 VSS.n1646 1.50266
R6466 VSS.n3906 VSS.n3905 1.5016
R6467 VSS.n299 VSS.n297 1.5005
R6468 VSS.n1552 VSS.n1551 1.5005
R6469 VSS.n3897 VSS.n3896 1.5005
R6470 VSS.n3902 VSS.n3901 1.5005
R6471 VSS.n1726 VSS.n1725 1.5005
R6472 VSS.n3838 VSS.n3837 1.5005
R6473 VSS.n3753 VSS.n3752 1.5005
R6474 VSS.n3805 VSS.n3804 1.5005
R6475 VSS.n3825 VSS.n3824 1.5005
R6476 VSS.n3769 VSS.n3768 1.5005
R6477 VSS.n3780 VSS.n3779 1.5005
R6478 VSS.n1542 VSS.n1541 1.5005
R6479 VSS.n5760 VSS.t506 1.463
R6480 VSS.n5760 VSS.n5759 1.463
R6481 VSS.n5871 VSS.t638 1.463
R6482 VSS.n5871 VSS.n5870 1.463
R6483 VSS.n5848 VSS.t710 1.463
R6484 VSS.n5848 VSS.n5847 1.463
R6485 VSS.n5845 VSS.t662 1.463
R6486 VSS.n5845 VSS.n5844 1.463
R6487 VSS.n5843 VSS.t651 1.463
R6488 VSS.n5843 VSS.n5842 1.463
R6489 VSS.n5856 VSS.t679 1.463
R6490 VSS.n5856 VSS.n5855 1.463
R6491 VSS.n5854 VSS.t226 1.463
R6492 VSS.n5854 VSS.n5853 1.463
R6493 VSS.n5864 VSS.t444 1.463
R6494 VSS.n5864 VSS.n5863 1.463
R6495 VSS.n4747 VSS.t462 1.463
R6496 VSS.n4747 VSS.n4746 1.463
R6497 VSS.n5800 VSS.t633 1.463
R6498 VSS.n5800 VSS.n5799 1.463
R6499 VSS.n5808 VSS.t419 1.463
R6500 VSS.n5808 VSS.n5807 1.463
R6501 VSS.n5762 VSS.t664 1.463
R6502 VSS.n5762 VSS.n5761 1.463
R6503 VSS.n5765 VSS.t627 1.463
R6504 VSS.n5765 VSS.n5764 1.463
R6505 VSS.n5767 VSS.t643 1.463
R6506 VSS.n5767 VSS.n5766 1.463
R6507 VSS.n5775 VSS.t687 1.463
R6508 VSS.n5775 VSS.n5774 1.463
R6509 VSS.n5777 VSS.t510 1.463
R6510 VSS.n5777 VSS.n5776 1.463
R6511 VSS.n5657 VSS.n5656 1.4595
R6512 VSS.n4688 VSS.n4687 1.45883
R6513 VSS.n1520 VSS.n1516 1.45883
R6514 VSS.n5530 VSS.n5529 1.43813
R6515 VSS.n1256 VSS.n1255 1.43195
R6516 VSS.n1170 VSS.n1169 1.43182
R6517 VSS.n1344 VSS.n1343 1.43182
R6518 VSS.n1282 VSS.n1281 1.43182
R6519 VSS.n1306 VSS.n1305 1.43182
R6520 VSS.n1300 VSS.n1299 1.43182
R6521 VSS.n4193 VSS.n4192 1.36161
R6522 VSS.n979 VSS.n978 1.33389
R6523 VSS.n991 VSS.n990 1.33389
R6524 VSS.n982 VSS.n981 1.33375
R6525 VSS.n98 VSS.n97 1.33375
R6526 VSS.n4348 VSS.n4347 1.33375
R6527 VSS.n4342 VSS.n4341 1.33375
R6528 VSS.n4333 VSS.n4332 1.33375
R6529 VSS.n4326 VSS.n4325 1.33375
R6530 VSS.n5323 VSS.n5322 1.32883
R6531 VSS.n565 VSS.n564 1.32883
R6532 VSS.n684 VSS.n683 1.32883
R6533 VSS.n5659 VSS.n5658 1.32883
R6534 VSS.n5629 VSS.n5628 1.32883
R6535 VSS.n5618 VSS.n5617 1.32883
R6536 VSS.n1017 VSS.n1016 1.32883
R6537 VSS.n672 VSS.n671 1.32869
R6538 VSS.n553 VSS.n552 1.32869
R6539 VSS.n5335 VSS.n5334 1.32869
R6540 VSS.n4751 VSS.n4750 1.32869
R6541 VSS.n5649 VSS.n5648 1.32869
R6542 VSS.n5621 VSS.n5620 1.32869
R6543 VSS.n5604 VSS.n5603 1.32869
R6544 VSS.n1020 VSS.n1019 1.32869
R6545 VSS.n5300 VSS.n5299 1.27022
R6546 VSS.n4405 VSS.n4404 1.26985
R6547 VSS.n1023 VSS.n1022 1.26929
R6548 VSS.n1000 VSS.n999 1.26929
R6549 VSS.n18 VSS.n17 1.26929
R6550 VSS.n6056 VSS.n6055 1.26929
R6551 VSS.n4158 VSS.n4149 1.26439
R6552 VSS.n4179 VSS.n4176 1.26439
R6553 VSS.n4966 VSS.n4946 1.22037
R6554 VSS.n5771 VSS.t654 1.19623
R6555 VSS.t502 VSS.n5817 1.19623
R6556 VSS.n4002 VSS.n3998 1.16717
R6557 VSS.n1764 VSS.n1763 1.16276
R6558 VSS.n1763 VSS.n1762 1.16276
R6559 VSS.n1762 VSS.n1761 1.16276
R6560 VSS.n1761 VSS.n1760 1.16276
R6561 VSS.n1760 VSS.n1759 1.16276
R6562 VSS.n1759 VSS.n1758 1.16276
R6563 VSS.n1758 VSS.n1757 1.16276
R6564 VSS.n1757 VSS.n1756 1.16276
R6565 VSS.n1756 VSS.n1755 1.16276
R6566 VSS.n1755 VSS.n1754 1.16276
R6567 VSS.n2468 VSS.n2467 1.16276
R6568 VSS.n2467 VSS.n2466 1.16276
R6569 VSS.n2466 VSS.n2465 1.16276
R6570 VSS.n2465 VSS.n2464 1.16276
R6571 VSS.n2464 VSS.n2463 1.16276
R6572 VSS.n2463 VSS.n2462 1.16276
R6573 VSS.n2462 VSS.n2461 1.16276
R6574 VSS.n2461 VSS.n2460 1.16276
R6575 VSS.n2460 VSS.n2459 1.16276
R6576 VSS.n2459 VSS.n2458 1.16276
R6577 VSS.n2382 VSS.n2381 1.16276
R6578 VSS.n2381 VSS.n2380 1.16276
R6579 VSS.n2380 VSS.n2379 1.16276
R6580 VSS.n2379 VSS.n2378 1.16276
R6581 VSS.n2378 VSS.n2377 1.16276
R6582 VSS.n2377 VSS.n2376 1.16276
R6583 VSS.n2376 VSS.n2375 1.16276
R6584 VSS.n2375 VSS.n2374 1.16276
R6585 VSS.n2374 VSS.n2373 1.16276
R6586 VSS.n2373 VSS.n2372 1.16276
R6587 VSS.n2265 VSS.n2264 1.16276
R6588 VSS.n2264 VSS.n2263 1.16276
R6589 VSS.n2263 VSS.n2262 1.16276
R6590 VSS.n2262 VSS.n2261 1.16276
R6591 VSS.n2261 VSS.n2260 1.16276
R6592 VSS.n2260 VSS.n2259 1.16276
R6593 VSS.n2259 VSS.n2258 1.16276
R6594 VSS.n2258 VSS.n2257 1.16276
R6595 VSS.n2257 VSS.n2256 1.16276
R6596 VSS.n2256 VSS.n2255 1.16276
R6597 VSS.n2158 VSS.n2157 1.16276
R6598 VSS.n2157 VSS.n2156 1.16276
R6599 VSS.n2156 VSS.n2155 1.16276
R6600 VSS.n2155 VSS.n2154 1.16276
R6601 VSS.n2154 VSS.n2153 1.16276
R6602 VSS.n2153 VSS.n2152 1.16276
R6603 VSS.n2152 VSS.n2151 1.16276
R6604 VSS.n2151 VSS.n2150 1.16276
R6605 VSS.n2150 VSS.n2149 1.16276
R6606 VSS.n2149 VSS.n2148 1.16276
R6607 VSS.n2061 VSS.n2060 1.16276
R6608 VSS.n2060 VSS.n2059 1.16276
R6609 VSS.n2059 VSS.n2058 1.16276
R6610 VSS.n2058 VSS.n2057 1.16276
R6611 VSS.n2057 VSS.n2056 1.16276
R6612 VSS.n2056 VSS.n2055 1.16276
R6613 VSS.n2055 VSS.n2054 1.16276
R6614 VSS.n2054 VSS.n2053 1.16276
R6615 VSS.n2053 VSS.n2052 1.16276
R6616 VSS.n2052 VSS.n2051 1.16276
R6617 VSS.n1991 VSS.n1990 1.16276
R6618 VSS.n1990 VSS.n1989 1.16276
R6619 VSS.n1989 VSS.n1988 1.16276
R6620 VSS.n1988 VSS.n1987 1.16276
R6621 VSS.n1987 VSS.n1986 1.16276
R6622 VSS.n1986 VSS.n1985 1.16276
R6623 VSS.n1985 VSS.n1984 1.16276
R6624 VSS.n1984 VSS.n1983 1.16276
R6625 VSS.n1983 VSS.n1982 1.16276
R6626 VSS.n1982 VSS.n1981 1.16276
R6627 VSS.n1836 VSS.n1835 1.16276
R6628 VSS.n1835 VSS.n1834 1.16276
R6629 VSS.n1834 VSS.n1833 1.16276
R6630 VSS.n1833 VSS.n1832 1.16276
R6631 VSS.n1832 VSS.n1831 1.16276
R6632 VSS.n1831 VSS.n1830 1.16276
R6633 VSS.n1830 VSS.n1829 1.16276
R6634 VSS.n1829 VSS.n1828 1.16276
R6635 VSS.n1828 VSS.n1827 1.16276
R6636 VSS.n1827 VSS.n1826 1.16276
R6637 VSS.n1802 VSS.n1801 1.16276
R6638 VSS.n1801 VSS.n1800 1.16276
R6639 VSS.n1800 VSS.n1799 1.16276
R6640 VSS.n1799 VSS.n1798 1.16276
R6641 VSS.n1798 VSS.n1797 1.16276
R6642 VSS.n1797 VSS.n1796 1.16276
R6643 VSS.n1796 VSS.n1795 1.16276
R6644 VSS.n1795 VSS.n1794 1.16276
R6645 VSS.n1794 VSS.n1793 1.16276
R6646 VSS.n1793 VSS.n1792 1.16276
R6647 VSS.n1781 VSS.n1780 1.16276
R6648 VSS.n1780 VSS.n1779 1.16276
R6649 VSS.n1779 VSS.n1778 1.16276
R6650 VSS.n1778 VSS.n1777 1.16276
R6651 VSS.n1777 VSS.n1776 1.16276
R6652 VSS.n1776 VSS.n1775 1.16276
R6653 VSS.n1775 VSS.n1774 1.16276
R6654 VSS.n1774 VSS.n1773 1.16276
R6655 VSS.n1773 VSS.n1772 1.16276
R6656 VSS.n1772 VSS.n1771 1.16276
R6657 VSS.n1753 VSS.n1752 1.16276
R6658 VSS.n1752 VSS.n1751 1.16276
R6659 VSS.n1751 VSS.n1750 1.16276
R6660 VSS.n1750 VSS.n1749 1.16276
R6661 VSS.n1749 VSS.n1748 1.16276
R6662 VSS.n1748 VSS.n1747 1.16276
R6663 VSS.n1747 VSS.n1746 1.16276
R6664 VSS.n1746 VSS.n1745 1.16276
R6665 VSS.n1745 VSS.n1744 1.16276
R6666 VSS.n1744 VSS.n1743 1.16276
R6667 VSS.n4974 VSS.n4907 1.15537
R6668 VSS.n3589 VSS.n3588 1.13934
R6669 VSS.n2487 VSS.n2486 1.12652
R6670 VSS.n353 VSS.n349 1.12642
R6671 VSS.n1447 VSS.n1446 1.1255
R6672 VSS.n318 VSS.n317 1.1255
R6673 VSS.n3822 VSS.n3821 1.1255
R6674 VSS.n3835 VSS.n3831 1.1255
R6675 VSS.n3750 VSS.n3749 1.1255
R6676 VSS.n3802 VSS.n3797 1.1255
R6677 VSS.n3766 VSS.n3761 1.1255
R6678 VSS.n3789 VSS.n3788 1.1255
R6679 VSS.n1742 VSS.n1741 1.1255
R6680 VSS.n3529 VSS.n3506 1.1255
R6681 VSS.n1770 VSS.n1769 1.1255
R6682 VSS.n1791 VSS.n1790 1.1255
R6683 VSS.n1825 VSS.n1824 1.1255
R6684 VSS.n1964 VSS.n1963 1.1255
R6685 VSS.n2026 VSS.n2024 1.1255
R6686 VSS.n2798 VSS.n2073 1.1255
R6687 VSS.n2853 VSS.n2852 1.1255
R6688 VSS.n2818 VSS.n2080 1.1255
R6689 VSS.n2020 VSS.n2007 1.1255
R6690 VSS.n2856 VSS.n2013 1.1255
R6691 VSS.n2048 VSS.n2047 1.1255
R6692 VSS.n2799 VSS.n2079 1.1255
R6693 VSS.n2017 VSS.n2002 1.1255
R6694 VSS.n1994 VSS.n1993 1.1255
R6695 VSS.n2779 VSS.n2102 1.1255
R6696 VSS.n2756 VSS.n2127 1.1255
R6697 VSS.n2188 VSS.n2169 1.1255
R6698 VSS.n2189 VSS.n2188 1.1255
R6699 VSS.n2774 VSS.n2108 1.1255
R6700 VSS.n2190 VSS.n2171 1.1255
R6701 VSS.n2137 VSS.n2115 1.1255
R6702 VSS.n2191 VSS.n2172 1.1255
R6703 VSS.n2704 VSS.n2234 1.1255
R6704 VSS.n2230 VSS.n2219 1.1255
R6705 VSS.n2691 VSS.n2247 1.1255
R6706 VSS.n2296 VSS.n2252 1.1255
R6707 VSS.n2306 VSS.n2275 1.1255
R6708 VSS.n2703 VSS.n2235 1.1255
R6709 VSS.n2297 VSS.n2253 1.1255
R6710 VSS.n2670 VSS.n2277 1.1255
R6711 VSS.n2640 VSS.n2639 1.1255
R6712 VSS.n2572 VSS.n2364 1.1255
R6713 VSS.n2575 VSS.n2395 1.1255
R6714 VSS.n2331 VSS.n2329 1.1255
R6715 VSS.n2329 VSS.n2325 1.1255
R6716 VSS.n2624 VSS.n2360 1.1255
R6717 VSS.n2577 VSS.n2576 1.1255
R6718 VSS.n2623 VSS.n2361 1.1255
R6719 VSS.n2578 VSS.n2399 1.1255
R6720 VSS.n2632 VSS.n2346 1.1255
R6721 VSS.n2544 VSS.n2429 1.1255
R6722 VSS.n2426 VSS.n2416 1.1255
R6723 VSS.n2530 VSS.n2438 1.1255
R6724 VSS.n2502 VSS.n2474 1.1255
R6725 VSS.n2483 VSS.n2475 1.1255
R6726 VSS.n2527 VSS.n2440 1.1255
R6727 VSS.n2488 VSS.n2479 1.1255
R6728 VSS.n2521 VSS.n2451 1.1255
R6729 VSS.n2418 VSS.n2416 1.1255
R6730 VSS.n2552 VSS.n2418 1.1255
R6731 VSS.n2502 VSS.n2501 1.1255
R6732 VSS.n2501 VSS.n2500 1.1255
R6733 VSS.n2436 VSS.n2434 1.1255
R6734 VSS.n2438 VSS.n2436 1.1255
R6735 VSS.n2411 VSS.n2410 1.1255
R6736 VSS.n2412 VSS.n2411 1.1255
R6737 VSS.n2477 VSS.n2475 1.1255
R6738 VSS.n2499 VSS.n2477 1.1255
R6739 VSS.n2526 VSS.n2525 1.1255
R6740 VSS.n2527 VSS.n2526 1.1255
R6741 VSS.n2497 VSS.n2479 1.1255
R6742 VSS.n2498 VSS.n2497 1.1255
R6743 VSS.n2522 VSS.n2447 1.1255
R6744 VSS.n2522 VSS.n2521 1.1255
R6745 VSS.n2648 VSS.n2325 1.1255
R6746 VSS.n2623 VSS.n2352 1.1255
R6747 VSS.n2319 VSS.n2318 1.1255
R6748 VSS.n2583 VSS.n2567 1.1255
R6749 VSS.n2576 VSS.n2394 1.1255
R6750 VSS.n2596 VSS.n2399 1.1255
R6751 VSS.n2600 VSS.n2395 1.1255
R6752 VSS.n2600 VSS.n2599 1.1255
R6753 VSS.n2625 VSS.n2359 1.1255
R6754 VSS.n2625 VSS.n2624 1.1255
R6755 VSS.n2366 VSS.n2364 1.1255
R6756 VSS.n2613 VSS.n2366 1.1255
R6757 VSS.n2597 VSS.n2596 1.1255
R6758 VSS.n2633 VSS.n2338 1.1255
R6759 VSS.n2633 VSS.n2632 1.1255
R6760 VSS.n2639 VSS.n2638 1.1255
R6761 VSS.n2598 VSS.n2394 1.1255
R6762 VSS.n2584 VSS.n2583 1.1255
R6763 VSS.n2638 VSS.n2637 1.1255
R6764 VSS.n2318 VSS.n2317 1.1255
R6765 VSS.n2367 VSS.n2352 1.1255
R6766 VSS.n2310 VSS.n2309 1.1255
R6767 VSS.n2684 VSS.n2252 1.1255
R6768 VSS.n2211 VSS.n2210 1.1255
R6769 VSS.n2683 VSS.n2253 1.1255
R6770 VSS.n2703 VSS.n2227 1.1255
R6771 VSS.n2672 VSS.n2275 1.1255
R6772 VSS.n2692 VSS.n2691 1.1255
R6773 VSS.n2713 VSS.n2219 1.1255
R6774 VSS.n2714 VSS.n2713 1.1255
R6775 VSS.n2693 VSS.n2692 1.1255
R6776 VSS.n2673 VSS.n2672 1.1255
R6777 VSS.n2227 VSS.n2226 1.1255
R6778 VSS.n2683 VSS.n2682 1.1255
R6779 VSS.n2671 VSS.n2274 1.1255
R6780 VSS.n2671 VSS.n2670 1.1255
R6781 VSS.n2705 VSS.n2704 1.1255
R6782 VSS.n2210 VSS.n2209 1.1255
R6783 VSS.n2706 VSS.n2705 1.1255
R6784 VSS.n2684 VSS.n2250 1.1255
R6785 VSS.n2316 VSS.n2310 1.1255
R6786 VSS.n2740 VSS.n2169 1.1255
R6787 VSS.n2737 VSS.n2172 1.1255
R6788 VSS.n2752 VSS.n2751 1.1255
R6789 VSS.n2768 VSS.n2115 1.1255
R6790 VSS.n2738 VSS.n2171 1.1255
R6791 VSS.n2774 VSS.n2773 1.1255
R6792 VSS.n2093 VSS.n2092 1.1255
R6793 VSS.n2760 VSS.n2125 1.1255
R6794 VSS.n2729 VSS.n2728 1.1255
R6795 VSS.n2159 VSS.n2126 1.1255
R6796 VSS.n2756 VSS.n2126 1.1255
R6797 VSS.n2781 VSS.n2780 1.1255
R6798 VSS.n2780 VSS.n2779 1.1255
R6799 VSS.n2761 VSS.n2760 1.1255
R6800 VSS.n2728 VSS.n2727 1.1255
R6801 VSS.n2092 VSS.n2091 1.1255
R6802 VSS.n2773 VSS.n2772 1.1255
R6803 VSS.n2739 VSS.n2738 1.1255
R6804 VSS.n2768 VSS.n2112 1.1255
R6805 VSS.n2751 VSS.n2750 1.1255
R6806 VSS.n2737 VSS.n2170 1.1255
R6807 VSS.n1993 VSS.n1992 1.1255
R6808 VSS.n2865 VSS.n2007 1.1255
R6809 VSS.n2852 VSS.n2851 1.1255
R6810 VSS.n2870 VSS.n2002 1.1255
R6811 VSS.n2079 VSS.n2074 1.1255
R6812 VSS.n2089 VSS.n2087 1.1255
R6813 VSS.n2820 VSS.n2819 1.1255
R6814 VSS.n2819 VSS.n2818 1.1255
R6815 VSS.n2032 VSS.n2011 1.1255
R6816 VSS.n2013 VSS.n2011 1.1255
R6817 VSS.n2050 VSS.n2048 1.1255
R6818 VSS.n2823 VSS.n2073 1.1255
R6819 VSS.n2823 VSS.n2822 1.1255
R6820 VSS.n2090 VSS.n2087 1.1255
R6821 VSS.n2836 VSS.n2050 1.1255
R6822 VSS.n2821 VSS.n2074 1.1255
R6823 VSS.n2871 VSS.n2870 1.1255
R6824 VSS.n2851 VSS.n2850 1.1255
R6825 VSS.n2849 VSS.n2028 1.1255
R6826 VSS.n2028 VSS.n2026 1.1255
R6827 VSS.n2865 VSS.n2864 1.1255
R6828 VSS.n1920 VSS.n1905 1.1255
R6829 VSS.n1945 VSS.n1944 1.1255
R6830 VSS.n1932 VSS.n1895 1.1255
R6831 VSS.n1923 VSS.n1896 1.1255
R6832 VSS.n1911 VSS.n1910 1.1255
R6833 VSS.n1947 VSS.n1946 1.1255
R6834 VSS.n1974 VSS.n1973 1.1255
R6835 VSS.n1954 VSS.n1886 1.1255
R6836 VSS.n1922 VSS.n1921 1.1255
R6837 VSS.n1979 VSS.n1879 1.1255
R6838 VSS.n3052 VSS.n1825 1.1255
R6839 VSS.n3027 VSS.n3022 1.1255
R6840 VSS.n3068 VSS.n3063 1.1255
R6841 VSS.n2961 VSS.n2959 1.1255
R6842 VSS.n2980 VSS.n2973 1.1255
R6843 VSS.n2981 VSS.n2980 1.1255
R6844 VSS.n2999 VSS.n2998 1.1255
R6845 VSS.n2998 VSS.n2997 1.1255
R6846 VSS.n2962 VSS.n2961 1.1255
R6847 VSS.n3014 VSS.n3011 1.1255
R6848 VSS.n3048 VSS.n3044 1.1255
R6849 VSS.n3049 VSS.n3048 1.1255
R6850 VSS.n3015 VSS.n3014 1.1255
R6851 VSS.n2984 VSS.n2983 1.1255
R6852 VSS.n2983 VSS.n2982 1.1255
R6853 VSS.n3037 VSS.n3036 1.1255
R6854 VSS.n3038 VSS.n3037 1.1255
R6855 VSS.n3069 VSS.n3068 1.1255
R6856 VSS.n3028 VSS.n3027 1.1255
R6857 VSS.n1812 VSS.n1808 1.1255
R6858 VSS.n3188 VSS.n1791 1.1255
R6859 VSS.n3102 VSS.n3097 1.1255
R6860 VSS.n3146 VSS.n3145 1.1255
R6861 VSS.n3186 VSS.n3181 1.1255
R6862 VSS.n3239 VSS.n3238 1.1255
R6863 VSS.n3115 VSS.n3110 1.1255
R6864 VSS.n3153 VSS.n3152 1.1255
R6865 VSS.n3089 VSS.n3087 1.1255
R6866 VSS.n3130 VSS.n3129 1.1255
R6867 VSS.n3170 VSS.n3165 1.1255
R6868 VSS.n3171 VSS.n3170 1.1255
R6869 VSS.n3131 VSS.n3130 1.1255
R6870 VSS.n3090 VSS.n3089 1.1255
R6871 VSS.n3198 VSS.n3197 1.1255
R6872 VSS.n3197 VSS.n3196 1.1255
R6873 VSS.n3154 VSS.n3153 1.1255
R6874 VSS.n3116 VSS.n3115 1.1255
R6875 VSS.n3240 VSS.n3239 1.1255
R6876 VSS.n3187 VSS.n3186 1.1255
R6877 VSS.n3147 VSS.n3146 1.1255
R6878 VSS.n3103 VSS.n3102 1.1255
R6879 VSS.n3359 VSS.n1770 1.1255
R6880 VSS.n3294 VSS.n3288 1.1255
R6881 VSS.n3335 VSS.n3328 1.1255
R6882 VSS.n3251 VSS.n3250 1.1255
R6883 VSS.n3298 VSS.n3297 1.1255
R6884 VSS.n3414 VSS.n3413 1.1255
R6885 VSS.n3413 VSS.n3412 1.1255
R6886 VSS.n3353 VSS.n3352 1.1255
R6887 VSS.n3354 VSS.n3353 1.1255
R6888 VSS.n3299 VSS.n3298 1.1255
R6889 VSS.n3252 VSS.n3251 1.1255
R6890 VSS.n3259 VSS.n3258 1.1255
R6891 VSS.n3258 VSS.n3257 1.1255
R6892 VSS.n3338 VSS.n3337 1.1255
R6893 VSS.n3314 VSS.n3311 1.1255
R6894 VSS.n3274 VSS.n3273 1.1255
R6895 VSS.n3339 VSS.n3338 1.1255
R6896 VSS.n3315 VSS.n3314 1.1255
R6897 VSS.n3275 VSS.n3274 1.1255
R6898 VSS.n3336 VSS.n3335 1.1255
R6899 VSS.n3295 VSS.n3294 1.1255
R6900 VSS.n3726 VSS.n1742 1.1255
R6901 VSS.n3662 VSS.n3657 1.1255
R6902 VSS.n3701 VSS.n3695 1.1255
R6903 VSS.n3647 VSS.n3646 1.1255
R6904 VSS.n3622 VSS.n3620 1.1255
R6905 VSS.n3636 VSS.n3631 1.1255
R6906 VSS.n3734 VSS.n3733 1.1255
R6907 VSS.n3721 VSS.n3717 1.1255
R6908 VSS.n3685 VSS.n3684 1.1255
R6909 VSS.n3684 VSS.n3683 1.1255
R6910 VSS.n3665 VSS.n3664 1.1255
R6911 VSS.n3709 VSS.n3708 1.1255
R6912 VSS.n3735 VSS.n3734 1.1255
R6913 VSS.n3710 VSS.n3709 1.1255
R6914 VSS.n3666 VSS.n3665 1.1255
R6915 VSS.n3637 VSS.n3636 1.1255
R6916 VSS.n3623 VSS.n3622 1.1255
R6917 VSS.n3722 VSS.n3721 1.1255
R6918 VSS.n3648 VSS.n3647 1.1255
R6919 VSS.n3702 VSS.n3701 1.1255
R6920 VSS.n3663 VSS.n3662 1.1255
R6921 VSS.n3790 VSS.n3789 1.1255
R6922 VSS.n3767 VSS.n3766 1.1255
R6923 VSS.n3751 VSS.n3750 1.1255
R6924 VSS.n3836 VSS.n3835 1.1255
R6925 VSS.n3803 VSS.n3802 1.1255
R6926 VSS.n3823 VSS.n3822 1.1255
R6927 VSS.n1642 VSS.n1641 1.1255
R6928 VSS.n1503 VSS.n1502 1.1234
R6929 VSS.n1814 VSS.n1813 1.12321
R6930 VSS.n1554 VSS.n1553 1.12277
R6931 VSS.n1544 VSS.n1543 1.12277
R6932 VSS.n5866 VSS.t253 1.10896
R6933 VSS.n5892 VSS.t457 1.10896
R6934 VSS.n316 VSS.n315 1.09796
R6935 VSS.n4012 VSS.n4011 1.06994
R6936 VSS.n4002 VSS.n4001 1.06994
R6937 VSS.n690 VSS.n688 1.03151
R6938 VSS.n916 VSS.n914 1.02489
R6939 VSS.n1397 VSS.n1395 1.02489
R6940 VSS.t136 VSS.t240 1.01328
R6941 VSS.n5119 VSS.n5117 1.01328
R6942 VSS.t233 VSS.t167 1.01328
R6943 VSS.t167 VSS.t142 1.01328
R6944 VSS.n1284 VSS.n1168 1.0102
R6945 VSS.n5794 VSS.n5793 0.999031
R6946 VSS.n4158 VSS.n4157 0.972722
R6947 VSS.n4179 VSS.n4178 0.972722
R6948 VSS.n27 VSS.n26 0.967979
R6949 VSS.n2915 VSS.n1980 0.96059
R6950 VSS.n4150 VSS.t737 0.93818
R6951 VSS.n1322 VSS.n1321 0.93818
R6952 VSS.n1511 VSS.n1510 0.931667
R6953 VSS.n889 VSS.n888 0.929276
R6954 VSS.n879 VSS.n878 0.928071
R6955 VSS.n1450 VSS.n1449 0.925894
R6956 VSS.n4335 VSS.n253 0.919029
R6957 VSS.n4419 VSS.n4355 0.919029
R6958 VSS.n1012 VSS.n1010 0.910283
R6959 VSS.n3086 VSS.n3085 0.900727
R6960 VSS.n2802 VSS.n2795 0.900647
R6961 VSS.n2663 VSS.n2662 0.900647
R6962 VSS.n2140 VSS.n2125 0.9005
R6963 VSS.n2753 VSS.n2752 0.9005
R6964 VSS.n3619 VSS.n3618 0.900467
R6965 VSS.n2958 VSS.n2957 0.900467
R6966 VSS.n2581 VSS.n2580 0.900467
R6967 VSS.n3407 VSS.n3406 0.900443
R6968 VSS.n3233 VSS.n3232 0.900443
R6969 VSS.n2657 VSS.n2656 0.900443
R6970 VSS.n2561 VSS.n2560 0.900442
R6971 VSS.n2880 VSS.n2879 0.900405
R6972 VSS.n2195 VSS.n2193 0.900387
R6973 VSS.n1909 VSS.n1908 0.900368
R6974 VSS.n2790 VSS.n2789 0.900365
R6975 VSS.n2723 VSS.n2722 0.900365
R6976 VSS.n1874 VSS.n1873 0.900347
R6977 VSS.n1556 VSS.n1555 0.900305
R6978 VSS.n1644 VSS.n1643 0.90028
R6979 VSS.n336 VSS.n335 0.898922
R6980 VSS.n1807 VSS.n1806 0.898321
R6981 VSS.n314 VSS.n308 0.897993
R6982 VSS.n1646 VSS.n1645 0.891062
R6983 VSS.n4193 VSS.n4189 0.8755
R6984 VSS.n564 VSS.n563 0.849401
R6985 VSS.n683 VSS.n682 0.849401
R6986 VSS.n5658 VSS.n5657 0.849401
R6987 VSS.n5334 VSS.n5333 0.849205
R6988 VSS.n978 VSS.n977 0.846031
R6989 VSS.n990 VSS.n989 0.846031
R6990 VSS.n4347 VSS.n4346 0.845835
R6991 VSS.n4332 VSS.n4331 0.845835
R6992 VSS.n882 VSS.n874 0.829906
R6993 VSS.n5816 VSS.n5815 0.801258
R6994 VSS.n4137 VSS.n4134 0.79929
R6995 VSS.n5858 VSS 0.793969
R6996 VSS.n5736 VSS.n5735 0.781777
R6997 VSS.n5744 VSS.n5743 0.781777
R6998 VSS.n1299 VSS.n1298 0.780455
R6999 VSS.n4688 VSS.n4685 0.778278
R7000 VSS.n1520 VSS.n1519 0.778278
R7001 VSS.n5782 VSS.n5781 0.772481
R7002 VSS.n315 VSS.n314 0.768418
R7003 VSS.n4203 VSS.n4201 0.726531
R7004 VSS.n5815 VSS.n5763 0.722141
R7005 VSS.n5894 VSS.n5893 0.715474
R7006 VSS.n5865 VSS.n4745 0.703683
R7007 VSS.n4107 VSS.n4106 0.69552
R7008 VSS.n4239 VSS.n4238 0.69552
R7009 VSS.n1033 VSS 0.683795
R7010 VSS.n1464 VSS.n1416 0.681056
R7011 VSS.n4980 VSS.n4979 0.66722
R7012 VSS.n4602 VSS.n4601 0.66701
R7013 VSS.n4591 VSS.n4590 0.66701
R7014 VSS.n4657 VSS.n4656 0.66701
R7015 VSS.n4670 VSS.n4669 0.66701
R7016 VSS.n4572 VSS.n4571 0.66701
R7017 VSS.n3893 VSS.n1719 0.652915
R7018 VSS.n4005 VSS.t536 0.65037
R7019 VSS.n3858 VSS.n1720 0.643803
R7020 VSS.n140 VSS.n137 0.642239
R7021 VSS.n183 VSS.n180 0.642239
R7022 VSS.n238 VSS.n235 0.642239
R7023 VSS.n5176 VSS.n5175 0.642239
R7024 VSS.n5202 VSS.n5201 0.642239
R7025 VSS.n4782 VSS.n4781 0.642239
R7026 VSS.n5859 VSS.n4745 0.618484
R7027 VSS.n2835 VSS.n2061 0.615498
R7028 VSS.n2161 VSS.n2158 0.614262
R7029 VSS.n4501 VSS.n4500 0.611348
R7030 VSS.n5531 VSS.n5530 0.610998
R7031 VSS.n2266 VSS.n2265 0.609999
R7032 VSS.n3431 VSS.n1764 0.609008
R7033 VSS.n3003 VSS.n1836 0.608439
R7034 VSS.n3703 VSS.n1753 0.606848
R7035 VSS.n2612 VSS.n2382 0.606843
R7036 VSS.n3156 VSS.n1802 0.606489
R7037 VSS.n3316 VSS.n1781 0.605607
R7038 VSS.n2896 VSS.n1991 0.601243
R7039 VSS.n235 VSS.n232 0.597879
R7040 VSS.n4781 VSS.n4780 0.597879
R7041 VSS.n137 VSS.n134 0.596788
R7042 VSS.n5201 VSS.n5200 0.596788
R7043 VSS.n180 VSS.n177 0.595696
R7044 VSS.n5175 VSS.n5174 0.595696
R7045 VSS.n2512 VSS.n2468 0.593624
R7046 VSS.n174 VSS.n173 0.587994
R7047 VSS.n5173 VSS.n5172 0.587128
R7048 VSS.n131 VSS.n130 0.586903
R7049 VSS.n5199 VSS.n5198 0.586037
R7050 VSS.n229 VSS.n228 0.585812
R7051 VSS.n4779 VSS.n4778 0.584946
R7052 VSS.n834 VSS.n833 0.583833
R7053 VSS.n5198 VSS.n5197 0.574718
R7054 VSS.n130 VSS.n127 0.574288
R7055 VSS.n4778 VSS.n4777 0.573627
R7056 VSS.n228 VSS.n225 0.573197
R7057 VSS.n3530 VSS.n3529 0.563
R7058 VSS.n2544 VSS.n2425 0.563
R7059 VSS.n2425 VSS.n2423 0.563
R7060 VSS.n2433 VSS.n2423 0.563
R7061 VSS.n3566 VSS.n3530 0.563
R7062 VSS.n3567 VSS.n3566 0.563
R7063 VSS.n1567 VSS.n1566 0.551597
R7064 VSS.n173 VSS.n170 0.550283
R7065 VSS.n5172 VSS.n5171 0.550283
R7066 VSS.n4363 VSS.n4362 0.54076
R7067 VSS.n3738 VSS.n1728 0.534462
R7068 VSS.n5895 VSS.n4744 0.508005
R7069 VSS.n4742 VSS.n4741 0.508005
R7070 VSS.n511 VSS.n510 0.505601
R7071 VSS.n4317 VSS.n4316 0.505601
R7072 VSS.n963 VSS.n962 0.502377
R7073 VSS.n4366 VSS.n4365 0.502362
R7074 VSS.n5269 VSS.n5268 0.502362
R7075 VSS.n4369 VSS.n4368 0.497425
R7076 VSS.n5272 VSS.n5271 0.497402
R7077 VSS.n4025 VSS.n4024 0.486611
R7078 VSS.n5830 VSS.n5745 0.477891
R7079 VSS.n3242 VSS.n3241 0.473104
R7080 VSS.n940 VSS.n939 0.472687
R7081 VSS.n4136 VSS.n4135 0.472687
R7082 VSS.n2660 VSS.n2659 0.467151
R7083 VSS.n3416 VSS.n3415 0.465504
R7084 VSS.n1328 VSS.n1327 0.459689
R7085 VSS.n4117 VSS.n4116 0.459689
R7086 VSS.n1369 VSS.n1368 0.459446
R7087 VSS.n1286 VSS.n1285 0.459446
R7088 VSS.n3842 VSS.n3841 0.459227
R7089 VSS.n2916 VSS.n2915 0.458913
R7090 VSS.n5831 VSS.n5738 0.458326
R7091 VSS.n2726 VSS.n2725 0.456584
R7092 VSS.n2793 VSS.n2792 0.451624
R7093 VSS.n2564 VSS.n2563 0.449946
R7094 VSS.n1403 VSS 0.449668
R7095 VSS.n3072 VSS.n3071 0.443676
R7096 VSS.n3574 VSS.n3573 0.441768
R7097 VSS.n66 VSS.n65 0.435547
R7098 VSS.n5106 VSS.n5105 0.434956
R7099 VSS.n4117 VSS.n4111 0.4313
R7100 VSS.n117 VSS.n116 0.427022
R7101 VSS.n4761 VSS.n4758 0.426043
R7102 VSS VSS.n1402 0.405813
R7103 VSS.n489 VSS.n488 0.402035
R7104 VSS.n4044 VSS.n4043 0.402035
R7105 VSS.n364 VSS.n363 0.402035
R7106 VSS.n504 VSS.n503 0.402035
R7107 VSS.n4309 VSS.n4308 0.402035
R7108 VSS.n4111 VSS.n4108 0.402035
R7109 VSS.n4275 VSS.n4274 0.402035
R7110 VSS.n4273 VSS.n4272 0.402035
R7111 VSS.n3914 VSS.n3913 0.402035
R7112 VSS.n4106 VSS.n4105 0.401791
R7113 VSS.n5475 VSS.n5472 0.393137
R7114 VSS.n4515 VSS.n4512 0.393137
R7115 VSS.n5539 VSS.n5538 0.391771
R7116 VSS.n735 VSS.n732 0.390642
R7117 VSS.n511 VSS.n504 0.390642
R7118 VSS.n773 VSS.n770 0.390642
R7119 VSS.n4312 VSS.n4309 0.390642
R7120 VSS.n28 VSS.n27 0.383479
R7121 VSS.n249 VSS.n248 0.383166
R7122 VSS.n4393 VSS.n4392 0.383166
R7123 VSS.n1014 VSS.n1013 0.383166
R7124 VSS.n49 VSS.n48 0.382921
R7125 VSS.n4416 VSS.n4415 0.382921
R7126 VSS.n4763 VSS.n4762 0.382921
R7127 VSS.n5120 VSS.n5119 0.382921
R7128 VSS.n5119 VSS.n5118 0.382921
R7129 VSS.n4560 VSS.n4510 0.376519
R7130 VSS.n4581 VSS.n87 0.376518
R7131 VSS.n5061 VSS.n5060 0.37489
R7132 VSS.n5075 VSS.n5048 0.374889
R7133 VSS.n5154 VSS.n5153 0.372135
R7134 VSS.n161 VSS.n148 0.372135
R7135 VSS.n4402 VSS.n4401 0.371392
R7136 VSS.n5297 VSS.n5296 0.371022
R7137 VSS.n4399 VSS.n4398 0.370645
R7138 VSS.n5294 VSS.n5293 0.370645
R7139 VSS.n5045 VSS.n5043 0.358977
R7140 VSS.n4613 VSS.n4610 0.358977
R7141 VSS.n4600 VSS.n63 0.356537
R7142 VSS.n5123 VSS.n5046 0.354994
R7143 VSS.n6063 VSS.n28 0.350926
R7144 VSS.n5872 VSS 0.347643
R7145 VSS.n5875 VSS 0.347643
R7146 VSS.n5801 VSS 0.347643
R7147 VSS VSS.n5806 0.347643
R7148 VSS.n5052 VSS.n5049 0.347591
R7149 VSS.n6060 VSS.n6058 0.342028
R7150 VSS.n147 VSS.n146 0.341179
R7151 VSS.n5152 VSS.n5151 0.340476
R7152 VSS.n106 VSS.n105 0.338978
R7153 VSS.n5633 VSS.n5312 0.331895
R7154 VSS.n5616 VSS.n5314 0.331895
R7155 VSS.n3980 VSS.n3977 0.327038
R7156 VSS.n5601 VSS.n5600 0.326081
R7157 VSS.n5098 VSS.n5047 0.321363
R7158 VSS.n4589 VSS.n76 0.320022
R7159 VSS.n5150 VSS.n5149 0.31827
R7160 VSS.n145 VSS.n144 0.318076
R7161 VSS.n4569 VSS.n4509 0.313628
R7162 VSS VSS.n2882 0.307487
R7163 VSS.n259 VSS.n257 0.302495
R7164 VSS.n5647 VSS.n5254 0.301198
R7165 VSS.n1167 VSS.n1166 0.3005
R7166 VSS.n4978 VSS.n4790 0.292445
R7167 VSS.n91 VSS.n90 0.291512
R7168 VSS.n4673 VSS.n58 0.290903
R7169 VSS.n4990 VSS.n4789 0.289506
R7170 VSS.n4970 VSS.n4908 0.288772
R7171 VSS.n4663 VSS.n59 0.287963
R7172 VSS.n57 VSS.n31 0.287229
R7173 VSS.n4949 VSS.n4948 0.285098
R7174 VSS.n4960 VSS.n4947 0.285098
R7175 VSS.n39 VSS.n33 0.283556
R7176 VSS.n47 VSS.n32 0.283556
R7177 VSS.n4275 VSS 0.281962
R7178 VSS.n5815 VSS.n5814 0.281211
R7179 VSS.n240 VSS.n239 0.2753
R7180 VSS.n5232 VSS.n4783 0.2753
R7181 VSS.n3877 VSS.n3876 0.274296
R7182 VSS.n221 VSS.n220 0.2729
R7183 VSS.n5203 VSS.n5185 0.2729
R7184 VSS.n184 VSS.n183 0.272046
R7185 VSS.n5177 VSS.n5176 0.27149
R7186 VSS.n241 VSS.n240 0.269479
R7187 VSS.n5234 VSS.n5232 0.269479
R7188 VSS.n3874 VSS.n3873 0.266088
R7189 VSS.n4503 VSS.n4502 0.254764
R7190 VSS.n220 VSS.n140 0.250935
R7191 VSS.n239 VSS.n238 0.250935
R7192 VSS.n5203 VSS.n5202 0.250935
R7193 VSS.n4783 VSS.n4782 0.250935
R7194 VSS.n5127 VSS.n5126 0.2505
R7195 VSS.n4606 VSS.n4605 0.2505
R7196 VSS.n142 VSS.n141 0.24562
R7197 VSS.n5084 VSS.n5081 0.244911
R7198 VSS.n952 VSS 0.243106
R7199 VSS.n5826 VSS.n5824 0.241879
R7200 VSS.n5303 VSS.n5302 0.241152
R7201 VSS.n5084 VSS.n5083 0.239887
R7202 VSS.n4376 VSS.n4357 0.235283
R7203 VSS.n4252 VSS.n4219 0.224214
R7204 VSS.n94 VSS.n88 0.213053
R7205 VSS.n86 VSS.n77 0.213053
R7206 VSS.n75 VSS.n64 0.213053
R7207 VSS.n5115 VSS.n5104 0.213053
R7208 VSS.n5094 VSS.n5088 0.213053
R7209 VSS.n5087 VSS.n5079 0.213053
R7210 VSS.n5091 VSS.n5090 0.211098
R7211 VSS.n4130 VSS.n908 0.205426
R7212 VSS.n5234 VSS.n5233 0.205144
R7213 VSS.n4873 VSS.n4872 0.205045
R7214 VSS.n5738 VSS.n5736 0.200065
R7215 VSS.n5745 VSS.n5744 0.200065
R7216 VSS.n143 VSS.n142 0.199702
R7217 VSS.n406 VSS.n360 0.1985
R7218 VSS.n4876 VSS.n4873 0.196574
R7219 VSS.n72 VSS.n71 0.196132
R7220 VSS.n5112 VSS.n5111 0.196132
R7221 VSS VSS.n1032 0.195846
R7222 VSS.n4050 VSS.n4031 0.193921
R7223 VSS.n4064 VSS.n1523 0.193087
R7224 VSS.n5756 VSS.n5752 0.188841
R7225 VSS.n413 VSS.n322 0.188079
R7226 VSS.n1174 VSS.n1171 0.188
R7227 VSS.n239 VSS.n221 0.1865
R7228 VSS.n5185 VSS.n4783 0.1865
R7229 VSS.n351 VSS.n350 0.185092
R7230 VSS.n220 VSS.n219 0.1805
R7231 VSS.n5204 VSS.n5203 0.1805
R7232 VSS.n4551 VSS.n4548 0.174181
R7233 VSS.n5511 VSS.n5508 0.17414
R7234 VSS.n4407 VSS.n4406 0.174137
R7235 VSS.n5303 VSS.n5301 0.172819
R7236 VSS.n83 VSS.n82 0.170926
R7237 VSS.n4120 VSS.n4119 0.169688
R7238 VSS.n21 VSS.n20 0.167572
R7239 VSS.n4311 VSS.n4310 0.164562
R7240 VSS.n3871 VSS.n3870 0.163308
R7241 VSS.n5153 VSS.n5152 0.163136
R7242 VSS.n148 VSS.n147 0.162433
R7243 VSS.n4205 VSS.n4203 0.161214
R7244 VSS.n954 VSS.n952 0.161214
R7245 VSS.n4121 VSS.n4120 0.161214
R7246 VSS.n4134 VSS.n4132 0.161214
R7247 VSS.n497 VSS.n493 0.160198
R7248 VSS.n5780 VSS.n5779 0.159119
R7249 VSS.n5859 VSS.n5858 0.157743
R7250 VSS.n4411 VSS.n4410 0.157329
R7251 VSS.n5308 VSS.n5306 0.15648
R7252 VSS.n5860 VSS.n5859 0.156251
R7253 VSS VSS.n4205 0.155589
R7254 VSS.n5287 VSS.n5282 0.155512
R7255 VSS.n4386 VSS.n4383 0.153637
R7256 VSS.n5151 VSS.n5150 0.153513
R7257 VSS.n4504 VSS.n4503 0.152808
R7258 VSS.n1293 VSS.n1290 0.15275
R7259 VSS.n146 VSS.n145 0.152738
R7260 VSS.n4556 VSS.n4555 0.152674
R7261 VSS.n4091 VSS.n4090 0.151571
R7262 VSS.n4129 VSS.n4127 0.151571
R7263 VSS.n961 VSS.n960 0.150768
R7264 VSS.n5000 VSS.n4994 0.150235
R7265 VSS.n4659 VSS.n4655 0.150235
R7266 VSS.n5019 VSS.n5016 0.148852
R7267 VSS.n5022 VSS.n5019 0.148852
R7268 VSS.n5025 VSS.n5022 0.148852
R7269 VSS.n5028 VSS.n5025 0.148852
R7270 VSS.n5031 VSS.n5028 0.148852
R7271 VSS.n5034 VSS.n5031 0.148852
R7272 VSS.n5037 VSS.n5034 0.148852
R7273 VSS.n5040 VSS.n5037 0.148852
R7274 VSS.n5043 VSS.n5040 0.148852
R7275 VSS.n5478 VSS.n5475 0.148852
R7276 VSS.n5481 VSS.n5478 0.148852
R7277 VSS.n5484 VSS.n5481 0.148852
R7278 VSS.n5487 VSS.n5484 0.148852
R7279 VSS.n5490 VSS.n5487 0.148852
R7280 VSS.n5493 VSS.n5490 0.148852
R7281 VSS.n5496 VSS.n5493 0.148852
R7282 VSS.n5499 VSS.n5496 0.148852
R7283 VSS.n5502 VSS.n5499 0.148852
R7284 VSS.n5505 VSS.n5502 0.148852
R7285 VSS.n4616 VSS.n4613 0.148852
R7286 VSS.n4619 VSS.n4616 0.148852
R7287 VSS.n4622 VSS.n4619 0.148852
R7288 VSS.n4625 VSS.n4622 0.148852
R7289 VSS.n4628 VSS.n4625 0.148852
R7290 VSS.n4631 VSS.n4628 0.148852
R7291 VSS.n4634 VSS.n4631 0.148852
R7292 VSS.n4637 VSS.n4634 0.148852
R7293 VSS.n4640 VSS.n4637 0.148852
R7294 VSS.n4545 VSS.n4542 0.148852
R7295 VSS.n4542 VSS.n4539 0.148852
R7296 VSS.n4539 VSS.n4536 0.148852
R7297 VSS.n4536 VSS.n4533 0.148852
R7298 VSS.n4533 VSS.n4530 0.148852
R7299 VSS.n4530 VSS.n4527 0.148852
R7300 VSS.n4527 VSS.n4524 0.148852
R7301 VSS.n4524 VSS.n4521 0.148852
R7302 VSS.n4521 VSS.n4518 0.148852
R7303 VSS.n4518 VSS.n4515 0.148852
R7304 VSS.n4119 VSS.n919 0.148402
R7305 VSS.n4391 VSS.n4389 0.147239
R7306 VSS.n167 VSS.n164 0.147239
R7307 VSS.n211 VSS.n208 0.147239
R7308 VSS.n214 VSS.n211 0.147239
R7309 VSS.n201 VSS.n198 0.147239
R7310 VSS.n204 VSS.n201 0.147239
R7311 VSS.n116 VSS.n113 0.147239
R7312 VSS.n251 VSS.n247 0.147239
R7313 VSS.n5160 VSS.n5157 0.147239
R7314 VSS.n5224 VSS.n5221 0.147239
R7315 VSS.n5227 VSS.n5224 0.147239
R7316 VSS.n5214 VSS.n5211 0.147239
R7317 VSS.n5217 VSS.n5214 0.147239
R7318 VSS.n4758 VSS.n4755 0.147239
R7319 VSS.n5252 VSS.n5250 0.147239
R7320 VSS.n5246 VSS.n5244 0.147239
R7321 VSS.n4427 VSS.n4424 0.147239
R7322 VSS.n4424 VSS.n4422 0.147239
R7323 VSS.n2883 VSS 0.145448
R7324 VSS.n5416 VSS.n5413 0.144304
R7325 VSS.n4433 VSS.n4430 0.144304
R7326 VSS.n5308 VSS.n5290 0.142348
R7327 VSS.n4414 VSS.n4413 0.142348
R7328 VSS.n4413 VSS.n4411 0.14137
R7329 VSS.n5508 VSS.n5505 0.139951
R7330 VSS.n4548 VSS.n4545 0.139951
R7331 VSS.n1302 VSS.n973 0.139082
R7332 VSS.n5279 VSS.n5278 0.137463
R7333 VSS.n4376 VSS.n4375 0.136472
R7334 VSS.n3739 VSS.n3738 0.133072
R7335 VSS.n290 VSS.n289 0.132286
R7336 VSS.n245 VSS.n244 0.131851
R7337 VSS.n5832 VSS.n5831 0.131118
R7338 VSS.n160 VSS.n157 0.130588
R7339 VSS.n109 VSS.n108 0.130302
R7340 VSS.n5144 VSS.n5141 0.130084
R7341 VSS.n5242 VSS.n5241 0.129374
R7342 VSS.n1374 VSS.n1371 0.12841
R7343 VSS.n1257 VSS.n1254 0.128
R7344 VSS.n5240 VSS.n5239 0.125349
R7345 VSS.n4171 VSS.n4170 0.12483
R7346 VSS.n107 VSS.n106 0.124421
R7347 VSS.n5280 VSS.n5279 0.123458
R7348 VSS.n244 VSS.n243 0.122817
R7349 VSS.n4430 VSS.n4427 0.122783
R7350 VSS.n5256 VSS.n5255 0.122669
R7351 VSS.n4377 VSS.n4376 0.122609
R7352 VSS.n1510 VSS.n1509 0.1225
R7353 VSS.n5304 VSS.n5303 0.12249
R7354 VSS.n5237 VSS.n5236 0.121959
R7355 VSS.n4379 VSS.n4378 0.121915
R7356 VSS.n5306 VSS.n5305 0.121915
R7357 VSS.n5282 VSS.n5281 0.121915
R7358 VSS.n4410 VSS.n4409 0.121915
R7359 VSS.n4381 VSS.n4380 0.121893
R7360 VSS.n106 VSS.n103 0.121804
R7361 VSS.n5239 VSS.n5238 0.121804
R7362 VSS.n4408 VSS.n4407 0.121641
R7363 VSS.n215 VSS.n191 0.120826
R7364 VSS.n4765 VSS.n4761 0.120826
R7365 VSS.n5071 VSS.n5068 0.119969
R7366 VSS.n5128 VSS.n5125 0.119969
R7367 VSS.n5065 VSS.n5063 0.119969
R7368 VSS.n4994 VSS.n4993 0.119969
R7369 VSS.n4989 VSS.n4986 0.119969
R7370 VSS.n4986 VSS.n4982 0.119969
R7371 VSS.n4965 VSS.n4963 0.119969
R7372 VSS.n4959 VSS.n4956 0.119969
R7373 VSS.n4956 VSS.n4952 0.119969
R7374 VSS.n5469 VSS.n5466 0.119969
R7375 VSS.n5472 VSS.n5469 0.119969
R7376 VSS.n4607 VSS.n4604 0.119969
R7377 VSS.n4566 VSS.n4563 0.119969
R7378 VSS.n4568 VSS.n4566 0.119969
R7379 VSS.n4577 VSS.n4574 0.119969
R7380 VSS.n38 VSS.n35 0.119969
R7381 VSS.n44 VSS.n41 0.119969
R7382 VSS.n46 VSS.n44 0.119969
R7383 VSS.n54 VSS.n51 0.119969
R7384 VSS.n56 VSS.n54 0.119969
R7385 VSS.n4679 VSS.n4676 0.119969
R7386 VSS.n4672 VSS.n4668 0.119969
R7387 VSS.n4668 VSS.n4665 0.119969
R7388 VSS.n4662 VSS.n4659 0.119969
R7389 VSS.n120 VSS.n117 0.119848
R7390 VSS.n5208 VSS.n5184 0.119848
R7391 VSS.n4165 VSS.n4164 0.119263
R7392 VSS.n888 VSS.n887 0.119263
R7393 VSS.n4557 VSS.n4554 0.119173
R7394 VSS.n5455 VSS.n5452 0.118921
R7395 VSS.n5452 VSS.n5449 0.118921
R7396 VSS.n5442 VSS.n5439 0.118921
R7397 VSS.n5439 VSS.n5436 0.118921
R7398 VSS.n5436 VSS.n5433 0.118921
R7399 VSS.n5433 VSS.n5430 0.118921
R7400 VSS.n5537 VSS.n5534 0.118921
R7401 VSS.n4446 VSS.n4443 0.118921
R7402 VSS.n4449 VSS.n4446 0.118921
R7403 VSS.n4452 VSS.n4449 0.118921
R7404 VSS.n4455 VSS.n4452 0.118921
R7405 VSS.n4458 VSS.n4455 0.118921
R7406 VSS.n4461 VSS.n4458 0.118921
R7407 VSS.n4464 VSS.n4461 0.118921
R7408 VSS.n4467 VSS.n4464 0.118921
R7409 VSS.n4474 VSS.n4471 0.118921
R7410 VSS.n4477 VSS.n4474 0.118921
R7411 VSS.n4480 VSS.n4477 0.118921
R7412 VSS.n4483 VSS.n4480 0.118921
R7413 VSS.n4486 VSS.n4483 0.118921
R7414 VSS.n108 VSS.n107 0.118335
R7415 VSS.n5241 VSS.n5240 0.118335
R7416 VSS.n4554 VSS.n4551 0.116783
R7417 VSS.n5427 VSS.n5426 0.116553
R7418 VSS.n5419 VSS.n5416 0.115403
R7419 VSS.n5514 VSS.n5513 0.115328
R7420 VSS.n4436 VSS.n4433 0.115214
R7421 VSS.n1340 VSS.n1338 0.113945
R7422 VSS.n1338 VSS.n1336 0.113945
R7423 VSS.n1332 VSS.n1330 0.113945
R7424 VSS.n1330 VSS.n1326 0.113945
R7425 VSS.n1326 VSS.n1324 0.113945
R7426 VSS.n1324 VSS.n1320 0.113945
R7427 VSS.n1320 VSS.n1316 0.113945
R7428 VSS.n1316 VSS.n1313 0.113945
R7429 VSS.n1308 VSS.n1307 0.113945
R7430 VSS.n1307 VSS.n1304 0.113945
R7431 VSS.n1377 VSS.n1374 0.113945
R7432 VSS.n1380 VSS.n1377 0.113945
R7433 VSS.n1384 VSS.n1380 0.113945
R7434 VSS.n1387 VSS.n1384 0.113945
R7435 VSS.n1391 VSS.n1387 0.113945
R7436 VSS.n4099 VSS.n4096 0.113945
R7437 VSS.n1301 VSS.n1297 0.113933
R7438 VSS.n5513 VSS.n5511 0.113776
R7439 VSS.n5066 VSS.n5065 0.113597
R7440 VSS.n874 VSS.n873 0.113103
R7441 VSS.n1290 VSS.n1288 0.113
R7442 VSS.n1297 VSS.n1293 0.113
R7443 VSS.n687 VSS.n685 0.113
R7444 VSS.n1259 VSS.n1257 0.113
R7445 VSS.n1262 VSS.n1259 0.113
R7446 VSS.n1265 VSS.n1262 0.113
R7447 VSS.n1268 VSS.n1265 0.113
R7448 VSS.n1271 VSS.n1268 0.113
R7449 VSS.n1274 VSS.n1271 0.113
R7450 VSS.n1277 VSS.n1274 0.113
R7451 VSS.n1280 VSS.n1277 0.113
R7452 VSS.n1283 VSS.n1280 0.113
R7453 VSS.n1178 VSS.n1174 0.113
R7454 VSS.n1181 VSS.n1178 0.113
R7455 VSS.n1184 VSS.n1181 0.113
R7456 VSS.n1187 VSS.n1184 0.113
R7457 VSS.n1190 VSS.n1187 0.113
R7458 VSS.n1193 VSS.n1190 0.113
R7459 VSS.n1196 VSS.n1193 0.113
R7460 VSS.n1199 VSS.n1196 0.113
R7461 VSS.n1203 VSS.n1199 0.113
R7462 VSS.n1206 VSS.n1203 0.113
R7463 VSS.n1209 VSS.n1206 0.113
R7464 VSS.n1212 VSS.n1209 0.113
R7465 VSS.n1215 VSS.n1212 0.113
R7466 VSS.n1218 VSS.n1215 0.113
R7467 VSS.n1221 VSS.n1218 0.113
R7468 VSS.n1224 VSS.n1221 0.113
R7469 VSS.n1228 VSS.n1224 0.113
R7470 VSS.n1231 VSS.n1228 0.113
R7471 VSS.n1234 VSS.n1231 0.113
R7472 VSS.n1237 VSS.n1234 0.113
R7473 VSS.n1240 VSS.n1237 0.113
R7474 VSS.n1243 VSS.n1240 0.113
R7475 VSS.n1246 VSS.n1243 0.113
R7476 VSS.n1249 VSS.n1246 0.113
R7477 VSS.n1251 VSS.n1249 0.113
R7478 VSS.n1254 VSS.n1251 0.113
R7479 VSS.n1345 VSS.n1342 0.113
R7480 VSS.n1347 VSS.n1345 0.113
R7481 VSS.n1350 VSS.n1347 0.113
R7482 VSS.n1352 VSS.n1350 0.113
R7483 VSS.n1355 VSS.n1352 0.113
R7484 VSS.n1357 VSS.n1355 0.113
R7485 VSS.n1360 VSS.n1357 0.113
R7486 VSS.n1362 VSS.n1360 0.113
R7487 VSS.n1365 VSS.n1362 0.113
R7488 VSS.n1367 VSS.n1365 0.113
R7489 VSS.n1371 VSS.n1367 0.113
R7490 VSS.n1164 VSS.n1161 0.112367
R7491 VSS.n5805 VSS.n5773 0.112006
R7492 VSS.n4414 VSS.n4379 0.111845
R7493 VSS.n4383 VSS.n4382 0.111448
R7494 VSS.n5258 VSS.n5257 0.111448
R7495 VSS.n491 VSS.n487 0.111156
R7496 VSS.n493 VSS.n491 0.111156
R7497 VSS.n487 VSS.n485 0.11043
R7498 VSS.n763 VSS.n760 0.110256
R7499 VSS.n760 VSS.n757 0.110256
R7500 VSS.n757 VSS.n754 0.110256
R7501 VSS.n4070 VSS.n4067 0.110256
R7502 VSS.n4083 VSS.n4070 0.110256
R7503 VSS.n4083 VSS.n4082 0.110256
R7504 VSS.n4082 VSS.n4079 0.110256
R7505 VSS.n4079 VSS.n4076 0.110256
R7506 VSS.n4076 VSS.n4073 0.110256
R7507 VSS.n366 VSS.n362 0.110256
R7508 VSS.n368 VSS.n366 0.110256
R7509 VSS.n371 VSS.n368 0.110256
R7510 VSS.n374 VSS.n371 0.110256
R7511 VSS.n377 VSS.n374 0.110256
R7512 VSS.n380 VSS.n377 0.110256
R7513 VSS.n383 VSS.n380 0.110256
R7514 VSS.n386 VSS.n383 0.110256
R7515 VSS.n389 VSS.n386 0.110256
R7516 VSS.n393 VSS.n389 0.110256
R7517 VSS.n396 VSS.n393 0.110256
R7518 VSS.n399 VSS.n396 0.110256
R7519 VSS.n402 VSS.n399 0.110256
R7520 VSS.n405 VSS.n402 0.110256
R7521 VSS.n412 VSS.n409 0.110256
R7522 VSS.n419 VSS.n416 0.110256
R7523 VSS.n422 VSS.n419 0.110256
R7524 VSS.n427 VSS.n422 0.110256
R7525 VSS.n430 VSS.n427 0.110256
R7526 VSS.n433 VSS.n430 0.110256
R7527 VSS.n436 VSS.n433 0.110256
R7528 VSS.n439 VSS.n436 0.110256
R7529 VSS.n442 VSS.n439 0.110256
R7530 VSS.n445 VSS.n442 0.110256
R7531 VSS.n448 VSS.n445 0.110256
R7532 VSS.n451 VSS.n448 0.110256
R7533 VSS.n454 VSS.n451 0.110256
R7534 VSS.n458 VSS.n454 0.110256
R7535 VSS.n461 VSS.n458 0.110256
R7536 VSS.n464 VSS.n461 0.110256
R7537 VSS.n473 VSS.n464 0.110256
R7538 VSS.n476 VSS.n473 0.110256
R7539 VSS.n479 VSS.n476 0.110256
R7540 VSS.n482 VSS.n479 0.110256
R7541 VSS.n485 VSS.n482 0.110256
R7542 VSS.n1534 VSS.n1531 0.110256
R7543 VSS.n1531 VSS.n1528 0.110256
R7544 VSS.n4037 VSS.n4034 0.110256
R7545 VSS.n3976 VSS.n3973 0.110256
R7546 VSS.n3973 VSS.n3970 0.110256
R7547 VSS.n3970 VSS.n3967 0.110256
R7548 VSS.n3967 VSS.n3964 0.110256
R7549 VSS.n3964 VSS.n3961 0.110256
R7550 VSS.n3961 VSS.n3958 0.110256
R7551 VSS.n3958 VSS.n3955 0.110256
R7552 VSS.n3955 VSS.n3952 0.110256
R7553 VSS.n3952 VSS.n3949 0.110256
R7554 VSS.n3949 VSS.n3946 0.110256
R7555 VSS.n3946 VSS.n3943 0.110256
R7556 VSS.n3943 VSS.n3940 0.110256
R7557 VSS.n3940 VSS.n3937 0.110256
R7558 VSS.n3937 VSS.n3934 0.110256
R7559 VSS.n3934 VSS.n3930 0.110256
R7560 VSS.n3930 VSS.n3927 0.110256
R7561 VSS.n3927 VSS.n3924 0.110256
R7562 VSS.n3924 VSS.n3921 0.110256
R7563 VSS.n3921 VSS.n3918 0.110256
R7564 VSS.n4046 VSS.n4042 0.110256
R7565 VSS.n4049 VSS.n4046 0.110256
R7566 VSS.n4057 VSS.n4053 0.110256
R7567 VSS.n4060 VSS.n4057 0.110256
R7568 VSS.n4063 VSS.n4060 0.110256
R7569 VSS.n728 VSS.n725 0.110256
R7570 VSS.n725 VSS.n722 0.110256
R7571 VSS.n722 VSS.n719 0.110256
R7572 VSS.n4280 VSS.n4278 0.110256
R7573 VSS.n4283 VSS.n4280 0.110256
R7574 VSS.n4286 VSS.n4283 0.110256
R7575 VSS.n4298 VSS.n4295 0.110256
R7576 VSS.n4295 VSS.n4292 0.110256
R7577 VSS.n4292 VSS.n4289 0.110256
R7578 VSS.n907 VSS.n905 0.110256
R7579 VSS.n905 VSS.n902 0.110256
R7580 VSS.n902 VSS.n899 0.110256
R7581 VSS.n899 VSS.n897 0.110256
R7582 VSS.n897 VSS.n895 0.110256
R7583 VSS.n895 VSS.n893 0.110256
R7584 VSS.n4226 VSS.n4223 0.110256
R7585 VSS.n4229 VSS.n4226 0.110256
R7586 VSS.n4232 VSS.n4229 0.110256
R7587 VSS.n4234 VSS.n4232 0.110256
R7588 VSS.n4237 VSS.n4234 0.110256
R7589 VSS.n4241 VSS.n4237 0.110256
R7590 VSS.n4244 VSS.n4241 0.110256
R7591 VSS.n4247 VSS.n4244 0.110256
R7592 VSS.n4251 VSS.n4247 0.110256
R7593 VSS.n4258 VSS.n4255 0.110256
R7594 VSS.n4261 VSS.n4258 0.110256
R7595 VSS.n4264 VSS.n4261 0.110256
R7596 VSS.n4267 VSS.n4264 0.110256
R7597 VSS.n4270 VSS.n4267 0.110256
R7598 VSS.n5781 VSS.n5780 0.110211
R7599 VSS.n243 VSS.n242 0.109357
R7600 VSS.n5236 VSS.n5235 0.109357
R7601 VSS.n6037 VSS 0.109087
R7602 VSS.n5259 VSS.n5258 0.108345
R7603 VSS.n5305 VSS.n5304 0.10833
R7604 VSS.n5281 VSS.n5280 0.10833
R7605 VSS.n4378 VSS.n4377 0.10833
R7606 VSS.n4409 VSS.n4408 0.10833
R7607 VSS.n4492 VSS.n4489 0.108109
R7608 VSS.n5520 VSS.n5517 0.108109
R7609 VSS.n4050 VSS.n4049 0.108061
R7610 VSS.n498 VSS.n497 0.108061
R7611 VSS.n1336 VSS.n1333 0.107895
R7612 VSS.n5287 VSS.n5286 0.10713
R7613 VSS.n5446 VSS.n5443 0.107079
R7614 VSS VSS.n358 0.107055
R7615 VSS.n4973 VSS.n4970 0.106429
R7616 VSS.n4299 VSS.n4298 0.105134
R7617 VSS.n5422 VSS.n5419 0.104711
R7618 VSS.n4439 VSS.n4436 0.104711
R7619 VSS.n252 VSS.n251 0.104196
R7620 VSS.n5250 VSS.n5247 0.104196
R7621 VSS.n5103 VSS.n5101 0.10383
R7622 VSS.n4596 VSS.n4593 0.103507
R7623 VSS.n5873 VSS 0.10345
R7624 VSS.n4610 VSS.n4608 0.103243
R7625 VSS.n5138 VSS.n5135 0.103217
R7626 VSS.n154 VSS.n151 0.103217
R7627 VSS.n4118 VSS.n4099 0.102601
R7628 VSS.n5129 VSS.n5045 0.102447
R7629 VSS.n4969 VSS.n4966 0.102447
R7630 VSS.n5135 VSS.n5132 0.102239
R7631 VSS.n5141 VSS.n5138 0.102239
R7632 VSS.n157 VSS.n154 0.102239
R7633 VSS.n151 VSS.n62 0.102239
R7634 VSS.n3846 VSS.n3845 0.100173
R7635 VSS.n187 VSS.n184 0.0999444
R7636 VSS.n240 VSS.n123 0.0999444
R7637 VSS.n5180 VSS.n5177 0.0999444
R7638 VSS.n5232 VSS.n5231 0.0999444
R7639 VSS VSS.n5816 0.0997784
R7640 VSS VSS.n5865 0.0997784
R7641 VSS.n5893 VSS 0.0997784
R7642 VSS VSS.n5763 0.0997784
R7643 VSS.n4584 VSS.n4581 0.0992611
R7644 VSS.n4382 VSS.n4381 0.0990345
R7645 VSS.n5257 VSS.n5256 0.0990345
R7646 VSS.n96 VSS.n95 0.0986818
R7647 VSS.n5078 VSS.n5075 0.0984646
R7648 VSS.n5066 VSS.n5059 0.0978681
R7649 VSS.n5006 VSS.n5003 0.0974231
R7650 VSS.n5013 VSS.n5010 0.0974231
R7651 VSS.n5016 VSS.n5013 0.0974231
R7652 VSS.n4643 VSS.n4640 0.0974231
R7653 VSS.n4646 VSS.n4643 0.0974231
R7654 VSS.n4652 VSS.n4649 0.0974231
R7655 VSS.n5410 VSS.n5409 0.0973478
R7656 VSS.n1165 VSS.n1164 0.0968905
R7657 VSS.n5010 VSS.n5006 0.0964341
R7658 VSS.n4649 VSS.n4646 0.0964341
R7659 VSS.n5290 VSS.n5287 0.0963696
R7660 VSS.n3915 VSS.n1534 0.0956219
R7661 VSS.n4963 VSS.n4960 0.0952788
R7662 VSS.n51 VSS.n47 0.0952788
R7663 VSS.n5054 VSS.n5053 0.0945909
R7664 VSS VSS.n5885 0.0945618
R7665 VSS.n5253 VSS.n5237 0.0945541
R7666 VSS.n4496 VSS.n4492 0.0942929
R7667 VSS.n5523 VSS.n5520 0.0941041
R7668 VSS.n4119 VSS.n4118 0.09365
R7669 VSS.n5235 VSS.n5234 0.0922143
R7670 VSS.n4560 VSS.n4559 0.0920929
R7671 VSS.n1031 VSS.n1030 0.0914091
R7672 VSS VSS.n0 0.0914091
R7673 VSS VSS.n6068 0.0914091
R7674 VSS.n6068 VSS.n6067 0.0914091
R7675 VSS.n6067 VSS.n6066 0.0914091
R7676 VSS.n6062 VSS.n6061 0.0914091
R7677 VSS.n242 VSS.n241 0.0913571
R7678 VSS.n1284 VSS.n1283 0.09125
R7679 VSS.n1024 VSS.n1012 0.0909545
R7680 VSS.n321 VSS.n320 0.0907679
R7681 VSS.n252 VSS.n109 0.0905
R7682 VSS.n5247 VSS.n5242 0.0905
R7683 VSS.n4978 VSS.n4977 0.0905
R7684 VSS.n4419 VSS.n4418 0.0905
R7685 VSS.n4676 VSS.n4673 0.0905
R7686 VSS.n4073 VSS.n908 0.0897683
R7687 VSS.n4042 VSS.n4040 0.0897683
R7688 VSS.n5132 VSS.n5129 0.0895217
R7689 VSS.n5123 VSS.n5122 0.0889071
R7690 VSS.n4608 VSS.n62 0.0885435
R7691 VSS.n4600 VSS.n4599 0.0881106
R7692 VSS.n5834 VSS.n5833 0.0877209
R7693 VSS.n5526 VSS.n5523 0.0873421
R7694 VSS.n4499 VSS.n4496 0.0873421
R7695 VSS.n1452 VSS.n1451 0.0862944
R7696 VSS.n1449 VSS.n1448 0.0862944
R7697 VSS.n5362 VSS.n5359 0.0854057
R7698 VSS.n5365 VSS.n5362 0.0854057
R7699 VSS.n5368 VSS.n5365 0.0854057
R7700 VSS.n5371 VSS.n5368 0.0854057
R7701 VSS.n5374 VSS.n5371 0.0854057
R7702 VSS.n5377 VSS.n5374 0.0854057
R7703 VSS.n5380 VSS.n5377 0.0854057
R7704 VSS.n5383 VSS.n5380 0.0854057
R7705 VSS.n5386 VSS.n5383 0.0854057
R7706 VSS.n5389 VSS.n5386 0.0854057
R7707 VSS.n5392 VSS.n5389 0.0854057
R7708 VSS.n5395 VSS.n5392 0.0854057
R7709 VSS.n5398 VSS.n5395 0.0854057
R7710 VSS.n5401 VSS.n5398 0.0854057
R7711 VSS.n5545 VSS.n5542 0.0854057
R7712 VSS.n5548 VSS.n5545 0.0854057
R7713 VSS.n5551 VSS.n5548 0.0854057
R7714 VSS.n5554 VSS.n5551 0.0854057
R7715 VSS.n5561 VSS.n5558 0.0854057
R7716 VSS.n5564 VSS.n5561 0.0854057
R7717 VSS.n5567 VSS.n5564 0.0854057
R7718 VSS.n5569 VSS.n5567 0.0854057
R7719 VSS.n5577 VSS.n5573 0.0854057
R7720 VSS.n5580 VSS.n5577 0.0854057
R7721 VSS.n5583 VSS.n5580 0.0854057
R7722 VSS.n5586 VSS.n5583 0.0854057
R7723 VSS.n5589 VSS.n5586 0.0854057
R7724 VSS.n5596 VSS.n5593 0.0854057
R7725 VSS.n5599 VSS.n5596 0.0854057
R7726 VSS.n1032 VSS.n1031 0.0850455
R7727 VSS.n4360 VSS.n4358 0.0846795
R7728 VSS.n5262 VSS.n5259 0.0846304
R7729 VSS.n5359 VSS.n5356 0.0843639
R7730 VSS.n4559 VSS.n4557 0.0841283
R7731 VSS.n39 VSS.n38 0.0841283
R7732 VSS.n5095 VSS.n5078 0.0838349
R7733 VSS.n4760 VSS.n4759 0.0838333
R7734 VSS.n5098 VSS.n5097 0.0837469
R7735 VSS.n4589 VSS.n4588 0.0832732
R7736 VSS.n5463 VSS.n5459 0.0832014
R7737 VSS.n5356 VSS.n5353 0.0830864
R7738 VSS VSS.n5861 0.083054
R7739 VSS.n4585 VSS.n4584 0.0830384
R7740 VSS.n4345 VSS.n4343 0.0828171
R7741 VSS.n1161 VSS.n1158 0.0828171
R7742 VSS.n1158 VSS.n1155 0.0828171
R7743 VSS.n1155 VSS.n1152 0.0828171
R7744 VSS.n1152 VSS.n1149 0.0828171
R7745 VSS.n1149 VSS.n1146 0.0828171
R7746 VSS.n1146 VSS.n1143 0.0828171
R7747 VSS.n1143 VSS.n1140 0.0828171
R7748 VSS.n1140 VSS.n1137 0.0828171
R7749 VSS.n1137 VSS.n1134 0.0828171
R7750 VSS.n1134 VSS.n1131 0.0828171
R7751 VSS.n1131 VSS.n1128 0.0828171
R7752 VSS.n1128 VSS.n1125 0.0828171
R7753 VSS.n1125 VSS.n1122 0.0828171
R7754 VSS.n1122 VSS.n1119 0.0828171
R7755 VSS.n1119 VSS.n1116 0.0828171
R7756 VSS.n1116 VSS.n1113 0.0828171
R7757 VSS.n1113 VSS.n1110 0.0828171
R7758 VSS.n1110 VSS.n1107 0.0828171
R7759 VSS.n1107 VSS.n1104 0.0828171
R7760 VSS.n1104 VSS.n1101 0.0828171
R7761 VSS.n1101 VSS.n1098 0.0828171
R7762 VSS.n1098 VSS.n1095 0.0828171
R7763 VSS.n1095 VSS.n1092 0.0828171
R7764 VSS.n1092 VSS.n1089 0.0828171
R7765 VSS.n1089 VSS.n1086 0.0828171
R7766 VSS.n1086 VSS.n1083 0.0828171
R7767 VSS.n1083 VSS.n1080 0.0828171
R7768 VSS.n1080 VSS.n1076 0.0828171
R7769 VSS.n1076 VSS.n1073 0.0828171
R7770 VSS.n1073 VSS.n1070 0.0828171
R7771 VSS.n1070 VSS.n1067 0.0828171
R7772 VSS.n1067 VSS.n1064 0.0828171
R7773 VSS.n1064 VSS.n1061 0.0828171
R7774 VSS.n1061 VSS.n1058 0.0828171
R7775 VSS.n1058 VSS.n1055 0.0828171
R7776 VSS.n1055 VSS.n1052 0.0828171
R7777 VSS.n1052 VSS.n1049 0.0828171
R7778 VSS.n1049 VSS.n1046 0.0828171
R7779 VSS.n1046 VSS.n1043 0.0828171
R7780 VSS.n1043 VSS.n1040 0.0828171
R7781 VSS.n1040 VSS.n1037 0.0828171
R7782 VSS.n713 VSS.n710 0.0828171
R7783 VSS.n710 VSS.n707 0.0828171
R7784 VSS.n707 VSS.n704 0.0828171
R7785 VSS.n700 VSS.n697 0.0828171
R7786 VSS.n697 VSS.n694 0.0828171
R7787 VSS.n691 VSS.n687 0.0828171
R7788 VSS.n685 VSS.n681 0.0828171
R7789 VSS.n681 VSS.n678 0.0828171
R7790 VSS.n678 VSS.n675 0.0828171
R7791 VSS.n675 VSS.n673 0.0828171
R7792 VSS.n673 VSS.n670 0.0828171
R7793 VSS.n670 VSS.n667 0.0828171
R7794 VSS.n667 VSS.n664 0.0828171
R7795 VSS.n664 VSS.n661 0.0828171
R7796 VSS.n661 VSS.n658 0.0828171
R7797 VSS.n658 VSS.n655 0.0828171
R7798 VSS.n655 VSS.n652 0.0828171
R7799 VSS.n652 VSS.n649 0.0828171
R7800 VSS.n649 VSS.n646 0.0828171
R7801 VSS.n646 VSS.n643 0.0828171
R7802 VSS.n643 VSS.n640 0.0828171
R7803 VSS.n640 VSS.n637 0.0828171
R7804 VSS.n637 VSS.n634 0.0828171
R7805 VSS.n634 VSS.n631 0.0828171
R7806 VSS.n631 VSS.n628 0.0828171
R7807 VSS.n628 VSS.n625 0.0828171
R7808 VSS.n625 VSS.n622 0.0828171
R7809 VSS.n622 VSS.n619 0.0828171
R7810 VSS.n619 VSS.n616 0.0828171
R7811 VSS.n616 VSS.n613 0.0828171
R7812 VSS.n613 VSS.n610 0.0828171
R7813 VSS.n610 VSS.n607 0.0828171
R7814 VSS.n607 VSS.n604 0.0828171
R7815 VSS.n604 VSS.n601 0.0828171
R7816 VSS.n601 VSS.n598 0.0828171
R7817 VSS.n598 VSS.n595 0.0828171
R7818 VSS.n595 VSS.n593 0.0828171
R7819 VSS.n593 VSS.n589 0.0828171
R7820 VSS.n589 VSS.n586 0.0828171
R7821 VSS.n586 VSS.n583 0.0828171
R7822 VSS.n583 VSS.n580 0.0828171
R7823 VSS.n580 VSS.n577 0.0828171
R7824 VSS.n577 VSS.n574 0.0828171
R7825 VSS.n574 VSS.n571 0.0828171
R7826 VSS.n571 VSS.n566 0.0828171
R7827 VSS.n566 VSS.n562 0.0828171
R7828 VSS.n562 VSS.n559 0.0828171
R7829 VSS.n559 VSS.n556 0.0828171
R7830 VSS.n556 VSS.n554 0.0828171
R7831 VSS.n554 VSS.n551 0.0828171
R7832 VSS.n551 VSS.n548 0.0828171
R7833 VSS.n548 VSS.n545 0.0828171
R7834 VSS.n545 VSS.n542 0.0828171
R7835 VSS.n542 VSS.n539 0.0828171
R7836 VSS.n539 VSS.n536 0.0828171
R7837 VSS.n536 VSS.n533 0.0828171
R7838 VSS.n533 VSS.n530 0.0828171
R7839 VSS.n530 VSS.n526 0.0828171
R7840 VSS.n526 VSS.n523 0.0828171
R7841 VSS.n523 VSS.n520 0.0828171
R7842 VSS.n520 VSS.n517 0.0828171
R7843 VSS.n517 VSS.n514 0.0828171
R7844 VSS.n5321 VSS.n5317 0.0828171
R7845 VSS.n5324 VSS.n5321 0.0828171
R7846 VSS.n5326 VSS.n5324 0.0828171
R7847 VSS.n5329 VSS.n5326 0.0828171
R7848 VSS.n5332 VSS.n5329 0.0828171
R7849 VSS.n5336 VSS.n5332 0.0828171
R7850 VSS.n5341 VSS.n5336 0.0828171
R7851 VSS.n5344 VSS.n5341 0.0828171
R7852 VSS.n5347 VSS.n5344 0.0828171
R7853 VSS.n5350 VSS.n5347 0.0828171
R7854 VSS.n5353 VSS.n5350 0.0828171
R7855 VSS.n787 VSS.n784 0.0828171
R7856 VSS.n784 VSS.n781 0.0828171
R7857 VSS.n781 VSS.n778 0.0828171
R7858 VSS.n778 VSS.n775 0.0828171
R7859 VSS.n751 VSS.n748 0.0828171
R7860 VSS.n748 VSS.n745 0.0828171
R7861 VSS.n745 VSS.n742 0.0828171
R7862 VSS.n742 VSS.n739 0.0828171
R7863 VSS.n992 VSS.n988 0.0828171
R7864 VSS.n988 VSS.n985 0.0828171
R7865 VSS.n985 VSS.n983 0.0828171
R7866 VSS.n983 VSS.n980 0.0828171
R7867 VSS.n980 VSS.n976 0.0828171
R7868 VSS.n976 VSS.n99 0.0828171
R7869 VSS.n4354 VSS.n4351 0.0828171
R7870 VSS.n4351 VSS.n4349 0.0828171
R7871 VSS.n4349 VSS.n4345 0.0828171
R7872 VSS.n4343 VSS.n4340 0.0828171
R7873 VSS.n4340 VSS.n4337 0.0828171
R7874 VSS.n4334 VSS.n4330 0.0828171
R7875 VSS.n4327 VSS.n4324 0.0828171
R7876 VSS.n4324 VSS.n4321 0.0828171
R7877 VSS.n4321 VSS.n4319 0.0828171
R7878 VSS.n4319 VSS.n4315 0.0828171
R7879 VSS.n1008 VSS.n1005 0.0828171
R7880 VSS.n1005 VSS.n1002 0.0828171
R7881 VSS.n1002 VSS.n998 0.0828171
R7882 VSS.n998 VSS.n995 0.0828171
R7883 VSS.n15 VSS.n5 0.0828171
R7884 VSS.n15 VSS.n14 0.0828171
R7885 VSS.n14 VSS.n11 0.0828171
R7886 VSS.n11 VSS.n8 0.0828171
R7887 VSS.n6053 VSS.n6052 0.0828171
R7888 VSS.n6052 VSS.n6049 0.0828171
R7889 VSS.n6049 VSS.n6046 0.0828171
R7890 VSS.n6046 VSS.n6043 0.0828171
R7891 VSS.n6043 VSS.n6040 0.0828171
R7892 VSS.n6036 VSS.n6032 0.0828171
R7893 VSS.n6032 VSS.n6029 0.0828171
R7894 VSS.n6029 VSS.n6025 0.0828171
R7895 VSS.n6025 VSS.n6022 0.0828171
R7896 VSS.n6022 VSS.n6019 0.0828171
R7897 VSS.n6019 VSS.n6015 0.0828171
R7898 VSS.n6015 VSS.n6012 0.0828171
R7899 VSS.n6012 VSS.n6009 0.0828171
R7900 VSS.n6009 VSS.n6006 0.0828171
R7901 VSS.n6006 VSS.n6003 0.0828171
R7902 VSS.n6003 VSS.n6000 0.0828171
R7903 VSS.n6000 VSS.n5997 0.0828171
R7904 VSS.n5997 VSS.n5994 0.0828171
R7905 VSS.n5994 VSS.n5991 0.0828171
R7906 VSS.n5991 VSS.n5988 0.0828171
R7907 VSS.n5988 VSS.n5985 0.0828171
R7908 VSS.n5985 VSS.n5982 0.0828171
R7909 VSS.n5982 VSS.n5979 0.0828171
R7910 VSS.n5979 VSS.n5976 0.0828171
R7911 VSS.n5976 VSS.n5973 0.0828171
R7912 VSS.n5973 VSS.n5969 0.0828171
R7913 VSS.n5969 VSS.n5966 0.0828171
R7914 VSS.n5966 VSS.n5963 0.0828171
R7915 VSS.n5963 VSS.n5960 0.0828171
R7916 VSS.n5960 VSS.n5957 0.0828171
R7917 VSS.n5957 VSS.n5954 0.0828171
R7918 VSS.n5954 VSS.n5950 0.0828171
R7919 VSS.n5950 VSS.n5947 0.0828171
R7920 VSS.n5947 VSS.n5943 0.0828171
R7921 VSS.n5943 VSS.n5940 0.0828171
R7922 VSS.n5940 VSS.n5937 0.0828171
R7923 VSS.n5937 VSS.n5934 0.0828171
R7924 VSS.n5934 VSS.n5931 0.0828171
R7925 VSS.n5931 VSS.n5928 0.0828171
R7926 VSS.n5928 VSS.n5925 0.0828171
R7927 VSS.n5925 VSS.n5922 0.0828171
R7928 VSS.n5922 VSS.n5919 0.0828171
R7929 VSS.n5919 VSS.n5916 0.0828171
R7930 VSS.n5916 VSS.n5913 0.0828171
R7931 VSS.n5913 VSS.n5910 0.0828171
R7932 VSS.n5910 VSS.n5907 0.0828171
R7933 VSS.n5907 VSS.n5904 0.0828171
R7934 VSS.n5904 VSS.n5901 0.0828171
R7935 VSS.n4749 VSS.n4740 0.0828171
R7936 VSS.n4752 VSS.n4749 0.0828171
R7937 VSS.n5714 VSS.n4752 0.0828171
R7938 VSS.n5714 VSS.n5713 0.0828171
R7939 VSS.n5713 VSS.n5710 0.0828171
R7940 VSS.n5710 VSS.n5707 0.0828171
R7941 VSS.n5707 VSS.n5704 0.0828171
R7942 VSS.n5704 VSS.n5701 0.0828171
R7943 VSS.n5701 VSS.n5698 0.0828171
R7944 VSS.n5698 VSS.n5695 0.0828171
R7945 VSS.n5695 VSS.n5691 0.0828171
R7946 VSS.n5691 VSS.n5688 0.0828171
R7947 VSS.n5688 VSS.n5685 0.0828171
R7948 VSS.n5685 VSS.n5682 0.0828171
R7949 VSS.n5682 VSS.n5679 0.0828171
R7950 VSS.n5679 VSS.n5676 0.0828171
R7951 VSS.n5676 VSS.n5673 0.0828171
R7952 VSS.n5673 VSS.n5670 0.0828171
R7953 VSS.n5670 VSS.n5663 0.0828171
R7954 VSS.n5663 VSS.n5660 0.0828171
R7955 VSS.n5660 VSS.n5655 0.0828171
R7956 VSS.n5655 VSS.n5652 0.0828171
R7957 VSS.n5652 VSS.n5650 0.0828171
R7958 VSS.n5646 VSS.n5643 0.0828171
R7959 VSS.n5643 VSS.n5641 0.0828171
R7960 VSS.n5641 VSS.n5638 0.0828171
R7961 VSS.n5638 VSS.n5636 0.0828171
R7962 VSS.n5632 VSS.n5630 0.0828171
R7963 VSS.n5630 VSS.n5627 0.0828171
R7964 VSS.n5627 VSS.n5624 0.0828171
R7965 VSS.n5624 VSS.n5622 0.0828171
R7966 VSS.n5622 VSS.n5619 0.0828171
R7967 VSS.n5615 VSS.n5612 0.0828171
R7968 VSS.n5612 VSS.n5609 0.0828171
R7969 VSS.n5609 VSS.n5607 0.0828171
R7970 VSS.n5607 VSS.n5605 0.0828171
R7971 VSS.n5409 VSS.n5406 0.0826739
R7972 VSS.n4599 VSS.n4597 0.082242
R7973 VSS.n704 VSS.n701 0.0817195
R7974 VSS.n188 VSS.n167 0.0816957
R7975 VSS.n271 VSS.n270 0.0816607
R7976 VSS.n4872 VSS.n4871 0.0815383
R7977 VSS.n5122 VSS.n5116 0.0814455
R7978 VSS.n6040 VSS.n6037 0.0811707
R7979 VSS.n5072 VSS.n5071 0.0809425
R7980 VSS.n955 VSS.n954 0.0808571
R7981 VSS.n4132 VSS.n4130 0.0808571
R7982 VSS.n4219 VSS.n4207 0.0808571
R7983 VSS.n5181 VSS.n5160 0.0807174
R7984 VSS.n4328 VSS 0.0803113
R7985 VSS.n4500 VSS.n4499 0.0802368
R7986 VSS.n4578 VSS.n4577 0.080146
R7987 VSS.n307 VSS.n306 0.079766
R7988 VSS.n5531 VSS.n5526 0.0794474
R7989 VSS.n313 VSS.n312 0.0794283
R7990 VSS VSS.n950 0.07925
R7991 VSS.n4040 VSS.n4037 0.0787927
R7992 VSS.n5896 VSS.n4740 0.0784268
R7993 VSS.n4990 VSS.n4989 0.0777566
R7994 VSS.n4064 VSS.n4063 0.0773293
R7995 VSS.n5088 VSS.n5087 0.0770957
R7996 VSS.n5538 VSS.n5455 0.077079
R7997 VSS.n4665 VSS.n4663 0.0769602
R7998 VSS.n5570 VSS.n5569 0.0769151
R7999 VSS.n5462 VSS.n5460 0.076587
R8000 VSS.n4328 VSS.n4327 0.0762317
R8001 VSS.n4092 VSS 0.0760357
R8002 VSS.n4130 VSS 0.0760357
R8003 VSS.n908 VSS.n907 0.0758658
R8004 VSS.n5221 VSS.n5218 0.0758261
R8005 VSS.n1333 VSS.n938 0.0755
R8006 VSS VSS.n955 0.0752321
R8007 VSS.n882 VSS.n879 0.0752
R8008 VSS.n205 VSS.n204 0.0748478
R8009 VSS.n5605 VSS.n5602 0.0745854
R8010 VSS VSS.n5446 0.0739211
R8011 VSS.n5253 VSS.n5252 0.0738696
R8012 VSS VSS.n4467 0.0731316
R8013 VSS.n276 VSS.n275 0.0728214
R8014 VSS.n4680 VSS.n57 0.0721814
R8015 VSS.n1304 VSS.n1302 0.0715924
R8016 VSS.n4574 VSS.n4570 0.071385
R8017 VSS.n5802 VSS 0.0710963
R8018 VSS.n6064 VSS.n6063 0.0709545
R8019 VSS.n4974 VSS.n4973 0.0705885
R8020 VSS.n337 VSS.n333 0.0704107
R8021 VSS.n360 VSS.n359 0.0704107
R8022 VSS.n4219 VSS.n4218 0.0704107
R8023 VSS.n3977 VSS.n3976 0.0700122
R8024 VSS.n4299 VSS.n4286 0.0700122
R8025 VSS.n5616 VSS.n5615 0.0696463
R8026 VSS.n4507 VSS.n4506 0.0687418
R8027 VSS.n5058 VSS.n5057 0.0687418
R8028 VSS.n4118 VSS.n1340 0.0685672
R8029 VSS.n3918 VSS.n3915 0.0685488
R8030 VSS.n5636 VSS.n5633 0.0685488
R8031 VSS.n5872 VSS.n5862 0.068
R8032 VSS.n5876 VSS.n5875 0.068
R8033 VSS.n5801 VSS.n5797 0.068
R8034 VSS.n5806 VSS.n5772 0.068
R8035 VSS.n1309 VSS.n1308 0.0678109
R8036 VSS.n5538 VSS.n5537 0.0676053
R8037 VSS.n75 VSS.n66 0.0675213
R8038 VSS.n5115 VSS.n5106 0.0675213
R8039 VSS.n5423 VSS.n5422 0.0673304
R8040 VSS.n4440 VSS.n4439 0.067297
R8041 VSS.n5517 VSS.n5514 0.0670217
R8042 VSS.n85 VSS.n84 0.0666326
R8043 VSS.n5093 VSS.n5092 0.0661354
R8044 VSS.n5795 VSS.n5794 0.066046
R8045 VSS.n4093 VSS.n4092 0.0656429
R8046 VSS.n4278 VSS.n4276 0.0656219
R8047 VSS.n5542 VSS.n5539 0.0655943
R8048 VSS.n5593 VSS.n5590 0.0655943
R8049 VSS.n74 VSS.n73 0.0649262
R8050 VSS.n5114 VSS.n5113 0.0644344
R8051 VSS.n80 VSS.n79 0.0640294
R8052 VSS.n4096 VSS.n4093 0.0640294
R8053 VSS.n1309 VSS.n955 0.0639286
R8054 VSS.n5814 VSS.n5813 0.0636651
R8055 VSS.n5094 VSS.n5093 0.0636492
R8056 VSS.n86 VSS.n85 0.0636492
R8057 VSS.n5059 VSS.n5058 0.0633022
R8058 VSS.n4508 VSS.n4507 0.0633022
R8059 VSS.n75 VSS.n74 0.062959
R8060 VSS.n5115 VSS.n5114 0.062959
R8061 VSS.n729 VSS.n728 0.0626951
R8062 VSS.n5087 VSS.n5086 0.0622838
R8063 VSS.n94 VSS.n93 0.0622838
R8064 VSS.n4411 VSS.n4391 0.0621304
R8065 VSS.n5265 VSS.n5264 0.0618391
R8066 VSS.n310 VSS.n309 0.0616009
R8067 VSS.n302 VSS.n301 0.0616009
R8068 VSS.n4570 VSS.n4508 0.0613736
R8069 VSS.n4578 VSS.n94 0.0611892
R8070 VSS.n208 VSS.n205 0.0611522
R8071 VSS.n4252 VSS.n4251 0.0605
R8072 VSS.n5157 VSS.n5154 0.0603902
R8073 VSS.n5218 VSS.n5217 0.0601739
R8074 VSS.n929 VSS.n926 0.0596608
R8075 VSS.n931 VSS.n929 0.0596608
R8076 VSS.n932 VSS.n931 0.0596608
R8077 VSS.n937 VSS 0.0596608
R8078 VSS.n945 VSS.n942 0.0596608
R8079 VSS.n947 VSS.n945 0.0596608
R8080 VSS.n4849 VSS.n4846 0.0596608
R8081 VSS.n4852 VSS.n4849 0.0596608
R8082 VSS.n4853 VSS.n4852 0.0596608
R8083 VSS VSS.n4853 0.0596608
R8084 VSS.n4861 VSS.n4858 0.0596608
R8085 VSS.n4864 VSS.n4861 0.0596608
R8086 VSS.n4867 VSS.n4864 0.0596608
R8087 VSS.n4811 VSS.n4808 0.0596608
R8088 VSS.n4814 VSS.n4811 0.0596608
R8089 VSS.n4815 VSS.n4814 0.0596608
R8090 VSS VSS.n4815 0.0596608
R8091 VSS.n4823 VSS.n4820 0.0596608
R8092 VSS.n4826 VSS.n4823 0.0596608
R8093 VSS.n4829 VSS.n4826 0.0596608
R8094 VSS.n4883 VSS.n4880 0.0596608
R8095 VSS.n4886 VSS.n4883 0.0596608
R8096 VSS.n4887 VSS.n4886 0.0596608
R8097 VSS VSS.n4887 0.0596608
R8098 VSS.n4895 VSS.n4892 0.0596608
R8099 VSS.n4900 VSS.n4895 0.0596608
R8100 VSS.n4903 VSS.n4900 0.0596608
R8101 VSS.n4924 VSS.n4921 0.0596608
R8102 VSS.n4927 VSS.n4924 0.0596608
R8103 VSS.n4928 VSS.n4927 0.0596608
R8104 VSS VSS.n4928 0.0596608
R8105 VSS.n4936 VSS.n4933 0.0596608
R8106 VSS.n4939 VSS.n4936 0.0596608
R8107 VSS.n4942 VSS.n4939 0.0596608
R8108 VSS.n4143 VSS.n4140 0.0596608
R8109 VSS.n4145 VSS.n4143 0.0596608
R8110 VSS.n164 VSS.n161 0.0594119
R8111 VSS.n5849 VSS.n5846 0.0587734
R8112 VSS.n767 VSS.n763 0.0583049
R8113 VSS.n4020 VSS.n4019 0.0574719
R8114 VSS.n4422 VSS.n4419 0.0572391
R8115 VSS.n5003 VSS.n5000 0.0568736
R8116 VSS.n4655 VSS.n4652 0.0568736
R8117 VSS.n5602 VSS.n5599 0.0559717
R8118 VSS.n406 VSS.n405 0.055378
R8119 VSS.n409 VSS.n406 0.055378
R8120 VSS.n413 VSS.n412 0.055378
R8121 VSS.n416 VSS.n413 0.055378
R8122 VSS.n5184 VSS.n5181 0.0552826
R8123 VSS.n932 VSS.n922 0.0552552
R8124 VSS.n4858 VSS.n4836 0.0552552
R8125 VSS.n4820 VSS.n4799 0.0552552
R8126 VSS.n4892 VSS.n4793 0.0552552
R8127 VSS.n4933 VSS.n4911 0.0552552
R8128 VSS VSS.n218 0.0549444
R8129 VSS.n5207 VSS 0.0543889
R8130 VSS.n191 VSS.n188 0.0543043
R8131 VSS.n4008 VSS.n4007 0.0536953
R8132 VSS VSS.n4147 0.0533671
R8133 VSS.n4184 VSS.n4181 0.0533671
R8134 VSS.n4443 VSS.n4440 0.0530777
R8135 VSS.n5426 VSS.n5423 0.0530398
R8136 VSS.n1037 VSS.n1034 0.0526341
R8137 VSS.n4019 VSS.n4016 0.0521084
R8138 VSS.n4007 VSS.n4004 0.0521084
R8139 VSS.n5085 VSS.n5084 0.0514211
R8140 VSS.n4873 VSS.n4833 0.0513891
R8141 VSS.n5254 VSS.n4765 0.0513696
R8142 VSS.n4197 VSS.n4195 0.0508497
R8143 VSS.n4355 VSS.n99 0.050439
R8144 VSS.n4093 VSS.n1391 0.050416
R8145 VSS.n4255 VSS.n4252 0.0502561
R8146 VSS.n701 VSS.n700 0.0498902
R8147 VSS.n4335 VSS.n4334 0.0498902
R8148 VSS.n4977 VSS.n4974 0.0498805
R8149 VSS.n885 VSS.n884 0.0496753
R8150 VSS.n1030 VSS.n1029 0.0486818
R8151 VSS.n6061 VSS.n6060 0.0486818
R8152 VSS.n5555 VSS.n5554 0.0486132
R8153 VSS.n4030 VSS.n4027 0.0483322
R8154 VSS.n4313 VSS.n787 0.0476951
R8155 VSS.n1313 VSS.n1309 0.0466345
R8156 VSS.n4471 VSS 0.0462895
R8157 VSS VSS.n5204 0.0460556
R8158 VSS.n6066 VSS.n6065 0.0459545
R8159 VSS.n6065 VSS.n6064 0.0459545
R8160 VSS.n4276 VSS.n4270 0.0458659
R8161 VSS.n5783 VSS.n5782 0.0457506
R8162 VSS.n93 VSS.n92 0.0457432
R8163 VSS.n219 VSS 0.0455
R8164 VSS.n5449 VSS 0.0455
R8165 VSS.n5309 VSS.n5308 0.0455
R8166 VSS.n5086 VSS.n5085 0.0452568
R8167 VSS.n5813 VSS 0.0450872
R8168 VSS.n73 VSS.n68 0.04425
R8169 VSS.n5113 VSS.n5108 0.04425
R8170 VSS.n1650 VSS.n1649 0.044243
R8171 VSS.n950 VSS.n948 0.0439266
R8172 VSS.n4877 VSS.n4876 0.0439266
R8173 VSS.n4918 VSS.n4917 0.0439266
R8174 VSS.n4138 VSS.n4137 0.0439266
R8175 VSS.n5247 VSS.n5246 0.0435435
R8176 VSS.n4663 VSS.n4662 0.0435088
R8177 VSS.n1029 VSS.n0 0.0432273
R8178 VSS.n1302 VSS.n1301 0.0428529
R8179 VSS.n4993 VSS.n4990 0.0427124
R8180 VSS.n82 VSS.n81 0.0426277
R8181 VSS.n1505 VSS.n1408 0.0425561
R8182 VSS.n5647 VSS.n5646 0.0422073
R8183 VSS.n5650 VSS.n5647 0.0411098
R8184 VSS.n1687 VSS.n1673 0.0404721
R8185 VSS.n4580 VSS.n4578 0.040323
R8186 VSS.n1523 VSS.n1522 0.0401503
R8187 VSS.n5074 VSS.n5072 0.0395266
R8188 VSS.n1034 VSS.n1008 0.0394634
R8189 VSS.n4389 VSS.n4386 0.0386522
R8190 VSS.n4067 VSS.n4064 0.0385488
R8191 VSS.n5779 VSS.n5778 0.0377928
R8192 VSS.n5804 VSS.n5803 0.037656
R8193 VSS.n938 VSS.n937 0.0376329
R8194 VSS.n5443 VSS.n5442 0.0376053
R8195 VSS.n5558 VSS.n5555 0.0372925
R8196 VSS.n6065 VSS.n21 0.0372105
R8197 VSS.n1564 VSS.n1563 0.0368785
R8198 VSS.n1568 VSS.n1567 0.0368564
R8199 VSS.n775 VSS.n774 0.0367195
R8200 VSS.n5309 VSS.n5262 0.0366957
R8201 VSS.n4952 VSS.n4949 0.0363407
R8202 VSS.n41 VSS.n39 0.0363407
R8203 VSS.n1404 VSS.n1403 0.0357448
R8204 VSS.n4375 VSS.n4374 0.0352779
R8205 VSS.n5278 VSS.n5277 0.0352465
R8206 VSS.n924 VSS.n919 0.0351154
R8207 VSS.n3981 VSS.n3980 0.0351154
R8208 VSS.n4871 VSS.n4868 0.0351154
R8209 VSS.n4833 VSS.n4830 0.0351154
R8210 VSS.n4907 VSS.n4904 0.0351154
R8211 VSS.n4946 VSS.n4943 0.0351154
R8212 VSS.n4185 VSS.n4184 0.0351154
R8213 VSS.n4201 VSS.n4198 0.0351154
R8214 VSS.n4680 VSS.n4679 0.0347478
R8215 VSS.n3994 VSS.n3993 0.034486
R8216 VSS.n4125 VSS.n912 0.0334464
R8217 VSS.n739 VSS.n736 0.0334268
R8218 VSS.n4337 VSS.n4335 0.0334268
R8219 VSS.n4569 VSS.n4568 0.0331549
R8220 VSS.n4355 VSS.n4354 0.032878
R8221 VSS.n4146 VSS.n4145 0.0325979
R8222 VSS.n4604 VSS.n4600 0.0323584
R8223 VSS.n3071 VSS.n1815 0.0323182
R8224 VSS.n1645 VSS.n1579 0.0320446
R8225 VSS.n1551 VSS.n1550 0.032
R8226 VSS.n1726 VSS.n1721 0.032
R8227 VSS.n1541 VSS.n1540 0.032
R8228 VSS.n4031 VSS.n4030 0.0319685
R8229 VSS.n4699 VSS.n4695 0.0318333
R8230 VSS.n4703 VSS.n4699 0.0318333
R8231 VSS.n4713 VSS.n4703 0.0318333
R8232 VSS.n4719 VSS 0.0318333
R8233 VSS.n4723 VSS.n4719 0.0318333
R8234 VSS.n4727 VSS.n4723 0.0318333
R8235 VSS.n4731 VSS.n4727 0.0318333
R8236 VSS.n5125 VSS.n5123 0.0315619
R8237 VSS.n1558 VSS.n1557 0.0309839
R8238 VSS.n5828 VSS.n5827 0.0308614
R8239 VSS.n314 VSS.n313 0.0305726
R8240 VSS.n1679 VSS.n1678 0.0302848
R8241 VSS.n4982 VSS.n4978 0.029969
R8242 VSS.n4673 VSS.n4672 0.029969
R8243 VSS.n1664 VSS.n1663 0.0299134
R8244 VSS.n4713 VSS.n4708 0.0295
R8245 VSS.n887 VSS.n886 0.0292629
R8246 VSS.n1586 VSS.n1585 0.0291175
R8247 VSS.n2439 VSS.n2429 0.0289279
R8248 VSS.n4153 VSS.n788 0.0288217
R8249 VSS.n966 VSS.n964 0.028625
R8250 VSS.n286 VSS.n283 0.028625
R8251 VSS.n330 VSS.n327 0.028625
R8252 VSS.n3506 VSS.n3500 0.028625
R8253 VSS.n4089 VSS.n4088 0.028625
R8254 VSS.n4126 VSS.n4125 0.028625
R8255 VSS.n4215 VSS.n4212 0.028625
R8256 VSS.n1165 VSS.n992 0.0284878
R8257 VSS.n872 VSS.n871 0.0284
R8258 VSS.n4563 VSS.n4560 0.0283761
R8259 VSS.n886 VSS.n885 0.0283351
R8260 VSS.n5755 VSS.n5746 0.0282695
R8261 VSS.n4031 VSS.n3984 0.0281923
R8262 VSS.n5430 VSS.n5427 0.0281316
R8263 VSS.n1613 VSS.n1612 0.0276659
R8264 VSS.n5063 VSS.n5061 0.0275796
R8265 VSS.n873 VSS.n872 0.0275
R8266 VSS.n1574 VSS.n1573 0.0274585
R8267 VSS.n90 VSS.n89 0.0273085
R8268 VSS.n5083 VSS.n5082 0.0273085
R8269 VSS.n253 VSS.n101 0.026913
R8270 VSS.n1677 VSS.n1676 0.0266
R8271 VSS.n1682 VSS.n1681 0.0266
R8272 VSS.n4370 VSS.n4369 0.0265939
R8273 VSS.n1502 VSS.n1409 0.0265748
R8274 VSS.n1448 VSS.n1447 0.0265748
R8275 VSS.n5804 VSS.n5796 0.0265092
R8276 VSS.n5803 VSS.n5802 0.0265092
R8277 VSS.n5882 VSS.n5881 0.0264481
R8278 VSS.n2803 VSS.n2082 0.0262358
R8279 VSS.n5274 VSS.n5272 0.0261799
R8280 VSS.n1899 VSS.n1898 0.0261034
R8281 VSS.n312 VSS.n311 0.0260963
R8282 VSS.n4368 VSS.n4367 0.0259717
R8283 VSS.n5271 VSS.n5270 0.0259717
R8284 VSS.n1703 VSS.n1702 0.0258911
R8285 VSS.n1446 VSS.n1445 0.0257336
R8286 VSS.n1447 VSS.n1408 0.0257336
R8287 VSS.n1547 VSS.n1546 0.0257
R8288 VSS.n1723 VSS.n1722 0.0257
R8289 VSS.n1537 VSS.n1536 0.0257
R8290 VSS.n1434 VSS.n1431 0.0256748
R8291 VSS.n1440 VSS.n1437 0.0256748
R8292 VSS.n1497 VSS.n1494 0.0256748
R8293 VSS.n1491 VSS.n1488 0.0256748
R8294 VSS.n806 VSS.n803 0.0256748
R8295 VSS.n812 VSS.n809 0.0256748
R8296 VSS.n818 VSS.n815 0.0256748
R8297 VSS.n846 VSS.n843 0.0256748
R8298 VSS.n853 VSS.n850 0.0256748
R8299 VSS.n1596 VSS.n1595 0.0255922
R8300 VSS.n2179 VSS.n2143 0.0254833
R8301 VSS.n1582 VSS.n1581 0.0253848
R8302 VSS.n2805 VSS.n2088 0.0253328
R8303 VSS.n2307 VSS.n2284 0.0253328
R8304 VSS.n311 VSS.n310 0.0252706
R8305 VSS.n308 VSS.n307 0.0252706
R8306 VSS.n4960 VSS.n4959 0.0251903
R8307 VSS.n47 VSS.n46 0.0251903
R8308 VSS.n2797 VSS.n2796 0.0251823
R8309 VSS.n1914 VSS.n1913 0.0251724
R8310 VSS.n926 VSS.n924 0.0250455
R8311 VSS.n1501 VSS.n1475 0.0250455
R8312 VSS.n3984 VSS.n3981 0.0250455
R8313 VSS.n4868 VSS.n4867 0.0250455
R8314 VSS.n4830 VSS.n4829 0.0250455
R8315 VSS.n4904 VSS.n4903 0.0250455
R8316 VSS.n4943 VSS.n4942 0.0250455
R8317 VSS.n4198 VSS.n4197 0.0250455
R8318 VSS.n2429 VSS.n2413 0.0249978
R8319 VSS.n1570 VSS 0.0247376
R8320 VSS.n820 VSS.n819 0.0247308
R8321 VSS.n5277 VSS.n5263 0.0247308
R8322 VSS.n335 VSS.n334 0.024574
R8323 VSS.n2808 VSS.n2807 0.0244298
R8324 VSS.n1811 VSS.n1810 0.0243636
R8325 VSS.n1625 VSS.n1624 0.0241406
R8326 VSS.n694 VSS.n691 0.0240976
R8327 VSS.n5901 VSS.n5898 0.0240976
R8328 VSS.n5413 VSS.n5410 0.0239783
R8329 VSS.n1806 VSS.n1805 0.0236818
R8330 VSS.n1808 VSS.n1804 0.0236818
R8331 VSS.n1606 VSS.n1605 0.0235184
R8332 VSS.n4737 VSS.n4732 0.0235
R8333 VSS.n5267 VSS.n5266 0.0234789
R8334 VSS VSS.n5879 0.0234091
R8335 VSS.n3583 VSS.n3582 0.0233924
R8336 VSS.n161 VSS.n160 0.0232368
R8337 VSS VSS.n5835 0.0231603
R8338 VSS.n4364 VSS.n4363 0.0230525
R8339 VSS.n5254 VSS.n5253 0.023
R8340 VSS.n3505 VSS.n3504 0.0228692
R8341 VSS.n2956 VSS.n2955 0.0228692
R8342 VSS.n5154 VSS.n5144 0.0227632
R8343 VSS.n942 VSS.n938 0.022528
R8344 VSS.n2486 VSS.n2485 0.0225087
R8345 VSS.n1715 VSS.n1714 0.0221201
R8346 VSS.n4398 VSS.n4397 0.0220702
R8347 VSS.n1637 VSS.n1636 0.0220668
R8348 VSS.n5075 VSS.n5074 0.0220044
R8349 VSS.n346 VSS.n343 0.0217195
R8350 VSS.n273 VSS.n272 0.0213929
R8351 VSS.n4401 VSS.n4400 0.0213264
R8352 VSS.n5293 VSS.n5292 0.0213264
R8353 VSS.n5296 VSS.n5295 0.0213264
R8354 VSS.n4374 VSS.n4373 0.0212692
R8355 VSS.n4581 VSS.n4580 0.021208
R8356 VSS.n4506 VSS.n96 0.0209545
R8357 VSS.n5057 VSS.n5054 0.0209545
R8358 VSS.n6063 VSS.n6062 0.0209545
R8359 VSS.n4365 VSS.n4364 0.0208774
R8360 VSS.n2915 VSS.n2914 0.020815
R8361 VSS.n349 VSS.n347 0.0207174
R8362 VSS.n317 VSS.n268 0.0207174
R8363 VSS.n1461 VSS 0.0206399
R8364 VSS.n2141 VSS.n2131 0.0205167
R8365 VSS.n2294 VSS.n2293 0.0205167
R8366 VSS.n4593 VSS.n4589 0.0204115
R8367 VSS.n2574 VSS.n2573 0.0203837
R8368 VSS.n300 VSS.n299 0.0203165
R8369 VSS.n5539 VSS.n5401 0.0203113
R8370 VSS.n5590 VSS.n5589 0.0203113
R8371 VSS.n2543 VSS.n2430 0.0201507
R8372 VSS.n245 VSS.n120 0.0200652
R8373 VSS.n349 VSS.n348 0.0200652
R8374 VSS.n317 VSS.n316 0.0200652
R8375 VSS.n5530 VSS.n5528 0.0200447
R8376 VSS.n5268 VSS.n5267 0.0200283
R8377 VSS.n4166 VSS.n4165 0.0199845
R8378 VSS.n5793 VSS.n5792 0.0198944
R8379 VSS.n3499 VSS.n3498 0.0198605
R8380 VSS.n4404 VSS.n4403 0.0198388
R8381 VSS.n297 VSS.n276 0.0197857
R8382 VSS.n4502 VSS.n4501 0.0197025
R8383 VSS.n5101 VSS.n5098 0.019615
R8384 VSS.n144 VSS.n143 0.0196091
R8385 VSS.n2591 VSS.n2404 0.0195988
R8386 VSS.n353 VSS.n352 0.0195947
R8387 VSS.n5197 VSS.n5196 0.019555
R8388 VSS.n4777 VSS.n4776 0.019555
R8389 VSS.n2541 VSS.n2431 0.0193646
R8390 VSS.n5149 VSS.n5148 0.0193395
R8391 VSS.n127 VSS.n126 0.0191251
R8392 VSS.n225 VSS.n224 0.0191251
R8393 VSS.n5299 VSS.n5298 0.019095
R8394 VSS.n247 VSS.n245 0.019087
R8395 VSS.n3457 VSS.n3456 0.0190756
R8396 VSS.n4163 VSS.n4162 0.0190567
R8397 VSS.n2721 VSS.n2213 0.0190117
R8398 VSS.n291 VSS.n290 0.0189821
R8399 VSS.n5874 VSS.n5850 0.0189532
R8400 VSS.n3617 VSS.n3616 0.0189448
R8401 VSS.n355 VSS.n354 0.0188673
R8402 VSS.n2589 VSS.n2405 0.018814
R8403 VSS.n5200 VSS.n5199 0.0186836
R8404 VSS.n4780 VSS.n4779 0.0186836
R8405 VSS.n5174 VSS.n5173 0.0186836
R8406 VSS.n306 VSS.n305 0.0186651
R8407 VSS.n5787 VSS.n5786 0.0186268
R8408 VSS.n2539 VSS.n2432 0.0185786
R8409 VSS.n3989 VSS.n3988 0.0185
R8410 VSS.n883 VSS.n882 0.0185
R8411 VSS.n4406 VSS.n4405 0.018485
R8412 VSS.n5298 VSS.n5297 0.0184602
R8413 VSS.n1444 VSS.n1443 0.0184371
R8414 VSS.n3446 VSS.n3445 0.0182907
R8415 VSS.n2732 VSS.n2731 0.0182592
R8416 VSS.n4173 VSS.n4172 0.0181289
R8417 VSS.n4386 VSS.n4385 0.0181087
R8418 VSS.n2719 VSS.n2214 0.0181087
R8419 VSS.n5301 VSS.n5300 0.0181073
R8420 VSS.n4403 VSS.n4402 0.0180867
R8421 VSS.n2587 VSS.n2408 0.0180291
R8422 VSS.n5129 VSS.n5128 0.0180221
R8423 VSS.n4966 VSS.n4965 0.0180221
R8424 VSS.n5789 VSS 0.017993
R8425 VSS.n304 VSS.n303 0.0178394
R8426 VSS.n134 VSS.n131 0.0178182
R8427 VSS.n177 VSS.n174 0.0178182
R8428 VSS.n232 VSS.n229 0.0178182
R8429 VSS.n1425 VSS.n1424 0.0178077
R8430 VSS.n1482 VSS.n1481 0.0178077
R8431 VSS.n797 VSS.n796 0.0178077
R8432 VSS.n863 VSS.n862 0.0178077
R8433 VSS.n2855 VSS.n2021 0.0178077
R8434 VSS.n2292 VSS.n2212 0.0176572
R8435 VSS.n3502 VSS.n3501 0.0176366
R8436 VSS.n1549 VSS.n1548 0.0175923
R8437 VSS.n1539 VSS.n1538 0.0175923
R8438 VSS.n3990 VSS.n3987 0.0175
R8439 VSS.n870 VSS.n856 0.017493
R8440 VSS.n972 VSS.n967 0.0174458
R8441 VSS.n967 VSS.n966 0.0173807
R8442 VSS.n272 VSS.n271 0.017375
R8443 VSS.n275 VSS.n274 0.017375
R8444 VSS.n2570 VSS.n2569 0.017375
R8445 VSS.n2201 VSS.n2194 0.0173562
R8446 VSS.n4608 VSS.n4607 0.0172257
R8447 VSS.n2717 VSS.n2215 0.0172057
R8448 VSS.n971 VSS.n968 0.0171955
R8449 VSS.n253 VSS.n252 0.0171304
R8450 VSS.n264 VSS.n263 0.0170306
R8451 VSS.n3071 VSS.n3070 0.0167984
R8452 VSS.n2855 VSS.n2854 0.0167542
R8453 VSS.n1407 VSS.n1406 0.0165
R8454 VSS.n2021 VSS.n1995 0.0164532
R8455 VSS.n2207 VSS.n2206 0.0164532
R8456 VSS.n4570 VSS.n4569 0.0164292
R8457 VSS.n4170 VSS.n4169 0.0162732
R8458 VSS.n948 VSS.n947 0.0162343
R8459 VSS.n4846 VSS.n4843 0.0162343
R8460 VSS.n4808 VSS.n4805 0.0162343
R8461 VSS.n4880 VSS.n4877 0.0162343
R8462 VSS.n4921 VSS.n4918 0.0162343
R8463 VSS.n4140 VSS.n4138 0.0162343
R8464 VSS.n2545 VSS.n2428 0.0162205
R8465 VSS.n5211 VSS.n5208 0.0161522
R8466 VSS.n318 VSS.n267 0.0161122
R8467 VSS.n3402 VSS.n3401 0.0160669
R8468 VSS.n736 VSS.n713 0.0158659
R8469 VSS.n5295 VSS.n5294 0.015852
R8470 VSS.n877 VSS.n876 0.0158
R8471 VSS.n1469 VSS 0.0156049
R8472 VSS.n1853 VSS.n1852 0.0155517
R8473 VSS.n1512 VSS.n1407 0.0155
R8474 VSS.n2547 VSS.n2424 0.0154345
R8475 VSS.n2184 VSS.n2129 0.0153997
R8476 VSS.n5270 VSS.n5269 0.015398
R8477 VSS.n2302 VSS.n2301 0.0152492
R8478 VSS.n215 VSS.n214 0.0151739
R8479 VSS.n4400 VSS.n4399 0.0151082
R8480 VSS.n5292 VSS.n5291 0.0151082
R8481 VSS.n2828 VSS.n2068 0.0150987
R8482 VSS.n3586 VSS.n3585 0.0150203
R8483 VSS.n3393 VSS.n3392 0.0148895
R8484 VSS.n5068 VSS.n5066 0.0148363
R8485 VSS.n5275 VSS.n5265 0.0148234
R8486 VSS.n4371 VSS.n4360 0.0148073
R8487 VSS.n5633 VSS.n5632 0.0147683
R8488 VSS.n4397 VSS.n4396 0.0147345
R8489 VSS.n840 VSS.n789 0.0146608
R8490 VSS.n2550 VSS.n2549 0.0146485
R8491 VSS.n3611 VSS.n3610 0.0146279
R8492 VSS.n1893 VSS.n1892 0.0146207
R8493 VSS.n4367 VSS.n4366 0.014549
R8494 VSS.n2746 VSS.n2745 0.0144967
R8495 VSS.n1872 VSS.n1871 0.0144655
R8496 VSS.n358 VSS.n357 0.0144024
R8497 VSS.n2678 VSS.n2677 0.0143462
R8498 VSS.n2830 VSS.n2065 0.0141957
R8499 VSS.n5830 VSS.n5829 0.0141817
R8500 VSS.n296 VSS 0.0141607
R8501 VSS.n319 VSS.n262 0.0141607
R8502 VSS.n1505 VSS.n1504 0.0141607
R8503 VSS.n5796 VSS.n5795 0.0141239
R8504 VSS.n3525 VSS.n3524 0.0141047
R8505 VSS.n2878 VSS.n1996 0.0140452
R8506 VSS.n4970 VSS.n4969 0.0140398
R8507 VSS.n57 VSS.n56 0.0140398
R8508 VSS.n1660 VSS.n1659 0.0140123
R8509 VSS.n1690 VSS.n1689 0.0140123
R8510 VSS.n1668 VSS.n1667 0.0140123
R8511 VSS.n1453 VSS.n1452 0.0139579
R8512 VSS.n4691 VSS.n4690 0.0138333
R8513 VSS.n2518 VSS.n2453 0.0137314
R8514 VSS.n1930 VSS.n1929 0.0136897
R8515 VSS.n5619 VSS.n5616 0.0136707
R8516 VSS.n2166 VSS.n2163 0.0135936
R8517 VSS.n1877 VSS.n1876 0.0135345
R8518 VSS.n4695 VSS.n4691 0.0135
R8519 VSS.n4169 VSS.n4168 0.0134897
R8520 VSS.n2271 VSS.n2268 0.0134431
R8521 VSS.n3487 VSS.n3486 0.0133198
R8522 VSS.n2833 VSS.n2832 0.0132926
R8523 VSS.n1815 VSS.n1814 0.0132273
R8524 VSS.n2944 VSS.n2943 0.013189
R8525 VSS.n2876 VSS.n1997 0.0131421
R8526 VSS.n4161 VSS.n4160 0.0130874
R8527 VSS.n2516 VSS.n2454 0.0129454
R8528 VSS.n1977 VSS.n1976 0.0126034
R8529 VSS.n3850 VSS.n3849 0.0125737
R8530 VSS.n774 VSS.n751 0.0125732
R8531 VSS.n3559 VSS.n3558 0.0125349
R8532 VSS.n3990 VSS.n3989 0.0125
R8533 VSS.n4175 VSS.n4174 0.012458
R8534 VSS.n267 VSS.n266 0.0124388
R8535 VSS.n83 VSS.n78 0.0124337
R8536 VSS.n5095 VSS.n5094 0.0124337
R8537 VSS.n4505 VSS.n4504 0.0123681
R8538 VSS.n72 VSS.n69 0.0123033
R8539 VSS.n5116 VSS.n5115 0.0123033
R8540 VSS.n1454 VSS.n1453 0.0122757
R8541 VSS.n2874 VSS.n1998 0.0122391
R8542 VSS.n876 VSS.n875 0.0122
R8543 VSS.n2514 VSS.n2456 0.0121594
R8544 VSS.n81 VSS.n80 0.0119894
R8545 VSS.n4585 VSS.n86 0.0119365
R8546 VSS.n5091 VSS.n5089 0.0119365
R8547 VSS.n5056 VSS.n5055 0.0118736
R8548 VSS.n4027 VSS.n4026 0.0118287
R8549 VSS.n4597 VSS.n75 0.0118115
R8550 VSS.n5112 VSS.n5109 0.0118115
R8551 VSS.n2788 VSS.n2095 0.0117876
R8552 VSS.n360 VSS.n337 0.01175
R8553 VSS.n2605 VSS.n2389 0.0116192
R8554 VSS.n352 VSS.n351 0.0115204
R8555 VSS.n71 VSS.n70 0.0113172
R8556 VSS.n5111 VSS.n5110 0.0113172
R8557 VSS.n3996 VSS.n3995 0.0111993
R8558 VSS.n2809 VSS.n2086 0.0111355
R8559 VSS.n964 VSS.n961 0.0109464
R8560 VSS.n289 VSS.n286 0.0109464
R8561 VSS.n320 VSS.n319 0.0109464
R8562 VSS.n4218 VSS.n4215 0.0109464
R8563 VSS.n2786 VSS.n2096 0.0108846
R8564 VSS.n2607 VSS.n2386 0.0108343
R8565 VSS.n4172 VSS.n4171 0.0107062
R8566 VSS.n1653 VSS.n1652 0.0106256
R8567 VSS.n2655 VSS.n2321 0.0105727
R8568 VSS.n1472 VSS.n1469 0.0105699
R8569 VSS.n3993 VSS.n1523 0.0105699
R8570 VSS.n4187 VSS.n4186 0.0105699
R8571 VSS.n2139 VSS.n2138 0.0104331
R8572 VSS.n2700 VSS.n2237 0.0104331
R8573 VSS.n1684 VSS.n1683 0.0102906
R8574 VSS.n973 VSS.n972 0.0101429
R8575 VSS.n1506 VSS.n1505 0.0101429
R8576 VSS.n333 VSS.n330 0.0101429
R8577 VSS.n4090 VSS.n4089 0.0101429
R8578 VSS.n4127 VSS.n4126 0.0101429
R8579 VSS.n3867 VSS.n3866 0.0100852
R8580 VSS.n3588 VSS.n3587 0.0100494
R8581 VSS.n2610 VSS.n2609 0.0100494
R8582 VSS.n343 VSS.n322 0.0100122
R8583 VSS.n5786 VSS.n5785 0.010007
R8584 VSS.n2784 VSS.n2097 0.00998161
R8585 VSS.n5116 VSS.n5103 0.00997368
R8586 VSS.n1522 VSS.n1521 0.00994056
R8587 VSS.n1514 VSS.n1513 0.00994056
R8588 VSS.n3885 VSS.n3884 0.00989535
R8589 VSS.n3809 VSS.n3808 0.00982401
R8590 VSS.n2653 VSS.n2322 0.00978779
R8591 VSS.n4164 VSS.n4163 0.00977835
R8592 VSS.n4173 VSS.n4166 0.00977835
R8593 VSS.n2964 VSS.n2963 0.00974419
R8594 VSS.n356 VSS.n355 0.00968367
R8595 VSS.n2131 VSS.n2130 0.0096806
R8596 VSS.n1577 VSS 0.00958911
R8597 VSS.n881 VSS.n880 0.00958707
R8598 VSS.n2766 VSS.n2765 0.0095301
R8599 VSS.n2698 VSS.n2238 0.0095301
R8600 VSS.n2332 VSS.n2320 0.00952616
R8601 VSS.n4597 VSS.n4596 0.0095
R8602 VSS.n3585 VSS.n3584 0.00939535
R8603 VSS.n4186 VSS.n4185 0.00931119
R8604 VSS.n4195 VSS.n4194 0.00931119
R8605 VSS.n3384 VSS.n3383 0.00926454
R8606 VSS.n68 VSS.n67 0.00925
R8607 VSS.n5108 VSS.n5107 0.00925
R8608 VSS.n4588 VSS.n4585 0.00902632
R8609 VSS.n2651 VSS.n2323 0.00900291
R8610 VSS.n5573 VSS.n5570 0.00899057
R8611 VSS.n3516 VSS.n3515 0.00887209
R8612 VSS.n4732 VSS.n4731 0.00883333
R8613 VSS.n1405 VSS.n1404 0.00868182
R8614 VSS.n870 VSS.n869 0.00868182
R8615 VSS.n4160 VSS.n4159 0.00868182
R8616 VSS.n4180 VSS.n4175 0.00868182
R8617 VSS.n2130 VSS.n2094 0.00862709
R8618 VSS.n2119 VSS.n2116 0.00862709
R8619 VSS.n2295 VSS.n2294 0.00862709
R8620 VSS.n2696 VSS.n2241 0.00862709
R8621 VSS.n3858 VSS.n3857 0.0086106
R8622 VSS.n2630 VSS.n2629 0.00861047
R8623 VSS.n5097 VSS.n5095 0.00855263
R8624 VSS.n2886 VSS.n2885 0.00855063
R8625 VSS.n3284 VSS.n3283 0.00847965
R8626 VSS.n3569 VSS.n3568 0.00840698
R8627 VSS.n2538 VSS.n2537 0.00838571
R8628 VSS.n1553 VSS.n1552 0.00836872
R8629 VSS.n1725 VSS.n1724 0.00836872
R8630 VSS.n1543 VSS.n1542 0.00836872
R8631 VSS.n1428 VSS.n1425 0.00836713
R8632 VSS.n1485 VSS.n1482 0.00836713
R8633 VSS.n800 VSS.n797 0.00836713
R8634 VSS.n866 VSS.n863 0.00836713
R8635 VSS.n2569 VSS.n2332 0.00834884
R8636 VSS.n3773 VSS.n3772 0.00833217
R8637 VSS.n198 VSS.n195 0.00832609
R8638 VSS.n2586 VSS.n2585 0.0082907
R8639 VSS.n3473 VSS.n3472 0.00808721
R8640 VSS.n3228 VSS.n3227 0.00808721
R8641 VSS.n4004 VSS.n4003 0.00805245
R8642 VSS.n3995 VSS.n3994 0.00805245
R8643 VSS.n3905 VSS.n3904 0.0080419
R8644 VSS.n1673 VSS.n1650 0.0080419
R8645 VSS.n2796 VSS.n2022 0.00802508
R8646 VSS.n1288 VSS.n1284 0.008
R8647 VSS.n3625 VSS.n3624 0.00797826
R8648 VSS.n1168 VSS.n1165 0.00795562
R8649 VSS.n1866 VSS.n1865 0.00794828
R8650 VSS.n305 VSS.n304 0.00793119
R8651 VSS.n303 VSS.n302 0.00793119
R8652 VSS.n265 VSS.n264 0.00784694
R8653 VSS.n2349 VSS.n2347 0.00782558
R8654 VSS.n357 VSS.n346 0.00781707
R8655 VSS.n1663 VSS.n1662 0.0077905
R8656 VSS.n1709 VSS.n1708 0.0077905
R8657 VSS.n3897 VSS.n1718 0.0077905
R8658 VSS.n1649 VSS.n1648 0.0077905
R8659 VSS.n274 VSS.n273 0.00773214
R8660 VSS.n2857 VSS.n2015 0.00772408
R8661 VSS.n3290 VSS.n3289 0.00769477
R8662 VSS.n5534 VSS.n5531 0.00760526
R8663 VSS.n2232 VSS.n2231 0.00757358
R8664 VSS.n1508 VSS.n1507 0.00757142
R8665 VSS.n1662 VSS.n1657 0.00753911
R8666 VSS.n1669 VSS.n1664 0.00753911
R8667 VSS.n1697 VSS.n1696 0.00753911
R8668 VSS.n2716 VSS.n2715 0.00748113
R8669 VSS.n1504 VSS.n1503 0.00743371
R8670 VSS VSS.n4008 0.00742308
R8671 VSS.n4003 VSS.n3996 0.00742308
R8672 VSS.n882 VSS.n881 0.00735714
R8673 VSS.n5228 VSS.n5227 0.00734783
R8674 VSS.n1611 VSS.n1610 0.00734332
R8675 VSS.n1641 VSS.n1640 0.00734332
R8676 VSS.n2208 VSS.n2198 0.0073277
R8677 VSS.n3545 VSS.n3544 0.00730233
R8678 VSS.n1671 VSS.n1670 0.00728771
R8679 VSS.n1713 VSS.n1712 0.00728771
R8680 VSS.n1813 VSS.n1812 0.00726364
R8681 VSS.n1609 VSS.n1608 0.00713594
R8682 VSS.n1639 VSS.n1638 0.00713594
R8683 VSS.n767 VSS.n766 0.00708537
R8684 VSS.n4330 VSS.n4328 0.00708537
R8685 VSS.n2356 VSS.n2354 0.0070407
R8686 VSS.n3907 VSS.n1691 0.00703631
R8687 VSS.n1701 VSS.n1700 0.00703631
R8688 VSS.n1705 VSS.n1704 0.00703631
R8689 VSS.n3803 VSS.n3794 0.00701869
R8690 VSS.n1961 VSS.n1960 0.00701724
R8691 VSS.n5113 VSS.n5112 0.00689344
R8692 VSS.n1032 VSS.n1024 0.00686364
R8693 VSS.n1862 VSS.n1861 0.00686207
R8694 VSS.n2859 VSS.n2012 0.00682107
R8695 VSS.n4500 VSS.n4486 0.00681579
R8696 VSS.n3779 VSS.n3778 0.00680841
R8697 VSS.n4161 VSS.n4146 0.00679371
R8698 VSS.n4159 VSS.n4147 0.00679371
R8699 VSS.n4174 VSS.n788 0.00679371
R8700 VSS.n4181 VSS.n4180 0.00679371
R8701 VSS.n1686 VSS.n1680 0.00678492
R8702 VSS.n1693 VSS.n1692 0.00678492
R8703 VSS.n2929 VSS.n2928 0.00677907
R8704 VSS.n5792 VSS 0.00671127
R8705 VSS.n3358 VSS.n3357 0.00668497
R8706 VSS.n2551 VSS.n2421 0.00667143
R8707 VSS.n2038 VSS.n2016 0.00667057
R8708 VSS.n2711 VSS.n2710 0.00667057
R8709 VSS.n5827 VSS 0.00664458
R8710 VSS.n1869 VSS.n1868 0.00655172
R8711 VSS.n1333 VSS.n1332 0.00655042
R8712 VSS.n5898 VSS.n5896 0.00653659
R8713 VSS VSS.n5755 0.00652231
R8714 VSS.n1557 VSS.n1556 0.00651383
R8715 VSS.n1584 VSS.n1583 0.00651383
R8716 VSS.n1509 VSS.n1508 0.0065
R8717 VSS.n736 VSS.n735 0.0064434
R8718 VSS.n701 VSS.n511 0.0064434
R8719 VSS.n774 VSS.n773 0.0064434
R8720 VSS.n4313 VSS.n4312 0.0064434
R8721 VSS.n73 VSS.n72 0.00640164
R8722 VSS.n2019 VSS.n2018 0.00636957
R8723 VSS.n1644 VSS.n1582 0.00630645
R8724 VSS.n1642 VSS.n1607 0.00630645
R8725 VSS.n301 VSS.n300 0.00627982
R8726 VSS.n3602 VSS.n3601 0.00625581
R8727 VSS.n2573 VSS.n2571 0.00625581
R8728 VSS.n1979 VSS.n1978 0.00624138
R8729 VSS.n1974 VSS.n1968 0.00624138
R8730 VSS.n1964 VSS.n1958 0.00624138
R8731 VSS.n1954 VSS.n1953 0.00624138
R8732 VSS.n1932 VSS.n1931 0.00624138
R8733 VSS.n1911 VSS.n1906 0.00624138
R8734 VSS.n1402 VSS.n912 0.00622751
R8735 VSS.n2834 VSS.n2062 0.00618562
R8736 VSS.n1565 VSS.n1564 0.00617757
R8737 VSS.n3797 VSS.n3796 0.00617757
R8738 VSS.n3820 VSS.n3819 0.00617757
R8739 VSS.n3802 VSS.n3801 0.00617757
R8740 VSS.n3767 VSS.n3758 0.00617757
R8741 VSS.n3319 VSS.n3318 0.00616474
R8742 VSS.n4194 VSS.n4187 0.00616434
R8743 VSS.n960 VSS 0.006125
R8744 VSS.n291 VSS 0.006125
R8745 VSS.n4207 VSS 0.006125
R8746 VSS.n2168 VSS.n2162 0.00610386
R8747 VSS.n1975 VSS.n1974 0.00608621
R8748 VSS.n1965 VSS.n1964 0.00608621
R8749 VSS.n1957 VSS.n1956 0.00608621
R8750 VSS.n1955 VSS.n1954 0.00608621
R8751 VSS.n1912 VSS.n1911 0.00608621
R8752 VSS.n2875 VSS.n1993 0.00606856
R8753 VSS.n2870 VSS.n2869 0.00606856
R8754 VSS.n2865 VSS.n2008 0.00606856
R8755 VSS.n2035 VSS.n2011 0.00606856
R8756 VSS.n2063 VSS.n2050 0.00606856
R8757 VSS.n2794 VSS.n2087 0.00606856
R8758 VSS.n2785 VSS.n2092 0.00606856
R8759 VSS.n2768 VSS.n2767 0.00606856
R8760 VSS.n2728 VSS.n2197 0.00606856
R8761 VSS.n2718 VSS.n2210 0.00606856
R8762 VSS.n2713 VSS.n2712 0.00606856
R8763 VSS.n2661 VSS.n2310 0.00606856
R8764 VSS.n3651 VSS.n3650 0.00606522
R8765 VSS.n3506 VSS.n3505 0.00599419
R8766 VSS.n1822 VSS.n1821 0.00599419
R8767 VSS.n5092 VSS.n5091 0.00596961
R8768 VSS.n3788 VSS.n3787 0.00596729
R8769 VSS.n3789 VSS.n3785 0.00596729
R8770 VSS.n3752 VSS.n3743 0.00596729
R8771 VSS.n1884 VSS.n1883 0.00593103
R8772 VSS.n2881 VSS.n1993 0.00591806
R8773 VSS.n2870 VSS.n2000 0.00591806
R8774 VSS.n2866 VSS.n2865 0.00591806
R8775 VSS.n2862 VSS.n2861 0.00591806
R8776 VSS.n2860 VSS.n2011 0.00591806
R8777 VSS.n2806 VSS.n2087 0.00591806
R8778 VSS.n2791 VSS.n2092 0.00591806
R8779 VSS.n2780 VSS.n2099 0.00591806
R8780 VSS.n2728 VSS.n2196 0.00591806
R8781 VSS.n2724 VSS.n2210 0.00591806
R8782 VSS.n2713 VSS.n2217 0.00591806
R8783 VSS.n2692 VSS.n2244 0.00591806
R8784 VSS.n2273 VSS.n2267 0.0059088
R8785 VSS.n1621 VSS.n1620 0.0058917
R8786 VSS.n1633 VSS.n1632 0.0058917
R8787 VSS.n1675 VSS.n1674 0.00588013
R8788 VSS.n2933 VSS.n2932 0.00586337
R8789 VSS.n825 VSS.n789 0.00584965
R8790 VSS.n3434 VSS.n3433 0.00584884
R8791 VSS.n1873 VSS.n1872 0.00577586
R8792 VSS.n1870 VSS.n1869 0.00577586
R8793 VSS.n1867 VSS.n1866 0.00577586
R8794 VSS.n1864 VSS.n1862 0.00577586
R8795 VSS.n1854 VSS.n1853 0.00577586
R8796 VSS.n1879 VSS.n1878 0.00577586
R8797 VSS.n1973 VSS.n1972 0.00577586
R8798 VSS.n1963 VSS.n1962 0.00577586
R8799 VSS.n1886 VSS.n1885 0.00577586
R8800 VSS.n1895 VSS.n1894 0.00577586
R8801 VSS.n2040 VSS.n2036 0.00576756
R8802 VSS.n2223 VSS.n2220 0.00576756
R8803 VSS.n2873 VSS.n2872 0.00571739
R8804 VSS.n1617 VSS.n1616 0.00568433
R8805 VSS.n1629 VSS.n1628 0.00568433
R8806 VSS.n1871 VSS.n1870 0.00562069
R8807 VSS.n1868 VSS.n1867 0.00562069
R8808 VSS.n1865 VSS.n1864 0.00562069
R8809 VSS.n1908 VSS.n1907 0.00562069
R8810 VSS.n1971 VSS.n1970 0.00562069
R8811 VSS.n2879 VSS.n2878 0.00561706
R8812 VSS.n2018 VSS.n2017 0.00561706
R8813 VSS.n2020 VSS.n2015 0.00561706
R8814 VSS.n2856 VSS.n2016 0.00561706
R8815 VSS.n2068 VSS.n2047 0.00561706
R8816 VSS.n2877 VSS.n1994 0.00561706
R8817 VSS.n2004 VSS.n2002 0.00561706
R8818 VSS.n2014 VSS.n2007 0.00561706
R8819 VSS.n2031 VSS.n2013 0.00561706
R8820 VSS.n2067 VSS.n2048 0.00561706
R8821 VSS.n2143 VSS.n2142 0.00561706
R8822 VSS.n2789 VSS.n2788 0.00561706
R8823 VSS.n2138 VSS.n2137 0.00561706
R8824 VSS.n2753 VSS.n2129 0.00561706
R8825 VSS.n2787 VSS.n2093 0.00561706
R8826 VSS.n2117 VSS.n2115 0.00561706
R8827 VSS.n2722 VSS.n2721 0.00561706
R8828 VSS.n2231 VSS.n2230 0.00561706
R8829 VSS.n2720 VSS.n2211 0.00561706
R8830 VSS.n2221 VSS.n2219 0.00561706
R8831 VSS.n2925 VSS.n2924 0.00560174
R8832 VSS.n3828 VSS.n3827 0.00554673
R8833 VSS.n1455 VSS.n1444 0.00553496
R8834 VSS.n1462 VSS.n1461 0.00553496
R8835 VSS.n1521 VSS.n1514 0.00553496
R8836 VSS.n3894 VSS.n3893 0.00552326
R8837 VSS.n4690 VSS.n4689 0.0055
R8838 VSS.n84 VSS.n83 0.00547238
R8839 VSS.n3691 VSS.n3690 0.00547093
R8840 VSS.n2017 VSS.n1996 0.00546656
R8841 VSS.n2020 VSS.n2019 0.00546656
R8842 VSS.n2857 VSS.n2856 0.00546656
R8843 VSS.n2803 VSS.n2802 0.00546656
R8844 VSS.n2002 VSS.n2001 0.00546656
R8845 VSS.n2868 VSS.n2867 0.00546656
R8846 VSS.n2007 VSS.n2005 0.00546656
R8847 VSS.n2858 VSS.n2013 0.00546656
R8848 VSS.n2804 VSS.n2089 0.00546656
R8849 VSS.n2142 VSS.n2141 0.00546656
R8850 VSS.n2102 VSS.n2095 0.00546656
R8851 VSS.n2140 VSS.n2139 0.00546656
R8852 VSS.n2140 VSS.n2127 0.00546656
R8853 VSS.n2754 VSS.n2753 0.00546656
R8854 VSS.n2731 VSS.n2193 0.00546656
R8855 VSS.n2779 VSS.n2101 0.00546656
R8856 VSS.n2730 VSS.n2729 0.00546656
R8857 VSS.n2230 VSS.n2213 0.00546656
R8858 VSS.n2247 VSS.n2237 0.00546656
R8859 VSS.n2219 VSS.n2218 0.00546656
R8860 VSS.n2691 VSS.n2246 0.00546656
R8861 VSS.n1808 VSS.n1807 0.00546429
R8862 VSS.n2512 VSS.n2511 0.00541429
R8863 VSS.n4418 VSS.n4414 0.0053913
R8864 VSS.n3004 VSS.n3003 0.00538372
R8865 VSS.n2422 VSS.n2418 0.00534716
R8866 VSS.n2540 VSS.n2423 0.00534716
R8867 VSS.n3622 VSS.n3621 0.00534012
R8868 VSS.n3503 VSS.n3502 0.00534012
R8869 VSS.n3561 VSS.n3560 0.00534012
R8870 VSS.n3542 VSS.n3541 0.00534012
R8871 VSS.n1770 VSS.n1766 0.00534012
R8872 VSS.n3274 VSS.n3267 0.00534012
R8873 VSS.n3239 VSS.n3205 0.00534012
R8874 VSS.n3197 VSS.n3193 0.00534012
R8875 VSS.n3170 VSS.n3169 0.00534012
R8876 VSS.n3130 VSS.n3123 0.00534012
R8877 VSS.n3089 VSS.n3088 0.00534012
R8878 VSS.n3068 VSS.n3067 0.00534012
R8879 VSS.n1825 VSS.n1819 0.00534012
R8880 VSS.n3048 VSS.n3047 0.00534012
R8881 VSS.n3014 VSS.n3013 0.00534012
R8882 VSS.n2961 VSS.n2960 0.00534012
R8883 VSS.n2652 VSS.n2318 0.00534012
R8884 VSS.n2633 VSS.n2341 0.00534012
R8885 VSS.n2384 VSS.n2366 0.00534012
R8886 VSS.n2583 VSS.n2582 0.00534012
R8887 VSS.n3761 VSS.n3760 0.00533645
R8888 VSS.n3766 VSS.n3765 0.00533645
R8889 VSS.n3833 VSS.n3832 0.00533645
R8890 VSS.n3813 VSS.n3812 0.00533645
R8891 VSS.n297 VSS.n296 0.00532143
R8892 VSS.n359 VSS 0.00532143
R8893 VSS VSS.n4091 0.00532143
R8894 VSS VSS.n4129 0.00532143
R8895 VSS.n1810 VSS.n1809 0.00527273
R8896 VSS.n2562 VSS.n2411 0.00521616
R8897 VSS.n2548 VSS.n2423 0.00521616
R8898 VSS.n3684 VSS.n3670 0.0052093
R8899 VSS.n3622 VSS.n3576 0.0052093
R8900 VSS.n3439 VSS.n3438 0.0052093
R8901 VSS.n3444 VSS.n3443 0.0052093
R8902 VSS.n3566 VSS.n3447 0.0052093
R8903 VSS.n3543 VSS.n3542 0.0052093
R8904 VSS.n3413 VSS.n3362 0.0052093
R8905 VSS.n3413 VSS.n3366 0.0052093
R8906 VSS.n3274 VSS.n3263 0.0052093
R8907 VSS.n3239 VSS.n3201 0.0052093
R8908 VSS.n3115 VSS.n3114 0.0052093
R8909 VSS.n3068 VSS.n3056 0.0052093
R8910 VSS.n1818 VSS.n1817 0.0052093
R8911 VSS.n2961 VSS.n2918 0.0052093
R8912 VSS.n2658 VSS.n2318 0.0052093
R8913 VSS.n2325 VSS.n2324 0.0052093
R8914 VSS.n2583 VSS.n2565 0.0052093
R8915 VSS.n2757 VSS.n2125 0.00516555
R8916 VSS.n2164 VSS.n2144 0.00516555
R8917 VSS.n2748 VSS.n2747 0.00516555
R8918 VSS.n3749 VSS.n3747 0.00512617
R8919 VSS.n3750 VSS.n3746 0.00512617
R8920 VSS.n3817 VSS.n3816 0.00512617
R8921 VSS.n5276 VSS.n5275 0.00511538
R8922 VSS.n4372 VSS.n4371 0.00511538
R8923 VSS.n318 VSS.n265 0.00509184
R8924 VSS.n3593 VSS.n3592 0.00507849
R8925 VSS.n1572 VSS.n1571 0.00506221
R8926 VSS.n1592 VSS.n1591 0.00506221
R8927 VSS.n1602 VSS.n1601 0.00506221
R8928 VSS.n5896 VSS.n5895 0.00504545
R8929 VSS.n2124 VSS.n2118 0.00501505
R8930 VSS.n2752 VSS.n2128 0.00501505
R8931 VSS.n2764 VSS.n2763 0.00501505
R8932 VSS.n1952 VSS.n1951 0.005
R8933 VSS.n2428 VSS.n2426 0.00495415
R8934 VSS.n2544 VSS.n2543 0.00495415
R8935 VSS.n2427 VSS.n2416 0.00495415
R8936 VSS.n2542 VSS.n2425 0.00495415
R8937 VSS.n3595 VSS.n3594 0.00494767
R8938 VSS.n3604 VSS.n3603 0.00494767
R8939 VSS.n3717 VSS.n3716 0.00494767
R8940 VSS.n3721 VSS.n3720 0.00494767
R8941 VSS.n3498 VSS.n3497 0.00494767
R8942 VSS.n3526 VSS.n3525 0.00494767
R8943 VSS.n3517 VSS.n3516 0.00494767
R8944 VSS.n3514 VSS.n3513 0.00494767
R8945 VSS.n3455 VSS.n3454 0.00494767
R8946 VSS.n3489 VSS.n3488 0.00494767
R8947 VSS.n3475 VSS.n3474 0.00494767
R8948 VSS.n3470 VSS.n3469 0.00494767
R8949 VSS.n3441 VSS.n3440 0.00494767
R8950 VSS.n3547 VSS.n3546 0.00494767
R8951 VSS.n3406 VSS.n3405 0.00494767
R8952 VSS.n3403 VSS.n3402 0.00494767
R8953 VSS.n3382 VSS.n3381 0.00494767
R8954 VSS.n3412 VSS.n3411 0.00494767
R8955 VSS.n1769 VSS.n1768 0.00494767
R8956 VSS.n3273 VSS.n3272 0.00494767
R8957 VSS.n3232 VSS.n3231 0.00494767
R8958 VSS.n3229 VSS.n3228 0.00494767
R8959 VSS.n3219 VSS.n3218 0.00494767
R8960 VSS.n3075 VSS.n3074 0.00494767
R8961 VSS.n3079 VSS.n3078 0.00494767
R8962 VSS.n3238 VSS.n3237 0.00494767
R8963 VSS.n3196 VSS.n3195 0.00494767
R8964 VSS.n3165 VSS.n3164 0.00494767
R8965 VSS.n3129 VSS.n3128 0.00494767
R8966 VSS.n3110 VSS.n3109 0.00494767
R8967 VSS.n2924 VSS.n2923 0.00494767
R8968 VSS.n2928 VSS.n2927 0.00494767
R8969 VSS.n2932 VSS.n2931 0.00494767
R8970 VSS.n2943 VSS.n2942 0.00494767
R8971 VSS.n3063 VSS.n3062 0.00494767
R8972 VSS.n1824 VSS.n1823 0.00494767
R8973 VSS.n3044 VSS.n3043 0.00494767
R8974 VSS.n3011 VSS.n3010 0.00494767
R8975 VSS.n2656 VSS.n2655 0.00494767
R8976 VSS.n2642 VSS.n2331 0.00494767
R8977 VSS.n2630 VSS.n2346 0.00494767
R8978 VSS.n2572 VSS.n2389 0.00494767
R8979 VSS.n2654 VSS.n2319 0.00494767
R8980 VSS.n2632 VSS.n2631 0.00494767
R8981 VSS.n2388 VSS.n2364 0.00494767
R8982 VSS VSS.n922 0.00490559
R8983 VSS.n1431 VSS.n1428 0.00490559
R8984 VSS.n1437 VSS.n1434 0.00490559
R8985 VSS.n1443 VSS.n1440 0.00490559
R8986 VSS.n1475 VSS.n1472 0.00490559
R8987 VSS.n1500 VSS.n1497 0.00490559
R8988 VSS.n1494 VSS.n1491 0.00490559
R8989 VSS.n1488 VSS.n1485 0.00490559
R8990 VSS.n4013 VSS 0.00490559
R8991 VSS.n803 VSS.n800 0.00490559
R8992 VSS.n809 VSS.n806 0.00490559
R8993 VSS.n815 VSS.n812 0.00490559
R8994 VSS.n819 VSS.n818 0.00490559
R8995 VSS.n843 VSS.n840 0.00490559
R8996 VSS.n856 VSS.n853 0.00490559
R8997 VSS.n869 VSS.n866 0.00490559
R8998 VSS VSS.n4836 0.00490559
R8999 VSS VSS.n4799 0.00490559
R9000 VSS VSS.n4793 0.00490559
R9001 VSS VSS.n4911 0.00490559
R9002 VSS VSS.n4153 0.00490559
R9003 VSS.n322 VSS.n321 0.00489024
R9004 VSS.n2034 VSS.n2030 0.00486455
R9005 VSS.n1512 VSS.n1511 0.00486421
R9006 VSS.n1569 VSS.n1559 0.00485484
R9007 VSS.n1576 VSS.n1575 0.00485484
R9008 VSS.n1590 VSS.n1589 0.00485484
R9009 VSS.n1600 VSS.n1599 0.00485484
R9010 VSS.n2545 VSS.n2544 0.00482314
R9011 VSS.n2546 VSS.n2425 0.00482314
R9012 VSS.n3594 VSS.n3593 0.00481686
R9013 VSS.n3603 VSS.n3602 0.00481686
R9014 VSS.n3618 VSS.n3617 0.00481686
R9015 VSS.n3620 VSS.n3578 0.00481686
R9016 VSS.n3636 VSS.n3635 0.00481686
R9017 VSS.n3529 VSS.n3499 0.00481686
R9018 VSS.n3515 VSS.n3514 0.00481686
R9019 VSS.n3530 VSS.n3458 0.00481686
R9020 VSS.n3471 VSS.n3470 0.00481686
R9021 VSS.n3404 VSS.n3403 0.00481686
R9022 VSS.n3383 VSS.n3382 0.00481686
R9023 VSS.n3380 VSS.n3379 0.00481686
R9024 VSS.n3273 VSS.n3268 0.00481686
R9025 VSS.n3230 VSS.n3229 0.00481686
R9026 VSS.n3218 VSS.n3217 0.00481686
R9027 VSS.n3217 VSS.n3216 0.00481686
R9028 VSS.n3078 VSS.n3076 0.00481686
R9029 VSS.n3082 VSS.n3080 0.00481686
R9030 VSS.n2923 VSS.n2921 0.00481686
R9031 VSS.n2927 VSS.n2925 0.00481686
R9032 VSS.n2931 VSS.n2929 0.00481686
R9033 VSS.n2957 VSS.n2956 0.00481686
R9034 VSS.n3063 VSS.n3058 0.00481686
R9035 VSS.n3061 VSS.n3060 0.00481686
R9036 VSS.n2959 VSS.n2920 0.00481686
R9037 VSS.n2331 VSS.n2321 0.00481686
R9038 VSS.n2641 VSS.n2640 0.00481686
R9039 VSS.n2580 VSS.n2404 0.00481686
R9040 VSS.n2329 VSS.n2328 0.00481686
R9041 VSS.n2644 VSS.n2329 0.00481686
R9042 VSS.n2567 VSS.n2566 0.00481686
R9043 VSS.n2895 VSS.n2894 0.0048038
R9044 VSS.n3844 VSS.n3842 0.00476036
R9045 VSS.n3872 VSS.n3871 0.00476036
R9046 VSS.n3875 VSS.n3874 0.00476036
R9047 VSS.n2611 VSS.n2383 0.00474419
R9048 VSS.n2132 VSS.n2108 0.00471405
R9049 VSS.n2760 VSS.n2759 0.00471405
R9050 VSS.n1967 VSS.n1966 0.00468966
R9051 VSS.n3683 VSS.n3682 0.00468605
R9052 VSS.n3697 VSS.n3696 0.00468605
R9053 VSS.n3647 VSS.n3641 0.00468605
R9054 VSS.n3378 VSS.n3377 0.00468605
R9055 VSS.n3249 VSS.n3248 0.00468605
R9056 VSS.n3245 VSS.n3244 0.00468605
R9057 VSS.n3215 VSS.n3214 0.00468605
R9058 VSS.n2639 VSS.n2334 0.00468605
R9059 VSS.n2006 VSS.n2003 0.00456355
R9060 VSS.n2137 VSS.n2136 0.00456355
R9061 VSS.n2751 VSS.n2146 0.00456355
R9062 VSS.n1454 VSS.n1450 0.00456316
R9063 VSS.n2783 VSS.n2782 0.00455797
R9064 VSS.n3564 VSS.n3563 0.00455523
R9065 VSS.n2914 VSS.n2913 0.00444937
R9066 VSS.n2555 VSS.n2417 0.00443013
R9067 VSS.n3615 VSS.n3614 0.00442442
R9068 VSS.n3631 VSS.n3630 0.00442442
R9069 VSS.n3083 VSS.n3082 0.00442442
R9070 VSS.n2646 VSS.n2325 0.00442442
R9071 VSS.n2485 VSS.n2484 0.00429913
R9072 VSS.n2519 VSS.n2518 0.00429913
R9073 VSS.n3592 VSS.n3591 0.0042936
R9074 VSS.n3613 VSS.n3612 0.0042936
R9075 VSS.n1737 VSS.n1736 0.0042936
R9076 VSS.n3646 VSS.n3645 0.0042936
R9077 VSS.n3684 VSS.n3676 0.0042936
R9078 VSS.n3512 VSS.n3511 0.0042936
R9079 VSS.n3463 VSS.n3462 0.0042936
R9080 VSS.n3535 VSS.n3534 0.0042936
R9081 VSS.n3227 VSS.n3226 0.0042936
R9082 VSS.n3225 VSS.n3224 0.0042936
R9083 VSS.n3085 VSS.n3084 0.0042936
R9084 VSS.n3046 VSS.n3045 0.0042936
R9085 VSS.n2571 VSS.n2570 0.0042936
R9086 VSS.n2629 VSS.n2348 0.0042936
R9087 VSS.n2361 VSS.n2360 0.0042936
R9088 VSS.n2624 VSS.n2623 0.0042936
R9089 VSS.n2638 VSS.n2336 0.0042936
R9090 VSS.n2625 VSS.n2352 0.0042936
R9091 VSS.n2650 VSS.n2649 0.00427907
R9092 VSS.n826 VSS.n825 0.00427622
R9093 VSS.n850 VSS.n847 0.00427622
R9094 VSS.n2774 VSS.n2109 0.00426254
R9095 VSS.n3662 VSS.n3661 0.00416279
R9096 VSS.n3496 VSS.n3495 0.00416279
R9097 VSS.n3452 VSS.n3451 0.00416279
R9098 VSS.n92 VSS.n91 0.00414865
R9099 VSS.n2134 VSS.n2115 0.00411204
R9100 VSS.n2239 VSS.n2227 0.00411204
R9101 VSS.n3587 VSS.n3586 0.00403198
R9102 VSS.n3597 VSS.n3596 0.00403198
R9103 VSS.n3599 VSS.n3598 0.00403198
R9104 VSS.n3601 VSS.n3600 0.00403198
R9105 VSS.n3231 VSS.n3230 0.00403198
R9106 VSS.n3163 VSS.n3162 0.00403198
R9107 VSS.n3097 VSS.n3096 0.00403198
R9108 VSS.n3066 VSS.n3065 0.00403198
R9109 VSS.n2640 VSS.n2333 0.00403198
R9110 VSS.n2122 VSS.n2121 0.00397826
R9111 VSS.n4168 VSS.n4167 0.00396895
R9112 VSS.n5277 VSS.n5276 0.00396154
R9113 VSS.n2705 VSS.n2224 0.00396154
R9114 VSS.n2517 VSS.n2452 0.00390611
R9115 VSS.n2515 VSS.n2455 0.00390611
R9116 VSS.n3731 VSS.n3730 0.00390116
R9117 VSS.n1739 VSS.n1738 0.00390116
R9118 VSS.n3728 VSS.n3727 0.00390116
R9119 VSS.n1733 VSS.n1732 0.00390116
R9120 VSS.n3466 VSS.n3465 0.00390116
R9121 VSS.n3460 VSS.n3459 0.00390116
R9122 VSS.n3538 VSS.n3537 0.00390116
R9123 VSS.n3532 VSS.n3531 0.00390116
R9124 VSS.n1788 VSS.n1787 0.00390116
R9125 VSS.n1784 VSS.n1783 0.00390116
R9126 VSS.n2346 VSS.n2345 0.00390116
R9127 VSS.n2628 VSS.n2627 0.00390116
R9128 VSS.n2355 VSS.n2351 0.00390116
R9129 VSS.n2616 VSS.n2365 0.00390116
R9130 VSS.n2695 VSS.n2694 0.00389623
R9131 VSS.n3847 VSS.n3846 0.00381797
R9132 VSS.n3849 VSS.n3848 0.00381797
R9133 VSS.n3868 VSS.n3867 0.00381797
R9134 VSS.n3870 VSS.n3869 0.00381797
R9135 VSS.n2773 VSS.n2110 0.00381104
R9136 VSS.n2737 VSS.n2736 0.00381104
R9137 VSS.n3609 VSS.n3608 0.00377035
R9138 VSS.n3657 VSS.n3656 0.00377035
R9139 VSS.n3504 VSS.n3503 0.00377035
R9140 VSS.n3528 VSS.n3527 0.00377035
R9141 VSS.n3524 VSS.n3523 0.00377035
R9142 VSS.n3522 VSS.n3521 0.00377035
R9143 VSS.n3519 VSS.n3518 0.00377035
R9144 VSS.n3492 VSS.n3491 0.00377035
R9145 VSS.n3482 VSS.n3481 0.00377035
R9146 VSS.n5066 VSS.n5052 0.00371429
R9147 VSS.n3277 VSS.n3276 0.00367919
R9148 VSS.n3780 VSS.n3774 0.00367016
R9149 VSS.n3807 VSS.n3806 0.00367016
R9150 VSS.n2106 VSS.n2102 0.00366054
R9151 VSS.n2769 VSS.n2768 0.00366054
R9152 VSS.n2182 VSS.n2169 0.00366054
R9153 VSS.n2701 VSS.n2235 0.00366054
R9154 VSS.n2285 VSS.n2247 0.00366054
R9155 VSS.n2703 VSS.n2702 0.00366054
R9156 VSS.n4026 VSS.n4020 0.00364685
R9157 VSS.n4016 VSS.n4013 0.00364685
R9158 VSS.n2559 VSS.n2414 0.0036441
R9159 VSS.n2558 VSS.n2557 0.0036441
R9160 VSS.n3607 VSS.n3606 0.00363953
R9161 VSS.n3693 VSS.n3692 0.00363953
R9162 VSS.n3699 VSS.n3698 0.00363953
R9163 VSS.n3213 VSS.n3211 0.00363953
R9164 VSS.n3102 VSS.n3101 0.00363953
R9165 VSS.n2639 VSS.n2335 0.00363953
R9166 VSS.n3896 VSS.n3895 0.00356977
R9167 VSS.n3425 VSS.n3424 0.00352326
R9168 VSS.n2108 VSS.n2107 0.00351003
R9169 VSS.n2234 VSS.n2233 0.00351003
R9170 VSS.n2704 VSS.n2229 0.00351003
R9171 VSS.n2683 VSS.n2254 0.00351003
R9172 VSS.n2672 VSS.n2272 0.00351003
R9173 VSS.n1731 VSS.n1730 0.00350872
R9174 VSS.n3513 VSS.n3512 0.00350872
R9175 VSS.n3554 VSS.n3553 0.00350872
R9176 VSS.n3385 VSS.n3384 0.00350872
R9177 VSS.n2620 VSS.n2363 0.00350872
R9178 VSS.n2632 VSS.n2342 0.00350872
R9179 VSS.n2619 VSS.n2618 0.00350872
R9180 VSS.n3893 VSS.n3892 0.00347674
R9181 VSS.n732 VSS.n729 0.0034717
R9182 VSS.n504 VSS.n498 0.0034717
R9183 VSS.n770 VSS.n767 0.0034717
R9184 VSS.n4276 VSS.n4275 0.0034717
R9185 VSS.n4309 VSS.n4299 0.0034717
R9186 VSS.n1948 VSS.n1947 0.00344828
R9187 VSS.n2357 VSS.n2353 0.00340698
R9188 VSS.n3485 VSS.n3484 0.00337791
R9189 VSS.n3477 VSS.n3476 0.00337791
R9190 VSS.n3557 VSS.n3556 0.00337791
R9191 VSS.n3549 VSS.n3548 0.00337791
R9192 VSS.n2851 VSS.n2027 0.00335953
R9193 VSS.n2191 VSS.n2176 0.00335953
R9194 VSS.n2174 VSS.n2172 0.00335953
R9195 VSS.n2777 VSS.n2776 0.00335953
R9196 VSS.n3753 VSS.n3740 0.0032972
R9197 VSS.n3771 VSS.n3770 0.0032972
R9198 VSS.n3886 VSS.n3885 0.0032907
R9199 VSS.n3892 VSS.n3891 0.0032907
R9200 VSS.n3915 VSS.n3914 0.00327533
R9201 VSS.n3845 VSS.n3844 0.00324751
R9202 VSS.n3876 VSS.n3875 0.00324751
R9203 VSS.n3873 VSS.n3872 0.00324751
R9204 VSS.n3236 VSS.n3235 0.00324709
R9205 VSS.n3168 VSS.n3167 0.00324709
R9206 VSS.n2638 VSS.n2337 0.00324709
R9207 VSS.n1804 VSS.n1803 0.00322727
R9208 VSS.n2189 VSS.n2178 0.00320903
R9209 VSS.n2779 VSS.n2778 0.00320903
R9210 VSS.n2188 VSS.n2187 0.00320903
R9211 VSS.n2691 VSS.n2690 0.00320903
R9212 VSS.n3878 VSS.n3877 0.00319767
R9213 VSS.n3884 VSS.n3883 0.00319767
R9214 VSS.n3889 VSS.n3888 0.00319767
R9215 VSS.n2873 VSS.n1992 0.00317559
R9216 VSS.n2871 VSS.n1999 0.00317559
R9217 VSS.n2864 VSS.n2863 0.00317559
R9218 VSS.n2033 VSS.n2032 0.00317559
R9219 VSS.n2793 VSS.n2090 0.00317559
R9220 VSS.n3852 VSS.n3851 0.00317281
R9221 VSS.n3856 VSS.n3855 0.00317281
R9222 VSS.n3861 VSS.n3860 0.00317281
R9223 VSS.n3865 VSS.n3864 0.00317281
R9224 VSS.n4689 VSS.n4681 0.00316667
R9225 VSS.n3191 VSS.n3190 0.00315896
R9226 VSS.n878 VSS.n877 0.00313878
R9227 VSS.n1861 VSS.n1860 0.00313793
R9228 VSS.n1859 VSS.n1858 0.00313793
R9229 VSS.n1858 VSS.n1856 0.00313793
R9230 VSS.n1856 VSS.n1855 0.00313793
R9231 VSS.n1852 VSS.n1851 0.00313793
R9232 VSS.n1849 VSS.n1848 0.00313793
R9233 VSS.n1846 VSS.n1845 0.00313793
R9234 VSS.n1947 VSS.n1945 0.00313793
R9235 VSS.n1923 VSS.n1922 0.00313793
R9236 VSS.n2526 VSS.n2444 0.00312009
R9237 VSS.n3286 VSS.n3285 0.00311628
R9238 VSS.n3292 VSS.n3291 0.00311628
R9239 VSS.n3220 VSS.n3219 0.00311628
R9240 VSS.n3076 VSS.n3075 0.00311628
R9241 VSS.n3129 VSS.n3124 0.00311628
R9242 VSS.n2634 VSS.n2633 0.00311628
R9243 VSS.n2882 VSS.n1992 0.0031087
R9244 VSS.n2872 VSS.n2871 0.0031087
R9245 VSS.n2864 VSS.n2009 0.0031087
R9246 VSS.n2032 VSS.n2010 0.0031087
R9247 VSS.n2090 VSS.n2086 0.0031087
R9248 VSS.n3881 VSS.n3880 0.00310465
R9249 VSS.n2783 VSS.n2091 0.00307649
R9250 VSS.n2121 VSS.n2112 0.00307649
R9251 VSS.n2727 VSS.n2726 0.00307649
R9252 VSS.n2854 VSS.n2022 0.00305853
R9253 VSS.n2800 VSS.n2797 0.00305853
R9254 VSS.n2038 VSS.n2023 0.00305853
R9255 VSS.n2853 VSS.n2024 0.00305853
R9256 VSS.n2843 VSS.n2024 0.00305853
R9257 VSS.n2843 VSS.n2842 0.00305853
R9258 VSS.n2828 VSS.n2827 0.00305853
R9259 VSS.n2799 VSS.n2798 0.00305853
R9260 VSS.n2816 VSS.n2815 0.00305853
R9261 VSS.n2852 VSS.n2026 0.00305853
R9262 VSS.n2079 VSS.n2073 0.00305853
R9263 VSS.n2851 VSS.n2028 0.00305853
R9264 VSS.n2823 VSS.n2074 0.00305853
R9265 VSS.n2775 VSS.n2774 0.00305853
R9266 VSS.n2295 VSS.n2284 0.00305853
R9267 VSS.n2297 VSS.n2296 0.00305853
R9268 VSS.n2300 VSS.n2297 0.00305853
R9269 VSS.n2301 VSS.n2300 0.00305853
R9270 VSS.n2306 VSS.n2305 0.00305853
R9271 VSS.n2253 VSS.n2252 0.00305853
R9272 VSS.n2299 VSS.n2253 0.00305853
R9273 VSS.n2304 VSS.n2275 0.00305853
R9274 VSS.n2684 VSS.n2683 0.00305853
R9275 VSS.n3810 VSS.n3809 0.00301748
R9276 VSS.n3841 VSS.n3840 0.00301748
R9277 VSS.n2716 VSS.n2209 0.00301572
R9278 VSS.n2714 VSS.n2216 0.00301572
R9279 VSS.n2660 VSS.n2316 0.00301572
R9280 VSS.n2792 VSS.n2091 0.00301208
R9281 VSS.n2782 VSS.n2781 0.00301208
R9282 VSS.n2727 VSS.n2208 0.00301208
R9283 VSS.n2534 VSS.n2436 0.00298908
R9284 VSS.n3144 VSS.n3143 0.00298547
R9285 VSS.n3037 VSS.n3031 0.00298547
R9286 VSS.n2579 VSS.n2568 0.00298547
R9287 VSS.n2604 VSS.n2390 0.00298547
R9288 VSS.n2578 VSS.n2577 0.00298547
R9289 VSS.n2592 VSS.n2591 0.00298547
R9290 VSS.n2576 VSS.n2399 0.00298547
R9291 VSS.n2596 VSS.n2394 0.00298547
R9292 VSS.n1860 VSS.n1859 0.00298276
R9293 VSS.n1855 VSS.n1854 0.00298276
R9294 VSS.n1920 VSS.n1919 0.00298276
R9295 VSS.n4506 VSS.n4505 0.00297253
R9296 VSS.n5057 VSS.n5056 0.00297253
R9297 VSS.n2725 VSS.n2209 0.00295283
R9298 VSS.n2715 VSS.n2714 0.00295283
R9299 VSS.n2694 VSS.n2693 0.00295283
R9300 VSS.n3838 VSS.n3826 0.00292424
R9301 VSS.n2795 VSS.n2089 0.00292012
R9302 VSS.n2662 VSS.n2309 0.00292012
R9303 VSS.n2853 VSS.n2023 0.00290803
R9304 VSS.n2842 VSS.n2047 0.00290803
R9305 VSS.n2852 VSS.n2025 0.00290803
R9306 VSS.n2819 VSS.n2078 0.00290803
R9307 VSS.n2308 VSS.n2307 0.00290803
R9308 VSS.n2296 VSS.n2291 0.00290803
R9309 VSS.n2305 VSS.n2302 0.00290803
R9310 VSS.n2306 VSS.n2277 0.00290803
R9311 VSS.n2664 VSS.n2283 0.00290803
R9312 VSS.n2290 VSS.n2252 0.00290803
R9313 VSS.n2670 VSS.n2275 0.00290803
R9314 VSS.n2672 VSS.n2671 0.00290803
R9315 VSS.n2863 VSS.n2010 0.00290803
R9316 VSS.n3589 VSS.n3580 0.0028968
R9317 VSS.n3509 VSS.n3508 0.0028968
R9318 VSS.n3859 VSS.n3858 0.00289631
R9319 VSS.n3590 VSS.n3589 0.00289361
R9320 VSS.n3510 VSS.n3509 0.00289361
R9321 VSS.n299 VSS.n298 0.00287973
R9322 VSS.n3392 VSS.n3391 0.00285465
R9323 VSS.n3314 VSS.n3304 0.00285465
R9324 VSS.n2835 VSS.n2834 0.00284114
R9325 VSS.n4162 VSS.n889 0.00283689
R9326 VSS.n4708 VSS 0.00283333
R9327 VSS.n1924 VSS.n1923 0.00282759
R9328 VSS.n2650 VSS.n2317 0.00282558
R9329 VSS.n2353 VSS.n2338 0.00282558
R9330 VSS.n2584 VSS.n2564 0.00282558
R9331 VSS.n3069 VSS.n3054 0.00282558
R9332 VSS.n3052 VSS.n3051 0.00282558
R9333 VSS.n3049 VSS.n3041 0.00282558
R9334 VSS.n3015 VSS.n3004 0.00282558
R9335 VSS.n2962 VSS.n2916 0.00282558
R9336 VSS.n3435 VSS.n3434 0.00282558
R9337 VSS.n3423 VSS.n3422 0.00282558
R9338 VSS.n3623 VSS.n3574 0.00281884
R9339 VSS.n3240 VSS.n3200 0.00281214
R9340 VSS.n3198 VSS.n3191 0.00281214
R9341 VSS.n3171 VSS.n3158 0.00281214
R9342 VSS.n3131 VSS.n3118 0.00281214
R9343 VSS.n3090 VSS.n3072 0.00281214
R9344 VSS.n3359 VSS.n3358 0.00281214
R9345 VSS.n3275 VSS.n3262 0.00281214
R9346 VSS.n4374 VSS.n4372 0.00280769
R9347 VSS.n3087 VSS.n3086 0.00278682
R9348 VSS.n2552 VSS.n2551 0.00278571
R9349 VSS.n2538 VSS.n2433 0.00278571
R9350 VSS.n2659 VSS.n2317 0.00276744
R9351 VSS.n2649 VSS.n2648 0.00276744
R9352 VSS.n2585 VSS.n2584 0.00276744
R9353 VSS.n3070 VSS.n3069 0.00276744
R9354 VSS.n3053 VSS.n3052 0.00276744
R9355 VSS.n3050 VSS.n3049 0.00276744
R9356 VSS.n2963 VSS.n2962 0.00276744
R9357 VSS.n3573 VSS.n3572 0.00276744
R9358 VSS.n3572 VSS.n3571 0.00276744
R9359 VSS.n3570 VSS.n3569 0.00276744
R9360 VSS.n3568 VSS.n3567 0.00276744
R9361 VSS.n3424 VSS.n3423 0.00276744
R9362 VSS.n3723 VSS.n3722 0.00276087
R9363 VSS.n3686 VSS.n3685 0.00276087
R9364 VSS.n3624 VSS.n3623 0.00276087
R9365 VSS.n2824 VSS.n2823 0.00275752
R9366 VSS.n2780 VSS.n2100 0.00275752
R9367 VSS.n2692 VSS.n2245 0.00275752
R9368 VSS.n3241 VSS.n3240 0.00275434
R9369 VSS.n3199 VSS.n3198 0.00275434
R9370 VSS.n3117 VSS.n3116 0.00275434
R9371 VSS.n3415 VSS.n3414 0.00275434
R9372 VSS.n3276 VSS.n3275 0.00275434
R9373 VSS.n2563 VSS.n2410 0.00272857
R9374 VSS.n2433 VSS.n2421 0.00272857
R9375 VSS.n2484 VSS.n2439 0.00272707
R9376 VSS.n2531 VSS.n2430 0.00272707
R9377 VSS.n2450 VSS.n2440 0.00272707
R9378 VSS.n2527 VSS.n2442 0.00272707
R9379 VSS.n2497 VSS.n2496 0.00272707
R9380 VSS.n3468 VSS.n3467 0.00272384
R9381 VSS.n3130 VSS.n3119 0.00272384
R9382 VSS.n2934 VSS.n2933 0.00272384
R9383 VSS.n2938 VSS.n2936 0.00272384
R9384 VSS.n2939 VSS.n2938 0.00272384
R9385 VSS.n2940 VSS.n2939 0.00272384
R9386 VSS.n2945 VSS.n2944 0.00272384
R9387 VSS.n2950 VSS.n2948 0.00272384
R9388 VSS.n2954 VSS.n2953 0.00272384
R9389 VSS.n1980 VSS.n1979 0.00270985
R9390 VSS.n1456 VSS.n1455 0.0027028
R9391 VSS.n1456 VSS.n1417 0.0027028
R9392 VSS.n1462 VSS.n1417 0.0027028
R9393 VSS VSS.n1414 0.0027028
R9394 VSS VSS.n1414 0.0027028
R9395 VSS VSS.n835 0.0027028
R9396 VSS.n835 VSS 0.0027028
R9397 VSS.n2225 VSS.n2216 0.00270126
R9398 VSS.n729 VSS.n716 0.00269512
R9399 VSS.n4053 VSS.n4050 0.00269512
R9400 VSS.n2749 VSS.n2162 0.00269002
R9401 VSS.n1882 VSS.n1881 0.00267241
R9402 VSS.n1944 VSS.n1943 0.00267241
R9403 VSS.n1941 VSS.n1940 0.00267241
R9404 VSS.n1891 VSS.n1890 0.00267241
R9405 VSS.n1903 VSS.n1902 0.00267241
R9406 VSS.n1950 VSS.n1949 0.00267241
R9407 VSS.n1935 VSS.n1934 0.00267241
R9408 VSS.n1928 VSS.n1927 0.00267241
R9409 VSS.n1918 VSS.n1917 0.00267241
R9410 VSS.n4111 VSS.n908 0.00266
R9411 VSS.n3437 VSS.n3436 0.00265116
R9412 VSS.n3426 VSS.n3425 0.00265116
R9413 VSS.n2762 VSS.n2122 0.0026256
R9414 VSS.n2039 VSS.n2037 0.00260702
R9415 VSS.n2845 VSS.n2026 0.00260702
R9416 VSS.n2841 VSS.n2046 0.00260702
R9417 VSS.n2829 VSS.n2066 0.00260702
R9418 VSS.n2814 VSS.n2081 0.00260702
R9419 VSS.n2042 VSS.n2041 0.00260702
R9420 VSS.n2839 VSS.n2049 0.00260702
R9421 VSS.n2831 VSS.n2064 0.00260702
R9422 VSS.n2812 VSS.n2084 0.00260702
R9423 VSS.n2773 VSS.n2104 0.00260702
R9424 VSS.n2298 VSS.n2269 0.00260702
R9425 VSS.n2689 VSS.n2688 0.00260702
R9426 VSS.n2685 VSS.n2684 0.00260702
R9427 VSS.n2680 VSS.n2679 0.00260702
R9428 VSS.n2531 VSS.n2530 0.00259607
R9429 VSS.n2505 VSS.n2504 0.00259607
R9430 VSS.n2532 VSS.n2438 0.00259607
R9431 VSS.n2479 VSS.n2475 0.00259607
R9432 VSS.n2501 VSS.n2476 0.00259607
R9433 VSS.n2497 VSS.n2477 0.00259607
R9434 VSS.n3388 VSS.n3387 0.00259302
R9435 VSS.n3222 VSS.n3221 0.00259302
R9436 VSS.n3136 VSS.n3135 0.00259302
R9437 VSS.n2936 VSS.n2934 0.00259302
R9438 VSS.n2942 VSS.n2940 0.00259302
R9439 VSS.n3036 VSS.n3035 0.00259302
R9440 VSS.n2980 VSS.n2979 0.00259302
R9441 VSS.n2603 VSS.n2602 0.00259302
R9442 VSS.n2590 VSS.n2402 0.00259302
R9443 VSS.n2393 VSS.n2392 0.00259302
R9444 VSS.n2588 VSS.n2407 0.00259302
R9445 VSS.n3051 VSS.n3050 0.00259302
R9446 VSS.n3637 VSS.n3626 0.00258696
R9447 VSS.n3116 VSS.n3105 0.00258092
R9448 VSS.n3414 VSS.n3361 0.00258092
R9449 VSS.n2553 VSS.n2420 0.00255714
R9450 VSS.n5894 VSS.n4745 0.00254563
R9451 VSS.n1812 VSS.n1811 0.00254545
R9452 VSS.n3649 VSS.n3648 0.00252899
R9453 VSS.n2912 VSS.n2911 0.00252532
R9454 VSS.n2909 VSS.n2908 0.00252532
R9455 VSS.n2906 VSS.n2905 0.00252532
R9456 VSS.n2884 VSS.n2883 0.00252532
R9457 VSS.n3154 VSS.n3147 0.00252312
R9458 VSS.n3104 VSS.n3103 0.00252312
R9459 VSS.n3360 VSS.n3359 0.00252312
R9460 VSS.n3261 VSS.n3260 0.00252312
R9461 VSS.n3259 VSS.n3252 0.00252312
R9462 VSS.n3243 VSS.n3242 0.00252312
R9463 VSS.n1847 VSS.n1846 0.00251724
R9464 VSS.n1905 VSS.n1904 0.00251724
R9465 VSS.n2913 VSS.n2912 0.00247468
R9466 VSS.n2910 VSS.n2909 0.00247468
R9467 VSS.n2907 VSS.n2906 0.00247468
R9468 VSS.n2897 VSS.n2896 0.00247468
R9469 VSS.n2885 VSS.n2884 0.00247468
R9470 VSS.n3722 VSS.n3713 0.00247101
R9471 VSS.n3391 VSS.n3390 0.00246221
R9472 VSS.n3307 VSS.n3306 0.00246221
R9473 VSS.n3311 VSS.n3308 0.00246221
R9474 VSS.n3303 VSS.n3302 0.00246221
R9475 VSS.n3204 VSS.n3203 0.00246221
R9476 VSS.n2998 VSS.n2990 0.00246221
R9477 VSS.n2816 VSS.n2080 0.00245652
R9478 VSS.n2840 VSS.n2048 0.00245652
R9479 VSS.n2818 VSS.n2817 0.00245652
R9480 VSS.n2179 VSS.n2177 0.00245652
R9481 VSS.n2107 VSS.n2106 0.00245652
R9482 VSS.n2185 VSS.n2184 0.00245652
R9483 VSS.n2190 VSS.n2189 0.00245652
R9484 VSS.n2733 VSS.n2176 0.00245652
R9485 VSS.n2105 VSS.n2103 0.00245652
R9486 VSS.n2188 VSS.n2171 0.00245652
R9487 VSS.n2738 VSS.n2169 0.00245652
R9488 VSS.n2293 VSS.n2292 0.00245652
R9489 VSS.n2233 VSS.n2232 0.00245652
R9490 VSS.n2235 VSS.n2234 0.00245652
R9491 VSS.n2701 VSS.n2700 0.00245652
R9492 VSS.n2286 VSS.n2285 0.00245652
R9493 VSS.n2704 VSS.n2703 0.00245652
R9494 VSS.n2287 VSS.n2248 0.00245652
R9495 VSS.n2303 VSS.n2270 0.00245652
R9496 VSS.n2666 VSS.n2665 0.00245652
R9497 VSS.n2705 VSS.n2227 0.00245652
R9498 VSS.n2676 VSS.n2675 0.00245652
R9499 VSS.n2668 VSS.n2667 0.00245652
R9500 VSS.n2313 VSS.n2279 0.00245652
R9501 VSS.n5877 VSS.n5846 0.00244245
R9502 VSS.n5850 VSS.n5849 0.00244245
R9503 VSS.n5874 VSS.n5873 0.00244245
R9504 VSS.n5861 VSS.n5860 0.00244245
R9505 VSS.n2033 VSS.n2029 0.0024398
R9506 VSS VSS.n826 0.00238811
R9507 VSS.n1850 VSS.n1849 0.00236207
R9508 VSS.n3687 VSS.n3686 0.00235507
R9509 VSS.n2489 VSS.n2488 0.00233406
R9510 VSS.n2533 VSS.n2437 0.00233406
R9511 VSS.n2481 VSS.n2479 0.00233406
R9512 VSS.n2535 VSS.n2435 0.00233406
R9513 VSS.n3381 VSS.n3380 0.0023314
R9514 VSS.n3294 VSS.n3293 0.0023314
R9515 VSS.n3127 VSS.n3126 0.0023314
R9516 VSS.n3170 VSS.n3160 0.0023314
R9517 VSS.n3034 VSS.n3033 0.0023314
R9518 VSS.n3022 VSS.n3021 0.0023314
R9519 VSS.n2993 VSS.n2992 0.0023314
R9520 VSS.n2971 VSS.n2970 0.0023314
R9521 VSS.n3030 VSS.n3029 0.0023314
R9522 VSS.n2987 VSS.n2986 0.0023314
R9523 VSS.n2978 VSS.n2977 0.0023314
R9524 VSS.n2596 VSS.n2595 0.0023314
R9525 VSS.n2908 VSS.n2907 0.00232278
R9526 VSS.n2798 VSS.n2069 0.00230602
R9527 VSS.n2073 VSS.n2070 0.00230602
R9528 VSS.n2114 VSS.n2113 0.00230602
R9529 VSS.n2009 VSS.n1999 0.00230602
R9530 VSS.n2761 VSS.n2123 0.00230354
R9531 VSS.n3663 VSS.n3652 0.0022971
R9532 VSS.n2491 VSS.n2490 0.00224426
R9533 VSS.n2648 VSS.n2647 0.00224419
R9534 VSS.n5274 VSS.n5273 0.00224148
R9535 VSS.n1879 VSS.n1874 0.00222181
R9536 VSS.n1945 VSS.n1938 0.0022069
R9537 VSS.n2530 VSS.n2529 0.00220306
R9538 VSS.n2504 VSS.n2474 0.00220306
R9539 VSS.n2506 VSS.n2473 0.00220306
R9540 VSS.n2503 VSS.n2502 0.00220306
R9541 VSS.n2492 VSS.n2482 0.00220306
R9542 VSS.n2508 VSS.n2471 0.00220306
R9543 VSS.n3400 VSS.n3399 0.00220058
R9544 VSS.n3397 VSS.n3396 0.00220058
R9545 VSS.n3394 VSS.n3393 0.00220058
R9546 VSS.n3221 VSS.n3220 0.00220058
R9547 VSS.n3177 VSS.n3176 0.00220058
R9548 VSS.n3138 VSS.n3137 0.00220058
R9549 VSS.n2953 VSS.n2952 0.00220058
R9550 VSS.n3011 VSS.n3008 0.00220058
R9551 VSS.n2973 VSS.n2972 0.00220058
R9552 VSS.n2340 VSS.n2339 0.00220058
R9553 VSS.n2601 VSS.n2600 0.00220058
R9554 VSS.n1643 VSS.n1642 0.0022002
R9555 VSS.n2242 VSS.n2226 0.00219811
R9556 VSS.n2790 VSS.n2093 0.00219111
R9557 VSS.n2723 VSS.n2211 0.00219111
R9558 VSS.n2637 VSS.n2326 0.00218605
R9559 VSS.n2358 VSS.n2357 0.00218605
R9560 VSS.n2367 VSS.n2359 0.00218605
R9561 VSS.n2614 VSS.n2371 0.00218605
R9562 VSS.n3041 VSS.n3040 0.00218605
R9563 VSS.n3421 VSS.n3420 0.00218605
R9564 VSS.n3419 VSS.n3418 0.00218605
R9565 VSS.n3417 VSS.n3416 0.00218605
R9566 VSS.n3737 VSS.n3736 0.00218116
R9567 VSS.n3735 VSS.n3726 0.00218116
R9568 VSS.n3725 VSS.n3724 0.00218116
R9569 VSS.n3685 VSS.n3669 0.00218116
R9570 VSS.n3190 VSS.n3189 0.0021763
R9571 VSS.n3188 VSS.n3187 0.0021763
R9572 VSS.n5181 VSS.n5180 0.00216667
R9573 VSS.n5218 VSS.n4786 0.00216667
R9574 VSS.n5208 VSS.n5207 0.00216667
R9575 VSS.n5231 VSS.n5228 0.00216667
R9576 VSS.n2513 VSS.n2457 0.00215714
R9577 VSS.n2847 VSS.n2028 0.00215552
R9578 VSS.n2282 VSS.n2277 0.00215552
R9579 VSS.n5791 VSS.n5789 0.00214789
R9580 VSS.n6037 VSS.n6036 0.00214634
R9581 VSS.n2707 VSS.n2706 0.00213522
R9582 VSS.n3667 VSS.n3666 0.00212319
R9583 VSS.n3157 VSS.n3156 0.0021185
R9584 VSS.n2111 VSS.n2098 0.00211031
R9585 VSS.n2203 VSS.n2170 0.00211031
R9586 VSS.n2451 VSS.n2450 0.00207205
R9587 VSS.n3401 VSS.n3400 0.00206977
R9588 VSS.n3398 VSS.n3397 0.00206977
R9589 VSS.n3395 VSS.n3394 0.00206977
R9590 VSS.n3335 VSS.n3334 0.00206977
R9591 VSS.n2948 VSS.n2946 0.00206977
R9592 VSS.n2997 VSS.n2996 0.00206977
R9593 VSS.n3054 VSS.n3053 0.00206977
R9594 VSS.n3688 VSS.n3687 0.00206522
R9595 VSS.n2561 VSS.n2412 0.0020629
R9596 VSS.n3449 VSS.n3448 0.00206165
R9597 VSS.n3412 VSS.n3407 0.00206165
R9598 VSS.n3238 VSS.n3233 0.00206165
R9599 VSS.n2657 VSS.n2319 0.00206165
R9600 VSS.n1910 VSS.n1909 0.0020532
R9601 VSS.n1933 VSS.n1932 0.00205172
R9602 VSS.n2488 VSS.n2487 0.00204803
R9603 VSS.n2487 VSS.n2483 0.00204706
R9604 VSS.n2741 VSS.n2740 0.00204589
R9605 VSS.n2729 VSS.n2195 0.00202155
R9606 VSS.n2838 VSS.n2050 0.00200502
R9607 VSS.n2180 VSS.n2165 0.00200502
R9608 VSS.n2735 VSS.n2734 0.00200502
R9609 VSS.n2744 VSS.n2743 0.00200502
R9610 VSS.n2199 VSS.n2173 0.00200502
R9611 VSS.n2664 VSS.n2663 0.00200502
R9612 VSS.n2228 VSS.n2222 0.00200502
R9613 VSS.n2699 VSS.n2236 0.00200502
R9614 VSS.n2709 VSS.n2708 0.00200502
R9615 VSS.n2697 VSS.n2240 0.00200502
R9616 VSS.n2880 VSS.n1994 0.00199156
R9617 VSS.n2850 VSS.n2043 0.00197157
R9618 VSS.n2905 VSS.n2904 0.00196835
R9619 VSS.n3433 VSS.n3432 0.00195349
R9620 VSS.n1559 VSS.n1558 0.00195161
R9621 VSS.n1571 VSS.n1569 0.00195161
R9622 VSS.n1573 VSS.n1572 0.00195161
R9623 VSS.n1575 VSS.n1574 0.00195161
R9624 VSS.n1581 VSS.n1580 0.00195161
R9625 VSS.n1591 VSS.n1590 0.00195161
R9626 VSS.n1601 VSS.n1600 0.00195161
R9627 VSS.n2682 VSS.n2681 0.00194654
R9628 VSS.n2674 VSS.n2673 0.00194654
R9629 VSS.n3173 VSS.n3172 0.00194509
R9630 VSS.n3555 VSS.n3554 0.00193895
R9631 VSS.n3551 VSS.n3550 0.00193895
R9632 VSS.n3540 VSS.n3539 0.00193895
R9633 VSS.n3386 VSS.n3385 0.00193895
R9634 VSS.n3288 VSS.n3287 0.00193895
R9635 VSS.n3353 VSS.n3345 0.00193895
R9636 VSS.n3027 VSS.n3026 0.00193895
R9637 VSS.n2578 VSS.n2403 0.00193895
R9638 VSS.n2401 VSS.n2399 0.00193895
R9639 VSS.n2772 VSS.n2771 0.00191707
R9640 VSS.n5312 VSS.n5309 0.00189535
R9641 VSS.n5406 VSS.n5314 0.00189535
R9642 VSS.n3620 VSS.n3619 0.00188813
R9643 VSS.n2959 VSS.n2958 0.00188813
R9644 VSS.n2581 VSS.n2567 0.00188813
R9645 VSS.n3103 VSS.n3092 0.00188728
R9646 VSS.n2911 VSS.n2910 0.00186709
R9647 VSS.n356 VSS.n353 0.00185388
R9648 VSS.n2770 VSS.n2112 0.00185266
R9649 VSS.n3431 VSS.n3430 0.00183721
R9650 VSS.n3724 VSS.n3723 0.00183333
R9651 VSS.n3091 VSS.n3090 0.00182948
R9652 VSS.n3278 VSS.n3277 0.00182948
R9653 VSS.n4370 VSS.n4361 0.0018278
R9654 VSS.n2525 VSS.n2524 0.00181429
R9655 VSS.n2560 VSS.n2559 0.00181004
R9656 VSS.n2441 VSS.n2438 0.00181004
R9657 VSS.n3701 VSS.n3700 0.00180814
R9658 VSS.n3389 VSS.n3388 0.00180814
R9659 VSS.n3350 VSS.n3349 0.00180814
R9660 VSS.n3324 VSS.n3323 0.00180814
R9661 VSS.n3344 VSS.n3343 0.00180814
R9662 VSS.n3331 VSS.n3330 0.00180814
R9663 VSS.n3211 VSS.n3210 0.00180814
R9664 VSS.n3179 VSS.n3178 0.00180814
R9665 VSS.n3142 VSS.n3141 0.00180814
R9666 VSS.n3100 VSS.n3099 0.00180814
R9667 VSS.n3014 VSS.n3006 0.00180814
R9668 VSS.n2572 VSS.n2363 0.00180814
R9669 VSS.n2575 VSS.n2390 0.00180814
R9670 VSS.n2395 VSS.n2391 0.00180814
R9671 VSS.n2612 VSS.n2611 0.00177907
R9672 VSS.n3039 VSS.n3038 0.00177907
R9673 VSS.n3428 VSS.n3427 0.00177907
R9674 VSS.n3133 VSS.n3132 0.00177168
R9675 VSS.n3299 VSS.n3296 0.00177168
R9676 VSS.n2820 VSS.n2077 0.0017709
R9677 VSS.n3760 VSS.n3759 0.00176168
R9678 VSS.n3836 VSS.n3829 0.00176168
R9679 VSS.n1513 VSS.n1405 0.00175874
R9680 VSS.n2536 VSS.n2434 0.00175714
R9681 VSS.n1579 VSS.n1577 0.00174752
R9682 VSS.n1619 VSS.n1618 0.00174424
R9683 VSS.n1631 VSS.n1630 0.00174424
R9684 VSS.n2637 VSS.n2636 0.00172093
R9685 VSS.n3712 VSS.n3711 0.00171739
R9686 VSS.n3158 VSS.n3157 0.00171387
R9687 VSS.n2670 VSS.n2669 0.00170401
R9688 VSS.n2822 VSS.n2076 0.00170401
R9689 VSS.n2312 VSS.n2311 0.00169497
R9690 VSS.n2426 VSS.n2414 0.00167904
R9691 VSS.n2521 VSS.n2449 0.00167904
R9692 VSS.n3584 VSS.n3583 0.00167733
R9693 VSS.n3606 VSS.n3605 0.00167733
R9694 VSS.n3608 VSS.n3607 0.00167733
R9695 VSS.n3610 VSS.n3609 0.00167733
R9696 VSS.n3709 VSS.n3705 0.00167733
R9697 VSS.n3529 VSS.n3528 0.00167733
R9698 VSS.n3396 VSS.n3395 0.00167733
R9699 VSS.n3348 VSS.n3347 0.00167733
R9700 VSS.n3328 VSS.n3327 0.00167733
R9701 VSS.n3326 VSS.n3325 0.00167733
R9702 VSS.n3342 VSS.n3341 0.00167733
R9703 VSS.n3333 VSS.n3332 0.00167733
R9704 VSS.n2635 VSS.n2338 0.00166279
R9705 VSS.n2771 VSS.n2770 0.00165942
R9706 VSS.n2161 VSS.n2160 0.00165942
R9707 VSS.n3316 VSS.n3315 0.00165607
R9708 VSS.n2498 VSS.n2478 0.00164286
R9709 VSS.n2043 VSS.n2029 0.00163712
R9710 VSS.n2850 VSS.n2849 0.00163712
R9711 VSS.n2837 VSS.n2044 0.00163712
R9712 VSS.n2075 VSS.n2062 0.00163712
R9713 VSS.n2822 VSS.n2821 0.00163712
R9714 VSS.n2810 VSS.n2077 0.00163712
R9715 VSS.n3749 VSS.n3748 0.00163084
R9716 VSS.n2903 VSS.n2902 0.00161392
R9717 VSS.n188 VSS.n187 0.00161111
R9718 VSS.n218 VSS.n215 0.00161111
R9719 VSS.n205 VSS.n194 0.00161111
R9720 VSS.n195 VSS.n123 0.00161111
R9721 VSS.n2636 VSS.n2635 0.00160465
R9722 VSS.n2397 VSS.n2396 0.00160465
R9723 VSS.n2598 VSS.n2597 0.00160465
R9724 VSS.n2586 VSS.n2409 0.00160465
R9725 VSS.n2981 VSS.n2966 0.00160465
R9726 VSS.n3710 VSS.n3703 0.00160145
R9727 VSS.n4315 VSS.n4313 0.00159756
R9728 VSS.n2500 VSS.n2469 0.00158571
R9729 VSS.n2687 VSS.n2243 0.00156918
R9730 VSS.n2681 VSS.n2267 0.00156918
R9731 VSS.n2283 VSS.n2282 0.00155351
R9732 VSS.n2280 VSS.n2278 0.00155351
R9733 VSS.n2309 VSS.n2281 0.00155351
R9734 VSS.n3746 VSS.n3745 0.0015514
R9735 VSS.n3816 VSS.n3815 0.0015514
R9736 VSS.n3818 VSS.n3817 0.0015514
R9737 VSS.n3824 VSS.n3814 0.0015514
R9738 VSS.n2522 VSS.n2448 0.00154803
R9739 VSS.n1742 VSS.n1734 0.00154651
R9740 VSS.n3527 VSS.n3526 0.00154651
R9741 VSS.n3523 VSS.n3522 0.00154651
R9742 VSS.n3483 VSS.n3482 0.00154651
R9743 VSS.n3534 VSS.n3533 0.00154651
R9744 VSS.n3405 VSS.n3404 0.00154651
R9745 VSS.n3399 VSS.n3398 0.00154651
R9746 VSS.n3390 VSS.n3389 0.00154651
R9747 VSS.n3352 VSS.n3351 0.00154651
R9748 VSS.n3271 VSS.n3270 0.00154651
R9749 VSS.n3080 VSS.n3079 0.00154651
R9750 VSS.n3186 VSS.n3185 0.00154651
R9751 VSS.n3122 VSS.n3121 0.00154651
R9752 VSS.n2613 VSS.n2612 0.00154651
R9753 VSS.n3000 VSS.n2999 0.00154651
R9754 VSS.n3318 VSS.n3317 0.00154046
R9755 VSS.n1587 VSS.n1586 0.00153687
R9756 VSS.n1589 VSS.n1588 0.00153687
R9757 VSS.n1597 VSS.n1596 0.00153687
R9758 VSS.n1599 VSS.n1598 0.00153687
R9759 VSS.n1607 VSS.n1606 0.00153687
R9760 VSS.n2674 VSS.n2273 0.00150629
R9761 VSS.n2673 VSS.n2274 0.00150629
R9762 VSS.n2315 VSS.n2312 0.00150629
R9763 VSS.n1694 VSS.n1693 0.00150559
R9764 VSS.n1699 VSS.n1698 0.00150559
R9765 VSS.n1704 VSS.n1703 0.00150559
R9766 VSS.n1706 VSS.n1705 0.00150559
R9767 VSS.n2597 VSS.n2398 0.00148837
R9768 VSS.n3040 VSS.n3039 0.00148837
R9769 VSS.n3038 VSS.n3028 0.00148837
R9770 VSS.n3017 VSS.n3016 0.00148837
R9771 VSS.n3002 VSS.n3001 0.00148837
R9772 VSS.n2999 VSS.n2984 0.00148837
R9773 VSS.n2966 VSS.n2965 0.00148837
R9774 VSS.n3132 VSS.n3131 0.00148266
R9775 VSS.n3295 VSS.n3278 0.00148266
R9776 VSS.n2537 VSS.n2536 0.00147143
R9777 VSS.n2781 VSS.n2098 0.00146618
R9778 VSS.n2889 VSS.n2888 0.00146203
R9779 VSS.n1654 VSS.n1651 0.00145031
R9780 VSS.n1685 VSS.n1682 0.00144995
R9781 VSS.n1685 VSS.n1684 0.00144995
R9782 VSS.n1654 VSS.n1653 0.0014496
R9783 VSS VSS.n820 0.00144406
R9784 VSS.n2693 VSS.n2243 0.0014434
R9785 VSS.n2266 VSS.n2250 0.0014434
R9786 VSS.n1937 VSS.n1936 0.00143104
R9787 VSS.n2599 VSS.n2397 0.00143023
R9788 VSS.n3092 VSS.n3091 0.00142485
R9789 VSS.n3300 VSS.n3299 0.00142485
R9790 VSS.n2415 VSS.n2412 0.00141703
R9791 VSS.n2445 VSS.n2436 0.00141703
R9792 VSS.n2526 VSS.n2443 0.00141703
R9793 VSS.n3600 VSS.n3599 0.0014157
R9794 VSS.n3695 VSS.n3694 0.0014157
R9795 VSS.n3734 VSS.n3729 0.0014157
R9796 VSS.n3536 VSS.n3535 0.0014157
R9797 VSS.n3387 VSS.n3386 0.0014157
R9798 VSS.n1791 VSS.n1785 0.0014157
R9799 VSS.n2345 VSS.n2333 0.0014157
R9800 VSS.n2344 VSS.n2343 0.0014157
R9801 VSS.n2617 VSS.n2364 0.0014157
R9802 VSS.n2626 VSS.n2625 0.0014157
R9803 VSS.n2510 VSS.n2469 0.00141429
R9804 VSS.n2499 VSS.n2498 0.00141429
R9805 VSS.n2892 VSS.n2891 0.00141139
R9806 VSS.n2846 VSS.n2045 0.00140301
R9807 VSS.n2136 VSS.n2132 0.00140301
R9808 VSS.n2135 VSS.n2133 0.00140301
R9809 VSS.n2772 VSS.n2111 0.00140177
R9810 VSS.n1554 VSS.n1545 0.0014
R9811 VSS.n1552 VSS.n1547 0.0014
R9812 VSS.n1551 VSS.n1549 0.0014
R9813 VSS.n1667 VSS.n1666 0.0014
R9814 VSS.n1689 VSS.n1688 0.0014
R9815 VSS.n1659 VSS.n1658 0.0014
R9816 VSS.n1677 VSS.n1675 0.0014
R9817 VSS.n1727 VSS.n1726 0.0014
R9818 VSS.n1725 VSS.n1723 0.0014
R9819 VSS.n1561 VSS.n1560 0.0014
R9820 VSS.n1541 VSS.n1539 0.0014
R9821 VSS.n1542 VSS.n1537 0.0014
R9822 VSS.n1544 VSS.n1535 0.0014
R9823 VSS.n2686 VSS.n2250 0.0013805
R9824 VSS.n3429 VSS.n3428 0.00137209
R9825 VSS.n3200 VSS.n3199 0.00136705
R9826 VSS.n3336 VSS.n3321 0.00136705
R9827 VSS.n2904 VSS.n2903 0.00136076
R9828 VSS.n2902 VSS.n2901 0.00136076
R9829 VSS.n2899 VSS.n2898 0.00136076
R9830 VSS.n2894 VSS.n2893 0.00136076
R9831 VSS.n2891 VSS.n2890 0.00136076
R9832 VSS.n2888 VSS.n2887 0.00136076
R9833 VSS.n3765 VSS.n3764 0.00134112
R9834 VSS.n3763 VSS.n3762 0.00134112
R9835 VSS.n3834 VSS.n3833 0.00134112
R9836 VSS.n3743 VSS.n3742 0.00134112
R9837 VSS.n3812 VSS.n3811 0.00134112
R9838 VSS.n3814 VSS.n3813 0.00134112
R9839 VSS.n3825 VSS.n3810 0.00133916
R9840 VSS.n3840 VSS.n3839 0.00133916
R9841 VSS.n2742 VSS.n2168 0.00133736
R9842 VSS.n2740 VSS.n2739 0.00133736
R9843 VSS.n2204 VSS.n2203 0.00133736
R9844 VSS.n1614 VSS.n1613 0.00132949
R9845 VSS.n1616 VSS.n1615 0.00132949
R9846 VSS.n1623 VSS.n1622 0.00132949
R9847 VSS.n1626 VSS.n1625 0.00132949
R9848 VSS.n1628 VSS.n1627 0.00132949
R9849 VSS.n1635 VSS.n1634 0.00132949
R9850 VSS.n1638 VSS.n1637 0.00132949
R9851 VSS.n1585 VSS.n1584 0.00132949
R9852 VSS.n1593 VSS.n1592 0.00132949
R9853 VSS.n1595 VSS.n1594 0.00132949
R9854 VSS.n1603 VSS.n1602 0.00132949
R9855 VSS.n1605 VSS.n1604 0.00132949
R9856 VSS.n2707 VSS.n2225 0.00131761
R9857 VSS.n2706 VSS.n2226 0.00131761
R9858 VSS.n2695 VSS.n2242 0.00131761
R9859 VSS.n3432 VSS.n3431 0.00131395
R9860 VSS.n3172 VSS.n3171 0.00130925
R9861 VSS.n3355 VSS.n3354 0.00130925
R9862 VSS.n2848 VSS.n2044 0.00130268
R9863 VSS.n2556 VSS.n2416 0.00128603
R9864 VSS.n2523 VSS.n2522 0.00128603
R9865 VSS.n3596 VSS.n3595 0.00128488
R9866 VSS.n3598 VSS.n3597 0.00128488
R9867 VSS.n3708 VSS.n3707 0.00128488
R9868 VSS.n3655 VSS.n3654 0.00128488
R9869 VSS.n3660 VSS.n3659 0.00128488
R9870 VSS.n3495 VSS.n3494 0.00128488
R9871 VSS.n3530 VSS.n3493 0.00128488
R9872 VSS.n3025 VSS.n3024 0.00128488
R9873 VSS.n2621 VSS.n2620 0.00128488
R9874 VSS.n5514 VSS.n5463 0.00127586
R9875 VSS.n1680 VSS.n1679 0.00125419
R9876 VSS.n1695 VSS.n1694 0.00125419
R9877 VSS.n1700 VSS.n1699 0.00125419
R9878 VSS.n1702 VSS.n1701 0.00125419
R9879 VSS.n1711 VSS.n1710 0.00125419
R9880 VSS.n1712 VSS.n1711 0.00125419
R9881 VSS.n1714 VSS.n1713 0.00125419
R9882 VSS.n1716 VSS.n1715 0.00125419
R9883 VSS.n1718 VSS.n1717 0.00125419
R9884 VSS.n3904 VSS.n3903 0.00125419
R9885 VSS.n3908 VSS.n1687 0.00125419
R9886 VSS.n3702 VSS.n3688 0.00125362
R9887 VSS.n2671 VSS.n2276 0.00125251
R9888 VSS.n3134 VSS.n3133 0.00125145
R9889 VSS.n3356 VSS.n3355 0.00125145
R9890 VSS.n3339 VSS.n3336 0.00125145
R9891 VSS.n3320 VSS.n3319 0.00125145
R9892 VSS.n2849 VSS.n2848 0.00123579
R9893 VSS.n5883 VSS.n5882 0.0012013
R9894 VSS.n5879 VSS.n5878 0.0012013
R9895 VSS.n3018 VSS.n3017 0.00119767
R9896 VSS.n3711 VSS.n3710 0.00119565
R9897 VSS.n3357 VSS.n3356 0.00119364
R9898 VSS.n3354 VSS.n3339 0.00119364
R9899 VSS.n3321 VSS.n3320 0.00119364
R9900 VSS.n2837 VSS.n2836 0.0011689
R9901 VSS.n2519 VSS.n2451 0.00115502
R9902 VSS.n2521 VSS.n2520 0.00115502
R9903 VSS.n3591 VSS.n3590 0.00115407
R9904 VSS.n1741 VSS.n1740 0.00115407
R9905 VSS.n3675 VSS.n3674 0.00115407
R9906 VSS.n3497 VSS.n3496 0.00115407
R9907 VSS.n3520 VSS.n3519 0.00115407
R9908 VSS.n3508 VSS.n3507 0.00115407
R9909 VSS.n3490 VSS.n3489 0.00115407
R9910 VSS.n3479 VSS.n3478 0.00115407
R9911 VSS.n3462 VSS.n3461 0.00115407
R9912 VSS.n3311 VSS.n3310 0.00115407
R9913 VSS.n3224 VSS.n3222 0.00115407
R9914 VSS.n3181 VSS.n3180 0.00115407
R9915 VSS.n2621 VSS.n2361 0.00115407
R9916 VSS.n2623 VSS.n2622 0.00115407
R9917 VSS.n2369 VSS.n2352 0.00115407
R9918 VSS.n3879 VSS.n3878 0.00115116
R9919 VSS.n3883 VSS.n3882 0.00115116
R9920 VSS.n3851 VSS.n3850 0.00114516
R9921 VSS.n3857 VSS.n3856 0.00114516
R9922 VSS.n3860 VSS.n3859 0.00114516
R9923 VSS.n3866 VSS.n3865 0.00114516
R9924 VSS.n3028 VSS.n3018 0.00113953
R9925 VSS.n3422 VSS.n3421 0.00113953
R9926 VSS.n3418 VSS.n3417 0.00113953
R9927 VSS.n3726 VSS.n3725 0.00113768
R9928 VSS.n3187 VSS.n3174 0.00113584
R9929 VSS.n3784 VSS.n3783 0.00113084
R9930 VSS.n3758 VSS.n3757 0.00113084
R9931 VSS.n3757 VSS.n3756 0.00113084
R9932 VSS.n3756 VSS.n3755 0.00113084
R9933 VSS.n3829 VSS.n3828 0.00113084
R9934 VSS.n1501 VSS.n1500 0.00112937
R9935 VSS.n847 VSS.n846 0.00112937
R9936 VSS.n2457 VSS.n2447 0.00112857
R9937 VSS.n1612 VSS.n1611 0.00112212
R9938 VSS.n1615 VSS.n1614 0.00112212
R9939 VSS.n1622 VSS.n1621 0.00112212
R9940 VSS.n1624 VSS.n1623 0.00112212
R9941 VSS.n1627 VSS.n1626 0.00112212
R9942 VSS.n1634 VSS.n1633 0.00112212
R9943 VSS.n1636 VSS.n1635 0.00112212
R9944 VSS.n1594 VSS.n1593 0.00112212
R9945 VSS.n1604 VSS.n1603 0.00112212
R9946 VSS.n1851 VSS.n1850 0.00112069
R9947 VSS.n1848 VSS.n1847 0.00112069
R9948 VSS.n1845 VSS.n1844 0.00112069
R9949 VSS.n1922 VSS.n1920 0.00112069
R9950 VSS.n2900 VSS.n2899 0.00110759
R9951 VSS.n2801 VSS.n2800 0.00110201
R9952 VSS.n2827 VSS.n2069 0.00110201
R9953 VSS.n2799 VSS.n2080 0.00110201
R9954 VSS.n2815 VSS.n2082 0.00110201
R9955 VSS.n2818 VSS.n2079 0.00110201
R9956 VSS.n2819 VSS.n2074 0.00110201
R9957 VSS.n2145 VSS.n2126 0.00110201
R9958 VSS.n2291 VSS.n2286 0.00110201
R9959 VSS.n2314 VSS.n2310 0.00110201
R9960 VSS.n2647 VSS.n2326 0.0010814
R9961 VSS.n2359 VSS.n2358 0.0010814
R9962 VSS.n3016 VSS.n3015 0.0010814
R9963 VSS.n3420 VSS.n3419 0.0010814
R9964 VSS.n2750 VSS.n2161 0.00107971
R9965 VSS.n3736 VSS.n3735 0.00107971
R9966 VSS.n3189 VSS.n3188 0.00107803
R9967 VSS.n2525 VSS.n2446 0.00107143
R9968 VSS.n3740 VSS.n3739 0.00105944
R9969 VSS.n3772 VSS.n3771 0.00105944
R9970 VSS.n3887 VSS.n3886 0.00105814
R9971 VSS.n3891 VSS.n3890 0.00105814
R9972 VSS.n2901 VSS.n2900 0.00105696
R9973 VSS.n3854 VSS.n3853 0.00105299
R9974 VSS.n3863 VSS.n3862 0.00105299
R9975 VSS.n2529 VSS.n2440 0.00102402
R9976 VSS.n2505 VSS.n2453 0.00102402
R9977 VSS.n2483 VSS.n2474 0.00102402
R9978 VSS.n2493 VSS.n2489 0.00102402
R9979 VSS.n2528 VSS.n2527 0.00102402
R9980 VSS.n2502 VSS.n2475 0.00102402
R9981 VSS.n2419 VSS.n2411 0.00102402
R9982 VSS.n2501 VSS.n2477 0.00102402
R9983 VSS.n3582 VSS.n3581 0.00102326
R9984 VSS.n3580 VSS.n3579 0.00102326
R9985 VSS.n3612 VSS.n3611 0.00102326
R9986 VSS.n3614 VSS.n3613 0.00102326
R9987 VSS.n3616 VSS.n3615 0.00102326
R9988 VSS.n3733 VSS.n3732 0.00102326
R9989 VSS.n3679 VSS.n3678 0.00102326
R9990 VSS.n3521 VSS.n3520 0.00102326
R9991 VSS.n3511 VSS.n3510 0.00102326
R9992 VSS.n3464 VSS.n3463 0.00102326
R9993 VSS.n3288 VSS.n3282 0.00102326
R9994 VSS.n3226 VSS.n3225 0.00102326
R9995 VSS.n3084 VSS.n3083 0.00102326
R9996 VSS.n1790 VSS.n1789 0.00102326
R9997 VSS.n3095 VSS.n3094 0.00102326
R9998 VSS.n3184 VSS.n3183 0.00102326
R9999 VSS.n2946 VSS.n2945 0.00102326
R10000 VSS.n2952 VSS.n2950 0.00102326
R10001 VSS.n2955 VSS.n2954 0.00102326
R10002 VSS.n2574 VSS.n2568 0.00102326
R10003 VSS.n2360 VSS.n2348 0.00102326
R10004 VSS.n2605 VSS.n2604 0.00102326
R10005 VSS.n2577 VSS.n2575 0.00102326
R10006 VSS.n2592 VSS.n2403 0.00102326
R10007 VSS.n2624 VSS.n2350 0.00102326
R10008 VSS.n2576 VSS.n2395 0.00102326
R10009 VSS.n2645 VSS.n2327 0.00102326
R10010 VSS.n2615 VSS.n2366 0.00102326
R10011 VSS.n2600 VSS.n2394 0.00102326
R10012 VSS.n3669 VSS.n3668 0.00102174
R10013 VSS.n3666 VSS.n3663 0.00102174
R10014 VSS.n3652 VSS.n3651 0.00102174
R10015 VSS.n2898 VSS.n2897 0.00100633
R10016 VSS.n2687 VSS.n2686 0.00100314
R10017 VSS.n1670 VSS.n1669 0.00100279
R10018 VSS.n1707 VSS.n1706 0.00100279
R10019 VSS.n3902 VSS.n3898 0.00100279
R10020 VSS VSS.n5880 0.000967532
R10021 VSS.n3769 VSS.n3754 0.0009662
R10022 VSS.n1878 VSS.n1877 0.000965517
R10023 VSS.n1876 VSS.n1875 0.000965517
R10024 VSS.n1972 VSS.n1971 0.000965517
R10025 VSS.n1970 VSS.n1969 0.000965517
R10026 VSS.n1962 VSS.n1961 0.000965517
R10027 VSS.n1960 VSS.n1959 0.000965517
R10028 VSS.n1885 VSS.n1884 0.000965517
R10029 VSS.n1883 VSS.n1882 0.000965517
R10030 VSS.n1881 VSS.n1880 0.000965517
R10031 VSS.n1943 VSS.n1942 0.000965517
R10032 VSS.n1942 VSS.n1941 0.000965517
R10033 VSS.n1940 VSS.n1939 0.000965517
R10034 VSS.n1894 VSS.n1893 0.000965517
R10035 VSS.n1892 VSS.n1891 0.000965517
R10036 VSS.n1890 VSS.n1889 0.000965517
R10037 VSS.n1888 VSS.n1887 0.000965517
R10038 VSS.n1904 VSS.n1903 0.000965517
R10039 VSS.n1902 VSS.n1901 0.000965517
R10040 VSS.n1900 VSS.n1899 0.000965517
R10041 VSS.n1898 VSS.n1897 0.000965517
R10042 VSS.n1978 VSS.n1977 0.000965517
R10043 VSS.n1976 VSS.n1975 0.000965517
R10044 VSS.n1968 VSS.n1967 0.000965517
R10045 VSS.n1966 VSS.n1965 0.000965517
R10046 VSS.n1958 VSS.n1957 0.000965517
R10047 VSS.n1956 VSS.n1955 0.000965517
R10048 VSS.n1953 VSS.n1952 0.000965517
R10049 VSS.n1951 VSS.n1950 0.000965517
R10050 VSS.n1949 VSS.n1948 0.000965517
R10051 VSS.n1938 VSS.n1937 0.000965517
R10052 VSS.n1936 VSS.n1935 0.000965517
R10053 VSS.n1934 VSS.n1933 0.000965517
R10054 VSS.n1931 VSS.n1930 0.000965517
R10055 VSS.n1929 VSS.n1928 0.000965517
R10056 VSS.n1927 VSS.n1926 0.000965517
R10057 VSS.n1925 VSS.n1924 0.000965517
R10058 VSS.n1919 VSS.n1918 0.000965517
R10059 VSS.n1917 VSS.n1916 0.000965517
R10060 VSS.n1915 VSS.n1914 0.000965517
R10061 VSS.n1913 VSS.n1912 0.000965517
R10062 VSS.n3703 VSS.n3702 0.000963768
R10063 VSS.n3118 VSS.n3117 0.000962428
R10064 VSS.n2877 VSS.n2876 0.000951505
R10065 VSS.n2001 VSS.n1997 0.000951505
R10066 VSS.n2868 VSS.n2004 0.000951505
R10067 VSS.n2867 VSS.n2005 0.000951505
R10068 VSS.n2014 VSS.n2012 0.000951505
R10069 VSS.n2859 VSS.n2858 0.000951505
R10070 VSS.n2036 VSS.n2031 0.000951505
R10071 VSS.n2040 VSS.n2039 0.000951505
R10072 VSS.n2037 VSS.n2025 0.000951505
R10073 VSS.n2845 VSS.n2844 0.000951505
R10074 VSS.n2844 VSS.n2046 0.000951505
R10075 VSS.n2841 VSS.n2840 0.000951505
R10076 VSS.n2067 VSS.n2065 0.000951505
R10077 VSS.n2830 VSS.n2829 0.000951505
R10078 VSS.n2826 VSS.n2066 0.000951505
R10079 VSS.n2825 VSS.n2070 0.000951505
R10080 VSS.n2817 VSS.n2081 0.000951505
R10081 VSS.n2814 VSS.n2813 0.000951505
R10082 VSS.n2088 VSS.n2083 0.000951505
R10083 VSS.n2805 VSS.n2804 0.000951505
R10084 VSS.n2875 VSS.n2874 0.000951505
R10085 VSS.n2000 VSS.n1998 0.000951505
R10086 VSS.n2869 VSS.n2003 0.000951505
R10087 VSS.n2866 VSS.n2006 0.000951505
R10088 VSS.n2862 VSS.n2008 0.000951505
R10089 VSS.n2861 VSS.n2860 0.000951505
R10090 VSS.n2035 VSS.n2034 0.000951505
R10091 VSS.n2041 VSS.n2030 0.000951505
R10092 VSS.n2042 VSS.n2027 0.000951505
R10093 VSS.n2847 VSS.n2846 0.000951505
R10094 VSS.n2049 VSS.n2045 0.000951505
R10095 VSS.n2839 VSS.n2838 0.000951505
R10096 VSS.n2833 VSS.n2063 0.000951505
R10097 VSS.n2832 VSS.n2831 0.000951505
R10098 VSS.n2071 VSS.n2064 0.000951505
R10099 VSS.n2824 VSS.n2072 0.000951505
R10100 VSS.n2084 VSS.n2078 0.000951505
R10101 VSS.n2812 VSS.n2811 0.000951505
R10102 VSS.n2808 VSS.n2085 0.000951505
R10103 VSS.n2807 VSS.n2806 0.000951505
R10104 VSS.n2787 VSS.n2786 0.000951505
R10105 VSS.n2101 VSS.n2096 0.000951505
R10106 VSS.n2778 VSS.n2103 0.000951505
R10107 VSS.n2775 VSS.n2105 0.000951505
R10108 VSS.n2133 VSS.n2109 0.000951505
R10109 VSS.n2135 VSS.n2134 0.000951505
R10110 VSS.n2766 VSS.n2117 0.000951505
R10111 VSS.n2765 VSS.n2118 0.000951505
R10112 VSS.n2125 VSS.n2124 0.000951505
R10113 VSS.n2755 VSS.n2128 0.000951505
R10114 VSS.n2752 VSS.n2144 0.000951505
R10115 VSS.n2746 VSS.n2164 0.000951505
R10116 VSS.n2745 VSS.n2165 0.000951505
R10117 VSS.n2735 VSS.n2174 0.000951505
R10118 VSS.n2730 VSS.n2194 0.000951505
R10119 VSS.n2785 VSS.n2784 0.000951505
R10120 VSS.n2099 VSS.n2097 0.000951505
R10121 VSS.n2777 VSS.n2100 0.000951505
R10122 VSS.n2776 VSS.n2104 0.000951505
R10123 VSS.n2113 VSS.n2110 0.000951505
R10124 VSS.n2769 VSS.n2114 0.000951505
R10125 VSS.n2767 VSS.n2116 0.000951505
R10126 VSS.n2764 VSS.n2119 0.000951505
R10127 VSS.n2763 VSS.n2120 0.000951505
R10128 VSS.n2760 VSS.n2120 0.000951505
R10129 VSS.n2759 VSS.n2758 0.000951505
R10130 VSS.n2146 VSS.n2145 0.000951505
R10131 VSS.n2751 VSS.n2147 0.000951505
R10132 VSS.n2748 VSS.n2147 0.000951505
R10133 VSS.n2747 VSS.n2163 0.000951505
R10134 VSS.n2744 VSS.n2166 0.000951505
R10135 VSS.n2736 VSS.n2173 0.000951505
R10136 VSS.n2207 VSS.n2196 0.000951505
R10137 VSS.n2720 VSS.n2719 0.000951505
R10138 VSS.n2218 VSS.n2214 0.000951505
R10139 VSS.n2711 VSS.n2221 0.000951505
R10140 VSS.n2710 VSS.n2222 0.000951505
R10141 VSS.n2229 VSS.n2228 0.000951505
R10142 VSS.n2702 VSS.n2236 0.000951505
R10143 VSS.n2699 VSS.n2698 0.000951505
R10144 VSS.n2246 VSS.n2238 0.000951505
R10145 VSS.n2690 VSS.n2248 0.000951505
R10146 VSS.n2299 VSS.n2298 0.000951505
R10147 VSS.n2678 VSS.n2269 0.000951505
R10148 VSS.n2677 VSS.n2270 0.000951505
R10149 VSS.n2304 VSS.n2303 0.000951505
R10150 VSS.n2669 VSS.n2278 0.000951505
R10151 VSS.n2666 VSS.n2280 0.000951505
R10152 VSS.n2665 VSS.n2281 0.000951505
R10153 VSS.n2718 VSS.n2717 0.000951505
R10154 VSS.n2217 VSS.n2215 0.000951505
R10155 VSS.n2712 VSS.n2220 0.000951505
R10156 VSS.n2709 VSS.n2223 0.000951505
R10157 VSS.n2708 VSS.n2224 0.000951505
R10158 VSS.n2240 VSS.n2239 0.000951505
R10159 VSS.n2697 VSS.n2696 0.000951505
R10160 VSS.n2244 VSS.n2241 0.000951505
R10161 VSS.n2689 VSS.n2245 0.000951505
R10162 VSS.n2688 VSS.n2249 0.000951505
R10163 VSS.n2685 VSS.n2251 0.000951505
R10164 VSS.n2680 VSS.n2254 0.000951505
R10165 VSS.n2679 VSS.n2268 0.000951505
R10166 VSS.n2676 VSS.n2271 0.000951505
R10167 VSS.n2675 VSS.n2272 0.000951505
R10168 VSS.n2668 VSS.n2276 0.000951505
R10169 VSS.n2667 VSS.n2279 0.000951505
R10170 VSS.n2314 VSS.n2313 0.000951505
R10171 VSS.n2160 VSS.n2159 0.000950886
R10172 VSS.n1563 VSS.n1562 0.000920561
R10173 VSS.n3787 VSS.n3786 0.000920561
R10174 VSS.n3796 VSS.n3795 0.000920561
R10175 VSS.n3831 VSS.n3830 0.000920561
R10176 VSS.n3764 VSS.n3763 0.000920561
R10177 VSS.n3783 VSS.n3782 0.000920561
R10178 VSS.n3785 VSS.n3784 0.000920561
R10179 VSS.n3801 VSS.n3800 0.000920561
R10180 VSS.n3800 VSS.n3799 0.000920561
R10181 VSS.n3799 VSS.n3798 0.000920561
R10182 VSS.n3835 VSS.n3834 0.000920561
R10183 VSS.n3742 VSS.n3741 0.000920561
R10184 VSS.n3776 VSS.n3775 0.000920561
R10185 VSS.n3777 VSS.n3776 0.000920561
R10186 VSS.n3778 VSS.n3777 0.000920561
R10187 VSS.n3794 VSS.n3793 0.000920561
R10188 VSS.n3792 VSS.n3791 0.000920561
R10189 VSS.n1588 VSS.n1587 0.000914747
R10190 VSS.n1598 VSS.n1597 0.000914747
R10191 VSS.n1034 VSS.n1033 0.000914747
R10192 VSS.n3156 VSS.n3155 0.000904624
R10193 VSS.n2446 VSS.n2434 0.0009
R10194 VSS.n2558 VSS.n2415 0.000893013
R10195 VSS.n2557 VSS.n2556 0.000893013
R10196 VSS.n2427 VSS.n2424 0.000893013
R10197 VSS.n2547 VSS.n2546 0.000893013
R10198 VSS.n2542 VSS.n2541 0.000893013
R10199 VSS.n2437 VSS.n2431 0.000893013
R10200 VSS.n2533 VSS.n2532 0.000893013
R10201 VSS.n2528 VSS.n2441 0.000893013
R10202 VSS.n2449 VSS.n2442 0.000893013
R10203 VSS.n2520 VSS.n2452 0.000893013
R10204 VSS.n2517 VSS.n2516 0.000893013
R10205 VSS.n2472 VSS.n2454 0.000893013
R10206 VSS.n2507 VSS.n2506 0.000893013
R10207 VSS.n2503 VSS.n2473 0.000893013
R10208 VSS.n2495 VSS.n2481 0.000893013
R10209 VSS.n2494 VSS.n2482 0.000893013
R10210 VSS.n2419 VSS.n2417 0.000893013
R10211 VSS.n2555 VSS.n2554 0.000893013
R10212 VSS.n2554 VSS.n2418 0.000893013
R10213 VSS.n2550 VSS.n2422 0.000893013
R10214 VSS.n2549 VSS.n2548 0.000893013
R10215 VSS.n2540 VSS.n2539 0.000893013
R10216 VSS.n2435 VSS.n2432 0.000893013
R10217 VSS.n2535 VSS.n2534 0.000893013
R10218 VSS.n2445 VSS.n2443 0.000893013
R10219 VSS.n2523 VSS.n2444 0.000893013
R10220 VSS.n2455 VSS.n2448 0.000893013
R10221 VSS.n2515 VSS.n2514 0.000893013
R10222 VSS.n2470 VSS.n2456 0.000893013
R10223 VSS.n2509 VSS.n2508 0.000893013
R10224 VSS.n2476 VSS.n2471 0.000893013
R10225 VSS.n2496 VSS.n2480 0.000893013
R10226 VSS.n3732 VSS.n3731 0.000892442
R10227 VSS.n1740 VSS.n1739 0.000892442
R10228 VSS.n1738 VSS.n1737 0.000892442
R10229 VSS.n1736 VSS.n1735 0.000892442
R10230 VSS.n3716 VSS.n3715 0.000892442
R10231 VSS.n3715 VSS.n3714 0.000892442
R10232 VSS.n3707 VSS.n3706 0.000892442
R10233 VSS.n3694 VSS.n3693 0.000892442
R10234 VSS.n3692 VSS.n3691 0.000892442
R10235 VSS.n3690 VSS.n3689 0.000892442
R10236 VSS.n3678 VSS.n3677 0.000892442
R10237 VSS.n3656 VSS.n3655 0.000892442
R10238 VSS.n3654 VSS.n3653 0.000892442
R10239 VSS.n3643 VSS.n3642 0.000892442
R10240 VSS.n3645 VSS.n3644 0.000892442
R10241 VSS.n3630 VSS.n3629 0.000892442
R10242 VSS.n3628 VSS.n3627 0.000892442
R10243 VSS.n3578 VSS.n3577 0.000892442
R10244 VSS.n3729 VSS.n3728 0.000892442
R10245 VSS.n1734 VSS.n1733 0.000892442
R10246 VSS.n1732 VSS.n1731 0.000892442
R10247 VSS.n1730 VSS.n1729 0.000892442
R10248 VSS.n3720 VSS.n3719 0.000892442
R10249 VSS.n3719 VSS.n3718 0.000892442
R10250 VSS.n3705 VSS.n3704 0.000892442
R10251 VSS.n3700 VSS.n3699 0.000892442
R10252 VSS.n3698 VSS.n3697 0.000892442
R10253 VSS.n3676 VSS.n3675 0.000892442
R10254 VSS.n3661 VSS.n3660 0.000892442
R10255 VSS.n3659 VSS.n3658 0.000892442
R10256 VSS.n3639 VSS.n3638 0.000892442
R10257 VSS.n3641 VSS.n3640 0.000892442
R10258 VSS.n3635 VSS.n3634 0.000892442
R10259 VSS.n3633 VSS.n3632 0.000892442
R10260 VSS.n3576 VSS.n3575 0.000892442
R10261 VSS.n3518 VSS.n3517 0.000892442
R10262 VSS.n3450 VSS.n3449 0.000892442
R10263 VSS.n3451 VSS.n3450 0.000892442
R10264 VSS.n3453 VSS.n3452 0.000892442
R10265 VSS.n3456 VSS.n3455 0.000892442
R10266 VSS.n3458 VSS.n3457 0.000892442
R10267 VSS.n3493 VSS.n3492 0.000892442
R10268 VSS.n3491 VSS.n3490 0.000892442
R10269 VSS.n3488 VSS.n3487 0.000892442
R10270 VSS.n3486 VSS.n3485 0.000892442
R10271 VSS.n3484 VSS.n3483 0.000892442
R10272 VSS.n3480 VSS.n3479 0.000892442
R10273 VSS.n3478 VSS.n3477 0.000892442
R10274 VSS.n3476 VSS.n3475 0.000892442
R10275 VSS.n3474 VSS.n3473 0.000892442
R10276 VSS.n3472 VSS.n3471 0.000892442
R10277 VSS.n3469 VSS.n3468 0.000892442
R10278 VSS.n3467 VSS.n3466 0.000892442
R10279 VSS.n3465 VSS.n3464 0.000892442
R10280 VSS.n3461 VSS.n3460 0.000892442
R10281 VSS.n3440 VSS.n3439 0.000892442
R10282 VSS.n3445 VSS.n3444 0.000892442
R10283 VSS.n3447 VSS.n3446 0.000892442
R10284 VSS.n3566 VSS.n3565 0.000892442
R10285 VSS.n3565 VSS.n3564 0.000892442
R10286 VSS.n3563 VSS.n3562 0.000892442
R10287 VSS.n3560 VSS.n3559 0.000892442
R10288 VSS.n3558 VSS.n3557 0.000892442
R10289 VSS.n3556 VSS.n3555 0.000892442
R10290 VSS.n3550 VSS.n3549 0.000892442
R10291 VSS.n3548 VSS.n3547 0.000892442
R10292 VSS.n3546 VSS.n3545 0.000892442
R10293 VSS.n3544 VSS.n3543 0.000892442
R10294 VSS.n3541 VSS.n3540 0.000892442
R10295 VSS.n3539 VSS.n3538 0.000892442
R10296 VSS.n3537 VSS.n3536 0.000892442
R10297 VSS.n3533 VSS.n3532 0.000892442
R10298 VSS.n3411 VSS.n3410 0.000892442
R10299 VSS.n3409 VSS.n3408 0.000892442
R10300 VSS.n1768 VSS.n1767 0.000892442
R10301 VSS.n3347 VSS.n3346 0.000892442
R10302 VSS.n3349 VSS.n3348 0.000892442
R10303 VSS.n3351 VSS.n3350 0.000892442
R10304 VSS.n3327 VSS.n3326 0.000892442
R10305 VSS.n3325 VSS.n3324 0.000892442
R10306 VSS.n3323 VSS.n3322 0.000892442
R10307 VSS.n3306 VSS.n3305 0.000892442
R10308 VSS.n3308 VSS.n3307 0.000892442
R10309 VSS.n3310 VSS.n3309 0.000892442
R10310 VSS.n3282 VSS.n3281 0.000892442
R10311 VSS.n3287 VSS.n3286 0.000892442
R10312 VSS.n3285 VSS.n3284 0.000892442
R10313 VSS.n3272 VSS.n3271 0.000892442
R10314 VSS.n3270 VSS.n3269 0.000892442
R10315 VSS.n1766 VSS.n1765 0.000892442
R10316 VSS.n3341 VSS.n3340 0.000892442
R10317 VSS.n3343 VSS.n3342 0.000892442
R10318 VSS.n3345 VSS.n3344 0.000892442
R10319 VSS.n3334 VSS.n3333 0.000892442
R10320 VSS.n3332 VSS.n3331 0.000892442
R10321 VSS.n3330 VSS.n3329 0.000892442
R10322 VSS.n3302 VSS.n3301 0.000892442
R10323 VSS.n3304 VSS.n3303 0.000892442
R10324 VSS.n3313 VSS.n3312 0.000892442
R10325 VSS.n3280 VSS.n3279 0.000892442
R10326 VSS.n3293 VSS.n3292 0.000892442
R10327 VSS.n3291 VSS.n3290 0.000892442
R10328 VSS.n3267 VSS.n3266 0.000892442
R10329 VSS.n3265 VSS.n3264 0.000892442
R10330 VSS.n3254 VSS.n3253 0.000892442
R10331 VSS.n3246 VSS.n3245 0.000892442
R10332 VSS.n3237 VSS.n3236 0.000892442
R10333 VSS.n3235 VSS.n3234 0.000892442
R10334 VSS.n3195 VSS.n3194 0.000892442
R10335 VSS.n1787 VSS.n1786 0.000892442
R10336 VSS.n1789 VSS.n1788 0.000892442
R10337 VSS.n3180 VSS.n3179 0.000892442
R10338 VSS.n3178 VSS.n3177 0.000892442
R10339 VSS.n3176 VSS.n3175 0.000892442
R10340 VSS.n3164 VSS.n3163 0.000892442
R10341 VSS.n3162 VSS.n3161 0.000892442
R10342 VSS.n3143 VSS.n3142 0.000892442
R10343 VSS.n3128 VSS.n3127 0.000892442
R10344 VSS.n3126 VSS.n3125 0.000892442
R10345 VSS.n3109 VSS.n3108 0.000892442
R10346 VSS.n3107 VSS.n3106 0.000892442
R10347 VSS.n3096 VSS.n3095 0.000892442
R10348 VSS.n3094 VSS.n3093 0.000892442
R10349 VSS.n3205 VSS.n3204 0.000892442
R10350 VSS.n3203 VSS.n3202 0.000892442
R10351 VSS.n3193 VSS.n3192 0.000892442
R10352 VSS.n1783 VSS.n1782 0.000892442
R10353 VSS.n1785 VSS.n1784 0.000892442
R10354 VSS.n3185 VSS.n3184 0.000892442
R10355 VSS.n3183 VSS.n3182 0.000892442
R10356 VSS.n3160 VSS.n3159 0.000892442
R10357 VSS.n3169 VSS.n3168 0.000892442
R10358 VSS.n3167 VSS.n3166 0.000892442
R10359 VSS.n3149 VSS.n3148 0.000892442
R10360 VSS.n3139 VSS.n3138 0.000892442
R10361 VSS.n3137 VSS.n3136 0.000892442
R10362 VSS.n3123 VSS.n3122 0.000892442
R10363 VSS.n3121 VSS.n3120 0.000892442
R10364 VSS.n3101 VSS.n3100 0.000892442
R10365 VSS.n3099 VSS.n3098 0.000892442
R10366 VSS.n3058 VSS.n3057 0.000892442
R10367 VSS.n3062 VSS.n3061 0.000892442
R10368 VSS.n3060 VSS.n3059 0.000892442
R10369 VSS.n1823 VSS.n1822 0.000892442
R10370 VSS.n1821 VSS.n1820 0.000892442
R10371 VSS.n3043 VSS.n3042 0.000892442
R10372 VSS.n3033 VSS.n3032 0.000892442
R10373 VSS.n3035 VSS.n3034 0.000892442
R10374 VSS.n3021 VSS.n3020 0.000892442
R10375 VSS.n3020 VSS.n3019 0.000892442
R10376 VSS.n3008 VSS.n3007 0.000892442
R10377 VSS.n3010 VSS.n3009 0.000892442
R10378 VSS.n2992 VSS.n2991 0.000892442
R10379 VSS.n2994 VSS.n2993 0.000892442
R10380 VSS.n2996 VSS.n2995 0.000892442
R10381 VSS.n2972 VSS.n2971 0.000892442
R10382 VSS.n2970 VSS.n2969 0.000892442
R10383 VSS.n2968 VSS.n2967 0.000892442
R10384 VSS.n2920 VSS.n2919 0.000892442
R10385 VSS.n3056 VSS.n3055 0.000892442
R10386 VSS.n3067 VSS.n3066 0.000892442
R10387 VSS.n3065 VSS.n3064 0.000892442
R10388 VSS.n1819 VSS.n1818 0.000892442
R10389 VSS.n1817 VSS.n1816 0.000892442
R10390 VSS.n3047 VSS.n3046 0.000892442
R10391 VSS.n3031 VSS.n3030 0.000892442
R10392 VSS.n3026 VSS.n3025 0.000892442
R10393 VSS.n3024 VSS.n3023 0.000892442
R10394 VSS.n3006 VSS.n3005 0.000892442
R10395 VSS.n3013 VSS.n3012 0.000892442
R10396 VSS.n2986 VSS.n2985 0.000892442
R10397 VSS.n2988 VSS.n2987 0.000892442
R10398 VSS.n2990 VSS.n2989 0.000892442
R10399 VSS.n2979 VSS.n2978 0.000892442
R10400 VSS.n2977 VSS.n2976 0.000892442
R10401 VSS.n2975 VSS.n2974 0.000892442
R10402 VSS.n2918 VSS.n2917 0.000892442
R10403 VSS.n2654 VSS.n2653 0.000892442
R10404 VSS.n2328 VSS.n2322 0.000892442
R10405 VSS.n2343 VSS.n2335 0.000892442
R10406 VSS.n2344 VSS.n2342 0.000892442
R10407 VSS.n2631 VSS.n2347 0.000892442
R10408 VSS.n2628 VSS.n2349 0.000892442
R10409 VSS.n2627 VSS.n2350 0.000892442
R10410 VSS.n2622 VSS.n2362 0.000892442
R10411 VSS.n2619 VSS.n2362 0.000892442
R10412 VSS.n2618 VSS.n2617 0.000892442
R10413 VSS.n2388 VSS.n2386 0.000892442
R10414 VSS.n2607 VSS.n2606 0.000892442
R10415 VSS.n2603 VSS.n2387 0.000892442
R10416 VSS.n2602 VSS.n2391 0.000892442
R10417 VSS.n2594 VSS.n2401 0.000892442
R10418 VSS.n2593 VSS.n2402 0.000892442
R10419 VSS.n2590 VSS.n2589 0.000892442
R10420 VSS.n2566 VSS.n2405 0.000892442
R10421 VSS.n2652 VSS.n2651 0.000892442
R10422 VSS.n2324 VSS.n2323 0.000892442
R10423 VSS.n2646 VSS.n2645 0.000892442
R10424 VSS.n2336 VSS.n2327 0.000892442
R10425 VSS.n2339 VSS.n2337 0.000892442
R10426 VSS.n2634 VSS.n2340 0.000892442
R10427 VSS.n2354 VSS.n2341 0.000892442
R10428 VSS.n2356 VSS.n2355 0.000892442
R10429 VSS.n2626 VSS.n2351 0.000892442
R10430 VSS.n2369 VSS.n2368 0.000892442
R10431 VSS.n2368 VSS.n2365 0.000892442
R10432 VSS.n2616 VSS.n2615 0.000892442
R10433 VSS.n2610 VSS.n2384 0.000892442
R10434 VSS.n2609 VSS.n2608 0.000892442
R10435 VSS.n2392 VSS.n2385 0.000892442
R10436 VSS.n2601 VSS.n2393 0.000892442
R10437 VSS.n2595 VSS.n2400 0.000892442
R10438 VSS.n2407 VSS.n2406 0.000892442
R10439 VSS.n2588 VSS.n2587 0.000892442
R10440 VSS.n2565 VSS.n2408 0.000892442
R10441 VSS.n2762 VSS.n2761 0.000886473
R10442 VSS.n2750 VSS.n2749 0.000886473
R10443 VSS.n2371 VSS.n2370 0.000848837
R10444 VSS.n3713 VSS.n3712 0.000847826
R10445 VSS.n2524 VSS.n2447 0.000842857
R10446 VSS.n2836 VSS.n2835 0.000834448
R10447 VSS.n2159 VSS.n2123 0.000822061
R10448 VSS.n2311 VSS.n2274 0.000814465
R10449 VSS.n2192 VSS.n2177 0.000801003
R10450 VSS.n2185 VSS.n2178 0.000801003
R10451 VSS.n2191 VSS.n2190 0.000801003
R10452 VSS.n2733 VSS.n2732 0.000801003
R10453 VSS.n2757 VSS.n2756 0.000801003
R10454 VSS.n2183 VSS.n2180 0.000801003
R10455 VSS.n2187 VSS.n2186 0.000801003
R10456 VSS.n2172 VSS.n2171 0.000801003
R10457 VSS.n2734 VSS.n2175 0.000801003
R10458 VSS.n2201 VSS.n2200 0.000801003
R10459 VSS.n2758 VSS.n2126 0.000801003
R10460 VSS.n2743 VSS.n2167 0.000801003
R10461 VSS.n2182 VSS.n2181 0.000801003
R10462 VSS.n2738 VSS.n2737 0.000801003
R10463 VSS.n2202 VSS.n2199 0.000801003
R10464 VSS.n2206 VSS.n2205 0.000801003
R10465 VSS.n2289 VSS.n2288 0.000801003
R10466 VSS.n2251 VSS.n2249 0.000801003
R10467 VSS.n2370 VSS.n2367 0.000790698
R10468 VSS.n3147 VSS.n3134 0.000789017
R10469 VSS.n3252 VSS.n3243 0.000789017
R10470 VSS.n3895 VSS.n3894 0.00077907
R10471 VSS.n2076 VSS.n2075 0.000767559
R10472 VSS.n2821 VSS.n2820 0.000767559
R10473 VSS.n2810 VSS.n2809 0.000767559
R10474 VSS.n3682 VSS.n3681 0.000761628
R10475 VSS.n3680 VSS.n3679 0.000761628
R10476 VSS.n3673 VSS.n3672 0.000761628
R10477 VSS.n3454 VSS.n3453 0.000761628
R10478 VSS.n3442 VSS.n3441 0.000761628
R10479 VSS.n3562 VSS.n3561 0.000761628
R10480 VSS.n3553 VSS.n3552 0.000761628
R10481 VSS.n3379 VSS.n3378 0.000761628
R10482 VSS.n3410 VSS.n3409 0.000761628
R10483 VSS.n3257 VSS.n3256 0.000761628
R10484 VSS.n3250 VSS.n3249 0.000761628
R10485 VSS.n3365 VSS.n3364 0.000761628
R10486 VSS.n3314 VSS.n3313 0.000761628
R10487 VSS.n3266 VSS.n3265 0.000761628
R10488 VSS.n3251 VSS.n3246 0.000761628
R10489 VSS.n3216 VSS.n3215 0.000761628
R10490 VSS.n3152 VSS.n3151 0.000761628
R10491 VSS.n3145 VSS.n3144 0.000761628
R10492 VSS.n3108 VSS.n3107 0.000761628
R10493 VSS.n3146 VSS.n3139 0.000761628
R10494 VSS.n3113 VSS.n3112 0.000761628
R10495 VSS.n2642 VSS.n2641 0.000761628
R10496 VSS.n2643 VSS.n2330 0.000761628
R10497 VSS.n5785 VSS 0.000753521
R10498 VSS VSS.n5791 0.000753521
R10499 VSS.n2316 VSS.n2315 0.000751572
R10500 VSS.n1657 VSS.n1656 0.000751397
R10501 VSS.n1672 VSS.n1671 0.000751397
R10502 VSS.n1696 VSS.n1695 0.000751397
R10503 VSS.n1698 VSS.n1697 0.000751397
R10504 VSS.n1708 VSS.n1707 0.000751397
R10505 VSS.n1710 VSS.n1709 0.000751397
R10506 VSS.n1717 VSS.n1716 0.000751397
R10507 VSS.n3898 VSS.n3897 0.000751397
R10508 VSS.n3905 VSS.n3902 0.000751397
R10509 VSS.n4118 VSS.n4117 0.00074
R10510 VSS.n5881 VSS 0.000733766
R10511 VSS.n5880 VSS 0.000733766
R10512 VSS.n2614 VSS.n2613 0.000732558
R10513 VSS.n2396 VSS.n2383 0.000732558
R10514 VSS.n2599 VSS.n2598 0.000732558
R10515 VSS.n2409 VSS.n2398 0.000732558
R10516 VSS.n3001 VSS.n3000 0.000732558
R10517 VSS.n2984 VSS.n2981 0.000732558
R10518 VSS.n2965 VSS.n2964 0.000732558
R10519 VSS.n3650 VSS.n3649 0.000731884
R10520 VSS.n3648 VSS.n3637 0.000731884
R10521 VSS.n3626 VSS.n3625 0.000731884
R10522 VSS.n3174 VSS.n3173 0.000731214
R10523 VSS.n3155 VSS.n3154 0.000731214
R10524 VSS.n3105 VSS.n3104 0.000731214
R10525 VSS.n3361 VSS.n3360 0.000731214
R10526 VSS.n3260 VSS.n3259 0.000731214
R10527 VSS.n2420 VSS.n2410 0.000728571
R10528 VSS.n2511 VSS.n2510 0.000728571
R10529 VSS.n2500 VSS.n2499 0.000728571
R10530 VSS.n5831 VSS.n5830 0.000713777
R10531 VSS.n5833 VSS.n5832 0.000713777
R10532 VSS.n5835 VSS.n5834 0.000713777
R10533 VSS.n5885 VSS.n5884 0.000713777
R10534 VSS.n3821 VSS.n3820 0.00071028
R10535 VSS.n3745 VSS.n3744 0.00071028
R10536 VSS.n3822 VSS.n3818 0.00071028
R10537 VSS.n3752 VSS.n3751 0.00071028
R10538 VSS.n3768 VSS.n3767 0.00071028
R10539 VSS.n3804 VSS.n3790 0.00071028
R10540 VSS.n3804 VSS.n3803 0.00071028
R10541 VSS.n3793 VSS.n3792 0.00071028
R10542 VSS.n3824 VSS.n3823 0.00071028
R10543 VSS.n3837 VSS.n3836 0.00071028
R10544 VSS.n1610 VSS.n1609 0.000707373
R10545 VSS.n1618 VSS.n1617 0.000707373
R10546 VSS.n1620 VSS.n1619 0.000707373
R10547 VSS.n1630 VSS.n1629 0.000707373
R10548 VSS.n1632 VSS.n1631 0.000707373
R10549 VSS.n1641 VSS.n1639 0.000707373
R10550 VSS.n2893 VSS.n2892 0.000702532
R10551 VSS.n2890 VSS.n2889 0.000702532
R10552 VSS.n2887 VSS.n2886 0.000702532
R10553 VSS.n3774 VSS.n3773 0.00068648
R10554 VSS.n3808 VSS.n3807 0.00068648
R10555 VSS.n3901 VSS.n3899 0.000686047
R10556 VSS.n3567 VSS.n3437 0.000674419
R10557 VSS.n3427 VSS.n3426 0.000674419
R10558 VSS.n2553 VSS.n2552 0.000671429
R10559 VSS.n2513 VSS.n2512 0.000671429
R10560 VSS.n1889 VSS.n1888 0.000655172
R10561 VSS.n1901 VSS.n1900 0.000655172
R10562 VSS.n1926 VSS.n1925 0.000655172
R10563 VSS.n1916 VSS.n1915 0.000655172
R10564 VSS.n2826 VSS.n2825 0.000650502
R10565 VSS.n2813 VSS.n2083 0.000650502
R10566 VSS.n2072 VSS.n2071 0.000650502
R10567 VSS.n2811 VSS.n2085 0.000650502
R10568 VSS.n2754 VSS.n2127 0.000650502
R10569 VSS.n2756 VSS.n2755 0.000650502
R10570 VSS.n2186 VSS.n2183 0.000650502
R10571 VSS.n2200 VSS.n2175 0.000650502
R10572 VSS.n2181 VSS.n2167 0.000650502
R10573 VSS.n2205 VSS.n2202 0.000650502
R10574 VSS.n2288 VSS.n2287 0.000650502
R10575 VSS.n2290 VSS.n2289 0.000650502
R10576 VSS.n2507 VSS.n2472 0.000631004
R10577 VSS.n2495 VSS.n2494 0.000631004
R10578 VSS.n2509 VSS.n2470 0.000631004
R10579 VSS.n2490 VSS.n2480 0.000631004
R10580 VSS.n3605 VSS.n3604 0.000630814
R10581 VSS.n3681 VSS.n3680 0.000630814
R10582 VSS.n3644 VSS.n3643 0.000630814
R10583 VSS.n3629 VSS.n3628 0.000630814
R10584 VSS.n3674 VSS.n3673 0.000630814
R10585 VSS.n3672 VSS.n3671 0.000630814
R10586 VSS.n3640 VSS.n3639 0.000630814
R10587 VSS.n3634 VSS.n3633 0.000630814
R10588 VSS.n3481 VSS.n3480 0.000630814
R10589 VSS.n3443 VSS.n3442 0.000630814
R10590 VSS.n3552 VSS.n3551 0.000630814
R10591 VSS.n3377 VSS.n3376 0.000630814
R10592 VSS.n3257 VSS.n3255 0.000630814
R10593 VSS.n3250 VSS.n3247 0.000630814
R10594 VSS.n3366 VSS.n3365 0.000630814
R10595 VSS.n3364 VSS.n3363 0.000630814
R10596 VSS.n3294 VSS.n3280 0.000630814
R10597 VSS.n3258 VSS.n3254 0.000630814
R10598 VSS.n3214 VSS.n3213 0.000630814
R10599 VSS.n3152 VSS.n3150 0.000630814
R10600 VSS.n3145 VSS.n3140 0.000630814
R10601 VSS.n3153 VSS.n3149 0.000630814
R10602 VSS.n3114 VSS.n3113 0.000630814
R10603 VSS.n3112 VSS.n3111 0.000630814
R10604 VSS.n2995 VSS.n2994 0.000630814
R10605 VSS.n2969 VSS.n2968 0.000630814
R10606 VSS.n2989 VSS.n2988 0.000630814
R10607 VSS.n2976 VSS.n2975 0.000630814
R10608 VSS.n2644 VSS.n2643 0.000630814
R10609 VSS.n2334 VSS.n2330 0.000630814
R10610 VSS.n2606 VSS.n2387 0.000630814
R10611 VSS.n2594 VSS.n2593 0.000630814
R10612 VSS.n2608 VSS.n2385 0.000630814
R10613 VSS.n2406 VSS.n2400 0.000630814
R10614 VSS.n2742 VSS.n2741 0.000628824
R10615 VSS.n2739 VSS.n2170 0.000628824
R10616 VSS.n2204 VSS.n2198 0.000628824
R10617 VSS.n2682 VSS.n2266 0.000625786
R10618 VSS.n3436 VSS.n3435 0.000616279
R10619 VSS.n3430 VSS.n3429 0.000616279
R10620 VSS.n3668 VSS.n3667 0.000615942
R10621 VSS.n3315 VSS.n3300 0.000615607
R10622 VSS.n3262 VSS.n3261 0.000615607
R10623 VSS.n3754 VSS.n3753 0.00059324
R10624 VSS.n3770 VSS.n3769 0.00059324
R10625 VSS.n3781 VSS.n3780 0.00059324
R10626 VSS.n3805 VSS.n3781 0.00059324
R10627 VSS.n3806 VSS.n3805 0.00059324
R10628 VSS.n3826 VSS.n3825 0.00059324
R10629 VSS.n3839 VSS.n3838 0.00059324
R10630 VSS.n3880 VSS.n3879 0.000593023
R10631 VSS.n3882 VSS.n3881 0.000593023
R10632 VSS.n3888 VSS.n3887 0.000593023
R10633 VSS.n3890 VSS.n3889 0.000593023
R10634 VSS.n3901 VSS.n3900 0.000593023
R10635 VSS.n3848 VSS.n3847 0.000592166
R10636 VSS.n3853 VSS.n3852 0.000592166
R10637 VSS.n3855 VSS.n3854 0.000592166
R10638 VSS.n3862 VSS.n3861 0.000592166
R10639 VSS.n3864 VSS.n3863 0.000592166
R10640 VSS.n3869 VSS.n3868 0.000592166
R10641 VSS.n3003 VSS.n3002 0.00055814
R10642 VSS.n3571 VSS.n3570 0.00055814
R10643 VSS.n3317 VSS.n3316 0.000557804
R10644 VSS.n3296 VSS.n3295 0.000557804
R10645 VSS.n2896 VSS.n2895 0.000550633
R10646 PFD_T2_0.INV_mag_1.IN.n25 PFD_T2_0.INV_mag_1.IN.t0 226.316
R10647 PFD_T2_0.INV_mag_1.IN.n6 PFD_T2_0.INV_mag_1.IN.t26 116.993
R10648 PFD_T2_0.INV_mag_1.IN.n30 PFD_T2_0.INV_mag_1.IN.t32 33.8279
R10649 PFD_T2_0.INV_mag_1.IN.n31 PFD_T2_0.INV_mag_1.IN.n30 30.2144
R10650 PFD_T2_0.INV_mag_1.IN.t28 PFD_T2_0.INV_mag_1.IN.n3 25.0458
R10651 PFD_T2_0.INV_mag_1.IN.n28 PFD_T2_0.INV_mag_1.IN.n27 16.5048
R10652 PFD_T2_0.INV_mag_1.IN.n29 PFD_T2_0.INV_mag_1.IN.n28 16.5048
R10653 PFD_T2_0.INV_mag_1.IN.n3 PFD_T2_0.INV_mag_1.IN.t23 15.3305
R10654 PFD_T2_0.INV_mag_1.IN.n4 PFD_T2_0.INV_mag_1.IN.t29 15.1914
R10655 PFD_T2_0.INV_mag_1.IN.n3 PFD_T2_0.INV_mag_1.IN.n31 12.8616
R10656 PFD_T2_0.INV_mag_1.IN.n4 PFD_T2_0.INV_mag_1.IN.t21 12.6987
R10657 PFD_T2_0.INV_mag_1.IN.n5 PFD_T2_0.INV_mag_1.IN.t28 12.1515
R10658 PFD_T2_0.INV_mag_1.IN.t19 PFD_T2_0.INV_mag_1.IN.n6 11.3159
R10659 PFD_T2_0.INV_mag_1.IN.n25 PFD_T2_0.INV_mag_1.IN.t2 10.9468
R10660 PFD_T2_0.INV_mag_1.IN.n6 PFD_T2_0.INV_mag_1.IN.t17 10.2935
R10661 PFD_T2_0.INV_mag_1.IN.n0 PFD_T2_0.INV_mag_1.IN.n4 10.261
R10662 PFD_T2_0.INV_mag_1.IN.n27 PFD_T2_0.INV_mag_1.IN.t33 9.4175
R10663 PFD_T2_0.INV_mag_1.IN.n28 PFD_T2_0.INV_mag_1.IN.t20 9.4175
R10664 PFD_T2_0.INV_mag_1.IN.t23 PFD_T2_0.INV_mag_1.IN.n29 9.4175
R10665 PFD_T2_0.INV_mag_1.IN.n27 PFD_T2_0.INV_mag_1.IN.t22 9.1985
R10666 PFD_T2_0.INV_mag_1.IN.n28 PFD_T2_0.INV_mag_1.IN.t27 9.1985
R10667 PFD_T2_0.INV_mag_1.IN.n29 PFD_T2_0.INV_mag_1.IN.t30 9.1985
R10668 PFD_T2_0.INV_mag_1.IN.n3 PFD_T2_0.INV_mag_1.IN.t24 8.05323
R10669 PFD_T2_0.INV_mag_1.IN.n15 PFD_T2_0.INV_mag_1.IN.n14 6.76657
R10670 PFD_T2_0.INV_mag_1.IN.n1 PFD_T2_0.INV_mag_1.IN.n26 6.46231
R10671 PFD_T2_0.INV_mag_1.IN.n15 PFD_T2_0.INV_mag_1.IN.n12 5.58741
R10672 PFD_T2_0.INV_mag_1.IN.n22 PFD_T2_0.INV_mag_1.IN.n10 5.17308
R10673 PFD_T2_0.INV_mag_1.IN.n1 PFD_T2_0.INV_mag_1.IN.n25 4.73858
R10674 PFD_T2_0.INV_mag_1.IN.n30 PFD_T2_0.INV_mag_1.IN.t25 3.6505
R10675 PFD_T2_0.INV_mag_1.IN.n31 PFD_T2_0.INV_mag_1.IN.t18 3.6505
R10676 PFD_T2_0.INV_mag_1.IN.n8 PFD_T2_0.INV_mag_1.IN.t13 3.6405
R10677 PFD_T2_0.INV_mag_1.IN.n8 PFD_T2_0.INV_mag_1.IN.n7 3.6405
R10678 PFD_T2_0.INV_mag_1.IN.n10 PFD_T2_0.INV_mag_1.IN.t14 3.6405
R10679 PFD_T2_0.INV_mag_1.IN.n10 PFD_T2_0.INV_mag_1.IN.n9 3.6405
R10680 PFD_T2_0.INV_mag_1.IN.n20 PFD_T2_0.INV_mag_1.IN.t4 3.6405
R10681 PFD_T2_0.INV_mag_1.IN.n20 PFD_T2_0.INV_mag_1.IN.n19 3.6405
R10682 PFD_T2_0.INV_mag_1.IN.n12 PFD_T2_0.INV_mag_1.IN.t16 3.6405
R10683 PFD_T2_0.INV_mag_1.IN.n12 PFD_T2_0.INV_mag_1.IN.n11 3.6405
R10684 PFD_T2_0.INV_mag_1.IN.n17 PFD_T2_0.INV_mag_1.IN.t5 3.6405
R10685 PFD_T2_0.INV_mag_1.IN.n17 PFD_T2_0.INV_mag_1.IN.n16 3.6405
R10686 PFD_T2_0.INV_mag_1.IN.n24 PFD_T2_0.INV_mag_1.IN.t3 3.6405
R10687 PFD_T2_0.INV_mag_1.IN.n24 PFD_T2_0.INV_mag_1.IN.n23 3.6405
R10688 PFD_T2_0.INV_mag_1.IN.n14 PFD_T2_0.INV_mag_1.IN.t12 3.2765
R10689 PFD_T2_0.INV_mag_1.IN.n14 PFD_T2_0.INV_mag_1.IN.n13 3.2765
R10690 PFD_T2_0.INV_mag_1.IN.n2 PFD_T2_0.INV_mag_1.IN.n22 3.17603
R10691 PFD_T2_0.INV_mag_1.IN.n22 PFD_T2_0.INV_mag_1.IN.n21 3.15378
R10692 PFD_T2_0.INV_mag_1.IN.n1 PFD_T2_0.INV_mag_1.IN.n24 2.94791
R10693 PFD_T2_0.INV_mag_1.IN.n18 PFD_T2_0.INV_mag_1.IN.n17 2.92863
R10694 PFD_T2_0.INV_mag_1.IN.n21 PFD_T2_0.INV_mag_1.IN.n20 2.6005
R10695 PFD_T2_0.INV_mag_1.IN.n2 PFD_T2_0.INV_mag_1.IN.n8 2.6005
R10696 PFD_T2_0.INV_mag_1.IN.n18 PFD_T2_0.INV_mag_1.IN.n15 2.26925
R10697 PFD_T2_0.INV_mag_1.IN PFD_T2_0.INV_mag_1.IN.n0 6.76224
R10698 PFD_T2_0.INV_mag_1.IN PFD_T2_0.INV_mag_1.IN.t19 4.69745
R10699 PFD_T2_0.INV_mag_1.IN.n0 PFD_T2_0.INV_mag_1.IN.n5 2.6584
R10700 PFD_T2_0.INV_mag_1.IN.n2 PFD_T2_0.INV_mag_1.IN.n1 1.0806
R10701 PFD_T2_0.INV_mag_1.IN.n5 PFD_T2_0.INV_mag_1.IN.n2 1.06506
R10702 PFD_T2_0.INV_mag_1.IN.n21 PFD_T2_0.INV_mag_1.IN.n18 1.00114
R10703 PFD_T2_0.INV_mag_1.OUT.n0 PFD_T2_0.INV_mag_1.OUT.t9 29.3524
R10704 PFD_T2_0.INV_mag_1.OUT.n2 PFD_T2_0.INV_mag_1.OUT.t4 23.3605
R10705 PFD_T2_0.INV_mag_1.OUT.n3 PFD_T2_0.INV_mag_1.OUT.n0 16.8716
R10706 PFD_T2_0.INV_mag_1.OUT.n4 PFD_T2_0.INV_mag_1.OUT.t3 12.4111
R10707 PFD_T2_0.INV_mag_1.OUT.n0 PFD_T2_0.INV_mag_1.OUT.t6 9.0525
R10708 PFD_T2_0.INV_mag_1.OUT.n3 PFD_T2_0.INV_mag_1.OUT.t8 9.0525
R10709 PFD_T2_0.INV_mag_1.OUT.t3 PFD_T2_0.INV_mag_1.OUT.n3 9.0525
R10710 PFD_T2_0.INV_mag_1.OUT.n0 PFD_T2_0.INV_mag_1.OUT.t5 9.0525
R10711 PFD_T2_0.INV_mag_1.OUT.n2 PFD_T2_0.INV_mag_1.OUT.t7 8.7605
R10712 PFD_T2_0.INV_mag_1.OUT PFD_T2_0.INV_mag_1.OUT.n5 6.74425
R10713 PFD_T2_0.INV_mag_1.OUT PFD_T2_0.INV_mag_1.OUT.n1 5.41686
R10714 PFD_T2_0.INV_mag_1.OUT.n7 PFD_T2_0.INV_mag_1.OUT.t1 3.6405
R10715 PFD_T2_0.INV_mag_1.OUT.n7 PFD_T2_0.INV_mag_1.OUT.n6 3.6405
R10716 PFD_T2_0.INV_mag_1.OUT.n1 PFD_T2_0.INV_mag_1.OUT.n2 9.03264
R10717 PFD_T2_0.INV_mag_1.OUT PFD_T2_0.INV_mag_1.OUT.n7 3.34789
R10718 PFD_T2_0.INV_mag_1.OUT.n1 PFD_T2_0.INV_mag_1.OUT.n4 1.1347
R10719 PFD_T2_0.Buffer_V_2_0.IN.n1 PFD_T2_0.Buffer_V_2_0.IN.t11 13.2135
R10720 PFD_T2_0.Buffer_V_2_0.IN.n2 PFD_T2_0.Buffer_V_2_0.IN.n1 12.5844
R10721 PFD_T2_0.Buffer_V_2_0.IN.n1 PFD_T2_0.Buffer_V_2_0.IN.t13 9.8555
R10722 PFD_T2_0.Buffer_V_2_0.IN.n2 PFD_T2_0.Buffer_V_2_0.IN.t12 9.71737
R10723 PFD_T2_0.Buffer_V_2_0.IN.n16 PFD_T2_0.Buffer_V_2_0.IN.n7 6.60246
R10724 PFD_T2_0.Buffer_V_2_0.IN.n0 PFD_T2_0.Buffer_V_2_0.IN.n18 4.10693
R10725 PFD_T2_0.Buffer_V_2_0.IN.n0 PFD_T2_0.Buffer_V_2_0.IN.n2 3.78915
R10726 PFD_T2_0.Buffer_V_2_0.IN.n11 PFD_T2_0.Buffer_V_2_0.IN.t2 3.6405
R10727 PFD_T2_0.Buffer_V_2_0.IN.n11 PFD_T2_0.Buffer_V_2_0.IN.n10 3.6405
R10728 PFD_T2_0.Buffer_V_2_0.IN.n13 PFD_T2_0.Buffer_V_2_0.IN.t3 3.6405
R10729 PFD_T2_0.Buffer_V_2_0.IN.n13 PFD_T2_0.Buffer_V_2_0.IN.n12 3.6405
R10730 PFD_T2_0.Buffer_V_2_0.IN.n14 PFD_T2_0.Buffer_V_2_0.IN.n11 3.54941
R10731 PFD_T2_0.Buffer_V_2_0.IN.n15 PFD_T2_0.Buffer_V_2_0.IN.n9 3.33833
R10732 PFD_T2_0.Buffer_V_2_0.IN.n17 PFD_T2_0.Buffer_V_2_0.IN.n6 3.33833
R10733 PFD_T2_0.Buffer_V_2_0.IN.n9 PFD_T2_0.Buffer_V_2_0.IN.t5 3.2765
R10734 PFD_T2_0.Buffer_V_2_0.IN.n9 PFD_T2_0.Buffer_V_2_0.IN.n8 3.2765
R10735 PFD_T2_0.Buffer_V_2_0.IN.n4 PFD_T2_0.Buffer_V_2_0.IN.t10 3.2765
R10736 PFD_T2_0.Buffer_V_2_0.IN.n4 PFD_T2_0.Buffer_V_2_0.IN.n3 3.2765
R10737 PFD_T2_0.Buffer_V_2_0.IN.n6 PFD_T2_0.Buffer_V_2_0.IN.t9 3.2765
R10738 PFD_T2_0.Buffer_V_2_0.IN.n6 PFD_T2_0.Buffer_V_2_0.IN.n5 3.2765
R10739 PFD_T2_0.Buffer_V_2_0.IN.n14 PFD_T2_0.Buffer_V_2_0.IN.n13 2.78441
R10740 PFD_T2_0.Buffer_V_2_0.IN.n18 PFD_T2_0.Buffer_V_2_0.IN.n4 1.8538
R10741 PFD_T2_0.Buffer_V_2_0.IN.n18 PFD_T2_0.Buffer_V_2_0.IN.n17 0.78641
R10742 PFD_T2_0.Buffer_V_2_0.IN.n16 PFD_T2_0.Buffer_V_2_0.IN.n15 0.524848
R10743 PFD_T2_0.Buffer_V_2_0.IN.n15 PFD_T2_0.Buffer_V_2_0.IN.n14 0.358543
R10744 PFD_T2_0.Buffer_V_2_0.IN.n17 PFD_T2_0.Buffer_V_2_0.IN.n16 0.274413
R10745 PFD_T2_0.Buffer_V_2_0.IN PFD_T2_0.Buffer_V_2_0.IN.n0 0.264033
R10746 PFD_T2_0.INV_mag_0.IN.n6 PFD_T2_0.INV_mag_0.IN.t14 219.017
R10747 PFD_T2_0.INV_mag_0.IN.n3 PFD_T2_0.INV_mag_0.IN.t28 116.993
R10748 PFD_T2_0.INV_mag_0.IN.n25 PFD_T2_0.INV_mag_0.IN.t23 33.8279
R10749 PFD_T2_0.INV_mag_0.IN.n26 PFD_T2_0.INV_mag_0.IN.n25 30.2144
R10750 PFD_T2_0.INV_mag_0.IN.t20 PFD_T2_0.INV_mag_0.IN.n1 25.0458
R10751 PFD_T2_0.INV_mag_0.IN.n28 PFD_T2_0.INV_mag_0.IN.n27 16.5048
R10752 PFD_T2_0.INV_mag_0.IN.n29 PFD_T2_0.INV_mag_0.IN.n28 16.5048
R10753 PFD_T2_0.INV_mag_0.IN.n1 PFD_T2_0.INV_mag_0.IN.t24 15.3305
R10754 PFD_T2_0.INV_mag_0.IN.n4 PFD_T2_0.INV_mag_0.IN.t25 15.2644
R10755 PFD_T2_0.INV_mag_0.IN.n1 PFD_T2_0.INV_mag_0.IN.n26 12.8616
R10756 PFD_T2_0.INV_mag_0.IN.n4 PFD_T2_0.INV_mag_0.IN.t17 12.7717
R10757 PFD_T2_0.INV_mag_0.IN.n0 PFD_T2_0.INV_mag_0.IN.t20 12.0785
R10758 PFD_T2_0.INV_mag_0.IN.t18 PFD_T2_0.INV_mag_0.IN.n3 11.3197
R10759 PFD_T2_0.INV_mag_0.IN.n6 PFD_T2_0.INV_mag_0.IN.t12 10.8543
R10760 PFD_T2_0.INV_mag_0.IN.n3 PFD_T2_0.INV_mag_0.IN.t29 10.2935
R10761 PFD_T2_0.INV_mag_0.IN.n27 PFD_T2_0.INV_mag_0.IN.t21 9.4175
R10762 PFD_T2_0.INV_mag_0.IN.n28 PFD_T2_0.INV_mag_0.IN.t31 9.4175
R10763 PFD_T2_0.INV_mag_0.IN.t24 PFD_T2_0.INV_mag_0.IN.n29 9.4175
R10764 PFD_T2_0.INV_mag_0.IN.n27 PFD_T2_0.INV_mag_0.IN.t33 9.1985
R10765 PFD_T2_0.INV_mag_0.IN.n28 PFD_T2_0.INV_mag_0.IN.t26 9.1985
R10766 PFD_T2_0.INV_mag_0.IN.n29 PFD_T2_0.INV_mag_0.IN.t19 9.1985
R10767 PFD_T2_0.INV_mag_0.IN.n30 PFD_T2_0.INV_mag_0.IN.n4 8.99637
R10768 PFD_T2_0.INV_mag_0.IN.n1 PFD_T2_0.INV_mag_0.IN.t32 8.05323
R10769 PFD_T2_0.INV_mag_0.IN.n17 PFD_T2_0.INV_mag_0.IN.n16 6.76657
R10770 PFD_T2_0.INV_mag_0.IN.n2 PFD_T2_0.INV_mag_0.IN.n5 6.46389
R10771 PFD_T2_0.INV_mag_0.IN.n22 PFD_T2_0.INV_mag_0.IN.n10 5.77603
R10772 PFD_T2_0.INV_mag_0.IN.n17 PFD_T2_0.INV_mag_0.IN.n14 5.58741
R10773 PFD_T2_0.INV_mag_0.IN PFD_T2_0.INV_mag_0.IN.n30 5.21028
R10774 PFD_T2_0.INV_mag_0.IN.n2 PFD_T2_0.INV_mag_0.IN.n6 4.7386
R10775 PFD_T2_0.INV_mag_0.IN PFD_T2_0.INV_mag_0.IN.t18 4.69432
R10776 PFD_T2_0.INV_mag_0.IN.n25 PFD_T2_0.INV_mag_0.IN.t30 3.6505
R10777 PFD_T2_0.INV_mag_0.IN.n26 PFD_T2_0.INV_mag_0.IN.t22 3.6505
R10778 PFD_T2_0.INV_mag_0.IN.n14 PFD_T2_0.INV_mag_0.IN.t1 3.6405
R10779 PFD_T2_0.INV_mag_0.IN.n14 PFD_T2_0.INV_mag_0.IN.n13 3.6405
R10780 PFD_T2_0.INV_mag_0.IN.n12 PFD_T2_0.INV_mag_0.IN.t3 3.6405
R10781 PFD_T2_0.INV_mag_0.IN.n12 PFD_T2_0.INV_mag_0.IN.n11 3.6405
R10782 PFD_T2_0.INV_mag_0.IN.n24 PFD_T2_0.INV_mag_0.IN.t2 3.6405
R10783 PFD_T2_0.INV_mag_0.IN.n24 PFD_T2_0.INV_mag_0.IN.n23 3.6405
R10784 PFD_T2_0.INV_mag_0.IN.n8 PFD_T2_0.INV_mag_0.IN.t13 3.6405
R10785 PFD_T2_0.INV_mag_0.IN.n8 PFD_T2_0.INV_mag_0.IN.n7 3.6405
R10786 PFD_T2_0.INV_mag_0.IN.n10 PFD_T2_0.INV_mag_0.IN.t4 3.6405
R10787 PFD_T2_0.INV_mag_0.IN.n10 PFD_T2_0.INV_mag_0.IN.n9 3.6405
R10788 PFD_T2_0.INV_mag_0.IN.n19 PFD_T2_0.INV_mag_0.IN.t0 3.6405
R10789 PFD_T2_0.INV_mag_0.IN.n19 PFD_T2_0.INV_mag_0.IN.n18 3.6405
R10790 PFD_T2_0.INV_mag_0.IN.n16 PFD_T2_0.INV_mag_0.IN.t16 3.2765
R10791 PFD_T2_0.INV_mag_0.IN.n16 PFD_T2_0.INV_mag_0.IN.n15 3.2765
R10792 PFD_T2_0.INV_mag_0.IN.n22 PFD_T2_0.INV_mag_0.IN.n21 3.15378
R10793 PFD_T2_0.INV_mag_0.IN.n2 PFD_T2_0.INV_mag_0.IN.n8 2.94651
R10794 PFD_T2_0.INV_mag_0.IN.n20 PFD_T2_0.INV_mag_0.IN.n19 2.92863
R10795 PFD_T2_0.INV_mag_0.IN.n0 PFD_T2_0.INV_mag_0.IN.n24 2.6005
R10796 PFD_T2_0.INV_mag_0.IN.n21 PFD_T2_0.INV_mag_0.IN.n12 2.6005
R10797 PFD_T2_0.INV_mag_0.IN.n0 PFD_T2_0.INV_mag_0.IN.n22 2.57308
R10798 PFD_T2_0.INV_mag_0.IN.n20 PFD_T2_0.INV_mag_0.IN.n17 2.26925
R10799 PFD_T2_0.INV_mag_0.IN.n21 PFD_T2_0.INV_mag_0.IN.n20 1.00114
R10800 PFD_T2_0.INV_mag_0.IN.n30 PFD_T2_0.INV_mag_0.IN.n0 3.21412
R10801 PFD_T2_0.INV_mag_0.IN.n0 PFD_T2_0.INV_mag_0.IN.n2 2.10654
R10802 a_24437_9224.n3 a_24437_9224.n2 7.21994
R10803 a_24437_9224.n2 a_24437_9224.t2 7.21316
R10804 a_24437_9224.n1 a_24437_9224.t0 3.6405
R10805 a_24437_9224.n1 a_24437_9224.n0 3.6405
R10806 a_24437_9224.n2 a_24437_9224.n1 2.76192
R10807 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n21 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t41 23.6945
R10808 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n22 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t51 23.6945
R10809 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n22 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n21 18.8035
R10810 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n19 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n16 15.8172
R10811 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n25 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n24 15.8172
R10812 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n24 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n16 15.8172
R10813 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t56 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n19 14.8925
R10814 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t42 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n16 14.8925
R10815 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n24 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t49 14.8925
R10816 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n23 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n17 12.2457
R10817 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n23 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n18 12.2457
R10818 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n20 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n18 12.2457
R10819 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n26 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t37 11.6285
R10820 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n9 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t34 9.07373
R10821 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n9 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t55 8.94903
R10822 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t50 8.91906
R10823 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t32 8.91906
R10824 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t54 8.91906
R10825 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t41 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n20 8.9065
R10826 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t57 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n18 8.9065
R10827 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n23 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t36 8.9065
R10828 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t51 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n17 8.9065
R10829 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t43 8.88175
R10830 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n9 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t48 8.78051
R10831 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t44 8.78051
R10832 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n9 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t38 8.76753
R10833 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n9 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t58 8.76753
R10834 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n13 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t24 8.71893
R10835 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t52 8.71324
R10836 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t46 8.71324
R10837 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n19 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t53 8.6145
R10838 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n16 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t40 8.6145
R10839 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n24 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t45 8.6145
R10840 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n25 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t31 8.59715
R10841 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t35 8.50259
R10842 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t47 8.38837
R10843 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n20 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t56 8.3225
R10844 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n18 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t42 8.3225
R10845 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t49 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n23 8.3225
R10846 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n17 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t37 8.3225
R10847 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n9 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t33 8.30411
R10848 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t39 7.40199
R10849 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n8 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t2 6.43598
R10850 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n36 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n14 6.42121
R10851 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n8 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t29 6.39767
R10852 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t3 6.02861
R10853 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n33 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n32 5.82997
R10854 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n5 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n45 8.13848
R10855 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n36 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n35 5.23266
R10856 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n50 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t7 4.93756
R10857 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n40 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t14 4.89657
R10858 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n10 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n51 4.89332
R10859 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n13 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t25 4.76585
R10860 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n14 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n29 4.70534
R10861 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n14 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n28 4.70317
R10862 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n26 4.60939
R10863 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n55 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n6 4.53389
R10864 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n6 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n54 4.22351
R10865 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n43 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n42 4.04842
R10866 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n52 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t15 4.00791
R10867 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n57 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n56 3.96274
R10868 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n37 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n27 3.95313
R10869 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n13 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t19 3.94347
R10870 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n6 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t18 3.80888
R10871 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n33 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n31 3.77407
R10872 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n8 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n59 3.75742
R10873 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n27 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN 3.73676
R10874 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n59 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n58 3.65936
R10875 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n21 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t57 3.6505
R10876 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t36 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n22 3.6505
R10877 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n49 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t12 3.6405
R10878 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n49 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n48 3.6405
R10879 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n1 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t6 3.6405
R10880 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n1 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n46 3.6405
R10881 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n0 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t5 3.6405
R10882 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n0 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n39 3.6405
R10883 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n35 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n34 3.47613
R10884 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n31 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n30 3.47611
R10885 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n14 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n33 3.35867
R10886 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n12 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n36 3.3208
R10887 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n59 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t0 3.31708
R10888 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n12 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n13 3.31211
R10889 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n26 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n25 3.1807
R10890 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n8 3.15957
R10891 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n37 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n12 3.14573
R10892 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n15 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n50 2.97396
R10893 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n31 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t22 2.86261
R10894 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n35 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t27 2.8626
R10895 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n12 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN 2.7938
R10896 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n55 2.75901
R10897 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n2 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n15 2.62313
R10898 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n27 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN 2.36584
R10899 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n11 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n37 2.35267
R10900 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n44 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n43 2.24883
R10901 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n53 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n52 2.24559
R10902 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n11 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n2 2.03424
R10903 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n9 1.9805
R10904 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n10 1.86182
R10905 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n55 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n53 1.85837
R10906 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n8 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n7 1.81023
R10907 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n15 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n41 1.78522
R10908 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n5 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n49 4.56052
R10909 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n2 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n38 3.16799
R10910 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n3 2.93012
R10911 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n15 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n5 2.786
R10912 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n38 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n0 2.75194
R10913 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n47 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n1 2.75094
R10914 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n11 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n4 2.62258
R10915 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n5 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n47 1.77011
R10916 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n5 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n44 1.76105
R10917 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n57 1.5089
R10918 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n41 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n40 1.495
R10919 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n7 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n11 1.47485
R10920 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n2 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t12 15.4917
R10921 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n4 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t14 15.3942
R10922 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n5 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t16 14.904
R10923 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n9 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t15 14.7749
R10924 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n3 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t21 13.6019
R10925 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n9 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t18 13.5312
R10926 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n7 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t19 13.4877
R10927 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n5 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t20 13.227
R10928 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n6 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t13 13.1835
R10929 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n2 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t17 8.17943
R10930 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n0 4.7425
R10931 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n25 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t7 3.6405
R10932 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n25 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n24 3.6405
R10933 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n16 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t5 3.6405
R10934 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n16 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n15 3.6405
R10935 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n14 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t9 3.6405
R10936 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n14 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n13 3.6405
R10937 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n23 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t11 3.6405
R10938 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n23 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n22 3.6405
R10939 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n27 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n21 3.50463
R10940 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n28 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n19 3.50463
R10941 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n21 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t1 3.2765
R10942 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n21 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n20 3.2765
R10943 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n19 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t0 3.2765
R10944 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n19 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n18 3.2765
R10945 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n17 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n14 3.06224
R10946 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n26 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n23 3.06224
R10947 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n17 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n16 2.6005
R10948 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n26 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n25 2.6005
R10949 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n1 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT 2.28587
R10950 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n12 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n1 2.2505
R10951 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n8 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n4 1.5982
R10952 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n10 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n8 1.18336
R10953 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n11 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n10 0.961395
R10954 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n1 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n11 0.806561
R10955 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n28 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n27 0.798761
R10956 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n0 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT 0.65726
R10957 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n1 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n0 0.56461
R10958 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n28 0.539611
R10959 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n3 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n2 0.381495
R10960 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n10 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n9 0.37501
R10961 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n4 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n3 0.355126
R10962 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n7 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n6 0.31227
R10963 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n6 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n5 0.298874
R10964 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n8 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n7 0.233052
R10965 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n28 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n17 0.18637
R10966 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n27 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n26 0.18637
R10967 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n12 0.185454
R10968 VCTRL2.n124 VCTRL2.n123 10.0043
R10969 VCTRL2.n124 VCTRL2.n61 9.34779
R10970 VCTRL2.n53 VCTRL2.t66 8.213
R10971 VCTRL2.n26 VCTRL2.t30 8.213
R10972 VCTRL2.n112 VCTRL2.t12 8.16955
R10973 VCTRL2.n99 VCTRL2.t36 8.16955
R10974 VCTRL2.n33 VCTRL2.t23 8.16955
R10975 VCTRL2.n18 VCTRL2.t16 8.16955
R10976 VCTRL2.n22 VCTRL2.t24 8.16955
R10977 VCTRL2.n58 VCTRL2.t34 8.16955
R10978 VCTRL2.n88 VCTRL2.t22 8.1261
R10979 VCTRL2.n81 VCTRL2.t26 8.1261
R10980 VCTRL2.n95 VCTRL2.t17 8.1261
R10981 VCTRL2.n117 VCTRL2.t0 8.1261
R10982 VCTRL2.n44 VCTRL2.t11 8.1261
R10983 VCTRL2.n13 VCTRL2.t67 8.1261
R10984 VCTRL2.n75 VCTRL2.t9 8.08264
R10985 VCTRL2.n67 VCTRL2.t72 8.08264
R10986 VCTRL2.n49 VCTRL2.t15 7.51776
R10987 VCTRL2.n24 VCTRL2.t70 7.51776
R10988 VCTRL2.n108 VCTRL2.t13 7.47431
R10989 VCTRL2.n97 VCTRL2.t44 7.47431
R10990 VCTRL2.n56 VCTRL2.t74 7.47431
R10991 VCTRL2.n29 VCTRL2.t60 7.47431
R10992 VCTRL2.n15 VCTRL2.t54 7.47431
R10993 VCTRL2.n51 VCTRL2.t2 7.47431
R10994 VCTRL2.n20 VCTRL2.t61 7.47431
R10995 VCTRL2.n25 VCTRL2.t48 7.47431
R10996 VCTRL2.n85 VCTRL2.t49 7.43086
R10997 VCTRL2.n78 VCTRL2.t59 7.43086
R10998 VCTRL2.n111 VCTRL2.t1 7.43086
R10999 VCTRL2.n92 VCTRL2.t75 7.43086
R11000 VCTRL2.n115 VCTRL2.t19 7.43086
R11001 VCTRL2.n98 VCTRL2.t27 7.43086
R11002 VCTRL2.n30 VCTRL2.t38 7.43086
R11003 VCTRL2.n16 VCTRL2.t32 7.43086
R11004 VCTRL2.n41 VCTRL2.t45 7.43086
R11005 VCTRL2.n5 VCTRL2.t18 7.43086
R11006 VCTRL2.n21 VCTRL2.t39 7.43086
R11007 VCTRL2.n57 VCTRL2.t51 7.43086
R11008 VCTRL2.n87 VCTRL2.t33 7.3874
R11009 VCTRL2.n80 VCTRL2.t40 7.3874
R11010 VCTRL2.n72 VCTRL2.t8 7.3874
R11011 VCTRL2.n65 VCTRL2.t31 7.3874
R11012 VCTRL2.n93 VCTRL2.t57 7.3874
R11013 VCTRL2.n116 VCTRL2.t7 7.3874
R11014 VCTRL2.n42 VCTRL2.t25 7.3874
R11015 VCTRL2.n11 VCTRL2.t3 7.3874
R11016 VCTRL2.n74 VCTRL2.t73 7.34395
R11017 VCTRL2.n66 VCTRL2.t14 7.34395
R11018 VCTRL2.n76 VCTRL2.t62 7.3005
R11019 VCTRL2.n68 VCTRL2.t42 7.3005
R11020 VCTRL2.n96 VCTRL2.t76 7.25705
R11021 VCTRL2.n89 VCTRL2.t79 7.25705
R11022 VCTRL2.n82 VCTRL2.t4 7.25705
R11023 VCTRL2.t9 VCTRL2.n74 7.25705
R11024 VCTRL2.t72 VCTRL2.n66 7.25705
R11025 VCTRL2.n118 VCTRL2.t52 7.25705
R11026 VCTRL2.n45 VCTRL2.t28 7.25705
R11027 VCTRL2.n14 VCTRL2.t6 7.25705
R11028 VCTRL2.n100 VCTRL2.t10 7.2136
R11029 VCTRL2.t22 VCTRL2.n87 7.2136
R11030 VCTRL2.t26 VCTRL2.n80 7.2136
R11031 VCTRL2.t73 VCTRL2.n72 7.2136
R11032 VCTRL2.t14 VCTRL2.n65 7.2136
R11033 VCTRL2.n113 VCTRL2.t69 7.2136
R11034 VCTRL2.t17 VCTRL2.n93 7.2136
R11035 VCTRL2.t0 VCTRL2.n116 7.2136
R11036 VCTRL2.n34 VCTRL2.t41 7.2136
R11037 VCTRL2.n19 VCTRL2.t35 7.2136
R11038 VCTRL2.t11 VCTRL2.n42 7.2136
R11039 VCTRL2.t67 VCTRL2.n11 7.2136
R11040 VCTRL2.n23 VCTRL2.t43 7.2136
R11041 VCTRL2.n59 VCTRL2.t55 7.2136
R11042 VCTRL2.t33 VCTRL2.n85 7.17014
R11043 VCTRL2.t40 VCTRL2.n78 7.17014
R11044 VCTRL2.t12 VCTRL2.n111 7.17014
R11045 VCTRL2.t57 VCTRL2.n92 7.17014
R11046 VCTRL2.t7 VCTRL2.n115 7.17014
R11047 VCTRL2.t36 VCTRL2.n98 7.17014
R11048 VCTRL2.t23 VCTRL2.n30 7.17014
R11049 VCTRL2.t16 VCTRL2.n16 7.17014
R11050 VCTRL2.t25 VCTRL2.n41 7.17014
R11051 VCTRL2.t3 VCTRL2.n5 7.17014
R11052 VCTRL2.n54 VCTRL2.t5 7.17014
R11053 VCTRL2.t24 VCTRL2.n21 7.17014
R11054 VCTRL2.t34 VCTRL2.n57 7.17014
R11055 VCTRL2.n27 VCTRL2.t50 7.17014
R11056 VCTRL2.t1 VCTRL2.n108 7.12669
R11057 VCTRL2.t27 VCTRL2.n97 7.12669
R11058 VCTRL2.t38 VCTRL2.n29 7.12669
R11059 VCTRL2.t32 VCTRL2.n15 7.12669
R11060 VCTRL2.t66 VCTRL2.n51 7.12669
R11061 VCTRL2.t39 VCTRL2.n20 7.12669
R11062 VCTRL2.t51 VCTRL2.n56 7.12669
R11063 VCTRL2.t30 VCTRL2.n25 7.12669
R11064 VCTRL2.t2 VCTRL2.n49 7.08324
R11065 VCTRL2.n54 VCTRL2.t20 7.08324
R11066 VCTRL2.t48 VCTRL2.n24 7.08324
R11067 VCTRL2.n27 VCTRL2.t71 7.08324
R11068 VCTRL2.n113 VCTRL2.t53 7.03979
R11069 VCTRL2.n100 VCTRL2.t78 7.03979
R11070 VCTRL2.n34 VCTRL2.t63 7.03979
R11071 VCTRL2.n19 VCTRL2.t56 7.03979
R11072 VCTRL2.n23 VCTRL2.t64 7.03979
R11073 VCTRL2.n59 VCTRL2.t77 7.03979
R11074 VCTRL2.n96 VCTRL2.t58 6.99633
R11075 VCTRL2.n89 VCTRL2.t65 6.99633
R11076 VCTRL2.n82 VCTRL2.t68 6.99633
R11077 VCTRL2.n118 VCTRL2.t37 6.99633
R11078 VCTRL2.n45 VCTRL2.t47 6.99633
R11079 VCTRL2.n14 VCTRL2.t21 6.99633
R11080 VCTRL2.n76 VCTRL2.t46 6.95288
R11081 VCTRL2.n68 VCTRL2.t29 6.95288
R11082 VCTRL2.t46 VCTRL2.n75 6.51836
R11083 VCTRL2.t29 VCTRL2.n67 6.51836
R11084 VCTRL2.t58 VCTRL2.n95 6.4749
R11085 VCTRL2.t65 VCTRL2.n88 6.4749
R11086 VCTRL2.t68 VCTRL2.n81 6.4749
R11087 VCTRL2.t37 VCTRL2.n117 6.4749
R11088 VCTRL2.t47 VCTRL2.n44 6.4749
R11089 VCTRL2.t21 VCTRL2.n13 6.4749
R11090 VCTRL2.t53 VCTRL2.n112 6.43145
R11091 VCTRL2.t78 VCTRL2.n99 6.43145
R11092 VCTRL2.t63 VCTRL2.n33 6.43145
R11093 VCTRL2.t56 VCTRL2.n18 6.43145
R11094 VCTRL2.t64 VCTRL2.n22 6.43145
R11095 VCTRL2.t77 VCTRL2.n58 6.43145
R11096 VCTRL2.t20 VCTRL2.n53 6.388
R11097 VCTRL2.t71 VCTRL2.n26 6.388
R11098 VCTRL2.n28 VCTRL2.n27 4.03166
R11099 VCTRL2.n101 VCTRL2.n100 4.0306
R11100 VCTRL2.n119 VCTRL2.n118 3.63007
R11101 VCTRL2.n60 VCTRL2.n59 3.62933
R11102 VCTRL2.n11 VCTRL2.n10 3.62499
R11103 VCTRL2.n102 VCTRL2.n89 3.62466
R11104 VCTRL2.n88 VCTRL2.n83 3.62466
R11105 VCTRL2.n108 VCTRL2.n107 3.62466
R11106 VCTRL2.n5 VCTRL2.n4 3.62466
R11107 VCTRL2.n41 VCTRL2.n40 3.62466
R11108 VCTRL2.n28 VCTRL2.n23 3.62466
R11109 VCTRL2.n36 VCTRL2.n19 3.62466
R11110 VCTRL2.n47 VCTRL2.n14 3.62466
R11111 VCTRL2.n85 VCTRL2.n84 3.62466
R11112 VCTRL2.n87 VCTRL2.n86 3.62466
R11113 VCTRL2.n112 VCTRL2.n106 3.62466
R11114 VCTRL2.n114 VCTRL2.n113 3.62466
R11115 VCTRL2.n111 VCTRL2.n110 3.62466
R11116 VCTRL2.n18 VCTRL2.n17 3.62466
R11117 VCTRL2.n44 VCTRL2.n43 3.62466
R11118 VCTRL2.n46 VCTRL2.n45 3.62466
R11119 VCTRL2.n13 VCTRL2.n12 3.62466
R11120 VCTRL2.n101 VCTRL2.n96 3.62462
R11121 VCTRL2.n103 VCTRL2.n82 3.62462
R11122 VCTRL2.n78 VCTRL2.n77 3.62462
R11123 VCTRL2.n80 VCTRL2.n79 3.62462
R11124 VCTRL2.n75 VCTRL2.n70 3.62462
R11125 VCTRL2.n104 VCTRL2.n76 3.62462
R11126 VCTRL2.n72 VCTRL2.n71 3.62462
R11127 VCTRL2.n74 VCTRL2.n73 3.62462
R11128 VCTRL2.n67 VCTRL2.n63 3.62462
R11129 VCTRL2.n105 VCTRL2.n68 3.62462
R11130 VCTRL2.n65 VCTRL2.n64 3.62462
R11131 VCTRL2.n93 VCTRL2.n90 3.62462
R11132 VCTRL2.n92 VCTRL2.n91 3.62462
R11133 VCTRL2.n95 VCTRL2.n94 3.62462
R11134 VCTRL2.n33 VCTRL2.n32 3.62462
R11135 VCTRL2.n35 VCTRL2.n34 3.62462
R11136 VCTRL2.n49 VCTRL2.n48 3.62462
R11137 VCTRL2.n53 VCTRL2.n52 3.62462
R11138 VCTRL2.n55 VCTRL2.n54 3.62462
R11139 VCTRL2.n51 VCTRL2.n50 3.62462
R11140 VCTRL2.n122 VCTRL2.n121 2.2505
R11141 VCTRL2.n3 VCTRL2.n2 2.2505
R11142 VCTRL2.n125 VCTRL2.n124 1.5049
R11143 VCTRL2 VCTRL2.n0 1.16594
R11144 VCTRL2 VCTRL2.n62 1.16341
R11145 VCTRL2.n122 VCTRL2.n119 1.05045
R11146 VCTRL2.n61 VCTRL2.n60 0.984409
R11147 VCTRL2.n120 VCTRL2 0.936261
R11148 VCTRL2.n1 VCTRL2 0.936261
R11149 VCTRL2.n125 VCTRL2 0.61117
R11150 VCTRL2.n119 VCTRL2.n114 0.442081
R11151 VCTRL2.n60 VCTRL2.n55 0.441056
R11152 VCTRL2.n8 VCTRL2.n7 0.404715
R11153 VCTRL2.n36 VCTRL2.n35 0.404715
R11154 VCTRL2.n103 VCTRL2.n102 0.404539
R11155 VCTRL2.n39 VCTRL2.n38 0.404539
R11156 VCTRL2.n46 VCTRL2.n36 0.401155
R11157 VCTRL2.n9 VCTRL2.n8 0.401155
R11158 VCTRL2.n40 VCTRL2.n39 0.401155
R11159 VCTRL2.n104 VCTRL2.n103 0.400353
R11160 VCTRL2.n70 VCTRL2.n69 0.400178
R11161 VCTRL2.n47 VCTRL2.n46 0.398905
R11162 VCTRL2.n10 VCTRL2.n9 0.398484
R11163 VCTRL2.n55 VCTRL2.n47 0.397919
R11164 VCTRL2.n114 VCTRL2.n105 0.397919
R11165 VCTRL2.n105 VCTRL2.n104 0.397753
R11166 VCTRL2.n110 VCTRL2.n109 0.397744
R11167 VCTRL2.n7 VCTRL2.n6 0.389969
R11168 VCTRL2.n102 VCTRL2.n101 0.389723
R11169 VCTRL2.n38 VCTRL2.n37 0.389723
R11170 VCTRL2.n35 VCTRL2.n28 0.389547
R11171 VCTRL2.n32 VCTRL2.n31 0.389547
R11172 VCTRL2 VCTRL2.n125 0.10046
R11173 VCTRL2.n123 VCTRL2.n62 0.0698976
R11174 VCTRL2.n3 VCTRL2.n0 0.0695909
R11175 VCTRL2.n121 VCTRL2 0.0362534
R11176 VCTRL2.n2 VCTRL2 0.0362534
R11177 VCTRL2.n123 VCTRL2.n122 0.0124277
R11178 VCTRL2.n61 VCTRL2.n3 0.00395428
R11179 VCTRL2.n121 VCTRL2.n120 0.00173288
R11180 VCTRL2.n2 VCTRL2.n1 0.00173288
R11181 a_25706_n567.n90 a_25706_n567.n89 9.67588
R11182 a_25706_n567.n42 a_25706_n567.n41 3.74413
R11183 a_25706_n567.n26 a_25706_n567.n25 3.74025
R11184 a_25706_n567.n8 a_25706_n567.n12 3.72928
R11185 a_25706_n567.n9 a_25706_n567.n14 3.71799
R11186 a_25706_n567.n7 a_25706_n567.n6 3.60834
R11187 a_25706_n567.n21 a_25706_n567.t38 3.2765
R11188 a_25706_n567.n21 a_25706_n567.n20 3.2765
R11189 a_25706_n567.n23 a_25706_n567.t31 3.2765
R11190 a_25706_n567.n23 a_25706_n567.n22 3.2765
R11191 a_25706_n567.n70 a_25706_n567.t46 3.2765
R11192 a_25706_n567.n70 a_25706_n567.n69 3.2765
R11193 a_25706_n567.n67 a_25706_n567.t54 3.2765
R11194 a_25706_n567.n67 a_25706_n567.n66 3.2765
R11195 a_25706_n567.n63 a_25706_n567.t48 3.2765
R11196 a_25706_n567.n63 a_25706_n567.n62 3.2765
R11197 a_25706_n567.n60 a_25706_n567.t41 3.2765
R11198 a_25706_n567.n60 a_25706_n567.n59 3.2765
R11199 a_25706_n567.n56 a_25706_n567.t59 3.2765
R11200 a_25706_n567.n56 a_25706_n567.n55 3.2765
R11201 a_25706_n567.n87 a_25706_n567.t52 3.2765
R11202 a_25706_n567.n87 a_25706_n567.n86 3.2765
R11203 a_25706_n567.n84 a_25706_n567.t43 3.2765
R11204 a_25706_n567.n84 a_25706_n567.n83 3.2765
R11205 a_25706_n567.n80 a_25706_n567.t57 3.2765
R11206 a_25706_n567.n80 a_25706_n567.n79 3.2765
R11207 a_25706_n567.n77 a_25706_n567.t51 3.2765
R11208 a_25706_n567.n77 a_25706_n567.n76 3.2765
R11209 a_25706_n567.n73 a_25706_n567.t42 3.2765
R11210 a_25706_n567.n73 a_25706_n567.n72 3.2765
R11211 a_25706_n567.n36 a_25706_n567.t35 3.2765
R11212 a_25706_n567.n36 a_25706_n567.n35 3.2765
R11213 a_25706_n567.n34 a_25706_n567.t4 3.2765
R11214 a_25706_n567.n34 a_25706_n567.n33 3.2765
R11215 a_25706_n567.n30 a_25706_n567.t34 3.2765
R11216 a_25706_n567.n30 a_25706_n567.n29 3.2765
R11217 a_25706_n567.n28 a_25706_n567.t16 3.2765
R11218 a_25706_n567.n28 a_25706_n567.n27 3.2765
R11219 a_25706_n567.n19 a_25706_n567.t13 3.2765
R11220 a_25706_n567.n19 a_25706_n567.n18 3.2765
R11221 a_25706_n567.n12 a_25706_n567.t6 3.2765
R11222 a_25706_n567.n12 a_25706_n567.n11 3.2765
R11223 a_25706_n567.n16 a_25706_n567.t1 3.2765
R11224 a_25706_n567.n16 a_25706_n567.n15 3.2765
R11225 a_25706_n567.n14 a_25706_n567.t33 3.2765
R11226 a_25706_n567.n14 a_25706_n567.n13 3.2765
R11227 a_25706_n567.n4 a_25706_n567.t21 3.2765
R11228 a_25706_n567.n4 a_25706_n567.n3 3.2765
R11229 a_25706_n567.n39 a_25706_n567.t22 3.2765
R11230 a_25706_n567.n39 a_25706_n567.n38 3.2765
R11231 a_25706_n567.n46 a_25706_n567.t27 3.2765
R11232 a_25706_n567.n46 a_25706_n567.n45 3.2765
R11233 a_25706_n567.n44 a_25706_n567.t8 3.2765
R11234 a_25706_n567.n44 a_25706_n567.n43 3.2765
R11235 a_25706_n567.n41 a_25706_n567.t0 3.2765
R11236 a_25706_n567.n41 a_25706_n567.n40 3.2765
R11237 a_25706_n567.n49 a_25706_n567.t15 3.2765
R11238 a_25706_n567.n49 a_25706_n567.n48 3.2765
R11239 a_25706_n567.n2 a_25706_n567.t25 3.2765
R11240 a_25706_n567.n2 a_25706_n567.n1 3.2765
R11241 a_25706_n567.n52 a_25706_n567.t17 3.2765
R11242 a_25706_n567.n52 a_25706_n567.n51 3.2765
R11243 a_25706_n567.n25 a_25706_n567.t9 3.2765
R11244 a_25706_n567.n25 a_25706_n567.n24 3.2765
R11245 a_25706_n567.n94 a_25706_n567.t32 3.2765
R11246 a_25706_n567.n95 a_25706_n567.n94 3.2765
R11247 a_25706_n567.n74 a_25706_n567.n73 3.1505
R11248 a_25706_n567.n78 a_25706_n567.n77 3.1505
R11249 a_25706_n567.n81 a_25706_n567.n80 3.1505
R11250 a_25706_n567.n85 a_25706_n567.n84 3.1505
R11251 a_25706_n567.n88 a_25706_n567.n87 3.1505
R11252 a_25706_n567.n57 a_25706_n567.n56 3.1505
R11253 a_25706_n567.n61 a_25706_n567.n60 3.1505
R11254 a_25706_n567.n64 a_25706_n567.n63 3.1505
R11255 a_25706_n567.n68 a_25706_n567.n67 3.1505
R11256 a_25706_n567.n71 a_25706_n567.n70 3.1505
R11257 a_25706_n567.n47 a_25706_n567.n46 3.1505
R11258 a_25706_n567.n50 a_25706_n567.n49 3.1505
R11259 a_25706_n567.n53 a_25706_n567.n52 3.1505
R11260 a_25706_n567.n5 a_25706_n567.n4 3.1505
R11261 a_25706_n567.n31 a_25706_n567.n30 3.1505
R11262 a_25706_n567.n37 a_25706_n567.n36 3.1505
R11263 a_25706_n567.n92 a_25706_n567.n23 3.1505
R11264 a_25706_n567.n94 a_25706_n567.n93 3.1505
R11265 a_25706_n567.n17 a_25706_n567.n10 2.34866
R11266 a_25706_n567.n8 a_25706_n567.n19 1.8475
R11267 a_25706_n567.n42 a_25706_n567.n44 1.84743
R11268 a_25706_n567.n6 a_25706_n567.n2 1.84743
R11269 a_25706_n567.n26 a_25706_n567.n28 1.8474
R11270 a_25706_n567.n0 a_25706_n567.n39 1.84737
R11271 a_25706_n567.n32 a_25706_n567.n34 1.84737
R11272 a_25706_n567.n7 a_25706_n567.n21 1.84737
R11273 a_25706_n567.n10 a_25706_n567.n16 1.84618
R11274 a_25706_n567.n8 a_25706_n567.n17 1.48093
R11275 a_25706_n567.n54 a_25706_n567.n53 0.899822
R11276 a_25706_n567.n92 a_25706_n567.n91 0.899822
R11277 a_25706_n567.n81 a_25706_n567.n78 0.758798
R11278 a_25706_n567.n64 a_25706_n567.n61 0.758798
R11279 a_25706_n567.n89 a_25706_n567.n71 0.724996
R11280 a_25706_n567.n88 a_25706_n567.n85 0.7205
R11281 a_25706_n567.n71 a_25706_n567.n68 0.7205
R11282 a_25706_n567.n89 a_25706_n567.n88 0.636952
R11283 a_25706_n567.n93 a_25706_n567.n8 0.618999
R11284 a_25706_n567.n50 a_25706_n567.n0 0.607482
R11285 a_25706_n567.n37 a_25706_n567.n32 0.604163
R11286 a_25706_n567.n7 a_25706_n567.n92 0.60198
R11287 a_25706_n567.n93 a_25706_n567.n7 0.601843
R11288 a_25706_n567.n32 a_25706_n567.n31 0.598752
R11289 a_25706_n567.n31 a_25706_n567.n26 0.597003
R11290 a_25706_n567.n0 a_25706_n567.n47 0.595434
R11291 a_25706_n567.n47 a_25706_n567.n42 0.593116
R11292 a_25706_n567.n6 a_25706_n567.n5 0.593116
R11293 a_25706_n567.n75 a_25706_n567.n74 0.555819
R11294 a_25706_n567.n58 a_25706_n567.n57 0.555819
R11295 a_25706_n567.n85 a_25706_n567.n82 0.551989
R11296 a_25706_n567.n68 a_25706_n567.n65 0.551989
R11297 a_25706_n567.n90 a_25706_n567.n54 0.3917
R11298 a_25706_n567.n82 a_25706_n567.n81 0.283904
R11299 a_25706_n567.n65 a_25706_n567.n64 0.283904
R11300 a_25706_n567.n78 a_25706_n567.n75 0.280074
R11301 a_25706_n567.n61 a_25706_n567.n58 0.280074
R11302 a_25706_n567.n91 a_25706_n567.n90 0.2621
R11303 a_25706_n567.n54 a_25706_n567.n50 0.247022
R11304 a_25706_n567.n91 a_25706_n567.n37 0.247022
R11305 a_25706_n567.n10 a_25706_n567.n9 0.0460206
R11306 DN_INPUT.t0 DN_INPUT.t3 44.058
R11307 DN_INPUT.n0 DN_INPUT.t1 38.8649
R11308 DN_INPUT.t1 DN_INPUT.t0 28.6791
R11309 DN_INPUT.n0 DN_INPUT.t2 7.3005
R11310 DN_INPUT DN_INPUT.n0 5.27587
R11311 a_27875_9714.t6 a_27875_9714.t7 44.058
R11312 a_27875_9714.n1 a_27875_9714.t8 34.6465
R11313 a_27875_9714.n1 a_27875_9714.t6 15.1219
R11314 a_27875_9714.n5 a_27875_9714.t3 5.29595
R11315 a_27875_9714.n2 a_27875_9714.n0 4.97104
R11316 a_27875_9714.n2 a_27875_9714.n1 4.16767
R11317 a_27875_9714.n5 a_27875_9714.n4 3.01333
R11318 a_27875_9714.n7 a_27875_9714.n6 3.01333
R11319 a_27875_9714.n4 a_27875_9714.t4 1.6255
R11320 a_27875_9714.n4 a_27875_9714.n3 1.6255
R11321 a_27875_9714.n7 a_27875_9714.t0 1.6255
R11322 a_27875_9714.n8 a_27875_9714.n7 1.6255
R11323 a_27875_9714.n6 a_27875_9714.n5 0.845717
R11324 a_27875_9714.n6 a_27875_9714.n2 0.423109
R11325 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n9 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n8 15.8172
R11326 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n11 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n10 15.8172
R11327 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n10 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n9 15.8172
R11328 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n9 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t37 14.8925
R11329 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n10 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t43 14.8925
R11330 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n17 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n16 12.2457
R11331 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n16 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n14 12.2457
R11332 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n14 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n12 12.2457
R11333 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n18 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t58 11.6285
R11334 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n52 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t41 9.5787
R11335 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n49 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t45 9.55768
R11336 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n12 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t56 8.9065
R11337 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n14 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t42 8.9065
R11338 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n16 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t47 8.9065
R11339 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n17 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t35 8.9065
R11340 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n64 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n60 8.86038
R11341 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n9 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t33 8.6145
R11342 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n8 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t46 8.6145
R11343 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n10 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t39 8.6145
R11344 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n11 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t54 8.59715
R11345 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n52 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t52 8.57144
R11346 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n53 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t57 8.57144
R11347 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n54 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t50 8.57144
R11348 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n31 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t0 8.54728
R11349 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n5 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t38 8.52112
R11350 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n0 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t53 8.52112
R11351 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n2 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t32 8.52112
R11352 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n7 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t48 8.52112
R11353 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n51 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t55 8.51092
R11354 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n50 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t34 8.51092
R11355 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n49 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t31 8.51092
R11356 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n0 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t40 8.35286
R11357 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n12 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t49 8.3225
R11358 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t58 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n17 8.3225
R11359 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n7 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t36 8.31073
R11360 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n2 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t44 8.31073
R11361 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n5 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t51 8.31073
R11362 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n22 7.05764
R11363 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t27 6.83153
R11364 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n31 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t29 6.78441
R11365 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n35 6.45366
R11366 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n29 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n28 6.20932
R11367 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n21 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t23 5.87174
R11368 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n76 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t16 5.30249
R11369 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n42 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n41 5.28839
R11370 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n1 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t15 4.92134
R11371 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n58 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t9 4.89657
R11372 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n44 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t12 4.89616
R11373 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n73 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n36 4.87698
R11374 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n6 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n57 4.63042
R11375 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n70 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n56 4.63037
R11376 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n45 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n1 4.22693
R11377 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n18 4.223
R11378 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n46 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n42 4.02972
R11379 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n34 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n33 4.0288
R11380 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n74 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n73 3.96222
R11381 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t42 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n13 3.6505
R11382 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t47 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n15 3.6505
R11383 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n62 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t5 3.6405
R11384 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n62 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n61 3.6405
R11385 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n78 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t13 3.6405
R11386 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n78 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n79 3.6405
R11387 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n38 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t10 3.6405
R11388 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n38 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n37 3.6405
R11389 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n33 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t28 3.6405
R11390 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n33 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n32 3.6405
R11391 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n67 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t6 3.6405
R11392 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n67 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n66 3.6405
R11393 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n24 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n23 3.47613
R11394 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n20 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n19 3.47609
R11395 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n26 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n25 3.47601
R11396 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n21 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n20 3.39857
R11397 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n45 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n77 3.27464
R11398 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n18 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n11 3.1807
R11399 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n75 3.16877
R11400 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n47 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n76 2.96981
R11401 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n26 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t18 2.8627
R11402 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n20 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t22 2.86263
R11403 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n24 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t25 2.8626
R11404 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n69 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n68 2.60609
R11405 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n24 2.48343
R11406 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n30 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN 2.30073
R11407 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n75 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN 2.29178
R11408 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n27 2.24606
R11409 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n6 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n69 2.24505
R11410 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n68 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n67 4.81682
R11411 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n64 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n63 3.77141
R11412 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n1 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n44 2.52627
R11413 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n65 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n59 1.8072
R11414 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n48 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n40 1.76824
R11415 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n63 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n62 1.65829
R11416 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n39 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n38 1.65829
R11417 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n55 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n51 1.6131
R11418 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n55 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n54 1.57488
R11419 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n44 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n43 1.53436
R11420 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n71 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n70 1.51602
R11421 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n59 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n58 1.49487
R11422 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n36 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n34 1.32452
R11423 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n77 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n78 1.25757
R11424 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n40 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n39 1.12313
R11425 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n4 1.05601
R11426 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n30 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n29 1.01067
R11427 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n50 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n49 0.996664
R11428 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n0 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n5 0.992966
R11429 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n21 0.983287
R11430 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n27 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n26 0.982856
R11431 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n2 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n0 0.975705
R11432 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n72 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n71 0.968726
R11433 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n73 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n72 0.955885
R11434 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n53 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n52 0.953514
R11435 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n29 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n3 0.911933
R11436 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n46 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n45 0.856289
R11437 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n48 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n47 0.843442
R11438 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n68 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n65 0.8015
R11439 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n70 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n6 0.741046
R11440 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n34 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n31 0.710717
R11441 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n71 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n7 0.698938
R11442 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n72 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n48 0.656959
R11443 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n47 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n46 0.398395
R11444 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n65 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n64 0.3875
R11445 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n54 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n53 0.364199
R11446 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n74 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n30 0.362023
R11447 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n7 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n2 0.359267
R11448 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n51 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n50 0.323514
R11449 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n5 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n55 0.321048
R11450 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n75 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n74 0.271283
R11451 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n36 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN 0.147028
R11452 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n73 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n72 15.8172
R11453 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n74 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n73 15.8172
R11454 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n75 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n74 15.8172
R11455 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n73 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t50 14.8925
R11456 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n74 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t43 14.8925
R11457 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n81 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n80 12.2457
R11458 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n80 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n78 12.2457
R11459 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n78 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n76 12.2457
R11460 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n82 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t37 11.6285
R11461 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n36 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t35 9.07401
R11462 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n40 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t45 8.94931
R11463 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n35 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t32 8.91612
R11464 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n34 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t58 8.91612
R11465 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n32 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t40 8.91612
R11466 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n76 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t53 8.9065
R11467 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n78 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t47 8.9065
R11468 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n80 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t36 8.9065
R11469 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n81 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t57 8.9065
R11470 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n30 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t54 8.88203
R11471 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n38 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t42 8.78079
R11472 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n41 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t39 8.78079
R11473 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n37 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t46 8.76459
R11474 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n36 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t44 8.76459
R11475 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n11 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n9 8.71932
R11476 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n31 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t55 8.71352
R11477 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n2 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t51 8.71352
R11478 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n73 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t49 8.6145
R11479 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n72 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t56 8.6145
R11480 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n74 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t38 8.6145
R11481 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n75 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t31 8.59715
R11482 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n53 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t1 8.51681
R11483 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n0 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t41 8.50287
R11484 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t52 8.38543
R11485 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n76 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t33 8.3225
R11486 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t37 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n81 8.3225
R11487 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n39 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t34 8.30117
R11488 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n7 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n6 8.23463
R11489 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n30 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t48 7.39905
R11490 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n26 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n25 6.43594
R11491 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n20 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n19 6.42269
R11492 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n5 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n27 6.3977
R11493 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n1 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n33 6.02773
R11494 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n17 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t18 5.83006
R11495 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n66 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n52 5.43818
R11496 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n20 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n14 5.23259
R11497 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n65 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n64 4.89653
R11498 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n42 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t10 4.89315
R11499 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t26 4.88822
R11500 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n11 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n10 4.72831
R11501 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n18 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t17 4.70462
R11502 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n19 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t20 4.70346
R11503 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n49 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n48 4.53146
R11504 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n82 4.22145
R11505 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n55 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t11 4.04969
R11506 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n59 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n60 4.00854
R11507 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n44 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n43 4.00757
R11508 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n29 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t12 4.00481
R11509 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n12 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n8 3.90715
R11510 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n71 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n70 3.79925
R11511 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n17 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n16 3.77445
R11512 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n47 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n46 3.76989
R11513 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n26 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n24 3.76191
R11514 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n24 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t27 3.7183
R11515 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t47 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n77 3.6505
R11516 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t36 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n79 3.6505
R11517 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n62 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t6 3.6405
R11518 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n62 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n61 3.6405
R11519 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n57 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t14 3.6405
R11520 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n57 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n56 3.6405
R11521 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n52 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t7 3.6405
R11522 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n52 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n51 3.6405
R11523 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n14 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t19 3.47629
R11524 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n16 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t16 3.47627
R11525 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n21 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n20 3.3208
R11526 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n47 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t3 3.26228
R11527 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n24 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n23 3.25601
R11528 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n82 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n75 3.1807
R11529 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n5 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN 3.15982
R11530 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n70 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n22 3.14573
R11531 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n59 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n58 2.8959
R11532 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n18 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n17 2.88663
R11533 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n16 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n15 2.86148
R11534 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n14 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n13 2.86147
R11535 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n21 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n12 2.83772
R11536 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n49 2.75932
R11537 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n66 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n7 2.62155
R11538 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n71 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN 2.36584
R11539 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n70 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n69 2.35159
R11540 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n22 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN 2.30603
R11541 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n45 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n44 2.2491
R11542 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n54 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n55 2.24586
R11543 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n68 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n67 2.03309
R11544 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n71 1.93478
R11545 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n49 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n45 1.85135
R11546 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n7 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n63 1.79127
R11547 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n53 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n54 1.76701
R11548 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n58 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n57 1.65928
R11549 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n7 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n53 1.6295
R11550 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n50 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n29 1.50938
R11551 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n63 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n65 1.495
R11552 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n69 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n28 1.47463
R11553 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n60 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n62 1.25653
R11554 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n67 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n66 1.22576
R11555 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n0 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n4 1.19023
R11556 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n53 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n59 1.1585
R11557 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n42 1.1379
R11558 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n48 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n47 1.00671
R11559 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n28 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n5 0.931417
R11560 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n5 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n26 0.878898
R11561 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n68 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n50 0.836865
R11562 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n39 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n38 0.650226
R11563 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n69 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n68 0.597881
R11564 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n22 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n21 0.488268
R11565 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n2 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n32 0.487486
R11566 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n12 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n11 0.477758
R11567 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n19 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n18 0.472393
R11568 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n50 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n0 0.415098
R11569 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n2 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n1 0.384677
R11570 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n3 0.384538
R11571 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n41 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n40 0.345705
R11572 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n31 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n30 0.345705
R11573 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n41 0.34324
R11574 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n37 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n36 0.342007
R11575 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n35 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n34 0.342007
R11576 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n34 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n2 0.33461
R11577 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n38 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n37 0.325979
R11578 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n40 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n39 0.318582
R11579 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n32 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n31 0.312418
R11580 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n0 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n35 0.312418
R11581 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n23 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t18 23.6945
R11582 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t20 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n24 23.6945
R11583 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n24 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n23 18.8035
R11584 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n21 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n19 15.8172
R11585 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n21 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n20 15.8172
R11586 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n20 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n16 15.8172
R11587 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n19 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t13 14.8925
R11588 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t21 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n21 14.8925
R11589 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n20 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t16 14.8925
R11590 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n25 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n17 12.2457
R11591 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n22 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n17 12.2457
R11592 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n22 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n18 12.2457
R11593 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n26 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t15 11.6285
R11594 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n18 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t18 8.9065
R11595 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t17 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n22 8.9065
R11596 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t22 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n17 8.9065
R11597 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n25 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t20 8.9065
R11598 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n21 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t19 8.6145
R11599 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n19 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t23 8.6145
R11600 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n20 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t14 8.6145
R11601 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n16 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t12 8.59715
R11602 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t13 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n18 8.3225
R11603 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n22 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t21 8.3225
R11604 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t16 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n17 8.3225
R11605 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t15 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n25 8.3225
R11606 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n26 4.223
R11607 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n23 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t17 3.6505
R11608 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n24 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t22 3.6505
R11609 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n11 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t7 3.6405
R11610 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n11 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n10 3.6405
R11611 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n5 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t9 3.6405
R11612 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n5 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n4 3.6405
R11613 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n7 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t4 3.6405
R11614 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n7 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n6 3.6405
R11615 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n13 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t6 3.6405
R11616 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n13 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n12 3.6405
R11617 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n15 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n1 3.50463
R11618 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n9 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n3 3.50463
R11619 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n1 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t1 3.2765
R11620 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n1 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n0 3.2765
R11621 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n3 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t3 3.2765
R11622 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n3 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n2 3.2765
R11623 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n26 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n16 3.1807
R11624 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n8 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n7 3.06224
R11625 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n14 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n11 3.06224
R11626 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n8 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n5 2.6005
R11627 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n14 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n13 2.6005
R11628 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n15 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n9 0.798761
R11629 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n15 0.562022
R11630 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n9 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n8 0.18637
R11631 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n15 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n14 0.18637
R11632 mux_magic_3.OR_magic_0.A.t5 mux_magic_3.OR_magic_0.A.t7 44.6331
R11633 mux_magic_3.OR_magic_0.A.t4 mux_magic_3.OR_magic_0.A.t6 31.5469
R11634 mux_magic_3.OR_magic_0.A.t6 mux_magic_3.OR_magic_0.A.t3 28.6791
R11635 mux_magic_3.OR_magic_0.A.n0 mux_magic_3.OR_magic_0.A.t5 19.3585
R11636 mux_magic_3.OR_magic_0.A.n0 mux_magic_3.OR_magic_0.A.t4 12.1889
R11637 mux_magic_3.OR_magic_0.A mux_magic_3.OR_magic_0.A.n1 5.0317
R11638 mux_magic_3.OR_magic_0.A mux_magic_3.OR_magic_0.A.n0 4.23754
R11639 mux_magic_3.OR_magic_0.A mux_magic_3.OR_magic_0.A.n3 3.36245
R11640 mux_magic_3.OR_magic_0.A.n3 mux_magic_3.OR_magic_0.A.t1 1.6255
R11641 mux_magic_3.OR_magic_0.A.n3 mux_magic_3.OR_magic_0.A.n2 1.6255
R11642 a_21443_9476.t6 a_21443_9476.t8 31.5469
R11643 a_21443_9476.n2 a_21443_9476.t6 13.227
R11644 a_21443_9476.n2 a_21443_9476.t7 13.138
R11645 a_21443_9476.n0 a_21443_9476.t0 6.53038
R11646 a_21443_9476.n0 a_21443_9476.n2 4.33404
R11647 a_21443_9476.n6 a_21443_9476.n3 4.2255
R11648 a_21443_9476.n8 a_21443_9476.n7 4.2255
R11649 a_21443_9476.n6 a_21443_9476.n5 3.81956
R11650 a_21443_9476.n0 a_21443_9476.n1 2.62675
R11651 a_21443_9476.n5 a_21443_9476.t5 1.6255
R11652 a_21443_9476.n5 a_21443_9476.n4 1.6255
R11653 a_21443_9476.n7 a_21443_9476.n6 0.947457
R11654 a_21443_9476.n7 a_21443_9476.n0 0.600587
R11655 a_43528_12082.t0 a_43528_12082.t1 12.9675
R11656 a_43828_11460.t0 a_43828_11460.t1 12.9675
R11657 mux_magic_2.AND2_magic_0.A.t12 mux_magic_2.AND2_magic_0.A.t9 144.929
R11658 mux_magic_2.AND2_magic_0.A.t10 mux_magic_2.AND2_magic_0.A.t11 44.058
R11659 mux_magic_2.AND2_magic_0.A.n2 mux_magic_2.AND2_magic_0.A.t12 14.7309
R11660 mux_magic_2.AND2_magic_0.A.n2 mux_magic_2.AND2_magic_0.A.t10 13.9487
R11661 mux_magic_2.AND2_magic_0.A mux_magic_2.AND2_magic_0.A.n2 9.83788
R11662 mux_magic_2.AND2_magic_0.A.n1 mux_magic_2.AND2_magic_0.A.n4 4.99061
R11663 mux_magic_2.AND2_magic_0.A mux_magic_2.AND2_magic_0.A.n11 4.5405
R11664 mux_magic_2.AND2_magic_0.A.n1 mux_magic_2.AND2_magic_0.A.n3 4.2255
R11665 mux_magic_2.AND2_magic_0.A.n0 mux_magic_2.AND2_magic_0.A.n10 3.52811
R11666 mux_magic_2.AND2_magic_0.A.n0 mux_magic_2.AND2_magic_0.A.n6 3.30485
R11667 mux_magic_2.AND2_magic_0.A.n0 mux_magic_2.AND2_magic_0.A.n8 2.6005
R11668 mux_magic_2.AND2_magic_0.A.n6 mux_magic_2.AND2_magic_0.A.t6 1.6255
R11669 mux_magic_2.AND2_magic_0.A.n6 mux_magic_2.AND2_magic_0.A.n5 1.6255
R11670 mux_magic_2.AND2_magic_0.A.n8 mux_magic_2.AND2_magic_0.A.t3 1.6255
R11671 mux_magic_2.AND2_magic_0.A.n8 mux_magic_2.AND2_magic_0.A.n7 1.6255
R11672 mux_magic_2.AND2_magic_0.A.n10 mux_magic_2.AND2_magic_0.A.t0 1.463
R11673 mux_magic_2.AND2_magic_0.A.n10 mux_magic_2.AND2_magic_0.A.n9 1.463
R11674 mux_magic_2.AND2_magic_0.A.n1 mux_magic_2.AND2_magic_0.A.n0 1.19985
R11675 mux_magic_2.AND2_magic_0.A mux_magic_2.AND2_magic_0.A.n1 0.819535
R11676 a_20097_11741.n3 a_20097_11741.n1 6.04375
R11677 a_20097_11741.n3 a_20097_11741.n2 1.55052
R11678 a_20097_11741.n1 a_20097_11741.t3 1.463
R11679 a_20097_11741.n1 a_20097_11741.n0 1.463
R11680 a_20097_11741.t0 a_20097_11741.n3 1.3335
R11681 a_19897_11741.t7 a_19897_11741.t8 44.058
R11682 a_19897_11741.n3 a_19897_11741.t6 34.6465
R11683 a_19897_11741.n3 a_19897_11741.t7 15.1219
R11684 a_19897_11741.n6 a_19897_11741.t2 5.29595
R11685 a_19897_11741.n4 a_19897_11741.n2 4.97104
R11686 a_19897_11741.n4 a_19897_11741.n3 4.16767
R11687 a_19897_11741.n5 a_19897_11741.n1 3.01333
R11688 a_19897_11741.n7 a_19897_11741.n6 3.01333
R11689 a_19897_11741.n1 a_19897_11741.t5 1.6255
R11690 a_19897_11741.n1 a_19897_11741.n0 1.6255
R11691 a_19897_11741.n7 a_19897_11741.t0 1.6255
R11692 a_19897_11741.n8 a_19897_11741.n7 1.6255
R11693 a_19897_11741.n6 a_19897_11741.n5 0.845717
R11694 a_19897_11741.n5 a_19897_11741.n4 0.423109
R11695 a_25557_8739.n0 a_25557_8739.t3 24.1084
R11696 a_25557_8739.n1 a_25557_8739.t5 12.5565
R11697 a_25557_8739.n0 a_25557_8739.t4 8.6145
R11698 a_25557_8739.n2 a_25557_8739.t0 6.71215
R11699 a_25557_8739.n2 a_25557_8739.n1 4.46748
R11700 a_25557_8739.n3 a_25557_8739.t1 3.6405
R11701 a_25557_8739.n4 a_25557_8739.n3 3.6405
R11702 a_25557_8739.n3 a_25557_8739.n2 2.83724
R11703 a_25557_8739.n1 a_25557_8739.n0 1.8985
R11704 a_34443_2598.n69 a_34443_2598.n51 9.67588
R11705 a_34443_2598.n4 a_34443_2598.n89 3.7286
R11706 a_34443_2598.n15 a_34443_2598.n14 3.71799
R11707 a_34443_2598.n2 a_34443_2598.n59 3.71473
R11708 a_34443_2598.n1 a_34443_2598.n75 3.70973
R11709 a_34443_2598.n87 a_34443_2598.t23 3.2765
R11710 a_34443_2598.n87 a_34443_2598.n86 3.2765
R11711 a_34443_2598.n12 a_34443_2598.t6 3.2765
R11712 a_34443_2598.n12 a_34443_2598.n11 3.2765
R11713 a_34443_2598.n9 a_34443_2598.t28 3.2765
R11714 a_34443_2598.n9 a_34443_2598.n8 3.2765
R11715 a_34443_2598.n7 a_34443_2598.t20 3.2765
R11716 a_34443_2598.n7 a_34443_2598.n6 3.2765
R11717 a_34443_2598.n66 a_34443_2598.t8 3.2765
R11718 a_34443_2598.n66 a_34443_2598.n65 3.2765
R11719 a_34443_2598.n53 a_34443_2598.t12 3.2765
R11720 a_34443_2598.n53 a_34443_2598.n52 3.2765
R11721 a_34443_2598.n55 a_34443_2598.t24 3.2765
R11722 a_34443_2598.n55 a_34443_2598.n54 3.2765
R11723 a_34443_2598.n80 a_34443_2598.t38 3.2765
R11724 a_34443_2598.n80 a_34443_2598.n79 3.2765
R11725 a_34443_2598.n71 a_34443_2598.t32 3.2765
R11726 a_34443_2598.n71 a_34443_2598.n70 3.2765
R11727 a_34443_2598.n18 a_34443_2598.t42 3.2765
R11728 a_34443_2598.n18 a_34443_2598.n17 3.2765
R11729 a_34443_2598.n20 a_34443_2598.t58 3.2765
R11730 a_34443_2598.n20 a_34443_2598.n19 3.2765
R11731 a_34443_2598.n26 a_34443_2598.t50 3.2765
R11732 a_34443_2598.n26 a_34443_2598.n25 3.2765
R11733 a_34443_2598.n22 a_34443_2598.t43 3.2765
R11734 a_34443_2598.n22 a_34443_2598.n21 3.2765
R11735 a_34443_2598.n24 a_34443_2598.t47 3.2765
R11736 a_34443_2598.n24 a_34443_2598.n23 3.2765
R11737 a_34443_2598.n39 a_34443_2598.t55 3.2765
R11738 a_34443_2598.n39 a_34443_2598.n38 3.2765
R11739 a_34443_2598.n41 a_34443_2598.t59 3.2765
R11740 a_34443_2598.n41 a_34443_2598.n40 3.2765
R11741 a_34443_2598.n43 a_34443_2598.t40 3.2765
R11742 a_34443_2598.n43 a_34443_2598.n42 3.2765
R11743 a_34443_2598.n35 a_34443_2598.t56 3.2765
R11744 a_34443_2598.n35 a_34443_2598.n34 3.2765
R11745 a_34443_2598.n37 a_34443_2598.t44 3.2765
R11746 a_34443_2598.n37 a_34443_2598.n36 3.2765
R11747 a_34443_2598.n84 a_34443_2598.t1 3.2765
R11748 a_34443_2598.n84 a_34443_2598.n83 3.2765
R11749 a_34443_2598.n73 a_34443_2598.t4 3.2765
R11750 a_34443_2598.n73 a_34443_2598.n72 3.2765
R11751 a_34443_2598.n77 a_34443_2598.t30 3.2765
R11752 a_34443_2598.n77 a_34443_2598.n76 3.2765
R11753 a_34443_2598.n75 a_34443_2598.t36 3.2765
R11754 a_34443_2598.n75 a_34443_2598.n74 3.2765
R11755 a_34443_2598.n57 a_34443_2598.t33 3.2765
R11756 a_34443_2598.n57 a_34443_2598.n56 3.2765
R11757 a_34443_2598.n61 a_34443_2598.t10 3.2765
R11758 a_34443_2598.n61 a_34443_2598.n60 3.2765
R11759 a_34443_2598.n59 a_34443_2598.t22 3.2765
R11760 a_34443_2598.n59 a_34443_2598.n58 3.2765
R11761 a_34443_2598.n14 a_34443_2598.t18 3.2765
R11762 a_34443_2598.n14 a_34443_2598.n13 3.2765
R11763 a_34443_2598.n91 a_34443_2598.t0 3.2765
R11764 a_34443_2598.n91 a_34443_2598.n90 3.2765
R11765 a_34443_2598.n89 a_34443_2598.t11 3.2765
R11766 a_34443_2598.n89 a_34443_2598.n88 3.2765
R11767 a_34443_2598.n93 a_34443_2598.t13 3.2765
R11768 a_34443_2598.n94 a_34443_2598.n93 3.2765
R11769 a_34443_2598.n49 a_34443_2598.n37 3.1505
R11770 a_34443_2598.n50 a_34443_2598.n35 3.1505
R11771 a_34443_2598.n44 a_34443_2598.n43 3.1505
R11772 a_34443_2598.n46 a_34443_2598.n41 3.1505
R11773 a_34443_2598.n47 a_34443_2598.n39 3.1505
R11774 a_34443_2598.n29 a_34443_2598.n24 3.1505
R11775 a_34443_2598.n30 a_34443_2598.n22 3.1505
R11776 a_34443_2598.n27 a_34443_2598.n26 3.1505
R11777 a_34443_2598.n32 a_34443_2598.n20 3.1505
R11778 a_34443_2598.n33 a_34443_2598.n18 3.1505
R11779 a_34443_2598.n85 a_34443_2598.n84 3.1505
R11780 a_34443_2598.n81 a_34443_2598.n71 3.1505
R11781 a_34443_2598.n78 a_34443_2598.n73 3.1505
R11782 a_34443_2598.n62 a_34443_2598.n57 3.1505
R11783 a_34443_2598.n64 a_34443_2598.n53 3.1505
R11784 a_34443_2598.n67 a_34443_2598.n66 3.1505
R11785 a_34443_2598.n10 a_34443_2598.n9 3.1505
R11786 a_34443_2598.n92 a_34443_2598.n87 3.1505
R11787 a_34443_2598.n4 a_34443_2598.n91 1.84747
R11788 a_34443_2598.n2 a_34443_2598.n61 1.84743
R11789 a_34443_2598.n1 a_34443_2598.n77 1.84737
R11790 a_34443_2598.n0 a_34443_2598.n80 1.84737
R11791 a_34443_2598.n63 a_34443_2598.n55 1.84737
R11792 a_34443_2598.n5 a_34443_2598.n7 1.84732
R11793 a_34443_2598.n93 a_34443_2598.n3 1.84728
R11794 a_34443_2598.n16 a_34443_2598.n12 1.84618
R11795 a_34443_2598.n85 a_34443_2598.n82 0.899822
R11796 a_34443_2598.n68 a_34443_2598.n67 0.899822
R11797 a_34443_2598.n47 a_34443_2598.n46 0.758798
R11798 a_34443_2598.n30 a_34443_2598.n29 0.758798
R11799 a_34443_2598.n51 a_34443_2598.n50 0.724996
R11800 a_34443_2598.n50 a_34443_2598.n49 0.7205
R11801 a_34443_2598.n33 a_34443_2598.n32 0.7205
R11802 a_34443_2598.n51 a_34443_2598.n33 0.636952
R11803 a_34443_2598.n16 a_34443_2598.n10 0.622339
R11804 a_34443_2598.n64 a_34443_2598.n63 0.607482
R11805 a_34443_2598.n81 a_34443_2598.n0 0.604163
R11806 a_34443_2598.n3 a_34443_2598.n85 0.602337
R11807 a_34443_2598.n63 a_34443_2598.n62 0.595434
R11808 a_34443_2598.n45 a_34443_2598.n44 0.555819
R11809 a_34443_2598.n28 a_34443_2598.n27 0.555819
R11810 a_34443_2598.n49 a_34443_2598.n48 0.551989
R11811 a_34443_2598.n32 a_34443_2598.n31 0.551989
R11812 a_34443_2598.n69 a_34443_2598.n68 0.378745
R11813 a_34443_2598.n48 a_34443_2598.n47 0.283904
R11814 a_34443_2598.n31 a_34443_2598.n30 0.283904
R11815 a_34443_2598.n46 a_34443_2598.n45 0.280074
R11816 a_34443_2598.n29 a_34443_2598.n28 0.280074
R11817 a_34443_2598.n82 a_34443_2598.n69 0.248582
R11818 a_34443_2598.n82 a_34443_2598.n81 0.247022
R11819 a_34443_2598.n68 a_34443_2598.n64 0.247022
R11820 a_34443_2598.n16 a_34443_2598.n15 0.0460206
R11821 a_34443_2598.n5 a_34443_2598.n3 3.58925
R11822 a_34443_2598.n78 a_34443_2598.n1 0.627536
R11823 a_34443_2598.n62 a_34443_2598.n2 0.622521
R11824 a_34443_2598.n92 a_34443_2598.n4 0.619689
R11825 a_34443_2598.n10 a_34443_2598.n5 0.609769
R11826 a_34443_2598.n3 a_34443_2598.n92 0.602476
R11827 a_34443_2598.n0 a_34443_2598.n78 0.598753
R11828 RES_74k_1.P.n98 RES_74k_1.P.n97 9.42182
R11829 RES_74k_1.P.n103 RES_74k_1.P.n102 9.3792
R11830 RES_74k_1.P.n110 RES_74k_1.P.n109 9.07899
R11831 RES_74k_1.P.n103 RES_74k_1.P.t39 8.84311
R11832 RES_74k_1.P.n106 RES_74k_1.P.t37 8.83779
R11833 RES_74k_1.P.n105 RES_74k_1.P.n104 8.83029
R11834 RES_74k_1.P.n100 RES_74k_1.P.n99 8.83029
R11835 RES_74k_1.P.n98 RES_74k_1.P.t35 8.79474
R11836 RES_74k_1.P.n101 RES_74k_1.P.t32 8.76273
R11837 RES_74k_1.P.n112 RES_74k_1.P.n111 8.5505
R11838 RES_74k_1.P.n110 RES_74k_1.P.t75 8.5505
R11839 RES_74k_1.P.n113 RES_74k_1.P.t77 8.03277
R11840 RES_74k_1.P.n116 RES_74k_1.P.n115 6.73062
R11841 RES_74k_1.P.n20 RES_74k_1.P.t24 6.45834
R11842 RES_74k_1.P.n92 RES_74k_1.P.t82 6.1905
R11843 RES_74k_1.P.n46 RES_74k_1.P.t81 6.1905
R11844 RES_74k_1.P.n45 RES_74k_1.P.t9 6.1905
R11845 RES_74k_1.P.n44 RES_74k_1.P.t8 6.1905
R11846 RES_74k_1.P.n43 RES_74k_1.P.t45 6.1905
R11847 RES_74k_1.P.n42 RES_74k_1.P.t44 6.1905
R11848 RES_74k_1.P.n41 RES_74k_1.P.t102 6.1905
R11849 RES_74k_1.P.n40 RES_74k_1.P.t101 6.1905
R11850 RES_74k_1.P.n39 RES_74k_1.P.t5 6.1905
R11851 RES_74k_1.P.n38 RES_74k_1.P.t4 6.1905
R11852 RES_74k_1.P.n36 RES_74k_1.P.t69 6.1905
R11853 RES_74k_1.P.n20 RES_74k_1.P.t41 6.1905
R11854 RES_74k_1.P.n21 RES_74k_1.P.t3 6.1905
R11855 RES_74k_1.P.n22 RES_74k_1.P.t51 6.1905
R11856 RES_74k_1.P.n23 RES_74k_1.P.t67 6.1905
R11857 RES_74k_1.P.n24 RES_74k_1.P.t80 6.1905
R11858 RES_74k_1.P.n25 RES_74k_1.P.t108 6.1905
R11859 RES_74k_1.P.n26 RES_74k_1.P.t23 6.1905
R11860 RES_74k_1.P.n27 RES_74k_1.P.t57 6.1905
R11861 RES_74k_1.P.n28 RES_74k_1.P.t19 6.1905
R11862 RES_74k_1.P.n29 RES_74k_1.P.t88 6.1905
R11863 RES_74k_1.P.n30 RES_74k_1.P.t49 6.1905
R11864 RES_74k_1.P.n31 RES_74k_1.P.t1 6.1905
R11865 RES_74k_1.P.n32 RES_74k_1.P.t92 6.1905
R11866 RES_74k_1.P.n33 RES_74k_1.P.t43 6.1905
R11867 RES_74k_1.P.n34 RES_74k_1.P.t100 6.1905
R11868 RES_74k_1.P.n35 RES_74k_1.P.t53 6.1905
R11869 RES_74k_1.P.n66 RES_74k_1.P.t25 6.1905
R11870 RES_74k_1.P.n67 RES_74k_1.P.t46 6.1905
R11871 RES_74k_1.P.n68 RES_74k_1.P.t47 6.1905
R11872 RES_74k_1.P.n69 RES_74k_1.P.t97 6.1905
R11873 RES_74k_1.P.n70 RES_74k_1.P.t98 6.1905
R11874 RES_74k_1.P.n71 RES_74k_1.P.t64 6.1905
R11875 RES_74k_1.P.n72 RES_74k_1.P.t65 6.1905
R11876 RES_74k_1.P.n73 RES_74k_1.P.t89 6.1905
R11877 RES_74k_1.P.n64 RES_74k_1.P.t90 6.1905
R11878 RES_74k_1.P.n63 RES_74k_1.P.t84 6.1905
R11879 RES_74k_1.P.n62 RES_74k_1.P.t61 6.1905
R11880 RES_74k_1.P.n61 RES_74k_1.P.t13 6.1905
R11881 RES_74k_1.P.n60 RES_74k_1.P.t71 6.1905
R11882 RES_74k_1.P.n59 RES_74k_1.P.t86 6.1905
R11883 RES_74k_1.P.n58 RES_74k_1.P.t94 6.1905
R11884 RES_74k_1.P.n57 RES_74k_1.P.t21 6.1905
R11885 RES_74k_1.P.n56 RES_74k_1.P.t74 6.1905
R11886 RES_74k_1.P.n55 RES_74k_1.P.t55 6.1905
R11887 RES_74k_1.P.n54 RES_74k_1.P.t31 6.1905
R11888 RES_74k_1.P.n53 RES_74k_1.P.t17 6.1905
R11889 RES_74k_1.P.n52 RES_74k_1.P.t7 6.1905
R11890 RES_74k_1.P.n51 RES_74k_1.P.t63 6.1905
R11891 RES_74k_1.P.n50 RES_74k_1.P.t11 6.1905
R11892 RES_74k_1.P.n49 RES_74k_1.P.t29 6.1905
R11893 RES_74k_1.P.n48 RES_74k_1.P.t15 6.1905
R11894 RES_74k_1.P.n47 RES_74k_1.P.t96 6.1905
R11895 RES_74k_1.P.n89 RES_74k_1.P.t83 6.1905
R11896 RES_74k_1.P.n65 RES_74k_1.P.t95 6.1905
R11897 RES_74k_1.P.n74 RES_74k_1.P.t14 6.1905
R11898 RES_74k_1.P.n75 RES_74k_1.P.t28 6.1905
R11899 RES_74k_1.P.n76 RES_74k_1.P.t10 6.1905
R11900 RES_74k_1.P.n77 RES_74k_1.P.t62 6.1905
R11901 RES_74k_1.P.n78 RES_74k_1.P.t6 6.1905
R11902 RES_74k_1.P.n79 RES_74k_1.P.t16 6.1905
R11903 RES_74k_1.P.n80 RES_74k_1.P.t30 6.1905
R11904 RES_74k_1.P.n81 RES_74k_1.P.t54 6.1905
R11905 RES_74k_1.P.n82 RES_74k_1.P.t73 6.1905
R11906 RES_74k_1.P.n83 RES_74k_1.P.t20 6.1905
R11907 RES_74k_1.P.n84 RES_74k_1.P.t93 6.1905
R11908 RES_74k_1.P.n85 RES_74k_1.P.t85 6.1905
R11909 RES_74k_1.P.n86 RES_74k_1.P.t70 6.1905
R11910 RES_74k_1.P.n87 RES_74k_1.P.t12 6.1905
R11911 RES_74k_1.P.n88 RES_74k_1.P.t60 6.1905
R11912 RES_74k_1.P.n3 RES_74k_1.P.t40 6.1905
R11913 RES_74k_1.P.n4 RES_74k_1.P.t2 6.1905
R11914 RES_74k_1.P.n5 RES_74k_1.P.t50 6.1905
R11915 RES_74k_1.P.n6 RES_74k_1.P.t66 6.1905
R11916 RES_74k_1.P.n7 RES_74k_1.P.t79 6.1905
R11917 RES_74k_1.P.n8 RES_74k_1.P.t107 6.1905
R11918 RES_74k_1.P.n9 RES_74k_1.P.t22 6.1905
R11919 RES_74k_1.P.n10 RES_74k_1.P.t56 6.1905
R11920 RES_74k_1.P.n11 RES_74k_1.P.t18 6.1905
R11921 RES_74k_1.P.n12 RES_74k_1.P.t87 6.1905
R11922 RES_74k_1.P.n13 RES_74k_1.P.t48 6.1905
R11923 RES_74k_1.P.n14 RES_74k_1.P.t0 6.1905
R11924 RES_74k_1.P.n15 RES_74k_1.P.t91 6.1905
R11925 RES_74k_1.P.n16 RES_74k_1.P.t42 6.1905
R11926 RES_74k_1.P.n17 RES_74k_1.P.t99 6.1905
R11927 RES_74k_1.P.n18 RES_74k_1.P.t52 6.1905
R11928 RES_74k_1.P.n19 RES_74k_1.P.t68 6.1905
R11929 RES_74k_1.P.n135 RES_74k_1.P.t105 5.81586
R11930 RES_74k_1.P.n143 RES_74k_1.P.n140 5.10148
R11931 RES_74k_1.P.n139 RES_74k_1.P.n138 5.10115
R11932 RES_74k_1.P.n137 RES_74k_1.P.n136 5.08021
R11933 RES_74k_1.P.n143 RES_74k_1.P.n142 4.66166
R11934 RES_74k_1.P.n93 RES_74k_1.P.t72 3.49604
R11935 RES_74k_1.P.n130 RES_74k_1.P.n129 3.47886
R11936 RES_74k_1.P.n135 RES_74k_1.P.n134 2.85093
R11937 RES_74k_1.P.n94 RES_74k_1.P.n93 2.52714
R11938 RES_74k_1.P.n119 RES_74k_1.P.t109 2.38861
R11939 RES_74k_1.P.n120 RES_74k_1.P.t112 2.38861
R11940 RES_74k_1.P.n0 RES_74k_1.P.t110 2.38861
R11941 RES_74k_1.P.n114 RES_74k_1.P 2.35224
R11942 RES_74k_1.P RES_74k_1.P.n94 2.3422
R11943 RES_74k_1.P.n0 RES_74k_1.P.n122 2.29444
R11944 RES_74k_1.P.n0 RES_74k_1.P.n121 2.29444
R11945 RES_74k_1.P.n291 RES_74k_1.P.n289 2.29119
R11946 RES_74k_1.P.n310 RES_74k_1.P.n150 2.29119
R11947 RES_74k_1.P.n148 RES_74k_1.P.n299 2.28464
R11948 RES_74k_1.P.n118 RES_74k_1.P.n117 2.25183
R11949 RES_74k_1.P.n131 RES_74k_1.P.n130 2.25092
R11950 RES_74k_1.P.n242 RES_74k_1.P.n286 2.2505
R11951 RES_74k_1.P.n241 RES_74k_1.P.n240 2.2505
R11952 RES_74k_1.P.n239 RES_74k_1.P.n238 2.2505
R11953 RES_74k_1.P.n237 RES_74k_1.P.n236 2.2505
R11954 RES_74k_1.P.n234 RES_74k_1.P.n235 2.2505
R11955 RES_74k_1.P.n229 RES_74k_1.P.n230 2.2505
R11956 RES_74k_1.P.n119 RES_74k_1.P.t114 2.2505
R11957 RES_74k_1.P.n120 RES_74k_1.P.t113 2.2505
R11958 RES_74k_1.P.n0 RES_74k_1.P.t111 2.2505
R11959 RES_74k_1.P.n147 RES_74k_1.P.n191 2.2505
R11960 RES_74k_1.P.n146 RES_74k_1.P.n199 2.2505
R11961 RES_74k_1.P.n129 RES_74k_1.P.n128 2.2505
R11962 RES_74k_1.P.n96 RES_74k_1.P.n95 2.2505
R11963 RES_74k_1.P.n134 RES_74k_1.P.t106 2.16717
R11964 RES_74k_1.P.n134 RES_74k_1.P.n133 2.16717
R11965 RES_74k_1.P.n142 RES_74k_1.P.t26 1.9505
R11966 RES_74k_1.P.n142 RES_74k_1.P.n141 1.9505
R11967 RES_74k_1.P.n107 RES_74k_1.P.n106 1.92684
R11968 RES_74k_1.P.n132 RES_74k_1.P.n131 1.90259
R11969 RES_74k_1.P RES_74k_1.P.n132 1.70729
R11970 RES_74k_1.P.n108 RES_74k_1.P.n107 1.50147
R11971 RES_74k_1.P.n188 RES_74k_1.P.n186 1.5005
R11972 RES_74k_1.P.n196 RES_74k_1.P.n194 1.5005
R11973 RES_74k_1.P.n296 RES_74k_1.P.n297 1.5005
R11974 RES_74k_1.P.n152 RES_74k_1.P.n157 1.5005
R11975 RES_74k_1.P.n114 RES_74k_1.P.n113 1.40626
R11976 RES_74k_1.P.n90 RES_74k_1.P.n63 1.2155
R11977 RES_74k_1.P.n37 RES_74k_1.P.n19 1.2155
R11978 RES_74k_1.P.n64 RES_74k_1.P.n73 1.20532
R11979 RES_74k_1.P.n72 RES_74k_1.P.n71 1.20532
R11980 RES_74k_1.P.n70 RES_74k_1.P.n69 1.20532
R11981 RES_74k_1.P.n68 RES_74k_1.P.n67 1.20532
R11982 RES_74k_1.P.n39 RES_74k_1.P.n38 1.20532
R11983 RES_74k_1.P.n41 RES_74k_1.P.n40 1.20532
R11984 RES_74k_1.P.n43 RES_74k_1.P.n42 1.20532
R11985 RES_74k_1.P.n45 RES_74k_1.P.n44 1.20532
R11986 RES_74k_1.P.n91 RES_74k_1.P.n46 1.19574
R11987 RES_74k_1.P.n223 RES_74k_1.P.n218 1.15852
R11988 RES_74k_1.P.n286 RES_74k_1.P.n163 1.1255
R11989 RES_74k_1.P.n243 RES_74k_1.P.n206 1.1255
R11990 RES_74k_1.P.n235 RES_74k_1.P.n171 1.1255
R11991 RES_74k_1.P.n307 RES_74k_1.P.n159 1.1255
R11992 RES_74k_1.P.n202 RES_74k_1.P.n203 1.1255
R11993 RES_74k_1.P.n126 RES_74k_1.P.n124 1.1255
R11994 RES_74k_1.P.n145 RES_74k_1.P.n180 1.1255
R11995 RES_74k_1.P.n176 RES_74k_1.P.n177 1.1255
R11996 RES_74k_1.P.n171 RES_74k_1.P.n172 1.1255
R11997 RES_74k_1.P.n165 RES_74k_1.P.n166 1.1255
R11998 RES_74k_1.P.n163 RES_74k_1.P.n164 1.1255
R11999 RES_74k_1.P.n191 RES_74k_1.P.n189 1.12277
R12000 RES_74k_1.P.n199 RES_74k_1.P.n197 1.12277
R12001 RES_74k_1.P.n299 RES_74k_1.P.n300 1.12277
R12002 RES_74k_1.P.n150 RES_74k_1.P.n149 1.12277
R12003 RES_74k_1.P.n112 RES_74k_1.P.n110 1.1179
R12004 RES_74k_1.P.n291 RES_74k_1.P.n219 1.09572
R12005 RES_74k_1.P.n132 RES_74k_1.P 1.06348
R12006 RES_74k_1.P.n310 RES_74k_1.P.n242 0.963384
R12007 RES_74k_1.P.n232 RES_74k_1.P.n229 0.888704
R12008 RES_74k_1.P.n115 RES_74k_1.P.n108 0.859311
R12009 RES_74k_1.P.n128 RES_74k_1.P.n127 0.750314
R12010 RES_74k_1.P.n117 RES_74k_1.P.n123 0.677022
R12011 RES_74k_1.P.n148 RES_74k_1.P.n146 0.660845
R12012 RES_74k_1.P.n137 RES_74k_1.P.n135 0.644196
R12013 RES_74k_1.P.n63 RES_74k_1.P.n62 0.587457
R12014 RES_74k_1.P.n62 RES_74k_1.P.n61 0.587457
R12015 RES_74k_1.P.n61 RES_74k_1.P.n60 0.587457
R12016 RES_74k_1.P.n60 RES_74k_1.P.n59 0.587457
R12017 RES_74k_1.P.n59 RES_74k_1.P.n58 0.587457
R12018 RES_74k_1.P.n58 RES_74k_1.P.n57 0.587457
R12019 RES_74k_1.P.n57 RES_74k_1.P.n56 0.587457
R12020 RES_74k_1.P.n56 RES_74k_1.P.n55 0.587457
R12021 RES_74k_1.P.n55 RES_74k_1.P.n54 0.587457
R12022 RES_74k_1.P.n54 RES_74k_1.P.n53 0.587457
R12023 RES_74k_1.P.n53 RES_74k_1.P.n52 0.587457
R12024 RES_74k_1.P.n52 RES_74k_1.P.n51 0.587457
R12025 RES_74k_1.P.n51 RES_74k_1.P.n50 0.587457
R12026 RES_74k_1.P.n50 RES_74k_1.P.n49 0.587457
R12027 RES_74k_1.P.n49 RES_74k_1.P.n48 0.587457
R12028 RES_74k_1.P.n48 RES_74k_1.P.n47 0.587457
R12029 RES_74k_1.P.n89 RES_74k_1.P.n88 0.587457
R12030 RES_74k_1.P.n88 RES_74k_1.P.n87 0.587457
R12031 RES_74k_1.P.n87 RES_74k_1.P.n86 0.587457
R12032 RES_74k_1.P.n86 RES_74k_1.P.n85 0.587457
R12033 RES_74k_1.P.n85 RES_74k_1.P.n84 0.587457
R12034 RES_74k_1.P.n84 RES_74k_1.P.n83 0.587457
R12035 RES_74k_1.P.n83 RES_74k_1.P.n82 0.587457
R12036 RES_74k_1.P.n82 RES_74k_1.P.n81 0.587457
R12037 RES_74k_1.P.n81 RES_74k_1.P.n80 0.587457
R12038 RES_74k_1.P.n80 RES_74k_1.P.n79 0.587457
R12039 RES_74k_1.P.n79 RES_74k_1.P.n78 0.587457
R12040 RES_74k_1.P.n78 RES_74k_1.P.n77 0.587457
R12041 RES_74k_1.P.n77 RES_74k_1.P.n76 0.587457
R12042 RES_74k_1.P.n76 RES_74k_1.P.n75 0.587457
R12043 RES_74k_1.P.n75 RES_74k_1.P.n74 0.587457
R12044 RES_74k_1.P.n74 RES_74k_1.P.n65 0.587457
R12045 RES_74k_1.P.n19 RES_74k_1.P.n18 0.587457
R12046 RES_74k_1.P.n18 RES_74k_1.P.n17 0.587457
R12047 RES_74k_1.P.n17 RES_74k_1.P.n16 0.587457
R12048 RES_74k_1.P.n16 RES_74k_1.P.n15 0.587457
R12049 RES_74k_1.P.n15 RES_74k_1.P.n14 0.587457
R12050 RES_74k_1.P.n14 RES_74k_1.P.n13 0.587457
R12051 RES_74k_1.P.n13 RES_74k_1.P.n12 0.587457
R12052 RES_74k_1.P.n12 RES_74k_1.P.n11 0.587457
R12053 RES_74k_1.P.n11 RES_74k_1.P.n10 0.587457
R12054 RES_74k_1.P.n10 RES_74k_1.P.n9 0.587457
R12055 RES_74k_1.P.n9 RES_74k_1.P.n8 0.587457
R12056 RES_74k_1.P.n8 RES_74k_1.P.n7 0.587457
R12057 RES_74k_1.P.n7 RES_74k_1.P.n6 0.587457
R12058 RES_74k_1.P.n6 RES_74k_1.P.n5 0.587457
R12059 RES_74k_1.P.n5 RES_74k_1.P.n4 0.587457
R12060 RES_74k_1.P.n4 RES_74k_1.P.n3 0.587457
R12061 RES_74k_1.P.n36 RES_74k_1.P.n35 0.587457
R12062 RES_74k_1.P.n35 RES_74k_1.P.n34 0.587457
R12063 RES_74k_1.P.n34 RES_74k_1.P.n33 0.587457
R12064 RES_74k_1.P.n33 RES_74k_1.P.n32 0.587457
R12065 RES_74k_1.P.n32 RES_74k_1.P.n31 0.587457
R12066 RES_74k_1.P.n31 RES_74k_1.P.n30 0.587457
R12067 RES_74k_1.P.n30 RES_74k_1.P.n29 0.587457
R12068 RES_74k_1.P.n29 RES_74k_1.P.n28 0.587457
R12069 RES_74k_1.P.n28 RES_74k_1.P.n27 0.587457
R12070 RES_74k_1.P.n27 RES_74k_1.P.n26 0.587457
R12071 RES_74k_1.P.n26 RES_74k_1.P.n25 0.587457
R12072 RES_74k_1.P.n25 RES_74k_1.P.n24 0.587457
R12073 RES_74k_1.P.n24 RES_74k_1.P.n23 0.587457
R12074 RES_74k_1.P.n23 RES_74k_1.P.n22 0.587457
R12075 RES_74k_1.P.n22 RES_74k_1.P.n21 0.587457
R12076 RES_74k_1.P.n21 RES_74k_1.P.n20 0.587457
R12077 RES_74k_1.P.n100 RES_74k_1.P.n98 0.576883
R12078 RES_74k_1.P.n101 RES_74k_1.P.n100 0.571972
R12079 RES_74k_1.P.n106 RES_74k_1.P.n105 0.550283
R12080 RES_74k_1.P.n105 RES_74k_1.P.n103 0.544413
R12081 RES_74k_1.P.n93 RES_74k_1.P.n92 0.54333
R12082 RES_74k_1.P.n129 RES_74k_1.P.n147 0.472288
R12083 RES_74k_1.P.n113 RES_74k_1.P.n112 0.454295
R12084 RES_74k_1.P.n139 RES_74k_1.P.n137 0.45084
R12085 RES_74k_1.P.n115 RES_74k_1.P.n114 0.321541
R12086 RES_74k_1.P.n144 RES_74k_1.P.n143 0.309585
R12087 RES_74k_1.P.n144 RES_74k_1.P.n139 0.274999
R12088 RES_74k_1.P.n73 RES_74k_1.P.n72 0.274015
R12089 RES_74k_1.P.n71 RES_74k_1.P.n70 0.274015
R12090 RES_74k_1.P.n69 RES_74k_1.P.n68 0.274015
R12091 RES_74k_1.P.n67 RES_74k_1.P.n66 0.274015
R12092 RES_74k_1.P.n40 RES_74k_1.P.n39 0.274015
R12093 RES_74k_1.P.n42 RES_74k_1.P.n41 0.274015
R12094 RES_74k_1.P.n44 RES_74k_1.P.n43 0.274015
R12095 RES_74k_1.P.n46 RES_74k_1.P.n45 0.274015
R12096 RES_74k_1.P.n65 RES_74k_1.P.n64 0.268344
R12097 RES_74k_1.P.n38 RES_74k_1.P.n37 0.264431
R12098 RES_74k_1.P.n91 RES_74k_1.P.n90 0.254848
R12099 RES_74k_1.P.n96 RES_74k_1.P.n94 0.140594
R12100 RES_74k_1.P.n107 RES_74k_1.P.n101 0.112274
R12101 RES_74k_1.P RES_74k_1.P.n108 0.11163
R12102 RES_74k_1.P.n123 RES_74k_1.P.n120 0.0995566
R12103 RES_74k_1.P RES_74k_1.P.n144 0.0936034
R12104 RES_74k_1.P.n117 RES_74k_1.P.n119 0.0692209
R12105 RES_74k_1.P.n118 RES_74k_1.P.n307 0.0665262
R12106 RES_74k_1.P.n95 RES_74k_1.P 0.0488962
R12107 RES_74k_1.P.n116 RES_74k_1.P.n96 0.0412547
R12108 RES_74k_1.P.n213 RES_74k_1.P.n228 0.0366935
R12109 RES_74k_1.P.n186 RES_74k_1.P.n185 0.032
R12110 RES_74k_1.P.n194 RES_74k_1.P.n193 0.032
R12111 RES_74k_1.P.n297 RES_74k_1.P.n298 0.032
R12112 RES_74k_1.P.n157 RES_74k_1.P.n156 0.032
R12113 RES_74k_1.P.n234 RES_74k_1.P 0.0315619
R12114 RES_74k_1.P.n90 RES_74k_1.P.n89 0.0298478
R12115 RES_74k_1.P.n37 RES_74k_1.P.n36 0.0298478
R12116 RES_74k_1.P.n92 RES_74k_1.P.n91 0.0298478
R12117 RES_74k_1.P.n183 RES_74k_1.P.n190 0.0257
R12118 RES_74k_1.P.n175 RES_74k_1.P.n198 0.0257
R12119 RES_74k_1.P.n292 RES_74k_1.P.n301 0.0257
R12120 RES_74k_1.P.n154 RES_74k_1.P.n153 0.0257
R12121 RES_74k_1.P.n216 RES_74k_1.P.n225 0.0256613
R12122 RES_74k_1.P.n277 RES_74k_1.P.n279 0.0241947
R12123 RES_74k_1.P.n268 RES_74k_1.P.n244 0.0224027
R12124 RES_74k_1.P.n214 RES_74k_1.P.n224 0.0219839
R12125 RES_74k_1.P.n249 RES_74k_1.P.n257 0.0216062
R12126 RES_74k_1.P.n204 RES_74k_1.P.n205 0.0210088
R12127 RES_74k_1.P.n261 RES_74k_1.P.n253 0.0198142
R12128 RES_74k_1.P.n200 RES_74k_1.P.n179 0.0184204
R12129 RES_74k_1.P.n184 RES_74k_1.P.n182 0.0175923
R12130 RES_74k_1.P.n192 RES_74k_1.P.n174 0.0175923
R12131 RES_74k_1.P.n293 RES_74k_1.P.n294 0.0175923
R12132 RES_74k_1.P.n155 RES_74k_1.P.n158 0.0175923
R12133 RES_74k_1.P.n147 RES_74k_1.P.n148 0.0108448
R12134 RES_74k_1.P.n189 RES_74k_1.P.n188 0.00836872
R12135 RES_74k_1.P.n197 RES_74k_1.P.n196 0.00836872
R12136 RES_74k_1.P.n300 RES_74k_1.P.n296 0.00836872
R12137 RES_74k_1.P.n149 RES_74k_1.P.n152 0.00836872
R12138 RES_74k_1.P.n168 RES_74k_1.P.n252 0.00667257
R12139 RES_74k_1.P.n272 RES_74k_1.P.n237 0.00607522
R12140 RES_74k_1.P.n273 RES_74k_1.P.n176 0.00607522
R12141 RES_74k_1.P.n239 RES_74k_1.P.n255 0.00587611
R12142 RES_74k_1.P.n165 RES_74k_1.P.n256 0.00587611
R12143 RES_74k_1.P.n146 RES_74k_1.P.n310 0.00567241
R12144 RES_74k_1.P.n229 RES_74k_1.P.n291 0.00563308
R12145 RES_74k_1.P.n124 RES_74k_1.P.n125 0.00558246
R12146 RES_74k_1.P.n211 RES_74k_1.P.n222 0.00495161
R12147 RES_74k_1.P.n215 RES_74k_1.P.n208 0.00475806
R12148 RES_74k_1.P.n212 RES_74k_1.P.n226 0.00475806
R12149 RES_74k_1.P.n220 RES_74k_1.P.n227 0.00456452
R12150 RES_74k_1.P.n181 RES_74k_1.P.n306 0.00443013
R12151 RES_74k_1.P.n209 RES_74k_1.P.n217 0.00437097
R12152 RES_74k_1.P.n275 RES_74k_1.P.n249 0.00428319
R12153 RES_74k_1.P.n170 RES_74k_1.P.n284 0.00428319
R12154 RES_74k_1.P.n242 RES_74k_1.P.n234 0.00428319
R12155 RES_74k_1.P.n210 RES_74k_1.P.n221 0.00417742
R12156 RES_74k_1.P.n266 RES_74k_1.P.n241 0.00368584
R12157 RES_74k_1.P.n201 RES_74k_1.P.n285 0.00368584
R12158 RES_74k_1.P.n267 RES_74k_1.P.n243 0.00368584
R12159 RES_74k_1.P.n145 RES_74k_1.P.n309 0.0036441
R12160 RES_74k_1.P.n233 RES_74k_1.P.n281 0.00348673
R12161 RES_74k_1.P.n161 RES_74k_1.P.n262 0.00348673
R12162 RES_74k_1.P.n202 RES_74k_1.P.n282 0.00348673
R12163 RES_74k_1.P.n247 RES_74k_1.P.n274 0.00348673
R12164 RES_74k_1.P.n164 RES_74k_1.P.n248 0.00328761
R12165 RES_74k_1.P.n287 RES_74k_1.P.n250 0.00328761
R12166 RES_74k_1.P.n127 RES_74k_1.P.n126 0.00327501
R12167 RES_74k_1.P.n241 RES_74k_1.P.n233 0.0030885
R12168 RES_74k_1.P.n279 RES_74k_1.P.n266 0.0030885
R12169 RES_74k_1.P.n173 RES_74k_1.P.n288 0.0030885
R12170 RES_74k_1.P.n243 RES_74k_1.P.n202 0.0030885
R12171 RES_74k_1.P.n240 RES_74k_1.P.n232 0.0030885
R12172 RES_74k_1.P.n307 RES_74k_1.P.n145 0.00285808
R12173 RES_74k_1.P.n286 RES_74k_1.P.n259 0.00249115
R12174 RES_74k_1.P.n245 RES_74k_1.P.n169 0.00249115
R12175 RES_74k_1.P.n163 RES_74k_1.P.n260 0.00249115
R12176 RES_74k_1.P.n235 RES_74k_1.P.n275 0.00229204
R12177 RES_74k_1.P.n207 RES_74k_1.P.n246 0.00229204
R12178 RES_74k_1.P.n280 RES_74k_1.P.n263 0.00229204
R12179 RES_74k_1.P.n171 RES_74k_1.P.n276 0.00229204
R12180 RES_74k_1.P.n217 RES_74k_1.P.n214 0.00224194
R12181 RES_74k_1.P.n283 RES_74k_1.P.n265 0.00209292
R12182 RES_74k_1.P.n302 RES_74k_1.P.n304 0.00207205
R12183 RES_74k_1.P RES_74k_1.P.n236 0.00189381
R12184 RES_74k_1.P.n305 RES_74k_1.P.n308 0.00187555
R12185 RES_74k_1.P.n218 RES_74k_1.P.n210 0.00187097
R12186 RES_74k_1.P.n218 RES_74k_1.P.n209 0.00187029
R12187 RES_74k_1.P.n219 RES_74k_1.P.n213 0.00185484
R12188 RES_74k_1.P.n225 RES_74k_1.P.n220 0.00185484
R12189 RES_74k_1.P.n227 RES_74k_1.P.n212 0.00185484
R12190 RES_74k_1.P.n228 RES_74k_1.P.n223 0.00166129
R12191 RES_74k_1.P.n224 RES_74k_1.P.n215 0.00166129
R12192 RES_74k_1.P.n208 RES_74k_1.P.n211 0.00166129
R12193 RES_74k_1.P.n222 RES_74k_1.P.n216 0.00166129
R12194 RES_74k_1.P.n282 RES_74k_1.P.n283 0.00149557
R12195 RES_74k_1.P.n250 RES_74k_1.P.n261 0.00149557
R12196 RES_74k_1.P.n276 RES_74k_1.P.n287 0.00149557
R12197 RES_74k_1.P.n309 RES_74k_1.P.n305 0.00148253
R12198 RES_74k_1.P.n191 RES_74k_1.P.n187 0.0014
R12199 RES_74k_1.P.n188 RES_74k_1.P.n183 0.0014
R12200 RES_74k_1.P.n186 RES_74k_1.P.n184 0.0014
R12201 RES_74k_1.P.n199 RES_74k_1.P.n195 0.0014
R12202 RES_74k_1.P.n196 RES_74k_1.P.n175 0.0014
R12203 RES_74k_1.P.n194 RES_74k_1.P.n192 0.0014
R12204 RES_74k_1.P.n230 RES_74k_1.P.n231 0.0014
R12205 RES_74k_1.P.n289 RES_74k_1.P.n290 0.0014
R12206 RES_74k_1.P.n299 RES_74k_1.P.n295 0.0014
R12207 RES_74k_1.P.n296 RES_74k_1.P.n292 0.0014
R12208 RES_74k_1.P.n297 RES_74k_1.P.n293 0.0014
R12209 RES_74k_1.P.n157 RES_74k_1.P.n155 0.0014
R12210 RES_74k_1.P.n152 RES_74k_1.P.n154 0.0014
R12211 RES_74k_1.P.n150 RES_74k_1.P.n151 0.0014
R12212 RES_74k_1.P.n284 RES_74k_1.P.n207 0.00129646
R12213 RES_74k_1.P.n262 RES_74k_1.P.n200 0.00129646
R12214 RES_74k_1.P.n288 RES_74k_1.P.n161 0.00129646
R12215 RES_74k_1.P.n263 RES_74k_1.P.n267 0.00129646
R12216 RES_74k_1.P.n244 RES_74k_1.P.n280 0.00129646
R12217 RES_74k_1.P.n278 RES_74k_1.P.n251 0.00129646
R12218 RES_74k_1.P.n260 RES_74k_1.P.n247 0.00129646
R12219 RES_74k_1.P.n306 RES_74k_1.P.n302 0.00128603
R12220 RES_74k_1.P.n169 RES_74k_1.P.n264 0.00109734
R12221 RES_74k_1.P.n205 RES_74k_1.P.n245 0.00109734
R12222 RES_74k_1.P.n269 RES_74k_1.P.n178 0.00109734
R12223 RES_74k_1.P.n248 RES_74k_1.P.n201 0.00109734
R12224 RES_74k_1.P.n270 RES_74k_1.P.n258 0.00109734
R12225 RES_74k_1.P.n167 RES_74k_1.P.n254 0.00089823
R12226 RES_74k_1.P.n131 RES_74k_1.P.n116 0.000852941
R12227 RES_74k_1.P.n255 RES_74k_1.P.n277 0.000699115
R12228 RES_74k_1.P.n237 RES_74k_1.P.n239 0.000699115
R12229 RES_74k_1.P.n257 RES_74k_1.P.n272 0.000699115
R12230 RES_74k_1.P.n203 RES_74k_1.P.n170 0.000699115
R12231 RES_74k_1.P.n206 RES_74k_1.P.n160 0.000699115
R12232 RES_74k_1.P.n178 RES_74k_1.P.n204 0.000699115
R12233 RES_74k_1.P.n252 RES_74k_1.P.n269 0.000699115
R12234 RES_74k_1.P.n166 RES_74k_1.P.n168 0.000699115
R12235 RES_74k_1.P.n254 RES_74k_1.P.n271 0.000699115
R12236 RES_74k_1.P.n179 RES_74k_1.P.n167 0.000699115
R12237 RES_74k_1.P.n172 RES_74k_1.P.n173 0.000699115
R12238 RES_74k_1.P.n164 RES_74k_1.P.n162 0.000699115
R12239 RES_74k_1.P.n251 RES_74k_1.P.n268 0.000699115
R12240 RES_74k_1.P.n256 RES_74k_1.P.n278 0.000699115
R12241 RES_74k_1.P.n176 RES_74k_1.P.n165 0.000699115
R12242 RES_74k_1.P.n258 RES_74k_1.P.n273 0.000699115
R12243 RES_74k_1.P.n253 RES_74k_1.P.n270 0.000699115
R12244 RES_74k_1.P.n126 RES_74k_1.P.n118 0.000696507
R12245 RES_74k_1.P.n180 RES_74k_1.P.n181 0.000696507
R12246 RES_74k_1.P.n159 RES_74k_1.P.n303 0.000696507
R12247 RES_74k_1.P.n0 RES_74k_1.P.n1 2.63208
R12248 RES_74k_1.P.n0 RES_74k_1.P.n2 2.63208
R12249 RES_74k_1.P.n123 RES_74k_1.P.n0 0.741958
R12250 A_MUX_0.Tr_Gate_1.CLK.n2 A_MUX_0.Tr_Gate_1.CLK.t21 45.6363
R12251 A_MUX_0.Tr_Gate_1.CLK.n4 A_MUX_0.Tr_Gate_1.CLK.t13 29.6446
R12252 A_MUX_0.Tr_Gate_1.CLK.t17 A_MUX_0.Tr_Gate_1.CLK.n5 29.6446
R12253 A_MUX_0.Tr_Gate_1.CLK.n6 A_MUX_0.Tr_Gate_1.CLK.t15 24.6117
R12254 A_MUX_0.Tr_Gate_1.CLK.n5 A_MUX_0.Tr_Gate_1.CLK.n4 22.2047
R12255 A_MUX_0.Tr_Gate_1.CLK.t21 A_MUX_0.Tr_Gate_1.CLK.t16 22.1925
R12256 A_MUX_0.Tr_Gate_1.CLK.n3 A_MUX_0.Tr_Gate_1.CLK.n2 20.9314
R12257 A_MUX_0.Tr_Gate_1.CLK A_MUX_0.Tr_Gate_1.CLK.t17 18.5231
R12258 A_MUX_0.Tr_Gate_1.CLK.n6 A_MUX_0.Tr_Gate_1.CLK.t18 6.1325
R12259 A_MUX_0.Tr_Gate_1.CLK.n4 A_MUX_0.Tr_Gate_1.CLK.t19 6.1325
R12260 A_MUX_0.Tr_Gate_1.CLK.n5 A_MUX_0.Tr_Gate_1.CLK.t14 6.1325
R12261 A_MUX_0.Tr_Gate_1.CLK.n2 A_MUX_0.Tr_Gate_1.CLK.t20 6.1325
R12262 A_MUX_0.Tr_Gate_1.CLK.n3 A_MUX_0.Tr_Gate_1.CLK.t12 6.1325
R12263 A_MUX_0.Tr_Gate_1.CLK A_MUX_0.Tr_Gate_1.CLK.n3 5.28481
R12264 A_MUX_0.Tr_Gate_1.CLK A_MUX_0.Tr_Gate_1.CLK.n6 4.89628
R12265 A_MUX_0.Tr_Gate_1.CLK.n18 A_MUX_0.Tr_Gate_1.CLK.t1 3.6405
R12266 A_MUX_0.Tr_Gate_1.CLK.n18 A_MUX_0.Tr_Gate_1.CLK.n17 3.6405
R12267 A_MUX_0.Tr_Gate_1.CLK.n10 A_MUX_0.Tr_Gate_1.CLK.t4 3.6405
R12268 A_MUX_0.Tr_Gate_1.CLK.n10 A_MUX_0.Tr_Gate_1.CLK.n9 3.6405
R12269 A_MUX_0.Tr_Gate_1.CLK.n8 A_MUX_0.Tr_Gate_1.CLK.t3 3.6405
R12270 A_MUX_0.Tr_Gate_1.CLK.n8 A_MUX_0.Tr_Gate_1.CLK.n7 3.6405
R12271 A_MUX_0.Tr_Gate_1.CLK.n16 A_MUX_0.Tr_Gate_1.CLK.t0 3.6405
R12272 A_MUX_0.Tr_Gate_1.CLK.n16 A_MUX_0.Tr_Gate_1.CLK.n15 3.6405
R12273 A_MUX_0.Tr_Gate_1.CLK.n0 A_MUX_0.Tr_Gate_1.CLK.n14 3.50463
R12274 A_MUX_0.Tr_Gate_1.CLK.n1 A_MUX_0.Tr_Gate_1.CLK.n12 3.50463
R12275 A_MUX_0.Tr_Gate_1.CLK.n14 A_MUX_0.Tr_Gate_1.CLK.t2 3.2765
R12276 A_MUX_0.Tr_Gate_1.CLK.n14 A_MUX_0.Tr_Gate_1.CLK.n13 3.2765
R12277 A_MUX_0.Tr_Gate_1.CLK.n12 A_MUX_0.Tr_Gate_1.CLK.t5 3.2765
R12278 A_MUX_0.Tr_Gate_1.CLK.n12 A_MUX_0.Tr_Gate_1.CLK.n11 3.2765
R12279 A_MUX_0.Tr_Gate_1.CLK.n1 A_MUX_0.Tr_Gate_1.CLK.n8 3.06224
R12280 A_MUX_0.Tr_Gate_1.CLK.n0 A_MUX_0.Tr_Gate_1.CLK.n16 3.06224
R12281 A_MUX_0.Tr_Gate_1.CLK.n1 A_MUX_0.Tr_Gate_1.CLK.n10 2.6005
R12282 A_MUX_0.Tr_Gate_1.CLK.n0 A_MUX_0.Tr_Gate_1.CLK.n18 2.6005
R12283 A_MUX_0.Tr_Gate_1.CLK.n1 A_MUX_0.Tr_Gate_1.CLK 1.62988
R12284 A_MUX_0.Tr_Gate_1.CLK.n1 A_MUX_0.Tr_Gate_1.CLK.n0 0.98463
R12285 VCO_DFF_C_0.VCTRL.n4 VCO_DFF_C_0.VCTRL.t20 27.5268
R12286 VCO_DFF_C_0.VCTRL.n17 VCO_DFF_C_0.VCTRL.t17 27.5268
R12287 VCO_DFF_C_0.VCTRL.n19 VCO_DFF_C_0.VCTRL.t24 25.3421
R12288 VCO_DFF_C_0.VCTRL.n7 VCO_DFF_C_0.VCTRL.t32 25.3421
R12289 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCTRL.n16 9.02002
R12290 VCO_DFF_C_0.VCTRL.n21 VCO_DFF_C_0.VCTRL.t34 8.86359
R12291 VCO_DFF_C_0.VCTRL.n9 VCO_DFF_C_0.VCTRL.t21 8.86319
R12292 VCO_DFF_C_0.VCTRL.n30 VCO_DFF_C_0.VCTRL 8.47187
R12293 VCO_DFF_C_0.VCTRL.n11 VCO_DFF_C_0.VCTRL.t31 7.92693
R12294 VCO_DFF_C_0.VCTRL.n24 VCO_DFF_C_0.VCTRL.t28 7.92677
R12295 VCO_DFF_C_0.VCTRL.n8 VCO_DFF_C_0.VCTRL.t16 7.79605
R12296 VCO_DFF_C_0.VCTRL.n22 VCO_DFF_C_0.VCTRL.t19 7.79604
R12297 VCO_DFF_C_0.VCTRL.n5 VCO_DFF_C_0.VCTRL.t30 7.57548
R12298 VCO_DFF_C_0.VCTRL.n18 VCO_DFF_C_0.VCTRL.t26 7.54055
R12299 VCO_DFF_C_0.VCTRL.n6 VCO_DFF_C_0.VCTRL.t27 7.49426
R12300 VCO_DFF_C_0.VCTRL.n23 VCO_DFF_C_0.VCTRL.t29 7.49403
R12301 VCO_DFF_C_0.VCTRL.n0 VCO_DFF_C_0.VCTRL.t3 6.74387
R12302 VCO_DFF_C_0.VCTRL.n1 VCO_DFF_C_0.VCTRL.n48 6.74326
R12303 VCO_DFF_C_0.VCTRL.n12 VCO_DFF_C_0.VCTRL.t23 6.73304
R12304 VCO_DFF_C_0.VCTRL.n25 VCO_DFF_C_0.VCTRL.t18 6.73175
R12305 VCO_DFF_C_0.VCTRL.n1 VCO_DFF_C_0.VCTRL.n49 5.1005
R12306 VCO_DFF_C_0.VCTRL.n0 VCO_DFF_C_0.VCTRL.t0 5.1005
R12307 VCO_DFF_C_0.VCTRL.n5 VCO_DFF_C_0.VCTRL.n4 4.72106
R12308 VCO_DFF_C_0.VCTRL.n18 VCO_DFF_C_0.VCTRL.n17 4.72106
R12309 VCO_DFF_C_0.VCTRL.n10 VCO_DFF_C_0.VCTRL.n7 3.90288
R12310 VCO_DFF_C_0.VCTRL.n20 VCO_DFF_C_0.VCTRL.n19 3.90053
R12311 VCO_DFF_C_0.VCTRL.n46 VCO_DFF_C_0.VCTRL.n43 3.57508
R12312 VCO_DFF_C_0.VCTRL.n34 VCO_DFF_C_0.VCTRL.n37 3.56654
R12313 VCO_DFF_C_0.VCTRL.n1 VCO_DFF_C_0.VCTRL.t9 3.40075
R12314 VCO_DFF_C_0.VCTRL.n0 VCO_DFF_C_0.VCTRL.n38 3.40011
R12315 VCO_DFF_C_0.VCTRL.n39 VCO_DFF_C_0.VCTRL.t2 3.00158
R12316 VCO_DFF_C_0.VCTRL.n50 VCO_DFF_C_0.VCTRL.n47 3.00032
R12317 VCO_DFF_C_0.VCTRL.n15 VCO_DFF_C_0.VCTRL 2.50091
R12318 VCO_DFF_C_0.VCTRL.n28 VCO_DFF_C_0.VCTRL 2.46425
R12319 VCO_DFF_C_0.VCTRL.n35 VCO_DFF_C_0.VCTRL.n33 2.41287
R12320 VCO_DFF_C_0.VCTRL.n52 VCO_DFF_C_0.VCTRL.n41 2.36206
R12321 VCO_DFF_C_0.VCTRL.n16 VCO_DFF_C_0.VCTRL 2.32969
R12322 VCO_DFF_C_0.VCTRL.n41 VCO_DFF_C_0.VCTRL.n40 2.30849
R12323 VCO_DFF_C_0.VCTRL.n3 VCO_DFF_C_0.VCTRL.n35 2.26352
R12324 VCO_DFF_C_0.VCTRL.n19 VCO_DFF_C_0.VCTRL.t22 2.17312
R12325 VCO_DFF_C_0.VCTRL.n4 VCO_DFF_C_0.VCTRL.t35 2.17312
R12326 VCO_DFF_C_0.VCTRL.n7 VCO_DFF_C_0.VCTRL.t25 2.17312
R12327 VCO_DFF_C_0.VCTRL.n17 VCO_DFF_C_0.VCTRL.t33 2.17312
R12328 VCO_DFF_C_0.VCTRL.n37 VCO_DFF_C_0.VCTRL.t13 2.16717
R12329 VCO_DFF_C_0.VCTRL.n37 VCO_DFF_C_0.VCTRL.n36 2.16717
R12330 VCO_DFF_C_0.VCTRL.n33 VCO_DFF_C_0.VCTRL.t12 2.16717
R12331 VCO_DFF_C_0.VCTRL.n33 VCO_DFF_C_0.VCTRL.n32 2.16717
R12332 VCO_DFF_C_0.VCTRL.n45 VCO_DFF_C_0.VCTRL.t4 2.16717
R12333 VCO_DFF_C_0.VCTRL.n45 VCO_DFF_C_0.VCTRL.n44 2.16717
R12334 VCO_DFF_C_0.VCTRL.n43 VCO_DFF_C_0.VCTRL.t7 2.16717
R12335 VCO_DFF_C_0.VCTRL.n43 VCO_DFF_C_0.VCTRL.n42 2.16717
R12336 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCTRL.n28 1.89901
R12337 VCO_DFF_C_0.VCTRL.n26 VCO_DFF_C_0.VCTRL.n25 1.896
R12338 VCO_DFF_C_0.VCTRL.n13 VCO_DFF_C_0.VCTRL.n12 1.89145
R12339 VCO_DFF_C_0.VCTRL.n51 VCO_DFF_C_0.VCTRL.n50 1.84797
R12340 VCO_DFF_C_0.VCTRL.n3 VCO_DFF_C_0.VCTRL.n39 1.82978
R12341 VCO_DFF_C_0.VCTRL.n27 VCO_DFF_C_0.VCTRL.n26 1.5395
R12342 VCO_DFF_C_0.VCTRL.n14 VCO_DFF_C_0.VCTRL.n13 1.5395
R12343 VCO_DFF_C_0.VCTRL.n29 VCO_DFF_C_0.VCTRL 1.4706
R12344 VCO_DFF_C_0.VCTRL.n2 VCO_DFF_C_0.VCTRL 0.663665
R12345 VCO_DFF_C_0.VCTRL.n2 VCO_DFF_C_0.VCTRL.n31 1.25555
R12346 VCO_DFF_C_0.VCTRL.n46 VCO_DFF_C_0.VCTRL.n45 1.25233
R12347 VCO_DFF_C_0.VCTRL.n51 VCO_DFF_C_0.VCTRL.n46 1.12574
R12348 VCO_DFF_C_0.VCTRL.n11 VCO_DFF_C_0.VCTRL.n10 1.05913
R12349 VCO_DFF_C_0.VCTRL.n13 VCO_DFF_C_0.VCTRL.n6 0.957464
R12350 VCO_DFF_C_0.VCTRL.n26 VCO_DFF_C_0.VCTRL.n23 0.95722
R12351 VCO_DFF_C_0.VCTRL.n16 VCO_DFF_C_0.VCTRL.n15 0.798473
R12352 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCTRL.n52 0.751569
R12353 VCO_DFF_C_0.VCTRL.n9 VCO_DFF_C_0.VCTRL.n8 0.749817
R12354 VCO_DFF_C_0.VCTRL.n22 VCO_DFF_C_0.VCTRL.n21 0.749568
R12355 VCO_DFF_C_0.VCTRL.n40 VCO_DFF_C_0.VCTRL 0.736653
R12356 VCO_DFF_C_0.VCTRL.n23 VCO_DFF_C_0.VCTRL.n22 0.622921
R12357 VCO_DFF_C_0.VCTRL.n8 VCO_DFF_C_0.VCTRL.n6 0.622675
R12358 VCO_DFF_C_0.VCTRL.n21 VCO_DFF_C_0.VCTRL.n20 0.602194
R12359 VCO_DFF_C_0.VCTRL.n10 VCO_DFF_C_0.VCTRL.n9 0.602194
R12360 VCO_DFF_C_0.VCTRL.n50 VCO_DFF_C_0.VCTRL.n1 0.558374
R12361 VCO_DFF_C_0.VCTRL.n39 VCO_DFF_C_0.VCTRL.n0 0.558372
R12362 VCO_DFF_C_0.VCTRL.n29 VCO_DFF_C_0.VCTRL 0.550625
R12363 VCO_DFF_C_0.VCTRL.n12 VCO_DFF_C_0.VCTRL.n11 0.453053
R12364 VCO_DFF_C_0.VCTRL.n25 VCO_DFF_C_0.VCTRL.n24 0.451515
R12365 VCO_DFF_C_0.VCTRL.n15 VCO_DFF_C_0.VCTRL.n14 0.43025
R12366 VCO_DFF_C_0.VCTRL.n28 VCO_DFF_C_0.VCTRL.n27 0.43025
R12367 VCO_DFF_C_0.VCTRL.n40 VCO_DFF_C_0.VCTRL.n3 0.394824
R12368 VCO_DFF_C_0.VCTRL.n52 VCO_DFF_C_0.VCTRL.n51 0.33941
R12369 VCO_DFF_C_0.VCTRL.n14 VCO_DFF_C_0.VCTRL.n5 0.266
R12370 VCO_DFF_C_0.VCTRL.n27 VCO_DFF_C_0.VCTRL.n18 0.266
R12371 VCO_DFF_C_0.VCTRL.n41 VCO_DFF_C_0.VCTRL.n2 0.25987
R12372 VCO_DFF_C_0.VCTRL.n31 VCO_DFF_C_0.VCTRL.n30 0.23889
R12373 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCTRL.n29 0.195324
R12374 VCO_DFF_C_0.VCTRL.n35 VCO_DFF_C_0.VCTRL.n34 0.145661
R12375 a_22967_8787.n0 a_22967_8787.t14 33.8126
R12376 a_22967_8787.n1 a_22967_8787.n0 30.3299
R12377 a_22967_8787.n2 a_22967_8787.n1 30.3299
R12378 a_22967_8787.n3 a_22967_8787.n2 30.3299
R12379 a_22967_8787.n4 a_22967_8787.n3 30.3299
R12380 a_22967_8787.n5 a_22967_8787.n4 30.3299
R12381 a_22967_8787.n6 a_22967_8787.n5 30.3299
R12382 a_22967_8787.n7 a_22967_8787.n6 30.3299
R12383 a_22967_8787.n8 a_22967_8787.n7 30.3299
R12384 a_22967_8787.n12 a_22967_8787.t7 26.2202
R12385 a_22967_8787.n9 a_22967_8787.t6 12.8368
R12386 a_22967_8787.n9 a_22967_8787.n8 12.0257
R12387 a_22967_8787.n13 a_22967_8787.n12 8.40022
R12388 a_22967_8787.n14 a_22967_8787.n9 5.21471
R12389 a_22967_8787.n12 a_22967_8787.t15 3.6505
R12390 a_22967_8787.n0 a_22967_8787.t4 3.6505
R12391 a_22967_8787.n1 a_22967_8787.t11 3.6505
R12392 a_22967_8787.n2 a_22967_8787.t5 3.6505
R12393 a_22967_8787.n3 a_22967_8787.t12 3.6505
R12394 a_22967_8787.n4 a_22967_8787.t9 3.6505
R12395 a_22967_8787.n5 a_22967_8787.t16 3.6505
R12396 a_22967_8787.n6 a_22967_8787.t10 3.6505
R12397 a_22967_8787.n7 a_22967_8787.t13 3.6505
R12398 a_22967_8787.n8 a_22967_8787.t8 3.6505
R12399 a_22967_8787.n15 a_22967_8787.t3 3.6405
R12400 a_22967_8787.n16 a_22967_8787.n15 3.6405
R12401 a_22967_8787.n14 a_22967_8787.n13 3.38778
R12402 a_22967_8787.n11 a_22967_8787.t1 3.38774
R12403 a_22967_8787.n11 a_22967_8787.n10 2.97656
R12404 a_22967_8787.n13 a_22967_8787.n11 2.47435
R12405 a_22967_8787.n15 a_22967_8787.n14 1.25578
R12406 a_21443_8068.n5 a_21443_8068.n4 5.71637
R12407 a_21443_8068.n6 a_21443_8068.t2 4.95333
R12408 a_21443_8068.n7 a_21443_8068.n1 3.54746
R12409 a_21443_8068.n5 a_21443_8068.n3 2.6005
R12410 a_21443_8068.n8 a_21443_8068.n7 2.6005
R12411 a_21443_8068.n1 a_21443_8068.t4 1.6255
R12412 a_21443_8068.n1 a_21443_8068.n0 1.6255
R12413 a_21443_8068.n3 a_21443_8068.t6 1.6255
R12414 a_21443_8068.n3 a_21443_8068.n2 1.6255
R12415 a_21443_8068.n8 a_21443_8068.t5 1.6255
R12416 a_21443_8068.n9 a_21443_8068.n8 1.6255
R12417 a_21443_8068.n6 a_21443_8068.n5 0.728326
R12418 a_21443_8068.n7 a_21443_8068.n6 0.552239
R12419 VCO_DFF_C_0.VCO_C_0.OUTB.n20 VCO_DFF_C_0.VCO_C_0.OUTB.t47 45.6363
R12420 VCO_DFF_C_0.VCO_C_0.OUTB.n26 VCO_DFF_C_0.VCO_C_0.OUTB.t35 45.6363
R12421 VCO_DFF_C_0.VCO_C_0.OUTB.n23 VCO_DFF_C_0.VCO_C_0.OUTB.t48 29.6446
R12422 VCO_DFF_C_0.VCO_C_0.OUTB.t51 VCO_DFF_C_0.VCO_C_0.OUTB.n24 29.6446
R12423 VCO_DFF_C_0.VCO_C_0.OUTB.n29 VCO_DFF_C_0.VCO_C_0.OUTB.t43 29.6446
R12424 VCO_DFF_C_0.VCO_C_0.OUTB.t41 VCO_DFF_C_0.VCO_C_0.OUTB.n30 29.6446
R12425 VCO_DFF_C_0.VCO_C_0.OUTB.n19 VCO_DFF_C_0.VCO_C_0.OUTB.t33 24.6117
R12426 VCO_DFF_C_0.VCO_C_0.OUTB.n28 VCO_DFF_C_0.VCO_C_0.OUTB.t32 24.6117
R12427 VCO_DFF_C_0.VCO_C_0.OUTB.n40 VCO_DFF_C_0.VCO_C_0.OUTB.t28 23.6945
R12428 VCO_DFF_C_0.VCO_C_0.OUTB.t16 VCO_DFF_C_0.VCO_C_0.OUTB.n41 23.6945
R12429 VCO_DFF_C_0.VCO_C_0.OUTB.n24 VCO_DFF_C_0.VCO_C_0.OUTB.n23 22.2047
R12430 VCO_DFF_C_0.VCO_C_0.OUTB.n30 VCO_DFF_C_0.VCO_C_0.OUTB.n29 22.2047
R12431 VCO_DFF_C_0.VCO_C_0.OUTB.t47 VCO_DFF_C_0.VCO_C_0.OUTB.t15 22.1925
R12432 VCO_DFF_C_0.VCO_C_0.OUTB.t35 VCO_DFF_C_0.VCO_C_0.OUTB.t46 22.1925
R12433 VCO_DFF_C_0.VCO_C_0.OUTB.n21 VCO_DFF_C_0.VCO_C_0.OUTB.n20 20.9314
R12434 VCO_DFF_C_0.VCO_C_0.OUTB.n27 VCO_DFF_C_0.VCO_C_0.OUTB.n26 20.9314
R12435 VCO_DFF_C_0.VCO_C_0.OUTB.n41 VCO_DFF_C_0.VCO_C_0.OUTB.n40 18.8035
R12436 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.OUTB.t41 18.5191
R12437 VCO_DFF_C_0.VCO_C_0.OUTB.n25 VCO_DFF_C_0.VCO_C_0.OUTB.t51 17.9055
R12438 VCO_DFF_C_0.VCO_C_0.OUTB.n38 VCO_DFF_C_0.VCO_C_0.OUTB.n36 15.8172
R12439 VCO_DFF_C_0.VCO_C_0.OUTB.n38 VCO_DFF_C_0.VCO_C_0.OUTB.n37 15.8172
R12440 VCO_DFF_C_0.VCO_C_0.OUTB.n37 VCO_DFF_C_0.VCO_C_0.OUTB.n33 15.8172
R12441 VCO_DFF_C_0.VCO_C_0.OUTB.n46 VCO_DFF_C_0.VCO_C_0.OUTB.t14 15.4917
R12442 VCO_DFF_C_0.VCO_C_0.OUTB.n48 VCO_DFF_C_0.VCO_C_0.OUTB.t18 15.3942
R12443 VCO_DFF_C_0.VCO_C_0.OUTB.n49 VCO_DFF_C_0.VCO_C_0.OUTB.t38 14.9265
R12444 VCO_DFF_C_0.VCO_C_0.OUTB.n36 VCO_DFF_C_0.VCO_C_0.OUTB.t52 14.8925
R12445 VCO_DFF_C_0.VCO_C_0.OUTB.t27 VCO_DFF_C_0.VCO_C_0.OUTB.n38 14.8925
R12446 VCO_DFF_C_0.VCO_C_0.OUTB.n37 VCO_DFF_C_0.VCO_C_0.OUTB.t17 14.8925
R12447 VCO_DFF_C_0.VCO_C_0.OUTB.n53 VCO_DFF_C_0.VCO_C_0.OUTB.t31 14.7749
R12448 VCO_DFF_C_0.VCO_C_0.OUTB.n47 VCO_DFF_C_0.VCO_C_0.OUTB.t50 13.6019
R12449 VCO_DFF_C_0.VCO_C_0.OUTB.n53 VCO_DFF_C_0.VCO_C_0.OUTB.t23 13.5312
R12450 VCO_DFF_C_0.VCO_C_0.OUTB.n51 VCO_DFF_C_0.VCO_C_0.OUTB.t42 13.4877
R12451 VCO_DFF_C_0.VCO_C_0.OUTB.n49 VCO_DFF_C_0.VCO_C_0.OUTB.t30 13.227
R12452 VCO_DFF_C_0.VCO_C_0.OUTB.n50 VCO_DFF_C_0.VCO_C_0.OUTB.t26 13.1835
R12453 VCO_DFF_C_0.VCO_C_0.OUTB.n42 VCO_DFF_C_0.VCO_C_0.OUTB.n34 12.2457
R12454 VCO_DFF_C_0.VCO_C_0.OUTB.n39 VCO_DFF_C_0.VCO_C_0.OUTB.n34 12.2457
R12455 VCO_DFF_C_0.VCO_C_0.OUTB.n39 VCO_DFF_C_0.VCO_C_0.OUTB.n35 12.2457
R12456 VCO_DFF_C_0.VCO_C_0.OUTB.n43 VCO_DFF_C_0.VCO_C_0.OUTB.t36 11.6285
R12457 VCO_DFF_C_0.VCO_C_0.OUTB.n45 VCO_DFF_C_0.VCO_C_0.OUTB.n2 9.0064
R12458 VCO_DFF_C_0.VCO_C_0.OUTB.n35 VCO_DFF_C_0.VCO_C_0.OUTB.t28 8.9065
R12459 VCO_DFF_C_0.VCO_C_0.OUTB.t49 VCO_DFF_C_0.VCO_C_0.OUTB.n39 8.9065
R12460 VCO_DFF_C_0.VCO_C_0.OUTB.t37 VCO_DFF_C_0.VCO_C_0.OUTB.n34 8.9065
R12461 VCO_DFF_C_0.VCO_C_0.OUTB.n42 VCO_DFF_C_0.VCO_C_0.OUTB.t16 8.9065
R12462 VCO_DFF_C_0.VCO_C_0.OUTB.n38 VCO_DFF_C_0.VCO_C_0.OUTB.t24 8.6145
R12463 VCO_DFF_C_0.VCO_C_0.OUTB.n36 VCO_DFF_C_0.VCO_C_0.OUTB.t45 8.6145
R12464 VCO_DFF_C_0.VCO_C_0.OUTB.n37 VCO_DFF_C_0.VCO_C_0.OUTB.t13 8.6145
R12465 VCO_DFF_C_0.VCO_C_0.OUTB.n33 VCO_DFF_C_0.VCO_C_0.OUTB.t34 8.59715
R12466 VCO_DFF_C_0.VCO_C_0.OUTB.t52 VCO_DFF_C_0.VCO_C_0.OUTB.n35 8.3225
R12467 VCO_DFF_C_0.VCO_C_0.OUTB.n39 VCO_DFF_C_0.VCO_C_0.OUTB.t27 8.3225
R12468 VCO_DFF_C_0.VCO_C_0.OUTB.t17 VCO_DFF_C_0.VCO_C_0.OUTB.n34 8.3225
R12469 VCO_DFF_C_0.VCO_C_0.OUTB.t36 VCO_DFF_C_0.VCO_C_0.OUTB.n42 8.3225
R12470 VCO_DFF_C_0.VCO_C_0.OUTB.n2 VCO_DFF_C_0.VCO_C_0.OUTB.n25 8.24338
R12471 VCO_DFF_C_0.VCO_C_0.OUTB.n46 VCO_DFF_C_0.VCO_C_0.OUTB.t53 8.1387
R12472 VCO_DFF_C_0.VCO_C_0.OUTB.n23 VCO_DFF_C_0.VCO_C_0.OUTB.t40 6.1325
R12473 VCO_DFF_C_0.VCO_C_0.OUTB.n24 VCO_DFF_C_0.VCO_C_0.OUTB.t44 6.1325
R12474 VCO_DFF_C_0.VCO_C_0.OUTB.n19 VCO_DFF_C_0.VCO_C_0.OUTB.t22 6.1325
R12475 VCO_DFF_C_0.VCO_C_0.OUTB.n20 VCO_DFF_C_0.VCO_C_0.OUTB.t21 6.1325
R12476 VCO_DFF_C_0.VCO_C_0.OUTB.n21 VCO_DFF_C_0.VCO_C_0.OUTB.t12 6.1325
R12477 VCO_DFF_C_0.VCO_C_0.OUTB.n28 VCO_DFF_C_0.VCO_C_0.OUTB.t39 6.1325
R12478 VCO_DFF_C_0.VCO_C_0.OUTB.n29 VCO_DFF_C_0.VCO_C_0.OUTB.t25 6.1325
R12479 VCO_DFF_C_0.VCO_C_0.OUTB.n30 VCO_DFF_C_0.VCO_C_0.OUTB.t19 6.1325
R12480 VCO_DFF_C_0.VCO_C_0.OUTB.n26 VCO_DFF_C_0.VCO_C_0.OUTB.t20 6.1325
R12481 VCO_DFF_C_0.VCO_C_0.OUTB.n27 VCO_DFF_C_0.VCO_C_0.OUTB.t29 6.1325
R12482 VCO_DFF_C_0.VCO_C_0.OUTB.n32 VCO_DFF_C_0.VCO_C_0.OUTB.n27 5.5044
R12483 VCO_DFF_C_0.VCO_C_0.OUTB.n22 VCO_DFF_C_0.VCO_C_0.OUTB.n21 5.38991
R12484 VCO_DFF_C_0.VCO_C_0.OUTB.n22 VCO_DFF_C_0.VCO_C_0.OUTB.n19 4.83094
R12485 VCO_DFF_C_0.VCO_C_0.OUTB.n31 VCO_DFF_C_0.VCO_C_0.OUTB.n28 4.83094
R12486 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.OUTB.n43 4.223
R12487 VCO_DFF_C_0.VCO_C_0.OUTB.n40 VCO_DFF_C_0.VCO_C_0.OUTB.t49 3.6505
R12488 VCO_DFF_C_0.VCO_C_0.OUTB.n41 VCO_DFF_C_0.VCO_C_0.OUTB.t37 3.6505
R12489 VCO_DFF_C_0.VCO_C_0.OUTB.n14 VCO_DFF_C_0.VCO_C_0.OUTB.t8 3.6405
R12490 VCO_DFF_C_0.VCO_C_0.OUTB.n14 VCO_DFF_C_0.VCO_C_0.OUTB.n13 3.6405
R12491 VCO_DFF_C_0.VCO_C_0.OUTB.n8 VCO_DFF_C_0.VCO_C_0.OUTB.t10 3.6405
R12492 VCO_DFF_C_0.VCO_C_0.OUTB.n8 VCO_DFF_C_0.VCO_C_0.OUTB.n7 3.6405
R12493 VCO_DFF_C_0.VCO_C_0.OUTB.n10 VCO_DFF_C_0.VCO_C_0.OUTB.t6 3.6405
R12494 VCO_DFF_C_0.VCO_C_0.OUTB.n10 VCO_DFF_C_0.VCO_C_0.OUTB.n9 3.6405
R12495 VCO_DFF_C_0.VCO_C_0.OUTB.n16 VCO_DFF_C_0.VCO_C_0.OUTB.t5 3.6405
R12496 VCO_DFF_C_0.VCO_C_0.OUTB.n16 VCO_DFF_C_0.VCO_C_0.OUTB.n15 3.6405
R12497 VCO_DFF_C_0.VCO_C_0.OUTB.n18 VCO_DFF_C_0.VCO_C_0.OUTB.n4 3.50463
R12498 VCO_DFF_C_0.VCO_C_0.OUTB.n12 VCO_DFF_C_0.VCO_C_0.OUTB.n6 3.50463
R12499 VCO_DFF_C_0.VCO_C_0.OUTB.n4 VCO_DFF_C_0.VCO_C_0.OUTB.t1 3.2765
R12500 VCO_DFF_C_0.VCO_C_0.OUTB.n4 VCO_DFF_C_0.VCO_C_0.OUTB.n3 3.2765
R12501 VCO_DFF_C_0.VCO_C_0.OUTB.n6 VCO_DFF_C_0.VCO_C_0.OUTB.t3 3.2765
R12502 VCO_DFF_C_0.VCO_C_0.OUTB.n6 VCO_DFF_C_0.VCO_C_0.OUTB.n5 3.2765
R12503 VCO_DFF_C_0.VCO_C_0.OUTB.n43 VCO_DFF_C_0.VCO_C_0.OUTB.n33 3.1807
R12504 VCO_DFF_C_0.VCO_C_0.OUTB.n11 VCO_DFF_C_0.VCO_C_0.OUTB.n10 3.06224
R12505 VCO_DFF_C_0.VCO_C_0.OUTB.n17 VCO_DFF_C_0.VCO_C_0.OUTB.n14 3.06224
R12506 VCO_DFF_C_0.VCO_C_0.OUTB.n2 VCO_DFF_C_0.VCO_C_0.OUTB.n44 2.82705
R12507 VCO_DFF_C_0.VCO_C_0.OUTB.n11 VCO_DFF_C_0.VCO_C_0.OUTB.n8 2.6005
R12508 VCO_DFF_C_0.VCO_C_0.OUTB.n17 VCO_DFF_C_0.VCO_C_0.OUTB.n16 2.6005
R12509 VCO_DFF_C_0.VCO_C_0.OUTB.n2 VCO_DFF_C_0.VCO_C_0.OUTB 2.36547
R12510 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.OUTB.n56 2.30807
R12511 VCO_DFF_C_0.VCO_C_0.OUTB.n0 VCO_DFF_C_0.VCO_C_0.OUTB.n1 1.10603
R12512 VCO_DFF_C_0.VCO_C_0.OUTB.n56 VCO_DFF_C_0.VCO_C_0.OUTB.n55 2.2505
R12513 VCO_DFF_C_0.VCO_C_0.OUTB.n52 VCO_DFF_C_0.VCO_C_0.OUTB.n48 1.5982
R12514 VCO_DFF_C_0.VCO_C_0.OUTB.n54 VCO_DFF_C_0.VCO_C_0.OUTB.n52 1.18336
R12515 VCO_DFF_C_0.VCO_C_0.OUTB.n55 VCO_DFF_C_0.VCO_C_0.OUTB.n54 0.977746
R12516 VCO_DFF_C_0.VCO_C_0.OUTB.n18 VCO_DFF_C_0.VCO_C_0.OUTB.n12 0.798761
R12517 VCO_DFF_C_0.VCO_C_0.OUTB.n45 VCO_DFF_C_0.VCO_C_0.OUTB.n0 0.66931
R12518 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.OUTB.n22 0.658318
R12519 VCO_DFF_C_0.VCO_C_0.OUTB.n31 VCO_DFF_C_0.VCO_C_0.OUTB 0.637045
R12520 VCO_DFF_C_0.VCO_C_0.OUTB.n25 VCO_DFF_C_0.VCO_C_0.OUTB 0.6125
R12521 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.OUTB.n18 0.562022
R12522 VCO_DFF_C_0.VCO_C_0.OUTB.n32 VCO_DFF_C_0.VCO_C_0.OUTB.n31 0.458758
R12523 VCO_DFF_C_0.VCO_C_0.OUTB.n47 VCO_DFF_C_0.VCO_C_0.OUTB.n46 0.381495
R12524 VCO_DFF_C_0.VCO_C_0.OUTB.n54 VCO_DFF_C_0.VCO_C_0.OUTB.n53 0.37501
R12525 VCO_DFF_C_0.VCO_C_0.OUTB.n48 VCO_DFF_C_0.VCO_C_0.OUTB.n47 0.355126
R12526 VCO_DFF_C_0.VCO_C_0.OUTB.n51 VCO_DFF_C_0.VCO_C_0.OUTB.n50 0.31227
R12527 VCO_DFF_C_0.VCO_C_0.OUTB.n50 VCO_DFF_C_0.VCO_C_0.OUTB.n49 0.298874
R12528 VCO_DFF_C_0.VCO_C_0.OUTB.n56 VCO_DFF_C_0.VCO_C_0.OUTB.n0 0.281082
R12529 VCO_DFF_C_0.VCO_C_0.OUTB.n44 VCO_DFF_C_0.VCO_C_0.OUTB.n32 0.238532
R12530 VCO_DFF_C_0.VCO_C_0.OUTB.n52 VCO_DFF_C_0.VCO_C_0.OUTB.n51 0.233052
R12531 VCO_DFF_C_0.VCO_C_0.OUTB.n12 VCO_DFF_C_0.VCO_C_0.OUTB.n11 0.18637
R12532 VCO_DFF_C_0.VCO_C_0.OUTB.n18 VCO_DFF_C_0.VCO_C_0.OUTB.n17 0.18637
R12533 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.OUTB.n1 0.203752
R12534 VCO_DFF_C_0.VCO_C_0.OUTB.n55 VCO_DFF_C_0.VCO_C_0.OUTB.n45 0.137564
R12535 VCO_DFF_C_0.VCO_C_0.OUTB.n44 VCO_DFF_C_0.VCO_C_0.OUTB 0.104622
R12536 VCO_DFF_C_0.VCO_C_0.OUTB.n1 VCO_DFF_C_0.VCO_C_0.OUTB 0.147946
R12537 S6.t5 S6.t9 144.929
R12538 S6.t2 S6.t11 44.058
R12539 S6.n1 S6.t12 25.9486
R12540 S6.t12 S6 16.1689
R12541 S6.n4 S6.n3 15.8172
R12542 S6.n5 S6.n4 15.8172
R12543 S6.n0 S6.t5 14.796
R12544 S6.n6 S6.t1 14.4701
R12545 S6.n0 S6.t2 13.8835
R12546 S6.n2 S6.n1 13.2388
R12547 S6.n2 S6.t3 12.7103
R12548 S6.n3 S6.t7 11.7326
R12549 S6.n3 S6.t4 11.7326
R12550 S6.n4 S6.t8 11.7326
R12551 S6.n4 S6.t6 11.7326
R12552 S6.n5 S6.t10 11.7326
R12553 S6.t1 S6.n5 11.7326
R12554 S6 S6.n0 9.83788
R12555 S6.n1 S6.t0 7.3005
R12556 S6 S6.n6 4.18916
R12557 S6.n6 S6.n2 1.49961
R12558 mux_magic_3.AND2_magic_0.A.t9 mux_magic_3.AND2_magic_0.A.t11 144.929
R12559 mux_magic_3.AND2_magic_0.A.t12 mux_magic_3.AND2_magic_0.A.t10 44.058
R12560 mux_magic_3.AND2_magic_0.A.n0 mux_magic_3.AND2_magic_0.A.t9 14.796
R12561 mux_magic_3.AND2_magic_0.A.n0 mux_magic_3.AND2_magic_0.A.t12 13.8835
R12562 mux_magic_3.AND2_magic_0.A mux_magic_3.AND2_magic_0.A.n0 9.83788
R12563 mux_magic_3.AND2_magic_0.A.n11 mux_magic_3.AND2_magic_0.A.n2 4.99061
R12564 mux_magic_3.AND2_magic_0.A.n14 mux_magic_3.AND2_magic_0.A.n1 4.5405
R12565 mux_magic_3.AND2_magic_0.A.n13 mux_magic_3.AND2_magic_0.A.n12 4.2255
R12566 mux_magic_3.AND2_magic_0.A.n10 mux_magic_3.AND2_magic_0.A.n4 3.52811
R12567 mux_magic_3.AND2_magic_0.A.n9 mux_magic_3.AND2_magic_0.A.n6 3.30485
R12568 mux_magic_3.AND2_magic_0.A.n9 mux_magic_3.AND2_magic_0.A.n8 2.6005
R12569 mux_magic_3.AND2_magic_0.A.n6 mux_magic_3.AND2_magic_0.A.t6 1.6255
R12570 mux_magic_3.AND2_magic_0.A.n6 mux_magic_3.AND2_magic_0.A.n5 1.6255
R12571 mux_magic_3.AND2_magic_0.A.n8 mux_magic_3.AND2_magic_0.A.t4 1.6255
R12572 mux_magic_3.AND2_magic_0.A.n8 mux_magic_3.AND2_magic_0.A.n7 1.6255
R12573 mux_magic_3.AND2_magic_0.A.n4 mux_magic_3.AND2_magic_0.A.t2 1.463
R12574 mux_magic_3.AND2_magic_0.A.n4 mux_magic_3.AND2_magic_0.A.n3 1.463
R12575 mux_magic_3.AND2_magic_0.A.n11 mux_magic_3.AND2_magic_0.A.n10 0.8105
R12576 mux_magic_3.AND2_magic_0.A.n13 mux_magic_3.AND2_magic_0.A.n11 0.389848
R12577 mux_magic_3.AND2_magic_0.A.n10 mux_magic_3.AND2_magic_0.A.n9 0.389848
R12578 mux_magic_3.AND2_magic_0.A.n14 mux_magic_3.AND2_magic_0.A.n13 0.256804
R12579 mux_magic_3.AND2_magic_0.A mux_magic_3.AND2_magic_0.A.n14 0.173882
R12580 mux_magic_1.OR_magic_0.B.t7 mux_magic_1.OR_magic_0.B.t3 44.6331
R12581 mux_magic_1.OR_magic_0.B.t5 mux_magic_1.OR_magic_0.B.t7 43.4094
R12582 mux_magic_1.OR_magic_0.B.t4 mux_magic_1.OR_magic_0.B.t5 31.5469
R12583 mux_magic_1.OR_magic_0.B.n0 mux_magic_1.OR_magic_0.B.t4 15.0567
R12584 mux_magic_1.OR_magic_0.B.n0 mux_magic_1.OR_magic_0.B.t6 13.6228
R12585 mux_magic_1.OR_magic_0.B mux_magic_1.OR_magic_0.B.n1 5.03757
R12586 mux_magic_1.OR_magic_0.B mux_magic_1.OR_magic_0.B.n0 4.2675
R12587 mux_magic_1.OR_magic_0.B mux_magic_1.OR_magic_0.B.n3 3.36521
R12588 mux_magic_1.OR_magic_0.B.n3 mux_magic_1.OR_magic_0.B.t1 1.6255
R12589 mux_magic_1.OR_magic_0.B.n3 mux_magic_1.OR_magic_0.B.n2 1.6255
R12590 a_29415_9553.t6 a_29415_9553.t7 31.5469
R12591 a_29415_9553.n2 a_29415_9553.t6 13.227
R12592 a_29415_9553.n2 a_29415_9553.t8 13.138
R12593 a_29415_9553.n0 a_29415_9553.t5 6.53038
R12594 a_29415_9553.n0 a_29415_9553.n2 4.33404
R12595 a_29415_9553.n4 a_29415_9553.n3 4.2255
R12596 a_29415_9553.n6 a_29415_9553.n5 4.2255
R12597 a_29415_9553.n8 a_29415_9553.n6 3.81956
R12598 a_29415_9553.n0 a_29415_9553.n1 2.62675
R12599 a_29415_9553.t0 a_29415_9553.n8 1.6255
R12600 a_29415_9553.n8 a_29415_9553.n7 1.6255
R12601 a_29415_9553.n6 a_29415_9553.n4 0.947457
R12602 a_29415_9553.n4 a_29415_9553.n0 0.600587
R12603 a_29415_8145.n9 a_29415_8145.n8 5.71637
R12604 a_29415_8145.n5 a_29415_8145.t4 4.95333
R12605 a_29415_8145.n4 a_29415_8145.n1 3.54746
R12606 a_29415_8145.n4 a_29415_8145.n3 2.6005
R12607 a_29415_8145.n8 a_29415_8145.n7 2.6005
R12608 a_29415_8145.n7 a_29415_8145.t0 1.6255
R12609 a_29415_8145.n7 a_29415_8145.n6 1.6255
R12610 a_29415_8145.n1 a_29415_8145.t2 1.6255
R12611 a_29415_8145.n1 a_29415_8145.n0 1.6255
R12612 a_29415_8145.n3 a_29415_8145.t1 1.6255
R12613 a_29415_8145.n3 a_29415_8145.n2 1.6255
R12614 a_29415_8145.n8 a_29415_8145.n5 0.728326
R12615 a_29415_8145.n5 a_29415_8145.n4 0.552239
R12616 OUT.n7 OUT.t27 23.6945
R12617 OUT.t31 OUT.n8 23.6945
R12618 OUT.n34 OUT.t20 23.6945
R12619 OUT.t15 OUT.n35 23.6945
R12620 OUT.n8 OUT.n7 18.8035
R12621 OUT.n35 OUT.n34 18.8035
R12622 OUT.n5 OUT.n3 15.8172
R12623 OUT.n4 OUT.n0 15.8172
R12624 OUT.n5 OUT.n4 15.8172
R12625 OUT.n32 OUT.n30 15.8172
R12626 OUT.n32 OUT.n31 15.8172
R12627 OUT.n31 OUT.n27 15.8172
R12628 OUT.n3 OUT.t16 14.8925
R12629 OUT.t22 OUT.n5 14.8925
R12630 OUT.n4 OUT.t35 14.8925
R12631 OUT.n30 OUT.t34 14.8925
R12632 OUT.t21 OUT.n32 14.8925
R12633 OUT.n31 OUT.t32 14.8925
R12634 OUT.n9 OUT.n1 12.2457
R12635 OUT.n6 OUT.n1 12.2457
R12636 OUT.n6 OUT.n2 12.2457
R12637 OUT.n36 OUT.n28 12.2457
R12638 OUT.n33 OUT.n28 12.2457
R12639 OUT.n33 OUT.n29 12.2457
R12640 OUT.n10 OUT.t23 11.6285
R12641 OUT.n37 OUT.t28 11.6285
R12642 OUT.n2 OUT.t27 8.9065
R12643 OUT.t29 OUT.n6 8.9065
R12644 OUT.t18 OUT.n1 8.9065
R12645 OUT.n9 OUT.t31 8.9065
R12646 OUT.n29 OUT.t20 8.9065
R12647 OUT.t33 OUT.n33 8.9065
R12648 OUT.t19 OUT.n28 8.9065
R12649 OUT.n36 OUT.t15 8.9065
R12650 OUT.n5 OUT.t25 8.6145
R12651 OUT.n3 OUT.t17 8.6145
R12652 OUT.n4 OUT.t14 8.6145
R12653 OUT.n32 OUT.t30 8.6145
R12654 OUT.n30 OUT.t24 8.6145
R12655 OUT.n31 OUT.t12 8.6145
R12656 OUT.n0 OUT.t26 8.59715
R12657 OUT.n27 OUT.t13 8.59715
R12658 OUT.t16 OUT.n2 8.3225
R12659 OUT.n6 OUT.t22 8.3225
R12660 OUT.t35 OUT.n1 8.3225
R12661 OUT.t23 OUT.n9 8.3225
R12662 OUT.t34 OUT.n29 8.3225
R12663 OUT.n33 OUT.t21 8.3225
R12664 OUT.t32 OUT.n28 8.3225
R12665 OUT.t28 OUT.n36 8.3225
R12666 OUT.n40 OUT 4.9636
R12667 OUT OUT.n10 4.223
R12668 OUT OUT.n37 4.223
R12669 OUT.n7 OUT.t29 3.6505
R12670 OUT.n8 OUT.t18 3.6505
R12671 OUT.n34 OUT.t33 3.6505
R12672 OUT.n35 OUT.t19 3.6505
R12673 OUT.n14 OUT.t11 3.6405
R12674 OUT.n14 OUT.n13 3.6405
R12675 OUT.n12 OUT.t2 3.6405
R12676 OUT.n12 OUT.n11 3.6405
R12677 OUT.n21 OUT.t7 3.6405
R12678 OUT.n21 OUT.n20 3.6405
R12679 OUT.n19 OUT.t1 3.6405
R12680 OUT.n19 OUT.n18 3.6405
R12681 OUT.n26 OUT.n17 3.50463
R12682 OUT.n25 OUT.n24 3.50463
R12683 OUT.n17 OUT.t0 3.2765
R12684 OUT.n17 OUT.n16 3.2765
R12685 OUT.n24 OUT.t8 3.2765
R12686 OUT.n24 OUT.n23 3.2765
R12687 OUT.n10 OUT.n0 3.1807
R12688 OUT.n37 OUT.n27 3.1807
R12689 OUT.n15 OUT.n12 3.06224
R12690 OUT.n22 OUT.n19 3.06224
R12691 OUT.n15 OUT.n14 2.6005
R12692 OUT.n22 OUT.n21 2.6005
R12693 OUT OUT.n40 1.41493
R12694 OUT.n38 OUT 1.24006
R12695 OUT.n26 OUT.n25 0.798761
R12696 OUT.n39 OUT.n38 0.611422
R12697 OUT OUT.n26 0.562022
R12698 OUT.n38 OUT 0.247022
R12699 OUT.n40 OUT.n39 0.202264
R12700 OUT.n39 OUT 0.19218
R12701 OUT.n26 OUT.n15 0.18637
R12702 OUT.n25 OUT.n22 0.18637
R12703 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n18 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t12 5.81586
R12704 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n26 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n23 5.10148
R12705 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n22 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n21 5.10116
R12706 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n20 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n19 5.08021
R12707 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n26 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n25 4.66166
R12708 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n10 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t7 3.6405
R12709 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n10 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n9 3.6405
R12710 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n3 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t8 3.6405
R12711 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n3 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n2 3.6405
R12712 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n5 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t5 3.6405
R12713 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n5 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n4 3.6405
R12714 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n12 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t11 3.6405
R12715 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n12 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n11 3.6405
R12716 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n14 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n8 3.50463
R12717 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n15 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n1 3.50463
R12718 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n8 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t2 3.2765
R12719 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n8 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n7 3.2765
R12720 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n1 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t0 3.2765
R12721 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n1 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n0 3.2765
R12722 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n6 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n5 3.06224
R12723 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n13 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n12 3.06224
R12724 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n18 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n17 2.85093
R12725 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n6 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n3 2.6005
R12726 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n13 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n10 2.6005
R12727 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n27 2.36593
R12728 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n17 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t15 2.16717
R12729 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n17 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n16 2.16717
R12730 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n25 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t17 1.9505
R12731 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n25 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n24 1.9505
R12732 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n15 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n14 0.798761
R12733 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n20 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n18 0.644196
R12734 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n15 0.562022
R12735 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n22 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n20 0.450839
R12736 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n27 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n26 0.358498
R12737 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n27 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n22 0.229792
R12738 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n15 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n6 0.18637
R12739 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n14 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n13 0.18637
R12740 a_43828_11254.t0 a_43828_11254.t1 12.9675
R12741 a_43528_10632.t0 a_43528_10632.t1 12.9675
R12742 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n7 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t18 23.6945
R12743 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n8 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t22 23.6945
R12744 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n8 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n7 18.8035
R12745 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n5 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n2 15.8172
R12746 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n11 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n10 15.8172
R12747 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n10 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n2 15.8172
R12748 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t27 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n5 14.8925
R12749 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t25 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n2 14.8925
R12750 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n10 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t23 14.8925
R12751 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n9 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n3 12.2457
R12752 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n9 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n4 12.2457
R12753 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n6 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n4 12.2457
R12754 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n12 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t19 11.6285
R12755 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t18 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n6 8.9065
R12756 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t21 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n4 8.9065
R12757 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n9 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t17 8.9065
R12758 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t22 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n3 8.9065
R12759 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n5 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t16 8.6145
R12760 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n2 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t26 8.6145
R12761 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n10 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t24 8.6145
R12762 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n11 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t20 8.59715
R12763 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n6 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t27 8.3225
R12764 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n4 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t25 8.3225
R12765 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t23 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n9 8.3225
R12766 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n3 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t19 8.3225
R12767 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n1 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t3 6.74566
R12768 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n0 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t10 6.74332
R12769 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n0 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t11 5.1005
R12770 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n1 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t2 5.1005
R12771 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n12 4.223
R12772 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n7 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t21 3.6505
R12773 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t17 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n8 3.6505
R12774 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n19 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n16 3.57508
R12775 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n28 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n27 3.5743
R12776 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n0 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n13 3.40011
R12777 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n1 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n22 3.40001
R12778 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n12 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n11 3.1807
R12779 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n23 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t1 3.00159
R12780 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n14 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t8 3.00158
R12781 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n20 2.58112
R12782 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n29 2.58112
R12783 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n18 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t5 2.16717
R12784 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n18 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n17 2.16717
R12785 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n16 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t6 2.16717
R12786 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n16 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n15 2.16717
R12787 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n25 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t15 2.16717
R12788 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n25 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n24 2.16717
R12789 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n27 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t12 2.16717
R12790 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n27 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n26 2.16717
R12791 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n20 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n14 1.84821
R12792 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n29 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n23 1.84725
R12793 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n19 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n18 1.25233
R12794 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n28 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n25 1.25225
R12795 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n29 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n28 1.12575
R12796 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n20 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n19 1.12554
R12797 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n21 0.784521
R12798 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n21 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT 0.689881
R12799 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n23 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n1 0.55941
R12800 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n14 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n0 0.558372
R12801 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n21 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT 0.25925
R12802 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n29 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t57 23.6945
R12803 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n30 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t40 23.6945
R12804 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n30 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n29 18.8035
R12805 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n27 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n24 15.8172
R12806 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n32 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n24 15.8172
R12807 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n33 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n32 15.8172
R12808 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t41 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n27 14.8925
R12809 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t45 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n24 14.8925
R12810 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n32 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t49 14.8925
R12811 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n31 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n25 12.2457
R12812 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n31 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n26 12.2457
R12813 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n28 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n26 12.2457
R12814 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n34 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t43 11.6285
R12815 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n37 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t51 9.57577
R12816 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n40 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t54 9.55796
R12817 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n66 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t9 9.31704
R12818 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n50 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n44 8.94165
R12819 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t57 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n28 8.9065
R12820 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t52 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n26 8.9065
R12821 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n31 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t33 8.9065
R12822 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t40 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n25 8.9065
R12823 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n27 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t32 8.6145
R12824 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n24 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t37 8.6145
R12825 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n32 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t44 8.6145
R12826 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n33 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t34 8.59715
R12827 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n11 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n10 8.59228
R12828 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n37 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t31 8.56851
R12829 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n38 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t39 8.56851
R12830 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n39 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t38 8.56851
R12831 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t42 8.5214
R12832 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n0 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t35 8.5214
R12833 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n1 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t56 8.5214
R12834 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n6 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t58 8.5214
R12835 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n42 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t47 8.5112
R12836 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n41 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t48 8.5112
R12837 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n40 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t36 8.5112
R12838 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n0 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t53 8.34992
R12839 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n28 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t41 8.3225
R12840 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n26 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t45 8.3225
R12841 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t49 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n31 8.3225
R12842 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n25 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t43 8.3225
R12843 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n67 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n72 8.65114
R12844 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n6 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t50 8.30779
R12845 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n1 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t46 8.30779
R12846 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t55 8.30779
R12847 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n64 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n62 7.40037
R12848 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t26 7.05758
R12849 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n2 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n21 6.80072
R12850 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n11 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n9 6.73941
R12851 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t17 6.45366
R12852 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n22 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t22 6.2092
R12853 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n16 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n15 5.83551
R12854 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n45 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t11 4.89657
R12855 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n64 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n63 4.88218
R12856 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n71 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n70 4.87529
R12857 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n5 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t10 4.6632
R12858 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n55 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t3 4.63112
R12859 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n49 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n48 5.42442
R12860 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n68 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n58 4.54362
R12861 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n34 4.223
R12862 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n65 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n61 4.01867
R12863 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n12 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n8 3.9838
R12864 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n70 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n36 3.96161
R12865 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n65 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n64 3.87403
R12866 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n29 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t52 3.6505
R12867 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t33 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n30 3.6505
R12868 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n48 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t2 3.6405
R12869 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n48 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n47 3.6405
R12870 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n8 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t16 3.6405
R12871 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n8 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n7 3.6405
R12872 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n58 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t7 3.6405
R12873 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n58 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n57 3.6405
R12874 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n60 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t8 3.6405
R12875 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n60 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n59 3.6405
R12876 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n52 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t0 3.6405
R12877 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n52 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n51 3.6405
R12878 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n18 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t30 3.47629
R12879 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n14 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t29 3.47625
R12880 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n20 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t27 3.47617
R12881 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n16 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n14 3.39849
R12882 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n34 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n33 3.1807
R12883 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n20 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n19 2.86157
R12884 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n14 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n13 2.8615
R12885 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n18 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n17 2.86147
R12886 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n18 2.48336
R12887 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n2 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n20 2.47781
R12888 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n35 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN 2.35499
R12889 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n23 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN 2.30073
R12890 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n5 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n54 2.24532
R12891 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n53 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n52 4.81789
R12892 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n54 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n53 2.21522
R12893 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n49 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n46 1.7262
R12894 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n43 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n42 1.61187
R12895 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n43 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n39 1.57365
R12896 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n56 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n55 1.51564
R12897 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n35 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN 1.51518
R12898 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n46 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n45 1.49463
R12899 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n71 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n12 1.36952
R12900 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n61 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n60 1.25753
R12901 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n2 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n3 1.05601
R12902 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n23 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n22 1.01067
R12903 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n41 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n40 0.996664
R12904 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n0 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n4 0.992966
R12905 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n16 0.983287
R12906 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n1 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n0 0.975705
R12907 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n69 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n56 0.969569
R12908 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n70 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n69 0.955885
R12909 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n38 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n37 0.953514
R12910 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n22 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n2 0.907492
R12911 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n66 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n65 0.856289
R12912 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n68 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n67 0.843096
R12913 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n53 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n50 0.8015
R12914 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n12 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n11 0.800717
R12915 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n55 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n5 0.741058
R12916 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n56 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n6 0.69855
R12917 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n69 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n68 0.656716
R12918 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n67 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n66 0.398395
R12919 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n50 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n49 0.3875
R12920 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n39 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n38 0.364199
R12921 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n36 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n23 0.362368
R12922 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n6 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n1 0.359267
R12923 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n42 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n41 0.323514
R12924 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n43 0.319815
R12925 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n36 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n35 0.193979
R12926 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n71 0.147028
R12927 a_22879_10704.n1 a_22879_10704.t2 7.58276
R12928 a_22879_10704.n3 a_22879_10704.n1 7.16556
R12929 a_22879_10704.n1 a_22879_10704.n0 6.4265
R12930 a_22879_10704.n3 a_22879_10704.n2 3.4179
R12931 a_22879_10704.t1 a_22879_10704.n3 2.93981
R12932 mux_magic_1.AND2_magic_0.A.t11 mux_magic_1.AND2_magic_0.A.t12 144.929
R12933 mux_magic_1.AND2_magic_0.A.t9 mux_magic_1.AND2_magic_0.A.t10 44.058
R12934 mux_magic_1.AND2_magic_0.A.n2 mux_magic_1.AND2_magic_0.A.t11 14.796
R12935 mux_magic_1.AND2_magic_0.A.n2 mux_magic_1.AND2_magic_0.A.t9 13.8835
R12936 mux_magic_1.AND2_magic_0.A mux_magic_1.AND2_magic_0.A.n2 9.83788
R12937 mux_magic_1.AND2_magic_0.A.n1 mux_magic_1.AND2_magic_0.A.n4 4.99061
R12938 mux_magic_1.AND2_magic_0.A mux_magic_1.AND2_magic_0.A.n3 4.5405
R12939 mux_magic_1.AND2_magic_0.A.n1 mux_magic_1.AND2_magic_0.A.n11 4.2255
R12940 mux_magic_1.AND2_magic_0.A.n0 mux_magic_1.AND2_magic_0.A.n6 3.52811
R12941 mux_magic_1.AND2_magic_0.A.n0 mux_magic_1.AND2_magic_0.A.n10 3.30485
R12942 mux_magic_1.AND2_magic_0.A.n0 mux_magic_1.AND2_magic_0.A.n8 2.6005
R12943 mux_magic_1.AND2_magic_0.A.n8 mux_magic_1.AND2_magic_0.A.t7 1.6255
R12944 mux_magic_1.AND2_magic_0.A.n8 mux_magic_1.AND2_magic_0.A.n7 1.6255
R12945 mux_magic_1.AND2_magic_0.A.n10 mux_magic_1.AND2_magic_0.A.t5 1.6255
R12946 mux_magic_1.AND2_magic_0.A.n10 mux_magic_1.AND2_magic_0.A.n9 1.6255
R12947 mux_magic_1.AND2_magic_0.A.n6 mux_magic_1.AND2_magic_0.A.t4 1.463
R12948 mux_magic_1.AND2_magic_0.A.n6 mux_magic_1.AND2_magic_0.A.n5 1.463
R12949 mux_magic_1.AND2_magic_0.A.n1 mux_magic_1.AND2_magic_0.A.n0 1.19985
R12950 mux_magic_1.AND2_magic_0.A mux_magic_1.AND2_magic_0.A.n1 0.819535
R12951 a_27875_8520.t6 a_27875_8520.t7 44.058
R12952 a_27875_8520.n3 a_27875_8520.t8 34.6465
R12953 a_27875_8520.n3 a_27875_8520.t6 15.1219
R12954 a_27875_8520.n6 a_27875_8520.t2 5.29595
R12955 a_27875_8520.n4 a_27875_8520.n2 4.97104
R12956 a_27875_8520.n4 a_27875_8520.n3 4.16767
R12957 a_27875_8520.n5 a_27875_8520.n1 3.01333
R12958 a_27875_8520.n7 a_27875_8520.n6 3.01333
R12959 a_27875_8520.n1 a_27875_8520.t4 1.6255
R12960 a_27875_8520.n1 a_27875_8520.n0 1.6255
R12961 a_27875_8520.n7 a_27875_8520.t0 1.6255
R12962 a_27875_8520.n8 a_27875_8520.n7 1.6255
R12963 a_27875_8520.n6 a_27875_8520.n5 0.845717
R12964 a_27875_8520.n5 a_27875_8520.n4 0.423109
R12965 a_19897_10547.t6 a_19897_10547.t7 44.058
R12966 a_19897_10547.n3 a_19897_10547.t8 34.6465
R12967 a_19897_10547.n3 a_19897_10547.t6 15.1219
R12968 a_19897_10547.n6 a_19897_10547.t0 5.29595
R12969 a_19897_10547.n4 a_19897_10547.n2 4.97104
R12970 a_19897_10547.n4 a_19897_10547.n3 4.16767
R12971 a_19897_10547.n5 a_19897_10547.n1 3.01333
R12972 a_19897_10547.n7 a_19897_10547.n6 3.01333
R12973 a_19897_10547.n1 a_19897_10547.t4 1.6255
R12974 a_19897_10547.n1 a_19897_10547.n0 1.6255
R12975 a_19897_10547.n7 a_19897_10547.t3 1.6255
R12976 a_19897_10547.n8 a_19897_10547.n7 1.6255
R12977 a_19897_10547.n6 a_19897_10547.n5 0.845717
R12978 a_19897_10547.n5 a_19897_10547.n4 0.423109
R12979 mux_magic_2.OR_magic_0.B.t4 mux_magic_2.OR_magic_0.B.t7 44.6331
R12980 mux_magic_2.OR_magic_0.B.t3 mux_magic_2.OR_magic_0.B.t4 43.4094
R12981 mux_magic_2.OR_magic_0.B.t5 mux_magic_2.OR_magic_0.B.t3 31.5469
R12982 mux_magic_2.OR_magic_0.B.n0 mux_magic_2.OR_magic_0.B.t5 15.0567
R12983 mux_magic_2.OR_magic_0.B.n0 mux_magic_2.OR_magic_0.B.t6 13.6228
R12984 mux_magic_2.OR_magic_0.B mux_magic_2.OR_magic_0.B.n1 5.03757
R12985 mux_magic_2.OR_magic_0.B mux_magic_2.OR_magic_0.B.n0 4.2675
R12986 mux_magic_2.OR_magic_0.B mux_magic_2.OR_magic_0.B.n3 3.36521
R12987 mux_magic_2.OR_magic_0.B.n3 mux_magic_2.OR_magic_0.B.t1 1.6255
R12988 mux_magic_2.OR_magic_0.B.n3 mux_magic_2.OR_magic_0.B.n2 1.6255
R12989 PFD_T2_0.INV_mag_0.OUT.n4 PFD_T2_0.INV_mag_0.OUT.n3 34.5741
R12990 PFD_T2_0.INV_mag_0.OUT.n3 PFD_T2_0.INV_mag_0.OUT.t8 33.8279
R12991 PFD_T2_0.INV_mag_0.OUT.n0 PFD_T2_0.INV_mag_0.OUT.t3 30.6524
R12992 PFD_T2_0.INV_mag_0.OUT.n1 PFD_T2_0.INV_mag_0.OUT.t4 30.6524
R12993 PFD_T2_0.INV_mag_0.OUT.n0 PFD_T2_0.INV_mag_0.OUT.t7 9.5635
R12994 PFD_T2_0.INV_mag_0.OUT.n1 PFD_T2_0.INV_mag_0.OUT.t5 9.5635
R12995 PFD_T2_0.INV_mag_0.OUT.n5 PFD_T2_0.INV_mag_0.OUT.n4 9.26523
R12996 PFD_T2_0.INV_mag_0.OUT PFD_T2_0.INV_mag_0.OUT.n6 6.74425
R12997 PFD_T2_0.INV_mag_0.OUT.n4 PFD_T2_0.INV_mag_0.OUT.t9 6.5705
R12998 PFD_T2_0.INV_mag_0.OUT.n2 PFD_T2_0.INV_mag_0.OUT.n0 5.32623
R12999 PFD_T2_0.INV_mag_0.OUT.n2 PFD_T2_0.INV_mag_0.OUT.n1 4.78052
R13000 PFD_T2_0.INV_mag_0.OUT PFD_T2_0.INV_mag_0.OUT.n5 4.4032
R13001 PFD_T2_0.INV_mag_0.OUT.n3 PFD_T2_0.INV_mag_0.OUT.t6 3.6505
R13002 PFD_T2_0.INV_mag_0.OUT.n8 PFD_T2_0.INV_mag_0.OUT.t1 3.6405
R13003 PFD_T2_0.INV_mag_0.OUT.n8 PFD_T2_0.INV_mag_0.OUT.n7 3.6405
R13004 PFD_T2_0.INV_mag_0.OUT.n5 PFD_T2_0.INV_mag_0.OUT.n2 3.38996
R13005 PFD_T2_0.INV_mag_0.OUT PFD_T2_0.INV_mag_0.OUT.n8 3.35938
R13006 a_22966_11778.n2 a_22966_11778.t11 33.8126
R13007 a_22966_11778.n3 a_22966_11778.n2 30.3299
R13008 a_22966_11778.n4 a_22966_11778.n3 30.3299
R13009 a_22966_11778.n5 a_22966_11778.n4 30.3299
R13010 a_22966_11778.n6 a_22966_11778.n5 30.3299
R13011 a_22966_11778.n7 a_22966_11778.n6 30.3299
R13012 a_22966_11778.n8 a_22966_11778.n7 30.3299
R13013 a_22966_11778.n9 a_22966_11778.n8 30.3299
R13014 a_22966_11778.n10 a_22966_11778.n9 30.3299
R13015 a_22966_11778.n13 a_22966_11778.t14 26.2932
R13016 a_22966_11778.n11 a_22966_11778.t9 12.8368
R13017 a_22966_11778.n11 a_22966_11778.n10 12.0257
R13018 a_22966_11778.n14 a_22966_11778.n13 8.47283
R13019 a_22966_11778.n12 a_22966_11778.n11 5.21433
R13020 a_22966_11778.n2 a_22966_11778.t4 3.6505
R13021 a_22966_11778.n3 a_22966_11778.t10 3.6505
R13022 a_22966_11778.n4 a_22966_11778.t15 3.6505
R13023 a_22966_11778.n5 a_22966_11778.t6 3.6505
R13024 a_22966_11778.n6 a_22966_11778.t16 3.6505
R13025 a_22966_11778.n7 a_22966_11778.t7 3.6505
R13026 a_22966_11778.n8 a_22966_11778.t12 3.6505
R13027 a_22966_11778.n9 a_22966_11778.t8 3.6505
R13028 a_22966_11778.n10 a_22966_11778.t13 3.6505
R13029 a_22966_11778.n13 a_22966_11778.t5 3.6505
R13030 a_22966_11778.n1 a_22966_11778.t2 3.6405
R13031 a_22966_11778.n1 a_22966_11778.n0 3.6405
R13032 a_22966_11778.n14 a_22966_11778.n12 3.50583
R13033 a_22966_11778.n15 a_22966_11778.t0 3.38777
R13034 a_22966_11778.n16 a_22966_11778.n15 2.97653
R13035 a_22966_11778.n15 a_22966_11778.n14 2.47455
R13036 a_22966_11778.n12 a_22966_11778.n1 1.25598
R13037 S3.t5 S3.t12 144.929
R13038 S3.t0 S3.t1 44.058
R13039 S3.n1 S3.t9 25.9486
R13040 S3.t9 S3 16.1689
R13041 S3.n4 S3.n3 15.8172
R13042 S3.n5 S3.n4 15.8172
R13043 S3.n0 S3.t5 14.796
R13044 S3.n6 S3.t3 14.4701
R13045 S3.n0 S3.t0 13.8835
R13046 S3.n2 S3.n1 13.2388
R13047 S3.n2 S3.t6 12.7103
R13048 S3.n3 S3.t7 11.7326
R13049 S3.n3 S3.t4 11.7326
R13050 S3.n4 S3.t10 11.7326
R13051 S3.n4 S3.t8 11.7326
R13052 S3.n5 S3.t11 11.7326
R13053 S3.t3 S3.n5 11.7326
R13054 S3 S3.n0 9.83788
R13055 S3.n1 S3.t2 7.3005
R13056 S3 S3.n6 4.18916
R13057 S3.n6 S3.n2 1.49961
R13058 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n9 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t13 14.1829
R13059 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n8 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t12 13.9657
R13060 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n2 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t20 13.3574
R13061 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n1 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t17 13.1401
R13062 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n1 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t14 12.9025
R13063 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n3 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t16 12.6187
R13064 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n4 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t21 8.77788
R13065 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n5 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t19 8.64752
R13066 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n5 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t15 8.56062
R13067 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n4 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t18 8.43026
R13068 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n6 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n5 6.11825
R13069 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n6 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n4 5.88354
R13070 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n11 4.64372
R13071 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n22 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t8 3.6405
R13072 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n22 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n21 3.6405
R13073 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n15 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t6 3.6405
R13074 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n15 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n14 3.6405
R13075 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n17 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t5 3.6405
R13076 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n17 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n16 3.6405
R13077 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n24 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t7 3.6405
R13078 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n24 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n23 3.6405
R13079 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n26 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n20 3.50463
R13080 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n27 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n13 3.50463
R13081 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n20 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t2 3.2765
R13082 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n20 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n19 3.2765
R13083 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n13 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t1 3.2765
R13084 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n13 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n12 3.2765
R13085 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n18 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n17 3.06224
R13086 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n25 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n24 3.06224
R13087 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n18 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n15 2.6005
R13088 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n25 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n22 2.6005
R13089 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n11 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT 2.32194
R13090 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n0 2.31638
R13091 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n0 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n10 2.2505
R13092 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n8 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n7 1.58291
R13093 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n7 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n3 1.47586
R13094 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n10 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n9 1.33917
R13095 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n9 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n8 1.23958
R13096 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n27 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n26 0.798761
R13097 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n27 0.562022
R13098 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n7 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n6 0.448735
R13099 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n3 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n2 0.386992
R13100 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n2 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n1 0.340685
R13101 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n27 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n18 0.18637
R13102 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n26 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n25 0.18637
R13103 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n11 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n0 0.130397
R13104 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n26 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t23 45.6363
R13105 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n22 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t30 45.6363
R13106 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n17 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t15 29.6446
R13107 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t16 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n18 29.6446
R13108 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n19 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t20 29.6446
R13109 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t19 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n20 29.6446
R13110 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n16 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t21 24.6117
R13111 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n21 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t28 24.6117
R13112 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n18 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n17 22.2047
R13113 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n20 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n19 22.2047
R13114 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t23 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t29 22.1925
R13115 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t30 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t18 22.1925
R13116 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t16 21.8613
R13117 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n27 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n26 20.9314
R13118 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n23 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n22 20.9314
R13119 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n25 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t19 17.8613
R13120 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n28 10.8592
R13121 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n25 8.94379
R13122 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n16 8.87094
R13123 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n26 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t27 6.1325
R13124 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n27 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t25 6.1325
R13125 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n17 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t31 6.1325
R13126 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n18 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t14 6.1325
R13127 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n16 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t13 6.1325
R13128 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n19 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t17 6.1325
R13129 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n20 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t22 6.1325
R13130 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n21 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t12 6.1325
R13131 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n22 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t24 6.1325
R13132 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n23 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t26 6.1325
R13133 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n24 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n23 5.38991
R13134 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n28 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n27 5.12094
R13135 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n24 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n21 4.83094
R13136 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n10 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t7 3.6405
R13137 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n10 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n9 3.6405
R13138 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n3 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t9 3.6405
R13139 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n3 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n2 3.6405
R13140 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n5 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t5 3.6405
R13141 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n5 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n4 3.6405
R13142 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n12 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t11 3.6405
R13143 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n12 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n11 3.6405
R13144 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n14 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n8 3.50463
R13145 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n15 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n1 3.50463
R13146 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n8 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t1 3.2765
R13147 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n8 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n7 3.2765
R13148 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n1 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t2 3.2765
R13149 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n1 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n0 3.2765
R13150 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n6 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n5 3.06224
R13151 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n13 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n12 3.06224
R13152 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n6 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n3 2.6005
R13153 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n13 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n10 2.6005
R13154 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n28 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK 1.07267
R13155 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n15 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n14 0.798761
R13156 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n24 0.658318
R13157 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n25 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK 0.628846
R13158 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n15 0.562022
R13159 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n15 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n6 0.18637
R13160 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n14 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n13 0.18637
R13161 a_44716_n517.n0 a_44716_n517.t6 29.2961
R13162 a_44716_n517.n1 a_44716_n517.n0 21.9292
R13163 a_44716_n517.n2 a_44716_n517.n1 18.1271
R13164 a_44716_n517.n2 a_44716_n517.t7 11.1695
R13165 a_44716_n517.n0 a_44716_n517.t8 6.1325
R13166 a_44716_n517.n1 a_44716_n517.t9 6.1325
R13167 a_44716_n517.n6 a_44716_n517.n5 4.93252
R13168 a_44716_n517.n6 a_44716_n517.t1 4.70348
R13169 a_44716_n517.n8 a_44716_n517.n2 4.6311
R13170 a_44716_n517.n9 a_44716_n517.n8 2.85093
R13171 a_44716_n517.n4 a_44716_n517.t2 2.16717
R13172 a_44716_n517.n4 a_44716_n517.n3 2.16717
R13173 a_44716_n517.n9 a_44716_n517.t3 2.16717
R13174 a_44716_n517.n10 a_44716_n517.n9 2.16717
R13175 a_44716_n517.n7 a_44716_n517.n6 1.58582
R13176 a_44716_n517.n7 a_44716_n517.n4 1.24371
R13177 a_44716_n517.n8 a_44716_n517.n7 0.971051
R13178 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n21 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t16 23.6945
R13179 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n22 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t22 23.6945
R13180 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n22 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n21 18.8035
R13181 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n19 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n16 15.8172
R13182 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n24 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n16 15.8172
R13183 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n25 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n24 15.8172
R13184 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t18 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n19 14.8925
R13185 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t20 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n16 14.8925
R13186 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n24 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t23 14.8925
R13187 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n23 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n17 12.2457
R13188 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n23 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n18 12.2457
R13189 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n20 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n18 12.2457
R13190 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n26 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t13 11.6285
R13191 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t16 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n20 8.9065
R13192 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t17 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n18 8.9065
R13193 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n23 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t15 8.9065
R13194 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t22 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n17 8.9065
R13195 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n19 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t19 8.6145
R13196 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n16 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t21 8.6145
R13197 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n24 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t12 8.6145
R13198 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n25 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t14 8.59715
R13199 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n20 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t18 8.3225
R13200 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n18 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t20 8.3225
R13201 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t23 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n23 8.3225
R13202 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n17 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t13 8.3225
R13203 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n26 4.223
R13204 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n21 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t17 3.6505
R13205 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t15 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n22 3.6505
R13206 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n12 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t8 3.6405
R13207 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n12 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n11 3.6405
R13208 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n1 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t5 3.6405
R13209 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n1 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n0 3.6405
R13210 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t7 3.6405
R13211 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n2 3.6405
R13212 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n10 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t10 3.6405
R13213 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n10 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n9 3.6405
R13214 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n14 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n8 3.50463
R13215 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n15 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n6 3.50463
R13216 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n8 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t2 3.2765
R13217 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n8 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n7 3.2765
R13218 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n6 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t1 3.2765
R13219 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n6 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n5 3.2765
R13220 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n26 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n25 3.1807
R13221 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n1 3.06224
R13222 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n13 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n10 3.06224
R13223 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n3 2.6005
R13224 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n13 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n12 2.6005
R13225 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n15 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n14 0.798761
R13226 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n15 0.562022
R13227 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n15 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n4 0.18637
R13228 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n14 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n13 0.18637
R13229 VCO_DFF_C_0.VCO_C_0.OUT.n24 VCO_DFF_C_0.VCO_C_0.OUT.t14 14.1829
R13230 VCO_DFF_C_0.VCO_C_0.OUT.n23 VCO_DFF_C_0.VCO_C_0.OUT.t21 13.9657
R13231 VCO_DFF_C_0.VCO_C_0.OUT.n17 VCO_DFF_C_0.VCO_C_0.OUT.t18 13.3574
R13232 VCO_DFF_C_0.VCO_C_0.OUT.n16 VCO_DFF_C_0.VCO_C_0.OUT.t15 13.1401
R13233 VCO_DFF_C_0.VCO_C_0.OUT.n16 VCO_DFF_C_0.VCO_C_0.OUT.t16 12.9025
R13234 VCO_DFF_C_0.VCO_C_0.OUT.n18 VCO_DFF_C_0.VCO_C_0.OUT.t17 12.6187
R13235 VCO_DFF_C_0.VCO_C_0.OUT.n20 VCO_DFF_C_0.VCO_C_0.OUT.t20 8.77788
R13236 VCO_DFF_C_0.VCO_C_0.OUT.n19 VCO_DFF_C_0.VCO_C_0.OUT.t12 8.64752
R13237 VCO_DFF_C_0.VCO_C_0.OUT.n19 VCO_DFF_C_0.VCO_C_0.OUT.t19 8.56062
R13238 VCO_DFF_C_0.VCO_C_0.OUT.n20 VCO_DFF_C_0.VCO_C_0.OUT.t13 8.43026
R13239 VCO_DFF_C_0.VCO_C_0.OUT.n21 VCO_DFF_C_0.VCO_C_0.OUT.n19 6.11825
R13240 VCO_DFF_C_0.VCO_C_0.OUT.n21 VCO_DFF_C_0.VCO_C_0.OUT.n20 5.88354
R13241 VCO_DFF_C_0.VCO_C_0.OUT.n10 VCO_DFF_C_0.VCO_C_0.OUT.t5 3.6405
R13242 VCO_DFF_C_0.VCO_C_0.OUT.n10 VCO_DFF_C_0.VCO_C_0.OUT.n9 3.6405
R13243 VCO_DFF_C_0.VCO_C_0.OUT.n3 VCO_DFF_C_0.VCO_C_0.OUT.t6 3.6405
R13244 VCO_DFF_C_0.VCO_C_0.OUT.n3 VCO_DFF_C_0.VCO_C_0.OUT.n2 3.6405
R13245 VCO_DFF_C_0.VCO_C_0.OUT.n1 VCO_DFF_C_0.VCO_C_0.OUT.t8 3.6405
R13246 VCO_DFF_C_0.VCO_C_0.OUT.n1 VCO_DFF_C_0.VCO_C_0.OUT.n0 3.6405
R13247 VCO_DFF_C_0.VCO_C_0.OUT.n12 VCO_DFF_C_0.VCO_C_0.OUT.t11 3.6405
R13248 VCO_DFF_C_0.VCO_C_0.OUT.n12 VCO_DFF_C_0.VCO_C_0.OUT.n11 3.6405
R13249 VCO_DFF_C_0.VCO_C_0.OUT.n14 VCO_DFF_C_0.VCO_C_0.OUT.n8 3.50463
R13250 VCO_DFF_C_0.VCO_C_0.OUT.n15 VCO_DFF_C_0.VCO_C_0.OUT.n6 3.50463
R13251 VCO_DFF_C_0.VCO_C_0.OUT.n8 VCO_DFF_C_0.VCO_C_0.OUT.t2 3.2765
R13252 VCO_DFF_C_0.VCO_C_0.OUT.n8 VCO_DFF_C_0.VCO_C_0.OUT.n7 3.2765
R13253 VCO_DFF_C_0.VCO_C_0.OUT.n6 VCO_DFF_C_0.VCO_C_0.OUT.t0 3.2765
R13254 VCO_DFF_C_0.VCO_C_0.OUT.n6 VCO_DFF_C_0.VCO_C_0.OUT.n5 3.2765
R13255 VCO_DFF_C_0.VCO_C_0.OUT.n4 VCO_DFF_C_0.VCO_C_0.OUT.n1 3.06224
R13256 VCO_DFF_C_0.VCO_C_0.OUT.n13 VCO_DFF_C_0.VCO_C_0.OUT.n10 3.06224
R13257 VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.OUT.n24 2.91964
R13258 VCO_DFF_C_0.VCO_C_0.OUT.n4 VCO_DFF_C_0.VCO_C_0.OUT.n3 2.6005
R13259 VCO_DFF_C_0.VCO_C_0.OUT.n13 VCO_DFF_C_0.VCO_C_0.OUT.n12 2.6005
R13260 VCO_DFF_C_0.VCO_C_0.OUT.n23 VCO_DFF_C_0.VCO_C_0.OUT.n22 1.58291
R13261 VCO_DFF_C_0.VCO_C_0.OUT.n22 VCO_DFF_C_0.VCO_C_0.OUT.n18 1.47586
R13262 VCO_DFF_C_0.VCO_C_0.OUT.n24 VCO_DFF_C_0.VCO_C_0.OUT.n23 1.23958
R13263 VCO_DFF_C_0.VCO_C_0.OUT.n15 VCO_DFF_C_0.VCO_C_0.OUT.n14 0.798761
R13264 VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.OUT.n15 0.561439
R13265 VCO_DFF_C_0.VCO_C_0.OUT.n22 VCO_DFF_C_0.VCO_C_0.OUT.n21 0.448735
R13266 VCO_DFF_C_0.VCO_C_0.OUT.n18 VCO_DFF_C_0.VCO_C_0.OUT.n17 0.386992
R13267 VCO_DFF_C_0.VCO_C_0.OUT.n17 VCO_DFF_C_0.VCO_C_0.OUT.n16 0.340685
R13268 VCO_DFF_C_0.VCO_C_0.OUT.n15 VCO_DFF_C_0.VCO_C_0.OUT.n4 0.18637
R13269 VCO_DFF_C_0.VCO_C_0.OUT.n14 VCO_DFF_C_0.VCO_C_0.OUT.n13 0.18637
R13270 a_22880_9797.t1 a_22880_9797.n3 7.58276
R13271 a_22880_9797.n3 a_22880_9797.n1 7.1657
R13272 a_22880_9797.n3 a_22880_9797.n2 6.4265
R13273 a_22880_9797.n1 a_22880_9797.n0 3.41789
R13274 a_22880_9797.n1 a_22880_9797.t2 2.93982
R13275 ITAIL1.n5 ITAIL1.n4 28.0418
R13276 ITAIL1.n3 ITAIL1.n2 14.6005
R13277 ITAIL1.n1 ITAIL1.n0 7.61735
R13278 ITAIL1.n1 ITAIL1.t7 7.20135
R13279 ITAIL1.n8 ITAIL1.n7 6.82463
R13280 ITAIL1.n10 ITAIL1.t4 6.77907
R13281 ITAIL1.n5 ITAIL1.t0 6.71389
R13282 ITAIL1.n2 ITAIL1.t11 6.51836
R13283 ITAIL1.n2 ITAIL1.t2 6.51836
R13284 ITAIL1.n3 ITAIL1.t10 6.51836
R13285 ITAIL1.n10 ITAIL1.t12 6.25764
R13286 ITAIL1.n4 ITAIL1.t6 6.25764
R13287 ITAIL1.n6 ITAIL1.t13 6.19246
R13288 ITAIL1.n11 ITAIL1.t5 5.89613
R13289 ITAIL1.n11 ITAIL1.n10 4.23548
R13290 ITAIL1.n8 ITAIL1.n6 4.21461
R13291 ITAIL1.n13 ITAIL1 2.59768
R13292 ITAIL1 ITAIL1.n13 2.36014
R13293 ITAIL1.n9 ITAIL1.n8 1.42665
R13294 ITAIL1.n12 ITAIL1.n11 1.13763
R13295 ITAIL1.n13 ITAIL1.n12 0.501708
R13296 ITAIL1.n12 ITAIL1.n9 0.474918
R13297 ITAIL1.n4 ITAIL1.n3 0.261214
R13298 ITAIL1.n9 ITAIL1.n1 0.2105
R13299 ITAIL1.n6 ITAIL1.n5 0.130857
R13300 UP.n1 UP.n0 14.6005
R13301 UP.n3 UP.n2 12.8446
R13302 UP.n0 UP.t3 6.51836
R13303 UP.n0 UP.t7 6.51836
R13304 UP.n1 UP.t5 6.51836
R13305 UP.n3 UP.t4 6.388
R13306 UP.n2 UP.t6 6.19246
R13307 UP.n10 UP.n9 5.47387
R13308 UP.n4 UP.n3 5.03263
R13309 UP.n11 UP.n7 4.65398
R13310 UP.n10 UP.n8 4.2255
R13311 UP.n5 UP 2.32152
R13312 UP.n6 UP 2.0124
R13313 UP UP.n4 1.20571
R13314 UP.n6 UP.n5 0.85728
R13315 UP.n12 UP.n6 0.515191
R13316 UP.n11 UP.n10 0.427022
R13317 UP.n2 UP.n1 0.326393
R13318 UP.n12 UP 0.283382
R13319 UP UP.n11 0.257096
R13320 UP.n5 UP.n4 0.124995
R13321 UP UP.n12 0.00534345
R13322 a_31940_9626.n3 a_31940_9626.n2 10.1602
R13323 a_31940_9626.n1 a_31940_9626.n0 5.4005
R13324 a_31940_9626.n1 a_31940_9626.t2 5.4005
R13325 a_31940_9626.n7 a_31940_9626.n6 5.4005
R13326 a_31940_9626.n7 a_31940_9626.t6 5.4005
R13327 a_31940_9626.n5 a_31940_9626.n4 5.4005
R13328 a_31940_9626.n5 a_31940_9626.t5 5.4005
R13329 a_31940_9626.n10 a_31940_9626.t0 5.4005
R13330 a_31940_9626.n11 a_31940_9626.n10 5.4005
R13331 a_31940_9626.n8 a_31940_9626.n5 3.51269
R13332 a_31940_9626.n10 a_31940_9626.n9 3.31203
R13333 a_31940_9626.n3 a_31940_9626.n1 3.28072
R13334 a_31940_9626.n8 a_31940_9626.n7 3.1505
R13335 a_31940_9626.n9 a_31940_9626.n3 1.46985
R13336 a_31940_9626.n9 a_31940_9626.n8 1.03855
R13337 DIV_OUT.t3 DIV_OUT.t2 44.058
R13338 DIV_OUT.n0 DIV_OUT.t0 38.8649
R13339 DIV_OUT.t0 DIV_OUT.t3 28.6791
R13340 DIV_OUT.n0 DIV_OUT.t1 7.3005
R13341 DIV_OUT DIV_OUT.n0 5.27587
R13342 a_20103_8443.n3 a_20103_8443.n2 6.04536
R13343 a_20103_8443.n2 a_20103_8443.n1 1.5502
R13344 a_20103_8443.t2 a_20103_8443.n3 1.463
R13345 a_20103_8443.n3 a_20103_8443.n0 1.463
R13346 a_20103_8443.n2 a_20103_8443.t0 1.33385
R13347 a_44728_10426.t0 a_44728_10426.t1 12.9675
R13348 a_44428_9804.t0 a_44428_9804.t1 12.9675
R13349 S4.n16 S4.t18 45.6363
R13350 S4.n12 S4.t13 29.6446
R13351 S4.t14 S4.n13 29.6446
R13352 S4.n11 S4.t20 24.6117
R13353 S4.n5 S4.t6 23.6945
R13354 S4.n6 S4.t12 23.6945
R13355 S4.n13 S4.n12 22.2047
R13356 S4.t18 S4.t3 22.1925
R13357 S4.n17 S4.n16 20.9314
R13358 S4.n6 S4.n5 18.8035
R13359 S4 S4.t14 18.5175
R13360 S4.n3 S4.n0 15.8172
R13361 S4.n9 S4.n8 15.8172
R13362 S4.n8 S4.n0 15.8172
R13363 S4.t9 S4.n3 14.8925
R13364 S4.t15 S4.n0 14.8925
R13365 S4.n8 S4.t4 14.8925
R13366 S4.n7 S4.n1 12.2457
R13367 S4.n7 S4.n2 12.2457
R13368 S4.n4 S4.n2 12.2457
R13369 S4.n10 S4.t16 11.6285
R13370 S4.t6 S4.n4 8.9065
R13371 S4.t11 S4.n2 8.9065
R13372 S4.n7 S4.t0 8.9065
R13373 S4.t12 S4.n1 8.9065
R13374 S4.n3 S4.t10 8.6145
R13375 S4.n0 S4.t17 8.6145
R13376 S4.n8 S4.t5 8.6145
R13377 S4.n9 S4.t19 8.59715
R13378 S4.n4 S4.t9 8.3225
R13379 S4.n2 S4.t15 8.3225
R13380 S4.t4 S4.n7 8.3225
R13381 S4.n1 S4.t16 8.3225
R13382 S4.n11 S4.t7 6.1325
R13383 S4.n12 S4.t1 6.1325
R13384 S4.n13 S4.t2 6.1325
R13385 S4.n16 S4.t8 6.1325
R13386 S4.n17 S4.t21 6.1325
R13387 S4.n18 S4.n17 4.86779
R13388 S4.n14 S4.n11 4.79907
R13389 S4 S4.n10 4.223
R13390 S4.n5 S4.t11 3.6505
R13391 S4.t0 S4.n6 3.6505
R13392 S4.n10 S4.n9 3.1807
R13393 S4.n19 S4.n18 2.65123
R13394 S4.n14 S4 0.640368
R13395 S4.n15 S4 0.1655
R13396 S4.n18 S4.n15 0.109537
R13397 S4.n19 S4 0.0733182
R13398 S4.n15 S4.n14 0.0592755
R13399 S4 S4.n19 0.0318393
R13400 a_42628_9598.t0 a_42628_9598.t1 12.9675
R13401 a_42928_8976.t0 a_42928_8976.t1 12.9675
R13402 a_44728_12082.t0 a_44728_12082.t1 12.9675
R13403 a_44428_11460.t0 a_44428_11460.t1 12.9675
R13404 a_20103_9637.n2 a_20103_9637.n1 6.04392
R13405 a_20103_9637.n3 a_20103_9637.n2 1.55019
R13406 a_20103_9637.n1 a_20103_9637.t0 1.463
R13407 a_20103_9637.n1 a_20103_9637.n0 1.463
R13408 a_20103_9637.n2 a_20103_9637.t2 1.33386
R13409 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n3 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n2 5.81586
R13410 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n8 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t0 5.10148
R13411 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n5 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t1 5.1005
R13412 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n4 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t16 5.08021
R13413 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n8 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n7 4.66266
R13414 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n19 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t10 3.6405
R13415 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n19 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n18 3.6405
R13416 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n21 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t5 3.6405
R13417 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n21 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n20 3.6405
R13418 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n12 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t6 3.6405
R13419 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n12 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n11 3.6405
R13420 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n14 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t15 3.6405
R13421 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n14 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n13 3.6405
R13422 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n23 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n17 3.50463
R13423 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n24 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n10 3.50463
R13424 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n17 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t13 3.2765
R13425 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n17 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n16 3.2765
R13426 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n10 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t9 3.2765
R13427 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n10 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n9 3.2765
R13428 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n22 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n21 3.06224
R13429 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n15 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n14 3.06224
R13430 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n3 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n1 2.85093
R13431 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n22 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n19 2.6005
R13432 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n15 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n12 2.6005
R13433 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n1 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t19 2.16717
R13434 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n1 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n0 2.16717
R13435 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n7 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t2 1.9505
R13436 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n7 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n6 1.9505
R13437 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n24 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n23 0.798761
R13438 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n4 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n3 0.644196
R13439 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n24 0.562022
R13440 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n5 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n4 0.447229
R13441 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n5 0.392597
R13442 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n8 0.308628
R13443 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n23 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n22 0.18637
R13444 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n24 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n15 0.18637
R13445 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n27 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t27 23.6945
R13446 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n28 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t16 23.6945
R13447 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n28 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n27 18.8035
R13448 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n25 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n22 15.8172
R13449 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n31 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n30 15.8172
R13450 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n30 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n22 15.8172
R13451 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t26 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n25 14.8925
R13452 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t25 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n22 14.8925
R13453 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n30 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t22 14.8925
R13454 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n29 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n23 12.2457
R13455 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n29 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n24 12.2457
R13456 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n26 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n24 12.2457
R13457 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n32 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t20 11.6285
R13458 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t27 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n26 8.9065
R13459 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t18 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n24 8.9065
R13460 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n29 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t24 8.9065
R13461 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t16 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n23 8.9065
R13462 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n25 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t23 8.6145
R13463 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n22 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t21 8.6145
R13464 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n30 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t19 8.6145
R13465 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n31 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t17 8.59715
R13466 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n26 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t26 8.3225
R13467 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n24 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t25 8.3225
R13468 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t22 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n29 8.3225
R13469 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n23 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t20 8.3225
R13470 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n33 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN 6.97731
R13471 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n0 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n18 6.74326
R13472 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n1 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n7 6.74324
R13473 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n0 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n19 5.1005
R13474 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n1 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n8 5.1005
R13475 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n32 4.21749
R13476 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n27 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t18 3.6505
R13477 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t24 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n28 3.6505
R13478 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n6 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n3 3.57508
R13479 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n16 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n15 3.5743
R13480 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n1 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t5 3.40075
R13481 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n0 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t0 3.40065
R13482 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n32 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n31 3.1807
R13483 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n10 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n9 3.00095
R13484 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n20 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n17 3.00034
R13485 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n21 2.58093
R13486 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n11 2.58093
R13487 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n13 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t11 2.16717
R13488 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n13 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n12 2.16717
R13489 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n15 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t8 2.16717
R13490 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n15 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n14 2.16717
R13491 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n5 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t13 2.16717
R13492 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n5 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n4 2.16717
R13493 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n3 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t14 2.16717
R13494 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n3 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n2 2.16717
R13495 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n11 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n10 1.84762
R13496 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n21 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n20 1.847
R13497 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n6 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n5 1.25233
R13498 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n16 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n13 1.25225
R13499 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n21 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n16 1.12594
R13500 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n11 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n6 1.12574
R13501 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n33 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN 0.812356
R13502 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n33 0.728851
R13503 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n20 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n0 0.559412
R13504 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n10 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n1 0.557726
R13505 a_21437_10708.t8 a_21437_10708.t7 31.5469
R13506 a_21437_10708.n4 a_21437_10708.t8 13.2715
R13507 a_21437_10708.n4 a_21437_10708.t6 13.0934
R13508 a_21437_10708.n0 a_21437_10708.t5 6.52735
R13509 a_21437_10708.n0 a_21437_10708.n4 4.33404
R13510 a_21437_10708.n6 a_21437_10708.n1 4.2255
R13511 a_21437_10708.n5 a_21437_10708.n2 4.2255
R13512 a_21437_10708.n8 a_21437_10708.n6 3.81956
R13513 a_21437_10708.n0 a_21437_10708.n3 2.62633
R13514 a_21437_10708.t0 a_21437_10708.n8 1.6255
R13515 a_21437_10708.n8 a_21437_10708.n7 1.6255
R13516 a_21437_10708.n6 a_21437_10708.n5 0.947457
R13517 a_21437_10708.n5 a_21437_10708.n0 0.602634
R13518 PFD_T2_0.FIN.n0 PFD_T2_0.FIN.t5 12.4835
R13519 PFD_T2_0.FIN.n2 PFD_T2_0.FIN.t4 11.5345
R13520 PFD_T2_0.FIN.n0 PFD_T2_0.FIN.t3 11.4615
R13521 PFD_T2_0.FIN.n1 PFD_T2_0.FIN.t6 11.4615
R13522 PFD_T2_0.FIN.n1 PFD_T2_0.FIN.n0 10.6935
R13523 PFD_T2_0.FIN.n5 PFD_T2_0.FIN.n4 5.47387
R13524 PFD_T2_0.FIN PFD_T2_0.FIN.n2 5.24808
R13525 PFD_T2_0.FIN.n7 PFD_T2_0.FIN.n6 4.65398
R13526 PFD_T2_0.FIN.n5 PFD_T2_0.FIN.n3 4.2255
R13527 PFD_T2_0.FIN.n2 PFD_T2_0.FIN.n1 0.9495
R13528 PFD_T2_0.FIN PFD_T2_0.FIN.n7 0.44667
R13529 PFD_T2_0.FIN.n7 PFD_T2_0.FIN.n5 0.427022
R13530 a_41879_1284.n2 a_41879_1284.t6 29.3691
R13531 a_41879_1284.n3 a_41879_1284.n2 21.9292
R13532 a_41879_1284.n4 a_41879_1284.n3 18.1271
R13533 a_41879_1284.n4 a_41879_1284.t8 11.2425
R13534 a_41879_1284.n7 a_41879_1284.t0 10.2135
R13535 a_41879_1284.n2 a_41879_1284.t7 6.1325
R13536 a_41879_1284.n3 a_41879_1284.t9 6.1325
R13537 a_41879_1284.n7 a_41879_1284.n6 4.68398
R13538 a_41879_1284.n5 a_41879_1284.n4 4.6302
R13539 a_41879_1284.n5 a_41879_1284.n1 2.85093
R13540 a_41879_1284.n1 a_41879_1284.t2 2.16717
R13541 a_41879_1284.n1 a_41879_1284.n0 2.16717
R13542 a_41879_1284.n9 a_41879_1284.t3 2.16717
R13543 a_41879_1284.n10 a_41879_1284.n9 2.16717
R13544 a_41879_1284.n8 a_41879_1284.n7 1.58618
R13545 a_41879_1284.n9 a_41879_1284.n8 1.24388
R13546 a_41879_1284.n8 a_41879_1284.n5 0.97169
R13547 S2.t1 S2.t0 144.929
R13548 S2.t6 S2.t2 44.058
R13549 S2.n4 S2.t10 25.8834
R13550 S2.t10 S2 16.2341
R13551 S2.n1 S2.n0 15.8172
R13552 S2.n2 S2.n1 15.8172
R13553 S2.n3 S2.t1 14.7309
R13554 S2.n6 S2.t4 14.5353
R13555 S2.n3 S2.t6 13.9487
R13556 S2.n5 S2.n4 13.2388
R13557 S2.n5 S2.t11 12.6451
R13558 S2.n0 S2.t7 11.7326
R13559 S2.n0 S2.t3 11.7326
R13560 S2.n1 S2.t12 11.7326
R13561 S2.n1 S2.t9 11.7326
R13562 S2.n2 S2.t8 11.7326
R13563 S2.t4 S2.n2 11.7326
R13564 S2 S2.n3 9.83788
R13565 S2.n4 S2.t5 7.3005
R13566 S2 S2.n6 4.18916
R13567 S2.n6 S2.n5 1.49961
R13568 a_27922_10564.n3 a_27922_10564.n1 6.04375
R13569 a_27922_10564.n3 a_27922_10564.n2 1.55052
R13570 a_27922_10564.n1 a_27922_10564.t3 1.463
R13571 a_27922_10564.n1 a_27922_10564.n0 1.463
R13572 a_27922_10564.t0 a_27922_10564.n3 1.3335
R13573 a_27722_10564.t8 a_27722_10564.t7 44.058
R13574 a_27722_10564.n3 a_27722_10564.t6 34.6465
R13575 a_27722_10564.n3 a_27722_10564.t8 15.1219
R13576 a_27722_10564.n6 a_27722_10564.t2 5.29595
R13577 a_27722_10564.n4 a_27722_10564.n2 4.97104
R13578 a_27722_10564.n4 a_27722_10564.n3 4.16767
R13579 a_27722_10564.n5 a_27722_10564.n1 3.01333
R13580 a_27722_10564.n8 a_27722_10564.n6 3.01333
R13581 a_27722_10564.n1 a_27722_10564.t4 1.6255
R13582 a_27722_10564.n1 a_27722_10564.n0 1.6255
R13583 a_27722_10564.t1 a_27722_10564.n8 1.6255
R13584 a_27722_10564.n8 a_27722_10564.n7 1.6255
R13585 a_27722_10564.n6 a_27722_10564.n5 0.845717
R13586 a_27722_10564.n5 a_27722_10564.n4 0.423109
R13587 S1.t1 S1.t7 144.929
R13588 S1.t9 S1.t11 44.058
R13589 S1.n4 S1.t6 25.8834
R13590 S1.t6 S1 16.2341
R13591 S1.n1 S1.n0 15.8172
R13592 S1.n2 S1.n1 15.8172
R13593 S1.n3 S1.t1 14.7309
R13594 S1.n6 S1.t3 14.5353
R13595 S1.n3 S1.t9 13.9487
R13596 S1.n5 S1.n4 13.2388
R13597 S1.n5 S1.t12 12.6451
R13598 S1.n0 S1.t2 11.7326
R13599 S1.n0 S1.t10 11.7326
R13600 S1.n1 S1.t8 11.7326
R13601 S1.n1 S1.t4 11.7326
R13602 S1.n2 S1.t5 11.7326
R13603 S1.t3 S1.n2 11.7326
R13604 S1 S1.n3 9.83788
R13605 S1.n4 S1.t0 7.3005
R13606 S1 S1.n6 4.18916
R13607 S1.n6 S1.n5 1.49961
R13608 a_44428_11254.t0 a_44428_11254.t1 12.9675
R13609 a_44728_10632.t0 a_44728_10632.t1 12.9675
R13610 PRE_SCALAR.t0 PRE_SCALAR.t2 44.058
R13611 PRE_SCALAR.n0 PRE_SCALAR.t1 38.8649
R13612 PRE_SCALAR.t1 PRE_SCALAR.t0 28.6791
R13613 PRE_SCALAR.n0 PRE_SCALAR.t3 7.3005
R13614 PRE_SCALAR PRE_SCALAR.n0 5.27587
R13615 mux_magic_0.AND2_magic_0.A.t10 mux_magic_0.AND2_magic_0.A.t9 144.929
R13616 mux_magic_0.AND2_magic_0.A.t12 mux_magic_0.AND2_magic_0.A.t11 44.058
R13617 mux_magic_0.AND2_magic_0.A.n0 mux_magic_0.AND2_magic_0.A.t10 14.7309
R13618 mux_magic_0.AND2_magic_0.A.n0 mux_magic_0.AND2_magic_0.A.t12 13.9487
R13619 mux_magic_0.AND2_magic_0.A mux_magic_0.AND2_magic_0.A.n0 9.83788
R13620 mux_magic_0.AND2_magic_0.A.n11 mux_magic_0.AND2_magic_0.A.n2 4.99061
R13621 mux_magic_0.AND2_magic_0.A.n14 mux_magic_0.AND2_magic_0.A.n1 4.5405
R13622 mux_magic_0.AND2_magic_0.A.n13 mux_magic_0.AND2_magic_0.A.n12 4.2255
R13623 mux_magic_0.AND2_magic_0.A.n10 mux_magic_0.AND2_magic_0.A.n9 3.52811
R13624 mux_magic_0.AND2_magic_0.A.n7 mux_magic_0.AND2_magic_0.A.n4 3.30485
R13625 mux_magic_0.AND2_magic_0.A.n7 mux_magic_0.AND2_magic_0.A.n6 2.6005
R13626 mux_magic_0.AND2_magic_0.A.n4 mux_magic_0.AND2_magic_0.A.t3 1.6255
R13627 mux_magic_0.AND2_magic_0.A.n4 mux_magic_0.AND2_magic_0.A.n3 1.6255
R13628 mux_magic_0.AND2_magic_0.A.n6 mux_magic_0.AND2_magic_0.A.t4 1.6255
R13629 mux_magic_0.AND2_magic_0.A.n6 mux_magic_0.AND2_magic_0.A.n5 1.6255
R13630 mux_magic_0.AND2_magic_0.A.n9 mux_magic_0.AND2_magic_0.A.t2 1.463
R13631 mux_magic_0.AND2_magic_0.A.n9 mux_magic_0.AND2_magic_0.A.n8 1.463
R13632 mux_magic_0.AND2_magic_0.A.n11 mux_magic_0.AND2_magic_0.A.n10 0.8105
R13633 mux_magic_0.AND2_magic_0.A.n10 mux_magic_0.AND2_magic_0.A.n7 0.389848
R13634 mux_magic_0.AND2_magic_0.A.n13 mux_magic_0.AND2_magic_0.A.n11 0.389848
R13635 mux_magic_0.AND2_magic_0.A.n14 mux_magic_0.AND2_magic_0.A.n13 0.256804
R13636 mux_magic_0.AND2_magic_0.A mux_magic_0.AND2_magic_0.A.n14 0.173882
R13637 a_27922_11758.n3 a_27922_11758.n1 6.04375
R13638 a_27922_11758.n3 a_27922_11758.n2 1.55052
R13639 a_27922_11758.n1 a_27922_11758.t3 1.463
R13640 a_27922_11758.n1 a_27922_11758.n0 1.463
R13641 a_27922_11758.t0 a_27922_11758.n3 1.3335
R13642 a_27722_11758.t7 a_27722_11758.t8 44.058
R13643 a_27722_11758.n3 a_27722_11758.t6 34.6465
R13644 a_27722_11758.n3 a_27722_11758.t7 15.1219
R13645 a_27722_11758.n6 a_27722_11758.t0 5.29595
R13646 a_27722_11758.n4 a_27722_11758.n2 4.97104
R13647 a_27722_11758.n4 a_27722_11758.n3 4.16767
R13648 a_27722_11758.n5 a_27722_11758.n1 3.01333
R13649 a_27722_11758.n8 a_27722_11758.n6 3.01333
R13650 a_27722_11758.n1 a_27722_11758.t4 1.6255
R13651 a_27722_11758.n1 a_27722_11758.n0 1.6255
R13652 a_27722_11758.t3 a_27722_11758.n8 1.6255
R13653 a_27722_11758.n8 a_27722_11758.n7 1.6255
R13654 a_27722_11758.n6 a_27722_11758.n5 0.845717
R13655 a_27722_11758.n5 a_27722_11758.n4 0.423109
R13656 ITAIL.n7 ITAIL.t10 10.9054
R13657 ITAIL.n0 ITAIL.t17 10.8613
R13658 ITAIL.n17 ITAIL.t23 10.773
R13659 ITAIL.n13 ITAIL.t26 10.6003
R13660 ITAIL.n0 ITAIL.t0 10.5984
R13661 ITAIL.n17 ITAIL.t8 10.5336
R13662 ITAIL.n7 ITAIL.t18 10.5336
R13663 ITAIL.n1 ITAIL.t21 10.5334
R13664 ITAIL.n35 ITAIL.t22 10.533
R13665 ITAIL.n34 ITAIL.t4 10.5098
R13666 ITAIL.n18 ITAIL.t27 10.4686
R13667 ITAIL.n16 ITAIL.t12 10.0514
R13668 ITAIL.n10 ITAIL.t2 9.72546
R13669 ITAIL.n4 ITAIL.t6 9.65907
R13670 ITAIL.n36 ITAIL.t14 9.29485
R13671 ITAIL.n37 ITAIL.t19 8.47237
R13672 ITAIL.n29 ITAIL.t7 8.17686
R13673 ITAIL.n24 ITAIL.t13 8.07837
R13674 ITAIL.n25 ITAIL.n23 7.98962
R13675 ITAIL.n30 ITAIL.n28 7.84993
R13676 ITAIL.n29 ITAIL.t1 7.79699
R13677 ITAIL.n32 ITAIL.n26 7.73548
R13678 ITAIL.n24 ITAIL.t9 7.72811
R13679 ITAIL.n31 ITAIL.n27 7.58076
R13680 ITAIL.n39 ITAIL.n38 3.7682
R13681 ITAIL.n32 ITAIL.n31 1.75757
R13682 ITAIL.n20 ITAIL.n16 1.50725
R13683 ITAIL.n11 ITAIL.n10 1.50717
R13684 ITAIL.n6 ITAIL.n5 1.49748
R13685 ITAIL.n39 ITAIL 1.10761
R13686 ITAIL.n31 ITAIL.n30 0.661924
R13687 ITAIL.n14 ITAIL.n6 0.490305
R13688 ITAIL.n21 ITAIL.n14 0.446994
R13689 ITAIL.n37 ITAIL.n36 0.413008
R13690 ITAIL.n1 ITAIL.n0 0.390708
R13691 ITAIL.n36 ITAIL.n35 0.375243
R13692 ITAIL.n18 ITAIL.n17 0.365503
R13693 ITAIL.n19 ITAIL.n18 0.357915
R13694 ITAIL.n2 ITAIL.n1 0.357771
R13695 ITAIL.n13 ITAIL.n12 0.356995
R13696 ITAIL.n8 ITAIL.n7 0.341087
R13697 ITAIL.n33 ITAIL.n32 0.31096
R13698 ITAIL.n25 ITAIL.n24 0.301864
R13699 ITAIL.n30 ITAIL.n29 0.285711
R13700 ITAIL.n38 ITAIL.n22 0.278
R13701 ITAIL.n38 ITAIL.n37 0.244031
R13702 ITAIL.n33 ITAIL.n25 0.2255
R13703 ITAIL.n35 ITAIL.n34 0.201238
R13704 ITAIL.n34 ITAIL.n33 0.1493
R13705 ITAIL ITAIL.n39 0.0489615
R13706 ITAIL.n11 ITAIL.n8 0.028981
R13707 ITAIL.n14 ITAIL.n13 0.0236995
R13708 ITAIL.n21 ITAIL.n20 0.017375
R13709 ITAIL.n12 ITAIL.n11 0.0163348
R13710 ITAIL.n20 ITAIL.n19 0.0150187
R13711 ITAIL.n6 ITAIL.n3 0.013491
R13712 ITAIL.n3 ITAIL.n2 0.0117754
R13713 ITAIL.n22 ITAIL.n21 0.003875
R13714 ITAIL.n16 ITAIL.n15 0.00243623
R13715 ITAIL.n10 ITAIL.n9 0.00242648
R13716 ITAIL.n5 ITAIL.n4 0.00155882
R13717 mux_magic_0.OR_magic_0.A.t5 mux_magic_0.OR_magic_0.A.t3 44.6331
R13718 mux_magic_0.OR_magic_0.A.t7 mux_magic_0.OR_magic_0.A.t4 31.5469
R13719 mux_magic_0.OR_magic_0.A.t4 mux_magic_0.OR_magic_0.A.t6 28.6791
R13720 mux_magic_0.OR_magic_0.A.n0 mux_magic_0.OR_magic_0.A.t5 19.4237
R13721 mux_magic_0.OR_magic_0.A.n0 mux_magic_0.OR_magic_0.A.t7 12.1237
R13722 mux_magic_0.OR_magic_0.A mux_magic_0.OR_magic_0.A.n1 5.0317
R13723 mux_magic_0.OR_magic_0.A mux_magic_0.OR_magic_0.A.n0 4.23754
R13724 mux_magic_0.OR_magic_0.A mux_magic_0.OR_magic_0.A.n3 3.36245
R13725 mux_magic_0.OR_magic_0.A.n3 mux_magic_0.OR_magic_0.A.t1 1.6255
R13726 mux_magic_0.OR_magic_0.A.n3 mux_magic_0.OR_magic_0.A.n2 1.6255
R13727 a_29262_12133.n7 a_29262_12133.n0 5.71637
R13728 a_29262_12133.n6 a_29262_12133.t1 4.95333
R13729 a_29262_12133.n5 a_29262_12133.n4 3.54746
R13730 a_29262_12133.n5 a_29262_12133.n2 2.6005
R13731 a_29262_12133.n8 a_29262_12133.n7 2.6005
R13732 a_29262_12133.n2 a_29262_12133.t4 1.6255
R13733 a_29262_12133.n2 a_29262_12133.n1 1.6255
R13734 a_29262_12133.n4 a_29262_12133.t7 1.6255
R13735 a_29262_12133.n4 a_29262_12133.n3 1.6255
R13736 a_29262_12133.n8 a_29262_12133.t6 1.6255
R13737 a_29262_12133.n9 a_29262_12133.n8 1.6255
R13738 a_29262_12133.n7 a_29262_12133.n6 0.728326
R13739 a_29262_12133.n6 a_29262_12133.n5 0.552239
R13740 a_23836_10693.t2 a_23836_10693.n5 6.64563
R13741 a_23836_10693.n5 a_23836_10693.t3 6.61433
R13742 a_23836_10693.n4 a_23836_10693.n3 3.36963
R13743 a_23836_10693.n4 a_23836_10693.n1 3.33833
R13744 a_23836_10693.n3 a_23836_10693.t0 3.2765
R13745 a_23836_10693.n3 a_23836_10693.n2 3.2765
R13746 a_23836_10693.n1 a_23836_10693.t4 3.2765
R13747 a_23836_10693.n1 a_23836_10693.n0 3.2765
R13748 a_23836_10693.n5 a_23836_10693.n4 0.781777
R13749 a_45928_10426.t0 a_45928_10426.t1 12.9675
R13750 a_46228_9804.t0 a_46228_9804.t1 12.9675
R13751 a_44428_9598.t0 a_44428_9598.t1 12.9675
R13752 a_44128_8976.t0 a_44128_8976.t1 12.9675
R13753 a_42763_5679.n5 a_42763_5679.t9 29.2961
R13754 a_42763_5679.n6 a_42763_5679.n5 21.9292
R13755 a_42763_5679.n7 a_42763_5679.n6 18.1271
R13756 a_42763_5679.n7 a_42763_5679.t8 11.1695
R13757 a_42763_5679.n3 a_42763_5679.t0 10.2143
R13758 a_42763_5679.n5 a_42763_5679.t7 6.1325
R13759 a_42763_5679.n6 a_42763_5679.t6 6.1325
R13760 a_42763_5679.n3 a_42763_5679.n2 4.68517
R13761 a_42763_5679.n8 a_42763_5679.n7 4.6311
R13762 a_42763_5679.n10 a_42763_5679.n8 2.85093
R13763 a_42763_5679.n1 a_42763_5679.t2 2.16717
R13764 a_42763_5679.n1 a_42763_5679.n0 2.16717
R13765 a_42763_5679.t5 a_42763_5679.n10 2.16717
R13766 a_42763_5679.n10 a_42763_5679.n9 2.16717
R13767 a_42763_5679.n4 a_42763_5679.n3 1.58582
R13768 a_42763_5679.n4 a_42763_5679.n1 1.24371
R13769 a_42763_5679.n8 a_42763_5679.n4 0.971051
R13770 a_45928_8770.t0 a_45928_8770.t1 12.9675
R13771 a_45628_8148.t0 a_45628_8148.t1 12.9675
R13772 OUTB.n27 OUTB 6.6528
R13773 OUTB.n6 OUTB.n5 5.81586
R13774 OUTB.n2 OUTB.t15 5.10151
R13775 OUTB.n8 OUTB.t12 5.1005
R13776 OUTB.n7 OUTB.t17 5.08021
R13777 OUTB.n2 OUTB.n1 4.66164
R13778 OUTB.n13 OUTB.t11 3.6405
R13779 OUTB.n13 OUTB.n12 3.6405
R13780 OUTB.n15 OUTB.t7 3.6405
R13781 OUTB.n15 OUTB.n14 3.6405
R13782 OUTB.n20 OUTB.t4 3.6405
R13783 OUTB.n20 OUTB.n19 3.6405
R13784 OUTB.n22 OUTB.t10 3.6405
R13785 OUTB.n22 OUTB.n21 3.6405
R13786 OUTB.n25 OUTB.n11 3.50463
R13787 OUTB.n24 OUTB.n18 3.50463
R13788 OUTB.n11 OUTB.t2 3.2765
R13789 OUTB.n11 OUTB.n10 3.2765
R13790 OUTB.n18 OUTB.t3 3.2765
R13791 OUTB.n18 OUTB.n17 3.2765
R13792 OUTB.n16 OUTB.n15 3.06224
R13793 OUTB.n23 OUTB.n22 3.06224
R13794 OUTB.n6 OUTB.n4 2.85093
R13795 OUTB.n16 OUTB.n13 2.6005
R13796 OUTB.n23 OUTB.n20 2.6005
R13797 OUTB.n4 OUTB.t18 2.16717
R13798 OUTB.n4 OUTB.n3 2.16717
R13799 OUTB.n1 OUTB.t14 1.9505
R13800 OUTB.n1 OUTB.n0 1.9505
R13801 OUTB.n27 OUTB.n26 1.47848
R13802 OUTB OUTB.n27 1.06887
R13803 OUTB.n25 OUTB.n24 0.798761
R13804 OUTB.n7 OUTB.n6 0.644196
R13805 OUTB OUTB.n25 0.562022
R13806 OUTB.n8 OUTB.n7 0.447229
R13807 OUTB.n9 OUTB.n2 0.308586
R13808 OUTB.n9 OUTB.n8 0.277162
R13809 OUTB.n25 OUTB.n16 0.18637
R13810 OUTB.n24 OUTB.n23 0.18637
R13811 OUTB.n26 OUTB 0.161224
R13812 OUTB OUTB.n9 0.115935
R13813 OUTB.n26 OUTB 0.0483126
R13814 a_42628_8770.t0 a_42628_8770.t1 10.2205
R13815 a_42628_8148.t0 a_42628_8148.t1 12.9675
R13816 a_31732_10267.n13 a_31732_10267.n12 10.0413
R13817 a_31732_10267.n5 a_31732_10267.t5 8.81226
R13818 a_31732_10267.n12 a_31732_10267.n0 8.80202
R13819 a_31732_10267.n4 a_31732_10267.t3 8.78441
R13820 a_31732_10267.n10 a_31732_10267.t1 8.6005
R13821 a_31732_10267.n8 a_31732_10267.n6 8.15323
R13822 a_31732_10267.n8 a_31732_10267.n7 8.13693
R13823 a_31732_10267.n9 a_31732_10267.t6 8.0091
R13824 a_31732_10267.n1 a_31732_10267.t8 5.72901
R13825 a_31732_10267.n1 a_31732_10267.t11 5.2005
R13826 a_31732_10267.n2 a_31732_10267.t10 5.2005
R13827 a_31732_10267.n3 a_31732_10267.t9 5.2005
R13828 a_31732_10267.n10 a_31732_10267.n9 2.91981
R13829 a_31732_10267.n12 a_31732_10267.n11 2.34763
R13830 a_31732_10267.n11 a_31732_10267.n5 2.1305
R13831 a_31732_10267.n4 a_31732_10267.n3 1.88322
R13832 a_31732_10267.n5 a_31732_10267.n4 1.10344
R13833 a_31732_10267.n2 a_31732_10267.n1 0.529011
R13834 a_31732_10267.n3 a_31732_10267.n2 0.529011
R13835 a_31732_10267.n11 a_31732_10267.n10 0.294424
R13836 a_31732_10267.n9 a_31732_10267.n8 0.219455
R13837 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n20 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t23 23.6945
R13838 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t21 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n21 23.6945
R13839 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n21 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n20 18.8035
R13840 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n18 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n16 15.8172
R13841 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n18 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n17 15.8172
R13842 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n17 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n13 15.8172
R13843 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n16 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t30 14.8925
R13844 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t22 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n18 14.8925
R13845 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n17 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t20 14.8925
R13846 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n22 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n14 12.2457
R13847 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n19 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n14 12.2457
R13848 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n19 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n15 12.2457
R13849 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n23 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t26 11.6285
R13850 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n15 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t23 8.9065
R13851 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t31 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n19 8.9065
R13852 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t28 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n14 8.9065
R13853 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n22 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t21 8.9065
R13854 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n18 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t25 8.6145
R13855 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n16 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t24 8.6145
R13856 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n17 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t27 8.6145
R13857 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n13 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t29 8.59715
R13858 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t30 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n15 8.3225
R13859 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n19 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t22 8.3225
R13860 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t20 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n14 8.3225
R13861 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t26 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n22 8.3225
R13862 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n24 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n12 5.24044
R13863 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n7 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n4 5.10151
R13864 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n9 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n3 5.10119
R13865 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n10 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n2 5.08021
R13866 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n7 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n6 4.66164
R13867 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n23 4.223
R13868 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n20 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t31 3.6505
R13869 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n21 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t28 3.6505
R13870 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n37 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t12 3.6405
R13871 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n37 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n36 3.6405
R13872 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n28 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t9 3.6405
R13873 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n28 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n27 3.6405
R13874 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n26 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t8 3.6405
R13875 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n26 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n25 3.6405
R13876 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n35 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t11 3.6405
R13877 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n35 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n34 3.6405
R13878 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n39 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n33 3.50463
R13879 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n40 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n31 3.50463
R13880 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n12 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t18 3.40711
R13881 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n33 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t6 3.2765
R13882 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n33 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n32 3.2765
R13883 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n31 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t4 3.2765
R13884 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n31 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n30 3.2765
R13885 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n23 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n13 3.1807
R13886 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n29 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n26 3.06224
R13887 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n38 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n35 3.06224
R13888 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n11 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n1 2.85093
R13889 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n29 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n28 2.6005
R13890 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n38 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n37 2.6005
R13891 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n8 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT 2.36593
R13892 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n1 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t17 2.16717
R13893 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n1 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n0 2.16717
R13894 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n24 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT 2.01183
R13895 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n6 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t3 1.9505
R13896 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n6 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n5 1.9505
R13897 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n12 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n11 1.0205
R13898 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n40 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n39 0.798761
R13899 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n11 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n10 0.644196
R13900 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n40 0.562022
R13901 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n10 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n9 0.450799
R13902 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n8 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n7 0.358456
R13903 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n24 0.278326
R13904 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n9 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n8 0.229792
R13905 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n40 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n29 0.18637
R13906 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n39 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n38 0.18637
R13907 PFD_T2_0.FDIV.n1 PFD_T2_0.FDIV.n0 13.9524
R13908 PFD_T2_0.FDIV.n0 PFD_T2_0.FDIV.t4 12.4105
R13909 PFD_T2_0.FDIV.n0 PFD_T2_0.FDIV.t6 11.5345
R13910 PFD_T2_0.FDIV PFD_T2_0.FDIV.n1 8.49358
R13911 PFD_T2_0.FDIV.n1 PFD_T2_0.FDIV.t3 8.1035
R13912 PFD_T2_0.FDIV.n1 PFD_T2_0.FDIV.t5 7.6655
R13913 PFD_T2_0.FDIV.n5 PFD_T2_0.FDIV.n3 5.47387
R13914 PFD_T2_0.FDIV.n6 PFD_T2_0.FDIV.n2 4.65398
R13915 PFD_T2_0.FDIV.n5 PFD_T2_0.FDIV.n4 4.2255
R13916 PFD_T2_0.FDIV.n6 PFD_T2_0.FDIV.n5 0.427022
R13917 PFD_T2_0.FDIV PFD_T2_0.FDIV.n6 0.421777
R13918 a_24436_11277.n1 a_24436_11277.t0 7.21081
R13919 a_24436_11277.n1 a_24436_11277.n0 7.15165
R13920 a_24436_11277.n2 a_24436_11277.t2 3.6405
R13921 a_24436_11277.n3 a_24436_11277.n2 3.6405
R13922 a_24436_11277.n2 a_24436_11277.n1 2.77149
R13923 a_45158_5339.n0 a_45158_5339.t8 29.2961
R13924 a_45158_5339.n1 a_45158_5339.n0 21.9292
R13925 a_45158_5339.n2 a_45158_5339.n1 18.1271
R13926 a_45158_5339.n2 a_45158_5339.t6 11.1695
R13927 a_45158_5339.n0 a_45158_5339.t7 6.1325
R13928 a_45158_5339.n1 a_45158_5339.t9 6.1325
R13929 a_45158_5339.n6 a_45158_5339.n5 4.93252
R13930 a_45158_5339.n6 a_45158_5339.t0 4.70348
R13931 a_45158_5339.n8 a_45158_5339.n2 4.6311
R13932 a_45158_5339.n10 a_45158_5339.n8 2.85093
R13933 a_45158_5339.n4 a_45158_5339.t4 2.16717
R13934 a_45158_5339.n4 a_45158_5339.n3 2.16717
R13935 a_45158_5339.t5 a_45158_5339.n10 2.16717
R13936 a_45158_5339.n10 a_45158_5339.n9 2.16717
R13937 a_45158_5339.n7 a_45158_5339.n6 1.58582
R13938 a_45158_5339.n7 a_45158_5339.n4 1.24371
R13939 a_45158_5339.n8 a_45158_5339.n7 0.971051
R13940 mux_magic_0.OR_magic_0.B.t6 mux_magic_0.OR_magic_0.B.t5 44.6331
R13941 mux_magic_0.OR_magic_0.B.t4 mux_magic_0.OR_magic_0.B.t6 43.4094
R13942 mux_magic_0.OR_magic_0.B.t7 mux_magic_0.OR_magic_0.B.t4 31.5469
R13943 mux_magic_0.OR_magic_0.B.n0 mux_magic_0.OR_magic_0.B.t7 15.0567
R13944 mux_magic_0.OR_magic_0.B.n0 mux_magic_0.OR_magic_0.B.t3 13.6228
R13945 mux_magic_0.OR_magic_0.B mux_magic_0.OR_magic_0.B.n1 5.03757
R13946 mux_magic_0.OR_magic_0.B mux_magic_0.OR_magic_0.B.n0 4.2675
R13947 mux_magic_0.OR_magic_0.B mux_magic_0.OR_magic_0.B.n3 3.36521
R13948 mux_magic_0.OR_magic_0.B.n3 mux_magic_0.OR_magic_0.B.t2 1.6255
R13949 mux_magic_0.OR_magic_0.B.n3 mux_magic_0.OR_magic_0.B.n2 1.6255
R13950 a_45328_12082.t0 a_45328_12082.t1 12.9675
R13951 a_45628_11460.t0 a_45628_11460.t1 12.9675
R13952 a_44128_8770.t0 a_44128_8770.t1 12.9675
R13953 a_43828_8148.t0 a_43828_8148.t1 12.9675
R13954 a_31468_10271.t8 a_31468_10271.t7 17.9898
R13955 a_31468_10271.t9 a_31468_10271.t8 17.9898
R13956 a_31468_10271.t6 a_31468_10271.t9 17.9898
R13957 a_31468_10271.n1 a_31468_10271.t6 13.0554
R13958 a_31468_10271.n0 a_31468_10271.n5 8.89703
R13959 a_31468_10271.n1 a_31468_10271.n2 8.71168
R13960 a_31468_10271.n0 a_31468_10271.n6 8.60182
R13961 a_31468_10271.n0 a_31468_10271.n3 8.6005
R13962 a_31468_10271.n7 a_31468_10271.n1 8.6005
R13963 a_31468_10271.n0 a_31468_10271.n4 8.5505
R13964 a_31468_10271.n1 a_31468_10271.n0 2.08339
R13965 DN.t7 DN.t5 12.5148
R13966 DN.n3 DN.t7 10.2564
R13967 DN.n0 DN.t4 10.1117
R13968 DN.n1 DN.t6 9.54068
R13969 DN.n2 DN.t8 9.4755
R13970 DN.n0 DN.t3 9.4755
R13971 DN.n7 DN.n5 5.47387
R13972 DN.n9 DN.n8 4.65398
R13973 DN.n7 DN.n6 4.2255
R13974 DN.n4 DN 1.15322
R13975 DN.n4 DN 0.960106
R13976 DN.n2 DN.n1 0.50481
R13977 DN.n1 DN.n0 0.501707
R13978 DN.n9 DN.n7 0.427022
R13979 DN.n3 DN.n2 0.332569
R13980 DN DN.n9 0.257096
R13981 DN DN.n3 0.2505
R13982 DN DN.n4 0.0373182
R13983 a_45628_11254.t0 a_45628_11254.t1 12.9675
R13984 a_45328_10632.t0 a_45328_10632.t1 12.9675
R13985 F_IN.t3 F_IN.t1 44.058
R13986 F_IN.n0 F_IN.t0 38.8649
R13987 F_IN.t0 F_IN.t3 28.6791
R13988 F_IN.n0 F_IN.t2 7.3005
R13989 F_IN F_IN.n0 5.27587
R13990 F_IN.n1 F_IN 2.72439
R13991 F_IN.n1 F_IN 1.4172
R13992 F_IN F_IN.n1 0.00465837
R13993 a_20097_10547.n2 a_20097_10547.n1 6.04407
R13994 a_20097_10547.n1 a_20097_10547.n0 1.55018
R13995 a_20097_10547.n2 a_20097_10547.t2 1.463
R13996 a_20097_10547.n3 a_20097_10547.n2 1.463
R13997 a_20097_10547.n1 a_20097_10547.t0 1.33387
R13998 a_22880_10947.n3 a_22880_10947.n2 6.53021
R13999 a_22880_10947.n2 a_22880_10947.t2 6.47121
R14000 a_22880_10947.n1 a_22880_10947.t0 3.35758
R14001 a_22880_10947.n1 a_22880_10947.n0 3.01392
R14002 a_22880_10947.n2 a_22880_10947.n1 2.46725
R14003 a_19903_8443.t6 a_19903_8443.t7 44.058
R14004 a_19903_8443.n3 a_19903_8443.t8 34.6465
R14005 a_19903_8443.n3 a_19903_8443.t6 15.1219
R14006 a_19903_8443.n6 a_19903_8443.t3 5.29595
R14007 a_19903_8443.n4 a_19903_8443.n2 4.97104
R14008 a_19903_8443.n4 a_19903_8443.n3 4.16767
R14009 a_19903_8443.n5 a_19903_8443.n1 3.01333
R14010 a_19903_8443.n8 a_19903_8443.n6 3.01333
R14011 a_19903_8443.n1 a_19903_8443.t5 1.6255
R14012 a_19903_8443.n1 a_19903_8443.n0 1.6255
R14013 a_19903_8443.t1 a_19903_8443.n8 1.6255
R14014 a_19903_8443.n8 a_19903_8443.n7 1.6255
R14015 a_19903_8443.n6 a_19903_8443.n5 0.845717
R14016 a_19903_8443.n5 a_19903_8443.n4 0.423109
R14017 mux_magic_3.OR_magic_0.B.t6 mux_magic_3.OR_magic_0.B.t7 44.6331
R14018 mux_magic_3.OR_magic_0.B.t5 mux_magic_3.OR_magic_0.B.t6 43.4094
R14019 mux_magic_3.OR_magic_0.B.t3 mux_magic_3.OR_magic_0.B.t5 31.5469
R14020 mux_magic_3.OR_magic_0.B.n0 mux_magic_3.OR_magic_0.B.t3 15.0567
R14021 mux_magic_3.OR_magic_0.B.n0 mux_magic_3.OR_magic_0.B.t4 13.6228
R14022 mux_magic_3.OR_magic_0.B mux_magic_3.OR_magic_0.B.n1 5.03757
R14023 mux_magic_3.OR_magic_0.B mux_magic_3.OR_magic_0.B.n0 4.2675
R14024 mux_magic_3.OR_magic_0.B mux_magic_3.OR_magic_0.B.n3 3.36521
R14025 mux_magic_3.OR_magic_0.B.n3 mux_magic_3.OR_magic_0.B.t1 1.6255
R14026 mux_magic_3.OR_magic_0.B.n3 mux_magic_3.OR_magic_0.B.n2 1.6255
R14027 mux_magic_2.OR_magic_0.A.t3 mux_magic_2.OR_magic_0.A.t6 44.6331
R14028 mux_magic_2.OR_magic_0.A.t5 mux_magic_2.OR_magic_0.A.t7 31.5469
R14029 mux_magic_2.OR_magic_0.A.t7 mux_magic_2.OR_magic_0.A.t4 28.6791
R14030 mux_magic_2.OR_magic_0.A.n0 mux_magic_2.OR_magic_0.A.t3 19.4237
R14031 mux_magic_2.OR_magic_0.A.n0 mux_magic_2.OR_magic_0.A.t5 12.1237
R14032 mux_magic_2.OR_magic_0.A mux_magic_2.OR_magic_0.A.n1 5.0317
R14033 mux_magic_2.OR_magic_0.A mux_magic_2.OR_magic_0.A.n0 4.23754
R14034 mux_magic_2.OR_magic_0.A mux_magic_2.OR_magic_0.A.n3 3.36245
R14035 mux_magic_2.OR_magic_0.A.n3 mux_magic_2.OR_magic_0.A.t1 1.6255
R14036 mux_magic_2.OR_magic_0.A.n3 mux_magic_2.OR_magic_0.A.n2 1.6255
R14037 a_21437_12116.n3 a_21437_12116.n0 5.71637
R14038 a_21437_12116.n4 a_21437_12116.t7 4.95333
R14039 a_21437_12116.n7 a_21437_12116.n6 3.54746
R14040 a_21437_12116.n3 a_21437_12116.n2 2.6005
R14041 a_21437_12116.n9 a_21437_12116.n7 2.6005
R14042 a_21437_12116.n6 a_21437_12116.t1 1.6255
R14043 a_21437_12116.n6 a_21437_12116.n5 1.6255
R14044 a_21437_12116.n2 a_21437_12116.t2 1.6255
R14045 a_21437_12116.n2 a_21437_12116.n1 1.6255
R14046 a_21437_12116.t3 a_21437_12116.n9 1.6255
R14047 a_21437_12116.n9 a_21437_12116.n8 1.6255
R14048 a_21437_12116.n4 a_21437_12116.n3 0.728326
R14049 a_21437_12116.n7 a_21437_12116.n4 0.552239
R14050 a_29262_10725.t6 a_29262_10725.t8 31.5469
R14051 a_29262_10725.n5 a_29262_10725.t6 13.2715
R14052 a_29262_10725.n5 a_29262_10725.t7 13.0934
R14053 a_29262_10725.n4 a_29262_10725.t0 6.52735
R14054 a_29262_10725.n6 a_29262_10725.n5 4.33404
R14055 a_29262_10725.n7 a_29262_10725.n2 4.2255
R14056 a_29262_10725.n9 a_29262_10725.n8 4.2255
R14057 a_29262_10725.n8 a_29262_10725.n1 3.81956
R14058 a_29262_10725.n4 a_29262_10725.n3 2.62633
R14059 a_29262_10725.n1 a_29262_10725.t4 1.6255
R14060 a_29262_10725.n1 a_29262_10725.n0 1.6255
R14061 a_29262_10725.n8 a_29262_10725.n7 0.947457
R14062 a_29262_10725.n7 a_29262_10725.n6 0.368326
R14063 a_29262_10725.n6 a_29262_10725.n4 0.234808
R14064 a_22881_9554.n1 a_22881_9554.n0 6.53012
R14065 a_22881_9554.n1 a_22881_9554.t3 6.47102
R14066 a_22881_9554.t1 a_22881_9554.n3 3.35684
R14067 a_22881_9554.n3 a_22881_9554.n2 3.01376
R14068 a_22881_9554.n3 a_22881_9554.n1 2.46742
R14069 PFD_T2_0.DOWN.t6 PFD_T2_0.DOWN.t5 44.058
R14070 PFD_T2_0.DOWN.n0 PFD_T2_0.DOWN.t3 38.8649
R14071 PFD_T2_0.DOWN.t3 PFD_T2_0.DOWN.t6 28.6791
R14072 PFD_T2_0.DOWN.n0 PFD_T2_0.DOWN.t4 7.3005
R14073 PFD_T2_0.DOWN.n4 PFD_T2_0.DOWN.n1 6.76498
R14074 PFD_T2_0.DOWN PFD_T2_0.DOWN.n0 5.38424
R14075 PFD_T2_0.DOWN.n3 PFD_T2_0.DOWN.t2 3.6405
R14076 PFD_T2_0.DOWN.n3 PFD_T2_0.DOWN.n2 3.6405
R14077 PFD_T2_0.DOWN.n4 PFD_T2_0.DOWN.n3 2.78441
R14078 PFD_T2_0.DOWN PFD_T2_0.DOWN.n4 0.471261
R14079 a_42628_11460.t0 a_42628_11460.t1 12.9675
R14080 a_46528_12082.t0 a_46528_12082.t1 12.9675
R14081 a_46228_11460.t0 a_46228_11460.t1 12.9675
R14082 a_19903_9637.t6 a_19903_9637.t7 44.058
R14083 a_19903_9637.n1 a_19903_9637.t8 34.6465
R14084 a_19903_9637.n1 a_19903_9637.t6 15.1219
R14085 a_19903_9637.n5 a_19903_9637.t5 5.29595
R14086 a_19903_9637.n2 a_19903_9637.n0 4.97104
R14087 a_19903_9637.n2 a_19903_9637.n1 4.16767
R14088 a_19903_9637.n5 a_19903_9637.n4 3.01333
R14089 a_19903_9637.n8 a_19903_9637.n6 3.01333
R14090 a_19903_9637.n4 a_19903_9637.t2 1.6255
R14091 a_19903_9637.n4 a_19903_9637.n3 1.6255
R14092 a_19903_9637.t1 a_19903_9637.n8 1.6255
R14093 a_19903_9637.n8 a_19903_9637.n7 1.6255
R14094 a_19903_9637.n6 a_19903_9637.n5 0.845717
R14095 a_19903_9637.n6 a_19903_9637.n2 0.423109
R14096 a_45328_10426.t0 a_45328_10426.t1 12.9675
R14097 a_45628_9804.t0 a_45628_9804.t1 12.9675
R14098 PFD_T2_0.Buffer_V_2_1.IN.n3 PFD_T2_0.Buffer_V_2_1.IN.t13 13.1405
R14099 PFD_T2_0.Buffer_V_2_1.IN.n4 PFD_T2_0.Buffer_V_2_1.IN.n3 12.4464
R14100 PFD_T2_0.Buffer_V_2_1.IN.n3 PFD_T2_0.Buffer_V_2_1.IN.t12 9.9285
R14101 PFD_T2_0.Buffer_V_2_1.IN.n22 PFD_T2_0.Buffer_V_2_1.IN.t11 9.7095
R14102 PFD_T2_0.Buffer_V_2_1.IN.n19 PFD_T2_0.Buffer_V_2_1.IN.n18 6.60246
R14103 PFD_T2_0.Buffer_V_2_1.IN.n1 PFD_T2_0.Buffer_V_2_1.IN.n5 4.5005
R14104 PFD_T2_0.Buffer_V_2_1.IN.n1 PFD_T2_0.Buffer_V_2_1.IN.n23 4.25602
R14105 PFD_T2_0.Buffer_V_2_1.IN.n1 PFD_T2_0.Buffer_V_2_1.IN.n2 4.22422
R14106 PFD_T2_0.Buffer_V_2_1.IN.n11 PFD_T2_0.Buffer_V_2_1.IN.t3 3.6405
R14107 PFD_T2_0.Buffer_V_2_1.IN.n11 PFD_T2_0.Buffer_V_2_1.IN.n10 3.6405
R14108 PFD_T2_0.Buffer_V_2_1.IN.n13 PFD_T2_0.Buffer_V_2_1.IN.t4 3.6405
R14109 PFD_T2_0.Buffer_V_2_1.IN.n13 PFD_T2_0.Buffer_V_2_1.IN.n12 3.6405
R14110 PFD_T2_0.Buffer_V_2_1.IN.n14 PFD_T2_0.Buffer_V_2_1.IN.n13 3.54941
R14111 PFD_T2_0.Buffer_V_2_1.IN.n17 PFD_T2_0.Buffer_V_2_1.IN.n16 3.33833
R14112 PFD_T2_0.Buffer_V_2_1.IN.n20 PFD_T2_0.Buffer_V_2_1.IN.n9 3.33833
R14113 PFD_T2_0.Buffer_V_2_1.IN.n16 PFD_T2_0.Buffer_V_2_1.IN.t8 3.2765
R14114 PFD_T2_0.Buffer_V_2_1.IN.n16 PFD_T2_0.Buffer_V_2_1.IN.n15 3.2765
R14115 PFD_T2_0.Buffer_V_2_1.IN.n9 PFD_T2_0.Buffer_V_2_1.IN.t0 3.2765
R14116 PFD_T2_0.Buffer_V_2_1.IN.n9 PFD_T2_0.Buffer_V_2_1.IN.n8 3.2765
R14117 PFD_T2_0.Buffer_V_2_1.IN.n0 PFD_T2_0.Buffer_V_2_1.IN.t1 3.2238
R14118 PFD_T2_0.Buffer_V_2_1.IN.n14 PFD_T2_0.Buffer_V_2_1.IN.n11 2.78441
R14119 PFD_T2_0.Buffer_V_2_1.IN.n7 PFD_T2_0.Buffer_V_2_1.IN.n6 1.9535
R14120 PFD_T2_0.Buffer_V_2_1.IN.n2 PFD_T2_0.Buffer_V_2_1.IN.n0 1.82827
R14121 PFD_T2_0.Buffer_V_2_1.IN.n0 PFD_T2_0.Buffer_V_2_1.IN.n7 1.37516
R14122 PFD_T2_0.Buffer_V_2_1.IN.n2 PFD_T2_0.Buffer_V_2_1.IN.n20 0.891537
R14123 PFD_T2_0.Buffer_V_2_1.IN.n23 PFD_T2_0.Buffer_V_2_1.IN.n21 0.729844
R14124 PFD_T2_0.Buffer_V_2_1.IN.n23 PFD_T2_0.Buffer_V_2_1.IN.n22 0.587069
R14125 PFD_T2_0.Buffer_V_2_1.IN.n19 PFD_T2_0.Buffer_V_2_1.IN.n17 0.524848
R14126 PFD_T2_0.Buffer_V_2_1.IN.n5 PFD_T2_0.Buffer_V_2_1.IN.n4 0.5115
R14127 PFD_T2_0.Buffer_V_2_1.IN.n17 PFD_T2_0.Buffer_V_2_1.IN.n14 0.358543
R14128 PFD_T2_0.Buffer_V_2_1.IN.n20 PFD_T2_0.Buffer_V_2_1.IN.n19 0.274413
R14129 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.Buffer_V_2_1.IN.n1 0.271564
R14130 a_43828_9598.t0 a_43828_9598.t1 12.9675
R14131 a_43528_8976.t0 a_43528_8976.t1 12.9675
R14132 VCTRL_IN.n3 VCTRL_IN.n2 5.81586
R14133 VCTRL_IN.n5 VCTRL_IN.t3 5.10208
R14134 VCTRL_IN.n8 VCTRL_IN.t1 5.10194
R14135 VCTRL_IN.n4 VCTRL_IN.t5 5.08021
R14136 VCTRL_IN.n8 VCTRL_IN.n7 4.66114
R14137 VCTRL_IN.n3 VCTRL_IN.n1 2.85093
R14138 VCTRL_IN.n1 VCTRL_IN.t6 2.16717
R14139 VCTRL_IN.n1 VCTRL_IN.n0 2.16717
R14140 VCTRL_IN.n7 VCTRL_IN.t0 1.9505
R14141 VCTRL_IN.n7 VCTRL_IN.n6 1.9505
R14142 VCTRL_IN.n4 VCTRL_IN.n3 0.644196
R14143 VCTRL_IN.n5 VCTRL_IN.n4 0.449473
R14144 VCTRL_IN.n9 VCTRL_IN.n8 0.21214
R14145 VCTRL_IN.n9 VCTRL_IN.n5 0.198571
R14146 VCTRL_IN VCTRL_IN.n9 0.0718949
R14147 a_42628_11254.t0 a_42628_11254.t1 12.9675
R14148 a_42628_10426.t0 a_42628_10426.t1 10.2205
R14149 a_46228_11254.t0 a_46228_11254.t1 12.9675
R14150 a_46528_10632.t0 a_46528_10632.t1 12.9675
R14151 mux_magic_1.OR_magic_0.A.t3 mux_magic_1.OR_magic_0.A.t6 44.6331
R14152 mux_magic_1.OR_magic_0.A.t5 mux_magic_1.OR_magic_0.A.t4 31.5469
R14153 mux_magic_1.OR_magic_0.A.t4 mux_magic_1.OR_magic_0.A.t7 28.6791
R14154 mux_magic_1.OR_magic_0.A.n0 mux_magic_1.OR_magic_0.A.t3 19.3585
R14155 mux_magic_1.OR_magic_0.A.n0 mux_magic_1.OR_magic_0.A.t5 12.1889
R14156 mux_magic_1.OR_magic_0.A mux_magic_1.OR_magic_0.A.n1 5.0317
R14157 mux_magic_1.OR_magic_0.A mux_magic_1.OR_magic_0.A.n0 4.23754
R14158 mux_magic_1.OR_magic_0.A mux_magic_1.OR_magic_0.A.n3 3.36245
R14159 mux_magic_1.OR_magic_0.A.n3 mux_magic_1.OR_magic_0.A.t1 1.6255
R14160 mux_magic_1.OR_magic_0.A.n3 mux_magic_1.OR_magic_0.A.n2 1.6255
R14161 a_23837_9553.n2 a_23837_9553.t0 6.64563
R14162 a_23837_9553.n2 a_23837_9553.t4 6.61433
R14163 a_23837_9553.n5 a_23837_9553.n3 3.36963
R14164 a_23837_9553.n3 a_23837_9553.n1 3.33833
R14165 a_23837_9553.n1 a_23837_9553.t3 3.2765
R14166 a_23837_9553.n1 a_23837_9553.n0 3.2765
R14167 a_23837_9553.t2 a_23837_9553.n5 3.2765
R14168 a_23837_9553.n5 a_23837_9553.n4 3.2765
R14169 a_23837_9553.n3 a_23837_9553.n2 0.781777
R14170 a_45028_9598.t0 a_45028_9598.t1 12.9675
R14171 a_45328_8976.t0 a_45328_8976.t1 12.9675
R14172 a_28075_8520.n2 a_28075_8520.n1 6.04392
R14173 a_28075_8520.n3 a_28075_8520.n2 1.55019
R14174 a_28075_8520.n1 a_28075_8520.t0 1.463
R14175 a_28075_8520.n1 a_28075_8520.n0 1.463
R14176 a_28075_8520.n2 a_28075_8520.t2 1.33386
R14177 a_46528_8770.t0 a_46528_8770.t1 12.9675
R14178 a_43528_8770.t0 a_43528_8770.t1 12.9675
R14179 a_28075_9714.n2 a_28075_9714.n1 6.04536
R14180 a_28075_9714.n1 a_28075_9714.n0 1.5502
R14181 a_28075_9714.n2 a_28075_9714.t2 1.463
R14182 a_28075_9714.n3 a_28075_9714.n2 1.463
R14183 a_28075_9714.n1 a_28075_9714.t0 1.33385
R14184 a_44716_1837.n3 a_44716_1837.t8 29.3691
R14185 a_44716_1837.n4 a_44716_1837.n3 21.9292
R14186 a_44716_1837.n5 a_44716_1837.n4 18.1271
R14187 a_44716_1837.n5 a_44716_1837.t9 11.2425
R14188 a_44716_1837.n8 a_44716_1837.n7 10.1038
R14189 a_44716_1837.n3 a_44716_1837.t6 6.1325
R14190 a_44716_1837.n4 a_44716_1837.t7 6.1325
R14191 a_44716_1837.n8 a_44716_1837.t0 4.70149
R14192 a_44716_1837.n6 a_44716_1837.n5 4.6302
R14193 a_44716_1837.n6 a_44716_1837.n2 2.85093
R14194 a_44716_1837.n2 a_44716_1837.t2 2.16717
R14195 a_44716_1837.n2 a_44716_1837.n1 2.16717
R14196 a_44716_1837.t5 a_44716_1837.n10 2.16717
R14197 a_44716_1837.n10 a_44716_1837.n0 2.16717
R14198 a_44716_1837.n9 a_44716_1837.n8 1.58618
R14199 a_44716_1837.n10 a_44716_1837.n9 1.24388
R14200 a_44716_1837.n9 a_44716_1837.n6 0.97169
R14201 a_43228_11460.t0 a_43228_11460.t1 12.9675
R14202 a_41879_n196.n5 a_41879_n196.t8 29.2961
R14203 a_41879_n196.n6 a_41879_n196.n5 21.9292
R14204 a_41879_n196.n7 a_41879_n196.n6 18.1271
R14205 a_41879_n196.n7 a_41879_n196.t6 11.1695
R14206 a_41879_n196.n3 a_41879_n196.t0 10.2143
R14207 a_41879_n196.n5 a_41879_n196.t9 6.1325
R14208 a_41879_n196.n6 a_41879_n196.t7 6.1325
R14209 a_41879_n196.n3 a_41879_n196.n2 4.68517
R14210 a_41879_n196.n8 a_41879_n196.n7 4.6311
R14211 a_41879_n196.n10 a_41879_n196.n8 2.85093
R14212 a_41879_n196.n1 a_41879_n196.t2 2.16717
R14213 a_41879_n196.n1 a_41879_n196.n0 2.16717
R14214 a_41879_n196.t5 a_41879_n196.n10 2.16717
R14215 a_41879_n196.n10 a_41879_n196.n9 2.16717
R14216 a_41879_n196.n4 a_41879_n196.n3 1.58582
R14217 a_41879_n196.n4 a_41879_n196.n1 1.24371
R14218 a_41879_n196.n8 a_41879_n196.n4 0.971051
R14219 a_43228_11254.t0 a_43228_11254.t1 12.9675
R14220 a_44728_8770.t0 a_44728_8770.t1 12.9675
R14221 a_45028_8148.t0 a_45028_8148.t1 12.9675
R14222 UP_INPUT.t2 UP_INPUT.t1 44.058
R14223 UP_INPUT.n0 UP_INPUT.t0 38.8649
R14224 UP_INPUT.t0 UP_INPUT.t2 28.6791
R14225 UP_INPUT.n0 UP_INPUT.t3 7.3005
R14226 UP_INPUT UP_INPUT.n0 5.27587
R14227 PFD_T2_0.UP.t6 PFD_T2_0.UP.t4 44.058
R14228 PFD_T2_0.UP.n0 PFD_T2_0.UP.t3 38.8649
R14229 PFD_T2_0.UP.t3 PFD_T2_0.UP.t6 28.6791
R14230 PFD_T2_0.UP.n0 PFD_T2_0.UP.t5 7.3005
R14231 PFD_T2_0.UP PFD_T2_0.UP.n1 6.76498
R14232 PFD_T2_0.UP PFD_T2_0.UP.n0 5.27587
R14233 PFD_T2_0.UP.n3 PFD_T2_0.UP.t2 3.6405
R14234 PFD_T2_0.UP.n3 PFD_T2_0.UP.n2 3.6405
R14235 PFD_T2_0.UP PFD_T2_0.UP.n3 2.78441
R14236 a_44128_12082.t0 a_44128_12082.t1 12.9675
R14237 a_25556_11637.n0 a_25556_11637.t5 24.1814
R14238 a_25556_11637.n1 a_25556_11637.t4 12.4835
R14239 a_25556_11637.n0 a_25556_11637.t3 8.6875
R14240 a_25556_11637.n2 a_25556_11637.t0 6.71215
R14241 a_25556_11637.n2 a_25556_11637.n1 4.46748
R14242 a_25556_11637.n3 a_25556_11637.t1 3.6405
R14243 a_25556_11637.n4 a_25556_11637.n3 3.6405
R14244 a_25556_11637.n3 a_25556_11637.n2 2.83724
R14245 a_25556_11637.n1 a_25556_11637.n0 1.8985
R14246 a_44128_10632.t0 a_44128_10632.t1 12.9675
R14247 a_46528_10426.t0 a_46528_10426.t1 12.9675
R14248 a_42928_10426.t0 a_42928_10426.t1 12.9675
R14249 a_43228_9804.t0 a_43228_9804.t1 12.9675
R14250 a_44728_8976.t0 a_44728_8976.t1 12.9675
R14251 a_46228_9598.t0 a_46228_9598.t1 12.9675
R14252 a_45928_8976.t0 a_45928_8976.t1 12.9675
R14253 a_45028_11460.t0 a_45028_11460.t1 12.9675
R14254 a_44428_8148.t0 a_44428_8148.t1 12.9675
R14255 a_45028_11254.t0 a_45028_11254.t1 12.9675
R14256 a_45928_12082.t0 a_45928_12082.t1 12.9675
R14257 a_42628_9804.t0 a_42628_9804.t1 12.9675
R14258 a_45928_10632.t0 a_45928_10632.t1 12.9675
R14259 a_44128_10426.t0 a_44128_10426.t1 12.9675
R14260 a_43828_9804.t0 a_43828_9804.t1 12.9675
R14261 a_45628_9598.t0 a_45628_9598.t1 12.9675
R14262 a_42928_12082.t0 a_42928_12082.t1 12.9675
R14263 a_42928_10632.t0 a_42928_10632.t1 12.9675
R14264 a_45328_8770.t0 a_45328_8770.t1 12.9675
R14265 a_46828_9598.t0 a_46828_9598.t1 10.2205
R14266 a_43528_10426.t0 a_43528_10426.t1 12.9675
R14267 a_45028_9804.t0 a_45028_9804.t1 12.9675
R14268 a_46528_8976.t0 a_46528_8976.t1 12.9675
R14269 a_43228_9598.t0 a_43228_9598.t1 12.9675
R14270 a_46228_8148.t0 a_46228_8148.t1 12.9675
R14271 a_46828_11254.t0 a_46828_11254.t1 10.2205
C0 A_MUX_0.Tr_Gate_1.CLK VDD 1.93f
C1 RES_74k_1.P VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT 5.27e-19
C2 PFD_T2_0.INV_mag_1.IN PFD_T2_0.FDIV 0.149f
C3 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT 1.64f
C4 mux_magic_2.AND2_magic_0.A S1 0.421f
C5 mux_magic_3.OR_magic_0.A DIV_OUT 0.00118f
C6 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN VDD 0.921f
C7 VCO_DFF_C_0.VCTRL DN 0.109f
C8 RES_74k_1.P S4 0.0112f
C9 PFD_T2_0.INV_mag_0.IN PFD_T2_0.FDIV 3.6e-22
C10 VCO_DFF_C_0.VCO_C_0.OUTB OUTB 0.725f
C11 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN m1_30034_1474# 0.103f
C12 mux_magic_1.AND2_magic_0.A UP_INPUT 7.89e-20
C13 VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.OUTB 1.64f
C14 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VDD 14.9f
C15 PFD_T2_0.INV_mag_1.OUT S2 0.0248f
C16 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.OUTB 0.618f
C17 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VDD 3.8f
C18 PFD_T2_0.DOWN DN_INPUT 0.0322f
C19 RES_74k_1.M m1_53234_16109# 0.782f
C20 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT 1.21f
C21 PFD_T2_0.INV_mag_1.IN mux_magic_3.OR_magic_0.A 2.08e-19
C22 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VDD 0.795f
C23 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN 0.488f
C24 S2 S3 0.0293f
C25 F_IN S6 0.00677f
C26 mux_magic_0.OR_magic_0.B mux_magic_1.OR_magic_0.A 8.13e-19
C27 mux_magic_1.OR_magic_0.A UP 3.03e-19
C28 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_0.IN 1.57f
C29 VCO_DFF_C_0.VCTRL VCTRL_IN 1.25f
C30 mux_magic_3.OR_magic_0.B S3 0.00168f
C31 RES_74k_1.P VDD 23.1f
C32 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT 0.0107f
C33 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_2.IN 0.915f
C34 PFD_T2_0.INV_mag_1.IN S2 0.00119f
C35 RES_74k_1.P A_MUX_0.Tr_Gate_1.CLK 0.496f
C36 mux_magic_2.OR_magic_0.B mux_magic_3.OR_magic_0.A 3.55e-21
C37 PFD_T2_0.Buffer_V_2_0.IN PFD_T2_0.DOWN 0.014f
C38 mux_magic_1.AND2_magic_0.A VDD 1.31f
C39 PFD_T2_0.INV_mag_1.OUT UP_INPUT 0.0197f
C40 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT 1.21f
C41 PFD_T2_0.INV_mag_0.IN S2 0.0531f
C42 VCO_DFF_C_0.VCO_C_0.OUT VCTRL2 0.0145f
C43 mux_magic_0.OR_magic_0.B mux_magic_1.OR_magic_0.B 4.14e-20
C44 PFD_T2_0.UP S2 0.193f
C45 mux_magic_2.OR_magic_0.A mux_magic_3.OR_magic_0.A 0.00129f
C46 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCTRL2 0.344f
C47 mux_magic_1.OR_magic_0.B UP 5.42e-19
C48 PFD_T2_0.INV_mag_1.IN mux_magic_3.OR_magic_0.B 4.1e-19
C49 S6 DIV_OUT 0.272f
C50 VDD ITAIL1 0.775f
C51 VDD PRE_SCALAR 0.922f
C52 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN 0.624f
C53 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN m1_33892_1807# 0.00112f
C54 UP_INPUT S3 8.12e-19
C55 VDD F_IN 0.364f
C56 PFD_T2_0.FIN S2 9.45e-19
C57 mux_magic_1.OR_magic_0.A PFD_T2_0.DOWN 0.00118f
C58 PFD_T2_0.INV_mag_1.OUT PFD_T2_0.INV_mag_0.OUT 0.479f
C59 mux_magic_0.OR_magic_0.A mux_magic_1.OR_magic_0.B 9.11e-20
C60 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT OUTB 0.0234f
C61 mux_magic_2.OR_magic_0.B S2 0.00863f
C62 VCO_DFF_C_0.VCO_C_0.OUTB OUT 0.00703f
C63 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.OUTB 0.0222f
C64 S4 OUTB 0.0286f
C65 PFD_T2_0.Buffer_V_2_1.IN S2 0.0205f
C66 mux_magic_2.OR_magic_0.A S2 0.00163f
C67 mux_magic_2.OR_magic_0.B mux_magic_3.OR_magic_0.B 0.00142f
C68 PFD_T2_0.INV_mag_1.OUT VDD 0.708f
C69 mux_magic_0.AND2_magic_0.A S2 0.428f
C70 PFD_T2_0.INV_mag_0.IN UP_INPUT 4.06e-19
C71 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.OUT 0.385f
C72 PFD_T2_0.UP UP_INPUT 0.13f
C73 mux_magic_2.OR_magic_0.A mux_magic_3.OR_magic_0.B 3.55e-21
C74 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_4.IN 0.00342f
C75 mux_magic_1.OR_magic_0.B DN 0.00106f
C76 VDD DIV_OUT 0.892f
C77 mux_magic_0.OR_magic_0.B ITAIL 5.71e-19
C78 mux_magic_1.OR_magic_0.B DN_INPUT 0.00118f
C79 UP ITAIL 0.634f
C80 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT 3.61e-20
C81 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_5.IN 3.46e-19
C82 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_3.IN 3.19f
C83 VDD S3 2.39f
C84 PFD_T2_0.INV_mag_1.IN PFD_T2_0.INV_mag_0.OUT 0.218f
C85 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VDD 2.87f
C86 mux_magic_2.OR_magic_0.B UP_INPUT 1.47e-19
C87 mux_magic_0.OR_magic_0.A S2 1.1e-20
C88 PFD_T2_0.FDIV mux_magic_3.AND2_magic_0.A 8.78e-21
C89 PFD_T2_0.INV_mag_0.IN PFD_T2_0.INV_mag_0.OUT 0.318f
C90 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN 7.97e-19
C91 PFD_T2_0.FDIV PFD_T2_0.Buffer_V_2_0.IN 0.00947f
C92 RES_74k_1.P ITAIL1 1.67f
C93 PFD_T2_0.Buffer_V_2_1.IN UP_INPUT 1.54e-20
C94 VCO_DFF_C_0.VCTRL VCTRL2 0.227f
C95 VDD OUTB 0.781f
C96 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT 0.765f
C97 PFD_T2_0.INV_mag_1.IN VDD 5f
C98 A_MUX_0.Tr_Gate_1.CLK OUTB 0.00188f
C99 PFD_T2_0.FIN PFD_T2_0.INV_mag_0.OUT 0.0515f
C100 PFD_T2_0.DOWN S2 1.31e-20
C101 VCO_DFF_C_0.VCO_C_0.OUT VDD 0.723f
C102 mux_magic_0.AND2_magic_0.A UP_INPUT 0.0788f
C103 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VDD 12.5f
C104 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT 0.306f
C105 PFD_T2_0.INV_mag_0.IN VDD 4.75f
C106 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.OUTB 0.915f
C107 mux_magic_0.OR_magic_0.B UP_INPUT 0.00118f
C108 VCO_DFF_C_0.VCO_C_0.OUTB VCTRL_IN 0.00272f
C109 PFD_T2_0.UP VDD 0.977f
C110 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT 0.419f
C111 ITAIL DN 0.0315f
C112 S2 DN_INPUT 0.785f
C113 mux_magic_3.OR_magic_0.A mux_magic_3.AND2_magic_0.A 0.00108f
C114 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT OUT 0.577f
C115 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.INV_mag_0.OUT 0.00184f
C116 PRE_SCALAR F_IN 0.0271f
C117 PFD_T2_0.FIN VDD 0.785f
C118 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK OUTB 0.493f
C119 mux_magic_2.OR_magic_0.B VDD 1.19f
C120 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.OUT 9.22e-19
C121 VCO_DFF_C_0.VCTRL S4 0.523f
C122 mux_magic_1.OR_magic_0.B mux_magic_1.OR_magic_0.A 0.178f
C123 m1_33892_1807# VDD 0.0434f
C124 PFD_T2_0.Buffer_V_2_1.IN VDD 1.18f
C125 mux_magic_2.OR_magic_0.A VDD 1.23f
C126 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_4.IN 0.13f
C127 m1_30034_1474# VDD 0.0163f
C128 mux_magic_1.AND2_magic_0.A S3 0.425f
C129 PFD_T2_0.DOWN UP_INPUT 0.00739f
C130 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_5.IN 0.391f
C131 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT 0.02f
C132 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT 0.389f
C133 mux_magic_0.AND2_magic_0.A VDD 1.32f
C134 mux_magic_0.OR_magic_0.B VDD 1.2f
C135 VDD UP 0.998f
C136 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN m1_33892_1807# 0.106f
C137 UP_INPUT DN_INPUT 0.95f
C138 RES_74k_1.P OUTB 0.168f
C139 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCTRL2 0.321f
C140 S1 S6 0.0283f
C141 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VDD 2.74f
C142 mux_magic_0.OR_magic_0.A VDD 1.24f
C143 PFD_T2_0.INV_mag_0.OUT PFD_T2_0.DOWN 7.95e-19
C144 mux_magic_2.AND2_magic_0.A VDD 1.3f
C145 VDD OUT 4.42f
C146 VCO_DFF_C_0.VCTRL VDD 12.8f
C147 A_MUX_0.Tr_Gate_1.CLK VCO_DFF_C_0.VCTRL 0.422f
C148 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.OUTB 0.348f
C149 PFD_T2_0.INV_mag_0.OUT DN_INPUT 0.142f
C150 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN OUT 0.382f
C151 mux_magic_3.AND2_magic_0.A S6 0.425f
C152 PFD_T2_0.INV_mag_1.OUT S3 6.87e-19
C153 PFD_T2_0.DOWN VDD 1.07f
C154 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN 0.546f
C155 S4 VCTRL_IN 0.548f
C156 mux_magic_3.OR_magic_0.B PFD_T2_0.FDIV 1.24e-20
C157 VDD DN 2.35f
C158 VCO_DFF_C_0.VCO_C_0.OUTB VCTRL2 0.00407f
C159 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_2.IN 1.63f
C160 VDD DN_INPUT 0.853f
C161 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK OUT 0.00102f
C162 VDD S1 1.8f
C163 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_4.IN 0.00756f
C164 PFD_T2_0.INV_mag_1.IN PFD_T2_0.INV_mag_1.OUT 0.229f
C165 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT 0.0108f
C166 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.IN 0.388f
C167 mux_magic_2.OR_magic_0.B F_IN 0.00118f
C168 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT 0.00912f
C169 PFD_T2_0.INV_mag_0.OUT PFD_T2_0.Buffer_V_2_0.IN 0.187f
C170 RES_74k_1.P UP 0.00276f
C171 PFD_T2_0.INV_mag_0.IN PFD_T2_0.INV_mag_1.OUT 0.405f
C172 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT 0.403f
C173 mux_magic_2.OR_magic_0.A PRE_SCALAR 0.00118f
C174 PFD_T2_0.UP PFD_T2_0.INV_mag_1.OUT 0.0222f
C175 mux_magic_3.AND2_magic_0.A VDD 1.29f
C176 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT OUTB 0.00852f
C177 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VDD 0.958f
C178 mux_magic_3.OR_magic_0.B mux_magic_3.OR_magic_0.A 0.178f
C179 VCO_DFF_C_0.VCO_C_0.OUTB S4 0.0152f
C180 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCTRL2 0.0917f
C181 RES_74k_1.P OUT 0.0217f
C182 RES_74k_1.P VCO_DFF_C_0.VCTRL 1.41f
C183 PFD_T2_0.Buffer_V_2_0.IN VDD 1.3f
C184 UP ITAIL1 0.079f
C185 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VDD 14.8f
C186 RES_74k_1.M VDD 0.826f
C187 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.OUTB 0.00204f
C188 VDD VCTRL_IN 0.112f
C189 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VDD 2.15f
C190 PFD_T2_0.INV_mag_0.OUT PFD_T2_0.FDIV 0.0514f
C191 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.INV_mag_1.OUT 0.135f
C192 mux_magic_2.AND2_magic_0.A PRE_SCALAR 0.574f
C193 PFD_T2_0.DOWN mux_magic_1.AND2_magic_0.A 0.408f
C194 mux_magic_2.AND2_magic_0.A F_IN 0.0189f
C195 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT 0.00977f
C196 PFD_T2_0.INV_mag_0.IN PFD_T2_0.INV_mag_1.IN 1.33f
C197 mux_magic_3.OR_magic_0.A S6 1.1e-20
C198 mux_magic_1.OR_magic_0.A VDD 1.24f
C199 RES_74k_1.P DN 1.07e-19
C200 PFD_T2_0.UP PFD_T2_0.INV_mag_1.IN 4.12e-19
C201 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.OUT 0.791f
C202 mux_magic_1.AND2_magic_0.A DN 8.78e-21
C203 PFD_T2_0.FDIV VDD 0.84f
C204 mux_magic_1.AND2_magic_0.A DN_INPUT 0.0174f
C205 PFD_T2_0.FIN PFD_T2_0.INV_mag_1.IN 0.0083f
C206 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT 7.5e-19
C207 PFD_T2_0.UP PFD_T2_0.INV_mag_0.IN 1.06e-19
C208 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_4.IN 2.23e-19
C209 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.IN 3.46e-19
C210 VCO_DFF_C_0.VCO_C_0.OUTB VDD 5.93f
C211 PFD_T2_0.FIN PFD_T2_0.INV_mag_0.IN 0.141f
C212 DN ITAIL1 5.59e-19
C213 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.IN 0.809f
C214 S2 UP_INPUT 0.34f
C215 mux_magic_1.OR_magic_0.B VDD 1.19f
C216 mux_magic_2.OR_magic_0.B PFD_T2_0.INV_mag_0.IN 3.92e-19
C217 S1 PRE_SCALAR 0.426f
C218 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.INV_mag_1.IN 0.0388f
C219 S1 F_IN 0.515f
C220 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT 0.403f
C221 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.INV_mag_0.IN 0.428f
C222 mux_magic_2.OR_magic_0.A PFD_T2_0.INV_mag_0.IN 2.07e-19
C223 mux_magic_2.OR_magic_0.B PFD_T2_0.FIN 3.02e-21
C224 PFD_T2_0.INV_mag_1.OUT PFD_T2_0.DOWN 0.0184f
C225 mux_magic_3.OR_magic_0.A VDD 1.23f
C226 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN m1_30034_1474# 0.00112f
C227 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCTRL2 0.0273f
C228 PFD_T2_0.UP PFD_T2_0.Buffer_V_2_1.IN 0.00913f
C229 RES_74k_1.P RES_74k_1.M 0.231f
C230 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.OUTB 0.0179f
C231 RES_74k_1.P VCTRL_IN 4.84e-20
C232 PFD_T2_0.INV_mag_0.OUT S2 1.77e-20
C233 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT OUT 0.0191f
C234 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK 0.703f
C235 PFD_T2_0.FIN PFD_T2_0.Buffer_V_2_1.IN 0.00931f
C236 PFD_T2_0.INV_mag_1.OUT DN_INPUT 0.216f
C237 mux_magic_0.AND2_magic_0.A PFD_T2_0.UP 0.376f
C238 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VDD 12.6f
C239 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN OUTB 1.27f
C240 mux_magic_3.AND2_magic_0.A F_IN 5.44e-19
C241 mux_magic_2.OR_magic_0.A mux_magic_2.OR_magic_0.B 0.178f
C242 PFD_T2_0.DOWN S3 0.203f
C243 OUTB OUT 0.5f
C244 VCO_DFF_C_0.VCTRL OUTB 0.0294f
C245 VDD S2 3f
C246 mux_magic_1.OR_magic_0.A mux_magic_1.AND2_magic_0.A 0.00108f
C247 VDD ITAIL 6.65f
C248 S3 DN_INPUT 0.214f
C249 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.OUT 0.0471f
C250 PFD_T2_0.UP mux_magic_0.OR_magic_0.A 0.00118f
C251 VDD VCTRL2 1.23f
C252 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_5.IN 3.31f
C253 mux_magic_0.AND2_magic_0.A PFD_T2_0.Buffer_V_2_1.IN 2.76e-20
C254 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN 10.3f
C255 PFD_T2_0.INV_mag_1.IN PFD_T2_0.DOWN 0.0028f
C256 mux_magic_2.AND2_magic_0.A PFD_T2_0.FIN 8.78e-21
C257 mux_magic_3.OR_magic_0.B VDD 1.19f
C258 PFD_T2_0.INV_mag_1.OUT PFD_T2_0.Buffer_V_2_0.IN 0.0183f
C259 PFD_T2_0.INV_mag_0.OUT UP_INPUT 8.05e-19
C260 mux_magic_3.AND2_magic_0.A DIV_OUT 0.51f
C261 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.IN 0.674f
C262 PFD_T2_0.INV_mag_1.IN DN_INPUT 0.0154f
C263 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VDD 2.59f
C264 mux_magic_0.AND2_magic_0.A UP 8.78e-21
C265 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCTRL2 0.108f
C266 mux_magic_2.AND2_magic_0.A mux_magic_2.OR_magic_0.A 0.00108f
C267 VCO_DFF_C_0.VCTRL m1_33892_1807# 5.46e-20
C268 PFD_T2_0.INV_mag_0.IN DN_INPUT 0.0495f
C269 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT 0.381f
C270 mux_magic_0.OR_magic_0.B UP 0.0203f
C271 VDD S4 2.92f
C272 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN 1.27f
C273 PFD_T2_0.UP DN_INPUT 0.0335f
C274 PFD_T2_0.Buffer_V_2_0.IN S3 0.00109f
C275 mux_magic_0.AND2_magic_0.A mux_magic_0.OR_magic_0.A 0.00108f
C276 A_MUX_0.Tr_Gate_1.CLK S4 0.403f
C277 VDD UP_INPUT 0.694f
C278 VCO_DFF_C_0.VCTRL m1_30034_1474# 0.0168f
C279 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCTRL2 0.198f
C280 VDD S6 1.81f
C281 mux_magic_0.OR_magic_0.A mux_magic_0.OR_magic_0.B 0.178f
C282 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VDD 2.16f
C283 mux_magic_0.OR_magic_0.A UP 0.00973f
C284 mux_magic_2.OR_magic_0.B DN_INPUT 7.17e-19
C285 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VDD 0.893f
C286 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT 0.39f
C287 PFD_T2_0.INV_mag_1.IN PFD_T2_0.Buffer_V_2_0.IN 0.595f
C288 mux_magic_1.OR_magic_0.A S3 1.1e-20
C289 RES_74k_1.P ITAIL 1.83f
C290 PFD_T2_0.Buffer_V_2_1.IN DN_INPUT 0.0136f
C291 mux_magic_2.OR_magic_0.A DN_INPUT 2.66e-20
C292 PFD_T2_0.INV_mag_0.OUT VDD 0.674f
C293 VCTRL_IN OUTB 0.0234f
C294 mux_magic_2.OR_magic_0.A S1 1.1e-20
C295 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.OUT 1.19f
C296 PFD_T2_0.INV_mag_0.IN PFD_T2_0.Buffer_V_2_0.IN 0.0412f
C297 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN 10.4f
C298 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_4.IN 0.4f
C299 mux_magic_0.AND2_magic_0.A DN_INPUT 2.16e-19
C300 VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT 5.91e-19
C301 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT 0.00409f
C302 UP DN 0.547f
C303 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_2.IN 1.2f
C304 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT 0.652f
C305 ITAIL ITAIL1 0.0176f
.ends

