magic
tech gf180mcuD
magscale 1 10
timestamp 1713971361
<< checkpaint >>
rect -3420 -2036 16830 9134
<< nwell >>
rect 6621 2240 6774 2933
rect 6663 516 6799 1207
<< pwell >>
rect 6552 2040 6848 2177
rect 5665 1329 6864 1466
<< psubdiff >>
rect -1321 6670 14510 6671
rect -1321 6663 14820 6670
rect -1321 6639 14821 6663
rect -1321 6623 14739 6639
rect -1321 6577 -1261 6623
rect -1215 6577 -1111 6623
rect -1065 6577 -961 6623
rect -915 6577 -811 6623
rect -765 6577 -661 6623
rect -615 6577 -511 6623
rect -465 6577 -361 6623
rect -315 6577 -211 6623
rect -165 6577 -61 6623
rect -15 6577 89 6623
rect 135 6577 239 6623
rect 285 6577 389 6623
rect 435 6577 539 6623
rect 585 6577 689 6623
rect 735 6577 839 6623
rect 885 6577 989 6623
rect 1035 6577 1139 6623
rect 1185 6577 1289 6623
rect 1335 6577 1439 6623
rect 1485 6577 1589 6623
rect 1635 6577 1739 6623
rect 1785 6577 1889 6623
rect 1935 6577 2039 6623
rect 2085 6577 2189 6623
rect 2235 6577 2339 6623
rect 2385 6577 2489 6623
rect 2535 6577 2639 6623
rect 2685 6577 2789 6623
rect 2835 6577 2939 6623
rect 2985 6577 3089 6623
rect 3135 6577 3239 6623
rect 3285 6577 3389 6623
rect 3435 6577 3539 6623
rect 3585 6577 3689 6623
rect 3735 6577 3839 6623
rect 3885 6577 3989 6623
rect 4035 6577 4139 6623
rect 4185 6577 4289 6623
rect 4335 6577 4439 6623
rect 4485 6577 4589 6623
rect 4635 6577 4739 6623
rect 4785 6577 4889 6623
rect 4935 6577 5039 6623
rect 5085 6577 5189 6623
rect 5235 6577 5339 6623
rect 5385 6577 5489 6623
rect 5535 6577 5639 6623
rect 5685 6577 5789 6623
rect 5835 6577 5939 6623
rect 5985 6577 6089 6623
rect 6135 6577 6239 6623
rect 6285 6577 6389 6623
rect 6435 6577 6539 6623
rect 6585 6577 6689 6623
rect 6735 6577 6839 6623
rect 6885 6577 6989 6623
rect 7035 6577 7139 6623
rect 7185 6577 7289 6623
rect 7335 6577 7439 6623
rect 7485 6577 7589 6623
rect 7635 6577 7739 6623
rect 7785 6577 7889 6623
rect 7935 6577 8039 6623
rect 8085 6577 8189 6623
rect 8235 6577 8339 6623
rect 8385 6577 8489 6623
rect 8535 6577 8639 6623
rect 8685 6577 8789 6623
rect 8835 6577 8939 6623
rect 8985 6577 9089 6623
rect 9135 6577 9239 6623
rect 9285 6577 9389 6623
rect 9435 6577 9539 6623
rect 9585 6577 9689 6623
rect 9735 6577 9839 6623
rect 9885 6577 9989 6623
rect 10035 6577 10139 6623
rect 10185 6577 10289 6623
rect 10335 6577 10439 6623
rect 10485 6577 10589 6623
rect 10635 6577 10739 6623
rect 10785 6577 10889 6623
rect 10935 6577 11039 6623
rect 11085 6577 11189 6623
rect 11235 6577 11339 6623
rect 11385 6577 11489 6623
rect 11535 6577 11639 6623
rect 11685 6577 11789 6623
rect 11835 6577 11939 6623
rect 11985 6577 12089 6623
rect 12135 6577 12239 6623
rect 12285 6577 12389 6623
rect 12435 6577 12539 6623
rect 12585 6577 12689 6623
rect 12735 6577 12839 6623
rect 12885 6577 12989 6623
rect 13035 6577 13139 6623
rect 13185 6577 13289 6623
rect 13335 6577 13439 6623
rect 13485 6577 13589 6623
rect 13635 6577 13739 6623
rect 13785 6577 13889 6623
rect 13935 6577 14039 6623
rect 14085 6577 14189 6623
rect 14235 6577 14339 6623
rect 14385 6616 14739 6623
rect 14385 6577 14544 6616
rect -1321 6570 14544 6577
rect 14590 6593 14739 6616
rect 14785 6593 14821 6639
rect 14590 6570 14821 6593
rect -1321 6543 14821 6570
rect -1321 6542 14510 6543
rect -1321 6506 -1192 6542
rect 14690 6530 14821 6543
rect -1321 6460 -1286 6506
rect -1240 6460 -1192 6506
rect -1321 6356 -1192 6460
rect -1321 6310 -1286 6356
rect -1240 6310 -1192 6356
rect -1321 6206 -1192 6310
rect -1321 6160 -1286 6206
rect -1240 6160 -1192 6206
rect -1321 6056 -1192 6160
rect -1321 6010 -1286 6056
rect -1240 6010 -1192 6056
rect -1321 5906 -1192 6010
rect -1321 5860 -1286 5906
rect -1240 5860 -1192 5906
rect -1321 5756 -1192 5860
rect -1321 5710 -1286 5756
rect -1240 5710 -1192 5756
rect -1321 5606 -1192 5710
rect -1321 5560 -1286 5606
rect -1240 5560 -1192 5606
rect -1321 5456 -1192 5560
rect -1321 5410 -1286 5456
rect -1240 5410 -1192 5456
rect -1321 5306 -1192 5410
rect -1321 5260 -1286 5306
rect -1240 5260 -1192 5306
rect -1321 5156 -1192 5260
rect -1321 5110 -1286 5156
rect -1240 5110 -1192 5156
rect -1321 5006 -1192 5110
rect -1321 4960 -1286 5006
rect -1240 4960 -1192 5006
rect -1321 4856 -1192 4960
rect -1321 4810 -1286 4856
rect -1240 4810 -1192 4856
rect -1321 4706 -1192 4810
rect -1321 4660 -1286 4706
rect -1240 4660 -1192 4706
rect -1321 4556 -1192 4660
rect -1321 4510 -1286 4556
rect -1240 4510 -1192 4556
rect -1321 4406 -1192 4510
rect -1321 4360 -1286 4406
rect -1240 4360 -1192 4406
rect -1321 4256 -1192 4360
rect -1321 4210 -1286 4256
rect -1240 4210 -1192 4256
rect -1321 4106 -1192 4210
rect -1321 4060 -1286 4106
rect -1240 4060 -1192 4106
rect -1321 3956 -1192 4060
rect -1321 3910 -1286 3956
rect -1240 3910 -1192 3956
rect -1321 3806 -1192 3910
rect -1321 3760 -1286 3806
rect -1240 3760 -1192 3806
rect -1321 3656 -1192 3760
rect -1321 3610 -1286 3656
rect -1240 3610 -1192 3656
rect -1321 3506 -1192 3610
rect -1321 3460 -1286 3506
rect -1240 3460 -1192 3506
rect -1321 3356 -1192 3460
rect -1321 3310 -1286 3356
rect -1240 3310 -1192 3356
rect -1321 3206 -1192 3310
rect -1321 3160 -1286 3206
rect -1240 3160 -1192 3206
rect -1321 3056 -1192 3160
rect -1321 3010 -1286 3056
rect -1240 3010 -1192 3056
rect -1321 2906 -1192 3010
rect -1321 2860 -1286 2906
rect -1240 2860 -1192 2906
rect -1321 2756 -1192 2860
rect -1321 2710 -1286 2756
rect -1240 2710 -1192 2756
rect -1321 2606 -1192 2710
rect -1321 2560 -1286 2606
rect -1240 2560 -1192 2606
rect -1321 2456 -1192 2560
rect -1321 2410 -1286 2456
rect -1240 2410 -1192 2456
rect -1321 2306 -1192 2410
rect -1321 2260 -1286 2306
rect -1240 2260 -1192 2306
rect -1321 2156 -1192 2260
rect -1321 2110 -1286 2156
rect -1240 2110 -1192 2156
rect -1321 2006 -1192 2110
rect -1321 1960 -1286 2006
rect -1240 1960 -1192 2006
rect -1321 1856 -1192 1960
rect -1321 1810 -1286 1856
rect -1240 1810 -1192 1856
rect -1321 1706 -1192 1810
rect -1321 1660 -1286 1706
rect -1240 1660 -1192 1706
rect -1321 1556 -1192 1660
rect -1321 1510 -1286 1556
rect -1240 1510 -1192 1556
rect -1321 1406 -1192 1510
rect -1321 1360 -1286 1406
rect -1240 1360 -1192 1406
rect -1321 1256 -1192 1360
rect -1321 1210 -1286 1256
rect -1240 1210 -1192 1256
rect -1321 1106 -1192 1210
rect -1321 1060 -1286 1106
rect -1240 1060 -1192 1106
rect -1321 956 -1192 1060
rect -1321 910 -1286 956
rect -1240 910 -1192 956
rect -1321 806 -1192 910
rect -1321 760 -1286 806
rect -1240 760 -1192 806
rect -1321 656 -1192 760
rect -1321 610 -1286 656
rect -1240 610 -1192 656
rect -1321 506 -1192 610
rect -1321 460 -1286 506
rect -1240 460 -1192 506
rect -1321 356 -1192 460
rect -1321 310 -1286 356
rect -1240 310 -1192 356
rect -1321 206 -1192 310
rect -1321 160 -1286 206
rect -1240 160 -1192 206
rect -1321 116 -1192 160
rect 14692 6489 14821 6530
rect 14692 6443 14739 6489
rect 14785 6443 14821 6489
rect 14692 6339 14821 6443
rect 14692 6293 14739 6339
rect 14785 6293 14821 6339
rect 14692 6189 14821 6293
rect 14692 6143 14739 6189
rect 14785 6143 14821 6189
rect 14692 6039 14821 6143
rect 14692 5993 14739 6039
rect 14785 5993 14821 6039
rect 14692 5889 14821 5993
rect 14692 5843 14739 5889
rect 14785 5843 14821 5889
rect 14692 5739 14821 5843
rect 14692 5693 14739 5739
rect 14785 5693 14821 5739
rect 14692 5589 14821 5693
rect 14692 5543 14739 5589
rect 14785 5543 14821 5589
rect 14692 5439 14821 5543
rect 14692 5393 14739 5439
rect 14785 5393 14821 5439
rect 14692 5289 14821 5393
rect 14692 5243 14739 5289
rect 14785 5243 14821 5289
rect 14692 5139 14821 5243
rect 14692 5093 14739 5139
rect 14785 5093 14821 5139
rect 14692 4989 14821 5093
rect 14692 4943 14739 4989
rect 14785 4943 14821 4989
rect 14692 4839 14821 4943
rect 14692 4793 14739 4839
rect 14785 4793 14821 4839
rect 14692 4689 14821 4793
rect 14692 4643 14739 4689
rect 14785 4643 14821 4689
rect 14692 4539 14821 4643
rect 14692 4493 14739 4539
rect 14785 4493 14821 4539
rect 14692 4389 14821 4493
rect 14692 4343 14739 4389
rect 14785 4343 14821 4389
rect 14692 4239 14821 4343
rect 14692 4193 14739 4239
rect 14785 4193 14821 4239
rect 14692 4089 14821 4193
rect 14692 4043 14739 4089
rect 14785 4043 14821 4089
rect 14692 3939 14821 4043
rect 14692 3893 14739 3939
rect 14785 3893 14821 3939
rect 14692 3789 14821 3893
rect 14692 3743 14739 3789
rect 14785 3743 14821 3789
rect 14692 3639 14821 3743
rect 14692 3593 14739 3639
rect 14785 3593 14821 3639
rect 14692 3489 14821 3593
rect 14692 3443 14739 3489
rect 14785 3443 14821 3489
rect 14692 3339 14821 3443
rect 14692 3293 14739 3339
rect 14785 3293 14821 3339
rect 14692 3189 14821 3293
rect 14692 3143 14739 3189
rect 14785 3143 14821 3189
rect 14692 3039 14821 3143
rect 14692 2993 14739 3039
rect 14785 2993 14821 3039
rect 14692 2889 14821 2993
rect 14692 2843 14739 2889
rect 14785 2843 14821 2889
rect 14692 2739 14821 2843
rect 14692 2693 14739 2739
rect 14785 2693 14821 2739
rect 14692 2589 14821 2693
rect 14692 2543 14739 2589
rect 14785 2543 14821 2589
rect 14692 2439 14821 2543
rect 14692 2393 14739 2439
rect 14785 2393 14821 2439
rect 14692 2289 14821 2393
rect 14692 2243 14739 2289
rect 14785 2243 14821 2289
rect 14692 2139 14821 2243
rect 14692 2093 14739 2139
rect 14785 2093 14821 2139
rect 14692 1989 14821 2093
rect 14692 1943 14739 1989
rect 14785 1943 14821 1989
rect 14692 1839 14821 1943
rect 14692 1793 14739 1839
rect 14785 1793 14821 1839
rect 14692 1689 14821 1793
rect 14692 1643 14739 1689
rect 14785 1643 14821 1689
rect 14692 1539 14821 1643
rect 14692 1493 14739 1539
rect 14785 1493 14821 1539
rect 14692 1389 14821 1493
rect 14692 1343 14739 1389
rect 14785 1343 14821 1389
rect 14692 1239 14821 1343
rect 14692 1193 14739 1239
rect 14785 1193 14821 1239
rect 14692 1089 14821 1193
rect 14692 1043 14739 1089
rect 14785 1043 14821 1089
rect 14692 939 14821 1043
rect 14692 893 14739 939
rect 14785 893 14821 939
rect 14692 789 14821 893
rect 14692 743 14739 789
rect 14785 743 14821 789
rect 14692 639 14821 743
rect 14692 593 14739 639
rect 14785 593 14821 639
rect 14692 489 14821 593
rect 14692 443 14739 489
rect 14785 443 14821 489
rect 14692 339 14821 443
rect 14692 293 14739 339
rect 14785 293 14821 339
rect 14692 189 14821 293
rect 14692 143 14739 189
rect 14785 143 14821 189
rect -1321 108 14510 116
rect 14692 108 14821 143
rect -1321 79 14821 108
rect -1321 56 -1091 79
rect -1321 10 -1286 56
rect -1240 33 -1091 56
rect -1045 33 -941 79
rect -895 33 -791 79
rect -745 33 -641 79
rect -595 33 -491 79
rect -445 33 -341 79
rect -295 33 -191 79
rect -145 33 -41 79
rect 5 33 109 79
rect 155 33 259 79
rect 305 33 409 79
rect 455 33 559 79
rect 605 33 709 79
rect 755 33 859 79
rect 905 33 1009 79
rect 1055 33 1159 79
rect 1205 33 1309 79
rect 1355 33 1459 79
rect 1505 33 1609 79
rect 1655 33 1759 79
rect 1805 33 1909 79
rect 1955 33 2059 79
rect 2105 33 2209 79
rect 2255 33 2359 79
rect 2405 33 2509 79
rect 2555 33 2659 79
rect 2705 33 2809 79
rect 2855 33 2959 79
rect 3005 33 3109 79
rect 3155 33 3259 79
rect 3305 33 3409 79
rect 3455 33 3559 79
rect 3605 33 3709 79
rect 3755 33 3859 79
rect 3905 33 4009 79
rect 4055 33 4159 79
rect 4205 33 4309 79
rect 4355 33 4459 79
rect 4505 33 4609 79
rect 4655 33 4759 79
rect 4805 33 4909 79
rect 4955 33 5059 79
rect 5105 33 5209 79
rect 5255 33 5359 79
rect 5405 33 5509 79
rect 5555 33 5659 79
rect 5705 33 5809 79
rect 5855 33 5959 79
rect 6005 33 6109 79
rect 6155 33 6259 79
rect 6305 33 6409 79
rect 6455 33 6559 79
rect 6605 33 6709 79
rect 6755 33 6859 79
rect 6905 33 7009 79
rect 7055 33 7159 79
rect 7205 33 7309 79
rect 7355 33 7459 79
rect 7505 33 7609 79
rect 7655 33 7759 79
rect 7805 33 7909 79
rect 7955 33 8059 79
rect 8105 33 8209 79
rect 8255 33 8359 79
rect 8405 33 8509 79
rect 8555 33 8659 79
rect 8705 33 8809 79
rect 8855 33 8959 79
rect 9005 33 9109 79
rect 9155 33 9259 79
rect 9305 33 9409 79
rect 9455 33 9559 79
rect 9605 33 9709 79
rect 9755 33 9859 79
rect 9905 33 10009 79
rect 10055 33 10159 79
rect 10205 33 10309 79
rect 10355 33 10459 79
rect 10505 33 10609 79
rect 10655 33 10759 79
rect 10805 33 10909 79
rect 10955 33 11059 79
rect 11105 33 11209 79
rect 11255 33 11359 79
rect 11405 33 11509 79
rect 11555 33 11659 79
rect 11705 33 11809 79
rect 11855 33 11959 79
rect 12005 33 12109 79
rect 12155 33 12259 79
rect 12305 33 12409 79
rect 12455 33 12559 79
rect 12605 33 12709 79
rect 12755 33 12859 79
rect 12905 33 13009 79
rect 13055 33 13159 79
rect 13205 33 13309 79
rect 13355 33 13459 79
rect 13505 33 13609 79
rect 13655 33 13759 79
rect 13805 33 13909 79
rect 13955 33 14059 79
rect 14105 33 14209 79
rect 14255 33 14359 79
rect 14405 72 14821 79
rect 14405 33 14564 72
rect -1240 26 14564 33
rect 14610 26 14714 72
rect 14760 26 14821 72
rect -1240 10 14821 26
rect -1321 -13 14821 10
rect 14510 -21 14821 -13
<< psubdiffcont >>
rect -1261 6577 -1215 6623
rect -1111 6577 -1065 6623
rect -961 6577 -915 6623
rect -811 6577 -765 6623
rect -661 6577 -615 6623
rect -511 6577 -465 6623
rect -361 6577 -315 6623
rect -211 6577 -165 6623
rect -61 6577 -15 6623
rect 89 6577 135 6623
rect 239 6577 285 6623
rect 389 6577 435 6623
rect 539 6577 585 6623
rect 689 6577 735 6623
rect 839 6577 885 6623
rect 989 6577 1035 6623
rect 1139 6577 1185 6623
rect 1289 6577 1335 6623
rect 1439 6577 1485 6623
rect 1589 6577 1635 6623
rect 1739 6577 1785 6623
rect 1889 6577 1935 6623
rect 2039 6577 2085 6623
rect 2189 6577 2235 6623
rect 2339 6577 2385 6623
rect 2489 6577 2535 6623
rect 2639 6577 2685 6623
rect 2789 6577 2835 6623
rect 2939 6577 2985 6623
rect 3089 6577 3135 6623
rect 3239 6577 3285 6623
rect 3389 6577 3435 6623
rect 3539 6577 3585 6623
rect 3689 6577 3735 6623
rect 3839 6577 3885 6623
rect 3989 6577 4035 6623
rect 4139 6577 4185 6623
rect 4289 6577 4335 6623
rect 4439 6577 4485 6623
rect 4589 6577 4635 6623
rect 4739 6577 4785 6623
rect 4889 6577 4935 6623
rect 5039 6577 5085 6623
rect 5189 6577 5235 6623
rect 5339 6577 5385 6623
rect 5489 6577 5535 6623
rect 5639 6577 5685 6623
rect 5789 6577 5835 6623
rect 5939 6577 5985 6623
rect 6089 6577 6135 6623
rect 6239 6577 6285 6623
rect 6389 6577 6435 6623
rect 6539 6577 6585 6623
rect 6689 6577 6735 6623
rect 6839 6577 6885 6623
rect 6989 6577 7035 6623
rect 7139 6577 7185 6623
rect 7289 6577 7335 6623
rect 7439 6577 7485 6623
rect 7589 6577 7635 6623
rect 7739 6577 7785 6623
rect 7889 6577 7935 6623
rect 8039 6577 8085 6623
rect 8189 6577 8235 6623
rect 8339 6577 8385 6623
rect 8489 6577 8535 6623
rect 8639 6577 8685 6623
rect 8789 6577 8835 6623
rect 8939 6577 8985 6623
rect 9089 6577 9135 6623
rect 9239 6577 9285 6623
rect 9389 6577 9435 6623
rect 9539 6577 9585 6623
rect 9689 6577 9735 6623
rect 9839 6577 9885 6623
rect 9989 6577 10035 6623
rect 10139 6577 10185 6623
rect 10289 6577 10335 6623
rect 10439 6577 10485 6623
rect 10589 6577 10635 6623
rect 10739 6577 10785 6623
rect 10889 6577 10935 6623
rect 11039 6577 11085 6623
rect 11189 6577 11235 6623
rect 11339 6577 11385 6623
rect 11489 6577 11535 6623
rect 11639 6577 11685 6623
rect 11789 6577 11835 6623
rect 11939 6577 11985 6623
rect 12089 6577 12135 6623
rect 12239 6577 12285 6623
rect 12389 6577 12435 6623
rect 12539 6577 12585 6623
rect 12689 6577 12735 6623
rect 12839 6577 12885 6623
rect 12989 6577 13035 6623
rect 13139 6577 13185 6623
rect 13289 6577 13335 6623
rect 13439 6577 13485 6623
rect 13589 6577 13635 6623
rect 13739 6577 13785 6623
rect 13889 6577 13935 6623
rect 14039 6577 14085 6623
rect 14189 6577 14235 6623
rect 14339 6577 14385 6623
rect 14544 6570 14590 6616
rect 14739 6593 14785 6639
rect -1286 6460 -1240 6506
rect -1286 6310 -1240 6356
rect -1286 6160 -1240 6206
rect -1286 6010 -1240 6056
rect -1286 5860 -1240 5906
rect -1286 5710 -1240 5756
rect -1286 5560 -1240 5606
rect -1286 5410 -1240 5456
rect -1286 5260 -1240 5306
rect -1286 5110 -1240 5156
rect -1286 4960 -1240 5006
rect -1286 4810 -1240 4856
rect -1286 4660 -1240 4706
rect -1286 4510 -1240 4556
rect -1286 4360 -1240 4406
rect -1286 4210 -1240 4256
rect -1286 4060 -1240 4106
rect -1286 3910 -1240 3956
rect -1286 3760 -1240 3806
rect -1286 3610 -1240 3656
rect -1286 3460 -1240 3506
rect -1286 3310 -1240 3356
rect -1286 3160 -1240 3206
rect -1286 3010 -1240 3056
rect -1286 2860 -1240 2906
rect -1286 2710 -1240 2756
rect -1286 2560 -1240 2606
rect -1286 2410 -1240 2456
rect -1286 2260 -1240 2306
rect -1286 2110 -1240 2156
rect -1286 1960 -1240 2006
rect -1286 1810 -1240 1856
rect -1286 1660 -1240 1706
rect -1286 1510 -1240 1556
rect -1286 1360 -1240 1406
rect -1286 1210 -1240 1256
rect -1286 1060 -1240 1106
rect -1286 910 -1240 956
rect -1286 760 -1240 806
rect -1286 610 -1240 656
rect -1286 460 -1240 506
rect -1286 310 -1240 356
rect -1286 160 -1240 206
rect 14739 6443 14785 6489
rect 14739 6293 14785 6339
rect 14739 6143 14785 6189
rect 14739 5993 14785 6039
rect 14739 5843 14785 5889
rect 14739 5693 14785 5739
rect 14739 5543 14785 5589
rect 14739 5393 14785 5439
rect 14739 5243 14785 5289
rect 14739 5093 14785 5139
rect 14739 4943 14785 4989
rect 14739 4793 14785 4839
rect 14739 4643 14785 4689
rect 14739 4493 14785 4539
rect 14739 4343 14785 4389
rect 14739 4193 14785 4239
rect 14739 4043 14785 4089
rect 14739 3893 14785 3939
rect 14739 3743 14785 3789
rect 14739 3593 14785 3639
rect 14739 3443 14785 3489
rect 14739 3293 14785 3339
rect 14739 3143 14785 3189
rect 14739 2993 14785 3039
rect 14739 2843 14785 2889
rect 14739 2693 14785 2739
rect 14739 2543 14785 2589
rect 14739 2393 14785 2439
rect 14739 2243 14785 2289
rect 14739 2093 14785 2139
rect 14739 1943 14785 1989
rect 14739 1793 14785 1839
rect 14739 1643 14785 1689
rect 14739 1493 14785 1539
rect 14739 1343 14785 1389
rect 14739 1193 14785 1239
rect 14739 1043 14785 1089
rect 14739 893 14785 939
rect 14739 743 14785 789
rect 14739 593 14785 639
rect 14739 443 14785 489
rect 14739 293 14785 339
rect 14739 143 14785 189
rect -1286 10 -1240 56
rect -1091 33 -1045 79
rect -941 33 -895 79
rect -791 33 -745 79
rect -641 33 -595 79
rect -491 33 -445 79
rect -341 33 -295 79
rect -191 33 -145 79
rect -41 33 5 79
rect 109 33 155 79
rect 259 33 305 79
rect 409 33 455 79
rect 559 33 605 79
rect 709 33 755 79
rect 859 33 905 79
rect 1009 33 1055 79
rect 1159 33 1205 79
rect 1309 33 1355 79
rect 1459 33 1505 79
rect 1609 33 1655 79
rect 1759 33 1805 79
rect 1909 33 1955 79
rect 2059 33 2105 79
rect 2209 33 2255 79
rect 2359 33 2405 79
rect 2509 33 2555 79
rect 2659 33 2705 79
rect 2809 33 2855 79
rect 2959 33 3005 79
rect 3109 33 3155 79
rect 3259 33 3305 79
rect 3409 33 3455 79
rect 3559 33 3605 79
rect 3709 33 3755 79
rect 3859 33 3905 79
rect 4009 33 4055 79
rect 4159 33 4205 79
rect 4309 33 4355 79
rect 4459 33 4505 79
rect 4609 33 4655 79
rect 4759 33 4805 79
rect 4909 33 4955 79
rect 5059 33 5105 79
rect 5209 33 5255 79
rect 5359 33 5405 79
rect 5509 33 5555 79
rect 5659 33 5705 79
rect 5809 33 5855 79
rect 5959 33 6005 79
rect 6109 33 6155 79
rect 6259 33 6305 79
rect 6409 33 6455 79
rect 6559 33 6605 79
rect 6709 33 6755 79
rect 6859 33 6905 79
rect 7009 33 7055 79
rect 7159 33 7205 79
rect 7309 33 7355 79
rect 7459 33 7505 79
rect 7609 33 7655 79
rect 7759 33 7805 79
rect 7909 33 7955 79
rect 8059 33 8105 79
rect 8209 33 8255 79
rect 8359 33 8405 79
rect 8509 33 8555 79
rect 8659 33 8705 79
rect 8809 33 8855 79
rect 8959 33 9005 79
rect 9109 33 9155 79
rect 9259 33 9305 79
rect 9409 33 9455 79
rect 9559 33 9605 79
rect 9709 33 9755 79
rect 9859 33 9905 79
rect 10009 33 10055 79
rect 10159 33 10205 79
rect 10309 33 10355 79
rect 10459 33 10505 79
rect 10609 33 10655 79
rect 10759 33 10805 79
rect 10909 33 10955 79
rect 11059 33 11105 79
rect 11209 33 11255 79
rect 11359 33 11405 79
rect 11509 33 11555 79
rect 11659 33 11705 79
rect 11809 33 11855 79
rect 11959 33 12005 79
rect 12109 33 12155 79
rect 12259 33 12305 79
rect 12409 33 12455 79
rect 12559 33 12605 79
rect 12709 33 12755 79
rect 12859 33 12905 79
rect 13009 33 13055 79
rect 13159 33 13205 79
rect 13309 33 13355 79
rect 13459 33 13505 79
rect 13609 33 13655 79
rect 13759 33 13805 79
rect 13909 33 13955 79
rect 14059 33 14105 79
rect 14209 33 14255 79
rect 14359 33 14405 79
rect 14564 26 14610 72
rect 14714 26 14760 72
<< metal1 >>
rect 6422 7084 6566 7134
rect 6422 7032 6476 7084
rect 6528 7041 6566 7084
rect 6528 7032 6761 7041
rect 6422 6995 6761 7032
rect 6423 6937 6761 6995
rect 6423 6877 6565 6937
rect 6423 6825 6475 6877
rect 6527 6825 6565 6877
rect 6423 6786 6565 6825
rect 14510 6680 14830 6681
rect -1330 6639 14830 6680
rect -1330 6623 14739 6639
rect -1330 6577 -1261 6623
rect -1215 6577 -1111 6623
rect -1065 6577 -961 6623
rect -915 6577 -811 6623
rect -765 6577 -661 6623
rect -615 6577 -511 6623
rect -465 6577 -361 6623
rect -315 6577 -211 6623
rect -165 6577 -61 6623
rect -15 6577 89 6623
rect 135 6577 239 6623
rect 285 6577 389 6623
rect 435 6577 539 6623
rect 585 6577 689 6623
rect 735 6577 839 6623
rect 885 6577 989 6623
rect 1035 6577 1139 6623
rect 1185 6577 1289 6623
rect 1335 6577 1439 6623
rect 1485 6577 1589 6623
rect 1635 6577 1739 6623
rect 1785 6577 1889 6623
rect 1935 6577 2039 6623
rect 2085 6577 2189 6623
rect 2235 6577 2339 6623
rect 2385 6577 2489 6623
rect 2535 6577 2639 6623
rect 2685 6577 2789 6623
rect 2835 6577 2939 6623
rect 2985 6577 3089 6623
rect 3135 6577 3239 6623
rect 3285 6577 3389 6623
rect 3435 6577 3539 6623
rect 3585 6577 3689 6623
rect 3735 6577 3839 6623
rect 3885 6577 3989 6623
rect 4035 6577 4139 6623
rect 4185 6577 4289 6623
rect 4335 6577 4439 6623
rect 4485 6577 4589 6623
rect 4635 6577 4739 6623
rect 4785 6577 4889 6623
rect 4935 6577 5039 6623
rect 5085 6577 5189 6623
rect 5235 6577 5339 6623
rect 5385 6577 5489 6623
rect 5535 6577 5639 6623
rect 5685 6577 5789 6623
rect 5835 6577 5939 6623
rect 5985 6577 6089 6623
rect 6135 6577 6239 6623
rect 6285 6577 6389 6623
rect 6435 6577 6539 6623
rect 6585 6577 6689 6623
rect 6735 6577 6839 6623
rect 6885 6577 6989 6623
rect 7035 6577 7139 6623
rect 7185 6577 7289 6623
rect 7335 6577 7439 6623
rect 7485 6577 7589 6623
rect 7635 6577 7739 6623
rect 7785 6577 7889 6623
rect 7935 6577 8039 6623
rect 8085 6577 8189 6623
rect 8235 6577 8339 6623
rect 8385 6577 8489 6623
rect 8535 6577 8639 6623
rect 8685 6577 8789 6623
rect 8835 6577 8939 6623
rect 8985 6577 9089 6623
rect 9135 6577 9239 6623
rect 9285 6577 9389 6623
rect 9435 6577 9539 6623
rect 9585 6577 9689 6623
rect 9735 6577 9839 6623
rect 9885 6577 9989 6623
rect 10035 6577 10139 6623
rect 10185 6577 10289 6623
rect 10335 6577 10439 6623
rect 10485 6577 10589 6623
rect 10635 6577 10739 6623
rect 10785 6577 10889 6623
rect 10935 6577 11039 6623
rect 11085 6577 11189 6623
rect 11235 6577 11339 6623
rect 11385 6577 11489 6623
rect 11535 6577 11639 6623
rect 11685 6577 11789 6623
rect 11835 6577 11939 6623
rect 11985 6577 12089 6623
rect 12135 6577 12239 6623
rect 12285 6577 12389 6623
rect 12435 6577 12539 6623
rect 12585 6577 12689 6623
rect 12735 6577 12839 6623
rect 12885 6577 12989 6623
rect 13035 6577 13139 6623
rect 13185 6577 13289 6623
rect 13335 6577 13439 6623
rect 13485 6577 13589 6623
rect 13635 6577 13739 6623
rect 13785 6577 13889 6623
rect 13935 6577 14039 6623
rect 14085 6577 14189 6623
rect 14235 6577 14339 6623
rect 14385 6616 14739 6623
rect 14385 6577 14544 6616
rect -1330 6570 14544 6577
rect 14590 6593 14739 6616
rect 14785 6593 14830 6639
rect 14590 6570 14830 6593
rect -1330 6517 14830 6570
rect -1330 6516 14510 6517
rect -1330 6506 -1166 6516
rect -1330 6460 -1286 6506
rect -1240 6460 -1166 6506
rect -1330 6356 -1166 6460
rect -1330 6310 -1286 6356
rect -1240 6310 -1166 6356
rect -1330 6206 -1166 6310
rect -1330 6160 -1286 6206
rect -1240 6160 -1166 6206
rect -1330 6056 -1166 6160
rect -1330 6010 -1286 6056
rect -1240 6010 -1166 6056
rect -1330 5906 -1166 6010
rect -1330 5860 -1286 5906
rect -1240 5860 -1166 5906
rect -1330 5756 -1166 5860
rect -1330 5710 -1286 5756
rect -1240 5710 -1166 5756
rect -1330 5606 -1166 5710
rect -1330 5560 -1286 5606
rect -1240 5560 -1166 5606
rect -1330 5456 -1166 5560
rect -1330 5410 -1286 5456
rect -1240 5410 -1166 5456
rect -1330 5306 -1166 5410
rect -1330 5260 -1286 5306
rect -1240 5260 -1166 5306
rect -1330 5156 -1166 5260
rect -1330 5110 -1286 5156
rect -1240 5110 -1166 5156
rect -1330 5006 -1166 5110
rect -1330 4960 -1286 5006
rect -1240 4960 -1166 5006
rect -1330 4856 -1166 4960
rect -1330 4810 -1286 4856
rect -1240 4810 -1166 4856
rect -1330 4706 -1166 4810
rect -1330 4660 -1286 4706
rect -1240 4660 -1166 4706
rect -1330 4556 -1166 4660
rect -1330 4510 -1286 4556
rect -1240 4510 -1166 4556
rect 4532 4523 4612 6336
rect 5169 4829 5261 6516
rect 14666 6489 14830 6517
rect 14666 6443 14739 6489
rect 14785 6443 14830 6489
rect 14666 6339 14830 6443
rect 14666 6293 14739 6339
rect 14785 6293 14830 6339
rect 14666 6189 14830 6293
rect 14666 6143 14739 6189
rect 14785 6143 14830 6189
rect 7806 6062 7862 6071
rect 7791 6039 7879 6062
rect 14666 6039 14830 6143
rect 7730 5979 7927 6039
rect 14666 5993 14739 6039
rect 14785 5993 14830 6039
rect 7791 5932 7879 5979
rect 7791 5930 7808 5932
rect 6615 5791 7065 5908
rect 7792 5880 7808 5930
rect 7860 5880 7879 5932
rect 7792 5865 7879 5880
rect 14666 5889 14830 5993
rect 7797 5805 7870 5865
rect 14666 5843 14739 5889
rect 14785 5843 14830 5889
rect 14666 5805 14830 5843
rect 5338 5266 5564 5267
rect 5338 5252 5672 5266
rect 5338 5251 5674 5252
rect 5337 5243 5674 5251
rect 5337 5242 5495 5243
rect 5337 5190 5365 5242
rect 5417 5191 5495 5242
rect 5547 5191 5674 5243
rect 5417 5190 5674 5191
rect 5337 5183 5674 5190
rect 6596 5247 6755 5270
rect 6596 5195 6692 5247
rect 6744 5195 6755 5247
rect 5337 5161 5672 5183
rect 6596 5182 6755 5195
rect 5337 5160 5563 5161
rect 6573 4844 6673 4873
rect 5169 4737 5696 4829
rect 6573 4792 6600 4844
rect 6652 4792 6673 4844
rect 6573 4762 6673 4792
rect -1330 4406 -1166 4510
rect 4280 4502 4612 4523
rect 4280 4450 4484 4502
rect 4536 4450 4612 4502
rect 4280 4438 4612 4450
rect 4280 4414 4558 4438
rect -1330 4360 -1286 4406
rect -1240 4360 -1166 4406
rect 5171 4405 5258 4413
rect 5496 4405 5631 4411
rect -1330 4256 -1166 4360
rect -1330 4210 -1286 4256
rect -1240 4210 -1166 4256
rect 4942 4404 5641 4405
rect 4942 4352 5187 4404
rect 5239 4399 5641 4404
rect 5239 4395 5673 4399
rect 5239 4352 5513 4395
rect 4942 4343 5513 4352
rect 5565 4343 5673 4395
rect 6711 4353 6792 4365
rect 6711 4350 6727 4353
rect 4942 4339 5673 4343
rect 4942 4333 5641 4339
rect 4942 4223 5014 4333
rect 5496 4327 5631 4333
rect 6596 4304 6727 4350
rect 6711 4301 6727 4304
rect 6779 4301 6792 4353
rect 6711 4289 6792 4301
rect -1330 4106 -1166 4210
rect 4934 4214 5021 4223
rect 4934 4162 4950 4214
rect 5002 4162 5021 4214
rect 4934 4147 5021 4162
rect 4942 4124 5014 4147
rect -1330 4060 -1286 4106
rect -1240 4060 -1166 4106
rect -1330 3956 -1166 4060
rect -1330 3910 -1286 3956
rect -1240 3910 -1166 3956
rect -1330 3806 -1166 3910
rect 4151 3905 5664 4003
rect -1330 3760 -1286 3806
rect -1240 3760 -1166 3806
rect 6948 3781 7065 5791
rect 7795 5796 7882 5805
rect 7795 5744 7811 5796
rect 7863 5744 7882 5796
rect 7795 5729 7882 5744
rect 14510 5739 14830 5805
rect 7797 5650 7870 5729
rect 14510 5693 14739 5739
rect 14785 5693 14830 5739
rect 14510 5676 14830 5693
rect 7795 5641 7882 5650
rect 7795 5589 7811 5641
rect 7863 5589 7882 5641
rect 7795 5574 7882 5589
rect 14666 5589 14830 5676
rect 7797 5495 7870 5574
rect 14666 5543 14739 5589
rect 14785 5543 14830 5589
rect 14666 5526 14830 5543
rect 7795 5486 7882 5495
rect 7795 5434 7811 5486
rect 7863 5434 7882 5486
rect 7795 5419 7882 5434
rect 13573 5439 14830 5526
rect 13573 5424 14739 5439
rect 7797 5370 7870 5419
rect 14666 5393 14739 5424
rect 14785 5393 14830 5439
rect 14666 5289 14830 5393
rect 14666 5243 14739 5289
rect 14785 5243 14830 5289
rect 14666 5139 14830 5243
rect 14666 5093 14739 5139
rect 14785 5093 14830 5139
rect 14666 5005 14830 5093
rect 14510 4989 14830 5005
rect 14510 4943 14739 4989
rect 14785 4943 14830 4989
rect 7299 4859 7399 4875
rect 7536 4863 7636 4879
rect 14510 4876 14830 4943
rect 7536 4859 7655 4863
rect 7766 4859 7866 4873
rect 7275 4848 8004 4859
rect 7275 4844 7566 4848
rect 7275 4792 7329 4844
rect 7381 4796 7566 4844
rect 7618 4842 8004 4848
rect 7618 4796 7796 4842
rect 7381 4792 7796 4796
rect 7275 4790 7796 4792
rect 7848 4790 8004 4842
rect 7275 4777 8004 4790
rect 14666 4839 14830 4876
rect 14666 4793 14739 4839
rect 14785 4793 14830 4839
rect 7299 4764 7399 4777
rect 7536 4768 7636 4777
rect 7766 4775 7885 4777
rect 7766 4762 7866 4775
rect 14666 4689 14830 4793
rect 14666 4643 14739 4689
rect 14785 4643 14830 4689
rect 14666 4539 14830 4643
rect 14666 4507 14739 4539
rect 13573 4493 14739 4507
rect 14785 4493 14830 4539
rect 13573 4405 14830 4493
rect 14666 4389 14830 4405
rect 7165 4361 7762 4369
rect 7152 4353 7762 4361
rect 7152 4352 7351 4353
rect 7152 4300 7168 4352
rect 7220 4313 7351 4352
rect 7220 4300 7239 4313
rect 7152 4285 7239 4300
rect 7335 4301 7351 4313
rect 7403 4313 7557 4353
rect 7403 4301 7422 4313
rect 7335 4286 7422 4301
rect 7541 4301 7557 4313
rect 7609 4313 7762 4353
rect 7609 4301 7628 4313
rect 7541 4286 7628 4301
rect 7706 4239 7762 4313
rect 14666 4343 14739 4389
rect 14785 4343 14830 4389
rect 14666 4239 14830 4343
rect 7685 4229 7777 4239
rect 7685 4177 7704 4229
rect 7756 4177 7777 4229
rect 14666 4205 14739 4239
rect 7685 4137 7777 4177
rect 14510 4193 14739 4205
rect 14785 4193 14830 4239
rect 14510 4089 14830 4193
rect 14510 4076 14739 4089
rect 14666 4043 14739 4076
rect 14785 4043 14830 4089
rect 7780 4023 7782 4042
rect 7780 4019 7839 4023
rect 7779 3967 7839 4019
rect 7779 3956 7782 3967
rect -1330 3656 -1166 3760
rect -1330 3610 -1286 3656
rect -1240 3610 -1166 3656
rect 4521 3746 4676 3781
rect 5247 3746 5365 3758
rect 4521 3732 5365 3746
rect 4521 3680 5279 3732
rect 5331 3680 5365 3732
rect 4521 3666 5365 3680
rect 4521 3647 4676 3666
rect 5247 3658 5365 3666
rect -1330 3506 -1166 3610
rect -1330 3460 -1286 3506
rect -1240 3460 -1166 3506
rect -1330 3356 -1166 3460
rect -1330 3310 -1286 3356
rect -1240 3310 -1166 3356
rect -1330 3206 -1166 3310
rect -1330 3160 -1286 3206
rect -1240 3160 -1166 3206
rect -1330 3056 -1166 3160
rect -1330 3010 -1286 3056
rect -1240 3010 -1166 3056
rect -1330 2906 -1166 3010
rect 6122 2965 6303 3670
rect 6542 3664 7065 3781
rect 14666 3939 14830 4043
rect 14666 3893 14739 3939
rect 14785 3893 14830 3939
rect 14666 3789 14830 3893
rect 14666 3743 14739 3789
rect 14785 3743 14830 3789
rect 14666 3639 14830 3743
rect 14666 3593 14739 3639
rect 14785 3593 14830 3639
rect 14666 3489 14830 3593
rect 14666 3443 14739 3489
rect 14785 3443 14830 3489
rect 14666 3339 14830 3443
rect 14666 3293 14739 3339
rect 14785 3293 14830 3339
rect 14666 3189 14830 3293
rect 14666 3143 14739 3189
rect 14785 3143 14830 3189
rect 7669 3012 8726 3113
rect 14666 3039 14830 3143
rect 7669 3008 7770 3012
rect -1330 2860 -1286 2906
rect -1240 2860 -1166 2906
rect -1330 2756 -1166 2860
rect 6614 2858 6819 2933
rect 7670 2911 7770 3008
rect 14666 2993 14739 3039
rect 14785 2993 14830 3039
rect 14666 2889 14830 2993
rect 14666 2843 14739 2889
rect 14785 2843 14830 2889
rect -1330 2710 -1286 2756
rect -1240 2710 -1166 2756
rect -1330 2606 -1166 2710
rect 7994 2788 8093 2807
rect 7994 2736 8023 2788
rect 8075 2736 8093 2788
rect 7994 2638 8093 2736
rect 14666 2739 14830 2843
rect 14666 2693 14739 2739
rect 14785 2693 14830 2739
rect 7994 2629 8098 2638
rect -1330 2560 -1286 2606
rect -1240 2574 -1166 2606
rect -1240 2560 -690 2574
rect -1330 2456 -690 2560
rect -1330 2410 -1286 2456
rect -1240 2445 -690 2456
rect -1240 2410 -1166 2445
rect -1330 2306 -1166 2410
rect -1330 2260 -1286 2306
rect -1240 2260 -1166 2306
rect 5116 2343 5172 2628
rect 7994 2577 8028 2629
rect 8080 2577 8098 2629
rect 7994 2564 8098 2577
rect 14666 2589 14830 2693
rect 7994 2489 8093 2564
rect 7994 2437 8012 2489
rect 8064 2437 8093 2489
rect 7994 2412 8093 2437
rect 14666 2543 14739 2589
rect 14785 2543 14830 2589
rect 14666 2439 14830 2543
rect 5517 2343 5564 2349
rect 5116 2326 5564 2343
rect 7994 2332 8080 2412
rect 5116 2287 5617 2326
rect 5517 2279 5617 2287
rect -1330 2156 -1166 2260
rect 6555 2240 6849 2286
rect 7818 2275 8080 2332
rect 7818 2223 7901 2275
rect 7953 2246 8080 2275
rect 14666 2393 14739 2439
rect 14785 2393 14830 2439
rect 14666 2289 14830 2393
rect 7953 2223 7985 2246
rect 7818 2177 7985 2223
rect 14666 2243 14739 2289
rect 14785 2243 14830 2289
rect -1330 2110 -1286 2156
rect -1240 2110 -1166 2156
rect -1330 2006 -1166 2110
rect -1330 1960 -1286 2006
rect -1240 1960 -1166 2006
rect -1330 1856 -1166 1960
rect 14666 2139 14830 2243
rect 14666 2093 14739 2139
rect 14785 2093 14830 2139
rect 14666 1989 14830 2093
rect 14666 1943 14739 1989
rect 14785 1943 14830 1989
rect 4830 1880 5888 1934
rect -1330 1810 -1286 1856
rect -1240 1810 -1166 1856
rect -1330 1774 -1166 1810
rect 6577 1799 6815 1876
rect 14666 1839 14830 1943
rect -1330 1706 -690 1774
rect -1330 1660 -1286 1706
rect -1240 1660 -690 1706
rect -1330 1645 -690 1660
rect 6667 1651 6766 1799
rect 14666 1793 14739 1839
rect 14785 1793 14830 1839
rect 14666 1689 14830 1793
rect -1330 1556 -1166 1645
rect 6617 1574 6855 1651
rect 14666 1643 14739 1689
rect 14785 1643 14830 1689
rect -1330 1510 -1286 1556
rect -1240 1510 -1166 1556
rect 4833 1514 5891 1568
rect 14666 1539 14830 1643
rect -1330 1406 -1166 1510
rect -1330 1360 -1286 1406
rect -1240 1360 -1166 1406
rect -1330 1256 -1166 1360
rect 14666 1493 14739 1539
rect 14785 1493 14830 1539
rect 14666 1389 14830 1493
rect 14666 1343 14739 1389
rect 14785 1343 14830 1389
rect 7843 1267 7971 1290
rect 8053 1267 8146 1288
rect 8222 1267 8315 1283
rect 8380 1267 8473 1283
rect -1330 1210 -1286 1256
rect -1240 1210 -1166 1256
rect 7796 1259 8525 1267
rect 7796 1258 8072 1259
rect -1330 1106 -1166 1210
rect 6600 1209 6647 1222
rect -1330 1060 -1286 1106
rect -1240 1060 -1166 1106
rect -1330 974 -1166 1060
rect 5124 1118 5629 1174
rect 6600 1163 6855 1209
rect 7796 1206 7895 1258
rect 7947 1207 8072 1258
rect 8124 1254 8525 1259
rect 8124 1207 8241 1254
rect 7947 1206 8241 1207
rect 7796 1202 8241 1206
rect 8293 1202 8399 1254
rect 8451 1202 8525 1254
rect 7796 1192 8525 1202
rect 14666 1239 14830 1343
rect 14666 1193 14739 1239
rect 14785 1193 14830 1239
rect 7843 1184 7971 1192
rect 8053 1186 8146 1192
rect 8222 1181 8315 1192
rect 8380 1181 8473 1192
rect 6600 1151 6647 1163
rect -1330 956 -690 974
rect -1330 910 -1286 956
rect -1240 910 -690 956
rect -1330 845 -690 910
rect -1330 806 -1166 845
rect -1330 760 -1286 806
rect -1240 760 -1166 806
rect -1330 656 -1166 760
rect -1330 610 -1286 656
rect -1240 610 -1166 656
rect -1330 506 -1166 610
rect -1330 460 -1286 506
rect -1240 460 -1166 506
rect -1330 356 -1166 460
rect -1330 310 -1286 356
rect -1240 310 -1166 356
rect -1330 206 -1166 310
rect -1330 160 -1286 206
rect -1240 160 -1166 206
rect -1330 128 -1166 160
rect -712 128 -594 651
rect 88 128 206 651
rect 888 128 1006 698
rect 1688 128 1806 698
rect 5124 594 5180 1118
rect 13599 1095 14510 1171
rect 14666 1089 14830 1193
rect 14666 1043 14739 1089
rect 14785 1043 14830 1089
rect 14666 939 14830 1043
rect 14666 893 14739 939
rect 14785 893 14830 939
rect 7811 763 8731 869
rect 14666 789 14830 893
rect 5026 593 5180 594
rect 14666 743 14739 789
rect 14785 743 14830 789
rect 14666 639 14830 743
rect 14666 593 14739 639
rect 14785 593 14830 639
rect 5026 507 5189 593
rect 6651 516 6828 582
rect 5026 504 5152 507
rect 14666 489 14830 593
rect 14666 443 14739 489
rect 14785 443 14830 489
rect 14666 339 14830 443
rect 14666 293 14739 339
rect 14785 293 14830 339
rect 14666 189 14830 293
rect 14666 143 14739 189
rect 14785 143 14830 189
rect 14666 134 14830 143
rect 14510 128 14830 134
rect -1330 79 14830 128
rect -1330 56 -1091 79
rect -1330 10 -1286 56
rect -1240 33 -1091 56
rect -1045 33 -941 79
rect -895 33 -791 79
rect -745 33 -641 79
rect -595 33 -491 79
rect -445 33 -341 79
rect -295 33 -191 79
rect -145 33 -41 79
rect 5 33 109 79
rect 155 33 259 79
rect 305 33 409 79
rect 455 33 559 79
rect 605 33 709 79
rect 755 33 859 79
rect 905 33 1009 79
rect 1055 33 1159 79
rect 1205 33 1309 79
rect 1355 33 1459 79
rect 1505 33 1609 79
rect 1655 33 1759 79
rect 1805 33 1909 79
rect 1955 33 2059 79
rect 2105 33 2209 79
rect 2255 33 2359 79
rect 2405 33 2509 79
rect 2555 33 2659 79
rect 2705 33 2809 79
rect 2855 33 2959 79
rect 3005 33 3109 79
rect 3155 33 3259 79
rect 3305 33 3409 79
rect 3455 33 3559 79
rect 3605 33 3709 79
rect 3755 33 3859 79
rect 3905 33 4009 79
rect 4055 33 4159 79
rect 4205 33 4309 79
rect 4355 33 4459 79
rect 4505 33 4609 79
rect 4655 33 4759 79
rect 4805 33 4909 79
rect 4955 33 5059 79
rect 5105 33 5209 79
rect 5255 33 5359 79
rect 5405 33 5509 79
rect 5555 33 5659 79
rect 5705 33 5809 79
rect 5855 33 5959 79
rect 6005 33 6109 79
rect 6155 33 6259 79
rect 6305 33 6409 79
rect 6455 33 6559 79
rect 6605 33 6709 79
rect 6755 33 6859 79
rect 6905 33 7009 79
rect 7055 33 7159 79
rect 7205 33 7309 79
rect 7355 33 7459 79
rect 7505 33 7609 79
rect 7655 33 7759 79
rect 7805 33 7909 79
rect 7955 33 8059 79
rect 8105 33 8209 79
rect 8255 33 8359 79
rect 8405 33 8509 79
rect 8555 33 8659 79
rect 8705 33 8809 79
rect 8855 33 8959 79
rect 9005 33 9109 79
rect 9155 33 9259 79
rect 9305 33 9409 79
rect 9455 33 9559 79
rect 9605 33 9709 79
rect 9755 33 9859 79
rect 9905 33 10009 79
rect 10055 33 10159 79
rect 10205 33 10309 79
rect 10355 33 10459 79
rect 10505 33 10609 79
rect 10655 33 10759 79
rect 10805 33 10909 79
rect 10955 33 11059 79
rect 11105 33 11209 79
rect 11255 33 11359 79
rect 11405 33 11509 79
rect 11555 33 11659 79
rect 11705 33 11809 79
rect 11855 33 11959 79
rect 12005 33 12109 79
rect 12155 33 12259 79
rect 12305 33 12409 79
rect 12455 33 12559 79
rect 12605 33 12709 79
rect 12755 33 12859 79
rect 12905 33 13009 79
rect 13055 33 13159 79
rect 13205 33 13309 79
rect 13355 33 13459 79
rect 13505 33 13609 79
rect 13655 33 13759 79
rect 13805 33 13909 79
rect 13955 33 14059 79
rect 14105 33 14209 79
rect 14255 33 14359 79
rect 14405 72 14830 79
rect 14405 33 14564 72
rect -1240 26 14564 33
rect 14610 26 14714 72
rect 14760 26 14830 72
rect -1240 10 14830 26
rect -1330 -30 14830 10
rect -1330 -31 14510 -30
rect 3957 -35 14510 -31
rect 4112 -36 14510 -35
<< via1 >>
rect 6476 7032 6528 7084
rect 6475 6825 6527 6877
rect 7808 5880 7860 5932
rect 5365 5190 5417 5242
rect 5495 5191 5547 5243
rect 6692 5195 6744 5247
rect 6600 4792 6652 4844
rect 4484 4450 4536 4502
rect 5187 4352 5239 4404
rect 5513 4343 5565 4395
rect 6727 4301 6779 4353
rect 4950 4162 5002 4214
rect 7811 5744 7863 5796
rect 7811 5589 7863 5641
rect 7811 5434 7863 5486
rect 7329 4792 7381 4844
rect 7566 4796 7618 4848
rect 7796 4790 7848 4842
rect 7168 4300 7220 4352
rect 7351 4301 7403 4353
rect 7557 4301 7609 4353
rect 7704 4177 7756 4229
rect 5279 3680 5331 3732
rect 8023 2736 8075 2788
rect 8028 2577 8080 2629
rect 8012 2437 8064 2489
rect 7901 2223 7953 2275
rect 7895 1206 7947 1258
rect 8072 1207 8124 1259
rect 8241 1202 8293 1254
rect 8399 1202 8451 1254
<< metal2 >>
rect 6422 7084 6566 7134
rect 6422 7032 6476 7084
rect 6528 7032 6566 7084
rect 6422 6995 6566 7032
rect 6423 6877 6565 6995
rect 6423 6825 6475 6877
rect 6527 6825 6565 6877
rect 6423 6786 6565 6825
rect 6447 6448 6551 6786
rect -928 6344 13865 6448
rect -928 2984 -824 6344
rect 4206 6014 4377 6083
rect 7791 6039 7879 6062
rect 4308 5252 4377 6014
rect 7730 5979 7927 6039
rect 7791 5932 7879 5979
rect 7791 5930 7808 5932
rect 7792 5880 7808 5930
rect 7860 5880 7879 5932
rect 7792 5865 7879 5880
rect 7806 5805 7862 5865
rect 7795 5796 7882 5805
rect 7795 5744 7811 5796
rect 7863 5744 7882 5796
rect 7795 5729 7882 5744
rect 7806 5650 7862 5729
rect 7795 5641 7882 5650
rect 7795 5589 7811 5641
rect 7863 5589 7882 5641
rect 7795 5574 7882 5589
rect 7806 5495 7862 5574
rect 7795 5486 7882 5495
rect 7795 5434 7811 5486
rect 7863 5434 7882 5486
rect 7795 5419 7882 5434
rect 5483 5252 5569 5259
rect 4308 5243 5569 5252
rect 4308 5242 5495 5243
rect 4308 5190 5365 5242
rect 5417 5191 5495 5242
rect 5547 5191 5569 5243
rect 5417 5190 5569 5191
rect 4308 5183 5569 5190
rect 6677 5249 6750 5260
rect 7806 5249 7862 5419
rect 6677 5247 7862 5249
rect 6677 5195 6692 5247
rect 6744 5195 7862 5247
rect 6677 5193 7862 5195
rect 6677 5184 6750 5193
rect 5340 5177 5569 5183
rect 5340 5176 5512 5177
rect 5340 5175 5441 5176
rect 6573 4859 6673 4873
rect 7299 4859 7399 4875
rect 7536 4863 7636 4879
rect 7524 4859 7636 4863
rect 7766 4859 7866 4873
rect 6573 4848 7866 4859
rect 6573 4844 7566 4848
rect 6573 4792 6600 4844
rect 6652 4792 7329 4844
rect 7381 4796 7566 4844
rect 7618 4842 7866 4848
rect 7618 4796 7796 4842
rect 7381 4792 7796 4796
rect 6573 4790 7796 4792
rect 7848 4790 7866 4842
rect 6573 4777 7866 4790
rect 6573 4762 6673 4777
rect 7299 4764 7399 4777
rect 7536 4768 7636 4777
rect 7754 4775 7866 4777
rect 7766 4762 7866 4775
rect 4280 4502 4558 4523
rect 4280 4450 4484 4502
rect 4536 4450 4558 4502
rect 4280 4414 4558 4450
rect 5171 4411 5258 4413
rect 5170 4404 5258 4411
rect 5170 4399 5187 4404
rect 4946 4352 5187 4399
rect 5239 4399 5258 4404
rect 5496 4399 5582 4407
rect 5239 4395 5582 4399
rect 5239 4352 5513 4395
rect 4946 4343 5513 4352
rect 5565 4343 5582 4395
rect 4946 4339 5582 4343
rect 4946 4223 5006 4339
rect 5171 4337 5258 4339
rect 5496 4327 5582 4339
rect 6711 4355 6792 4365
rect 7152 4359 7239 4361
rect 7335 4360 7422 4362
rect 7541 4360 7628 4362
rect 7151 4355 7239 4359
rect 7334 4355 7422 4360
rect 7540 4355 7628 4360
rect 6711 4353 7769 4355
rect 6711 4301 6727 4353
rect 6779 4352 7351 4353
rect 6779 4301 7168 4352
rect 6711 4300 7168 4301
rect 7220 4301 7351 4352
rect 7403 4301 7557 4353
rect 7609 4301 7769 4353
rect 7220 4300 7769 4301
rect 6711 4299 7769 4300
rect 6711 4289 6792 4299
rect 7151 4290 7239 4299
rect 7334 4291 7422 4299
rect 7540 4291 7628 4299
rect 7152 4285 7239 4290
rect 7335 4286 7422 4291
rect 7541 4286 7628 4291
rect 7713 4239 7769 4299
rect 7685 4229 7777 4239
rect 4934 4221 5021 4223
rect 4933 4214 5021 4221
rect 4933 4162 4950 4214
rect 5002 4162 5021 4214
rect 4933 4152 5021 4162
rect 4934 4147 5021 4152
rect 7685 4177 7704 4229
rect 7756 4177 7777 4229
rect 4946 3037 5006 4147
rect 7685 4137 7777 4177
rect 7710 4029 7770 4137
rect 7779 4029 7782 4042
rect 7710 3963 7859 4029
rect 7779 3956 7782 3963
rect 5247 3732 5365 3758
rect 5247 3680 5279 3732
rect 5331 3680 5365 3732
rect 5247 3658 5365 3680
rect 12842 3729 12946 3782
rect 13761 3729 13865 6344
rect 5265 3567 5345 3658
rect 12842 3625 13865 3729
rect 5265 3487 6770 3567
rect -928 2880 32 2984
rect 6690 1819 6770 3487
rect 8011 2797 8119 3598
rect 8009 2788 8119 2797
rect 8009 2736 8023 2788
rect 8075 2736 8119 2788
rect 8009 2723 8119 2736
rect 8011 2629 8119 2723
rect 8011 2577 8028 2629
rect 8080 2577 8119 2629
rect 8011 2498 8119 2577
rect 7998 2489 8119 2498
rect 7998 2437 8012 2489
rect 8064 2437 8119 2489
rect 7998 2424 8119 2437
rect 8011 2319 8119 2424
rect 7861 2275 8119 2319
rect 7861 2223 7901 2275
rect 7953 2223 8119 2275
rect 7861 2195 8119 2223
rect 7861 2183 8015 2195
rect 8533 1819 8613 2272
rect 6690 1739 8613 1819
rect 7843 1267 7971 1290
rect 8053 1267 8146 1288
rect 8222 1267 8315 1283
rect 8380 1267 8473 1283
rect 7843 1259 8598 1267
rect 7843 1258 8072 1259
rect 7843 1206 7895 1258
rect 7947 1207 8072 1258
rect 8124 1254 8598 1259
rect 8124 1207 8241 1254
rect 7947 1206 8241 1207
rect 7843 1202 8241 1206
rect 8293 1202 8399 1254
rect 8451 1202 8598 1254
rect 7843 1197 8598 1202
rect 7843 1184 7971 1197
rect 8053 1186 8146 1197
rect 8222 1181 8315 1197
rect 8380 1181 8598 1197
rect 5026 593 5152 594
rect 5026 575 5189 593
rect 5005 519 5189 575
rect 5026 507 5189 519
rect 8528 582 8598 1181
rect 8528 512 8683 582
rect 5026 504 5175 507
rect 5119 490 5175 504
<< metal3 >>
rect 7730 5979 7927 6039
rect 7779 3989 7780 4019
use DelayCell_mag  DelayCell_mag_0
timestamp 1713971361
transform -1 0 8828 0 1 643
box 3309 -332 9664 5505
use DelayCell_mag  DelayCell_mag_1
timestamp 1713971361
transform 1 0 4062 0 -1 5952
box 3309 -332 9664 5505
use INV_2  INV_2_0
timestamp 1713185578
transform 1 0 5578 0 -1 4306
box 21 -485 1081 648
use INV_2  INV_2_1
timestamp 1713185578
transform -1 0 6684 0 -1 1123
box 21 -485 1081 648
use INV_2  INV_2_2
timestamp 1713185578
transform -1 0 7854 0 1 2284
box 21 -485 1081 648
use INV_2  INV_2_3
timestamp 1713185578
transform -1 0 7880 0 -1 1165
box 21 -485 1081 648
use INV_2  INV_2_4
timestamp 1713185578
transform -1 0 6645 0 1 2323
box 21 -485 1081 648
use INV_2  INV_2_5
timestamp 1713185578
transform 1 0 5578 0 1 5260
box 21 -485 1081 648
<< labels >>
flabel metal1 s 4567 6296 4567 6296 0 FreeSans 2500 0 0 0 VCTRL
port 1 nsew
flabel metal1 s 5215 6405 5215 6405 0 FreeSans 2500 0 0 0 VSS
port 2 nsew
flabel metal1 s 14055 1135 14055 1135 0 FreeSans 2500 0 0 0 VDD
port 3 nsew
flabel metal1 s 5144 780 5144 780 0 FreeSans 2500 0 0 0 OUTB
port 4 nsew
flabel metal1 s 5235 2311 5235 2311 0 FreeSans 2500 0 0 0 OUT
port 5 nsew
flabel metal1 s 6645 6983 6645 6983 0 FreeSans 2500 0 0 0 VCTRL2
port 6 nsew
<< end >>
