magic
tech gf180mcuC
magscale 1 10
timestamp 1714558796
<< nwell >>
rect 10048 3568 11290 3621
rect 10048 3547 12019 3568
rect 7342 3322 12019 3547
rect 7342 3245 11387 3322
rect 10048 3118 11290 3245
rect 7429 3113 11290 3118
rect 10048 2895 11290 3113
rect 279 2330 1941 2743
rect 279 2154 4730 2330
rect 140 2083 4730 2154
rect 110 2019 166 2020
rect 279 2002 4730 2083
<< nsubdiff >>
rect 11250 3385 11932 3502
rect 453 2154 822 2171
rect 140 2100 822 2154
rect 140 2083 509 2100
<< metal1 >>
rect 1453 4969 1466 5014
rect 12029 3912 12188 3981
rect 12063 3909 12188 3912
rect 11144 3419 11225 3456
rect 11190 3392 11225 3419
rect -125 1389 -47 3374
rect 48 2955 91 2994
rect 7157 2497 7274 2724
rect 12119 2627 12188 3909
rect 11927 2558 12188 2627
rect 854 2174 880 2211
rect 854 2148 882 2174
rect 854 2133 880 2148
rect 110 2019 166 2020
rect 12 1600 71 1652
rect -125 1388 28 1389
rect -125 1283 66 1388
<< metal3 >>
rect 1472 622 1530 5018
rect 1473 621 1490 622
use CLK_div_10_mag  CLK_div_10_mag_0
timestamp 1714558667
transform 1 0 0 0 1 0
box -40 0 12197 3533
use CLK_div_10_mag  CLK_div_10_mag_1
timestamp 1714558667
transform -1 0 12072 0 -1 5567
box -40 0 12197 3533
<< labels >>
flabel metal1 -78 2965 -78 2965 0 FreeSans 320 0 0 0 VSS
port 0 nsew
flabel metal1 7204 2612 7204 2612 0 FreeSans 320 0 0 0 VDD
port 1 nsew
flabel metal1 40 1612 40 1612 0 FreeSans 320 0 0 0 CLK
port 2 nsew
flabel metal1 68 2973 68 2973 0 FreeSans 320 0 0 0 Vdiv100
port 3 nsew
flabel metal1 1459 4985 1459 4985 0 FreeSans 320 0 0 0 RST
port 4 nsew
<< end >>
