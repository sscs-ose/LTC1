magic
tech gf180mcuC
magscale 1 10
timestamp 1683999746
<< nwell >>
rect -118 526 286 631
rect -32 292 31 526
<< psubdiff >>
rect -80 -95 236 -82
rect -80 -141 -67 -95
rect 223 -141 236 -95
rect -80 -154 236 -141
<< nsubdiff >>
rect -80 594 243 607
rect -80 538 -65 594
rect 229 538 243 594
rect -80 525 243 538
<< psubdiffcont >>
rect -67 -141 223 -95
<< nsubdiffcont >>
rect -65 538 229 594
<< polysilicon >>
rect 56 200 112 248
rect 18 187 112 200
rect 18 141 31 187
rect 87 141 112 187
rect 18 128 112 141
rect 56 103 112 128
<< polycontact >>
rect 31 141 87 187
<< metal1 >>
rect -118 594 286 631
rect -118 538 -65 594
rect 229 538 286 594
rect -118 525 286 538
rect -32 292 31 525
rect -118 187 93 200
rect -118 141 31 187
rect 87 141 93 187
rect -118 128 93 141
rect 139 189 202 450
rect 139 131 286 189
rect -34 -69 33 60
rect 139 14 202 131
rect -118 -95 286 -69
rect -118 -141 -67 -95
rect 223 -141 286 -95
rect -118 -175 286 -141
use nmos_3p3_DDNVWA  nmos_3p3_DDNVWA_0
timestamp 1683999746
transform 1 0 84 0 1 37
box -144 -97 144 97
use pmos_3p3_MQGBLR  pmos_3p3_MQGBLR_0
timestamp 1683999746
transform 1 0 84 0 1 372
box -202 -210 202 210
<< labels >>
flabel nsubdiffcont 82 566 82 566 0 FreeSans 640 0 0 0 VDD
port 0 nsew
flabel psubdiffcont 80 -120 80 -120 0 FreeSans 640 0 0 0 VSS
port 1 nsew
flabel metal1 -106 158 -106 158 0 FreeSans 640 0 0 0 IN
port 2 nsew
flabel metal1 276 159 276 159 0 FreeSans 640 0 0 0 OUT
port 3 nsew
<< end >>
