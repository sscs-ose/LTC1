magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1052 -1316 1052 1316
<< metal2 >>
rect -52 311 52 316
rect -52 283 -47 311
rect -19 283 19 311
rect 47 283 52 311
rect -52 245 52 283
rect -52 217 -47 245
rect -19 217 19 245
rect 47 217 52 245
rect -52 179 52 217
rect -52 151 -47 179
rect -19 151 19 179
rect 47 151 52 179
rect -52 113 52 151
rect -52 85 -47 113
rect -19 85 19 113
rect 47 85 52 113
rect -52 47 52 85
rect -52 19 -47 47
rect -19 19 19 47
rect 47 19 52 47
rect -52 -19 52 19
rect -52 -47 -47 -19
rect -19 -47 19 -19
rect 47 -47 52 -19
rect -52 -85 52 -47
rect -52 -113 -47 -85
rect -19 -113 19 -85
rect 47 -113 52 -85
rect -52 -151 52 -113
rect -52 -179 -47 -151
rect -19 -179 19 -151
rect 47 -179 52 -151
rect -52 -217 52 -179
rect -52 -245 -47 -217
rect -19 -245 19 -217
rect 47 -245 52 -217
rect -52 -283 52 -245
rect -52 -311 -47 -283
rect -19 -311 19 -283
rect 47 -311 52 -283
rect -52 -316 52 -311
<< via2 >>
rect -47 283 -19 311
rect 19 283 47 311
rect -47 217 -19 245
rect 19 217 47 245
rect -47 151 -19 179
rect 19 151 47 179
rect -47 85 -19 113
rect 19 85 47 113
rect -47 19 -19 47
rect 19 19 47 47
rect -47 -47 -19 -19
rect 19 -47 47 -19
rect -47 -113 -19 -85
rect 19 -113 47 -85
rect -47 -179 -19 -151
rect 19 -179 47 -151
rect -47 -245 -19 -217
rect 19 -245 47 -217
rect -47 -311 -19 -283
rect 19 -311 47 -283
<< metal3 >>
rect -52 311 52 316
rect -52 283 -47 311
rect -19 283 19 311
rect 47 283 52 311
rect -52 245 52 283
rect -52 217 -47 245
rect -19 217 19 245
rect 47 217 52 245
rect -52 179 52 217
rect -52 151 -47 179
rect -19 151 19 179
rect 47 151 52 179
rect -52 113 52 151
rect -52 85 -47 113
rect -19 85 19 113
rect 47 85 52 113
rect -52 47 52 85
rect -52 19 -47 47
rect -19 19 19 47
rect 47 19 52 47
rect -52 -19 52 19
rect -52 -47 -47 -19
rect -19 -47 19 -19
rect 47 -47 52 -19
rect -52 -85 52 -47
rect -52 -113 -47 -85
rect -19 -113 19 -85
rect 47 -113 52 -85
rect -52 -151 52 -113
rect -52 -179 -47 -151
rect -19 -179 19 -151
rect 47 -179 52 -151
rect -52 -217 52 -179
rect -52 -245 -47 -217
rect -19 -245 19 -217
rect 47 -245 52 -217
rect -52 -283 52 -245
rect -52 -311 -47 -283
rect -19 -311 19 -283
rect 47 -311 52 -283
rect -52 -316 52 -311
<< end >>
