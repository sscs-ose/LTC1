magic
tech gf180mcuD
magscale 1 10
timestamp 1713971361
<< checkpaint >>
rect -2791 -2040 7078 4784
<< pwell >>
rect -496 30 1706 2551
rect 1759 316 5030 2395
<< ndiff >>
rect 92 739 105 798
<< psubdiff >>
rect 1693 2600 1777 2602
rect -541 2580 1777 2600
rect -541 2579 134 2580
rect -541 2533 -521 2579
rect -475 2534 134 2579
rect 180 2534 284 2580
rect 330 2534 434 2580
rect 480 2534 584 2580
rect 630 2534 734 2580
rect 780 2534 884 2580
rect 930 2534 1034 2580
rect 1080 2534 1184 2580
rect 1230 2534 1334 2580
rect 1380 2534 1777 2580
rect -475 2533 1777 2534
rect -541 2530 1777 2533
rect -541 2516 1709 2530
rect -541 2391 -457 2516
rect -541 2345 -525 2391
rect -479 2345 -457 2391
rect -541 2241 -457 2345
rect 1693 2484 1709 2516
rect 1755 2484 1777 2530
rect 1693 2422 1777 2484
rect 1693 2399 5075 2422
rect 1693 2398 2173 2399
rect 1693 2380 1860 2398
rect 1693 2334 1709 2380
rect 1755 2352 1860 2380
rect 1906 2352 1964 2398
rect 2010 2352 2069 2398
rect 2115 2353 2173 2398
rect 2219 2353 2323 2399
rect 2369 2353 2473 2399
rect 2519 2353 2623 2399
rect 2669 2353 2773 2399
rect 2819 2353 2923 2399
rect 2969 2353 3073 2399
rect 3119 2353 3223 2399
rect 3269 2353 3373 2399
rect 3419 2353 3523 2399
rect 3569 2353 3673 2399
rect 3719 2353 3823 2399
rect 3869 2353 3973 2399
rect 4019 2353 4123 2399
rect 4169 2353 4273 2399
rect 4319 2353 4423 2399
rect 4469 2353 4573 2399
rect 4619 2383 5075 2399
rect 4619 2353 5010 2383
rect 2115 2352 5010 2353
rect 1755 2338 5010 2352
rect 1755 2334 1777 2338
rect -541 2195 -525 2241
rect -479 2195 -457 2241
rect -541 2091 -457 2195
rect -541 2045 -525 2091
rect -479 2045 -457 2091
rect 1693 2230 1777 2334
rect 1693 2184 1709 2230
rect 1755 2184 1777 2230
rect 4991 2337 5010 2338
rect 5056 2337 5075 2383
rect 4991 2233 5075 2337
rect 1693 2080 1777 2184
rect 4991 2187 5010 2233
rect 5056 2187 5075 2233
rect 4991 2083 5075 2187
rect -541 1941 -457 2045
rect 1693 2034 1709 2080
rect 1755 2034 1777 2080
rect -541 1895 -525 1941
rect -479 1895 -457 1941
rect -541 1791 -457 1895
rect -541 1745 -525 1791
rect -479 1745 -457 1791
rect 1693 1930 1777 2034
rect 4991 2037 5010 2083
rect 5056 2037 5075 2083
rect 1693 1884 1709 1930
rect 1755 1884 1777 1930
rect -541 1641 -457 1745
rect 1693 1780 1777 1884
rect 1693 1734 1709 1780
rect 1755 1734 1777 1780
rect -541 1595 -525 1641
rect -479 1595 -457 1641
rect -541 1491 -457 1595
rect 1693 1630 1777 1734
rect 1693 1584 1709 1630
rect 1755 1584 1777 1630
rect -541 1445 -525 1491
rect -479 1445 -457 1491
rect -541 1341 -457 1445
rect -541 1295 -525 1341
rect -479 1295 -457 1341
rect -541 1191 -457 1295
rect 1693 1480 1777 1584
rect 1693 1434 1709 1480
rect 1755 1434 1777 1480
rect 1693 1330 1777 1434
rect 1693 1284 1709 1330
rect 1755 1284 1777 1330
rect -541 1145 -525 1191
rect -479 1145 -457 1191
rect 1693 1180 1777 1284
rect -541 1041 -457 1145
rect -541 995 -525 1041
rect -479 995 -457 1041
rect -541 891 -457 995
rect 1693 1134 1709 1180
rect 1755 1134 1777 1180
rect -541 845 -525 891
rect -479 845 -457 891
rect -541 741 -457 845
rect 1693 1030 1777 1134
rect 1693 984 1709 1030
rect 1755 984 1777 1030
rect 1693 880 1777 984
rect 1693 834 1709 880
rect 1755 834 1777 880
rect -541 695 -525 741
rect -479 695 -457 741
rect 1693 730 1777 834
rect 4991 1933 5075 2037
rect 4991 1887 5010 1933
rect 5056 1887 5075 1933
rect 4991 1783 5075 1887
rect 4991 1737 5010 1783
rect 5056 1737 5075 1783
rect 4991 1633 5075 1737
rect 4991 1587 5010 1633
rect 5056 1587 5075 1633
rect 4991 1483 5075 1587
rect 4991 1437 5010 1483
rect 5056 1437 5075 1483
rect 4991 1333 5075 1437
rect 4991 1287 5010 1333
rect 5056 1287 5075 1333
rect 4991 1183 5075 1287
rect 4991 1137 5010 1183
rect 5056 1137 5075 1183
rect 4991 1033 5075 1137
rect 4991 987 5010 1033
rect 5056 987 5075 1033
rect 4991 883 5075 987
rect 4991 837 5010 883
rect 5056 837 5075 883
rect -541 591 -457 695
rect -541 545 -525 591
rect -479 545 -457 591
rect 1693 684 1709 730
rect 1755 684 1777 730
rect -541 441 -457 545
rect -541 395 -525 441
rect -479 395 -457 441
rect 1693 580 1777 684
rect 4991 733 5075 837
rect 4991 687 5010 733
rect 5056 687 5075 733
rect 1693 534 1709 580
rect 1755 534 1777 580
rect -541 291 -457 395
rect 1693 430 1777 534
rect 1693 384 1709 430
rect 1755 384 1777 430
rect 1693 343 1777 384
rect 4991 583 5075 687
rect 4991 537 5010 583
rect 5056 537 5075 583
rect 4991 433 5075 537
rect 4991 387 5010 433
rect 5056 387 5075 433
rect 4991 343 5075 387
rect -541 245 -525 291
rect -479 245 -457 291
rect -541 141 -457 245
rect 1693 326 5075 343
rect 1693 325 2278 326
rect 1693 279 1730 325
rect 1776 279 1840 325
rect 1886 279 1950 325
rect 1996 279 2059 325
rect 2105 279 2169 325
rect 2215 280 2278 325
rect 2324 280 2428 326
rect 2474 280 2578 326
rect 2624 280 2728 326
rect 2774 280 2878 326
rect 2924 280 3028 326
rect 3074 280 3178 326
rect 3224 280 3328 326
rect 3374 280 3478 326
rect 3524 280 3628 326
rect 3674 280 3778 326
rect 3824 280 3928 326
rect 3974 280 4078 326
rect 4124 280 4228 326
rect 4274 280 4378 326
rect 4424 280 4528 326
rect 4574 325 4948 326
rect 4574 323 4801 325
rect 4574 280 4660 323
rect 2215 279 4660 280
rect 1693 277 4660 279
rect 4706 279 4801 323
rect 4847 280 4948 325
rect 4994 280 5075 326
rect 4847 279 5075 280
rect 4706 277 5075 279
rect 1693 259 5075 277
rect 1693 176 1785 259
rect -541 95 -525 141
rect -479 95 -457 141
rect -541 46 -457 95
rect 1693 130 1710 176
rect 1756 130 1785 176
rect 1693 46 1785 130
rect -541 30 1785 46
rect -541 -16 -158 30
rect -112 -16 -8 30
rect 38 -16 142 30
rect 188 -16 292 30
rect 338 -16 442 30
rect 488 -16 592 30
rect 638 -16 742 30
rect 788 -16 892 30
rect 938 -16 1042 30
rect 1088 -16 1192 30
rect 1238 -16 1342 30
rect 1388 -16 1483 30
rect 1529 -16 1673 30
rect 1719 -16 1785 30
rect -541 -33 1785 -16
<< psubdiffcont >>
rect -521 2533 -475 2579
rect 134 2534 180 2580
rect 284 2534 330 2580
rect 434 2534 480 2580
rect 584 2534 630 2580
rect 734 2534 780 2580
rect 884 2534 930 2580
rect 1034 2534 1080 2580
rect 1184 2534 1230 2580
rect 1334 2534 1380 2580
rect -525 2345 -479 2391
rect 1709 2484 1755 2530
rect 1709 2334 1755 2380
rect 1860 2352 1906 2398
rect 1964 2352 2010 2398
rect 2069 2352 2115 2398
rect 2173 2353 2219 2399
rect 2323 2353 2369 2399
rect 2473 2353 2519 2399
rect 2623 2353 2669 2399
rect 2773 2353 2819 2399
rect 2923 2353 2969 2399
rect 3073 2353 3119 2399
rect 3223 2353 3269 2399
rect 3373 2353 3419 2399
rect 3523 2353 3569 2399
rect 3673 2353 3719 2399
rect 3823 2353 3869 2399
rect 3973 2353 4019 2399
rect 4123 2353 4169 2399
rect 4273 2353 4319 2399
rect 4423 2353 4469 2399
rect 4573 2353 4619 2399
rect -525 2195 -479 2241
rect -525 2045 -479 2091
rect 1709 2184 1755 2230
rect 5010 2337 5056 2383
rect 5010 2187 5056 2233
rect 1709 2034 1755 2080
rect -525 1895 -479 1941
rect -525 1745 -479 1791
rect 5010 2037 5056 2083
rect 1709 1884 1755 1930
rect 1709 1734 1755 1780
rect -525 1595 -479 1641
rect 1709 1584 1755 1630
rect -525 1445 -479 1491
rect -525 1295 -479 1341
rect 1709 1434 1755 1480
rect 1709 1284 1755 1330
rect -525 1145 -479 1191
rect -525 995 -479 1041
rect 1709 1134 1755 1180
rect -525 845 -479 891
rect 1709 984 1755 1030
rect 1709 834 1755 880
rect -525 695 -479 741
rect 5010 1887 5056 1933
rect 5010 1737 5056 1783
rect 5010 1587 5056 1633
rect 5010 1437 5056 1483
rect 5010 1287 5056 1333
rect 5010 1137 5056 1183
rect 5010 987 5056 1033
rect 5010 837 5056 883
rect -525 545 -479 591
rect 1709 684 1755 730
rect -525 395 -479 441
rect 5010 687 5056 733
rect 1709 534 1755 580
rect 1709 384 1755 430
rect 5010 537 5056 583
rect 5010 387 5056 433
rect -525 245 -479 291
rect 1730 279 1776 325
rect 1840 279 1886 325
rect 1950 279 1996 325
rect 2059 279 2105 325
rect 2169 279 2215 325
rect 2278 280 2324 326
rect 2428 280 2474 326
rect 2578 280 2624 326
rect 2728 280 2774 326
rect 2878 280 2924 326
rect 3028 280 3074 326
rect 3178 280 3224 326
rect 3328 280 3374 326
rect 3478 280 3524 326
rect 3628 280 3674 326
rect 3778 280 3824 326
rect 3928 280 3974 326
rect 4078 280 4124 326
rect 4228 280 4274 326
rect 4378 280 4424 326
rect 4528 280 4574 326
rect 4660 277 4706 323
rect 4801 279 4847 325
rect 4948 280 4994 326
rect -525 95 -479 141
rect 1710 130 1756 176
rect -158 -16 -112 30
rect -8 -16 38 30
rect 142 -16 188 30
rect 292 -16 338 30
rect 442 -16 488 30
rect 592 -16 638 30
rect 742 -16 788 30
rect 892 -16 938 30
rect 1042 -16 1088 30
rect 1192 -16 1238 30
rect 1342 -16 1388 30
rect 1483 -16 1529 30
rect 1673 -16 1719 30
<< polysilicon >>
rect 116 2246 284 2274
rect 116 2200 176 2246
rect 222 2200 284 2246
rect -286 2177 -118 2191
rect -286 2131 -234 2177
rect -188 2131 -118 2177
rect -286 2080 -118 2131
rect 116 2125 284 2200
rect 932 2241 1100 2273
rect 932 2195 985 2241
rect 1031 2195 1100 2241
rect 932 2124 1100 2195
rect 1333 2179 1501 2193
rect 1333 2133 1385 2179
rect 1431 2133 1501 2179
rect 1333 2102 1501 2133
rect 1945 2180 2113 2194
rect 1945 2134 1997 2180
rect 2043 2134 2113 2180
rect 1945 2082 2113 2134
rect 4651 2178 4819 2192
rect 4651 2132 4703 2178
rect 4749 2132 4819 2178
rect 4651 2081 4819 2132
rect -286 1936 -118 1980
rect 388 1878 555 1950
rect 116 1837 283 1859
rect 116 1791 178 1837
rect 224 1791 283 1837
rect 388 1832 439 1878
rect 485 1832 555 1878
rect 388 1805 555 1832
rect 659 1876 827 1943
rect 659 1830 723 1876
rect 769 1830 827 1876
rect 1945 1938 2113 1983
rect 659 1803 827 1830
rect 932 1832 1100 1861
rect -286 1743 -118 1757
rect -286 1697 -234 1743
rect -188 1697 -118 1743
rect -286 1646 -118 1697
rect 116 1675 283 1791
rect 932 1786 987 1832
rect 1033 1786 1100 1832
rect 932 1683 1100 1786
rect 2345 1889 2513 1945
rect 1332 1744 1500 1758
rect 1332 1698 1384 1744
rect 1430 1698 1500 1744
rect 1332 1647 1500 1698
rect 1945 1851 2113 1865
rect 1945 1805 1997 1851
rect 2043 1805 2113 1851
rect 1945 1753 2113 1805
rect 2345 1843 2396 1889
rect 2442 1843 2513 1889
rect 1945 1609 2113 1654
rect -286 1502 -118 1546
rect 388 1420 556 1504
rect 388 1374 447 1420
rect 493 1374 556 1420
rect -288 1347 -120 1361
rect -288 1301 -236 1347
rect -190 1301 -120 1347
rect -288 1250 -120 1301
rect 388 1286 556 1374
rect 660 1425 828 1510
rect 1332 1503 1500 1547
rect 660 1379 713 1425
rect 759 1379 828 1425
rect 660 1292 828 1379
rect 2345 1579 2513 1843
rect 2345 1533 2406 1579
rect 2452 1533 2513 1579
rect 1332 1347 1500 1361
rect 1332 1301 1384 1347
rect 1430 1301 1500 1347
rect 1332 1250 1500 1301
rect 1945 1516 2113 1530
rect 1945 1470 1997 1516
rect 2043 1470 2113 1516
rect 1945 1418 2113 1470
rect 1945 1274 2113 1319
rect 2345 1226 2513 1533
rect -288 1106 -120 1150
rect 116 1048 284 1112
rect 116 1002 181 1048
rect 227 1002 284 1048
rect 116 983 284 1002
rect 932 1039 1100 1112
rect 1332 1106 1500 1150
rect 932 993 988 1039
rect 1034 993 1100 1039
rect 388 955 556 984
rect -290 911 -122 925
rect -290 865 -238 911
rect -192 865 -122 911
rect -290 814 -122 865
rect 388 909 449 955
rect 495 909 556 955
rect 388 850 556 909
rect 659 956 828 976
rect 932 965 1100 993
rect 1945 1180 2113 1194
rect 1945 1134 1997 1180
rect 2043 1134 2113 1180
rect 1945 1082 2113 1134
rect 2345 1180 2409 1226
rect 2455 1180 2513 1226
rect 659 910 729 956
rect 775 910 828 956
rect 659 841 828 910
rect 1332 911 1500 925
rect 1332 865 1384 911
rect 1430 865 1500 911
rect 1332 814 1500 865
rect 1945 938 2113 983
rect 2345 891 2513 1180
rect 1945 844 2113 858
rect 1945 798 1997 844
rect 2043 798 2113 844
rect 1945 746 2113 798
rect 2345 845 2409 891
rect 2455 845 2513 891
rect 2345 782 2513 845
rect 2617 1888 2785 1948
rect 2617 1842 2671 1888
rect 2717 1842 2785 1888
rect 2617 1578 2785 1842
rect 2617 1532 2681 1578
rect 2727 1532 2785 1578
rect 2617 1225 2785 1532
rect 2617 1179 2684 1225
rect 2730 1179 2785 1225
rect 2617 890 2785 1179
rect 2617 844 2684 890
rect 2730 844 2785 890
rect 2617 785 2785 844
rect 2889 1888 3057 1951
rect 2889 1842 2937 1888
rect 2983 1842 3057 1888
rect 2889 1578 3057 1842
rect 2889 1532 2947 1578
rect 2993 1532 3057 1578
rect 2889 1225 3057 1532
rect 2889 1179 2950 1225
rect 2996 1179 3057 1225
rect 2889 890 3057 1179
rect 2889 844 2950 890
rect 2996 844 3057 890
rect 2889 788 3057 844
rect 3161 1888 3329 1950
rect 3161 1842 3210 1888
rect 3256 1842 3329 1888
rect 3161 1578 3329 1842
rect 3161 1532 3220 1578
rect 3266 1532 3329 1578
rect 3161 1225 3329 1532
rect 3161 1179 3223 1225
rect 3269 1179 3329 1225
rect 3161 890 3329 1179
rect 3161 844 3223 890
rect 3269 844 3329 890
rect 3161 787 3329 844
rect 3433 1887 3601 1950
rect 3433 1841 3482 1887
rect 3528 1841 3601 1887
rect 3433 1577 3601 1841
rect 3433 1531 3492 1577
rect 3538 1531 3601 1577
rect 3433 1224 3601 1531
rect 3433 1178 3495 1224
rect 3541 1178 3601 1224
rect 3433 889 3601 1178
rect 3433 843 3495 889
rect 3541 843 3601 889
rect 3433 787 3601 843
rect 3705 1887 3873 1948
rect 3705 1841 3752 1887
rect 3798 1841 3873 1887
rect 3705 1577 3873 1841
rect 3705 1531 3762 1577
rect 3808 1531 3873 1577
rect 3705 1224 3873 1531
rect 3705 1178 3765 1224
rect 3811 1178 3873 1224
rect 3705 889 3873 1178
rect 3705 843 3765 889
rect 3811 843 3873 889
rect 3705 785 3873 843
rect 3977 1889 4145 1947
rect 3977 1843 4021 1889
rect 4067 1843 4145 1889
rect 3977 1579 4145 1843
rect 3977 1533 4031 1579
rect 4077 1533 4145 1579
rect 3977 1226 4145 1533
rect 3977 1180 4034 1226
rect 4080 1180 4145 1226
rect 3977 891 4145 1180
rect 3977 845 4034 891
rect 4080 845 4145 891
rect 3977 784 4145 845
rect 4249 1888 4417 1948
rect 4651 1937 4819 1981
rect 4249 1842 4324 1888
rect 4370 1842 4417 1888
rect 4249 1578 4417 1842
rect 4650 1850 4818 1864
rect 4650 1804 4702 1850
rect 4748 1804 4818 1850
rect 4650 1753 4818 1804
rect 4650 1609 4818 1653
rect 4249 1532 4334 1578
rect 4380 1532 4417 1578
rect 4249 1225 4417 1532
rect 4651 1514 4819 1528
rect 4651 1468 4703 1514
rect 4749 1468 4819 1514
rect 4651 1417 4819 1468
rect 4651 1273 4819 1317
rect 4249 1179 4337 1225
rect 4383 1179 4417 1225
rect 4249 890 4417 1179
rect 4649 1179 4817 1193
rect 4649 1133 4701 1179
rect 4747 1133 4817 1179
rect 4649 1082 4817 1133
rect 4649 938 4817 982
rect 4249 844 4337 890
rect 4383 844 4417 890
rect 4249 785 4417 844
rect 4650 843 4818 857
rect 4650 797 4702 843
rect 4748 797 4818 843
rect 4650 746 4818 797
rect -290 670 -122 714
rect 116 628 284 673
rect 116 582 170 628
rect 216 582 284 628
rect 932 632 1100 674
rect 1332 670 1500 714
rect 116 553 284 582
rect 388 572 555 590
rect -290 535 -122 549
rect -290 489 -238 535
rect -192 489 -122 535
rect -290 438 -122 489
rect 388 526 437 572
rect 483 526 555 572
rect 388 472 555 526
rect 660 583 828 597
rect 660 537 715 583
rect 761 537 828 583
rect 932 586 998 632
rect 1044 586 1100 632
rect 932 554 1100 586
rect 1945 602 2113 647
rect 4650 602 4818 646
rect 660 476 828 537
rect 1332 536 1500 550
rect 1332 490 1384 536
rect 1430 490 1500 536
rect 1332 439 1500 490
rect -290 294 -122 338
rect 115 235 284 303
rect 115 189 173 235
rect 219 189 284 235
rect 115 171 284 189
rect 932 235 1100 298
rect 1332 295 1500 339
rect 932 189 990 235
rect 1036 189 1100 235
rect 932 174 1100 189
<< polycontact >>
rect 176 2200 222 2246
rect -234 2131 -188 2177
rect 985 2195 1031 2241
rect 1385 2133 1431 2179
rect 1997 2134 2043 2180
rect 4703 2132 4749 2178
rect 178 1791 224 1837
rect 439 1832 485 1878
rect 723 1830 769 1876
rect -234 1697 -188 1743
rect 987 1786 1033 1832
rect 1384 1698 1430 1744
rect 1997 1805 2043 1851
rect 2396 1843 2442 1889
rect 447 1374 493 1420
rect -236 1301 -190 1347
rect 713 1379 759 1425
rect 2406 1533 2452 1579
rect 1384 1301 1430 1347
rect 1997 1470 2043 1516
rect 181 1002 227 1048
rect 988 993 1034 1039
rect -238 865 -192 911
rect 449 909 495 955
rect 1997 1134 2043 1180
rect 2409 1180 2455 1226
rect 729 910 775 956
rect 1384 865 1430 911
rect 1997 798 2043 844
rect 2409 845 2455 891
rect 2671 1842 2717 1888
rect 2681 1532 2727 1578
rect 2684 1179 2730 1225
rect 2684 844 2730 890
rect 2937 1842 2983 1888
rect 2947 1532 2993 1578
rect 2950 1179 2996 1225
rect 2950 844 2996 890
rect 3210 1842 3256 1888
rect 3220 1532 3266 1578
rect 3223 1179 3269 1225
rect 3223 844 3269 890
rect 3482 1841 3528 1887
rect 3492 1531 3538 1577
rect 3495 1178 3541 1224
rect 3495 843 3541 889
rect 3752 1841 3798 1887
rect 3762 1531 3808 1577
rect 3765 1178 3811 1224
rect 3765 843 3811 889
rect 4021 1843 4067 1889
rect 4031 1533 4077 1579
rect 4034 1180 4080 1226
rect 4034 845 4080 891
rect 4324 1842 4370 1888
rect 4702 1804 4748 1850
rect 4334 1532 4380 1578
rect 4703 1468 4749 1514
rect 4337 1179 4383 1225
rect 4701 1133 4747 1179
rect 4337 844 4383 890
rect 4702 797 4748 843
rect 170 582 216 628
rect -238 489 -192 535
rect 437 526 483 572
rect 715 537 761 583
rect 998 586 1044 632
rect 1384 490 1430 536
rect 173 189 219 235
rect 990 189 1036 235
<< metal1 >>
rect 289 2716 375 2748
rect 289 2664 308 2716
rect 360 2664 375 2716
rect 1251 2739 1345 2784
rect 1251 2687 1274 2739
rect 1326 2687 1345 2739
rect 1251 2677 1345 2687
rect 4169 2726 4394 2755
rect 4169 2725 4324 2726
rect 289 2655 375 2664
rect 4169 2673 4189 2725
rect 4241 2674 4324 2725
rect 4376 2674 4394 2726
rect 4241 2673 4394 2674
rect -554 2580 1793 2602
rect -554 2579 134 2580
rect -554 2533 -521 2579
rect -475 2534 134 2579
rect 180 2534 284 2580
rect 330 2534 434 2580
rect 480 2534 584 2580
rect 630 2534 734 2580
rect 780 2534 884 2580
rect 930 2534 1034 2580
rect 1080 2534 1184 2580
rect 1230 2534 1334 2580
rect 1380 2534 1793 2580
rect 4169 2599 4394 2673
rect 4169 2547 4194 2599
rect 4246 2596 4394 2599
rect 4246 2547 4321 2596
rect 4169 2544 4321 2547
rect 4373 2544 4394 2596
rect 4169 2536 4394 2544
rect -475 2533 1793 2534
rect -554 2530 1793 2533
rect -554 2511 1709 2530
rect -554 2391 -441 2511
rect 1680 2484 1709 2511
rect 1755 2484 1793 2530
rect 1680 2425 1793 2484
rect -554 2345 -525 2391
rect -479 2345 -441 2391
rect -707 2277 -626 2292
rect -770 2275 -626 2277
rect -770 2223 -693 2275
rect -641 2223 -626 2275
rect -770 2221 -626 2223
rect -707 2206 -626 2221
rect -554 2241 -441 2345
rect -101 2406 -21 2415
rect 566 2406 631 2409
rect 1265 2406 1336 2420
rect -101 2403 1336 2406
rect -101 2351 -86 2403
rect -34 2351 572 2403
rect 624 2351 1278 2403
rect 1330 2351 1336 2403
rect -101 2348 1336 2351
rect -101 2344 -21 2348
rect 566 2344 631 2348
rect 1265 2334 1336 2348
rect 1680 2399 5078 2425
rect 1680 2398 2173 2399
rect 1680 2380 1860 2398
rect 1680 2334 1709 2380
rect 1755 2352 1860 2380
rect 1906 2352 1964 2398
rect 2010 2352 2069 2398
rect 2115 2353 2173 2398
rect 2219 2353 2323 2399
rect 2369 2353 2473 2399
rect 2519 2353 2623 2399
rect 2669 2353 2773 2399
rect 2819 2353 2923 2399
rect 2969 2353 3073 2399
rect 3119 2353 3223 2399
rect 3269 2353 3373 2399
rect 3419 2353 3523 2399
rect 3569 2353 3673 2399
rect 3719 2353 3823 2399
rect 3869 2353 3973 2399
rect 4019 2353 4123 2399
rect 4169 2353 4273 2399
rect 4319 2353 4423 2399
rect 4469 2353 4573 2399
rect 4619 2383 5078 2399
rect 4619 2353 5010 2383
rect 2115 2352 5010 2353
rect 1755 2337 5010 2352
rect 5056 2337 5078 2383
rect 1755 2334 5078 2337
rect 1680 2333 5078 2334
rect -554 2195 -525 2241
rect -479 2195 -441 2241
rect -554 2190 -441 2195
rect 155 2250 242 2268
rect 155 2198 173 2250
rect 225 2198 242 2250
rect -554 2177 -44 2190
rect 155 2180 242 2198
rect 964 2245 1051 2263
rect 964 2193 982 2245
rect 1034 2193 1051 2245
rect -554 2140 -234 2177
rect -554 2091 -441 2140
rect -554 2045 -525 2091
rect -479 2045 -441 2091
rect -554 1941 -441 2045
rect -361 1980 -314 2140
rect -246 2131 -234 2140
rect -188 2140 -44 2177
rect -188 2131 -176 2140
rect -246 2119 -176 2131
rect -91 1982 -44 2140
rect 312 2130 903 2178
rect 964 2175 1051 2193
rect 1680 2230 1793 2333
rect 2313 2235 2475 2333
rect 2729 2235 2891 2333
rect 3069 2235 3231 2333
rect 3608 2235 3770 2333
rect 4154 2235 4316 2333
rect 1680 2192 1709 2230
rect 1258 2184 1709 2192
rect 1755 2184 1793 2230
rect 2270 2191 4493 2235
rect 4986 2233 5078 2333
rect 4986 2191 5010 2233
rect 1258 2179 1793 2184
rect 26 2061 104 2083
rect 313 2080 359 2130
rect 26 2009 38 2061
rect 90 2009 104 2061
rect 26 1981 104 2009
rect -554 1895 -525 1941
rect -479 1895 -441 1941
rect -554 1791 -441 1895
rect -554 1745 -525 1791
rect -479 1756 -441 1791
rect 157 1841 244 1859
rect 157 1789 175 1841
rect 227 1789 244 1841
rect 157 1771 244 1789
rect 312 1765 359 2080
rect 585 2061 655 2083
rect 585 2009 589 2061
rect 641 2009 655 2061
rect 585 1985 655 2009
rect 419 1882 505 1900
rect 419 1830 436 1882
rect 488 1830 505 1882
rect 419 1812 505 1830
rect 702 1880 789 1898
rect 702 1828 720 1880
rect 772 1828 789 1880
rect 702 1811 789 1828
rect 856 1765 903 2130
rect 1258 2142 1385 2179
rect 1123 2061 1203 2084
rect 1123 2009 1138 2061
rect 1190 2009 1203 2061
rect 1123 1981 1203 2009
rect 1258 1982 1305 2142
rect 1373 2133 1385 2142
rect 1431 2144 1793 2179
rect 1431 2142 1575 2144
rect 1431 2133 1443 2142
rect 1373 2121 1443 2133
rect 1528 1984 1575 2142
rect 1680 2080 1793 2144
rect 1680 2034 1709 2080
rect 1755 2034 1793 2080
rect 1680 1997 1793 2034
rect 1870 2180 2187 2190
rect 1870 2143 1997 2180
rect 1870 1997 1917 2143
rect 1985 2134 1997 2143
rect 2043 2143 2187 2180
rect 2043 2134 2055 2143
rect 1985 2122 2055 2134
rect 2140 2096 2187 2143
rect 2115 2081 2187 2096
rect 2270 2187 5010 2191
rect 5056 2187 5078 2233
rect 2270 2178 5078 2187
rect 2270 2160 4703 2178
rect 2115 2069 2188 2081
rect 2115 2019 2187 2069
rect 2115 1997 2188 2019
rect 1680 1969 2188 1997
rect 2270 1969 2316 2160
rect 1680 1930 2316 1969
rect 1680 1884 1709 1930
rect 1755 1884 2316 1930
rect 1680 1858 2316 1884
rect 1680 1857 2187 1858
rect 966 1836 1053 1854
rect 966 1784 984 1836
rect 1036 1784 1053 1836
rect 966 1766 1053 1784
rect 1680 1780 1793 1857
rect -479 1745 -44 1756
rect -554 1743 -44 1745
rect -554 1707 -234 1743
rect -554 1641 -441 1707
rect -554 1595 -525 1641
rect -479 1595 -441 1641
rect -554 1491 -441 1595
rect -361 1706 -234 1707
rect -361 1546 -314 1706
rect -246 1697 -234 1706
rect -188 1706 -44 1743
rect -188 1697 -176 1706
rect -246 1685 -176 1697
rect -91 1548 -44 1706
rect 312 1719 903 1765
rect 1680 1756 1709 1780
rect 1532 1754 1709 1756
rect 32 1625 105 1647
rect 32 1573 38 1625
rect 90 1573 105 1625
rect -554 1445 -525 1491
rect -479 1445 -441 1491
rect -554 1360 -441 1445
rect -554 1347 -46 1360
rect -554 1341 -236 1347
rect -554 1295 -525 1341
rect -479 1311 -236 1341
rect -479 1295 -441 1311
rect -554 1191 -441 1295
rect -554 1145 -525 1191
rect -479 1145 -441 1191
rect -363 1310 -236 1311
rect -363 1150 -316 1310
rect -248 1301 -236 1310
rect -190 1310 -46 1347
rect -190 1301 -178 1310
rect -248 1289 -178 1301
rect -93 1152 -46 1310
rect 32 1250 105 1573
rect 31 1228 105 1250
rect 31 1176 37 1228
rect 89 1176 105 1228
rect 31 1157 105 1176
rect 32 1147 105 1157
rect -554 1041 -441 1145
rect 312 1075 359 1719
rect 569 1625 657 1646
rect 569 1573 589 1625
rect 641 1573 657 1625
rect 569 1546 657 1573
rect 426 1424 513 1442
rect 426 1372 444 1424
rect 496 1372 513 1424
rect 426 1354 513 1372
rect 692 1429 779 1447
rect 692 1377 710 1429
rect 762 1377 779 1429
rect 692 1359 779 1377
rect 585 1229 655 1249
rect 585 1177 589 1229
rect 641 1177 655 1229
rect 585 1150 655 1177
rect 856 1075 903 1719
rect 1257 1744 1709 1754
rect 1257 1707 1384 1744
rect 1123 1625 1195 1652
rect 1123 1573 1138 1625
rect 1190 1573 1195 1625
rect 1123 1249 1195 1573
rect 1257 1547 1304 1707
rect 1372 1698 1384 1707
rect 1430 1734 1709 1744
rect 1755 1734 1793 1780
rect 1430 1710 1793 1734
rect 1430 1707 1574 1710
rect 1430 1698 1442 1707
rect 1372 1686 1442 1698
rect 1527 1645 1574 1707
rect 1680 1660 1793 1710
rect 1870 1851 2187 1857
rect 1870 1814 1997 1851
rect 1870 1660 1917 1814
rect 1985 1805 1997 1814
rect 2043 1814 2187 1851
rect 2043 1805 2055 1814
rect 1985 1793 2055 1805
rect 2140 1752 2187 1814
rect 2140 1740 2188 1752
rect 2140 1730 2187 1740
rect 2119 1660 2189 1730
rect 1680 1650 2189 1660
rect 1680 1648 2200 1650
rect 2270 1648 2316 1858
rect 2378 1892 2458 1905
rect 2378 1840 2392 1892
rect 2444 1840 2458 1892
rect 2378 1826 2458 1840
rect 2542 1747 2588 2080
rect 2655 1893 2735 1907
rect 2655 1841 2669 1893
rect 2721 1841 2735 1893
rect 2655 1827 2735 1841
rect 2526 1735 2608 1747
rect 2526 1683 2541 1735
rect 2593 1683 2608 1735
rect 2526 1670 2608 1683
rect 1527 1634 1575 1645
rect 1527 1560 1574 1634
rect 1680 1630 2316 1648
rect 1680 1584 1709 1630
rect 1755 1584 2316 1630
rect 1527 1549 1575 1560
rect 1680 1537 2316 1584
rect 1680 1520 2200 1537
rect 1680 1480 1793 1520
rect 1680 1434 1709 1480
rect 1755 1434 1793 1480
rect 1680 1357 1793 1434
rect 1257 1347 1793 1357
rect 1257 1310 1384 1347
rect 1100 1217 1196 1249
rect 1100 1165 1117 1217
rect 1169 1165 1196 1217
rect 1100 1143 1196 1165
rect 1257 1150 1304 1310
rect 1372 1301 1384 1310
rect 1430 1330 1793 1347
rect 1430 1311 1709 1330
rect 1430 1310 1574 1311
rect 1430 1301 1442 1310
rect 1372 1289 1442 1301
rect 1527 1248 1574 1310
rect 1680 1284 1709 1311
rect 1755 1328 1793 1330
rect 1870 1516 2200 1520
rect 1870 1479 1997 1516
rect 1870 1328 1917 1479
rect 1985 1470 1997 1479
rect 2043 1503 2200 1516
rect 2043 1479 2187 1503
rect 2043 1470 2055 1479
rect 1985 1458 2055 1470
rect 2140 1417 2187 1479
rect 2140 1405 2188 1417
rect 2270 1413 2316 1537
rect 2388 1582 2468 1595
rect 2388 1530 2402 1582
rect 2454 1530 2468 1582
rect 2388 1516 2468 1530
rect 2140 1362 2187 1405
rect 2241 1387 2345 1413
rect 2119 1328 2189 1362
rect 1755 1284 2189 1328
rect 2241 1335 2265 1387
rect 2317 1335 2345 1387
rect 2241 1307 2345 1335
rect 1680 1248 2189 1284
rect 2270 1248 2316 1307
rect 1527 1237 1575 1248
rect 1527 1163 1574 1237
rect 1680 1188 2316 1248
rect 1680 1180 1793 1188
rect 1527 1152 1575 1163
rect -554 995 -525 1041
rect -479 995 -441 1041
rect -554 924 -441 995
rect 160 1052 247 1070
rect 160 1000 178 1052
rect 230 1000 247 1052
rect 160 982 247 1000
rect 312 1029 903 1075
rect 1680 1134 1709 1180
rect 1755 1134 1793 1180
rect -554 911 -48 924
rect -554 891 -238 911
rect -554 845 -525 891
rect -479 875 -238 891
rect -479 845 -441 875
rect -554 741 -441 845
rect -554 695 -525 741
rect -479 695 -441 741
rect -365 874 -238 875
rect -365 714 -318 874
rect -250 865 -238 874
rect -192 874 -48 911
rect -192 865 -180 874
rect -250 853 -180 865
rect -95 716 -48 874
rect 24 793 105 813
rect 24 741 38 793
rect 90 741 105 793
rect 24 713 105 741
rect -554 591 -441 695
rect -554 545 -525 591
rect -479 548 -441 591
rect 149 632 236 650
rect 149 580 167 632
rect 219 580 236 632
rect 149 562 236 580
rect -479 545 -48 548
rect -554 535 -48 545
rect -554 499 -238 535
rect -554 441 -441 499
rect -554 395 -525 441
rect -479 395 -441 441
rect -554 291 -441 395
rect -365 498 -238 499
rect -365 338 -318 498
rect -250 489 -238 498
rect -192 498 -48 535
rect -192 489 -180 498
rect -250 477 -180 489
rect -95 340 -48 498
rect 26 417 104 437
rect 26 365 38 417
rect 90 365 104 417
rect 26 338 104 365
rect -554 245 -525 291
rect -479 245 -441 291
rect 312 284 359 1029
rect 428 959 515 977
rect 428 907 446 959
rect 498 907 515 959
rect 428 889 515 907
rect 708 960 795 978
rect 708 908 726 960
rect 778 908 795 960
rect 708 890 795 908
rect 582 793 654 814
rect 582 741 589 793
rect 641 741 654 793
rect 582 714 654 741
rect 416 576 503 594
rect 416 524 434 576
rect 486 524 503 576
rect 416 506 503 524
rect 694 587 781 605
rect 694 535 712 587
rect 764 535 781 587
rect 694 517 781 535
rect 580 417 655 438
rect 580 365 589 417
rect 641 365 655 417
rect 580 338 655 365
rect 856 284 903 1029
rect 967 1043 1054 1061
rect 967 991 985 1043
rect 1037 991 1054 1043
rect 967 973 1054 991
rect 1680 1030 1793 1134
rect 1680 984 1709 1030
rect 1755 989 1793 1030
rect 1870 1180 2316 1188
rect 1870 1143 1997 1180
rect 1870 989 1917 1143
rect 1985 1134 1997 1143
rect 2043 1143 2316 1180
rect 2391 1229 2471 1242
rect 2391 1177 2405 1229
rect 2457 1177 2471 1229
rect 2391 1163 2471 1177
rect 2043 1134 2055 1143
rect 2113 1137 2316 1143
rect 1985 1122 2055 1134
rect 2140 1081 2187 1137
rect 2140 1069 2188 1081
rect 2140 1011 2187 1069
rect 2130 989 2200 1011
rect 1755 984 2200 989
rect 1680 945 2200 984
rect 2270 945 2316 1137
rect 2542 1084 2588 1670
rect 2665 1583 2745 1597
rect 2665 1531 2679 1583
rect 2731 1531 2745 1583
rect 2665 1517 2745 1531
rect 2814 1425 2860 2160
rect 2919 1893 2999 1907
rect 2919 1841 2934 1893
rect 2986 1841 2999 1893
rect 2919 1827 2999 1841
rect 3086 1758 3132 2080
rect 3194 1894 3274 1908
rect 3194 1842 3208 1894
rect 3260 1842 3274 1894
rect 3194 1828 3274 1842
rect 3048 1733 3152 1758
rect 3048 1681 3072 1733
rect 3124 1681 3152 1733
rect 3048 1652 3152 1681
rect 2929 1583 3009 1597
rect 2929 1531 2944 1583
rect 2996 1531 3009 1583
rect 2929 1517 3009 1531
rect 2786 1392 2890 1425
rect 2786 1340 2815 1392
rect 2867 1340 2890 1392
rect 2786 1319 2890 1340
rect 2668 1230 2748 1244
rect 2668 1178 2682 1230
rect 2734 1178 2748 1230
rect 2668 1164 2748 1178
rect 2516 1055 2620 1084
rect 2516 1003 2540 1055
rect 2592 1003 2620 1055
rect 2516 978 2620 1003
rect 1680 922 2316 945
rect 1528 921 2316 922
rect 1257 911 2316 921
rect 1257 874 1384 911
rect 1122 793 1203 815
rect 1122 741 1138 793
rect 1190 741 1203 793
rect 1122 715 1203 741
rect 1257 714 1304 874
rect 1372 865 1384 874
rect 1430 880 2316 911
rect 1430 876 1709 880
rect 1430 874 1574 876
rect 1430 865 1442 874
rect 1372 853 1442 865
rect 1527 812 1574 874
rect 1680 834 1709 876
rect 1755 849 2316 880
rect 1755 834 1793 849
rect 1527 801 1575 812
rect 1527 727 1574 801
rect 1680 730 1793 834
rect 1527 716 1575 727
rect 1680 684 1709 730
rect 1755 684 1793 730
rect 977 636 1064 654
rect 977 584 995 636
rect 1047 584 1064 636
rect 977 566 1064 584
rect 1680 580 1793 684
rect 1870 844 2316 849
rect 1870 807 1997 844
rect 1870 647 1917 807
rect 1985 798 1997 807
rect 2043 834 2316 844
rect 2043 807 2187 834
rect 2043 798 2055 807
rect 1985 786 2055 798
rect 2140 745 2187 807
rect 2140 733 2188 745
rect 2270 744 2316 834
rect 2391 894 2471 907
rect 2391 842 2405 894
rect 2457 842 2471 894
rect 2391 828 2471 842
rect 2140 660 2187 733
rect 2245 714 2349 744
rect 2245 662 2270 714
rect 2322 662 2349 714
rect 2140 649 2188 660
rect 2142 648 2188 649
rect 2245 638 2349 662
rect 1680 546 1709 580
rect 1257 536 1709 546
rect 1257 499 1384 536
rect 1119 417 1193 438
rect 1119 365 1128 417
rect 1180 365 1193 417
rect 1119 337 1193 365
rect 1257 339 1304 499
rect 1372 490 1384 499
rect 1430 534 1709 536
rect 1755 534 1793 580
rect 1430 500 1793 534
rect 1430 499 1574 500
rect 1430 490 1442 499
rect 1372 478 1442 490
rect 1527 437 1574 499
rect 1527 426 1575 437
rect 1680 430 1793 500
rect 1527 352 1574 426
rect 1680 384 1709 430
rect 1755 384 1793 430
rect 1527 341 1575 352
rect 1680 347 1793 384
rect 2270 347 2316 638
rect 2542 570 2588 978
rect 2668 895 2748 909
rect 2668 843 2682 895
rect 2734 843 2748 895
rect 2668 829 2748 843
rect 2814 751 2860 1319
rect 2932 1230 3012 1244
rect 2932 1178 2947 1230
rect 2999 1178 3012 1230
rect 2932 1164 3012 1178
rect 3086 1083 3132 1652
rect 3204 1584 3284 1598
rect 3204 1532 3218 1584
rect 3270 1532 3284 1584
rect 3204 1518 3284 1532
rect 3358 1424 3404 2160
rect 3465 1893 3545 1907
rect 3465 1841 3480 1893
rect 3532 1841 3545 1893
rect 3465 1827 3545 1841
rect 3630 1761 3676 2080
rect 3736 1891 3816 1906
rect 3736 1839 3750 1891
rect 3802 1839 3816 1891
rect 3736 1826 3816 1839
rect 3597 1736 3701 1761
rect 3597 1684 3624 1736
rect 3676 1684 3701 1736
rect 3597 1655 3701 1684
rect 3475 1583 3555 1597
rect 3475 1531 3490 1583
rect 3542 1531 3555 1583
rect 3475 1517 3555 1531
rect 3333 1392 3437 1424
rect 3333 1340 3360 1392
rect 3412 1340 3437 1392
rect 3333 1318 3437 1340
rect 3207 1231 3287 1245
rect 3207 1179 3221 1231
rect 3273 1179 3287 1231
rect 3207 1165 3287 1179
rect 3057 1050 3161 1083
rect 3057 998 3080 1050
rect 3132 998 3161 1050
rect 3057 977 3161 998
rect 2932 895 3012 909
rect 2932 843 2947 895
rect 2999 843 3012 895
rect 2932 829 3012 843
rect 2790 723 2894 751
rect 2790 671 2815 723
rect 2867 671 2894 723
rect 2790 645 2894 671
rect 3086 570 3132 977
rect 3207 896 3287 910
rect 3207 844 3221 896
rect 3273 844 3287 896
rect 3207 830 3287 844
rect 3358 754 3404 1318
rect 3478 1230 3558 1244
rect 3478 1178 3493 1230
rect 3545 1178 3558 1230
rect 3478 1164 3558 1178
rect 3630 1095 3676 1655
rect 3746 1581 3826 1596
rect 3746 1529 3760 1581
rect 3812 1529 3826 1581
rect 3746 1516 3826 1529
rect 3902 1423 3948 2160
rect 4446 2132 4703 2160
rect 4749 2132 5078 2178
rect 4446 2086 5078 2132
rect 4010 1893 4090 1907
rect 4010 1841 4018 1893
rect 4070 1841 4090 1893
rect 4010 1827 4090 1841
rect 4174 1755 4220 2080
rect 4446 2072 4493 2086
rect 4305 1892 4385 1907
rect 4305 1840 4321 1892
rect 4373 1840 4385 1892
rect 4305 1827 4385 1840
rect 4446 1859 4492 2072
rect 4576 1981 4623 2086
rect 4846 2083 5078 2086
rect 4846 2080 5010 2083
rect 4846 1983 4893 2080
rect 4986 2037 5010 2080
rect 5056 2037 5078 2083
rect 4986 1933 5078 2037
rect 4986 1887 5010 1933
rect 5056 1887 5078 1933
rect 4986 1863 5078 1887
rect 4575 1859 5078 1863
rect 4446 1850 5078 1859
rect 4446 1804 4702 1850
rect 4748 1804 5078 1850
rect 4446 1783 5078 1804
rect 4446 1766 5010 1783
rect 4143 1734 4248 1755
rect 4143 1682 4167 1734
rect 4219 1682 4248 1734
rect 4143 1659 4248 1682
rect 4020 1583 4100 1597
rect 4020 1531 4028 1583
rect 4080 1531 4100 1583
rect 4020 1517 4100 1531
rect 3880 1392 3984 1423
rect 3880 1340 3909 1392
rect 3961 1340 3984 1392
rect 3880 1317 3984 1340
rect 3749 1228 3829 1243
rect 3749 1176 3763 1228
rect 3815 1176 3829 1228
rect 3749 1163 3829 1176
rect 3601 1065 3705 1095
rect 3601 1013 3625 1065
rect 3677 1013 3705 1065
rect 3601 989 3705 1013
rect 3478 895 3558 909
rect 3478 843 3493 895
rect 3545 843 3558 895
rect 3478 829 3558 843
rect 3342 728 3446 754
rect 3342 676 3369 728
rect 3421 676 3446 728
rect 3342 648 3446 676
rect 3630 570 3676 989
rect 3749 893 3829 908
rect 3749 841 3763 893
rect 3815 841 3829 893
rect 3749 828 3829 841
rect 3902 755 3948 1317
rect 4023 1230 4103 1244
rect 4023 1178 4031 1230
rect 4083 1178 4103 1230
rect 4023 1164 4103 1178
rect 4174 1093 4220 1659
rect 4315 1582 4395 1597
rect 4315 1530 4331 1582
rect 4383 1530 4395 1582
rect 4315 1517 4395 1530
rect 4446 1593 4492 1766
rect 4575 1653 4622 1766
rect 4845 1746 5010 1766
rect 4845 1655 4892 1746
rect 4986 1737 5010 1746
rect 5056 1737 5078 1783
rect 4986 1633 5078 1737
rect 4986 1593 5010 1633
rect 4446 1587 5010 1593
rect 5056 1587 5078 1633
rect 4446 1514 5078 1587
rect 4446 1500 4703 1514
rect 4446 1425 4492 1500
rect 4576 1477 4703 1500
rect 4425 1396 4529 1425
rect 4425 1344 4449 1396
rect 4501 1344 4529 1396
rect 4425 1319 4529 1344
rect 4446 1248 4492 1319
rect 4576 1317 4623 1477
rect 4691 1468 4703 1477
rect 4749 1500 5078 1514
rect 4749 1477 4893 1500
rect 4749 1468 4761 1477
rect 4691 1456 4761 1468
rect 4846 1319 4893 1477
rect 4986 1483 5078 1500
rect 4986 1437 5010 1483
rect 5056 1437 5078 1483
rect 4986 1333 5078 1437
rect 4986 1287 5010 1333
rect 5056 1287 5078 1333
rect 4986 1248 5078 1287
rect 4318 1229 4398 1244
rect 4318 1177 4334 1229
rect 4386 1177 4398 1229
rect 4318 1164 4398 1177
rect 4446 1183 5078 1248
rect 4446 1179 5010 1183
rect 4446 1155 4701 1179
rect 4153 1065 4257 1093
rect 4153 1013 4179 1065
rect 4231 1013 4257 1065
rect 4153 987 4257 1013
rect 4023 895 4103 909
rect 4023 843 4031 895
rect 4083 843 4103 895
rect 4023 829 4103 843
rect 3874 728 3978 755
rect 3874 676 3900 728
rect 3952 676 3978 728
rect 3874 649 3978 676
rect 3902 648 3948 649
rect 4174 570 4220 987
rect 4446 912 4492 1155
rect 4574 1142 4701 1155
rect 4574 982 4621 1142
rect 4689 1133 4701 1142
rect 4747 1155 5010 1179
rect 4747 1142 4891 1155
rect 4747 1133 4759 1142
rect 4689 1121 4759 1133
rect 4844 984 4891 1142
rect 4986 1137 5010 1155
rect 5056 1137 5078 1183
rect 4986 1033 5078 1137
rect 4986 987 5010 1033
rect 5056 987 5078 1033
rect 4986 912 5078 987
rect 4318 894 4398 909
rect 4318 842 4334 894
rect 4386 842 4398 894
rect 4318 829 4398 842
rect 4446 883 5078 912
rect 4446 843 5010 883
rect 4446 831 4702 843
rect 4444 819 4702 831
rect 4444 758 4492 819
rect 4575 806 4702 819
rect 4420 728 4524 758
rect 4420 676 4445 728
rect 4497 676 4524 728
rect 4420 652 4524 676
rect 2542 533 4220 570
rect 2542 495 3409 533
rect 3389 481 3409 495
rect 3461 495 4220 533
rect 4444 648 4492 652
rect 3461 481 3483 495
rect 3389 472 3483 481
rect 4444 347 4491 648
rect 4575 646 4622 806
rect 4690 797 4702 806
rect 4748 837 5010 843
rect 5056 837 5078 883
rect 4748 819 5078 837
rect 4748 806 4892 819
rect 4748 797 4760 806
rect 4690 785 4760 797
rect 4845 648 4892 806
rect 4986 733 5078 819
rect 4986 687 5010 733
rect 5056 687 5078 733
rect 4986 583 5078 687
rect 4986 537 5010 583
rect 5056 537 5078 583
rect 4986 433 5078 537
rect 4986 387 5010 433
rect 5056 387 5078 433
rect 4986 347 5078 387
rect -726 229 -647 245
rect -791 227 -647 229
rect -791 175 -713 227
rect -661 175 -647 227
rect -791 173 -647 175
rect -726 162 -647 173
rect -554 141 -441 245
rect 152 239 239 257
rect 152 187 170 239
rect 222 187 239 239
rect 312 238 903 284
rect 1680 326 5078 347
rect 1680 325 2278 326
rect 1680 279 1730 325
rect 1776 279 1840 325
rect 1886 279 1950 325
rect 1996 279 2059 325
rect 2105 279 2169 325
rect 2215 280 2278 325
rect 2324 280 2428 326
rect 2474 280 2578 326
rect 2624 280 2728 326
rect 2774 280 2878 326
rect 2924 280 3028 326
rect 3074 280 3178 326
rect 3224 280 3328 326
rect 3374 280 3478 326
rect 3524 280 3628 326
rect 3674 280 3778 326
rect 3824 280 3928 326
rect 3974 280 4078 326
rect 4124 280 4228 326
rect 4274 280 4378 326
rect 4424 280 4528 326
rect 4574 325 4948 326
rect 4574 323 4801 325
rect 4574 280 4660 323
rect 2215 279 4660 280
rect 1680 277 4660 279
rect 4706 279 4801 323
rect 4847 280 4948 325
rect 4994 280 5078 326
rect 4847 279 5078 280
rect 4706 277 5078 279
rect 969 239 1056 257
rect 152 171 239 187
rect 560 179 610 238
rect 969 187 987 239
rect 1039 187 1056 239
rect -554 95 -525 141
rect -479 95 -441 141
rect 544 163 627 179
rect 969 173 1056 187
rect 1680 255 5078 277
rect 1680 176 1796 255
rect 544 111 559 163
rect 611 111 627 163
rect 544 97 627 111
rect 1680 130 1710 176
rect 1756 130 1796 176
rect -554 51 -441 95
rect 1680 51 1796 130
rect -554 30 1796 51
rect -554 -16 -158 30
rect -112 -16 -8 30
rect 38 -16 142 30
rect 188 -16 292 30
rect 338 -16 442 30
rect 488 -16 592 30
rect 638 -16 742 30
rect 788 -16 892 30
rect 938 -16 1042 30
rect 1088 -16 1192 30
rect 1238 -16 1342 30
rect 1388 -16 1483 30
rect 1529 -16 1673 30
rect 1719 -16 1796 30
rect -554 -40 1796 -16
<< via1 >>
rect 308 2664 360 2716
rect 1274 2687 1326 2739
rect 4189 2673 4241 2725
rect 4324 2674 4376 2726
rect 4194 2547 4246 2599
rect 4321 2544 4373 2596
rect -693 2223 -641 2275
rect -86 2351 -34 2403
rect 572 2351 624 2403
rect 1278 2351 1330 2403
rect 173 2246 225 2250
rect 173 2200 176 2246
rect 176 2200 222 2246
rect 222 2200 225 2246
rect 173 2198 225 2200
rect 982 2241 1034 2245
rect 982 2195 985 2241
rect 985 2195 1031 2241
rect 1031 2195 1034 2241
rect 982 2193 1034 2195
rect 38 2009 90 2061
rect 175 1837 227 1841
rect 175 1791 178 1837
rect 178 1791 224 1837
rect 224 1791 227 1837
rect 175 1789 227 1791
rect 589 2009 641 2061
rect 436 1878 488 1882
rect 436 1832 439 1878
rect 439 1832 485 1878
rect 485 1832 488 1878
rect 436 1830 488 1832
rect 720 1876 772 1880
rect 720 1830 723 1876
rect 723 1830 769 1876
rect 769 1830 772 1876
rect 720 1828 772 1830
rect 1138 2009 1190 2061
rect 984 1832 1036 1836
rect 984 1786 987 1832
rect 987 1786 1033 1832
rect 1033 1786 1036 1832
rect 984 1784 1036 1786
rect 38 1573 90 1625
rect 37 1176 89 1228
rect 589 1573 641 1625
rect 444 1420 496 1424
rect 444 1374 447 1420
rect 447 1374 493 1420
rect 493 1374 496 1420
rect 444 1372 496 1374
rect 710 1425 762 1429
rect 710 1379 713 1425
rect 713 1379 759 1425
rect 759 1379 762 1425
rect 710 1377 762 1379
rect 589 1177 641 1229
rect 1138 1573 1190 1625
rect 2392 1889 2444 1892
rect 2392 1843 2396 1889
rect 2396 1843 2442 1889
rect 2442 1843 2444 1889
rect 2392 1840 2444 1843
rect 2669 1888 2721 1893
rect 2669 1842 2671 1888
rect 2671 1842 2717 1888
rect 2717 1842 2721 1888
rect 2669 1841 2721 1842
rect 2541 1683 2593 1735
rect 1117 1165 1169 1217
rect 2402 1579 2454 1582
rect 2402 1533 2406 1579
rect 2406 1533 2452 1579
rect 2452 1533 2454 1579
rect 2402 1530 2454 1533
rect 2265 1335 2317 1387
rect 178 1048 230 1052
rect 178 1002 181 1048
rect 181 1002 227 1048
rect 227 1002 230 1048
rect 178 1000 230 1002
rect 38 741 90 793
rect 167 628 219 632
rect 167 582 170 628
rect 170 582 216 628
rect 216 582 219 628
rect 167 580 219 582
rect 38 365 90 417
rect 446 955 498 959
rect 446 909 449 955
rect 449 909 495 955
rect 495 909 498 955
rect 446 907 498 909
rect 726 956 778 960
rect 726 910 729 956
rect 729 910 775 956
rect 775 910 778 956
rect 726 908 778 910
rect 589 741 641 793
rect 434 572 486 576
rect 434 526 437 572
rect 437 526 483 572
rect 483 526 486 572
rect 434 524 486 526
rect 712 583 764 587
rect 712 537 715 583
rect 715 537 761 583
rect 761 537 764 583
rect 712 535 764 537
rect 589 365 641 417
rect 985 1039 1037 1043
rect 985 993 988 1039
rect 988 993 1034 1039
rect 1034 993 1037 1039
rect 985 991 1037 993
rect 2405 1226 2457 1229
rect 2405 1180 2409 1226
rect 2409 1180 2455 1226
rect 2455 1180 2457 1226
rect 2405 1177 2457 1180
rect 2679 1578 2731 1583
rect 2679 1532 2681 1578
rect 2681 1532 2727 1578
rect 2727 1532 2731 1578
rect 2679 1531 2731 1532
rect 2934 1888 2986 1893
rect 2934 1842 2937 1888
rect 2937 1842 2983 1888
rect 2983 1842 2986 1888
rect 2934 1841 2986 1842
rect 3208 1888 3260 1894
rect 3208 1842 3210 1888
rect 3210 1842 3256 1888
rect 3256 1842 3260 1888
rect 3072 1681 3124 1733
rect 2944 1578 2996 1583
rect 2944 1532 2947 1578
rect 2947 1532 2993 1578
rect 2993 1532 2996 1578
rect 2944 1531 2996 1532
rect 2815 1340 2867 1392
rect 2682 1225 2734 1230
rect 2682 1179 2684 1225
rect 2684 1179 2730 1225
rect 2730 1179 2734 1225
rect 2682 1178 2734 1179
rect 2540 1003 2592 1055
rect 1138 741 1190 793
rect 995 632 1047 636
rect 995 586 998 632
rect 998 586 1044 632
rect 1044 586 1047 632
rect 995 584 1047 586
rect 2405 891 2457 894
rect 2405 845 2409 891
rect 2409 845 2455 891
rect 2455 845 2457 891
rect 2405 842 2457 845
rect 2270 662 2322 714
rect 1128 365 1180 417
rect 2682 890 2734 895
rect 2682 844 2684 890
rect 2684 844 2730 890
rect 2730 844 2734 890
rect 2682 843 2734 844
rect 2947 1225 2999 1230
rect 2947 1179 2950 1225
rect 2950 1179 2996 1225
rect 2996 1179 2999 1225
rect 2947 1178 2999 1179
rect 3218 1578 3270 1584
rect 3218 1532 3220 1578
rect 3220 1532 3266 1578
rect 3266 1532 3270 1578
rect 3480 1887 3532 1893
rect 3480 1841 3482 1887
rect 3482 1841 3528 1887
rect 3528 1841 3532 1887
rect 3750 1887 3802 1891
rect 3750 1841 3752 1887
rect 3752 1841 3798 1887
rect 3798 1841 3802 1887
rect 3750 1839 3802 1841
rect 3624 1684 3676 1736
rect 3490 1577 3542 1583
rect 3490 1531 3492 1577
rect 3492 1531 3538 1577
rect 3538 1531 3542 1577
rect 3360 1340 3412 1392
rect 3221 1225 3273 1231
rect 3221 1179 3223 1225
rect 3223 1179 3269 1225
rect 3269 1179 3273 1225
rect 3080 998 3132 1050
rect 2947 890 2999 895
rect 2947 844 2950 890
rect 2950 844 2996 890
rect 2996 844 2999 890
rect 2947 843 2999 844
rect 2815 671 2867 723
rect 3221 890 3273 896
rect 3221 844 3223 890
rect 3223 844 3269 890
rect 3269 844 3273 890
rect 3493 1224 3545 1230
rect 3493 1178 3495 1224
rect 3495 1178 3541 1224
rect 3541 1178 3545 1224
rect 3760 1577 3812 1581
rect 3760 1531 3762 1577
rect 3762 1531 3808 1577
rect 3808 1531 3812 1577
rect 3760 1529 3812 1531
rect 4018 1889 4070 1893
rect 4018 1843 4021 1889
rect 4021 1843 4067 1889
rect 4067 1843 4070 1889
rect 4018 1841 4070 1843
rect 4321 1888 4373 1892
rect 4321 1842 4324 1888
rect 4324 1842 4370 1888
rect 4370 1842 4373 1888
rect 4321 1840 4373 1842
rect 4167 1682 4219 1734
rect 4028 1579 4080 1583
rect 4028 1533 4031 1579
rect 4031 1533 4077 1579
rect 4077 1533 4080 1579
rect 4028 1531 4080 1533
rect 3909 1340 3961 1392
rect 3763 1224 3815 1228
rect 3763 1178 3765 1224
rect 3765 1178 3811 1224
rect 3811 1178 3815 1224
rect 3763 1176 3815 1178
rect 3625 1013 3677 1065
rect 3493 889 3545 895
rect 3493 843 3495 889
rect 3495 843 3541 889
rect 3541 843 3545 889
rect 3369 676 3421 728
rect 3763 889 3815 893
rect 3763 843 3765 889
rect 3765 843 3811 889
rect 3811 843 3815 889
rect 3763 841 3815 843
rect 4031 1226 4083 1230
rect 4031 1180 4034 1226
rect 4034 1180 4080 1226
rect 4080 1180 4083 1226
rect 4031 1178 4083 1180
rect 4331 1578 4383 1582
rect 4331 1532 4334 1578
rect 4334 1532 4380 1578
rect 4380 1532 4383 1578
rect 4331 1530 4383 1532
rect 4449 1344 4501 1396
rect 4334 1225 4386 1229
rect 4334 1179 4337 1225
rect 4337 1179 4383 1225
rect 4383 1179 4386 1225
rect 4334 1177 4386 1179
rect 4179 1013 4231 1065
rect 4031 891 4083 895
rect 4031 845 4034 891
rect 4034 845 4080 891
rect 4080 845 4083 891
rect 4031 843 4083 845
rect 3900 676 3952 728
rect 4334 890 4386 894
rect 4334 844 4337 890
rect 4337 844 4383 890
rect 4383 844 4386 890
rect 4334 842 4386 844
rect 4445 676 4497 728
rect 3409 481 3461 533
rect -713 175 -661 227
rect 170 235 222 239
rect 170 189 173 235
rect 173 189 219 235
rect 219 189 222 235
rect 170 187 222 189
rect 987 235 1039 239
rect 987 189 990 235
rect 990 189 1036 235
rect 1036 189 1039 235
rect 987 187 1039 189
rect 559 111 611 163
<< metal2 >>
rect 1251 2739 1345 2756
rect 289 2716 375 2731
rect 289 2664 308 2716
rect 360 2664 375 2716
rect 1251 2687 1274 2739
rect 1326 2687 1345 2739
rect 1251 2677 1345 2687
rect 4169 2726 4394 2755
rect 4169 2725 4324 2726
rect 289 2655 375 2664
rect -101 2403 -21 2415
rect -101 2351 -86 2403
rect -34 2351 -21 2403
rect -101 2344 -21 2351
rect -707 2277 -626 2292
rect -707 2221 -695 2277
rect -639 2221 -626 2277
rect -707 2206 -626 2221
rect -89 1628 -31 2344
rect 155 2252 242 2268
rect 155 2196 171 2252
rect 227 2196 242 2252
rect 155 2180 242 2196
rect 35 2083 104 2138
rect 26 2061 104 2083
rect 26 2009 38 2061
rect 90 2009 104 2061
rect 26 1995 104 2009
rect 305 1995 363 2655
rect 1271 2420 1329 2677
rect 4169 2673 4189 2725
rect 4241 2674 4324 2725
rect 4376 2674 4394 2726
rect 4241 2673 4394 2674
rect 4169 2599 4394 2673
rect 4169 2547 4194 2599
rect 4246 2596 4394 2599
rect 4246 2547 4321 2596
rect 4169 2544 4321 2547
rect 4373 2544 4394 2596
rect 4169 2536 4394 2544
rect 557 2403 654 2418
rect 557 2351 572 2403
rect 624 2351 654 2403
rect 557 2336 654 2351
rect 1265 2403 1336 2420
rect 1265 2351 1278 2403
rect 1330 2351 1336 2403
rect 26 1981 363 1995
rect 585 2083 642 2336
rect 1265 2334 1336 2351
rect 964 2247 1051 2263
rect 964 2191 980 2247
rect 1036 2191 1051 2247
rect 964 2175 1051 2191
rect 585 2061 655 2083
rect 585 2009 589 2061
rect 641 2009 655 2061
rect 1123 2061 1203 2084
rect 1123 2059 1138 2061
rect 585 1985 655 2009
rect 852 2009 1138 2059
rect 1190 2009 1203 2061
rect 852 2001 1203 2009
rect 35 1937 363 1981
rect 157 1843 244 1859
rect 157 1787 173 1843
rect 229 1787 244 1843
rect 157 1771 244 1787
rect 25 1628 101 1640
rect -89 1625 101 1628
rect -89 1573 38 1625
rect 90 1573 101 1625
rect -89 1570 101 1573
rect 24 1554 101 1570
rect 305 1618 363 1937
rect 419 1884 505 1900
rect 419 1828 434 1884
rect 490 1828 505 1884
rect 419 1812 505 1828
rect 702 1882 789 1898
rect 702 1826 718 1882
rect 774 1826 789 1882
rect 702 1810 789 1826
rect 569 1625 657 1646
rect 569 1618 589 1625
rect 305 1573 589 1618
rect 641 1618 657 1625
rect 852 1618 910 2001
rect 1123 1981 1203 2001
rect 966 1838 1053 1854
rect 966 1782 982 1838
rect 1038 1782 1053 1838
rect 966 1766 1053 1782
rect 641 1573 910 1618
rect 305 1560 910 1573
rect 1122 1629 1206 1641
rect 1271 1629 1329 2334
rect 2378 1894 2458 1905
rect 2655 1894 2735 1907
rect 2919 1894 2999 1907
rect 3194 1894 3274 1908
rect 4319 1907 4375 2536
rect 3465 1894 3545 1907
rect 3736 1894 3816 1906
rect 4010 1894 4090 1907
rect 4305 1894 4385 1907
rect 2378 1893 3208 1894
rect 2378 1892 2669 1893
rect 2378 1840 2392 1892
rect 2444 1841 2669 1892
rect 2721 1841 2934 1893
rect 2986 1842 3208 1893
rect 3260 1893 4385 1894
rect 3260 1842 3480 1893
rect 2986 1841 3480 1842
rect 3532 1891 4018 1893
rect 3532 1841 3750 1891
rect 2444 1840 3750 1841
rect 2378 1839 3750 1840
rect 3802 1841 4018 1891
rect 4070 1892 4385 1893
rect 4070 1841 4321 1892
rect 3802 1840 4321 1841
rect 4373 1840 4385 1892
rect 3802 1839 4385 1840
rect 2378 1838 4385 1839
rect 2378 1826 2458 1838
rect 2655 1827 2735 1838
rect 2919 1827 2999 1838
rect 3194 1828 3274 1838
rect 3465 1827 3545 1838
rect 3736 1826 3816 1838
rect 4010 1827 4090 1838
rect 4305 1827 4385 1838
rect 3048 1747 3152 1758
rect 3597 1747 3701 1761
rect 4155 1755 4232 1756
rect 4143 1747 4248 1755
rect 2526 1736 4248 1747
rect 2526 1735 3624 1736
rect 2526 1683 2541 1735
rect 2593 1733 3624 1735
rect 2593 1683 3072 1733
rect 2526 1681 3072 1683
rect 3124 1684 3624 1733
rect 3676 1734 4248 1736
rect 3676 1684 4167 1734
rect 3124 1682 4167 1684
rect 4219 1682 4248 1734
rect 3124 1681 4248 1682
rect 2526 1670 4248 1681
rect 3048 1652 3152 1670
rect 3597 1655 3701 1670
rect 4143 1659 4248 1670
rect 1122 1625 1329 1629
rect 1122 1573 1138 1625
rect 1190 1573 1329 1625
rect 1122 1571 1329 1573
rect 2388 1584 2468 1595
rect 2665 1584 2745 1597
rect 2929 1584 3009 1597
rect 3204 1584 3284 1598
rect 3475 1584 3555 1597
rect 3746 1584 3826 1596
rect 4020 1584 4100 1597
rect 4315 1584 4395 1597
rect 2388 1583 3218 1584
rect 2388 1582 2679 1583
rect 569 1546 657 1560
rect 1122 1552 1206 1571
rect 426 1426 513 1442
rect 426 1370 442 1426
rect 498 1370 513 1426
rect 426 1354 513 1370
rect 581 1250 638 1546
rect 2388 1530 2402 1582
rect 2454 1531 2679 1582
rect 2731 1531 2944 1583
rect 2996 1532 3218 1583
rect 3270 1583 4395 1584
rect 3270 1532 3490 1583
rect 2996 1531 3490 1532
rect 3542 1581 4028 1583
rect 3542 1531 3760 1581
rect 2454 1530 3760 1531
rect 2388 1529 3760 1530
rect 3812 1531 4028 1581
rect 4080 1582 4395 1583
rect 4080 1531 4331 1582
rect 3812 1530 4331 1531
rect 4383 1530 4395 1582
rect 3812 1529 4395 1530
rect 2388 1528 4395 1529
rect 2388 1516 2468 1528
rect 2665 1517 2745 1528
rect 2929 1517 3009 1528
rect 3204 1518 3284 1528
rect 3475 1517 3555 1528
rect 3746 1516 3826 1528
rect 4020 1517 4100 1528
rect 4315 1517 4395 1528
rect 695 1431 779 1447
rect 695 1375 708 1431
rect 764 1375 779 1431
rect 2327 1413 4529 1427
rect 695 1359 779 1375
rect 2241 1396 4529 1413
rect 2241 1392 4449 1396
rect 2241 1387 2815 1392
rect 2241 1335 2265 1387
rect 2317 1340 2815 1387
rect 2867 1340 3360 1392
rect 3412 1340 3909 1392
rect 3961 1344 4449 1392
rect 4501 1344 4529 1396
rect 3961 1340 4529 1344
rect 2317 1335 4529 1340
rect 2241 1307 4529 1335
rect 2327 1306 4529 1307
rect 31 1231 103 1250
rect -171 1228 103 1231
rect -171 1176 37 1228
rect 89 1176 103 1228
rect 569 1249 638 1250
rect 569 1229 655 1249
rect 569 1221 589 1229
rect -171 1173 103 1176
rect -171 423 -113 1173
rect 31 1157 103 1173
rect 307 1177 589 1221
rect 641 1221 655 1229
rect 1100 1222 1196 1249
rect 2391 1231 2471 1242
rect 2668 1231 2748 1244
rect 2932 1231 3012 1244
rect 3207 1231 3287 1245
rect 3478 1231 3558 1244
rect 3749 1231 3829 1243
rect 4023 1231 4103 1244
rect 4318 1231 4398 1244
rect 2391 1230 3221 1231
rect 2391 1229 2682 1230
rect 641 1177 910 1221
rect 307 1165 910 1177
rect 160 1054 247 1070
rect 160 998 176 1054
rect 232 998 247 1054
rect 160 982 247 998
rect 307 870 363 1165
rect 569 1150 655 1165
rect 569 1149 634 1150
rect 428 961 515 977
rect 428 905 444 961
rect 500 905 515 961
rect 428 889 515 905
rect 708 962 795 978
rect 708 906 724 962
rect 780 906 795 962
rect 708 890 795 906
rect 23 811 363 870
rect 24 793 105 811
rect 24 741 38 793
rect 90 741 105 793
rect 24 713 105 741
rect 582 793 654 814
rect 582 741 589 793
rect 641 741 654 793
rect 582 714 654 741
rect 854 788 910 1165
rect 1100 1217 1431 1222
rect 1100 1165 1117 1217
rect 1169 1165 1431 1217
rect 1100 1160 1431 1165
rect 2391 1177 2405 1229
rect 2457 1178 2682 1229
rect 2734 1178 2947 1230
rect 2999 1179 3221 1230
rect 3273 1230 4398 1231
rect 3273 1179 3493 1230
rect 2999 1178 3493 1179
rect 3545 1228 4031 1230
rect 3545 1178 3763 1228
rect 2457 1177 3763 1178
rect 2391 1176 3763 1177
rect 3815 1178 4031 1228
rect 4083 1229 4398 1230
rect 4083 1178 4334 1229
rect 3815 1177 4334 1178
rect 4386 1177 4398 1229
rect 3815 1176 4398 1177
rect 2391 1175 4398 1176
rect 2391 1163 2471 1175
rect 2668 1164 2748 1175
rect 2932 1164 3012 1175
rect 3207 1165 3287 1175
rect 3478 1164 3558 1175
rect 3749 1163 3829 1175
rect 4023 1164 4103 1175
rect 4318 1164 4398 1175
rect 1100 1143 1196 1160
rect 967 1045 1054 1061
rect 967 989 983 1045
rect 1039 989 1054 1045
rect 967 973 1054 989
rect 1122 793 1203 815
rect 1122 788 1138 793
rect 854 741 1138 788
rect 1190 741 1203 793
rect 854 732 1203 741
rect 303 658 654 714
rect 149 634 236 650
rect 149 578 165 634
rect 221 578 236 634
rect 149 562 236 578
rect 26 423 104 437
rect -171 419 104 423
rect 303 419 359 658
rect 416 578 503 594
rect 416 522 432 578
rect 488 522 503 578
rect 416 506 503 522
rect 694 589 781 605
rect 694 533 710 589
rect 766 533 781 589
rect 694 517 781 533
rect -171 417 359 419
rect -171 365 38 417
rect 90 365 359 417
rect 26 363 359 365
rect 580 417 655 438
rect 580 365 589 417
rect 641 407 655 417
rect 855 407 911 732
rect 1122 715 1203 732
rect 977 638 1064 654
rect 977 582 993 638
rect 1049 582 1064 638
rect 977 566 1064 582
rect 641 365 911 407
rect 26 338 104 363
rect 580 351 911 365
rect 1119 421 1193 438
rect 1369 421 1431 1160
rect 2516 1067 2620 1084
rect 3057 1067 3161 1083
rect 3601 1067 3705 1095
rect 4153 1067 4257 1093
rect 2516 1065 4257 1067
rect 2516 1055 3625 1065
rect 2516 1003 2540 1055
rect 2592 1050 3625 1055
rect 2592 1003 3080 1050
rect 2516 998 3080 1003
rect 3132 1013 3625 1050
rect 3677 1013 4179 1065
rect 4231 1013 4257 1065
rect 3132 998 4257 1013
rect 2516 990 4257 998
rect 2516 978 2620 990
rect 3057 977 3161 990
rect 3601 989 3705 990
rect 4153 987 4257 990
rect 2391 896 2471 907
rect 2668 896 2748 909
rect 2932 896 3012 909
rect 3207 896 3287 910
rect 3478 896 3558 909
rect 3749 896 3829 908
rect 4023 896 4103 909
rect 4318 896 4398 909
rect 2391 895 3221 896
rect 2391 894 2682 895
rect 2391 842 2405 894
rect 2457 843 2682 894
rect 2734 843 2947 895
rect 2999 844 3221 895
rect 3273 895 4398 896
rect 3273 844 3493 895
rect 2999 843 3493 844
rect 3545 893 4031 895
rect 3545 843 3763 893
rect 2457 842 3763 843
rect 2391 841 3763 842
rect 3815 843 4031 893
rect 4083 894 4398 895
rect 4083 843 4334 894
rect 3815 842 4334 843
rect 4386 842 4398 894
rect 3815 841 4398 842
rect 2391 840 4398 841
rect 2391 828 2471 840
rect 2668 829 2748 840
rect 2932 829 3012 840
rect 3207 830 3287 840
rect 3478 829 3558 840
rect 3749 828 3829 840
rect 4023 829 4103 840
rect 4318 829 4398 840
rect 2245 735 2349 744
rect 2790 735 2894 751
rect 3342 735 3446 754
rect 3874 735 3978 755
rect 4420 735 4524 758
rect 2245 728 4532 735
rect 2245 723 3369 728
rect 2245 714 2815 723
rect 2245 662 2270 714
rect 2322 671 2815 714
rect 2867 676 3369 723
rect 3421 676 3900 728
rect 3952 676 4445 728
rect 4497 676 4532 728
rect 2867 671 4532 676
rect 2322 662 4532 671
rect 2245 649 4532 662
rect 2245 638 2349 649
rect 2790 645 2894 649
rect 3342 648 3446 649
rect 3389 533 3483 550
rect 3389 481 3409 533
rect 3461 481 3483 533
rect 3389 472 3483 481
rect 1119 417 1431 421
rect 1119 365 1128 417
rect 1180 365 1431 417
rect 1119 359 1431 365
rect 580 338 655 351
rect 1119 337 1193 359
rect -726 229 -647 245
rect -726 173 -715 229
rect -659 173 -647 229
rect -726 162 -647 173
rect 152 241 239 257
rect 152 185 168 241
rect 224 185 239 241
rect 152 171 239 185
rect 969 241 1056 257
rect 969 185 985 241
rect 1041 185 1056 241
rect 544 163 627 179
rect 969 173 1056 185
rect 544 111 559 163
rect 611 111 627 163
rect 544 110 627 111
rect 3406 110 3464 472
rect 544 97 3464 110
rect 555 52 3464 97
<< via2 >>
rect -695 2275 -639 2277
rect -695 2223 -693 2275
rect -693 2223 -641 2275
rect -641 2223 -639 2275
rect -695 2221 -639 2223
rect 171 2250 227 2252
rect 171 2198 173 2250
rect 173 2198 225 2250
rect 225 2198 227 2250
rect 171 2196 227 2198
rect 980 2245 1036 2247
rect 980 2193 982 2245
rect 982 2193 1034 2245
rect 1034 2193 1036 2245
rect 980 2191 1036 2193
rect 173 1841 229 1843
rect 173 1789 175 1841
rect 175 1789 227 1841
rect 227 1789 229 1841
rect 173 1787 229 1789
rect 434 1882 490 1884
rect 434 1830 436 1882
rect 436 1830 488 1882
rect 488 1830 490 1882
rect 434 1828 490 1830
rect 718 1880 774 1882
rect 718 1828 720 1880
rect 720 1828 772 1880
rect 772 1828 774 1880
rect 718 1826 774 1828
rect 982 1836 1038 1838
rect 982 1784 984 1836
rect 984 1784 1036 1836
rect 1036 1784 1038 1836
rect 982 1782 1038 1784
rect 442 1424 498 1426
rect 442 1372 444 1424
rect 444 1372 496 1424
rect 496 1372 498 1424
rect 442 1370 498 1372
rect 708 1429 764 1431
rect 708 1377 710 1429
rect 710 1377 762 1429
rect 762 1377 764 1429
rect 708 1375 764 1377
rect 176 1052 232 1054
rect 176 1000 178 1052
rect 178 1000 230 1052
rect 230 1000 232 1052
rect 176 998 232 1000
rect 444 959 500 961
rect 444 907 446 959
rect 446 907 498 959
rect 498 907 500 959
rect 444 905 500 907
rect 724 960 780 962
rect 724 908 726 960
rect 726 908 778 960
rect 778 908 780 960
rect 724 906 780 908
rect 983 1043 1039 1045
rect 983 991 985 1043
rect 985 991 1037 1043
rect 1037 991 1039 1043
rect 983 989 1039 991
rect 165 632 221 634
rect 165 580 167 632
rect 167 580 219 632
rect 219 580 221 632
rect 165 578 221 580
rect 432 576 488 578
rect 432 524 434 576
rect 434 524 486 576
rect 486 524 488 576
rect 432 522 488 524
rect 710 587 766 589
rect 710 535 712 587
rect 712 535 764 587
rect 764 535 766 587
rect 710 533 766 535
rect 993 636 1049 638
rect 993 584 995 636
rect 995 584 1047 636
rect 1047 584 1049 636
rect 993 582 1049 584
rect -715 227 -659 229
rect -715 175 -713 227
rect -713 175 -661 227
rect -661 175 -659 227
rect -715 173 -659 175
rect 168 239 224 241
rect 168 187 170 239
rect 170 187 222 239
rect 222 187 224 239
rect 168 185 224 187
rect 985 239 1041 241
rect 985 187 987 239
rect 987 187 1039 239
rect 1039 187 1041 239
rect 985 185 1041 187
<< metal3 >>
rect -707 2277 -626 2292
rect -707 2221 -695 2277
rect -639 2252 1272 2277
rect -639 2221 171 2252
rect -707 2206 -626 2221
rect 155 2196 171 2221
rect 227 2247 1272 2252
rect 227 2221 980 2247
rect 227 2196 242 2221
rect 155 2180 242 2196
rect 964 2191 980 2221
rect 1036 2221 1272 2247
rect 1036 2191 1051 2221
rect 964 2175 1051 2191
rect 408 1884 524 1907
rect -87 1868 51 1869
rect 408 1868 434 1884
rect -87 1843 434 1868
rect -87 1813 173 1843
rect -87 1060 -31 1813
rect 35 1812 173 1813
rect 157 1787 173 1812
rect 229 1828 434 1843
rect 490 1868 524 1884
rect 692 1882 808 1905
rect 692 1868 718 1882
rect 490 1828 718 1868
rect 229 1826 718 1828
rect 774 1868 808 1882
rect 774 1838 1100 1868
rect 774 1826 982 1838
rect 229 1812 982 1826
rect 229 1787 244 1812
rect 702 1810 789 1812
rect 157 1771 244 1787
rect 966 1782 982 1812
rect 1038 1812 1100 1838
rect 1038 1782 1053 1812
rect 966 1766 1053 1782
rect 1216 1453 1272 2221
rect 388 1431 1272 1453
rect 388 1426 708 1431
rect 388 1370 442 1426
rect 498 1375 708 1426
rect 764 1375 1272 1431
rect 498 1370 1272 1375
rect 388 1351 1272 1370
rect 127 1060 273 1088
rect -87 1054 273 1060
rect -87 998 176 1054
rect 232 1021 273 1054
rect 946 1048 1092 1090
rect 946 1045 1093 1048
rect 946 1022 983 1045
rect 691 1021 983 1022
rect 232 998 983 1021
rect -87 989 983 998
rect 1039 992 1093 1045
rect 1039 989 1092 992
rect -87 966 1092 989
rect -87 965 950 966
rect -726 229 -647 245
rect -87 229 -31 965
rect 411 961 569 965
rect 411 905 444 961
rect 500 905 569 961
rect 411 882 569 905
rect 691 962 849 965
rect 691 906 724 962
rect 780 906 849 962
rect 691 883 849 906
rect 149 639 238 652
rect 977 639 1066 656
rect 1216 639 1272 1351
rect 116 638 1272 639
rect 116 634 993 638
rect 116 582 165 634
rect 149 578 165 582
rect 221 589 993 634
rect 221 583 710 589
rect 221 582 278 583
rect 221 578 238 582
rect 149 562 238 578
rect 403 578 528 583
rect 403 522 432 578
rect 488 522 528 578
rect 682 563 710 583
rect 403 506 528 522
rect 694 533 710 563
rect 766 583 993 589
rect 766 563 791 583
rect 977 582 993 583
rect 1049 583 1272 638
rect 1049 582 1066 583
rect 977 566 1066 582
rect 766 533 781 563
rect 694 517 781 533
rect 145 241 248 266
rect 145 229 168 241
rect -726 173 -715 229
rect -659 185 168 229
rect 224 229 248 241
rect 961 241 1063 264
rect 961 229 985 241
rect 224 185 985 229
rect 1041 229 1063 241
rect 1041 185 1100 229
rect -659 173 1100 185
rect -726 162 -647 173
rect 115 171 302 173
use nmos_3p3_AG6HDQ  nmos_3p3_AG6HDQ_0
timestamp 1713185578
transform 1 0 1016 0 1 388
box -196 -118 196 118
use nmos_3p3_AG6HDQ  nmos_3p3_AG6HDQ_1
timestamp 1713185578
transform 1 0 200 0 1 388
box -196 -118 196 118
use nmos_3p3_AG6HDQ  nmos_3p3_AG6HDQ_2
timestamp 1713185578
transform 1 0 1016 0 1 1596
box -196 -118 196 118
use nmos_3p3_AG6HDQ  nmos_3p3_AG6HDQ_3
timestamp 1713185578
transform 1 0 200 0 1 1596
box -196 -118 196 118
use nmos_3p3_AG6HDQ  nmos_3p3_AG6HDQ_4
timestamp 1713185578
transform 1 0 200 0 1 764
box -196 -118 196 118
use nmos_3p3_AG6HDQ  nmos_3p3_AG6HDQ_5
timestamp 1713185578
transform 1 0 1016 0 1 764
box -196 -118 196 118
use nmos_3p3_AG6HDQ  nmos_3p3_AG6HDQ_6
timestamp 1713185578
transform 1 0 200 0 1 1200
box -196 -118 196 118
use nmos_3p3_AG6HDQ  nmos_3p3_AG6HDQ_7
timestamp 1713185578
transform 1 0 1016 0 1 1200
box -196 -118 196 118
use nmos_3p3_AG6HDQ  nmos_3p3_AG6HDQ_8
timestamp 1713185578
transform 1 0 200 0 1 2032
box -196 -118 196 118
use nmos_3p3_AG6HDQ  nmos_3p3_AG6HDQ_9
timestamp 1713185578
transform 1 0 1016 0 1 2032
box -196 -118 196 118
use nmos_3p3_AG6HDQ  nmos_3p3_AG6HDQ_10
timestamp 1713185578
transform 1 0 1416 0 1 764
box -196 -118 196 118
use nmos_3p3_AG6HDQ  nmos_3p3_AG6HDQ_11
timestamp 1713185578
transform 1 0 1416 0 1 1200
box -196 -118 196 118
use nmos_3p3_AG6HDQ  nmos_3p3_AG6HDQ_12
timestamp 1713185578
transform 1 0 1416 0 1 1596
box -196 -118 196 118
use nmos_3p3_AG6HDQ  nmos_3p3_AG6HDQ_13
timestamp 1713185578
transform 1 0 1416 0 1 388
box -196 -118 196 118
use nmos_3p3_AG6HDQ  nmos_3p3_AG6HDQ_14
timestamp 1713185578
transform 1 0 4734 0 1 696
box -196 -118 196 118
use nmos_3p3_AG6HDQ  nmos_3p3_AG6HDQ_15
timestamp 1713185578
transform 1 0 2029 0 1 2032
box -196 -118 196 118
use nmos_3p3_AG6HDQ  nmos_3p3_AG6HDQ_16
timestamp 1713185578
transform 1 0 2029 0 1 696
box -196 -118 196 118
use nmos_3p3_AG6HDQ  nmos_3p3_AG6HDQ_17
timestamp 1713185578
transform 1 0 2029 0 1 1703
box -196 -118 196 118
use nmos_3p3_AG6HDQ  nmos_3p3_AG6HDQ_18
timestamp 1713185578
transform 1 0 2029 0 1 1368
box -196 -118 196 118
use nmos_3p3_AG6HDQ  nmos_3p3_AG6HDQ_19
timestamp 1713185578
transform 1 0 2029 0 1 1032
box -196 -118 196 118
use nmos_3p3_AG6HDQ  nmos_3p3_AG6HDQ_20
timestamp 1713185578
transform 1 0 4735 0 1 2032
box -196 -118 196 118
use nmos_3p3_AG6HDQ  nmos_3p3_AG6HDQ_21
timestamp 1713185578
transform 1 0 4734 0 1 1704
box -196 -118 196 118
use nmos_3p3_AG6HDQ  nmos_3p3_AG6HDQ_22
timestamp 1713185578
transform 1 0 4735 0 1 1368
box -196 -118 196 118
use nmos_3p3_AG6HDQ  nmos_3p3_AG6HDQ_23
timestamp 1713185578
transform 1 0 4733 0 1 1032
box -196 -118 196 118
use nmos_3p3_AG6HDQ  nmos_3p3_AG6HDQ_24
timestamp 1713185578
transform 1 0 -202 0 1 2031
box -196 -118 196 118
use nmos_3p3_AG6HDQ  nmos_3p3_AG6HDQ_25
timestamp 1713185578
transform 1 0 -206 0 1 388
box -196 -118 196 118
use nmos_3p3_AG6HDQ  nmos_3p3_AG6HDQ_26
timestamp 1713185578
transform 1 0 -202 0 1 1596
box -196 -118 196 118
use nmos_3p3_AG6HDQ  nmos_3p3_AG6HDQ_27
timestamp 1713185578
transform 1 0 -204 0 1 1200
box -196 -118 196 118
use nmos_3p3_AG6HDQ  nmos_3p3_AG6HDQ_28
timestamp 1713185578
transform 1 0 -206 0 1 764
box -196 -118 196 118
use nmos_3p3_AG6HDQ  nmos_3p3_AG6HDQ_29
timestamp 1713185578
transform 1 0 1417 0 1 2032
box -196 -118 196 118
use nmos_3p3_FG6HDQ  nmos_3p3_FG6HDQ_0
timestamp 1713185578
transform 1 0 3381 0 1 2032
box -1148 -118 1148 118
use nmos_3p3_FG6HDQ  nmos_3p3_FG6HDQ_1
timestamp 1713185578
transform 1 0 3381 0 1 1032
box -1148 -118 1148 118
use nmos_3p3_FG6HDQ  nmos_3p3_FG6HDQ_2
timestamp 1713185578
transform 1 0 3381 0 1 696
box -1148 -118 1148 118
use nmos_3p3_FG6HDQ  nmos_3p3_FG6HDQ_3
timestamp 1713185578
transform 1 0 3381 0 1 1368
box -1148 -118 1148 118
use nmos_3p3_FG6HDQ  nmos_3p3_FG6HDQ_4
timestamp 1713185578
transform 1 0 3381 0 1 1704
box -1148 -118 1148 118
use nmos_3p3_VB6HDQ  nmos_3p3_VB6HDQ_0
timestamp 1713185578
transform 1 0 608 0 1 388
box -332 -118 332 118
use nmos_3p3_VB6HDQ  nmos_3p3_VB6HDQ_1
timestamp 1713185578
transform 1 0 608 0 1 1596
box -332 -118 332 118
use nmos_3p3_VB6HDQ  nmos_3p3_VB6HDQ_2
timestamp 1713185578
transform 1 0 608 0 1 764
box -332 -118 332 118
use nmos_3p3_VB6HDQ  nmos_3p3_VB6HDQ_3
timestamp 1713185578
transform 1 0 608 0 1 1200
box -332 -118 332 118
use nmos_3p3_VB6HDQ  nmos_3p3_VB6HDQ_4
timestamp 1713185578
transform 1 0 608 0 1 2032
box -332 -118 332 118
<< labels >>
flabel metal1 s 1294 2771 1294 2771 0 FreeSans 750 0 0 0 M9
port 1 nsew
flabel metal1 s 328 2738 328 2738 0 FreeSans 750 0 0 0 M8
port 2 nsew
flabel metal1 s -738 2248 -738 2248 0 FreeSans 750 0 0 0 GM8
port 3 nsew
flabel metal1 s -758 200 -758 200 0 FreeSans 750 0 0 0 GM9
port 4 nsew
flabel metal1 s 3138 2279 3138 2279 0 FreeSans 750 0 0 0 VSS
port 5 nsew
flabel metal1 s 4260 2568 4260 2568 0 FreeSans 750 0 0 0 VCTRL2
port 6 nsew
<< end >>
