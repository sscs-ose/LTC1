magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -4495 -2195 4495 2195
<< psubdiff >>
rect -2495 173 2495 195
rect -2495 -173 -2473 173
rect 2473 -173 2495 173
rect -2495 -195 2495 -173
<< psubdiffcont >>
rect -2473 -173 2473 173
<< metal1 >>
rect -2484 173 2484 184
rect -2484 -173 -2473 173
rect 2473 -173 2484 173
rect -2484 -184 2484 -173
<< end >>
