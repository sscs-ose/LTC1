** sch_path: /home/shahid/GF180Projects/Top_test/top/xschem/pex_dec_3x8_updated_TB_ibr.sym
**.subckt pex_dec_3x8_updated_TB_ibr
V1 VDD VSS 3.3
.save i(v1)
V2 VSS GND 0
.save i(v2)
V3 IN1 VSS pulse(3.3 0 0 100p 100p 200n 400n)
.save i(v3)
V4 IN2 VSS pulse(3.3 0 0 100p 100p 100n 200n)
.save i(v4)
V5 IN3 VSS pulse(3.3 0 0 100p 100p 50n 100n)
.save i(v5)
x2 IN1 VSS VDD D0 D1 D2 D3 D4 D5 D6 D7 IN3 IN2 pex_dec_3x8_ibr_mag
**** begin user architecture code

.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical



.include pex_dec_3x8_ibr_mag.spice
.control
save all
tran 50p 500n
plot v(IN1) v(IN2)+3.5 v(IN3)+7 v(D0)+10.5 v(D1)+14 v(D2)+17.5 v(D3)+21 v(D4)+24.5 v(D5)+28
+ v(D6)+31.5 v(D7)+35



*write test_nfet_03v3.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
