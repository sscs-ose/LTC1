** sch_path: /home/shahid/Videos/opamp_xschem/Folded_Cascode_Amplifier/RES_TEST.sch
**.subckt RES_TEST VDD VOUT_N VOUT_P VIN_N VIN_P VOUT_OPAMP_N VOUT_OPAMP_P
*.iopin VDD
*.opin VOUT_N
*.opin VOUT_P
*.ipin VIN_N
*.ipin VIN_P
*.opin VOUT_OPAMP_N
*.opin VOUT_OPAMP_P
XR37 net7 VIN_P VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR1 net1 VIN_N VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR2 net8 net7 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR3 net2 net1 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR4 R7_R3_P net8 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR5 R7_R3_N net2 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR6 net9 R7_R3_P VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR7 net3 R7_R3_N VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR8 net10 net9 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR9 net4 net3 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR10 net12 net10 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR11 net48 net4 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR12 net11 net12 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR13 net5 net48 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR14 net13 net11 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR15 net6 net5 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR16 net14 net13 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR17 net15 net6 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR18 R7_R10_R8_P net14 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR19 R7_R10_R8_N net15 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR20 net20 R7_R10_R8_P VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR21 net16 R7_R10_R8_N VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR22 net21 net20 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR23 net17 net16 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR24 net23 net21 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR25 net47 net17 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR26 net22 net23 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR27 net18 net47 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR28 net24 net22 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR29 net19 net18 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR30 net25 net24 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR31 net26 net19 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR32 net27 net25 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR33 net28 net26 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR34 VOUT_OPAMP_P net27 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR35 VOUT_OPAMP_N net28 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR36 net29 R7_R10_R8_N VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR38 net30 net29 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR39 net46 net30 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR40 net31 net46 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR41 net32 net31 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR42 net33 net32 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR43 net34 net33 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR44 net45 net34 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR45 net35 net42 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR46 net36 net35 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR47 net38 net36 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR48 net37 net38 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR49 net39 net37 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR50 net40 net39 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR51 net41 net40 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR52 R7_R10_R8_P net41 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR53 net43 VOUT_N VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR54 net42 net43 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR55 net44 net45 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR56 VOUT_P net44 VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR57 VOUT_OPAMP_P VOUT_OPAMP_P VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR58 VOUT_OPAMP_N VOUT_OPAMP_N VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR59 VOUT_OPAMP_P VOUT_OPAMP_P VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR60 VOUT_OPAMP_N VOUT_OPAMP_N VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XC1 R7_R3_P R7_R3_N cap_mim_2f0_m4m5_noshield c_width=16.2e-6 c_length=15e-6 m=1
XC2 R7_R3_P R7_R3_N cap_mim_2f0_m4m5_noshield c_width=16.2e-6 c_length=15e-6 m=1
XC3 R7_R3_P R7_R3_N cap_mim_2f0_m4m5_noshield c_width=16.2e-6 c_length=15e-6 m=1
XC4 R7_R10_R8_N R7_R10_R8_P cap_mim_2f0_m4m5_noshield c_width=16.2e-6 c_length=15e-6 m=1
XC5 VOUT_N VOUT_OPAMP_P cap_mim_2f0_m4m5_noshield c_width=16e-6 c_length=15.2e-6 m=1
XC6 VOUT_P VOUT_OPAMP_N cap_mim_2f0_m4m5_noshield c_width=16e-6 c_length=15.2e-6 m=1
XR61 VDD VDD VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR62 VDD VDD VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR63 VDD VDD VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR64 VDD VDD VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR65 VDD VDD VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR66 VDD VDD VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR67 VDD VDD VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR68 VDD VDD VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR69 VDD VDD VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR70 VDD VDD VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR71 VDD VDD VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XR72 VDD VDD VDD ppolyf_u r_width=1e-6 r_length=2.3e-6 m=1
XC7 R7_R10_R8_N R7_R10_R8_P cap_mim_2f0_m4m5_noshield c_width=16.2e-6 c_length=15e-6 m=1
XC8 VOUT_P VOUT_OPAMP_N cap_mim_2f0_m4m5_noshield c_width=16e-6 c_length=15.2e-6 m=1
XC9 VOUT_N VOUT_OPAMP_P cap_mim_2f0_m4m5_noshield c_width=16e-6 c_length=15.2e-6 m=1
XC10 R7_R3_P R7_R3_N cap_mim_2f0_m4m5_noshield c_width=16.2e-6 c_length=15e-6 m=1
XC11 R7_R3_P R7_R3_N cap_mim_2f0_m4m5_noshield c_width=16.2e-6 c_length=15e-6 m=1
XC12 R7_R3_P R7_R3_N cap_mim_2f0_m4m5_noshield c_width=16.2e-6 c_length=15e-6 m=1
**.ends
.end
