* NGSPICE file created from resistor_PGA_new.ext - technology: gf180mcuC

.subckt ppolyf_u_W5AMT6 a_3240_n202# a_2280_n202# a_1320_n202# a_1320_100# a_n280_100#
+ a_n600_100# a_n1240_n202# a_n3160_n202# a_n4120_n202# a_1960_100# a_n1240_100# a_n2200_n202#
+ a_680_n202# a_n1880_100# a_2920_100# a_n2200_100# a_n2840_100# a_3560_100# a_40_n202#
+ a_n600_n202# a_n3480_100# a_n3800_100# a_3560_n202# a_2600_n202# a_1640_n202# a_n1560_n202#
+ a_n3480_n202# a_1000_100# a_680_100# a_n2520_n202# a_40_100# a_1640_100# a_n920_100#
+ a_1000_n202# a_n1560_100# a_2600_100# a_2280_100# w_n4304_n386# a_360_n202# a_n2520_100#
+ a_3240_100# a_3880_n202# a_n920_n202# a_3880_100# a_2920_n202# a_1960_n202# a_n3160_100#
+ a_n1880_n202# a_n2840_n202# a_n3800_n202# a_360_100# a_n280_n202# a_n4120_100#
X0 a_680_100# a_680_n202# w_n4304_n386# ppolyf_u r_width=1.2u r_length=1u
X1 a_3880_100# a_3880_n202# w_n4304_n386# ppolyf_u r_width=1.2u r_length=1u
X2 a_n2840_100# a_n2840_n202# w_n4304_n386# ppolyf_u r_width=1.2u r_length=1u
X3 a_2280_100# a_2280_n202# w_n4304_n386# ppolyf_u r_width=1.2u r_length=1u
X4 a_n1240_100# a_n1240_n202# w_n4304_n386# ppolyf_u r_width=1.2u r_length=1u
X5 a_1640_100# a_1640_n202# w_n4304_n386# ppolyf_u r_width=1.2u r_length=1u
X6 a_n280_100# a_n280_n202# w_n4304_n386# ppolyf_u r_width=1.2u r_length=1u
X7 a_n4120_100# a_n4120_n202# w_n4304_n386# ppolyf_u r_width=1.2u r_length=1u
X8 a_40_100# a_40_n202# w_n4304_n386# ppolyf_u r_width=1.2u r_length=1u
X9 a_n1880_100# a_n1880_n202# w_n4304_n386# ppolyf_u r_width=1.2u r_length=1u
X10 a_n3160_100# a_n3160_n202# w_n4304_n386# ppolyf_u r_width=1.2u r_length=1u
X11 a_360_100# a_360_n202# w_n4304_n386# ppolyf_u r_width=1.2u r_length=1u
X12 a_3560_100# a_3560_n202# w_n4304_n386# ppolyf_u r_width=1.2u r_length=1u
X13 a_n2520_100# a_n2520_n202# w_n4304_n386# ppolyf_u r_width=1.2u r_length=1u
X14 a_2920_100# a_2920_n202# w_n4304_n386# ppolyf_u r_width=1.2u r_length=1u
X15 a_1320_100# a_1320_n202# w_n4304_n386# ppolyf_u r_width=1.2u r_length=1u
X16 a_n3800_100# a_n3800_n202# w_n4304_n386# ppolyf_u r_width=1.2u r_length=1u
X17 a_n920_100# a_n920_n202# w_n4304_n386# ppolyf_u r_width=1.2u r_length=1u
X18 a_n2200_100# a_n2200_n202# w_n4304_n386# ppolyf_u r_width=1.2u r_length=1u
X19 a_n1560_100# a_n1560_n202# w_n4304_n386# ppolyf_u r_width=1.2u r_length=1u
X20 a_1960_100# a_1960_n202# w_n4304_n386# ppolyf_u r_width=1.2u r_length=1u
X21 a_n600_100# a_n600_n202# w_n4304_n386# ppolyf_u r_width=1.2u r_length=1u
X22 a_3240_100# a_3240_n202# w_n4304_n386# ppolyf_u r_width=1.2u r_length=1u
X23 a_2600_100# a_2600_n202# w_n4304_n386# ppolyf_u r_width=1.2u r_length=1u
X24 a_1000_100# a_1000_n202# w_n4304_n386# ppolyf_u r_width=1.2u r_length=1u
X25 a_n3480_100# a_n3480_n202# w_n4304_n386# ppolyf_u r_width=1.2u r_length=1u
.ends

.subckt resistor_PGA_new A B C D E F G H VDD
Xppolyf_u_W5AMT6_2 m1_12869_13281# m1_12454_14253# m1_12454_14253# m1_11494_14585#
+ m1_9748_14562# m1_9574_14585# m1_8069_13933# E VDD m1_12134_14585# m1_9254_14585#
+ m1_7109_13933# m1_10854_14253# m1_8294_14585# m1_13094_14585# m1_8294_14585# m1_7334_14585#
+ D m1_9989_14253# m1_9029_13281# G E m1_12869_13933# m1_11909_13933# m1_10949_13933#
+ m1_8614_14253# m1_6469_14253# m1_11174_14585# m1_11174_14585# m1_8614_14253# m1_9748_14562#
+ m1_12134_14585# m1_9254_14585# m1_10949_14253# m1_8934_14905# m1_13094_14585# m1_12774_14905#
+ VDD m1_10309_14253# m1_7654_14585# F VDD m1_9669_13933# VDD m1_13734_13933# m1_11909_14253#
+ m1_7334_14585# m1_8069_14253# m1_7109_14253# E m1_9574_14585# m1_9029_13933# VDD
+ ppolyf_u_W5AMT6
Xppolyf_u_W5AMT6_3 m1_13414_13601# m1_13414_13601# m1_11494_13601# m1_12454_13933#
+ m1_9669_13933# m1_9349_13933# m1_9254_13601# m1_7334_13601# VDD m1_11909_13933#
+ m1_8069_14253# m1_8294_13601# m1_11174_13601# m1_8069_13933# m1_12869_13933# m1_7109_14253#
+ m1_7109_13933# m1_13734_13933# m1_9770_13579# m1_9574_13601# A E F m1_13094_13601#
+ m1_12134_13601# m1_9574_13601# m1_7654_13601# m1_10949_13933# m1_9989_14253# m1_7654_13601#
+ m1_10854_14253# m1_10949_14253# m1_9029_13933# m1_11174_13601# m1_8614_13933# m1_11909_14253#
+ m1_12454_13933# VDD m1_11494_13601# m1_8614_13933# B VDD m1_9254_13601# VDD m1_13094_13601#
+ m1_12134_13601# E m1_8294_13601# m1_7334_13601# E m1_9989_14905# m1_9770_13579#
+ VDD ppolyf_u_W5AMT6
Xppolyf_u_W5AMT6_0 m1_13414_12949# m1_13414_12949# m1_11494_12949# m1_11269_13281#
+ m1_9400_13269# m1_9400_13269# m1_9254_12949# m1_7334_12949# VDD m1_11909_13281#
+ m1_8934_13281# m1_8294_12949# m1_11174_12949# m1_8069_13281# m1_12869_13281# m1_6469_14905#
+ m1_8934_13281# H m1_9731_12925# m1_9574_12949# G G H m1_13094_12949# m1_12134_12949#
+ m1_9574_12949# m1_7654_12949# m1_12774_13281# m1_10309_14253# m1_7654_12949# m1_10534_13281#
+ m1_10309_14905# m1_9029_13281# m1_11174_12949# m1_8389_13281# m1_12774_13281# m1_12229_13281#
+ VDD m1_11494_12949# m1_7429_13281# H VDD m1_9254_12949# VDD m1_13094_12949# m1_12134_12949#
+ m1_6469_14253# m1_8294_12949# m1_7334_12949# G m1_10534_13281# m1_9731_12925# VDD
+ ppolyf_u_W5AMT6
Xppolyf_u_W5AMT6_1 m1_11909_13281# m1_12454_14905# m1_11326_14886# m1_11269_13281#
+ m1_9749_15222# m1_9574_15237# m1_8934_14905# C VDD m1_12134_15237# m1_9254_15237#
+ m1_7486_14886# m1_9029_14905# m1_8294_15237# m1_13094_15237# m1_8294_15237# m1_7334_15237#
+ B m1_9989_14905# m1_8069_13281# C A B m1_12774_14905# m1_11326_14886# m1_8614_14905#
+ m1_6469_14905# m1_11174_15237# m1_11174_15237# m1_7486_14886# m1_9749_15222# m1_12134_15237#
+ m1_9254_15237# m1_11494_14585# m1_8389_13281# m1_13094_15237# m1_12229_13281# VDD
+ m1_10309_14905# m1_7429_13281# B VDD m1_9029_14905# VDD D m1_12454_14905# m1_7334_15237#
+ m1_8614_14905# m1_7654_14585# A m1_9574_15237# m1_9349_13933# VDD ppolyf_u_W5AMT6
.ends

