magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2478 -8178 2478 8178
<< nwell >>
rect -478 -6178 478 6178
<< nsubdiff >>
rect -395 6073 395 6095
rect -395 -6073 -373 6073
rect 373 -6073 395 6073
rect -395 -6095 395 -6073
<< nsubdiffcont >>
rect -373 -6073 373 6073
<< metal1 >>
rect -384 6073 384 6084
rect -384 -6073 -373 6073
rect 373 -6073 384 6073
rect -384 -6084 384 -6073
<< end >>
