magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -6662 -2786 6662 2786
<< psubdiff >>
rect -4662 764 4662 786
rect -4662 718 -4640 764
rect -4594 718 -4526 764
rect -4480 718 -4412 764
rect -4366 718 -4298 764
rect -4252 718 -4184 764
rect -4138 718 -4070 764
rect -4024 718 -3956 764
rect -3910 718 -3842 764
rect -3796 718 -3728 764
rect -3682 718 -3614 764
rect -3568 718 -3500 764
rect -3454 718 -3386 764
rect -3340 718 -3272 764
rect -3226 718 -3158 764
rect -3112 718 -3044 764
rect -2998 718 -2930 764
rect -2884 718 -2816 764
rect -2770 718 -2702 764
rect -2656 718 -2588 764
rect -2542 718 -2474 764
rect -2428 718 -2360 764
rect -2314 718 -2246 764
rect -2200 718 -2132 764
rect -2086 718 -2018 764
rect -1972 718 -1904 764
rect -1858 718 -1790 764
rect -1744 718 -1676 764
rect -1630 718 -1562 764
rect -1516 718 -1448 764
rect -1402 718 -1334 764
rect -1288 718 -1220 764
rect -1174 718 -1106 764
rect -1060 718 -992 764
rect -946 718 -878 764
rect -832 718 -764 764
rect -718 718 -650 764
rect -604 718 -536 764
rect -490 718 -422 764
rect -376 718 -308 764
rect -262 718 -194 764
rect -148 718 -80 764
rect -34 718 34 764
rect 80 718 148 764
rect 194 718 262 764
rect 308 718 376 764
rect 422 718 490 764
rect 536 718 604 764
rect 650 718 718 764
rect 764 718 832 764
rect 878 718 946 764
rect 992 718 1060 764
rect 1106 718 1174 764
rect 1220 718 1288 764
rect 1334 718 1402 764
rect 1448 718 1516 764
rect 1562 718 1630 764
rect 1676 718 1744 764
rect 1790 718 1858 764
rect 1904 718 1972 764
rect 2018 718 2086 764
rect 2132 718 2200 764
rect 2246 718 2314 764
rect 2360 718 2428 764
rect 2474 718 2542 764
rect 2588 718 2656 764
rect 2702 718 2770 764
rect 2816 718 2884 764
rect 2930 718 2998 764
rect 3044 718 3112 764
rect 3158 718 3226 764
rect 3272 718 3340 764
rect 3386 718 3454 764
rect 3500 718 3568 764
rect 3614 718 3682 764
rect 3728 718 3796 764
rect 3842 718 3910 764
rect 3956 718 4024 764
rect 4070 718 4138 764
rect 4184 718 4252 764
rect 4298 718 4366 764
rect 4412 718 4480 764
rect 4526 718 4594 764
rect 4640 718 4662 764
rect -4662 650 4662 718
rect -4662 604 -4640 650
rect -4594 604 -4526 650
rect -4480 604 -4412 650
rect -4366 604 -4298 650
rect -4252 604 -4184 650
rect -4138 604 -4070 650
rect -4024 604 -3956 650
rect -3910 604 -3842 650
rect -3796 604 -3728 650
rect -3682 604 -3614 650
rect -3568 604 -3500 650
rect -3454 604 -3386 650
rect -3340 604 -3272 650
rect -3226 604 -3158 650
rect -3112 604 -3044 650
rect -2998 604 -2930 650
rect -2884 604 -2816 650
rect -2770 604 -2702 650
rect -2656 604 -2588 650
rect -2542 604 -2474 650
rect -2428 604 -2360 650
rect -2314 604 -2246 650
rect -2200 604 -2132 650
rect -2086 604 -2018 650
rect -1972 604 -1904 650
rect -1858 604 -1790 650
rect -1744 604 -1676 650
rect -1630 604 -1562 650
rect -1516 604 -1448 650
rect -1402 604 -1334 650
rect -1288 604 -1220 650
rect -1174 604 -1106 650
rect -1060 604 -992 650
rect -946 604 -878 650
rect -832 604 -764 650
rect -718 604 -650 650
rect -604 604 -536 650
rect -490 604 -422 650
rect -376 604 -308 650
rect -262 604 -194 650
rect -148 604 -80 650
rect -34 604 34 650
rect 80 604 148 650
rect 194 604 262 650
rect 308 604 376 650
rect 422 604 490 650
rect 536 604 604 650
rect 650 604 718 650
rect 764 604 832 650
rect 878 604 946 650
rect 992 604 1060 650
rect 1106 604 1174 650
rect 1220 604 1288 650
rect 1334 604 1402 650
rect 1448 604 1516 650
rect 1562 604 1630 650
rect 1676 604 1744 650
rect 1790 604 1858 650
rect 1904 604 1972 650
rect 2018 604 2086 650
rect 2132 604 2200 650
rect 2246 604 2314 650
rect 2360 604 2428 650
rect 2474 604 2542 650
rect 2588 604 2656 650
rect 2702 604 2770 650
rect 2816 604 2884 650
rect 2930 604 2998 650
rect 3044 604 3112 650
rect 3158 604 3226 650
rect 3272 604 3340 650
rect 3386 604 3454 650
rect 3500 604 3568 650
rect 3614 604 3682 650
rect 3728 604 3796 650
rect 3842 604 3910 650
rect 3956 604 4024 650
rect 4070 604 4138 650
rect 4184 604 4252 650
rect 4298 604 4366 650
rect 4412 604 4480 650
rect 4526 604 4594 650
rect 4640 604 4662 650
rect -4662 536 4662 604
rect -4662 490 -4640 536
rect -4594 490 -4526 536
rect -4480 490 -4412 536
rect -4366 490 -4298 536
rect -4252 490 -4184 536
rect -4138 490 -4070 536
rect -4024 490 -3956 536
rect -3910 490 -3842 536
rect -3796 490 -3728 536
rect -3682 490 -3614 536
rect -3568 490 -3500 536
rect -3454 490 -3386 536
rect -3340 490 -3272 536
rect -3226 490 -3158 536
rect -3112 490 -3044 536
rect -2998 490 -2930 536
rect -2884 490 -2816 536
rect -2770 490 -2702 536
rect -2656 490 -2588 536
rect -2542 490 -2474 536
rect -2428 490 -2360 536
rect -2314 490 -2246 536
rect -2200 490 -2132 536
rect -2086 490 -2018 536
rect -1972 490 -1904 536
rect -1858 490 -1790 536
rect -1744 490 -1676 536
rect -1630 490 -1562 536
rect -1516 490 -1448 536
rect -1402 490 -1334 536
rect -1288 490 -1220 536
rect -1174 490 -1106 536
rect -1060 490 -992 536
rect -946 490 -878 536
rect -832 490 -764 536
rect -718 490 -650 536
rect -604 490 -536 536
rect -490 490 -422 536
rect -376 490 -308 536
rect -262 490 -194 536
rect -148 490 -80 536
rect -34 490 34 536
rect 80 490 148 536
rect 194 490 262 536
rect 308 490 376 536
rect 422 490 490 536
rect 536 490 604 536
rect 650 490 718 536
rect 764 490 832 536
rect 878 490 946 536
rect 992 490 1060 536
rect 1106 490 1174 536
rect 1220 490 1288 536
rect 1334 490 1402 536
rect 1448 490 1516 536
rect 1562 490 1630 536
rect 1676 490 1744 536
rect 1790 490 1858 536
rect 1904 490 1972 536
rect 2018 490 2086 536
rect 2132 490 2200 536
rect 2246 490 2314 536
rect 2360 490 2428 536
rect 2474 490 2542 536
rect 2588 490 2656 536
rect 2702 490 2770 536
rect 2816 490 2884 536
rect 2930 490 2998 536
rect 3044 490 3112 536
rect 3158 490 3226 536
rect 3272 490 3340 536
rect 3386 490 3454 536
rect 3500 490 3568 536
rect 3614 490 3682 536
rect 3728 490 3796 536
rect 3842 490 3910 536
rect 3956 490 4024 536
rect 4070 490 4138 536
rect 4184 490 4252 536
rect 4298 490 4366 536
rect 4412 490 4480 536
rect 4526 490 4594 536
rect 4640 490 4662 536
rect -4662 422 4662 490
rect -4662 376 -4640 422
rect -4594 376 -4526 422
rect -4480 376 -4412 422
rect -4366 376 -4298 422
rect -4252 376 -4184 422
rect -4138 376 -4070 422
rect -4024 376 -3956 422
rect -3910 376 -3842 422
rect -3796 376 -3728 422
rect -3682 376 -3614 422
rect -3568 376 -3500 422
rect -3454 376 -3386 422
rect -3340 376 -3272 422
rect -3226 376 -3158 422
rect -3112 376 -3044 422
rect -2998 376 -2930 422
rect -2884 376 -2816 422
rect -2770 376 -2702 422
rect -2656 376 -2588 422
rect -2542 376 -2474 422
rect -2428 376 -2360 422
rect -2314 376 -2246 422
rect -2200 376 -2132 422
rect -2086 376 -2018 422
rect -1972 376 -1904 422
rect -1858 376 -1790 422
rect -1744 376 -1676 422
rect -1630 376 -1562 422
rect -1516 376 -1448 422
rect -1402 376 -1334 422
rect -1288 376 -1220 422
rect -1174 376 -1106 422
rect -1060 376 -992 422
rect -946 376 -878 422
rect -832 376 -764 422
rect -718 376 -650 422
rect -604 376 -536 422
rect -490 376 -422 422
rect -376 376 -308 422
rect -262 376 -194 422
rect -148 376 -80 422
rect -34 376 34 422
rect 80 376 148 422
rect 194 376 262 422
rect 308 376 376 422
rect 422 376 490 422
rect 536 376 604 422
rect 650 376 718 422
rect 764 376 832 422
rect 878 376 946 422
rect 992 376 1060 422
rect 1106 376 1174 422
rect 1220 376 1288 422
rect 1334 376 1402 422
rect 1448 376 1516 422
rect 1562 376 1630 422
rect 1676 376 1744 422
rect 1790 376 1858 422
rect 1904 376 1972 422
rect 2018 376 2086 422
rect 2132 376 2200 422
rect 2246 376 2314 422
rect 2360 376 2428 422
rect 2474 376 2542 422
rect 2588 376 2656 422
rect 2702 376 2770 422
rect 2816 376 2884 422
rect 2930 376 2998 422
rect 3044 376 3112 422
rect 3158 376 3226 422
rect 3272 376 3340 422
rect 3386 376 3454 422
rect 3500 376 3568 422
rect 3614 376 3682 422
rect 3728 376 3796 422
rect 3842 376 3910 422
rect 3956 376 4024 422
rect 4070 376 4138 422
rect 4184 376 4252 422
rect 4298 376 4366 422
rect 4412 376 4480 422
rect 4526 376 4594 422
rect 4640 376 4662 422
rect -4662 308 4662 376
rect -4662 262 -4640 308
rect -4594 262 -4526 308
rect -4480 262 -4412 308
rect -4366 262 -4298 308
rect -4252 262 -4184 308
rect -4138 262 -4070 308
rect -4024 262 -3956 308
rect -3910 262 -3842 308
rect -3796 262 -3728 308
rect -3682 262 -3614 308
rect -3568 262 -3500 308
rect -3454 262 -3386 308
rect -3340 262 -3272 308
rect -3226 262 -3158 308
rect -3112 262 -3044 308
rect -2998 262 -2930 308
rect -2884 262 -2816 308
rect -2770 262 -2702 308
rect -2656 262 -2588 308
rect -2542 262 -2474 308
rect -2428 262 -2360 308
rect -2314 262 -2246 308
rect -2200 262 -2132 308
rect -2086 262 -2018 308
rect -1972 262 -1904 308
rect -1858 262 -1790 308
rect -1744 262 -1676 308
rect -1630 262 -1562 308
rect -1516 262 -1448 308
rect -1402 262 -1334 308
rect -1288 262 -1220 308
rect -1174 262 -1106 308
rect -1060 262 -992 308
rect -946 262 -878 308
rect -832 262 -764 308
rect -718 262 -650 308
rect -604 262 -536 308
rect -490 262 -422 308
rect -376 262 -308 308
rect -262 262 -194 308
rect -148 262 -80 308
rect -34 262 34 308
rect 80 262 148 308
rect 194 262 262 308
rect 308 262 376 308
rect 422 262 490 308
rect 536 262 604 308
rect 650 262 718 308
rect 764 262 832 308
rect 878 262 946 308
rect 992 262 1060 308
rect 1106 262 1174 308
rect 1220 262 1288 308
rect 1334 262 1402 308
rect 1448 262 1516 308
rect 1562 262 1630 308
rect 1676 262 1744 308
rect 1790 262 1858 308
rect 1904 262 1972 308
rect 2018 262 2086 308
rect 2132 262 2200 308
rect 2246 262 2314 308
rect 2360 262 2428 308
rect 2474 262 2542 308
rect 2588 262 2656 308
rect 2702 262 2770 308
rect 2816 262 2884 308
rect 2930 262 2998 308
rect 3044 262 3112 308
rect 3158 262 3226 308
rect 3272 262 3340 308
rect 3386 262 3454 308
rect 3500 262 3568 308
rect 3614 262 3682 308
rect 3728 262 3796 308
rect 3842 262 3910 308
rect 3956 262 4024 308
rect 4070 262 4138 308
rect 4184 262 4252 308
rect 4298 262 4366 308
rect 4412 262 4480 308
rect 4526 262 4594 308
rect 4640 262 4662 308
rect -4662 194 4662 262
rect -4662 148 -4640 194
rect -4594 148 -4526 194
rect -4480 148 -4412 194
rect -4366 148 -4298 194
rect -4252 148 -4184 194
rect -4138 148 -4070 194
rect -4024 148 -3956 194
rect -3910 148 -3842 194
rect -3796 148 -3728 194
rect -3682 148 -3614 194
rect -3568 148 -3500 194
rect -3454 148 -3386 194
rect -3340 148 -3272 194
rect -3226 148 -3158 194
rect -3112 148 -3044 194
rect -2998 148 -2930 194
rect -2884 148 -2816 194
rect -2770 148 -2702 194
rect -2656 148 -2588 194
rect -2542 148 -2474 194
rect -2428 148 -2360 194
rect -2314 148 -2246 194
rect -2200 148 -2132 194
rect -2086 148 -2018 194
rect -1972 148 -1904 194
rect -1858 148 -1790 194
rect -1744 148 -1676 194
rect -1630 148 -1562 194
rect -1516 148 -1448 194
rect -1402 148 -1334 194
rect -1288 148 -1220 194
rect -1174 148 -1106 194
rect -1060 148 -992 194
rect -946 148 -878 194
rect -832 148 -764 194
rect -718 148 -650 194
rect -604 148 -536 194
rect -490 148 -422 194
rect -376 148 -308 194
rect -262 148 -194 194
rect -148 148 -80 194
rect -34 148 34 194
rect 80 148 148 194
rect 194 148 262 194
rect 308 148 376 194
rect 422 148 490 194
rect 536 148 604 194
rect 650 148 718 194
rect 764 148 832 194
rect 878 148 946 194
rect 992 148 1060 194
rect 1106 148 1174 194
rect 1220 148 1288 194
rect 1334 148 1402 194
rect 1448 148 1516 194
rect 1562 148 1630 194
rect 1676 148 1744 194
rect 1790 148 1858 194
rect 1904 148 1972 194
rect 2018 148 2086 194
rect 2132 148 2200 194
rect 2246 148 2314 194
rect 2360 148 2428 194
rect 2474 148 2542 194
rect 2588 148 2656 194
rect 2702 148 2770 194
rect 2816 148 2884 194
rect 2930 148 2998 194
rect 3044 148 3112 194
rect 3158 148 3226 194
rect 3272 148 3340 194
rect 3386 148 3454 194
rect 3500 148 3568 194
rect 3614 148 3682 194
rect 3728 148 3796 194
rect 3842 148 3910 194
rect 3956 148 4024 194
rect 4070 148 4138 194
rect 4184 148 4252 194
rect 4298 148 4366 194
rect 4412 148 4480 194
rect 4526 148 4594 194
rect 4640 148 4662 194
rect -4662 80 4662 148
rect -4662 34 -4640 80
rect -4594 34 -4526 80
rect -4480 34 -4412 80
rect -4366 34 -4298 80
rect -4252 34 -4184 80
rect -4138 34 -4070 80
rect -4024 34 -3956 80
rect -3910 34 -3842 80
rect -3796 34 -3728 80
rect -3682 34 -3614 80
rect -3568 34 -3500 80
rect -3454 34 -3386 80
rect -3340 34 -3272 80
rect -3226 34 -3158 80
rect -3112 34 -3044 80
rect -2998 34 -2930 80
rect -2884 34 -2816 80
rect -2770 34 -2702 80
rect -2656 34 -2588 80
rect -2542 34 -2474 80
rect -2428 34 -2360 80
rect -2314 34 -2246 80
rect -2200 34 -2132 80
rect -2086 34 -2018 80
rect -1972 34 -1904 80
rect -1858 34 -1790 80
rect -1744 34 -1676 80
rect -1630 34 -1562 80
rect -1516 34 -1448 80
rect -1402 34 -1334 80
rect -1288 34 -1220 80
rect -1174 34 -1106 80
rect -1060 34 -992 80
rect -946 34 -878 80
rect -832 34 -764 80
rect -718 34 -650 80
rect -604 34 -536 80
rect -490 34 -422 80
rect -376 34 -308 80
rect -262 34 -194 80
rect -148 34 -80 80
rect -34 34 34 80
rect 80 34 148 80
rect 194 34 262 80
rect 308 34 376 80
rect 422 34 490 80
rect 536 34 604 80
rect 650 34 718 80
rect 764 34 832 80
rect 878 34 946 80
rect 992 34 1060 80
rect 1106 34 1174 80
rect 1220 34 1288 80
rect 1334 34 1402 80
rect 1448 34 1516 80
rect 1562 34 1630 80
rect 1676 34 1744 80
rect 1790 34 1858 80
rect 1904 34 1972 80
rect 2018 34 2086 80
rect 2132 34 2200 80
rect 2246 34 2314 80
rect 2360 34 2428 80
rect 2474 34 2542 80
rect 2588 34 2656 80
rect 2702 34 2770 80
rect 2816 34 2884 80
rect 2930 34 2998 80
rect 3044 34 3112 80
rect 3158 34 3226 80
rect 3272 34 3340 80
rect 3386 34 3454 80
rect 3500 34 3568 80
rect 3614 34 3682 80
rect 3728 34 3796 80
rect 3842 34 3910 80
rect 3956 34 4024 80
rect 4070 34 4138 80
rect 4184 34 4252 80
rect 4298 34 4366 80
rect 4412 34 4480 80
rect 4526 34 4594 80
rect 4640 34 4662 80
rect -4662 -34 4662 34
rect -4662 -80 -4640 -34
rect -4594 -80 -4526 -34
rect -4480 -80 -4412 -34
rect -4366 -80 -4298 -34
rect -4252 -80 -4184 -34
rect -4138 -80 -4070 -34
rect -4024 -80 -3956 -34
rect -3910 -80 -3842 -34
rect -3796 -80 -3728 -34
rect -3682 -80 -3614 -34
rect -3568 -80 -3500 -34
rect -3454 -80 -3386 -34
rect -3340 -80 -3272 -34
rect -3226 -80 -3158 -34
rect -3112 -80 -3044 -34
rect -2998 -80 -2930 -34
rect -2884 -80 -2816 -34
rect -2770 -80 -2702 -34
rect -2656 -80 -2588 -34
rect -2542 -80 -2474 -34
rect -2428 -80 -2360 -34
rect -2314 -80 -2246 -34
rect -2200 -80 -2132 -34
rect -2086 -80 -2018 -34
rect -1972 -80 -1904 -34
rect -1858 -80 -1790 -34
rect -1744 -80 -1676 -34
rect -1630 -80 -1562 -34
rect -1516 -80 -1448 -34
rect -1402 -80 -1334 -34
rect -1288 -80 -1220 -34
rect -1174 -80 -1106 -34
rect -1060 -80 -992 -34
rect -946 -80 -878 -34
rect -832 -80 -764 -34
rect -718 -80 -650 -34
rect -604 -80 -536 -34
rect -490 -80 -422 -34
rect -376 -80 -308 -34
rect -262 -80 -194 -34
rect -148 -80 -80 -34
rect -34 -80 34 -34
rect 80 -80 148 -34
rect 194 -80 262 -34
rect 308 -80 376 -34
rect 422 -80 490 -34
rect 536 -80 604 -34
rect 650 -80 718 -34
rect 764 -80 832 -34
rect 878 -80 946 -34
rect 992 -80 1060 -34
rect 1106 -80 1174 -34
rect 1220 -80 1288 -34
rect 1334 -80 1402 -34
rect 1448 -80 1516 -34
rect 1562 -80 1630 -34
rect 1676 -80 1744 -34
rect 1790 -80 1858 -34
rect 1904 -80 1972 -34
rect 2018 -80 2086 -34
rect 2132 -80 2200 -34
rect 2246 -80 2314 -34
rect 2360 -80 2428 -34
rect 2474 -80 2542 -34
rect 2588 -80 2656 -34
rect 2702 -80 2770 -34
rect 2816 -80 2884 -34
rect 2930 -80 2998 -34
rect 3044 -80 3112 -34
rect 3158 -80 3226 -34
rect 3272 -80 3340 -34
rect 3386 -80 3454 -34
rect 3500 -80 3568 -34
rect 3614 -80 3682 -34
rect 3728 -80 3796 -34
rect 3842 -80 3910 -34
rect 3956 -80 4024 -34
rect 4070 -80 4138 -34
rect 4184 -80 4252 -34
rect 4298 -80 4366 -34
rect 4412 -80 4480 -34
rect 4526 -80 4594 -34
rect 4640 -80 4662 -34
rect -4662 -148 4662 -80
rect -4662 -194 -4640 -148
rect -4594 -194 -4526 -148
rect -4480 -194 -4412 -148
rect -4366 -194 -4298 -148
rect -4252 -194 -4184 -148
rect -4138 -194 -4070 -148
rect -4024 -194 -3956 -148
rect -3910 -194 -3842 -148
rect -3796 -194 -3728 -148
rect -3682 -194 -3614 -148
rect -3568 -194 -3500 -148
rect -3454 -194 -3386 -148
rect -3340 -194 -3272 -148
rect -3226 -194 -3158 -148
rect -3112 -194 -3044 -148
rect -2998 -194 -2930 -148
rect -2884 -194 -2816 -148
rect -2770 -194 -2702 -148
rect -2656 -194 -2588 -148
rect -2542 -194 -2474 -148
rect -2428 -194 -2360 -148
rect -2314 -194 -2246 -148
rect -2200 -194 -2132 -148
rect -2086 -194 -2018 -148
rect -1972 -194 -1904 -148
rect -1858 -194 -1790 -148
rect -1744 -194 -1676 -148
rect -1630 -194 -1562 -148
rect -1516 -194 -1448 -148
rect -1402 -194 -1334 -148
rect -1288 -194 -1220 -148
rect -1174 -194 -1106 -148
rect -1060 -194 -992 -148
rect -946 -194 -878 -148
rect -832 -194 -764 -148
rect -718 -194 -650 -148
rect -604 -194 -536 -148
rect -490 -194 -422 -148
rect -376 -194 -308 -148
rect -262 -194 -194 -148
rect -148 -194 -80 -148
rect -34 -194 34 -148
rect 80 -194 148 -148
rect 194 -194 262 -148
rect 308 -194 376 -148
rect 422 -194 490 -148
rect 536 -194 604 -148
rect 650 -194 718 -148
rect 764 -194 832 -148
rect 878 -194 946 -148
rect 992 -194 1060 -148
rect 1106 -194 1174 -148
rect 1220 -194 1288 -148
rect 1334 -194 1402 -148
rect 1448 -194 1516 -148
rect 1562 -194 1630 -148
rect 1676 -194 1744 -148
rect 1790 -194 1858 -148
rect 1904 -194 1972 -148
rect 2018 -194 2086 -148
rect 2132 -194 2200 -148
rect 2246 -194 2314 -148
rect 2360 -194 2428 -148
rect 2474 -194 2542 -148
rect 2588 -194 2656 -148
rect 2702 -194 2770 -148
rect 2816 -194 2884 -148
rect 2930 -194 2998 -148
rect 3044 -194 3112 -148
rect 3158 -194 3226 -148
rect 3272 -194 3340 -148
rect 3386 -194 3454 -148
rect 3500 -194 3568 -148
rect 3614 -194 3682 -148
rect 3728 -194 3796 -148
rect 3842 -194 3910 -148
rect 3956 -194 4024 -148
rect 4070 -194 4138 -148
rect 4184 -194 4252 -148
rect 4298 -194 4366 -148
rect 4412 -194 4480 -148
rect 4526 -194 4594 -148
rect 4640 -194 4662 -148
rect -4662 -262 4662 -194
rect -4662 -308 -4640 -262
rect -4594 -308 -4526 -262
rect -4480 -308 -4412 -262
rect -4366 -308 -4298 -262
rect -4252 -308 -4184 -262
rect -4138 -308 -4070 -262
rect -4024 -308 -3956 -262
rect -3910 -308 -3842 -262
rect -3796 -308 -3728 -262
rect -3682 -308 -3614 -262
rect -3568 -308 -3500 -262
rect -3454 -308 -3386 -262
rect -3340 -308 -3272 -262
rect -3226 -308 -3158 -262
rect -3112 -308 -3044 -262
rect -2998 -308 -2930 -262
rect -2884 -308 -2816 -262
rect -2770 -308 -2702 -262
rect -2656 -308 -2588 -262
rect -2542 -308 -2474 -262
rect -2428 -308 -2360 -262
rect -2314 -308 -2246 -262
rect -2200 -308 -2132 -262
rect -2086 -308 -2018 -262
rect -1972 -308 -1904 -262
rect -1858 -308 -1790 -262
rect -1744 -308 -1676 -262
rect -1630 -308 -1562 -262
rect -1516 -308 -1448 -262
rect -1402 -308 -1334 -262
rect -1288 -308 -1220 -262
rect -1174 -308 -1106 -262
rect -1060 -308 -992 -262
rect -946 -308 -878 -262
rect -832 -308 -764 -262
rect -718 -308 -650 -262
rect -604 -308 -536 -262
rect -490 -308 -422 -262
rect -376 -308 -308 -262
rect -262 -308 -194 -262
rect -148 -308 -80 -262
rect -34 -308 34 -262
rect 80 -308 148 -262
rect 194 -308 262 -262
rect 308 -308 376 -262
rect 422 -308 490 -262
rect 536 -308 604 -262
rect 650 -308 718 -262
rect 764 -308 832 -262
rect 878 -308 946 -262
rect 992 -308 1060 -262
rect 1106 -308 1174 -262
rect 1220 -308 1288 -262
rect 1334 -308 1402 -262
rect 1448 -308 1516 -262
rect 1562 -308 1630 -262
rect 1676 -308 1744 -262
rect 1790 -308 1858 -262
rect 1904 -308 1972 -262
rect 2018 -308 2086 -262
rect 2132 -308 2200 -262
rect 2246 -308 2314 -262
rect 2360 -308 2428 -262
rect 2474 -308 2542 -262
rect 2588 -308 2656 -262
rect 2702 -308 2770 -262
rect 2816 -308 2884 -262
rect 2930 -308 2998 -262
rect 3044 -308 3112 -262
rect 3158 -308 3226 -262
rect 3272 -308 3340 -262
rect 3386 -308 3454 -262
rect 3500 -308 3568 -262
rect 3614 -308 3682 -262
rect 3728 -308 3796 -262
rect 3842 -308 3910 -262
rect 3956 -308 4024 -262
rect 4070 -308 4138 -262
rect 4184 -308 4252 -262
rect 4298 -308 4366 -262
rect 4412 -308 4480 -262
rect 4526 -308 4594 -262
rect 4640 -308 4662 -262
rect -4662 -376 4662 -308
rect -4662 -422 -4640 -376
rect -4594 -422 -4526 -376
rect -4480 -422 -4412 -376
rect -4366 -422 -4298 -376
rect -4252 -422 -4184 -376
rect -4138 -422 -4070 -376
rect -4024 -422 -3956 -376
rect -3910 -422 -3842 -376
rect -3796 -422 -3728 -376
rect -3682 -422 -3614 -376
rect -3568 -422 -3500 -376
rect -3454 -422 -3386 -376
rect -3340 -422 -3272 -376
rect -3226 -422 -3158 -376
rect -3112 -422 -3044 -376
rect -2998 -422 -2930 -376
rect -2884 -422 -2816 -376
rect -2770 -422 -2702 -376
rect -2656 -422 -2588 -376
rect -2542 -422 -2474 -376
rect -2428 -422 -2360 -376
rect -2314 -422 -2246 -376
rect -2200 -422 -2132 -376
rect -2086 -422 -2018 -376
rect -1972 -422 -1904 -376
rect -1858 -422 -1790 -376
rect -1744 -422 -1676 -376
rect -1630 -422 -1562 -376
rect -1516 -422 -1448 -376
rect -1402 -422 -1334 -376
rect -1288 -422 -1220 -376
rect -1174 -422 -1106 -376
rect -1060 -422 -992 -376
rect -946 -422 -878 -376
rect -832 -422 -764 -376
rect -718 -422 -650 -376
rect -604 -422 -536 -376
rect -490 -422 -422 -376
rect -376 -422 -308 -376
rect -262 -422 -194 -376
rect -148 -422 -80 -376
rect -34 -422 34 -376
rect 80 -422 148 -376
rect 194 -422 262 -376
rect 308 -422 376 -376
rect 422 -422 490 -376
rect 536 -422 604 -376
rect 650 -422 718 -376
rect 764 -422 832 -376
rect 878 -422 946 -376
rect 992 -422 1060 -376
rect 1106 -422 1174 -376
rect 1220 -422 1288 -376
rect 1334 -422 1402 -376
rect 1448 -422 1516 -376
rect 1562 -422 1630 -376
rect 1676 -422 1744 -376
rect 1790 -422 1858 -376
rect 1904 -422 1972 -376
rect 2018 -422 2086 -376
rect 2132 -422 2200 -376
rect 2246 -422 2314 -376
rect 2360 -422 2428 -376
rect 2474 -422 2542 -376
rect 2588 -422 2656 -376
rect 2702 -422 2770 -376
rect 2816 -422 2884 -376
rect 2930 -422 2998 -376
rect 3044 -422 3112 -376
rect 3158 -422 3226 -376
rect 3272 -422 3340 -376
rect 3386 -422 3454 -376
rect 3500 -422 3568 -376
rect 3614 -422 3682 -376
rect 3728 -422 3796 -376
rect 3842 -422 3910 -376
rect 3956 -422 4024 -376
rect 4070 -422 4138 -376
rect 4184 -422 4252 -376
rect 4298 -422 4366 -376
rect 4412 -422 4480 -376
rect 4526 -422 4594 -376
rect 4640 -422 4662 -376
rect -4662 -490 4662 -422
rect -4662 -536 -4640 -490
rect -4594 -536 -4526 -490
rect -4480 -536 -4412 -490
rect -4366 -536 -4298 -490
rect -4252 -536 -4184 -490
rect -4138 -536 -4070 -490
rect -4024 -536 -3956 -490
rect -3910 -536 -3842 -490
rect -3796 -536 -3728 -490
rect -3682 -536 -3614 -490
rect -3568 -536 -3500 -490
rect -3454 -536 -3386 -490
rect -3340 -536 -3272 -490
rect -3226 -536 -3158 -490
rect -3112 -536 -3044 -490
rect -2998 -536 -2930 -490
rect -2884 -536 -2816 -490
rect -2770 -536 -2702 -490
rect -2656 -536 -2588 -490
rect -2542 -536 -2474 -490
rect -2428 -536 -2360 -490
rect -2314 -536 -2246 -490
rect -2200 -536 -2132 -490
rect -2086 -536 -2018 -490
rect -1972 -536 -1904 -490
rect -1858 -536 -1790 -490
rect -1744 -536 -1676 -490
rect -1630 -536 -1562 -490
rect -1516 -536 -1448 -490
rect -1402 -536 -1334 -490
rect -1288 -536 -1220 -490
rect -1174 -536 -1106 -490
rect -1060 -536 -992 -490
rect -946 -536 -878 -490
rect -832 -536 -764 -490
rect -718 -536 -650 -490
rect -604 -536 -536 -490
rect -490 -536 -422 -490
rect -376 -536 -308 -490
rect -262 -536 -194 -490
rect -148 -536 -80 -490
rect -34 -536 34 -490
rect 80 -536 148 -490
rect 194 -536 262 -490
rect 308 -536 376 -490
rect 422 -536 490 -490
rect 536 -536 604 -490
rect 650 -536 718 -490
rect 764 -536 832 -490
rect 878 -536 946 -490
rect 992 -536 1060 -490
rect 1106 -536 1174 -490
rect 1220 -536 1288 -490
rect 1334 -536 1402 -490
rect 1448 -536 1516 -490
rect 1562 -536 1630 -490
rect 1676 -536 1744 -490
rect 1790 -536 1858 -490
rect 1904 -536 1972 -490
rect 2018 -536 2086 -490
rect 2132 -536 2200 -490
rect 2246 -536 2314 -490
rect 2360 -536 2428 -490
rect 2474 -536 2542 -490
rect 2588 -536 2656 -490
rect 2702 -536 2770 -490
rect 2816 -536 2884 -490
rect 2930 -536 2998 -490
rect 3044 -536 3112 -490
rect 3158 -536 3226 -490
rect 3272 -536 3340 -490
rect 3386 -536 3454 -490
rect 3500 -536 3568 -490
rect 3614 -536 3682 -490
rect 3728 -536 3796 -490
rect 3842 -536 3910 -490
rect 3956 -536 4024 -490
rect 4070 -536 4138 -490
rect 4184 -536 4252 -490
rect 4298 -536 4366 -490
rect 4412 -536 4480 -490
rect 4526 -536 4594 -490
rect 4640 -536 4662 -490
rect -4662 -604 4662 -536
rect -4662 -650 -4640 -604
rect -4594 -650 -4526 -604
rect -4480 -650 -4412 -604
rect -4366 -650 -4298 -604
rect -4252 -650 -4184 -604
rect -4138 -650 -4070 -604
rect -4024 -650 -3956 -604
rect -3910 -650 -3842 -604
rect -3796 -650 -3728 -604
rect -3682 -650 -3614 -604
rect -3568 -650 -3500 -604
rect -3454 -650 -3386 -604
rect -3340 -650 -3272 -604
rect -3226 -650 -3158 -604
rect -3112 -650 -3044 -604
rect -2998 -650 -2930 -604
rect -2884 -650 -2816 -604
rect -2770 -650 -2702 -604
rect -2656 -650 -2588 -604
rect -2542 -650 -2474 -604
rect -2428 -650 -2360 -604
rect -2314 -650 -2246 -604
rect -2200 -650 -2132 -604
rect -2086 -650 -2018 -604
rect -1972 -650 -1904 -604
rect -1858 -650 -1790 -604
rect -1744 -650 -1676 -604
rect -1630 -650 -1562 -604
rect -1516 -650 -1448 -604
rect -1402 -650 -1334 -604
rect -1288 -650 -1220 -604
rect -1174 -650 -1106 -604
rect -1060 -650 -992 -604
rect -946 -650 -878 -604
rect -832 -650 -764 -604
rect -718 -650 -650 -604
rect -604 -650 -536 -604
rect -490 -650 -422 -604
rect -376 -650 -308 -604
rect -262 -650 -194 -604
rect -148 -650 -80 -604
rect -34 -650 34 -604
rect 80 -650 148 -604
rect 194 -650 262 -604
rect 308 -650 376 -604
rect 422 -650 490 -604
rect 536 -650 604 -604
rect 650 -650 718 -604
rect 764 -650 832 -604
rect 878 -650 946 -604
rect 992 -650 1060 -604
rect 1106 -650 1174 -604
rect 1220 -650 1288 -604
rect 1334 -650 1402 -604
rect 1448 -650 1516 -604
rect 1562 -650 1630 -604
rect 1676 -650 1744 -604
rect 1790 -650 1858 -604
rect 1904 -650 1972 -604
rect 2018 -650 2086 -604
rect 2132 -650 2200 -604
rect 2246 -650 2314 -604
rect 2360 -650 2428 -604
rect 2474 -650 2542 -604
rect 2588 -650 2656 -604
rect 2702 -650 2770 -604
rect 2816 -650 2884 -604
rect 2930 -650 2998 -604
rect 3044 -650 3112 -604
rect 3158 -650 3226 -604
rect 3272 -650 3340 -604
rect 3386 -650 3454 -604
rect 3500 -650 3568 -604
rect 3614 -650 3682 -604
rect 3728 -650 3796 -604
rect 3842 -650 3910 -604
rect 3956 -650 4024 -604
rect 4070 -650 4138 -604
rect 4184 -650 4252 -604
rect 4298 -650 4366 -604
rect 4412 -650 4480 -604
rect 4526 -650 4594 -604
rect 4640 -650 4662 -604
rect -4662 -718 4662 -650
rect -4662 -764 -4640 -718
rect -4594 -764 -4526 -718
rect -4480 -764 -4412 -718
rect -4366 -764 -4298 -718
rect -4252 -764 -4184 -718
rect -4138 -764 -4070 -718
rect -4024 -764 -3956 -718
rect -3910 -764 -3842 -718
rect -3796 -764 -3728 -718
rect -3682 -764 -3614 -718
rect -3568 -764 -3500 -718
rect -3454 -764 -3386 -718
rect -3340 -764 -3272 -718
rect -3226 -764 -3158 -718
rect -3112 -764 -3044 -718
rect -2998 -764 -2930 -718
rect -2884 -764 -2816 -718
rect -2770 -764 -2702 -718
rect -2656 -764 -2588 -718
rect -2542 -764 -2474 -718
rect -2428 -764 -2360 -718
rect -2314 -764 -2246 -718
rect -2200 -764 -2132 -718
rect -2086 -764 -2018 -718
rect -1972 -764 -1904 -718
rect -1858 -764 -1790 -718
rect -1744 -764 -1676 -718
rect -1630 -764 -1562 -718
rect -1516 -764 -1448 -718
rect -1402 -764 -1334 -718
rect -1288 -764 -1220 -718
rect -1174 -764 -1106 -718
rect -1060 -764 -992 -718
rect -946 -764 -878 -718
rect -832 -764 -764 -718
rect -718 -764 -650 -718
rect -604 -764 -536 -718
rect -490 -764 -422 -718
rect -376 -764 -308 -718
rect -262 -764 -194 -718
rect -148 -764 -80 -718
rect -34 -764 34 -718
rect 80 -764 148 -718
rect 194 -764 262 -718
rect 308 -764 376 -718
rect 422 -764 490 -718
rect 536 -764 604 -718
rect 650 -764 718 -718
rect 764 -764 832 -718
rect 878 -764 946 -718
rect 992 -764 1060 -718
rect 1106 -764 1174 -718
rect 1220 -764 1288 -718
rect 1334 -764 1402 -718
rect 1448 -764 1516 -718
rect 1562 -764 1630 -718
rect 1676 -764 1744 -718
rect 1790 -764 1858 -718
rect 1904 -764 1972 -718
rect 2018 -764 2086 -718
rect 2132 -764 2200 -718
rect 2246 -764 2314 -718
rect 2360 -764 2428 -718
rect 2474 -764 2542 -718
rect 2588 -764 2656 -718
rect 2702 -764 2770 -718
rect 2816 -764 2884 -718
rect 2930 -764 2998 -718
rect 3044 -764 3112 -718
rect 3158 -764 3226 -718
rect 3272 -764 3340 -718
rect 3386 -764 3454 -718
rect 3500 -764 3568 -718
rect 3614 -764 3682 -718
rect 3728 -764 3796 -718
rect 3842 -764 3910 -718
rect 3956 -764 4024 -718
rect 4070 -764 4138 -718
rect 4184 -764 4252 -718
rect 4298 -764 4366 -718
rect 4412 -764 4480 -718
rect 4526 -764 4594 -718
rect 4640 -764 4662 -718
rect -4662 -786 4662 -764
<< psubdiffcont >>
rect -4640 718 -4594 764
rect -4526 718 -4480 764
rect -4412 718 -4366 764
rect -4298 718 -4252 764
rect -4184 718 -4138 764
rect -4070 718 -4024 764
rect -3956 718 -3910 764
rect -3842 718 -3796 764
rect -3728 718 -3682 764
rect -3614 718 -3568 764
rect -3500 718 -3454 764
rect -3386 718 -3340 764
rect -3272 718 -3226 764
rect -3158 718 -3112 764
rect -3044 718 -2998 764
rect -2930 718 -2884 764
rect -2816 718 -2770 764
rect -2702 718 -2656 764
rect -2588 718 -2542 764
rect -2474 718 -2428 764
rect -2360 718 -2314 764
rect -2246 718 -2200 764
rect -2132 718 -2086 764
rect -2018 718 -1972 764
rect -1904 718 -1858 764
rect -1790 718 -1744 764
rect -1676 718 -1630 764
rect -1562 718 -1516 764
rect -1448 718 -1402 764
rect -1334 718 -1288 764
rect -1220 718 -1174 764
rect -1106 718 -1060 764
rect -992 718 -946 764
rect -878 718 -832 764
rect -764 718 -718 764
rect -650 718 -604 764
rect -536 718 -490 764
rect -422 718 -376 764
rect -308 718 -262 764
rect -194 718 -148 764
rect -80 718 -34 764
rect 34 718 80 764
rect 148 718 194 764
rect 262 718 308 764
rect 376 718 422 764
rect 490 718 536 764
rect 604 718 650 764
rect 718 718 764 764
rect 832 718 878 764
rect 946 718 992 764
rect 1060 718 1106 764
rect 1174 718 1220 764
rect 1288 718 1334 764
rect 1402 718 1448 764
rect 1516 718 1562 764
rect 1630 718 1676 764
rect 1744 718 1790 764
rect 1858 718 1904 764
rect 1972 718 2018 764
rect 2086 718 2132 764
rect 2200 718 2246 764
rect 2314 718 2360 764
rect 2428 718 2474 764
rect 2542 718 2588 764
rect 2656 718 2702 764
rect 2770 718 2816 764
rect 2884 718 2930 764
rect 2998 718 3044 764
rect 3112 718 3158 764
rect 3226 718 3272 764
rect 3340 718 3386 764
rect 3454 718 3500 764
rect 3568 718 3614 764
rect 3682 718 3728 764
rect 3796 718 3842 764
rect 3910 718 3956 764
rect 4024 718 4070 764
rect 4138 718 4184 764
rect 4252 718 4298 764
rect 4366 718 4412 764
rect 4480 718 4526 764
rect 4594 718 4640 764
rect -4640 604 -4594 650
rect -4526 604 -4480 650
rect -4412 604 -4366 650
rect -4298 604 -4252 650
rect -4184 604 -4138 650
rect -4070 604 -4024 650
rect -3956 604 -3910 650
rect -3842 604 -3796 650
rect -3728 604 -3682 650
rect -3614 604 -3568 650
rect -3500 604 -3454 650
rect -3386 604 -3340 650
rect -3272 604 -3226 650
rect -3158 604 -3112 650
rect -3044 604 -2998 650
rect -2930 604 -2884 650
rect -2816 604 -2770 650
rect -2702 604 -2656 650
rect -2588 604 -2542 650
rect -2474 604 -2428 650
rect -2360 604 -2314 650
rect -2246 604 -2200 650
rect -2132 604 -2086 650
rect -2018 604 -1972 650
rect -1904 604 -1858 650
rect -1790 604 -1744 650
rect -1676 604 -1630 650
rect -1562 604 -1516 650
rect -1448 604 -1402 650
rect -1334 604 -1288 650
rect -1220 604 -1174 650
rect -1106 604 -1060 650
rect -992 604 -946 650
rect -878 604 -832 650
rect -764 604 -718 650
rect -650 604 -604 650
rect -536 604 -490 650
rect -422 604 -376 650
rect -308 604 -262 650
rect -194 604 -148 650
rect -80 604 -34 650
rect 34 604 80 650
rect 148 604 194 650
rect 262 604 308 650
rect 376 604 422 650
rect 490 604 536 650
rect 604 604 650 650
rect 718 604 764 650
rect 832 604 878 650
rect 946 604 992 650
rect 1060 604 1106 650
rect 1174 604 1220 650
rect 1288 604 1334 650
rect 1402 604 1448 650
rect 1516 604 1562 650
rect 1630 604 1676 650
rect 1744 604 1790 650
rect 1858 604 1904 650
rect 1972 604 2018 650
rect 2086 604 2132 650
rect 2200 604 2246 650
rect 2314 604 2360 650
rect 2428 604 2474 650
rect 2542 604 2588 650
rect 2656 604 2702 650
rect 2770 604 2816 650
rect 2884 604 2930 650
rect 2998 604 3044 650
rect 3112 604 3158 650
rect 3226 604 3272 650
rect 3340 604 3386 650
rect 3454 604 3500 650
rect 3568 604 3614 650
rect 3682 604 3728 650
rect 3796 604 3842 650
rect 3910 604 3956 650
rect 4024 604 4070 650
rect 4138 604 4184 650
rect 4252 604 4298 650
rect 4366 604 4412 650
rect 4480 604 4526 650
rect 4594 604 4640 650
rect -4640 490 -4594 536
rect -4526 490 -4480 536
rect -4412 490 -4366 536
rect -4298 490 -4252 536
rect -4184 490 -4138 536
rect -4070 490 -4024 536
rect -3956 490 -3910 536
rect -3842 490 -3796 536
rect -3728 490 -3682 536
rect -3614 490 -3568 536
rect -3500 490 -3454 536
rect -3386 490 -3340 536
rect -3272 490 -3226 536
rect -3158 490 -3112 536
rect -3044 490 -2998 536
rect -2930 490 -2884 536
rect -2816 490 -2770 536
rect -2702 490 -2656 536
rect -2588 490 -2542 536
rect -2474 490 -2428 536
rect -2360 490 -2314 536
rect -2246 490 -2200 536
rect -2132 490 -2086 536
rect -2018 490 -1972 536
rect -1904 490 -1858 536
rect -1790 490 -1744 536
rect -1676 490 -1630 536
rect -1562 490 -1516 536
rect -1448 490 -1402 536
rect -1334 490 -1288 536
rect -1220 490 -1174 536
rect -1106 490 -1060 536
rect -992 490 -946 536
rect -878 490 -832 536
rect -764 490 -718 536
rect -650 490 -604 536
rect -536 490 -490 536
rect -422 490 -376 536
rect -308 490 -262 536
rect -194 490 -148 536
rect -80 490 -34 536
rect 34 490 80 536
rect 148 490 194 536
rect 262 490 308 536
rect 376 490 422 536
rect 490 490 536 536
rect 604 490 650 536
rect 718 490 764 536
rect 832 490 878 536
rect 946 490 992 536
rect 1060 490 1106 536
rect 1174 490 1220 536
rect 1288 490 1334 536
rect 1402 490 1448 536
rect 1516 490 1562 536
rect 1630 490 1676 536
rect 1744 490 1790 536
rect 1858 490 1904 536
rect 1972 490 2018 536
rect 2086 490 2132 536
rect 2200 490 2246 536
rect 2314 490 2360 536
rect 2428 490 2474 536
rect 2542 490 2588 536
rect 2656 490 2702 536
rect 2770 490 2816 536
rect 2884 490 2930 536
rect 2998 490 3044 536
rect 3112 490 3158 536
rect 3226 490 3272 536
rect 3340 490 3386 536
rect 3454 490 3500 536
rect 3568 490 3614 536
rect 3682 490 3728 536
rect 3796 490 3842 536
rect 3910 490 3956 536
rect 4024 490 4070 536
rect 4138 490 4184 536
rect 4252 490 4298 536
rect 4366 490 4412 536
rect 4480 490 4526 536
rect 4594 490 4640 536
rect -4640 376 -4594 422
rect -4526 376 -4480 422
rect -4412 376 -4366 422
rect -4298 376 -4252 422
rect -4184 376 -4138 422
rect -4070 376 -4024 422
rect -3956 376 -3910 422
rect -3842 376 -3796 422
rect -3728 376 -3682 422
rect -3614 376 -3568 422
rect -3500 376 -3454 422
rect -3386 376 -3340 422
rect -3272 376 -3226 422
rect -3158 376 -3112 422
rect -3044 376 -2998 422
rect -2930 376 -2884 422
rect -2816 376 -2770 422
rect -2702 376 -2656 422
rect -2588 376 -2542 422
rect -2474 376 -2428 422
rect -2360 376 -2314 422
rect -2246 376 -2200 422
rect -2132 376 -2086 422
rect -2018 376 -1972 422
rect -1904 376 -1858 422
rect -1790 376 -1744 422
rect -1676 376 -1630 422
rect -1562 376 -1516 422
rect -1448 376 -1402 422
rect -1334 376 -1288 422
rect -1220 376 -1174 422
rect -1106 376 -1060 422
rect -992 376 -946 422
rect -878 376 -832 422
rect -764 376 -718 422
rect -650 376 -604 422
rect -536 376 -490 422
rect -422 376 -376 422
rect -308 376 -262 422
rect -194 376 -148 422
rect -80 376 -34 422
rect 34 376 80 422
rect 148 376 194 422
rect 262 376 308 422
rect 376 376 422 422
rect 490 376 536 422
rect 604 376 650 422
rect 718 376 764 422
rect 832 376 878 422
rect 946 376 992 422
rect 1060 376 1106 422
rect 1174 376 1220 422
rect 1288 376 1334 422
rect 1402 376 1448 422
rect 1516 376 1562 422
rect 1630 376 1676 422
rect 1744 376 1790 422
rect 1858 376 1904 422
rect 1972 376 2018 422
rect 2086 376 2132 422
rect 2200 376 2246 422
rect 2314 376 2360 422
rect 2428 376 2474 422
rect 2542 376 2588 422
rect 2656 376 2702 422
rect 2770 376 2816 422
rect 2884 376 2930 422
rect 2998 376 3044 422
rect 3112 376 3158 422
rect 3226 376 3272 422
rect 3340 376 3386 422
rect 3454 376 3500 422
rect 3568 376 3614 422
rect 3682 376 3728 422
rect 3796 376 3842 422
rect 3910 376 3956 422
rect 4024 376 4070 422
rect 4138 376 4184 422
rect 4252 376 4298 422
rect 4366 376 4412 422
rect 4480 376 4526 422
rect 4594 376 4640 422
rect -4640 262 -4594 308
rect -4526 262 -4480 308
rect -4412 262 -4366 308
rect -4298 262 -4252 308
rect -4184 262 -4138 308
rect -4070 262 -4024 308
rect -3956 262 -3910 308
rect -3842 262 -3796 308
rect -3728 262 -3682 308
rect -3614 262 -3568 308
rect -3500 262 -3454 308
rect -3386 262 -3340 308
rect -3272 262 -3226 308
rect -3158 262 -3112 308
rect -3044 262 -2998 308
rect -2930 262 -2884 308
rect -2816 262 -2770 308
rect -2702 262 -2656 308
rect -2588 262 -2542 308
rect -2474 262 -2428 308
rect -2360 262 -2314 308
rect -2246 262 -2200 308
rect -2132 262 -2086 308
rect -2018 262 -1972 308
rect -1904 262 -1858 308
rect -1790 262 -1744 308
rect -1676 262 -1630 308
rect -1562 262 -1516 308
rect -1448 262 -1402 308
rect -1334 262 -1288 308
rect -1220 262 -1174 308
rect -1106 262 -1060 308
rect -992 262 -946 308
rect -878 262 -832 308
rect -764 262 -718 308
rect -650 262 -604 308
rect -536 262 -490 308
rect -422 262 -376 308
rect -308 262 -262 308
rect -194 262 -148 308
rect -80 262 -34 308
rect 34 262 80 308
rect 148 262 194 308
rect 262 262 308 308
rect 376 262 422 308
rect 490 262 536 308
rect 604 262 650 308
rect 718 262 764 308
rect 832 262 878 308
rect 946 262 992 308
rect 1060 262 1106 308
rect 1174 262 1220 308
rect 1288 262 1334 308
rect 1402 262 1448 308
rect 1516 262 1562 308
rect 1630 262 1676 308
rect 1744 262 1790 308
rect 1858 262 1904 308
rect 1972 262 2018 308
rect 2086 262 2132 308
rect 2200 262 2246 308
rect 2314 262 2360 308
rect 2428 262 2474 308
rect 2542 262 2588 308
rect 2656 262 2702 308
rect 2770 262 2816 308
rect 2884 262 2930 308
rect 2998 262 3044 308
rect 3112 262 3158 308
rect 3226 262 3272 308
rect 3340 262 3386 308
rect 3454 262 3500 308
rect 3568 262 3614 308
rect 3682 262 3728 308
rect 3796 262 3842 308
rect 3910 262 3956 308
rect 4024 262 4070 308
rect 4138 262 4184 308
rect 4252 262 4298 308
rect 4366 262 4412 308
rect 4480 262 4526 308
rect 4594 262 4640 308
rect -4640 148 -4594 194
rect -4526 148 -4480 194
rect -4412 148 -4366 194
rect -4298 148 -4252 194
rect -4184 148 -4138 194
rect -4070 148 -4024 194
rect -3956 148 -3910 194
rect -3842 148 -3796 194
rect -3728 148 -3682 194
rect -3614 148 -3568 194
rect -3500 148 -3454 194
rect -3386 148 -3340 194
rect -3272 148 -3226 194
rect -3158 148 -3112 194
rect -3044 148 -2998 194
rect -2930 148 -2884 194
rect -2816 148 -2770 194
rect -2702 148 -2656 194
rect -2588 148 -2542 194
rect -2474 148 -2428 194
rect -2360 148 -2314 194
rect -2246 148 -2200 194
rect -2132 148 -2086 194
rect -2018 148 -1972 194
rect -1904 148 -1858 194
rect -1790 148 -1744 194
rect -1676 148 -1630 194
rect -1562 148 -1516 194
rect -1448 148 -1402 194
rect -1334 148 -1288 194
rect -1220 148 -1174 194
rect -1106 148 -1060 194
rect -992 148 -946 194
rect -878 148 -832 194
rect -764 148 -718 194
rect -650 148 -604 194
rect -536 148 -490 194
rect -422 148 -376 194
rect -308 148 -262 194
rect -194 148 -148 194
rect -80 148 -34 194
rect 34 148 80 194
rect 148 148 194 194
rect 262 148 308 194
rect 376 148 422 194
rect 490 148 536 194
rect 604 148 650 194
rect 718 148 764 194
rect 832 148 878 194
rect 946 148 992 194
rect 1060 148 1106 194
rect 1174 148 1220 194
rect 1288 148 1334 194
rect 1402 148 1448 194
rect 1516 148 1562 194
rect 1630 148 1676 194
rect 1744 148 1790 194
rect 1858 148 1904 194
rect 1972 148 2018 194
rect 2086 148 2132 194
rect 2200 148 2246 194
rect 2314 148 2360 194
rect 2428 148 2474 194
rect 2542 148 2588 194
rect 2656 148 2702 194
rect 2770 148 2816 194
rect 2884 148 2930 194
rect 2998 148 3044 194
rect 3112 148 3158 194
rect 3226 148 3272 194
rect 3340 148 3386 194
rect 3454 148 3500 194
rect 3568 148 3614 194
rect 3682 148 3728 194
rect 3796 148 3842 194
rect 3910 148 3956 194
rect 4024 148 4070 194
rect 4138 148 4184 194
rect 4252 148 4298 194
rect 4366 148 4412 194
rect 4480 148 4526 194
rect 4594 148 4640 194
rect -4640 34 -4594 80
rect -4526 34 -4480 80
rect -4412 34 -4366 80
rect -4298 34 -4252 80
rect -4184 34 -4138 80
rect -4070 34 -4024 80
rect -3956 34 -3910 80
rect -3842 34 -3796 80
rect -3728 34 -3682 80
rect -3614 34 -3568 80
rect -3500 34 -3454 80
rect -3386 34 -3340 80
rect -3272 34 -3226 80
rect -3158 34 -3112 80
rect -3044 34 -2998 80
rect -2930 34 -2884 80
rect -2816 34 -2770 80
rect -2702 34 -2656 80
rect -2588 34 -2542 80
rect -2474 34 -2428 80
rect -2360 34 -2314 80
rect -2246 34 -2200 80
rect -2132 34 -2086 80
rect -2018 34 -1972 80
rect -1904 34 -1858 80
rect -1790 34 -1744 80
rect -1676 34 -1630 80
rect -1562 34 -1516 80
rect -1448 34 -1402 80
rect -1334 34 -1288 80
rect -1220 34 -1174 80
rect -1106 34 -1060 80
rect -992 34 -946 80
rect -878 34 -832 80
rect -764 34 -718 80
rect -650 34 -604 80
rect -536 34 -490 80
rect -422 34 -376 80
rect -308 34 -262 80
rect -194 34 -148 80
rect -80 34 -34 80
rect 34 34 80 80
rect 148 34 194 80
rect 262 34 308 80
rect 376 34 422 80
rect 490 34 536 80
rect 604 34 650 80
rect 718 34 764 80
rect 832 34 878 80
rect 946 34 992 80
rect 1060 34 1106 80
rect 1174 34 1220 80
rect 1288 34 1334 80
rect 1402 34 1448 80
rect 1516 34 1562 80
rect 1630 34 1676 80
rect 1744 34 1790 80
rect 1858 34 1904 80
rect 1972 34 2018 80
rect 2086 34 2132 80
rect 2200 34 2246 80
rect 2314 34 2360 80
rect 2428 34 2474 80
rect 2542 34 2588 80
rect 2656 34 2702 80
rect 2770 34 2816 80
rect 2884 34 2930 80
rect 2998 34 3044 80
rect 3112 34 3158 80
rect 3226 34 3272 80
rect 3340 34 3386 80
rect 3454 34 3500 80
rect 3568 34 3614 80
rect 3682 34 3728 80
rect 3796 34 3842 80
rect 3910 34 3956 80
rect 4024 34 4070 80
rect 4138 34 4184 80
rect 4252 34 4298 80
rect 4366 34 4412 80
rect 4480 34 4526 80
rect 4594 34 4640 80
rect -4640 -80 -4594 -34
rect -4526 -80 -4480 -34
rect -4412 -80 -4366 -34
rect -4298 -80 -4252 -34
rect -4184 -80 -4138 -34
rect -4070 -80 -4024 -34
rect -3956 -80 -3910 -34
rect -3842 -80 -3796 -34
rect -3728 -80 -3682 -34
rect -3614 -80 -3568 -34
rect -3500 -80 -3454 -34
rect -3386 -80 -3340 -34
rect -3272 -80 -3226 -34
rect -3158 -80 -3112 -34
rect -3044 -80 -2998 -34
rect -2930 -80 -2884 -34
rect -2816 -80 -2770 -34
rect -2702 -80 -2656 -34
rect -2588 -80 -2542 -34
rect -2474 -80 -2428 -34
rect -2360 -80 -2314 -34
rect -2246 -80 -2200 -34
rect -2132 -80 -2086 -34
rect -2018 -80 -1972 -34
rect -1904 -80 -1858 -34
rect -1790 -80 -1744 -34
rect -1676 -80 -1630 -34
rect -1562 -80 -1516 -34
rect -1448 -80 -1402 -34
rect -1334 -80 -1288 -34
rect -1220 -80 -1174 -34
rect -1106 -80 -1060 -34
rect -992 -80 -946 -34
rect -878 -80 -832 -34
rect -764 -80 -718 -34
rect -650 -80 -604 -34
rect -536 -80 -490 -34
rect -422 -80 -376 -34
rect -308 -80 -262 -34
rect -194 -80 -148 -34
rect -80 -80 -34 -34
rect 34 -80 80 -34
rect 148 -80 194 -34
rect 262 -80 308 -34
rect 376 -80 422 -34
rect 490 -80 536 -34
rect 604 -80 650 -34
rect 718 -80 764 -34
rect 832 -80 878 -34
rect 946 -80 992 -34
rect 1060 -80 1106 -34
rect 1174 -80 1220 -34
rect 1288 -80 1334 -34
rect 1402 -80 1448 -34
rect 1516 -80 1562 -34
rect 1630 -80 1676 -34
rect 1744 -80 1790 -34
rect 1858 -80 1904 -34
rect 1972 -80 2018 -34
rect 2086 -80 2132 -34
rect 2200 -80 2246 -34
rect 2314 -80 2360 -34
rect 2428 -80 2474 -34
rect 2542 -80 2588 -34
rect 2656 -80 2702 -34
rect 2770 -80 2816 -34
rect 2884 -80 2930 -34
rect 2998 -80 3044 -34
rect 3112 -80 3158 -34
rect 3226 -80 3272 -34
rect 3340 -80 3386 -34
rect 3454 -80 3500 -34
rect 3568 -80 3614 -34
rect 3682 -80 3728 -34
rect 3796 -80 3842 -34
rect 3910 -80 3956 -34
rect 4024 -80 4070 -34
rect 4138 -80 4184 -34
rect 4252 -80 4298 -34
rect 4366 -80 4412 -34
rect 4480 -80 4526 -34
rect 4594 -80 4640 -34
rect -4640 -194 -4594 -148
rect -4526 -194 -4480 -148
rect -4412 -194 -4366 -148
rect -4298 -194 -4252 -148
rect -4184 -194 -4138 -148
rect -4070 -194 -4024 -148
rect -3956 -194 -3910 -148
rect -3842 -194 -3796 -148
rect -3728 -194 -3682 -148
rect -3614 -194 -3568 -148
rect -3500 -194 -3454 -148
rect -3386 -194 -3340 -148
rect -3272 -194 -3226 -148
rect -3158 -194 -3112 -148
rect -3044 -194 -2998 -148
rect -2930 -194 -2884 -148
rect -2816 -194 -2770 -148
rect -2702 -194 -2656 -148
rect -2588 -194 -2542 -148
rect -2474 -194 -2428 -148
rect -2360 -194 -2314 -148
rect -2246 -194 -2200 -148
rect -2132 -194 -2086 -148
rect -2018 -194 -1972 -148
rect -1904 -194 -1858 -148
rect -1790 -194 -1744 -148
rect -1676 -194 -1630 -148
rect -1562 -194 -1516 -148
rect -1448 -194 -1402 -148
rect -1334 -194 -1288 -148
rect -1220 -194 -1174 -148
rect -1106 -194 -1060 -148
rect -992 -194 -946 -148
rect -878 -194 -832 -148
rect -764 -194 -718 -148
rect -650 -194 -604 -148
rect -536 -194 -490 -148
rect -422 -194 -376 -148
rect -308 -194 -262 -148
rect -194 -194 -148 -148
rect -80 -194 -34 -148
rect 34 -194 80 -148
rect 148 -194 194 -148
rect 262 -194 308 -148
rect 376 -194 422 -148
rect 490 -194 536 -148
rect 604 -194 650 -148
rect 718 -194 764 -148
rect 832 -194 878 -148
rect 946 -194 992 -148
rect 1060 -194 1106 -148
rect 1174 -194 1220 -148
rect 1288 -194 1334 -148
rect 1402 -194 1448 -148
rect 1516 -194 1562 -148
rect 1630 -194 1676 -148
rect 1744 -194 1790 -148
rect 1858 -194 1904 -148
rect 1972 -194 2018 -148
rect 2086 -194 2132 -148
rect 2200 -194 2246 -148
rect 2314 -194 2360 -148
rect 2428 -194 2474 -148
rect 2542 -194 2588 -148
rect 2656 -194 2702 -148
rect 2770 -194 2816 -148
rect 2884 -194 2930 -148
rect 2998 -194 3044 -148
rect 3112 -194 3158 -148
rect 3226 -194 3272 -148
rect 3340 -194 3386 -148
rect 3454 -194 3500 -148
rect 3568 -194 3614 -148
rect 3682 -194 3728 -148
rect 3796 -194 3842 -148
rect 3910 -194 3956 -148
rect 4024 -194 4070 -148
rect 4138 -194 4184 -148
rect 4252 -194 4298 -148
rect 4366 -194 4412 -148
rect 4480 -194 4526 -148
rect 4594 -194 4640 -148
rect -4640 -308 -4594 -262
rect -4526 -308 -4480 -262
rect -4412 -308 -4366 -262
rect -4298 -308 -4252 -262
rect -4184 -308 -4138 -262
rect -4070 -308 -4024 -262
rect -3956 -308 -3910 -262
rect -3842 -308 -3796 -262
rect -3728 -308 -3682 -262
rect -3614 -308 -3568 -262
rect -3500 -308 -3454 -262
rect -3386 -308 -3340 -262
rect -3272 -308 -3226 -262
rect -3158 -308 -3112 -262
rect -3044 -308 -2998 -262
rect -2930 -308 -2884 -262
rect -2816 -308 -2770 -262
rect -2702 -308 -2656 -262
rect -2588 -308 -2542 -262
rect -2474 -308 -2428 -262
rect -2360 -308 -2314 -262
rect -2246 -308 -2200 -262
rect -2132 -308 -2086 -262
rect -2018 -308 -1972 -262
rect -1904 -308 -1858 -262
rect -1790 -308 -1744 -262
rect -1676 -308 -1630 -262
rect -1562 -308 -1516 -262
rect -1448 -308 -1402 -262
rect -1334 -308 -1288 -262
rect -1220 -308 -1174 -262
rect -1106 -308 -1060 -262
rect -992 -308 -946 -262
rect -878 -308 -832 -262
rect -764 -308 -718 -262
rect -650 -308 -604 -262
rect -536 -308 -490 -262
rect -422 -308 -376 -262
rect -308 -308 -262 -262
rect -194 -308 -148 -262
rect -80 -308 -34 -262
rect 34 -308 80 -262
rect 148 -308 194 -262
rect 262 -308 308 -262
rect 376 -308 422 -262
rect 490 -308 536 -262
rect 604 -308 650 -262
rect 718 -308 764 -262
rect 832 -308 878 -262
rect 946 -308 992 -262
rect 1060 -308 1106 -262
rect 1174 -308 1220 -262
rect 1288 -308 1334 -262
rect 1402 -308 1448 -262
rect 1516 -308 1562 -262
rect 1630 -308 1676 -262
rect 1744 -308 1790 -262
rect 1858 -308 1904 -262
rect 1972 -308 2018 -262
rect 2086 -308 2132 -262
rect 2200 -308 2246 -262
rect 2314 -308 2360 -262
rect 2428 -308 2474 -262
rect 2542 -308 2588 -262
rect 2656 -308 2702 -262
rect 2770 -308 2816 -262
rect 2884 -308 2930 -262
rect 2998 -308 3044 -262
rect 3112 -308 3158 -262
rect 3226 -308 3272 -262
rect 3340 -308 3386 -262
rect 3454 -308 3500 -262
rect 3568 -308 3614 -262
rect 3682 -308 3728 -262
rect 3796 -308 3842 -262
rect 3910 -308 3956 -262
rect 4024 -308 4070 -262
rect 4138 -308 4184 -262
rect 4252 -308 4298 -262
rect 4366 -308 4412 -262
rect 4480 -308 4526 -262
rect 4594 -308 4640 -262
rect -4640 -422 -4594 -376
rect -4526 -422 -4480 -376
rect -4412 -422 -4366 -376
rect -4298 -422 -4252 -376
rect -4184 -422 -4138 -376
rect -4070 -422 -4024 -376
rect -3956 -422 -3910 -376
rect -3842 -422 -3796 -376
rect -3728 -422 -3682 -376
rect -3614 -422 -3568 -376
rect -3500 -422 -3454 -376
rect -3386 -422 -3340 -376
rect -3272 -422 -3226 -376
rect -3158 -422 -3112 -376
rect -3044 -422 -2998 -376
rect -2930 -422 -2884 -376
rect -2816 -422 -2770 -376
rect -2702 -422 -2656 -376
rect -2588 -422 -2542 -376
rect -2474 -422 -2428 -376
rect -2360 -422 -2314 -376
rect -2246 -422 -2200 -376
rect -2132 -422 -2086 -376
rect -2018 -422 -1972 -376
rect -1904 -422 -1858 -376
rect -1790 -422 -1744 -376
rect -1676 -422 -1630 -376
rect -1562 -422 -1516 -376
rect -1448 -422 -1402 -376
rect -1334 -422 -1288 -376
rect -1220 -422 -1174 -376
rect -1106 -422 -1060 -376
rect -992 -422 -946 -376
rect -878 -422 -832 -376
rect -764 -422 -718 -376
rect -650 -422 -604 -376
rect -536 -422 -490 -376
rect -422 -422 -376 -376
rect -308 -422 -262 -376
rect -194 -422 -148 -376
rect -80 -422 -34 -376
rect 34 -422 80 -376
rect 148 -422 194 -376
rect 262 -422 308 -376
rect 376 -422 422 -376
rect 490 -422 536 -376
rect 604 -422 650 -376
rect 718 -422 764 -376
rect 832 -422 878 -376
rect 946 -422 992 -376
rect 1060 -422 1106 -376
rect 1174 -422 1220 -376
rect 1288 -422 1334 -376
rect 1402 -422 1448 -376
rect 1516 -422 1562 -376
rect 1630 -422 1676 -376
rect 1744 -422 1790 -376
rect 1858 -422 1904 -376
rect 1972 -422 2018 -376
rect 2086 -422 2132 -376
rect 2200 -422 2246 -376
rect 2314 -422 2360 -376
rect 2428 -422 2474 -376
rect 2542 -422 2588 -376
rect 2656 -422 2702 -376
rect 2770 -422 2816 -376
rect 2884 -422 2930 -376
rect 2998 -422 3044 -376
rect 3112 -422 3158 -376
rect 3226 -422 3272 -376
rect 3340 -422 3386 -376
rect 3454 -422 3500 -376
rect 3568 -422 3614 -376
rect 3682 -422 3728 -376
rect 3796 -422 3842 -376
rect 3910 -422 3956 -376
rect 4024 -422 4070 -376
rect 4138 -422 4184 -376
rect 4252 -422 4298 -376
rect 4366 -422 4412 -376
rect 4480 -422 4526 -376
rect 4594 -422 4640 -376
rect -4640 -536 -4594 -490
rect -4526 -536 -4480 -490
rect -4412 -536 -4366 -490
rect -4298 -536 -4252 -490
rect -4184 -536 -4138 -490
rect -4070 -536 -4024 -490
rect -3956 -536 -3910 -490
rect -3842 -536 -3796 -490
rect -3728 -536 -3682 -490
rect -3614 -536 -3568 -490
rect -3500 -536 -3454 -490
rect -3386 -536 -3340 -490
rect -3272 -536 -3226 -490
rect -3158 -536 -3112 -490
rect -3044 -536 -2998 -490
rect -2930 -536 -2884 -490
rect -2816 -536 -2770 -490
rect -2702 -536 -2656 -490
rect -2588 -536 -2542 -490
rect -2474 -536 -2428 -490
rect -2360 -536 -2314 -490
rect -2246 -536 -2200 -490
rect -2132 -536 -2086 -490
rect -2018 -536 -1972 -490
rect -1904 -536 -1858 -490
rect -1790 -536 -1744 -490
rect -1676 -536 -1630 -490
rect -1562 -536 -1516 -490
rect -1448 -536 -1402 -490
rect -1334 -536 -1288 -490
rect -1220 -536 -1174 -490
rect -1106 -536 -1060 -490
rect -992 -536 -946 -490
rect -878 -536 -832 -490
rect -764 -536 -718 -490
rect -650 -536 -604 -490
rect -536 -536 -490 -490
rect -422 -536 -376 -490
rect -308 -536 -262 -490
rect -194 -536 -148 -490
rect -80 -536 -34 -490
rect 34 -536 80 -490
rect 148 -536 194 -490
rect 262 -536 308 -490
rect 376 -536 422 -490
rect 490 -536 536 -490
rect 604 -536 650 -490
rect 718 -536 764 -490
rect 832 -536 878 -490
rect 946 -536 992 -490
rect 1060 -536 1106 -490
rect 1174 -536 1220 -490
rect 1288 -536 1334 -490
rect 1402 -536 1448 -490
rect 1516 -536 1562 -490
rect 1630 -536 1676 -490
rect 1744 -536 1790 -490
rect 1858 -536 1904 -490
rect 1972 -536 2018 -490
rect 2086 -536 2132 -490
rect 2200 -536 2246 -490
rect 2314 -536 2360 -490
rect 2428 -536 2474 -490
rect 2542 -536 2588 -490
rect 2656 -536 2702 -490
rect 2770 -536 2816 -490
rect 2884 -536 2930 -490
rect 2998 -536 3044 -490
rect 3112 -536 3158 -490
rect 3226 -536 3272 -490
rect 3340 -536 3386 -490
rect 3454 -536 3500 -490
rect 3568 -536 3614 -490
rect 3682 -536 3728 -490
rect 3796 -536 3842 -490
rect 3910 -536 3956 -490
rect 4024 -536 4070 -490
rect 4138 -536 4184 -490
rect 4252 -536 4298 -490
rect 4366 -536 4412 -490
rect 4480 -536 4526 -490
rect 4594 -536 4640 -490
rect -4640 -650 -4594 -604
rect -4526 -650 -4480 -604
rect -4412 -650 -4366 -604
rect -4298 -650 -4252 -604
rect -4184 -650 -4138 -604
rect -4070 -650 -4024 -604
rect -3956 -650 -3910 -604
rect -3842 -650 -3796 -604
rect -3728 -650 -3682 -604
rect -3614 -650 -3568 -604
rect -3500 -650 -3454 -604
rect -3386 -650 -3340 -604
rect -3272 -650 -3226 -604
rect -3158 -650 -3112 -604
rect -3044 -650 -2998 -604
rect -2930 -650 -2884 -604
rect -2816 -650 -2770 -604
rect -2702 -650 -2656 -604
rect -2588 -650 -2542 -604
rect -2474 -650 -2428 -604
rect -2360 -650 -2314 -604
rect -2246 -650 -2200 -604
rect -2132 -650 -2086 -604
rect -2018 -650 -1972 -604
rect -1904 -650 -1858 -604
rect -1790 -650 -1744 -604
rect -1676 -650 -1630 -604
rect -1562 -650 -1516 -604
rect -1448 -650 -1402 -604
rect -1334 -650 -1288 -604
rect -1220 -650 -1174 -604
rect -1106 -650 -1060 -604
rect -992 -650 -946 -604
rect -878 -650 -832 -604
rect -764 -650 -718 -604
rect -650 -650 -604 -604
rect -536 -650 -490 -604
rect -422 -650 -376 -604
rect -308 -650 -262 -604
rect -194 -650 -148 -604
rect -80 -650 -34 -604
rect 34 -650 80 -604
rect 148 -650 194 -604
rect 262 -650 308 -604
rect 376 -650 422 -604
rect 490 -650 536 -604
rect 604 -650 650 -604
rect 718 -650 764 -604
rect 832 -650 878 -604
rect 946 -650 992 -604
rect 1060 -650 1106 -604
rect 1174 -650 1220 -604
rect 1288 -650 1334 -604
rect 1402 -650 1448 -604
rect 1516 -650 1562 -604
rect 1630 -650 1676 -604
rect 1744 -650 1790 -604
rect 1858 -650 1904 -604
rect 1972 -650 2018 -604
rect 2086 -650 2132 -604
rect 2200 -650 2246 -604
rect 2314 -650 2360 -604
rect 2428 -650 2474 -604
rect 2542 -650 2588 -604
rect 2656 -650 2702 -604
rect 2770 -650 2816 -604
rect 2884 -650 2930 -604
rect 2998 -650 3044 -604
rect 3112 -650 3158 -604
rect 3226 -650 3272 -604
rect 3340 -650 3386 -604
rect 3454 -650 3500 -604
rect 3568 -650 3614 -604
rect 3682 -650 3728 -604
rect 3796 -650 3842 -604
rect 3910 -650 3956 -604
rect 4024 -650 4070 -604
rect 4138 -650 4184 -604
rect 4252 -650 4298 -604
rect 4366 -650 4412 -604
rect 4480 -650 4526 -604
rect 4594 -650 4640 -604
rect -4640 -764 -4594 -718
rect -4526 -764 -4480 -718
rect -4412 -764 -4366 -718
rect -4298 -764 -4252 -718
rect -4184 -764 -4138 -718
rect -4070 -764 -4024 -718
rect -3956 -764 -3910 -718
rect -3842 -764 -3796 -718
rect -3728 -764 -3682 -718
rect -3614 -764 -3568 -718
rect -3500 -764 -3454 -718
rect -3386 -764 -3340 -718
rect -3272 -764 -3226 -718
rect -3158 -764 -3112 -718
rect -3044 -764 -2998 -718
rect -2930 -764 -2884 -718
rect -2816 -764 -2770 -718
rect -2702 -764 -2656 -718
rect -2588 -764 -2542 -718
rect -2474 -764 -2428 -718
rect -2360 -764 -2314 -718
rect -2246 -764 -2200 -718
rect -2132 -764 -2086 -718
rect -2018 -764 -1972 -718
rect -1904 -764 -1858 -718
rect -1790 -764 -1744 -718
rect -1676 -764 -1630 -718
rect -1562 -764 -1516 -718
rect -1448 -764 -1402 -718
rect -1334 -764 -1288 -718
rect -1220 -764 -1174 -718
rect -1106 -764 -1060 -718
rect -992 -764 -946 -718
rect -878 -764 -832 -718
rect -764 -764 -718 -718
rect -650 -764 -604 -718
rect -536 -764 -490 -718
rect -422 -764 -376 -718
rect -308 -764 -262 -718
rect -194 -764 -148 -718
rect -80 -764 -34 -718
rect 34 -764 80 -718
rect 148 -764 194 -718
rect 262 -764 308 -718
rect 376 -764 422 -718
rect 490 -764 536 -718
rect 604 -764 650 -718
rect 718 -764 764 -718
rect 832 -764 878 -718
rect 946 -764 992 -718
rect 1060 -764 1106 -718
rect 1174 -764 1220 -718
rect 1288 -764 1334 -718
rect 1402 -764 1448 -718
rect 1516 -764 1562 -718
rect 1630 -764 1676 -718
rect 1744 -764 1790 -718
rect 1858 -764 1904 -718
rect 1972 -764 2018 -718
rect 2086 -764 2132 -718
rect 2200 -764 2246 -718
rect 2314 -764 2360 -718
rect 2428 -764 2474 -718
rect 2542 -764 2588 -718
rect 2656 -764 2702 -718
rect 2770 -764 2816 -718
rect 2884 -764 2930 -718
rect 2998 -764 3044 -718
rect 3112 -764 3158 -718
rect 3226 -764 3272 -718
rect 3340 -764 3386 -718
rect 3454 -764 3500 -718
rect 3568 -764 3614 -718
rect 3682 -764 3728 -718
rect 3796 -764 3842 -718
rect 3910 -764 3956 -718
rect 4024 -764 4070 -718
rect 4138 -764 4184 -718
rect 4252 -764 4298 -718
rect 4366 -764 4412 -718
rect 4480 -764 4526 -718
rect 4594 -764 4640 -718
<< metal1 >>
rect -4651 764 4651 775
rect -4651 718 -4640 764
rect -4594 718 -4526 764
rect -4480 718 -4412 764
rect -4366 718 -4298 764
rect -4252 718 -4184 764
rect -4138 718 -4070 764
rect -4024 718 -3956 764
rect -3910 718 -3842 764
rect -3796 718 -3728 764
rect -3682 718 -3614 764
rect -3568 718 -3500 764
rect -3454 718 -3386 764
rect -3340 718 -3272 764
rect -3226 718 -3158 764
rect -3112 718 -3044 764
rect -2998 718 -2930 764
rect -2884 718 -2816 764
rect -2770 718 -2702 764
rect -2656 718 -2588 764
rect -2542 718 -2474 764
rect -2428 718 -2360 764
rect -2314 718 -2246 764
rect -2200 718 -2132 764
rect -2086 718 -2018 764
rect -1972 718 -1904 764
rect -1858 718 -1790 764
rect -1744 718 -1676 764
rect -1630 718 -1562 764
rect -1516 718 -1448 764
rect -1402 718 -1334 764
rect -1288 718 -1220 764
rect -1174 718 -1106 764
rect -1060 718 -992 764
rect -946 718 -878 764
rect -832 718 -764 764
rect -718 718 -650 764
rect -604 718 -536 764
rect -490 718 -422 764
rect -376 718 -308 764
rect -262 718 -194 764
rect -148 718 -80 764
rect -34 718 34 764
rect 80 718 148 764
rect 194 718 262 764
rect 308 718 376 764
rect 422 718 490 764
rect 536 718 604 764
rect 650 718 718 764
rect 764 718 832 764
rect 878 718 946 764
rect 992 718 1060 764
rect 1106 718 1174 764
rect 1220 718 1288 764
rect 1334 718 1402 764
rect 1448 718 1516 764
rect 1562 718 1630 764
rect 1676 718 1744 764
rect 1790 718 1858 764
rect 1904 718 1972 764
rect 2018 718 2086 764
rect 2132 718 2200 764
rect 2246 718 2314 764
rect 2360 718 2428 764
rect 2474 718 2542 764
rect 2588 718 2656 764
rect 2702 718 2770 764
rect 2816 718 2884 764
rect 2930 718 2998 764
rect 3044 718 3112 764
rect 3158 718 3226 764
rect 3272 718 3340 764
rect 3386 718 3454 764
rect 3500 718 3568 764
rect 3614 718 3682 764
rect 3728 718 3796 764
rect 3842 718 3910 764
rect 3956 718 4024 764
rect 4070 718 4138 764
rect 4184 718 4252 764
rect 4298 718 4366 764
rect 4412 718 4480 764
rect 4526 718 4594 764
rect 4640 718 4651 764
rect -4651 650 4651 718
rect -4651 604 -4640 650
rect -4594 604 -4526 650
rect -4480 604 -4412 650
rect -4366 604 -4298 650
rect -4252 604 -4184 650
rect -4138 604 -4070 650
rect -4024 604 -3956 650
rect -3910 604 -3842 650
rect -3796 604 -3728 650
rect -3682 604 -3614 650
rect -3568 604 -3500 650
rect -3454 604 -3386 650
rect -3340 604 -3272 650
rect -3226 604 -3158 650
rect -3112 604 -3044 650
rect -2998 604 -2930 650
rect -2884 604 -2816 650
rect -2770 604 -2702 650
rect -2656 604 -2588 650
rect -2542 604 -2474 650
rect -2428 604 -2360 650
rect -2314 604 -2246 650
rect -2200 604 -2132 650
rect -2086 604 -2018 650
rect -1972 604 -1904 650
rect -1858 604 -1790 650
rect -1744 604 -1676 650
rect -1630 604 -1562 650
rect -1516 604 -1448 650
rect -1402 604 -1334 650
rect -1288 604 -1220 650
rect -1174 604 -1106 650
rect -1060 604 -992 650
rect -946 604 -878 650
rect -832 604 -764 650
rect -718 604 -650 650
rect -604 604 -536 650
rect -490 604 -422 650
rect -376 604 -308 650
rect -262 604 -194 650
rect -148 604 -80 650
rect -34 604 34 650
rect 80 604 148 650
rect 194 604 262 650
rect 308 604 376 650
rect 422 604 490 650
rect 536 604 604 650
rect 650 604 718 650
rect 764 604 832 650
rect 878 604 946 650
rect 992 604 1060 650
rect 1106 604 1174 650
rect 1220 604 1288 650
rect 1334 604 1402 650
rect 1448 604 1516 650
rect 1562 604 1630 650
rect 1676 604 1744 650
rect 1790 604 1858 650
rect 1904 604 1972 650
rect 2018 604 2086 650
rect 2132 604 2200 650
rect 2246 604 2314 650
rect 2360 604 2428 650
rect 2474 604 2542 650
rect 2588 604 2656 650
rect 2702 604 2770 650
rect 2816 604 2884 650
rect 2930 604 2998 650
rect 3044 604 3112 650
rect 3158 604 3226 650
rect 3272 604 3340 650
rect 3386 604 3454 650
rect 3500 604 3568 650
rect 3614 604 3682 650
rect 3728 604 3796 650
rect 3842 604 3910 650
rect 3956 604 4024 650
rect 4070 604 4138 650
rect 4184 604 4252 650
rect 4298 604 4366 650
rect 4412 604 4480 650
rect 4526 604 4594 650
rect 4640 604 4651 650
rect -4651 536 4651 604
rect -4651 490 -4640 536
rect -4594 490 -4526 536
rect -4480 490 -4412 536
rect -4366 490 -4298 536
rect -4252 490 -4184 536
rect -4138 490 -4070 536
rect -4024 490 -3956 536
rect -3910 490 -3842 536
rect -3796 490 -3728 536
rect -3682 490 -3614 536
rect -3568 490 -3500 536
rect -3454 490 -3386 536
rect -3340 490 -3272 536
rect -3226 490 -3158 536
rect -3112 490 -3044 536
rect -2998 490 -2930 536
rect -2884 490 -2816 536
rect -2770 490 -2702 536
rect -2656 490 -2588 536
rect -2542 490 -2474 536
rect -2428 490 -2360 536
rect -2314 490 -2246 536
rect -2200 490 -2132 536
rect -2086 490 -2018 536
rect -1972 490 -1904 536
rect -1858 490 -1790 536
rect -1744 490 -1676 536
rect -1630 490 -1562 536
rect -1516 490 -1448 536
rect -1402 490 -1334 536
rect -1288 490 -1220 536
rect -1174 490 -1106 536
rect -1060 490 -992 536
rect -946 490 -878 536
rect -832 490 -764 536
rect -718 490 -650 536
rect -604 490 -536 536
rect -490 490 -422 536
rect -376 490 -308 536
rect -262 490 -194 536
rect -148 490 -80 536
rect -34 490 34 536
rect 80 490 148 536
rect 194 490 262 536
rect 308 490 376 536
rect 422 490 490 536
rect 536 490 604 536
rect 650 490 718 536
rect 764 490 832 536
rect 878 490 946 536
rect 992 490 1060 536
rect 1106 490 1174 536
rect 1220 490 1288 536
rect 1334 490 1402 536
rect 1448 490 1516 536
rect 1562 490 1630 536
rect 1676 490 1744 536
rect 1790 490 1858 536
rect 1904 490 1972 536
rect 2018 490 2086 536
rect 2132 490 2200 536
rect 2246 490 2314 536
rect 2360 490 2428 536
rect 2474 490 2542 536
rect 2588 490 2656 536
rect 2702 490 2770 536
rect 2816 490 2884 536
rect 2930 490 2998 536
rect 3044 490 3112 536
rect 3158 490 3226 536
rect 3272 490 3340 536
rect 3386 490 3454 536
rect 3500 490 3568 536
rect 3614 490 3682 536
rect 3728 490 3796 536
rect 3842 490 3910 536
rect 3956 490 4024 536
rect 4070 490 4138 536
rect 4184 490 4252 536
rect 4298 490 4366 536
rect 4412 490 4480 536
rect 4526 490 4594 536
rect 4640 490 4651 536
rect -4651 422 4651 490
rect -4651 376 -4640 422
rect -4594 376 -4526 422
rect -4480 376 -4412 422
rect -4366 376 -4298 422
rect -4252 376 -4184 422
rect -4138 376 -4070 422
rect -4024 376 -3956 422
rect -3910 376 -3842 422
rect -3796 376 -3728 422
rect -3682 376 -3614 422
rect -3568 376 -3500 422
rect -3454 376 -3386 422
rect -3340 376 -3272 422
rect -3226 376 -3158 422
rect -3112 376 -3044 422
rect -2998 376 -2930 422
rect -2884 376 -2816 422
rect -2770 376 -2702 422
rect -2656 376 -2588 422
rect -2542 376 -2474 422
rect -2428 376 -2360 422
rect -2314 376 -2246 422
rect -2200 376 -2132 422
rect -2086 376 -2018 422
rect -1972 376 -1904 422
rect -1858 376 -1790 422
rect -1744 376 -1676 422
rect -1630 376 -1562 422
rect -1516 376 -1448 422
rect -1402 376 -1334 422
rect -1288 376 -1220 422
rect -1174 376 -1106 422
rect -1060 376 -992 422
rect -946 376 -878 422
rect -832 376 -764 422
rect -718 376 -650 422
rect -604 376 -536 422
rect -490 376 -422 422
rect -376 376 -308 422
rect -262 376 -194 422
rect -148 376 -80 422
rect -34 376 34 422
rect 80 376 148 422
rect 194 376 262 422
rect 308 376 376 422
rect 422 376 490 422
rect 536 376 604 422
rect 650 376 718 422
rect 764 376 832 422
rect 878 376 946 422
rect 992 376 1060 422
rect 1106 376 1174 422
rect 1220 376 1288 422
rect 1334 376 1402 422
rect 1448 376 1516 422
rect 1562 376 1630 422
rect 1676 376 1744 422
rect 1790 376 1858 422
rect 1904 376 1972 422
rect 2018 376 2086 422
rect 2132 376 2200 422
rect 2246 376 2314 422
rect 2360 376 2428 422
rect 2474 376 2542 422
rect 2588 376 2656 422
rect 2702 376 2770 422
rect 2816 376 2884 422
rect 2930 376 2998 422
rect 3044 376 3112 422
rect 3158 376 3226 422
rect 3272 376 3340 422
rect 3386 376 3454 422
rect 3500 376 3568 422
rect 3614 376 3682 422
rect 3728 376 3796 422
rect 3842 376 3910 422
rect 3956 376 4024 422
rect 4070 376 4138 422
rect 4184 376 4252 422
rect 4298 376 4366 422
rect 4412 376 4480 422
rect 4526 376 4594 422
rect 4640 376 4651 422
rect -4651 308 4651 376
rect -4651 262 -4640 308
rect -4594 262 -4526 308
rect -4480 262 -4412 308
rect -4366 262 -4298 308
rect -4252 262 -4184 308
rect -4138 262 -4070 308
rect -4024 262 -3956 308
rect -3910 262 -3842 308
rect -3796 262 -3728 308
rect -3682 262 -3614 308
rect -3568 262 -3500 308
rect -3454 262 -3386 308
rect -3340 262 -3272 308
rect -3226 262 -3158 308
rect -3112 262 -3044 308
rect -2998 262 -2930 308
rect -2884 262 -2816 308
rect -2770 262 -2702 308
rect -2656 262 -2588 308
rect -2542 262 -2474 308
rect -2428 262 -2360 308
rect -2314 262 -2246 308
rect -2200 262 -2132 308
rect -2086 262 -2018 308
rect -1972 262 -1904 308
rect -1858 262 -1790 308
rect -1744 262 -1676 308
rect -1630 262 -1562 308
rect -1516 262 -1448 308
rect -1402 262 -1334 308
rect -1288 262 -1220 308
rect -1174 262 -1106 308
rect -1060 262 -992 308
rect -946 262 -878 308
rect -832 262 -764 308
rect -718 262 -650 308
rect -604 262 -536 308
rect -490 262 -422 308
rect -376 262 -308 308
rect -262 262 -194 308
rect -148 262 -80 308
rect -34 262 34 308
rect 80 262 148 308
rect 194 262 262 308
rect 308 262 376 308
rect 422 262 490 308
rect 536 262 604 308
rect 650 262 718 308
rect 764 262 832 308
rect 878 262 946 308
rect 992 262 1060 308
rect 1106 262 1174 308
rect 1220 262 1288 308
rect 1334 262 1402 308
rect 1448 262 1516 308
rect 1562 262 1630 308
rect 1676 262 1744 308
rect 1790 262 1858 308
rect 1904 262 1972 308
rect 2018 262 2086 308
rect 2132 262 2200 308
rect 2246 262 2314 308
rect 2360 262 2428 308
rect 2474 262 2542 308
rect 2588 262 2656 308
rect 2702 262 2770 308
rect 2816 262 2884 308
rect 2930 262 2998 308
rect 3044 262 3112 308
rect 3158 262 3226 308
rect 3272 262 3340 308
rect 3386 262 3454 308
rect 3500 262 3568 308
rect 3614 262 3682 308
rect 3728 262 3796 308
rect 3842 262 3910 308
rect 3956 262 4024 308
rect 4070 262 4138 308
rect 4184 262 4252 308
rect 4298 262 4366 308
rect 4412 262 4480 308
rect 4526 262 4594 308
rect 4640 262 4651 308
rect -4651 194 4651 262
rect -4651 148 -4640 194
rect -4594 148 -4526 194
rect -4480 148 -4412 194
rect -4366 148 -4298 194
rect -4252 148 -4184 194
rect -4138 148 -4070 194
rect -4024 148 -3956 194
rect -3910 148 -3842 194
rect -3796 148 -3728 194
rect -3682 148 -3614 194
rect -3568 148 -3500 194
rect -3454 148 -3386 194
rect -3340 148 -3272 194
rect -3226 148 -3158 194
rect -3112 148 -3044 194
rect -2998 148 -2930 194
rect -2884 148 -2816 194
rect -2770 148 -2702 194
rect -2656 148 -2588 194
rect -2542 148 -2474 194
rect -2428 148 -2360 194
rect -2314 148 -2246 194
rect -2200 148 -2132 194
rect -2086 148 -2018 194
rect -1972 148 -1904 194
rect -1858 148 -1790 194
rect -1744 148 -1676 194
rect -1630 148 -1562 194
rect -1516 148 -1448 194
rect -1402 148 -1334 194
rect -1288 148 -1220 194
rect -1174 148 -1106 194
rect -1060 148 -992 194
rect -946 148 -878 194
rect -832 148 -764 194
rect -718 148 -650 194
rect -604 148 -536 194
rect -490 148 -422 194
rect -376 148 -308 194
rect -262 148 -194 194
rect -148 148 -80 194
rect -34 148 34 194
rect 80 148 148 194
rect 194 148 262 194
rect 308 148 376 194
rect 422 148 490 194
rect 536 148 604 194
rect 650 148 718 194
rect 764 148 832 194
rect 878 148 946 194
rect 992 148 1060 194
rect 1106 148 1174 194
rect 1220 148 1288 194
rect 1334 148 1402 194
rect 1448 148 1516 194
rect 1562 148 1630 194
rect 1676 148 1744 194
rect 1790 148 1858 194
rect 1904 148 1972 194
rect 2018 148 2086 194
rect 2132 148 2200 194
rect 2246 148 2314 194
rect 2360 148 2428 194
rect 2474 148 2542 194
rect 2588 148 2656 194
rect 2702 148 2770 194
rect 2816 148 2884 194
rect 2930 148 2998 194
rect 3044 148 3112 194
rect 3158 148 3226 194
rect 3272 148 3340 194
rect 3386 148 3454 194
rect 3500 148 3568 194
rect 3614 148 3682 194
rect 3728 148 3796 194
rect 3842 148 3910 194
rect 3956 148 4024 194
rect 4070 148 4138 194
rect 4184 148 4252 194
rect 4298 148 4366 194
rect 4412 148 4480 194
rect 4526 148 4594 194
rect 4640 148 4651 194
rect -4651 80 4651 148
rect -4651 34 -4640 80
rect -4594 34 -4526 80
rect -4480 34 -4412 80
rect -4366 34 -4298 80
rect -4252 34 -4184 80
rect -4138 34 -4070 80
rect -4024 34 -3956 80
rect -3910 34 -3842 80
rect -3796 34 -3728 80
rect -3682 34 -3614 80
rect -3568 34 -3500 80
rect -3454 34 -3386 80
rect -3340 34 -3272 80
rect -3226 34 -3158 80
rect -3112 34 -3044 80
rect -2998 34 -2930 80
rect -2884 34 -2816 80
rect -2770 34 -2702 80
rect -2656 34 -2588 80
rect -2542 34 -2474 80
rect -2428 34 -2360 80
rect -2314 34 -2246 80
rect -2200 34 -2132 80
rect -2086 34 -2018 80
rect -1972 34 -1904 80
rect -1858 34 -1790 80
rect -1744 34 -1676 80
rect -1630 34 -1562 80
rect -1516 34 -1448 80
rect -1402 34 -1334 80
rect -1288 34 -1220 80
rect -1174 34 -1106 80
rect -1060 34 -992 80
rect -946 34 -878 80
rect -832 34 -764 80
rect -718 34 -650 80
rect -604 34 -536 80
rect -490 34 -422 80
rect -376 34 -308 80
rect -262 34 -194 80
rect -148 34 -80 80
rect -34 34 34 80
rect 80 34 148 80
rect 194 34 262 80
rect 308 34 376 80
rect 422 34 490 80
rect 536 34 604 80
rect 650 34 718 80
rect 764 34 832 80
rect 878 34 946 80
rect 992 34 1060 80
rect 1106 34 1174 80
rect 1220 34 1288 80
rect 1334 34 1402 80
rect 1448 34 1516 80
rect 1562 34 1630 80
rect 1676 34 1744 80
rect 1790 34 1858 80
rect 1904 34 1972 80
rect 2018 34 2086 80
rect 2132 34 2200 80
rect 2246 34 2314 80
rect 2360 34 2428 80
rect 2474 34 2542 80
rect 2588 34 2656 80
rect 2702 34 2770 80
rect 2816 34 2884 80
rect 2930 34 2998 80
rect 3044 34 3112 80
rect 3158 34 3226 80
rect 3272 34 3340 80
rect 3386 34 3454 80
rect 3500 34 3568 80
rect 3614 34 3682 80
rect 3728 34 3796 80
rect 3842 34 3910 80
rect 3956 34 4024 80
rect 4070 34 4138 80
rect 4184 34 4252 80
rect 4298 34 4366 80
rect 4412 34 4480 80
rect 4526 34 4594 80
rect 4640 34 4651 80
rect -4651 -34 4651 34
rect -4651 -80 -4640 -34
rect -4594 -80 -4526 -34
rect -4480 -80 -4412 -34
rect -4366 -80 -4298 -34
rect -4252 -80 -4184 -34
rect -4138 -80 -4070 -34
rect -4024 -80 -3956 -34
rect -3910 -80 -3842 -34
rect -3796 -80 -3728 -34
rect -3682 -80 -3614 -34
rect -3568 -80 -3500 -34
rect -3454 -80 -3386 -34
rect -3340 -80 -3272 -34
rect -3226 -80 -3158 -34
rect -3112 -80 -3044 -34
rect -2998 -80 -2930 -34
rect -2884 -80 -2816 -34
rect -2770 -80 -2702 -34
rect -2656 -80 -2588 -34
rect -2542 -80 -2474 -34
rect -2428 -80 -2360 -34
rect -2314 -80 -2246 -34
rect -2200 -80 -2132 -34
rect -2086 -80 -2018 -34
rect -1972 -80 -1904 -34
rect -1858 -80 -1790 -34
rect -1744 -80 -1676 -34
rect -1630 -80 -1562 -34
rect -1516 -80 -1448 -34
rect -1402 -80 -1334 -34
rect -1288 -80 -1220 -34
rect -1174 -80 -1106 -34
rect -1060 -80 -992 -34
rect -946 -80 -878 -34
rect -832 -80 -764 -34
rect -718 -80 -650 -34
rect -604 -80 -536 -34
rect -490 -80 -422 -34
rect -376 -80 -308 -34
rect -262 -80 -194 -34
rect -148 -80 -80 -34
rect -34 -80 34 -34
rect 80 -80 148 -34
rect 194 -80 262 -34
rect 308 -80 376 -34
rect 422 -80 490 -34
rect 536 -80 604 -34
rect 650 -80 718 -34
rect 764 -80 832 -34
rect 878 -80 946 -34
rect 992 -80 1060 -34
rect 1106 -80 1174 -34
rect 1220 -80 1288 -34
rect 1334 -80 1402 -34
rect 1448 -80 1516 -34
rect 1562 -80 1630 -34
rect 1676 -80 1744 -34
rect 1790 -80 1858 -34
rect 1904 -80 1972 -34
rect 2018 -80 2086 -34
rect 2132 -80 2200 -34
rect 2246 -80 2314 -34
rect 2360 -80 2428 -34
rect 2474 -80 2542 -34
rect 2588 -80 2656 -34
rect 2702 -80 2770 -34
rect 2816 -80 2884 -34
rect 2930 -80 2998 -34
rect 3044 -80 3112 -34
rect 3158 -80 3226 -34
rect 3272 -80 3340 -34
rect 3386 -80 3454 -34
rect 3500 -80 3568 -34
rect 3614 -80 3682 -34
rect 3728 -80 3796 -34
rect 3842 -80 3910 -34
rect 3956 -80 4024 -34
rect 4070 -80 4138 -34
rect 4184 -80 4252 -34
rect 4298 -80 4366 -34
rect 4412 -80 4480 -34
rect 4526 -80 4594 -34
rect 4640 -80 4651 -34
rect -4651 -148 4651 -80
rect -4651 -194 -4640 -148
rect -4594 -194 -4526 -148
rect -4480 -194 -4412 -148
rect -4366 -194 -4298 -148
rect -4252 -194 -4184 -148
rect -4138 -194 -4070 -148
rect -4024 -194 -3956 -148
rect -3910 -194 -3842 -148
rect -3796 -194 -3728 -148
rect -3682 -194 -3614 -148
rect -3568 -194 -3500 -148
rect -3454 -194 -3386 -148
rect -3340 -194 -3272 -148
rect -3226 -194 -3158 -148
rect -3112 -194 -3044 -148
rect -2998 -194 -2930 -148
rect -2884 -194 -2816 -148
rect -2770 -194 -2702 -148
rect -2656 -194 -2588 -148
rect -2542 -194 -2474 -148
rect -2428 -194 -2360 -148
rect -2314 -194 -2246 -148
rect -2200 -194 -2132 -148
rect -2086 -194 -2018 -148
rect -1972 -194 -1904 -148
rect -1858 -194 -1790 -148
rect -1744 -194 -1676 -148
rect -1630 -194 -1562 -148
rect -1516 -194 -1448 -148
rect -1402 -194 -1334 -148
rect -1288 -194 -1220 -148
rect -1174 -194 -1106 -148
rect -1060 -194 -992 -148
rect -946 -194 -878 -148
rect -832 -194 -764 -148
rect -718 -194 -650 -148
rect -604 -194 -536 -148
rect -490 -194 -422 -148
rect -376 -194 -308 -148
rect -262 -194 -194 -148
rect -148 -194 -80 -148
rect -34 -194 34 -148
rect 80 -194 148 -148
rect 194 -194 262 -148
rect 308 -194 376 -148
rect 422 -194 490 -148
rect 536 -194 604 -148
rect 650 -194 718 -148
rect 764 -194 832 -148
rect 878 -194 946 -148
rect 992 -194 1060 -148
rect 1106 -194 1174 -148
rect 1220 -194 1288 -148
rect 1334 -194 1402 -148
rect 1448 -194 1516 -148
rect 1562 -194 1630 -148
rect 1676 -194 1744 -148
rect 1790 -194 1858 -148
rect 1904 -194 1972 -148
rect 2018 -194 2086 -148
rect 2132 -194 2200 -148
rect 2246 -194 2314 -148
rect 2360 -194 2428 -148
rect 2474 -194 2542 -148
rect 2588 -194 2656 -148
rect 2702 -194 2770 -148
rect 2816 -194 2884 -148
rect 2930 -194 2998 -148
rect 3044 -194 3112 -148
rect 3158 -194 3226 -148
rect 3272 -194 3340 -148
rect 3386 -194 3454 -148
rect 3500 -194 3568 -148
rect 3614 -194 3682 -148
rect 3728 -194 3796 -148
rect 3842 -194 3910 -148
rect 3956 -194 4024 -148
rect 4070 -194 4138 -148
rect 4184 -194 4252 -148
rect 4298 -194 4366 -148
rect 4412 -194 4480 -148
rect 4526 -194 4594 -148
rect 4640 -194 4651 -148
rect -4651 -262 4651 -194
rect -4651 -308 -4640 -262
rect -4594 -308 -4526 -262
rect -4480 -308 -4412 -262
rect -4366 -308 -4298 -262
rect -4252 -308 -4184 -262
rect -4138 -308 -4070 -262
rect -4024 -308 -3956 -262
rect -3910 -308 -3842 -262
rect -3796 -308 -3728 -262
rect -3682 -308 -3614 -262
rect -3568 -308 -3500 -262
rect -3454 -308 -3386 -262
rect -3340 -308 -3272 -262
rect -3226 -308 -3158 -262
rect -3112 -308 -3044 -262
rect -2998 -308 -2930 -262
rect -2884 -308 -2816 -262
rect -2770 -308 -2702 -262
rect -2656 -308 -2588 -262
rect -2542 -308 -2474 -262
rect -2428 -308 -2360 -262
rect -2314 -308 -2246 -262
rect -2200 -308 -2132 -262
rect -2086 -308 -2018 -262
rect -1972 -308 -1904 -262
rect -1858 -308 -1790 -262
rect -1744 -308 -1676 -262
rect -1630 -308 -1562 -262
rect -1516 -308 -1448 -262
rect -1402 -308 -1334 -262
rect -1288 -308 -1220 -262
rect -1174 -308 -1106 -262
rect -1060 -308 -992 -262
rect -946 -308 -878 -262
rect -832 -308 -764 -262
rect -718 -308 -650 -262
rect -604 -308 -536 -262
rect -490 -308 -422 -262
rect -376 -308 -308 -262
rect -262 -308 -194 -262
rect -148 -308 -80 -262
rect -34 -308 34 -262
rect 80 -308 148 -262
rect 194 -308 262 -262
rect 308 -308 376 -262
rect 422 -308 490 -262
rect 536 -308 604 -262
rect 650 -308 718 -262
rect 764 -308 832 -262
rect 878 -308 946 -262
rect 992 -308 1060 -262
rect 1106 -308 1174 -262
rect 1220 -308 1288 -262
rect 1334 -308 1402 -262
rect 1448 -308 1516 -262
rect 1562 -308 1630 -262
rect 1676 -308 1744 -262
rect 1790 -308 1858 -262
rect 1904 -308 1972 -262
rect 2018 -308 2086 -262
rect 2132 -308 2200 -262
rect 2246 -308 2314 -262
rect 2360 -308 2428 -262
rect 2474 -308 2542 -262
rect 2588 -308 2656 -262
rect 2702 -308 2770 -262
rect 2816 -308 2884 -262
rect 2930 -308 2998 -262
rect 3044 -308 3112 -262
rect 3158 -308 3226 -262
rect 3272 -308 3340 -262
rect 3386 -308 3454 -262
rect 3500 -308 3568 -262
rect 3614 -308 3682 -262
rect 3728 -308 3796 -262
rect 3842 -308 3910 -262
rect 3956 -308 4024 -262
rect 4070 -308 4138 -262
rect 4184 -308 4252 -262
rect 4298 -308 4366 -262
rect 4412 -308 4480 -262
rect 4526 -308 4594 -262
rect 4640 -308 4651 -262
rect -4651 -376 4651 -308
rect -4651 -422 -4640 -376
rect -4594 -422 -4526 -376
rect -4480 -422 -4412 -376
rect -4366 -422 -4298 -376
rect -4252 -422 -4184 -376
rect -4138 -422 -4070 -376
rect -4024 -422 -3956 -376
rect -3910 -422 -3842 -376
rect -3796 -422 -3728 -376
rect -3682 -422 -3614 -376
rect -3568 -422 -3500 -376
rect -3454 -422 -3386 -376
rect -3340 -422 -3272 -376
rect -3226 -422 -3158 -376
rect -3112 -422 -3044 -376
rect -2998 -422 -2930 -376
rect -2884 -422 -2816 -376
rect -2770 -422 -2702 -376
rect -2656 -422 -2588 -376
rect -2542 -422 -2474 -376
rect -2428 -422 -2360 -376
rect -2314 -422 -2246 -376
rect -2200 -422 -2132 -376
rect -2086 -422 -2018 -376
rect -1972 -422 -1904 -376
rect -1858 -422 -1790 -376
rect -1744 -422 -1676 -376
rect -1630 -422 -1562 -376
rect -1516 -422 -1448 -376
rect -1402 -422 -1334 -376
rect -1288 -422 -1220 -376
rect -1174 -422 -1106 -376
rect -1060 -422 -992 -376
rect -946 -422 -878 -376
rect -832 -422 -764 -376
rect -718 -422 -650 -376
rect -604 -422 -536 -376
rect -490 -422 -422 -376
rect -376 -422 -308 -376
rect -262 -422 -194 -376
rect -148 -422 -80 -376
rect -34 -422 34 -376
rect 80 -422 148 -376
rect 194 -422 262 -376
rect 308 -422 376 -376
rect 422 -422 490 -376
rect 536 -422 604 -376
rect 650 -422 718 -376
rect 764 -422 832 -376
rect 878 -422 946 -376
rect 992 -422 1060 -376
rect 1106 -422 1174 -376
rect 1220 -422 1288 -376
rect 1334 -422 1402 -376
rect 1448 -422 1516 -376
rect 1562 -422 1630 -376
rect 1676 -422 1744 -376
rect 1790 -422 1858 -376
rect 1904 -422 1972 -376
rect 2018 -422 2086 -376
rect 2132 -422 2200 -376
rect 2246 -422 2314 -376
rect 2360 -422 2428 -376
rect 2474 -422 2542 -376
rect 2588 -422 2656 -376
rect 2702 -422 2770 -376
rect 2816 -422 2884 -376
rect 2930 -422 2998 -376
rect 3044 -422 3112 -376
rect 3158 -422 3226 -376
rect 3272 -422 3340 -376
rect 3386 -422 3454 -376
rect 3500 -422 3568 -376
rect 3614 -422 3682 -376
rect 3728 -422 3796 -376
rect 3842 -422 3910 -376
rect 3956 -422 4024 -376
rect 4070 -422 4138 -376
rect 4184 -422 4252 -376
rect 4298 -422 4366 -376
rect 4412 -422 4480 -376
rect 4526 -422 4594 -376
rect 4640 -422 4651 -376
rect -4651 -490 4651 -422
rect -4651 -536 -4640 -490
rect -4594 -536 -4526 -490
rect -4480 -536 -4412 -490
rect -4366 -536 -4298 -490
rect -4252 -536 -4184 -490
rect -4138 -536 -4070 -490
rect -4024 -536 -3956 -490
rect -3910 -536 -3842 -490
rect -3796 -536 -3728 -490
rect -3682 -536 -3614 -490
rect -3568 -536 -3500 -490
rect -3454 -536 -3386 -490
rect -3340 -536 -3272 -490
rect -3226 -536 -3158 -490
rect -3112 -536 -3044 -490
rect -2998 -536 -2930 -490
rect -2884 -536 -2816 -490
rect -2770 -536 -2702 -490
rect -2656 -536 -2588 -490
rect -2542 -536 -2474 -490
rect -2428 -536 -2360 -490
rect -2314 -536 -2246 -490
rect -2200 -536 -2132 -490
rect -2086 -536 -2018 -490
rect -1972 -536 -1904 -490
rect -1858 -536 -1790 -490
rect -1744 -536 -1676 -490
rect -1630 -536 -1562 -490
rect -1516 -536 -1448 -490
rect -1402 -536 -1334 -490
rect -1288 -536 -1220 -490
rect -1174 -536 -1106 -490
rect -1060 -536 -992 -490
rect -946 -536 -878 -490
rect -832 -536 -764 -490
rect -718 -536 -650 -490
rect -604 -536 -536 -490
rect -490 -536 -422 -490
rect -376 -536 -308 -490
rect -262 -536 -194 -490
rect -148 -536 -80 -490
rect -34 -536 34 -490
rect 80 -536 148 -490
rect 194 -536 262 -490
rect 308 -536 376 -490
rect 422 -536 490 -490
rect 536 -536 604 -490
rect 650 -536 718 -490
rect 764 -536 832 -490
rect 878 -536 946 -490
rect 992 -536 1060 -490
rect 1106 -536 1174 -490
rect 1220 -536 1288 -490
rect 1334 -536 1402 -490
rect 1448 -536 1516 -490
rect 1562 -536 1630 -490
rect 1676 -536 1744 -490
rect 1790 -536 1858 -490
rect 1904 -536 1972 -490
rect 2018 -536 2086 -490
rect 2132 -536 2200 -490
rect 2246 -536 2314 -490
rect 2360 -536 2428 -490
rect 2474 -536 2542 -490
rect 2588 -536 2656 -490
rect 2702 -536 2770 -490
rect 2816 -536 2884 -490
rect 2930 -536 2998 -490
rect 3044 -536 3112 -490
rect 3158 -536 3226 -490
rect 3272 -536 3340 -490
rect 3386 -536 3454 -490
rect 3500 -536 3568 -490
rect 3614 -536 3682 -490
rect 3728 -536 3796 -490
rect 3842 -536 3910 -490
rect 3956 -536 4024 -490
rect 4070 -536 4138 -490
rect 4184 -536 4252 -490
rect 4298 -536 4366 -490
rect 4412 -536 4480 -490
rect 4526 -536 4594 -490
rect 4640 -536 4651 -490
rect -4651 -604 4651 -536
rect -4651 -650 -4640 -604
rect -4594 -650 -4526 -604
rect -4480 -650 -4412 -604
rect -4366 -650 -4298 -604
rect -4252 -650 -4184 -604
rect -4138 -650 -4070 -604
rect -4024 -650 -3956 -604
rect -3910 -650 -3842 -604
rect -3796 -650 -3728 -604
rect -3682 -650 -3614 -604
rect -3568 -650 -3500 -604
rect -3454 -650 -3386 -604
rect -3340 -650 -3272 -604
rect -3226 -650 -3158 -604
rect -3112 -650 -3044 -604
rect -2998 -650 -2930 -604
rect -2884 -650 -2816 -604
rect -2770 -650 -2702 -604
rect -2656 -650 -2588 -604
rect -2542 -650 -2474 -604
rect -2428 -650 -2360 -604
rect -2314 -650 -2246 -604
rect -2200 -650 -2132 -604
rect -2086 -650 -2018 -604
rect -1972 -650 -1904 -604
rect -1858 -650 -1790 -604
rect -1744 -650 -1676 -604
rect -1630 -650 -1562 -604
rect -1516 -650 -1448 -604
rect -1402 -650 -1334 -604
rect -1288 -650 -1220 -604
rect -1174 -650 -1106 -604
rect -1060 -650 -992 -604
rect -946 -650 -878 -604
rect -832 -650 -764 -604
rect -718 -650 -650 -604
rect -604 -650 -536 -604
rect -490 -650 -422 -604
rect -376 -650 -308 -604
rect -262 -650 -194 -604
rect -148 -650 -80 -604
rect -34 -650 34 -604
rect 80 -650 148 -604
rect 194 -650 262 -604
rect 308 -650 376 -604
rect 422 -650 490 -604
rect 536 -650 604 -604
rect 650 -650 718 -604
rect 764 -650 832 -604
rect 878 -650 946 -604
rect 992 -650 1060 -604
rect 1106 -650 1174 -604
rect 1220 -650 1288 -604
rect 1334 -650 1402 -604
rect 1448 -650 1516 -604
rect 1562 -650 1630 -604
rect 1676 -650 1744 -604
rect 1790 -650 1858 -604
rect 1904 -650 1972 -604
rect 2018 -650 2086 -604
rect 2132 -650 2200 -604
rect 2246 -650 2314 -604
rect 2360 -650 2428 -604
rect 2474 -650 2542 -604
rect 2588 -650 2656 -604
rect 2702 -650 2770 -604
rect 2816 -650 2884 -604
rect 2930 -650 2998 -604
rect 3044 -650 3112 -604
rect 3158 -650 3226 -604
rect 3272 -650 3340 -604
rect 3386 -650 3454 -604
rect 3500 -650 3568 -604
rect 3614 -650 3682 -604
rect 3728 -650 3796 -604
rect 3842 -650 3910 -604
rect 3956 -650 4024 -604
rect 4070 -650 4138 -604
rect 4184 -650 4252 -604
rect 4298 -650 4366 -604
rect 4412 -650 4480 -604
rect 4526 -650 4594 -604
rect 4640 -650 4651 -604
rect -4651 -718 4651 -650
rect -4651 -764 -4640 -718
rect -4594 -764 -4526 -718
rect -4480 -764 -4412 -718
rect -4366 -764 -4298 -718
rect -4252 -764 -4184 -718
rect -4138 -764 -4070 -718
rect -4024 -764 -3956 -718
rect -3910 -764 -3842 -718
rect -3796 -764 -3728 -718
rect -3682 -764 -3614 -718
rect -3568 -764 -3500 -718
rect -3454 -764 -3386 -718
rect -3340 -764 -3272 -718
rect -3226 -764 -3158 -718
rect -3112 -764 -3044 -718
rect -2998 -764 -2930 -718
rect -2884 -764 -2816 -718
rect -2770 -764 -2702 -718
rect -2656 -764 -2588 -718
rect -2542 -764 -2474 -718
rect -2428 -764 -2360 -718
rect -2314 -764 -2246 -718
rect -2200 -764 -2132 -718
rect -2086 -764 -2018 -718
rect -1972 -764 -1904 -718
rect -1858 -764 -1790 -718
rect -1744 -764 -1676 -718
rect -1630 -764 -1562 -718
rect -1516 -764 -1448 -718
rect -1402 -764 -1334 -718
rect -1288 -764 -1220 -718
rect -1174 -764 -1106 -718
rect -1060 -764 -992 -718
rect -946 -764 -878 -718
rect -832 -764 -764 -718
rect -718 -764 -650 -718
rect -604 -764 -536 -718
rect -490 -764 -422 -718
rect -376 -764 -308 -718
rect -262 -764 -194 -718
rect -148 -764 -80 -718
rect -34 -764 34 -718
rect 80 -764 148 -718
rect 194 -764 262 -718
rect 308 -764 376 -718
rect 422 -764 490 -718
rect 536 -764 604 -718
rect 650 -764 718 -718
rect 764 -764 832 -718
rect 878 -764 946 -718
rect 992 -764 1060 -718
rect 1106 -764 1174 -718
rect 1220 -764 1288 -718
rect 1334 -764 1402 -718
rect 1448 -764 1516 -718
rect 1562 -764 1630 -718
rect 1676 -764 1744 -718
rect 1790 -764 1858 -718
rect 1904 -764 1972 -718
rect 2018 -764 2086 -718
rect 2132 -764 2200 -718
rect 2246 -764 2314 -718
rect 2360 -764 2428 -718
rect 2474 -764 2542 -718
rect 2588 -764 2656 -718
rect 2702 -764 2770 -718
rect 2816 -764 2884 -718
rect 2930 -764 2998 -718
rect 3044 -764 3112 -718
rect 3158 -764 3226 -718
rect 3272 -764 3340 -718
rect 3386 -764 3454 -718
rect 3500 -764 3568 -718
rect 3614 -764 3682 -718
rect 3728 -764 3796 -718
rect 3842 -764 3910 -718
rect 3956 -764 4024 -718
rect 4070 -764 4138 -718
rect 4184 -764 4252 -718
rect 4298 -764 4366 -718
rect 4412 -764 4480 -718
rect 4526 -764 4594 -718
rect 4640 -764 4651 -718
rect -4651 -775 4651 -764
<< end >>
