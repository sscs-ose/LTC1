magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2128 -3491 2128 3491
<< nwell >>
rect -128 -1491 128 1491
<< nsubdiff >>
rect -45 1386 45 1408
rect -45 -1386 -23 1386
rect 23 -1386 45 1386
rect -45 -1408 45 -1386
<< nsubdiffcont >>
rect -23 -1386 23 1386
<< metal1 >>
rect -34 1386 34 1397
rect -34 -1386 -23 1386
rect 23 -1386 34 1386
rect -34 -1397 34 -1386
<< end >>
