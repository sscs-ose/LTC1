magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2228 -8078 2228 8078
<< nwell >>
rect -228 -6078 228 6078
<< nsubdiff >>
rect -145 5945 145 5995
rect -145 -5945 -117 5945
rect 117 -5945 145 5945
rect -145 -5995 145 -5945
<< nsubdiffcont >>
rect -117 -5945 117 5945
<< metal1 >>
rect -134 5945 134 5984
rect -134 -5945 -117 5945
rect 117 -5945 134 5945
rect -134 -5984 134 -5945
<< end >>
