magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2045 -2515 2045 2515
<< psubdiff >>
rect -45 493 45 515
rect -45 -493 -23 493
rect 23 -493 45 493
rect -45 -515 45 -493
<< psubdiffcont >>
rect -23 -493 23 493
<< metal1 >>
rect -34 493 34 504
rect -34 -493 -23 493
rect 23 -493 34 493
rect -34 -504 34 -493
<< end >>
