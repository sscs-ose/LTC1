magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1349 -6068 1349 6068
<< metal3 >>
rect -349 5063 349 5068
rect -349 5035 -344 5063
rect -316 5035 -278 5063
rect -250 5035 -212 5063
rect -184 5035 -146 5063
rect -118 5035 -80 5063
rect -52 5035 -14 5063
rect 14 5035 52 5063
rect 80 5035 118 5063
rect 146 5035 184 5063
rect 212 5035 250 5063
rect 278 5035 316 5063
rect 344 5035 349 5063
rect -349 4997 349 5035
rect -349 4969 -344 4997
rect -316 4969 -278 4997
rect -250 4969 -212 4997
rect -184 4969 -146 4997
rect -118 4969 -80 4997
rect -52 4969 -14 4997
rect 14 4969 52 4997
rect 80 4969 118 4997
rect 146 4969 184 4997
rect 212 4969 250 4997
rect 278 4969 316 4997
rect 344 4969 349 4997
rect -349 4931 349 4969
rect -349 4903 -344 4931
rect -316 4903 -278 4931
rect -250 4903 -212 4931
rect -184 4903 -146 4931
rect -118 4903 -80 4931
rect -52 4903 -14 4931
rect 14 4903 52 4931
rect 80 4903 118 4931
rect 146 4903 184 4931
rect 212 4903 250 4931
rect 278 4903 316 4931
rect 344 4903 349 4931
rect -349 4865 349 4903
rect -349 4837 -344 4865
rect -316 4837 -278 4865
rect -250 4837 -212 4865
rect -184 4837 -146 4865
rect -118 4837 -80 4865
rect -52 4837 -14 4865
rect 14 4837 52 4865
rect 80 4837 118 4865
rect 146 4837 184 4865
rect 212 4837 250 4865
rect 278 4837 316 4865
rect 344 4837 349 4865
rect -349 4799 349 4837
rect -349 4771 -344 4799
rect -316 4771 -278 4799
rect -250 4771 -212 4799
rect -184 4771 -146 4799
rect -118 4771 -80 4799
rect -52 4771 -14 4799
rect 14 4771 52 4799
rect 80 4771 118 4799
rect 146 4771 184 4799
rect 212 4771 250 4799
rect 278 4771 316 4799
rect 344 4771 349 4799
rect -349 4733 349 4771
rect -349 4705 -344 4733
rect -316 4705 -278 4733
rect -250 4705 -212 4733
rect -184 4705 -146 4733
rect -118 4705 -80 4733
rect -52 4705 -14 4733
rect 14 4705 52 4733
rect 80 4705 118 4733
rect 146 4705 184 4733
rect 212 4705 250 4733
rect 278 4705 316 4733
rect 344 4705 349 4733
rect -349 4667 349 4705
rect -349 4639 -344 4667
rect -316 4639 -278 4667
rect -250 4639 -212 4667
rect -184 4639 -146 4667
rect -118 4639 -80 4667
rect -52 4639 -14 4667
rect 14 4639 52 4667
rect 80 4639 118 4667
rect 146 4639 184 4667
rect 212 4639 250 4667
rect 278 4639 316 4667
rect 344 4639 349 4667
rect -349 4601 349 4639
rect -349 4573 -344 4601
rect -316 4573 -278 4601
rect -250 4573 -212 4601
rect -184 4573 -146 4601
rect -118 4573 -80 4601
rect -52 4573 -14 4601
rect 14 4573 52 4601
rect 80 4573 118 4601
rect 146 4573 184 4601
rect 212 4573 250 4601
rect 278 4573 316 4601
rect 344 4573 349 4601
rect -349 4535 349 4573
rect -349 4507 -344 4535
rect -316 4507 -278 4535
rect -250 4507 -212 4535
rect -184 4507 -146 4535
rect -118 4507 -80 4535
rect -52 4507 -14 4535
rect 14 4507 52 4535
rect 80 4507 118 4535
rect 146 4507 184 4535
rect 212 4507 250 4535
rect 278 4507 316 4535
rect 344 4507 349 4535
rect -349 4469 349 4507
rect -349 4441 -344 4469
rect -316 4441 -278 4469
rect -250 4441 -212 4469
rect -184 4441 -146 4469
rect -118 4441 -80 4469
rect -52 4441 -14 4469
rect 14 4441 52 4469
rect 80 4441 118 4469
rect 146 4441 184 4469
rect 212 4441 250 4469
rect 278 4441 316 4469
rect 344 4441 349 4469
rect -349 4403 349 4441
rect -349 4375 -344 4403
rect -316 4375 -278 4403
rect -250 4375 -212 4403
rect -184 4375 -146 4403
rect -118 4375 -80 4403
rect -52 4375 -14 4403
rect 14 4375 52 4403
rect 80 4375 118 4403
rect 146 4375 184 4403
rect 212 4375 250 4403
rect 278 4375 316 4403
rect 344 4375 349 4403
rect -349 4337 349 4375
rect -349 4309 -344 4337
rect -316 4309 -278 4337
rect -250 4309 -212 4337
rect -184 4309 -146 4337
rect -118 4309 -80 4337
rect -52 4309 -14 4337
rect 14 4309 52 4337
rect 80 4309 118 4337
rect 146 4309 184 4337
rect 212 4309 250 4337
rect 278 4309 316 4337
rect 344 4309 349 4337
rect -349 4271 349 4309
rect -349 4243 -344 4271
rect -316 4243 -278 4271
rect -250 4243 -212 4271
rect -184 4243 -146 4271
rect -118 4243 -80 4271
rect -52 4243 -14 4271
rect 14 4243 52 4271
rect 80 4243 118 4271
rect 146 4243 184 4271
rect 212 4243 250 4271
rect 278 4243 316 4271
rect 344 4243 349 4271
rect -349 4205 349 4243
rect -349 4177 -344 4205
rect -316 4177 -278 4205
rect -250 4177 -212 4205
rect -184 4177 -146 4205
rect -118 4177 -80 4205
rect -52 4177 -14 4205
rect 14 4177 52 4205
rect 80 4177 118 4205
rect 146 4177 184 4205
rect 212 4177 250 4205
rect 278 4177 316 4205
rect 344 4177 349 4205
rect -349 4139 349 4177
rect -349 4111 -344 4139
rect -316 4111 -278 4139
rect -250 4111 -212 4139
rect -184 4111 -146 4139
rect -118 4111 -80 4139
rect -52 4111 -14 4139
rect 14 4111 52 4139
rect 80 4111 118 4139
rect 146 4111 184 4139
rect 212 4111 250 4139
rect 278 4111 316 4139
rect 344 4111 349 4139
rect -349 4073 349 4111
rect -349 4045 -344 4073
rect -316 4045 -278 4073
rect -250 4045 -212 4073
rect -184 4045 -146 4073
rect -118 4045 -80 4073
rect -52 4045 -14 4073
rect 14 4045 52 4073
rect 80 4045 118 4073
rect 146 4045 184 4073
rect 212 4045 250 4073
rect 278 4045 316 4073
rect 344 4045 349 4073
rect -349 4007 349 4045
rect -349 3979 -344 4007
rect -316 3979 -278 4007
rect -250 3979 -212 4007
rect -184 3979 -146 4007
rect -118 3979 -80 4007
rect -52 3979 -14 4007
rect 14 3979 52 4007
rect 80 3979 118 4007
rect 146 3979 184 4007
rect 212 3979 250 4007
rect 278 3979 316 4007
rect 344 3979 349 4007
rect -349 3941 349 3979
rect -349 3913 -344 3941
rect -316 3913 -278 3941
rect -250 3913 -212 3941
rect -184 3913 -146 3941
rect -118 3913 -80 3941
rect -52 3913 -14 3941
rect 14 3913 52 3941
rect 80 3913 118 3941
rect 146 3913 184 3941
rect 212 3913 250 3941
rect 278 3913 316 3941
rect 344 3913 349 3941
rect -349 3875 349 3913
rect -349 3847 -344 3875
rect -316 3847 -278 3875
rect -250 3847 -212 3875
rect -184 3847 -146 3875
rect -118 3847 -80 3875
rect -52 3847 -14 3875
rect 14 3847 52 3875
rect 80 3847 118 3875
rect 146 3847 184 3875
rect 212 3847 250 3875
rect 278 3847 316 3875
rect 344 3847 349 3875
rect -349 3809 349 3847
rect -349 3781 -344 3809
rect -316 3781 -278 3809
rect -250 3781 -212 3809
rect -184 3781 -146 3809
rect -118 3781 -80 3809
rect -52 3781 -14 3809
rect 14 3781 52 3809
rect 80 3781 118 3809
rect 146 3781 184 3809
rect 212 3781 250 3809
rect 278 3781 316 3809
rect 344 3781 349 3809
rect -349 3743 349 3781
rect -349 3715 -344 3743
rect -316 3715 -278 3743
rect -250 3715 -212 3743
rect -184 3715 -146 3743
rect -118 3715 -80 3743
rect -52 3715 -14 3743
rect 14 3715 52 3743
rect 80 3715 118 3743
rect 146 3715 184 3743
rect 212 3715 250 3743
rect 278 3715 316 3743
rect 344 3715 349 3743
rect -349 3677 349 3715
rect -349 3649 -344 3677
rect -316 3649 -278 3677
rect -250 3649 -212 3677
rect -184 3649 -146 3677
rect -118 3649 -80 3677
rect -52 3649 -14 3677
rect 14 3649 52 3677
rect 80 3649 118 3677
rect 146 3649 184 3677
rect 212 3649 250 3677
rect 278 3649 316 3677
rect 344 3649 349 3677
rect -349 3611 349 3649
rect -349 3583 -344 3611
rect -316 3583 -278 3611
rect -250 3583 -212 3611
rect -184 3583 -146 3611
rect -118 3583 -80 3611
rect -52 3583 -14 3611
rect 14 3583 52 3611
rect 80 3583 118 3611
rect 146 3583 184 3611
rect 212 3583 250 3611
rect 278 3583 316 3611
rect 344 3583 349 3611
rect -349 3545 349 3583
rect -349 3517 -344 3545
rect -316 3517 -278 3545
rect -250 3517 -212 3545
rect -184 3517 -146 3545
rect -118 3517 -80 3545
rect -52 3517 -14 3545
rect 14 3517 52 3545
rect 80 3517 118 3545
rect 146 3517 184 3545
rect 212 3517 250 3545
rect 278 3517 316 3545
rect 344 3517 349 3545
rect -349 3479 349 3517
rect -349 3451 -344 3479
rect -316 3451 -278 3479
rect -250 3451 -212 3479
rect -184 3451 -146 3479
rect -118 3451 -80 3479
rect -52 3451 -14 3479
rect 14 3451 52 3479
rect 80 3451 118 3479
rect 146 3451 184 3479
rect 212 3451 250 3479
rect 278 3451 316 3479
rect 344 3451 349 3479
rect -349 3413 349 3451
rect -349 3385 -344 3413
rect -316 3385 -278 3413
rect -250 3385 -212 3413
rect -184 3385 -146 3413
rect -118 3385 -80 3413
rect -52 3385 -14 3413
rect 14 3385 52 3413
rect 80 3385 118 3413
rect 146 3385 184 3413
rect 212 3385 250 3413
rect 278 3385 316 3413
rect 344 3385 349 3413
rect -349 3347 349 3385
rect -349 3319 -344 3347
rect -316 3319 -278 3347
rect -250 3319 -212 3347
rect -184 3319 -146 3347
rect -118 3319 -80 3347
rect -52 3319 -14 3347
rect 14 3319 52 3347
rect 80 3319 118 3347
rect 146 3319 184 3347
rect 212 3319 250 3347
rect 278 3319 316 3347
rect 344 3319 349 3347
rect -349 3281 349 3319
rect -349 3253 -344 3281
rect -316 3253 -278 3281
rect -250 3253 -212 3281
rect -184 3253 -146 3281
rect -118 3253 -80 3281
rect -52 3253 -14 3281
rect 14 3253 52 3281
rect 80 3253 118 3281
rect 146 3253 184 3281
rect 212 3253 250 3281
rect 278 3253 316 3281
rect 344 3253 349 3281
rect -349 3215 349 3253
rect -349 3187 -344 3215
rect -316 3187 -278 3215
rect -250 3187 -212 3215
rect -184 3187 -146 3215
rect -118 3187 -80 3215
rect -52 3187 -14 3215
rect 14 3187 52 3215
rect 80 3187 118 3215
rect 146 3187 184 3215
rect 212 3187 250 3215
rect 278 3187 316 3215
rect 344 3187 349 3215
rect -349 3149 349 3187
rect -349 3121 -344 3149
rect -316 3121 -278 3149
rect -250 3121 -212 3149
rect -184 3121 -146 3149
rect -118 3121 -80 3149
rect -52 3121 -14 3149
rect 14 3121 52 3149
rect 80 3121 118 3149
rect 146 3121 184 3149
rect 212 3121 250 3149
rect 278 3121 316 3149
rect 344 3121 349 3149
rect -349 3083 349 3121
rect -349 3055 -344 3083
rect -316 3055 -278 3083
rect -250 3055 -212 3083
rect -184 3055 -146 3083
rect -118 3055 -80 3083
rect -52 3055 -14 3083
rect 14 3055 52 3083
rect 80 3055 118 3083
rect 146 3055 184 3083
rect 212 3055 250 3083
rect 278 3055 316 3083
rect 344 3055 349 3083
rect -349 3017 349 3055
rect -349 2989 -344 3017
rect -316 2989 -278 3017
rect -250 2989 -212 3017
rect -184 2989 -146 3017
rect -118 2989 -80 3017
rect -52 2989 -14 3017
rect 14 2989 52 3017
rect 80 2989 118 3017
rect 146 2989 184 3017
rect 212 2989 250 3017
rect 278 2989 316 3017
rect 344 2989 349 3017
rect -349 2951 349 2989
rect -349 2923 -344 2951
rect -316 2923 -278 2951
rect -250 2923 -212 2951
rect -184 2923 -146 2951
rect -118 2923 -80 2951
rect -52 2923 -14 2951
rect 14 2923 52 2951
rect 80 2923 118 2951
rect 146 2923 184 2951
rect 212 2923 250 2951
rect 278 2923 316 2951
rect 344 2923 349 2951
rect -349 2885 349 2923
rect -349 2857 -344 2885
rect -316 2857 -278 2885
rect -250 2857 -212 2885
rect -184 2857 -146 2885
rect -118 2857 -80 2885
rect -52 2857 -14 2885
rect 14 2857 52 2885
rect 80 2857 118 2885
rect 146 2857 184 2885
rect 212 2857 250 2885
rect 278 2857 316 2885
rect 344 2857 349 2885
rect -349 2819 349 2857
rect -349 2791 -344 2819
rect -316 2791 -278 2819
rect -250 2791 -212 2819
rect -184 2791 -146 2819
rect -118 2791 -80 2819
rect -52 2791 -14 2819
rect 14 2791 52 2819
rect 80 2791 118 2819
rect 146 2791 184 2819
rect 212 2791 250 2819
rect 278 2791 316 2819
rect 344 2791 349 2819
rect -349 2753 349 2791
rect -349 2725 -344 2753
rect -316 2725 -278 2753
rect -250 2725 -212 2753
rect -184 2725 -146 2753
rect -118 2725 -80 2753
rect -52 2725 -14 2753
rect 14 2725 52 2753
rect 80 2725 118 2753
rect 146 2725 184 2753
rect 212 2725 250 2753
rect 278 2725 316 2753
rect 344 2725 349 2753
rect -349 2687 349 2725
rect -349 2659 -344 2687
rect -316 2659 -278 2687
rect -250 2659 -212 2687
rect -184 2659 -146 2687
rect -118 2659 -80 2687
rect -52 2659 -14 2687
rect 14 2659 52 2687
rect 80 2659 118 2687
rect 146 2659 184 2687
rect 212 2659 250 2687
rect 278 2659 316 2687
rect 344 2659 349 2687
rect -349 2621 349 2659
rect -349 2593 -344 2621
rect -316 2593 -278 2621
rect -250 2593 -212 2621
rect -184 2593 -146 2621
rect -118 2593 -80 2621
rect -52 2593 -14 2621
rect 14 2593 52 2621
rect 80 2593 118 2621
rect 146 2593 184 2621
rect 212 2593 250 2621
rect 278 2593 316 2621
rect 344 2593 349 2621
rect -349 2555 349 2593
rect -349 2527 -344 2555
rect -316 2527 -278 2555
rect -250 2527 -212 2555
rect -184 2527 -146 2555
rect -118 2527 -80 2555
rect -52 2527 -14 2555
rect 14 2527 52 2555
rect 80 2527 118 2555
rect 146 2527 184 2555
rect 212 2527 250 2555
rect 278 2527 316 2555
rect 344 2527 349 2555
rect -349 2489 349 2527
rect -349 2461 -344 2489
rect -316 2461 -278 2489
rect -250 2461 -212 2489
rect -184 2461 -146 2489
rect -118 2461 -80 2489
rect -52 2461 -14 2489
rect 14 2461 52 2489
rect 80 2461 118 2489
rect 146 2461 184 2489
rect 212 2461 250 2489
rect 278 2461 316 2489
rect 344 2461 349 2489
rect -349 2423 349 2461
rect -349 2395 -344 2423
rect -316 2395 -278 2423
rect -250 2395 -212 2423
rect -184 2395 -146 2423
rect -118 2395 -80 2423
rect -52 2395 -14 2423
rect 14 2395 52 2423
rect 80 2395 118 2423
rect 146 2395 184 2423
rect 212 2395 250 2423
rect 278 2395 316 2423
rect 344 2395 349 2423
rect -349 2357 349 2395
rect -349 2329 -344 2357
rect -316 2329 -278 2357
rect -250 2329 -212 2357
rect -184 2329 -146 2357
rect -118 2329 -80 2357
rect -52 2329 -14 2357
rect 14 2329 52 2357
rect 80 2329 118 2357
rect 146 2329 184 2357
rect 212 2329 250 2357
rect 278 2329 316 2357
rect 344 2329 349 2357
rect -349 2291 349 2329
rect -349 2263 -344 2291
rect -316 2263 -278 2291
rect -250 2263 -212 2291
rect -184 2263 -146 2291
rect -118 2263 -80 2291
rect -52 2263 -14 2291
rect 14 2263 52 2291
rect 80 2263 118 2291
rect 146 2263 184 2291
rect 212 2263 250 2291
rect 278 2263 316 2291
rect 344 2263 349 2291
rect -349 2225 349 2263
rect -349 2197 -344 2225
rect -316 2197 -278 2225
rect -250 2197 -212 2225
rect -184 2197 -146 2225
rect -118 2197 -80 2225
rect -52 2197 -14 2225
rect 14 2197 52 2225
rect 80 2197 118 2225
rect 146 2197 184 2225
rect 212 2197 250 2225
rect 278 2197 316 2225
rect 344 2197 349 2225
rect -349 2159 349 2197
rect -349 2131 -344 2159
rect -316 2131 -278 2159
rect -250 2131 -212 2159
rect -184 2131 -146 2159
rect -118 2131 -80 2159
rect -52 2131 -14 2159
rect 14 2131 52 2159
rect 80 2131 118 2159
rect 146 2131 184 2159
rect 212 2131 250 2159
rect 278 2131 316 2159
rect 344 2131 349 2159
rect -349 2093 349 2131
rect -349 2065 -344 2093
rect -316 2065 -278 2093
rect -250 2065 -212 2093
rect -184 2065 -146 2093
rect -118 2065 -80 2093
rect -52 2065 -14 2093
rect 14 2065 52 2093
rect 80 2065 118 2093
rect 146 2065 184 2093
rect 212 2065 250 2093
rect 278 2065 316 2093
rect 344 2065 349 2093
rect -349 2027 349 2065
rect -349 1999 -344 2027
rect -316 1999 -278 2027
rect -250 1999 -212 2027
rect -184 1999 -146 2027
rect -118 1999 -80 2027
rect -52 1999 -14 2027
rect 14 1999 52 2027
rect 80 1999 118 2027
rect 146 1999 184 2027
rect 212 1999 250 2027
rect 278 1999 316 2027
rect 344 1999 349 2027
rect -349 1961 349 1999
rect -349 1933 -344 1961
rect -316 1933 -278 1961
rect -250 1933 -212 1961
rect -184 1933 -146 1961
rect -118 1933 -80 1961
rect -52 1933 -14 1961
rect 14 1933 52 1961
rect 80 1933 118 1961
rect 146 1933 184 1961
rect 212 1933 250 1961
rect 278 1933 316 1961
rect 344 1933 349 1961
rect -349 1895 349 1933
rect -349 1867 -344 1895
rect -316 1867 -278 1895
rect -250 1867 -212 1895
rect -184 1867 -146 1895
rect -118 1867 -80 1895
rect -52 1867 -14 1895
rect 14 1867 52 1895
rect 80 1867 118 1895
rect 146 1867 184 1895
rect 212 1867 250 1895
rect 278 1867 316 1895
rect 344 1867 349 1895
rect -349 1829 349 1867
rect -349 1801 -344 1829
rect -316 1801 -278 1829
rect -250 1801 -212 1829
rect -184 1801 -146 1829
rect -118 1801 -80 1829
rect -52 1801 -14 1829
rect 14 1801 52 1829
rect 80 1801 118 1829
rect 146 1801 184 1829
rect 212 1801 250 1829
rect 278 1801 316 1829
rect 344 1801 349 1829
rect -349 1763 349 1801
rect -349 1735 -344 1763
rect -316 1735 -278 1763
rect -250 1735 -212 1763
rect -184 1735 -146 1763
rect -118 1735 -80 1763
rect -52 1735 -14 1763
rect 14 1735 52 1763
rect 80 1735 118 1763
rect 146 1735 184 1763
rect 212 1735 250 1763
rect 278 1735 316 1763
rect 344 1735 349 1763
rect -349 1697 349 1735
rect -349 1669 -344 1697
rect -316 1669 -278 1697
rect -250 1669 -212 1697
rect -184 1669 -146 1697
rect -118 1669 -80 1697
rect -52 1669 -14 1697
rect 14 1669 52 1697
rect 80 1669 118 1697
rect 146 1669 184 1697
rect 212 1669 250 1697
rect 278 1669 316 1697
rect 344 1669 349 1697
rect -349 1631 349 1669
rect -349 1603 -344 1631
rect -316 1603 -278 1631
rect -250 1603 -212 1631
rect -184 1603 -146 1631
rect -118 1603 -80 1631
rect -52 1603 -14 1631
rect 14 1603 52 1631
rect 80 1603 118 1631
rect 146 1603 184 1631
rect 212 1603 250 1631
rect 278 1603 316 1631
rect 344 1603 349 1631
rect -349 1565 349 1603
rect -349 1537 -344 1565
rect -316 1537 -278 1565
rect -250 1537 -212 1565
rect -184 1537 -146 1565
rect -118 1537 -80 1565
rect -52 1537 -14 1565
rect 14 1537 52 1565
rect 80 1537 118 1565
rect 146 1537 184 1565
rect 212 1537 250 1565
rect 278 1537 316 1565
rect 344 1537 349 1565
rect -349 1499 349 1537
rect -349 1471 -344 1499
rect -316 1471 -278 1499
rect -250 1471 -212 1499
rect -184 1471 -146 1499
rect -118 1471 -80 1499
rect -52 1471 -14 1499
rect 14 1471 52 1499
rect 80 1471 118 1499
rect 146 1471 184 1499
rect 212 1471 250 1499
rect 278 1471 316 1499
rect 344 1471 349 1499
rect -349 1433 349 1471
rect -349 1405 -344 1433
rect -316 1405 -278 1433
rect -250 1405 -212 1433
rect -184 1405 -146 1433
rect -118 1405 -80 1433
rect -52 1405 -14 1433
rect 14 1405 52 1433
rect 80 1405 118 1433
rect 146 1405 184 1433
rect 212 1405 250 1433
rect 278 1405 316 1433
rect 344 1405 349 1433
rect -349 1367 349 1405
rect -349 1339 -344 1367
rect -316 1339 -278 1367
rect -250 1339 -212 1367
rect -184 1339 -146 1367
rect -118 1339 -80 1367
rect -52 1339 -14 1367
rect 14 1339 52 1367
rect 80 1339 118 1367
rect 146 1339 184 1367
rect 212 1339 250 1367
rect 278 1339 316 1367
rect 344 1339 349 1367
rect -349 1301 349 1339
rect -349 1273 -344 1301
rect -316 1273 -278 1301
rect -250 1273 -212 1301
rect -184 1273 -146 1301
rect -118 1273 -80 1301
rect -52 1273 -14 1301
rect 14 1273 52 1301
rect 80 1273 118 1301
rect 146 1273 184 1301
rect 212 1273 250 1301
rect 278 1273 316 1301
rect 344 1273 349 1301
rect -349 1235 349 1273
rect -349 1207 -344 1235
rect -316 1207 -278 1235
rect -250 1207 -212 1235
rect -184 1207 -146 1235
rect -118 1207 -80 1235
rect -52 1207 -14 1235
rect 14 1207 52 1235
rect 80 1207 118 1235
rect 146 1207 184 1235
rect 212 1207 250 1235
rect 278 1207 316 1235
rect 344 1207 349 1235
rect -349 1169 349 1207
rect -349 1141 -344 1169
rect -316 1141 -278 1169
rect -250 1141 -212 1169
rect -184 1141 -146 1169
rect -118 1141 -80 1169
rect -52 1141 -14 1169
rect 14 1141 52 1169
rect 80 1141 118 1169
rect 146 1141 184 1169
rect 212 1141 250 1169
rect 278 1141 316 1169
rect 344 1141 349 1169
rect -349 1103 349 1141
rect -349 1075 -344 1103
rect -316 1075 -278 1103
rect -250 1075 -212 1103
rect -184 1075 -146 1103
rect -118 1075 -80 1103
rect -52 1075 -14 1103
rect 14 1075 52 1103
rect 80 1075 118 1103
rect 146 1075 184 1103
rect 212 1075 250 1103
rect 278 1075 316 1103
rect 344 1075 349 1103
rect -349 1037 349 1075
rect -349 1009 -344 1037
rect -316 1009 -278 1037
rect -250 1009 -212 1037
rect -184 1009 -146 1037
rect -118 1009 -80 1037
rect -52 1009 -14 1037
rect 14 1009 52 1037
rect 80 1009 118 1037
rect 146 1009 184 1037
rect 212 1009 250 1037
rect 278 1009 316 1037
rect 344 1009 349 1037
rect -349 971 349 1009
rect -349 943 -344 971
rect -316 943 -278 971
rect -250 943 -212 971
rect -184 943 -146 971
rect -118 943 -80 971
rect -52 943 -14 971
rect 14 943 52 971
rect 80 943 118 971
rect 146 943 184 971
rect 212 943 250 971
rect 278 943 316 971
rect 344 943 349 971
rect -349 905 349 943
rect -349 877 -344 905
rect -316 877 -278 905
rect -250 877 -212 905
rect -184 877 -146 905
rect -118 877 -80 905
rect -52 877 -14 905
rect 14 877 52 905
rect 80 877 118 905
rect 146 877 184 905
rect 212 877 250 905
rect 278 877 316 905
rect 344 877 349 905
rect -349 839 349 877
rect -349 811 -344 839
rect -316 811 -278 839
rect -250 811 -212 839
rect -184 811 -146 839
rect -118 811 -80 839
rect -52 811 -14 839
rect 14 811 52 839
rect 80 811 118 839
rect 146 811 184 839
rect 212 811 250 839
rect 278 811 316 839
rect 344 811 349 839
rect -349 773 349 811
rect -349 745 -344 773
rect -316 745 -278 773
rect -250 745 -212 773
rect -184 745 -146 773
rect -118 745 -80 773
rect -52 745 -14 773
rect 14 745 52 773
rect 80 745 118 773
rect 146 745 184 773
rect 212 745 250 773
rect 278 745 316 773
rect 344 745 349 773
rect -349 707 349 745
rect -349 679 -344 707
rect -316 679 -278 707
rect -250 679 -212 707
rect -184 679 -146 707
rect -118 679 -80 707
rect -52 679 -14 707
rect 14 679 52 707
rect 80 679 118 707
rect 146 679 184 707
rect 212 679 250 707
rect 278 679 316 707
rect 344 679 349 707
rect -349 641 349 679
rect -349 613 -344 641
rect -316 613 -278 641
rect -250 613 -212 641
rect -184 613 -146 641
rect -118 613 -80 641
rect -52 613 -14 641
rect 14 613 52 641
rect 80 613 118 641
rect 146 613 184 641
rect 212 613 250 641
rect 278 613 316 641
rect 344 613 349 641
rect -349 575 349 613
rect -349 547 -344 575
rect -316 547 -278 575
rect -250 547 -212 575
rect -184 547 -146 575
rect -118 547 -80 575
rect -52 547 -14 575
rect 14 547 52 575
rect 80 547 118 575
rect 146 547 184 575
rect 212 547 250 575
rect 278 547 316 575
rect 344 547 349 575
rect -349 509 349 547
rect -349 481 -344 509
rect -316 481 -278 509
rect -250 481 -212 509
rect -184 481 -146 509
rect -118 481 -80 509
rect -52 481 -14 509
rect 14 481 52 509
rect 80 481 118 509
rect 146 481 184 509
rect 212 481 250 509
rect 278 481 316 509
rect 344 481 349 509
rect -349 443 349 481
rect -349 415 -344 443
rect -316 415 -278 443
rect -250 415 -212 443
rect -184 415 -146 443
rect -118 415 -80 443
rect -52 415 -14 443
rect 14 415 52 443
rect 80 415 118 443
rect 146 415 184 443
rect 212 415 250 443
rect 278 415 316 443
rect 344 415 349 443
rect -349 377 349 415
rect -349 349 -344 377
rect -316 349 -278 377
rect -250 349 -212 377
rect -184 349 -146 377
rect -118 349 -80 377
rect -52 349 -14 377
rect 14 349 52 377
rect 80 349 118 377
rect 146 349 184 377
rect 212 349 250 377
rect 278 349 316 377
rect 344 349 349 377
rect -349 311 349 349
rect -349 283 -344 311
rect -316 283 -278 311
rect -250 283 -212 311
rect -184 283 -146 311
rect -118 283 -80 311
rect -52 283 -14 311
rect 14 283 52 311
rect 80 283 118 311
rect 146 283 184 311
rect 212 283 250 311
rect 278 283 316 311
rect 344 283 349 311
rect -349 245 349 283
rect -349 217 -344 245
rect -316 217 -278 245
rect -250 217 -212 245
rect -184 217 -146 245
rect -118 217 -80 245
rect -52 217 -14 245
rect 14 217 52 245
rect 80 217 118 245
rect 146 217 184 245
rect 212 217 250 245
rect 278 217 316 245
rect 344 217 349 245
rect -349 179 349 217
rect -349 151 -344 179
rect -316 151 -278 179
rect -250 151 -212 179
rect -184 151 -146 179
rect -118 151 -80 179
rect -52 151 -14 179
rect 14 151 52 179
rect 80 151 118 179
rect 146 151 184 179
rect 212 151 250 179
rect 278 151 316 179
rect 344 151 349 179
rect -349 113 349 151
rect -349 85 -344 113
rect -316 85 -278 113
rect -250 85 -212 113
rect -184 85 -146 113
rect -118 85 -80 113
rect -52 85 -14 113
rect 14 85 52 113
rect 80 85 118 113
rect 146 85 184 113
rect 212 85 250 113
rect 278 85 316 113
rect 344 85 349 113
rect -349 47 349 85
rect -349 19 -344 47
rect -316 19 -278 47
rect -250 19 -212 47
rect -184 19 -146 47
rect -118 19 -80 47
rect -52 19 -14 47
rect 14 19 52 47
rect 80 19 118 47
rect 146 19 184 47
rect 212 19 250 47
rect 278 19 316 47
rect 344 19 349 47
rect -349 -19 349 19
rect -349 -47 -344 -19
rect -316 -47 -278 -19
rect -250 -47 -212 -19
rect -184 -47 -146 -19
rect -118 -47 -80 -19
rect -52 -47 -14 -19
rect 14 -47 52 -19
rect 80 -47 118 -19
rect 146 -47 184 -19
rect 212 -47 250 -19
rect 278 -47 316 -19
rect 344 -47 349 -19
rect -349 -85 349 -47
rect -349 -113 -344 -85
rect -316 -113 -278 -85
rect -250 -113 -212 -85
rect -184 -113 -146 -85
rect -118 -113 -80 -85
rect -52 -113 -14 -85
rect 14 -113 52 -85
rect 80 -113 118 -85
rect 146 -113 184 -85
rect 212 -113 250 -85
rect 278 -113 316 -85
rect 344 -113 349 -85
rect -349 -151 349 -113
rect -349 -179 -344 -151
rect -316 -179 -278 -151
rect -250 -179 -212 -151
rect -184 -179 -146 -151
rect -118 -179 -80 -151
rect -52 -179 -14 -151
rect 14 -179 52 -151
rect 80 -179 118 -151
rect 146 -179 184 -151
rect 212 -179 250 -151
rect 278 -179 316 -151
rect 344 -179 349 -151
rect -349 -217 349 -179
rect -349 -245 -344 -217
rect -316 -245 -278 -217
rect -250 -245 -212 -217
rect -184 -245 -146 -217
rect -118 -245 -80 -217
rect -52 -245 -14 -217
rect 14 -245 52 -217
rect 80 -245 118 -217
rect 146 -245 184 -217
rect 212 -245 250 -217
rect 278 -245 316 -217
rect 344 -245 349 -217
rect -349 -283 349 -245
rect -349 -311 -344 -283
rect -316 -311 -278 -283
rect -250 -311 -212 -283
rect -184 -311 -146 -283
rect -118 -311 -80 -283
rect -52 -311 -14 -283
rect 14 -311 52 -283
rect 80 -311 118 -283
rect 146 -311 184 -283
rect 212 -311 250 -283
rect 278 -311 316 -283
rect 344 -311 349 -283
rect -349 -349 349 -311
rect -349 -377 -344 -349
rect -316 -377 -278 -349
rect -250 -377 -212 -349
rect -184 -377 -146 -349
rect -118 -377 -80 -349
rect -52 -377 -14 -349
rect 14 -377 52 -349
rect 80 -377 118 -349
rect 146 -377 184 -349
rect 212 -377 250 -349
rect 278 -377 316 -349
rect 344 -377 349 -349
rect -349 -415 349 -377
rect -349 -443 -344 -415
rect -316 -443 -278 -415
rect -250 -443 -212 -415
rect -184 -443 -146 -415
rect -118 -443 -80 -415
rect -52 -443 -14 -415
rect 14 -443 52 -415
rect 80 -443 118 -415
rect 146 -443 184 -415
rect 212 -443 250 -415
rect 278 -443 316 -415
rect 344 -443 349 -415
rect -349 -481 349 -443
rect -349 -509 -344 -481
rect -316 -509 -278 -481
rect -250 -509 -212 -481
rect -184 -509 -146 -481
rect -118 -509 -80 -481
rect -52 -509 -14 -481
rect 14 -509 52 -481
rect 80 -509 118 -481
rect 146 -509 184 -481
rect 212 -509 250 -481
rect 278 -509 316 -481
rect 344 -509 349 -481
rect -349 -547 349 -509
rect -349 -575 -344 -547
rect -316 -575 -278 -547
rect -250 -575 -212 -547
rect -184 -575 -146 -547
rect -118 -575 -80 -547
rect -52 -575 -14 -547
rect 14 -575 52 -547
rect 80 -575 118 -547
rect 146 -575 184 -547
rect 212 -575 250 -547
rect 278 -575 316 -547
rect 344 -575 349 -547
rect -349 -613 349 -575
rect -349 -641 -344 -613
rect -316 -641 -278 -613
rect -250 -641 -212 -613
rect -184 -641 -146 -613
rect -118 -641 -80 -613
rect -52 -641 -14 -613
rect 14 -641 52 -613
rect 80 -641 118 -613
rect 146 -641 184 -613
rect 212 -641 250 -613
rect 278 -641 316 -613
rect 344 -641 349 -613
rect -349 -679 349 -641
rect -349 -707 -344 -679
rect -316 -707 -278 -679
rect -250 -707 -212 -679
rect -184 -707 -146 -679
rect -118 -707 -80 -679
rect -52 -707 -14 -679
rect 14 -707 52 -679
rect 80 -707 118 -679
rect 146 -707 184 -679
rect 212 -707 250 -679
rect 278 -707 316 -679
rect 344 -707 349 -679
rect -349 -745 349 -707
rect -349 -773 -344 -745
rect -316 -773 -278 -745
rect -250 -773 -212 -745
rect -184 -773 -146 -745
rect -118 -773 -80 -745
rect -52 -773 -14 -745
rect 14 -773 52 -745
rect 80 -773 118 -745
rect 146 -773 184 -745
rect 212 -773 250 -745
rect 278 -773 316 -745
rect 344 -773 349 -745
rect -349 -811 349 -773
rect -349 -839 -344 -811
rect -316 -839 -278 -811
rect -250 -839 -212 -811
rect -184 -839 -146 -811
rect -118 -839 -80 -811
rect -52 -839 -14 -811
rect 14 -839 52 -811
rect 80 -839 118 -811
rect 146 -839 184 -811
rect 212 -839 250 -811
rect 278 -839 316 -811
rect 344 -839 349 -811
rect -349 -877 349 -839
rect -349 -905 -344 -877
rect -316 -905 -278 -877
rect -250 -905 -212 -877
rect -184 -905 -146 -877
rect -118 -905 -80 -877
rect -52 -905 -14 -877
rect 14 -905 52 -877
rect 80 -905 118 -877
rect 146 -905 184 -877
rect 212 -905 250 -877
rect 278 -905 316 -877
rect 344 -905 349 -877
rect -349 -943 349 -905
rect -349 -971 -344 -943
rect -316 -971 -278 -943
rect -250 -971 -212 -943
rect -184 -971 -146 -943
rect -118 -971 -80 -943
rect -52 -971 -14 -943
rect 14 -971 52 -943
rect 80 -971 118 -943
rect 146 -971 184 -943
rect 212 -971 250 -943
rect 278 -971 316 -943
rect 344 -971 349 -943
rect -349 -1009 349 -971
rect -349 -1037 -344 -1009
rect -316 -1037 -278 -1009
rect -250 -1037 -212 -1009
rect -184 -1037 -146 -1009
rect -118 -1037 -80 -1009
rect -52 -1037 -14 -1009
rect 14 -1037 52 -1009
rect 80 -1037 118 -1009
rect 146 -1037 184 -1009
rect 212 -1037 250 -1009
rect 278 -1037 316 -1009
rect 344 -1037 349 -1009
rect -349 -1075 349 -1037
rect -349 -1103 -344 -1075
rect -316 -1103 -278 -1075
rect -250 -1103 -212 -1075
rect -184 -1103 -146 -1075
rect -118 -1103 -80 -1075
rect -52 -1103 -14 -1075
rect 14 -1103 52 -1075
rect 80 -1103 118 -1075
rect 146 -1103 184 -1075
rect 212 -1103 250 -1075
rect 278 -1103 316 -1075
rect 344 -1103 349 -1075
rect -349 -1141 349 -1103
rect -349 -1169 -344 -1141
rect -316 -1169 -278 -1141
rect -250 -1169 -212 -1141
rect -184 -1169 -146 -1141
rect -118 -1169 -80 -1141
rect -52 -1169 -14 -1141
rect 14 -1169 52 -1141
rect 80 -1169 118 -1141
rect 146 -1169 184 -1141
rect 212 -1169 250 -1141
rect 278 -1169 316 -1141
rect 344 -1169 349 -1141
rect -349 -1207 349 -1169
rect -349 -1235 -344 -1207
rect -316 -1235 -278 -1207
rect -250 -1235 -212 -1207
rect -184 -1235 -146 -1207
rect -118 -1235 -80 -1207
rect -52 -1235 -14 -1207
rect 14 -1235 52 -1207
rect 80 -1235 118 -1207
rect 146 -1235 184 -1207
rect 212 -1235 250 -1207
rect 278 -1235 316 -1207
rect 344 -1235 349 -1207
rect -349 -1273 349 -1235
rect -349 -1301 -344 -1273
rect -316 -1301 -278 -1273
rect -250 -1301 -212 -1273
rect -184 -1301 -146 -1273
rect -118 -1301 -80 -1273
rect -52 -1301 -14 -1273
rect 14 -1301 52 -1273
rect 80 -1301 118 -1273
rect 146 -1301 184 -1273
rect 212 -1301 250 -1273
rect 278 -1301 316 -1273
rect 344 -1301 349 -1273
rect -349 -1339 349 -1301
rect -349 -1367 -344 -1339
rect -316 -1367 -278 -1339
rect -250 -1367 -212 -1339
rect -184 -1367 -146 -1339
rect -118 -1367 -80 -1339
rect -52 -1367 -14 -1339
rect 14 -1367 52 -1339
rect 80 -1367 118 -1339
rect 146 -1367 184 -1339
rect 212 -1367 250 -1339
rect 278 -1367 316 -1339
rect 344 -1367 349 -1339
rect -349 -1405 349 -1367
rect -349 -1433 -344 -1405
rect -316 -1433 -278 -1405
rect -250 -1433 -212 -1405
rect -184 -1433 -146 -1405
rect -118 -1433 -80 -1405
rect -52 -1433 -14 -1405
rect 14 -1433 52 -1405
rect 80 -1433 118 -1405
rect 146 -1433 184 -1405
rect 212 -1433 250 -1405
rect 278 -1433 316 -1405
rect 344 -1433 349 -1405
rect -349 -1471 349 -1433
rect -349 -1499 -344 -1471
rect -316 -1499 -278 -1471
rect -250 -1499 -212 -1471
rect -184 -1499 -146 -1471
rect -118 -1499 -80 -1471
rect -52 -1499 -14 -1471
rect 14 -1499 52 -1471
rect 80 -1499 118 -1471
rect 146 -1499 184 -1471
rect 212 -1499 250 -1471
rect 278 -1499 316 -1471
rect 344 -1499 349 -1471
rect -349 -1537 349 -1499
rect -349 -1565 -344 -1537
rect -316 -1565 -278 -1537
rect -250 -1565 -212 -1537
rect -184 -1565 -146 -1537
rect -118 -1565 -80 -1537
rect -52 -1565 -14 -1537
rect 14 -1565 52 -1537
rect 80 -1565 118 -1537
rect 146 -1565 184 -1537
rect 212 -1565 250 -1537
rect 278 -1565 316 -1537
rect 344 -1565 349 -1537
rect -349 -1603 349 -1565
rect -349 -1631 -344 -1603
rect -316 -1631 -278 -1603
rect -250 -1631 -212 -1603
rect -184 -1631 -146 -1603
rect -118 -1631 -80 -1603
rect -52 -1631 -14 -1603
rect 14 -1631 52 -1603
rect 80 -1631 118 -1603
rect 146 -1631 184 -1603
rect 212 -1631 250 -1603
rect 278 -1631 316 -1603
rect 344 -1631 349 -1603
rect -349 -1669 349 -1631
rect -349 -1697 -344 -1669
rect -316 -1697 -278 -1669
rect -250 -1697 -212 -1669
rect -184 -1697 -146 -1669
rect -118 -1697 -80 -1669
rect -52 -1697 -14 -1669
rect 14 -1697 52 -1669
rect 80 -1697 118 -1669
rect 146 -1697 184 -1669
rect 212 -1697 250 -1669
rect 278 -1697 316 -1669
rect 344 -1697 349 -1669
rect -349 -1735 349 -1697
rect -349 -1763 -344 -1735
rect -316 -1763 -278 -1735
rect -250 -1763 -212 -1735
rect -184 -1763 -146 -1735
rect -118 -1763 -80 -1735
rect -52 -1763 -14 -1735
rect 14 -1763 52 -1735
rect 80 -1763 118 -1735
rect 146 -1763 184 -1735
rect 212 -1763 250 -1735
rect 278 -1763 316 -1735
rect 344 -1763 349 -1735
rect -349 -1801 349 -1763
rect -349 -1829 -344 -1801
rect -316 -1829 -278 -1801
rect -250 -1829 -212 -1801
rect -184 -1829 -146 -1801
rect -118 -1829 -80 -1801
rect -52 -1829 -14 -1801
rect 14 -1829 52 -1801
rect 80 -1829 118 -1801
rect 146 -1829 184 -1801
rect 212 -1829 250 -1801
rect 278 -1829 316 -1801
rect 344 -1829 349 -1801
rect -349 -1867 349 -1829
rect -349 -1895 -344 -1867
rect -316 -1895 -278 -1867
rect -250 -1895 -212 -1867
rect -184 -1895 -146 -1867
rect -118 -1895 -80 -1867
rect -52 -1895 -14 -1867
rect 14 -1895 52 -1867
rect 80 -1895 118 -1867
rect 146 -1895 184 -1867
rect 212 -1895 250 -1867
rect 278 -1895 316 -1867
rect 344 -1895 349 -1867
rect -349 -1933 349 -1895
rect -349 -1961 -344 -1933
rect -316 -1961 -278 -1933
rect -250 -1961 -212 -1933
rect -184 -1961 -146 -1933
rect -118 -1961 -80 -1933
rect -52 -1961 -14 -1933
rect 14 -1961 52 -1933
rect 80 -1961 118 -1933
rect 146 -1961 184 -1933
rect 212 -1961 250 -1933
rect 278 -1961 316 -1933
rect 344 -1961 349 -1933
rect -349 -1999 349 -1961
rect -349 -2027 -344 -1999
rect -316 -2027 -278 -1999
rect -250 -2027 -212 -1999
rect -184 -2027 -146 -1999
rect -118 -2027 -80 -1999
rect -52 -2027 -14 -1999
rect 14 -2027 52 -1999
rect 80 -2027 118 -1999
rect 146 -2027 184 -1999
rect 212 -2027 250 -1999
rect 278 -2027 316 -1999
rect 344 -2027 349 -1999
rect -349 -2065 349 -2027
rect -349 -2093 -344 -2065
rect -316 -2093 -278 -2065
rect -250 -2093 -212 -2065
rect -184 -2093 -146 -2065
rect -118 -2093 -80 -2065
rect -52 -2093 -14 -2065
rect 14 -2093 52 -2065
rect 80 -2093 118 -2065
rect 146 -2093 184 -2065
rect 212 -2093 250 -2065
rect 278 -2093 316 -2065
rect 344 -2093 349 -2065
rect -349 -2131 349 -2093
rect -349 -2159 -344 -2131
rect -316 -2159 -278 -2131
rect -250 -2159 -212 -2131
rect -184 -2159 -146 -2131
rect -118 -2159 -80 -2131
rect -52 -2159 -14 -2131
rect 14 -2159 52 -2131
rect 80 -2159 118 -2131
rect 146 -2159 184 -2131
rect 212 -2159 250 -2131
rect 278 -2159 316 -2131
rect 344 -2159 349 -2131
rect -349 -2197 349 -2159
rect -349 -2225 -344 -2197
rect -316 -2225 -278 -2197
rect -250 -2225 -212 -2197
rect -184 -2225 -146 -2197
rect -118 -2225 -80 -2197
rect -52 -2225 -14 -2197
rect 14 -2225 52 -2197
rect 80 -2225 118 -2197
rect 146 -2225 184 -2197
rect 212 -2225 250 -2197
rect 278 -2225 316 -2197
rect 344 -2225 349 -2197
rect -349 -2263 349 -2225
rect -349 -2291 -344 -2263
rect -316 -2291 -278 -2263
rect -250 -2291 -212 -2263
rect -184 -2291 -146 -2263
rect -118 -2291 -80 -2263
rect -52 -2291 -14 -2263
rect 14 -2291 52 -2263
rect 80 -2291 118 -2263
rect 146 -2291 184 -2263
rect 212 -2291 250 -2263
rect 278 -2291 316 -2263
rect 344 -2291 349 -2263
rect -349 -2329 349 -2291
rect -349 -2357 -344 -2329
rect -316 -2357 -278 -2329
rect -250 -2357 -212 -2329
rect -184 -2357 -146 -2329
rect -118 -2357 -80 -2329
rect -52 -2357 -14 -2329
rect 14 -2357 52 -2329
rect 80 -2357 118 -2329
rect 146 -2357 184 -2329
rect 212 -2357 250 -2329
rect 278 -2357 316 -2329
rect 344 -2357 349 -2329
rect -349 -2395 349 -2357
rect -349 -2423 -344 -2395
rect -316 -2423 -278 -2395
rect -250 -2423 -212 -2395
rect -184 -2423 -146 -2395
rect -118 -2423 -80 -2395
rect -52 -2423 -14 -2395
rect 14 -2423 52 -2395
rect 80 -2423 118 -2395
rect 146 -2423 184 -2395
rect 212 -2423 250 -2395
rect 278 -2423 316 -2395
rect 344 -2423 349 -2395
rect -349 -2461 349 -2423
rect -349 -2489 -344 -2461
rect -316 -2489 -278 -2461
rect -250 -2489 -212 -2461
rect -184 -2489 -146 -2461
rect -118 -2489 -80 -2461
rect -52 -2489 -14 -2461
rect 14 -2489 52 -2461
rect 80 -2489 118 -2461
rect 146 -2489 184 -2461
rect 212 -2489 250 -2461
rect 278 -2489 316 -2461
rect 344 -2489 349 -2461
rect -349 -2527 349 -2489
rect -349 -2555 -344 -2527
rect -316 -2555 -278 -2527
rect -250 -2555 -212 -2527
rect -184 -2555 -146 -2527
rect -118 -2555 -80 -2527
rect -52 -2555 -14 -2527
rect 14 -2555 52 -2527
rect 80 -2555 118 -2527
rect 146 -2555 184 -2527
rect 212 -2555 250 -2527
rect 278 -2555 316 -2527
rect 344 -2555 349 -2527
rect -349 -2593 349 -2555
rect -349 -2621 -344 -2593
rect -316 -2621 -278 -2593
rect -250 -2621 -212 -2593
rect -184 -2621 -146 -2593
rect -118 -2621 -80 -2593
rect -52 -2621 -14 -2593
rect 14 -2621 52 -2593
rect 80 -2621 118 -2593
rect 146 -2621 184 -2593
rect 212 -2621 250 -2593
rect 278 -2621 316 -2593
rect 344 -2621 349 -2593
rect -349 -2659 349 -2621
rect -349 -2687 -344 -2659
rect -316 -2687 -278 -2659
rect -250 -2687 -212 -2659
rect -184 -2687 -146 -2659
rect -118 -2687 -80 -2659
rect -52 -2687 -14 -2659
rect 14 -2687 52 -2659
rect 80 -2687 118 -2659
rect 146 -2687 184 -2659
rect 212 -2687 250 -2659
rect 278 -2687 316 -2659
rect 344 -2687 349 -2659
rect -349 -2725 349 -2687
rect -349 -2753 -344 -2725
rect -316 -2753 -278 -2725
rect -250 -2753 -212 -2725
rect -184 -2753 -146 -2725
rect -118 -2753 -80 -2725
rect -52 -2753 -14 -2725
rect 14 -2753 52 -2725
rect 80 -2753 118 -2725
rect 146 -2753 184 -2725
rect 212 -2753 250 -2725
rect 278 -2753 316 -2725
rect 344 -2753 349 -2725
rect -349 -2791 349 -2753
rect -349 -2819 -344 -2791
rect -316 -2819 -278 -2791
rect -250 -2819 -212 -2791
rect -184 -2819 -146 -2791
rect -118 -2819 -80 -2791
rect -52 -2819 -14 -2791
rect 14 -2819 52 -2791
rect 80 -2819 118 -2791
rect 146 -2819 184 -2791
rect 212 -2819 250 -2791
rect 278 -2819 316 -2791
rect 344 -2819 349 -2791
rect -349 -2857 349 -2819
rect -349 -2885 -344 -2857
rect -316 -2885 -278 -2857
rect -250 -2885 -212 -2857
rect -184 -2885 -146 -2857
rect -118 -2885 -80 -2857
rect -52 -2885 -14 -2857
rect 14 -2885 52 -2857
rect 80 -2885 118 -2857
rect 146 -2885 184 -2857
rect 212 -2885 250 -2857
rect 278 -2885 316 -2857
rect 344 -2885 349 -2857
rect -349 -2923 349 -2885
rect -349 -2951 -344 -2923
rect -316 -2951 -278 -2923
rect -250 -2951 -212 -2923
rect -184 -2951 -146 -2923
rect -118 -2951 -80 -2923
rect -52 -2951 -14 -2923
rect 14 -2951 52 -2923
rect 80 -2951 118 -2923
rect 146 -2951 184 -2923
rect 212 -2951 250 -2923
rect 278 -2951 316 -2923
rect 344 -2951 349 -2923
rect -349 -2989 349 -2951
rect -349 -3017 -344 -2989
rect -316 -3017 -278 -2989
rect -250 -3017 -212 -2989
rect -184 -3017 -146 -2989
rect -118 -3017 -80 -2989
rect -52 -3017 -14 -2989
rect 14 -3017 52 -2989
rect 80 -3017 118 -2989
rect 146 -3017 184 -2989
rect 212 -3017 250 -2989
rect 278 -3017 316 -2989
rect 344 -3017 349 -2989
rect -349 -3055 349 -3017
rect -349 -3083 -344 -3055
rect -316 -3083 -278 -3055
rect -250 -3083 -212 -3055
rect -184 -3083 -146 -3055
rect -118 -3083 -80 -3055
rect -52 -3083 -14 -3055
rect 14 -3083 52 -3055
rect 80 -3083 118 -3055
rect 146 -3083 184 -3055
rect 212 -3083 250 -3055
rect 278 -3083 316 -3055
rect 344 -3083 349 -3055
rect -349 -3121 349 -3083
rect -349 -3149 -344 -3121
rect -316 -3149 -278 -3121
rect -250 -3149 -212 -3121
rect -184 -3149 -146 -3121
rect -118 -3149 -80 -3121
rect -52 -3149 -14 -3121
rect 14 -3149 52 -3121
rect 80 -3149 118 -3121
rect 146 -3149 184 -3121
rect 212 -3149 250 -3121
rect 278 -3149 316 -3121
rect 344 -3149 349 -3121
rect -349 -3187 349 -3149
rect -349 -3215 -344 -3187
rect -316 -3215 -278 -3187
rect -250 -3215 -212 -3187
rect -184 -3215 -146 -3187
rect -118 -3215 -80 -3187
rect -52 -3215 -14 -3187
rect 14 -3215 52 -3187
rect 80 -3215 118 -3187
rect 146 -3215 184 -3187
rect 212 -3215 250 -3187
rect 278 -3215 316 -3187
rect 344 -3215 349 -3187
rect -349 -3253 349 -3215
rect -349 -3281 -344 -3253
rect -316 -3281 -278 -3253
rect -250 -3281 -212 -3253
rect -184 -3281 -146 -3253
rect -118 -3281 -80 -3253
rect -52 -3281 -14 -3253
rect 14 -3281 52 -3253
rect 80 -3281 118 -3253
rect 146 -3281 184 -3253
rect 212 -3281 250 -3253
rect 278 -3281 316 -3253
rect 344 -3281 349 -3253
rect -349 -3319 349 -3281
rect -349 -3347 -344 -3319
rect -316 -3347 -278 -3319
rect -250 -3347 -212 -3319
rect -184 -3347 -146 -3319
rect -118 -3347 -80 -3319
rect -52 -3347 -14 -3319
rect 14 -3347 52 -3319
rect 80 -3347 118 -3319
rect 146 -3347 184 -3319
rect 212 -3347 250 -3319
rect 278 -3347 316 -3319
rect 344 -3347 349 -3319
rect -349 -3385 349 -3347
rect -349 -3413 -344 -3385
rect -316 -3413 -278 -3385
rect -250 -3413 -212 -3385
rect -184 -3413 -146 -3385
rect -118 -3413 -80 -3385
rect -52 -3413 -14 -3385
rect 14 -3413 52 -3385
rect 80 -3413 118 -3385
rect 146 -3413 184 -3385
rect 212 -3413 250 -3385
rect 278 -3413 316 -3385
rect 344 -3413 349 -3385
rect -349 -3451 349 -3413
rect -349 -3479 -344 -3451
rect -316 -3479 -278 -3451
rect -250 -3479 -212 -3451
rect -184 -3479 -146 -3451
rect -118 -3479 -80 -3451
rect -52 -3479 -14 -3451
rect 14 -3479 52 -3451
rect 80 -3479 118 -3451
rect 146 -3479 184 -3451
rect 212 -3479 250 -3451
rect 278 -3479 316 -3451
rect 344 -3479 349 -3451
rect -349 -3517 349 -3479
rect -349 -3545 -344 -3517
rect -316 -3545 -278 -3517
rect -250 -3545 -212 -3517
rect -184 -3545 -146 -3517
rect -118 -3545 -80 -3517
rect -52 -3545 -14 -3517
rect 14 -3545 52 -3517
rect 80 -3545 118 -3517
rect 146 -3545 184 -3517
rect 212 -3545 250 -3517
rect 278 -3545 316 -3517
rect 344 -3545 349 -3517
rect -349 -3583 349 -3545
rect -349 -3611 -344 -3583
rect -316 -3611 -278 -3583
rect -250 -3611 -212 -3583
rect -184 -3611 -146 -3583
rect -118 -3611 -80 -3583
rect -52 -3611 -14 -3583
rect 14 -3611 52 -3583
rect 80 -3611 118 -3583
rect 146 -3611 184 -3583
rect 212 -3611 250 -3583
rect 278 -3611 316 -3583
rect 344 -3611 349 -3583
rect -349 -3649 349 -3611
rect -349 -3677 -344 -3649
rect -316 -3677 -278 -3649
rect -250 -3677 -212 -3649
rect -184 -3677 -146 -3649
rect -118 -3677 -80 -3649
rect -52 -3677 -14 -3649
rect 14 -3677 52 -3649
rect 80 -3677 118 -3649
rect 146 -3677 184 -3649
rect 212 -3677 250 -3649
rect 278 -3677 316 -3649
rect 344 -3677 349 -3649
rect -349 -3715 349 -3677
rect -349 -3743 -344 -3715
rect -316 -3743 -278 -3715
rect -250 -3743 -212 -3715
rect -184 -3743 -146 -3715
rect -118 -3743 -80 -3715
rect -52 -3743 -14 -3715
rect 14 -3743 52 -3715
rect 80 -3743 118 -3715
rect 146 -3743 184 -3715
rect 212 -3743 250 -3715
rect 278 -3743 316 -3715
rect 344 -3743 349 -3715
rect -349 -3781 349 -3743
rect -349 -3809 -344 -3781
rect -316 -3809 -278 -3781
rect -250 -3809 -212 -3781
rect -184 -3809 -146 -3781
rect -118 -3809 -80 -3781
rect -52 -3809 -14 -3781
rect 14 -3809 52 -3781
rect 80 -3809 118 -3781
rect 146 -3809 184 -3781
rect 212 -3809 250 -3781
rect 278 -3809 316 -3781
rect 344 -3809 349 -3781
rect -349 -3847 349 -3809
rect -349 -3875 -344 -3847
rect -316 -3875 -278 -3847
rect -250 -3875 -212 -3847
rect -184 -3875 -146 -3847
rect -118 -3875 -80 -3847
rect -52 -3875 -14 -3847
rect 14 -3875 52 -3847
rect 80 -3875 118 -3847
rect 146 -3875 184 -3847
rect 212 -3875 250 -3847
rect 278 -3875 316 -3847
rect 344 -3875 349 -3847
rect -349 -3913 349 -3875
rect -349 -3941 -344 -3913
rect -316 -3941 -278 -3913
rect -250 -3941 -212 -3913
rect -184 -3941 -146 -3913
rect -118 -3941 -80 -3913
rect -52 -3941 -14 -3913
rect 14 -3941 52 -3913
rect 80 -3941 118 -3913
rect 146 -3941 184 -3913
rect 212 -3941 250 -3913
rect 278 -3941 316 -3913
rect 344 -3941 349 -3913
rect -349 -3979 349 -3941
rect -349 -4007 -344 -3979
rect -316 -4007 -278 -3979
rect -250 -4007 -212 -3979
rect -184 -4007 -146 -3979
rect -118 -4007 -80 -3979
rect -52 -4007 -14 -3979
rect 14 -4007 52 -3979
rect 80 -4007 118 -3979
rect 146 -4007 184 -3979
rect 212 -4007 250 -3979
rect 278 -4007 316 -3979
rect 344 -4007 349 -3979
rect -349 -4045 349 -4007
rect -349 -4073 -344 -4045
rect -316 -4073 -278 -4045
rect -250 -4073 -212 -4045
rect -184 -4073 -146 -4045
rect -118 -4073 -80 -4045
rect -52 -4073 -14 -4045
rect 14 -4073 52 -4045
rect 80 -4073 118 -4045
rect 146 -4073 184 -4045
rect 212 -4073 250 -4045
rect 278 -4073 316 -4045
rect 344 -4073 349 -4045
rect -349 -4111 349 -4073
rect -349 -4139 -344 -4111
rect -316 -4139 -278 -4111
rect -250 -4139 -212 -4111
rect -184 -4139 -146 -4111
rect -118 -4139 -80 -4111
rect -52 -4139 -14 -4111
rect 14 -4139 52 -4111
rect 80 -4139 118 -4111
rect 146 -4139 184 -4111
rect 212 -4139 250 -4111
rect 278 -4139 316 -4111
rect 344 -4139 349 -4111
rect -349 -4177 349 -4139
rect -349 -4205 -344 -4177
rect -316 -4205 -278 -4177
rect -250 -4205 -212 -4177
rect -184 -4205 -146 -4177
rect -118 -4205 -80 -4177
rect -52 -4205 -14 -4177
rect 14 -4205 52 -4177
rect 80 -4205 118 -4177
rect 146 -4205 184 -4177
rect 212 -4205 250 -4177
rect 278 -4205 316 -4177
rect 344 -4205 349 -4177
rect -349 -4243 349 -4205
rect -349 -4271 -344 -4243
rect -316 -4271 -278 -4243
rect -250 -4271 -212 -4243
rect -184 -4271 -146 -4243
rect -118 -4271 -80 -4243
rect -52 -4271 -14 -4243
rect 14 -4271 52 -4243
rect 80 -4271 118 -4243
rect 146 -4271 184 -4243
rect 212 -4271 250 -4243
rect 278 -4271 316 -4243
rect 344 -4271 349 -4243
rect -349 -4309 349 -4271
rect -349 -4337 -344 -4309
rect -316 -4337 -278 -4309
rect -250 -4337 -212 -4309
rect -184 -4337 -146 -4309
rect -118 -4337 -80 -4309
rect -52 -4337 -14 -4309
rect 14 -4337 52 -4309
rect 80 -4337 118 -4309
rect 146 -4337 184 -4309
rect 212 -4337 250 -4309
rect 278 -4337 316 -4309
rect 344 -4337 349 -4309
rect -349 -4375 349 -4337
rect -349 -4403 -344 -4375
rect -316 -4403 -278 -4375
rect -250 -4403 -212 -4375
rect -184 -4403 -146 -4375
rect -118 -4403 -80 -4375
rect -52 -4403 -14 -4375
rect 14 -4403 52 -4375
rect 80 -4403 118 -4375
rect 146 -4403 184 -4375
rect 212 -4403 250 -4375
rect 278 -4403 316 -4375
rect 344 -4403 349 -4375
rect -349 -4441 349 -4403
rect -349 -4469 -344 -4441
rect -316 -4469 -278 -4441
rect -250 -4469 -212 -4441
rect -184 -4469 -146 -4441
rect -118 -4469 -80 -4441
rect -52 -4469 -14 -4441
rect 14 -4469 52 -4441
rect 80 -4469 118 -4441
rect 146 -4469 184 -4441
rect 212 -4469 250 -4441
rect 278 -4469 316 -4441
rect 344 -4469 349 -4441
rect -349 -4507 349 -4469
rect -349 -4535 -344 -4507
rect -316 -4535 -278 -4507
rect -250 -4535 -212 -4507
rect -184 -4535 -146 -4507
rect -118 -4535 -80 -4507
rect -52 -4535 -14 -4507
rect 14 -4535 52 -4507
rect 80 -4535 118 -4507
rect 146 -4535 184 -4507
rect 212 -4535 250 -4507
rect 278 -4535 316 -4507
rect 344 -4535 349 -4507
rect -349 -4573 349 -4535
rect -349 -4601 -344 -4573
rect -316 -4601 -278 -4573
rect -250 -4601 -212 -4573
rect -184 -4601 -146 -4573
rect -118 -4601 -80 -4573
rect -52 -4601 -14 -4573
rect 14 -4601 52 -4573
rect 80 -4601 118 -4573
rect 146 -4601 184 -4573
rect 212 -4601 250 -4573
rect 278 -4601 316 -4573
rect 344 -4601 349 -4573
rect -349 -4639 349 -4601
rect -349 -4667 -344 -4639
rect -316 -4667 -278 -4639
rect -250 -4667 -212 -4639
rect -184 -4667 -146 -4639
rect -118 -4667 -80 -4639
rect -52 -4667 -14 -4639
rect 14 -4667 52 -4639
rect 80 -4667 118 -4639
rect 146 -4667 184 -4639
rect 212 -4667 250 -4639
rect 278 -4667 316 -4639
rect 344 -4667 349 -4639
rect -349 -4705 349 -4667
rect -349 -4733 -344 -4705
rect -316 -4733 -278 -4705
rect -250 -4733 -212 -4705
rect -184 -4733 -146 -4705
rect -118 -4733 -80 -4705
rect -52 -4733 -14 -4705
rect 14 -4733 52 -4705
rect 80 -4733 118 -4705
rect 146 -4733 184 -4705
rect 212 -4733 250 -4705
rect 278 -4733 316 -4705
rect 344 -4733 349 -4705
rect -349 -4771 349 -4733
rect -349 -4799 -344 -4771
rect -316 -4799 -278 -4771
rect -250 -4799 -212 -4771
rect -184 -4799 -146 -4771
rect -118 -4799 -80 -4771
rect -52 -4799 -14 -4771
rect 14 -4799 52 -4771
rect 80 -4799 118 -4771
rect 146 -4799 184 -4771
rect 212 -4799 250 -4771
rect 278 -4799 316 -4771
rect 344 -4799 349 -4771
rect -349 -4837 349 -4799
rect -349 -4865 -344 -4837
rect -316 -4865 -278 -4837
rect -250 -4865 -212 -4837
rect -184 -4865 -146 -4837
rect -118 -4865 -80 -4837
rect -52 -4865 -14 -4837
rect 14 -4865 52 -4837
rect 80 -4865 118 -4837
rect 146 -4865 184 -4837
rect 212 -4865 250 -4837
rect 278 -4865 316 -4837
rect 344 -4865 349 -4837
rect -349 -4903 349 -4865
rect -349 -4931 -344 -4903
rect -316 -4931 -278 -4903
rect -250 -4931 -212 -4903
rect -184 -4931 -146 -4903
rect -118 -4931 -80 -4903
rect -52 -4931 -14 -4903
rect 14 -4931 52 -4903
rect 80 -4931 118 -4903
rect 146 -4931 184 -4903
rect 212 -4931 250 -4903
rect 278 -4931 316 -4903
rect 344 -4931 349 -4903
rect -349 -4969 349 -4931
rect -349 -4997 -344 -4969
rect -316 -4997 -278 -4969
rect -250 -4997 -212 -4969
rect -184 -4997 -146 -4969
rect -118 -4997 -80 -4969
rect -52 -4997 -14 -4969
rect 14 -4997 52 -4969
rect 80 -4997 118 -4969
rect 146 -4997 184 -4969
rect 212 -4997 250 -4969
rect 278 -4997 316 -4969
rect 344 -4997 349 -4969
rect -349 -5035 349 -4997
rect -349 -5063 -344 -5035
rect -316 -5063 -278 -5035
rect -250 -5063 -212 -5035
rect -184 -5063 -146 -5035
rect -118 -5063 -80 -5035
rect -52 -5063 -14 -5035
rect 14 -5063 52 -5035
rect 80 -5063 118 -5035
rect 146 -5063 184 -5035
rect 212 -5063 250 -5035
rect 278 -5063 316 -5035
rect 344 -5063 349 -5035
rect -349 -5068 349 -5063
<< via3 >>
rect -344 5035 -316 5063
rect -278 5035 -250 5063
rect -212 5035 -184 5063
rect -146 5035 -118 5063
rect -80 5035 -52 5063
rect -14 5035 14 5063
rect 52 5035 80 5063
rect 118 5035 146 5063
rect 184 5035 212 5063
rect 250 5035 278 5063
rect 316 5035 344 5063
rect -344 4969 -316 4997
rect -278 4969 -250 4997
rect -212 4969 -184 4997
rect -146 4969 -118 4997
rect -80 4969 -52 4997
rect -14 4969 14 4997
rect 52 4969 80 4997
rect 118 4969 146 4997
rect 184 4969 212 4997
rect 250 4969 278 4997
rect 316 4969 344 4997
rect -344 4903 -316 4931
rect -278 4903 -250 4931
rect -212 4903 -184 4931
rect -146 4903 -118 4931
rect -80 4903 -52 4931
rect -14 4903 14 4931
rect 52 4903 80 4931
rect 118 4903 146 4931
rect 184 4903 212 4931
rect 250 4903 278 4931
rect 316 4903 344 4931
rect -344 4837 -316 4865
rect -278 4837 -250 4865
rect -212 4837 -184 4865
rect -146 4837 -118 4865
rect -80 4837 -52 4865
rect -14 4837 14 4865
rect 52 4837 80 4865
rect 118 4837 146 4865
rect 184 4837 212 4865
rect 250 4837 278 4865
rect 316 4837 344 4865
rect -344 4771 -316 4799
rect -278 4771 -250 4799
rect -212 4771 -184 4799
rect -146 4771 -118 4799
rect -80 4771 -52 4799
rect -14 4771 14 4799
rect 52 4771 80 4799
rect 118 4771 146 4799
rect 184 4771 212 4799
rect 250 4771 278 4799
rect 316 4771 344 4799
rect -344 4705 -316 4733
rect -278 4705 -250 4733
rect -212 4705 -184 4733
rect -146 4705 -118 4733
rect -80 4705 -52 4733
rect -14 4705 14 4733
rect 52 4705 80 4733
rect 118 4705 146 4733
rect 184 4705 212 4733
rect 250 4705 278 4733
rect 316 4705 344 4733
rect -344 4639 -316 4667
rect -278 4639 -250 4667
rect -212 4639 -184 4667
rect -146 4639 -118 4667
rect -80 4639 -52 4667
rect -14 4639 14 4667
rect 52 4639 80 4667
rect 118 4639 146 4667
rect 184 4639 212 4667
rect 250 4639 278 4667
rect 316 4639 344 4667
rect -344 4573 -316 4601
rect -278 4573 -250 4601
rect -212 4573 -184 4601
rect -146 4573 -118 4601
rect -80 4573 -52 4601
rect -14 4573 14 4601
rect 52 4573 80 4601
rect 118 4573 146 4601
rect 184 4573 212 4601
rect 250 4573 278 4601
rect 316 4573 344 4601
rect -344 4507 -316 4535
rect -278 4507 -250 4535
rect -212 4507 -184 4535
rect -146 4507 -118 4535
rect -80 4507 -52 4535
rect -14 4507 14 4535
rect 52 4507 80 4535
rect 118 4507 146 4535
rect 184 4507 212 4535
rect 250 4507 278 4535
rect 316 4507 344 4535
rect -344 4441 -316 4469
rect -278 4441 -250 4469
rect -212 4441 -184 4469
rect -146 4441 -118 4469
rect -80 4441 -52 4469
rect -14 4441 14 4469
rect 52 4441 80 4469
rect 118 4441 146 4469
rect 184 4441 212 4469
rect 250 4441 278 4469
rect 316 4441 344 4469
rect -344 4375 -316 4403
rect -278 4375 -250 4403
rect -212 4375 -184 4403
rect -146 4375 -118 4403
rect -80 4375 -52 4403
rect -14 4375 14 4403
rect 52 4375 80 4403
rect 118 4375 146 4403
rect 184 4375 212 4403
rect 250 4375 278 4403
rect 316 4375 344 4403
rect -344 4309 -316 4337
rect -278 4309 -250 4337
rect -212 4309 -184 4337
rect -146 4309 -118 4337
rect -80 4309 -52 4337
rect -14 4309 14 4337
rect 52 4309 80 4337
rect 118 4309 146 4337
rect 184 4309 212 4337
rect 250 4309 278 4337
rect 316 4309 344 4337
rect -344 4243 -316 4271
rect -278 4243 -250 4271
rect -212 4243 -184 4271
rect -146 4243 -118 4271
rect -80 4243 -52 4271
rect -14 4243 14 4271
rect 52 4243 80 4271
rect 118 4243 146 4271
rect 184 4243 212 4271
rect 250 4243 278 4271
rect 316 4243 344 4271
rect -344 4177 -316 4205
rect -278 4177 -250 4205
rect -212 4177 -184 4205
rect -146 4177 -118 4205
rect -80 4177 -52 4205
rect -14 4177 14 4205
rect 52 4177 80 4205
rect 118 4177 146 4205
rect 184 4177 212 4205
rect 250 4177 278 4205
rect 316 4177 344 4205
rect -344 4111 -316 4139
rect -278 4111 -250 4139
rect -212 4111 -184 4139
rect -146 4111 -118 4139
rect -80 4111 -52 4139
rect -14 4111 14 4139
rect 52 4111 80 4139
rect 118 4111 146 4139
rect 184 4111 212 4139
rect 250 4111 278 4139
rect 316 4111 344 4139
rect -344 4045 -316 4073
rect -278 4045 -250 4073
rect -212 4045 -184 4073
rect -146 4045 -118 4073
rect -80 4045 -52 4073
rect -14 4045 14 4073
rect 52 4045 80 4073
rect 118 4045 146 4073
rect 184 4045 212 4073
rect 250 4045 278 4073
rect 316 4045 344 4073
rect -344 3979 -316 4007
rect -278 3979 -250 4007
rect -212 3979 -184 4007
rect -146 3979 -118 4007
rect -80 3979 -52 4007
rect -14 3979 14 4007
rect 52 3979 80 4007
rect 118 3979 146 4007
rect 184 3979 212 4007
rect 250 3979 278 4007
rect 316 3979 344 4007
rect -344 3913 -316 3941
rect -278 3913 -250 3941
rect -212 3913 -184 3941
rect -146 3913 -118 3941
rect -80 3913 -52 3941
rect -14 3913 14 3941
rect 52 3913 80 3941
rect 118 3913 146 3941
rect 184 3913 212 3941
rect 250 3913 278 3941
rect 316 3913 344 3941
rect -344 3847 -316 3875
rect -278 3847 -250 3875
rect -212 3847 -184 3875
rect -146 3847 -118 3875
rect -80 3847 -52 3875
rect -14 3847 14 3875
rect 52 3847 80 3875
rect 118 3847 146 3875
rect 184 3847 212 3875
rect 250 3847 278 3875
rect 316 3847 344 3875
rect -344 3781 -316 3809
rect -278 3781 -250 3809
rect -212 3781 -184 3809
rect -146 3781 -118 3809
rect -80 3781 -52 3809
rect -14 3781 14 3809
rect 52 3781 80 3809
rect 118 3781 146 3809
rect 184 3781 212 3809
rect 250 3781 278 3809
rect 316 3781 344 3809
rect -344 3715 -316 3743
rect -278 3715 -250 3743
rect -212 3715 -184 3743
rect -146 3715 -118 3743
rect -80 3715 -52 3743
rect -14 3715 14 3743
rect 52 3715 80 3743
rect 118 3715 146 3743
rect 184 3715 212 3743
rect 250 3715 278 3743
rect 316 3715 344 3743
rect -344 3649 -316 3677
rect -278 3649 -250 3677
rect -212 3649 -184 3677
rect -146 3649 -118 3677
rect -80 3649 -52 3677
rect -14 3649 14 3677
rect 52 3649 80 3677
rect 118 3649 146 3677
rect 184 3649 212 3677
rect 250 3649 278 3677
rect 316 3649 344 3677
rect -344 3583 -316 3611
rect -278 3583 -250 3611
rect -212 3583 -184 3611
rect -146 3583 -118 3611
rect -80 3583 -52 3611
rect -14 3583 14 3611
rect 52 3583 80 3611
rect 118 3583 146 3611
rect 184 3583 212 3611
rect 250 3583 278 3611
rect 316 3583 344 3611
rect -344 3517 -316 3545
rect -278 3517 -250 3545
rect -212 3517 -184 3545
rect -146 3517 -118 3545
rect -80 3517 -52 3545
rect -14 3517 14 3545
rect 52 3517 80 3545
rect 118 3517 146 3545
rect 184 3517 212 3545
rect 250 3517 278 3545
rect 316 3517 344 3545
rect -344 3451 -316 3479
rect -278 3451 -250 3479
rect -212 3451 -184 3479
rect -146 3451 -118 3479
rect -80 3451 -52 3479
rect -14 3451 14 3479
rect 52 3451 80 3479
rect 118 3451 146 3479
rect 184 3451 212 3479
rect 250 3451 278 3479
rect 316 3451 344 3479
rect -344 3385 -316 3413
rect -278 3385 -250 3413
rect -212 3385 -184 3413
rect -146 3385 -118 3413
rect -80 3385 -52 3413
rect -14 3385 14 3413
rect 52 3385 80 3413
rect 118 3385 146 3413
rect 184 3385 212 3413
rect 250 3385 278 3413
rect 316 3385 344 3413
rect -344 3319 -316 3347
rect -278 3319 -250 3347
rect -212 3319 -184 3347
rect -146 3319 -118 3347
rect -80 3319 -52 3347
rect -14 3319 14 3347
rect 52 3319 80 3347
rect 118 3319 146 3347
rect 184 3319 212 3347
rect 250 3319 278 3347
rect 316 3319 344 3347
rect -344 3253 -316 3281
rect -278 3253 -250 3281
rect -212 3253 -184 3281
rect -146 3253 -118 3281
rect -80 3253 -52 3281
rect -14 3253 14 3281
rect 52 3253 80 3281
rect 118 3253 146 3281
rect 184 3253 212 3281
rect 250 3253 278 3281
rect 316 3253 344 3281
rect -344 3187 -316 3215
rect -278 3187 -250 3215
rect -212 3187 -184 3215
rect -146 3187 -118 3215
rect -80 3187 -52 3215
rect -14 3187 14 3215
rect 52 3187 80 3215
rect 118 3187 146 3215
rect 184 3187 212 3215
rect 250 3187 278 3215
rect 316 3187 344 3215
rect -344 3121 -316 3149
rect -278 3121 -250 3149
rect -212 3121 -184 3149
rect -146 3121 -118 3149
rect -80 3121 -52 3149
rect -14 3121 14 3149
rect 52 3121 80 3149
rect 118 3121 146 3149
rect 184 3121 212 3149
rect 250 3121 278 3149
rect 316 3121 344 3149
rect -344 3055 -316 3083
rect -278 3055 -250 3083
rect -212 3055 -184 3083
rect -146 3055 -118 3083
rect -80 3055 -52 3083
rect -14 3055 14 3083
rect 52 3055 80 3083
rect 118 3055 146 3083
rect 184 3055 212 3083
rect 250 3055 278 3083
rect 316 3055 344 3083
rect -344 2989 -316 3017
rect -278 2989 -250 3017
rect -212 2989 -184 3017
rect -146 2989 -118 3017
rect -80 2989 -52 3017
rect -14 2989 14 3017
rect 52 2989 80 3017
rect 118 2989 146 3017
rect 184 2989 212 3017
rect 250 2989 278 3017
rect 316 2989 344 3017
rect -344 2923 -316 2951
rect -278 2923 -250 2951
rect -212 2923 -184 2951
rect -146 2923 -118 2951
rect -80 2923 -52 2951
rect -14 2923 14 2951
rect 52 2923 80 2951
rect 118 2923 146 2951
rect 184 2923 212 2951
rect 250 2923 278 2951
rect 316 2923 344 2951
rect -344 2857 -316 2885
rect -278 2857 -250 2885
rect -212 2857 -184 2885
rect -146 2857 -118 2885
rect -80 2857 -52 2885
rect -14 2857 14 2885
rect 52 2857 80 2885
rect 118 2857 146 2885
rect 184 2857 212 2885
rect 250 2857 278 2885
rect 316 2857 344 2885
rect -344 2791 -316 2819
rect -278 2791 -250 2819
rect -212 2791 -184 2819
rect -146 2791 -118 2819
rect -80 2791 -52 2819
rect -14 2791 14 2819
rect 52 2791 80 2819
rect 118 2791 146 2819
rect 184 2791 212 2819
rect 250 2791 278 2819
rect 316 2791 344 2819
rect -344 2725 -316 2753
rect -278 2725 -250 2753
rect -212 2725 -184 2753
rect -146 2725 -118 2753
rect -80 2725 -52 2753
rect -14 2725 14 2753
rect 52 2725 80 2753
rect 118 2725 146 2753
rect 184 2725 212 2753
rect 250 2725 278 2753
rect 316 2725 344 2753
rect -344 2659 -316 2687
rect -278 2659 -250 2687
rect -212 2659 -184 2687
rect -146 2659 -118 2687
rect -80 2659 -52 2687
rect -14 2659 14 2687
rect 52 2659 80 2687
rect 118 2659 146 2687
rect 184 2659 212 2687
rect 250 2659 278 2687
rect 316 2659 344 2687
rect -344 2593 -316 2621
rect -278 2593 -250 2621
rect -212 2593 -184 2621
rect -146 2593 -118 2621
rect -80 2593 -52 2621
rect -14 2593 14 2621
rect 52 2593 80 2621
rect 118 2593 146 2621
rect 184 2593 212 2621
rect 250 2593 278 2621
rect 316 2593 344 2621
rect -344 2527 -316 2555
rect -278 2527 -250 2555
rect -212 2527 -184 2555
rect -146 2527 -118 2555
rect -80 2527 -52 2555
rect -14 2527 14 2555
rect 52 2527 80 2555
rect 118 2527 146 2555
rect 184 2527 212 2555
rect 250 2527 278 2555
rect 316 2527 344 2555
rect -344 2461 -316 2489
rect -278 2461 -250 2489
rect -212 2461 -184 2489
rect -146 2461 -118 2489
rect -80 2461 -52 2489
rect -14 2461 14 2489
rect 52 2461 80 2489
rect 118 2461 146 2489
rect 184 2461 212 2489
rect 250 2461 278 2489
rect 316 2461 344 2489
rect -344 2395 -316 2423
rect -278 2395 -250 2423
rect -212 2395 -184 2423
rect -146 2395 -118 2423
rect -80 2395 -52 2423
rect -14 2395 14 2423
rect 52 2395 80 2423
rect 118 2395 146 2423
rect 184 2395 212 2423
rect 250 2395 278 2423
rect 316 2395 344 2423
rect -344 2329 -316 2357
rect -278 2329 -250 2357
rect -212 2329 -184 2357
rect -146 2329 -118 2357
rect -80 2329 -52 2357
rect -14 2329 14 2357
rect 52 2329 80 2357
rect 118 2329 146 2357
rect 184 2329 212 2357
rect 250 2329 278 2357
rect 316 2329 344 2357
rect -344 2263 -316 2291
rect -278 2263 -250 2291
rect -212 2263 -184 2291
rect -146 2263 -118 2291
rect -80 2263 -52 2291
rect -14 2263 14 2291
rect 52 2263 80 2291
rect 118 2263 146 2291
rect 184 2263 212 2291
rect 250 2263 278 2291
rect 316 2263 344 2291
rect -344 2197 -316 2225
rect -278 2197 -250 2225
rect -212 2197 -184 2225
rect -146 2197 -118 2225
rect -80 2197 -52 2225
rect -14 2197 14 2225
rect 52 2197 80 2225
rect 118 2197 146 2225
rect 184 2197 212 2225
rect 250 2197 278 2225
rect 316 2197 344 2225
rect -344 2131 -316 2159
rect -278 2131 -250 2159
rect -212 2131 -184 2159
rect -146 2131 -118 2159
rect -80 2131 -52 2159
rect -14 2131 14 2159
rect 52 2131 80 2159
rect 118 2131 146 2159
rect 184 2131 212 2159
rect 250 2131 278 2159
rect 316 2131 344 2159
rect -344 2065 -316 2093
rect -278 2065 -250 2093
rect -212 2065 -184 2093
rect -146 2065 -118 2093
rect -80 2065 -52 2093
rect -14 2065 14 2093
rect 52 2065 80 2093
rect 118 2065 146 2093
rect 184 2065 212 2093
rect 250 2065 278 2093
rect 316 2065 344 2093
rect -344 1999 -316 2027
rect -278 1999 -250 2027
rect -212 1999 -184 2027
rect -146 1999 -118 2027
rect -80 1999 -52 2027
rect -14 1999 14 2027
rect 52 1999 80 2027
rect 118 1999 146 2027
rect 184 1999 212 2027
rect 250 1999 278 2027
rect 316 1999 344 2027
rect -344 1933 -316 1961
rect -278 1933 -250 1961
rect -212 1933 -184 1961
rect -146 1933 -118 1961
rect -80 1933 -52 1961
rect -14 1933 14 1961
rect 52 1933 80 1961
rect 118 1933 146 1961
rect 184 1933 212 1961
rect 250 1933 278 1961
rect 316 1933 344 1961
rect -344 1867 -316 1895
rect -278 1867 -250 1895
rect -212 1867 -184 1895
rect -146 1867 -118 1895
rect -80 1867 -52 1895
rect -14 1867 14 1895
rect 52 1867 80 1895
rect 118 1867 146 1895
rect 184 1867 212 1895
rect 250 1867 278 1895
rect 316 1867 344 1895
rect -344 1801 -316 1829
rect -278 1801 -250 1829
rect -212 1801 -184 1829
rect -146 1801 -118 1829
rect -80 1801 -52 1829
rect -14 1801 14 1829
rect 52 1801 80 1829
rect 118 1801 146 1829
rect 184 1801 212 1829
rect 250 1801 278 1829
rect 316 1801 344 1829
rect -344 1735 -316 1763
rect -278 1735 -250 1763
rect -212 1735 -184 1763
rect -146 1735 -118 1763
rect -80 1735 -52 1763
rect -14 1735 14 1763
rect 52 1735 80 1763
rect 118 1735 146 1763
rect 184 1735 212 1763
rect 250 1735 278 1763
rect 316 1735 344 1763
rect -344 1669 -316 1697
rect -278 1669 -250 1697
rect -212 1669 -184 1697
rect -146 1669 -118 1697
rect -80 1669 -52 1697
rect -14 1669 14 1697
rect 52 1669 80 1697
rect 118 1669 146 1697
rect 184 1669 212 1697
rect 250 1669 278 1697
rect 316 1669 344 1697
rect -344 1603 -316 1631
rect -278 1603 -250 1631
rect -212 1603 -184 1631
rect -146 1603 -118 1631
rect -80 1603 -52 1631
rect -14 1603 14 1631
rect 52 1603 80 1631
rect 118 1603 146 1631
rect 184 1603 212 1631
rect 250 1603 278 1631
rect 316 1603 344 1631
rect -344 1537 -316 1565
rect -278 1537 -250 1565
rect -212 1537 -184 1565
rect -146 1537 -118 1565
rect -80 1537 -52 1565
rect -14 1537 14 1565
rect 52 1537 80 1565
rect 118 1537 146 1565
rect 184 1537 212 1565
rect 250 1537 278 1565
rect 316 1537 344 1565
rect -344 1471 -316 1499
rect -278 1471 -250 1499
rect -212 1471 -184 1499
rect -146 1471 -118 1499
rect -80 1471 -52 1499
rect -14 1471 14 1499
rect 52 1471 80 1499
rect 118 1471 146 1499
rect 184 1471 212 1499
rect 250 1471 278 1499
rect 316 1471 344 1499
rect -344 1405 -316 1433
rect -278 1405 -250 1433
rect -212 1405 -184 1433
rect -146 1405 -118 1433
rect -80 1405 -52 1433
rect -14 1405 14 1433
rect 52 1405 80 1433
rect 118 1405 146 1433
rect 184 1405 212 1433
rect 250 1405 278 1433
rect 316 1405 344 1433
rect -344 1339 -316 1367
rect -278 1339 -250 1367
rect -212 1339 -184 1367
rect -146 1339 -118 1367
rect -80 1339 -52 1367
rect -14 1339 14 1367
rect 52 1339 80 1367
rect 118 1339 146 1367
rect 184 1339 212 1367
rect 250 1339 278 1367
rect 316 1339 344 1367
rect -344 1273 -316 1301
rect -278 1273 -250 1301
rect -212 1273 -184 1301
rect -146 1273 -118 1301
rect -80 1273 -52 1301
rect -14 1273 14 1301
rect 52 1273 80 1301
rect 118 1273 146 1301
rect 184 1273 212 1301
rect 250 1273 278 1301
rect 316 1273 344 1301
rect -344 1207 -316 1235
rect -278 1207 -250 1235
rect -212 1207 -184 1235
rect -146 1207 -118 1235
rect -80 1207 -52 1235
rect -14 1207 14 1235
rect 52 1207 80 1235
rect 118 1207 146 1235
rect 184 1207 212 1235
rect 250 1207 278 1235
rect 316 1207 344 1235
rect -344 1141 -316 1169
rect -278 1141 -250 1169
rect -212 1141 -184 1169
rect -146 1141 -118 1169
rect -80 1141 -52 1169
rect -14 1141 14 1169
rect 52 1141 80 1169
rect 118 1141 146 1169
rect 184 1141 212 1169
rect 250 1141 278 1169
rect 316 1141 344 1169
rect -344 1075 -316 1103
rect -278 1075 -250 1103
rect -212 1075 -184 1103
rect -146 1075 -118 1103
rect -80 1075 -52 1103
rect -14 1075 14 1103
rect 52 1075 80 1103
rect 118 1075 146 1103
rect 184 1075 212 1103
rect 250 1075 278 1103
rect 316 1075 344 1103
rect -344 1009 -316 1037
rect -278 1009 -250 1037
rect -212 1009 -184 1037
rect -146 1009 -118 1037
rect -80 1009 -52 1037
rect -14 1009 14 1037
rect 52 1009 80 1037
rect 118 1009 146 1037
rect 184 1009 212 1037
rect 250 1009 278 1037
rect 316 1009 344 1037
rect -344 943 -316 971
rect -278 943 -250 971
rect -212 943 -184 971
rect -146 943 -118 971
rect -80 943 -52 971
rect -14 943 14 971
rect 52 943 80 971
rect 118 943 146 971
rect 184 943 212 971
rect 250 943 278 971
rect 316 943 344 971
rect -344 877 -316 905
rect -278 877 -250 905
rect -212 877 -184 905
rect -146 877 -118 905
rect -80 877 -52 905
rect -14 877 14 905
rect 52 877 80 905
rect 118 877 146 905
rect 184 877 212 905
rect 250 877 278 905
rect 316 877 344 905
rect -344 811 -316 839
rect -278 811 -250 839
rect -212 811 -184 839
rect -146 811 -118 839
rect -80 811 -52 839
rect -14 811 14 839
rect 52 811 80 839
rect 118 811 146 839
rect 184 811 212 839
rect 250 811 278 839
rect 316 811 344 839
rect -344 745 -316 773
rect -278 745 -250 773
rect -212 745 -184 773
rect -146 745 -118 773
rect -80 745 -52 773
rect -14 745 14 773
rect 52 745 80 773
rect 118 745 146 773
rect 184 745 212 773
rect 250 745 278 773
rect 316 745 344 773
rect -344 679 -316 707
rect -278 679 -250 707
rect -212 679 -184 707
rect -146 679 -118 707
rect -80 679 -52 707
rect -14 679 14 707
rect 52 679 80 707
rect 118 679 146 707
rect 184 679 212 707
rect 250 679 278 707
rect 316 679 344 707
rect -344 613 -316 641
rect -278 613 -250 641
rect -212 613 -184 641
rect -146 613 -118 641
rect -80 613 -52 641
rect -14 613 14 641
rect 52 613 80 641
rect 118 613 146 641
rect 184 613 212 641
rect 250 613 278 641
rect 316 613 344 641
rect -344 547 -316 575
rect -278 547 -250 575
rect -212 547 -184 575
rect -146 547 -118 575
rect -80 547 -52 575
rect -14 547 14 575
rect 52 547 80 575
rect 118 547 146 575
rect 184 547 212 575
rect 250 547 278 575
rect 316 547 344 575
rect -344 481 -316 509
rect -278 481 -250 509
rect -212 481 -184 509
rect -146 481 -118 509
rect -80 481 -52 509
rect -14 481 14 509
rect 52 481 80 509
rect 118 481 146 509
rect 184 481 212 509
rect 250 481 278 509
rect 316 481 344 509
rect -344 415 -316 443
rect -278 415 -250 443
rect -212 415 -184 443
rect -146 415 -118 443
rect -80 415 -52 443
rect -14 415 14 443
rect 52 415 80 443
rect 118 415 146 443
rect 184 415 212 443
rect 250 415 278 443
rect 316 415 344 443
rect -344 349 -316 377
rect -278 349 -250 377
rect -212 349 -184 377
rect -146 349 -118 377
rect -80 349 -52 377
rect -14 349 14 377
rect 52 349 80 377
rect 118 349 146 377
rect 184 349 212 377
rect 250 349 278 377
rect 316 349 344 377
rect -344 283 -316 311
rect -278 283 -250 311
rect -212 283 -184 311
rect -146 283 -118 311
rect -80 283 -52 311
rect -14 283 14 311
rect 52 283 80 311
rect 118 283 146 311
rect 184 283 212 311
rect 250 283 278 311
rect 316 283 344 311
rect -344 217 -316 245
rect -278 217 -250 245
rect -212 217 -184 245
rect -146 217 -118 245
rect -80 217 -52 245
rect -14 217 14 245
rect 52 217 80 245
rect 118 217 146 245
rect 184 217 212 245
rect 250 217 278 245
rect 316 217 344 245
rect -344 151 -316 179
rect -278 151 -250 179
rect -212 151 -184 179
rect -146 151 -118 179
rect -80 151 -52 179
rect -14 151 14 179
rect 52 151 80 179
rect 118 151 146 179
rect 184 151 212 179
rect 250 151 278 179
rect 316 151 344 179
rect -344 85 -316 113
rect -278 85 -250 113
rect -212 85 -184 113
rect -146 85 -118 113
rect -80 85 -52 113
rect -14 85 14 113
rect 52 85 80 113
rect 118 85 146 113
rect 184 85 212 113
rect 250 85 278 113
rect 316 85 344 113
rect -344 19 -316 47
rect -278 19 -250 47
rect -212 19 -184 47
rect -146 19 -118 47
rect -80 19 -52 47
rect -14 19 14 47
rect 52 19 80 47
rect 118 19 146 47
rect 184 19 212 47
rect 250 19 278 47
rect 316 19 344 47
rect -344 -47 -316 -19
rect -278 -47 -250 -19
rect -212 -47 -184 -19
rect -146 -47 -118 -19
rect -80 -47 -52 -19
rect -14 -47 14 -19
rect 52 -47 80 -19
rect 118 -47 146 -19
rect 184 -47 212 -19
rect 250 -47 278 -19
rect 316 -47 344 -19
rect -344 -113 -316 -85
rect -278 -113 -250 -85
rect -212 -113 -184 -85
rect -146 -113 -118 -85
rect -80 -113 -52 -85
rect -14 -113 14 -85
rect 52 -113 80 -85
rect 118 -113 146 -85
rect 184 -113 212 -85
rect 250 -113 278 -85
rect 316 -113 344 -85
rect -344 -179 -316 -151
rect -278 -179 -250 -151
rect -212 -179 -184 -151
rect -146 -179 -118 -151
rect -80 -179 -52 -151
rect -14 -179 14 -151
rect 52 -179 80 -151
rect 118 -179 146 -151
rect 184 -179 212 -151
rect 250 -179 278 -151
rect 316 -179 344 -151
rect -344 -245 -316 -217
rect -278 -245 -250 -217
rect -212 -245 -184 -217
rect -146 -245 -118 -217
rect -80 -245 -52 -217
rect -14 -245 14 -217
rect 52 -245 80 -217
rect 118 -245 146 -217
rect 184 -245 212 -217
rect 250 -245 278 -217
rect 316 -245 344 -217
rect -344 -311 -316 -283
rect -278 -311 -250 -283
rect -212 -311 -184 -283
rect -146 -311 -118 -283
rect -80 -311 -52 -283
rect -14 -311 14 -283
rect 52 -311 80 -283
rect 118 -311 146 -283
rect 184 -311 212 -283
rect 250 -311 278 -283
rect 316 -311 344 -283
rect -344 -377 -316 -349
rect -278 -377 -250 -349
rect -212 -377 -184 -349
rect -146 -377 -118 -349
rect -80 -377 -52 -349
rect -14 -377 14 -349
rect 52 -377 80 -349
rect 118 -377 146 -349
rect 184 -377 212 -349
rect 250 -377 278 -349
rect 316 -377 344 -349
rect -344 -443 -316 -415
rect -278 -443 -250 -415
rect -212 -443 -184 -415
rect -146 -443 -118 -415
rect -80 -443 -52 -415
rect -14 -443 14 -415
rect 52 -443 80 -415
rect 118 -443 146 -415
rect 184 -443 212 -415
rect 250 -443 278 -415
rect 316 -443 344 -415
rect -344 -509 -316 -481
rect -278 -509 -250 -481
rect -212 -509 -184 -481
rect -146 -509 -118 -481
rect -80 -509 -52 -481
rect -14 -509 14 -481
rect 52 -509 80 -481
rect 118 -509 146 -481
rect 184 -509 212 -481
rect 250 -509 278 -481
rect 316 -509 344 -481
rect -344 -575 -316 -547
rect -278 -575 -250 -547
rect -212 -575 -184 -547
rect -146 -575 -118 -547
rect -80 -575 -52 -547
rect -14 -575 14 -547
rect 52 -575 80 -547
rect 118 -575 146 -547
rect 184 -575 212 -547
rect 250 -575 278 -547
rect 316 -575 344 -547
rect -344 -641 -316 -613
rect -278 -641 -250 -613
rect -212 -641 -184 -613
rect -146 -641 -118 -613
rect -80 -641 -52 -613
rect -14 -641 14 -613
rect 52 -641 80 -613
rect 118 -641 146 -613
rect 184 -641 212 -613
rect 250 -641 278 -613
rect 316 -641 344 -613
rect -344 -707 -316 -679
rect -278 -707 -250 -679
rect -212 -707 -184 -679
rect -146 -707 -118 -679
rect -80 -707 -52 -679
rect -14 -707 14 -679
rect 52 -707 80 -679
rect 118 -707 146 -679
rect 184 -707 212 -679
rect 250 -707 278 -679
rect 316 -707 344 -679
rect -344 -773 -316 -745
rect -278 -773 -250 -745
rect -212 -773 -184 -745
rect -146 -773 -118 -745
rect -80 -773 -52 -745
rect -14 -773 14 -745
rect 52 -773 80 -745
rect 118 -773 146 -745
rect 184 -773 212 -745
rect 250 -773 278 -745
rect 316 -773 344 -745
rect -344 -839 -316 -811
rect -278 -839 -250 -811
rect -212 -839 -184 -811
rect -146 -839 -118 -811
rect -80 -839 -52 -811
rect -14 -839 14 -811
rect 52 -839 80 -811
rect 118 -839 146 -811
rect 184 -839 212 -811
rect 250 -839 278 -811
rect 316 -839 344 -811
rect -344 -905 -316 -877
rect -278 -905 -250 -877
rect -212 -905 -184 -877
rect -146 -905 -118 -877
rect -80 -905 -52 -877
rect -14 -905 14 -877
rect 52 -905 80 -877
rect 118 -905 146 -877
rect 184 -905 212 -877
rect 250 -905 278 -877
rect 316 -905 344 -877
rect -344 -971 -316 -943
rect -278 -971 -250 -943
rect -212 -971 -184 -943
rect -146 -971 -118 -943
rect -80 -971 -52 -943
rect -14 -971 14 -943
rect 52 -971 80 -943
rect 118 -971 146 -943
rect 184 -971 212 -943
rect 250 -971 278 -943
rect 316 -971 344 -943
rect -344 -1037 -316 -1009
rect -278 -1037 -250 -1009
rect -212 -1037 -184 -1009
rect -146 -1037 -118 -1009
rect -80 -1037 -52 -1009
rect -14 -1037 14 -1009
rect 52 -1037 80 -1009
rect 118 -1037 146 -1009
rect 184 -1037 212 -1009
rect 250 -1037 278 -1009
rect 316 -1037 344 -1009
rect -344 -1103 -316 -1075
rect -278 -1103 -250 -1075
rect -212 -1103 -184 -1075
rect -146 -1103 -118 -1075
rect -80 -1103 -52 -1075
rect -14 -1103 14 -1075
rect 52 -1103 80 -1075
rect 118 -1103 146 -1075
rect 184 -1103 212 -1075
rect 250 -1103 278 -1075
rect 316 -1103 344 -1075
rect -344 -1169 -316 -1141
rect -278 -1169 -250 -1141
rect -212 -1169 -184 -1141
rect -146 -1169 -118 -1141
rect -80 -1169 -52 -1141
rect -14 -1169 14 -1141
rect 52 -1169 80 -1141
rect 118 -1169 146 -1141
rect 184 -1169 212 -1141
rect 250 -1169 278 -1141
rect 316 -1169 344 -1141
rect -344 -1235 -316 -1207
rect -278 -1235 -250 -1207
rect -212 -1235 -184 -1207
rect -146 -1235 -118 -1207
rect -80 -1235 -52 -1207
rect -14 -1235 14 -1207
rect 52 -1235 80 -1207
rect 118 -1235 146 -1207
rect 184 -1235 212 -1207
rect 250 -1235 278 -1207
rect 316 -1235 344 -1207
rect -344 -1301 -316 -1273
rect -278 -1301 -250 -1273
rect -212 -1301 -184 -1273
rect -146 -1301 -118 -1273
rect -80 -1301 -52 -1273
rect -14 -1301 14 -1273
rect 52 -1301 80 -1273
rect 118 -1301 146 -1273
rect 184 -1301 212 -1273
rect 250 -1301 278 -1273
rect 316 -1301 344 -1273
rect -344 -1367 -316 -1339
rect -278 -1367 -250 -1339
rect -212 -1367 -184 -1339
rect -146 -1367 -118 -1339
rect -80 -1367 -52 -1339
rect -14 -1367 14 -1339
rect 52 -1367 80 -1339
rect 118 -1367 146 -1339
rect 184 -1367 212 -1339
rect 250 -1367 278 -1339
rect 316 -1367 344 -1339
rect -344 -1433 -316 -1405
rect -278 -1433 -250 -1405
rect -212 -1433 -184 -1405
rect -146 -1433 -118 -1405
rect -80 -1433 -52 -1405
rect -14 -1433 14 -1405
rect 52 -1433 80 -1405
rect 118 -1433 146 -1405
rect 184 -1433 212 -1405
rect 250 -1433 278 -1405
rect 316 -1433 344 -1405
rect -344 -1499 -316 -1471
rect -278 -1499 -250 -1471
rect -212 -1499 -184 -1471
rect -146 -1499 -118 -1471
rect -80 -1499 -52 -1471
rect -14 -1499 14 -1471
rect 52 -1499 80 -1471
rect 118 -1499 146 -1471
rect 184 -1499 212 -1471
rect 250 -1499 278 -1471
rect 316 -1499 344 -1471
rect -344 -1565 -316 -1537
rect -278 -1565 -250 -1537
rect -212 -1565 -184 -1537
rect -146 -1565 -118 -1537
rect -80 -1565 -52 -1537
rect -14 -1565 14 -1537
rect 52 -1565 80 -1537
rect 118 -1565 146 -1537
rect 184 -1565 212 -1537
rect 250 -1565 278 -1537
rect 316 -1565 344 -1537
rect -344 -1631 -316 -1603
rect -278 -1631 -250 -1603
rect -212 -1631 -184 -1603
rect -146 -1631 -118 -1603
rect -80 -1631 -52 -1603
rect -14 -1631 14 -1603
rect 52 -1631 80 -1603
rect 118 -1631 146 -1603
rect 184 -1631 212 -1603
rect 250 -1631 278 -1603
rect 316 -1631 344 -1603
rect -344 -1697 -316 -1669
rect -278 -1697 -250 -1669
rect -212 -1697 -184 -1669
rect -146 -1697 -118 -1669
rect -80 -1697 -52 -1669
rect -14 -1697 14 -1669
rect 52 -1697 80 -1669
rect 118 -1697 146 -1669
rect 184 -1697 212 -1669
rect 250 -1697 278 -1669
rect 316 -1697 344 -1669
rect -344 -1763 -316 -1735
rect -278 -1763 -250 -1735
rect -212 -1763 -184 -1735
rect -146 -1763 -118 -1735
rect -80 -1763 -52 -1735
rect -14 -1763 14 -1735
rect 52 -1763 80 -1735
rect 118 -1763 146 -1735
rect 184 -1763 212 -1735
rect 250 -1763 278 -1735
rect 316 -1763 344 -1735
rect -344 -1829 -316 -1801
rect -278 -1829 -250 -1801
rect -212 -1829 -184 -1801
rect -146 -1829 -118 -1801
rect -80 -1829 -52 -1801
rect -14 -1829 14 -1801
rect 52 -1829 80 -1801
rect 118 -1829 146 -1801
rect 184 -1829 212 -1801
rect 250 -1829 278 -1801
rect 316 -1829 344 -1801
rect -344 -1895 -316 -1867
rect -278 -1895 -250 -1867
rect -212 -1895 -184 -1867
rect -146 -1895 -118 -1867
rect -80 -1895 -52 -1867
rect -14 -1895 14 -1867
rect 52 -1895 80 -1867
rect 118 -1895 146 -1867
rect 184 -1895 212 -1867
rect 250 -1895 278 -1867
rect 316 -1895 344 -1867
rect -344 -1961 -316 -1933
rect -278 -1961 -250 -1933
rect -212 -1961 -184 -1933
rect -146 -1961 -118 -1933
rect -80 -1961 -52 -1933
rect -14 -1961 14 -1933
rect 52 -1961 80 -1933
rect 118 -1961 146 -1933
rect 184 -1961 212 -1933
rect 250 -1961 278 -1933
rect 316 -1961 344 -1933
rect -344 -2027 -316 -1999
rect -278 -2027 -250 -1999
rect -212 -2027 -184 -1999
rect -146 -2027 -118 -1999
rect -80 -2027 -52 -1999
rect -14 -2027 14 -1999
rect 52 -2027 80 -1999
rect 118 -2027 146 -1999
rect 184 -2027 212 -1999
rect 250 -2027 278 -1999
rect 316 -2027 344 -1999
rect -344 -2093 -316 -2065
rect -278 -2093 -250 -2065
rect -212 -2093 -184 -2065
rect -146 -2093 -118 -2065
rect -80 -2093 -52 -2065
rect -14 -2093 14 -2065
rect 52 -2093 80 -2065
rect 118 -2093 146 -2065
rect 184 -2093 212 -2065
rect 250 -2093 278 -2065
rect 316 -2093 344 -2065
rect -344 -2159 -316 -2131
rect -278 -2159 -250 -2131
rect -212 -2159 -184 -2131
rect -146 -2159 -118 -2131
rect -80 -2159 -52 -2131
rect -14 -2159 14 -2131
rect 52 -2159 80 -2131
rect 118 -2159 146 -2131
rect 184 -2159 212 -2131
rect 250 -2159 278 -2131
rect 316 -2159 344 -2131
rect -344 -2225 -316 -2197
rect -278 -2225 -250 -2197
rect -212 -2225 -184 -2197
rect -146 -2225 -118 -2197
rect -80 -2225 -52 -2197
rect -14 -2225 14 -2197
rect 52 -2225 80 -2197
rect 118 -2225 146 -2197
rect 184 -2225 212 -2197
rect 250 -2225 278 -2197
rect 316 -2225 344 -2197
rect -344 -2291 -316 -2263
rect -278 -2291 -250 -2263
rect -212 -2291 -184 -2263
rect -146 -2291 -118 -2263
rect -80 -2291 -52 -2263
rect -14 -2291 14 -2263
rect 52 -2291 80 -2263
rect 118 -2291 146 -2263
rect 184 -2291 212 -2263
rect 250 -2291 278 -2263
rect 316 -2291 344 -2263
rect -344 -2357 -316 -2329
rect -278 -2357 -250 -2329
rect -212 -2357 -184 -2329
rect -146 -2357 -118 -2329
rect -80 -2357 -52 -2329
rect -14 -2357 14 -2329
rect 52 -2357 80 -2329
rect 118 -2357 146 -2329
rect 184 -2357 212 -2329
rect 250 -2357 278 -2329
rect 316 -2357 344 -2329
rect -344 -2423 -316 -2395
rect -278 -2423 -250 -2395
rect -212 -2423 -184 -2395
rect -146 -2423 -118 -2395
rect -80 -2423 -52 -2395
rect -14 -2423 14 -2395
rect 52 -2423 80 -2395
rect 118 -2423 146 -2395
rect 184 -2423 212 -2395
rect 250 -2423 278 -2395
rect 316 -2423 344 -2395
rect -344 -2489 -316 -2461
rect -278 -2489 -250 -2461
rect -212 -2489 -184 -2461
rect -146 -2489 -118 -2461
rect -80 -2489 -52 -2461
rect -14 -2489 14 -2461
rect 52 -2489 80 -2461
rect 118 -2489 146 -2461
rect 184 -2489 212 -2461
rect 250 -2489 278 -2461
rect 316 -2489 344 -2461
rect -344 -2555 -316 -2527
rect -278 -2555 -250 -2527
rect -212 -2555 -184 -2527
rect -146 -2555 -118 -2527
rect -80 -2555 -52 -2527
rect -14 -2555 14 -2527
rect 52 -2555 80 -2527
rect 118 -2555 146 -2527
rect 184 -2555 212 -2527
rect 250 -2555 278 -2527
rect 316 -2555 344 -2527
rect -344 -2621 -316 -2593
rect -278 -2621 -250 -2593
rect -212 -2621 -184 -2593
rect -146 -2621 -118 -2593
rect -80 -2621 -52 -2593
rect -14 -2621 14 -2593
rect 52 -2621 80 -2593
rect 118 -2621 146 -2593
rect 184 -2621 212 -2593
rect 250 -2621 278 -2593
rect 316 -2621 344 -2593
rect -344 -2687 -316 -2659
rect -278 -2687 -250 -2659
rect -212 -2687 -184 -2659
rect -146 -2687 -118 -2659
rect -80 -2687 -52 -2659
rect -14 -2687 14 -2659
rect 52 -2687 80 -2659
rect 118 -2687 146 -2659
rect 184 -2687 212 -2659
rect 250 -2687 278 -2659
rect 316 -2687 344 -2659
rect -344 -2753 -316 -2725
rect -278 -2753 -250 -2725
rect -212 -2753 -184 -2725
rect -146 -2753 -118 -2725
rect -80 -2753 -52 -2725
rect -14 -2753 14 -2725
rect 52 -2753 80 -2725
rect 118 -2753 146 -2725
rect 184 -2753 212 -2725
rect 250 -2753 278 -2725
rect 316 -2753 344 -2725
rect -344 -2819 -316 -2791
rect -278 -2819 -250 -2791
rect -212 -2819 -184 -2791
rect -146 -2819 -118 -2791
rect -80 -2819 -52 -2791
rect -14 -2819 14 -2791
rect 52 -2819 80 -2791
rect 118 -2819 146 -2791
rect 184 -2819 212 -2791
rect 250 -2819 278 -2791
rect 316 -2819 344 -2791
rect -344 -2885 -316 -2857
rect -278 -2885 -250 -2857
rect -212 -2885 -184 -2857
rect -146 -2885 -118 -2857
rect -80 -2885 -52 -2857
rect -14 -2885 14 -2857
rect 52 -2885 80 -2857
rect 118 -2885 146 -2857
rect 184 -2885 212 -2857
rect 250 -2885 278 -2857
rect 316 -2885 344 -2857
rect -344 -2951 -316 -2923
rect -278 -2951 -250 -2923
rect -212 -2951 -184 -2923
rect -146 -2951 -118 -2923
rect -80 -2951 -52 -2923
rect -14 -2951 14 -2923
rect 52 -2951 80 -2923
rect 118 -2951 146 -2923
rect 184 -2951 212 -2923
rect 250 -2951 278 -2923
rect 316 -2951 344 -2923
rect -344 -3017 -316 -2989
rect -278 -3017 -250 -2989
rect -212 -3017 -184 -2989
rect -146 -3017 -118 -2989
rect -80 -3017 -52 -2989
rect -14 -3017 14 -2989
rect 52 -3017 80 -2989
rect 118 -3017 146 -2989
rect 184 -3017 212 -2989
rect 250 -3017 278 -2989
rect 316 -3017 344 -2989
rect -344 -3083 -316 -3055
rect -278 -3083 -250 -3055
rect -212 -3083 -184 -3055
rect -146 -3083 -118 -3055
rect -80 -3083 -52 -3055
rect -14 -3083 14 -3055
rect 52 -3083 80 -3055
rect 118 -3083 146 -3055
rect 184 -3083 212 -3055
rect 250 -3083 278 -3055
rect 316 -3083 344 -3055
rect -344 -3149 -316 -3121
rect -278 -3149 -250 -3121
rect -212 -3149 -184 -3121
rect -146 -3149 -118 -3121
rect -80 -3149 -52 -3121
rect -14 -3149 14 -3121
rect 52 -3149 80 -3121
rect 118 -3149 146 -3121
rect 184 -3149 212 -3121
rect 250 -3149 278 -3121
rect 316 -3149 344 -3121
rect -344 -3215 -316 -3187
rect -278 -3215 -250 -3187
rect -212 -3215 -184 -3187
rect -146 -3215 -118 -3187
rect -80 -3215 -52 -3187
rect -14 -3215 14 -3187
rect 52 -3215 80 -3187
rect 118 -3215 146 -3187
rect 184 -3215 212 -3187
rect 250 -3215 278 -3187
rect 316 -3215 344 -3187
rect -344 -3281 -316 -3253
rect -278 -3281 -250 -3253
rect -212 -3281 -184 -3253
rect -146 -3281 -118 -3253
rect -80 -3281 -52 -3253
rect -14 -3281 14 -3253
rect 52 -3281 80 -3253
rect 118 -3281 146 -3253
rect 184 -3281 212 -3253
rect 250 -3281 278 -3253
rect 316 -3281 344 -3253
rect -344 -3347 -316 -3319
rect -278 -3347 -250 -3319
rect -212 -3347 -184 -3319
rect -146 -3347 -118 -3319
rect -80 -3347 -52 -3319
rect -14 -3347 14 -3319
rect 52 -3347 80 -3319
rect 118 -3347 146 -3319
rect 184 -3347 212 -3319
rect 250 -3347 278 -3319
rect 316 -3347 344 -3319
rect -344 -3413 -316 -3385
rect -278 -3413 -250 -3385
rect -212 -3413 -184 -3385
rect -146 -3413 -118 -3385
rect -80 -3413 -52 -3385
rect -14 -3413 14 -3385
rect 52 -3413 80 -3385
rect 118 -3413 146 -3385
rect 184 -3413 212 -3385
rect 250 -3413 278 -3385
rect 316 -3413 344 -3385
rect -344 -3479 -316 -3451
rect -278 -3479 -250 -3451
rect -212 -3479 -184 -3451
rect -146 -3479 -118 -3451
rect -80 -3479 -52 -3451
rect -14 -3479 14 -3451
rect 52 -3479 80 -3451
rect 118 -3479 146 -3451
rect 184 -3479 212 -3451
rect 250 -3479 278 -3451
rect 316 -3479 344 -3451
rect -344 -3545 -316 -3517
rect -278 -3545 -250 -3517
rect -212 -3545 -184 -3517
rect -146 -3545 -118 -3517
rect -80 -3545 -52 -3517
rect -14 -3545 14 -3517
rect 52 -3545 80 -3517
rect 118 -3545 146 -3517
rect 184 -3545 212 -3517
rect 250 -3545 278 -3517
rect 316 -3545 344 -3517
rect -344 -3611 -316 -3583
rect -278 -3611 -250 -3583
rect -212 -3611 -184 -3583
rect -146 -3611 -118 -3583
rect -80 -3611 -52 -3583
rect -14 -3611 14 -3583
rect 52 -3611 80 -3583
rect 118 -3611 146 -3583
rect 184 -3611 212 -3583
rect 250 -3611 278 -3583
rect 316 -3611 344 -3583
rect -344 -3677 -316 -3649
rect -278 -3677 -250 -3649
rect -212 -3677 -184 -3649
rect -146 -3677 -118 -3649
rect -80 -3677 -52 -3649
rect -14 -3677 14 -3649
rect 52 -3677 80 -3649
rect 118 -3677 146 -3649
rect 184 -3677 212 -3649
rect 250 -3677 278 -3649
rect 316 -3677 344 -3649
rect -344 -3743 -316 -3715
rect -278 -3743 -250 -3715
rect -212 -3743 -184 -3715
rect -146 -3743 -118 -3715
rect -80 -3743 -52 -3715
rect -14 -3743 14 -3715
rect 52 -3743 80 -3715
rect 118 -3743 146 -3715
rect 184 -3743 212 -3715
rect 250 -3743 278 -3715
rect 316 -3743 344 -3715
rect -344 -3809 -316 -3781
rect -278 -3809 -250 -3781
rect -212 -3809 -184 -3781
rect -146 -3809 -118 -3781
rect -80 -3809 -52 -3781
rect -14 -3809 14 -3781
rect 52 -3809 80 -3781
rect 118 -3809 146 -3781
rect 184 -3809 212 -3781
rect 250 -3809 278 -3781
rect 316 -3809 344 -3781
rect -344 -3875 -316 -3847
rect -278 -3875 -250 -3847
rect -212 -3875 -184 -3847
rect -146 -3875 -118 -3847
rect -80 -3875 -52 -3847
rect -14 -3875 14 -3847
rect 52 -3875 80 -3847
rect 118 -3875 146 -3847
rect 184 -3875 212 -3847
rect 250 -3875 278 -3847
rect 316 -3875 344 -3847
rect -344 -3941 -316 -3913
rect -278 -3941 -250 -3913
rect -212 -3941 -184 -3913
rect -146 -3941 -118 -3913
rect -80 -3941 -52 -3913
rect -14 -3941 14 -3913
rect 52 -3941 80 -3913
rect 118 -3941 146 -3913
rect 184 -3941 212 -3913
rect 250 -3941 278 -3913
rect 316 -3941 344 -3913
rect -344 -4007 -316 -3979
rect -278 -4007 -250 -3979
rect -212 -4007 -184 -3979
rect -146 -4007 -118 -3979
rect -80 -4007 -52 -3979
rect -14 -4007 14 -3979
rect 52 -4007 80 -3979
rect 118 -4007 146 -3979
rect 184 -4007 212 -3979
rect 250 -4007 278 -3979
rect 316 -4007 344 -3979
rect -344 -4073 -316 -4045
rect -278 -4073 -250 -4045
rect -212 -4073 -184 -4045
rect -146 -4073 -118 -4045
rect -80 -4073 -52 -4045
rect -14 -4073 14 -4045
rect 52 -4073 80 -4045
rect 118 -4073 146 -4045
rect 184 -4073 212 -4045
rect 250 -4073 278 -4045
rect 316 -4073 344 -4045
rect -344 -4139 -316 -4111
rect -278 -4139 -250 -4111
rect -212 -4139 -184 -4111
rect -146 -4139 -118 -4111
rect -80 -4139 -52 -4111
rect -14 -4139 14 -4111
rect 52 -4139 80 -4111
rect 118 -4139 146 -4111
rect 184 -4139 212 -4111
rect 250 -4139 278 -4111
rect 316 -4139 344 -4111
rect -344 -4205 -316 -4177
rect -278 -4205 -250 -4177
rect -212 -4205 -184 -4177
rect -146 -4205 -118 -4177
rect -80 -4205 -52 -4177
rect -14 -4205 14 -4177
rect 52 -4205 80 -4177
rect 118 -4205 146 -4177
rect 184 -4205 212 -4177
rect 250 -4205 278 -4177
rect 316 -4205 344 -4177
rect -344 -4271 -316 -4243
rect -278 -4271 -250 -4243
rect -212 -4271 -184 -4243
rect -146 -4271 -118 -4243
rect -80 -4271 -52 -4243
rect -14 -4271 14 -4243
rect 52 -4271 80 -4243
rect 118 -4271 146 -4243
rect 184 -4271 212 -4243
rect 250 -4271 278 -4243
rect 316 -4271 344 -4243
rect -344 -4337 -316 -4309
rect -278 -4337 -250 -4309
rect -212 -4337 -184 -4309
rect -146 -4337 -118 -4309
rect -80 -4337 -52 -4309
rect -14 -4337 14 -4309
rect 52 -4337 80 -4309
rect 118 -4337 146 -4309
rect 184 -4337 212 -4309
rect 250 -4337 278 -4309
rect 316 -4337 344 -4309
rect -344 -4403 -316 -4375
rect -278 -4403 -250 -4375
rect -212 -4403 -184 -4375
rect -146 -4403 -118 -4375
rect -80 -4403 -52 -4375
rect -14 -4403 14 -4375
rect 52 -4403 80 -4375
rect 118 -4403 146 -4375
rect 184 -4403 212 -4375
rect 250 -4403 278 -4375
rect 316 -4403 344 -4375
rect -344 -4469 -316 -4441
rect -278 -4469 -250 -4441
rect -212 -4469 -184 -4441
rect -146 -4469 -118 -4441
rect -80 -4469 -52 -4441
rect -14 -4469 14 -4441
rect 52 -4469 80 -4441
rect 118 -4469 146 -4441
rect 184 -4469 212 -4441
rect 250 -4469 278 -4441
rect 316 -4469 344 -4441
rect -344 -4535 -316 -4507
rect -278 -4535 -250 -4507
rect -212 -4535 -184 -4507
rect -146 -4535 -118 -4507
rect -80 -4535 -52 -4507
rect -14 -4535 14 -4507
rect 52 -4535 80 -4507
rect 118 -4535 146 -4507
rect 184 -4535 212 -4507
rect 250 -4535 278 -4507
rect 316 -4535 344 -4507
rect -344 -4601 -316 -4573
rect -278 -4601 -250 -4573
rect -212 -4601 -184 -4573
rect -146 -4601 -118 -4573
rect -80 -4601 -52 -4573
rect -14 -4601 14 -4573
rect 52 -4601 80 -4573
rect 118 -4601 146 -4573
rect 184 -4601 212 -4573
rect 250 -4601 278 -4573
rect 316 -4601 344 -4573
rect -344 -4667 -316 -4639
rect -278 -4667 -250 -4639
rect -212 -4667 -184 -4639
rect -146 -4667 -118 -4639
rect -80 -4667 -52 -4639
rect -14 -4667 14 -4639
rect 52 -4667 80 -4639
rect 118 -4667 146 -4639
rect 184 -4667 212 -4639
rect 250 -4667 278 -4639
rect 316 -4667 344 -4639
rect -344 -4733 -316 -4705
rect -278 -4733 -250 -4705
rect -212 -4733 -184 -4705
rect -146 -4733 -118 -4705
rect -80 -4733 -52 -4705
rect -14 -4733 14 -4705
rect 52 -4733 80 -4705
rect 118 -4733 146 -4705
rect 184 -4733 212 -4705
rect 250 -4733 278 -4705
rect 316 -4733 344 -4705
rect -344 -4799 -316 -4771
rect -278 -4799 -250 -4771
rect -212 -4799 -184 -4771
rect -146 -4799 -118 -4771
rect -80 -4799 -52 -4771
rect -14 -4799 14 -4771
rect 52 -4799 80 -4771
rect 118 -4799 146 -4771
rect 184 -4799 212 -4771
rect 250 -4799 278 -4771
rect 316 -4799 344 -4771
rect -344 -4865 -316 -4837
rect -278 -4865 -250 -4837
rect -212 -4865 -184 -4837
rect -146 -4865 -118 -4837
rect -80 -4865 -52 -4837
rect -14 -4865 14 -4837
rect 52 -4865 80 -4837
rect 118 -4865 146 -4837
rect 184 -4865 212 -4837
rect 250 -4865 278 -4837
rect 316 -4865 344 -4837
rect -344 -4931 -316 -4903
rect -278 -4931 -250 -4903
rect -212 -4931 -184 -4903
rect -146 -4931 -118 -4903
rect -80 -4931 -52 -4903
rect -14 -4931 14 -4903
rect 52 -4931 80 -4903
rect 118 -4931 146 -4903
rect 184 -4931 212 -4903
rect 250 -4931 278 -4903
rect 316 -4931 344 -4903
rect -344 -4997 -316 -4969
rect -278 -4997 -250 -4969
rect -212 -4997 -184 -4969
rect -146 -4997 -118 -4969
rect -80 -4997 -52 -4969
rect -14 -4997 14 -4969
rect 52 -4997 80 -4969
rect 118 -4997 146 -4969
rect 184 -4997 212 -4969
rect 250 -4997 278 -4969
rect 316 -4997 344 -4969
rect -344 -5063 -316 -5035
rect -278 -5063 -250 -5035
rect -212 -5063 -184 -5035
rect -146 -5063 -118 -5035
rect -80 -5063 -52 -5035
rect -14 -5063 14 -5035
rect 52 -5063 80 -5035
rect 118 -5063 146 -5035
rect 184 -5063 212 -5035
rect 250 -5063 278 -5035
rect 316 -5063 344 -5035
<< metal4 >>
rect -349 5063 349 5068
rect -349 5035 -344 5063
rect -316 5035 -278 5063
rect -250 5035 -212 5063
rect -184 5035 -146 5063
rect -118 5035 -80 5063
rect -52 5035 -14 5063
rect 14 5035 52 5063
rect 80 5035 118 5063
rect 146 5035 184 5063
rect 212 5035 250 5063
rect 278 5035 316 5063
rect 344 5035 349 5063
rect -349 4997 349 5035
rect -349 4969 -344 4997
rect -316 4969 -278 4997
rect -250 4969 -212 4997
rect -184 4969 -146 4997
rect -118 4969 -80 4997
rect -52 4969 -14 4997
rect 14 4969 52 4997
rect 80 4969 118 4997
rect 146 4969 184 4997
rect 212 4969 250 4997
rect 278 4969 316 4997
rect 344 4969 349 4997
rect -349 4931 349 4969
rect -349 4903 -344 4931
rect -316 4903 -278 4931
rect -250 4903 -212 4931
rect -184 4903 -146 4931
rect -118 4903 -80 4931
rect -52 4903 -14 4931
rect 14 4903 52 4931
rect 80 4903 118 4931
rect 146 4903 184 4931
rect 212 4903 250 4931
rect 278 4903 316 4931
rect 344 4903 349 4931
rect -349 4865 349 4903
rect -349 4837 -344 4865
rect -316 4837 -278 4865
rect -250 4837 -212 4865
rect -184 4837 -146 4865
rect -118 4837 -80 4865
rect -52 4837 -14 4865
rect 14 4837 52 4865
rect 80 4837 118 4865
rect 146 4837 184 4865
rect 212 4837 250 4865
rect 278 4837 316 4865
rect 344 4837 349 4865
rect -349 4799 349 4837
rect -349 4771 -344 4799
rect -316 4771 -278 4799
rect -250 4771 -212 4799
rect -184 4771 -146 4799
rect -118 4771 -80 4799
rect -52 4771 -14 4799
rect 14 4771 52 4799
rect 80 4771 118 4799
rect 146 4771 184 4799
rect 212 4771 250 4799
rect 278 4771 316 4799
rect 344 4771 349 4799
rect -349 4733 349 4771
rect -349 4705 -344 4733
rect -316 4705 -278 4733
rect -250 4705 -212 4733
rect -184 4705 -146 4733
rect -118 4705 -80 4733
rect -52 4705 -14 4733
rect 14 4705 52 4733
rect 80 4705 118 4733
rect 146 4705 184 4733
rect 212 4705 250 4733
rect 278 4705 316 4733
rect 344 4705 349 4733
rect -349 4667 349 4705
rect -349 4639 -344 4667
rect -316 4639 -278 4667
rect -250 4639 -212 4667
rect -184 4639 -146 4667
rect -118 4639 -80 4667
rect -52 4639 -14 4667
rect 14 4639 52 4667
rect 80 4639 118 4667
rect 146 4639 184 4667
rect 212 4639 250 4667
rect 278 4639 316 4667
rect 344 4639 349 4667
rect -349 4601 349 4639
rect -349 4573 -344 4601
rect -316 4573 -278 4601
rect -250 4573 -212 4601
rect -184 4573 -146 4601
rect -118 4573 -80 4601
rect -52 4573 -14 4601
rect 14 4573 52 4601
rect 80 4573 118 4601
rect 146 4573 184 4601
rect 212 4573 250 4601
rect 278 4573 316 4601
rect 344 4573 349 4601
rect -349 4535 349 4573
rect -349 4507 -344 4535
rect -316 4507 -278 4535
rect -250 4507 -212 4535
rect -184 4507 -146 4535
rect -118 4507 -80 4535
rect -52 4507 -14 4535
rect 14 4507 52 4535
rect 80 4507 118 4535
rect 146 4507 184 4535
rect 212 4507 250 4535
rect 278 4507 316 4535
rect 344 4507 349 4535
rect -349 4469 349 4507
rect -349 4441 -344 4469
rect -316 4441 -278 4469
rect -250 4441 -212 4469
rect -184 4441 -146 4469
rect -118 4441 -80 4469
rect -52 4441 -14 4469
rect 14 4441 52 4469
rect 80 4441 118 4469
rect 146 4441 184 4469
rect 212 4441 250 4469
rect 278 4441 316 4469
rect 344 4441 349 4469
rect -349 4403 349 4441
rect -349 4375 -344 4403
rect -316 4375 -278 4403
rect -250 4375 -212 4403
rect -184 4375 -146 4403
rect -118 4375 -80 4403
rect -52 4375 -14 4403
rect 14 4375 52 4403
rect 80 4375 118 4403
rect 146 4375 184 4403
rect 212 4375 250 4403
rect 278 4375 316 4403
rect 344 4375 349 4403
rect -349 4337 349 4375
rect -349 4309 -344 4337
rect -316 4309 -278 4337
rect -250 4309 -212 4337
rect -184 4309 -146 4337
rect -118 4309 -80 4337
rect -52 4309 -14 4337
rect 14 4309 52 4337
rect 80 4309 118 4337
rect 146 4309 184 4337
rect 212 4309 250 4337
rect 278 4309 316 4337
rect 344 4309 349 4337
rect -349 4271 349 4309
rect -349 4243 -344 4271
rect -316 4243 -278 4271
rect -250 4243 -212 4271
rect -184 4243 -146 4271
rect -118 4243 -80 4271
rect -52 4243 -14 4271
rect 14 4243 52 4271
rect 80 4243 118 4271
rect 146 4243 184 4271
rect 212 4243 250 4271
rect 278 4243 316 4271
rect 344 4243 349 4271
rect -349 4205 349 4243
rect -349 4177 -344 4205
rect -316 4177 -278 4205
rect -250 4177 -212 4205
rect -184 4177 -146 4205
rect -118 4177 -80 4205
rect -52 4177 -14 4205
rect 14 4177 52 4205
rect 80 4177 118 4205
rect 146 4177 184 4205
rect 212 4177 250 4205
rect 278 4177 316 4205
rect 344 4177 349 4205
rect -349 4139 349 4177
rect -349 4111 -344 4139
rect -316 4111 -278 4139
rect -250 4111 -212 4139
rect -184 4111 -146 4139
rect -118 4111 -80 4139
rect -52 4111 -14 4139
rect 14 4111 52 4139
rect 80 4111 118 4139
rect 146 4111 184 4139
rect 212 4111 250 4139
rect 278 4111 316 4139
rect 344 4111 349 4139
rect -349 4073 349 4111
rect -349 4045 -344 4073
rect -316 4045 -278 4073
rect -250 4045 -212 4073
rect -184 4045 -146 4073
rect -118 4045 -80 4073
rect -52 4045 -14 4073
rect 14 4045 52 4073
rect 80 4045 118 4073
rect 146 4045 184 4073
rect 212 4045 250 4073
rect 278 4045 316 4073
rect 344 4045 349 4073
rect -349 4007 349 4045
rect -349 3979 -344 4007
rect -316 3979 -278 4007
rect -250 3979 -212 4007
rect -184 3979 -146 4007
rect -118 3979 -80 4007
rect -52 3979 -14 4007
rect 14 3979 52 4007
rect 80 3979 118 4007
rect 146 3979 184 4007
rect 212 3979 250 4007
rect 278 3979 316 4007
rect 344 3979 349 4007
rect -349 3941 349 3979
rect -349 3913 -344 3941
rect -316 3913 -278 3941
rect -250 3913 -212 3941
rect -184 3913 -146 3941
rect -118 3913 -80 3941
rect -52 3913 -14 3941
rect 14 3913 52 3941
rect 80 3913 118 3941
rect 146 3913 184 3941
rect 212 3913 250 3941
rect 278 3913 316 3941
rect 344 3913 349 3941
rect -349 3875 349 3913
rect -349 3847 -344 3875
rect -316 3847 -278 3875
rect -250 3847 -212 3875
rect -184 3847 -146 3875
rect -118 3847 -80 3875
rect -52 3847 -14 3875
rect 14 3847 52 3875
rect 80 3847 118 3875
rect 146 3847 184 3875
rect 212 3847 250 3875
rect 278 3847 316 3875
rect 344 3847 349 3875
rect -349 3809 349 3847
rect -349 3781 -344 3809
rect -316 3781 -278 3809
rect -250 3781 -212 3809
rect -184 3781 -146 3809
rect -118 3781 -80 3809
rect -52 3781 -14 3809
rect 14 3781 52 3809
rect 80 3781 118 3809
rect 146 3781 184 3809
rect 212 3781 250 3809
rect 278 3781 316 3809
rect 344 3781 349 3809
rect -349 3743 349 3781
rect -349 3715 -344 3743
rect -316 3715 -278 3743
rect -250 3715 -212 3743
rect -184 3715 -146 3743
rect -118 3715 -80 3743
rect -52 3715 -14 3743
rect 14 3715 52 3743
rect 80 3715 118 3743
rect 146 3715 184 3743
rect 212 3715 250 3743
rect 278 3715 316 3743
rect 344 3715 349 3743
rect -349 3677 349 3715
rect -349 3649 -344 3677
rect -316 3649 -278 3677
rect -250 3649 -212 3677
rect -184 3649 -146 3677
rect -118 3649 -80 3677
rect -52 3649 -14 3677
rect 14 3649 52 3677
rect 80 3649 118 3677
rect 146 3649 184 3677
rect 212 3649 250 3677
rect 278 3649 316 3677
rect 344 3649 349 3677
rect -349 3611 349 3649
rect -349 3583 -344 3611
rect -316 3583 -278 3611
rect -250 3583 -212 3611
rect -184 3583 -146 3611
rect -118 3583 -80 3611
rect -52 3583 -14 3611
rect 14 3583 52 3611
rect 80 3583 118 3611
rect 146 3583 184 3611
rect 212 3583 250 3611
rect 278 3583 316 3611
rect 344 3583 349 3611
rect -349 3545 349 3583
rect -349 3517 -344 3545
rect -316 3517 -278 3545
rect -250 3517 -212 3545
rect -184 3517 -146 3545
rect -118 3517 -80 3545
rect -52 3517 -14 3545
rect 14 3517 52 3545
rect 80 3517 118 3545
rect 146 3517 184 3545
rect 212 3517 250 3545
rect 278 3517 316 3545
rect 344 3517 349 3545
rect -349 3479 349 3517
rect -349 3451 -344 3479
rect -316 3451 -278 3479
rect -250 3451 -212 3479
rect -184 3451 -146 3479
rect -118 3451 -80 3479
rect -52 3451 -14 3479
rect 14 3451 52 3479
rect 80 3451 118 3479
rect 146 3451 184 3479
rect 212 3451 250 3479
rect 278 3451 316 3479
rect 344 3451 349 3479
rect -349 3413 349 3451
rect -349 3385 -344 3413
rect -316 3385 -278 3413
rect -250 3385 -212 3413
rect -184 3385 -146 3413
rect -118 3385 -80 3413
rect -52 3385 -14 3413
rect 14 3385 52 3413
rect 80 3385 118 3413
rect 146 3385 184 3413
rect 212 3385 250 3413
rect 278 3385 316 3413
rect 344 3385 349 3413
rect -349 3347 349 3385
rect -349 3319 -344 3347
rect -316 3319 -278 3347
rect -250 3319 -212 3347
rect -184 3319 -146 3347
rect -118 3319 -80 3347
rect -52 3319 -14 3347
rect 14 3319 52 3347
rect 80 3319 118 3347
rect 146 3319 184 3347
rect 212 3319 250 3347
rect 278 3319 316 3347
rect 344 3319 349 3347
rect -349 3281 349 3319
rect -349 3253 -344 3281
rect -316 3253 -278 3281
rect -250 3253 -212 3281
rect -184 3253 -146 3281
rect -118 3253 -80 3281
rect -52 3253 -14 3281
rect 14 3253 52 3281
rect 80 3253 118 3281
rect 146 3253 184 3281
rect 212 3253 250 3281
rect 278 3253 316 3281
rect 344 3253 349 3281
rect -349 3215 349 3253
rect -349 3187 -344 3215
rect -316 3187 -278 3215
rect -250 3187 -212 3215
rect -184 3187 -146 3215
rect -118 3187 -80 3215
rect -52 3187 -14 3215
rect 14 3187 52 3215
rect 80 3187 118 3215
rect 146 3187 184 3215
rect 212 3187 250 3215
rect 278 3187 316 3215
rect 344 3187 349 3215
rect -349 3149 349 3187
rect -349 3121 -344 3149
rect -316 3121 -278 3149
rect -250 3121 -212 3149
rect -184 3121 -146 3149
rect -118 3121 -80 3149
rect -52 3121 -14 3149
rect 14 3121 52 3149
rect 80 3121 118 3149
rect 146 3121 184 3149
rect 212 3121 250 3149
rect 278 3121 316 3149
rect 344 3121 349 3149
rect -349 3083 349 3121
rect -349 3055 -344 3083
rect -316 3055 -278 3083
rect -250 3055 -212 3083
rect -184 3055 -146 3083
rect -118 3055 -80 3083
rect -52 3055 -14 3083
rect 14 3055 52 3083
rect 80 3055 118 3083
rect 146 3055 184 3083
rect 212 3055 250 3083
rect 278 3055 316 3083
rect 344 3055 349 3083
rect -349 3017 349 3055
rect -349 2989 -344 3017
rect -316 2989 -278 3017
rect -250 2989 -212 3017
rect -184 2989 -146 3017
rect -118 2989 -80 3017
rect -52 2989 -14 3017
rect 14 2989 52 3017
rect 80 2989 118 3017
rect 146 2989 184 3017
rect 212 2989 250 3017
rect 278 2989 316 3017
rect 344 2989 349 3017
rect -349 2951 349 2989
rect -349 2923 -344 2951
rect -316 2923 -278 2951
rect -250 2923 -212 2951
rect -184 2923 -146 2951
rect -118 2923 -80 2951
rect -52 2923 -14 2951
rect 14 2923 52 2951
rect 80 2923 118 2951
rect 146 2923 184 2951
rect 212 2923 250 2951
rect 278 2923 316 2951
rect 344 2923 349 2951
rect -349 2885 349 2923
rect -349 2857 -344 2885
rect -316 2857 -278 2885
rect -250 2857 -212 2885
rect -184 2857 -146 2885
rect -118 2857 -80 2885
rect -52 2857 -14 2885
rect 14 2857 52 2885
rect 80 2857 118 2885
rect 146 2857 184 2885
rect 212 2857 250 2885
rect 278 2857 316 2885
rect 344 2857 349 2885
rect -349 2819 349 2857
rect -349 2791 -344 2819
rect -316 2791 -278 2819
rect -250 2791 -212 2819
rect -184 2791 -146 2819
rect -118 2791 -80 2819
rect -52 2791 -14 2819
rect 14 2791 52 2819
rect 80 2791 118 2819
rect 146 2791 184 2819
rect 212 2791 250 2819
rect 278 2791 316 2819
rect 344 2791 349 2819
rect -349 2753 349 2791
rect -349 2725 -344 2753
rect -316 2725 -278 2753
rect -250 2725 -212 2753
rect -184 2725 -146 2753
rect -118 2725 -80 2753
rect -52 2725 -14 2753
rect 14 2725 52 2753
rect 80 2725 118 2753
rect 146 2725 184 2753
rect 212 2725 250 2753
rect 278 2725 316 2753
rect 344 2725 349 2753
rect -349 2687 349 2725
rect -349 2659 -344 2687
rect -316 2659 -278 2687
rect -250 2659 -212 2687
rect -184 2659 -146 2687
rect -118 2659 -80 2687
rect -52 2659 -14 2687
rect 14 2659 52 2687
rect 80 2659 118 2687
rect 146 2659 184 2687
rect 212 2659 250 2687
rect 278 2659 316 2687
rect 344 2659 349 2687
rect -349 2621 349 2659
rect -349 2593 -344 2621
rect -316 2593 -278 2621
rect -250 2593 -212 2621
rect -184 2593 -146 2621
rect -118 2593 -80 2621
rect -52 2593 -14 2621
rect 14 2593 52 2621
rect 80 2593 118 2621
rect 146 2593 184 2621
rect 212 2593 250 2621
rect 278 2593 316 2621
rect 344 2593 349 2621
rect -349 2555 349 2593
rect -349 2527 -344 2555
rect -316 2527 -278 2555
rect -250 2527 -212 2555
rect -184 2527 -146 2555
rect -118 2527 -80 2555
rect -52 2527 -14 2555
rect 14 2527 52 2555
rect 80 2527 118 2555
rect 146 2527 184 2555
rect 212 2527 250 2555
rect 278 2527 316 2555
rect 344 2527 349 2555
rect -349 2489 349 2527
rect -349 2461 -344 2489
rect -316 2461 -278 2489
rect -250 2461 -212 2489
rect -184 2461 -146 2489
rect -118 2461 -80 2489
rect -52 2461 -14 2489
rect 14 2461 52 2489
rect 80 2461 118 2489
rect 146 2461 184 2489
rect 212 2461 250 2489
rect 278 2461 316 2489
rect 344 2461 349 2489
rect -349 2423 349 2461
rect -349 2395 -344 2423
rect -316 2395 -278 2423
rect -250 2395 -212 2423
rect -184 2395 -146 2423
rect -118 2395 -80 2423
rect -52 2395 -14 2423
rect 14 2395 52 2423
rect 80 2395 118 2423
rect 146 2395 184 2423
rect 212 2395 250 2423
rect 278 2395 316 2423
rect 344 2395 349 2423
rect -349 2357 349 2395
rect -349 2329 -344 2357
rect -316 2329 -278 2357
rect -250 2329 -212 2357
rect -184 2329 -146 2357
rect -118 2329 -80 2357
rect -52 2329 -14 2357
rect 14 2329 52 2357
rect 80 2329 118 2357
rect 146 2329 184 2357
rect 212 2329 250 2357
rect 278 2329 316 2357
rect 344 2329 349 2357
rect -349 2291 349 2329
rect -349 2263 -344 2291
rect -316 2263 -278 2291
rect -250 2263 -212 2291
rect -184 2263 -146 2291
rect -118 2263 -80 2291
rect -52 2263 -14 2291
rect 14 2263 52 2291
rect 80 2263 118 2291
rect 146 2263 184 2291
rect 212 2263 250 2291
rect 278 2263 316 2291
rect 344 2263 349 2291
rect -349 2225 349 2263
rect -349 2197 -344 2225
rect -316 2197 -278 2225
rect -250 2197 -212 2225
rect -184 2197 -146 2225
rect -118 2197 -80 2225
rect -52 2197 -14 2225
rect 14 2197 52 2225
rect 80 2197 118 2225
rect 146 2197 184 2225
rect 212 2197 250 2225
rect 278 2197 316 2225
rect 344 2197 349 2225
rect -349 2159 349 2197
rect -349 2131 -344 2159
rect -316 2131 -278 2159
rect -250 2131 -212 2159
rect -184 2131 -146 2159
rect -118 2131 -80 2159
rect -52 2131 -14 2159
rect 14 2131 52 2159
rect 80 2131 118 2159
rect 146 2131 184 2159
rect 212 2131 250 2159
rect 278 2131 316 2159
rect 344 2131 349 2159
rect -349 2093 349 2131
rect -349 2065 -344 2093
rect -316 2065 -278 2093
rect -250 2065 -212 2093
rect -184 2065 -146 2093
rect -118 2065 -80 2093
rect -52 2065 -14 2093
rect 14 2065 52 2093
rect 80 2065 118 2093
rect 146 2065 184 2093
rect 212 2065 250 2093
rect 278 2065 316 2093
rect 344 2065 349 2093
rect -349 2027 349 2065
rect -349 1999 -344 2027
rect -316 1999 -278 2027
rect -250 1999 -212 2027
rect -184 1999 -146 2027
rect -118 1999 -80 2027
rect -52 1999 -14 2027
rect 14 1999 52 2027
rect 80 1999 118 2027
rect 146 1999 184 2027
rect 212 1999 250 2027
rect 278 1999 316 2027
rect 344 1999 349 2027
rect -349 1961 349 1999
rect -349 1933 -344 1961
rect -316 1933 -278 1961
rect -250 1933 -212 1961
rect -184 1933 -146 1961
rect -118 1933 -80 1961
rect -52 1933 -14 1961
rect 14 1933 52 1961
rect 80 1933 118 1961
rect 146 1933 184 1961
rect 212 1933 250 1961
rect 278 1933 316 1961
rect 344 1933 349 1961
rect -349 1895 349 1933
rect -349 1867 -344 1895
rect -316 1867 -278 1895
rect -250 1867 -212 1895
rect -184 1867 -146 1895
rect -118 1867 -80 1895
rect -52 1867 -14 1895
rect 14 1867 52 1895
rect 80 1867 118 1895
rect 146 1867 184 1895
rect 212 1867 250 1895
rect 278 1867 316 1895
rect 344 1867 349 1895
rect -349 1829 349 1867
rect -349 1801 -344 1829
rect -316 1801 -278 1829
rect -250 1801 -212 1829
rect -184 1801 -146 1829
rect -118 1801 -80 1829
rect -52 1801 -14 1829
rect 14 1801 52 1829
rect 80 1801 118 1829
rect 146 1801 184 1829
rect 212 1801 250 1829
rect 278 1801 316 1829
rect 344 1801 349 1829
rect -349 1763 349 1801
rect -349 1735 -344 1763
rect -316 1735 -278 1763
rect -250 1735 -212 1763
rect -184 1735 -146 1763
rect -118 1735 -80 1763
rect -52 1735 -14 1763
rect 14 1735 52 1763
rect 80 1735 118 1763
rect 146 1735 184 1763
rect 212 1735 250 1763
rect 278 1735 316 1763
rect 344 1735 349 1763
rect -349 1697 349 1735
rect -349 1669 -344 1697
rect -316 1669 -278 1697
rect -250 1669 -212 1697
rect -184 1669 -146 1697
rect -118 1669 -80 1697
rect -52 1669 -14 1697
rect 14 1669 52 1697
rect 80 1669 118 1697
rect 146 1669 184 1697
rect 212 1669 250 1697
rect 278 1669 316 1697
rect 344 1669 349 1697
rect -349 1631 349 1669
rect -349 1603 -344 1631
rect -316 1603 -278 1631
rect -250 1603 -212 1631
rect -184 1603 -146 1631
rect -118 1603 -80 1631
rect -52 1603 -14 1631
rect 14 1603 52 1631
rect 80 1603 118 1631
rect 146 1603 184 1631
rect 212 1603 250 1631
rect 278 1603 316 1631
rect 344 1603 349 1631
rect -349 1565 349 1603
rect -349 1537 -344 1565
rect -316 1537 -278 1565
rect -250 1537 -212 1565
rect -184 1537 -146 1565
rect -118 1537 -80 1565
rect -52 1537 -14 1565
rect 14 1537 52 1565
rect 80 1537 118 1565
rect 146 1537 184 1565
rect 212 1537 250 1565
rect 278 1537 316 1565
rect 344 1537 349 1565
rect -349 1499 349 1537
rect -349 1471 -344 1499
rect -316 1471 -278 1499
rect -250 1471 -212 1499
rect -184 1471 -146 1499
rect -118 1471 -80 1499
rect -52 1471 -14 1499
rect 14 1471 52 1499
rect 80 1471 118 1499
rect 146 1471 184 1499
rect 212 1471 250 1499
rect 278 1471 316 1499
rect 344 1471 349 1499
rect -349 1433 349 1471
rect -349 1405 -344 1433
rect -316 1405 -278 1433
rect -250 1405 -212 1433
rect -184 1405 -146 1433
rect -118 1405 -80 1433
rect -52 1405 -14 1433
rect 14 1405 52 1433
rect 80 1405 118 1433
rect 146 1405 184 1433
rect 212 1405 250 1433
rect 278 1405 316 1433
rect 344 1405 349 1433
rect -349 1367 349 1405
rect -349 1339 -344 1367
rect -316 1339 -278 1367
rect -250 1339 -212 1367
rect -184 1339 -146 1367
rect -118 1339 -80 1367
rect -52 1339 -14 1367
rect 14 1339 52 1367
rect 80 1339 118 1367
rect 146 1339 184 1367
rect 212 1339 250 1367
rect 278 1339 316 1367
rect 344 1339 349 1367
rect -349 1301 349 1339
rect -349 1273 -344 1301
rect -316 1273 -278 1301
rect -250 1273 -212 1301
rect -184 1273 -146 1301
rect -118 1273 -80 1301
rect -52 1273 -14 1301
rect 14 1273 52 1301
rect 80 1273 118 1301
rect 146 1273 184 1301
rect 212 1273 250 1301
rect 278 1273 316 1301
rect 344 1273 349 1301
rect -349 1235 349 1273
rect -349 1207 -344 1235
rect -316 1207 -278 1235
rect -250 1207 -212 1235
rect -184 1207 -146 1235
rect -118 1207 -80 1235
rect -52 1207 -14 1235
rect 14 1207 52 1235
rect 80 1207 118 1235
rect 146 1207 184 1235
rect 212 1207 250 1235
rect 278 1207 316 1235
rect 344 1207 349 1235
rect -349 1169 349 1207
rect -349 1141 -344 1169
rect -316 1141 -278 1169
rect -250 1141 -212 1169
rect -184 1141 -146 1169
rect -118 1141 -80 1169
rect -52 1141 -14 1169
rect 14 1141 52 1169
rect 80 1141 118 1169
rect 146 1141 184 1169
rect 212 1141 250 1169
rect 278 1141 316 1169
rect 344 1141 349 1169
rect -349 1103 349 1141
rect -349 1075 -344 1103
rect -316 1075 -278 1103
rect -250 1075 -212 1103
rect -184 1075 -146 1103
rect -118 1075 -80 1103
rect -52 1075 -14 1103
rect 14 1075 52 1103
rect 80 1075 118 1103
rect 146 1075 184 1103
rect 212 1075 250 1103
rect 278 1075 316 1103
rect 344 1075 349 1103
rect -349 1037 349 1075
rect -349 1009 -344 1037
rect -316 1009 -278 1037
rect -250 1009 -212 1037
rect -184 1009 -146 1037
rect -118 1009 -80 1037
rect -52 1009 -14 1037
rect 14 1009 52 1037
rect 80 1009 118 1037
rect 146 1009 184 1037
rect 212 1009 250 1037
rect 278 1009 316 1037
rect 344 1009 349 1037
rect -349 971 349 1009
rect -349 943 -344 971
rect -316 943 -278 971
rect -250 943 -212 971
rect -184 943 -146 971
rect -118 943 -80 971
rect -52 943 -14 971
rect 14 943 52 971
rect 80 943 118 971
rect 146 943 184 971
rect 212 943 250 971
rect 278 943 316 971
rect 344 943 349 971
rect -349 905 349 943
rect -349 877 -344 905
rect -316 877 -278 905
rect -250 877 -212 905
rect -184 877 -146 905
rect -118 877 -80 905
rect -52 877 -14 905
rect 14 877 52 905
rect 80 877 118 905
rect 146 877 184 905
rect 212 877 250 905
rect 278 877 316 905
rect 344 877 349 905
rect -349 839 349 877
rect -349 811 -344 839
rect -316 811 -278 839
rect -250 811 -212 839
rect -184 811 -146 839
rect -118 811 -80 839
rect -52 811 -14 839
rect 14 811 52 839
rect 80 811 118 839
rect 146 811 184 839
rect 212 811 250 839
rect 278 811 316 839
rect 344 811 349 839
rect -349 773 349 811
rect -349 745 -344 773
rect -316 745 -278 773
rect -250 745 -212 773
rect -184 745 -146 773
rect -118 745 -80 773
rect -52 745 -14 773
rect 14 745 52 773
rect 80 745 118 773
rect 146 745 184 773
rect 212 745 250 773
rect 278 745 316 773
rect 344 745 349 773
rect -349 707 349 745
rect -349 679 -344 707
rect -316 679 -278 707
rect -250 679 -212 707
rect -184 679 -146 707
rect -118 679 -80 707
rect -52 679 -14 707
rect 14 679 52 707
rect 80 679 118 707
rect 146 679 184 707
rect 212 679 250 707
rect 278 679 316 707
rect 344 679 349 707
rect -349 641 349 679
rect -349 613 -344 641
rect -316 613 -278 641
rect -250 613 -212 641
rect -184 613 -146 641
rect -118 613 -80 641
rect -52 613 -14 641
rect 14 613 52 641
rect 80 613 118 641
rect 146 613 184 641
rect 212 613 250 641
rect 278 613 316 641
rect 344 613 349 641
rect -349 575 349 613
rect -349 547 -344 575
rect -316 547 -278 575
rect -250 547 -212 575
rect -184 547 -146 575
rect -118 547 -80 575
rect -52 547 -14 575
rect 14 547 52 575
rect 80 547 118 575
rect 146 547 184 575
rect 212 547 250 575
rect 278 547 316 575
rect 344 547 349 575
rect -349 509 349 547
rect -349 481 -344 509
rect -316 481 -278 509
rect -250 481 -212 509
rect -184 481 -146 509
rect -118 481 -80 509
rect -52 481 -14 509
rect 14 481 52 509
rect 80 481 118 509
rect 146 481 184 509
rect 212 481 250 509
rect 278 481 316 509
rect 344 481 349 509
rect -349 443 349 481
rect -349 415 -344 443
rect -316 415 -278 443
rect -250 415 -212 443
rect -184 415 -146 443
rect -118 415 -80 443
rect -52 415 -14 443
rect 14 415 52 443
rect 80 415 118 443
rect 146 415 184 443
rect 212 415 250 443
rect 278 415 316 443
rect 344 415 349 443
rect -349 377 349 415
rect -349 349 -344 377
rect -316 349 -278 377
rect -250 349 -212 377
rect -184 349 -146 377
rect -118 349 -80 377
rect -52 349 -14 377
rect 14 349 52 377
rect 80 349 118 377
rect 146 349 184 377
rect 212 349 250 377
rect 278 349 316 377
rect 344 349 349 377
rect -349 311 349 349
rect -349 283 -344 311
rect -316 283 -278 311
rect -250 283 -212 311
rect -184 283 -146 311
rect -118 283 -80 311
rect -52 283 -14 311
rect 14 283 52 311
rect 80 283 118 311
rect 146 283 184 311
rect 212 283 250 311
rect 278 283 316 311
rect 344 283 349 311
rect -349 245 349 283
rect -349 217 -344 245
rect -316 217 -278 245
rect -250 217 -212 245
rect -184 217 -146 245
rect -118 217 -80 245
rect -52 217 -14 245
rect 14 217 52 245
rect 80 217 118 245
rect 146 217 184 245
rect 212 217 250 245
rect 278 217 316 245
rect 344 217 349 245
rect -349 179 349 217
rect -349 151 -344 179
rect -316 151 -278 179
rect -250 151 -212 179
rect -184 151 -146 179
rect -118 151 -80 179
rect -52 151 -14 179
rect 14 151 52 179
rect 80 151 118 179
rect 146 151 184 179
rect 212 151 250 179
rect 278 151 316 179
rect 344 151 349 179
rect -349 113 349 151
rect -349 85 -344 113
rect -316 85 -278 113
rect -250 85 -212 113
rect -184 85 -146 113
rect -118 85 -80 113
rect -52 85 -14 113
rect 14 85 52 113
rect 80 85 118 113
rect 146 85 184 113
rect 212 85 250 113
rect 278 85 316 113
rect 344 85 349 113
rect -349 47 349 85
rect -349 19 -344 47
rect -316 19 -278 47
rect -250 19 -212 47
rect -184 19 -146 47
rect -118 19 -80 47
rect -52 19 -14 47
rect 14 19 52 47
rect 80 19 118 47
rect 146 19 184 47
rect 212 19 250 47
rect 278 19 316 47
rect 344 19 349 47
rect -349 -19 349 19
rect -349 -47 -344 -19
rect -316 -47 -278 -19
rect -250 -47 -212 -19
rect -184 -47 -146 -19
rect -118 -47 -80 -19
rect -52 -47 -14 -19
rect 14 -47 52 -19
rect 80 -47 118 -19
rect 146 -47 184 -19
rect 212 -47 250 -19
rect 278 -47 316 -19
rect 344 -47 349 -19
rect -349 -85 349 -47
rect -349 -113 -344 -85
rect -316 -113 -278 -85
rect -250 -113 -212 -85
rect -184 -113 -146 -85
rect -118 -113 -80 -85
rect -52 -113 -14 -85
rect 14 -113 52 -85
rect 80 -113 118 -85
rect 146 -113 184 -85
rect 212 -113 250 -85
rect 278 -113 316 -85
rect 344 -113 349 -85
rect -349 -151 349 -113
rect -349 -179 -344 -151
rect -316 -179 -278 -151
rect -250 -179 -212 -151
rect -184 -179 -146 -151
rect -118 -179 -80 -151
rect -52 -179 -14 -151
rect 14 -179 52 -151
rect 80 -179 118 -151
rect 146 -179 184 -151
rect 212 -179 250 -151
rect 278 -179 316 -151
rect 344 -179 349 -151
rect -349 -217 349 -179
rect -349 -245 -344 -217
rect -316 -245 -278 -217
rect -250 -245 -212 -217
rect -184 -245 -146 -217
rect -118 -245 -80 -217
rect -52 -245 -14 -217
rect 14 -245 52 -217
rect 80 -245 118 -217
rect 146 -245 184 -217
rect 212 -245 250 -217
rect 278 -245 316 -217
rect 344 -245 349 -217
rect -349 -283 349 -245
rect -349 -311 -344 -283
rect -316 -311 -278 -283
rect -250 -311 -212 -283
rect -184 -311 -146 -283
rect -118 -311 -80 -283
rect -52 -311 -14 -283
rect 14 -311 52 -283
rect 80 -311 118 -283
rect 146 -311 184 -283
rect 212 -311 250 -283
rect 278 -311 316 -283
rect 344 -311 349 -283
rect -349 -349 349 -311
rect -349 -377 -344 -349
rect -316 -377 -278 -349
rect -250 -377 -212 -349
rect -184 -377 -146 -349
rect -118 -377 -80 -349
rect -52 -377 -14 -349
rect 14 -377 52 -349
rect 80 -377 118 -349
rect 146 -377 184 -349
rect 212 -377 250 -349
rect 278 -377 316 -349
rect 344 -377 349 -349
rect -349 -415 349 -377
rect -349 -443 -344 -415
rect -316 -443 -278 -415
rect -250 -443 -212 -415
rect -184 -443 -146 -415
rect -118 -443 -80 -415
rect -52 -443 -14 -415
rect 14 -443 52 -415
rect 80 -443 118 -415
rect 146 -443 184 -415
rect 212 -443 250 -415
rect 278 -443 316 -415
rect 344 -443 349 -415
rect -349 -481 349 -443
rect -349 -509 -344 -481
rect -316 -509 -278 -481
rect -250 -509 -212 -481
rect -184 -509 -146 -481
rect -118 -509 -80 -481
rect -52 -509 -14 -481
rect 14 -509 52 -481
rect 80 -509 118 -481
rect 146 -509 184 -481
rect 212 -509 250 -481
rect 278 -509 316 -481
rect 344 -509 349 -481
rect -349 -547 349 -509
rect -349 -575 -344 -547
rect -316 -575 -278 -547
rect -250 -575 -212 -547
rect -184 -575 -146 -547
rect -118 -575 -80 -547
rect -52 -575 -14 -547
rect 14 -575 52 -547
rect 80 -575 118 -547
rect 146 -575 184 -547
rect 212 -575 250 -547
rect 278 -575 316 -547
rect 344 -575 349 -547
rect -349 -613 349 -575
rect -349 -641 -344 -613
rect -316 -641 -278 -613
rect -250 -641 -212 -613
rect -184 -641 -146 -613
rect -118 -641 -80 -613
rect -52 -641 -14 -613
rect 14 -641 52 -613
rect 80 -641 118 -613
rect 146 -641 184 -613
rect 212 -641 250 -613
rect 278 -641 316 -613
rect 344 -641 349 -613
rect -349 -679 349 -641
rect -349 -707 -344 -679
rect -316 -707 -278 -679
rect -250 -707 -212 -679
rect -184 -707 -146 -679
rect -118 -707 -80 -679
rect -52 -707 -14 -679
rect 14 -707 52 -679
rect 80 -707 118 -679
rect 146 -707 184 -679
rect 212 -707 250 -679
rect 278 -707 316 -679
rect 344 -707 349 -679
rect -349 -745 349 -707
rect -349 -773 -344 -745
rect -316 -773 -278 -745
rect -250 -773 -212 -745
rect -184 -773 -146 -745
rect -118 -773 -80 -745
rect -52 -773 -14 -745
rect 14 -773 52 -745
rect 80 -773 118 -745
rect 146 -773 184 -745
rect 212 -773 250 -745
rect 278 -773 316 -745
rect 344 -773 349 -745
rect -349 -811 349 -773
rect -349 -839 -344 -811
rect -316 -839 -278 -811
rect -250 -839 -212 -811
rect -184 -839 -146 -811
rect -118 -839 -80 -811
rect -52 -839 -14 -811
rect 14 -839 52 -811
rect 80 -839 118 -811
rect 146 -839 184 -811
rect 212 -839 250 -811
rect 278 -839 316 -811
rect 344 -839 349 -811
rect -349 -877 349 -839
rect -349 -905 -344 -877
rect -316 -905 -278 -877
rect -250 -905 -212 -877
rect -184 -905 -146 -877
rect -118 -905 -80 -877
rect -52 -905 -14 -877
rect 14 -905 52 -877
rect 80 -905 118 -877
rect 146 -905 184 -877
rect 212 -905 250 -877
rect 278 -905 316 -877
rect 344 -905 349 -877
rect -349 -943 349 -905
rect -349 -971 -344 -943
rect -316 -971 -278 -943
rect -250 -971 -212 -943
rect -184 -971 -146 -943
rect -118 -971 -80 -943
rect -52 -971 -14 -943
rect 14 -971 52 -943
rect 80 -971 118 -943
rect 146 -971 184 -943
rect 212 -971 250 -943
rect 278 -971 316 -943
rect 344 -971 349 -943
rect -349 -1009 349 -971
rect -349 -1037 -344 -1009
rect -316 -1037 -278 -1009
rect -250 -1037 -212 -1009
rect -184 -1037 -146 -1009
rect -118 -1037 -80 -1009
rect -52 -1037 -14 -1009
rect 14 -1037 52 -1009
rect 80 -1037 118 -1009
rect 146 -1037 184 -1009
rect 212 -1037 250 -1009
rect 278 -1037 316 -1009
rect 344 -1037 349 -1009
rect -349 -1075 349 -1037
rect -349 -1103 -344 -1075
rect -316 -1103 -278 -1075
rect -250 -1103 -212 -1075
rect -184 -1103 -146 -1075
rect -118 -1103 -80 -1075
rect -52 -1103 -14 -1075
rect 14 -1103 52 -1075
rect 80 -1103 118 -1075
rect 146 -1103 184 -1075
rect 212 -1103 250 -1075
rect 278 -1103 316 -1075
rect 344 -1103 349 -1075
rect -349 -1141 349 -1103
rect -349 -1169 -344 -1141
rect -316 -1169 -278 -1141
rect -250 -1169 -212 -1141
rect -184 -1169 -146 -1141
rect -118 -1169 -80 -1141
rect -52 -1169 -14 -1141
rect 14 -1169 52 -1141
rect 80 -1169 118 -1141
rect 146 -1169 184 -1141
rect 212 -1169 250 -1141
rect 278 -1169 316 -1141
rect 344 -1169 349 -1141
rect -349 -1207 349 -1169
rect -349 -1235 -344 -1207
rect -316 -1235 -278 -1207
rect -250 -1235 -212 -1207
rect -184 -1235 -146 -1207
rect -118 -1235 -80 -1207
rect -52 -1235 -14 -1207
rect 14 -1235 52 -1207
rect 80 -1235 118 -1207
rect 146 -1235 184 -1207
rect 212 -1235 250 -1207
rect 278 -1235 316 -1207
rect 344 -1235 349 -1207
rect -349 -1273 349 -1235
rect -349 -1301 -344 -1273
rect -316 -1301 -278 -1273
rect -250 -1301 -212 -1273
rect -184 -1301 -146 -1273
rect -118 -1301 -80 -1273
rect -52 -1301 -14 -1273
rect 14 -1301 52 -1273
rect 80 -1301 118 -1273
rect 146 -1301 184 -1273
rect 212 -1301 250 -1273
rect 278 -1301 316 -1273
rect 344 -1301 349 -1273
rect -349 -1339 349 -1301
rect -349 -1367 -344 -1339
rect -316 -1367 -278 -1339
rect -250 -1367 -212 -1339
rect -184 -1367 -146 -1339
rect -118 -1367 -80 -1339
rect -52 -1367 -14 -1339
rect 14 -1367 52 -1339
rect 80 -1367 118 -1339
rect 146 -1367 184 -1339
rect 212 -1367 250 -1339
rect 278 -1367 316 -1339
rect 344 -1367 349 -1339
rect -349 -1405 349 -1367
rect -349 -1433 -344 -1405
rect -316 -1433 -278 -1405
rect -250 -1433 -212 -1405
rect -184 -1433 -146 -1405
rect -118 -1433 -80 -1405
rect -52 -1433 -14 -1405
rect 14 -1433 52 -1405
rect 80 -1433 118 -1405
rect 146 -1433 184 -1405
rect 212 -1433 250 -1405
rect 278 -1433 316 -1405
rect 344 -1433 349 -1405
rect -349 -1471 349 -1433
rect -349 -1499 -344 -1471
rect -316 -1499 -278 -1471
rect -250 -1499 -212 -1471
rect -184 -1499 -146 -1471
rect -118 -1499 -80 -1471
rect -52 -1499 -14 -1471
rect 14 -1499 52 -1471
rect 80 -1499 118 -1471
rect 146 -1499 184 -1471
rect 212 -1499 250 -1471
rect 278 -1499 316 -1471
rect 344 -1499 349 -1471
rect -349 -1537 349 -1499
rect -349 -1565 -344 -1537
rect -316 -1565 -278 -1537
rect -250 -1565 -212 -1537
rect -184 -1565 -146 -1537
rect -118 -1565 -80 -1537
rect -52 -1565 -14 -1537
rect 14 -1565 52 -1537
rect 80 -1565 118 -1537
rect 146 -1565 184 -1537
rect 212 -1565 250 -1537
rect 278 -1565 316 -1537
rect 344 -1565 349 -1537
rect -349 -1603 349 -1565
rect -349 -1631 -344 -1603
rect -316 -1631 -278 -1603
rect -250 -1631 -212 -1603
rect -184 -1631 -146 -1603
rect -118 -1631 -80 -1603
rect -52 -1631 -14 -1603
rect 14 -1631 52 -1603
rect 80 -1631 118 -1603
rect 146 -1631 184 -1603
rect 212 -1631 250 -1603
rect 278 -1631 316 -1603
rect 344 -1631 349 -1603
rect -349 -1669 349 -1631
rect -349 -1697 -344 -1669
rect -316 -1697 -278 -1669
rect -250 -1697 -212 -1669
rect -184 -1697 -146 -1669
rect -118 -1697 -80 -1669
rect -52 -1697 -14 -1669
rect 14 -1697 52 -1669
rect 80 -1697 118 -1669
rect 146 -1697 184 -1669
rect 212 -1697 250 -1669
rect 278 -1697 316 -1669
rect 344 -1697 349 -1669
rect -349 -1735 349 -1697
rect -349 -1763 -344 -1735
rect -316 -1763 -278 -1735
rect -250 -1763 -212 -1735
rect -184 -1763 -146 -1735
rect -118 -1763 -80 -1735
rect -52 -1763 -14 -1735
rect 14 -1763 52 -1735
rect 80 -1763 118 -1735
rect 146 -1763 184 -1735
rect 212 -1763 250 -1735
rect 278 -1763 316 -1735
rect 344 -1763 349 -1735
rect -349 -1801 349 -1763
rect -349 -1829 -344 -1801
rect -316 -1829 -278 -1801
rect -250 -1829 -212 -1801
rect -184 -1829 -146 -1801
rect -118 -1829 -80 -1801
rect -52 -1829 -14 -1801
rect 14 -1829 52 -1801
rect 80 -1829 118 -1801
rect 146 -1829 184 -1801
rect 212 -1829 250 -1801
rect 278 -1829 316 -1801
rect 344 -1829 349 -1801
rect -349 -1867 349 -1829
rect -349 -1895 -344 -1867
rect -316 -1895 -278 -1867
rect -250 -1895 -212 -1867
rect -184 -1895 -146 -1867
rect -118 -1895 -80 -1867
rect -52 -1895 -14 -1867
rect 14 -1895 52 -1867
rect 80 -1895 118 -1867
rect 146 -1895 184 -1867
rect 212 -1895 250 -1867
rect 278 -1895 316 -1867
rect 344 -1895 349 -1867
rect -349 -1933 349 -1895
rect -349 -1961 -344 -1933
rect -316 -1961 -278 -1933
rect -250 -1961 -212 -1933
rect -184 -1961 -146 -1933
rect -118 -1961 -80 -1933
rect -52 -1961 -14 -1933
rect 14 -1961 52 -1933
rect 80 -1961 118 -1933
rect 146 -1961 184 -1933
rect 212 -1961 250 -1933
rect 278 -1961 316 -1933
rect 344 -1961 349 -1933
rect -349 -1999 349 -1961
rect -349 -2027 -344 -1999
rect -316 -2027 -278 -1999
rect -250 -2027 -212 -1999
rect -184 -2027 -146 -1999
rect -118 -2027 -80 -1999
rect -52 -2027 -14 -1999
rect 14 -2027 52 -1999
rect 80 -2027 118 -1999
rect 146 -2027 184 -1999
rect 212 -2027 250 -1999
rect 278 -2027 316 -1999
rect 344 -2027 349 -1999
rect -349 -2065 349 -2027
rect -349 -2093 -344 -2065
rect -316 -2093 -278 -2065
rect -250 -2093 -212 -2065
rect -184 -2093 -146 -2065
rect -118 -2093 -80 -2065
rect -52 -2093 -14 -2065
rect 14 -2093 52 -2065
rect 80 -2093 118 -2065
rect 146 -2093 184 -2065
rect 212 -2093 250 -2065
rect 278 -2093 316 -2065
rect 344 -2093 349 -2065
rect -349 -2131 349 -2093
rect -349 -2159 -344 -2131
rect -316 -2159 -278 -2131
rect -250 -2159 -212 -2131
rect -184 -2159 -146 -2131
rect -118 -2159 -80 -2131
rect -52 -2159 -14 -2131
rect 14 -2159 52 -2131
rect 80 -2159 118 -2131
rect 146 -2159 184 -2131
rect 212 -2159 250 -2131
rect 278 -2159 316 -2131
rect 344 -2159 349 -2131
rect -349 -2197 349 -2159
rect -349 -2225 -344 -2197
rect -316 -2225 -278 -2197
rect -250 -2225 -212 -2197
rect -184 -2225 -146 -2197
rect -118 -2225 -80 -2197
rect -52 -2225 -14 -2197
rect 14 -2225 52 -2197
rect 80 -2225 118 -2197
rect 146 -2225 184 -2197
rect 212 -2225 250 -2197
rect 278 -2225 316 -2197
rect 344 -2225 349 -2197
rect -349 -2263 349 -2225
rect -349 -2291 -344 -2263
rect -316 -2291 -278 -2263
rect -250 -2291 -212 -2263
rect -184 -2291 -146 -2263
rect -118 -2291 -80 -2263
rect -52 -2291 -14 -2263
rect 14 -2291 52 -2263
rect 80 -2291 118 -2263
rect 146 -2291 184 -2263
rect 212 -2291 250 -2263
rect 278 -2291 316 -2263
rect 344 -2291 349 -2263
rect -349 -2329 349 -2291
rect -349 -2357 -344 -2329
rect -316 -2357 -278 -2329
rect -250 -2357 -212 -2329
rect -184 -2357 -146 -2329
rect -118 -2357 -80 -2329
rect -52 -2357 -14 -2329
rect 14 -2357 52 -2329
rect 80 -2357 118 -2329
rect 146 -2357 184 -2329
rect 212 -2357 250 -2329
rect 278 -2357 316 -2329
rect 344 -2357 349 -2329
rect -349 -2395 349 -2357
rect -349 -2423 -344 -2395
rect -316 -2423 -278 -2395
rect -250 -2423 -212 -2395
rect -184 -2423 -146 -2395
rect -118 -2423 -80 -2395
rect -52 -2423 -14 -2395
rect 14 -2423 52 -2395
rect 80 -2423 118 -2395
rect 146 -2423 184 -2395
rect 212 -2423 250 -2395
rect 278 -2423 316 -2395
rect 344 -2423 349 -2395
rect -349 -2461 349 -2423
rect -349 -2489 -344 -2461
rect -316 -2489 -278 -2461
rect -250 -2489 -212 -2461
rect -184 -2489 -146 -2461
rect -118 -2489 -80 -2461
rect -52 -2489 -14 -2461
rect 14 -2489 52 -2461
rect 80 -2489 118 -2461
rect 146 -2489 184 -2461
rect 212 -2489 250 -2461
rect 278 -2489 316 -2461
rect 344 -2489 349 -2461
rect -349 -2527 349 -2489
rect -349 -2555 -344 -2527
rect -316 -2555 -278 -2527
rect -250 -2555 -212 -2527
rect -184 -2555 -146 -2527
rect -118 -2555 -80 -2527
rect -52 -2555 -14 -2527
rect 14 -2555 52 -2527
rect 80 -2555 118 -2527
rect 146 -2555 184 -2527
rect 212 -2555 250 -2527
rect 278 -2555 316 -2527
rect 344 -2555 349 -2527
rect -349 -2593 349 -2555
rect -349 -2621 -344 -2593
rect -316 -2621 -278 -2593
rect -250 -2621 -212 -2593
rect -184 -2621 -146 -2593
rect -118 -2621 -80 -2593
rect -52 -2621 -14 -2593
rect 14 -2621 52 -2593
rect 80 -2621 118 -2593
rect 146 -2621 184 -2593
rect 212 -2621 250 -2593
rect 278 -2621 316 -2593
rect 344 -2621 349 -2593
rect -349 -2659 349 -2621
rect -349 -2687 -344 -2659
rect -316 -2687 -278 -2659
rect -250 -2687 -212 -2659
rect -184 -2687 -146 -2659
rect -118 -2687 -80 -2659
rect -52 -2687 -14 -2659
rect 14 -2687 52 -2659
rect 80 -2687 118 -2659
rect 146 -2687 184 -2659
rect 212 -2687 250 -2659
rect 278 -2687 316 -2659
rect 344 -2687 349 -2659
rect -349 -2725 349 -2687
rect -349 -2753 -344 -2725
rect -316 -2753 -278 -2725
rect -250 -2753 -212 -2725
rect -184 -2753 -146 -2725
rect -118 -2753 -80 -2725
rect -52 -2753 -14 -2725
rect 14 -2753 52 -2725
rect 80 -2753 118 -2725
rect 146 -2753 184 -2725
rect 212 -2753 250 -2725
rect 278 -2753 316 -2725
rect 344 -2753 349 -2725
rect -349 -2791 349 -2753
rect -349 -2819 -344 -2791
rect -316 -2819 -278 -2791
rect -250 -2819 -212 -2791
rect -184 -2819 -146 -2791
rect -118 -2819 -80 -2791
rect -52 -2819 -14 -2791
rect 14 -2819 52 -2791
rect 80 -2819 118 -2791
rect 146 -2819 184 -2791
rect 212 -2819 250 -2791
rect 278 -2819 316 -2791
rect 344 -2819 349 -2791
rect -349 -2857 349 -2819
rect -349 -2885 -344 -2857
rect -316 -2885 -278 -2857
rect -250 -2885 -212 -2857
rect -184 -2885 -146 -2857
rect -118 -2885 -80 -2857
rect -52 -2885 -14 -2857
rect 14 -2885 52 -2857
rect 80 -2885 118 -2857
rect 146 -2885 184 -2857
rect 212 -2885 250 -2857
rect 278 -2885 316 -2857
rect 344 -2885 349 -2857
rect -349 -2923 349 -2885
rect -349 -2951 -344 -2923
rect -316 -2951 -278 -2923
rect -250 -2951 -212 -2923
rect -184 -2951 -146 -2923
rect -118 -2951 -80 -2923
rect -52 -2951 -14 -2923
rect 14 -2951 52 -2923
rect 80 -2951 118 -2923
rect 146 -2951 184 -2923
rect 212 -2951 250 -2923
rect 278 -2951 316 -2923
rect 344 -2951 349 -2923
rect -349 -2989 349 -2951
rect -349 -3017 -344 -2989
rect -316 -3017 -278 -2989
rect -250 -3017 -212 -2989
rect -184 -3017 -146 -2989
rect -118 -3017 -80 -2989
rect -52 -3017 -14 -2989
rect 14 -3017 52 -2989
rect 80 -3017 118 -2989
rect 146 -3017 184 -2989
rect 212 -3017 250 -2989
rect 278 -3017 316 -2989
rect 344 -3017 349 -2989
rect -349 -3055 349 -3017
rect -349 -3083 -344 -3055
rect -316 -3083 -278 -3055
rect -250 -3083 -212 -3055
rect -184 -3083 -146 -3055
rect -118 -3083 -80 -3055
rect -52 -3083 -14 -3055
rect 14 -3083 52 -3055
rect 80 -3083 118 -3055
rect 146 -3083 184 -3055
rect 212 -3083 250 -3055
rect 278 -3083 316 -3055
rect 344 -3083 349 -3055
rect -349 -3121 349 -3083
rect -349 -3149 -344 -3121
rect -316 -3149 -278 -3121
rect -250 -3149 -212 -3121
rect -184 -3149 -146 -3121
rect -118 -3149 -80 -3121
rect -52 -3149 -14 -3121
rect 14 -3149 52 -3121
rect 80 -3149 118 -3121
rect 146 -3149 184 -3121
rect 212 -3149 250 -3121
rect 278 -3149 316 -3121
rect 344 -3149 349 -3121
rect -349 -3187 349 -3149
rect -349 -3215 -344 -3187
rect -316 -3215 -278 -3187
rect -250 -3215 -212 -3187
rect -184 -3215 -146 -3187
rect -118 -3215 -80 -3187
rect -52 -3215 -14 -3187
rect 14 -3215 52 -3187
rect 80 -3215 118 -3187
rect 146 -3215 184 -3187
rect 212 -3215 250 -3187
rect 278 -3215 316 -3187
rect 344 -3215 349 -3187
rect -349 -3253 349 -3215
rect -349 -3281 -344 -3253
rect -316 -3281 -278 -3253
rect -250 -3281 -212 -3253
rect -184 -3281 -146 -3253
rect -118 -3281 -80 -3253
rect -52 -3281 -14 -3253
rect 14 -3281 52 -3253
rect 80 -3281 118 -3253
rect 146 -3281 184 -3253
rect 212 -3281 250 -3253
rect 278 -3281 316 -3253
rect 344 -3281 349 -3253
rect -349 -3319 349 -3281
rect -349 -3347 -344 -3319
rect -316 -3347 -278 -3319
rect -250 -3347 -212 -3319
rect -184 -3347 -146 -3319
rect -118 -3347 -80 -3319
rect -52 -3347 -14 -3319
rect 14 -3347 52 -3319
rect 80 -3347 118 -3319
rect 146 -3347 184 -3319
rect 212 -3347 250 -3319
rect 278 -3347 316 -3319
rect 344 -3347 349 -3319
rect -349 -3385 349 -3347
rect -349 -3413 -344 -3385
rect -316 -3413 -278 -3385
rect -250 -3413 -212 -3385
rect -184 -3413 -146 -3385
rect -118 -3413 -80 -3385
rect -52 -3413 -14 -3385
rect 14 -3413 52 -3385
rect 80 -3413 118 -3385
rect 146 -3413 184 -3385
rect 212 -3413 250 -3385
rect 278 -3413 316 -3385
rect 344 -3413 349 -3385
rect -349 -3451 349 -3413
rect -349 -3479 -344 -3451
rect -316 -3479 -278 -3451
rect -250 -3479 -212 -3451
rect -184 -3479 -146 -3451
rect -118 -3479 -80 -3451
rect -52 -3479 -14 -3451
rect 14 -3479 52 -3451
rect 80 -3479 118 -3451
rect 146 -3479 184 -3451
rect 212 -3479 250 -3451
rect 278 -3479 316 -3451
rect 344 -3479 349 -3451
rect -349 -3517 349 -3479
rect -349 -3545 -344 -3517
rect -316 -3545 -278 -3517
rect -250 -3545 -212 -3517
rect -184 -3545 -146 -3517
rect -118 -3545 -80 -3517
rect -52 -3545 -14 -3517
rect 14 -3545 52 -3517
rect 80 -3545 118 -3517
rect 146 -3545 184 -3517
rect 212 -3545 250 -3517
rect 278 -3545 316 -3517
rect 344 -3545 349 -3517
rect -349 -3583 349 -3545
rect -349 -3611 -344 -3583
rect -316 -3611 -278 -3583
rect -250 -3611 -212 -3583
rect -184 -3611 -146 -3583
rect -118 -3611 -80 -3583
rect -52 -3611 -14 -3583
rect 14 -3611 52 -3583
rect 80 -3611 118 -3583
rect 146 -3611 184 -3583
rect 212 -3611 250 -3583
rect 278 -3611 316 -3583
rect 344 -3611 349 -3583
rect -349 -3649 349 -3611
rect -349 -3677 -344 -3649
rect -316 -3677 -278 -3649
rect -250 -3677 -212 -3649
rect -184 -3677 -146 -3649
rect -118 -3677 -80 -3649
rect -52 -3677 -14 -3649
rect 14 -3677 52 -3649
rect 80 -3677 118 -3649
rect 146 -3677 184 -3649
rect 212 -3677 250 -3649
rect 278 -3677 316 -3649
rect 344 -3677 349 -3649
rect -349 -3715 349 -3677
rect -349 -3743 -344 -3715
rect -316 -3743 -278 -3715
rect -250 -3743 -212 -3715
rect -184 -3743 -146 -3715
rect -118 -3743 -80 -3715
rect -52 -3743 -14 -3715
rect 14 -3743 52 -3715
rect 80 -3743 118 -3715
rect 146 -3743 184 -3715
rect 212 -3743 250 -3715
rect 278 -3743 316 -3715
rect 344 -3743 349 -3715
rect -349 -3781 349 -3743
rect -349 -3809 -344 -3781
rect -316 -3809 -278 -3781
rect -250 -3809 -212 -3781
rect -184 -3809 -146 -3781
rect -118 -3809 -80 -3781
rect -52 -3809 -14 -3781
rect 14 -3809 52 -3781
rect 80 -3809 118 -3781
rect 146 -3809 184 -3781
rect 212 -3809 250 -3781
rect 278 -3809 316 -3781
rect 344 -3809 349 -3781
rect -349 -3847 349 -3809
rect -349 -3875 -344 -3847
rect -316 -3875 -278 -3847
rect -250 -3875 -212 -3847
rect -184 -3875 -146 -3847
rect -118 -3875 -80 -3847
rect -52 -3875 -14 -3847
rect 14 -3875 52 -3847
rect 80 -3875 118 -3847
rect 146 -3875 184 -3847
rect 212 -3875 250 -3847
rect 278 -3875 316 -3847
rect 344 -3875 349 -3847
rect -349 -3913 349 -3875
rect -349 -3941 -344 -3913
rect -316 -3941 -278 -3913
rect -250 -3941 -212 -3913
rect -184 -3941 -146 -3913
rect -118 -3941 -80 -3913
rect -52 -3941 -14 -3913
rect 14 -3941 52 -3913
rect 80 -3941 118 -3913
rect 146 -3941 184 -3913
rect 212 -3941 250 -3913
rect 278 -3941 316 -3913
rect 344 -3941 349 -3913
rect -349 -3979 349 -3941
rect -349 -4007 -344 -3979
rect -316 -4007 -278 -3979
rect -250 -4007 -212 -3979
rect -184 -4007 -146 -3979
rect -118 -4007 -80 -3979
rect -52 -4007 -14 -3979
rect 14 -4007 52 -3979
rect 80 -4007 118 -3979
rect 146 -4007 184 -3979
rect 212 -4007 250 -3979
rect 278 -4007 316 -3979
rect 344 -4007 349 -3979
rect -349 -4045 349 -4007
rect -349 -4073 -344 -4045
rect -316 -4073 -278 -4045
rect -250 -4073 -212 -4045
rect -184 -4073 -146 -4045
rect -118 -4073 -80 -4045
rect -52 -4073 -14 -4045
rect 14 -4073 52 -4045
rect 80 -4073 118 -4045
rect 146 -4073 184 -4045
rect 212 -4073 250 -4045
rect 278 -4073 316 -4045
rect 344 -4073 349 -4045
rect -349 -4111 349 -4073
rect -349 -4139 -344 -4111
rect -316 -4139 -278 -4111
rect -250 -4139 -212 -4111
rect -184 -4139 -146 -4111
rect -118 -4139 -80 -4111
rect -52 -4139 -14 -4111
rect 14 -4139 52 -4111
rect 80 -4139 118 -4111
rect 146 -4139 184 -4111
rect 212 -4139 250 -4111
rect 278 -4139 316 -4111
rect 344 -4139 349 -4111
rect -349 -4177 349 -4139
rect -349 -4205 -344 -4177
rect -316 -4205 -278 -4177
rect -250 -4205 -212 -4177
rect -184 -4205 -146 -4177
rect -118 -4205 -80 -4177
rect -52 -4205 -14 -4177
rect 14 -4205 52 -4177
rect 80 -4205 118 -4177
rect 146 -4205 184 -4177
rect 212 -4205 250 -4177
rect 278 -4205 316 -4177
rect 344 -4205 349 -4177
rect -349 -4243 349 -4205
rect -349 -4271 -344 -4243
rect -316 -4271 -278 -4243
rect -250 -4271 -212 -4243
rect -184 -4271 -146 -4243
rect -118 -4271 -80 -4243
rect -52 -4271 -14 -4243
rect 14 -4271 52 -4243
rect 80 -4271 118 -4243
rect 146 -4271 184 -4243
rect 212 -4271 250 -4243
rect 278 -4271 316 -4243
rect 344 -4271 349 -4243
rect -349 -4309 349 -4271
rect -349 -4337 -344 -4309
rect -316 -4337 -278 -4309
rect -250 -4337 -212 -4309
rect -184 -4337 -146 -4309
rect -118 -4337 -80 -4309
rect -52 -4337 -14 -4309
rect 14 -4337 52 -4309
rect 80 -4337 118 -4309
rect 146 -4337 184 -4309
rect 212 -4337 250 -4309
rect 278 -4337 316 -4309
rect 344 -4337 349 -4309
rect -349 -4375 349 -4337
rect -349 -4403 -344 -4375
rect -316 -4403 -278 -4375
rect -250 -4403 -212 -4375
rect -184 -4403 -146 -4375
rect -118 -4403 -80 -4375
rect -52 -4403 -14 -4375
rect 14 -4403 52 -4375
rect 80 -4403 118 -4375
rect 146 -4403 184 -4375
rect 212 -4403 250 -4375
rect 278 -4403 316 -4375
rect 344 -4403 349 -4375
rect -349 -4441 349 -4403
rect -349 -4469 -344 -4441
rect -316 -4469 -278 -4441
rect -250 -4469 -212 -4441
rect -184 -4469 -146 -4441
rect -118 -4469 -80 -4441
rect -52 -4469 -14 -4441
rect 14 -4469 52 -4441
rect 80 -4469 118 -4441
rect 146 -4469 184 -4441
rect 212 -4469 250 -4441
rect 278 -4469 316 -4441
rect 344 -4469 349 -4441
rect -349 -4507 349 -4469
rect -349 -4535 -344 -4507
rect -316 -4535 -278 -4507
rect -250 -4535 -212 -4507
rect -184 -4535 -146 -4507
rect -118 -4535 -80 -4507
rect -52 -4535 -14 -4507
rect 14 -4535 52 -4507
rect 80 -4535 118 -4507
rect 146 -4535 184 -4507
rect 212 -4535 250 -4507
rect 278 -4535 316 -4507
rect 344 -4535 349 -4507
rect -349 -4573 349 -4535
rect -349 -4601 -344 -4573
rect -316 -4601 -278 -4573
rect -250 -4601 -212 -4573
rect -184 -4601 -146 -4573
rect -118 -4601 -80 -4573
rect -52 -4601 -14 -4573
rect 14 -4601 52 -4573
rect 80 -4601 118 -4573
rect 146 -4601 184 -4573
rect 212 -4601 250 -4573
rect 278 -4601 316 -4573
rect 344 -4601 349 -4573
rect -349 -4639 349 -4601
rect -349 -4667 -344 -4639
rect -316 -4667 -278 -4639
rect -250 -4667 -212 -4639
rect -184 -4667 -146 -4639
rect -118 -4667 -80 -4639
rect -52 -4667 -14 -4639
rect 14 -4667 52 -4639
rect 80 -4667 118 -4639
rect 146 -4667 184 -4639
rect 212 -4667 250 -4639
rect 278 -4667 316 -4639
rect 344 -4667 349 -4639
rect -349 -4705 349 -4667
rect -349 -4733 -344 -4705
rect -316 -4733 -278 -4705
rect -250 -4733 -212 -4705
rect -184 -4733 -146 -4705
rect -118 -4733 -80 -4705
rect -52 -4733 -14 -4705
rect 14 -4733 52 -4705
rect 80 -4733 118 -4705
rect 146 -4733 184 -4705
rect 212 -4733 250 -4705
rect 278 -4733 316 -4705
rect 344 -4733 349 -4705
rect -349 -4771 349 -4733
rect -349 -4799 -344 -4771
rect -316 -4799 -278 -4771
rect -250 -4799 -212 -4771
rect -184 -4799 -146 -4771
rect -118 -4799 -80 -4771
rect -52 -4799 -14 -4771
rect 14 -4799 52 -4771
rect 80 -4799 118 -4771
rect 146 -4799 184 -4771
rect 212 -4799 250 -4771
rect 278 -4799 316 -4771
rect 344 -4799 349 -4771
rect -349 -4837 349 -4799
rect -349 -4865 -344 -4837
rect -316 -4865 -278 -4837
rect -250 -4865 -212 -4837
rect -184 -4865 -146 -4837
rect -118 -4865 -80 -4837
rect -52 -4865 -14 -4837
rect 14 -4865 52 -4837
rect 80 -4865 118 -4837
rect 146 -4865 184 -4837
rect 212 -4865 250 -4837
rect 278 -4865 316 -4837
rect 344 -4865 349 -4837
rect -349 -4903 349 -4865
rect -349 -4931 -344 -4903
rect -316 -4931 -278 -4903
rect -250 -4931 -212 -4903
rect -184 -4931 -146 -4903
rect -118 -4931 -80 -4903
rect -52 -4931 -14 -4903
rect 14 -4931 52 -4903
rect 80 -4931 118 -4903
rect 146 -4931 184 -4903
rect 212 -4931 250 -4903
rect 278 -4931 316 -4903
rect 344 -4931 349 -4903
rect -349 -4969 349 -4931
rect -349 -4997 -344 -4969
rect -316 -4997 -278 -4969
rect -250 -4997 -212 -4969
rect -184 -4997 -146 -4969
rect -118 -4997 -80 -4969
rect -52 -4997 -14 -4969
rect 14 -4997 52 -4969
rect 80 -4997 118 -4969
rect 146 -4997 184 -4969
rect 212 -4997 250 -4969
rect 278 -4997 316 -4969
rect 344 -4997 349 -4969
rect -349 -5035 349 -4997
rect -349 -5063 -344 -5035
rect -316 -5063 -278 -5035
rect -250 -5063 -212 -5035
rect -184 -5063 -146 -5035
rect -118 -5063 -80 -5035
rect -52 -5063 -14 -5035
rect 14 -5063 52 -5035
rect 80 -5063 118 -5035
rect 146 -5063 184 -5035
rect 212 -5063 250 -5035
rect 278 -5063 316 -5035
rect 344 -5063 349 -5035
rect -349 -5068 349 -5063
<< end >>
