magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2083 -9815 10992 5035
<< isosubstrate >>
rect 2390 -6738 8471 -6737
rect 5759 -7815 8471 -6738
<< nwell >>
rect -83 53 8471 3035
rect 5925 -7651 7121 -6737
<< nsubdiff >>
rect 8234 2930 8388 2952
rect 8234 2862 8320 2930
rect 8298 2696 8320 2862
rect 8366 2696 8388 2930
rect 8298 2272 8388 2696
rect 8298 226 8320 2272
rect 8234 158 8320 226
rect 8366 158 8388 2272
rect 8234 136 8388 158
<< nsubdiffcont >>
rect 8320 2696 8366 2930
rect 8320 158 8366 2272
<< polysilicon >>
rect 6922 -7404 7092 -7264
rect 7477 -7404 7774 -7264
<< metal1 >>
rect 79 2873 165 2941
rect 8223 2930 8377 2941
rect 8223 2873 8320 2930
rect 8309 2696 8320 2873
rect 8366 2696 8377 2930
rect 8309 2669 8377 2696
rect 406 2166 474 2602
rect 7678 2446 8992 2602
rect 406 1606 474 2042
rect 7678 1886 7746 2322
rect 8309 2272 8377 2338
rect 406 1046 474 1482
rect 7678 1326 7746 1762
rect 406 486 474 922
rect 7678 766 7746 1202
rect 8309 215 8320 2272
rect 79 147 165 215
rect 8223 158 8320 215
rect 8366 158 8377 2272
rect 8223 147 8377 158
rect 6019 -7113 6087 -7027
rect 8309 -7113 8377 -7027
rect 6019 -7250 6878 -7174
rect 7818 -7250 8377 -7174
rect 6278 -7494 8118 -7418
rect 8309 -7643 8377 -7440
rect 8836 -7516 8992 2446
<< metal2 >>
rect 7938 -7516 8992 -7440
use M1_NWELL_CDNS_40661953145231  M1_NWELL_CDNS_40661953145231_0
timestamp 1713338890
transform 1 0 45 0 -1 1544
box -128 -1491 128 1491
use M1_NWELL_CDNS_40661953145273  M1_NWELL_CDNS_40661953145273_0
timestamp 1713338890
transform 0 -1 6053 -1 0 -7335
box -316 -128 316 128
use M1_NWELL_CDNS_40661953145315  M1_NWELL_CDNS_40661953145315_0
timestamp 1713338890
transform 0 -1 6523 -1 0 -6993
box -128 -598 128 598
use M1_NWELL_CDNS_40661953145316  M1_NWELL_CDNS_40661953145316_0
timestamp 1713338890
transform 1 0 4194 0 -1 181
box -4123 -128 4123 128
use M1_NWELL_CDNS_40661953145316  M1_NWELL_CDNS_40661953145316_1
timestamp 1713338890
transform 1 0 4194 0 -1 2907
box -4123 -128 4123 128
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_0
timestamp 1713338890
transform 0 -1 7003 1 0 -7334
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_1
timestamp 1713338890
transform 0 -1 7566 1 0 -7334
box -42 -89 42 89
use M1_PSUB_CDNS_69033583165609  M1_PSUB_CDNS_69033583165609_0
timestamp 1713338890
transform 0 1 7873 -1 0 -7677
box -45 -515 45 515
use M1_PSUB_CDNS_69033583165609  M1_PSUB_CDNS_69033583165609_1
timestamp 1713338890
transform 0 1 7873 -1 0 -6993
box -45 -515 45 515
use M1_PSUB_CDNS_69033583165621  M1_PSUB_CDNS_69033583165621_0
timestamp 1713338890
transform 0 1 8343 -1 0 -7335
box -233 -45 233 45
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_0
timestamp 1713338890
transform 1 0 8028 0 1 -7478
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_1
timestamp 1713338890
transform 1 0 8902 0 1 -7478
box -90 -38 90 38
use nmos_6p0_CDNS_4066195314530  nmos_6p0_CDNS_4066195314530_0
timestamp 1713338890
transform 0 -1 8118 -1 0 -7264
box -88 -44 228 344
use pmos_6p0_CDNS_4066195314512  pmos_6p0_CDNS_4066195314512_0
timestamp 1713338890
transform 0 -1 6878 -1 0 -7264
box -208 -120 348 720
use ppolyf_u_CDNS_4066195314532  ppolyf_u_CDNS_4066195314532_0
timestamp 1713338890
transform -1 0 5208 0 1 484
box 0 0 4804 160
use ppolyf_u_CDNS_4066195314533  ppolyf_u_CDNS_4066195314533_0
timestamp 1713338890
transform 1 0 404 0 1 764
box 0 0 7344 160
use ppolyf_u_CDNS_4066195314533  ppolyf_u_CDNS_4066195314533_1
timestamp 1713338890
transform -1 0 7748 0 1 1044
box 0 0 7344 160
use ppolyf_u_CDNS_4066195314533  ppolyf_u_CDNS_4066195314533_2
timestamp 1713338890
transform 1 0 404 0 1 1324
box 0 0 7344 160
use ppolyf_u_CDNS_4066195314533  ppolyf_u_CDNS_4066195314533_3
timestamp 1713338890
transform 1 0 404 0 1 2444
box 0 0 7344 160
use ppolyf_u_CDNS_4066195314533  ppolyf_u_CDNS_4066195314533_4
timestamp 1713338890
transform 1 0 404 0 1 2164
box 0 0 7344 160
use ppolyf_u_CDNS_4066195314533  ppolyf_u_CDNS_4066195314533_5
timestamp 1713338890
transform 1 0 404 0 1 1884
box 0 0 7344 160
use ppolyf_u_CDNS_4066195314533  ppolyf_u_CDNS_4066195314533_6
timestamp 1713338890
transform -1 0 7748 0 1 1604
box 0 0 7344 160
<< labels >>
rlabel metal1 s 7561 -7333 7561 -7333 4 PD
port 1 nsew
rlabel metal1 s 7110 -7333 7110 -7333 4 PU_B
port 2 nsew
rlabel metal1 s 8343 -7192 8343 -7192 4 DVSS
port 3 nsew
rlabel metal1 s 6048 -7005 6048 -7005 4 DVDD
port 4 nsew
rlabel metal1 s 5175 575 5175 575 4 A
port 5 nsew
<< end >>
