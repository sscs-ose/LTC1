magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -9001 -2045 9001 2045
<< psubdiff >>
rect -7001 23 7001 45
rect -7001 -23 -6979 23
rect 6979 -23 7001 23
rect -7001 -45 7001 -23
<< psubdiffcont >>
rect -6979 -23 6979 23
<< metal1 >>
rect -6990 23 6990 34
rect -6990 -23 -6979 23
rect 6979 -23 6990 23
rect -6990 -34 6990 -23
<< end >>
