* NGSPICE file created from CLK_div_108_mag_flat.ext - technology: gf180mcuC

.subckt pex_CLK_div_108_mag VSS VDD RST Vdiv108 CLK
X0 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_2.JK_FF_mag_1.K.t3 a_10058_1318# VSS.t247 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1 a_8733_1362# CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t221 VSS.t220 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 a_8169_1362# VSS.t125 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X3 VSS JK_FF_mag_0.nand2_mag_1.IN2 a_9803_3948# VSS.t105 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X4 a_2486_1354# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t149 VSS.t148 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X5 a_7759_221# RST.t0 a_7599_221# VSS.t217 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X6 a_3805_213# CLK_div_3_mag_0.CLK.t2 a_3645_213# VSS.t195 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X7 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_2.Q1 VDD.t101 VDD.t100 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X8 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_1512_213# VSS.t241 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X9 VDD CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VDD.t202 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X10 VDD JK_FF_mag_1.QB JK_FF_mag_1.nand3_mag_0.OUT VDD.t151 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X11 a_10058_1318# CLK_div_3_mag_2.CLK.t2 a_9898_1318# VSS.t216 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X12 a_5118_3858# CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VSS.t113 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X13 a_8169_1362# CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t270 VSS.t269 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X14 a_8320_2831# JK_FF_mag_1.QB JK_FF_mag_1.nand3_mag_0.OUT VSS.t91 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X15 VDD CLK_div_3_mag_2.CLK.t3 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT VDD.t356 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X16 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VDD.t3 VDD.t2 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X17 VSS JK_FF_mag_0.CLK JK_FF_mag_0.nand2_mag_3.IN1 VSS.t18 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X18 a_2640_257# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t151 VSS.t150 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X19 a_3836_4955# CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t1 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X20 VSS CLK.t0 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VSS.t114 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X21 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD.t420 VDD.t419 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X22 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_2.Q1 VDD.t99 VDD.t98 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X23 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t415 VDD.t414 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X24 VDD CLK_div_3_mag_0.CLK.t3 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t184 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X25 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t117 VDD.t116 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X26 a_1537_3858# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t0 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X27 VDD Vdiv108.t3 JK_FF_mag_1.nand3_mag_2.OUT VDD.t130 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X28 VDD VDD.t295 JK_FF_mag_0.nand3_mag_0.OUT VDD.t24 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X29 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t349 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X30 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_2.Q1 a_7035_221# VSS.t57 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X31 a_8326_3928# Vdiv108.t4 JK_FF_mag_1.nand3_mag_2.OUT VSS.t30 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X32 VSS VDD.t437 a_11655_3948# VSS.t165 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X33 VDD RST.t1 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT VDD.t70 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X34 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VDD.t306 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X35 CLK_div_3_mag_2.or_2_mag_0.IN2 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN VDD.t8 VDD.t7 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X36 a_4400_4955# CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VSS.t186 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X37 VDD CLK_div_3_mag_1.Q1.t3 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VDD.t255 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X38 VDD CLK_div_3_mag_1.JK_FF_mag_1.K.t2 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VDD.t258 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X39 VDD CLK_div_3_mag_0.JK_FF_mag_1.K.t3 CLK_div_3_mag_0.Q0 VDD.t366 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X40 a_5124_4955# CLK_div_3_mag_1.Q1.t4 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VSS.t157 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X41 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_2.CLK.t4 VDD.t359 VDD.t7 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X42 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t168 VDD.t167 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X43 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.CLK.t4 VSS.t146 VSS.t145 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X44 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT a_10622_1362# VSS.t74 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X45 a_2101_3858# CLK_div_3_mag_1.JK_FF_mag_1.K.t3 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VSS.t113 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X46 VDD CLK_div_3_mag_2.CLK.t5 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT VDD.t80 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X47 a_10052_221# CLK_div_3_mag_2.CLK.t6 a_9892_221# VSS.t44 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X48 VDD CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.CLK.t0 VDD.t252 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X49 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t355 VDD.t354 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X50 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD.t324 VDD.t323 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X51 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.JK_FF_mag_1.K.t4 VDD.t235 VDD.t234 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X52 VDD VDD.t291 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VDD.t292 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X53 VSS CLK.t1 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VSS.t117 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X54 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 a_7759_221# VSS.t268 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X55 a_9898_1318# CLK_div_3_mag_2.Q1 VSS.t56 VSS.t55 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X56 VSS VDD.t439 a_2267_4955# VSS.t168 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X57 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT RST.t2 VDD.t69 VDD.t68 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X58 a_409_3858# CLK_div_3_mag_1.JK_FF_mag_1.K.t5 CLK_div_3_mag_1.Q0.t1 VSS.t0 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X59 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_2.CLK.t7 VDD.t84 VDD.t83 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X60 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_2.JK_FF_mag_1.K.t4 VDD.t403 VDD.t402 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X61 VDD CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t334 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X62 a_3811_1310# CLK_div_3_mag_0.CLK.t5 a_3651_1310# VSS.t147 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X63 a_1352_213# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS.t67 VSS.t66 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X64 VDD CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_3_mag_2.Q1 VDD.t104 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X65 CLK_div_3_mag_2.Q0 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t338 VDD.t337 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X66 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 a_11340_265# VSS.t199 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X67 a_1543_4955# RST.t3 a_1383_4955# VSS.t218 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X68 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_2.JK_FF_mag_1.QB VDD.t103 VDD.t102 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X69 CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_2.Q0 a_11307_2697# VDD.t9 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X70 JK_FF_mag_0.CLK CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN VDD.t330 VDD.t329 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X71 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT VDD.t120 VDD.t119 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X72 a_10776_221# RST.t4 a_10616_221# VSS.t219 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X73 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_2.Q0 VDD.t408 VDD.t407 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X74 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK.t2 VDD.t198 VDD.t197 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X75 a_2267_4955# CLK.t3 a_2107_4955# VSS.t120 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X76 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD.t424 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X77 VSS CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.CLK.t1 VSS.t162 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X78 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t79 VDD.t78 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X79 a_1383_4955# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VSS.t276 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X80 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t416 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X81 a_7041_1318# CLK_div_3_mag_2.CLK.t8 a_6881_1318# VSS.t45 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X82 CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t230 VDD.t229 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X83 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_4529_213# VSS.t215 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X84 VSS CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_819_4955# VSS.t271 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X85 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_1.K.t1 VDD.t429 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X86 VDD CLK_div_3_mag_1.or_2_mag_0.IN2 a_852_2291# VDD.t300 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X87 VDD CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_1.QB VDD.t382 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X88 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t77 VDD.t76 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X89 VSS CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_255_4955# VSS.t279 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X90 JK_FF_mag_0.Q JK_FF_mag_0.QB VDD.t222 VDD.t221 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X91 a_6881_1318# CLK_div_3_mag_2.JK_FF_mag_1.K.t5 VSS.t246 VSS.t245 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X92 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_2.JK_FF_mag_1.QB a_7041_1318# VSS.t59 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X93 a_9803_3948# JK_FF_mag_0.QB JK_FF_mag_0.Q.t1 VSS.t127 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X94 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_2.Q0 a_10052_221# VSS.t252 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X95 VSS CLK.t4 a_1825_2759# VSS.t121 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X96 VDD CLK_div_3_mag_0.CLK.t6 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t181 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X97 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t374 VDD.t373 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X98 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t317 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X99 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_4375_1354# VSS.t212 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X100 VSS CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN VSS.t181 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X101 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.Q0 VDD.t18 VDD.t17 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X102 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT VDD.t166 VDD.t165 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X103 VSS CLK_div_3_mag_2.Q0 CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN VSS.t249 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X104 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_1.K.t4 a_5503_1354# VSS.t226 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X105 VDD JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand2_mag_1.IN2 VDD.t24 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X106 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.CLK.t7 VDD.t180 VDD.t179 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X107 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t353 VDD.t352 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X108 a_4375_1354# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS.t102 VSS.t101 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X109 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 a_10776_221# VSS.t43 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X110 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand3_mag_1.OUT VDD.t228 VDD.t24 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X111 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_2.Q1 a_10334_2461# VSS.t54 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X112 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.Q1 VDD.t381 VDD.t380 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X113 VSS JK_FF_mag_0.nand3_mag_1.IN1 a_10367_3948# VSS.t109 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X114 a_10931_3948# JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.IN1 VSS.t140 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X115 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.Q0 a_5060_2689# VDD.t16 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X116 a_2076_257# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS.t194 VSS.t193 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X117 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.CLK VDD.t25 VDD.t24 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X118 a_11655_3948# JK_FF_mag_0.CLK a_11495_3948# VSS.t17 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X119 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_1.Q1.t2 VDD.t409 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X120 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_0.nand2_mag_3.IN1 VDD.t28 VDD.t24 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X121 VDD JK_FF_mag_1.nand2_mag_1.IN2 Vdiv108.t0 VDD.t140 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X122 a_788_213# CLK_div_3_mag_0.CLK.t8 a_628_213# VSS.t89 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X123 VDD CLK_div_3_mag_2.Q1 CLK_div_3_mag_2.JK_FF_mag_1.QB VDD.t95 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X124 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VDD.t1 VDD.t0 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X125 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_1.Q0.t3 VSS.t61 VSS.t60 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X126 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t37 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X127 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_2.CLK.t9 VSS.t47 VSS.t46 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X128 VSS CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_3426_3858# VSS.t0 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X129 a_3990_3858# CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t0 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X130 a_10367_3948# JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand2_mag_1.IN2 VSS.t22 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X131 VDD JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.nand3_mag_1.IN1 VDD.t24 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X132 a_5060_2689# CLK_div_3_mag_0.or_2_mag_0.IN2 VDD.t118 VDD.t16 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X133 VSS JK_FF_mag_1.nand2_mag_1.IN2 a_6628_2831# VSS.t79 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X134 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t41 VDD.t40 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X135 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t348 VDD.t347 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X136 CLK_div_3_mag_2.Q0 CLK_div_3_mag_2.JK_FF_mag_1.K.t6 a_11750_1362# VSS.t244 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X137 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t394 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X138 VDD JK_FF_mag_0.QB JK_FF_mag_0.nand3_mag_0.OUT VDD.t24 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X139 a_10622_1362# CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT VSS.t223 VSS.t222 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X140 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT a_7605_1362# VSS.t100 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X141 VSS CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_4554_3858# VSS.t0 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X142 VSS JK_FF_mag_0.nand3_mag_0.OUT a_10931_3948# VSS.t204 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X143 a_11495_3948# JK_FF_mag_0.QB JK_FF_mag_0.nand3_mag_0.OUT VSS.t126 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X144 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.Q0 a_3805_213# VSS.t15 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X145 VDD VDD.t287 JK_FF_mag_0.nand3_mag_2.OUT VDD.t288 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X146 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t320 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X147 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t393 VDD.t392 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X148 a_3651_1310# CLK_div_3_mag_0.Q1 VSS.t236 VSS.t235 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X149 a_8887_265# CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t142 VSS.t141 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X150 VDD CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t216 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X151 CLK_div_3_mag_2.Q1 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t361 VDD.t360 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X152 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t428 VDD.t427 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X153 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.Q1 VDD.t379 VDD.t378 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X154 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT VDD.t299 VDD.t298 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X155 VDD JK_FF_mag_1.nand3_mag_2.OUT JK_FF_mag_1.nand3_mag_1.OUT VDD.t339 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X156 a_11307_2697# CLK_div_3_mag_2.or_2_mag_0.IN2 VDD.t10 VDD.t9 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X157 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.Q1 a_2640_257# VSS.t234 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X158 VDD CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_1.K.t0 VDD.t13 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X159 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t284 VDD.t286 VDD.t285 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X160 VDD CLK_div_3_mag_1.Q0.t4 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VDD.t107 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X161 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.CLK VDD.t23 VDD.t22 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X162 VDD JK_FF_mag_1.nand2_mag_4.IN2 JK_FF_mag_1.QB VDD.t231 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X163 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t49 VDD.t48 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X164 a_2107_4955# CLK_div_3_mag_1.Q0.t5 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VSS.t62 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X165 VDD JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand2_mag_4.IN2 VDD.t225 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X166 VSS JK_FF_mag_1.nand3_mag_2.OUT a_7762_3928# VSS.t30 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X167 VDD RST.t5 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD.t65 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X168 VSS JK_FF_mag_1.nand2_mag_4.IN2 a_6474_3928# VSS.t77 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X169 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.QB VDD.t388 VDD.t387 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X170 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t314 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X171 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t413 VDD.t412 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X172 VSS VDD.t441 a_11661_5045# VSS.t171 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X173 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VDD.t435 VDD.t434 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X174 JK_FF_mag_1.nand3_mag_1.OUT RST.t6 VDD.t64 VDD.t63 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X175 a_7762_3928# RST.t7 a_7602_3928# VSS.t30 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X176 JK_FF_mag_1.QB Vdiv108.t5 VDD.t196 VDD.t195 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X177 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT VDD.t125 VDD.t124 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X178 a_819_4955# CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t282 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X179 a_5657_257# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t231 VSS.t230 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X180 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_2076_257# VSS.t191 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X181 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.Q0.t6 VDD.t111 VDD.t110 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X182 a_6474_3928# Vdiv108.t6 JK_FF_mag_1.QB VSS.t77 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X183 a_852_2291# CLK_div_3_mag_1.Q0.t7 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN VDD.t112 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X184 VDD CLK_div_3_mag_0.CLK.t9 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t176 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X185 a_11661_5045# JK_FF_mag_0.CLK a_11501_5045# VSS.t16 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X186 JK_FF_mag_0.CLK CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN VSS.t197 VSS.t196 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X187 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t12 VDD.t11 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X188 a_255_4955# CLK_div_3_mag_1.Q0.t8 CLK_div_3_mag_1.JK_FF_mag_1.K VSS.t63 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X189 VSS JK_FF_mag_0.nand3_mag_1.OUT a_10213_5045# VSS.t137 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X190 a_8323_265# CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT VSS.t99 VSS.t98 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X191 a_7599_221# CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT VSS.t180 VSS.t179 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X192 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.Q1 a_788_213# VSS.t233 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X193 a_3645_213# VDD.t442 VSS.t175 VSS.t174 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X194 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t34 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X195 VDD CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t375 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X196 a_1825_2759# CLK_div_3_mag_1.Q1.t5 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN VSS.t158 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X197 VDD CLK.t5 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN VDD.t199 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X198 a_4939_1354# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t214 VSS.t213 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X199 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t241 VDD.t240 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X200 a_1512_213# RST.t8 a_1352_213# VSS.t128 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X201 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.QB a_794_1310# VSS.t238 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X202 VDD CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t121 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X203 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.or_2_mag_0.IN2 VSS.t69 VSS.t68 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X204 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.CLK.t10 VDD.t175 VDD.t174 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X205 CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_3_mag_2.Q1 a_8887_265# VSS.t53 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X206 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_4939_1354# VSS.t27 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X207 VDD JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.QB VDD.t50 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X208 a_794_1310# CLK_div_3_mag_0.CLK.t11 a_634_1310# VSS.t132 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X209 a_5503_1354# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t29 VSS.t28 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X210 a_5093_257# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS.t211 VSS.t210 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X211 a_4369_213# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS.t10 VSS.t9 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X212 VDD CLK_div_3_mag_2.Q0 CLK_div_3_mag_2.JK_FF_mag_1.K.t1 VDD.t404 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X213 a_10334_2461# CLK_div_3_mag_2.CLK.t10 VSS.t49 VSS.t48 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X214 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.CLK.t12 VSS.t134 VSS.t133 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X215 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT VDD.t281 VDD.t283 VDD.t282 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X216 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT VDD.t224 VDD.t223 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X217 VDD JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_1.nand3_mag_1.IN1 VDD.t154 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X218 CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_2.or_2_mag_0.IN2 VSS.t8 VSS.t7 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X219 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_1358_1354# VSS.t192 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X220 Vdiv108 JK_FF_mag_1.QB VDD.t150 VDD.t149 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X221 a_1922_1354# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t240 VSS.t239 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X222 VSS JK_FF_mag_0.nand2_mag_4.IN2 a_9649_5045# VSS.t36 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X223 VDD CLK_div_3_mag_1.JK_FF_mag_1.K.t6 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VDD.t202 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X224 VDD JK_FF_mag_0.CLK JK_FF_mag_0.nand2_mag_3.IN1 VDD.t19 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X225 VSS JK_FF_mag_1.nand3_mag_0.OUT a_7756_2831# VSS.t92 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X226 VDD VDD.t277 JK_FF_mag_1.nand3_mag_0.OUT VDD.t278 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X227 a_11904_265# CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t278 VSS.t277 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X228 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 a_11186_1362# VSS.t198 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X229 a_3426_3858# CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.Q1.t0 VSS.t0 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X230 VSS CLK_div_3_mag_1.JK_FF_mag_1.K.t7 a_5278_3858# VSS.t113 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X231 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t303 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X232 VDD CLK.t6 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VDD.t202 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X233 a_6628_2831# JK_FF_mag_1.QB Vdiv108.t1 VSS.t90 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X234 VDD JK_FF_mag_0.Q.t3 JK_FF_mag_1.nand2_mag_3.IN1 VDD.t137 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X235 a_11750_1362# CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t201 VSS.t200 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X236 CLK_div_3_mag_2.Q1 CLK_div_3_mag_2.JK_FF_mag_1.QB a_8733_1362# VSS.t58 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X237 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VDD.t313 VDD.t312 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X238 VSS VDD.t444 a_8480_2831# VSS.t176 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X239 CLK_div_3_mag_2.or_2_mag_0.IN2 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN VSS.t6 VSS.t5 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X240 VDD JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand2_mag_1.IN2 VDD.t45 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X241 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.Q0 a_5657_257# VSS.t14 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X242 a_7605_1362# CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT VSS.t71 VSS.t70 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X243 VSS CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_3990_3858# VSS.t0 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X244 a_4554_3858# CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t0 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X245 VSS JK_FF_mag_1.nand3_mag_1.IN1 a_7192_2831# VSS.t31 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X246 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand3_mag_1.OUT VDD.t161 VDD.t160 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X247 a_1358_1354# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS.t35 VSS.t34 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X248 JK_FF_mag_0.nand3_mag_1.OUT RST.t9 VDD.t61 VDD.t60 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X249 VDD RST.t10 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t58 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X250 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK.t7 VDD.t205 VDD.t202 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X251 a_7756_2831# JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand3_mag_1.IN1 VSS.t97 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X252 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_0.Q.t4 VDD.t33 VDD.t32 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X253 VDD CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.Q1 VDD.t385 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X254 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_1922_1354# VSS.t190 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X255 a_11186_1362# CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t42 VSS.t41 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X256 a_5278_3858# CLK.t8 a_5118_3858# VSS.t113 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X257 JK_FF_mag_1.nand2_mag_1.IN2 JK_FF_mag_1.nand2_mag_3.IN1 VDD.t136 VDD.t135 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X258 a_8480_2831# JK_FF_mag_0.Q.t5 a_8320_2831# VSS.t85 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X259 JK_FF_mag_1.nand2_mag_4.IN2 JK_FF_mag_1.nand2_mag_3.IN1 VDD.t134 VDD.t133 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X260 a_7192_2831# JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.nand2_mag_1.IN2 VSS.t78 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X261 a_11340_265# CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT VSS.t73 VSS.t72 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X262 a_6875_221# VDD.t445 VSS.t258 VSS.t257 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X263 VDD CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t213 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X264 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t309 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X265 VDD JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand3_mag_1.OUT VDD.t190 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X266 VDD VDD.t273 JK_FF_mag_1.nand3_mag_2.OUT VDD.t274 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X267 VSS JK_FF_mag_0.Q.t6 JK_FF_mag_1.nand2_mag_3.IN1 VSS.t86 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X268 a_10616_221# CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT VSS.t136 VSS.t135 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X269 VSS CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_3836_4955# VSS.t187 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X270 a_7038_3928# JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.nand2_mag_4.IN2 VSS.t77 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X271 VSS VDD.t447 a_8486_3928# VSS.t30 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X272 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t237 VDD.t236 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X273 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_2.CLK.t11 VSS.t51 VSS.t50 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X274 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VDD.t143 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X275 VDD JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.nand3_mag_1.OUT VDD.t344 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X276 VDD JK_FF_mag_0.Q.t7 JK_FF_mag_0.nand3_mag_2.OUT VDD.t146 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X277 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t113 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X278 VSS CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_4560_4955# VSS.t82 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X279 a_10937_5045# RST.t11 a_10777_5045# VSS.t129 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X280 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_1.QB VDD.t4 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X281 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand2_mag_3.IN1 VDD.t27 VDD.t26 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X282 VSS CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS.t11 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X283 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.K.t5 VDD.t370 VDD.t369 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X284 VDD VDD.t269 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VDD.t270 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X285 VSS CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_1537_3858# VSS.t0 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X286 VDD CLK_div_3_mag_1.Q1.t6 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VDD.t245 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X287 JK_FF_mag_1.nand3_mag_2.OUT JK_FF_mag_0.Q.t8 VDD.t127 VDD.t126 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X288 VSS CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_3272_4955# VSS.t2 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X289 VDD CLK.t9 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VDD.t206 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X290 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_2.CLK.t12 VDD.t86 VDD.t85 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X291 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_5093_257# VSS.t26 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X292 VSS VDD.t449 a_5284_4955# VSS.t261 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X293 VSS CLK_div_3_mag_1.Q1.t7 a_2261_3858# VSS.t113 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X294 a_8486_3928# JK_FF_mag_0.Q.t9 a_8326_3928# VSS.t30 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X295 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t421 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X296 VDD JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand2_mag_4.IN2 VDD.t157 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X297 VDD JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand3_mag_1.OUT VDD.t42 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X298 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.Q1 a_4087_2453# VSS.t232 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X299 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT RST.t12 VDD.t57 VDD.t56 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X300 VSS CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_973_3858# VSS.t0 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X301 VSS JK_FF_mag_1.nand3_mag_1.OUT a_7038_3928# VSS.t77 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X302 a_7602_3928# JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand3_mag_1.OUT VSS.t30 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X303 a_4529_213# RST.t13 a_4369_213# VSS.t130 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X304 a_4560_4955# RST.t14 a_4400_4955# VSS.t131 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X305 a_10777_5045# JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand3_mag_1.OUT VSS.t108 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X306 CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.Q1.t8 VDD.t249 VDD.t248 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X307 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.CLK.t13 VDD.t173 VDD.t172 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X308 VDD CLK_div_3_mag_2.CLK.t13 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT VDD.t87 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X309 a_3272_4955# CLK_div_3_mag_1.Q1.t9 CLK_div_3_mag_1.JK_FF_mag_1.QB VSS.t161 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X310 VSS JK_FF_mag_0.nand3_mag_2.OUT a_10937_5045# VSS.t207 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X311 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK.t10 VDD.t210 VDD.t209 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X312 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK.t11 VDD.t212 VDD.t211 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X313 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.K.t6 VDD.t372 VDD.t371 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X314 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t239 VDD.t238 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X315 a_5284_4955# CLK.t12 a_5124_4955# VSS.t112 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X316 a_11501_5045# JK_FF_mag_0.Q.t10 JK_FF_mag_0.nand3_mag_2.OUT VSS.t75 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X317 VDD CLK_div_3_mag_2.Q1 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN VDD.t7 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X318 a_10213_5045# JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand2_mag_4.IN2 VSS.t21 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X319 a_2261_3858# CLK.t13 a_2101_3858# VSS.t113 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X320 a_4087_2453# CLK_div_3_mag_0.CLK.t14 VSS.t104 VSS.t103 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X321 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_1.Q0.t0 VDD.t73 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X322 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VDD.t433 VDD.t432 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X323 VDD CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_1.or_2_mag_0.IN2 VDD.t242 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X324 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_1.Q1.t10 VDD.t251 VDD.t250 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X325 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.Q0 a_11904_265# VSS.t248 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X326 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD.t29 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X327 VSS CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 a_409_3858# VSS.t0 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X328 a_973_3858# CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t0 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X329 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.K.t7 a_3811_1310# VSS.t227 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X330 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT VDD.t266 VDD.t268 VDD.t267 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X331 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t263 VDD.t265 VDD.t264 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X332 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_2.JK_FF_mag_1.K.t7 VDD.t400 VDD.t399 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X333 VDD CLK_div_3_mag_2.JK_FF_mag_1.K.t8 CLK_div_3_mag_2.Q0 VDD.t397 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X334 VSS CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_1543_4955# VSS.t23 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X335 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS.t153 VSS.t152 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X336 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT VDD.t363 VDD.t362 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X337 VDD RST.t15 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT VDD.t53 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X338 VDD CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t162 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X339 VDD CLK_div_3_mag_0.CLK.t15 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t169 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X340 a_7035_221# CLK_div_3_mag_2.CLK.t14 a_6875_221# VSS.t52 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X341 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t391 VDD.t390 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X342 JK_FF_mag_0.QB JK_FF_mag_0.Q.t11 VDD.t129 VDD.t128 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X343 VDD CLK_div_3_mag_2.CLK.t15 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT VDD.t90 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X344 a_634_1310# CLK_div_3_mag_0.JK_FF_mag_1.K.t8 VSS.t229 VSS.t228 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X345 VSS CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_1.or_2_mag_0.IN2 VSS.t154 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X346 VDD CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t331 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X347 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_1.QB a_2486_1354# VSS.t237 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X348 a_9892_221# VDD.t450 VSS.t265 VSS.t264 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X349 a_628_213# VDD.t451 VSS.t267 VSS.t266 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X350 a_9649_5045# JK_FF_mag_0.Q.t12 JK_FF_mag_0.QB VSS.t76 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X351 VDD JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_0.Q.t0 VDD.t187 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X352 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 a_8323_265# VSS.t124 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
R0 CLK_div_3_mag_2.JK_FF_mag_1.K.n4 CLK_div_3_mag_2.JK_FF_mag_1.K.t3 37.1986
R1 CLK_div_3_mag_2.JK_FF_mag_1.K.n3 CLK_div_3_mag_2.JK_FF_mag_1.K.t6 31.528
R2 CLK_div_3_mag_2.JK_FF_mag_1.K.n2 CLK_div_3_mag_2.JK_FF_mag_1.K.t4 30.5184
R3 CLK_div_3_mag_2.JK_FF_mag_1.K.n2 CLK_div_3_mag_2.JK_FF_mag_1.K.t5 24.7029
R4 CLK_div_3_mag_2.JK_FF_mag_1.K.n4 CLK_div_3_mag_2.JK_FF_mag_1.K.t7 17.6614
R5 CLK_div_3_mag_2.JK_FF_mag_1.K.n3 CLK_div_3_mag_2.JK_FF_mag_1.K.t8 15.3826
R6 CLK_div_3_mag_2.JK_FF_mag_1.K.n0 CLK_div_3_mag_2.JK_FF_mag_1.K 12.0843
R7 CLK_div_3_mag_2.JK_FF_mag_1.K.n0 CLK_div_3_mag_2.JK_FF_mag_1.K.n3 9.86691
R8 CLK_div_3_mag_2.JK_FF_mag_1.K.n5 CLK_div_3_mag_2.JK_FF_mag_1.K 6.09789
R9 CLK_div_3_mag_2.JK_FF_mag_1.K.n1 CLK_div_3_mag_2.JK_FF_mag_1.K.n7 2.99416
R10 CLK_div_3_mag_2.JK_FF_mag_1.K.n7 CLK_div_3_mag_2.JK_FF_mag_1.K.t1 2.2755
R11 CLK_div_3_mag_2.JK_FF_mag_1.K.n7 CLK_div_3_mag_2.JK_FF_mag_1.K.n6 2.2755
R12 CLK_div_3_mag_2.JK_FF_mag_1.K.n1 CLK_div_3_mag_2.JK_FF_mag_1.K.n5 2.2505
R13 CLK_div_3_mag_2.JK_FF_mag_1.K.n0 CLK_div_3_mag_2.JK_FF_mag_1.K 2.24173
R14 CLK_div_3_mag_2.JK_FF_mag_1.K.n5 CLK_div_3_mag_2.JK_FF_mag_1.K.n0 1.93723
R15 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_1.K.n2 1.81225
R16 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_1.K.n4 1.43709
R17 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_1.K.n1 0.281955
R18 VSS.n95 VSS.n94 97420.2
R19 VSS.n114 VSS.n113 89849.5
R20 VSS.n134 VSS.n133 43844.2
R21 VSS.n103 VSS.n102 31806.2
R22 VSS.n103 VSS.n97 26438.2
R23 VSS.n205 VSS.t18 24327.3
R24 VSS.n129 VSS.t152 22790.4
R25 VSS.n76 VSS.t154 22790.4
R26 VSS.n112 VSS.n111 20600.7
R27 VSS.n133 VSS.n112 16688.2
R28 VSS.t90 VSS.t224 10317.7
R29 VSS.n204 VSS.t248 7248.49
R30 VSS.t171 VSS.n25 7216.19
R31 VSS.n304 VSS.t266 6442.66
R32 VSS.t103 VSS.n129 6161.91
R33 VSS.t121 VSS.n76 5632.67
R34 VSS.t127 VSS.n34 5216.28
R35 VSS.n205 VSS.n204 4665.29
R36 VSS.t68 VSS.n131 4526.01
R37 VSS.n131 VSS.t232 4340.6
R38 VSS.n132 VSS.t11 4253.36
R39 VSS.t181 VSS.n82 4137.27
R40 VSS.n133 VSS.n97 3907.3
R41 VSS.n60 VSS.n59 3893.61
R42 VSS.n284 VSS.n283 3893.61
R43 VSS.n257 VSS.n256 3730.25
R44 VSS.t176 VSS.t86 3492.02
R45 VSS.t92 VSS.t91 3492.02
R46 VSS.t78 VSS.t79 3492.02
R47 VSS.n133 VSS.t31 3396.94
R48 VSS.n117 VSS.n114 3278.96
R49 VSS.n198 VSS.t58 3278.56
R50 VSS.t5 VSS.t7 2781.65
R51 VSS.n257 VSS.t14 2637.2
R52 VSS.t257 VSS.n257 2624.81
R53 VSS.n204 VSS.t244 2581.72
R54 VSS.t207 VSS.t75 2319.79
R55 VSS.t36 VSS.t21 2319.79
R56 VSS.t28 VSS.t27 2307.56
R57 VSS.t213 VSS.t212 2307.56
R58 VSS.t101 VSS.t227 2307.56
R59 VSS.t148 VSS.t190 2307.56
R60 VSS.t239 VSS.t192 2307.56
R61 VSS.t34 VSS.t238 2307.56
R62 VSS.t200 VSS.t198 2307.56
R63 VSS.t41 VSS.t74 2307.56
R64 VSS.t222 VSS.t247 2307.56
R65 VSS.t55 VSS.t46 2307.56
R66 VSS.t220 VSS.t125 2307.56
R67 VSS.t269 VSS.t100 2307.56
R68 VSS.t70 VSS.t59 2307.56
R69 VSS.t204 VSS.t126 2307.56
R70 VSS.t109 VSS.t140 2307.56
R71 VSS.t105 VSS.t22 2307.56
R72 VSS.t174 VSS.n284 2124.81
R73 VSS.n284 VSS.t234 2119.78
R74 VSS.t264 VSS.n228 2098.85
R75 VSS.n59 VSS.t161 2095.66
R76 VSS.n228 VSS.t53 2093.89
R77 VSS.n59 VSS.t168 2090.7
R78 VSS.t26 VSS.t230 2029.37
R79 VSS.t15 VSS.t9 2029.37
R80 VSS.t191 VSS.t150 2029.37
R81 VSS.t233 VSS.t66 2029.37
R82 VSS.t199 VSS.t277 2004.58
R83 VSS.t252 VSS.t135 2004.58
R84 VSS.t124 VSS.t141 2004.58
R85 VSS.t57 VSS.t179 2004.58
R86 VSS.t82 VSS.t157 2001.52
R87 VSS.t2 VSS.t1 2001.52
R88 VSS.t23 VSS.t62 2001.52
R89 VSS.t279 VSS.t282 2001.52
R90 VSS.t11 VSS.t68 1832.21
R91 VSS.n282 VSS.t237 1713.53
R92 VSS.t196 VSS.n205 1601.22
R93 VSS.n130 VSS.t103 1570.47
R94 VSS.n283 VSS.n282 1565.03
R95 VSS.t85 VSS.t176 1382.98
R96 VSS.t91 VSS.t85 1382.98
R97 VSS.t97 VSS.t92 1382.98
R98 VSS.t31 VSS.t78 1382.98
R99 VSS.t79 VSS.t90 1382.98
R100 VSS.n54 VSS.t76 1347.25
R101 VSS.n304 VSS.t228 1199.47
R102 VSS.t165 VSS.n25 1199.47
R103 VSS.n256 VSS.t226 1153.78
R104 VSS.n83 VSS.t60 976.995
R105 VSS.t158 VSS.n93 957.056
R106 VSS.n136 VSS.n135 944.073
R107 VSS.n135 VSS.n134 936.184
R108 VSS.t75 VSS.t16 918.729
R109 VSS.t129 VSS.t108 918.729
R110 VSS.t227 VSS.t147 913.885
R111 VSS.t238 VSS.t132 913.885
R112 VSS.t247 VSS.t216 913.885
R113 VSS.t59 VSS.t45 913.885
R114 VSS.t126 VSS.t17 913.885
R115 VSS.t18 VSS.n176 858.178
R116 VSS.t130 VSS.t215 803.71
R117 VSS.t195 VSS.t15 803.71
R118 VSS.t128 VSS.t241 803.71
R119 VSS.t89 VSS.t233 803.71
R120 VSS.t219 VSS.t43 793.894
R121 VSS.t44 VSS.t252 793.894
R122 VSS.t217 VSS.t268 793.894
R123 VSS.t52 VSS.t57 793.894
R124 VSS.t157 VSS.t112 792.683
R125 VSS.t131 VSS.t186 792.683
R126 VSS.t62 VSS.t120 792.683
R127 VSS.t218 VSS.t276 792.683
R128 VSS.n208 VSS.t249 776.83
R129 VSS.n305 VSS.t145 741.9
R130 VSS.n83 VSS.t181 697.854
R131 VSS.n93 VSS.t121 638.038
R132 VSS.n254 VSS.t50 625
R133 VSS.n159 VSS.n54 614.241
R134 VSS.t7 VSS.n208 554.879
R135 VSS.t16 VSS.n45 551.237
R136 VSS.n47 VSS.t129 551.237
R137 VSS.t21 VSS.n49 551.237
R138 VSS.t76 VSS.n51 551.237
R139 VSS.t226 VSS.n252 548.331
R140 VSS.t27 VSS.n251 548.331
R141 VSS.t212 VSS.n250 548.331
R142 VSS.t147 VSS.n249 548.331
R143 VSS.t237 VSS.n281 548.331
R144 VSS.t190 VSS.n280 548.331
R145 VSS.t192 VSS.n279 548.331
R146 VSS.t244 VSS.n203 548.331
R147 VSS.t198 VSS.n202 548.331
R148 VSS.t74 VSS.n201 548.331
R149 VSS.t216 VSS.n200 548.331
R150 VSS.t58 VSS.n197 548.331
R151 VSS.t125 VSS.n196 548.331
R152 VSS.t100 VSS.n195 548.331
R153 VSS.t45 VSS.n194 548.331
R154 VSS.t17 VSS.n28 548.331
R155 VSS.t140 VSS.n30 548.331
R156 VSS.t22 VSS.n32 548.331
R157 VSS.n35 VSS.t127 548.331
R158 VSS.n212 VSS.t54 546.41
R159 VSS.n265 VSS.t14 482.226
R160 VSS.n266 VSS.t26 482.226
R161 VSS.n270 VSS.t130 482.226
R162 VSS.n285 VSS.t195 482.226
R163 VSS.n291 VSS.t234 482.226
R164 VSS.n292 VSS.t191 482.226
R165 VSS.n296 VSS.t128 482.226
R166 VSS.n297 VSS.t89 482.226
R167 VSS.n222 VSS.t248 476.337
R168 VSS.n223 VSS.t199 476.337
R169 VSS.n227 VSS.t219 476.337
R170 VSS.n229 VSS.t44 476.337
R171 VSS.n235 VSS.t53 476.337
R172 VSS.n236 VSS.t124 476.337
R173 VSS.n240 VSS.t217 476.337
R174 VSS.n258 VSS.t52 476.337
R175 VSS.t112 VSS.n2 475.611
R176 VSS.n4 VSS.t131 475.611
R177 VSS.t1 VSS.n6 475.611
R178 VSS.t161 VSS.n8 475.611
R179 VSS.t120 VSS.n11 475.611
R180 VSS.n13 VSS.t218 475.611
R181 VSS.t282 VSS.n15 475.611
R182 VSS.n17 VSS.t63 475.611
R183 VSS.n45 VSS.t171 367.491
R184 VSS.n47 VSS.t207 367.491
R185 VSS.n49 VSS.t137 367.491
R186 VSS.n51 VSS.t36 367.491
R187 VSS.n252 VSS.t28 365.555
R188 VSS.n251 VSS.t213 365.555
R189 VSS.n250 VSS.t101 365.555
R190 VSS.n249 VSS.t235 365.555
R191 VSS.n281 VSS.t148 365.555
R192 VSS.n280 VSS.t239 365.555
R193 VSS.n279 VSS.t34 365.555
R194 VSS.t228 VSS.n303 365.555
R195 VSS.n203 VSS.t200 365.555
R196 VSS.n202 VSS.t41 365.555
R197 VSS.n201 VSS.t222 365.555
R198 VSS.n200 VSS.t55 365.555
R199 VSS.n197 VSS.t220 365.555
R200 VSS.n196 VSS.t269 365.555
R201 VSS.n195 VSS.t70 365.555
R202 VSS.n194 VSS.t245 365.555
R203 VSS.n28 VSS.t165 365.555
R204 VSS.n30 VSS.t204 365.555
R205 VSS.n32 VSS.t109 365.555
R206 VSS.n35 VSS.t105 365.555
R207 VSS.n212 VSS.t48 364.274
R208 VSS.t230 VSS.n265 321.485
R209 VSS.n266 VSS.t210 321.485
R210 VSS.t9 VSS.n270 321.485
R211 VSS.n285 VSS.t174 321.485
R212 VSS.t150 VSS.n291 321.485
R213 VSS.n292 VSS.t193 321.485
R214 VSS.t66 VSS.n296 321.485
R215 VSS.n297 VSS.t266 321.485
R216 VSS.t277 VSS.n222 317.558
R217 VSS.n223 VSS.t72 317.558
R218 VSS.t135 VSS.n227 317.558
R219 VSS.n229 VSS.t264 317.558
R220 VSS.t141 VSS.n235 317.558
R221 VSS.n236 VSS.t98 317.558
R222 VSS.t179 VSS.n240 317.558
R223 VSS.n258 VSS.t257 317.558
R224 VSS.n2 VSS.t261 317.074
R225 VSS.n4 VSS.t82 317.074
R226 VSS.n6 VSS.t187 317.074
R227 VSS.n8 VSS.t2 317.074
R228 VSS.t168 VSS.n11 317.074
R229 VSS.n13 VSS.t23 317.074
R230 VSS.n15 VSS.t271 317.074
R231 VSS.n17 VSS.t279 317.074
R232 VSS.t232 VSS.n130 174.498
R233 VSS.n156 VSS.t114 132.601
R234 VSS.n283 VSS.n272 119.948
R235 VSS.n199 VSS.n198 119.948
R236 VSS.n130 VSS.n128 116.072
R237 VSS.n94 VSS.t158 109.663
R238 VSS.n159 VSS.n158 98.3817
R239 VSS.n133 VSS.t97 95.0803
R240 VSS.n158 VSS.n157 84.6938
R241 VSS.n157 VSS.n73 79.2822
R242 VSS.t224 VSS.n132 65.4367
R243 VSS.n85 VSS.t162 59.8164
R244 VSS.n73 VSS.n60 58.3607
R245 VSS.t0 VSS.t117 53.9561
R246 VSS.t86 VSS.n117 51.8622
R247 VSS.t117 VSS.n95 49.5516
R248 VSS.n206 VSS.t196 47.5615
R249 VSS.t114 VSS.n136 47.0524
R250 VSS.n272 VSS.t133 34.2711
R251 VSS.t46 VSS.n199 34.2711
R252 VSS.n209 VSS.t5 34.1511
R253 VSS.n256 VSS.n255 32.2586
R254 VSS.n305 VSS.n304 23.9328
R255 VSS.n176 VSS.n25 22.147
R256 VSS.n157 VSS.n96 21.4726
R257 VSS.n255 VSS.n254 20.1618
R258 VSS.n96 VSS.t113 19.2704
R259 VSS.t30 VSS.t77 18.8212
R260 VSS.t113 VSS.t0 12.113
R261 VSS.t77 VSS.n156 11.1218
R262 VSS.n271 VSS.t134 9.3736
R263 VSS.n185 VSS.t47 9.3736
R264 VSS.n253 VSS.t51 9.3736
R265 VSS.n75 VSS.n74 9.37275
R266 VSS.n116 VSS.n115 9.37275
R267 VSS.n175 VSS.n26 9.37275
R268 VSS.n155 VSS.n137 9.37275
R269 VSS.n126 VSS.t153 9.36521
R270 VSS.n211 VSS.t6 9.36521
R271 VSS.n217 VSS.n207 9.3221
R272 VSS.n215 VSS.t8 9.3221
R273 VSS.n122 VSS.n120 9.3221
R274 VSS.n124 VSS.t69 9.3221
R275 VSS.n79 VSS.n78 9.30652
R276 VSS.n307 VSS.t146 9.30652
R277 VSS.n218 VSS.t197 9.30652
R278 VSS.n121 VSS.t225 9.30652
R279 VSS.n87 VSS.n84 9.29578
R280 VSS.n88 VSS.t61 9.29271
R281 VSS.n90 VSS.n80 9.29271
R282 VSS VSS.t104 7.30633
R283 VSS VSS.t49 7.30633
R284 VSS VSS.n77 7.23092
R285 VSS.n143 VSS.n141 7.19156
R286 VSS.n145 VSS.n140 7.19156
R287 VSS.n147 VSS.n139 7.19156
R288 VSS.n71 VSS.n70 7.19156
R289 VSS.n68 VSS.n67 7.19156
R290 VSS.n65 VSS.n64 7.19156
R291 VSS.n37 VSS.n33 7.19156
R292 VSS.n39 VSS.n31 7.19156
R293 VSS.n41 VSS.n29 7.19156
R294 VSS.n151 VSS.n150 7.19156
R295 VSS.n56 VSS.n55 7.19156
R296 VSS.n110 VSS.n109 7.19156
R297 VSS.n107 VSS.n98 7.19156
R298 VSS.n105 VSS.n99 7.19156
R299 VSS.n242 VSS.t29 7.19156
R300 VSS.n244 VSS.t214 7.19156
R301 VSS.n246 VSS.t102 7.19156
R302 VSS.n274 VSS.t149 7.19156
R303 VSS.n276 VSS.t240 7.19156
R304 VSS.n277 VSS.t35 7.19156
R305 VSS.n178 VSS.t201 7.19156
R306 VSS.n180 VSS.t42 7.19156
R307 VSS.n182 VSS.t223 7.19156
R308 VSS.n187 VSS.t221 7.19156
R309 VSS.n189 VSS.t270 7.19156
R310 VSS.n191 VSS.t71 7.19156
R311 VSS.n263 VSS.t231 7.18656
R312 VSS.n268 VSS.t211 7.18656
R313 VSS.n289 VSS.t151 7.18656
R314 VSS.n294 VSS.t194 7.18656
R315 VSS.n220 VSS.t278 7.17656
R316 VSS.n225 VSS.t73 7.17656
R317 VSS.n233 VSS.t142 7.17656
R318 VSS.n238 VSS.t99 7.17656
R319 VSS.n310 VSS.n16 7.16323
R320 VSS.n312 VSS.n14 7.16323
R321 VSS.n319 VSS.n7 7.16323
R322 VSS.n321 VSS.n5 7.16323
R323 VSS.n167 VSS.n50 7.14656
R324 VSS.n169 VSS.n48 7.14656
R325 VSS.n308 VSS.n307 6.33607
R326 VSS.n149 VSS.n138 5.91399
R327 VSS.n62 VSS.n61 5.91399
R328 VSS.n43 VSS.n27 5.91399
R329 VSS.n162 VSS.n160 5.91399
R330 VSS.n164 VSS.n53 5.91399
R331 VSS.n101 VSS.n100 5.91399
R332 VSS.n247 VSS.t236 5.91399
R333 VSS.n301 VSS.t229 5.91399
R334 VSS.n183 VSS.t56 5.91399
R335 VSS.n192 VSS.t246 5.91399
R336 VSS.n20 VSS.t10 5.90898
R337 VSS.n287 VSS.t175 5.90898
R338 VSS.n18 VSS.t67 5.90898
R339 VSS.n299 VSS.t267 5.90898
R340 VSS.n24 VSS.t136 5.89898
R341 VSS.n231 VSS.t265 5.89898
R342 VSS.n22 VSS.t180 5.89898
R343 VSS.n260 VSS.t258 5.89898
R344 VSS.n314 VSS.n12 5.88565
R345 VSS.n316 VSS.n10 5.88565
R346 VSS.n323 VSS.n3 5.88565
R347 VSS.n1 VSS.n0 5.88565
R348 VSS.n171 VSS.n46 5.86898
R349 VSS.n173 VSS.n44 5.86898
R350 VSS.n73 VSS.n72 5.2005
R351 VSS.n73 VSS.n69 5.2005
R352 VSS.n73 VSS.n66 5.2005
R353 VSS.n73 VSS.n63 5.2005
R354 VSS.n96 VSS.n75 5.2005
R355 VSS.n142 VSS.n73 5.2005
R356 VSS.n144 VSS.n73 5.2005
R357 VSS.n146 VSS.n73 5.2005
R358 VSS.n148 VSS.n73 5.2005
R359 VSS.n172 VSS.n45 5.2005
R360 VSS.n170 VSS.n47 5.2005
R361 VSS.n168 VSS.n49 5.2005
R362 VSS.n166 VSS.n51 5.2005
R363 VSS.n112 VSS.n108 5.2005
R364 VSS.n106 VSS.n97 5.2005
R365 VSS.n104 VSS.n103 5.2005
R366 VSS.n117 VSS.n116 5.2005
R367 VSS.n213 VSS.n212 5.2005
R368 VSS.n210 VSS.n209 5.2005
R369 VSS.n216 VSS.n208 5.2005
R370 VSS.n219 VSS.n206 5.2005
R371 VSS.n131 VSS.n127 5.2005
R372 VSS.n132 VSS.n118 5.2005
R373 VSS.n89 VSS.n83 5.2005
R374 VSS.n93 VSS.n92 5.2005
R375 VSS.n86 VSS.n85 5.2005
R376 VSS.n82 VSS.n81 5.2005
R377 VSS.n306 VSS.n305 5.2005
R378 VSS.n265 VSS.n264 5.2005
R379 VSS.n267 VSS.n266 5.2005
R380 VSS.n270 VSS.n269 5.2005
R381 VSS.n286 VSS.n285 5.2005
R382 VSS.n291 VSS.n290 5.2005
R383 VSS.n293 VSS.n292 5.2005
R384 VSS.n296 VSS.n295 5.2005
R385 VSS.n298 VSS.n297 5.2005
R386 VSS.n303 VSS.n302 5.2005
R387 VSS.n279 VSS.n278 5.2005
R388 VSS.n280 VSS.n275 5.2005
R389 VSS.n281 VSS.n273 5.2005
R390 VSS.n252 VSS.n241 5.2005
R391 VSS.n251 VSS.n243 5.2005
R392 VSS.n250 VSS.n245 5.2005
R393 VSS.n249 VSS.n248 5.2005
R394 VSS.n272 VSS.n271 5.2005
R395 VSS.n254 VSS.n253 5.2005
R396 VSS.n259 VSS.n258 5.2005
R397 VSS.n240 VSS.n239 5.2005
R398 VSS.n237 VSS.n236 5.2005
R399 VSS.n235 VSS.n234 5.2005
R400 VSS.n230 VSS.n229 5.2005
R401 VSS.n227 VSS.n226 5.2005
R402 VSS.n224 VSS.n223 5.2005
R403 VSS.n222 VSS.n221 5.2005
R404 VSS.n203 VSS.n177 5.2005
R405 VSS.n202 VSS.n179 5.2005
R406 VSS.n201 VSS.n181 5.2005
R407 VSS.n200 VSS.n184 5.2005
R408 VSS.n199 VSS.n185 5.2005
R409 VSS.n197 VSS.n186 5.2005
R410 VSS.n196 VSS.n188 5.2005
R411 VSS.n195 VSS.n190 5.2005
R412 VSS.n194 VSS.n193 5.2005
R413 VSS.n176 VSS.n175 5.2005
R414 VSS.n36 VSS.n35 5.2005
R415 VSS.n38 VSS.n32 5.2005
R416 VSS.n40 VSS.n30 5.2005
R417 VSS.n42 VSS.n28 5.2005
R418 VSS.n159 VSS.n58 5.2005
R419 VSS.n159 VSS.n57 5.2005
R420 VSS.n161 VSS.n159 5.2005
R421 VSS.n163 VSS.n159 5.2005
R422 VSS.n156 VSS.n155 5.2005
R423 VSS.n324 VSS.n2 5.2005
R424 VSS.n322 VSS.n4 5.2005
R425 VSS.n320 VSS.n6 5.2005
R426 VSS.n318 VSS.n8 5.2005
R427 VSS.n315 VSS.n11 5.2005
R428 VSS.n313 VSS.n13 5.2005
R429 VSS.n311 VSS.n15 5.2005
R430 VSS.n309 VSS.n17 5.2005
R431 VSS.n157 VSS.t30 3.42245
R432 VSS.n262 VSS 2.278
R433 VSS VSS.n308 1.06574
R434 VSS.n165 VSS.n52 0.93911
R435 VSS.n174 VSS.n173 0.937801
R436 VSS.n300 VSS.n299 0.930005
R437 VSS.n288 VSS.n19 0.843437
R438 VSS.n232 VSS.n23 0.838483
R439 VSS.n261 VSS.n21 0.838483
R440 VSS.n317 VSS.n9 0.832426
R441 VSS.n154 VSS.n153 0.832426
R442 VSS VSS.n165 0.677636
R443 VSS VSS.n152 0.376792
R444 VSS VSS.n145 0.343161
R445 VSS VSS.n143 0.343161
R446 VSS.n68 VSS 0.343161
R447 VSS.n71 VSS 0.343161
R448 VSS VSS.n39 0.343161
R449 VSS VSS.n37 0.343161
R450 VSS.n107 VSS 0.343161
R451 VSS.n110 VSS 0.343161
R452 VSS VSS.n242 0.343161
R453 VSS VSS.n244 0.343161
R454 VSS VSS.n274 0.343161
R455 VSS VSS.n276 0.343161
R456 VSS VSS.n178 0.343161
R457 VSS VSS.n180 0.343161
R458 VSS VSS.n187 0.343161
R459 VSS VSS.n189 0.343161
R460 VSS.n125 VSS.n124 0.309418
R461 VSS.n215 VSS.n214 0.309418
R462 VSS.n91 VSS.n90 0.300071
R463 VSS.n172 VSS.n171 0.292623
R464 VSS.n170 VSS.n169 0.292623
R465 VSS.n148 VSS 0.289491
R466 VSS VSS.n63 0.289491
R467 VSS.n42 VSS 0.289491
R468 VSS VSS.n104 0.289491
R469 VSS.n248 VSS 0.289491
R470 VSS.n302 VSS 0.289491
R471 VSS.n184 VSS 0.289491
R472 VSS.n193 VSS 0.289491
R473 VSS.n308 VSS 0.267286
R474 VSS.n125 VSS.n119 0.255008
R475 VSS.n214 VSS.n213 0.255008
R476 VSS.n92 VSS.n91 0.230643
R477 VSS.n269 VSS.n268 0.222068
R478 VSS.n286 VSS.n20 0.222068
R479 VSS.n295 VSS.n294 0.222068
R480 VSS.n298 VSS.n18 0.222068
R481 VSS.n226 VSS.n225 0.222068
R482 VSS.n230 VSS.n24 0.222068
R483 VSS.n239 VSS.n238 0.222068
R484 VSS.n259 VSS.n22 0.222068
R485 VSS.n324 VSS.n323 0.222068
R486 VSS.n322 VSS.n321 0.222068
R487 VSS.n315 VSS.n314 0.222068
R488 VSS.n313 VSS.n312 0.222068
R489 VSS VSS.n167 0.209159
R490 VSS VSS.n147 0.191234
R491 VSS.n65 VSS 0.191234
R492 VSS VSS.n41 0.191234
R493 VSS.n105 VSS 0.191234
R494 VSS VSS.n246 0.191234
R495 VSS.n277 VSS 0.191234
R496 VSS VSS.n182 0.191234
R497 VSS VSS.n191 0.191234
R498 VSS.n218 VSS.n217 0.168119
R499 VSS.n122 VSS.n121 0.168119
R500 VSS.n263 VSS 0.158763
R501 VSS.n289 VSS 0.158763
R502 VSS.n220 VSS 0.158763
R503 VSS.n233 VSS 0.158763
R504 VSS VSS.n319 0.158763
R505 VSS VSS.n310 0.158763
R506 VSS.n262 VSS.n261 0.150892
R507 VSS.n88 VSS.n87 0.147714
R508 VSS.n153 VSS 0.142364
R509 VSS.n126 VSS.n125 0.141461
R510 VSS.n214 VSS.n211 0.141461
R511 VSS VSS.n19 0.137685
R512 VSS.n300 VSS 0.137685
R513 VSS VSS.n23 0.137685
R514 VSS VSS.n21 0.137685
R515 VSS VSS.n9 0.137136
R516 VSS VSS.n52 0.137136
R517 VSS VSS.n174 0.137136
R518 VSS VSS.n154 0.137136
R519 VSS.n217 VSS.n216 0.136634
R520 VSS.n123 VSS.n122 0.136634
R521 VSS VSS.n262 0.135131
R522 VSS.n163 VSS.n162 0.123535
R523 VSS.n147 VSS.n146 0.118573
R524 VSS.n145 VSS.n144 0.118573
R525 VSS.n143 VSS.n142 0.118573
R526 VSS.n66 VSS.n65 0.118573
R527 VSS.n69 VSS.n68 0.118573
R528 VSS.n72 VSS.n71 0.118573
R529 VSS.n41 VSS.n40 0.118573
R530 VSS.n39 VSS.n38 0.118573
R531 VSS.n37 VSS.n36 0.118573
R532 VSS.n106 VSS.n105 0.118573
R533 VSS.n108 VSS.n107 0.118573
R534 VSS.n111 VSS.n110 0.118573
R535 VSS.n242 VSS.n241 0.118573
R536 VSS.n244 VSS.n243 0.118573
R537 VSS.n246 VSS.n245 0.118573
R538 VSS.n274 VSS.n273 0.118573
R539 VSS.n276 VSS.n275 0.118573
R540 VSS.n278 VSS.n277 0.118573
R541 VSS.n178 VSS.n177 0.118573
R542 VSS.n180 VSS.n179 0.118573
R543 VSS.n182 VSS.n181 0.118573
R544 VSS.n187 VSS.n186 0.118573
R545 VSS.n189 VSS.n188 0.118573
R546 VSS.n191 VSS.n190 0.118573
R547 VSS.n89 VSS.n88 0.116857
R548 VSS VSS.n215 0.115458
R549 VSS.n124 VSS 0.115458
R550 VSS.n149 VSS 0.115271
R551 VSS VSS.n62 0.115271
R552 VSS.n43 VSS 0.115271
R553 VSS VSS.n101 0.115271
R554 VSS VSS.n247 0.115271
R555 VSS VSS.n301 0.115271
R556 VSS VSS.n183 0.115271
R557 VSS VSS.n192 0.115271
R558 VSS.n154 VSS.n149 0.10206
R559 VSS.n62 VSS.n9 0.10206
R560 VSS.n174 VSS.n43 0.10206
R561 VSS.n101 VSS.n52 0.10206
R562 VSS.n247 VSS.n19 0.10206
R563 VSS.n301 VSS.n300 0.10206
R564 VSS.n183 VSS.n23 0.10206
R565 VSS.n192 VSS.n21 0.10206
R566 VSS.n90 VSS 0.0975714
R567 VSS.n151 VSS 0.0883824
R568 VSS.n288 VSS.n287 0.0870678
R569 VSS.n232 VSS.n231 0.0870678
R570 VSS.n153 VSS.n1 0.0866864
R571 VSS.n317 VSS.n316 0.0866864
R572 VSS.n91 VSS.n79 0.0855927
R573 VSS VSS.n317 0.0855424
R574 VSS.n261 VSS.n260 0.0853298
R575 VSS VSS.n288 0.085161
R576 VSS VSS.n232 0.085161
R577 VSS.n169 VSS.n168 0.0723994
R578 VSS.n167 VSS.n166 0.0723994
R579 VSS.n173 VSS 0.0703883
R580 VSS.n171 VSS 0.0703883
R581 VSS.n307 VSS.n306 0.0675755
R582 VSS.n81 VSS.n79 0.0667264
R583 VSS.n127 VSS.n126 0.0589274
R584 VSS.n211 VSS.n210 0.0589274
R585 VSS.n219 VSS.n218 0.0564843
R586 VSS.n121 VSS.n118 0.0564843
R587 VSS.n264 VSS.n263 0.0550339
R588 VSS.n268 VSS.n267 0.0550339
R589 VSS.n290 VSS.n289 0.0550339
R590 VSS.n294 VSS.n293 0.0550339
R591 VSS.n221 VSS.n220 0.0550339
R592 VSS.n225 VSS.n224 0.0550339
R593 VSS.n234 VSS.n233 0.0550339
R594 VSS.n238 VSS.n237 0.0550339
R595 VSS.n321 VSS.n320 0.0550339
R596 VSS.n319 VSS.n318 0.0550339
R597 VSS.n312 VSS.n311 0.0550339
R598 VSS.n310 VSS.n309 0.0550339
R599 VSS VSS.n20 0.0535085
R600 VSS.n287 VSS 0.0535085
R601 VSS VSS.n18 0.0535085
R602 VSS.n299 VSS 0.0535085
R603 VSS VSS.n24 0.0535085
R604 VSS.n231 VSS 0.0535085
R605 VSS VSS.n22 0.0535085
R606 VSS.n260 VSS 0.0535085
R607 VSS VSS.n1 0.0535085
R608 VSS.n323 VSS 0.0535085
R609 VSS.n316 VSS 0.0535085
R610 VSS.n314 VSS 0.0535085
R611 VSS.n87 VSS.n86 0.0506429
R612 VSS.n57 VSS.n56 0.0307824
R613 VSS.n164 VSS 0.0299353
R614 VSS.n162 VSS 0.0299353
R615 VSS.n152 VSS.n151 0.0168059
R616 VSS.n152 VSS.n58 0.0144765
R617 VSS.n146 VSS 0.00545413
R618 VSS.n144 VSS 0.00545413
R619 VSS.n142 VSS 0.00545413
R620 VSS VSS.n66 0.00545413
R621 VSS VSS.n69 0.00545413
R622 VSS.n72 VSS 0.00545413
R623 VSS.n40 VSS 0.00545413
R624 VSS.n38 VSS 0.00545413
R625 VSS.n36 VSS 0.00545413
R626 VSS VSS.n106 0.00545413
R627 VSS VSS.n108 0.00545413
R628 VSS.n111 VSS 0.00545413
R629 VSS.n241 VSS 0.00545413
R630 VSS.n243 VSS 0.00545413
R631 VSS.n245 VSS 0.00545413
R632 VSS.n273 VSS 0.00545413
R633 VSS.n275 VSS 0.00545413
R634 VSS.n278 VSS 0.00545413
R635 VSS.n177 VSS 0.00545413
R636 VSS.n179 VSS 0.00545413
R637 VSS.n181 VSS 0.00545413
R638 VSS.n186 VSS 0.00545413
R639 VSS.n188 VSS 0.00545413
R640 VSS.n190 VSS 0.00545413
R641 VSS VSS.n148 0.00380275
R642 VSS.n63 VSS 0.00380275
R643 VSS VSS.n42 0.00380275
R644 VSS.n104 VSS 0.00380275
R645 VSS.n119 VSS 0.00380275
R646 VSS.n248 VSS 0.00380275
R647 VSS.n302 VSS 0.00380275
R648 VSS.n213 VSS 0.00380275
R649 VSS.n184 VSS 0.00380275
R650 VSS.n193 VSS 0.00380275
R651 VSS.n216 VSS 0.00352521
R652 VSS VSS.n123 0.00352521
R653 VSS.n168 VSS 0.00351676
R654 VSS.n166 VSS 0.00351676
R655 VSS.n92 VSS 0.00307143
R656 VSS VSS.n89 0.00307143
R657 VSS.n165 VSS.n164 0.00282941
R658 VSS.n264 VSS 0.00278814
R659 VSS.n267 VSS 0.00278814
R660 VSS.n290 VSS 0.00278814
R661 VSS.n293 VSS 0.00278814
R662 VSS.n221 VSS 0.00278814
R663 VSS.n224 VSS 0.00278814
R664 VSS.n234 VSS 0.00278814
R665 VSS.n237 VSS 0.00278814
R666 VSS.n320 VSS 0.00278814
R667 VSS.n318 VSS 0.00278814
R668 VSS.n311 VSS 0.00278814
R669 VSS.n309 VSS 0.00278814
R670 VSS VSS.n172 0.00251117
R671 VSS VSS.n170 0.00251117
R672 VSS.n75 VSS 0.00219811
R673 VSS.n116 VSS 0.00219811
R674 VSS.n175 VSS 0.00219811
R675 VSS.n127 VSS 0.00219811
R676 VSS.n271 VSS 0.00219811
R677 VSS.n81 VSS 0.00219811
R678 VSS.n306 VSS 0.00219811
R679 VSS.n210 VSS 0.00219811
R680 VSS.n185 VSS 0.00219811
R681 VSS.n253 VSS 0.00219811
R682 VSS.n155 VSS 0.00219811
R683 VSS.n269 VSS 0.00202542
R684 VSS VSS.n286 0.00202542
R685 VSS.n295 VSS 0.00202542
R686 VSS VSS.n298 0.00202542
R687 VSS.n226 VSS 0.00202542
R688 VSS VSS.n230 0.00202542
R689 VSS.n239 VSS 0.00202542
R690 VSS VSS.n259 0.00202542
R691 VSS VSS.n324 0.00202542
R692 VSS VSS.n322 0.00202542
R693 VSS VSS.n315 0.00202542
R694 VSS VSS.n313 0.00202542
R695 VSS VSS.n219 0.00191732
R696 VSS.n118 VSS 0.00191732
R697 VSS.n86 VSS 0.00178571
R698 VSS VSS.n57 0.00177059
R699 VSS.n58 VSS 0.00177059
R700 VSS VSS.n163 0.00134706
R701 VSS VSS.n161 0.00134706
R702 RST.n9 RST.t3 37.2596
R703 RST.n38 RST.t4 37.1991
R704 RST.n25 RST.t13 37.1991
R705 RST.n61 RST.t7 36.935
R706 RST.n0 RST.t11 36.935
R707 RST.n47 RST.t0 36.935
R708 RST.n30 RST.t8 36.935
R709 RST.n16 RST.t14 36.935
R710 RST.n61 RST.t6 18.1962
R711 RST.n0 RST.t9 18.1962
R712 RST.n47 RST.t15 18.1962
R713 RST.n30 RST.t5 18.1962
R714 RST.n16 RST.t12 18.1962
R715 RST.n38 RST.t1 17.66
R716 RST.n25 RST.t10 17.66
R717 RST.n9 RST.t2 17.5947
R718 RST.n29 RST.n28 9.41979
R719 RST.n42 RST.n41 9.37665
R720 RST.n20 RST.n19 4.81648
R721 RST.n54 RST.n53 4.51217
R722 RST.n19 RST.n18 4.5005
R723 RST.n55 RST.n54 4.5005
R724 RST.n57 RST.n56 4.5005
R725 RST.n20 RST.n13 4.44014
R726 RST.n35 RST.n34 3.74791
R727 RST.n34 RST.n20 3.63633
R728 RST.n70 RST.n69 2.25327
R729 RST.n33 RST.n32 2.25296
R730 RST.n50 RST.n49 2.2505
R731 RST.n17 RST.n15 2.25022
R732 RST.n32 RST.n29 2.25014
R733 RST.n63 RST.n62 2.24906
R734 RST.n13 RST.n12 2.24196
R735 RST.n41 RST.n40 2.24157
R736 RST.n28 RST.n27 2.24157
R737 RST.n62 RST.n61 2.12658
R738 RST.n17 RST.n16 2.12393
R739 RST.n1 RST.n0 2.12207
R740 RST.n48 RST.n47 2.12175
R741 RST.n31 RST.n30 2.12075
R742 RST.n67 RST.n57 2.06412
R743 RST.n34 RST.n33 1.93664
R744 RST.n68 RST.n7 1.73035
R745 RST.n65 RST.n64 1.60789
R746 RST.n5 RST.n3 1.5005
R747 RST.n10 RST.n9 1.42168
R748 RST.n39 RST.n38 1.41552
R749 RST.n26 RST.n25 1.41552
R750 RST.n7 RST.n6 1.13388
R751 RST.n68 RST.n67 0.659395
R752 RST.n70 RST.n68 0.610028
R753 RST.n14 RST 0.0584663
R754 RST RST.n55 0.0455
R755 RST.n46 RST 0.0410354
R756 RST.n37 RST 0.0410354
R757 RST.n22 RST 0.0410354
R758 RST.n24 RST 0.0410354
R759 RST.n11 RST 0.0394837
R760 RST.n12 RST.n11 0.0377414
R761 RST.n59 RST 0.0363802
R762 RST.n3 RST.n2 0.0361897
R763 RST.n49 RST.n46 0.0361897
R764 RST.n40 RST.n37 0.0361897
R765 RST.n32 RST.n22 0.0361897
R766 RST.n27 RST.n24 0.0361897
R767 RST.n2 RST 0.0348285
R768 RST.n60 RST.n59 0.0346379
R769 RST.n19 RST 0.0293
R770 RST.n45 RST.n44 0.0257439
R771 RST.n29 RST 0.0244407
R772 RST.n13 RST.n8 0.0238218
R773 RST.n41 RST.n36 0.0230258
R774 RST.n28 RST.n23 0.0230258
R775 RST.n18 RST.n14 0.0196058
R776 RST.n43 RST.n42 0.0191585
R777 RST.n63 RST.n58 0.016866
R778 RST.n66 RST.n65 0.0147105
R779 RST.n52 RST.n35 0.0132559
R780 RST.n5 RST.n4 0.0131308
R781 RST.n3 RST.n1 0.00981034
R782 RST.n33 RST.n21 0.00906463
R783 RST.n64 RST.n63 0.00887538
R784 RST.n67 RST.n66 0.00713158
R785 RST.n57 RST.n35 0.00687795
R786 RST.n54 RST.n52 0.00687795
R787 RST.n6 RST.n5 0.00685294
R788 RST.n51 RST.n50 0.0055
R789 RST.n56 RST 0.0055
R790 RST.n49 RST.n48 0.00515517
R791 RST.n40 RST.n39 0.00515517
R792 RST.n32 RST.n31 0.00515517
R793 RST.n27 RST.n26 0.00515517
R794 RST.n62 RST.n60 0.00487597
R795 RST.n50 RST.n45 0.00383333
R796 RST.n12 RST.n10 0.00360345
R797 RST.n44 RST.n43 0.00269512
R798 RST.n18 RST.n17 0.00255119
R799 RST.n56 RST.n51 0.00216667
R800 RST.n15 RST 0.0017
R801 RST RST.n21 0.00153448
R802 RST RST.n70 0.000978723
R803 CLK_div_3_mag_0.CLK.n9 CLK_div_3_mag_0.CLK.t11 36.935
R804 CLK_div_3_mag_0.CLK.n8 CLK_div_3_mag_0.CLK.t8 36.935
R805 CLK_div_3_mag_0.CLK.n13 CLK_div_3_mag_0.CLK.t5 36.935
R806 CLK_div_3_mag_0.CLK.n12 CLK_div_3_mag_0.CLK.t2 36.935
R807 CLK_div_3_mag_0.CLK.n10 CLK_div_3_mag_0.CLK.t10 30.6315
R808 CLK_div_3_mag_0.CLK.n14 CLK_div_3_mag_0.CLK.t7 25.5364
R809 CLK_div_3_mag_0.CLK.n17 CLK_div_3_mag_0.CLK.t13 25.536
R810 CLK_div_3_mag_0.CLK.n10 CLK_div_3_mag_0.CLK.t14 21.7275
R811 CLK_div_3_mag_0.CLK.n9 CLK_div_3_mag_0.CLK.t9 18.1962
R812 CLK_div_3_mag_0.CLK.n8 CLK_div_3_mag_0.CLK.t6 18.1962
R813 CLK_div_3_mag_0.CLK.n13 CLK_div_3_mag_0.CLK.t3 18.1962
R814 CLK_div_3_mag_0.CLK.n12 CLK_div_3_mag_0.CLK.t15 18.1962
R815 CLK_div_3_mag_0.CLK.n14 CLK_div_3_mag_0.CLK.t12 14.0749
R816 CLK_div_3_mag_0.CLK.n17 CLK_div_3_mag_0.CLK.t4 14.0734
R817 CLK_div_3_mag_0.CLK.n7 CLK_div_3_mag_0.CLK.t1 9.29842
R818 CLK_div_3_mag_0.CLK.n0 CLK_div_3_mag_0.CLK.n11 7.41537
R819 CLK_div_3_mag_0.CLK.n16 CLK_div_3_mag_0.CLK.n15 5.37352
R820 CLK_div_3_mag_0.CLK.n7 CLK_div_3_mag_0.CLK.t0 5.05693
R821 CLK_div_3_mag_0.CLK.n4 CLK_div_3_mag_0.CLK.n8 2.13042
R822 CLK_div_3_mag_0.CLK.n2 CLK_div_3_mag_0.CLK.n1 1.11863
R823 CLK_div_3_mag_0.CLK.n5 CLK_div_3_mag_0.CLK.n12 2.13042
R824 CLK_div_3_mag_0.CLK CLK_div_3_mag_0.CLK.n3 0.0786548
R825 CLK_div_3_mag_0.CLK.n13 CLK_div_3_mag_0.CLK.n3 2.13151
R826 CLK_div_3_mag_0.CLK.n14 CLK_div_3_mag_0.CLK 1.4356
R827 CLK_div_3_mag_0.CLK.n6 CLK_div_3_mag_0.CLK.n17 1.43283
R828 CLK_div_3_mag_0.CLK.n0 CLK_div_3_mag_0.CLK.n3 1.11863
R829 CLK_div_3_mag_0.CLK.n2 CLK_div_3_mag_0.CLK.n9 2.13151
R830 CLK_div_3_mag_0.CLK.n11 CLK_div_3_mag_0.CLK.n10 1.80477
R831 CLK_div_3_mag_0.CLK.n1 CLK_div_3_mag_0.CLK.n4 2.63808
R832 CLK_div_3_mag_0.CLK.n0 CLK_div_3_mag_0.CLK.n5 2.51975
R833 CLK_div_3_mag_0.CLK.n11 CLK_div_3_mag_0.CLK 0.105737
R834 CLK_div_3_mag_0.CLK CLK_div_3_mag_0.CLK.n7 0.0833947
R835 CLK_div_3_mag_0.CLK.n2 CLK_div_3_mag_0.CLK 0.0786548
R836 CLK_div_3_mag_0.CLK.n4 CLK_div_3_mag_0.CLK 0.0807313
R837 CLK_div_3_mag_0.CLK.n5 CLK_div_3_mag_0.CLK 0.0807313
R838 CLK_div_3_mag_0.CLK CLK_div_3_mag_0.CLK.n6 0.132999
R839 CLK_div_3_mag_0.CLK.n6 CLK_div_3_mag_0.CLK.n16 1.1982
R840 CLK_div_3_mag_0.CLK.n15 CLK_div_3_mag_0.CLK 1.19627
R841 CLK_div_3_mag_0.CLK.n15 CLK_div_3_mag_0.CLK.n0 1.01264
R842 CLK_div_3_mag_0.CLK.n16 CLK_div_3_mag_0.CLK.n1 0.894314
R843 VDD.t187 VDD.n62 15263.4
R844 VDD.t0 VDD.t409 13138
R845 VDD.n167 VDD.t83 2309.15
R846 VDD.t216 VDD.t360 1131.65
R847 VDD.t162 VDD.t412 1131.65
R848 VDD.t119 VDD.t102 1131.65
R849 VDD.t40 VDD.t37 961.905
R850 VDD.t349 VDD.t352 961.905
R851 VDD.t167 VDD.t369 961.905
R852 VDD.t179 VDD.t380 961.905
R853 VDD VDD.n339 899.707
R854 VDD.t331 VDD.t427 765.152
R855 VDD.t76 VDD.t124 765.152
R856 VDD.t407 VDD.t223 765.152
R857 VDD.t213 VDD.t229 765.152
R858 VDD.t414 VDD.t165 765.152
R859 VDD.t100 VDD.t298 765.152
R860 VDD.t143 VDD.t255 765.152
R861 VDD.t306 VDD.t309 765.152
R862 VDD.t4 VDD.t2 765.152
R863 VDD.t258 VDD.t113 765.152
R864 VDD.t419 VDD.t421 765.152
R865 VDD.t432 VDD.t73 765.152
R866 VDD.t29 VDD.t107 765.152
R867 VDD.t424 VDD.t416 765.152
R868 VDD.t429 VDD.t434 765.152
R869 VDD.t317 VDD.t238 765.152
R870 VDD.t390 VDD.t323 765.152
R871 VDD.t378 VDD.t116 765.152
R872 VDD.t34 VDD.t373 765.152
R873 VDD.t354 VDD.t347 765.152
R874 VDD.t17 VDD.t11 765.152
R875 VDD.t339 VDD.t130 765.152
R876 VDD.t42 VDD.t157 765.152
R877 VDD.t231 VDD.t133 765.152
R878 VDD.t334 VDD.t337 765.152
R879 VDD.t78 VDD.t121 765.152
R880 VDD.t399 VDD.t362 765.152
R881 VDD.t344 VDD.t146 765.152
R882 VDD.t190 VDD.t225 765.152
R883 VDD.t50 VDD.t26 765.152
R884 VDD.n358 VDD.t314 675.778
R885 VDD.n490 VDD.n489 634.846
R886 VDD.n61 VDD.t19 468.392
R887 VDD.n109 VDD.n108 450.161
R888 VDD.t360 VDD.t104 448.18
R889 VDD.t412 VDD.t216 448.18
R890 VDD.t102 VDD.t80 448.18
R891 VDD.t80 VDD.t402 448.18
R892 VDD.n475 VDD.t119 434.175
R893 VDD VDD.n405 426.699
R894 VDD.n405 VDD.t245 386.365
R895 VDD.t369 VDD.t184 380.952
R896 VDD VDD.n169 365.748
R897 VDD.t48 VDD.t300 330.365
R898 VDD.t375 VDD.t312 320.125
R899 VDD.t320 VDD.t250 320.125
R900 VDD.t70 VDD.t76 303.031
R901 VDD.t356 VDD.t407 303.031
R902 VDD.t53 VDD.t414 303.031
R903 VDD.t87 VDD.t100 303.031
R904 VDD.t255 VDD.t209 303.031
R905 VDD.t56 VDD.t306 303.031
R906 VDD.t211 VDD.t258 303.031
R907 VDD.t107 VDD.t197 303.031
R908 VDD.t68 VDD.t424 303.031
R909 VDD.t65 VDD.t390 303.031
R910 VDD.t181 VDD.t378 303.031
R911 VDD.t58 VDD.t354 303.031
R912 VDD.t169 VDD.t17 303.031
R913 VDD.t130 VDD.t126 303.031
R914 VDD.t63 VDD.t42 303.031
R915 VDD.t90 VDD.t399 303.031
R916 VDD.t146 VDD.t22 303.031
R917 VDD.t60 VDD.t190 303.031
R918 VDD.n489 VDD.n109 292.675
R919 VDD.n292 VDD.t366 242.857
R920 VDD.n307 VDD.t37 242.857
R921 VDD.n308 VDD.t349 242.857
R922 VDD.n313 VDD.t184 242.857
R923 VDD.n359 VDD.t385 242.857
R924 VDD.n167 VDD.t149 229.731
R925 VDD.n339 VDD.t252 194.631
R926 VDD.n73 VDD.t404 193.183
R927 VDD.n75 VDD.t331 193.183
R928 VDD.n78 VDD.t70 193.183
R929 VDD.n81 VDD.t356 193.183
R930 VDD.n111 VDD.t95 193.183
R931 VDD.n113 VDD.t213 193.183
R932 VDD.n116 VDD.t53 193.183
R933 VDD.n119 VDD.t87 193.183
R934 VDD.n230 VDD.t382 193.183
R935 VDD.n232 VDD.t317 193.183
R936 VDD.n235 VDD.t65 193.183
R937 VDD.n238 VDD.t181 193.183
R938 VDD.n271 VDD.t13 193.183
R939 VDD.n273 VDD.t34 193.183
R940 VDD.n276 VDD.t58 193.183
R941 VDD.n279 VDD.t169 193.183
R942 VDD.n96 VDD.t397 193.183
R943 VDD.n97 VDD.t334 193.183
R944 VDD.n103 VDD.t121 193.183
R945 VDD.n104 VDD.t90 193.183
R946 VDD.t209 VDD.n208 191.288
R947 VDD.n209 VDD.t56 191.288
R948 VDD.t2 VDD.n217 191.288
R949 VDD.n218 VDD.t248 191.288
R950 VDD.n404 VDD.t211 191.288
R951 VDD.n403 VDD.t419 191.288
R952 VDD.n402 VDD.t432 191.288
R953 VDD.n401 VDD.t234 191.288
R954 VDD.t197 VDD.n386 191.288
R955 VDD.n387 VDD.t68 191.288
R956 VDD.t434 VDD.n395 191.288
R957 VDD.n396 VDD.t110 191.288
R958 VDD.t126 VDD.n444 191.288
R959 VDD.n445 VDD.t63 191.288
R960 VDD.t133 VDD.n453 191.288
R961 VDD.n454 VDD.t195 191.288
R962 VDD.t22 VDD.n19 191.288
R963 VDD.n20 VDD.t60 191.288
R964 VDD.t26 VDD.n28 191.288
R965 VDD.n29 VDD.t128 191.288
R966 VDD.n410 VDD.t325 179.715
R967 VDD.n425 VDD.n424 179.567
R968 VDD.n108 VDD.t85 173.633
R969 VDD.n337 VDD.t371 164.286
R970 VDD.n63 VDD.t221 159.306
R971 VDD.n147 VDD.t32 151.653
R972 VDD.n466 VDD.t135 151.653
R973 VDD.t149 VDD.n166 151.653
R974 VDD.t394 VDD.n172 149.114
R975 VDD.n476 VDD.n475 145.647
R976 VDD.n478 VDD.t151 139.641
R977 VDD.n153 VDD.t160 139.641
R978 VDD.n292 VDD.t40 138.095
R979 VDD.t352 VDD.n307 138.095
R980 VDD.n308 VDD.t167 138.095
R981 VDD.t380 VDD.n313 138.095
R982 VDD.n359 VDD.n358 123.486
R983 VDD.n425 VDD.t16 117.647
R984 VDD.n208 VDD.t270 111.743
R985 VDD.n209 VDD.t143 111.743
R986 VDD.n217 VDD.t309 111.743
R987 VDD.n218 VDD.t4 111.743
R988 VDD.t245 VDD.n404 111.743
R989 VDD.t113 VDD.n403 111.743
R990 VDD.t421 VDD.n402 111.743
R991 VDD.t73 VDD.n401 111.743
R992 VDD.n386 VDD.t292 111.743
R993 VDD.n387 VDD.t29 111.743
R994 VDD.n395 VDD.t416 111.743
R995 VDD.n396 VDD.t429 111.743
R996 VDD.n444 VDD.t274 111.743
R997 VDD.n445 VDD.t339 111.743
R998 VDD.n453 VDD.t157 111.743
R999 VDD.n454 VDD.t231 111.743
R1000 VDD.n19 VDD.t288 111.743
R1001 VDD.n20 VDD.t344 111.743
R1002 VDD.n28 VDD.t225 111.743
R1003 VDD.n29 VDD.t50 111.743
R1004 VDD.t427 VDD.n73 109.849
R1005 VDD.t124 VDD.n75 109.849
R1006 VDD.t223 VDD.n78 109.849
R1007 VDD.n81 VDD.t267 109.849
R1008 VDD.t229 VDD.n111 109.849
R1009 VDD.t165 VDD.n113 109.849
R1010 VDD.t298 VDD.n116 109.849
R1011 VDD.n119 VDD.t282 109.849
R1012 VDD.t238 VDD.n230 109.849
R1013 VDD.t323 VDD.n232 109.849
R1014 VDD.t116 VDD.n235 109.849
R1015 VDD.n238 VDD.t264 109.849
R1016 VDD.t373 VDD.n271 109.849
R1017 VDD.t347 VDD.n273 109.849
R1018 VDD.t11 VDD.n276 109.849
R1019 VDD.n279 VDD.t285 109.849
R1020 VDD.t337 VDD.n96 109.849
R1021 VDD.n97 VDD.t78 109.849
R1022 VDD.t362 VDD.n103 109.849
R1023 VDD.n104 VDD.t98 109.849
R1024 VDD.n37 VDD.n33 107.162
R1025 VDD.t409 VDD.n410 104.983
R1026 VDD.t303 VDD.t375 101.147
R1027 VDD.t174 VDD.t0 101.147
R1028 VDD.t314 VDD.t199 101.147
R1029 VDD.t250 VDD.t392 101.147
R1030 VDD.t312 VDD.n187 99.062
R1031 VDD.n349 VDD.t320 99.062
R1032 VDD.n169 VDD.t202 97.8092
R1033 VDD.n61 VDD 95.381
R1034 VDD.n63 VDD.t187 93.0604
R1035 VDD.n173 VDD.n169 92.8798
R1036 VDD.n336 VDD.t176 91.0719
R1037 VDD.n147 VDD.t278 88.5891
R1038 VDD.n476 VDD.t154 88.5891
R1039 VDD.n466 VDD.t45 88.5891
R1040 VDD.n166 VDD.t140 88.5891
R1041 VDD.n40 VDD.n39 82.9474
R1042 VDD.t16 VDD.t364 82.5598
R1043 VDD.n347 VDD.t112 80.3576
R1044 VDD.n423 VDD.n175 75.0412
R1045 VDD.n62 VDD.t24 70.5827
R1046 VDD.n173 VDD.n172 66.048
R1047 VDD.n424 VDD.n172 63.984
R1048 VDD.n405 VDD.t206 62.1896
R1049 VDD.n186 VDD.t394 61.5229
R1050 VDD.n348 VDD.t48 60.4802
R1051 VDD.n411 VDD.n188 56.3092
R1052 VDD.n357 VDD.n320 56.3092
R1053 VDD.t300 VDD.t387 51.7862
R1054 VDD.t176 VDD.t112 51.7862
R1055 VDD.t371 VDD.n336 51.7862
R1056 VDD.t7 VDD.t9 41.7316
R1057 VDD.t9 VDD.t329 39.1388
R1058 VDD.n120 VDD.t266 30.9379
R1059 VDD.n195 VDD.t291 30.9379
R1060 VDD.n241 VDD.t284 30.9379
R1061 VDD.n434 VDD.t273 30.9379
R1062 VDD.n436 VDD.t277 30.9379
R1063 VDD.n10 VDD.t287 30.9379
R1064 VDD.n11 VDD.t295 30.9379
R1065 VDD.n198 VDD.t269 30.2877
R1066 VDD.n125 VDD.t281 30.0062
R1067 VDD.n240 VDD.t263 30.0062
R1068 VDD.n346 VDD.n328 26.7837
R1069 VDD.n120 VDD.t450 24.5101
R1070 VDD.n199 VDD.t449 24.5101
R1071 VDD.n195 VDD.t439 24.5101
R1072 VDD.n241 VDD.t442 24.5101
R1073 VDD.n434 VDD.t447 24.5101
R1074 VDD.n436 VDD.t444 24.5101
R1075 VDD.n10 VDD.t441 24.5101
R1076 VDD.n11 VDD.t437 24.5101
R1077 VDD.n124 VDD.t445 24.4392
R1078 VDD.n246 VDD.t451 24.4392
R1079 VDD.n61 VDD.n33 22.154
R1080 VDD.n479 VDD.n148 19.8342
R1081 VDD.n467 VDD.n465 19.8342
R1082 VDD.n465 VDD.n163 19.829
R1083 VDD.n39 VDD.t7 17.002
R1084 VDD.n475 VDD.t162 14.0061
R1085 VDD.n62 VDD.n61 13.3957
R1086 VDD.n358 VDD.t236 13.2791
R1087 VDD.n467 VDD.n154 11.8712
R1088 VDD.n479 VDD.n477 11.8642
R1089 VDD VDD.t179 11.0624
R1090 VDD.t387 VDD.n347 10.7148
R1091 VDD.n197 VDD.n196 8.14083
R1092 VDD.n423 VDD.n174 8.03133
R1093 VDD.n200 VDD.n199 8.0005
R1094 VDD.n247 VDD.n246 8.0005
R1095 VDD.n458 VDD.t84 7.00657
R1096 VDD.n122 VDD.n121 6.98838
R1097 VDD.n243 VDD.n242 6.98838
R1098 VDD.n491 VDD.n488 6.76423
R1099 VDD.n82 VDD.n81 6.3005
R1100 VDD.n85 VDD.n78 6.3005
R1101 VDD.n88 VDD.n75 6.3005
R1102 VDD.n91 VDD.n73 6.3005
R1103 VDD.n132 VDD.n119 6.3005
R1104 VDD.n135 VDD.n116 6.3005
R1105 VDD.n138 VDD.n113 6.3005
R1106 VDD.n141 VDD.n111 6.3005
R1107 VDD.n410 VDD.n409 6.3005
R1108 VDD.n208 VDD.n207 6.3005
R1109 VDD.n210 VDD.n209 6.3005
R1110 VDD.n217 VDD.n216 6.3005
R1111 VDD.n219 VDD.n218 6.3005
R1112 VDD.n386 VDD.n385 6.3005
R1113 VDD.n388 VDD.n387 6.3005
R1114 VDD.n395 VDD.n394 6.3005
R1115 VDD.n397 VDD.n396 6.3005
R1116 VDD.n401 VDD.n400 6.3005
R1117 VDD.n402 VDD.n372 6.3005
R1118 VDD.n403 VDD.n368 6.3005
R1119 VDD.n404 VDD.n224 6.3005
R1120 VDD VDD.n337 6.3005
R1121 VDD.n251 VDD.n238 6.3005
R1122 VDD.n254 VDD.n235 6.3005
R1123 VDD.n257 VDD.n232 6.3005
R1124 VDD.n260 VDD.n230 6.3005
R1125 VDD.n280 VDD.n279 6.3005
R1126 VDD.n283 VDD.n276 6.3005
R1127 VDD.n286 VDD.n273 6.3005
R1128 VDD.n289 VDD.n271 6.3005
R1129 VDD.n360 VDD.n359 6.3005
R1130 VDD.n313 VDD.n312 6.3005
R1131 VDD.n309 VDD.n308 6.3005
R1132 VDD.n307 VDD.n306 6.3005
R1133 VDD.n293 VDD.n292 6.3005
R1134 VDD VDD.n425 6.3005
R1135 VDD.n455 VDD.n454 6.3005
R1136 VDD.n453 VDD.n452 6.3005
R1137 VDD.n446 VDD.n445 6.3005
R1138 VDD.n444 VDD.n443 6.3005
R1139 VDD VDD.n167 6.3005
R1140 VDD.n103 VDD.n102 6.3005
R1141 VDD.n98 VDD.n97 6.3005
R1142 VDD.n96 VDD.n95 6.3005
R1143 VDD.n30 VDD.n29 6.3005
R1144 VDD.n28 VDD.n27 6.3005
R1145 VDD.n21 VDD.n20 6.3005
R1146 VDD.n19 VDD.n18 6.3005
R1147 VDD.n64 VDD.n63 6.3005
R1148 VDD.n58 VDD.n33 6.3005
R1149 VDD.n39 VDD 6.3005
R1150 VDD.n54 VDD.n37 6.3005
R1151 VDD.n51 VDD.n33 6.3005
R1152 VDD VDD.n40 6.3005
R1153 VDD.n46 VDD.n33 6.3005
R1154 VDD.n45 VDD.n43 6.3005
R1155 VDD.n105 VDD.n104 6.3005
R1156 VDD VDD.n109 6.3005
R1157 VDD.n43 VDD.n40 6.18288
R1158 VDD.n418 VDD.t241 5.85907
R1159 VDD.n326 VDD.n325 5.85007
R1160 VDD.n488 VDD.n148 5.58865
R1161 VDD.n188 VDD.t303 5.21426
R1162 VDD.t199 VDD.n357 5.21426
R1163 VDD.t242 VDD.n348 5.21426
R1164 VDD.n82 VDD.t268 5.213
R1165 VDD.n385 VDD.n381 5.213
R1166 VDD.n280 VDD.t286 5.213
R1167 VDD.n66 VDD.n65 5.18745
R1168 VDD.n171 VDD.n170 5.16448
R1169 VDD.n101 VDD.t363 5.13287
R1170 VDD.n100 VDD.n68 5.13287
R1171 VDD.n99 VDD.t79 5.13287
R1172 VDD.n70 VDD.n69 5.13287
R1173 VDD.n94 VDD.t338 5.13287
R1174 VDD.n93 VDD.n71 5.13287
R1175 VDD.n84 VDD.t224 5.13287
R1176 VDD.n87 VDD.t125 5.13287
R1177 VDD.n89 VDD.n74 5.13287
R1178 VDD.n90 VDD.t428 5.13287
R1179 VDD.n92 VDD.n72 5.13287
R1180 VDD.n134 VDD.t299 5.13287
R1181 VDD.n137 VDD.t166 5.13287
R1182 VDD.n139 VDD.n112 5.13287
R1183 VDD.n140 VDD.t230 5.13287
R1184 VDD.n142 VDD.n110 5.13287
R1185 VDD.n485 VDD.n149 5.13287
R1186 VDD.n157 VDD.n155 5.13287
R1187 VDD.n472 VDD.t161 5.13287
R1188 VDD.n469 VDD.n159 5.13287
R1189 VDD.n164 VDD.t136 5.13287
R1190 VDD.n462 VDD.n165 5.13287
R1191 VDD.n459 VDD.t150 5.13287
R1192 VDD.n223 VDD.n222 5.13287
R1193 VDD.n193 VDD.n192 5.13287
R1194 VDD.n212 VDD.n189 5.13287
R1195 VDD.n215 VDD.t3 5.13287
R1196 VDD.n214 VDD.n213 5.13287
R1197 VDD.n220 VDD.t249 5.13287
R1198 VDD.n367 VDD.n225 5.13287
R1199 VDD.n370 VDD.t420 5.13287
R1200 VDD.n371 VDD.n369 5.13287
R1201 VDD.n374 VDD.t433 5.13287
R1202 VDD.n375 VDD.n373 5.13287
R1203 VDD.n399 VDD.t235 5.13287
R1204 VDD.n380 VDD.n379 5.13287
R1205 VDD.n390 VDD.n376 5.13287
R1206 VDD.n393 VDD.t435 5.13287
R1207 VDD.n392 VDD.n391 5.13287
R1208 VDD.n398 VDD.t111 5.13287
R1209 VDD.n342 VDD.t372 5.13287
R1210 VDD.n323 VDD.n322 5.13287
R1211 VDD.n352 VDD.t251 5.13287
R1212 VDD.n331 VDD.t49 5.13287
R1213 VDD.n351 VDD.n324 5.13287
R1214 VDD.n353 VDD.t393 5.13287
R1215 VDD.n361 VDD.t237 5.13287
R1216 VDD.n315 VDD.n228 5.13287
R1217 VDD.n253 VDD.t117 5.13287
R1218 VDD.n256 VDD.t324 5.13287
R1219 VDD.n258 VDD.n231 5.13287
R1220 VDD.n259 VDD.t239 5.13287
R1221 VDD.n261 VDD.n229 5.13287
R1222 VDD.n263 VDD.t381 5.13287
R1223 VDD.n310 VDD.t168 5.13287
R1224 VDD.n267 VDD.n266 5.13287
R1225 VDD.n305 VDD.t353 5.13287
R1226 VDD.n295 VDD.n268 5.13287
R1227 VDD.n294 VDD.t41 5.13287
R1228 VDD.n291 VDD.n269 5.13287
R1229 VDD.n282 VDD.t12 5.13287
R1230 VDD.n285 VDD.t348 5.13287
R1231 VDD.n287 VDD.n272 5.13287
R1232 VDD.n288 VDD.t374 5.13287
R1233 VDD.n290 VDD.n270 5.13287
R1234 VDD.n185 VDD.t175 5.13287
R1235 VDD.n416 VDD.n182 5.13287
R1236 VDD.n439 VDD.n433 5.13287
R1237 VDD.n432 VDD.n431 5.13287
R1238 VDD.n448 VDD.n428 5.13287
R1239 VDD.n451 VDD.t134 5.13287
R1240 VDD.n450 VDD.n449 5.13287
R1241 VDD.n456 VDD.t196 5.13287
R1242 VDD.n59 VDD.n57 5.13287
R1243 VDD.n32 VDD.t222 5.13287
R1244 VDD.n14 VDD.n9 5.13287
R1245 VDD.n8 VDD.n7 5.13287
R1246 VDD.n23 VDD.n4 5.13287
R1247 VDD.n26 VDD.t27 5.13287
R1248 VDD.n25 VDD.n24 5.13287
R1249 VDD.n31 VDD.t129 5.13287
R1250 VDD.n52 VDD.n38 5.13287
R1251 VDD.n50 VDD.t228 5.13287
R1252 VDD.n48 VDD.n41 5.13287
R1253 VDD.n44 VDD.t28 5.13287
R1254 VDD.n3 VDD.t359 5.13287
R1255 VDD.n47 VDD.n42 5.13287
R1256 VDD.n107 VDD.t99 5.13287
R1257 VDD.n146 VDD.n145 5.12339
R1258 VDD.n461 VDD.t403 5.12339
R1259 VDD.n470 VDD.t120 5.12339
R1260 VDD.n473 VDD.n158 5.12339
R1261 VDD.n156 VDD.t413 5.12339
R1262 VDD.n482 VDD.n150 5.12339
R1263 VDD.n484 VDD.t361 5.12339
R1264 VDD.n420 VDD.n180 5.11866
R1265 VDD.n417 VDD.t313 5.11866
R1266 VDD.n415 VDD.n183 5.11866
R1267 VDD.n408 VDD.t326 5.11866
R1268 VDD VDD.n34 5.11334
R1269 VDD VDD.t365 5.111
R1270 VDD VDD.t330 5.10321
R1271 VDD.n338 VDD.t173 5.09614
R1272 VDD.n492 VDD.n144 5.09407
R1273 VDD.n406 VDD.n221 5.09407
R1274 VDD.n341 VDD.n335 5.09407
R1275 VDD.n262 VDD.t180 5.09407
R1276 VDD.n427 VDD.n168 5.09407
R1277 VDD.n49 VDD.t8 5.09407
R1278 VDD.n299 VDD.n297 4.98388
R1279 VDD.n319 VDD.n318 4.95192
R1280 VDD.n301 VDD.t1 4.94512
R1281 VDD.n496 VDD.t86 4.93234
R1282 VDD.n131 VDD.t283 4.8755
R1283 VDD.n203 VDD.n202 4.8755
R1284 VDD.n250 VDD.t265 4.8755
R1285 VDD.n243 VDD.n239 4.51383
R1286 VDD.n246 VDD.n245 4.5005
R1287 VDD.n477 VDD.n154 4.47742
R1288 VDD.t240 VDD.n186 4.17151
R1289 VDD.n411 VDD.t174 4.17151
R1290 VDD.t392 VDD.n320 4.17151
R1291 VDD.n332 VDD.n329 4.12326
R1292 VDD.n421 VDD.t118 4.12326
R1293 VDD.n53 VDD.t10 4.12326
R1294 VDD.n437 VDD.n436 4.08796
R1295 VDD VDD.n10 4.08647
R1296 VDD.n435 VDD.n434 4.07925
R1297 VDD.n12 VDD.n11 4.0492
R1298 VDD.n126 VDD.n125 3.61662
R1299 VDD.n244 VDD.n240 3.61662
R1300 VDD.n13 VDD.n12 3.16779
R1301 VDD.n343 VDD.n328 3.1505
R1302 VDD.n336 VDD.n328 3.1505
R1303 VDD.n346 VDD.n345 3.1505
R1304 VDD.n347 VDD.n346 3.1505
R1305 VDD.n330 VDD.n327 3.1505
R1306 VDD.n348 VDD.n327 3.1505
R1307 VDD VDD.n350 3.1505
R1308 VDD.n350 VDD.n349 3.1505
R1309 VDD.n354 VDD.n321 3.1505
R1310 VDD.n321 VDD.n320 3.1505
R1311 VDD.n356 VDD.n355 3.1505
R1312 VDD.n357 VDD.n356 3.1505
R1313 VDD VDD.n181 3.1505
R1314 VDD.n187 VDD.n181 3.1505
R1315 VDD.n414 VDD.n184 3.1505
R1316 VDD.n188 VDD.n184 3.1505
R1317 VDD.n413 VDD.n412 3.1505
R1318 VDD.n412 VDD.n411 3.1505
R1319 VDD.n419 VDD.n175 3.1505
R1320 VDD.n186 VDD.n175 3.1505
R1321 VDD.n178 VDD.n174 3.1505
R1322 VDD.n174 VDD.n173 3.1505
R1323 VDD.n423 VDD.n422 3.1505
R1324 VDD.n424 VDD.n423 3.1505
R1325 VDD.n465 VDD.n463 3.1505
R1326 VDD.n465 VDD.n464 3.1505
R1327 VDD VDD.n491 3.1505
R1328 VDD.n491 VDD.n490 3.1505
R1329 VDD.n483 VDD.n148 3.1505
R1330 VDD.n148 VDD.n147 3.1505
R1331 VDD.n477 VDD.n474 3.1505
R1332 VDD.n477 VDD.n476 3.1505
R1333 VDD.n468 VDD.n467 3.1505
R1334 VDD.n467 VDD.n466 3.1505
R1335 VDD.n460 VDD.n163 3.1505
R1336 VDD.n166 VDD.n163 3.1505
R1337 VDD.n154 VDD.n153 3.1505
R1338 VDD.n480 VDD.n479 3.1505
R1339 VDD.n479 VDD.n478 3.1505
R1340 VDD.n488 VDD.n486 3.1505
R1341 VDD.n488 VDD.n487 3.1505
R1342 VDD.n438 VDD.n437 3.04332
R1343 VDD.n490 VDD.t137 3.0035
R1344 VDD.n13 VDD 2.99802
R1345 VDD.n438 VDD.n435 2.93635
R1346 VDD.n262 VDD.n261 2.87282
R1347 VDD.n2 VDD.n1 2.85787
R1348 VDD.n83 VDD.n80 2.85787
R1349 VDD.n86 VDD.n77 2.85787
R1350 VDD.n133 VDD.n118 2.85787
R1351 VDD.n136 VDD.n115 2.85787
R1352 VDD.n481 VDD.n152 2.85787
R1353 VDD.n206 VDD.n205 2.85787
R1354 VDD.n211 VDD.n191 2.85787
R1355 VDD.n366 VDD.n227 2.85787
R1356 VDD.n384 VDD.n383 2.85787
R1357 VDD.n389 VDD.n378 2.85787
R1358 VDD.n344 VDD.n334 2.85787
R1359 VDD.n252 VDD.n237 2.85787
R1360 VDD.n255 VDD.n234 2.85787
R1361 VDD.n311 VDD.n265 2.85787
R1362 VDD.n281 VDD.n278 2.85787
R1363 VDD.n284 VDD.n275 2.85787
R1364 VDD.n442 VDD.n441 2.85787
R1365 VDD.n447 VDD.n430 2.85787
R1366 VDD.n17 VDD.n16 2.85787
R1367 VDD.n22 VDD.n6 2.85787
R1368 VDD.n55 VDD.n36 2.85787
R1369 VDD.n162 VDD.n161 2.84839
R1370 VDD.n179 VDD.n177 2.84366
R1371 VDD.n362 VDD.n319 2.6555
R1372 VDD.n301 VDD.n300 2.543
R1373 VDD.n14 VDD.n13 2.28302
R1374 VDD.n1 VDD.t400 2.2755
R1375 VDD.n1 VDD.n0 2.2755
R1376 VDD.n80 VDD.t408 2.2755
R1377 VDD.n80 VDD.n79 2.2755
R1378 VDD.n77 VDD.t77 2.2755
R1379 VDD.n77 VDD.n76 2.2755
R1380 VDD.n118 VDD.t101 2.2755
R1381 VDD.n118 VDD.n117 2.2755
R1382 VDD.n115 VDD.t415 2.2755
R1383 VDD.n115 VDD.n114 2.2755
R1384 VDD.n152 VDD.t33 2.2755
R1385 VDD.n152 VDD.n151 2.2755
R1386 VDD.n205 VDD.t210 2.2755
R1387 VDD.n205 VDD.n204 2.2755
R1388 VDD.n191 VDD.t57 2.2755
R1389 VDD.n191 VDD.n190 2.2755
R1390 VDD.n227 VDD.t212 2.2755
R1391 VDD.n227 VDD.n226 2.2755
R1392 VDD.n383 VDD.t198 2.2755
R1393 VDD.n383 VDD.n382 2.2755
R1394 VDD.n378 VDD.t69 2.2755
R1395 VDD.n378 VDD.n377 2.2755
R1396 VDD.n334 VDD.t388 2.2755
R1397 VDD.n334 VDD.n333 2.2755
R1398 VDD.n237 VDD.t379 2.2755
R1399 VDD.n237 VDD.n236 2.2755
R1400 VDD.n234 VDD.t391 2.2755
R1401 VDD.n234 VDD.n233 2.2755
R1402 VDD.n265 VDD.t370 2.2755
R1403 VDD.n265 VDD.n264 2.2755
R1404 VDD.n278 VDD.t18 2.2755
R1405 VDD.n278 VDD.n277 2.2755
R1406 VDD.n275 VDD.t355 2.2755
R1407 VDD.n275 VDD.n274 2.2755
R1408 VDD.n177 VDD.t205 2.2755
R1409 VDD.n177 VDD.n176 2.2755
R1410 VDD.n441 VDD.t127 2.2755
R1411 VDD.n441 VDD.n440 2.2755
R1412 VDD.n430 VDD.t64 2.2755
R1413 VDD.n430 VDD.n429 2.2755
R1414 VDD.n161 VDD.t103 2.2755
R1415 VDD.n161 VDD.n160 2.2755
R1416 VDD.n16 VDD.t23 2.2755
R1417 VDD.n16 VDD.n15 2.2755
R1418 VDD.n6 VDD.t61 2.2755
R1419 VDD.n6 VDD.n5 2.2755
R1420 VDD.n36 VDD.t25 2.2755
R1421 VDD.n36 VDD.n35 2.2755
R1422 VDD.n439 VDD.n438 2.26327
R1423 VDD.n196 VDD.n195 2.11346
R1424 VDD.n121 VDD.n120 2.11318
R1425 VDD.n242 VDD.n241 2.11318
R1426 VDD.n187 VDD.t240 2.08601
R1427 VDD.n349 VDD.t242 2.08601
R1428 VDD.n304 VDD 1.92803
R1429 VDD.n198 VDD.n197 1.82345
R1430 VDD VDD.n223 1.81843
R1431 VDD.t252 VDD.n337 1.78621
R1432 VDD.n412 VDD.n184 1.62825
R1433 VDD.n356 VDD.n321 1.62825
R1434 VDD.n123 VDD.n122 1.54785
R1435 VDD.n245 VDD.n243 1.54785
R1436 VDD.n291 VDD.n290 1.24303
R1437 VDD.n93 VDD.n92 1.16167
R1438 VDD.n399 VDD.n398 1.16051
R1439 VDD.n32 VDD.n31 1.11953
R1440 VDD.n407 VDD.n220 1.0737
R1441 VDD.n143 VDD.n142 1.02091
R1442 VDD VDD.n457 0.993637
R1443 VDD.n125 VDD.n124 0.840632
R1444 VDD.n246 VDD.n240 0.840632
R1445 VDD.n340 VDD.n338 0.8375
R1446 VDD VDD.n107 0.631399
R1447 VDD.n43 VDD.n37 0.515698
R1448 VDD.n106 VDD 0.468962
R1449 VDD.n365 VDD 0.468385
R1450 VDD.n364 VDD.n316 0.453551
R1451 VDD.n315 VDD.n314 0.425188
R1452 VDD.n199 VDD.n198 0.404541
R1453 VDD.n300 VDD.n299 0.3805
R1454 VDD.n299 VDD.n298 0.3425
R1455 VDD.n132 VDD.n131 0.337997
R1456 VDD.n207 VDD.n203 0.337997
R1457 VDD.n251 VDD.n250 0.337997
R1458 VDD.n131 VDD.n130 0.328132
R1459 VDD.n203 VDD.n201 0.328132
R1460 VDD.n250 VDD.n249 0.328132
R1461 VDD VDD.n263 0.306125
R1462 VDD.n60 VDD.n59 0.2525
R1463 VDD.n87 VDD.n86 0.233919
R1464 VDD.n84 VDD.n83 0.233919
R1465 VDD.n137 VDD.n136 0.233919
R1466 VDD.n134 VDD.n133 0.233919
R1467 VDD.n206 VDD.n193 0.233919
R1468 VDD.n212 VDD.n211 0.233919
R1469 VDD.n384 VDD.n380 0.233919
R1470 VDD.n390 VDD.n389 0.233919
R1471 VDD.n256 VDD.n255 0.233919
R1472 VDD.n253 VDD.n252 0.233919
R1473 VDD.n285 VDD.n284 0.233919
R1474 VDD.n282 VDD.n281 0.233919
R1475 VDD.n442 VDD.n432 0.233919
R1476 VDD.n448 VDD.n447 0.233919
R1477 VDD.n17 VDD.n8 0.233919
R1478 VDD.n23 VDD.n22 0.233919
R1479 VDD.n295 VDD.n294 0.227375
R1480 VDD.n362 VDD.n361 0.202062
R1481 VDD.n319 VDD.n317 0.200877
R1482 VDD.n350 VDD.n327 0.200048
R1483 VDD VDD.n310 0.197375
R1484 VDD.n302 VDD.n301 0.192387
R1485 VDD.n497 VDD.n496 0.185237
R1486 VDD VDD.n67 0.183481
R1487 VDD.n311 VDD 0.1805
R1488 VDD.n293 VDD.n291 0.173
R1489 VDD.n306 VDD.n295 0.173
R1490 VDD.n309 VDD.n267 0.173
R1491 VDD.n181 VDD.n175 0.171541
R1492 VDD.n314 VDD.n262 0.1715
R1493 VDD VDD.n311 0.171125
R1494 VDD VDD.n364 0.169599
R1495 VDD VDD.n303 0.168064
R1496 VDD.n90 VDD.n89 0.141016
R1497 VDD.n94 VDD.n70 0.141016
R1498 VDD.n100 VDD.n99 0.141016
R1499 VDD.n140 VDD.n139 0.141016
R1500 VDD.n215 VDD.n214 0.141016
R1501 VDD.n393 VDD.n392 0.141016
R1502 VDD.n371 VDD.n370 0.141016
R1503 VDD.n375 VDD.n374 0.141016
R1504 VDD.n259 VDD.n258 0.141016
R1505 VDD.n288 VDD.n287 0.141016
R1506 VDD.n451 VDD.n450 0.141016
R1507 VDD.n26 VDD.n25 0.141016
R1508 VDD.n407 VDD.n406 0.139745
R1509 VDD.n457 VDD.n456 0.137919
R1510 VDD.n312 VDD.n263 0.129875
R1511 VDD.n408 VDD.n407 0.129213
R1512 VDD.n294 VDD 0.128
R1513 VDD VDD.n305 0.128
R1514 VDD.n310 VDD 0.128
R1515 VDD.n361 VDD 0.128
R1516 VDD.n316 VDD.n315 0.126125
R1517 VDD.n367 VDD 0.123016
R1518 VDD.n101 VDD 0.122435
R1519 VDD.n305 VDD.n304 0.1205
R1520 VDD VDD.n2 0.111984
R1521 VDD VDD.n366 0.111403
R1522 VDD.n196 VDD 0.107393
R1523 VDD.n304 VDD.n267 0.107375
R1524 VDD.n92 VDD.n91 0.107339
R1525 VDD.n89 VDD.n88 0.107339
R1526 VDD.n95 VDD.n93 0.107339
R1527 VDD.n98 VDD.n70 0.107339
R1528 VDD.n102 VDD.n100 0.107339
R1529 VDD.n142 VDD.n141 0.107339
R1530 VDD.n139 VDD.n138 0.107339
R1531 VDD.n216 VDD.n215 0.107339
R1532 VDD.n220 VDD.n219 0.107339
R1533 VDD.n394 VDD.n393 0.107339
R1534 VDD.n398 VDD.n397 0.107339
R1535 VDD.n370 VDD.n368 0.107339
R1536 VDD.n374 VDD.n372 0.107339
R1537 VDD.n400 VDD.n399 0.107339
R1538 VDD.n261 VDD.n260 0.107339
R1539 VDD.n258 VDD.n257 0.107339
R1540 VDD.n290 VDD.n289 0.107339
R1541 VDD.n287 VDD.n286 0.107339
R1542 VDD.n452 VDD.n451 0.107339
R1543 VDD.n456 VDD.n455 0.107339
R1544 VDD.n27 VDD.n26 0.107339
R1545 VDD.n31 VDD.n30 0.107339
R1546 VDD.n121 VDD 0.106795
R1547 VDD.n242 VDD 0.106795
R1548 VDD VDD.n206 0.106758
R1549 VDD.n211 VDD 0.106758
R1550 VDD VDD.n384 0.106758
R1551 VDD.n389 VDD 0.106758
R1552 VDD VDD.n442 0.106758
R1553 VDD.n447 VDD 0.106758
R1554 VDD VDD.n17 0.106758
R1555 VDD.n22 VDD 0.106758
R1556 VDD.n457 VDD.n427 0.106657
R1557 VDD.n86 VDD 0.106177
R1558 VDD.n83 VDD 0.106177
R1559 VDD.n136 VDD 0.106177
R1560 VDD.n133 VDD 0.106177
R1561 VDD.n255 VDD 0.106177
R1562 VDD.n252 VDD 0.106177
R1563 VDD.n284 VDD 0.106177
R1564 VDD.n281 VDD 0.106177
R1565 VDD.n364 VDD.n363 0.0842931
R1566 VDD.n409 VDD.n408 0.0841364
R1567 VDD.n85 VDD.n84 0.080629
R1568 VDD.n135 VDD.n134 0.080629
R1569 VDD.n210 VDD.n193 0.080629
R1570 VDD.n388 VDD.n380 0.080629
R1571 VDD.n254 VDD.n253 0.080629
R1572 VDD.n283 VDD.n282 0.080629
R1573 VDD.n443 VDD.n439 0.080629
R1574 VDD.n446 VDD.n432 0.080629
R1575 VDD.n18 VDD.n14 0.080629
R1576 VDD.n21 VDD.n8 0.080629
R1577 VDD VDD.n90 0.0794677
R1578 VDD VDD.n87 0.0794677
R1579 VDD VDD.n94 0.0794677
R1580 VDD.n99 VDD 0.0794677
R1581 VDD VDD.n101 0.0794677
R1582 VDD VDD.n140 0.0794677
R1583 VDD VDD.n137 0.0794677
R1584 VDD VDD.n259 0.0794677
R1585 VDD VDD.n256 0.0794677
R1586 VDD VDD.n288 0.0794677
R1587 VDD VDD.n285 0.0794677
R1588 VDD VDD.n212 0.0788871
R1589 VDD.n214 VDD 0.0788871
R1590 VDD VDD.n390 0.0788871
R1591 VDD.n392 VDD 0.0788871
R1592 VDD VDD.n367 0.0788871
R1593 VDD VDD.n371 0.0788871
R1594 VDD VDD.n375 0.0788871
R1595 VDD VDD.n448 0.0788871
R1596 VDD.n450 VDD 0.0788871
R1597 VDD VDD.n23 0.0788871
R1598 VDD.n25 VDD 0.0788871
R1599 VDD.n332 VDD.n331 0.078669
R1600 VDD.n344 VDD 0.0774014
R1601 VDD.n421 VDD.n420 0.0755
R1602 VDD.n351 VDD 0.0752887
R1603 VDD.n179 VDD 0.0746892
R1604 VDD.n129 VDD 0.0733571
R1605 VDD.n248 VDD 0.0733571
R1606 VDD VDD.n417 0.0726622
R1607 VDD.n406 VDD 0.0701226
R1608 VDD.n194 VDD 0.0690714
R1609 VDD.n426 VDD 0.0644908
R1610 VDD.n64 VDD.n32 0.0639483
R1611 VDD.n49 VDD.n48 0.0624822
R1612 VDD.n352 VDD.n351 0.0605
R1613 VDD.n314 VDD 0.0605
R1614 VDD.n460 VDD.n459 0.0590159
R1615 VDD.n55 VDD 0.0587712
R1616 VDD.n417 VDD.n416 0.0580676
R1617 VDD.n331 VDD 0.0579648
R1618 VDD.n486 VDD.n146 0.0575723
R1619 VDD.n107 VDD.n106 0.0562419
R1620 VDD.n298 VDD 0.0559545
R1621 VDD.n473 VDD.n472 0.0558357
R1622 VDD.n365 VDD.n223 0.0556613
R1623 VDD.n420 VDD 0.0552297
R1624 VDD.n481 VDD.n480 0.0545636
R1625 VDD.n468 VDD.n162 0.0545636
R1626 VDD VDD.n482 0.0542456
R1627 VDD VDD.n164 0.0539276
R1628 VDD.n60 VDD 0.0535198
R1629 VDD VDD.n426 0.0486123
R1630 VDD.n360 VDD.n316 0.047375
R1631 VDD.n130 VDD.n129 0.0471071
R1632 VDD.n201 VDD.n194 0.0471071
R1633 VDD.n249 VDD.n248 0.0471071
R1634 VDD VDD.n53 0.0447373
R1635 VDD VDD.n497 0.0438735
R1636 VDD VDD.n470 0.0437509
R1637 VDD VDD.n157 0.0434329
R1638 VDD.n353 VDD.n352 0.0427535
R1639 VDD.n323 VDD.n317 0.0419084
R1640 VDD.n300 VDD.n296 0.04175
R1641 VDD.n366 VDD.n365 0.0417258
R1642 VDD.n106 VDD.n2 0.0411452
R1643 VDD.n416 VDD.n415 0.0410405
R1644 VDD.n52 VDD 0.0410363
R1645 VDD.n343 VDD.n342 0.0407465
R1646 VDD.n51 VDD 0.0406311
R1647 VDD.n302 VDD.n185 0.0402297
R1648 VDD.n200 VDD.n197 0.0387493
R1649 VDD.n67 VDD.n3 0.0383305
R1650 VDD.n156 VDD 0.0377085
R1651 VDD.n469 VDD 0.0373905
R1652 VDD.n426 VDD.n171 0.0360046
R1653 VDD.n355 VDD.n323 0.035993
R1654 VDD.n354 VDD.n353 0.035993
R1655 VDD.n128 VDD.n127 0.0358571
R1656 VDD.n201 VDD.n200 0.0358571
R1657 VDD.n247 VDD.n239 0.0358571
R1658 VDD VDD.n60 0.0352781
R1659 VDD.n495 VDD.n494 0.0350652
R1660 VDD.n415 VDD.n414 0.0345541
R1661 VDD.n413 VDD.n185 0.0345541
R1662 VDD.n130 VDD.n128 0.03425
R1663 VDD.n249 VDD.n247 0.03425
R1664 VDD.n47 VDD 0.0325339
R1665 VDD VDD.n44 0.0310085
R1666 VDD.n157 VDD.n156 0.030394
R1667 VDD.n470 VDD.n469 0.030394
R1668 VDD.n56 VDD.n55 0.0300932
R1669 VDD.n340 VDD 0.0293152
R1670 VDD.n345 VDD.n344 0.0283873
R1671 VDD.n422 VDD.n179 0.0268514
R1672 VDD VDD.n340 0.0265156
R1673 VDD.n427 VDD 0.026125
R1674 VDD.n492 VDD 0.0256877
R1675 VDD.n58 VDD.n56 0.0238911
R1676 VDD.n46 VDD.n45 0.0236864
R1677 VDD.n493 VDD.n492 0.0235375
R1678 VDD.n484 VDD.n483 0.0233975
R1679 VDD.n463 VDD.n462 0.0233975
R1680 VDD VDD.n485 0.0227615
R1681 VDD.n461 VDD 0.0224435
R1682 VDD VDD.n146 0.0223089
R1683 VDD.n459 VDD.n458 0.0221254
R1684 VDD.n485 VDD.n484 0.0214894
R1685 VDD.n462 VDD.n461 0.0214894
R1686 VDD.n365 VDD.n224 0.0206923
R1687 VDD.n106 VDD.n105 0.0201154
R1688 VDD.n341 VDD 0.0197188
R1689 VDD.n178 VDD.n171 0.0179324
R1690 VDD.n53 VDD.n52 0.0172797
R1691 VDD.n497 VDD.n495 0.0156807
R1692 VDD VDD.n338 0.0153624
R1693 VDD VDD.n50 0.0146639
R1694 VDD.n12 VDD 0.0139888
R1695 VDD.n494 VDD.n493 0.0137082
R1696 VDD.n339 VDD.t172 0.0119124
R1697 VDD.n363 VDD.n317 0.0119085
R1698 VDD VDD.n332 0.0110634
R1699 VDD.n303 VDD.n302 0.0110405
R1700 VDD VDD.n421 0.0110405
R1701 VDD.n50 VDD.n49 0.0108279
R1702 VDD.n59 VDD 0.00985644
R1703 VDD.n48 VDD.n47 0.00965254
R1704 VDD.n44 VDD.n3 0.00965254
R1705 VDD.n437 VDD 0.00937324
R1706 VDD.n60 VDD.n56 0.00918812
R1707 VDD.n194 VDD 0.00907143
R1708 VDD.n298 VDD.n296 0.00731818
R1709 VDD.n435 VDD 0.00725
R1710 VDD.n67 VDD.n66 0.00716667
R1711 VDD.n494 VDD 0.00636957
R1712 VDD.n342 VDD.n341 0.00565625
R1713 VDD.n303 VDD.n296 0.0055
R1714 VDD.n482 VDD.n481 0.0049523
R1715 VDD.n164 VDD.n162 0.0049523
R1716 VDD.n129 VDD 0.00478571
R1717 VDD.n248 VDD 0.00478571
R1718 VDD VDD.n354 0.00430282
R1719 VDD.n414 VDD 0.00374324
R1720 VDD.n127 VDD.n126 0.00371429
R1721 VDD.n244 VDD.n239 0.00371429
R1722 VDD.n474 VDD.n473 0.00368021
R1723 VDD.n472 VDD.n471 0.00368021
R1724 VDD.n345 VDD 0.00345775
R1725 VDD.n422 VDD 0.00333784
R1726 VDD.n45 VDD 0.00294068
R1727 VDD.n66 VDD 0.00291379
R1728 VDD.n54 VDD 0.00263559
R1729 VDD.n330 VDD.n326 0.00261268
R1730 VDD.n493 VDD.n143 0.00259302
R1731 VDD VDD.n293 0.002375
R1732 VDD.n306 VDD 0.002375
R1733 VDD VDD.n309 0.002375
R1734 VDD.n312 VDD 0.002375
R1735 VDD VDD.n360 0.002375
R1736 VDD.n363 VDD.n362 0.002375
R1737 VDD.n216 VDD 0.00224194
R1738 VDD.n219 VDD 0.00224194
R1739 VDD.n394 VDD 0.00224194
R1740 VDD.n397 VDD 0.00224194
R1741 VDD.n368 VDD 0.00224194
R1742 VDD.n372 VDD 0.00224194
R1743 VDD.n400 VDD 0.00224194
R1744 VDD.n452 VDD 0.00224194
R1745 VDD.n455 VDD 0.00224194
R1746 VDD.n27 VDD 0.00224194
R1747 VDD.n30 VDD 0.00224194
R1748 VDD.n419 VDD.n418 0.00212162
R1749 VDD.n126 VDD.n123 0.00210714
R1750 VDD.n245 VDD.n244 0.00210714
R1751 VDD.n409 VDD 0.00186364
R1752 VDD VDD.n54 0.00172034
R1753 VDD VDD.n419 0.00171622
R1754 VDD VDD.n413 0.00171622
R1755 VDD.n91 VDD 0.00166129
R1756 VDD.n88 VDD 0.00166129
R1757 VDD VDD.n85 0.00166129
R1758 VDD VDD.n82 0.00166129
R1759 VDD.n95 VDD 0.00166129
R1760 VDD VDD.n98 0.00166129
R1761 VDD.n102 VDD 0.00166129
R1762 VDD.n141 VDD 0.00166129
R1763 VDD.n138 VDD 0.00166129
R1764 VDD VDD.n135 0.00166129
R1765 VDD VDD.n132 0.00166129
R1766 VDD.n260 VDD 0.00166129
R1767 VDD.n257 VDD 0.00166129
R1768 VDD VDD.n254 0.00166129
R1769 VDD VDD.n251 0.00166129
R1770 VDD.n289 VDD 0.00166129
R1771 VDD.n286 VDD 0.00166129
R1772 VDD VDD.n283 0.00166129
R1773 VDD VDD.n280 0.00166129
R1774 VDD VDD.n64 0.00153448
R1775 VDD.n474 VDD 0.00145406
R1776 VDD VDD.n468 0.00145406
R1777 VDD VDD.n460 0.00145406
R1778 VDD VDD.n46 0.00141525
R1779 VDD VDD.n51 0.00138525
R1780 VDD VDD.n343 0.00134507
R1781 VDD.n355 VDD 0.00134507
R1782 VDD VDD.n326 0.00134507
R1783 VDD VDD.n330 0.00134507
R1784 VDD.n418 VDD 0.00131081
R1785 VDD.n486 VDD 0.00113604
R1786 VDD.n480 VDD 0.00113604
R1787 VDD.n471 VDD 0.00113604
R1788 VDD.n463 VDD 0.00113604
R1789 VDD.n458 VDD 0.00113604
R1790 VDD.n207 VDD 0.00108064
R1791 VDD VDD.n210 0.00108064
R1792 VDD.n385 VDD 0.00108064
R1793 VDD VDD.n388 0.00108064
R1794 VDD.n443 VDD 0.00108064
R1795 VDD VDD.n446 0.00108064
R1796 VDD.n18 VDD 0.00108064
R1797 VDD VDD.n21 0.00108064
R1798 VDD.n224 VDD 0.00107692
R1799 VDD.n105 VDD 0.00107692
R1800 VDD VDD.n178 0.000905405
R1801 VDD.n483 VDD 0.000818021
R1802 VDD VDD.n58 0.000722772
R1803 CLK_div_3_mag_2.CLK.n13 CLK_div_3_mag_2.CLK.t14 36.935
R1804 CLK_div_3_mag_2.CLK.n12 CLK_div_3_mag_2.CLK.t8 36.935
R1805 CLK_div_3_mag_2.CLK.n7 CLK_div_3_mag_2.CLK.t2 36.935
R1806 CLK_div_3_mag_2.CLK.n6 CLK_div_3_mag_2.CLK.t6 36.935
R1807 CLK_div_3_mag_2.CLK.n4 CLK_div_3_mag_2.CLK.t4 30.6315
R1808 CLK_div_3_mag_2.CLK.n10 CLK_div_3_mag_2.CLK.t7 25.5364
R1809 CLK_div_3_mag_2.CLK.n8 CLK_div_3_mag_2.CLK.t12 25.5364
R1810 CLK_div_3_mag_2.CLK.n4 CLK_div_3_mag_2.CLK.t10 21.7275
R1811 CLK_div_3_mag_2.CLK.n13 CLK_div_3_mag_2.CLK.t13 18.1962
R1812 CLK_div_3_mag_2.CLK.n12 CLK_div_3_mag_2.CLK.t5 18.1962
R1813 CLK_div_3_mag_2.CLK.n7 CLK_div_3_mag_2.CLK.t15 18.1962
R1814 CLK_div_3_mag_2.CLK.n6 CLK_div_3_mag_2.CLK.t3 18.1962
R1815 CLK_div_3_mag_2.CLK.n10 CLK_div_3_mag_2.CLK.t11 14.0749
R1816 CLK_div_3_mag_2.CLK.n8 CLK_div_3_mag_2.CLK.t9 14.0749
R1817 CLK_div_3_mag_2.CLK.n17 CLK_div_3_mag_2.CLK.n16 9.33985
R1818 CLK_div_3_mag_2.CLK.n0 CLK_div_3_mag_2.CLK.n5 7.41537
R1819 CLK_div_3_mag_2.CLK.n11 CLK_div_3_mag_2.CLK.n9 5.37352
R1820 CLK_div_3_mag_2.CLK.n17 CLK_div_3_mag_2.CLK.n15 5.17836
R1821 CLK_div_3_mag_2.CLK CLK_div_3_mag_2.CLK.n14 4.53799
R1822 CLK_div_3_mag_2.CLK CLK_div_3_mag_2.CLK.n13 2.13042
R1823 CLK_div_3_mag_2.CLK CLK_div_3_mag_2.CLK.n3 0.0786548
R1824 CLK_div_3_mag_2.CLK.n7 CLK_div_3_mag_2.CLK.n3 2.13151
R1825 CLK_div_3_mag_2.CLK.n8 CLK_div_3_mag_2.CLK 1.4356
R1826 CLK_div_3_mag_2.CLK.n10 CLK_div_3_mag_2.CLK 1.4356
R1827 CLK_div_3_mag_2.CLK.n2 CLK_div_3_mag_2.CLK 0.0786553
R1828 CLK_div_3_mag_2.CLK.n2 CLK_div_3_mag_2.CLK.n12 2.13151
R1829 CLK_div_3_mag_2.CLK.n0 CLK_div_3_mag_2.CLK.n3 1.11863
R1830 CLK_div_3_mag_2.CLK.n2 CLK_div_3_mag_2.CLK.n1 1.11857
R1831 CLK_div_3_mag_2.CLK.n5 CLK_div_3_mag_2.CLK.n4 1.80477
R1832 CLK_div_3_mag_2.CLK.n0 CLK_div_3_mag_2.CLK 2.51975
R1833 CLK_div_3_mag_2.CLK CLK_div_3_mag_2.CLK.n6 2.13042
R1834 CLK_div_3_mag_2.CLK.n14 CLK_div_3_mag_2.CLK 1.77243
R1835 CLK_div_3_mag_2.CLK.n1 CLK_div_3_mag_2.CLK.n11 0.882595
R1836 CLK_div_3_mag_2.CLK.n17 CLK_div_3_mag_2.CLK 0.115328
R1837 CLK_div_3_mag_2.CLK.n5 CLK_div_3_mag_2.CLK 0.105737
R1838 CLK_div_3_mag_2.CLK.n11 CLK_div_3_mag_2.CLK 1.19627
R1839 CLK_div_3_mag_2.CLK.n9 CLK_div_3_mag_2.CLK 1.19627
R1840 CLK_div_3_mag_2.CLK.n9 CLK_div_3_mag_2.CLK.n0 1.01264
R1841 CLK_div_3_mag_2.CLK.n14 CLK_div_3_mag_2.CLK.n1 0.693045
R1842 CLK.n3 CLK.t12 36.935
R1843 CLK.n7 CLK.t8 36.935
R1844 CLK.n17 CLK.t13 36.935
R1845 CLK.n21 CLK.t3 36.935
R1846 CLK.n27 CLK.t5 30.5752
R1847 CLK.n34 CLK.t9 25.4744
R1848 CLK.n13 CLK.t6 25.4744
R1849 CLK.n27 CLK.t4 21.7814
R1850 CLK.n3 CLK.t10 18.1962
R1851 CLK.n7 CLK.t7 18.1962
R1852 CLK.n17 CLK.t11 18.1962
R1853 CLK.n21 CLK.t2 18.1962
R1854 CLK.n13 CLK.t0 14.1417
R1855 CLK.n34 CLK.t1 14.1417
R1856 CLK.n29 CLK.n28 7.41483
R1857 CLK.n39 CLK.n38 5.37091
R1858 CLK CLK.n0 2.27523
R1859 CLK.n40 CLK.n10 2.25253
R1860 CLK.n31 CLK.n20 2.25107
R1861 CLK.n37 CLK.n36 2.24352
R1862 CLK.n16 CLK.n15 2.24352
R1863 CLK.n24 CLK.n21 2.12464
R1864 CLK.n4 CLK.n3 2.12444
R1865 CLK.n8 CLK.n7 2.12188
R1866 CLK.n18 CLK.n17 2.12188
R1867 CLK.n28 CLK.n27 1.80883
R1868 CLK.n42 CLK.n41 1.66871
R1869 CLK.n40 CLK.n39 1.64153
R1870 CLK.n29 CLK.n26 1.59838
R1871 CLK.n5 CLK.n4 1.50528
R1872 CLK.n25 CLK.n24 1.50503
R1873 CLK.n14 CLK.n13 1.42118
R1874 CLK.n35 CLK.n34 1.42118
R1875 CLK CLK.n42 0.922951
R1876 CLK.n38 CLK.n31 0.882596
R1877 CLK.n33 CLK 0.1605
R1878 CLK.n30 CLK.n29 0.118826
R1879 CLK.n28 CLK 0.108371
R1880 CLK.n38 CLK.n37 0.0733415
R1881 CLK.n39 CLK.n16 0.0733415
R1882 CLK.n12 CLK 0.05925
R1883 CLK.n42 CLK.n6 0.0503214
R1884 CLK.n1 CLK 0.0457995
R1885 CLK.n9 CLK 0.0457995
R1886 CLK.n19 CLK 0.0457995
R1887 CLK.n22 CLK 0.0457995
R1888 CLK.n6 CLK.n5 0.0406786
R1889 CLK.n26 CLK.n25 0.0386356
R1890 CLK.n2 CLK.n1 0.0377414
R1891 CLK.n10 CLK.n9 0.0377414
R1892 CLK.n20 CLK.n19 0.0377414
R1893 CLK.n23 CLK.n22 0.0377414
R1894 CLK.n15 CLK.n12 0.03175
R1895 CLK.n36 CLK.n33 0.03175
R1896 CLK.n37 CLK.n32 0.0198632
R1897 CLK.n16 CLK.n11 0.0198632
R1898 CLK.n31 CLK.n30 0.0122182
R1899 CLK.n41 CLK.n40 0.0110646
R1900 CLK.n10 CLK.n8 0.00360345
R1901 CLK.n20 CLK.n18 0.00360345
R1902 CLK.n4 CLK.n2 0.00203744
R1903 CLK.n24 CLK.n23 0.00203726
R1904 CLK.n15 CLK.n14 0.00175
R1905 CLK.n36 CLK.n35 0.00175
R1906 Vdiv108.n1 Vdiv108.t4 36.935
R1907 Vdiv108.n3 Vdiv108.t6 31.4332
R1908 Vdiv108.n1 Vdiv108.t3 18.1962
R1909 Vdiv108.n3 Vdiv108.t5 15.3826
R1910 Vdiv108.n8 Vdiv108.t1 7.09905
R1911 Vdiv108.n4 Vdiv108.n3 6.86029
R1912 Vdiv108.n5 Vdiv108.n2 5.01077
R1913 Vdiv108.n8 Vdiv108.n7 3.25053
R1914 Vdiv108.n10 Vdiv108.n9 2.48821
R1915 Vdiv108.n7 Vdiv108.t0 2.2755
R1916 Vdiv108.n7 Vdiv108.n6 2.2755
R1917 Vdiv108 Vdiv108.n0 2.26091
R1918 Vdiv108.n2 Vdiv108.n1 2.13459
R1919 Vdiv108 Vdiv108.n10 1.64069
R1920 Vdiv108.n10 Vdiv108.n5 1.15502
R1921 Vdiv108.n5 Vdiv108.n4 1.12067
R1922 Vdiv108.n9 Vdiv108.n8 0.0905
R1923 Vdiv108.n4 Vdiv108 0.0857632
R1924 Vdiv108.n2 Vdiv108 0.0800273
R1925 Vdiv108.n9 Vdiv108 0.073625
R1926 CLK_div_3_mag_1.Q1.n5 CLK_div_3_mag_1.Q1.t4 36.935
R1927 CLK_div_3_mag_1.Q1.n2 CLK_div_3_mag_1.Q1.t5 31.4332
R1928 CLK_div_3_mag_1.Q1.n6 CLK_div_3_mag_1.Q1.t9 31.4332
R1929 CLK_div_3_mag_1.Q1.n3 CLK_div_3_mag_1.Q1.t6 30.4613
R1930 CLK_div_3_mag_1.Q1.n3 CLK_div_3_mag_1.Q1.t7 24.7562
R1931 CLK_div_3_mag_1.Q1.n5 CLK_div_3_mag_1.Q1.t3 18.1962
R1932 CLK_div_3_mag_1.Q1.n2 CLK_div_3_mag_1.Q1.t10 15.3826
R1933 CLK_div_3_mag_1.Q1.n6 CLK_div_3_mag_1.Q1.t8 15.3826
R1934 CLK_div_3_mag_1.Q1.n4 CLK_div_3_mag_1.Q1 8.5575
R1935 CLK_div_3_mag_1.Q1 CLK_div_3_mag_1.Q1.t0 7.09905
R1936 CLK_div_3_mag_1.Q1 CLK_div_3_mag_1.Q1.n6 6.86029
R1937 CLK_div_3_mag_1.Q1.n2 CLK_div_3_mag_1.Q1 5.69501
R1938 CLK_div_3_mag_1.Q1.n7 CLK_div_3_mag_1.Q1 5.01077
R1939 CLK_div_3_mag_1.Q1 CLK_div_3_mag_1.Q1.n1 3.25053
R1940 CLK_div_3_mag_1.Q1 CLK_div_3_mag_1.Q1.n8 2.43532
R1941 CLK_div_3_mag_1.Q1.n1 CLK_div_3_mag_1.Q1.t2 2.2755
R1942 CLK_div_3_mag_1.Q1.n1 CLK_div_3_mag_1.Q1.n0 2.2755
R1943 CLK_div_3_mag_1.Q1 CLK_div_3_mag_1.Q1.n5 2.13459
R1944 CLK_div_3_mag_1.Q1 CLK_div_3_mag_1.Q1.n3 1.81638
R1945 CLK_div_3_mag_1.Q1.n8 CLK_div_3_mag_1.Q1.n7 1.45395
R1946 CLK_div_3_mag_1.Q1.n8 CLK_div_3_mag_1.Q1.n4 1.23718
R1947 CLK_div_3_mag_1.Q1.n7 CLK_div_3_mag_1.Q1 1.12067
R1948 CLK_div_3_mag_1.Q1.n4 CLK_div_3_mag_1.Q1 0.976433
R1949 CLK_div_3_mag_1.JK_FF_mag_1.K.n3 CLK_div_3_mag_1.JK_FF_mag_1.K.t3 37.1981
R1950 CLK_div_3_mag_1.JK_FF_mag_1.K.n5 CLK_div_3_mag_1.JK_FF_mag_1.K.t5 31.4332
R1951 CLK_div_3_mag_1.JK_FF_mag_1.K.n4 CLK_div_3_mag_1.JK_FF_mag_1.K.t6 30.4613
R1952 CLK_div_3_mag_1.JK_FF_mag_1.K.n4 CLK_div_3_mag_1.JK_FF_mag_1.K.t7 24.7562
R1953 CLK_div_3_mag_1.JK_FF_mag_1.K.n3 CLK_div_3_mag_1.JK_FF_mag_1.K.t2 17.6611
R1954 CLK_div_3_mag_1.JK_FF_mag_1.K.n5 CLK_div_3_mag_1.JK_FF_mag_1.K.t4 15.3826
R1955 CLK_div_3_mag_1.JK_FF_mag_1.K.n0 CLK_div_3_mag_1.JK_FF_mag_1.K 12.0716
R1956 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.K.n5 7.62076
R1957 CLK_div_3_mag_1.JK_FF_mag_1.K.n6 CLK_div_3_mag_1.JK_FF_mag_1.K 6.09789
R1958 CLK_div_3_mag_1.JK_FF_mag_1.K.n7 CLK_div_3_mag_1.JK_FF_mag_1.K.n2 2.99416
R1959 CLK_div_3_mag_1.JK_FF_mag_1.K.n2 CLK_div_3_mag_1.JK_FF_mag_1.K.t1 2.2755
R1960 CLK_div_3_mag_1.JK_FF_mag_1.K.n2 CLK_div_3_mag_1.JK_FF_mag_1.K.n1 2.2755
R1961 CLK_div_3_mag_1.JK_FF_mag_1.K.n7 CLK_div_3_mag_1.JK_FF_mag_1.K.n6 2.2505
R1962 CLK_div_3_mag_1.JK_FF_mag_1.K.n0 CLK_div_3_mag_1.JK_FF_mag_1.K 2.24788
R1963 CLK_div_3_mag_1.JK_FF_mag_1.K.n6 CLK_div_3_mag_1.JK_FF_mag_1.K.n0 1.94903
R1964 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.K.n4 1.81638
R1965 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.K.n3 1.43706
R1966 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.K.n7 0.4325
R1967 CLK_div_3_mag_0.JK_FF_mag_1.K.n4 CLK_div_3_mag_0.JK_FF_mag_1.K.t7 37.1986
R1968 CLK_div_3_mag_0.JK_FF_mag_1.K.n3 CLK_div_3_mag_0.JK_FF_mag_1.K.t4 31.528
R1969 CLK_div_3_mag_0.JK_FF_mag_1.K.n2 CLK_div_3_mag_0.JK_FF_mag_1.K.t6 30.5184
R1970 CLK_div_3_mag_0.JK_FF_mag_1.K.n2 CLK_div_3_mag_0.JK_FF_mag_1.K.t8 24.7029
R1971 CLK_div_3_mag_0.JK_FF_mag_1.K.n4 CLK_div_3_mag_0.JK_FF_mag_1.K.t5 17.6614
R1972 CLK_div_3_mag_0.JK_FF_mag_1.K.n3 CLK_div_3_mag_0.JK_FF_mag_1.K.t3 15.3826
R1973 CLK_div_3_mag_0.JK_FF_mag_1.K.n0 CLK_div_3_mag_0.JK_FF_mag_1.K 12.0843
R1974 CLK_div_3_mag_0.JK_FF_mag_1.K.n0 CLK_div_3_mag_0.JK_FF_mag_1.K.n3 9.86691
R1975 CLK_div_3_mag_0.JK_FF_mag_1.K.n5 CLK_div_3_mag_0.JK_FF_mag_1.K 6.09789
R1976 CLK_div_3_mag_0.JK_FF_mag_1.K.n1 CLK_div_3_mag_0.JK_FF_mag_1.K.n7 2.99416
R1977 CLK_div_3_mag_0.JK_FF_mag_1.K.n7 CLK_div_3_mag_0.JK_FF_mag_1.K.t0 2.2755
R1978 CLK_div_3_mag_0.JK_FF_mag_1.K.n7 CLK_div_3_mag_0.JK_FF_mag_1.K.n6 2.2755
R1979 CLK_div_3_mag_0.JK_FF_mag_1.K.n1 CLK_div_3_mag_0.JK_FF_mag_1.K.n5 2.2505
R1980 CLK_div_3_mag_0.JK_FF_mag_1.K.n0 CLK_div_3_mag_0.JK_FF_mag_1.K 2.24173
R1981 CLK_div_3_mag_0.JK_FF_mag_1.K.n5 CLK_div_3_mag_0.JK_FF_mag_1.K.n0 1.93723
R1982 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.K.n2 1.81225
R1983 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.K.n4 1.43709
R1984 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.K.n1 0.281955
R1985 CLK_div_3_mag_1.Q0.n2 CLK_div_3_mag_1.Q0.t5 36.935
R1986 CLK_div_3_mag_1.Q0.n3 CLK_div_3_mag_1.Q0.t8 31.4332
R1987 CLK_div_3_mag_1.Q0.n5 CLK_div_3_mag_1.Q0.t7 29.8135
R1988 CLK_div_3_mag_1.Q0.n5 CLK_div_3_mag_1.Q0.t3 27.8352
R1989 CLK_div_3_mag_1.Q0.n2 CLK_div_3_mag_1.Q0.t4 18.1962
R1990 CLK_div_3_mag_1.Q0.n3 CLK_div_3_mag_1.Q0.t6 15.3826
R1991 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.Q0.t1 7.09905
R1992 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.Q0.n3 6.86029
R1993 CLK_div_3_mag_1.Q0.n4 CLK_div_3_mag_1.Q0 5.01077
R1994 CLK_div_3_mag_1.Q0.n6 CLK_div_3_mag_1.Q0 3.41843
R1995 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.Q0.n1 3.25053
R1996 CLK_div_3_mag_1.Q0.n1 CLK_div_3_mag_1.Q0.t0 2.2755
R1997 CLK_div_3_mag_1.Q0.n1 CLK_div_3_mag_1.Q0.n0 2.2755
R1998 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.Q0.n6 2.2505
R1999 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.Q0.n2 2.13459
R2000 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.Q0.n5 1.74998
R2001 CLK_div_3_mag_1.Q0.n6 CLK_div_3_mag_1.Q0.n4 1.50381
R2002 CLK_div_3_mag_1.Q0.n4 CLK_div_3_mag_1.Q0 1.12067
R2003 JK_FF_mag_0.Q.n3 JK_FF_mag_0.Q.t10 36.935
R2004 JK_FF_mag_0.Q.n7 JK_FF_mag_0.Q.t5 36.935
R2005 JK_FF_mag_0.Q.n6 JK_FF_mag_0.Q.t9 36.935
R2006 JK_FF_mag_0.Q.n4 JK_FF_mag_0.Q.t12 31.4332
R2007 JK_FF_mag_0.Q.n8 JK_FF_mag_0.Q.t3 25.4744
R2008 JK_FF_mag_0.Q.n3 JK_FF_mag_0.Q.t7 18.1962
R2009 JK_FF_mag_0.Q.n7 JK_FF_mag_0.Q.t4 18.1962
R2010 JK_FF_mag_0.Q.n6 JK_FF_mag_0.Q.t8 18.1962
R2011 JK_FF_mag_0.Q.n4 JK_FF_mag_0.Q.t11 15.3826
R2012 JK_FF_mag_0.Q.n8 JK_FF_mag_0.Q.t6 14.1417
R2013 JK_FF_mag_0.Q JK_FF_mag_0.Q.t1 7.09905
R2014 JK_FF_mag_0.Q JK_FF_mag_0.Q.n4 6.86029
R2015 JK_FF_mag_0.Q.n5 JK_FF_mag_0.Q 5.01077
R2016 JK_FF_mag_0.Q.n9 JK_FF_mag_0.Q 3.57531
R2017 JK_FF_mag_0.Q JK_FF_mag_0.Q.n2 3.25053
R2018 JK_FF_mag_0.Q.n2 JK_FF_mag_0.Q.t0 2.2755
R2019 JK_FF_mag_0.Q.n2 JK_FF_mag_0.Q.n1 2.2755
R2020 JK_FF_mag_0.Q JK_FF_mag_0.Q.n7 2.13265
R2021 JK_FF_mag_0.Q.n0 JK_FF_mag_0.Q 2.63776
R2022 JK_FF_mag_0.Q JK_FF_mag_0.Q.n9 2.3405
R2023 JK_FF_mag_0.Q JK_FF_mag_0.Q.n3 2.13459
R2024 JK_FF_mag_0.Q.n6 JK_FF_mag_0.Q 2.13261
R2025 JK_FF_mag_0.Q.n0 JK_FF_mag_0.Q 2.1039
R2026 JK_FF_mag_0.Q JK_FF_mag_0.Q.n8 1.59303
R2027 JK_FF_mag_0.Q.n9 JK_FF_mag_0.Q.n5 1.42999
R2028 JK_FF_mag_0.Q.n5 JK_FF_mag_0.Q 1.12067
R2029 JK_FF_mag_0.Q.n0 JK_FF_mag_0.Q 1.11863
C0 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 8.16e-20
C1 VDD a_4375_1354# 3.14e-19
C2 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 0.122f
C3 JK_FF_mag_1.nand2_mag_1.IN2 a_7192_2831# 0.069f
C4 a_9898_1318# a_10058_1318# 0.0504f
C5 CLK_div_3_mag_2.Q1 a_8887_265# 0.0157f
C6 Vdiv108 a_7038_3928# 0.00859f
C7 VDD CLK_div_3_mag_1.JK_FF_mag_1.K 2.48f
C8 RST a_4400_4955# 0.00135f
C9 JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 8.36e-22
C10 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.01e-20
C11 CLK_div_3_mag_2.Q1 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT 0.101f
C12 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_4369_213# 9.1e-19
C13 JK_FF_mag_0.nand2_mag_3.IN1 a_11307_2697# 0.00225f
C14 VDD CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 0.391f
C15 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_1.or_2_mag_0.IN2 5.32e-19
C16 CLK CLK_div_3_mag_0.Q0 0.00111f
C17 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0636f
C18 RST a_2101_3858# 0.00154f
C19 RST a_2107_4955# 0.00218f
C20 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_973_3858# 0.011f
C21 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand3_mag_1.OUT 0.16f
C22 JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 2.83e-19
C23 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 a_7035_221# 1.46e-19
C24 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 9.62e-20
C25 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.338f
C26 RST JK_FF_mag_1.nand3_mag_1.OUT 0.437f
C27 a_9892_221# a_10052_221# 0.0504f
C28 JK_FF_mag_1.nand2_mag_1.IN2 a_6628_2831# 0.00372f
C29 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT a_9892_221# 0.0202f
C30 Vdiv108 a_6474_3928# 0.0157f
C31 RST a_3836_4955# 5.68e-19
C32 Vdiv108 a_6628_2831# 0.069f
C33 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_5657_257# 0.00372f
C34 VDD a_1512_213# 9.21e-19
C35 VDD a_634_1310# 5.99e-19
C36 RST a_1537_3858# 3.39e-19
C37 CLK_div_3_mag_2.Q0 a_11904_265# 0.0157f
C38 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.or_2_mag_0.IN2 1.43e-20
C39 VDD CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT 0.661f
C40 CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C41 RST a_1543_4955# 0.00119f
C42 VDD JK_FF_mag_0.nand2_mag_4.IN2 0.391f
C43 JK_FF_mag_1.nand2_mag_3.IN1 a_8326_3928# 1.46e-19
C44 CLK_div_3_mag_0.Q0 a_5503_1354# 0.069f
C45 JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_1.K 0.00112f
C46 VDD CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 0.472f
C47 VDD a_3651_1310# 2.21e-19
C48 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand3_mag_2.OUT 0.0016f
C49 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_819_4955# 0.0036f
C50 JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_2.Q1 0.0127f
C51 CLK CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.471f
C52 CLK CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 2e-20
C53 CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 1.53e-19
C54 RST CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 0.515f
C55 Vdiv108 a_5278_3858# 8.04e-19
C56 RST a_7759_221# 0.00191f
C57 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00183f
C58 RST a_3272_4955# 0.00114f
C59 VDD JK_FF_mag_0.Q 2.38f
C60 CLK_div_3_mag_2.Q1 a_10616_221# 3.6e-22
C61 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.0445f
C62 JK_FF_mag_0.Q CLK_div_3_mag_2.JK_FF_mag_1.QB 1.35e-19
C63 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT a_7599_221# 9.1e-19
C64 VDD CLK_div_3_mag_1.JK_FF_mag_1.QB 0.881f
C65 RST CLK_div_3_mag_0.JK_FF_mag_1.K 0.478f
C66 VDD CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.471f
C67 CLK_div_3_mag_2.Q0 a_11340_265# 0.00859f
C68 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_5118_3858# 0.00119f
C69 RST CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.0034f
C70 JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 2.42e-20
C71 RST a_1383_4955# 0.00103f
C72 CLK_div_3_mag_2.Q0 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT 7.24e-19
C73 VDD CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 0.421f
C74 VDD a_9892_221# 0.00743f
C75 CLK_div_3_mag_0.Q1 a_2076_257# 0.00859f
C76 JK_FF_mag_1.nand2_mag_3.IN1 a_8320_2831# 0.00119f
C77 VDD a_2486_1354# 3.56e-19
C78 CLK_div_3_mag_0.Q1 a_794_1310# 2.79e-20
C79 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0175f
C80 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_1512_213# 0.0733f
C81 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 6.7e-19
C82 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 9.62e-20
C83 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 1.88e-20
C84 CLK_div_3_mag_2.or_2_mag_0.IN2 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 4.52e-20
C85 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.0894f
C86 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_409_3858# 4.52e-20
C87 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_1.QB 0.215f
C88 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C89 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 5.43e-19
C90 Vdiv108 a_5118_3858# 1.86e-20
C91 JK_FF_mag_1.nand3_mag_2.OUT JK_FF_mag_1.nand3_mag_1.OUT 0.121f
C92 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.QB 0.0373f
C93 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.nand2_mag_1.IN2 0.36f
C94 CLK_div_3_mag_0.JK_FF_mag_1.K a_4529_213# 0.00696f
C95 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.655f
C96 CLK_div_3_mag_2.Q1 a_10052_221# 1.86e-20
C97 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_1.K 0.00105f
C98 CLK_div_3_mag_2.Q1 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT 9.98e-19
C99 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 a_8887_265# 0.00372f
C100 CLK_div_3_mag_0.or_2_mag_0.IN2 a_5060_2689# 8.64e-19
C101 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_5284_4955# 0.0202f
C102 RST CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.226f
C103 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0948f
C104 RST a_10334_2461# 4.17e-19
C105 Vdiv108 JK_FF_mag_1.nand2_mag_3.IN1 0.0168f
C106 a_852_2291# CLK_div_3_mag_0.JK_FF_mag_1.QB 3.86e-19
C107 CLK_div_3_mag_2.Q0 a_10776_221# 0.0101f
C108 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_4554_3858# 1.43e-19
C109 VDD a_11307_2697# 0.165f
C110 VDD a_1922_1354# 3.14e-19
C111 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C112 JK_FF_mag_1.nand2_mag_3.IN1 a_7756_2831# 1.43e-19
C113 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C114 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 0.159f
C115 VDD JK_FF_mag_0.nand3_mag_1.OUT 0.998f
C116 a_5124_4955# a_5284_4955# 0.0504f
C117 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_0.Q0 0.0342f
C118 JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_2.Q0 0.0254f
C119 CLK CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 1.29f
C120 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_255_4955# 0.00372f
C121 RST a_1352_213# 8.64e-19
C122 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0894f
C123 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 4.7e-20
C124 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0854f
C125 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 4.44e-20
C126 CLK_div_3_mag_2.Q1 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 1.12e-19
C127 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 a_8169_1362# 0.0059f
C128 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_5124_4955# 0.0731f
C129 RST JK_FF_mag_1.QB 0.164f
C130 CLK_div_3_mag_2.Q0 a_10616_221# 0.0102f
C131 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_3990_3858# 0.011f
C132 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.0174f
C133 VDD a_4087_2453# 5.92e-19
C134 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C135 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.00169f
C136 JK_FF_mag_1.nand2_mag_3.IN1 a_7038_3928# 0.0036f
C137 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT a_10622_1362# 0.0202f
C138 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.765f
C139 VDD a_2640_257# 0.00142f
C140 CLK_div_3_mag_0.Q0 a_3811_1310# 2.79e-20
C141 CLK Vdiv108 0.0553f
C142 VDD a_1358_1354# 3.14e-19
C143 JK_FF_mag_1.nand2_mag_3.IN1 a_7192_2831# 0.011f
C144 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.802f
C145 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.QB 0.199f
C146 CLK_div_3_mag_2.Q1 CLK_div_3_mag_2.JK_FF_mag_1.QB 1.94f
C147 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 a_11750_1362# 0.00372f
C148 VDD CLK_div_3_mag_2.Q1 2.51f
C149 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.231f
C150 JK_FF_mag_0.nand3_mag_2.OUT a_11661_5045# 0.0202f
C151 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_4375_1354# 0.00378f
C152 CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_3_mag_0.JK_FF_mag_1.QB 8.53e-19
C153 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_1922_1354# 4.52e-20
C154 RST CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0734f
C155 JK_FF_mag_1.QB CLK_div_3_mag_2.JK_FF_mag_1.K 0.0125f
C156 RST JK_FF_mag_0.nand3_mag_2.OUT 0.0549f
C157 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 a_7605_1362# 0.0697f
C158 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_4560_4955# 9.1e-19
C159 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.K 0.69f
C160 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand3_mag_0.OUT 0.0622f
C161 RST a_8887_265# 0.00114f
C162 CLK_div_3_mag_2.Q0 a_10052_221# 0.00789f
C163 VDD CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 0.406f
C164 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_3426_3858# 0.00118f
C165 CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 0.0576f
C166 JK_FF_mag_0.Q JK_FF_mag_0.QB 1.99f
C167 CLK_div_3_mag_2.Q0 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT 0.338f
C168 CLK_div_3_mag_2.JK_FF_mag_1.K a_11904_265# 0.0811f
C169 VDD CLK_div_3_mag_0.Q1 2.48f
C170 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_5093_257# 0.0036f
C171 JK_FF_mag_1.nand2_mag_3.IN1 a_6628_2831# 0.00118f
C172 VDD a_11750_1362# 3.56e-19
C173 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.768f
C174 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.403f
C175 CLK CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 4.99e-21
C176 JK_FF_mag_0.QB CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 1.63e-20
C177 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand2_mag_1.IN2 8.16e-20
C178 RST CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT 0.00417f
C179 JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 4.87e-20
C180 CLK_div_3_mag_1.or_2_mag_0.IN2 a_852_2291# 8.64e-19
C181 CLK_div_3_mag_0.Q1 a_3645_213# 2.55e-20
C182 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 a_11186_1362# 0.069f
C183 JK_FF_mag_0.nand3_mag_2.OUT a_11501_5045# 0.0731f
C184 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_3811_1310# 0.0732f
C185 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_1358_1354# 0.0202f
C186 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.JK_FF_mag_1.K 0.00761f
C187 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.121f
C188 JK_FF_mag_1.QB CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 0.00208f
C189 JK_FF_mag_0.Q a_11495_3948# 2.79e-20
C190 a_5118_3858# a_5278_3858# 0.0504f
C191 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.Q1 3.97e-20
C192 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_4400_4955# 2.88e-20
C193 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.Q0 8.04e-19
C194 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 3.97e-21
C195 CLK_div_3_mag_0.JK_FF_mag_1.K a_5657_257# 0.0811f
C196 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C197 a_5060_2689# CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.132f
C198 CLK_div_3_mag_2.Q0 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 0.107f
C199 JK_FF_mag_0.Q JK_FF_mag_0.nand2_mag_1.IN2 0.11f
C200 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.nand3_mag_0.OUT 0.00183f
C201 JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 6.05e-20
C202 CLK_div_3_mag_2.JK_FF_mag_1.K a_11340_265# 0.00964f
C203 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 0.321f
C204 JK_FF_mag_1.nand3_mag_2.OUT JK_FF_mag_1.QB 0.103f
C205 VDD a_11186_1362# 3.14e-19
C206 RST a_10776_221# 0.00103f
C207 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT 0.352f
C208 VDD JK_FF_mag_0.nand3_mag_1.IN1 0.655f
C209 CLK_div_3_mag_1.or_2_mag_0.IN2 a_1825_2759# 7.48e-20
C210 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_5503_1354# 0.00372f
C211 JK_FF_mag_0.nand3_mag_2.OUT a_10937_5045# 9.1e-19
C212 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_3651_1310# 0.0203f
C213 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.QB 0.25f
C214 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_2.or_2_mag_0.IN2 0.124f
C215 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0343f
C216 VDD CLK_div_3_mag_2.Q0 1.27f
C217 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 8.58e-20
C218 RST JK_FF_mag_0.nand2_mag_3.IN1 0.219f
C219 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.653f
C220 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.995f
C221 RST a_2076_257# 0.0015f
C222 JK_FF_mag_0.Q a_8486_3928# 0.00166f
C223 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.QB 7.08e-20
C224 RST CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.103f
C225 CLK_div_3_mag_2.JK_FF_mag_1.K a_10776_221# 0.00696f
C226 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.0718f
C227 JK_FF_mag_1.nand2_mag_4.IN2 JK_FF_mag_1.nand3_mag_1.OUT 0.122f
C228 RST CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.207f
C229 JK_FF_mag_0.Q CLK_div_3_mag_2.or_2_mag_0.IN2 3.19e-19
C230 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_3645_213# 1.17e-20
C231 RST a_10616_221# 0.00119f
C232 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT 0.00183f
C233 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 2.34e-19
C234 a_973_3858# CLK_div_3_mag_1.or_2_mag_0.IN2 4.9e-20
C235 a_4400_4955# a_4560_4955# 0.0504f
C236 CLK a_5278_3858# 0.011f
C237 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 3.67e-20
C238 VDD a_3805_213# 0.00305f
C239 JK_FF_mag_0.nand2_mag_3.IN1 a_11501_5045# 1.46e-19
C240 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 4.44e-20
C241 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_4939_1354# 0.069f
C242 CLK_div_3_mag_2.or_2_mag_0.IN2 CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 0.0445f
C243 JK_FF_mag_0.nand3_mag_2.OUT a_10777_5045# 2.88e-20
C244 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 2.98e-19
C245 JK_FF_mag_1.QB CLK_div_3_mag_0.or_2_mag_0.IN2 5.72e-20
C246 CLK_div_3_mag_1.JK_FF_mag_1.K Vdiv108 0.172f
C247 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C248 JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_1.K 0.0257f
C249 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.198f
C250 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C251 a_3645_213# a_3805_213# 0.0504f
C252 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.359f
C253 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_3836_4955# 0.069f
C254 CLK a_1825_2759# 0.0103f
C255 a_2101_3858# a_2261_3858# 0.0504f
C256 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_4529_213# 8.64e-19
C257 CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 0.175f
C258 VDD CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 0.394f
C259 JK_FF_mag_1.nand2_mag_3.IN1 a_7041_1318# 3.41e-20
C260 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_794_1310# 0.0732f
C261 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 1.01e-20
C262 JK_FF_mag_0.nand2_mag_4.IN2 a_9803_3948# 4.52e-20
C263 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand3_mag_0.OUT 0.0893f
C264 JK_FF_mag_0.Q a_8326_3928# 0.00203f
C265 a_2107_4955# a_2267_4955# 0.0504f
C266 CLK_div_3_mag_2.JK_FF_mag_1.K a_10616_221# 0.00695f
C267 JK_FF_mag_0.Q a_8480_2831# 0.0101f
C268 RST a_10052_221# 0.00218f
C269 CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 1.99e-19
C270 JK_FF_mag_0.nand3_mag_1.OUT a_10931_3948# 0.0202f
C271 CLK a_5118_3858# 0.00939f
C272 RST CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT 0.0981f
C273 RST CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.278f
C274 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 7.08e-20
C275 CLK_div_3_mag_0.Q0 CLK_div_3_mag_2.Q1 8.2e-19
C276 JK_FF_mag_1.QB JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C277 CLK CLK_div_3_mag_1.or_2_mag_0.IN2 6.62e-20
C278 CLK_div_3_mag_2.or_2_mag_0.IN2 a_11307_2697# 8.64e-19
C279 JK_FF_mag_0.Q a_9803_3948# 0.069f
C280 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_3272_4955# 0.00372f
C281 CLK JK_FF_mag_1.nand2_mag_3.IN1 1.86e-20
C282 VDD JK_FF_mag_1.nand3_mag_1.IN1 0.655f
C283 CLK_div_3_mag_0.Q1 a_4369_213# 3.6e-22
C284 JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_2.or_2_mag_0.IN2 7.58e-20
C285 JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_1.QB 1.49e-19
C286 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT a_7035_221# 1.5e-20
C287 JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_2.Q1 8.13e-19
C288 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.JK_FF_mag_1.K 0.00205f
C289 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.Q0 0.0285f
C290 JK_FF_mag_0.Q a_8320_2831# 0.00939f
C291 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT 0.0881f
C292 JK_FF_mag_0.nand3_mag_1.OUT a_10367_3948# 4.52e-20
C293 a_409_3858# CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 4.94e-20
C294 a_11307_2697# CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 1.4e-19
C295 CLK a_4554_3858# 6.43e-21
C296 a_6881_1318# a_7041_1318# 0.0504f
C297 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.QB 0.21f
C298 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 3.67e-20
C299 CLK_div_3_mag_1.Q0 a_852_2291# 0.0134f
C300 JK_FF_mag_0.Q JK_FF_mag_1.nand2_mag_1.IN2 1.48e-20
C301 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 8.59e-20
C302 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.or_2_mag_0.IN2 0.0012f
C303 JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 1.18e-21
C304 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.QB 0.038f
C305 VDD a_11661_5045# 0.00108f
C306 JK_FF_mag_0.Q Vdiv108 0.157f
C307 a_5060_2689# CLK_div_3_mag_0.JK_FF_mag_1.K 0.00168f
C308 CLK_div_3_mag_1.JK_FF_mag_1.K a_6474_3928# 1.51e-20
C309 CLK_div_3_mag_2.Q1 CLK_div_3_mag_2.or_2_mag_0.IN2 0.0138f
C310 CLK_div_3_mag_1.JK_FF_mag_1.QB Vdiv108 1.18e-20
C311 VDD RST 3.81f
C312 JK_FF_mag_0.QB CLK_div_3_mag_2.Q0 0.00187f
C313 Vdiv108 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 2.48e-19
C314 RST CLK_div_3_mag_2.JK_FF_mag_1.QB 0.685f
C315 JK_FF_mag_0.Q a_7756_2831# 6.43e-21
C316 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 0.0725f
C317 RST a_3645_213# 0.00218f
C318 CLK_div_3_mag_0.JK_FF_mag_1.QB a_3811_1310# 1.41e-20
C319 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_4554_3858# 0.0697f
C320 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 8.16e-20
C321 CLK a_3990_3858# 6.06e-21
C322 CLK_div_3_mag_1.JK_FF_mag_1.K a_852_2291# 0.00168f
C323 a_10367_3948# CLK_div_3_mag_2.Q1 1.59e-20
C324 JK_FF_mag_0.nand2_mag_3.IN1 a_10213_5045# 0.0036f
C325 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_4369_213# 0.0203f
C326 JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 1.35e-20
C327 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.101f
C328 RST CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.313f
C329 JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 0.00176f
C330 JK_FF_mag_1.nand2_mag_4.IN2 JK_FF_mag_1.QB 0.199f
C331 CLK_div_3_mag_2.Q1 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT 0.338f
C332 CLK_div_3_mag_2.Q1 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 0.104f
C333 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C334 JK_FF_mag_1.QB CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.0025f
C335 VDD CLK_div_3_mag_2.JK_FF_mag_1.K 2.55f
C336 CLK_div_3_mag_1.JK_FF_mag_1.K a_5278_3858# 8.64e-19
C337 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0343f
C338 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 1.82e-19
C339 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_1.QB 3.28e-19
C340 CLK_div_3_mag_0.JK_FF_mag_1.QB a_1512_213# 0.00696f
C341 CLK CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.013f
C342 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.651f
C343 CLK CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.272f
C344 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.or_2_mag_0.IN2 0.0655f
C345 VDD JK_FF_mag_0.nand3_mag_0.OUT 0.745f
C346 CLK_div_3_mag_0.JK_FF_mag_1.QB a_3651_1310# 1.86e-20
C347 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_3990_3858# 0.0059f
C348 CLK a_3426_3858# 9.45e-19
C349 CLK_div_3_mag_0.Q0 a_3805_213# 0.00789f
C350 JK_FF_mag_0.nand3_mag_1.IN1 a_10931_3948# 0.0697f
C351 RST CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.345f
C352 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 0.122f
C353 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 a_11750_1362# 0.00118f
C354 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 0.122f
C355 CLK_div_3_mag_2.or_2_mag_0.IN2 a_11186_1362# 4.9e-20
C356 VDD a_10937_5045# 2.21e-19
C357 JK_FF_mag_1.QB a_5060_2689# 4.33e-20
C358 VDD CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 1.01f
C359 CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 0.21f
C360 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.00183f
C361 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT a_7759_221# 0.0733f
C362 a_1383_4955# a_1543_4955# 0.0504f
C363 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.or_2_mag_0.IN2 0.00761f
C364 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 a_409_3858# 0.00372f
C365 CLK_div_3_mag_2.or_2_mag_0.IN2 CLK_div_3_mag_2.Q0 0.0655f
C366 CLK_div_3_mag_0.JK_FF_mag_1.QB a_2486_1354# 0.0112f
C367 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C368 CLK CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 7.13e-22
C369 CLK_div_3_mag_1.JK_FF_mag_1.K a_973_3858# 2.96e-19
C370 VDD JK_FF_mag_1.nand3_mag_2.OUT 0.749f
C371 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0622f
C372 JK_FF_mag_0.nand3_mag_1.IN1 a_10367_3948# 0.0059f
C373 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 a_10776_221# 8.64e-19
C374 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0622f
C375 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 a_11186_1362# 0.011f
C376 CLK_div_3_mag_1.Q0 a_819_4955# 0.00859f
C377 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 9.52e-19
C378 JK_FF_mag_0.CLK CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 1.24e-19
C379 CLK_div_3_mag_1.Q0 CLK 0.149f
C380 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0129f
C381 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.Q1 1.25e-19
C382 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.359f
C383 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.JK_FF_mag_1.K 0.0103f
C384 JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 5.36e-22
C385 CLK_div_3_mag_2.Q0 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 0.0175f
C386 RST a_11655_3948# 1e-18
C387 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT a_7605_1362# 0.00378f
C388 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.QB 0.25f
C389 JK_FF_mag_0.Q JK_FF_mag_0.CLK 0.149f
C390 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.122f
C391 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.01e-20
C392 RST JK_FF_mag_0.QB 0.123f
C393 JK_FF_mag_0.CLK CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 0.131f
C394 CLK_div_3_mag_1.JK_FF_mag_1.K a_819_4955# 0.00964f
C395 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_5503_1354# 0.00118f
C396 RST a_4369_213# 0.00201f
C397 CLK CLK_div_3_mag_1.JK_FF_mag_1.K 2.12f
C398 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.JK_FF_mag_1.K 0.00967f
C399 CLK_div_3_mag_2.Q1 a_9898_1318# 0.00149f
C400 JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT 1.65e-19
C401 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 3.34e-19
C402 VDD a_10213_5045# 3.14e-19
C403 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 7.24e-19
C404 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0714f
C405 VDD CLK_div_3_mag_0.or_2_mag_0.IN2 0.494f
C406 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_5093_257# 0.00378f
C407 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 3.67e-20
C408 RST CLK_div_3_mag_0.Q0 0.16f
C409 RST a_11495_3948# 0.00108f
C410 VDD a_5657_257# 3.14e-19
C411 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT a_7041_1318# 0.0732f
C412 CLK_div_3_mag_1.JK_FF_mag_1.QB a_5118_3858# 0.00392f
C413 CLK_div_3_mag_0.JK_FF_mag_1.QB a_2640_257# 0.0811f
C414 CLK_div_3_mag_0.JK_FF_mag_1.QB a_1358_1354# 3.33e-19
C415 JK_FF_mag_0.QB CLK_div_3_mag_2.JK_FF_mag_1.K 3.27e-19
C416 JK_FF_mag_0.nand3_mag_0.OUT a_11655_3948# 0.0203f
C417 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.103f
C418 JK_FF_mag_1.QB CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 4.62e-20
C419 a_4369_213# a_4529_213# 0.0504f
C420 RST JK_FF_mag_0.nand2_mag_1.IN2 0.0387f
C421 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT 0.00169f
C422 JK_FF_mag_0.Q JK_FF_mag_1.nand2_mag_3.IN1 0.416f
C423 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_4939_1354# 0.011f
C424 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.K 8.58e-20
C425 a_1825_2759# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 7.3e-20
C426 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 5.8e-21
C427 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.12e-19
C428 JK_FF_mag_0.QB JK_FF_mag_0.nand3_mag_0.OUT 0.343f
C429 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 1.12e-19
C430 CLK_div_3_mag_2.Q1 a_6875_221# 0.00335f
C431 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.352f
C432 CLK_div_3_mag_2.Q1 a_8733_1362# 0.069f
C433 CLK_div_3_mag_0.Q0 a_4529_213# 0.0101f
C434 VDD JK_FF_mag_1.nand3_mag_0.OUT 0.746f
C435 VDD a_9649_5045# 3.14e-19
C436 JK_FF_mag_0.CLK JK_FF_mag_0.nand3_mag_1.OUT 6.64e-19
C437 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 0.122f
C438 CLK_div_3_mag_0.Q0 CLK_div_3_mag_2.JK_FF_mag_1.K 8.52e-20
C439 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.391f
C440 CLK_div_3_mag_2.Q0 a_10058_1318# 2.79e-20
C441 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.397f
C442 JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT 2.25e-20
C443 JK_FF_mag_0.QB a_10937_5045# 0.00695f
C444 RST a_10931_3948# 0.00237f
C445 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 a_8733_1362# 0.00372f
C446 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT a_6881_1318# 0.0203f
C447 CLK_div_3_mag_2.Q1 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 0.00335f
C448 CLK_div_3_mag_1.JK_FF_mag_1.QB a_4554_3858# 3.33e-19
C449 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_2267_4955# 0.0202f
C450 a_4554_3858# CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 7.41e-20
C451 JK_FF_mag_0.nand3_mag_0.OUT a_11495_3948# 0.0732f
C452 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_1.QB 1.94f
C453 RST CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.0233f
C454 RST a_8486_3928# 0.00312f
C455 RST CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00791f
C456 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C457 RST CLK_div_3_mag_2.or_2_mag_0.IN2 0.00261f
C458 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_4375_1354# 1.43e-19
C459 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C460 JK_FF_mag_0.QB JK_FF_mag_1.nand3_mag_2.OUT 3.32e-20
C461 VDD a_5284_4955# 0.0128f
C462 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.391f
C463 CLK CLK_div_3_mag_1.JK_FF_mag_1.QB 0.362f
C464 CLK CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 1.42e-19
C465 JK_FF_mag_0.CLK CLK_div_3_mag_2.Q1 2.53e-19
C466 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 6.11e-19
C467 RST a_10367_3948# 0.00278f
C468 CLK_div_3_mag_0.Q1 a_852_2291# 4.71e-21
C469 JK_FF_mag_0.QB a_10777_5045# 0.00696f
C470 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 a_8169_1362# 0.069f
C471 VDD CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 0.653f
C472 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_2107_4955# 0.0731f
C473 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.799f
C474 JK_FF_mag_0.nand3_mag_0.OUT a_10931_3948# 0.00378f
C475 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.JK_FF_mag_1.K 2.37f
C476 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 1.71e-20
C477 RST CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT 0.0981f
C478 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_5284_4955# 1.17e-20
C479 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C480 RST CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 0.00941f
C481 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C482 RST a_8326_3928# 0.00286f
C483 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_2267_4955# 1.17e-20
C484 CLK_div_3_mag_2.or_2_mag_0.IN2 CLK_div_3_mag_2.JK_FF_mag_1.K 0.00761f
C485 RST a_8480_2831# 0.00208f
C486 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_3811_1310# 0.00119f
C487 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C488 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.313f
C489 VDD a_409_3858# 3.56e-19
C490 JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_2.or_2_mag_0.IN2 4.5e-19
C491 VDD a_5124_4955# 0.00852f
C492 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.121f
C493 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.QB 0.0147f
C494 CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 1.43e-20
C495 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.00131f
C496 JK_FF_mag_1.nand3_mag_1.IN1 Vdiv108 0.00344f
C497 RST a_5093_257# 9.32e-19
C498 CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 2.81e-20
C499 VDD JK_FF_mag_1.nand2_mag_4.IN2 0.391f
C500 RST a_9803_3948# 0.0026f
C501 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT a_9892_221# 1.17e-20
C502 VDD CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.422f
C503 JK_FF_mag_0.QB a_10213_5045# 0.00964f
C504 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.393f
C505 JK_FF_mag_1.nand3_mag_1.IN1 a_7602_3928# 8.64e-19
C506 CLK a_1922_1354# 7.3e-20
C507 RST a_10622_1362# 1.9e-19
C508 JK_FF_mag_1.nand3_mag_1.IN1 a_7756_2831# 0.0697f
C509 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_1543_4955# 9.1e-19
C510 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 0.69f
C511 JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_2.Q1 4.62e-20
C512 CLK_div_3_mag_1.JK_FF_mag_1.QB a_3426_3858# 0.0112f
C513 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 1.53e-19
C514 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_5124_4955# 1.5e-20
C515 VDD a_7035_221# 0.00869f
C516 RST a_7762_3928# 0.0019f
C517 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 4.28e-21
C518 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_2107_4955# 1.5e-20
C519 JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 1.62e-20
C520 RST a_8320_2831# 0.00198f
C521 RST CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.136f
C522 JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 3.91e-20
C523 CLK_div_3_mag_2.Q1 a_7041_1318# 2.79e-20
C524 VDD a_4560_4955# 8.48e-19
C525 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.122f
C526 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.Q0 0.0655f
C527 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 1.88e-20
C528 JK_FF_mag_1.nand3_mag_2.OUT a_8486_3928# 0.0202f
C529 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.CLK 9.71e-20
C530 VDD a_255_4955# 3.14e-19
C531 RST JK_FF_mag_1.nand2_mag_1.IN2 0.00736f
C532 VDD a_2261_3858# 2.21e-19
C533 CLK_div_3_mag_2.Q1 a_7599_221# 0.0102f
C534 CLK_div_3_mag_0.Q0 a_5657_257# 0.0157f
C535 JK_FF_mag_0.QB a_9649_5045# 0.0811f
C536 a_8733_1362# CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 4.52e-20
C537 VDD a_5060_2689# 0.165f
C538 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.0435f
C539 JK_FF_mag_0.CLK CLK_div_3_mag_2.Q0 0.011f
C540 CLK_div_3_mag_2.JK_FF_mag_1.K a_10622_1362# 1.75e-19
C541 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT 0.00118f
C542 VDD a_2267_4955# 0.00743f
C543 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_1383_4955# 2.88e-20
C544 CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 3.24e-19
C545 RST Vdiv108 0.0576f
C546 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 3.67e-20
C547 RST a_10058_1318# 6.43e-19
C548 JK_FF_mag_1.nand3_mag_1.IN1 a_7192_2831# 0.0059f
C549 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_1537_3858# 0.0202f
C550 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_4560_4955# 0.0203f
C551 RST a_7602_3928# 0.00155f
C552 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_1543_4955# 0.0203f
C553 RST a_7756_2831# 0.00276f
C554 JK_FF_mag_0.nand2_mag_3.IN1 a_10334_2461# 2.95e-19
C555 JK_FF_mag_1.nand3_mag_2.OUT a_8326_3928# 0.0731f
C556 VDD a_4400_4955# 6.26e-19
C557 JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_2.JK_FF_mag_1.K 0.00701f
C558 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_2076_257# 0.0036f
C559 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_794_1310# 0.00119f
C560 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_4087_2453# 7.3e-20
C561 Vdiv108 CLK_div_3_mag_2.JK_FF_mag_1.K 0.0176f
C562 VDD a_2107_4955# 0.00305f
C563 CLK_div_3_mag_2.JK_FF_mag_1.K a_10058_1318# 0.00392f
C564 CLK CLK_div_3_mag_0.Q1 2.1e-19
C565 RST a_9898_1318# 7.78e-19
C566 VDD JK_FF_mag_1.nand3_mag_1.OUT 0.998f
C567 CLK CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.0215f
C568 JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_1.QB 4.62e-20
C569 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_4400_4955# 0.0733f
C570 RST CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00467f
C571 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.QB 3.28e-19
C572 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 6.11e-19
C573 a_8320_2831# CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 3.41e-20
C574 a_3651_1310# a_3811_1310# 0.0504f
C575 CLK_div_3_mag_2.Q1 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 4.33e-19
C576 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_1383_4955# 0.0733f
C577 VDD a_628_213# 0.0131f
C578 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 9.98e-19
C579 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0103f
C580 RST a_7192_2831# 0.00106f
C581 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.or_2_mag_0.IN2 1.82e-19
C582 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_3990_3858# 0.069f
C583 VDD a_3836_4955# 0.00107f
C584 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C585 JK_FF_mag_1.nand3_mag_2.OUT a_7762_3928# 9.1e-19
C586 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_788_213# 0.0731f
C587 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_973_3858# 0.0059f
C588 JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 3.91e-20
C589 CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 4.44e-20
C590 VDD a_1537_3858# 3.14e-19
C591 Vdiv108 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 4.62e-20
C592 VDD a_1543_4955# 2.21e-19
C593 RST CLK_div_3_mag_0.JK_FF_mag_1.QB 0.703f
C594 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.321f
C595 RST a_8733_1362# 0.00118f
C596 RST a_6875_221# 0.00187f
C597 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.Q1 3.22e-19
C598 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 5.8e-21
C599 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 4.28e-21
C600 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C601 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_3836_4955# 0.00378f
C602 VDD CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 1f
C603 JK_FF_mag_1.nand3_mag_2.OUT Vdiv108 0.338f
C604 RST a_6628_2831# 4.31e-19
C605 CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 0.214f
C606 JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 8.36e-22
C607 RST CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 0.313f
C608 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.nand2_mag_3.IN1 0.00118f
C609 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_3426_3858# 0.00372f
C610 VDD a_7759_221# 7.97e-19
C611 JK_FF_mag_0.Q JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C612 CLK_div_3_mag_2.JK_FF_mag_1.QB a_7759_221# 0.00696f
C613 JK_FF_mag_1.nand3_mag_2.OUT a_7602_3928# 2.88e-20
C614 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_2076_257# 0.069f
C615 CLK_div_3_mag_0.Q1 a_788_213# 0.00789f
C616 VDD a_3272_4955# 0.00107f
C617 JK_FF_mag_0.Q CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 0.00169f
C618 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_628_213# 1.17e-20
C619 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK 0.00254f
C620 CLK CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 6.77e-21
C621 VDD CLK_div_3_mag_0.JK_FF_mag_1.K 2.43f
C622 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.209f
C623 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C624 VDD CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.471f
C625 JK_FF_mag_0.CLK a_11661_5045# 0.00117f
C626 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT a_11186_1362# 4.52e-20
C627 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 3.34e-19
C628 RST a_8169_1362# 0.00149f
C629 JK_FF_mag_1.nand3_mag_0.OUT a_8480_2831# 0.0203f
C630 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.121f
C631 JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT 1.26e-20
C632 CLK_div_3_mag_2.Q1 a_8323_265# 0.00859f
C633 CLK_div_3_mag_0.Q0 a_7035_221# 1.24e-20
C634 a_6628_2831# CLK_div_3_mag_2.JK_FF_mag_1.K 4.41e-19
C635 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.or_2_mag_0.IN2 4.34e-20
C636 RST JK_FF_mag_0.CLK 0.00972f
C637 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand2_mag_3.IN1 0.233f
C638 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.104f
C639 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 8.58e-20
C640 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_1512_213# 8.64e-19
C641 CLK_div_3_mag_2.Q0 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 0.0343f
C642 CLK_div_3_mag_2.or_2_mag_0.IN2 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 1.82e-19
C643 CLK_div_3_mag_1.JK_FF_mag_1.K a_4087_2453# 5.05e-19
C644 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 4.28e-21
C645 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_3805_213# 0.0731f
C646 JK_FF_mag_0.Q CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 1.87e-21
C647 VDD CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 0.42f
C648 RST a_1825_2759# 4.83e-19
C649 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.01f
C650 Vdiv108 CLK_div_3_mag_0.or_2_mag_0.IN2 9.71e-19
C651 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_409_3858# 0.00118f
C652 VDD a_10334_2461# 5.92e-19
C653 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 1.88e-20
C654 CLK_div_3_mag_0.Q0 a_5060_2689# 0.0134f
C655 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.122f
C656 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 a_8733_1362# 0.00118f
C657 JK_FF_mag_0.CLK a_11501_5045# 0.00164f
C658 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN a_11307_2697# 3.25e-19
C659 RST a_7605_1362# 0.00232f
C660 JK_FF_mag_1.nand3_mag_0.OUT a_8320_2831# 0.0732f
C661 JK_FF_mag_0.CLK CLK_div_3_mag_2.JK_FF_mag_1.K 4.52e-19
C662 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand3_mag_1.OUT 0.122f
C663 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 9.62e-20
C664 JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 0.00169f
C665 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C666 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 0.231f
C667 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 5.43e-19
C668 a_10616_221# a_10776_221# 0.0504f
C669 RST CLK_div_3_mag_1.or_2_mag_0.IN2 9.28e-19
C670 JK_FF_mag_0.CLK JK_FF_mag_0.nand3_mag_0.OUT 0.267f
C671 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_5093_257# 0.069f
C672 VDD a_1352_213# 0.00114f
C673 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT 0.00183f
C674 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_0.Q1 0.0276f
C675 RST JK_FF_mag_1.nand2_mag_3.IN1 0.073f
C676 Vdiv108 JK_FF_mag_1.nand3_mag_0.OUT 7.24e-19
C677 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 8.58e-20
C678 VDD JK_FF_mag_1.QB 0.921f
C679 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C680 JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 2.25e-20
C681 JK_FF_mag_0.Q JK_FF_mag_0.nand3_mag_1.OUT 0.0345f
C682 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_1512_213# 2.88e-20
C683 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 a_8169_1362# 0.011f
C684 a_11307_2697# CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 0.132f
C685 a_11750_1362# CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 4.52e-20
C686 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_4939_1354# 4.52e-20
C687 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 3.81e-19
C688 JK_FF_mag_1.nand3_mag_0.OUT a_7756_2831# 0.00378f
C689 RST a_7041_1318# 0.00183f
C690 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C691 VDD a_11904_265# 3.14e-19
C692 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 a_10622_1362# 0.0697f
C693 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.159f
C694 CLK_div_3_mag_2.Q1 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT 7.24e-19
C695 RST a_7599_221# 0.0017f
C696 CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0012f
C697 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.Q0 0.00335f
C698 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT a_10776_221# 2.88e-20
C699 CLK_div_3_mag_2.Q1 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 0.305f
C700 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT a_7035_221# 0.0731f
C701 JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_1.K 0.223f
C702 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.394f
C703 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.00118f
C704 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_3805_213# 1.46e-19
C705 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_1922_1354# 0.0059f
C706 VDD JK_FF_mag_0.nand3_mag_2.OUT 0.746f
C707 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_4087_2453# 0.069f
C708 RST CLK 0.147f
C709 VDD a_8887_265# 0.00127f
C710 CLK_div_3_mag_0.Q1 a_1512_213# 0.0101f
C711 CLK_div_3_mag_2.JK_FF_mag_1.QB a_8887_265# 0.0811f
C712 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 a_7605_1362# 1.43e-19
C713 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_4375_1354# 0.0202f
C714 RST a_6881_1318# 0.00192f
C715 JK_FF_mag_0.Q CLK_div_3_mag_2.Q1 0.00787f
C716 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_1352_213# 0.0203f
C717 RST CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.126f
C718 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_2101_3858# 0.00119f
C719 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_5124_4955# 1.46e-19
C720 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT Vdiv108 2.14e-19
C721 VDD a_11340_265# 3.14e-19
C722 CLK_div_3_mag_0.Q1 a_3651_1310# 0.00149f
C723 RST a_3990_3858# 7.24e-19
C724 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_2107_4955# 1.46e-19
C725 VDD CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT 0.647f
C726 CLK_div_3_mag_0.JK_FF_mag_1.K a_4369_213# 0.00695f
C727 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.121f
C728 CLK_div_3_mag_2.Q1 CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 0.00139f
C729 CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT 2.81e-20
C730 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.K 0.0435f
C731 CLK_div_3_mag_2.Q0 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C732 CLK_div_3_mag_2.Q1 a_9892_221# 2.55e-20
C733 JK_FF_mag_0.Q CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 2e-19
C734 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 1.12e-19
C735 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT a_10616_221# 9.1e-19
C736 JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 5.2e-20
C737 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 a_8323_265# 0.069f
C738 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.313f
C739 JK_FF_mag_1.nand3_mag_1.OUT a_8486_3928# 1.17e-20
C740 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.399f
C741 JK_FF_mag_1.nand2_mag_4.IN2 JK_FF_mag_1.nand2_mag_1.IN2 8.16e-20
C742 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_1358_1354# 0.0697f
C743 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00147f
C744 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_1.K 2.37f
C745 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN JK_FF_mag_1.nand2_mag_1.IN2 1.64e-20
C746 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.666f
C747 RST CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 0.276f
C748 RST CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.196f
C749 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0576f
C750 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_4529_213# 2.88e-20
C751 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 a_7041_1318# 0.00119f
C752 JK_FF_mag_1.nand3_mag_2.OUT JK_FF_mag_1.nand2_mag_3.IN1 0.00118f
C753 CLK_div_3_mag_2.JK_FF_mag_1.K a_6881_1318# 8.64e-19
C754 Vdiv108 JK_FF_mag_1.nand2_mag_4.IN2 0.0635f
C755 RST CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.0054f
C756 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.305f
C757 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 8.16e-20
C758 CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.0576f
C759 JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 4.9e-22
C760 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.122f
C761 RST a_5503_1354# 6.6e-19
C762 Vdiv108 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.00224f
C763 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_1537_3858# 1.43e-19
C764 CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN a_11750_1362# 4.94e-20
C765 JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 0.00148f
C766 RST a_3426_3858# 0.00158f
C767 CLK_div_3_mag_0.Q1 a_2486_1354# 0.069f
C768 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.0622f
C769 CLK_div_3_mag_2.Q1 a_11307_2697# 6.83e-19
C770 JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 4.65e-20
C771 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT a_10052_221# 0.0731f
C772 JK_FF_mag_1.nand3_mag_1.OUT a_8326_3928# 1.5e-20
C773 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_2.Q0 8.04e-19
C774 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 0.23f
C775 VDD JK_FF_mag_0.nand2_mag_3.IN1 1.28f
C776 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00335f
C777 VDD a_2076_257# 0.00142f
C778 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.Q 0.00392f
C779 VDD a_794_1310# 2.65e-19
C780 Vdiv108 a_5060_2689# 0.00101f
C781 RST a_4939_1354# 6.6e-19
C782 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.653f
C783 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.739f
C784 JK_FF_mag_1.nand2_mag_4.IN2 a_7038_3928# 0.069f
C785 VDD a_10616_221# 2.21e-19
C786 RST CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.104f
C787 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 3.67e-20
C788 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.352f
C789 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 1.53e-19
C790 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN a_7192_2831# 2.85e-21
C791 JK_FF_mag_1.nand3_mag_1.OUT a_7762_3928# 0.0203f
C792 RST CLK_div_3_mag_1.Q0 0.0462f
C793 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT 0.121f
C794 CLK_div_3_mag_2.Q0 CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 0.209f
C795 RST a_8323_265# 5.68e-19
C796 CLK_div_3_mag_2.Q0 a_9892_221# 0.00335f
C797 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 6.11e-19
C798 JK_FF_mag_1.QB CLK_div_3_mag_0.Q0 0.0012f
C799 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT a_7759_221# 2.88e-20
C800 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 1.99e-19
C801 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C802 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 3.97e-21
C803 RST a_4375_1354# 5.8e-19
C804 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_3836_4955# 0.0036f
C805 CLK_div_3_mag_0.Q1 a_4087_2453# 0.01f
C806 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.QB 0.103f
C807 VDD a_10052_221# 0.00305f
C808 JK_FF_mag_1.nand2_mag_4.IN2 a_6474_3928# 0.00372f
C809 CLK_div_3_mag_0.Q1 a_2640_257# 0.0157f
C810 CLK_div_3_mag_2.Q1 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C811 Vdiv108 JK_FF_mag_1.nand3_mag_1.OUT 0.0343f
C812 VDD CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT 0.739f
C813 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.338f
C814 JK_FF_mag_1.nand2_mag_4.IN2 a_6628_2831# 4.52e-20
C815 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.nand3_mag_0.OUT 0.0886f
C816 CLK_div_3_mag_2.or_2_mag_0.IN2 a_10334_2461# 7.48e-20
C817 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.995f
C818 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_2076_257# 0.00378f
C819 a_6875_221# a_7035_221# 0.0504f
C820 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN a_6628_2831# 2.93e-20
C821 RST CLK_div_3_mag_1.JK_FF_mag_1.K 0.305f
C822 JK_FF_mag_1.nand3_mag_1.OUT a_7602_3928# 0.0733f
C823 CLK_div_3_mag_1.Q0 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 2.71e-20
C824 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand3_mag_1.OUT 0.768f
C825 JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT 0.00148f
C826 CLK_div_3_mag_2.Q0 a_11307_2697# 0.0134f
C827 JK_FF_mag_1.nand3_mag_1.OUT a_7756_2831# 0.0202f
C828 CLK CLK_div_3_mag_0.or_2_mag_0.IN2 1.1e-19
C829 CLK_div_3_mag_0.JK_FF_mag_1.K a_5093_257# 0.00964f
C830 RST CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 0.00239f
C831 RST a_3811_1310# 0.00141f
C832 VDD CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 0.399f
C833 JK_FF_mag_0.Q JK_FF_mag_1.nand3_mag_1.IN1 9.71e-20
C834 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.K 3.19e-19
C835 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_0.Q1 4.27e-19
C836 JK_FF_mag_1.nand3_mag_1.OUT a_7038_3928# 0.00378f
C837 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 a_8323_265# 0.0036f
C838 JK_FF_mag_1.nand3_mag_1.OUT a_7192_2831# 4.52e-20
C839 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_819_4955# 0.069f
C840 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 0.198f
C841 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.Q0 2.71e-20
C842 JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT 1.35e-20
C843 JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_2.Q1 0.00204f
C844 RST a_1512_213# 0.00218f
C845 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 2.98e-19
C846 CLK CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 7.33e-19
C847 RST CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT 0.0188f
C848 a_7756_2831# CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 3.85e-20
C849 RST JK_FF_mag_0.nand2_mag_4.IN2 0.00417f
C850 VDD CLK_div_3_mag_2.JK_FF_mag_1.QB 0.883f
C851 RST CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 0.00602f
C852 RST a_3651_1310# 0.00188f
C853 CLK_div_3_mag_2.Q1 CLK_div_3_mag_2.Q0 0.0285f
C854 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.QB 0.28f
C855 VDD a_3645_213# 0.00743f
C856 JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_2.or_2_mag_0.IN2 3.26e-21
C857 JK_FF_mag_0.Q a_11661_5045# 0.00335f
C858 CLK a_5284_4955# 0.00315f
C859 RST JK_FF_mag_0.Q 0.304f
C860 JK_FF_mag_1.nand2_mag_4.IN2 JK_FF_mag_1.nand2_mag_3.IN1 0.321f
C861 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 1f
C862 JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 3.68e-20
C863 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_634_1310# 0.0203f
C864 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT 0.0948f
C865 RST CLK_div_3_mag_1.JK_FF_mag_1.QB 0.598f
C866 JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 2.83e-19
C867 RST CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.00152f
C868 JK_FF_mag_0.nand2_mag_3.IN1 a_11495_3948# 0.00119f
C869 CLK_div_3_mag_2.Q0 a_11750_1362# 0.069f
C870 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C871 CLK_div_3_mag_0.or_2_mag_0.IN2 a_4939_1354# 4.9e-20
C872 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_2.JK_FF_mag_1.K 0.00384f
C873 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 5.32e-19
C874 RST a_9892_221# 0.00218f
C875 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00335f
C876 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 4.33e-19
C877 CLK CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.259f
C878 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C879 RST a_2486_1354# 0.00229f
C880 JK_FF_mag_1.QB a_7762_3928# 0.00695f
C881 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.0725f
C882 CLK_div_3_mag_2.Q1 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 0.0636f
C883 JK_FF_mag_1.QB a_8320_2831# 0.00392f
C884 JK_FF_mag_0.Q a_11501_5045# 0.00789f
C885 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.QB 0.00488f
C886 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1f
C887 JK_FF_mag_0.Q CLK_div_3_mag_2.JK_FF_mag_1.K 0.0251f
C888 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 a_11340_265# 0.0036f
C889 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT a_6875_221# 1.17e-20
C890 RST CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.264f
C891 CLK_div_3_mag_0.Q1 a_3805_213# 1.86e-20
C892 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 0.0894f
C893 CLK a_5124_4955# 0.00164f
C894 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 8.59e-20
C895 JK_FF_mag_1.QB JK_FF_mag_1.nand2_mag_1.IN2 0.0592f
C896 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 0.0854f
C897 JK_FF_mag_0.nand2_mag_3.IN1 a_10931_3948# 1.43e-19
C898 JK_FF_mag_0.Q JK_FF_mag_0.nand3_mag_0.OUT 8.96e-19
C899 CLK JK_FF_mag_1.nand2_mag_4.IN2 3.21e-20
C900 CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_2.JK_FF_mag_1.K 0.00205f
C901 a_5503_1354# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 4.52e-20
C902 CLK CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 6.4e-19
C903 Vdiv108 JK_FF_mag_1.QB 1.96f
C904 JK_FF_mag_0.nand3_mag_1.OUT a_11661_5045# 1.17e-20
C905 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.QB 3.28e-19
C906 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C907 CLK CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 5.57e-19
C908 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.00166f
C909 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 0.765f
C910 RST a_1922_1354# 0.00158f
C911 JK_FF_mag_1.QB a_7602_3928# 0.00696f
C912 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 a_7759_221# 8.64e-19
C913 RST JK_FF_mag_0.nand3_mag_1.OUT 0.427f
C914 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_0.or_2_mag_0.IN2 0.0107f
C915 JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_2.or_2_mag_0.IN2 0.00511f
C916 JK_FF_mag_1.QB a_7756_2831# 3.08e-19
C917 JK_FF_mag_0.Q a_10937_5045# 0.0102f
C918 JK_FF_mag_1.nand3_mag_1.OUT a_7605_1362# 3.85e-20
C919 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C920 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 9.52e-19
C921 JK_FF_mag_0.Q CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 6.3e-19
C922 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.122f
C923 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.122f
C924 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT a_10622_1362# 0.00378f
C925 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT a_8169_1362# 4.52e-20
C926 a_852_2291# CLK_div_3_mag_0.JK_FF_mag_1.K 0.00488f
C927 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN a_852_2291# 3.25e-19
C928 JK_FF_mag_0.nand2_mag_3.IN1 a_10367_3948# 0.011f
C929 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.JK_FF_mag_1.QB 5.46e-20
C930 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.21f
C931 CLK a_2261_3858# 0.0101f
C932 a_11307_2697# CLK_div_3_mag_2.JK_FF_mag_1.K 0.00168f
C933 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.nand3_mag_1.OUT 0.16f
C934 JK_FF_mag_0.Q JK_FF_mag_1.nand3_mag_2.OUT 0.235f
C935 JK_FF_mag_0.nand3_mag_1.OUT a_11501_5045# 1.5e-20
C936 RST a_4087_2453# 3.19e-19
C937 VDD a_11655_3948# 0.00478f
C938 CLK a_2267_4955# 0.00117f
C939 JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 1.07e-22
C940 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.321f
C941 RST a_1358_1354# 1.25e-19
C942 RST a_2640_257# 0.00114f
C943 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN a_5503_1354# 4.94e-20
C944 JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_1.K 1.77e-19
C945 RST CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.0566f
C946 JK_FF_mag_1.QB a_7038_3928# 0.00964f
C947 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_1.K 0.198f
C948 JK_FF_mag_1.QB a_7192_2831# 2.96e-19
C949 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_3805_213# 1.5e-20
C950 JK_FF_mag_0.Q a_10777_5045# 0.0101f
C951 VDD JK_FF_mag_0.QB 0.913f
C952 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.0854f
C953 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_3426_3858# 4.52e-20
C954 RST CLK_div_3_mag_2.Q1 0.12f
C955 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_0.OUT 0.0622f
C956 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN a_852_2291# 0.132f
C957 VDD a_4369_213# 2.21e-19
C958 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT a_10058_1318# 0.0732f
C959 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT a_7605_1362# 0.0202f
C960 JK_FF_mag_0.nand2_mag_4.IN2 a_10213_5045# 0.069f
C961 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.16f
C962 a_1825_2759# CLK_div_3_mag_0.JK_FF_mag_1.K 5.05e-19
C963 CLK_div_3_mag_0.JK_FF_mag_1.QB a_1352_213# 0.00695f
C964 JK_FF_mag_0.nand2_mag_3.IN1 a_9803_3948# 0.00118f
C965 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN a_1825_2759# 0.069f
C966 RST CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 0.00818f
C967 CLK a_2101_3858# 0.00939f
C968 VDD CLK_div_3_mag_0.Q0 1.3f
C969 JK_FF_mag_0.nand3_mag_1.OUT a_10937_5045# 0.0203f
C970 Vdiv108 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 1.09e-19
C971 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_2261_3858# 0.0203f
C972 CLK_div_3_mag_0.Q0 CLK_div_3_mag_2.JK_FF_mag_1.QB 3.93e-21
C973 CLK a_2107_4955# 0.00164f
C974 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_1358_1354# 0.00378f
C975 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00183f
C976 RST CLK_div_3_mag_0.Q1 0.379f
C977 JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 2.42e-20
C978 CLK JK_FF_mag_1.nand3_mag_1.OUT 1.29e-20
C979 JK_FF_mag_1.QB a_6474_3928# 0.0811f
C980 CLK_div_3_mag_1.Q0 a_409_3858# 0.069f
C981 CLK_div_3_mag_0.Q0 a_3645_213# 0.00335f
C982 RST CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.00557f
C983 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.99e-19
C984 JK_FF_mag_1.QB a_6628_2831# 0.0114f
C985 CLK_div_3_mag_2.Q1 CLK_div_3_mag_2.JK_FF_mag_1.K 0.363f
C986 JK_FF_mag_0.Q a_10213_5045# 0.00859f
C987 VDD JK_FF_mag_0.nand2_mag_1.IN2 0.402f
C988 JK_FF_mag_1.QB CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 1.49e-19
C989 CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_3_mag_0.JK_FF_mag_1.K 0.0107f
C990 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 a_10052_221# 1.46e-19
C991 CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.124f
C992 CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_0.or_2_mag_0.IN2 8.53e-19
C993 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT a_9898_1318# 0.0203f
C994 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT 9.52e-19
C995 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.or_2_mag_0.IN2 0.124f
C996 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_4400_4955# 8.64e-19
C997 JK_FF_mag_0.nand2_mag_4.IN2 a_9649_5045# 0.00372f
C998 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 1.01e-20
C999 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 8.58e-20
C1000 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.175f
C1001 CLK_div_3_mag_2.or_2_mag_0.IN2 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 3.81e-19
C1002 CLK a_1537_3858# 6.43e-21
C1003 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT a_7599_221# 0.0203f
C1004 JK_FF_mag_0.nand3_mag_1.OUT a_10777_5045# 0.0733f
C1005 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_2101_3858# 0.0732f
C1006 JK_FF_mag_1.QB a_8169_1362# 2.24e-20
C1007 VDD a_10931_3948# 3.14e-19
C1008 CLK_div_3_mag_0.JK_FF_mag_1.K a_7041_1318# 8.34e-21
C1009 CLK_div_3_mag_2.JK_FF_mag_1.K a_11750_1362# 0.012f
C1010 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 7.24e-19
C1011 a_7599_221# a_7759_221# 0.0504f
C1012 CLK_div_3_mag_1.JK_FF_mag_1.K a_409_3858# 0.012f
C1013 a_5060_2689# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.4e-19
C1014 CLK_div_3_mag_2.Q1 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 0.0177f
C1015 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_1.or_2_mag_0.IN2 0.0445f
C1016 JK_FF_mag_0.Q JK_FF_mag_1.nand3_mag_0.OUT 0.267f
C1017 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 1.08f
C1018 JK_FF_mag_0.nand3_mag_1.IN1 RST 0.253f
C1019 JK_FF_mag_0.Q a_9649_5045# 0.0157f
C1020 VDD a_8486_3928# 0.00108f
C1021 CLK_div_3_mag_1.Q0 a_255_4955# 0.0157f
C1022 CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 4.34e-20
C1023 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.647f
C1024 CLK_div_3_mag_1.JK_FF_mag_1.K JK_FF_mag_1.nand2_mag_4.IN2 6.03e-21
C1025 VDD CLK_div_3_mag_2.or_2_mag_0.IN2 0.495f
C1026 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.00967f
C1027 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C1028 RST CLK_div_3_mag_2.Q0 0.0447f
C1029 CLK_div_3_mag_1.Q0 a_2267_4955# 0.00335f
C1030 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 0.359f
C1031 CLK CLK_div_3_mag_0.JK_FF_mag_1.K 0.0194f
C1032 a_628_213# a_788_213# 0.0504f
C1033 RST CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.145f
C1034 RST CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.333f
C1035 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_1537_3858# 0.00378f
C1036 JK_FF_mag_0.nand3_mag_1.OUT a_10213_5045# 0.00378f
C1037 CLK CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.0983f
C1038 VDD a_10367_3948# 3.14e-19
C1039 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_2486_1354# 0.00372f
C1040 CLK_div_3_mag_0.JK_FF_mag_1.K a_6881_1318# 1.05e-20
C1041 CLK_div_3_mag_2.JK_FF_mag_1.K a_11186_1362# 2.96e-19
C1042 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0881f
C1043 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 6.02e-20
C1044 JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_1.K 1.64e-19
C1045 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.CLK 0.235f
C1046 VDD CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 1.08f
C1047 CLK_div_3_mag_1.JK_FF_mag_1.K a_255_4955# 0.0811f
C1048 VDD CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT 0.801f
C1049 CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT 0.103f
C1050 CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 7.08e-20
C1051 RST a_3805_213# 0.00218f
C1052 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C1053 VDD a_8480_2831# 0.00533f
C1054 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand3_mag_0.OUT 0.122f
C1055 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C1056 CLK_div_3_mag_1.JK_FF_mag_1.K a_5060_2689# 0.00488f
C1057 CLK_div_3_mag_1.Q0 a_2101_3858# 2.79e-20
C1058 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.QB 0.28f
C1059 CLK_div_3_mag_2.Q0 CLK_div_3_mag_2.JK_FF_mag_1.K 2.37f
C1060 CLK_div_3_mag_1.Q0 a_2107_4955# 0.00789f
C1061 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_4529_213# 0.0733f
C1062 CLK CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 7.03e-21
C1063 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 5.8e-21
C1064 CLK_div_3_mag_0.or_2_mag_0.IN2 a_4087_2453# 7.48e-20
C1065 RST CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 0.0576f
C1066 CLK CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 2.93e-19
C1067 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 1.88e-20
C1068 JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_2.Q0 3.94e-19
C1069 VDD a_5093_257# 3.14e-19
C1070 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_1.JK_FF_mag_1.QB 0.103f
C1071 VDD a_9803_3948# 3.56e-19
C1072 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_1922_1354# 0.069f
C1073 CLK_div_3_mag_0.JK_FF_mag_1.QB a_2076_257# 0.00964f
C1074 a_11495_3948# a_11655_3948# 0.0504f
C1075 CLK_div_3_mag_0.JK_FF_mag_1.QB a_794_1310# 0.00392f
C1076 CLK_div_3_mag_0.JK_FF_mag_1.K a_5503_1354# 0.012f
C1077 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 2.34e-19
C1078 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_5278_3858# 0.0203f
C1079 VDD a_10622_1362# 3.14e-19
C1080 JK_FF_mag_0.QB a_11495_3948# 0.00392f
C1081 VDD a_7762_3928# 2.21e-19
C1082 CLK_div_3_mag_1.JK_FF_mag_1.K a_2101_3858# 0.00392f
C1083 CLK_div_3_mag_0.Q0 a_4369_213# 0.0102f
C1084 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 1.02f
C1085 RST JK_FF_mag_1.nand3_mag_1.IN1 0.248f
C1086 CLK_div_3_mag_1.Q0 a_1543_4955# 0.0102f
C1087 JK_FF_mag_0.QB JK_FF_mag_0.nand2_mag_1.IN2 0.0592f
C1088 CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 5.46e-20
C1089 CLK JK_FF_mag_1.QB 0.00288f
C1090 VDD JK_FF_mag_1.nand2_mag_1.IN2 0.402f
C1091 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_1.QB 0.175f
C1092 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 3.34e-19
C1093 JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_2.JK_FF_mag_1.QB 1.49e-19
C1094 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.71e-20
C1095 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.or_2_mag_0.IN2 0.0138f
C1096 CLK_div_3_mag_0.JK_FF_mag_1.K a_4939_1354# 2.96e-19
C1097 JK_FF_mag_0.nand3_mag_1.IN1 a_10777_5045# 8.64e-19
C1098 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_1.or_2_mag_0.IN2 3.81e-19
C1099 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.159f
C1100 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.69f
C1101 JK_FF_mag_0.CLK JK_FF_mag_0.nand2_mag_3.IN1 0.421f
C1102 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_5118_3858# 0.0732f
C1103 VDD Vdiv108 1.17f
C1104 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT a_8323_265# 0.00378f
C1105 CLK_div_3_mag_2.JK_FF_mag_1.QB a_10058_1318# 1.41e-20
C1106 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 a_973_3858# 0.069f
C1107 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_788_213# 1.46e-19
C1108 JK_FF_mag_0.QB a_10931_3948# 3.12e-19
C1109 CLK_div_3_mag_1.JK_FF_mag_1.K a_1537_3858# 1.75e-19
C1110 CLK_div_3_mag_1.JK_FF_mag_1.QB a_4560_4955# 0.00695f
C1111 VDD a_7756_2831# 3.14e-19
C1112 JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_1.K 0.00244f
C1113 CLK_div_3_mag_1.Q0 CLK_div_3_mag_0.JK_FF_mag_1.K 0.0342f
C1114 CLK_div_3_mag_1.JK_FF_mag_1.K a_1543_4955# 0.00695f
C1115 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 8.04e-19
C1116 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 0.313f
C1117 CLK_div_3_mag_1.Q0 a_1383_4955# 0.0101f
C1118 CLK_div_3_mag_1.JK_FF_mag_1.QB a_2261_3858# 1.86e-20
C1119 JK_FF_mag_0.QB a_8486_3928# 1.36e-20
C1120 CLK_div_3_mag_1.JK_FF_mag_1.QB a_5060_2689# 3.86e-19
C1121 JK_FF_mag_0.QB CLK_div_3_mag_2.or_2_mag_0.IN2 1.03e-19
C1122 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_5060_2689# 3.25e-19
C1123 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.107f
C1124 CLK_div_3_mag_0.JK_FF_mag_1.K a_4375_1354# 1.75e-19
C1125 JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT 6.05e-20
C1126 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_4554_3858# 0.00378f
C1127 VDD a_9898_1318# 2.21e-19
C1128 CLK_div_3_mag_2.JK_FF_mag_1.QB a_9898_1318# 1.86e-20
C1129 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 0.208f
C1130 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 7.24e-19
C1131 a_11501_5045# a_11661_5045# 0.0504f
C1132 VDD a_7038_3928# 3.14e-19
C1133 JK_FF_mag_0.QB a_10367_3948# 2.96e-19
C1134 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.399f
C1135 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.K 0.107f
C1136 CLK_div_3_mag_1.JK_FF_mag_1.QB a_4400_4955# 0.00696f
C1137 CLK_div_3_mag_1.Q0 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 4.29e-20
C1138 VDD a_7192_2831# 3.14e-19
C1139 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.00384f
C1140 JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 4.87e-20
C1141 a_7192_2831# CLK_div_3_mag_2.JK_FF_mag_1.QB 2.24e-20
C1142 CLK_div_3_mag_2.Q1 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 6.7e-19
C1143 CLK CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 7.81e-19
C1144 CLK_div_3_mag_1.JK_FF_mag_1.K a_1383_4955# 0.00696f
C1145 JK_FF_mag_0.QB CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 5.36e-22
C1146 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 4.52e-20
C1147 RST a_4529_213# 0.00185f
C1148 CLK_div_3_mag_1.JK_FF_mag_1.QB a_2101_3858# 1.41e-20
C1149 JK_FF_mag_0.QB a_8326_3928# 1.07e-20
C1150 CLK CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.298f
C1151 RST CLK_div_3_mag_2.JK_FF_mag_1.K 0.318f
C1152 JK_FF_mag_0.Q JK_FF_mag_1.nand3_mag_1.OUT 6.64e-19
C1153 RST CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 9.92e-19
C1154 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand3_mag_2.OUT 0.00151f
C1155 CLK_div_3_mag_0.JK_FF_mag_1.K a_3811_1310# 0.00392f
C1156 VDD CLK_div_3_mag_0.JK_FF_mag_1.QB 0.879f
C1157 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT a_11340_265# 0.00378f
C1158 VDD a_8733_1362# 3.58e-19
C1159 VDD a_6875_221# 0.013f
C1160 RST JK_FF_mag_0.nand3_mag_0.OUT 0.0128f
C1161 CLK_div_3_mag_2.JK_FF_mag_1.QB a_8733_1362# 0.0112f
C1162 CLK_div_3_mag_0.Q0 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT 6.94e-19
C1163 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 0.00205f
C1164 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 0.0622f
C1165 JK_FF_mag_0.QB a_9803_3948# 0.0114f
C1166 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 0.0622f
C1167 VDD a_6474_3928# 3.14e-19
C1168 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 3.19e-19
C1169 JK_FF_mag_0.nand2_mag_1.IN2 a_10367_3948# 0.069f
C1170 CLK_div_3_mag_1.JK_FF_mag_1.QB a_3836_4955# 0.00964f
C1171 VDD a_6628_2831# 3.56e-19
C1172 VDD CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 0.659f
C1173 JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 4.9e-22
C1174 RST a_10937_5045# 0.00145f
C1175 CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 0.0135f
C1176 CLK_div_3_mag_0.JK_FF_mag_1.K a_634_1310# 8.64e-19
C1177 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.122f
C1178 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT 8.28e-21
C1179 CLK_div_3_mag_2.Q1 a_7035_221# 0.00789f
C1180 RST CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 0.19f
C1181 CLK_div_3_mag_0.Q0 a_5093_257# 0.00859f
C1182 VDD a_852_2291# 0.165f
C1183 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_1.or_2_mag_0.IN2 4.52e-20
C1184 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK 0.235f
C1185 JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_2.JK_FF_mag_1.K 2.85e-19
C1186 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_973_3858# 4.52e-20
C1187 CLK CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 1.64e-20
C1188 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.00139f
C1189 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT a_10776_221# 0.0733f
C1190 VDD a_8169_1362# 3.17e-19
C1191 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 a_11186_1362# 0.0059f
C1192 RST JK_FF_mag_1.nand3_mag_2.OUT 0.104f
C1193 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00169f
C1194 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 8.59e-20
C1195 VDD JK_FF_mag_0.CLK 1.66f
C1196 CLK_div_3_mag_1.JK_FF_mag_1.K JK_FF_mag_1.QB 0.00117f
C1197 JK_FF_mag_0.nand2_mag_1.IN2 a_9803_3948# 0.00372f
C1198 VDD a_5278_3858# 2.26e-19
C1199 JK_FF_mag_0.QB Vdiv108 1.89e-20
C1200 CLK_div_3_mag_1.JK_FF_mag_1.QB a_3272_4955# 0.0811f
C1201 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.Q0 4.29e-20
C1202 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.215f
C1203 RST a_10777_5045# 0.0015f
C1204 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.122f
C1205 JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 2e-21
C1206 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 0.0718f
C1207 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.JK_FF_mag_1.K 0.00384f
C1208 a_8326_3928# a_8486_3928# 0.0504f
C1209 CLK_div_3_mag_2.Q0 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 0.00335f
C1210 CLK_div_3_mag_2.or_2_mag_0.IN2 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 5.32e-19
C1211 VDD a_1825_2759# 5.92e-19
C1212 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN a_10334_2461# 0.069f
C1213 Vdiv108 CLK_div_3_mag_0.Q0 9.68e-19
C1214 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 a_11904_265# 0.00372f
C1215 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT a_10616_221# 0.0203f
C1216 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.71e-20
C1217 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.107f
C1218 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.00183f
C1219 CLK_div_3_mag_0.Q1 a_5060_2689# 6.83e-19
C1220 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_819_4955# 0.00378f
C1221 VDD a_7605_1362# 3.17e-19
C1222 CLK_div_3_mag_2.JK_FF_mag_1.QB a_7605_1362# 3.16e-19
C1223 CLK CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.00302f
C1224 VDD a_5118_3858# 2.65e-19
C1225 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand3_mag_0.OUT 0.122f
C1226 a_1352_213# a_1512_213# 0.0504f
C1227 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_628_213# 0.0202f
C1228 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 8.58e-20
C1229 JK_FF_mag_0.Q a_10334_2461# 1.13e-20
C1230 VDD CLK_div_3_mag_1.or_2_mag_0.IN2 0.494f
C1231 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00131f
C1232 RST a_10213_5045# 1.74e-19
C1233 VDD a_973_3858# 3.14e-19
C1234 VDD JK_FF_mag_1.nand2_mag_3.IN1 1.22f
C1235 JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_1.QB 0.00208f
C1236 RST a_5657_257# 9.58e-19
C1237 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 1.71e-20
C1238 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_2486_1354# 0.00118f
C1239 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 a_11340_265# 0.069f
C1240 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.0725f
C1241 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT a_10052_221# 1.5e-20
C1242 VDD a_7041_1318# 2.65e-19
C1243 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT 0.121f
C1244 CLK_div_3_mag_2.JK_FF_mag_1.QB a_7041_1318# 0.00392f
C1245 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_4939_1354# 0.0059f
C1246 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.107f
C1247 a_10777_5045# a_10937_5045# 0.0504f
C1248 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.0948f
C1249 VDD a_4554_3858# 3.18e-19
C1250 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.0622f
C1251 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C1252 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.231f
C1253 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 a_10622_1362# 1.43e-19
C1254 VDD a_7599_221# 0.00102f
C1255 JK_FF_mag_0.Q JK_FF_mag_1.QB 0.307f
C1256 Vdiv108 a_8486_3928# 0.00335f
C1257 CLK_div_3_mag_0.Q1 a_628_213# 0.00335f
C1258 CLK_div_3_mag_2.JK_FF_mag_1.QB a_7599_221# 0.00695f
C1259 CLK_div_3_mag_1.Q0 a_794_1310# 4.49e-20
C1260 RST JK_FF_mag_1.nand3_mag_0.OUT 0.0216f
C1261 RST a_9649_5045# 1.83e-19
C1262 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_1.Q0 0.338f
C1263 RST CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.00239f
C1264 RST CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0126f
C1265 CLK_div_3_mag_2.Q1 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 0.0343f
C1266 VDD a_819_4955# 3.14e-19
C1267 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_4554_3858# 0.0202f
C1268 a_8320_2831# a_8480_2831# 0.0504f
C1269 VDD CLK 2.5f
C1270 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_1922_1354# 0.011f
C1271 CLK_div_3_mag_2.Q1 a_7759_221# 0.0101f
C1272 CLK_div_3_mag_0.Q0 a_6875_221# 1.61e-20
C1273 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN a_1358_1354# 7.41e-20
C1274 VDD a_6881_1318# 2.25e-19
C1275 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C1276 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.739f
C1277 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_4375_1354# 0.0697f
C1278 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C1279 VDD a_3990_3858# 3.18e-19
C1280 JK_FF_mag_0.CLK a_11655_3948# 0.0101f
C1281 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 a_10058_1318# 0.00119f
C1282 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.Q 0.338f
C1283 Vdiv108 a_8326_3928# 0.00789f
C1284 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_3645_213# 0.0202f
C1285 JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_2.JK_FF_mag_1.K 0.00464f
C1286 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT 2.34e-19
C1287 CLK CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.00481f
C1288 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_1.JK_FF_mag_1.K 0.0881f
C1289 RST CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0254f
C1290 JK_FF_mag_0.CLK JK_FF_mag_0.QB 0.307f
C1291 a_2486_1354# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 4.52e-20
C1292 VDD CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 0.995f
C1293 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.0343f
C1294 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_1358_1354# 1.43e-19
C1295 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_3990_3858# 4.52e-20
C1296 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.66f
C1297 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00118f
C1298 RST CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 0.143f
C1299 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_1.K 0.362f
C1300 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.647f
C1301 RST CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.0545f
C1302 VDD a_5503_1354# 3.56e-19
C1303 CLK_div_3_mag_2.Q1 a_10334_2461# 0.01f
C1304 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.QB 3.24e-19
C1305 JK_FF_mag_0.CLK a_11495_3948# 0.00939f
C1306 VDD a_3426_3858# 3.59e-19
C1307 JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 1.65e-19
C1308 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 2.81e-20
C1309 VDD a_788_213# 0.00882f
C1310 Vdiv108 a_7762_3928# 0.0102f
C1311 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.765f
C1312 Vdiv108 a_8320_2831# 2.79e-20
C1313 CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C1314 a_7602_3928# a_7762_3928# 0.0504f
C1315 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 Vdiv108 0.00308f
C1316 JK_FF_mag_0.CLK JK_FF_mag_0.nand2_mag_1.IN2 1.48e-20
C1317 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand2_mag_3.IN1 0.321f
C1318 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_1537_3858# 0.0697f
C1319 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_1352_213# 9.1e-19
C1320 a_634_1310# a_794_1310# 0.0504f
C1321 RST JK_FF_mag_1.nand2_mag_4.IN2 0.00128f
C1322 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_1.K 0.23f
C1323 JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 0.00493f
C1324 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 0.0435f
C1325 JK_FF_mag_1.nand3_mag_2.OUT JK_FF_mag_1.nand3_mag_0.OUT 0.00183f
C1326 Vdiv108 JK_FF_mag_1.nand2_mag_1.IN2 0.107f
C1327 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0169f
C1328 RST CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.0582f
C1329 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_852_2291# 1.4e-19
C1330 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.nand3_mag_1.OUT 0.121f
C1331 VDD a_4939_1354# 3.14e-19
C1332 RST a_7035_221# 0.00187f
C1333 a_5118_3858# CLK_div_3_mag_0.Q0 4.49e-20
C1334 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.08f
C1335 JK_FF_mag_0.CLK a_10931_3948# 6.43e-21
C1336 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT a_6875_221# 0.0202f
C1337 JK_FF_mag_0.Q JK_FF_mag_0.nand2_mag_3.IN1 0.0261f
C1338 Vdiv108 a_7602_3928# 0.0101f
C1339 RST a_4560_4955# 8.64e-19
C1340 VDD CLK_div_3_mag_1.Q0 1.27f
C1341 JK_FF_mag_1.QB CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 1.49e-19
C1342 JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_2.JK_FF_mag_1.K 2.23e-19
C1343 VDD a_8323_265# 0.00127f
C1344 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.23f
C1345 CLK_div_3_mag_2.JK_FF_mag_1.QB a_8323_265# 0.00964f
C1346 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_2640_257# 0.00372f
C1347 JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 0.00461f
C1348 CLK_div_3_mag_0.Q1 a_1352_213# 0.0102f
C1349 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 6.02e-20
C1350 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 5.8e-21
C1351 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand3_mag_1.OUT 0.768f
C1352 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT 0.00154f
C1353 RST a_2261_3858# 0.00214f
C1354 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 4.28e-21
C1355 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_1383_4955# 8.64e-19
C1356 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 6.02e-20
C1357 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_788_213# 1.5e-20
C1358 RST a_2267_4955# 0.00218f
C1359 a_11904_265# VSS 0.0687f
C1360 a_11340_265# VSS 0.0688f
C1361 a_10776_221# VSS 0.0362f
C1362 a_10616_221# VSS 0.0901f
C1363 a_10052_221# VSS 0.0363f
C1364 a_9892_221# VSS 0.0901f
C1365 a_8887_265# VSS 0.0687f
C1366 a_8323_265# VSS 0.0688f
C1367 a_7759_221# VSS 0.0362f
C1368 a_7599_221# VSS 0.0901f
C1369 a_7035_221# VSS 0.0363f
C1370 a_6875_221# VSS 0.0901f
C1371 a_5657_257# VSS 0.0679f
C1372 a_5093_257# VSS 0.068f
C1373 a_4529_213# VSS 0.0349f
C1374 a_4369_213# VSS 0.0887f
C1375 a_3805_213# VSS 0.0349f
C1376 a_3645_213# VSS 0.0887f
C1377 a_2640_257# VSS 0.0679f
C1378 a_2076_257# VSS 0.068f
C1379 a_1512_213# VSS 0.0349f
C1380 a_1352_213# VSS 0.0887f
C1381 a_788_213# VSS 0.0349f
C1382 a_628_213# VSS 0.0887f
C1383 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.418f
C1384 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.547f
C1385 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.418f
C1386 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.527f
C1387 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.417f
C1388 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.542f
C1389 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.417f
C1390 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.522f
C1391 a_11750_1362# VSS 0.0676f
C1392 a_11186_1362# VSS 0.0676f
C1393 a_10622_1362# VSS 0.0676f
C1394 a_10058_1318# VSS 0.0343f
C1395 a_9898_1318# VSS 0.0881f
C1396 a_8733_1362# VSS 0.0676f
C1397 a_8169_1362# VSS 0.0676f
C1398 a_7605_1362# VSS 0.0676f
C1399 a_7041_1318# VSS 0.0343f
C1400 a_6881_1318# VSS 0.0881f
C1401 a_5503_1354# VSS 0.0676f
C1402 a_4939_1354# VSS 0.0676f
C1403 a_4375_1354# VSS 0.0676f
C1404 a_3811_1310# VSS 0.0343f
C1405 a_3651_1310# VSS 0.0881f
C1406 a_2486_1354# VSS 0.0676f
C1407 a_1922_1354# VSS 0.0676f
C1408 a_1358_1354# VSS 0.0676f
C1409 a_794_1310# VSS 0.0343f
C1410 a_634_1310# VSS 0.0891f
C1411 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.414f
C1412 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.691f
C1413 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.725f
C1414 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.816f
C1415 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C1416 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.41f
C1417 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.707f
C1418 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.721f
C1419 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.811f
C1420 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.505f
C1421 CLK_div_3_mag_2.JK_FF_mag_1.QB VSS 0.852f
C1422 CLK_div_3_mag_2.JK_FF_mag_1.K VSS 4.21f
C1423 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.414f
C1424 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.691f
C1425 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.725f
C1426 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.811f
C1427 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C1428 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.414f
C1429 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.697f
C1430 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.722f
C1431 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.808f
C1432 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.506f
C1433 CLK_div_3_mag_0.JK_FF_mag_1.QB VSS 0.855f
C1434 CLK_div_3_mag_0.JK_FF_mag_1.K VSS 4.46f
C1435 a_10334_2461# VSS 0.0676f
C1436 CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN VSS 0.594f
C1437 a_11307_2697# VSS 0.0247f
C1438 a_4087_2453# VSS 0.0676f
C1439 CLK_div_3_mag_2.Q0 VSS 1.97f
C1440 CLK_div_3_mag_2.or_2_mag_0.IN2 VSS 0.414f
C1441 a_8480_2831# VSS 0.0881f
C1442 a_8320_2831# VSS 0.0343f
C1443 a_7756_2831# VSS 0.0676f
C1444 a_7192_2831# VSS 0.0676f
C1445 a_6628_2831# VSS 0.0676f
C1446 JK_FF_mag_1.nand3_mag_0.OUT VSS 0.505f
C1447 JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.41f
C1448 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS 0.591f
C1449 a_5060_2689# VSS 0.0247f
C1450 a_852_2291# VSS 0.0261f
C1451 a_1825_2759# VSS 0.0726f
C1452 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN VSS 0.437f
C1453 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN VSS 0.429f
C1454 CLK_div_3_mag_2.Q1 VSS 1.74f
C1455 CLK_div_3_mag_0.Q0 VSS 1.7f
C1456 CLK_div_3_mag_0.or_2_mag_0.IN2 VSS 0.414f
C1457 CLK_div_3_mag_1.or_2_mag_0.IN2 VSS 0.419f
C1458 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN VSS 0.632f
C1459 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS 0.431f
C1460 CLK_div_3_mag_0.Q1 VSS 1.71f
C1461 a_11655_3948# VSS 0.0881f
C1462 a_11495_3948# VSS 0.0343f
C1463 a_10931_3948# VSS 0.0676f
C1464 a_10367_3948# VSS 0.0676f
C1465 a_9803_3948# VSS 0.0676f
C1466 JK_FF_mag_0.nand3_mag_0.OUT VSS 0.506f
C1467 JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.413f
C1468 a_8486_3928# VSS 0.0881f
C1469 a_8326_3928# VSS 0.0343f
C1470 a_7762_3928# VSS 0.0881f
C1471 a_7602_3928# VSS 0.0343f
C1472 a_7038_3928# VSS 0.0676f
C1473 a_6474_3928# VSS 0.0675f
C1474 a_5278_3858# VSS 0.0881f
C1475 a_5118_3858# VSS 0.0343f
C1476 a_4554_3858# VSS 0.0676f
C1477 a_3990_3858# VSS 0.0676f
C1478 a_3426_3858# VSS 0.0676f
C1479 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.506f
C1480 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.414f
C1481 JK_FF_mag_1.QB VSS 0.883f
C1482 JK_FF_mag_1.nand3_mag_1.OUT VSS 0.806f
C1483 JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.699f
C1484 JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.418f
C1485 a_2261_3858# VSS 0.0881f
C1486 a_2101_3858# VSS 0.0343f
C1487 a_1537_3858# VSS 0.0676f
C1488 a_973_3858# VSS 0.0676f
C1489 a_409_3858# VSS 0.0676f
C1490 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C1491 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.415f
C1492 Vdiv108 VSS 1.64f
C1493 JK_FF_mag_1.nand3_mag_2.OUT VSS 0.541f
C1494 JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.722f
C1495 a_11661_5045# VSS 0.0957f
C1496 a_11501_5045# VSS 0.0418f
C1497 a_10937_5045# VSS 0.0956f
C1498 a_10777_5045# VSS 0.0418f
C1499 a_10213_5045# VSS 0.0719f
C1500 a_9649_5045# VSS 0.0718f
C1501 a_5284_4955# VSS 0.0922f
C1502 a_5124_4955# VSS 0.0384f
C1503 a_4560_4955# VSS 0.0922f
C1504 a_4400_4955# VSS 0.0384f
C1505 a_3836_4955# VSS 0.0701f
C1506 a_3272_4955# VSS 0.07f
C1507 CLK_div_3_mag_1.JK_FF_mag_1.QB VSS 0.857f
C1508 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.819f
C1509 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.693f
C1510 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.42f
C1511 a_2267_4955# VSS 0.0922f
C1512 a_2107_4955# VSS 0.0384f
C1513 a_1543_4955# VSS 0.0922f
C1514 a_1383_4955# VSS 0.0384f
C1515 a_819_4955# VSS 0.0701f
C1516 a_255_4955# VSS 0.07f
C1517 CLK_div_3_mag_1.JK_FF_mag_1.K VSS 4.23f
C1518 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.823f
C1519 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.691f
C1520 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.42f
C1521 JK_FF_mag_0.QB VSS 0.899f
C1522 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.534f
C1523 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.722f
C1524 CLK VSS 2.9f
C1525 CLK_div_3_mag_1.Q0 VSS 2.78f
C1526 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.554f
C1527 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.726f
C1528 JK_FF_mag_0.nand3_mag_1.OUT VSS 0.828f
C1529 JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.733f
C1530 JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.422f
C1531 JK_FF_mag_0.CLK VSS 1.67f
C1532 JK_FF_mag_0.Q VSS 3.3f
C1533 JK_FF_mag_0.nand3_mag_2.OUT VSS 0.564f
C1534 RST VSS 7.08f
C1535 JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.721f
C1536 VDD VSS 0.125p
C1537 JK_FF_mag_0.Q.n0 VSS 0.234f
C1538 JK_FF_mag_0.Q.t1 VSS 0.0161f
C1539 JK_FF_mag_0.Q.t0 VSS 0.0133f
C1540 JK_FF_mag_0.Q.n1 VSS 0.0133f
C1541 JK_FF_mag_0.Q.n2 VSS 0.032f
C1542 JK_FF_mag_0.Q.t10 VSS 0.0297f
C1543 JK_FF_mag_0.Q.t7 VSS 0.0195f
C1544 JK_FF_mag_0.Q.n3 VSS 0.0527f
C1545 JK_FF_mag_0.Q.t12 VSS 0.0212f
C1546 JK_FF_mag_0.Q.t11 VSS 0.017f
C1547 JK_FF_mag_0.Q.n4 VSS 0.0494f
C1548 JK_FF_mag_0.Q.n5 VSS 0.389f
C1549 JK_FF_mag_0.Q.t9 VSS 0.0297f
C1550 JK_FF_mag_0.Q.t8 VSS 0.0195f
C1551 JK_FF_mag_0.Q.n6 VSS 0.0524f
C1552 JK_FF_mag_0.Q.t5 VSS 0.0297f
C1553 JK_FF_mag_0.Q.t4 VSS 0.0195f
C1554 JK_FF_mag_0.Q.n7 VSS 0.0524f
C1555 JK_FF_mag_0.Q.t3 VSS 0.0244f
C1556 JK_FF_mag_0.Q.t6 VSS 0.00633f
C1557 JK_FF_mag_0.Q.n8 VSS 0.0406f
C1558 JK_FF_mag_0.Q.n9 VSS 0.486f
C1559 CLK_div_3_mag_1.Q0.t1 VSS 0.025f
C1560 CLK_div_3_mag_1.Q0.t0 VSS 0.0206f
C1561 CLK_div_3_mag_1.Q0.n0 VSS 0.0206f
C1562 CLK_div_3_mag_1.Q0.n1 VSS 0.0494f
C1563 CLK_div_3_mag_1.Q0.t5 VSS 0.0459f
C1564 CLK_div_3_mag_1.Q0.t4 VSS 0.0302f
C1565 CLK_div_3_mag_1.Q0.n2 VSS 0.0814f
C1566 CLK_div_3_mag_1.Q0.t8 VSS 0.0329f
C1567 CLK_div_3_mag_1.Q0.t6 VSS 0.0263f
C1568 CLK_div_3_mag_1.Q0.n3 VSS 0.0764f
C1569 CLK_div_3_mag_1.Q0.n4 VSS 0.606f
C1570 CLK_div_3_mag_1.Q0.t7 VSS 0.0641f
C1571 CLK_div_3_mag_1.Q0.t3 VSS 0.0199f
C1572 CLK_div_3_mag_1.Q0.n5 VSS 0.0675f
C1573 CLK_div_3_mag_1.Q0.n6 VSS 0.447f
C1574 CLK_div_3_mag_0.JK_FF_mag_1.K.n0 VSS 2.09f
C1575 CLK_div_3_mag_0.JK_FF_mag_1.K.n1 VSS 0.202f
C1576 CLK_div_3_mag_0.JK_FF_mag_1.K.t6 VSS 0.0704f
C1577 CLK_div_3_mag_0.JK_FF_mag_1.K.t8 VSS 0.0546f
C1578 CLK_div_3_mag_0.JK_FF_mag_1.K.n2 VSS 0.139f
C1579 CLK_div_3_mag_0.JK_FF_mag_1.K.t3 VSS 0.0437f
C1580 CLK_div_3_mag_0.JK_FF_mag_1.K.t4 VSS 0.0547f
C1581 CLK_div_3_mag_0.JK_FF_mag_1.K.n3 VSS 0.141f
C1582 CLK_div_3_mag_0.JK_FF_mag_1.K.t7 VSS 0.0768f
C1583 CLK_div_3_mag_0.JK_FF_mag_1.K.t5 VSS 0.0489f
C1584 CLK_div_3_mag_0.JK_FF_mag_1.K.n4 VSS 0.136f
C1585 CLK_div_3_mag_0.JK_FF_mag_1.K.n5 VSS 1.17f
C1586 CLK_div_3_mag_0.JK_FF_mag_1.K.t0 VSS 0.0341f
C1587 CLK_div_3_mag_0.JK_FF_mag_1.K.n6 VSS 0.0341f
C1588 CLK_div_3_mag_0.JK_FF_mag_1.K.n7 VSS 0.0805f
C1589 CLK_div_3_mag_1.JK_FF_mag_1.K.n0 VSS 2.1f
C1590 CLK_div_3_mag_1.JK_FF_mag_1.K.t1 VSS 0.0349f
C1591 CLK_div_3_mag_1.JK_FF_mag_1.K.n1 VSS 0.0349f
C1592 CLK_div_3_mag_1.JK_FF_mag_1.K.n2 VSS 0.0745f
C1593 CLK_div_3_mag_1.JK_FF_mag_1.K.t3 VSS 0.0785f
C1594 CLK_div_3_mag_1.JK_FF_mag_1.K.t2 VSS 0.05f
C1595 CLK_div_3_mag_1.JK_FF_mag_1.K.n3 VSS 0.139f
C1596 CLK_div_3_mag_1.JK_FF_mag_1.K.t7 VSS 0.056f
C1597 CLK_div_3_mag_1.JK_FF_mag_1.K.t6 VSS 0.0719f
C1598 CLK_div_3_mag_1.JK_FF_mag_1.K.n4 VSS 0.143f
C1599 CLK_div_3_mag_1.JK_FF_mag_1.K.t5 VSS 0.0558f
C1600 CLK_div_3_mag_1.JK_FF_mag_1.K.t4 VSS 0.0447f
C1601 CLK_div_3_mag_1.JK_FF_mag_1.K.n5 VSS 0.133f
C1602 CLK_div_3_mag_1.JK_FF_mag_1.K.n6 VSS 1.19f
C1603 CLK_div_3_mag_1.JK_FF_mag_1.K.n7 VSS 0.218f
C1604 CLK_div_3_mag_1.Q1.t0 VSS 0.021f
C1605 CLK_div_3_mag_1.Q1.t2 VSS 0.0173f
C1606 CLK_div_3_mag_1.Q1.n0 VSS 0.0173f
C1607 CLK_div_3_mag_1.Q1.n1 VSS 0.0415f
C1608 CLK_div_3_mag_1.Q1.t5 VSS 0.0276f
C1609 CLK_div_3_mag_1.Q1.t10 VSS 0.0221f
C1610 CLK_div_3_mag_1.Q1.n2 VSS 0.0625f
C1611 CLK_div_3_mag_1.Q1.t7 VSS 0.0277f
C1612 CLK_div_3_mag_1.Q1.t6 VSS 0.0355f
C1613 CLK_div_3_mag_1.Q1.n3 VSS 0.0706f
C1614 CLK_div_3_mag_1.Q1.n4 VSS 0.321f
C1615 CLK_div_3_mag_1.Q1.t4 VSS 0.0385f
C1616 CLK_div_3_mag_1.Q1.t3 VSS 0.0254f
C1617 CLK_div_3_mag_1.Q1.n5 VSS 0.0684f
C1618 CLK_div_3_mag_1.Q1.t9 VSS 0.0276f
C1619 CLK_div_3_mag_1.Q1.t8 VSS 0.0221f
C1620 CLK_div_3_mag_1.Q1.n6 VSS 0.0642f
C1621 CLK_div_3_mag_1.Q1.n7 VSS 0.505f
C1622 CLK_div_3_mag_1.Q1.n8 VSS 0.209f
C1623 CLK.n0 VSS 0.0709f
C1624 CLK.n1 VSS 0.00877f
C1625 CLK.n2 VSS 0.00438f
C1626 CLK.t12 VSS 0.0528f
C1627 CLK.t10 VSS 0.0348f
C1628 CLK.n3 VSS 0.0933f
C1629 CLK.n4 VSS 0.0122f
C1630 CLK.n5 VSS 0.0151f
C1631 CLK.n6 VSS 0.00888f
C1632 CLK.t8 VSS 0.0528f
C1633 CLK.t7 VSS 0.0348f
C1634 CLK.n7 VSS 0.0933f
C1635 CLK.n8 VSS 0.0122f
C1636 CLK.n9 VSS 0.00877f
C1637 CLK.n10 VSS 0.00434f
C1638 CLK.n11 VSS 0.0188f
C1639 CLK.n12 VSS 0.0148f
C1640 CLK.t6 VSS 0.0436f
C1641 CLK.t0 VSS 0.0113f
C1642 CLK.n13 VSS 0.0722f
C1643 CLK.n14 VSS 0.0153f
C1644 CLK.n15 VSS 0.00533f
C1645 CLK.n16 VSS 0.0114f
C1646 CLK.t13 VSS 0.0528f
C1647 CLK.t11 VSS 0.0348f
C1648 CLK.n17 VSS 0.0933f
C1649 CLK.n18 VSS 0.0122f
C1650 CLK.n19 VSS 0.00877f
C1651 CLK.n20 VSS 0.00433f
C1652 CLK.t3 VSS 0.0528f
C1653 CLK.t2 VSS 0.0348f
C1654 CLK.n21 VSS 0.0933f
C1655 CLK.n22 VSS 0.00877f
C1656 CLK.n23 VSS 0.00438f
C1657 CLK.n24 VSS 0.0122f
C1658 CLK.n25 VSS 0.0172f
C1659 CLK.n26 VSS 0.163f
C1660 CLK.t4 VSS 0.0274f
C1661 CLK.t5 VSS 0.0489f
C1662 CLK.n27 VSS 0.0932f
C1663 CLK.n28 VSS 0.299f
C1664 CLK.n29 VSS 0.36f
C1665 CLK.n30 VSS 0.0135f
C1666 CLK.n31 VSS 0.101f
C1667 CLK.n32 VSS 0.0188f
C1668 CLK.n33 VSS 0.0314f
C1669 CLK.t9 VSS 0.0436f
C1670 CLK.t1 VSS 0.0113f
C1671 CLK.n34 VSS 0.0722f
C1672 CLK.n35 VSS 0.0153f
C1673 CLK.n36 VSS 0.00533f
C1674 CLK.n37 VSS 0.0114f
C1675 CLK.n38 VSS 0.667f
C1676 CLK.n39 VSS 0.709f
C1677 CLK.n40 VSS 0.0589f
C1678 CLK.n41 VSS 0.169f
C1679 CLK.n42 VSS 0.262f
C1680 CLK_div_3_mag_2.CLK.n0 VSS 0.456f
C1681 CLK_div_3_mag_2.CLK.n1 VSS 0.144f
C1682 CLK_div_3_mag_2.CLK.n2 VSS 0.0182f
C1683 CLK_div_3_mag_2.CLK.n3 VSS 0.0182f
C1684 CLK_div_3_mag_2.CLK.t10 VSS 0.023f
C1685 CLK_div_3_mag_2.CLK.t4 VSS 0.0414f
C1686 CLK_div_3_mag_2.CLK.n4 VSS 0.0788f
C1687 CLK_div_3_mag_2.CLK.n5 VSS 0.253f
C1688 CLK_div_3_mag_2.CLK.t3 VSS 0.0294f
C1689 CLK_div_3_mag_2.CLK.t6 VSS 0.0446f
C1690 CLK_div_3_mag_2.CLK.n6 VSS 0.0789f
C1691 CLK_div_3_mag_2.CLK.t15 VSS 0.0294f
C1692 CLK_div_3_mag_2.CLK.t2 VSS 0.0446f
C1693 CLK_div_3_mag_2.CLK.n7 VSS 0.0789f
C1694 CLK_div_3_mag_2.CLK.t12 VSS 0.0369f
C1695 CLK_div_3_mag_2.CLK.t9 VSS 0.00942f
C1696 CLK_div_3_mag_2.CLK.n8 VSS 0.0611f
C1697 CLK_div_3_mag_2.CLK.n9 VSS 0.588f
C1698 CLK_div_3_mag_2.CLK.t7 VSS 0.0369f
C1699 CLK_div_3_mag_2.CLK.t11 VSS 0.00942f
C1700 CLK_div_3_mag_2.CLK.n10 VSS 0.0611f
C1701 CLK_div_3_mag_2.CLK.n11 VSS 0.587f
C1702 CLK_div_3_mag_2.CLK.t5 VSS 0.0294f
C1703 CLK_div_3_mag_2.CLK.t8 VSS 0.0446f
C1704 CLK_div_3_mag_2.CLK.n12 VSS 0.0789f
C1705 CLK_div_3_mag_2.CLK.t13 VSS 0.0294f
C1706 CLK_div_3_mag_2.CLK.t14 VSS 0.0446f
C1707 CLK_div_3_mag_2.CLK.n13 VSS 0.0789f
C1708 CLK_div_3_mag_2.CLK.n14 VSS 1.18f
C1709 CLK_div_3_mag_2.CLK.n15 VSS 0.0501f
C1710 CLK_div_3_mag_2.CLK.n16 VSS 0.015f
C1711 CLK_div_3_mag_2.CLK.n17 VSS 0.173f
C1712 VDD.t99 VSS 0.00681f
C1713 VDD.t400 VSS 0.0028f
C1714 VDD.n0 VSS 0.0028f
C1715 VDD.n1 VSS 0.00611f
C1716 VDD.n2 VSS 0.022f
C1717 VDD.t359 VSS 0.00681f
C1718 VDD.n3 VSS 0.0269f
C1719 VDD.t222 VSS 0.0068f
C1720 VDD.t129 VSS 0.0068f
C1721 VDD.t225 VSS 0.0822f
C1722 VDD.n4 VSS 0.00681f
C1723 VDD.t61 VSS 0.0028f
C1724 VDD.n5 VSS 0.0028f
C1725 VDD.n6 VSS 0.00611f
C1726 VDD.n7 VSS 0.00681f
C1727 VDD.n8 VSS 0.0398f
C1728 VDD.t288 VSS 0.082f
C1729 VDD.n9 VSS 0.00681f
C1730 VDD.t441 VSS 0.00443f
C1731 VDD.t287 VSS 0.00584f
C1732 VDD.n10 VSS 0.0115f
C1733 VDD.t437 VSS 0.00443f
C1734 VDD.t295 VSS 0.00584f
C1735 VDD.n11 VSS 0.0114f
C1736 VDD.n12 VSS 0.0104f
C1737 VDD.n13 VSS 0.0434f
C1738 VDD.n14 VSS 0.0317f
C1739 VDD.t23 VSS 0.0028f
C1740 VDD.n15 VSS 0.0028f
C1741 VDD.n16 VSS 0.00611f
C1742 VDD.n17 VSS 0.0388f
C1743 VDD.n18 VSS 0.0211f
C1744 VDD.n19 VSS 0.0422f
C1745 VDD.t22 VSS 0.0463f
C1746 VDD.t146 VSS 0.1f
C1747 VDD.t344 VSS 0.0822f
C1748 VDD.t190 VSS 0.1f
C1749 VDD.t60 VSS 0.0463f
C1750 VDD.n20 VSS 0.0422f
C1751 VDD.n21 VSS 0.0211f
C1752 VDD.n22 VSS 0.0388f
C1753 VDD.n23 VSS 0.0396f
C1754 VDD.t27 VSS 0.0068f
C1755 VDD.n24 VSS 0.00681f
C1756 VDD.n25 VSS 0.0313f
C1757 VDD.n26 VSS 0.0337f
C1758 VDD.n27 VSS 0.0236f
C1759 VDD.n28 VSS 0.0422f
C1760 VDD.t26 VSS 0.0897f
C1761 VDD.t50 VSS 0.0822f
C1762 VDD.t128 VSS 0.0884f
C1763 VDD.n29 VSS 0.0422f
C1764 VDD.n30 VSS 0.0236f
C1765 VDD.n31 VSS 0.063f
C1766 VDD.n32 VSS 0.0991f
C1767 VDD.t24 VSS 0.364f
C1768 VDD.n33 VSS 0.205f
C1769 VDD.t19 VSS 0.0682f
C1770 VDD.n34 VSS 0.00697f
C1771 VDD.t330 VSS 0.00681f
C1772 VDD.t25 VSS 0.0028f
C1773 VDD.n35 VSS 0.0028f
C1774 VDD.n36 VSS 0.00611f
C1775 VDD.n37 VSS 0.151f
C1776 VDD.t10 VSS 0.0163f
C1777 VDD.n38 VSS 0.00681f
C1778 VDD.t329 VSS 0.174f
C1779 VDD.t9 VSS 0.153f
C1780 VDD.t7 VSS 0.0744f
C1781 VDD.n39 VSS 0.136f
C1782 VDD.n40 VSS 0.122f
C1783 VDD.t228 VSS 0.0068f
C1784 VDD.t8 VSS 0.00677f
C1785 VDD.n41 VSS 0.00681f
C1786 VDD.n42 VSS 0.0068f
C1787 VDD.n43 VSS 0.0223f
C1788 VDD.t28 VSS 0.0068f
C1789 VDD.n44 VSS 0.0244f
C1790 VDD.n45 VSS 0.0221f
C1791 VDD.n46 VSS 0.0216f
C1792 VDD.n47 VSS 0.0249f
C1793 VDD.n48 VSS 0.0352f
C1794 VDD.n49 VSS 0.0374f
C1795 VDD.n50 VSS 0.02f
C1796 VDD.n51 VSS 0.0281f
C1797 VDD.n52 VSS 0.0305f
C1798 VDD.n53 VSS 0.038f
C1799 VDD.n54 VSS 0.016f
C1800 VDD.n55 VSS 0.0369f
C1801 VDD.n56 VSS 0.0292f
C1802 VDD.n57 VSS 0.00681f
C1803 VDD.n58 VSS 0.0282f
C1804 VDD.n59 VSS 0.0176f
C1805 VDD.n60 VSS 0.0568f
C1806 VDD.n61 VSS 0.0738f
C1807 VDD.n62 VSS 0.108f
C1808 VDD.t187 VSS 0.0836f
C1809 VDD.t221 VSS 0.0836f
C1810 VDD.n63 VSS 0.0479f
C1811 VDD.n64 VSS 0.0302f
C1812 VDD.n65 VSS 0.00703f
C1813 VDD.n66 VSS 0.0322f
C1814 VDD.n67 VSS 0.0386f
C1815 VDD.t121 VSS 0.0898f
C1816 VDD.n68 VSS 0.0068f
C1817 VDD.t79 VSS 0.00681f
C1818 VDD.n69 VSS 0.0068f
C1819 VDD.n70 VSS 0.0337f
C1820 VDD.t397 VSS 0.0886f
C1821 VDD.n71 VSS 0.0068f
C1822 VDD.n72 VSS 0.0068f
C1823 VDD.t404 VSS 0.0886f
C1824 VDD.n73 VSS 0.0422f
C1825 VDD.t428 VSS 0.00681f
C1826 VDD.n74 VSS 0.0068f
C1827 VDD.t427 VSS 0.082f
C1828 VDD.t331 VSS 0.0898f
C1829 VDD.n75 VSS 0.0422f
C1830 VDD.t125 VSS 0.00681f
C1831 VDD.t77 VSS 0.0028f
C1832 VDD.n76 VSS 0.0028f
C1833 VDD.n77 VSS 0.00611f
C1834 VDD.t124 VSS 0.082f
C1835 VDD.t76 VSS 0.1f
C1836 VDD.t70 VSS 0.0465f
C1837 VDD.n78 VSS 0.0422f
C1838 VDD.t224 VSS 0.00681f
C1839 VDD.t408 VSS 0.0028f
C1840 VDD.n79 VSS 0.0028f
C1841 VDD.n80 VSS 0.00611f
C1842 VDD.t223 VSS 0.082f
C1843 VDD.t407 VSS 0.1f
C1844 VDD.t356 VSS 0.0465f
C1845 VDD.t267 VSS 0.0818f
C1846 VDD.n81 VSS 0.0422f
C1847 VDD.t268 VSS 0.00729f
C1848 VDD.n82 VSS 0.0524f
C1849 VDD.n83 VSS 0.0387f
C1850 VDD.n84 VSS 0.0398f
C1851 VDD.n85 VSS 0.0211f
C1852 VDD.n86 VSS 0.0387f
C1853 VDD.n87 VSS 0.0397f
C1854 VDD.n88 VSS 0.0235f
C1855 VDD.n89 VSS 0.0337f
C1856 VDD.n90 VSS 0.0313f
C1857 VDD.n91 VSS 0.0235f
C1858 VDD.n92 VSS 0.0641f
C1859 VDD.n93 VSS 0.0729f
C1860 VDD.t338 VSS 0.00681f
C1861 VDD.n94 VSS 0.0313f
C1862 VDD.n95 VSS 0.0235f
C1863 VDD.n96 VSS 0.0422f
C1864 VDD.t337 VSS 0.082f
C1865 VDD.t334 VSS 0.0898f
C1866 VDD.t78 VSS 0.082f
C1867 VDD.n97 VSS 0.0422f
C1868 VDD.n98 VSS 0.0235f
C1869 VDD.n99 VSS 0.0313f
C1870 VDD.n100 VSS 0.0337f
C1871 VDD.t363 VSS 0.00681f
C1872 VDD.n101 VSS 0.0297f
C1873 VDD.n102 VSS 0.0235f
C1874 VDD.n103 VSS 0.0422f
C1875 VDD.t362 VSS 0.082f
C1876 VDD.t399 VSS 0.1f
C1877 VDD.t90 VSS 0.0465f
C1878 VDD.t98 VSS 0.0463f
C1879 VDD.n104 VSS 0.0422f
C1880 VDD.n105 VSS 0.0156f
C1881 VDD.n106 VSS 0.053f
C1882 VDD.n107 VSS 0.0307f
C1883 VDD.t85 VSS 0.0633f
C1884 VDD.n108 VSS 0.0563f
C1885 VDD.n109 VSS 0.0427f
C1886 VDD.n110 VSS 0.0068f
C1887 VDD.t95 VSS 0.0886f
C1888 VDD.n111 VSS 0.0422f
C1889 VDD.t230 VSS 0.00681f
C1890 VDD.n112 VSS 0.0068f
C1891 VDD.t229 VSS 0.082f
C1892 VDD.t213 VSS 0.0898f
C1893 VDD.n113 VSS 0.0422f
C1894 VDD.t166 VSS 0.00681f
C1895 VDD.t415 VSS 0.0028f
C1896 VDD.n114 VSS 0.0028f
C1897 VDD.n115 VSS 0.00611f
C1898 VDD.t165 VSS 0.082f
C1899 VDD.t414 VSS 0.1f
C1900 VDD.t53 VSS 0.0465f
C1901 VDD.n116 VSS 0.0422f
C1902 VDD.t299 VSS 0.00681f
C1903 VDD.t101 VSS 0.0028f
C1904 VDD.n117 VSS 0.0028f
C1905 VDD.n118 VSS 0.00611f
C1906 VDD.t298 VSS 0.082f
C1907 VDD.t100 VSS 0.1f
C1908 VDD.t87 VSS 0.0465f
C1909 VDD.t282 VSS 0.0818f
C1910 VDD.n119 VSS 0.0422f
C1911 VDD.t283 VSS 0.00636f
C1912 VDD.t266 VSS 0.00584f
C1913 VDD.t450 VSS 0.00443f
C1914 VDD.n120 VSS 0.0114f
C1915 VDD.n121 VSS 0.064f
C1916 VDD.n122 VSS 0.0836f
C1917 VDD.n123 VSS 0.00149f
C1918 VDD.t445 VSS 0.00441f
C1919 VDD.n124 VSS 0.00598f
C1920 VDD.t281 VSS 0.00567f
C1921 VDD.n125 VSS 0.0056f
C1922 VDD.n126 VSS 5.65e-20
C1923 VDD.n127 VSS 0.00176f
C1924 VDD.n128 VSS 8.1e-19
C1925 VDD.n129 VSS 6.73e-19
C1926 VDD.n130 VSS 0.00506f
C1927 VDD.n131 VSS 0.0159f
C1928 VDD.n132 VSS 0.0388f
C1929 VDD.n133 VSS 0.0387f
C1930 VDD.n134 VSS 0.0398f
C1931 VDD.n135 VSS 0.0211f
C1932 VDD.n136 VSS 0.0387f
C1933 VDD.n137 VSS 0.0397f
C1934 VDD.n138 VSS 0.0235f
C1935 VDD.n139 VSS 0.0337f
C1936 VDD.n140 VSS 0.0313f
C1937 VDD.n141 VSS 0.0235f
C1938 VDD.n142 VSS 0.0588f
C1939 VDD.n143 VSS 0.0327f
C1940 VDD.n144 VSS 0.00677f
C1941 VDD.n145 VSS 0.00678f
C1942 VDD.n146 VSS 0.0365f
C1943 VDD.t278 VSS 0.047f
C1944 VDD.t32 VSS 0.0585f
C1945 VDD.n147 VSS 0.0358f
C1946 VDD.n148 VSS 0.0427f
C1947 VDD.n149 VSS 0.00681f
C1948 VDD.t361 VSS 0.00678f
C1949 VDD.n150 VSS 0.00678f
C1950 VDD.t33 VSS 0.0028f
C1951 VDD.n151 VSS 0.0028f
C1952 VDD.n152 VSS 0.00611f
C1953 VDD.t160 VSS 0.0217f
C1954 VDD.n153 VSS 0.0905f
C1955 VDD.n154 VSS 0.0427f
C1956 VDD.n155 VSS 0.00681f
C1957 VDD.t413 VSS 0.00678f
C1958 VDD.n156 VSS 0.0315f
C1959 VDD.n157 VSS 0.0334f
C1960 VDD.n158 VSS 0.00678f
C1961 VDD.t161 VSS 0.0068f
C1962 VDD.t120 VSS 0.00678f
C1963 VDD.n159 VSS 0.00681f
C1964 VDD.t103 VSS 0.0028f
C1965 VDD.n160 VSS 0.0028f
C1966 VDD.n161 VSS 0.00608f
C1967 VDD.n162 VSS 0.0256f
C1968 VDD.n163 VSS 0.0221f
C1969 VDD.t136 VSS 0.0068f
C1970 VDD.n164 VSS 0.0288f
C1971 VDD.n165 VSS 0.00681f
C1972 VDD.t403 VSS 0.00678f
C1973 VDD.t150 VSS 0.0068f
C1974 VDD.t84 VSS 0.0103f
C1975 VDD.t140 VSS 0.047f
C1976 VDD.n166 VSS 0.0358f
C1977 VDD.t149 VSS 0.0569f
C1978 VDD.t83 VSS 0.0937f
C1979 VDD.n167 VSS 0.0964f
C1980 VDD.n168 VSS 0.00677f
C1981 VDD.t202 VSS 0.214f
C1982 VDD.n169 VSS 0.0819f
C1983 VDD.n170 VSS 0.00695f
C1984 VDD.n171 VSS 0.0369f
C1985 VDD.n172 VSS 0.0872f
C1986 VDD.n173 VSS 0.0502f
C1987 VDD.n174 VSS 0.0205f
C1988 VDD.n175 VSS 0.0256f
C1989 VDD.t205 VSS 0.0028f
C1990 VDD.n176 VSS 0.0028f
C1991 VDD.n177 VSS 0.00607f
C1992 VDD.n178 VSS 0.00328f
C1993 VDD.n179 VSS 0.0265f
C1994 VDD.t118 VSS 0.0163f
C1995 VDD.n180 VSS 0.00677f
C1996 VDD.t241 VSS 0.00856f
C1997 VDD.n181 VSS 0.0238f
C1998 VDD.t313 VSS 0.00677f
C1999 VDD.n182 VSS 0.0068f
C2000 VDD.n183 VSS 0.00677f
C2001 VDD.n184 VSS 0.0112f
C2002 VDD.t175 VSS 0.00681f
C2003 VDD.n185 VSS 0.0252f
C2004 VDD.t394 VSS 0.0651f
C2005 VDD.n186 VSS 0.0203f
C2006 VDD.t240 VSS 0.00193f
C2007 VDD.n187 VSS 0.0313f
C2008 VDD.t312 VSS 0.13f
C2009 VDD.t375 VSS 0.13f
C2010 VDD.t303 VSS 0.0329f
C2011 VDD.n188 VSS 0.019f
C2012 VDD.t325 VSS 0.0941f
C2013 VDD.t326 VSS 0.00677f
C2014 VDD.t249 VSS 0.0068f
C2015 VDD.t309 VSS 0.0822f
C2016 VDD.n189 VSS 0.00681f
C2017 VDD.t57 VSS 0.0028f
C2018 VDD.n190 VSS 0.0028f
C2019 VDD.n191 VSS 0.00611f
C2020 VDD.n192 VSS 0.00681f
C2021 VDD.n193 VSS 0.0398f
C2022 VDD.t270 VSS 0.082f
C2023 VDD.n194 VSS 6.73e-19
C2024 VDD.t439 VSS 0.00443f
C2025 VDD.t291 VSS 0.00584f
C2026 VDD.n195 VSS 0.0114f
C2027 VDD.n196 VSS 0.0758f
C2028 VDD.n197 VSS 0.0748f
C2029 VDD.t449 VSS 0.00443f
C2030 VDD.t269 VSS 0.00572f
C2031 VDD.n198 VSS 0.00544f
C2032 VDD.n199 VSS 0.00607f
C2033 VDD.n200 VSS 9.61e-19
C2034 VDD.n201 VSS 0.00508f
C2035 VDD.n202 VSS 0.00636f
C2036 VDD.n203 VSS 0.0159f
C2037 VDD.t210 VSS 0.0028f
C2038 VDD.n204 VSS 0.0028f
C2039 VDD.n205 VSS 0.00611f
C2040 VDD.n206 VSS 0.0388f
C2041 VDD.n207 VSS 0.0389f
C2042 VDD.n208 VSS 0.0422f
C2043 VDD.t209 VSS 0.0463f
C2044 VDD.t255 VSS 0.1f
C2045 VDD.t143 VSS 0.0822f
C2046 VDD.t306 VSS 0.1f
C2047 VDD.t56 VSS 0.0463f
C2048 VDD.n209 VSS 0.0422f
C2049 VDD.n210 VSS 0.0211f
C2050 VDD.n211 VSS 0.0388f
C2051 VDD.n212 VSS 0.0396f
C2052 VDD.t3 VSS 0.0068f
C2053 VDD.n213 VSS 0.00681f
C2054 VDD.n214 VSS 0.0313f
C2055 VDD.n215 VSS 0.0337f
C2056 VDD.n216 VSS 0.0236f
C2057 VDD.n217 VSS 0.0422f
C2058 VDD.t2 VSS 0.0897f
C2059 VDD.t4 VSS 0.0822f
C2060 VDD.t248 VSS 0.0884f
C2061 VDD.n218 VSS 0.0422f
C2062 VDD.n219 VSS 0.0236f
C2063 VDD.n220 VSS 0.0602f
C2064 VDD.n221 VSS 0.00677f
C2065 VDD.n222 VSS 0.00681f
C2066 VDD.n223 VSS 0.03f
C2067 VDD.t206 VSS 0.0602f
C2068 VDD.n224 VSS 0.0157f
C2069 VDD.n225 VSS 0.00681f
C2070 VDD.t212 VSS 0.0028f
C2071 VDD.n226 VSS 0.0028f
C2072 VDD.n227 VSS 0.00611f
C2073 VDD.n228 VSS 0.0068f
C2074 VDD.t180 VSS 0.00677f
C2075 VDD.n229 VSS 0.0068f
C2076 VDD.t382 VSS 0.0886f
C2077 VDD.n230 VSS 0.0422f
C2078 VDD.t239 VSS 0.00681f
C2079 VDD.n231 VSS 0.0068f
C2080 VDD.t238 VSS 0.082f
C2081 VDD.t317 VSS 0.0898f
C2082 VDD.n232 VSS 0.0422f
C2083 VDD.t324 VSS 0.00681f
C2084 VDD.t391 VSS 0.0028f
C2085 VDD.n233 VSS 0.0028f
C2086 VDD.n234 VSS 0.00611f
C2087 VDD.t323 VSS 0.082f
C2088 VDD.t390 VSS 0.1f
C2089 VDD.t65 VSS 0.0465f
C2090 VDD.n235 VSS 0.0422f
C2091 VDD.t117 VSS 0.00681f
C2092 VDD.t379 VSS 0.0028f
C2093 VDD.n236 VSS 0.0028f
C2094 VDD.n237 VSS 0.00611f
C2095 VDD.t116 VSS 0.082f
C2096 VDD.t378 VSS 0.1f
C2097 VDD.t181 VSS 0.0465f
C2098 VDD.t264 VSS 0.0818f
C2099 VDD.n238 VSS 0.0422f
C2100 VDD.t265 VSS 0.00636f
C2101 VDD.n239 VSS 0.00176f
C2102 VDD.t263 VSS 0.00567f
C2103 VDD.n240 VSS 0.0056f
C2104 VDD.t284 VSS 0.00584f
C2105 VDD.t442 VSS 0.00443f
C2106 VDD.n241 VSS 0.0114f
C2107 VDD.n242 VSS 0.064f
C2108 VDD.n243 VSS 0.0836f
C2109 VDD.n244 VSS 5.65e-20
C2110 VDD.n245 VSS 0.00149f
C2111 VDD.t451 VSS 0.00441f
C2112 VDD.n246 VSS 0.00598f
C2113 VDD.n247 VSS 8.1e-19
C2114 VDD.n248 VSS 6.73e-19
C2115 VDD.n249 VSS 0.00506f
C2116 VDD.n250 VSS 0.0159f
C2117 VDD.n251 VSS 0.0388f
C2118 VDD.n252 VSS 0.0387f
C2119 VDD.n253 VSS 0.0398f
C2120 VDD.n254 VSS 0.0211f
C2121 VDD.n255 VSS 0.0387f
C2122 VDD.n256 VSS 0.0397f
C2123 VDD.n257 VSS 0.0235f
C2124 VDD.n258 VSS 0.0337f
C2125 VDD.n259 VSS 0.0313f
C2126 VDD.n260 VSS 0.0235f
C2127 VDD.n261 VSS 0.0777f
C2128 VDD.n262 VSS 0.0238f
C2129 VDD.t381 VSS 0.00681f
C2130 VDD.n263 VSS 0.0266f
C2131 VDD.t184 VSS 0.037f
C2132 VDD.t370 VSS 0.0028f
C2133 VDD.n264 VSS 0.0028f
C2134 VDD.n265 VSS 0.00611f
C2135 VDD.t168 VSS 0.00681f
C2136 VDD.n266 VSS 0.0068f
C2137 VDD.n267 VSS 0.0211f
C2138 VDD.t37 VSS 0.0715f
C2139 VDD.n268 VSS 0.0068f
C2140 VDD.t41 VSS 0.00681f
C2141 VDD.n269 VSS 0.0068f
C2142 VDD.n270 VSS 0.0068f
C2143 VDD.t13 VSS 0.0886f
C2144 VDD.n271 VSS 0.0422f
C2145 VDD.t374 VSS 0.00681f
C2146 VDD.n272 VSS 0.0068f
C2147 VDD.t373 VSS 0.082f
C2148 VDD.t34 VSS 0.0898f
C2149 VDD.n273 VSS 0.0422f
C2150 VDD.t348 VSS 0.00681f
C2151 VDD.t355 VSS 0.0028f
C2152 VDD.n274 VSS 0.0028f
C2153 VDD.n275 VSS 0.00611f
C2154 VDD.t347 VSS 0.082f
C2155 VDD.t354 VSS 0.1f
C2156 VDD.t58 VSS 0.0465f
C2157 VDD.n276 VSS 0.0422f
C2158 VDD.t12 VSS 0.00681f
C2159 VDD.t18 VSS 0.0028f
C2160 VDD.n277 VSS 0.0028f
C2161 VDD.n278 VSS 0.00611f
C2162 VDD.t11 VSS 0.082f
C2163 VDD.t17 VSS 0.1f
C2164 VDD.t169 VSS 0.0465f
C2165 VDD.t285 VSS 0.0818f
C2166 VDD.n279 VSS 0.0422f
C2167 VDD.t286 VSS 0.00729f
C2168 VDD.n280 VSS 0.0524f
C2169 VDD.n281 VSS 0.0387f
C2170 VDD.n282 VSS 0.0398f
C2171 VDD.n283 VSS 0.0211f
C2172 VDD.n284 VSS 0.0387f
C2173 VDD.n285 VSS 0.0397f
C2174 VDD.n286 VSS 0.0235f
C2175 VDD.n287 VSS 0.0337f
C2176 VDD.n288 VSS 0.0313f
C2177 VDD.n289 VSS 0.0235f
C2178 VDD.n290 VSS 0.0657f
C2179 VDD.n291 VSS 0.057f
C2180 VDD.t366 VSS 0.0715f
C2181 VDD.t40 VSS 0.0653f
C2182 VDD.n292 VSS 0.0364f
C2183 VDD.n293 VSS 0.0198f
C2184 VDD.n294 VSS 0.0238f
C2185 VDD.n295 VSS 0.0252f
C2186 VDD.t353 VSS 0.00681f
C2187 VDD.n296 VSS 0.00906f
C2188 VDD.n297 VSS 0.00647f
C2189 VDD.n298 VSS 0.0103f
C2190 VDD.n299 VSS 0.00968f
C2191 VDD.n300 VSS 0.00838f
C2192 VDD.t1 VSS 0.00644f
C2193 VDD.n301 VSS 0.00934f
C2194 VDD.n302 VSS 0.0113f
C2195 VDD.n303 VSS 0.0246f
C2196 VDD.n304 VSS 0.0937f
C2197 VDD.n305 VSS 0.0201f
C2198 VDD.n306 VSS 0.0198f
C2199 VDD.n307 VSS 0.0364f
C2200 VDD.t352 VSS 0.0653f
C2201 VDD.t349 VSS 0.0708f
C2202 VDD.t369 VSS 0.0797f
C2203 VDD.t167 VSS 0.0653f
C2204 VDD.n308 VSS 0.034f
C2205 VDD.n309 VSS 0.0198f
C2206 VDD.n310 VSS 0.0228f
C2207 VDD.n311 VSS 0.0204f
C2208 VDD.n312 VSS 0.0183f
C2209 VDD.n313 VSS 0.0364f
C2210 VDD.t380 VSS 0.0653f
C2211 VDD.t179 VSS 0.0948f
C2212 VDD.n314 VSS 0.0186f
C2213 VDD.n315 VSS 0.0304f
C2214 VDD.n316 VSS 0.0279f
C2215 VDD.n317 VSS 0.0111f
C2216 VDD.n318 VSS 0.00645f
C2217 VDD.n319 VSS 0.00958f
C2218 VDD.t237 VSS 0.00681f
C2219 VDD.t385 VSS 0.0715f
C2220 VDD.t236 VSS 0.0465f
C2221 VDD.n320 VSS 0.0187f
C2222 VDD.n321 VSS 0.011f
C2223 VDD.n322 VSS 0.00681f
C2224 VDD.n323 VSS 0.0247f
C2225 VDD.t393 VSS 0.00681f
C2226 VDD.t251 VSS 0.0068f
C2227 VDD.n324 VSS 0.0068f
C2228 VDD.n325 VSS 0.00854f
C2229 VDD.n326 VSS 0.014f
C2230 VDD.n327 VSS 0.0235f
C2231 VDD.t392 VSS 0.0326f
C2232 VDD.t250 VSS 0.13f
C2233 VDD.t320 VSS 0.13f
C2234 VDD.t112 VSS 0.0557f
C2235 VDD.n328 VSS -0.00162f
C2236 VDD.n329 VSS 0.0163f
C2237 VDD.t49 VSS 0.00681f
C2238 VDD.n330 VSS 5.01e-19
C2239 VDD.n331 VSS 0.0346f
C2240 VDD.n332 VSS 0.0332f
C2241 VDD.t388 VSS 0.0028f
C2242 VDD.n333 VSS 0.0028f
C2243 VDD.n334 VSS 0.00611f
C2244 VDD.t372 VSS 0.00681f
C2245 VDD.n335 VSS 0.00677f
C2246 VDD.t176 VSS 0.0603f
C2247 VDD.n336 VSS 0.0603f
C2248 VDD.t371 VSS 0.0911f
C2249 VDD.n337 VSS 0.079f
C2250 VDD.t173 VSS 0.00678f
C2251 VDD.n338 VSS 0.0162f
C2252 VDD.t172 VSS 0.0265f
C2253 VDD.t252 VSS 0.0829f
C2254 VDD.n339 VSS 0.0891f
C2255 VDD.n340 VSS 0.0323f
C2256 VDD.n341 VSS 0.026f
C2257 VDD.n342 VSS 0.0337f
C2258 VDD.n343 VSS 0.0118f
C2259 VDD.n344 VSS 0.0261f
C2260 VDD.n345 VSS 0.00523f
C2261 VDD.n346 VSS 0.00936f
C2262 VDD.n347 VSS 0.0384f
C2263 VDD.t387 VSS 0.0264f
C2264 VDD.t300 VSS 0.154f
C2265 VDD.t48 VSS 0.132f
C2266 VDD.n348 VSS 0.0203f
C2267 VDD.t242 VSS 0.00226f
C2268 VDD.n349 VSS 0.0313f
C2269 VDD.n350 VSS 0.0232f
C2270 VDD.n351 VSS 0.0343f
C2271 VDD.n352 VSS 0.0288f
C2272 VDD.n353 VSS 0.0248f
C2273 VDD.n354 VSS 0.00666f
C2274 VDD.n355 VSS 0.00616f
C2275 VDD.n356 VSS 0.0112f
C2276 VDD.n357 VSS 0.019f
C2277 VDD.t199 VSS 0.0329f
C2278 VDD.t314 VSS 0.139f
C2279 VDD.n358 VSS 0.0381f
C2280 VDD.n359 VSS 0.0525f
C2281 VDD.n360 VSS 0.0155f
C2282 VDD.n361 VSS 0.023f
C2283 VDD.n362 VSS 0.00716f
C2284 VDD.n363 VSS 0.00621f
C2285 VDD.n364 VSS 0.0212f
C2286 VDD.n365 VSS 0.053f
C2287 VDD.n366 VSS 0.022f
C2288 VDD.n367 VSS 0.0297f
C2289 VDD.n368 VSS 0.0236f
C2290 VDD.n369 VSS 0.00681f
C2291 VDD.t420 VSS 0.0068f
C2292 VDD.n370 VSS 0.0337f
C2293 VDD.n371 VSS 0.0313f
C2294 VDD.n372 VSS 0.0236f
C2295 VDD.t234 VSS 0.0884f
C2296 VDD.n373 VSS 0.00681f
C2297 VDD.t433 VSS 0.0068f
C2298 VDD.n374 VSS 0.0337f
C2299 VDD.n375 VSS 0.0313f
C2300 VDD.t235 VSS 0.0068f
C2301 VDD.t111 VSS 0.0068f
C2302 VDD.t416 VSS 0.0822f
C2303 VDD.n376 VSS 0.00681f
C2304 VDD.t69 VSS 0.0028f
C2305 VDD.n377 VSS 0.0028f
C2306 VDD.n378 VSS 0.00611f
C2307 VDD.n379 VSS 0.00681f
C2308 VDD.n380 VSS 0.0398f
C2309 VDD.t292 VSS 0.082f
C2310 VDD.n381 VSS 0.00729f
C2311 VDD.t198 VSS 0.0028f
C2312 VDD.n382 VSS 0.0028f
C2313 VDD.n383 VSS 0.00611f
C2314 VDD.n384 VSS 0.0388f
C2315 VDD.n385 VSS 0.0524f
C2316 VDD.n386 VSS 0.0422f
C2317 VDD.t197 VSS 0.0463f
C2318 VDD.t107 VSS 0.1f
C2319 VDD.t29 VSS 0.0822f
C2320 VDD.t424 VSS 0.1f
C2321 VDD.t68 VSS 0.0463f
C2322 VDD.n387 VSS 0.0422f
C2323 VDD.n388 VSS 0.0211f
C2324 VDD.n389 VSS 0.0388f
C2325 VDD.n390 VSS 0.0396f
C2326 VDD.t435 VSS 0.0068f
C2327 VDD.n391 VSS 0.00681f
C2328 VDD.n392 VSS 0.0313f
C2329 VDD.n393 VSS 0.0337f
C2330 VDD.n394 VSS 0.0236f
C2331 VDD.n395 VSS 0.0422f
C2332 VDD.t434 VSS 0.0897f
C2333 VDD.t429 VSS 0.0822f
C2334 VDD.t110 VSS 0.0884f
C2335 VDD.n396 VSS 0.0422f
C2336 VDD.n397 VSS 0.0236f
C2337 VDD.n398 VSS 0.064f
C2338 VDD.n399 VSS 0.0728f
C2339 VDD.n400 VSS 0.0236f
C2340 VDD.n401 VSS 0.0422f
C2341 VDD.t73 VSS 0.0822f
C2342 VDD.t432 VSS 0.0897f
C2343 VDD.n402 VSS 0.0422f
C2344 VDD.t421 VSS 0.0822f
C2345 VDD.t419 VSS 0.0897f
C2346 VDD.n403 VSS 0.0422f
C2347 VDD.t113 VSS 0.0822f
C2348 VDD.t258 VSS 0.1f
C2349 VDD.t211 VSS 0.0463f
C2350 VDD.n404 VSS 0.0422f
C2351 VDD.t245 VSS 0.0467f
C2352 VDD.n405 VSS 0.0632f
C2353 VDD.n406 VSS 0.0213f
C2354 VDD.n407 VSS 0.0479f
C2355 VDD.n408 VSS 0.0404f
C2356 VDD.n409 VSS 0.0263f
C2357 VDD.n410 VSS 0.044f
C2358 VDD.t409 VSS 0.122f
C2359 VDD.t0 VSS 0.101f
C2360 VDD.t174 VSS 0.0326f
C2361 VDD.n411 VSS 0.0187f
C2362 VDD.n412 VSS 0.011f
C2363 VDD.n413 VSS 0.00649f
C2364 VDD.n414 VSS 0.00687f
C2365 VDD.n415 VSS 0.025f
C2366 VDD.n416 VSS 0.0296f
C2367 VDD.n417 VSS 0.0351f
C2368 VDD.n418 VSS 0.014f
C2369 VDD.n419 VSS 5.23e-19
C2370 VDD.n420 VSS 0.0352f
C2371 VDD.n421 VSS 0.0339f
C2372 VDD.n422 VSS 0.00538f
C2373 VDD.n423 VSS 0.0446f
C2374 VDD.n424 VSS 0.0769f
C2375 VDD.t364 VSS 0.163f
C2376 VDD.t16 VSS 0.0632f
C2377 VDD.n425 VSS 0.103f
C2378 VDD.t365 VSS 0.00683f
C2379 VDD.n426 VSS 0.0454f
C2380 VDD.n427 VSS 0.0546f
C2381 VDD.t196 VSS 0.0068f
C2382 VDD.t157 VSS 0.0822f
C2383 VDD.n428 VSS 0.00681f
C2384 VDD.t64 VSS 0.0028f
C2385 VDD.n429 VSS 0.0028f
C2386 VDD.n430 VSS 0.00611f
C2387 VDD.n431 VSS 0.00681f
C2388 VDD.n432 VSS 0.0398f
C2389 VDD.t274 VSS 0.082f
C2390 VDD.n433 VSS 0.00681f
C2391 VDD.t447 VSS 0.00443f
C2392 VDD.t273 VSS 0.00584f
C2393 VDD.n434 VSS 0.0115f
C2394 VDD.n435 VSS 0.00866f
C2395 VDD.t444 VSS 0.00443f
C2396 VDD.t277 VSS 0.00584f
C2397 VDD.n436 VSS 0.0115f
C2398 VDD.n437 VSS 0.00778f
C2399 VDD.n438 VSS 0.0469f
C2400 VDD.n439 VSS 0.0318f
C2401 VDD.t127 VSS 0.0028f
C2402 VDD.n440 VSS 0.0028f
C2403 VDD.n441 VSS 0.00611f
C2404 VDD.n442 VSS 0.0388f
C2405 VDD.n443 VSS 0.0211f
C2406 VDD.n444 VSS 0.0422f
C2407 VDD.t126 VSS 0.0463f
C2408 VDD.t130 VSS 0.1f
C2409 VDD.t339 VSS 0.0822f
C2410 VDD.t42 VSS 0.1f
C2411 VDD.t63 VSS 0.0463f
C2412 VDD.n445 VSS 0.0422f
C2413 VDD.n446 VSS 0.0211f
C2414 VDD.n447 VSS 0.0388f
C2415 VDD.n448 VSS 0.0396f
C2416 VDD.t134 VSS 0.0068f
C2417 VDD.n449 VSS 0.00681f
C2418 VDD.n450 VSS 0.0313f
C2419 VDD.n451 VSS 0.0337f
C2420 VDD.n452 VSS 0.0236f
C2421 VDD.n453 VSS 0.0422f
C2422 VDD.t133 VSS 0.0897f
C2423 VDD.t231 VSS 0.0822f
C2424 VDD.t195 VSS 0.0884f
C2425 VDD.n454 VSS 0.0422f
C2426 VDD.n455 VSS 0.0236f
C2427 VDD.n456 VSS 0.031f
C2428 VDD.n457 VSS 0.0683f
C2429 VDD.n458 VSS 0.0168f
C2430 VDD.n459 VSS 0.0355f
C2431 VDD.n460 VSS 0.0178f
C2432 VDD.n461 VSS 0.0243f
C2433 VDD.n462 VSS 0.0248f
C2434 VDD.n463 VSS 0.00704f
C2435 VDD.n464 VSS 0.0905f
C2436 VDD.n465 VSS 0.051f
C2437 VDD.t45 VSS 0.0829f
C2438 VDD.t135 VSS 0.0793f
C2439 VDD.n466 VSS 0.0358f
C2440 VDD.n467 VSS 0.0505f
C2441 VDD.n468 VSS 0.0165f
C2442 VDD.n469 VSS 0.0316f
C2443 VDD.n470 VSS 0.0333f
C2444 VDD.n471 VSS 0.00114f
C2445 VDD.n472 VSS 0.029f
C2446 VDD.n473 VSS 0.0288f
C2447 VDD.n474 VSS 0.00124f
C2448 VDD.t154 VSS 0.0829f
C2449 VDD.t104 VSS 0.0677f
C2450 VDD.t360 VSS 0.0677f
C2451 VDD.t216 VSS 0.0677f
C2452 VDD.t412 VSS 0.0677f
C2453 VDD.t162 VSS 0.0491f
C2454 VDD.t402 VSS 0.0677f
C2455 VDD.t80 VSS 0.0384f
C2456 VDD.t102 VSS 0.0677f
C2457 VDD.t119 VSS 0.0671f
C2458 VDD.n475 VSS 0.0418f
C2459 VDD.n476 VSS 0.0349f
C2460 VDD.n477 VSS 0.0428f
C2461 VDD.t151 VSS 0.0567f
C2462 VDD.n478 VSS 0.0905f
C2463 VDD.n479 VSS 0.0505f
C2464 VDD.n480 VSS 0.0164f
C2465 VDD.n481 VSS 0.0258f
C2466 VDD.n482 VSS 0.0287f
C2467 VDD.n483 VSS 0.00695f
C2468 VDD.n484 VSS 0.0246f
C2469 VDD.n485 VSS 0.0246f
C2470 VDD.n486 VSS 0.0179f
C2471 VDD.n487 VSS 0.0905f
C2472 VDD.n488 VSS 0.0367f
C2473 VDD.n489 VSS 0.0577f
C2474 VDD.t137 VSS 0.0571f
C2475 VDD.n490 VSS 0.0733f
C2476 VDD.n491 VSS 0.0435f
C2477 VDD.n492 VSS 0.028f
C2478 VDD.n493 VSS 0.0117f
C2479 VDD.n494 VSS 0.00711f
C2480 VDD.n495 VSS 0.00778f
C2481 VDD.t86 VSS 0.00644f
C2482 VDD.n496 VSS 0.0104f
C2483 VDD.n497 VSS 0.00827f
C2484 CLK_div_3_mag_0.CLK.n0 VSS 0.453f
C2485 CLK_div_3_mag_0.CLK.n1 VSS 0.286f
C2486 CLK_div_3_mag_0.CLK.n2 VSS 0.0181f
C2487 CLK_div_3_mag_0.CLK.n3 VSS 0.0181f
C2488 CLK_div_3_mag_0.CLK.n4 VSS 0.123f
C2489 CLK_div_3_mag_0.CLK.n5 VSS 0.114f
C2490 CLK_div_3_mag_0.CLK.n6 VSS 0.0581f
C2491 CLK_div_3_mag_0.CLK.t1 VSS 0.0147f
C2492 CLK_div_3_mag_0.CLK.t0 VSS 0.0475f
C2493 CLK_div_3_mag_0.CLK.n7 VSS 0.176f
C2494 CLK_div_3_mag_0.CLK.t6 VSS 0.0292f
C2495 CLK_div_3_mag_0.CLK.t8 VSS 0.0443f
C2496 CLK_div_3_mag_0.CLK.n8 VSS 0.0783f
C2497 CLK_div_3_mag_0.CLK.t9 VSS 0.0292f
C2498 CLK_div_3_mag_0.CLK.t11 VSS 0.0443f
C2499 CLK_div_3_mag_0.CLK.n9 VSS 0.0784f
C2500 CLK_div_3_mag_0.CLK.t14 VSS 0.0229f
C2501 CLK_div_3_mag_0.CLK.t10 VSS 0.0411f
C2502 CLK_div_3_mag_0.CLK.n10 VSS 0.0782f
C2503 CLK_div_3_mag_0.CLK.n11 VSS 0.251f
C2504 CLK_div_3_mag_0.CLK.t15 VSS 0.0292f
C2505 CLK_div_3_mag_0.CLK.t2 VSS 0.0443f
C2506 CLK_div_3_mag_0.CLK.n12 VSS 0.0783f
C2507 CLK_div_3_mag_0.CLK.t3 VSS 0.0292f
C2508 CLK_div_3_mag_0.CLK.t5 VSS 0.0443f
C2509 CLK_div_3_mag_0.CLK.n13 VSS 0.0784f
C2510 CLK_div_3_mag_0.CLK.t7 VSS 0.0366f
C2511 CLK_div_3_mag_0.CLK.t12 VSS 0.00936f
C2512 CLK_div_3_mag_0.CLK.n14 VSS 0.0607f
C2513 CLK_div_3_mag_0.CLK.n15 VSS 0.584f
C2514 CLK_div_3_mag_0.CLK.n16 VSS 0.584f
C2515 CLK_div_3_mag_0.CLK.t4 VSS 0.00936f
C2516 CLK_div_3_mag_0.CLK.t13 VSS 0.0366f
C2517 CLK_div_3_mag_0.CLK.n17 VSS 0.0607f
C2518 RST.t11 VSS 0.0103f
C2519 RST.t9 VSS 0.00679f
C2520 RST.n0 VSS 0.0182f
C2521 RST.n1 VSS 0.00251f
C2522 RST.n2 VSS 0.00146f
C2523 RST.n3 VSS 9.36e-19
C2524 RST.n4 VSS 0.00316f
C2525 RST.n5 VSS 0.00137f
C2526 RST.n6 VSS 0.00521f
C2527 RST.n7 VSS 0.212f
C2528 RST.n8 VSS 0.00297f
C2529 RST.t3 VSS 0.0104f
C2530 RST.t2 VSS 0.0066f
C2531 RST.n9 VSS 0.0183f
C2532 RST.n10 VSS 0.00238f
C2533 RST.n11 VSS 0.00158f
C2534 RST.n12 VSS 8.39e-19
C2535 RST.n13 VSS 0.0386f
C2536 RST.n14 VSS 0.00106f
C2537 RST.n15 VSS 0.0032f
C2538 RST.t14 VSS 0.0103f
C2539 RST.t12 VSS 0.00679f
C2540 RST.n16 VSS 0.0182f
C2541 RST.n17 VSS 0.00238f
C2542 RST.n18 VSS 8.53e-19
C2543 RST.n19 VSS 0.0676f
C2544 RST.n20 VSS 0.349f
C2545 RST.n21 VSS 8.18e-19
C2546 RST.n22 VSS 0.00158f
C2547 RST.n23 VSS 0.00305f
C2548 RST.n24 VSS 0.00158f
C2549 RST.t13 VSS 0.0104f
C2550 RST.t10 VSS 0.00663f
C2551 RST.n25 VSS 0.0183f
C2552 RST.n26 VSS 0.00235f
C2553 RST.n27 VSS 8.39e-19
C2554 RST.n28 VSS 0.0979f
C2555 RST.n29 VSS 0.122f
C2556 RST.t5 VSS 0.00679f
C2557 RST.t8 VSS 0.0103f
C2558 RST.n30 VSS 0.0182f
C2559 RST.n31 VSS 0.00235f
C2560 RST.n32 VSS 8.54e-19
C2561 RST.n33 VSS 0.0542f
C2562 RST.n34 VSS 0.679f
C2563 RST.n35 VSS 0.312f
C2564 RST.n36 VSS 0.00305f
C2565 RST.n37 VSS 0.00158f
C2566 RST.t4 VSS 0.0104f
C2567 RST.t1 VSS 0.00663f
C2568 RST.n38 VSS 0.0183f
C2569 RST.n39 VSS 0.00235f
C2570 RST.n40 VSS 8.39e-19
C2571 RST.n41 VSS 0.0974f
C2572 RST.n42 VSS 0.122f
C2573 RST.n43 VSS 8.77e-19
C2574 RST.n44 VSS 0.00114f
C2575 RST.n45 VSS 0.00174f
C2576 RST.n46 VSS 0.00158f
C2577 RST.t15 VSS 0.00679f
C2578 RST.t0 VSS 0.0103f
C2579 RST.n47 VSS 0.0182f
C2580 RST.n48 VSS 0.00235f
C2581 RST.n49 VSS 8.39e-19
C2582 RST.n50 VSS 1.5e-19
C2583 RST.n51 VSS 1.2e-19
C2584 RST.n52 VSS 0.00191f
C2585 RST.n53 VSS 0.00171f
C2586 RST.n54 VSS 0.00491f
C2587 RST.n55 VSS 0.00152f
C2588 RST.n56 VSS 1.2e-19
C2589 RST.n57 VSS 0.206f
C2590 RST.n58 VSS 0.00503f
C2591 RST.n59 VSS 0.00145f
C2592 RST.n60 VSS 8.84e-19
C2593 RST.t7 VSS 0.0103f
C2594 RST.t6 VSS 0.00679f
C2595 RST.n61 VSS 0.0182f
C2596 RST.n62 VSS 0.00253f
C2597 RST.n63 VSS 0.00312f
C2598 RST.n64 VSS 0.00209f
C2599 RST.n65 VSS 0.00929f
C2600 RST.n66 VSS 0.00465f
C2601 RST.n67 VSS 0.354f
C2602 RST.n68 VSS 0.515f
C2603 RST.n69 VSS 0.0949f
C2604 RST.n70 VSS 0.0537f
C2605 CLK_div_3_mag_2.JK_FF_mag_1.K.n0 VSS 2.18f
C2606 CLK_div_3_mag_2.JK_FF_mag_1.K.n1 VSS 0.211f
C2607 CLK_div_3_mag_2.JK_FF_mag_1.K.t4 VSS 0.0734f
C2608 CLK_div_3_mag_2.JK_FF_mag_1.K.t5 VSS 0.057f
C2609 CLK_div_3_mag_2.JK_FF_mag_1.K.n2 VSS 0.146f
C2610 CLK_div_3_mag_2.JK_FF_mag_1.K.t8 VSS 0.0456f
C2611 CLK_div_3_mag_2.JK_FF_mag_1.K.t6 VSS 0.0571f
C2612 CLK_div_3_mag_2.JK_FF_mag_1.K.n3 VSS 0.147f
C2613 CLK_div_3_mag_2.JK_FF_mag_1.K.t3 VSS 0.0801f
C2614 CLK_div_3_mag_2.JK_FF_mag_1.K.t7 VSS 0.051f
C2615 CLK_div_3_mag_2.JK_FF_mag_1.K.n4 VSS 0.142f
C2616 CLK_div_3_mag_2.JK_FF_mag_1.K.n5 VSS 1.22f
C2617 CLK_div_3_mag_2.JK_FF_mag_1.K.t1 VSS 0.0356f
C2618 CLK_div_3_mag_2.JK_FF_mag_1.K.n6 VSS 0.0356f
C2619 CLK_div_3_mag_2.JK_FF_mag_1.K.n7 VSS 0.084f
.ends

