* NGSPICE file created from AND_2_In_Layout_flat.ext - technology: gf180mcuC

.subckt AND_2_Input_PEX VDD A OUT B VSS
X0 a_24_68# A.t0 a_168_68# VSS.t6 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X1 a_168_68# A.t1 a_24_68# VSS.t5 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X2 a_168_68# A.t2 VDD.t4 VDD.t3 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X3 a_24_68# B.t0 VSS.t4 VSS.t3 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X4 VDD B.t1 a_168_68# VDD.t0 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X5 VSS B.t2 a_24_68# VSS.t0 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X6 OUT a_168_68# VDD.t6 VDD.t5 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X7 OUT a_168_68# VSS.t8 VSS.t7 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
R0 A.n0 A.t2 33.763
R1 A.n1 A.n0 17.2076
R2 A.n1 A.t1 15.8587
R3 A.n0 A.t0 13.9487
R4 A A.n1 4.06507
R5 VSS.t0 VSS.n26 389.159
R6 VSS.n23 VSS.t6 241.91
R7 VSS.n27 VSS.t0 105.178
R8 VSS.n17 VSS.t5 94.6607
R9 VSS.n3 VSS.t7 42.0717
R10 VSS.n14 VSS.t3 42.0717
R11 VSS.n16 VSS.n15 9.13939
R12 VSS.n28 VSS.n16 9.13939
R13 VSS.n6 VSS.t8 7.04085
R14 VSS VSS.n16 5.2005
R15 VSS VSS.n16 5.2005
R16 VSS.n2 VSS.n1 3.76485
R17 VSS.n1 VSS.t4 3.2765
R18 VSS.n1 VSS.n0 3.2765
R19 VSS.n4 VSS.n3 2.6005
R20 VSS.n9 VSS.n8 2.6005
R21 VSS.n8 VSS.n7 2.6005
R22 VSS.n12 VSS.n11 2.6005
R23 VSS.n11 VSS.n10 2.6005
R24 VSS.n15 VSS.n13 2.6005
R25 VSS.n15 VSS.n14 2.6005
R26 VSS.n26 VSS.n16 2.6005
R27 VSS.n29 VSS.n28 2.6005
R28 VSS.n28 VSS.n27 2.6005
R29 VSS.n25 VSS.n24 2.6005
R30 VSS.n24 VSS.n23 2.6005
R31 VSS.n22 VSS.n21 2.6005
R32 VSS.n21 VSS.n20 2.6005
R33 VSS.n18 VSS.n17 2.6005
R34 VSS.n5 VSS.n4 1.64943
R35 VSS.n19 VSS.n18 1.64943
R36 VSS.n22 VSS.n19 0.559135
R37 VSS.n6 VSS.n5 0.541457
R38 VSS.n12 VSS.n9 0.0760357
R39 VSS.n13 VSS.n12 0.0760357
R40 VSS VSS.n29 0.0760357
R41 VSS.n29 VSS.n25 0.0760357
R42 VSS.n25 VSS.n22 0.0760357
R43 VSS.n13 VSS.n2 0.0712143
R44 VSS.n9 VSS.n6 0.0181786
R45 VSS VSS.n2 0.00532143
R46 VDD.t0 VDD.n5 179.732
R47 VDD.n3 VDD.t5 58.0931
R48 VDD.n8 VDD.t3 56.5038
R49 VDD.n6 VDD.n4 8.2255
R50 VDD.n12 VDD.n6 8.2255
R51 VDD VDD.n6 6.3005
R52 VDD VDD.n6 6.3005
R53 VDD.n7 VDD.t4 4.7492
R54 VDD.n5 VDD.n4 3.1505
R55 VDD.n6 VDD.t0 3.1505
R56 VDD.n13 VDD.n12 3.1505
R57 VDD.n12 VDD.n11 3.1505
R58 VDD.n10 VDD.n9 3.1505
R59 VDD.n2 VDD.n1 2.9292
R60 VDD.n4 VDD.n3 1.87106
R61 VDD.n1 VDD.t6 1.8205
R62 VDD.n1 VDD.n0 1.8205
R63 VDD.n3 VDD.n2 0.578642
R64 VDD.n9 VDD.n8 0.134373
R65 VDD VDD.n13 0.0760357
R66 VDD.n13 VDD.n10 0.0760357
R67 VDD VDD.n2 0.0647857
R68 VDD.n10 VDD.n7 0.0422857
R69 B B.n0 57.1693
R70 B.t2 B.t1 55.0112
R71 B.n0 B.t2 29.9826
R72 B.n0 B.t0 9.1255
R73 OUT.n2 OUT.n0 7.06041
R74 OUT.n2 OUT.n1 5.10528
R75 OUT OUT.n2 0.0533261
C0 VDD B 0.104f
C1 OUT a_168_68# 0.0558f
C2 OUT a_24_68# 0.0273f
C3 A B 0.0425f
C4 a_168_68# VDD 0.527f
C5 a_24_68# VDD 0.0116f
C6 A a_168_68# 0.123f
C7 A a_24_68# 0.0803f
C8 a_168_68# B 0.0713f
C9 a_24_68# B 0.0465f
C10 OUT VDD 0.149f
C11 A OUT 2.75e-19
C12 a_168_68# a_24_68# 0.361f
C13 A VDD 0.149f
C14 OUT B 0.0238f
.ends

