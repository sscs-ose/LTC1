magic
tech gf180mcuC
magscale 1 10
timestamp 1694601504
<< metal1 >>
rect 53 1041 171 1159
rect -87 371 -5 435
rect 276 359 532 477
rect 733 359 958 477
rect 39 -224 157 -106
use Inv_4x  Inv_4x_0
timestamp 1694581763
transform 1 0 447 0 1 -34
box -58 -203 511 1214
use Inv_4x  Inv_4x_1
timestamp 1694581763
transform 1 0 -117 0 1 -34
box -58 -203 511 1214
<< labels >>
flabel metal1 115 1088 115 1088 0 FreeSans 1600 0 0 0 VDD
port 0 nsew
flabel metal1 92 -176 92 -176 0 FreeSans 1600 0 0 0 VSS
port 1 nsew
flabel metal1 884 410 884 410 0 FreeSans 1600 0 0 0 OUT
port 2 nsew
flabel metal1 -50 404 -50 404 0 FreeSans 1600 0 0 0 IN
port 3 nsew
flabel metal1 385 407 385 407 0 FreeSans 1600 0 0 0 M
port 4 nsew
<< end >>
