magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -2332 -2118 2332 2118
<< pwell >>
rect -332 -118 332 118
<< nmos >>
rect -220 -50 -52 50
rect 52 -50 220 50
<< ndiff >>
rect -308 23 -220 50
rect -308 -23 -295 23
rect -249 -23 -220 23
rect -308 -50 -220 -23
rect -52 23 52 50
rect -52 -23 -23 23
rect 23 -23 52 23
rect -52 -50 52 -23
rect 220 23 308 50
rect 220 -23 249 23
rect 295 -23 308 23
rect 220 -50 308 -23
<< ndiffc >>
rect -295 -23 -249 23
rect -23 -23 23 23
rect 249 -23 295 23
<< polysilicon >>
rect -220 50 -52 94
rect 52 50 220 94
rect -220 -94 -52 -50
rect 52 -94 220 -50
<< metal1 >>
rect -295 23 -249 48
rect -295 -48 -249 -23
rect -23 23 23 48
rect -23 -48 23 -23
rect 249 23 295 48
rect 249 -48 295 -23
<< end >>
