magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1505 -1073 1505 1073
<< metal1 >>
rect -505 67 505 73
rect -505 41 -499 67
rect -473 41 -445 67
rect -419 41 -391 67
rect -365 41 -337 67
rect -311 41 -283 67
rect -257 41 -229 67
rect -203 41 -175 67
rect -149 41 -121 67
rect -95 41 -67 67
rect -41 41 -13 67
rect 13 41 41 67
rect 67 41 95 67
rect 121 41 149 67
rect 175 41 203 67
rect 229 41 257 67
rect 283 41 311 67
rect 337 41 365 67
rect 391 41 419 67
rect 445 41 473 67
rect 499 41 505 67
rect -505 13 505 41
rect -505 -13 -499 13
rect -473 -13 -445 13
rect -419 -13 -391 13
rect -365 -13 -337 13
rect -311 -13 -283 13
rect -257 -13 -229 13
rect -203 -13 -175 13
rect -149 -13 -121 13
rect -95 -13 -67 13
rect -41 -13 -13 13
rect 13 -13 41 13
rect 67 -13 95 13
rect 121 -13 149 13
rect 175 -13 203 13
rect 229 -13 257 13
rect 283 -13 311 13
rect 337 -13 365 13
rect 391 -13 419 13
rect 445 -13 473 13
rect 499 -13 505 13
rect -505 -41 505 -13
rect -505 -67 -499 -41
rect -473 -67 -445 -41
rect -419 -67 -391 -41
rect -365 -67 -337 -41
rect -311 -67 -283 -41
rect -257 -67 -229 -41
rect -203 -67 -175 -41
rect -149 -67 -121 -41
rect -95 -67 -67 -41
rect -41 -67 -13 -41
rect 13 -67 41 -41
rect 67 -67 95 -41
rect 121 -67 149 -41
rect 175 -67 203 -41
rect 229 -67 257 -41
rect 283 -67 311 -41
rect 337 -67 365 -41
rect 391 -67 419 -41
rect 445 -67 473 -41
rect 499 -67 505 -41
rect -505 -73 505 -67
<< via1 >>
rect -499 41 -473 67
rect -445 41 -419 67
rect -391 41 -365 67
rect -337 41 -311 67
rect -283 41 -257 67
rect -229 41 -203 67
rect -175 41 -149 67
rect -121 41 -95 67
rect -67 41 -41 67
rect -13 41 13 67
rect 41 41 67 67
rect 95 41 121 67
rect 149 41 175 67
rect 203 41 229 67
rect 257 41 283 67
rect 311 41 337 67
rect 365 41 391 67
rect 419 41 445 67
rect 473 41 499 67
rect -499 -13 -473 13
rect -445 -13 -419 13
rect -391 -13 -365 13
rect -337 -13 -311 13
rect -283 -13 -257 13
rect -229 -13 -203 13
rect -175 -13 -149 13
rect -121 -13 -95 13
rect -67 -13 -41 13
rect -13 -13 13 13
rect 41 -13 67 13
rect 95 -13 121 13
rect 149 -13 175 13
rect 203 -13 229 13
rect 257 -13 283 13
rect 311 -13 337 13
rect 365 -13 391 13
rect 419 -13 445 13
rect 473 -13 499 13
rect -499 -67 -473 -41
rect -445 -67 -419 -41
rect -391 -67 -365 -41
rect -337 -67 -311 -41
rect -283 -67 -257 -41
rect -229 -67 -203 -41
rect -175 -67 -149 -41
rect -121 -67 -95 -41
rect -67 -67 -41 -41
rect -13 -67 13 -41
rect 41 -67 67 -41
rect 95 -67 121 -41
rect 149 -67 175 -41
rect 203 -67 229 -41
rect 257 -67 283 -41
rect 311 -67 337 -41
rect 365 -67 391 -41
rect 419 -67 445 -41
rect 473 -67 499 -41
<< metal2 >>
rect -505 67 505 73
rect -505 41 -499 67
rect -473 41 -445 67
rect -419 41 -391 67
rect -365 41 -337 67
rect -311 41 -283 67
rect -257 41 -229 67
rect -203 41 -175 67
rect -149 41 -121 67
rect -95 41 -67 67
rect -41 41 -13 67
rect 13 41 41 67
rect 67 41 95 67
rect 121 41 149 67
rect 175 41 203 67
rect 229 41 257 67
rect 283 41 311 67
rect 337 41 365 67
rect 391 41 419 67
rect 445 41 473 67
rect 499 41 505 67
rect -505 13 505 41
rect -505 -13 -499 13
rect -473 -13 -445 13
rect -419 -13 -391 13
rect -365 -13 -337 13
rect -311 -13 -283 13
rect -257 -13 -229 13
rect -203 -13 -175 13
rect -149 -13 -121 13
rect -95 -13 -67 13
rect -41 -13 -13 13
rect 13 -13 41 13
rect 67 -13 95 13
rect 121 -13 149 13
rect 175 -13 203 13
rect 229 -13 257 13
rect 283 -13 311 13
rect 337 -13 365 13
rect 391 -13 419 13
rect 445 -13 473 13
rect 499 -13 505 13
rect -505 -41 505 -13
rect -505 -67 -499 -41
rect -473 -67 -445 -41
rect -419 -67 -391 -41
rect -365 -67 -337 -41
rect -311 -67 -283 -41
rect -257 -67 -229 -41
rect -203 -67 -175 -41
rect -149 -67 -121 -41
rect -95 -67 -67 -41
rect -41 -67 -13 -41
rect 13 -67 41 -41
rect 67 -67 95 -41
rect 121 -67 149 -41
rect 175 -67 203 -41
rect 229 -67 257 -41
rect 283 -67 311 -41
rect 337 -67 365 -41
rect 391 -67 419 -41
rect 445 -67 473 -41
rect 499 -67 505 -41
rect -505 -73 505 -67
<< end >>
