magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2913 -2975 2913 2975
<< psubdiff >>
rect -913 953 913 975
rect -913 907 -891 953
rect -845 907 -767 953
rect -721 907 -643 953
rect -597 907 -519 953
rect -473 907 -395 953
rect -349 907 -271 953
rect -225 907 -147 953
rect -101 907 -23 953
rect 23 907 101 953
rect 147 907 225 953
rect 271 907 349 953
rect 395 907 473 953
rect 519 907 597 953
rect 643 907 721 953
rect 767 907 845 953
rect 891 907 913 953
rect -913 829 913 907
rect -913 783 -891 829
rect -845 783 -767 829
rect -721 783 -643 829
rect -597 783 -519 829
rect -473 783 -395 829
rect -349 783 -271 829
rect -225 783 -147 829
rect -101 783 -23 829
rect 23 783 101 829
rect 147 783 225 829
rect 271 783 349 829
rect 395 783 473 829
rect 519 783 597 829
rect 643 783 721 829
rect 767 783 845 829
rect 891 783 913 829
rect -913 705 913 783
rect -913 659 -891 705
rect -845 659 -767 705
rect -721 659 -643 705
rect -597 659 -519 705
rect -473 659 -395 705
rect -349 659 -271 705
rect -225 659 -147 705
rect -101 659 -23 705
rect 23 659 101 705
rect 147 659 225 705
rect 271 659 349 705
rect 395 659 473 705
rect 519 659 597 705
rect 643 659 721 705
rect 767 659 845 705
rect 891 659 913 705
rect -913 581 913 659
rect -913 535 -891 581
rect -845 535 -767 581
rect -721 535 -643 581
rect -597 535 -519 581
rect -473 535 -395 581
rect -349 535 -271 581
rect -225 535 -147 581
rect -101 535 -23 581
rect 23 535 101 581
rect 147 535 225 581
rect 271 535 349 581
rect 395 535 473 581
rect 519 535 597 581
rect 643 535 721 581
rect 767 535 845 581
rect 891 535 913 581
rect -913 457 913 535
rect -913 411 -891 457
rect -845 411 -767 457
rect -721 411 -643 457
rect -597 411 -519 457
rect -473 411 -395 457
rect -349 411 -271 457
rect -225 411 -147 457
rect -101 411 -23 457
rect 23 411 101 457
rect 147 411 225 457
rect 271 411 349 457
rect 395 411 473 457
rect 519 411 597 457
rect 643 411 721 457
rect 767 411 845 457
rect 891 411 913 457
rect -913 333 913 411
rect -913 287 -891 333
rect -845 287 -767 333
rect -721 287 -643 333
rect -597 287 -519 333
rect -473 287 -395 333
rect -349 287 -271 333
rect -225 287 -147 333
rect -101 287 -23 333
rect 23 287 101 333
rect 147 287 225 333
rect 271 287 349 333
rect 395 287 473 333
rect 519 287 597 333
rect 643 287 721 333
rect 767 287 845 333
rect 891 287 913 333
rect -913 209 913 287
rect -913 163 -891 209
rect -845 163 -767 209
rect -721 163 -643 209
rect -597 163 -519 209
rect -473 163 -395 209
rect -349 163 -271 209
rect -225 163 -147 209
rect -101 163 -23 209
rect 23 163 101 209
rect 147 163 225 209
rect 271 163 349 209
rect 395 163 473 209
rect 519 163 597 209
rect 643 163 721 209
rect 767 163 845 209
rect 891 163 913 209
rect -913 85 913 163
rect -913 39 -891 85
rect -845 39 -767 85
rect -721 39 -643 85
rect -597 39 -519 85
rect -473 39 -395 85
rect -349 39 -271 85
rect -225 39 -147 85
rect -101 39 -23 85
rect 23 39 101 85
rect 147 39 225 85
rect 271 39 349 85
rect 395 39 473 85
rect 519 39 597 85
rect 643 39 721 85
rect 767 39 845 85
rect 891 39 913 85
rect -913 -39 913 39
rect -913 -85 -891 -39
rect -845 -85 -767 -39
rect -721 -85 -643 -39
rect -597 -85 -519 -39
rect -473 -85 -395 -39
rect -349 -85 -271 -39
rect -225 -85 -147 -39
rect -101 -85 -23 -39
rect 23 -85 101 -39
rect 147 -85 225 -39
rect 271 -85 349 -39
rect 395 -85 473 -39
rect 519 -85 597 -39
rect 643 -85 721 -39
rect 767 -85 845 -39
rect 891 -85 913 -39
rect -913 -163 913 -85
rect -913 -209 -891 -163
rect -845 -209 -767 -163
rect -721 -209 -643 -163
rect -597 -209 -519 -163
rect -473 -209 -395 -163
rect -349 -209 -271 -163
rect -225 -209 -147 -163
rect -101 -209 -23 -163
rect 23 -209 101 -163
rect 147 -209 225 -163
rect 271 -209 349 -163
rect 395 -209 473 -163
rect 519 -209 597 -163
rect 643 -209 721 -163
rect 767 -209 845 -163
rect 891 -209 913 -163
rect -913 -287 913 -209
rect -913 -333 -891 -287
rect -845 -333 -767 -287
rect -721 -333 -643 -287
rect -597 -333 -519 -287
rect -473 -333 -395 -287
rect -349 -333 -271 -287
rect -225 -333 -147 -287
rect -101 -333 -23 -287
rect 23 -333 101 -287
rect 147 -333 225 -287
rect 271 -333 349 -287
rect 395 -333 473 -287
rect 519 -333 597 -287
rect 643 -333 721 -287
rect 767 -333 845 -287
rect 891 -333 913 -287
rect -913 -411 913 -333
rect -913 -457 -891 -411
rect -845 -457 -767 -411
rect -721 -457 -643 -411
rect -597 -457 -519 -411
rect -473 -457 -395 -411
rect -349 -457 -271 -411
rect -225 -457 -147 -411
rect -101 -457 -23 -411
rect 23 -457 101 -411
rect 147 -457 225 -411
rect 271 -457 349 -411
rect 395 -457 473 -411
rect 519 -457 597 -411
rect 643 -457 721 -411
rect 767 -457 845 -411
rect 891 -457 913 -411
rect -913 -535 913 -457
rect -913 -581 -891 -535
rect -845 -581 -767 -535
rect -721 -581 -643 -535
rect -597 -581 -519 -535
rect -473 -581 -395 -535
rect -349 -581 -271 -535
rect -225 -581 -147 -535
rect -101 -581 -23 -535
rect 23 -581 101 -535
rect 147 -581 225 -535
rect 271 -581 349 -535
rect 395 -581 473 -535
rect 519 -581 597 -535
rect 643 -581 721 -535
rect 767 -581 845 -535
rect 891 -581 913 -535
rect -913 -659 913 -581
rect -913 -705 -891 -659
rect -845 -705 -767 -659
rect -721 -705 -643 -659
rect -597 -705 -519 -659
rect -473 -705 -395 -659
rect -349 -705 -271 -659
rect -225 -705 -147 -659
rect -101 -705 -23 -659
rect 23 -705 101 -659
rect 147 -705 225 -659
rect 271 -705 349 -659
rect 395 -705 473 -659
rect 519 -705 597 -659
rect 643 -705 721 -659
rect 767 -705 845 -659
rect 891 -705 913 -659
rect -913 -783 913 -705
rect -913 -829 -891 -783
rect -845 -829 -767 -783
rect -721 -829 -643 -783
rect -597 -829 -519 -783
rect -473 -829 -395 -783
rect -349 -829 -271 -783
rect -225 -829 -147 -783
rect -101 -829 -23 -783
rect 23 -829 101 -783
rect 147 -829 225 -783
rect 271 -829 349 -783
rect 395 -829 473 -783
rect 519 -829 597 -783
rect 643 -829 721 -783
rect 767 -829 845 -783
rect 891 -829 913 -783
rect -913 -907 913 -829
rect -913 -953 -891 -907
rect -845 -953 -767 -907
rect -721 -953 -643 -907
rect -597 -953 -519 -907
rect -473 -953 -395 -907
rect -349 -953 -271 -907
rect -225 -953 -147 -907
rect -101 -953 -23 -907
rect 23 -953 101 -907
rect 147 -953 225 -907
rect 271 -953 349 -907
rect 395 -953 473 -907
rect 519 -953 597 -907
rect 643 -953 721 -907
rect 767 -953 845 -907
rect 891 -953 913 -907
rect -913 -975 913 -953
<< psubdiffcont >>
rect -891 907 -845 953
rect -767 907 -721 953
rect -643 907 -597 953
rect -519 907 -473 953
rect -395 907 -349 953
rect -271 907 -225 953
rect -147 907 -101 953
rect -23 907 23 953
rect 101 907 147 953
rect 225 907 271 953
rect 349 907 395 953
rect 473 907 519 953
rect 597 907 643 953
rect 721 907 767 953
rect 845 907 891 953
rect -891 783 -845 829
rect -767 783 -721 829
rect -643 783 -597 829
rect -519 783 -473 829
rect -395 783 -349 829
rect -271 783 -225 829
rect -147 783 -101 829
rect -23 783 23 829
rect 101 783 147 829
rect 225 783 271 829
rect 349 783 395 829
rect 473 783 519 829
rect 597 783 643 829
rect 721 783 767 829
rect 845 783 891 829
rect -891 659 -845 705
rect -767 659 -721 705
rect -643 659 -597 705
rect -519 659 -473 705
rect -395 659 -349 705
rect -271 659 -225 705
rect -147 659 -101 705
rect -23 659 23 705
rect 101 659 147 705
rect 225 659 271 705
rect 349 659 395 705
rect 473 659 519 705
rect 597 659 643 705
rect 721 659 767 705
rect 845 659 891 705
rect -891 535 -845 581
rect -767 535 -721 581
rect -643 535 -597 581
rect -519 535 -473 581
rect -395 535 -349 581
rect -271 535 -225 581
rect -147 535 -101 581
rect -23 535 23 581
rect 101 535 147 581
rect 225 535 271 581
rect 349 535 395 581
rect 473 535 519 581
rect 597 535 643 581
rect 721 535 767 581
rect 845 535 891 581
rect -891 411 -845 457
rect -767 411 -721 457
rect -643 411 -597 457
rect -519 411 -473 457
rect -395 411 -349 457
rect -271 411 -225 457
rect -147 411 -101 457
rect -23 411 23 457
rect 101 411 147 457
rect 225 411 271 457
rect 349 411 395 457
rect 473 411 519 457
rect 597 411 643 457
rect 721 411 767 457
rect 845 411 891 457
rect -891 287 -845 333
rect -767 287 -721 333
rect -643 287 -597 333
rect -519 287 -473 333
rect -395 287 -349 333
rect -271 287 -225 333
rect -147 287 -101 333
rect -23 287 23 333
rect 101 287 147 333
rect 225 287 271 333
rect 349 287 395 333
rect 473 287 519 333
rect 597 287 643 333
rect 721 287 767 333
rect 845 287 891 333
rect -891 163 -845 209
rect -767 163 -721 209
rect -643 163 -597 209
rect -519 163 -473 209
rect -395 163 -349 209
rect -271 163 -225 209
rect -147 163 -101 209
rect -23 163 23 209
rect 101 163 147 209
rect 225 163 271 209
rect 349 163 395 209
rect 473 163 519 209
rect 597 163 643 209
rect 721 163 767 209
rect 845 163 891 209
rect -891 39 -845 85
rect -767 39 -721 85
rect -643 39 -597 85
rect -519 39 -473 85
rect -395 39 -349 85
rect -271 39 -225 85
rect -147 39 -101 85
rect -23 39 23 85
rect 101 39 147 85
rect 225 39 271 85
rect 349 39 395 85
rect 473 39 519 85
rect 597 39 643 85
rect 721 39 767 85
rect 845 39 891 85
rect -891 -85 -845 -39
rect -767 -85 -721 -39
rect -643 -85 -597 -39
rect -519 -85 -473 -39
rect -395 -85 -349 -39
rect -271 -85 -225 -39
rect -147 -85 -101 -39
rect -23 -85 23 -39
rect 101 -85 147 -39
rect 225 -85 271 -39
rect 349 -85 395 -39
rect 473 -85 519 -39
rect 597 -85 643 -39
rect 721 -85 767 -39
rect 845 -85 891 -39
rect -891 -209 -845 -163
rect -767 -209 -721 -163
rect -643 -209 -597 -163
rect -519 -209 -473 -163
rect -395 -209 -349 -163
rect -271 -209 -225 -163
rect -147 -209 -101 -163
rect -23 -209 23 -163
rect 101 -209 147 -163
rect 225 -209 271 -163
rect 349 -209 395 -163
rect 473 -209 519 -163
rect 597 -209 643 -163
rect 721 -209 767 -163
rect 845 -209 891 -163
rect -891 -333 -845 -287
rect -767 -333 -721 -287
rect -643 -333 -597 -287
rect -519 -333 -473 -287
rect -395 -333 -349 -287
rect -271 -333 -225 -287
rect -147 -333 -101 -287
rect -23 -333 23 -287
rect 101 -333 147 -287
rect 225 -333 271 -287
rect 349 -333 395 -287
rect 473 -333 519 -287
rect 597 -333 643 -287
rect 721 -333 767 -287
rect 845 -333 891 -287
rect -891 -457 -845 -411
rect -767 -457 -721 -411
rect -643 -457 -597 -411
rect -519 -457 -473 -411
rect -395 -457 -349 -411
rect -271 -457 -225 -411
rect -147 -457 -101 -411
rect -23 -457 23 -411
rect 101 -457 147 -411
rect 225 -457 271 -411
rect 349 -457 395 -411
rect 473 -457 519 -411
rect 597 -457 643 -411
rect 721 -457 767 -411
rect 845 -457 891 -411
rect -891 -581 -845 -535
rect -767 -581 -721 -535
rect -643 -581 -597 -535
rect -519 -581 -473 -535
rect -395 -581 -349 -535
rect -271 -581 -225 -535
rect -147 -581 -101 -535
rect -23 -581 23 -535
rect 101 -581 147 -535
rect 225 -581 271 -535
rect 349 -581 395 -535
rect 473 -581 519 -535
rect 597 -581 643 -535
rect 721 -581 767 -535
rect 845 -581 891 -535
rect -891 -705 -845 -659
rect -767 -705 -721 -659
rect -643 -705 -597 -659
rect -519 -705 -473 -659
rect -395 -705 -349 -659
rect -271 -705 -225 -659
rect -147 -705 -101 -659
rect -23 -705 23 -659
rect 101 -705 147 -659
rect 225 -705 271 -659
rect 349 -705 395 -659
rect 473 -705 519 -659
rect 597 -705 643 -659
rect 721 -705 767 -659
rect 845 -705 891 -659
rect -891 -829 -845 -783
rect -767 -829 -721 -783
rect -643 -829 -597 -783
rect -519 -829 -473 -783
rect -395 -829 -349 -783
rect -271 -829 -225 -783
rect -147 -829 -101 -783
rect -23 -829 23 -783
rect 101 -829 147 -783
rect 225 -829 271 -783
rect 349 -829 395 -783
rect 473 -829 519 -783
rect 597 -829 643 -783
rect 721 -829 767 -783
rect 845 -829 891 -783
rect -891 -953 -845 -907
rect -767 -953 -721 -907
rect -643 -953 -597 -907
rect -519 -953 -473 -907
rect -395 -953 -349 -907
rect -271 -953 -225 -907
rect -147 -953 -101 -907
rect -23 -953 23 -907
rect 101 -953 147 -907
rect 225 -953 271 -907
rect 349 -953 395 -907
rect 473 -953 519 -907
rect 597 -953 643 -907
rect 721 -953 767 -907
rect 845 -953 891 -907
<< metal1 >>
rect -902 953 902 964
rect -902 907 -891 953
rect -845 907 -767 953
rect -721 907 -643 953
rect -597 907 -519 953
rect -473 907 -395 953
rect -349 907 -271 953
rect -225 907 -147 953
rect -101 907 -23 953
rect 23 907 101 953
rect 147 907 225 953
rect 271 907 349 953
rect 395 907 473 953
rect 519 907 597 953
rect 643 907 721 953
rect 767 907 845 953
rect 891 907 902 953
rect -902 829 902 907
rect -902 783 -891 829
rect -845 783 -767 829
rect -721 783 -643 829
rect -597 783 -519 829
rect -473 783 -395 829
rect -349 783 -271 829
rect -225 783 -147 829
rect -101 783 -23 829
rect 23 783 101 829
rect 147 783 225 829
rect 271 783 349 829
rect 395 783 473 829
rect 519 783 597 829
rect 643 783 721 829
rect 767 783 845 829
rect 891 783 902 829
rect -902 705 902 783
rect -902 659 -891 705
rect -845 659 -767 705
rect -721 659 -643 705
rect -597 659 -519 705
rect -473 659 -395 705
rect -349 659 -271 705
rect -225 659 -147 705
rect -101 659 -23 705
rect 23 659 101 705
rect 147 659 225 705
rect 271 659 349 705
rect 395 659 473 705
rect 519 659 597 705
rect 643 659 721 705
rect 767 659 845 705
rect 891 659 902 705
rect -902 581 902 659
rect -902 535 -891 581
rect -845 535 -767 581
rect -721 535 -643 581
rect -597 535 -519 581
rect -473 535 -395 581
rect -349 535 -271 581
rect -225 535 -147 581
rect -101 535 -23 581
rect 23 535 101 581
rect 147 535 225 581
rect 271 535 349 581
rect 395 535 473 581
rect 519 535 597 581
rect 643 535 721 581
rect 767 535 845 581
rect 891 535 902 581
rect -902 457 902 535
rect -902 411 -891 457
rect -845 411 -767 457
rect -721 411 -643 457
rect -597 411 -519 457
rect -473 411 -395 457
rect -349 411 -271 457
rect -225 411 -147 457
rect -101 411 -23 457
rect 23 411 101 457
rect 147 411 225 457
rect 271 411 349 457
rect 395 411 473 457
rect 519 411 597 457
rect 643 411 721 457
rect 767 411 845 457
rect 891 411 902 457
rect -902 333 902 411
rect -902 287 -891 333
rect -845 287 -767 333
rect -721 287 -643 333
rect -597 287 -519 333
rect -473 287 -395 333
rect -349 287 -271 333
rect -225 287 -147 333
rect -101 287 -23 333
rect 23 287 101 333
rect 147 287 225 333
rect 271 287 349 333
rect 395 287 473 333
rect 519 287 597 333
rect 643 287 721 333
rect 767 287 845 333
rect 891 287 902 333
rect -902 209 902 287
rect -902 163 -891 209
rect -845 163 -767 209
rect -721 163 -643 209
rect -597 163 -519 209
rect -473 163 -395 209
rect -349 163 -271 209
rect -225 163 -147 209
rect -101 163 -23 209
rect 23 163 101 209
rect 147 163 225 209
rect 271 163 349 209
rect 395 163 473 209
rect 519 163 597 209
rect 643 163 721 209
rect 767 163 845 209
rect 891 163 902 209
rect -902 85 902 163
rect -902 39 -891 85
rect -845 39 -767 85
rect -721 39 -643 85
rect -597 39 -519 85
rect -473 39 -395 85
rect -349 39 -271 85
rect -225 39 -147 85
rect -101 39 -23 85
rect 23 39 101 85
rect 147 39 225 85
rect 271 39 349 85
rect 395 39 473 85
rect 519 39 597 85
rect 643 39 721 85
rect 767 39 845 85
rect 891 39 902 85
rect -902 -39 902 39
rect -902 -85 -891 -39
rect -845 -85 -767 -39
rect -721 -85 -643 -39
rect -597 -85 -519 -39
rect -473 -85 -395 -39
rect -349 -85 -271 -39
rect -225 -85 -147 -39
rect -101 -85 -23 -39
rect 23 -85 101 -39
rect 147 -85 225 -39
rect 271 -85 349 -39
rect 395 -85 473 -39
rect 519 -85 597 -39
rect 643 -85 721 -39
rect 767 -85 845 -39
rect 891 -85 902 -39
rect -902 -163 902 -85
rect -902 -209 -891 -163
rect -845 -209 -767 -163
rect -721 -209 -643 -163
rect -597 -209 -519 -163
rect -473 -209 -395 -163
rect -349 -209 -271 -163
rect -225 -209 -147 -163
rect -101 -209 -23 -163
rect 23 -209 101 -163
rect 147 -209 225 -163
rect 271 -209 349 -163
rect 395 -209 473 -163
rect 519 -209 597 -163
rect 643 -209 721 -163
rect 767 -209 845 -163
rect 891 -209 902 -163
rect -902 -287 902 -209
rect -902 -333 -891 -287
rect -845 -333 -767 -287
rect -721 -333 -643 -287
rect -597 -333 -519 -287
rect -473 -333 -395 -287
rect -349 -333 -271 -287
rect -225 -333 -147 -287
rect -101 -333 -23 -287
rect 23 -333 101 -287
rect 147 -333 225 -287
rect 271 -333 349 -287
rect 395 -333 473 -287
rect 519 -333 597 -287
rect 643 -333 721 -287
rect 767 -333 845 -287
rect 891 -333 902 -287
rect -902 -411 902 -333
rect -902 -457 -891 -411
rect -845 -457 -767 -411
rect -721 -457 -643 -411
rect -597 -457 -519 -411
rect -473 -457 -395 -411
rect -349 -457 -271 -411
rect -225 -457 -147 -411
rect -101 -457 -23 -411
rect 23 -457 101 -411
rect 147 -457 225 -411
rect 271 -457 349 -411
rect 395 -457 473 -411
rect 519 -457 597 -411
rect 643 -457 721 -411
rect 767 -457 845 -411
rect 891 -457 902 -411
rect -902 -535 902 -457
rect -902 -581 -891 -535
rect -845 -581 -767 -535
rect -721 -581 -643 -535
rect -597 -581 -519 -535
rect -473 -581 -395 -535
rect -349 -581 -271 -535
rect -225 -581 -147 -535
rect -101 -581 -23 -535
rect 23 -581 101 -535
rect 147 -581 225 -535
rect 271 -581 349 -535
rect 395 -581 473 -535
rect 519 -581 597 -535
rect 643 -581 721 -535
rect 767 -581 845 -535
rect 891 -581 902 -535
rect -902 -659 902 -581
rect -902 -705 -891 -659
rect -845 -705 -767 -659
rect -721 -705 -643 -659
rect -597 -705 -519 -659
rect -473 -705 -395 -659
rect -349 -705 -271 -659
rect -225 -705 -147 -659
rect -101 -705 -23 -659
rect 23 -705 101 -659
rect 147 -705 225 -659
rect 271 -705 349 -659
rect 395 -705 473 -659
rect 519 -705 597 -659
rect 643 -705 721 -659
rect 767 -705 845 -659
rect 891 -705 902 -659
rect -902 -783 902 -705
rect -902 -829 -891 -783
rect -845 -829 -767 -783
rect -721 -829 -643 -783
rect -597 -829 -519 -783
rect -473 -829 -395 -783
rect -349 -829 -271 -783
rect -225 -829 -147 -783
rect -101 -829 -23 -783
rect 23 -829 101 -783
rect 147 -829 225 -783
rect 271 -829 349 -783
rect 395 -829 473 -783
rect 519 -829 597 -783
rect 643 -829 721 -783
rect 767 -829 845 -783
rect 891 -829 902 -783
rect -902 -907 902 -829
rect -902 -953 -891 -907
rect -845 -953 -767 -907
rect -721 -953 -643 -907
rect -597 -953 -519 -907
rect -473 -953 -395 -907
rect -349 -953 -271 -907
rect -225 -953 -147 -907
rect -101 -953 -23 -907
rect 23 -953 101 -907
rect 147 -953 225 -907
rect 271 -953 349 -907
rect 395 -953 473 -907
rect 519 -953 597 -907
rect 643 -953 721 -907
rect 767 -953 845 -907
rect 891 -953 902 -907
rect -902 -964 902 -953
<< end >>
