magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1484 -1732 1484 1732
<< metal2 >>
rect -484 727 484 732
rect -484 699 -479 727
rect -451 699 -417 727
rect -389 699 -355 727
rect -327 699 -293 727
rect -265 699 -231 727
rect -203 699 -169 727
rect -141 699 -107 727
rect -79 699 -45 727
rect -17 699 17 727
rect 45 699 79 727
rect 107 699 141 727
rect 169 699 203 727
rect 231 699 265 727
rect 293 699 327 727
rect 355 699 389 727
rect 417 699 451 727
rect 479 699 484 727
rect -484 665 484 699
rect -484 637 -479 665
rect -451 637 -417 665
rect -389 637 -355 665
rect -327 637 -293 665
rect -265 637 -231 665
rect -203 637 -169 665
rect -141 637 -107 665
rect -79 637 -45 665
rect -17 637 17 665
rect 45 637 79 665
rect 107 637 141 665
rect 169 637 203 665
rect 231 637 265 665
rect 293 637 327 665
rect 355 637 389 665
rect 417 637 451 665
rect 479 637 484 665
rect -484 603 484 637
rect -484 575 -479 603
rect -451 575 -417 603
rect -389 575 -355 603
rect -327 575 -293 603
rect -265 575 -231 603
rect -203 575 -169 603
rect -141 575 -107 603
rect -79 575 -45 603
rect -17 575 17 603
rect 45 575 79 603
rect 107 575 141 603
rect 169 575 203 603
rect 231 575 265 603
rect 293 575 327 603
rect 355 575 389 603
rect 417 575 451 603
rect 479 575 484 603
rect -484 541 484 575
rect -484 513 -479 541
rect -451 513 -417 541
rect -389 513 -355 541
rect -327 513 -293 541
rect -265 513 -231 541
rect -203 513 -169 541
rect -141 513 -107 541
rect -79 513 -45 541
rect -17 513 17 541
rect 45 513 79 541
rect 107 513 141 541
rect 169 513 203 541
rect 231 513 265 541
rect 293 513 327 541
rect 355 513 389 541
rect 417 513 451 541
rect 479 513 484 541
rect -484 479 484 513
rect -484 451 -479 479
rect -451 451 -417 479
rect -389 451 -355 479
rect -327 451 -293 479
rect -265 451 -231 479
rect -203 451 -169 479
rect -141 451 -107 479
rect -79 451 -45 479
rect -17 451 17 479
rect 45 451 79 479
rect 107 451 141 479
rect 169 451 203 479
rect 231 451 265 479
rect 293 451 327 479
rect 355 451 389 479
rect 417 451 451 479
rect 479 451 484 479
rect -484 417 484 451
rect -484 389 -479 417
rect -451 389 -417 417
rect -389 389 -355 417
rect -327 389 -293 417
rect -265 389 -231 417
rect -203 389 -169 417
rect -141 389 -107 417
rect -79 389 -45 417
rect -17 389 17 417
rect 45 389 79 417
rect 107 389 141 417
rect 169 389 203 417
rect 231 389 265 417
rect 293 389 327 417
rect 355 389 389 417
rect 417 389 451 417
rect 479 389 484 417
rect -484 355 484 389
rect -484 327 -479 355
rect -451 327 -417 355
rect -389 327 -355 355
rect -327 327 -293 355
rect -265 327 -231 355
rect -203 327 -169 355
rect -141 327 -107 355
rect -79 327 -45 355
rect -17 327 17 355
rect 45 327 79 355
rect 107 327 141 355
rect 169 327 203 355
rect 231 327 265 355
rect 293 327 327 355
rect 355 327 389 355
rect 417 327 451 355
rect 479 327 484 355
rect -484 293 484 327
rect -484 265 -479 293
rect -451 265 -417 293
rect -389 265 -355 293
rect -327 265 -293 293
rect -265 265 -231 293
rect -203 265 -169 293
rect -141 265 -107 293
rect -79 265 -45 293
rect -17 265 17 293
rect 45 265 79 293
rect 107 265 141 293
rect 169 265 203 293
rect 231 265 265 293
rect 293 265 327 293
rect 355 265 389 293
rect 417 265 451 293
rect 479 265 484 293
rect -484 231 484 265
rect -484 203 -479 231
rect -451 203 -417 231
rect -389 203 -355 231
rect -327 203 -293 231
rect -265 203 -231 231
rect -203 203 -169 231
rect -141 203 -107 231
rect -79 203 -45 231
rect -17 203 17 231
rect 45 203 79 231
rect 107 203 141 231
rect 169 203 203 231
rect 231 203 265 231
rect 293 203 327 231
rect 355 203 389 231
rect 417 203 451 231
rect 479 203 484 231
rect -484 169 484 203
rect -484 141 -479 169
rect -451 141 -417 169
rect -389 141 -355 169
rect -327 141 -293 169
rect -265 141 -231 169
rect -203 141 -169 169
rect -141 141 -107 169
rect -79 141 -45 169
rect -17 141 17 169
rect 45 141 79 169
rect 107 141 141 169
rect 169 141 203 169
rect 231 141 265 169
rect 293 141 327 169
rect 355 141 389 169
rect 417 141 451 169
rect 479 141 484 169
rect -484 107 484 141
rect -484 79 -479 107
rect -451 79 -417 107
rect -389 79 -355 107
rect -327 79 -293 107
rect -265 79 -231 107
rect -203 79 -169 107
rect -141 79 -107 107
rect -79 79 -45 107
rect -17 79 17 107
rect 45 79 79 107
rect 107 79 141 107
rect 169 79 203 107
rect 231 79 265 107
rect 293 79 327 107
rect 355 79 389 107
rect 417 79 451 107
rect 479 79 484 107
rect -484 45 484 79
rect -484 17 -479 45
rect -451 17 -417 45
rect -389 17 -355 45
rect -327 17 -293 45
rect -265 17 -231 45
rect -203 17 -169 45
rect -141 17 -107 45
rect -79 17 -45 45
rect -17 17 17 45
rect 45 17 79 45
rect 107 17 141 45
rect 169 17 203 45
rect 231 17 265 45
rect 293 17 327 45
rect 355 17 389 45
rect 417 17 451 45
rect 479 17 484 45
rect -484 -17 484 17
rect -484 -45 -479 -17
rect -451 -45 -417 -17
rect -389 -45 -355 -17
rect -327 -45 -293 -17
rect -265 -45 -231 -17
rect -203 -45 -169 -17
rect -141 -45 -107 -17
rect -79 -45 -45 -17
rect -17 -45 17 -17
rect 45 -45 79 -17
rect 107 -45 141 -17
rect 169 -45 203 -17
rect 231 -45 265 -17
rect 293 -45 327 -17
rect 355 -45 389 -17
rect 417 -45 451 -17
rect 479 -45 484 -17
rect -484 -79 484 -45
rect -484 -107 -479 -79
rect -451 -107 -417 -79
rect -389 -107 -355 -79
rect -327 -107 -293 -79
rect -265 -107 -231 -79
rect -203 -107 -169 -79
rect -141 -107 -107 -79
rect -79 -107 -45 -79
rect -17 -107 17 -79
rect 45 -107 79 -79
rect 107 -107 141 -79
rect 169 -107 203 -79
rect 231 -107 265 -79
rect 293 -107 327 -79
rect 355 -107 389 -79
rect 417 -107 451 -79
rect 479 -107 484 -79
rect -484 -141 484 -107
rect -484 -169 -479 -141
rect -451 -169 -417 -141
rect -389 -169 -355 -141
rect -327 -169 -293 -141
rect -265 -169 -231 -141
rect -203 -169 -169 -141
rect -141 -169 -107 -141
rect -79 -169 -45 -141
rect -17 -169 17 -141
rect 45 -169 79 -141
rect 107 -169 141 -141
rect 169 -169 203 -141
rect 231 -169 265 -141
rect 293 -169 327 -141
rect 355 -169 389 -141
rect 417 -169 451 -141
rect 479 -169 484 -141
rect -484 -203 484 -169
rect -484 -231 -479 -203
rect -451 -231 -417 -203
rect -389 -231 -355 -203
rect -327 -231 -293 -203
rect -265 -231 -231 -203
rect -203 -231 -169 -203
rect -141 -231 -107 -203
rect -79 -231 -45 -203
rect -17 -231 17 -203
rect 45 -231 79 -203
rect 107 -231 141 -203
rect 169 -231 203 -203
rect 231 -231 265 -203
rect 293 -231 327 -203
rect 355 -231 389 -203
rect 417 -231 451 -203
rect 479 -231 484 -203
rect -484 -265 484 -231
rect -484 -293 -479 -265
rect -451 -293 -417 -265
rect -389 -293 -355 -265
rect -327 -293 -293 -265
rect -265 -293 -231 -265
rect -203 -293 -169 -265
rect -141 -293 -107 -265
rect -79 -293 -45 -265
rect -17 -293 17 -265
rect 45 -293 79 -265
rect 107 -293 141 -265
rect 169 -293 203 -265
rect 231 -293 265 -265
rect 293 -293 327 -265
rect 355 -293 389 -265
rect 417 -293 451 -265
rect 479 -293 484 -265
rect -484 -327 484 -293
rect -484 -355 -479 -327
rect -451 -355 -417 -327
rect -389 -355 -355 -327
rect -327 -355 -293 -327
rect -265 -355 -231 -327
rect -203 -355 -169 -327
rect -141 -355 -107 -327
rect -79 -355 -45 -327
rect -17 -355 17 -327
rect 45 -355 79 -327
rect 107 -355 141 -327
rect 169 -355 203 -327
rect 231 -355 265 -327
rect 293 -355 327 -327
rect 355 -355 389 -327
rect 417 -355 451 -327
rect 479 -355 484 -327
rect -484 -389 484 -355
rect -484 -417 -479 -389
rect -451 -417 -417 -389
rect -389 -417 -355 -389
rect -327 -417 -293 -389
rect -265 -417 -231 -389
rect -203 -417 -169 -389
rect -141 -417 -107 -389
rect -79 -417 -45 -389
rect -17 -417 17 -389
rect 45 -417 79 -389
rect 107 -417 141 -389
rect 169 -417 203 -389
rect 231 -417 265 -389
rect 293 -417 327 -389
rect 355 -417 389 -389
rect 417 -417 451 -389
rect 479 -417 484 -389
rect -484 -451 484 -417
rect -484 -479 -479 -451
rect -451 -479 -417 -451
rect -389 -479 -355 -451
rect -327 -479 -293 -451
rect -265 -479 -231 -451
rect -203 -479 -169 -451
rect -141 -479 -107 -451
rect -79 -479 -45 -451
rect -17 -479 17 -451
rect 45 -479 79 -451
rect 107 -479 141 -451
rect 169 -479 203 -451
rect 231 -479 265 -451
rect 293 -479 327 -451
rect 355 -479 389 -451
rect 417 -479 451 -451
rect 479 -479 484 -451
rect -484 -513 484 -479
rect -484 -541 -479 -513
rect -451 -541 -417 -513
rect -389 -541 -355 -513
rect -327 -541 -293 -513
rect -265 -541 -231 -513
rect -203 -541 -169 -513
rect -141 -541 -107 -513
rect -79 -541 -45 -513
rect -17 -541 17 -513
rect 45 -541 79 -513
rect 107 -541 141 -513
rect 169 -541 203 -513
rect 231 -541 265 -513
rect 293 -541 327 -513
rect 355 -541 389 -513
rect 417 -541 451 -513
rect 479 -541 484 -513
rect -484 -575 484 -541
rect -484 -603 -479 -575
rect -451 -603 -417 -575
rect -389 -603 -355 -575
rect -327 -603 -293 -575
rect -265 -603 -231 -575
rect -203 -603 -169 -575
rect -141 -603 -107 -575
rect -79 -603 -45 -575
rect -17 -603 17 -575
rect 45 -603 79 -575
rect 107 -603 141 -575
rect 169 -603 203 -575
rect 231 -603 265 -575
rect 293 -603 327 -575
rect 355 -603 389 -575
rect 417 -603 451 -575
rect 479 -603 484 -575
rect -484 -637 484 -603
rect -484 -665 -479 -637
rect -451 -665 -417 -637
rect -389 -665 -355 -637
rect -327 -665 -293 -637
rect -265 -665 -231 -637
rect -203 -665 -169 -637
rect -141 -665 -107 -637
rect -79 -665 -45 -637
rect -17 -665 17 -637
rect 45 -665 79 -637
rect 107 -665 141 -637
rect 169 -665 203 -637
rect 231 -665 265 -637
rect 293 -665 327 -637
rect 355 -665 389 -637
rect 417 -665 451 -637
rect 479 -665 484 -637
rect -484 -699 484 -665
rect -484 -727 -479 -699
rect -451 -727 -417 -699
rect -389 -727 -355 -699
rect -327 -727 -293 -699
rect -265 -727 -231 -699
rect -203 -727 -169 -699
rect -141 -727 -107 -699
rect -79 -727 -45 -699
rect -17 -727 17 -699
rect 45 -727 79 -699
rect 107 -727 141 -699
rect 169 -727 203 -699
rect 231 -727 265 -699
rect 293 -727 327 -699
rect 355 -727 389 -699
rect 417 -727 451 -699
rect 479 -727 484 -699
rect -484 -732 484 -727
<< via2 >>
rect -479 699 -451 727
rect -417 699 -389 727
rect -355 699 -327 727
rect -293 699 -265 727
rect -231 699 -203 727
rect -169 699 -141 727
rect -107 699 -79 727
rect -45 699 -17 727
rect 17 699 45 727
rect 79 699 107 727
rect 141 699 169 727
rect 203 699 231 727
rect 265 699 293 727
rect 327 699 355 727
rect 389 699 417 727
rect 451 699 479 727
rect -479 637 -451 665
rect -417 637 -389 665
rect -355 637 -327 665
rect -293 637 -265 665
rect -231 637 -203 665
rect -169 637 -141 665
rect -107 637 -79 665
rect -45 637 -17 665
rect 17 637 45 665
rect 79 637 107 665
rect 141 637 169 665
rect 203 637 231 665
rect 265 637 293 665
rect 327 637 355 665
rect 389 637 417 665
rect 451 637 479 665
rect -479 575 -451 603
rect -417 575 -389 603
rect -355 575 -327 603
rect -293 575 -265 603
rect -231 575 -203 603
rect -169 575 -141 603
rect -107 575 -79 603
rect -45 575 -17 603
rect 17 575 45 603
rect 79 575 107 603
rect 141 575 169 603
rect 203 575 231 603
rect 265 575 293 603
rect 327 575 355 603
rect 389 575 417 603
rect 451 575 479 603
rect -479 513 -451 541
rect -417 513 -389 541
rect -355 513 -327 541
rect -293 513 -265 541
rect -231 513 -203 541
rect -169 513 -141 541
rect -107 513 -79 541
rect -45 513 -17 541
rect 17 513 45 541
rect 79 513 107 541
rect 141 513 169 541
rect 203 513 231 541
rect 265 513 293 541
rect 327 513 355 541
rect 389 513 417 541
rect 451 513 479 541
rect -479 451 -451 479
rect -417 451 -389 479
rect -355 451 -327 479
rect -293 451 -265 479
rect -231 451 -203 479
rect -169 451 -141 479
rect -107 451 -79 479
rect -45 451 -17 479
rect 17 451 45 479
rect 79 451 107 479
rect 141 451 169 479
rect 203 451 231 479
rect 265 451 293 479
rect 327 451 355 479
rect 389 451 417 479
rect 451 451 479 479
rect -479 389 -451 417
rect -417 389 -389 417
rect -355 389 -327 417
rect -293 389 -265 417
rect -231 389 -203 417
rect -169 389 -141 417
rect -107 389 -79 417
rect -45 389 -17 417
rect 17 389 45 417
rect 79 389 107 417
rect 141 389 169 417
rect 203 389 231 417
rect 265 389 293 417
rect 327 389 355 417
rect 389 389 417 417
rect 451 389 479 417
rect -479 327 -451 355
rect -417 327 -389 355
rect -355 327 -327 355
rect -293 327 -265 355
rect -231 327 -203 355
rect -169 327 -141 355
rect -107 327 -79 355
rect -45 327 -17 355
rect 17 327 45 355
rect 79 327 107 355
rect 141 327 169 355
rect 203 327 231 355
rect 265 327 293 355
rect 327 327 355 355
rect 389 327 417 355
rect 451 327 479 355
rect -479 265 -451 293
rect -417 265 -389 293
rect -355 265 -327 293
rect -293 265 -265 293
rect -231 265 -203 293
rect -169 265 -141 293
rect -107 265 -79 293
rect -45 265 -17 293
rect 17 265 45 293
rect 79 265 107 293
rect 141 265 169 293
rect 203 265 231 293
rect 265 265 293 293
rect 327 265 355 293
rect 389 265 417 293
rect 451 265 479 293
rect -479 203 -451 231
rect -417 203 -389 231
rect -355 203 -327 231
rect -293 203 -265 231
rect -231 203 -203 231
rect -169 203 -141 231
rect -107 203 -79 231
rect -45 203 -17 231
rect 17 203 45 231
rect 79 203 107 231
rect 141 203 169 231
rect 203 203 231 231
rect 265 203 293 231
rect 327 203 355 231
rect 389 203 417 231
rect 451 203 479 231
rect -479 141 -451 169
rect -417 141 -389 169
rect -355 141 -327 169
rect -293 141 -265 169
rect -231 141 -203 169
rect -169 141 -141 169
rect -107 141 -79 169
rect -45 141 -17 169
rect 17 141 45 169
rect 79 141 107 169
rect 141 141 169 169
rect 203 141 231 169
rect 265 141 293 169
rect 327 141 355 169
rect 389 141 417 169
rect 451 141 479 169
rect -479 79 -451 107
rect -417 79 -389 107
rect -355 79 -327 107
rect -293 79 -265 107
rect -231 79 -203 107
rect -169 79 -141 107
rect -107 79 -79 107
rect -45 79 -17 107
rect 17 79 45 107
rect 79 79 107 107
rect 141 79 169 107
rect 203 79 231 107
rect 265 79 293 107
rect 327 79 355 107
rect 389 79 417 107
rect 451 79 479 107
rect -479 17 -451 45
rect -417 17 -389 45
rect -355 17 -327 45
rect -293 17 -265 45
rect -231 17 -203 45
rect -169 17 -141 45
rect -107 17 -79 45
rect -45 17 -17 45
rect 17 17 45 45
rect 79 17 107 45
rect 141 17 169 45
rect 203 17 231 45
rect 265 17 293 45
rect 327 17 355 45
rect 389 17 417 45
rect 451 17 479 45
rect -479 -45 -451 -17
rect -417 -45 -389 -17
rect -355 -45 -327 -17
rect -293 -45 -265 -17
rect -231 -45 -203 -17
rect -169 -45 -141 -17
rect -107 -45 -79 -17
rect -45 -45 -17 -17
rect 17 -45 45 -17
rect 79 -45 107 -17
rect 141 -45 169 -17
rect 203 -45 231 -17
rect 265 -45 293 -17
rect 327 -45 355 -17
rect 389 -45 417 -17
rect 451 -45 479 -17
rect -479 -107 -451 -79
rect -417 -107 -389 -79
rect -355 -107 -327 -79
rect -293 -107 -265 -79
rect -231 -107 -203 -79
rect -169 -107 -141 -79
rect -107 -107 -79 -79
rect -45 -107 -17 -79
rect 17 -107 45 -79
rect 79 -107 107 -79
rect 141 -107 169 -79
rect 203 -107 231 -79
rect 265 -107 293 -79
rect 327 -107 355 -79
rect 389 -107 417 -79
rect 451 -107 479 -79
rect -479 -169 -451 -141
rect -417 -169 -389 -141
rect -355 -169 -327 -141
rect -293 -169 -265 -141
rect -231 -169 -203 -141
rect -169 -169 -141 -141
rect -107 -169 -79 -141
rect -45 -169 -17 -141
rect 17 -169 45 -141
rect 79 -169 107 -141
rect 141 -169 169 -141
rect 203 -169 231 -141
rect 265 -169 293 -141
rect 327 -169 355 -141
rect 389 -169 417 -141
rect 451 -169 479 -141
rect -479 -231 -451 -203
rect -417 -231 -389 -203
rect -355 -231 -327 -203
rect -293 -231 -265 -203
rect -231 -231 -203 -203
rect -169 -231 -141 -203
rect -107 -231 -79 -203
rect -45 -231 -17 -203
rect 17 -231 45 -203
rect 79 -231 107 -203
rect 141 -231 169 -203
rect 203 -231 231 -203
rect 265 -231 293 -203
rect 327 -231 355 -203
rect 389 -231 417 -203
rect 451 -231 479 -203
rect -479 -293 -451 -265
rect -417 -293 -389 -265
rect -355 -293 -327 -265
rect -293 -293 -265 -265
rect -231 -293 -203 -265
rect -169 -293 -141 -265
rect -107 -293 -79 -265
rect -45 -293 -17 -265
rect 17 -293 45 -265
rect 79 -293 107 -265
rect 141 -293 169 -265
rect 203 -293 231 -265
rect 265 -293 293 -265
rect 327 -293 355 -265
rect 389 -293 417 -265
rect 451 -293 479 -265
rect -479 -355 -451 -327
rect -417 -355 -389 -327
rect -355 -355 -327 -327
rect -293 -355 -265 -327
rect -231 -355 -203 -327
rect -169 -355 -141 -327
rect -107 -355 -79 -327
rect -45 -355 -17 -327
rect 17 -355 45 -327
rect 79 -355 107 -327
rect 141 -355 169 -327
rect 203 -355 231 -327
rect 265 -355 293 -327
rect 327 -355 355 -327
rect 389 -355 417 -327
rect 451 -355 479 -327
rect -479 -417 -451 -389
rect -417 -417 -389 -389
rect -355 -417 -327 -389
rect -293 -417 -265 -389
rect -231 -417 -203 -389
rect -169 -417 -141 -389
rect -107 -417 -79 -389
rect -45 -417 -17 -389
rect 17 -417 45 -389
rect 79 -417 107 -389
rect 141 -417 169 -389
rect 203 -417 231 -389
rect 265 -417 293 -389
rect 327 -417 355 -389
rect 389 -417 417 -389
rect 451 -417 479 -389
rect -479 -479 -451 -451
rect -417 -479 -389 -451
rect -355 -479 -327 -451
rect -293 -479 -265 -451
rect -231 -479 -203 -451
rect -169 -479 -141 -451
rect -107 -479 -79 -451
rect -45 -479 -17 -451
rect 17 -479 45 -451
rect 79 -479 107 -451
rect 141 -479 169 -451
rect 203 -479 231 -451
rect 265 -479 293 -451
rect 327 -479 355 -451
rect 389 -479 417 -451
rect 451 -479 479 -451
rect -479 -541 -451 -513
rect -417 -541 -389 -513
rect -355 -541 -327 -513
rect -293 -541 -265 -513
rect -231 -541 -203 -513
rect -169 -541 -141 -513
rect -107 -541 -79 -513
rect -45 -541 -17 -513
rect 17 -541 45 -513
rect 79 -541 107 -513
rect 141 -541 169 -513
rect 203 -541 231 -513
rect 265 -541 293 -513
rect 327 -541 355 -513
rect 389 -541 417 -513
rect 451 -541 479 -513
rect -479 -603 -451 -575
rect -417 -603 -389 -575
rect -355 -603 -327 -575
rect -293 -603 -265 -575
rect -231 -603 -203 -575
rect -169 -603 -141 -575
rect -107 -603 -79 -575
rect -45 -603 -17 -575
rect 17 -603 45 -575
rect 79 -603 107 -575
rect 141 -603 169 -575
rect 203 -603 231 -575
rect 265 -603 293 -575
rect 327 -603 355 -575
rect 389 -603 417 -575
rect 451 -603 479 -575
rect -479 -665 -451 -637
rect -417 -665 -389 -637
rect -355 -665 -327 -637
rect -293 -665 -265 -637
rect -231 -665 -203 -637
rect -169 -665 -141 -637
rect -107 -665 -79 -637
rect -45 -665 -17 -637
rect 17 -665 45 -637
rect 79 -665 107 -637
rect 141 -665 169 -637
rect 203 -665 231 -637
rect 265 -665 293 -637
rect 327 -665 355 -637
rect 389 -665 417 -637
rect 451 -665 479 -637
rect -479 -727 -451 -699
rect -417 -727 -389 -699
rect -355 -727 -327 -699
rect -293 -727 -265 -699
rect -231 -727 -203 -699
rect -169 -727 -141 -699
rect -107 -727 -79 -699
rect -45 -727 -17 -699
rect 17 -727 45 -699
rect 79 -727 107 -699
rect 141 -727 169 -699
rect 203 -727 231 -699
rect 265 -727 293 -699
rect 327 -727 355 -699
rect 389 -727 417 -699
rect 451 -727 479 -699
<< metal3 >>
rect -484 727 484 732
rect -484 699 -479 727
rect -451 699 -417 727
rect -389 699 -355 727
rect -327 699 -293 727
rect -265 699 -231 727
rect -203 699 -169 727
rect -141 699 -107 727
rect -79 699 -45 727
rect -17 699 17 727
rect 45 699 79 727
rect 107 699 141 727
rect 169 699 203 727
rect 231 699 265 727
rect 293 699 327 727
rect 355 699 389 727
rect 417 699 451 727
rect 479 699 484 727
rect -484 665 484 699
rect -484 637 -479 665
rect -451 637 -417 665
rect -389 637 -355 665
rect -327 637 -293 665
rect -265 637 -231 665
rect -203 637 -169 665
rect -141 637 -107 665
rect -79 637 -45 665
rect -17 637 17 665
rect 45 637 79 665
rect 107 637 141 665
rect 169 637 203 665
rect 231 637 265 665
rect 293 637 327 665
rect 355 637 389 665
rect 417 637 451 665
rect 479 637 484 665
rect -484 603 484 637
rect -484 575 -479 603
rect -451 575 -417 603
rect -389 575 -355 603
rect -327 575 -293 603
rect -265 575 -231 603
rect -203 575 -169 603
rect -141 575 -107 603
rect -79 575 -45 603
rect -17 575 17 603
rect 45 575 79 603
rect 107 575 141 603
rect 169 575 203 603
rect 231 575 265 603
rect 293 575 327 603
rect 355 575 389 603
rect 417 575 451 603
rect 479 575 484 603
rect -484 541 484 575
rect -484 513 -479 541
rect -451 513 -417 541
rect -389 513 -355 541
rect -327 513 -293 541
rect -265 513 -231 541
rect -203 513 -169 541
rect -141 513 -107 541
rect -79 513 -45 541
rect -17 513 17 541
rect 45 513 79 541
rect 107 513 141 541
rect 169 513 203 541
rect 231 513 265 541
rect 293 513 327 541
rect 355 513 389 541
rect 417 513 451 541
rect 479 513 484 541
rect -484 479 484 513
rect -484 451 -479 479
rect -451 451 -417 479
rect -389 451 -355 479
rect -327 451 -293 479
rect -265 451 -231 479
rect -203 451 -169 479
rect -141 451 -107 479
rect -79 451 -45 479
rect -17 451 17 479
rect 45 451 79 479
rect 107 451 141 479
rect 169 451 203 479
rect 231 451 265 479
rect 293 451 327 479
rect 355 451 389 479
rect 417 451 451 479
rect 479 451 484 479
rect -484 417 484 451
rect -484 389 -479 417
rect -451 389 -417 417
rect -389 389 -355 417
rect -327 389 -293 417
rect -265 389 -231 417
rect -203 389 -169 417
rect -141 389 -107 417
rect -79 389 -45 417
rect -17 389 17 417
rect 45 389 79 417
rect 107 389 141 417
rect 169 389 203 417
rect 231 389 265 417
rect 293 389 327 417
rect 355 389 389 417
rect 417 389 451 417
rect 479 389 484 417
rect -484 355 484 389
rect -484 327 -479 355
rect -451 327 -417 355
rect -389 327 -355 355
rect -327 327 -293 355
rect -265 327 -231 355
rect -203 327 -169 355
rect -141 327 -107 355
rect -79 327 -45 355
rect -17 327 17 355
rect 45 327 79 355
rect 107 327 141 355
rect 169 327 203 355
rect 231 327 265 355
rect 293 327 327 355
rect 355 327 389 355
rect 417 327 451 355
rect 479 327 484 355
rect -484 293 484 327
rect -484 265 -479 293
rect -451 265 -417 293
rect -389 265 -355 293
rect -327 265 -293 293
rect -265 265 -231 293
rect -203 265 -169 293
rect -141 265 -107 293
rect -79 265 -45 293
rect -17 265 17 293
rect 45 265 79 293
rect 107 265 141 293
rect 169 265 203 293
rect 231 265 265 293
rect 293 265 327 293
rect 355 265 389 293
rect 417 265 451 293
rect 479 265 484 293
rect -484 231 484 265
rect -484 203 -479 231
rect -451 203 -417 231
rect -389 203 -355 231
rect -327 203 -293 231
rect -265 203 -231 231
rect -203 203 -169 231
rect -141 203 -107 231
rect -79 203 -45 231
rect -17 203 17 231
rect 45 203 79 231
rect 107 203 141 231
rect 169 203 203 231
rect 231 203 265 231
rect 293 203 327 231
rect 355 203 389 231
rect 417 203 451 231
rect 479 203 484 231
rect -484 169 484 203
rect -484 141 -479 169
rect -451 141 -417 169
rect -389 141 -355 169
rect -327 141 -293 169
rect -265 141 -231 169
rect -203 141 -169 169
rect -141 141 -107 169
rect -79 141 -45 169
rect -17 141 17 169
rect 45 141 79 169
rect 107 141 141 169
rect 169 141 203 169
rect 231 141 265 169
rect 293 141 327 169
rect 355 141 389 169
rect 417 141 451 169
rect 479 141 484 169
rect -484 107 484 141
rect -484 79 -479 107
rect -451 79 -417 107
rect -389 79 -355 107
rect -327 79 -293 107
rect -265 79 -231 107
rect -203 79 -169 107
rect -141 79 -107 107
rect -79 79 -45 107
rect -17 79 17 107
rect 45 79 79 107
rect 107 79 141 107
rect 169 79 203 107
rect 231 79 265 107
rect 293 79 327 107
rect 355 79 389 107
rect 417 79 451 107
rect 479 79 484 107
rect -484 45 484 79
rect -484 17 -479 45
rect -451 17 -417 45
rect -389 17 -355 45
rect -327 17 -293 45
rect -265 17 -231 45
rect -203 17 -169 45
rect -141 17 -107 45
rect -79 17 -45 45
rect -17 17 17 45
rect 45 17 79 45
rect 107 17 141 45
rect 169 17 203 45
rect 231 17 265 45
rect 293 17 327 45
rect 355 17 389 45
rect 417 17 451 45
rect 479 17 484 45
rect -484 -17 484 17
rect -484 -45 -479 -17
rect -451 -45 -417 -17
rect -389 -45 -355 -17
rect -327 -45 -293 -17
rect -265 -45 -231 -17
rect -203 -45 -169 -17
rect -141 -45 -107 -17
rect -79 -45 -45 -17
rect -17 -45 17 -17
rect 45 -45 79 -17
rect 107 -45 141 -17
rect 169 -45 203 -17
rect 231 -45 265 -17
rect 293 -45 327 -17
rect 355 -45 389 -17
rect 417 -45 451 -17
rect 479 -45 484 -17
rect -484 -79 484 -45
rect -484 -107 -479 -79
rect -451 -107 -417 -79
rect -389 -107 -355 -79
rect -327 -107 -293 -79
rect -265 -107 -231 -79
rect -203 -107 -169 -79
rect -141 -107 -107 -79
rect -79 -107 -45 -79
rect -17 -107 17 -79
rect 45 -107 79 -79
rect 107 -107 141 -79
rect 169 -107 203 -79
rect 231 -107 265 -79
rect 293 -107 327 -79
rect 355 -107 389 -79
rect 417 -107 451 -79
rect 479 -107 484 -79
rect -484 -141 484 -107
rect -484 -169 -479 -141
rect -451 -169 -417 -141
rect -389 -169 -355 -141
rect -327 -169 -293 -141
rect -265 -169 -231 -141
rect -203 -169 -169 -141
rect -141 -169 -107 -141
rect -79 -169 -45 -141
rect -17 -169 17 -141
rect 45 -169 79 -141
rect 107 -169 141 -141
rect 169 -169 203 -141
rect 231 -169 265 -141
rect 293 -169 327 -141
rect 355 -169 389 -141
rect 417 -169 451 -141
rect 479 -169 484 -141
rect -484 -203 484 -169
rect -484 -231 -479 -203
rect -451 -231 -417 -203
rect -389 -231 -355 -203
rect -327 -231 -293 -203
rect -265 -231 -231 -203
rect -203 -231 -169 -203
rect -141 -231 -107 -203
rect -79 -231 -45 -203
rect -17 -231 17 -203
rect 45 -231 79 -203
rect 107 -231 141 -203
rect 169 -231 203 -203
rect 231 -231 265 -203
rect 293 -231 327 -203
rect 355 -231 389 -203
rect 417 -231 451 -203
rect 479 -231 484 -203
rect -484 -265 484 -231
rect -484 -293 -479 -265
rect -451 -293 -417 -265
rect -389 -293 -355 -265
rect -327 -293 -293 -265
rect -265 -293 -231 -265
rect -203 -293 -169 -265
rect -141 -293 -107 -265
rect -79 -293 -45 -265
rect -17 -293 17 -265
rect 45 -293 79 -265
rect 107 -293 141 -265
rect 169 -293 203 -265
rect 231 -293 265 -265
rect 293 -293 327 -265
rect 355 -293 389 -265
rect 417 -293 451 -265
rect 479 -293 484 -265
rect -484 -327 484 -293
rect -484 -355 -479 -327
rect -451 -355 -417 -327
rect -389 -355 -355 -327
rect -327 -355 -293 -327
rect -265 -355 -231 -327
rect -203 -355 -169 -327
rect -141 -355 -107 -327
rect -79 -355 -45 -327
rect -17 -355 17 -327
rect 45 -355 79 -327
rect 107 -355 141 -327
rect 169 -355 203 -327
rect 231 -355 265 -327
rect 293 -355 327 -327
rect 355 -355 389 -327
rect 417 -355 451 -327
rect 479 -355 484 -327
rect -484 -389 484 -355
rect -484 -417 -479 -389
rect -451 -417 -417 -389
rect -389 -417 -355 -389
rect -327 -417 -293 -389
rect -265 -417 -231 -389
rect -203 -417 -169 -389
rect -141 -417 -107 -389
rect -79 -417 -45 -389
rect -17 -417 17 -389
rect 45 -417 79 -389
rect 107 -417 141 -389
rect 169 -417 203 -389
rect 231 -417 265 -389
rect 293 -417 327 -389
rect 355 -417 389 -389
rect 417 -417 451 -389
rect 479 -417 484 -389
rect -484 -451 484 -417
rect -484 -479 -479 -451
rect -451 -479 -417 -451
rect -389 -479 -355 -451
rect -327 -479 -293 -451
rect -265 -479 -231 -451
rect -203 -479 -169 -451
rect -141 -479 -107 -451
rect -79 -479 -45 -451
rect -17 -479 17 -451
rect 45 -479 79 -451
rect 107 -479 141 -451
rect 169 -479 203 -451
rect 231 -479 265 -451
rect 293 -479 327 -451
rect 355 -479 389 -451
rect 417 -479 451 -451
rect 479 -479 484 -451
rect -484 -513 484 -479
rect -484 -541 -479 -513
rect -451 -541 -417 -513
rect -389 -541 -355 -513
rect -327 -541 -293 -513
rect -265 -541 -231 -513
rect -203 -541 -169 -513
rect -141 -541 -107 -513
rect -79 -541 -45 -513
rect -17 -541 17 -513
rect 45 -541 79 -513
rect 107 -541 141 -513
rect 169 -541 203 -513
rect 231 -541 265 -513
rect 293 -541 327 -513
rect 355 -541 389 -513
rect 417 -541 451 -513
rect 479 -541 484 -513
rect -484 -575 484 -541
rect -484 -603 -479 -575
rect -451 -603 -417 -575
rect -389 -603 -355 -575
rect -327 -603 -293 -575
rect -265 -603 -231 -575
rect -203 -603 -169 -575
rect -141 -603 -107 -575
rect -79 -603 -45 -575
rect -17 -603 17 -575
rect 45 -603 79 -575
rect 107 -603 141 -575
rect 169 -603 203 -575
rect 231 -603 265 -575
rect 293 -603 327 -575
rect 355 -603 389 -575
rect 417 -603 451 -575
rect 479 -603 484 -575
rect -484 -637 484 -603
rect -484 -665 -479 -637
rect -451 -665 -417 -637
rect -389 -665 -355 -637
rect -327 -665 -293 -637
rect -265 -665 -231 -637
rect -203 -665 -169 -637
rect -141 -665 -107 -637
rect -79 -665 -45 -637
rect -17 -665 17 -637
rect 45 -665 79 -637
rect 107 -665 141 -637
rect 169 -665 203 -637
rect 231 -665 265 -637
rect 293 -665 327 -637
rect 355 -665 389 -637
rect 417 -665 451 -637
rect 479 -665 484 -637
rect -484 -699 484 -665
rect -484 -727 -479 -699
rect -451 -727 -417 -699
rect -389 -727 -355 -699
rect -327 -727 -293 -699
rect -265 -727 -231 -699
rect -203 -727 -169 -699
rect -141 -727 -107 -699
rect -79 -727 -45 -699
rect -17 -727 17 -699
rect 45 -727 79 -699
rect 107 -727 141 -699
rect 169 -727 203 -699
rect 231 -727 265 -699
rect 293 -727 327 -699
rect 355 -727 389 -699
rect 417 -727 451 -699
rect 479 -727 484 -699
rect -484 -732 484 -727
<< end >>
