magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -7678 -2728 7678 2728
<< nwell >>
rect -5678 -728 5678 728
<< nsubdiff >>
rect -5595 623 5595 645
rect -5595 -623 -5573 623
rect 5573 -623 5595 623
rect -5595 -645 5595 -623
<< nsubdiffcont >>
rect -5573 -623 5573 623
<< metal1 >>
rect -5584 623 5584 634
rect -5584 -623 -5573 623
rect 5573 -623 5584 623
rect -5584 -634 5584 -623
<< end >>
