magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1589 -1285 1589 1285
<< metal2 >>
rect -589 280 589 285
rect -589 252 -584 280
rect -556 252 -508 280
rect -480 252 -432 280
rect -404 252 -356 280
rect -328 252 -280 280
rect -252 252 -204 280
rect -176 252 -128 280
rect -100 252 -52 280
rect -24 252 24 280
rect 52 252 100 280
rect 128 252 176 280
rect 204 252 252 280
rect 280 252 328 280
rect 356 252 404 280
rect 432 252 480 280
rect 508 252 556 280
rect 584 252 589 280
rect -589 204 589 252
rect -589 176 -584 204
rect -556 176 -508 204
rect -480 176 -432 204
rect -404 176 -356 204
rect -328 176 -280 204
rect -252 176 -204 204
rect -176 176 -128 204
rect -100 176 -52 204
rect -24 176 24 204
rect 52 176 100 204
rect 128 176 176 204
rect 204 176 252 204
rect 280 176 328 204
rect 356 176 404 204
rect 432 176 480 204
rect 508 176 556 204
rect 584 176 589 204
rect -589 128 589 176
rect -589 100 -584 128
rect -556 100 -508 128
rect -480 100 -432 128
rect -404 100 -356 128
rect -328 100 -280 128
rect -252 100 -204 128
rect -176 100 -128 128
rect -100 100 -52 128
rect -24 100 24 128
rect 52 100 100 128
rect 128 100 176 128
rect 204 100 252 128
rect 280 100 328 128
rect 356 100 404 128
rect 432 100 480 128
rect 508 100 556 128
rect 584 100 589 128
rect -589 52 589 100
rect -589 24 -584 52
rect -556 24 -508 52
rect -480 24 -432 52
rect -404 24 -356 52
rect -328 24 -280 52
rect -252 24 -204 52
rect -176 24 -128 52
rect -100 24 -52 52
rect -24 24 24 52
rect 52 24 100 52
rect 128 24 176 52
rect 204 24 252 52
rect 280 24 328 52
rect 356 24 404 52
rect 432 24 480 52
rect 508 24 556 52
rect 584 24 589 52
rect -589 -24 589 24
rect -589 -52 -584 -24
rect -556 -52 -508 -24
rect -480 -52 -432 -24
rect -404 -52 -356 -24
rect -328 -52 -280 -24
rect -252 -52 -204 -24
rect -176 -52 -128 -24
rect -100 -52 -52 -24
rect -24 -52 24 -24
rect 52 -52 100 -24
rect 128 -52 176 -24
rect 204 -52 252 -24
rect 280 -52 328 -24
rect 356 -52 404 -24
rect 432 -52 480 -24
rect 508 -52 556 -24
rect 584 -52 589 -24
rect -589 -100 589 -52
rect -589 -128 -584 -100
rect -556 -128 -508 -100
rect -480 -128 -432 -100
rect -404 -128 -356 -100
rect -328 -128 -280 -100
rect -252 -128 -204 -100
rect -176 -128 -128 -100
rect -100 -128 -52 -100
rect -24 -128 24 -100
rect 52 -128 100 -100
rect 128 -128 176 -100
rect 204 -128 252 -100
rect 280 -128 328 -100
rect 356 -128 404 -100
rect 432 -128 480 -100
rect 508 -128 556 -100
rect 584 -128 589 -100
rect -589 -176 589 -128
rect -589 -204 -584 -176
rect -556 -204 -508 -176
rect -480 -204 -432 -176
rect -404 -204 -356 -176
rect -328 -204 -280 -176
rect -252 -204 -204 -176
rect -176 -204 -128 -176
rect -100 -204 -52 -176
rect -24 -204 24 -176
rect 52 -204 100 -176
rect 128 -204 176 -176
rect 204 -204 252 -176
rect 280 -204 328 -176
rect 356 -204 404 -176
rect 432 -204 480 -176
rect 508 -204 556 -176
rect 584 -204 589 -176
rect -589 -252 589 -204
rect -589 -280 -584 -252
rect -556 -280 -508 -252
rect -480 -280 -432 -252
rect -404 -280 -356 -252
rect -328 -280 -280 -252
rect -252 -280 -204 -252
rect -176 -280 -128 -252
rect -100 -280 -52 -252
rect -24 -280 24 -252
rect 52 -280 100 -252
rect 128 -280 176 -252
rect 204 -280 252 -252
rect 280 -280 328 -252
rect 356 -280 404 -252
rect 432 -280 480 -252
rect 508 -280 556 -252
rect 584 -280 589 -252
rect -589 -285 589 -280
<< via2 >>
rect -584 252 -556 280
rect -508 252 -480 280
rect -432 252 -404 280
rect -356 252 -328 280
rect -280 252 -252 280
rect -204 252 -176 280
rect -128 252 -100 280
rect -52 252 -24 280
rect 24 252 52 280
rect 100 252 128 280
rect 176 252 204 280
rect 252 252 280 280
rect 328 252 356 280
rect 404 252 432 280
rect 480 252 508 280
rect 556 252 584 280
rect -584 176 -556 204
rect -508 176 -480 204
rect -432 176 -404 204
rect -356 176 -328 204
rect -280 176 -252 204
rect -204 176 -176 204
rect -128 176 -100 204
rect -52 176 -24 204
rect 24 176 52 204
rect 100 176 128 204
rect 176 176 204 204
rect 252 176 280 204
rect 328 176 356 204
rect 404 176 432 204
rect 480 176 508 204
rect 556 176 584 204
rect -584 100 -556 128
rect -508 100 -480 128
rect -432 100 -404 128
rect -356 100 -328 128
rect -280 100 -252 128
rect -204 100 -176 128
rect -128 100 -100 128
rect -52 100 -24 128
rect 24 100 52 128
rect 100 100 128 128
rect 176 100 204 128
rect 252 100 280 128
rect 328 100 356 128
rect 404 100 432 128
rect 480 100 508 128
rect 556 100 584 128
rect -584 24 -556 52
rect -508 24 -480 52
rect -432 24 -404 52
rect -356 24 -328 52
rect -280 24 -252 52
rect -204 24 -176 52
rect -128 24 -100 52
rect -52 24 -24 52
rect 24 24 52 52
rect 100 24 128 52
rect 176 24 204 52
rect 252 24 280 52
rect 328 24 356 52
rect 404 24 432 52
rect 480 24 508 52
rect 556 24 584 52
rect -584 -52 -556 -24
rect -508 -52 -480 -24
rect -432 -52 -404 -24
rect -356 -52 -328 -24
rect -280 -52 -252 -24
rect -204 -52 -176 -24
rect -128 -52 -100 -24
rect -52 -52 -24 -24
rect 24 -52 52 -24
rect 100 -52 128 -24
rect 176 -52 204 -24
rect 252 -52 280 -24
rect 328 -52 356 -24
rect 404 -52 432 -24
rect 480 -52 508 -24
rect 556 -52 584 -24
rect -584 -128 -556 -100
rect -508 -128 -480 -100
rect -432 -128 -404 -100
rect -356 -128 -328 -100
rect -280 -128 -252 -100
rect -204 -128 -176 -100
rect -128 -128 -100 -100
rect -52 -128 -24 -100
rect 24 -128 52 -100
rect 100 -128 128 -100
rect 176 -128 204 -100
rect 252 -128 280 -100
rect 328 -128 356 -100
rect 404 -128 432 -100
rect 480 -128 508 -100
rect 556 -128 584 -100
rect -584 -204 -556 -176
rect -508 -204 -480 -176
rect -432 -204 -404 -176
rect -356 -204 -328 -176
rect -280 -204 -252 -176
rect -204 -204 -176 -176
rect -128 -204 -100 -176
rect -52 -204 -24 -176
rect 24 -204 52 -176
rect 100 -204 128 -176
rect 176 -204 204 -176
rect 252 -204 280 -176
rect 328 -204 356 -176
rect 404 -204 432 -176
rect 480 -204 508 -176
rect 556 -204 584 -176
rect -584 -280 -556 -252
rect -508 -280 -480 -252
rect -432 -280 -404 -252
rect -356 -280 -328 -252
rect -280 -280 -252 -252
rect -204 -280 -176 -252
rect -128 -280 -100 -252
rect -52 -280 -24 -252
rect 24 -280 52 -252
rect 100 -280 128 -252
rect 176 -280 204 -252
rect 252 -280 280 -252
rect 328 -280 356 -252
rect 404 -280 432 -252
rect 480 -280 508 -252
rect 556 -280 584 -252
<< metal3 >>
rect -589 280 589 285
rect -589 252 -584 280
rect -556 252 -508 280
rect -480 252 -432 280
rect -404 252 -356 280
rect -328 252 -280 280
rect -252 252 -204 280
rect -176 252 -128 280
rect -100 252 -52 280
rect -24 252 24 280
rect 52 252 100 280
rect 128 252 176 280
rect 204 252 252 280
rect 280 252 328 280
rect 356 252 404 280
rect 432 252 480 280
rect 508 252 556 280
rect 584 252 589 280
rect -589 204 589 252
rect -589 176 -584 204
rect -556 176 -508 204
rect -480 176 -432 204
rect -404 176 -356 204
rect -328 176 -280 204
rect -252 176 -204 204
rect -176 176 -128 204
rect -100 176 -52 204
rect -24 176 24 204
rect 52 176 100 204
rect 128 176 176 204
rect 204 176 252 204
rect 280 176 328 204
rect 356 176 404 204
rect 432 176 480 204
rect 508 176 556 204
rect 584 176 589 204
rect -589 128 589 176
rect -589 100 -584 128
rect -556 100 -508 128
rect -480 100 -432 128
rect -404 100 -356 128
rect -328 100 -280 128
rect -252 100 -204 128
rect -176 100 -128 128
rect -100 100 -52 128
rect -24 100 24 128
rect 52 100 100 128
rect 128 100 176 128
rect 204 100 252 128
rect 280 100 328 128
rect 356 100 404 128
rect 432 100 480 128
rect 508 100 556 128
rect 584 100 589 128
rect -589 52 589 100
rect -589 24 -584 52
rect -556 24 -508 52
rect -480 24 -432 52
rect -404 24 -356 52
rect -328 24 -280 52
rect -252 24 -204 52
rect -176 24 -128 52
rect -100 24 -52 52
rect -24 24 24 52
rect 52 24 100 52
rect 128 24 176 52
rect 204 24 252 52
rect 280 24 328 52
rect 356 24 404 52
rect 432 24 480 52
rect 508 24 556 52
rect 584 24 589 52
rect -589 -24 589 24
rect -589 -52 -584 -24
rect -556 -52 -508 -24
rect -480 -52 -432 -24
rect -404 -52 -356 -24
rect -328 -52 -280 -24
rect -252 -52 -204 -24
rect -176 -52 -128 -24
rect -100 -52 -52 -24
rect -24 -52 24 -24
rect 52 -52 100 -24
rect 128 -52 176 -24
rect 204 -52 252 -24
rect 280 -52 328 -24
rect 356 -52 404 -24
rect 432 -52 480 -24
rect 508 -52 556 -24
rect 584 -52 589 -24
rect -589 -100 589 -52
rect -589 -128 -584 -100
rect -556 -128 -508 -100
rect -480 -128 -432 -100
rect -404 -128 -356 -100
rect -328 -128 -280 -100
rect -252 -128 -204 -100
rect -176 -128 -128 -100
rect -100 -128 -52 -100
rect -24 -128 24 -100
rect 52 -128 100 -100
rect 128 -128 176 -100
rect 204 -128 252 -100
rect 280 -128 328 -100
rect 356 -128 404 -100
rect 432 -128 480 -100
rect 508 -128 556 -100
rect 584 -128 589 -100
rect -589 -176 589 -128
rect -589 -204 -584 -176
rect -556 -204 -508 -176
rect -480 -204 -432 -176
rect -404 -204 -356 -176
rect -328 -204 -280 -176
rect -252 -204 -204 -176
rect -176 -204 -128 -176
rect -100 -204 -52 -176
rect -24 -204 24 -176
rect 52 -204 100 -176
rect 128 -204 176 -176
rect 204 -204 252 -176
rect 280 -204 328 -176
rect 356 -204 404 -176
rect 432 -204 480 -176
rect 508 -204 556 -176
rect 584 -204 589 -176
rect -589 -252 589 -204
rect -589 -280 -584 -252
rect -556 -280 -508 -252
rect -480 -280 -432 -252
rect -404 -280 -356 -252
rect -328 -280 -280 -252
rect -252 -280 -204 -252
rect -176 -280 -128 -252
rect -100 -280 -52 -252
rect -24 -280 24 -252
rect 52 -280 100 -252
rect 128 -280 176 -252
rect 204 -280 252 -252
rect 280 -280 328 -252
rect 356 -280 404 -252
rect 432 -280 480 -252
rect 508 -280 556 -252
rect 584 -280 589 -252
rect -589 -285 589 -280
<< end >>
