magic
tech gf180mcuC
magscale 1 10
timestamp 1692948427
<< nwell >>
rect -3356 -2050 -1223 1494
<< nsubdiff >>
rect -3309 1441 -1257 1456
rect -3309 1394 -3294 1441
rect -3247 1395 -3199 1441
rect -3153 1395 -3105 1441
rect -3059 1395 -3011 1441
rect -2965 1395 -2917 1441
rect -2871 1395 -2823 1441
rect -2777 1395 -2729 1441
rect -2683 1395 -2635 1441
rect -2589 1395 -2541 1441
rect -2495 1395 -2447 1441
rect -2401 1395 -2353 1441
rect -2307 1395 -2259 1441
rect -2213 1395 -2165 1441
rect -2119 1395 -2071 1441
rect -2025 1395 -1977 1441
rect -1931 1395 -1883 1441
rect -1837 1395 -1789 1441
rect -1743 1395 -1695 1441
rect -1649 1395 -1601 1441
rect -1555 1395 -1507 1441
rect -1461 1395 -1413 1441
rect -1367 1395 -1319 1441
rect -3247 1394 -1319 1395
rect -1272 1394 -1257 1441
rect -3309 1380 -1257 1394
rect -3309 1346 -3233 1380
rect -3309 1300 -3294 1346
rect -3248 1300 -3233 1346
rect -3309 1252 -3233 1300
rect -1333 1346 -1257 1380
rect -1333 1300 -1318 1346
rect -1272 1300 -1257 1346
rect -3309 1206 -3294 1252
rect -3248 1206 -3233 1252
rect -3309 1158 -3233 1206
rect -1333 1252 -1257 1300
rect -1333 1206 -1318 1252
rect -1272 1206 -1257 1252
rect -3309 1112 -3294 1158
rect -3248 1112 -3233 1158
rect -3309 1064 -3233 1112
rect -3309 1018 -3294 1064
rect -3248 1018 -3233 1064
rect -3309 970 -3233 1018
rect -3309 924 -3294 970
rect -3248 924 -3233 970
rect -3309 876 -3233 924
rect -3309 830 -3294 876
rect -3248 830 -3233 876
rect -3309 782 -3233 830
rect -3309 736 -3294 782
rect -3248 736 -3233 782
rect -3309 688 -3233 736
rect -3309 642 -3294 688
rect -3248 642 -3233 688
rect -3309 594 -3233 642
rect -3309 548 -3294 594
rect -3248 548 -3233 594
rect -3309 500 -3233 548
rect -1333 1158 -1257 1206
rect -1333 1112 -1318 1158
rect -1272 1112 -1257 1158
rect -1333 1064 -1257 1112
rect -1333 1018 -1318 1064
rect -1272 1018 -1257 1064
rect -1333 970 -1257 1018
rect -1333 924 -1318 970
rect -1272 924 -1257 970
rect -1333 876 -1257 924
rect -1333 830 -1318 876
rect -1272 830 -1257 876
rect -1333 782 -1257 830
rect -1333 736 -1318 782
rect -1272 736 -1257 782
rect -1333 688 -1257 736
rect -1333 642 -1318 688
rect -1272 642 -1257 688
rect -1333 594 -1257 642
rect -1333 548 -1318 594
rect -1272 548 -1257 594
rect -3309 454 -3294 500
rect -3248 454 -3233 500
rect -1333 500 -1257 548
rect -3309 406 -3233 454
rect -1333 454 -1318 500
rect -1272 454 -1257 500
rect -3309 360 -3294 406
rect -3248 360 -3233 406
rect -3309 312 -3233 360
rect -3309 266 -3294 312
rect -3248 266 -3233 312
rect -3309 218 -3233 266
rect -3309 172 -3294 218
rect -3248 172 -3233 218
rect -3309 124 -3233 172
rect -3309 78 -3294 124
rect -3248 78 -3233 124
rect -3309 30 -3233 78
rect -3309 -16 -3294 30
rect -3248 -16 -3233 30
rect -3309 -64 -3233 -16
rect -3309 -110 -3294 -64
rect -3248 -110 -3233 -64
rect -3309 -158 -3233 -110
rect -3309 -204 -3294 -158
rect -3248 -204 -3233 -158
rect -3309 -252 -3233 -204
rect -1333 406 -1257 454
rect -1333 360 -1318 406
rect -1272 360 -1257 406
rect -1333 312 -1257 360
rect -1333 266 -1318 312
rect -1272 266 -1257 312
rect -1333 218 -1257 266
rect -1333 172 -1318 218
rect -1272 172 -1257 218
rect -1333 124 -1257 172
rect -1333 78 -1318 124
rect -1272 78 -1257 124
rect -1333 30 -1257 78
rect -1333 -16 -1318 30
rect -1272 -16 -1257 30
rect -1333 -64 -1257 -16
rect -1333 -110 -1318 -64
rect -1272 -110 -1257 -64
rect -1333 -158 -1257 -110
rect -1333 -204 -1318 -158
rect -1272 -204 -1257 -158
rect -3309 -298 -3294 -252
rect -3248 -298 -3233 -252
rect -1333 -252 -1257 -204
rect -3309 -346 -3233 -298
rect -3309 -392 -3294 -346
rect -3248 -392 -3233 -346
rect -3309 -440 -3233 -392
rect -3309 -486 -3294 -440
rect -3248 -486 -3233 -440
rect -3309 -534 -3233 -486
rect -3309 -580 -3294 -534
rect -3248 -580 -3233 -534
rect -3309 -628 -3233 -580
rect -3309 -674 -3294 -628
rect -3248 -674 -3233 -628
rect -3309 -722 -3233 -674
rect -3309 -768 -3294 -722
rect -3248 -768 -3233 -722
rect -3309 -816 -3233 -768
rect -3309 -862 -3294 -816
rect -3248 -862 -3233 -816
rect -3309 -910 -3233 -862
rect -3309 -956 -3294 -910
rect -3248 -956 -3233 -910
rect -1333 -298 -1318 -252
rect -1272 -298 -1257 -252
rect -1333 -346 -1257 -298
rect -1333 -392 -1318 -346
rect -1272 -392 -1257 -346
rect -1333 -440 -1257 -392
rect -1333 -486 -1318 -440
rect -1272 -486 -1257 -440
rect -1333 -534 -1257 -486
rect -1333 -580 -1318 -534
rect -1272 -580 -1257 -534
rect -1333 -628 -1257 -580
rect -1333 -674 -1318 -628
rect -1272 -674 -1257 -628
rect -1333 -722 -1257 -674
rect -1333 -768 -1318 -722
rect -1272 -768 -1257 -722
rect -1333 -816 -1257 -768
rect -1333 -862 -1318 -816
rect -1272 -862 -1257 -816
rect -1333 -910 -1257 -862
rect -3309 -1004 -3233 -956
rect -3309 -1050 -3294 -1004
rect -3248 -1050 -3233 -1004
rect -1333 -956 -1318 -910
rect -1272 -956 -1257 -910
rect -1333 -1004 -1257 -956
rect -3309 -1098 -3233 -1050
rect -3309 -1144 -3294 -1098
rect -3248 -1144 -3233 -1098
rect -3309 -1192 -3233 -1144
rect -3309 -1238 -3294 -1192
rect -3248 -1238 -3233 -1192
rect -3309 -1286 -3233 -1238
rect -3309 -1332 -3294 -1286
rect -3248 -1332 -3233 -1286
rect -3309 -1380 -3233 -1332
rect -3309 -1426 -3294 -1380
rect -3248 -1426 -3233 -1380
rect -3309 -1474 -3233 -1426
rect -3309 -1520 -3294 -1474
rect -3248 -1520 -3233 -1474
rect -3309 -1568 -3233 -1520
rect -3309 -1614 -3294 -1568
rect -3248 -1614 -3233 -1568
rect -3309 -1662 -3233 -1614
rect -3309 -1708 -3294 -1662
rect -3248 -1708 -3233 -1662
rect -3309 -1756 -3233 -1708
rect -3309 -1802 -3294 -1756
rect -3248 -1802 -3233 -1756
rect -3309 -1850 -3233 -1802
rect -3309 -1896 -3294 -1850
rect -3248 -1896 -3233 -1850
rect -3309 -1929 -3233 -1896
rect -1333 -1050 -1318 -1004
rect -1272 -1050 -1257 -1004
rect -1333 -1098 -1257 -1050
rect -1333 -1144 -1318 -1098
rect -1272 -1144 -1257 -1098
rect -1333 -1192 -1257 -1144
rect -1333 -1238 -1318 -1192
rect -1272 -1238 -1257 -1192
rect -1333 -1286 -1257 -1238
rect -1333 -1332 -1318 -1286
rect -1272 -1332 -1257 -1286
rect -1333 -1380 -1257 -1332
rect -1333 -1426 -1318 -1380
rect -1272 -1426 -1257 -1380
rect -1333 -1474 -1257 -1426
rect -1333 -1520 -1318 -1474
rect -1272 -1520 -1257 -1474
rect -1333 -1568 -1257 -1520
rect -1333 -1614 -1318 -1568
rect -1272 -1614 -1257 -1568
rect -1333 -1662 -1257 -1614
rect -1333 -1708 -1318 -1662
rect -1272 -1708 -1257 -1662
rect -1333 -1756 -1257 -1708
rect -1333 -1802 -1318 -1756
rect -1272 -1802 -1257 -1756
rect -1333 -1850 -1257 -1802
rect -1333 -1896 -1318 -1850
rect -1272 -1896 -1257 -1850
rect -1333 -1929 -1257 -1896
rect -3309 -1944 -1257 -1929
rect -3309 -1990 -3293 -1944
rect -3247 -1990 -3199 -1944
rect -3153 -1990 -3105 -1944
rect -3059 -1990 -3011 -1944
rect -2965 -1990 -2917 -1944
rect -2871 -1990 -2823 -1944
rect -2777 -1990 -2729 -1944
rect -2683 -1990 -2635 -1944
rect -2589 -1990 -2541 -1944
rect -2495 -1990 -2447 -1944
rect -2401 -1990 -2353 -1944
rect -2307 -1990 -2259 -1944
rect -2213 -1990 -2165 -1944
rect -2119 -1990 -2071 -1944
rect -2025 -1990 -1977 -1944
rect -1931 -1990 -1883 -1944
rect -1837 -1990 -1789 -1944
rect -1743 -1990 -1695 -1944
rect -1649 -1990 -1601 -1944
rect -1555 -1990 -1507 -1944
rect -1461 -1990 -1413 -1944
rect -1367 -1990 -1319 -1944
rect -1273 -1990 -1257 -1944
rect -3309 -2005 -1257 -1990
<< nsubdiffcont >>
rect -3294 1394 -3247 1441
rect -3199 1395 -3153 1441
rect -3105 1395 -3059 1441
rect -3011 1395 -2965 1441
rect -2917 1395 -2871 1441
rect -2823 1395 -2777 1441
rect -2729 1395 -2683 1441
rect -2635 1395 -2589 1441
rect -2541 1395 -2495 1441
rect -2447 1395 -2401 1441
rect -2353 1395 -2307 1441
rect -2259 1395 -2213 1441
rect -2165 1395 -2119 1441
rect -2071 1395 -2025 1441
rect -1977 1395 -1931 1441
rect -1883 1395 -1837 1441
rect -1789 1395 -1743 1441
rect -1695 1395 -1649 1441
rect -1601 1395 -1555 1441
rect -1507 1395 -1461 1441
rect -1413 1395 -1367 1441
rect -1319 1394 -1272 1441
rect -3294 1300 -3248 1346
rect -1318 1300 -1272 1346
rect -3294 1206 -3248 1252
rect -1318 1206 -1272 1252
rect -3294 1112 -3248 1158
rect -3294 1018 -3248 1064
rect -3294 924 -3248 970
rect -3294 830 -3248 876
rect -3294 736 -3248 782
rect -3294 642 -3248 688
rect -3294 548 -3248 594
rect -1318 1112 -1272 1158
rect -1318 1018 -1272 1064
rect -1318 924 -1272 970
rect -1318 830 -1272 876
rect -1318 736 -1272 782
rect -1318 642 -1272 688
rect -1318 548 -1272 594
rect -3294 454 -3248 500
rect -1318 454 -1272 500
rect -3294 360 -3248 406
rect -3294 266 -3248 312
rect -3294 172 -3248 218
rect -3294 78 -3248 124
rect -3294 -16 -3248 30
rect -3294 -110 -3248 -64
rect -3294 -204 -3248 -158
rect -1318 360 -1272 406
rect -1318 266 -1272 312
rect -1318 172 -1272 218
rect -1318 78 -1272 124
rect -1318 -16 -1272 30
rect -1318 -110 -1272 -64
rect -1318 -204 -1272 -158
rect -3294 -298 -3248 -252
rect -3294 -392 -3248 -346
rect -3294 -486 -3248 -440
rect -3294 -580 -3248 -534
rect -3294 -674 -3248 -628
rect -3294 -768 -3248 -722
rect -3294 -862 -3248 -816
rect -3294 -956 -3248 -910
rect -1318 -298 -1272 -252
rect -1318 -392 -1272 -346
rect -1318 -486 -1272 -440
rect -1318 -580 -1272 -534
rect -1318 -674 -1272 -628
rect -1318 -768 -1272 -722
rect -1318 -862 -1272 -816
rect -3294 -1050 -3248 -1004
rect -1318 -956 -1272 -910
rect -3294 -1144 -3248 -1098
rect -3294 -1238 -3248 -1192
rect -3294 -1332 -3248 -1286
rect -3294 -1426 -3248 -1380
rect -3294 -1520 -3248 -1474
rect -3294 -1614 -3248 -1568
rect -3294 -1708 -3248 -1662
rect -3294 -1802 -3248 -1756
rect -3294 -1896 -3248 -1850
rect -1318 -1050 -1272 -1004
rect -1318 -1144 -1272 -1098
rect -1318 -1238 -1272 -1192
rect -1318 -1332 -1272 -1286
rect -1318 -1426 -1272 -1380
rect -1318 -1520 -1272 -1474
rect -1318 -1614 -1272 -1568
rect -1318 -1708 -1272 -1662
rect -1318 -1802 -1272 -1756
rect -1318 -1896 -1272 -1850
rect -3293 -1990 -3247 -1944
rect -3199 -1990 -3153 -1944
rect -3105 -1990 -3059 -1944
rect -3011 -1990 -2965 -1944
rect -2917 -1990 -2871 -1944
rect -2823 -1990 -2777 -1944
rect -2729 -1990 -2683 -1944
rect -2635 -1990 -2589 -1944
rect -2541 -1990 -2495 -1944
rect -2447 -1990 -2401 -1944
rect -2353 -1990 -2307 -1944
rect -2259 -1990 -2213 -1944
rect -2165 -1990 -2119 -1944
rect -2071 -1990 -2025 -1944
rect -1977 -1990 -1931 -1944
rect -1883 -1990 -1837 -1944
rect -1789 -1990 -1743 -1944
rect -1695 -1990 -1649 -1944
rect -1601 -1990 -1555 -1944
rect -1507 -1990 -1461 -1944
rect -1413 -1990 -1367 -1944
rect -1319 -1990 -1273 -1944
<< polysilicon >>
rect -2679 1260 -1919 1276
rect -2679 1214 -2323 1260
rect -2277 1214 -1919 1260
rect -2679 1192 -1919 1214
rect -2679 507 -1919 517
rect -2895 504 -2783 505
rect -2895 458 -2864 504
rect -2818 458 -2783 504
rect -2895 457 -2783 458
rect -2679 461 -2428 507
rect -2382 504 -1919 507
rect -2382 461 -2215 504
rect -2679 457 -2215 461
rect -2167 457 -1919 504
rect -1815 504 -1703 505
rect -1815 458 -1782 504
rect -1736 458 -1703 504
rect -1815 457 -1703 458
rect -2679 444 -1919 457
rect -2895 -232 -2783 -231
rect -2895 -278 -2864 -232
rect -2818 -278 -2783 -232
rect -2895 -279 -2783 -278
rect -2679 -232 -1919 -219
rect -2679 -278 -2428 -232
rect -2382 -278 -2215 -232
rect -2679 -279 -2215 -278
rect -2167 -279 -1919 -232
rect -1815 -232 -1703 -231
rect -1815 -278 -1781 -232
rect -1735 -278 -1703 -232
rect -1815 -279 -1703 -278
rect -2679 -292 -1919 -279
rect -2895 -968 -2783 -967
rect -2895 -1014 -2863 -968
rect -2817 -1014 -2783 -968
rect -2895 -1015 -2783 -1014
rect -2679 -970 -1919 -955
rect -2679 -971 -2215 -970
rect -2679 -1017 -2428 -971
rect -2382 -1017 -2215 -971
rect -2167 -1017 -1919 -970
rect -1815 -968 -1703 -967
rect -1815 -1014 -1781 -968
rect -1735 -1014 -1703 -968
rect -1815 -1015 -1703 -1014
rect -2679 -1028 -1919 -1017
<< polycontact >>
rect -2323 1214 -2277 1260
rect -2864 458 -2818 504
rect -2428 461 -2382 507
rect -2215 457 -2167 504
rect -1782 458 -1736 504
rect -2864 -278 -2818 -232
rect -2428 -278 -2382 -232
rect -2215 -279 -2167 -232
rect -1781 -278 -1735 -232
rect -2863 -1014 -2817 -968
rect -2428 -1017 -2382 -971
rect -2215 -1017 -2167 -970
rect -1781 -1014 -1735 -968
<< metal1 >>
rect -3320 1441 -1246 1467
rect -3320 1394 -3294 1441
rect -3247 1395 -3199 1441
rect -3153 1395 -3105 1441
rect -3059 1395 -3011 1441
rect -2965 1395 -2917 1441
rect -2871 1395 -2823 1441
rect -2777 1395 -2729 1441
rect -2683 1395 -2635 1441
rect -2589 1395 -2541 1441
rect -2495 1395 -2447 1441
rect -2401 1395 -2353 1441
rect -2307 1395 -2259 1441
rect -2213 1395 -2165 1441
rect -2119 1395 -2071 1441
rect -2025 1395 -1977 1441
rect -1931 1395 -1883 1441
rect -1837 1395 -1789 1441
rect -1743 1395 -1695 1441
rect -1649 1395 -1601 1441
rect -1555 1395 -1507 1441
rect -1461 1395 -1413 1441
rect -1367 1395 -1319 1441
rect -3247 1394 -1319 1395
rect -1272 1394 -1246 1441
rect -3320 1369 -1246 1394
rect -3320 1346 -3222 1369
rect -3320 1300 -3294 1346
rect -3248 1300 -3222 1346
rect -3320 1252 -3222 1300
rect -3320 1206 -3294 1252
rect -3248 1206 -3222 1252
rect -3320 1158 -3222 1206
rect -3320 1112 -3294 1158
rect -3248 1112 -3222 1158
rect -3320 1064 -3222 1112
rect -3320 1018 -3294 1064
rect -3248 1018 -3222 1064
rect -3320 970 -3222 1018
rect -3320 924 -3294 970
rect -3248 924 -3222 970
rect -3320 876 -3222 924
rect -3320 830 -3294 876
rect -3248 830 -3222 876
rect -3320 782 -3222 830
rect -3320 736 -3294 782
rect -3248 736 -3222 782
rect -3320 688 -3222 736
rect -3320 642 -3294 688
rect -3248 642 -3222 688
rect -3320 594 -3222 642
rect -3320 548 -3294 594
rect -3248 548 -3222 594
rect -3320 500 -3222 548
rect -3320 454 -3294 500
rect -3248 454 -3222 500
rect -3320 406 -3222 454
rect -3320 360 -3294 406
rect -3248 360 -3222 406
rect -3320 312 -3222 360
rect -3320 266 -3294 312
rect -3248 266 -3222 312
rect -3320 218 -3222 266
rect -3320 172 -3294 218
rect -3248 172 -3222 218
rect -3320 124 -3222 172
rect -3320 78 -3294 124
rect -3248 78 -3222 124
rect -3320 30 -3222 78
rect -3320 -16 -3294 30
rect -3248 -16 -3222 30
rect -3320 -64 -3222 -16
rect -3320 -110 -3294 -64
rect -3248 -110 -3222 -64
rect -3320 -158 -3222 -110
rect -3320 -204 -3294 -158
rect -3248 -204 -3222 -158
rect -3320 -252 -3222 -204
rect -3320 -298 -3294 -252
rect -3248 -298 -3222 -252
rect -3320 -346 -3222 -298
rect -3320 -392 -3294 -346
rect -3248 -392 -3222 -346
rect -3320 -440 -3222 -392
rect -3320 -486 -3294 -440
rect -3248 -486 -3222 -440
rect -3320 -534 -3222 -486
rect -3320 -580 -3294 -534
rect -3248 -580 -3222 -534
rect -3320 -628 -3222 -580
rect -3320 -674 -3294 -628
rect -3248 -674 -3222 -628
rect -3320 -722 -3222 -674
rect -3320 -768 -3294 -722
rect -3248 -768 -3222 -722
rect -3320 -816 -3222 -768
rect -3320 -862 -3294 -816
rect -3248 -862 -3222 -816
rect -3320 -910 -3222 -862
rect -3320 -956 -3294 -910
rect -3248 -956 -3222 -910
rect -3320 -1004 -3222 -956
rect -3320 -1050 -3294 -1004
rect -3248 -1050 -3222 -1004
rect -3320 -1098 -3222 -1050
rect -3320 -1144 -3294 -1098
rect -3248 -1144 -3222 -1098
rect -3320 -1192 -3222 -1144
rect -3320 -1238 -3294 -1192
rect -3248 -1238 -3222 -1192
rect -3320 -1286 -3222 -1238
rect -3320 -1332 -3294 -1286
rect -3248 -1332 -3222 -1286
rect -3320 -1380 -3222 -1332
rect -3320 -1426 -3294 -1380
rect -3248 -1426 -3222 -1380
rect -3320 -1474 -3222 -1426
rect -3320 -1520 -3294 -1474
rect -3248 -1520 -3222 -1474
rect -3320 -1568 -3222 -1520
rect -3320 -1614 -3294 -1568
rect -3248 -1614 -3222 -1568
rect -3320 -1662 -3222 -1614
rect -2973 508 -2921 1149
rect -2757 508 -2705 1150
rect -2973 504 -2705 508
rect -2973 458 -2864 504
rect -2818 458 -2705 504
rect -2973 454 -2705 458
rect -2973 -228 -2921 454
rect -2757 -228 -2705 454
rect -2973 -232 -2705 -228
rect -2973 -278 -2864 -232
rect -2818 -278 -2705 -232
rect -2973 -282 -2705 -278
rect -2973 -964 -2921 -282
rect -2757 -964 -2705 -282
rect -2973 -968 -2705 -964
rect -2973 -1014 -2863 -968
rect -2817 -1014 -2705 -968
rect -2973 -1018 -2705 -1014
rect -2973 -1660 -2921 -1018
rect -3320 -1708 -3294 -1662
rect -3248 -1708 -3222 -1662
rect -3320 -1756 -3222 -1708
rect -3320 -1802 -3294 -1756
rect -3248 -1802 -3222 -1756
rect -2757 -1764 -2705 -1018
rect -3320 -1850 -3222 -1802
rect -2773 -1774 -2689 -1764
rect -2773 -1828 -2758 -1774
rect -2704 -1828 -2689 -1774
rect -2773 -1842 -2689 -1828
rect -3320 -1896 -3294 -1850
rect -3248 -1896 -3222 -1850
rect -3320 -1918 -3222 -1896
rect -2541 -1918 -2489 1369
rect -2431 1289 -2312 1320
rect -2431 1229 -2402 1289
rect -2342 1281 -2312 1289
rect -2342 1260 -2165 1281
rect -2342 1229 -2323 1260
rect -2431 1214 -2323 1229
rect -2277 1214 -2165 1260
rect -2431 1201 -2165 1214
rect -2431 507 -2379 1201
rect -2431 461 -2428 507
rect -2382 461 -2379 507
rect -2431 -232 -2379 461
rect -2431 -278 -2428 -232
rect -2382 -278 -2379 -232
rect -2431 -971 -2379 -278
rect -2431 -1017 -2428 -971
rect -2382 -1017 -2379 -971
rect -2431 -1032 -2379 -1017
rect -2325 -1764 -2273 1150
rect -2217 504 -2165 1201
rect -2217 457 -2215 504
rect -2167 457 -2165 504
rect -2217 -232 -2165 457
rect -2217 -279 -2215 -232
rect -2167 -279 -2165 -232
rect -2217 -970 -2165 -279
rect -2217 -1017 -2215 -970
rect -2167 -1017 -2165 -970
rect -2217 -1032 -2165 -1017
rect -2343 -1774 -2259 -1764
rect -2343 -1828 -2326 -1774
rect -2272 -1828 -2259 -1774
rect -2343 -1842 -2259 -1828
rect -2109 -1918 -2057 1369
rect -1344 1346 -1246 1369
rect -1344 1300 -1318 1346
rect -1272 1300 -1246 1346
rect -1344 1252 -1246 1300
rect -1344 1206 -1318 1252
rect -1272 1206 -1246 1252
rect -1344 1158 -1246 1206
rect -1893 507 -1841 1150
rect -1677 507 -1625 1150
rect -1893 504 -1625 507
rect -1893 458 -1782 504
rect -1736 458 -1625 504
rect -1893 453 -1625 458
rect -1893 -228 -1841 453
rect -1677 -228 -1625 453
rect -1893 -232 -1625 -228
rect -1893 -278 -1781 -232
rect -1735 -278 -1625 -232
rect -1893 -282 -1625 -278
rect -1893 -964 -1841 -282
rect -1677 -964 -1625 -282
rect -1893 -968 -1625 -964
rect -1893 -1014 -1781 -968
rect -1735 -1014 -1625 -968
rect -1893 -1018 -1625 -1014
rect -1893 -1766 -1841 -1018
rect -1677 -1659 -1625 -1018
rect -1344 1112 -1318 1158
rect -1272 1112 -1246 1158
rect -1344 1064 -1246 1112
rect -1344 1018 -1318 1064
rect -1272 1018 -1246 1064
rect -1344 970 -1246 1018
rect -1344 924 -1318 970
rect -1272 924 -1246 970
rect -1344 876 -1246 924
rect -1344 830 -1318 876
rect -1272 845 -1246 876
rect -1272 830 -980 845
rect -1344 782 -980 830
rect -1344 736 -1318 782
rect -1272 736 -980 782
rect -1344 708 -980 736
rect -1344 688 -1246 708
rect -1344 642 -1318 688
rect -1272 642 -1246 688
rect -1344 594 -1246 642
rect -1344 548 -1318 594
rect -1272 548 -1246 594
rect -1344 500 -1246 548
rect -1344 454 -1318 500
rect -1272 454 -1246 500
rect -1344 406 -1246 454
rect -1344 360 -1318 406
rect -1272 360 -1246 406
rect -1344 312 -1246 360
rect -1344 266 -1318 312
rect -1272 266 -1246 312
rect -1344 218 -1246 266
rect -1344 172 -1318 218
rect -1272 172 -1246 218
rect -1344 124 -1246 172
rect -1344 78 -1318 124
rect -1272 78 -1246 124
rect -1344 58 -1246 78
rect -1344 30 -980 58
rect -1344 -16 -1318 30
rect -1272 -16 -980 30
rect -1344 -64 -980 -16
rect -1344 -110 -1318 -64
rect -1272 -79 -980 -64
rect -1272 -110 -1246 -79
rect -1344 -158 -1246 -110
rect -1344 -204 -1318 -158
rect -1272 -204 -1246 -158
rect -1344 -252 -1246 -204
rect -1344 -298 -1318 -252
rect -1272 -298 -1246 -252
rect -1344 -346 -1246 -298
rect -1344 -392 -1318 -346
rect -1272 -392 -1246 -346
rect -1344 -440 -1246 -392
rect -1344 -486 -1318 -440
rect -1272 -486 -1246 -440
rect -1344 -534 -1246 -486
rect -1344 -580 -1318 -534
rect -1272 -580 -1246 -534
rect -1344 -614 -1246 -580
rect -1344 -628 -980 -614
rect -1344 -674 -1318 -628
rect -1272 -674 -980 -628
rect -1344 -722 -980 -674
rect -1344 -768 -1318 -722
rect -1272 -751 -980 -722
rect -1272 -768 -1246 -751
rect -1344 -816 -1246 -768
rect -1344 -862 -1318 -816
rect -1272 -862 -1246 -816
rect -1344 -910 -1246 -862
rect -1344 -956 -1318 -910
rect -1272 -956 -1246 -910
rect -1344 -1004 -1246 -956
rect -1344 -1050 -1318 -1004
rect -1272 -1050 -1246 -1004
rect -1344 -1098 -1246 -1050
rect -1344 -1144 -1318 -1098
rect -1272 -1144 -1246 -1098
rect -1344 -1192 -1246 -1144
rect -1344 -1238 -1318 -1192
rect -1272 -1238 -1246 -1192
rect -1344 -1286 -980 -1238
rect -1344 -1332 -1318 -1286
rect -1272 -1332 -980 -1286
rect -1344 -1375 -980 -1332
rect -1344 -1380 -1246 -1375
rect -1344 -1426 -1318 -1380
rect -1272 -1426 -1246 -1380
rect -1344 -1474 -1246 -1426
rect -1344 -1520 -1318 -1474
rect -1272 -1520 -1246 -1474
rect -1344 -1568 -1246 -1520
rect -1344 -1614 -1318 -1568
rect -1272 -1614 -1246 -1568
rect -1344 -1662 -1246 -1614
rect -1344 -1708 -1318 -1662
rect -1272 -1708 -1246 -1662
rect -1344 -1756 -1246 -1708
rect -1909 -1777 -1825 -1766
rect -1909 -1831 -1894 -1777
rect -1840 -1831 -1825 -1777
rect -1909 -1844 -1825 -1831
rect -1344 -1802 -1318 -1756
rect -1272 -1802 -1246 -1756
rect -1344 -1813 -1246 -1802
rect -1344 -1850 -980 -1813
rect -1344 -1896 -1318 -1850
rect -1272 -1896 -980 -1850
rect -1344 -1918 -980 -1896
rect -3320 -1944 -980 -1918
rect -3320 -1990 -3293 -1944
rect -3247 -1990 -3199 -1944
rect -3153 -1990 -3105 -1944
rect -3059 -1990 -3011 -1944
rect -2965 -1990 -2917 -1944
rect -2871 -1990 -2823 -1944
rect -2777 -1990 -2729 -1944
rect -2683 -1990 -2635 -1944
rect -2589 -1990 -2541 -1944
rect -2495 -1990 -2447 -1944
rect -2401 -1990 -2353 -1944
rect -2307 -1990 -2259 -1944
rect -2213 -1990 -2165 -1944
rect -2119 -1990 -2071 -1944
rect -2025 -1990 -1977 -1944
rect -1931 -1990 -1883 -1944
rect -1837 -1990 -1789 -1944
rect -1743 -1990 -1695 -1944
rect -1649 -1990 -1601 -1944
rect -1555 -1990 -1507 -1944
rect -1461 -1990 -1413 -1944
rect -1367 -1990 -1319 -1944
rect -1273 -1950 -980 -1944
rect -1273 -1990 -1246 -1950
rect -3320 -2016 -1246 -1990
rect -3472 -2206 -1779 -2187
rect -3472 -2262 -3452 -2206
rect -3396 -2262 -3341 -2206
rect -3285 -2208 -1779 -2206
rect -3285 -2212 -2327 -2208
rect -3285 -2262 -2759 -2212
rect -3472 -2268 -2759 -2262
rect -2703 -2264 -2327 -2212
rect -2271 -2216 -1779 -2208
rect -2271 -2264 -1895 -2216
rect -2703 -2268 -1895 -2264
rect -3472 -2272 -1895 -2268
rect -1839 -2272 -1779 -2216
rect -3472 -2309 -1779 -2272
rect -3472 -2316 -3250 -2309
rect -3472 -2372 -3453 -2316
rect -3397 -2372 -3342 -2316
rect -3286 -2372 -3250 -2316
rect -3472 -2404 -3250 -2372
rect -1536 -2430 -1372 -2016
<< via1 >>
rect -2758 -1828 -2704 -1774
rect -2402 1229 -2342 1289
rect -2326 -1828 -2272 -1774
rect -1894 -1831 -1840 -1777
rect -3452 -2262 -3396 -2206
rect -3341 -2262 -3285 -2206
rect -2759 -2268 -2703 -2212
rect -2327 -2264 -2271 -2208
rect -1895 -2272 -1839 -2216
rect -3453 -2372 -3397 -2316
rect -3342 -2372 -3286 -2316
<< metal2 >>
rect -2407 1360 -1010 1442
rect -2407 1320 -2312 1360
rect -2431 1289 -2312 1320
rect -2431 1229 -2402 1289
rect -2342 1229 -2312 1289
rect -2431 1201 -2312 1229
rect -2773 -1774 -2689 -1764
rect -2773 -1828 -2758 -1774
rect -2704 -1828 -2689 -1774
rect -2773 -1842 -2689 -1828
rect -2343 -1774 -2259 -1764
rect -2343 -1828 -2326 -1774
rect -2272 -1828 -2259 -1774
rect -2343 -1842 -2259 -1828
rect -1909 -1777 -1825 -1766
rect -1909 -1831 -1894 -1777
rect -1840 -1831 -1825 -1777
rect -3472 -2206 -3250 -2187
rect -3472 -2262 -3452 -2206
rect -3396 -2262 -3341 -2206
rect -3285 -2262 -3250 -2206
rect -2759 -2207 -2703 -1842
rect -2327 -2201 -2271 -1842
rect -1909 -1844 -1825 -1831
rect -3472 -2316 -3250 -2262
rect -2773 -2212 -2689 -2207
rect -2773 -2268 -2759 -2212
rect -2703 -2268 -2689 -2212
rect -2773 -2285 -2689 -2268
rect -2341 -2208 -2257 -2201
rect -1895 -2208 -1839 -1844
rect -2341 -2264 -2327 -2208
rect -2271 -2264 -2257 -2208
rect -2341 -2279 -2257 -2264
rect -1909 -2216 -1825 -2208
rect -1909 -2272 -1895 -2216
rect -1839 -2272 -1825 -2216
rect -1909 -2286 -1825 -2272
rect -3472 -2372 -3453 -2316
rect -3397 -2372 -3342 -2316
rect -3286 -2372 -3250 -2316
rect -3472 -2404 -3250 -2372
rect -3472 -2430 -3352 -2404
use pmos_3p3_9BLZD7  pmos_3p3_9BLZD7_0
timestamp 1692615943
transform 1 0 -2299 0 1 -255
box -554 -1534 554 1534
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_16
timestamp 1692615943
transform 1 0 -2839 0 1 -1359
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_17
timestamp 1692615943
transform 1 0 -1759 0 1 -1359
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_18
timestamp 1692615943
transform 1 0 -2839 0 1 113
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_19
timestamp 1692615943
transform 1 0 -2839 0 1 -623
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_20
timestamp 1692615943
transform 1 0 -2839 0 1 849
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_21
timestamp 1692615943
transform 1 0 -1759 0 1 849
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_22
timestamp 1692615943
transform 1 0 -1759 0 1 113
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_23
timestamp 1692615943
transform 1 0 -1759 0 1 -623
box -230 -430 230 430
<< labels >>
flabel metal1 -1062 792 -1062 792 0 FreeSans 1600 0 0 0 VDD
port 0 nsew
<< end >>
