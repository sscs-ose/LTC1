magic
tech gf180mcuC
magscale 1 10
timestamp 1714558667
<< nwell >>
rect 568 2111 741 2148
rect 457 2077 851 2111
rect 1185 2081 1411 2113
rect 1749 2097 1976 2113
rect -42 2019 167 2065
rect 568 1993 741 2077
rect 1293 1993 1357 2081
rect 1796 2040 1976 2097
rect 1855 1993 1911 2040
rect -134 1833 -78 1834
rect -134 1832 -24 1833
rect -134 1830 -77 1832
rect -134 1815 -69 1818
rect -140 1777 -77 1782
rect 1621 1777 1735 1822
rect -144 1760 -79 1763
rect 1679 1759 1735 1777
rect -166 1721 368 1722
rect -166 1714 421 1721
rect -166 1674 899 1714
rect 980 1702 1116 1706
rect 1126 1703 1182 1706
rect 1690 1703 1756 1706
rect 2277 1700 2316 1702
rect 365 1657 899 1674
rect 429 1648 441 1657
rect 462 1648 611 1657
rect 1038 1649 1214 1651
rect 1126 1648 1182 1649
rect 1680 1648 1746 1651
rect 2302 1648 2316 1700
rect 2277 1646 2316 1648
rect 566 896 732 1051
rect 980 820 1038 901
rect 1291 896 1457 1051
rect 1891 991 2139 1017
rect 2015 896 2065 991
rect 1037 813 1038 820
rect 980 732 1047 813
rect 2403 636 2463 657
rect 2375 633 2463 636
rect 368 550 373 605
rect 422 550 425 618
rect 506 608 605 609
rect 506 606 573 608
rect 1230 606 1297 609
rect 506 605 582 606
rect 1230 605 1306 606
rect 506 602 573 605
rect 1164 596 1180 601
rect 366 539 425 550
rect 1125 551 1180 596
rect 1679 554 1833 609
rect 1843 606 1911 609
rect 2375 601 2460 633
rect 1230 551 1297 554
rect 1679 551 1901 554
rect 1125 549 1178 551
rect 1679 550 1833 551
<< pwell >>
rect -238 1398 186 1592
rect 408 1241 2365 1509
rect 402 144 2523 412
<< pdiff >>
rect 1037 810 1047 813
rect 983 808 1047 810
rect 981 799 1047 808
rect 983 795 1047 799
rect 1035 756 1047 795
rect 984 741 1047 756
rect 1037 737 1047 741
rect 1038 736 1047 737
<< psubdiff >>
rect -227 1296 -10 1377
rect -86 1194 -10 1296
rect -86 1181 165 1194
rect 446 1181 818 1194
rect 1146 1181 1385 1194
rect 1748 1181 1946 1194
rect -86 1118 2004 1181
rect 393 27 2161 97
rect 470 21 820 27
rect 1186 21 1536 27
rect 1904 21 2097 27
<< nsubdiff >>
rect 63 2104 915 2113
rect 1185 2104 1411 2113
rect 1749 2104 1976 2113
rect 63 2093 1976 2104
rect 63 2091 2013 2093
rect -168 2049 2013 2091
rect -168 2040 1976 2049
rect -168 2039 1803 2040
rect -168 2019 167 2039
rect 1891 1014 2139 1017
rect 393 942 2452 1014
<< polysilicon >>
rect 512 1697 603 1706
rect 581 1653 603 1697
rect 512 1650 603 1653
rect 368 550 373 605
<< metal1 >>
rect 568 2111 741 2148
rect 457 2077 851 2111
rect 1185 2081 1411 2113
rect 1749 2097 1976 2113
rect -42 2019 167 2065
rect 568 1993 741 2077
rect 1293 1993 1357 2081
rect 1796 2040 1976 2097
rect 1855 1993 1911 2040
rect 2272 1993 2581 2148
rect -380 1633 -350 1650
rect -390 1586 -337 1633
rect 512 1702 613 1703
rect 512 1697 524 1702
rect 576 1697 611 1702
rect 512 1651 524 1653
rect 512 1648 535 1651
rect 587 1648 611 1697
rect 86 1563 139 1610
rect 770 1599 812 1610
rect 1319 1599 1379 1610
rect 730 1544 816 1599
rect 1319 1596 1381 1599
rect 1326 1544 1381 1596
rect 1884 1544 1940 1610
rect 2344 1588 2401 1591
rect 2344 1586 2345 1588
rect 2333 1536 2345 1551
rect 2397 1586 2401 1588
rect 2408 1544 2449 1599
rect 2397 1536 2449 1544
rect 2333 1535 2449 1536
rect 2333 1514 2334 1535
rect -227 1297 -10 1377
rect -227 1296 13 1297
rect -150 1290 -41 1296
rect -21 1290 13 1296
rect -150 1283 13 1290
rect -150 1206 14 1283
rect -150 1097 64 1206
rect 569 1194 732 1206
rect 1287 1194 1302 1206
rect 1846 1194 1873 1206
rect 446 1173 818 1194
rect 1146 1173 1385 1194
rect 1748 1173 1946 1194
rect 569 1097 732 1173
rect 1287 1097 1302 1173
rect 1846 1097 1873 1173
rect -150 109 -41 1097
rect 566 896 732 1051
rect 1291 896 1457 1051
rect 2495 1050 2581 1993
rect 1891 991 2139 1017
rect 2015 896 2065 991
rect 2467 916 2581 1050
rect 980 801 1047 813
rect 980 749 984 801
rect 1036 749 1047 801
rect 980 732 1047 749
rect 506 605 518 606
rect 368 603 373 605
rect 368 551 371 603
rect 570 605 582 606
rect 1230 605 1242 606
rect 1164 596 1180 601
rect 1125 551 1180 596
rect 1294 605 1306 606
rect 368 550 373 551
rect 1125 549 1178 551
rect 80 466 133 513
rect 761 502 804 513
rect 1489 502 1528 513
rect 739 447 807 502
rect 1463 447 1535 502
rect 2036 447 2092 513
rect 2282 500 2289 512
rect 2282 453 2287 500
rect 2273 448 2287 453
rect 2339 448 2444 458
rect 2469 452 2524 499
rect 2273 447 2444 448
rect -150 106 2 109
rect -150 0 4 106
rect 561 40 724 109
rect 1285 40 1448 109
rect 470 21 820 40
rect 1186 21 1536 40
rect 2006 36 2038 109
rect 1904 21 2097 36
rect 561 0 724 21
rect 1285 0 1448 21
rect 2006 0 2038 21
<< via1 >>
rect -132 1780 -80 1832
rect -243 1600 -191 1652
rect 377 1651 429 1703
rect 535 1645 587 1697
rect 1127 1651 1179 1703
rect 1691 1651 1743 1703
rect 2251 1648 2303 1700
rect 1274 1544 1326 1596
rect 2345 1536 2397 1588
rect 984 749 1036 801
rect 371 551 423 603
rect 518 554 570 606
rect 1242 554 1294 606
rect 1845 554 1897 606
rect 2408 549 2460 601
rect 2287 448 2339 500
<< metal2 >>
rect -134 1833 -78 1834
rect -144 1832 1735 1833
rect -144 1780 -132 1832
rect -80 1780 1735 1832
rect -144 1777 1735 1780
rect -245 1714 421 1721
rect -245 1712 429 1714
rect -245 1703 441 1712
rect 1679 1706 1735 1777
rect -245 1664 377 1703
rect -245 1652 -188 1664
rect -245 1600 -243 1652
rect -191 1600 -188 1652
rect 365 1651 377 1664
rect 429 1651 441 1703
rect 980 1703 1191 1706
rect 365 1648 441 1651
rect 523 1698 589 1699
rect 523 1697 720 1698
rect -245 1587 -188 1600
rect 366 618 422 1648
rect 523 1645 535 1697
rect 587 1645 720 1697
rect 523 1642 720 1645
rect 366 603 425 618
rect 506 606 605 609
rect 366 551 371 603
rect 423 551 425 603
rect 366 539 425 551
rect 505 554 518 606
rect 570 554 605 606
rect 505 551 605 554
rect 505 268 562 551
rect 664 381 720 1642
rect 980 1651 1127 1703
rect 1179 1651 1191 1703
rect 980 1649 1191 1651
rect 1679 1703 1778 1706
rect 1679 1651 1691 1703
rect 1743 1651 1778 1703
rect 980 801 1038 1649
rect 1679 1648 1778 1651
rect 2221 1700 2316 1702
rect 2221 1648 2251 1700
rect 2303 1648 2316 1700
rect 1273 1600 1329 1608
rect 1272 1596 1329 1600
rect 1272 1544 1274 1596
rect 1326 1544 1329 1596
rect 1272 1542 1329 1544
rect 980 749 984 801
rect 1036 749 1038 801
rect 980 737 1038 749
rect 1273 609 1329 1542
rect 1230 606 1329 609
rect 1230 554 1242 606
rect 1294 554 1329 606
rect 1230 551 1329 554
rect 1679 609 1735 1648
rect 2221 1646 2316 1648
rect 1679 606 1932 609
rect 1679 554 1845 606
rect 1897 554 1932 606
rect 1679 551 1932 554
rect 1679 550 1833 551
rect 2221 544 2277 1646
rect 2333 1588 2410 1591
rect 2333 1536 2345 1588
rect 2397 1536 2410 1588
rect 2333 1514 2410 1536
rect 2354 657 2410 1514
rect 2354 601 2463 657
rect 2405 549 2408 601
rect 2460 549 2463 601
rect 2221 500 2341 544
rect 2221 488 2287 500
rect 2285 448 2287 488
rect 2339 448 2341 500
rect 2285 381 2341 448
rect 664 325 2341 381
rect 2405 268 2463 549
rect 505 210 2463 268
use GF_INV_MAG  GF_INV_MAG_0
timestamp 1714558667
transform 1 0 -272 0 1 1458
box -118 -175 286 666
use nand2_mag  nand2_mag_0
timestamp 1714137641
transform 1 0 1364 0 1 1285
box -70 -188 521 863
use nand2_mag  nand2_mag_1
timestamp 1714137641
transform 1 0 1928 0 1 1285
box -70 -188 521 863
use nand2_mag  nand2_mag_2
timestamp 1714137641
transform 1 0 800 0 1 1285
box -70 -188 521 863
use nand2_mag  nand2_mag_3
timestamp 1714137641
transform 1 0 1518 0 1 188
box -70 -188 521 863
use nand2_mag  nand2_mag_4
timestamp 1714137641
transform 1 0 2082 0 1 188
box -70 -188 521 863
use nand3_mag  nand3_mag_0
timestamp 1714137641
transform 1 0 76 0 1 1285
box -70 -188 671 863
use nand3_mag  nand3_mag_1
timestamp 1714137641
transform 1 0 794 0 1 188
box -70 -188 671 863
use nand3_mag  nand3_mag_2
timestamp 1714137641
transform 1 0 70 0 1 188
box -70 -188 671 863
<< labels >>
flabel metal1 650 2060 650 2060 0 FreeSans 320 0 0 0 VDD
port 1 nsew
flabel metal1 630 1130 630 1130 0 FreeSans 320 0 0 0 VSS
port 2 nsew
flabel metal1 -370 1610 -370 1610 0 FreeSans 320 0 0 0 CLK
port 3 nsew
flabel metal1 1170 570 1170 570 0 FreeSans 320 0 0 0 RST
port 6 nsew
flabel metal1 2485 473 2485 473 0 FreeSans 480 0 0 0 QB
port 8 nsew
flabel metal1 2430 1560 2430 1560 0 FreeSans 320 0 0 0 Q
port 7 nsew
flabel metal1 94 506 94 506 0 FreeSans 640 0 0 0 J
port 9 nsew
flabel metal1 104 1597 104 1597 0 FreeSans 640 0 0 0 K
port 10 nsew
<< end >>
