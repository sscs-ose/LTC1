magic
tech gf180mcuC
magscale 1 10
timestamp 1692680230
<< pwell >>
rect -1660 -536 1660 536
<< nmos >>
rect -1548 68 -1492 468
rect -1388 68 -1332 468
rect -1228 68 -1172 468
rect -1068 68 -1012 468
rect -908 68 -852 468
rect -748 68 -692 468
rect -588 68 -532 468
rect -428 68 -372 468
rect -268 68 -212 468
rect -108 68 -52 468
rect 52 68 108 468
rect 212 68 268 468
rect 372 68 428 468
rect 532 68 588 468
rect 692 68 748 468
rect 852 68 908 468
rect 1012 68 1068 468
rect 1172 68 1228 468
rect 1332 68 1388 468
rect 1492 68 1548 468
rect -1548 -468 -1492 -68
rect -1388 -468 -1332 -68
rect -1228 -468 -1172 -68
rect -1068 -468 -1012 -68
rect -908 -468 -852 -68
rect -748 -468 -692 -68
rect -588 -468 -532 -68
rect -428 -468 -372 -68
rect -268 -468 -212 -68
rect -108 -468 -52 -68
rect 52 -468 108 -68
rect 212 -468 268 -68
rect 372 -468 428 -68
rect 532 -468 588 -68
rect 692 -468 748 -68
rect 852 -468 908 -68
rect 1012 -468 1068 -68
rect 1172 -468 1228 -68
rect 1332 -468 1388 -68
rect 1492 -468 1548 -68
<< ndiff >>
rect -1636 455 -1548 468
rect -1636 81 -1623 455
rect -1577 81 -1548 455
rect -1636 68 -1548 81
rect -1492 455 -1388 468
rect -1492 81 -1463 455
rect -1417 81 -1388 455
rect -1492 68 -1388 81
rect -1332 455 -1228 468
rect -1332 81 -1303 455
rect -1257 81 -1228 455
rect -1332 68 -1228 81
rect -1172 455 -1068 468
rect -1172 81 -1143 455
rect -1097 81 -1068 455
rect -1172 68 -1068 81
rect -1012 455 -908 468
rect -1012 81 -983 455
rect -937 81 -908 455
rect -1012 68 -908 81
rect -852 455 -748 468
rect -852 81 -823 455
rect -777 81 -748 455
rect -852 68 -748 81
rect -692 455 -588 468
rect -692 81 -663 455
rect -617 81 -588 455
rect -692 68 -588 81
rect -532 455 -428 468
rect -532 81 -503 455
rect -457 81 -428 455
rect -532 68 -428 81
rect -372 455 -268 468
rect -372 81 -343 455
rect -297 81 -268 455
rect -372 68 -268 81
rect -212 455 -108 468
rect -212 81 -183 455
rect -137 81 -108 455
rect -212 68 -108 81
rect -52 455 52 468
rect -52 81 -23 455
rect 23 81 52 455
rect -52 68 52 81
rect 108 455 212 468
rect 108 81 137 455
rect 183 81 212 455
rect 108 68 212 81
rect 268 455 372 468
rect 268 81 297 455
rect 343 81 372 455
rect 268 68 372 81
rect 428 455 532 468
rect 428 81 457 455
rect 503 81 532 455
rect 428 68 532 81
rect 588 455 692 468
rect 588 81 617 455
rect 663 81 692 455
rect 588 68 692 81
rect 748 455 852 468
rect 748 81 777 455
rect 823 81 852 455
rect 748 68 852 81
rect 908 455 1012 468
rect 908 81 937 455
rect 983 81 1012 455
rect 908 68 1012 81
rect 1068 455 1172 468
rect 1068 81 1097 455
rect 1143 81 1172 455
rect 1068 68 1172 81
rect 1228 455 1332 468
rect 1228 81 1257 455
rect 1303 81 1332 455
rect 1228 68 1332 81
rect 1388 455 1492 468
rect 1388 81 1417 455
rect 1463 81 1492 455
rect 1388 68 1492 81
rect 1548 455 1636 468
rect 1548 81 1577 455
rect 1623 81 1636 455
rect 1548 68 1636 81
rect -1636 -81 -1548 -68
rect -1636 -455 -1623 -81
rect -1577 -455 -1548 -81
rect -1636 -468 -1548 -455
rect -1492 -81 -1388 -68
rect -1492 -455 -1463 -81
rect -1417 -455 -1388 -81
rect -1492 -468 -1388 -455
rect -1332 -81 -1228 -68
rect -1332 -455 -1303 -81
rect -1257 -455 -1228 -81
rect -1332 -468 -1228 -455
rect -1172 -81 -1068 -68
rect -1172 -455 -1143 -81
rect -1097 -455 -1068 -81
rect -1172 -468 -1068 -455
rect -1012 -81 -908 -68
rect -1012 -455 -983 -81
rect -937 -455 -908 -81
rect -1012 -468 -908 -455
rect -852 -81 -748 -68
rect -852 -455 -823 -81
rect -777 -455 -748 -81
rect -852 -468 -748 -455
rect -692 -81 -588 -68
rect -692 -455 -663 -81
rect -617 -455 -588 -81
rect -692 -468 -588 -455
rect -532 -81 -428 -68
rect -532 -455 -503 -81
rect -457 -455 -428 -81
rect -532 -468 -428 -455
rect -372 -81 -268 -68
rect -372 -455 -343 -81
rect -297 -455 -268 -81
rect -372 -468 -268 -455
rect -212 -81 -108 -68
rect -212 -455 -183 -81
rect -137 -455 -108 -81
rect -212 -468 -108 -455
rect -52 -81 52 -68
rect -52 -455 -23 -81
rect 23 -455 52 -81
rect -52 -468 52 -455
rect 108 -81 212 -68
rect 108 -455 137 -81
rect 183 -455 212 -81
rect 108 -468 212 -455
rect 268 -81 372 -68
rect 268 -455 297 -81
rect 343 -455 372 -81
rect 268 -468 372 -455
rect 428 -81 532 -68
rect 428 -455 457 -81
rect 503 -455 532 -81
rect 428 -468 532 -455
rect 588 -81 692 -68
rect 588 -455 617 -81
rect 663 -455 692 -81
rect 588 -468 692 -455
rect 748 -81 852 -68
rect 748 -455 777 -81
rect 823 -455 852 -81
rect 748 -468 852 -455
rect 908 -81 1012 -68
rect 908 -455 937 -81
rect 983 -455 1012 -81
rect 908 -468 1012 -455
rect 1068 -81 1172 -68
rect 1068 -455 1097 -81
rect 1143 -455 1172 -81
rect 1068 -468 1172 -455
rect 1228 -81 1332 -68
rect 1228 -455 1257 -81
rect 1303 -455 1332 -81
rect 1228 -468 1332 -455
rect 1388 -81 1492 -68
rect 1388 -455 1417 -81
rect 1463 -455 1492 -81
rect 1388 -468 1492 -455
rect 1548 -81 1636 -68
rect 1548 -455 1577 -81
rect 1623 -455 1636 -81
rect 1548 -468 1636 -455
<< ndiffc >>
rect -1623 81 -1577 455
rect -1463 81 -1417 455
rect -1303 81 -1257 455
rect -1143 81 -1097 455
rect -983 81 -937 455
rect -823 81 -777 455
rect -663 81 -617 455
rect -503 81 -457 455
rect -343 81 -297 455
rect -183 81 -137 455
rect -23 81 23 455
rect 137 81 183 455
rect 297 81 343 455
rect 457 81 503 455
rect 617 81 663 455
rect 777 81 823 455
rect 937 81 983 455
rect 1097 81 1143 455
rect 1257 81 1303 455
rect 1417 81 1463 455
rect 1577 81 1623 455
rect -1623 -455 -1577 -81
rect -1463 -455 -1417 -81
rect -1303 -455 -1257 -81
rect -1143 -455 -1097 -81
rect -983 -455 -937 -81
rect -823 -455 -777 -81
rect -663 -455 -617 -81
rect -503 -455 -457 -81
rect -343 -455 -297 -81
rect -183 -455 -137 -81
rect -23 -455 23 -81
rect 137 -455 183 -81
rect 297 -455 343 -81
rect 457 -455 503 -81
rect 617 -455 663 -81
rect 777 -455 823 -81
rect 937 -455 983 -81
rect 1097 -455 1143 -81
rect 1257 -455 1303 -81
rect 1417 -455 1463 -81
rect 1577 -455 1623 -81
<< polysilicon >>
rect -1548 468 -1492 512
rect -1388 468 -1332 512
rect -1228 468 -1172 512
rect -1068 468 -1012 512
rect -908 468 -852 512
rect -748 468 -692 512
rect -588 468 -532 512
rect -428 468 -372 512
rect -268 468 -212 512
rect -108 468 -52 512
rect 52 468 108 512
rect 212 468 268 512
rect 372 468 428 512
rect 532 468 588 512
rect 692 468 748 512
rect 852 468 908 512
rect 1012 468 1068 512
rect 1172 468 1228 512
rect 1332 468 1388 512
rect 1492 468 1548 512
rect -1548 24 -1492 68
rect -1388 24 -1332 68
rect -1228 24 -1172 68
rect -1068 24 -1012 68
rect -908 24 -852 68
rect -748 24 -692 68
rect -588 24 -532 68
rect -428 24 -372 68
rect -268 24 -212 68
rect -108 24 -52 68
rect 52 24 108 68
rect 212 24 268 68
rect 372 24 428 68
rect 532 24 588 68
rect 692 24 748 68
rect 852 24 908 68
rect 1012 24 1068 68
rect 1172 24 1228 68
rect 1332 24 1388 68
rect 1492 24 1548 68
rect -1548 -68 -1492 -24
rect -1388 -68 -1332 -24
rect -1228 -68 -1172 -24
rect -1068 -68 -1012 -24
rect -908 -68 -852 -24
rect -748 -68 -692 -24
rect -588 -68 -532 -24
rect -428 -68 -372 -24
rect -268 -68 -212 -24
rect -108 -68 -52 -24
rect 52 -68 108 -24
rect 212 -68 268 -24
rect 372 -68 428 -24
rect 532 -68 588 -24
rect 692 -68 748 -24
rect 852 -68 908 -24
rect 1012 -68 1068 -24
rect 1172 -68 1228 -24
rect 1332 -68 1388 -24
rect 1492 -68 1548 -24
rect -1548 -512 -1492 -468
rect -1388 -512 -1332 -468
rect -1228 -512 -1172 -468
rect -1068 -512 -1012 -468
rect -908 -512 -852 -468
rect -748 -512 -692 -468
rect -588 -512 -532 -468
rect -428 -512 -372 -468
rect -268 -512 -212 -468
rect -108 -512 -52 -468
rect 52 -512 108 -468
rect 212 -512 268 -468
rect 372 -512 428 -468
rect 532 -512 588 -468
rect 692 -512 748 -468
rect 852 -512 908 -468
rect 1012 -512 1068 -468
rect 1172 -512 1228 -468
rect 1332 -512 1388 -468
rect 1492 -512 1548 -468
<< metal1 >>
rect -1623 455 -1577 466
rect -1623 70 -1577 81
rect -1463 455 -1417 466
rect -1463 70 -1417 81
rect -1303 455 -1257 466
rect -1303 70 -1257 81
rect -1143 455 -1097 466
rect -1143 70 -1097 81
rect -983 455 -937 466
rect -983 70 -937 81
rect -823 455 -777 466
rect -823 70 -777 81
rect -663 455 -617 466
rect -663 70 -617 81
rect -503 455 -457 466
rect -503 70 -457 81
rect -343 455 -297 466
rect -343 70 -297 81
rect -183 455 -137 466
rect -183 70 -137 81
rect -23 455 23 466
rect -23 70 23 81
rect 137 455 183 466
rect 137 70 183 81
rect 297 455 343 466
rect 297 70 343 81
rect 457 455 503 466
rect 457 70 503 81
rect 617 455 663 466
rect 617 70 663 81
rect 777 455 823 466
rect 777 70 823 81
rect 937 455 983 466
rect 937 70 983 81
rect 1097 455 1143 466
rect 1097 70 1143 81
rect 1257 455 1303 466
rect 1257 70 1303 81
rect 1417 455 1463 466
rect 1417 70 1463 81
rect 1577 455 1623 466
rect 1577 70 1623 81
rect -1623 -81 -1577 -70
rect -1623 -466 -1577 -455
rect -1463 -81 -1417 -70
rect -1463 -466 -1417 -455
rect -1303 -81 -1257 -70
rect -1303 -466 -1257 -455
rect -1143 -81 -1097 -70
rect -1143 -466 -1097 -455
rect -983 -81 -937 -70
rect -983 -466 -937 -455
rect -823 -81 -777 -70
rect -823 -466 -777 -455
rect -663 -81 -617 -70
rect -663 -466 -617 -455
rect -503 -81 -457 -70
rect -503 -466 -457 -455
rect -343 -81 -297 -70
rect -343 -466 -297 -455
rect -183 -81 -137 -70
rect -183 -466 -137 -455
rect -23 -81 23 -70
rect -23 -466 23 -455
rect 137 -81 183 -70
rect 137 -466 183 -455
rect 297 -81 343 -70
rect 297 -466 343 -455
rect 457 -81 503 -70
rect 457 -466 503 -455
rect 617 -81 663 -70
rect 617 -466 663 -455
rect 777 -81 823 -70
rect 777 -466 823 -455
rect 937 -81 983 -70
rect 937 -466 983 -455
rect 1097 -81 1143 -70
rect 1097 -466 1143 -455
rect 1257 -81 1303 -70
rect 1257 -466 1303 -455
rect 1417 -81 1463 -70
rect 1417 -466 1463 -455
rect 1577 -81 1623 -70
rect 1577 -466 1623 -455
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 2.0 l 0.280 m 2 nf 20 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
