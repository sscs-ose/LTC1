magic
tech gf180mcuC
magscale 1 10
timestamp 1694434822
<< nwell >>
rect -1104 -1148 1104 1148
<< nsubdiff >>
rect -1080 1052 1080 1124
rect -1080 -1052 -1008 1052
rect 1008 -1052 1080 1052
rect -1080 -1124 1080 -1052
<< polysilicon >>
rect -920 951 -680 964
rect -920 905 -907 951
rect -693 905 -680 951
rect -920 862 -680 905
rect -920 619 -680 662
rect -920 573 -907 619
rect -693 573 -680 619
rect -920 560 -680 573
rect -600 951 -360 964
rect -600 905 -587 951
rect -373 905 -360 951
rect -600 862 -360 905
rect -600 619 -360 662
rect -600 573 -587 619
rect -373 573 -360 619
rect -600 560 -360 573
rect -280 951 -40 964
rect -280 905 -267 951
rect -53 905 -40 951
rect -280 862 -40 905
rect -280 619 -40 662
rect -280 573 -267 619
rect -53 573 -40 619
rect -280 560 -40 573
rect 40 951 280 964
rect 40 905 53 951
rect 267 905 280 951
rect 40 862 280 905
rect 40 619 280 662
rect 40 573 53 619
rect 267 573 280 619
rect 40 560 280 573
rect 360 951 600 964
rect 360 905 373 951
rect 587 905 600 951
rect 360 862 600 905
rect 360 619 600 662
rect 360 573 373 619
rect 587 573 600 619
rect 360 560 600 573
rect 680 951 920 964
rect 680 905 693 951
rect 907 905 920 951
rect 680 862 920 905
rect 680 619 920 662
rect 680 573 693 619
rect 907 573 920 619
rect 680 560 920 573
rect -920 443 -680 456
rect -920 397 -907 443
rect -693 397 -680 443
rect -920 354 -680 397
rect -920 111 -680 154
rect -920 65 -907 111
rect -693 65 -680 111
rect -920 52 -680 65
rect -600 443 -360 456
rect -600 397 -587 443
rect -373 397 -360 443
rect -600 354 -360 397
rect -600 111 -360 154
rect -600 65 -587 111
rect -373 65 -360 111
rect -600 52 -360 65
rect -280 443 -40 456
rect -280 397 -267 443
rect -53 397 -40 443
rect -280 354 -40 397
rect -280 111 -40 154
rect -280 65 -267 111
rect -53 65 -40 111
rect -280 52 -40 65
rect 40 443 280 456
rect 40 397 53 443
rect 267 397 280 443
rect 40 354 280 397
rect 40 111 280 154
rect 40 65 53 111
rect 267 65 280 111
rect 40 52 280 65
rect 360 443 600 456
rect 360 397 373 443
rect 587 397 600 443
rect 360 354 600 397
rect 360 111 600 154
rect 360 65 373 111
rect 587 65 600 111
rect 360 52 600 65
rect 680 443 920 456
rect 680 397 693 443
rect 907 397 920 443
rect 680 354 920 397
rect 680 111 920 154
rect 680 65 693 111
rect 907 65 920 111
rect 680 52 920 65
rect -920 -65 -680 -52
rect -920 -111 -907 -65
rect -693 -111 -680 -65
rect -920 -154 -680 -111
rect -920 -397 -680 -354
rect -920 -443 -907 -397
rect -693 -443 -680 -397
rect -920 -456 -680 -443
rect -600 -65 -360 -52
rect -600 -111 -587 -65
rect -373 -111 -360 -65
rect -600 -154 -360 -111
rect -600 -397 -360 -354
rect -600 -443 -587 -397
rect -373 -443 -360 -397
rect -600 -456 -360 -443
rect -280 -65 -40 -52
rect -280 -111 -267 -65
rect -53 -111 -40 -65
rect -280 -154 -40 -111
rect -280 -397 -40 -354
rect -280 -443 -267 -397
rect -53 -443 -40 -397
rect -280 -456 -40 -443
rect 40 -65 280 -52
rect 40 -111 53 -65
rect 267 -111 280 -65
rect 40 -154 280 -111
rect 40 -397 280 -354
rect 40 -443 53 -397
rect 267 -443 280 -397
rect 40 -456 280 -443
rect 360 -65 600 -52
rect 360 -111 373 -65
rect 587 -111 600 -65
rect 360 -154 600 -111
rect 360 -397 600 -354
rect 360 -443 373 -397
rect 587 -443 600 -397
rect 360 -456 600 -443
rect 680 -65 920 -52
rect 680 -111 693 -65
rect 907 -111 920 -65
rect 680 -154 920 -111
rect 680 -397 920 -354
rect 680 -443 693 -397
rect 907 -443 920 -397
rect 680 -456 920 -443
rect -920 -573 -680 -560
rect -920 -619 -907 -573
rect -693 -619 -680 -573
rect -920 -662 -680 -619
rect -920 -905 -680 -862
rect -920 -951 -907 -905
rect -693 -951 -680 -905
rect -920 -964 -680 -951
rect -600 -573 -360 -560
rect -600 -619 -587 -573
rect -373 -619 -360 -573
rect -600 -662 -360 -619
rect -600 -905 -360 -862
rect -600 -951 -587 -905
rect -373 -951 -360 -905
rect -600 -964 -360 -951
rect -280 -573 -40 -560
rect -280 -619 -267 -573
rect -53 -619 -40 -573
rect -280 -662 -40 -619
rect -280 -905 -40 -862
rect -280 -951 -267 -905
rect -53 -951 -40 -905
rect -280 -964 -40 -951
rect 40 -573 280 -560
rect 40 -619 53 -573
rect 267 -619 280 -573
rect 40 -662 280 -619
rect 40 -905 280 -862
rect 40 -951 53 -905
rect 267 -951 280 -905
rect 40 -964 280 -951
rect 360 -573 600 -560
rect 360 -619 373 -573
rect 587 -619 600 -573
rect 360 -662 600 -619
rect 360 -905 600 -862
rect 360 -951 373 -905
rect 587 -951 600 -905
rect 360 -964 600 -951
rect 680 -573 920 -560
rect 680 -619 693 -573
rect 907 -619 920 -573
rect 680 -662 920 -619
rect 680 -905 920 -862
rect 680 -951 693 -905
rect 907 -951 920 -905
rect 680 -964 920 -951
<< polycontact >>
rect -907 905 -693 951
rect -907 573 -693 619
rect -587 905 -373 951
rect -587 573 -373 619
rect -267 905 -53 951
rect -267 573 -53 619
rect 53 905 267 951
rect 53 573 267 619
rect 373 905 587 951
rect 373 573 587 619
rect 693 905 907 951
rect 693 573 907 619
rect -907 397 -693 443
rect -907 65 -693 111
rect -587 397 -373 443
rect -587 65 -373 111
rect -267 397 -53 443
rect -267 65 -53 111
rect 53 397 267 443
rect 53 65 267 111
rect 373 397 587 443
rect 373 65 587 111
rect 693 397 907 443
rect 693 65 907 111
rect -907 -111 -693 -65
rect -907 -443 -693 -397
rect -587 -111 -373 -65
rect -587 -443 -373 -397
rect -267 -111 -53 -65
rect -267 -443 -53 -397
rect 53 -111 267 -65
rect 53 -443 267 -397
rect 373 -111 587 -65
rect 373 -443 587 -397
rect 693 -111 907 -65
rect 693 -443 907 -397
rect -907 -619 -693 -573
rect -907 -951 -693 -905
rect -587 -619 -373 -573
rect -587 -951 -373 -905
rect -267 -619 -53 -573
rect -267 -951 -53 -905
rect 53 -619 267 -573
rect 53 -951 267 -905
rect 373 -619 587 -573
rect 373 -951 587 -905
rect 693 -619 907 -573
rect 693 -951 907 -905
<< ppolyres >>
rect -920 662 -680 862
rect -600 662 -360 862
rect -280 662 -40 862
rect 40 662 280 862
rect 360 662 600 862
rect 680 662 920 862
rect -920 154 -680 354
rect -600 154 -360 354
rect -280 154 -40 354
rect 40 154 280 354
rect 360 154 600 354
rect 680 154 920 354
rect -920 -354 -680 -154
rect -600 -354 -360 -154
rect -280 -354 -40 -154
rect 40 -354 280 -154
rect 360 -354 600 -154
rect 680 -354 920 -154
rect -920 -862 -680 -662
rect -600 -862 -360 -662
rect -280 -862 -40 -662
rect 40 -862 280 -662
rect 360 -862 600 -662
rect 680 -862 920 -662
<< metal1 >>
rect -918 905 -907 951
rect -693 905 -682 951
rect -598 905 -587 951
rect -373 905 -362 951
rect -278 905 -267 951
rect -53 905 -42 951
rect 42 905 53 951
rect 267 905 278 951
rect 362 905 373 951
rect 587 905 598 951
rect 682 905 693 951
rect 907 905 918 951
rect -918 573 -907 619
rect -693 573 -682 619
rect -598 573 -587 619
rect -373 573 -362 619
rect -278 573 -267 619
rect -53 573 -42 619
rect 42 573 53 619
rect 267 573 278 619
rect 362 573 373 619
rect 587 573 598 619
rect 682 573 693 619
rect 907 573 918 619
rect -918 397 -907 443
rect -693 397 -682 443
rect -598 397 -587 443
rect -373 397 -362 443
rect -278 397 -267 443
rect -53 397 -42 443
rect 42 397 53 443
rect 267 397 278 443
rect 362 397 373 443
rect 587 397 598 443
rect 682 397 693 443
rect 907 397 918 443
rect -918 65 -907 111
rect -693 65 -682 111
rect -598 65 -587 111
rect -373 65 -362 111
rect -278 65 -267 111
rect -53 65 -42 111
rect 42 65 53 111
rect 267 65 278 111
rect 362 65 373 111
rect 587 65 598 111
rect 682 65 693 111
rect 907 65 918 111
rect -918 -111 -907 -65
rect -693 -111 -682 -65
rect -598 -111 -587 -65
rect -373 -111 -362 -65
rect -278 -111 -267 -65
rect -53 -111 -42 -65
rect 42 -111 53 -65
rect 267 -111 278 -65
rect 362 -111 373 -65
rect 587 -111 598 -65
rect 682 -111 693 -65
rect 907 -111 918 -65
rect -918 -443 -907 -397
rect -693 -443 -682 -397
rect -598 -443 -587 -397
rect -373 -443 -362 -397
rect -278 -443 -267 -397
rect -53 -443 -42 -397
rect 42 -443 53 -397
rect 267 -443 278 -397
rect 362 -443 373 -397
rect 587 -443 598 -397
rect 682 -443 693 -397
rect 907 -443 918 -397
rect -918 -619 -907 -573
rect -693 -619 -682 -573
rect -598 -619 -587 -573
rect -373 -619 -362 -573
rect -278 -619 -267 -573
rect -53 -619 -42 -573
rect 42 -619 53 -573
rect 267 -619 278 -573
rect 362 -619 373 -573
rect 587 -619 598 -573
rect 682 -619 693 -573
rect 907 -619 918 -573
rect -918 -951 -907 -905
rect -693 -951 -682 -905
rect -598 -951 -587 -905
rect -373 -951 -362 -905
rect -278 -951 -267 -905
rect -53 -951 -42 -905
rect 42 -951 53 -905
rect 267 -951 278 -905
rect 362 -951 373 -905
rect 587 -951 598 -905
rect 682 -951 693 -905
rect 907 -951 918 -905
<< properties >>
string FIXED_BBOX -1044 -1088 1044 1088
string gencell ppolyf_u
string library gf180mcu
string parameters w 1.2 l 1.0 m 4 nx 6 wmin 0.80 lmin 1.00 rho 315 val 278.761 dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 0 grc 0 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 0
<< end >>
