magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2045 -2562 2045 2562
<< psubdiff >>
rect -45 540 45 562
rect -45 -540 -23 540
rect 23 -540 45 540
rect -45 -562 45 -540
<< psubdiffcont >>
rect -23 -540 23 540
<< metal1 >>
rect -34 540 34 551
rect -34 -540 -23 540
rect 23 -540 34 540
rect -34 -551 34 -540
<< end >>
