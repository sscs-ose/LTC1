magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -3103 -2109 3103 2109
<< metal2 >>
rect -1103 99 1103 109
rect -1103 43 -1093 99
rect -1037 43 -951 99
rect -895 43 -809 99
rect -753 43 -667 99
rect -611 43 -525 99
rect -469 43 -383 99
rect -327 43 -241 99
rect -185 43 -99 99
rect -43 43 43 99
rect 99 43 185 99
rect 241 43 327 99
rect 383 43 469 99
rect 525 43 611 99
rect 667 43 753 99
rect 809 43 895 99
rect 951 43 1037 99
rect 1093 43 1103 99
rect -1103 -43 1103 43
rect -1103 -99 -1093 -43
rect -1037 -99 -951 -43
rect -895 -99 -809 -43
rect -753 -99 -667 -43
rect -611 -99 -525 -43
rect -469 -99 -383 -43
rect -327 -99 -241 -43
rect -185 -99 -99 -43
rect -43 -99 43 -43
rect 99 -99 185 -43
rect 241 -99 327 -43
rect 383 -99 469 -43
rect 525 -99 611 -43
rect 667 -99 753 -43
rect 809 -99 895 -43
rect 951 -99 1037 -43
rect 1093 -99 1103 -43
rect -1103 -109 1103 -99
<< via2 >>
rect -1093 43 -1037 99
rect -951 43 -895 99
rect -809 43 -753 99
rect -667 43 -611 99
rect -525 43 -469 99
rect -383 43 -327 99
rect -241 43 -185 99
rect -99 43 -43 99
rect 43 43 99 99
rect 185 43 241 99
rect 327 43 383 99
rect 469 43 525 99
rect 611 43 667 99
rect 753 43 809 99
rect 895 43 951 99
rect 1037 43 1093 99
rect -1093 -99 -1037 -43
rect -951 -99 -895 -43
rect -809 -99 -753 -43
rect -667 -99 -611 -43
rect -525 -99 -469 -43
rect -383 -99 -327 -43
rect -241 -99 -185 -43
rect -99 -99 -43 -43
rect 43 -99 99 -43
rect 185 -99 241 -43
rect 327 -99 383 -43
rect 469 -99 525 -43
rect 611 -99 667 -43
rect 753 -99 809 -43
rect 895 -99 951 -43
rect 1037 -99 1093 -43
<< metal3 >>
rect -1103 99 1103 109
rect -1103 43 -1093 99
rect -1037 43 -951 99
rect -895 43 -809 99
rect -753 43 -667 99
rect -611 43 -525 99
rect -469 43 -383 99
rect -327 43 -241 99
rect -185 43 -99 99
rect -43 43 43 99
rect 99 43 185 99
rect 241 43 327 99
rect 383 43 469 99
rect 525 43 611 99
rect 667 43 753 99
rect 809 43 895 99
rect 951 43 1037 99
rect 1093 43 1103 99
rect -1103 -43 1103 43
rect -1103 -99 -1093 -43
rect -1037 -99 -951 -43
rect -895 -99 -809 -43
rect -753 -99 -667 -43
rect -611 -99 -525 -43
rect -469 -99 -383 -43
rect -327 -99 -241 -43
rect -185 -99 -99 -43
rect -43 -99 43 -43
rect 99 -99 185 -43
rect 241 -99 327 -43
rect 383 -99 469 -43
rect 525 -99 611 -43
rect 667 -99 753 -43
rect 809 -99 895 -43
rect 951 -99 1037 -43
rect 1093 -99 1103 -43
rect -1103 -109 1103 -99
<< end >>
