magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1071 -1123 1071 1123
<< metal1 >>
rect -71 117 71 123
rect -71 -117 -65 117
rect 65 -117 71 117
rect -71 -123 71 -117
<< via1 >>
rect -65 -117 65 117
<< metal2 >>
rect -71 117 71 123
rect -71 -117 -65 117
rect 65 -117 71 117
rect -71 -123 71 -117
<< end >>
