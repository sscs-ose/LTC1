magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1679 -1316 1679 1316
<< metal1 >>
rect -679 310 679 316
rect -679 284 -673 310
rect -647 284 -607 310
rect -581 284 -541 310
rect -515 284 -475 310
rect -449 284 -409 310
rect -383 284 -343 310
rect -317 284 -277 310
rect -251 284 -211 310
rect -185 284 -145 310
rect -119 284 -79 310
rect -53 284 -13 310
rect 13 284 53 310
rect 79 284 119 310
rect 145 284 185 310
rect 211 284 251 310
rect 277 284 317 310
rect 343 284 383 310
rect 409 284 449 310
rect 475 284 515 310
rect 541 284 581 310
rect 607 284 647 310
rect 673 284 679 310
rect -679 244 679 284
rect -679 218 -673 244
rect -647 218 -607 244
rect -581 218 -541 244
rect -515 218 -475 244
rect -449 218 -409 244
rect -383 218 -343 244
rect -317 218 -277 244
rect -251 218 -211 244
rect -185 218 -145 244
rect -119 218 -79 244
rect -53 218 -13 244
rect 13 218 53 244
rect 79 218 119 244
rect 145 218 185 244
rect 211 218 251 244
rect 277 218 317 244
rect 343 218 383 244
rect 409 218 449 244
rect 475 218 515 244
rect 541 218 581 244
rect 607 218 647 244
rect 673 218 679 244
rect -679 178 679 218
rect -679 152 -673 178
rect -647 152 -607 178
rect -581 152 -541 178
rect -515 152 -475 178
rect -449 152 -409 178
rect -383 152 -343 178
rect -317 152 -277 178
rect -251 152 -211 178
rect -185 152 -145 178
rect -119 152 -79 178
rect -53 152 -13 178
rect 13 152 53 178
rect 79 152 119 178
rect 145 152 185 178
rect 211 152 251 178
rect 277 152 317 178
rect 343 152 383 178
rect 409 152 449 178
rect 475 152 515 178
rect 541 152 581 178
rect 607 152 647 178
rect 673 152 679 178
rect -679 112 679 152
rect -679 86 -673 112
rect -647 86 -607 112
rect -581 86 -541 112
rect -515 86 -475 112
rect -449 86 -409 112
rect -383 86 -343 112
rect -317 86 -277 112
rect -251 86 -211 112
rect -185 86 -145 112
rect -119 86 -79 112
rect -53 86 -13 112
rect 13 86 53 112
rect 79 86 119 112
rect 145 86 185 112
rect 211 86 251 112
rect 277 86 317 112
rect 343 86 383 112
rect 409 86 449 112
rect 475 86 515 112
rect 541 86 581 112
rect 607 86 647 112
rect 673 86 679 112
rect -679 46 679 86
rect -679 20 -673 46
rect -647 20 -607 46
rect -581 20 -541 46
rect -515 20 -475 46
rect -449 20 -409 46
rect -383 20 -343 46
rect -317 20 -277 46
rect -251 20 -211 46
rect -185 20 -145 46
rect -119 20 -79 46
rect -53 20 -13 46
rect 13 20 53 46
rect 79 20 119 46
rect 145 20 185 46
rect 211 20 251 46
rect 277 20 317 46
rect 343 20 383 46
rect 409 20 449 46
rect 475 20 515 46
rect 541 20 581 46
rect 607 20 647 46
rect 673 20 679 46
rect -679 -20 679 20
rect -679 -46 -673 -20
rect -647 -46 -607 -20
rect -581 -46 -541 -20
rect -515 -46 -475 -20
rect -449 -46 -409 -20
rect -383 -46 -343 -20
rect -317 -46 -277 -20
rect -251 -46 -211 -20
rect -185 -46 -145 -20
rect -119 -46 -79 -20
rect -53 -46 -13 -20
rect 13 -46 53 -20
rect 79 -46 119 -20
rect 145 -46 185 -20
rect 211 -46 251 -20
rect 277 -46 317 -20
rect 343 -46 383 -20
rect 409 -46 449 -20
rect 475 -46 515 -20
rect 541 -46 581 -20
rect 607 -46 647 -20
rect 673 -46 679 -20
rect -679 -86 679 -46
rect -679 -112 -673 -86
rect -647 -112 -607 -86
rect -581 -112 -541 -86
rect -515 -112 -475 -86
rect -449 -112 -409 -86
rect -383 -112 -343 -86
rect -317 -112 -277 -86
rect -251 -112 -211 -86
rect -185 -112 -145 -86
rect -119 -112 -79 -86
rect -53 -112 -13 -86
rect 13 -112 53 -86
rect 79 -112 119 -86
rect 145 -112 185 -86
rect 211 -112 251 -86
rect 277 -112 317 -86
rect 343 -112 383 -86
rect 409 -112 449 -86
rect 475 -112 515 -86
rect 541 -112 581 -86
rect 607 -112 647 -86
rect 673 -112 679 -86
rect -679 -152 679 -112
rect -679 -178 -673 -152
rect -647 -178 -607 -152
rect -581 -178 -541 -152
rect -515 -178 -475 -152
rect -449 -178 -409 -152
rect -383 -178 -343 -152
rect -317 -178 -277 -152
rect -251 -178 -211 -152
rect -185 -178 -145 -152
rect -119 -178 -79 -152
rect -53 -178 -13 -152
rect 13 -178 53 -152
rect 79 -178 119 -152
rect 145 -178 185 -152
rect 211 -178 251 -152
rect 277 -178 317 -152
rect 343 -178 383 -152
rect 409 -178 449 -152
rect 475 -178 515 -152
rect 541 -178 581 -152
rect 607 -178 647 -152
rect 673 -178 679 -152
rect -679 -218 679 -178
rect -679 -244 -673 -218
rect -647 -244 -607 -218
rect -581 -244 -541 -218
rect -515 -244 -475 -218
rect -449 -244 -409 -218
rect -383 -244 -343 -218
rect -317 -244 -277 -218
rect -251 -244 -211 -218
rect -185 -244 -145 -218
rect -119 -244 -79 -218
rect -53 -244 -13 -218
rect 13 -244 53 -218
rect 79 -244 119 -218
rect 145 -244 185 -218
rect 211 -244 251 -218
rect 277 -244 317 -218
rect 343 -244 383 -218
rect 409 -244 449 -218
rect 475 -244 515 -218
rect 541 -244 581 -218
rect 607 -244 647 -218
rect 673 -244 679 -218
rect -679 -284 679 -244
rect -679 -310 -673 -284
rect -647 -310 -607 -284
rect -581 -310 -541 -284
rect -515 -310 -475 -284
rect -449 -310 -409 -284
rect -383 -310 -343 -284
rect -317 -310 -277 -284
rect -251 -310 -211 -284
rect -185 -310 -145 -284
rect -119 -310 -79 -284
rect -53 -310 -13 -284
rect 13 -310 53 -284
rect 79 -310 119 -284
rect 145 -310 185 -284
rect 211 -310 251 -284
rect 277 -310 317 -284
rect 343 -310 383 -284
rect 409 -310 449 -284
rect 475 -310 515 -284
rect 541 -310 581 -284
rect 607 -310 647 -284
rect 673 -310 679 -284
rect -679 -316 679 -310
<< via1 >>
rect -673 284 -647 310
rect -607 284 -581 310
rect -541 284 -515 310
rect -475 284 -449 310
rect -409 284 -383 310
rect -343 284 -317 310
rect -277 284 -251 310
rect -211 284 -185 310
rect -145 284 -119 310
rect -79 284 -53 310
rect -13 284 13 310
rect 53 284 79 310
rect 119 284 145 310
rect 185 284 211 310
rect 251 284 277 310
rect 317 284 343 310
rect 383 284 409 310
rect 449 284 475 310
rect 515 284 541 310
rect 581 284 607 310
rect 647 284 673 310
rect -673 218 -647 244
rect -607 218 -581 244
rect -541 218 -515 244
rect -475 218 -449 244
rect -409 218 -383 244
rect -343 218 -317 244
rect -277 218 -251 244
rect -211 218 -185 244
rect -145 218 -119 244
rect -79 218 -53 244
rect -13 218 13 244
rect 53 218 79 244
rect 119 218 145 244
rect 185 218 211 244
rect 251 218 277 244
rect 317 218 343 244
rect 383 218 409 244
rect 449 218 475 244
rect 515 218 541 244
rect 581 218 607 244
rect 647 218 673 244
rect -673 152 -647 178
rect -607 152 -581 178
rect -541 152 -515 178
rect -475 152 -449 178
rect -409 152 -383 178
rect -343 152 -317 178
rect -277 152 -251 178
rect -211 152 -185 178
rect -145 152 -119 178
rect -79 152 -53 178
rect -13 152 13 178
rect 53 152 79 178
rect 119 152 145 178
rect 185 152 211 178
rect 251 152 277 178
rect 317 152 343 178
rect 383 152 409 178
rect 449 152 475 178
rect 515 152 541 178
rect 581 152 607 178
rect 647 152 673 178
rect -673 86 -647 112
rect -607 86 -581 112
rect -541 86 -515 112
rect -475 86 -449 112
rect -409 86 -383 112
rect -343 86 -317 112
rect -277 86 -251 112
rect -211 86 -185 112
rect -145 86 -119 112
rect -79 86 -53 112
rect -13 86 13 112
rect 53 86 79 112
rect 119 86 145 112
rect 185 86 211 112
rect 251 86 277 112
rect 317 86 343 112
rect 383 86 409 112
rect 449 86 475 112
rect 515 86 541 112
rect 581 86 607 112
rect 647 86 673 112
rect -673 20 -647 46
rect -607 20 -581 46
rect -541 20 -515 46
rect -475 20 -449 46
rect -409 20 -383 46
rect -343 20 -317 46
rect -277 20 -251 46
rect -211 20 -185 46
rect -145 20 -119 46
rect -79 20 -53 46
rect -13 20 13 46
rect 53 20 79 46
rect 119 20 145 46
rect 185 20 211 46
rect 251 20 277 46
rect 317 20 343 46
rect 383 20 409 46
rect 449 20 475 46
rect 515 20 541 46
rect 581 20 607 46
rect 647 20 673 46
rect -673 -46 -647 -20
rect -607 -46 -581 -20
rect -541 -46 -515 -20
rect -475 -46 -449 -20
rect -409 -46 -383 -20
rect -343 -46 -317 -20
rect -277 -46 -251 -20
rect -211 -46 -185 -20
rect -145 -46 -119 -20
rect -79 -46 -53 -20
rect -13 -46 13 -20
rect 53 -46 79 -20
rect 119 -46 145 -20
rect 185 -46 211 -20
rect 251 -46 277 -20
rect 317 -46 343 -20
rect 383 -46 409 -20
rect 449 -46 475 -20
rect 515 -46 541 -20
rect 581 -46 607 -20
rect 647 -46 673 -20
rect -673 -112 -647 -86
rect -607 -112 -581 -86
rect -541 -112 -515 -86
rect -475 -112 -449 -86
rect -409 -112 -383 -86
rect -343 -112 -317 -86
rect -277 -112 -251 -86
rect -211 -112 -185 -86
rect -145 -112 -119 -86
rect -79 -112 -53 -86
rect -13 -112 13 -86
rect 53 -112 79 -86
rect 119 -112 145 -86
rect 185 -112 211 -86
rect 251 -112 277 -86
rect 317 -112 343 -86
rect 383 -112 409 -86
rect 449 -112 475 -86
rect 515 -112 541 -86
rect 581 -112 607 -86
rect 647 -112 673 -86
rect -673 -178 -647 -152
rect -607 -178 -581 -152
rect -541 -178 -515 -152
rect -475 -178 -449 -152
rect -409 -178 -383 -152
rect -343 -178 -317 -152
rect -277 -178 -251 -152
rect -211 -178 -185 -152
rect -145 -178 -119 -152
rect -79 -178 -53 -152
rect -13 -178 13 -152
rect 53 -178 79 -152
rect 119 -178 145 -152
rect 185 -178 211 -152
rect 251 -178 277 -152
rect 317 -178 343 -152
rect 383 -178 409 -152
rect 449 -178 475 -152
rect 515 -178 541 -152
rect 581 -178 607 -152
rect 647 -178 673 -152
rect -673 -244 -647 -218
rect -607 -244 -581 -218
rect -541 -244 -515 -218
rect -475 -244 -449 -218
rect -409 -244 -383 -218
rect -343 -244 -317 -218
rect -277 -244 -251 -218
rect -211 -244 -185 -218
rect -145 -244 -119 -218
rect -79 -244 -53 -218
rect -13 -244 13 -218
rect 53 -244 79 -218
rect 119 -244 145 -218
rect 185 -244 211 -218
rect 251 -244 277 -218
rect 317 -244 343 -218
rect 383 -244 409 -218
rect 449 -244 475 -218
rect 515 -244 541 -218
rect 581 -244 607 -218
rect 647 -244 673 -218
rect -673 -310 -647 -284
rect -607 -310 -581 -284
rect -541 -310 -515 -284
rect -475 -310 -449 -284
rect -409 -310 -383 -284
rect -343 -310 -317 -284
rect -277 -310 -251 -284
rect -211 -310 -185 -284
rect -145 -310 -119 -284
rect -79 -310 -53 -284
rect -13 -310 13 -284
rect 53 -310 79 -284
rect 119 -310 145 -284
rect 185 -310 211 -284
rect 251 -310 277 -284
rect 317 -310 343 -284
rect 383 -310 409 -284
rect 449 -310 475 -284
rect 515 -310 541 -284
rect 581 -310 607 -284
rect 647 -310 673 -284
<< metal2 >>
rect -679 310 679 316
rect -679 284 -673 310
rect -647 284 -607 310
rect -581 284 -541 310
rect -515 284 -475 310
rect -449 284 -409 310
rect -383 284 -343 310
rect -317 284 -277 310
rect -251 284 -211 310
rect -185 284 -145 310
rect -119 284 -79 310
rect -53 284 -13 310
rect 13 284 53 310
rect 79 284 119 310
rect 145 284 185 310
rect 211 284 251 310
rect 277 284 317 310
rect 343 284 383 310
rect 409 284 449 310
rect 475 284 515 310
rect 541 284 581 310
rect 607 284 647 310
rect 673 284 679 310
rect -679 244 679 284
rect -679 218 -673 244
rect -647 218 -607 244
rect -581 218 -541 244
rect -515 218 -475 244
rect -449 218 -409 244
rect -383 218 -343 244
rect -317 218 -277 244
rect -251 218 -211 244
rect -185 218 -145 244
rect -119 218 -79 244
rect -53 218 -13 244
rect 13 218 53 244
rect 79 218 119 244
rect 145 218 185 244
rect 211 218 251 244
rect 277 218 317 244
rect 343 218 383 244
rect 409 218 449 244
rect 475 218 515 244
rect 541 218 581 244
rect 607 218 647 244
rect 673 218 679 244
rect -679 178 679 218
rect -679 152 -673 178
rect -647 152 -607 178
rect -581 152 -541 178
rect -515 152 -475 178
rect -449 152 -409 178
rect -383 152 -343 178
rect -317 152 -277 178
rect -251 152 -211 178
rect -185 152 -145 178
rect -119 152 -79 178
rect -53 152 -13 178
rect 13 152 53 178
rect 79 152 119 178
rect 145 152 185 178
rect 211 152 251 178
rect 277 152 317 178
rect 343 152 383 178
rect 409 152 449 178
rect 475 152 515 178
rect 541 152 581 178
rect 607 152 647 178
rect 673 152 679 178
rect -679 112 679 152
rect -679 86 -673 112
rect -647 86 -607 112
rect -581 86 -541 112
rect -515 86 -475 112
rect -449 86 -409 112
rect -383 86 -343 112
rect -317 86 -277 112
rect -251 86 -211 112
rect -185 86 -145 112
rect -119 86 -79 112
rect -53 86 -13 112
rect 13 86 53 112
rect 79 86 119 112
rect 145 86 185 112
rect 211 86 251 112
rect 277 86 317 112
rect 343 86 383 112
rect 409 86 449 112
rect 475 86 515 112
rect 541 86 581 112
rect 607 86 647 112
rect 673 86 679 112
rect -679 46 679 86
rect -679 20 -673 46
rect -647 20 -607 46
rect -581 20 -541 46
rect -515 20 -475 46
rect -449 20 -409 46
rect -383 20 -343 46
rect -317 20 -277 46
rect -251 20 -211 46
rect -185 20 -145 46
rect -119 20 -79 46
rect -53 20 -13 46
rect 13 20 53 46
rect 79 20 119 46
rect 145 20 185 46
rect 211 20 251 46
rect 277 20 317 46
rect 343 20 383 46
rect 409 20 449 46
rect 475 20 515 46
rect 541 20 581 46
rect 607 20 647 46
rect 673 20 679 46
rect -679 -20 679 20
rect -679 -46 -673 -20
rect -647 -46 -607 -20
rect -581 -46 -541 -20
rect -515 -46 -475 -20
rect -449 -46 -409 -20
rect -383 -46 -343 -20
rect -317 -46 -277 -20
rect -251 -46 -211 -20
rect -185 -46 -145 -20
rect -119 -46 -79 -20
rect -53 -46 -13 -20
rect 13 -46 53 -20
rect 79 -46 119 -20
rect 145 -46 185 -20
rect 211 -46 251 -20
rect 277 -46 317 -20
rect 343 -46 383 -20
rect 409 -46 449 -20
rect 475 -46 515 -20
rect 541 -46 581 -20
rect 607 -46 647 -20
rect 673 -46 679 -20
rect -679 -86 679 -46
rect -679 -112 -673 -86
rect -647 -112 -607 -86
rect -581 -112 -541 -86
rect -515 -112 -475 -86
rect -449 -112 -409 -86
rect -383 -112 -343 -86
rect -317 -112 -277 -86
rect -251 -112 -211 -86
rect -185 -112 -145 -86
rect -119 -112 -79 -86
rect -53 -112 -13 -86
rect 13 -112 53 -86
rect 79 -112 119 -86
rect 145 -112 185 -86
rect 211 -112 251 -86
rect 277 -112 317 -86
rect 343 -112 383 -86
rect 409 -112 449 -86
rect 475 -112 515 -86
rect 541 -112 581 -86
rect 607 -112 647 -86
rect 673 -112 679 -86
rect -679 -152 679 -112
rect -679 -178 -673 -152
rect -647 -178 -607 -152
rect -581 -178 -541 -152
rect -515 -178 -475 -152
rect -449 -178 -409 -152
rect -383 -178 -343 -152
rect -317 -178 -277 -152
rect -251 -178 -211 -152
rect -185 -178 -145 -152
rect -119 -178 -79 -152
rect -53 -178 -13 -152
rect 13 -178 53 -152
rect 79 -178 119 -152
rect 145 -178 185 -152
rect 211 -178 251 -152
rect 277 -178 317 -152
rect 343 -178 383 -152
rect 409 -178 449 -152
rect 475 -178 515 -152
rect 541 -178 581 -152
rect 607 -178 647 -152
rect 673 -178 679 -152
rect -679 -218 679 -178
rect -679 -244 -673 -218
rect -647 -244 -607 -218
rect -581 -244 -541 -218
rect -515 -244 -475 -218
rect -449 -244 -409 -218
rect -383 -244 -343 -218
rect -317 -244 -277 -218
rect -251 -244 -211 -218
rect -185 -244 -145 -218
rect -119 -244 -79 -218
rect -53 -244 -13 -218
rect 13 -244 53 -218
rect 79 -244 119 -218
rect 145 -244 185 -218
rect 211 -244 251 -218
rect 277 -244 317 -218
rect 343 -244 383 -218
rect 409 -244 449 -218
rect 475 -244 515 -218
rect 541 -244 581 -218
rect 607 -244 647 -218
rect 673 -244 679 -218
rect -679 -284 679 -244
rect -679 -310 -673 -284
rect -647 -310 -607 -284
rect -581 -310 -541 -284
rect -515 -310 -475 -284
rect -449 -310 -409 -284
rect -383 -310 -343 -284
rect -317 -310 -277 -284
rect -251 -310 -211 -284
rect -185 -310 -145 -284
rect -119 -310 -79 -284
rect -53 -310 -13 -284
rect 13 -310 53 -284
rect 79 -310 119 -284
rect 145 -310 185 -284
rect 211 -310 251 -284
rect 277 -310 317 -284
rect 343 -310 383 -284
rect 409 -310 449 -284
rect 475 -310 515 -284
rect 541 -310 581 -284
rect 607 -310 647 -284
rect 673 -310 679 -284
rect -679 -316 679 -310
<< end >>
