magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2128 -2739 2128 2739
<< nwell >>
rect -128 -739 128 739
<< nsubdiff >>
rect -45 634 45 656
rect -45 -634 -23 634
rect 23 -634 45 634
rect -45 -656 45 -634
<< nsubdiffcont >>
rect -23 -634 23 634
<< metal1 >>
rect -34 634 34 645
rect -34 -634 -23 634
rect 23 -634 34 634
rect -34 -645 34 -634
<< end >>
