magic
tech gf180mcuC
magscale 1 10
timestamp 1691266842
<< error_p >>
rect -503 -48 -457 48
rect -343 -48 -297 48
rect -183 -48 -137 48
rect -23 -48 23 48
rect 137 -48 183 48
rect 297 -48 343 48
rect 457 -48 503 48
<< pwell >>
rect -540 -118 540 118
<< nmos >>
rect -428 -50 -372 50
rect -268 -50 -212 50
rect -108 -50 -52 50
rect 52 -50 108 50
rect 212 -50 268 50
rect 372 -50 428 50
<< ndiff >>
rect -516 37 -428 50
rect -516 -37 -503 37
rect -457 -37 -428 37
rect -516 -50 -428 -37
rect -372 37 -268 50
rect -372 -37 -343 37
rect -297 -37 -268 37
rect -372 -50 -268 -37
rect -212 37 -108 50
rect -212 -37 -183 37
rect -137 -37 -108 37
rect -212 -50 -108 -37
rect -52 37 52 50
rect -52 -37 -23 37
rect 23 -37 52 37
rect -52 -50 52 -37
rect 108 37 212 50
rect 108 -37 137 37
rect 183 -37 212 37
rect 108 -50 212 -37
rect 268 37 372 50
rect 268 -37 297 37
rect 343 -37 372 37
rect 268 -50 372 -37
rect 428 37 516 50
rect 428 -37 457 37
rect 503 -37 516 37
rect 428 -50 516 -37
<< ndiffc >>
rect -503 -37 -457 37
rect -343 -37 -297 37
rect -183 -37 -137 37
rect -23 -37 23 37
rect 137 -37 183 37
rect 297 -37 343 37
rect 457 -37 503 37
<< polysilicon >>
rect -428 50 -372 94
rect -268 50 -212 94
rect -108 50 -52 94
rect 52 50 108 94
rect 212 50 268 94
rect 372 50 428 94
rect -428 -94 -372 -50
rect -268 -94 -212 -50
rect -108 -94 -52 -50
rect 52 -94 108 -50
rect 212 -94 268 -50
rect 372 -94 428 -50
<< metal1 >>
rect -503 37 -457 48
rect -503 -48 -457 -37
rect -343 37 -297 48
rect -343 -48 -297 -37
rect -183 37 -137 48
rect -183 -48 -137 -37
rect -23 37 23 48
rect -23 -48 23 -37
rect 137 37 183 48
rect 137 -48 183 -37
rect 297 37 343 48
rect 297 -48 343 -37
rect 457 37 503 48
rect 457 -48 503 -37
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 0.5 l 0.280 m 1 nf 6 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
