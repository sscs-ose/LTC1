magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2278 -4578 2278 4578
<< nwell >>
rect -278 -2578 278 2578
<< nsubdiff >>
rect -195 2473 195 2495
rect -195 -2473 -173 2473
rect 173 -2473 195 2473
rect -195 -2495 195 -2473
<< nsubdiffcont >>
rect -173 -2473 173 2473
<< metal1 >>
rect -184 2473 184 2484
rect -184 -2473 -173 2473
rect 173 -2473 184 2473
rect -184 -2484 184 -2473
<< end >>
