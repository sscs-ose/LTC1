* NGSPICE file created from CM_magic_flat.ext - technology: gf180mcuC

.subckt pex_CM_magic OUT ITAIL  VSS 
X0 a_212_68# ITAIL.t2 OUT.t0 VSS.t5 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X1 a_212_n254# ITAIL.t0 ITAIL.t1 VSS.t5 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X2 VSS a_212_n254# a_212_68# VSS.t0 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X3 VSS a_212_n254# a_212_n254# VSS.t0 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
R0 ITAIL.n0 ITAIL.t0 12.1185
R1 ITAIL.n0 ITAIL.t2 11.3885
R2 ITAIL.n1 ITAIL.n0 7.97734
R3 ITAIL.n1 ITAIL.t1 6.12613
R4 ITAIL ITAIL.n1 0.267833
R5 OUT OUT.t0 6.1505
R6 VSS.n3 VSS.t5 429.322
R7 VSS.n3 VSS.t0 389.199
R8 VSS.n2 VSS.n0 6.47193
R9 VSS.n2 VSS.n1 5.8805
R10 VSS.n6 VSS.n5 2.6005
R11 VSS.n5 VSS.n3 2.6005
R12 VSS.n5 VSS.n4 1.19368
R13 VSS.n6 VSS.n2 0.510276
R14 VSS VSS.n6 0.0138663
C0 ITAIL a_212_n254# 0.14f
C1 a_212_68# OUT 0.0401f
C2 OUT ITAIL 0.0602f
C3 a_212_68# ITAIL 0.00862f
C4 OUT a_212_n254# 8.81e-19
C5 a_212_68# a_212_n254# 0.0536f
.ends

