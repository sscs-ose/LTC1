magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2752 -2544 2752 2544
<< nwell >>
rect -752 -544 752 544
<< nsubdiff >>
rect -669 439 669 461
rect -669 393 -647 439
rect -601 393 -543 439
rect -497 393 -439 439
rect -393 393 -335 439
rect -289 393 -231 439
rect -185 393 -127 439
rect -81 393 -23 439
rect 23 393 81 439
rect 127 393 185 439
rect 231 393 289 439
rect 335 393 393 439
rect 439 393 497 439
rect 543 393 601 439
rect 647 393 669 439
rect -669 335 669 393
rect -669 289 -647 335
rect -601 289 -543 335
rect -497 289 -439 335
rect -393 289 -335 335
rect -289 289 -231 335
rect -185 289 -127 335
rect -81 289 -23 335
rect 23 289 81 335
rect 127 289 185 335
rect 231 289 289 335
rect 335 289 393 335
rect 439 289 497 335
rect 543 289 601 335
rect 647 289 669 335
rect -669 231 669 289
rect -669 185 -647 231
rect -601 185 -543 231
rect -497 185 -439 231
rect -393 185 -335 231
rect -289 185 -231 231
rect -185 185 -127 231
rect -81 185 -23 231
rect 23 185 81 231
rect 127 185 185 231
rect 231 185 289 231
rect 335 185 393 231
rect 439 185 497 231
rect 543 185 601 231
rect 647 185 669 231
rect -669 127 669 185
rect -669 81 -647 127
rect -601 81 -543 127
rect -497 81 -439 127
rect -393 81 -335 127
rect -289 81 -231 127
rect -185 81 -127 127
rect -81 81 -23 127
rect 23 81 81 127
rect 127 81 185 127
rect 231 81 289 127
rect 335 81 393 127
rect 439 81 497 127
rect 543 81 601 127
rect 647 81 669 127
rect -669 23 669 81
rect -669 -23 -647 23
rect -601 -23 -543 23
rect -497 -23 -439 23
rect -393 -23 -335 23
rect -289 -23 -231 23
rect -185 -23 -127 23
rect -81 -23 -23 23
rect 23 -23 81 23
rect 127 -23 185 23
rect 231 -23 289 23
rect 335 -23 393 23
rect 439 -23 497 23
rect 543 -23 601 23
rect 647 -23 669 23
rect -669 -81 669 -23
rect -669 -127 -647 -81
rect -601 -127 -543 -81
rect -497 -127 -439 -81
rect -393 -127 -335 -81
rect -289 -127 -231 -81
rect -185 -127 -127 -81
rect -81 -127 -23 -81
rect 23 -127 81 -81
rect 127 -127 185 -81
rect 231 -127 289 -81
rect 335 -127 393 -81
rect 439 -127 497 -81
rect 543 -127 601 -81
rect 647 -127 669 -81
rect -669 -185 669 -127
rect -669 -231 -647 -185
rect -601 -231 -543 -185
rect -497 -231 -439 -185
rect -393 -231 -335 -185
rect -289 -231 -231 -185
rect -185 -231 -127 -185
rect -81 -231 -23 -185
rect 23 -231 81 -185
rect 127 -231 185 -185
rect 231 -231 289 -185
rect 335 -231 393 -185
rect 439 -231 497 -185
rect 543 -231 601 -185
rect 647 -231 669 -185
rect -669 -289 669 -231
rect -669 -335 -647 -289
rect -601 -335 -543 -289
rect -497 -335 -439 -289
rect -393 -335 -335 -289
rect -289 -335 -231 -289
rect -185 -335 -127 -289
rect -81 -335 -23 -289
rect 23 -335 81 -289
rect 127 -335 185 -289
rect 231 -335 289 -289
rect 335 -335 393 -289
rect 439 -335 497 -289
rect 543 -335 601 -289
rect 647 -335 669 -289
rect -669 -393 669 -335
rect -669 -439 -647 -393
rect -601 -439 -543 -393
rect -497 -439 -439 -393
rect -393 -439 -335 -393
rect -289 -439 -231 -393
rect -185 -439 -127 -393
rect -81 -439 -23 -393
rect 23 -439 81 -393
rect 127 -439 185 -393
rect 231 -439 289 -393
rect 335 -439 393 -393
rect 439 -439 497 -393
rect 543 -439 601 -393
rect 647 -439 669 -393
rect -669 -461 669 -439
<< nsubdiffcont >>
rect -647 393 -601 439
rect -543 393 -497 439
rect -439 393 -393 439
rect -335 393 -289 439
rect -231 393 -185 439
rect -127 393 -81 439
rect -23 393 23 439
rect 81 393 127 439
rect 185 393 231 439
rect 289 393 335 439
rect 393 393 439 439
rect 497 393 543 439
rect 601 393 647 439
rect -647 289 -601 335
rect -543 289 -497 335
rect -439 289 -393 335
rect -335 289 -289 335
rect -231 289 -185 335
rect -127 289 -81 335
rect -23 289 23 335
rect 81 289 127 335
rect 185 289 231 335
rect 289 289 335 335
rect 393 289 439 335
rect 497 289 543 335
rect 601 289 647 335
rect -647 185 -601 231
rect -543 185 -497 231
rect -439 185 -393 231
rect -335 185 -289 231
rect -231 185 -185 231
rect -127 185 -81 231
rect -23 185 23 231
rect 81 185 127 231
rect 185 185 231 231
rect 289 185 335 231
rect 393 185 439 231
rect 497 185 543 231
rect 601 185 647 231
rect -647 81 -601 127
rect -543 81 -497 127
rect -439 81 -393 127
rect -335 81 -289 127
rect -231 81 -185 127
rect -127 81 -81 127
rect -23 81 23 127
rect 81 81 127 127
rect 185 81 231 127
rect 289 81 335 127
rect 393 81 439 127
rect 497 81 543 127
rect 601 81 647 127
rect -647 -23 -601 23
rect -543 -23 -497 23
rect -439 -23 -393 23
rect -335 -23 -289 23
rect -231 -23 -185 23
rect -127 -23 -81 23
rect -23 -23 23 23
rect 81 -23 127 23
rect 185 -23 231 23
rect 289 -23 335 23
rect 393 -23 439 23
rect 497 -23 543 23
rect 601 -23 647 23
rect -647 -127 -601 -81
rect -543 -127 -497 -81
rect -439 -127 -393 -81
rect -335 -127 -289 -81
rect -231 -127 -185 -81
rect -127 -127 -81 -81
rect -23 -127 23 -81
rect 81 -127 127 -81
rect 185 -127 231 -81
rect 289 -127 335 -81
rect 393 -127 439 -81
rect 497 -127 543 -81
rect 601 -127 647 -81
rect -647 -231 -601 -185
rect -543 -231 -497 -185
rect -439 -231 -393 -185
rect -335 -231 -289 -185
rect -231 -231 -185 -185
rect -127 -231 -81 -185
rect -23 -231 23 -185
rect 81 -231 127 -185
rect 185 -231 231 -185
rect 289 -231 335 -185
rect 393 -231 439 -185
rect 497 -231 543 -185
rect 601 -231 647 -185
rect -647 -335 -601 -289
rect -543 -335 -497 -289
rect -439 -335 -393 -289
rect -335 -335 -289 -289
rect -231 -335 -185 -289
rect -127 -335 -81 -289
rect -23 -335 23 -289
rect 81 -335 127 -289
rect 185 -335 231 -289
rect 289 -335 335 -289
rect 393 -335 439 -289
rect 497 -335 543 -289
rect 601 -335 647 -289
rect -647 -439 -601 -393
rect -543 -439 -497 -393
rect -439 -439 -393 -393
rect -335 -439 -289 -393
rect -231 -439 -185 -393
rect -127 -439 -81 -393
rect -23 -439 23 -393
rect 81 -439 127 -393
rect 185 -439 231 -393
rect 289 -439 335 -393
rect 393 -439 439 -393
rect 497 -439 543 -393
rect 601 -439 647 -393
<< metal1 >>
rect -658 439 658 450
rect -658 393 -647 439
rect -601 393 -543 439
rect -497 393 -439 439
rect -393 393 -335 439
rect -289 393 -231 439
rect -185 393 -127 439
rect -81 393 -23 439
rect 23 393 81 439
rect 127 393 185 439
rect 231 393 289 439
rect 335 393 393 439
rect 439 393 497 439
rect 543 393 601 439
rect 647 393 658 439
rect -658 335 658 393
rect -658 289 -647 335
rect -601 289 -543 335
rect -497 289 -439 335
rect -393 289 -335 335
rect -289 289 -231 335
rect -185 289 -127 335
rect -81 289 -23 335
rect 23 289 81 335
rect 127 289 185 335
rect 231 289 289 335
rect 335 289 393 335
rect 439 289 497 335
rect 543 289 601 335
rect 647 289 658 335
rect -658 231 658 289
rect -658 185 -647 231
rect -601 185 -543 231
rect -497 185 -439 231
rect -393 185 -335 231
rect -289 185 -231 231
rect -185 185 -127 231
rect -81 185 -23 231
rect 23 185 81 231
rect 127 185 185 231
rect 231 185 289 231
rect 335 185 393 231
rect 439 185 497 231
rect 543 185 601 231
rect 647 185 658 231
rect -658 127 658 185
rect -658 81 -647 127
rect -601 81 -543 127
rect -497 81 -439 127
rect -393 81 -335 127
rect -289 81 -231 127
rect -185 81 -127 127
rect -81 81 -23 127
rect 23 81 81 127
rect 127 81 185 127
rect 231 81 289 127
rect 335 81 393 127
rect 439 81 497 127
rect 543 81 601 127
rect 647 81 658 127
rect -658 23 658 81
rect -658 -23 -647 23
rect -601 -23 -543 23
rect -497 -23 -439 23
rect -393 -23 -335 23
rect -289 -23 -231 23
rect -185 -23 -127 23
rect -81 -23 -23 23
rect 23 -23 81 23
rect 127 -23 185 23
rect 231 -23 289 23
rect 335 -23 393 23
rect 439 -23 497 23
rect 543 -23 601 23
rect 647 -23 658 23
rect -658 -81 658 -23
rect -658 -127 -647 -81
rect -601 -127 -543 -81
rect -497 -127 -439 -81
rect -393 -127 -335 -81
rect -289 -127 -231 -81
rect -185 -127 -127 -81
rect -81 -127 -23 -81
rect 23 -127 81 -81
rect 127 -127 185 -81
rect 231 -127 289 -81
rect 335 -127 393 -81
rect 439 -127 497 -81
rect 543 -127 601 -81
rect 647 -127 658 -81
rect -658 -185 658 -127
rect -658 -231 -647 -185
rect -601 -231 -543 -185
rect -497 -231 -439 -185
rect -393 -231 -335 -185
rect -289 -231 -231 -185
rect -185 -231 -127 -185
rect -81 -231 -23 -185
rect 23 -231 81 -185
rect 127 -231 185 -185
rect 231 -231 289 -185
rect 335 -231 393 -185
rect 439 -231 497 -185
rect 543 -231 601 -185
rect 647 -231 658 -185
rect -658 -289 658 -231
rect -658 -335 -647 -289
rect -601 -335 -543 -289
rect -497 -335 -439 -289
rect -393 -335 -335 -289
rect -289 -335 -231 -289
rect -185 -335 -127 -289
rect -81 -335 -23 -289
rect 23 -335 81 -289
rect 127 -335 185 -289
rect 231 -335 289 -289
rect 335 -335 393 -289
rect 439 -335 497 -289
rect 543 -335 601 -289
rect 647 -335 658 -289
rect -658 -393 658 -335
rect -658 -439 -647 -393
rect -601 -439 -543 -393
rect -497 -439 -439 -393
rect -393 -439 -335 -393
rect -289 -439 -231 -393
rect -185 -439 -127 -393
rect -81 -439 -23 -393
rect 23 -439 81 -393
rect 127 -439 185 -393
rect 231 -439 289 -393
rect 335 -439 393 -393
rect 439 -439 497 -393
rect 543 -439 601 -393
rect 647 -439 658 -393
rect -658 -450 658 -439
<< end >>
