magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2089 -2042 2089 2042
<< polysilicon >>
rect -89 23 89 42
rect -89 -23 -70 23
rect 70 -23 89 23
rect -89 -42 89 -23
<< polycontact >>
rect -70 -23 70 23
<< metal1 >>
rect -81 23 81 34
rect -81 -23 -70 23
rect 70 -23 81 23
rect -81 -34 81 -23
<< end >>
