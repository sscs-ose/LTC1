magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1050 -1732 1050 1732
<< metal2 >>
rect -50 727 50 732
rect -50 699 -45 727
rect -17 699 17 727
rect 45 699 50 727
rect -50 665 50 699
rect -50 637 -45 665
rect -17 637 17 665
rect 45 637 50 665
rect -50 603 50 637
rect -50 575 -45 603
rect -17 575 17 603
rect 45 575 50 603
rect -50 541 50 575
rect -50 513 -45 541
rect -17 513 17 541
rect 45 513 50 541
rect -50 479 50 513
rect -50 451 -45 479
rect -17 451 17 479
rect 45 451 50 479
rect -50 417 50 451
rect -50 389 -45 417
rect -17 389 17 417
rect 45 389 50 417
rect -50 355 50 389
rect -50 327 -45 355
rect -17 327 17 355
rect 45 327 50 355
rect -50 293 50 327
rect -50 265 -45 293
rect -17 265 17 293
rect 45 265 50 293
rect -50 231 50 265
rect -50 203 -45 231
rect -17 203 17 231
rect 45 203 50 231
rect -50 169 50 203
rect -50 141 -45 169
rect -17 141 17 169
rect 45 141 50 169
rect -50 107 50 141
rect -50 79 -45 107
rect -17 79 17 107
rect 45 79 50 107
rect -50 45 50 79
rect -50 17 -45 45
rect -17 17 17 45
rect 45 17 50 45
rect -50 -17 50 17
rect -50 -45 -45 -17
rect -17 -45 17 -17
rect 45 -45 50 -17
rect -50 -79 50 -45
rect -50 -107 -45 -79
rect -17 -107 17 -79
rect 45 -107 50 -79
rect -50 -141 50 -107
rect -50 -169 -45 -141
rect -17 -169 17 -141
rect 45 -169 50 -141
rect -50 -203 50 -169
rect -50 -231 -45 -203
rect -17 -231 17 -203
rect 45 -231 50 -203
rect -50 -265 50 -231
rect -50 -293 -45 -265
rect -17 -293 17 -265
rect 45 -293 50 -265
rect -50 -327 50 -293
rect -50 -355 -45 -327
rect -17 -355 17 -327
rect 45 -355 50 -327
rect -50 -389 50 -355
rect -50 -417 -45 -389
rect -17 -417 17 -389
rect 45 -417 50 -389
rect -50 -451 50 -417
rect -50 -479 -45 -451
rect -17 -479 17 -451
rect 45 -479 50 -451
rect -50 -513 50 -479
rect -50 -541 -45 -513
rect -17 -541 17 -513
rect 45 -541 50 -513
rect -50 -575 50 -541
rect -50 -603 -45 -575
rect -17 -603 17 -575
rect 45 -603 50 -575
rect -50 -637 50 -603
rect -50 -665 -45 -637
rect -17 -665 17 -637
rect 45 -665 50 -637
rect -50 -699 50 -665
rect -50 -727 -45 -699
rect -17 -727 17 -699
rect 45 -727 50 -699
rect -50 -732 50 -727
<< via2 >>
rect -45 699 -17 727
rect 17 699 45 727
rect -45 637 -17 665
rect 17 637 45 665
rect -45 575 -17 603
rect 17 575 45 603
rect -45 513 -17 541
rect 17 513 45 541
rect -45 451 -17 479
rect 17 451 45 479
rect -45 389 -17 417
rect 17 389 45 417
rect -45 327 -17 355
rect 17 327 45 355
rect -45 265 -17 293
rect 17 265 45 293
rect -45 203 -17 231
rect 17 203 45 231
rect -45 141 -17 169
rect 17 141 45 169
rect -45 79 -17 107
rect 17 79 45 107
rect -45 17 -17 45
rect 17 17 45 45
rect -45 -45 -17 -17
rect 17 -45 45 -17
rect -45 -107 -17 -79
rect 17 -107 45 -79
rect -45 -169 -17 -141
rect 17 -169 45 -141
rect -45 -231 -17 -203
rect 17 -231 45 -203
rect -45 -293 -17 -265
rect 17 -293 45 -265
rect -45 -355 -17 -327
rect 17 -355 45 -327
rect -45 -417 -17 -389
rect 17 -417 45 -389
rect -45 -479 -17 -451
rect 17 -479 45 -451
rect -45 -541 -17 -513
rect 17 -541 45 -513
rect -45 -603 -17 -575
rect 17 -603 45 -575
rect -45 -665 -17 -637
rect 17 -665 45 -637
rect -45 -727 -17 -699
rect 17 -727 45 -699
<< metal3 >>
rect -50 727 50 732
rect -50 699 -45 727
rect -17 699 17 727
rect 45 699 50 727
rect -50 665 50 699
rect -50 637 -45 665
rect -17 637 17 665
rect 45 637 50 665
rect -50 603 50 637
rect -50 575 -45 603
rect -17 575 17 603
rect 45 575 50 603
rect -50 541 50 575
rect -50 513 -45 541
rect -17 513 17 541
rect 45 513 50 541
rect -50 479 50 513
rect -50 451 -45 479
rect -17 451 17 479
rect 45 451 50 479
rect -50 417 50 451
rect -50 389 -45 417
rect -17 389 17 417
rect 45 389 50 417
rect -50 355 50 389
rect -50 327 -45 355
rect -17 327 17 355
rect 45 327 50 355
rect -50 293 50 327
rect -50 265 -45 293
rect -17 265 17 293
rect 45 265 50 293
rect -50 231 50 265
rect -50 203 -45 231
rect -17 203 17 231
rect 45 203 50 231
rect -50 169 50 203
rect -50 141 -45 169
rect -17 141 17 169
rect 45 141 50 169
rect -50 107 50 141
rect -50 79 -45 107
rect -17 79 17 107
rect 45 79 50 107
rect -50 45 50 79
rect -50 17 -45 45
rect -17 17 17 45
rect 45 17 50 45
rect -50 -17 50 17
rect -50 -45 -45 -17
rect -17 -45 17 -17
rect 45 -45 50 -17
rect -50 -79 50 -45
rect -50 -107 -45 -79
rect -17 -107 17 -79
rect 45 -107 50 -79
rect -50 -141 50 -107
rect -50 -169 -45 -141
rect -17 -169 17 -141
rect 45 -169 50 -141
rect -50 -203 50 -169
rect -50 -231 -45 -203
rect -17 -231 17 -203
rect 45 -231 50 -203
rect -50 -265 50 -231
rect -50 -293 -45 -265
rect -17 -293 17 -265
rect 45 -293 50 -265
rect -50 -327 50 -293
rect -50 -355 -45 -327
rect -17 -355 17 -327
rect 45 -355 50 -327
rect -50 -389 50 -355
rect -50 -417 -45 -389
rect -17 -417 17 -389
rect 45 -417 50 -389
rect -50 -451 50 -417
rect -50 -479 -45 -451
rect -17 -479 17 -451
rect 45 -479 50 -451
rect -50 -513 50 -479
rect -50 -541 -45 -513
rect -17 -541 17 -513
rect 45 -541 50 -513
rect -50 -575 50 -541
rect -50 -603 -45 -575
rect -17 -603 17 -575
rect 45 -603 50 -575
rect -50 -637 50 -603
rect -50 -665 -45 -637
rect -17 -665 17 -637
rect 45 -665 50 -637
rect -50 -699 50 -665
rect -50 -727 -45 -699
rect -17 -727 17 -699
rect 45 -727 50 -699
rect -50 -732 50 -727
<< end >>
