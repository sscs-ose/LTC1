* NGSPICE file created from BIASING_CURRENT_MAGIC.ext - technology: gf180mcuC

.subckt nfet_03v3_CT75PZ a_n52_n240# a_152_n240# a_52_n284# a_n152_n284# a_n240_n240#
+ VSUBS
X0 a_n52_n240# a_n152_n284# a_n240_n240# VSUBS nfet_03v3 ad=0.624p pd=2.92u as=1.06p ps=5.68u w=2.4u l=0.5u
X1 a_152_n240# a_52_n284# a_n52_n240# VSUBS nfet_03v3 ad=1.06p pd=5.68u as=0.624p ps=2.92u w=2.4u l=0.5u
.ends

.subckt nfet_03v3_CTB5PZ a_50_n240# a_n50_n284# a_n138_n240# VSUBS
X0 a_50_n240# a_n50_n284# a_n138_n240# VSUBS nfet_03v3 ad=1.06p pd=5.68u as=1.06p ps=5.68u w=2.4u l=0.5u
.ends

.subckt BIASING_CURRENT_MAGIC IBIAS_BUF1 IBIAS_BUF2 IBIAS_FILTER IBIAS_PGA G_SINK_UP
+ G_SINK_DOWN VSS
Xnfet_03v3_CT75PZ_1 m1_1867_n835# IBIAS_PGA G_SINK_UP G_SINK_UP IBIAS_PGA VSS nfet_03v3_CT75PZ
Xnfet_03v3_CT75PZ_0 m1_1867_n835# VSS G_SINK_DOWN G_SINK_DOWN VSS VSS nfet_03v3_CT75PZ
Xnfet_03v3_CT75PZ_2 m1_214_n835# IBIAS_BUF1 G_SINK_UP G_SINK_UP IBIAS_BUF1 VSS nfet_03v3_CT75PZ
Xnfet_03v3_CT75PZ_3 m1_214_n835# VSS G_SINK_DOWN G_SINK_DOWN VSS VSS nfet_03v3_CT75PZ
Xnfet_03v3_CT75PZ_4 m1_765_n835# VSS G_SINK_DOWN G_SINK_DOWN VSS VSS nfet_03v3_CT75PZ
Xnfet_03v3_CT75PZ_5 m1_765_n835# IBIAS_BUF2 G_SINK_UP G_SINK_UP IBIAS_BUF2 VSS nfet_03v3_CT75PZ
Xnfet_03v3_CT75PZ_6 m1_1316_n835# VSS G_SINK_DOWN G_SINK_DOWN VSS VSS nfet_03v3_CT75PZ
Xnfet_03v3_CT75PZ_7 m1_1316_n835# IBIAS_FILTER G_SINK_UP G_SINK_UP IBIAS_FILTER VSS
+ nfet_03v3_CT75PZ
Xnfet_03v3_CTB5PZ_0 VSS VSS VSS VSS nfet_03v3_CTB5PZ
Xnfet_03v3_CTB5PZ_1 VSS VSS VSS VSS nfet_03v3_CTB5PZ
Xnfet_03v3_CTB5PZ_2 VSS VSS VSS VSS nfet_03v3_CTB5PZ
Xnfet_03v3_CTB5PZ_3 VSS VSS VSS VSS nfet_03v3_CTB5PZ
.ends

