* NGSPICE file created from VCO_DFF_C_flat.ext - technology: gf180mcuC

.subckt pex_VCO_DFF_C VDD VSS VCTRL VCTRL2 OUT OUTB 
X0 VDD VCO_C_0.INV_2_3.IN.t30 VCO_C_0.INV_2_2.IN.t6 VDD.t29 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X1 VDD VCTRL.t0 VCO_C_0.INV_2_3.IN.t26 VDD.t199 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X2 VDD VCO_C_0.INV_2_2.IN.t31 VCO_C_0.INV_2_3.IN.t17 VDD.t23 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X3 VDD VCO_C_0.INV_2_2.IN.t32 VCO_C_0.INV_2_3.IN.t16 VDD.t2 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X4 VSS.t361 VSS.t359 VSS.t361 VSS.t360 nfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X5 VCO_C_0.OUTB VCO_C_0.INV_2_1.IN.t12 VSS.t67 VSS.t66 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X6 VCO_C_0.INV_2_5.OUT VCO_C_0.INV_2_5.IN.t31 VDD.t338 VDD.t142 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X7 DFF_3_mag_0.INV_2_1.IN a_17597_1404.t6 DFF_3_mag_0.INV_2_5.OUT.t19 VDD.t56 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X8 VCO_C_0.INV_2_1.IN VCO_C_0.INV_2_3.IN.t31 VDD.t45 VDD.t43 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X9 VSS.t358 VSS.t357 VSS.t358 VSS.t293 nfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X10 VSS.t356 VSS.t354 VSS.t356 VSS.t355 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X11 VDD VCO_C_0.INV_2_4.IN.t12 VCO_C_0.OUT.t7 VDD.t93 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X12 VDD VCO_C_0.INV_2_5.IN.t32 VCO_C_0.INV_2_0.IN.t30 VDD.t136 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X13 VDD DFF_3_mag_0.INV_2_5.IN.t20 DFF_3_mag_0.INV_2_5.OUT.t11 VDD.t169 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X14 VCO_C_0.INV_2_1.IN VCO_C_0.INV_2_3.IN.t32 VDD.t44 VDD.t43 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X15 VCO_C_0.INV_2_3.IN VCO_C_0.INV_2_2.IN.t33 VDD.t289 VDD.t0 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X16 VSS.t353 VSS.t352 VSS.t353 VSS.t296 nfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X17 VCO_C_0.INV_2_0.IN VCO_C_0.INV_2_5.IN.t33 VDD.t350 VDD.t66 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X18 VDD VCO_C_0.INV_2_3.IN.t33 VCO_C_0.INV_2_2.IN.t7 VDD.t23 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X19 VCO_C_0.INV_2_5.IN VCTRL.t1 VDD.t393 VDD.t325 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X20 OUTB OUT.t12 VDD.t401 VDD.t119 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X21 VCO_C_0.INV_2_3.IN VCO_C_0.INV_2_5.OUT.t12 a_10161_4198.t11 VSS.t77 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X22 VCO_C_0.INV_2_0.IN VCO_C_0.INV_2_5.IN.t34 VDD.t351 VDD.t71 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X23 VDD OUT.t13 DFF_3_mag_0.INV_2_4.OUT.t11 VDD.t156 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X24 DFF_3_mag_0.INV_2_5.IN VCO_C_0.OUTB.t13 DFF_3_mag_0.INV_2_3.IN.t3 VSS.t217 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X25 DFF_3_mag_0.INV_2_1.IN VCO_C_0.OUTB.t14 DFF_3_mag_0.INV_2_5.OUT.t2 VSS.t30 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X26 DFF_3_mag_0.INV_2_4.OUT OUT.t14 VDD.t404 VDD.t161 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X27 DFF_3_mag_0.INV_2_1.IN a_17597_2884.t6 OUTB.t0 VDD.t56 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X28 VSS.t351 VSS.t349 VSS.t351 VSS.t350 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X29 DFF_3_mag_0.INV_2_3.IN a_20434_3437.t6 DFF_3_mag_0.INV_2_5.IN.t17 VDD.t132 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X30 DFF_3_mag_0.INV_2_5.OUT DFF_3_mag_0.INV_2_5.IN.t21 VSS.t92 VSS.t91 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X31 OUTB OUT.t15 VDD.t405 VDD.t48 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X32 VCO_C_0.INV_2_0.OUT VCO_C_0.INV_2_0.IN.t31 VDD.t296 VDD.t101 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X33 VDD OUT.t16 DFF_3_mag_0.INV_2_4.OUT.t9 VDD.t163 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X34 VSS.t348 VSS.t347 VSS.t348 VSS.t329 nfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X35 DFF_3_mag_0.INV_2_3.IN a_20434_1083.t6 DFF_3_mag_0.INV_2_4.OUT.t3 VDD.t123 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X36 VCO_C_0.INV_2_5.IN VCO_C_0.INV_2_0.IN.t32 VDD.t297 VDD.t66 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X37 VSS VCTRL2.t3 a_10161_4198.t58 VSS.t7 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X38 VCO_C_0.INV_2_3.IN VCO_C_0.INV_2_2.IN.t34 VDD.t288 VDD.t18 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X39 VCO_C_0.INV_2_3.IN VCTRL.t2 VDD.t394 VDD.t199 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X40 DFF_3_mag_0.INV_2_3.IN VCO_C_0.OUTB.t15 DFF_3_mag_0.INV_2_5.IN.t3 VSS.t27 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X41 DFF_3_mag_0.INV_2_0.OUT VCO_C_0.OUTB.t16 VSS.t29 VSS.t28 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X42 VCO_C_0.INV_2_5.OUT VCO_C_0.INV_2_5.IN.t35 VSS.t135 VSS.t129 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X43 VDD.t251 VDD.t249 VDD.t251 VDD.t250 pfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X44 VSS VCTRL2.t6 a_10161_4198.t32 VSS.t7 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X45 VDD.t248 VDD.t247 VDD.t248 VDD.t190 pfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X46 VSS.t346 VSS.t345 VSS.t346 VSS.t322 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X47 VSS VCTRL2.t8 a_1424_1033.t58 VSS.t172 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X48 VSS VCTRL2.t10 a_10161_4198.t34 VSS.t12 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X49 VDD.t246 VDD.t244 VDD.t246 VDD.t245 pfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X50 VDD OUT.t17 OUTB.t12 VDD.t113 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X51 VCO_C_0.INV_2_2.IN VCO_C_0.INV_2_3.IN.t34 VDD.t40 VDD.t18 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X52 VSS.t344 VSS.t342 VSS.t344 VSS.t343 nfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X53 DFF_3_mag_0.INV_2_5.IN DFF_3_mag_0.INV_2_1.IN.t16 VDD.t322 VDD.t320 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X54 DFF_3_mag_0.INV_2_1.IN VCO_C_0.OUTB.t17 DFF_3_mag_0.INV_2_5.OUT.t1 VSS.t30 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X55 VDD VCO_C_0.INV_2_3.IN.t35 VCO_C_0.INV_2_1.IN.t5 VDD.t26 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X56 VDD.t243 VDD.t242 VDD.t243 VDD.t205 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X57 VDD.t241 VDD.t240 VDD.t241 VDD.t202 pfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X58 VCO_C_0.INV_2_5.IN VCO_C_0.INV_2_0.IN.t33 VDD.t298 VDD.t145 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X59 VDD OUT.t18 OUTB.t11 VDD.t50 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X60 VDD VCO_C_0.OUTB.t18 a_20434_3437.t3 VDD.t53 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X61 VCO_C_0.OUTB VCO_C_0.INV_2_1.IN.t13 VDD.t80 VDD.t79 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X62 VSS.t341 VSS.t340 VSS.t341 VSS.t264 nfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X63 DFF_3_mag_0.INV_2_4.OUT a_20434_1083.t7 DFF_3_mag_0.INV_2_3.IN.t9 VDD.t127 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X64 VCO_C_0.INV_2_3.IN VCO_C_0.INV_2_2.IN.t35 VDD.t287 VDD.t16 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X65 VSS VCTRL2.t14 a_1424_1033.t54 VSS.t172 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X66 VDD.t239 VDD.t238 VDD.t239 VDD.t208 pfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X67 VCO_C_0.INV_2_1.IN VCO_C_0.INV_2_3.IN.t36 VSS.t37 VSS.t36 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X68 VSS VCO_C_0.OUTB.t20 a_17597_1404.t5 VSS.t31 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X69 OUTB OUT.t19 VSS.t80 VSS.t79 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X70 VCO_C_0.OUTB VCO_C_0.INV_2_1.IN.t14 VDD.t386 VDD.t385 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X71 VCO_C_0.INV_2_0.IN VCO_C_0.INV_2_5.IN.t36 VDD.t352 VDD.t145 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X72 VSS.t339 VSS.t338 VSS.t339 VSS.t264 nfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X73 VDD DFF_3_mag_0.INV_2_1.IN.t17 DFF_3_mag_0.INV_2_5.IN.t11 VDD.t317 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X74 VCO_C_0.INV_2_2.IN VCO_C_0.INV_2_3.IN.t37 VDD.t37 VDD.t16 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X75 VSS VCTRL2.t15 a_10161_4198.t22 VSS.t142 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X76 DFF_3_mag_0.INV_2_1.IN DFF_3_mag_0.INV_2_0.OUT.t12 OUTB.t5 VSS.t70 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X77 DFF_3_mag_0.INV_2_1.IN VCO_C_0.OUTB.t21 DFF_3_mag_0.INV_2_5.OUT.t0 VSS.t34 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X78 VCO_C_0.INV_2_0.OUT VCO_C_0.INV_2_0.IN.t34 VSS.t62 VSS.t61 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X79 VSS.t337 VSS.t336 VSS.t337 VSS.t296 nfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X80 VCO_C_0.INV_2_5.IN VCO_C_0.OUTB.t22 a_1424_1033.t8 VSS.t35 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X81 VDD DFF_3_mag_0.INV_2_5.IN.t22 DFF_3_mag_0.INV_2_5.OUT.t13 VDD.t84 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X82 VCO_C_0.INV_2_3.IN VCTRL.t3 VDD.t395 VDD.t330 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X83 VSS.t335 VSS.t333 VSS.t335 VSS.t334 nfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X84 OUT DFF_3_mag_0.INV_2_3.IN.t16 VDD.t414 VDD.t119 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X85 VSS DFF_3_mag_0.INV_2_1.IN.t18 DFF_3_mag_0.INV_2_5.IN.t16 VSS.t93 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X86 VDD VCO_C_0.OUTB.t23 DFF_3_mag_0.INV_2_0.OUT.t7 VDD.t180 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X87 VSS VCTRL2.t17 a_10161_4198.t23 VSS.t142 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X88 VDD VCO_C_0.INV_2_5.IN.t37 VCO_C_0.INV_2_0.IN.t26 VDD.t103 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X89 VDD.t237 VDD.t235 VDD.t237 VDD.t236 pfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X90 DFF_3_mag_0.INV_2_0.OUT VCO_C_0.OUTB.t24 VDD.t423 VDD.t58 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X91 VCO_C_0.INV_2_0.OUT VCO_C_0.INV_2_0.IN.t35 VDD.t102 VDD.t101 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X92 VSS OUT.t20 OUTB.t17 VSS.t81 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X93 VCO_C_0.INV_2_4.IN VCO_C_0.INV_2_2.IN.t36 VDD.t282 VDD.t268 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X94 VSS VCTRL2.t19 a_1424_1033.t51 VSS.t185 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X95 VSS VCO_C_0.INV_2_2.IN.t37 VCO_C_0.INV_2_4.IN.t11 VSS.t114 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X96 VDD VCO_C_0.INV_2_4.IN.t13 VCO_C_0.OUT.t6 VDD.t93 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X97 VDD DFF_3_mag_0.INV_2_0.OUT.t14 a_17597_2884.t4 VDD.t78 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X98 VDD VCO_C_0.INV_2_1.IN.t15 VCO_C_0.OUTB.t5 VDD.t61 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X99 VSS OUT.t21 OUTB.t16 VSS.t84 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X100 VCO_C_0.OUTB VCO_C_0.INV_2_1.IN.t16 VSS.t257 VSS.t256 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X101 VDD VCO_C_0.INV_2_0.IN.t36 VCO_C_0.INV_2_5.IN.t13 VDD.t103 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X102 VSS VCO_C_0.INV_2_2.IN.t38 VCO_C_0.INV_2_4.IN.t10 VSS.t111 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X103 VDD VCO_C_0.INV_2_5.IN.t38 VCO_C_0.INV_2_5.OUT.t6 VDD.t355 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X104 VDD.t234 VDD.t232 VDD.t234 VDD.t233 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X105 VCO_C_0.INV_2_5.OUT VCO_C_0.INV_2_5.IN.t39 VDD.t359 VDD.t358 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X106 VDD DFF_3_mag_0.INV_2_0.OUT.t15 a_20434_1083.t2 VDD.t127 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X107 VDD VCO_C_0.INV_2_4.IN.t14 VCO_C_0.OUT.t5 VDD.t96 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X108 VSS DFF_3_mag_0.INV_2_0.OUT.t16 a_17597_2884.t0 VSS.t40 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X109 VDD DFF_3_mag_0.INV_2_3.IN.t17 OUT.t5 VDD.t113 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X110 VCO_C_0.OUT VCO_C_0.INV_2_4.IN.t15 VDD.t155 VDD.t154 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X111 VDD VCO_C_0.INV_2_5.IN.t40 VCO_C_0.INV_2_0.IN.t25 VDD.t68 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X112 VSS DFF_3_mag_0.INV_2_0.OUT.t17 a_20434_1083.t0 VSS.t43 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X113 VDD VCO_C_0.INV_2_3.IN.t38 VCO_C_0.INV_2_1.IN.t4 VDD.t5 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X114 OUT DFF_3_mag_0.INV_2_3.IN.t18 VDD.t116 VDD.t48 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X115 VSS VCTRL2.t22 a_1424_1033.t49 VSS.t153 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X116 VCO_C_0.INV_2_0.IN VCO_C_0.OUT.t13 a_1424_1033.t18 VSS.t103 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X117 VDD DFF_3_mag_0.INV_2_3.IN.t19 OUT.t7 VDD.t50 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X118 VDD VCTRL.t4 VCO_C_0.INV_2_0.IN.t14 VDD.t245 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X119 VCO_C_0.INV_2_3.IN VCO_C_0.INV_2_5.OUT.t14 a_10161_4198.t59 VSS.t48 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X120 VSS VCO_C_0.INV_2_4.IN.t16 VCO_C_0.OUT.t11 VSS.t88 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X121 VCO_C_0.INV_2_0.OUT VCO_C_0.INV_2_0.IN.t37 VDD.t106 VDD.t64 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X122 DFF_3_mag_0.INV_2_3.IN a_20434_1083.t8 DFF_3_mag_0.INV_2_4.OUT.t17 VDD.t132 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X123 VSS VCTRL2.t24 a_1424_1033.t48 VSS.t153 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X124 DFF_3_mag_0.INV_2_5.IN a_20434_3437.t7 DFF_3_mag_0.INV_2_3.IN.t14 VDD.t53 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X125 VSS DFF_3_mag_0.INV_2_5.IN.t23 DFF_3_mag_0.INV_2_5.OUT.t14 VSS.t93 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X126 VCO_C_0.INV_2_0.IN VCO_C_0.OUT.t14 a_1424_1033.t17 VSS.t35 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X127 VCO_C_0.INV_2_2.IN VCO_C_0.INV_2_3.IN.t39 VDD.t34 VDD.t8 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X128 VDD.t231 VDD.t230 VDD.t231 VDD.t205 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X129 VCO_C_0.INV_2_5.IN VCO_C_0.INV_2_0.IN.t38 VDD.t107 VDD.t71 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X130 VDD VCTRL.t5 VCO_C_0.INV_2_0.IN.t13 VDD.t325 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X131 VDD VCO_C_0.INV_2_2.IN.t39 VCO_C_0.INV_2_3.IN.t15 VDD.t10 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X132 VSS.t332 VSS.t331 VSS.t332 VSS.t308 nfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X133 VCO_C_0.INV_2_3.IN VCO_C_0.INV_2_5.OUT.t15 a_10161_4198.t37 VSS.t77 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X134 DFF_3_mag_0.INV_2_0.OUT VCO_C_0.OUTB.t26 VSS.t371 VSS.t370 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X135 VCO_C_0.INV_2_5.OUT VCO_C_0.INV_2_5.IN.t41 VSS.t74 VSS.t61 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X136 DFF_3_mag_0.INV_2_1.IN a_17597_1404.t7 DFF_3_mag_0.INV_2_5.OUT.t18 VDD.t76 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X137 VCO_C_0.INV_2_2.IN VCO_C_0.INV_2_0.OUT.t15 a_10161_4198.t51 VSS.t77 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X138 VCO_C_0.INV_2_3.IN VCO_C_0.INV_2_2.IN.t40 VDD.t284 VDD.t8 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X139 VSS VCTRL2.t26 a_10161_4198.t19 VSS.t12 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X140 VDD VCO_C_0.INV_2_3.IN.t40 VCO_C_0.INV_2_2.IN.t13 VDD.t10 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X141 DFF_3_mag_0.INV_2_5.OUT VCO_C_0.OUTB.t27 DFF_3_mag_0.INV_2_1.IN.t0 VSS.t31 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X142 VCO_C_0.OUTB VCO_C_0.INV_2_1.IN.t17 VDD.t89 VDD.t79 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X143 VCO_C_0.INV_2_2.IN VCO_C_0.INV_2_0.OUT.t16 a_10161_4198.t50 VSS.t48 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X144 OUT DFF_3_mag_0.INV_2_3.IN.t20 VSS.t69 VSS.t68 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X145 VSS.t330 VSS.t328 VSS.t330 VSS.t329 nfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X146 VSS.t327 VSS.t326 VSS.t327 VSS.t78 nfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X147 VDD DFF_3_mag_0.INV_2_1.IN.t19 DFF_3_mag_0.INV_2_5.IN.t10 VDD.t180 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X148 VSS.t325 VSS.t324 VSS.t325 VSS.t267 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X149 VSS.t323 VSS.t321 VSS.t323 VSS.t322 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X150 DFF_3_mag_0.INV_2_1.IN a_17597_2884.t7 OUTB.t1 VDD.t76 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X151 VSS VCTRL2.t29 a_10161_4198.t21 VSS.t12 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X152 VDD VCO_C_0.INV_2_0.IN.t39 VCO_C_0.INV_2_5.IN.t15 VDD.t108 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X153 VSS VCTRL2.t30 a_1424_1033.t45 VSS.t172 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X154 VCO_C_0.INV_2_5.IN VCO_C_0.INV_2_0.IN.t40 VDD.t112 VDD.t111 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X155 VSS VCO_C_0.INV_2_3.IN.t41 VCO_C_0.INV_2_1.IN.t10 VSS.t136 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X156 VDD VCO_C_0.INV_2_2.IN.t41 VCO_C_0.INV_2_4.IN.t6 VDD.t259 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X157 VCO_C_0.INV_2_0.IN VCTRL.t6 VDD.t400 VDD.t325 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X158 VDD.t229 VDD.t227 VDD.t229 VDD.t228 pfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X159 VCO_C_0.INV_2_5.IN VCO_C_0.OUTB.t31 a_1424_1033.t5 VSS.t103 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X160 VDD VCTRL.t7 VCO_C_0.INV_2_2.IN.t14 VDD.t199 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X161 VSS.t320 VSS.t319 VSS.t320 VSS.t264 nfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X162 VDD VCO_C_0.INV_2_2.IN.t42 VCO_C_0.INV_2_4.IN.t5 VDD.t254 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X163 VSS VCTRL2.t33 a_10161_4198.t15 VSS.t142 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X164 VSS.t318 VSS.t317 VSS.t318 VSS.t296 nfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X165 VSS VCO_C_0.INV_2_0.IN.t41 VCO_C_0.INV_2_0.OUT.t0 VSS.t49 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X166 VDD VCO_C_0.INV_2_3.IN.t42 VCO_C_0.INV_2_2.IN.t1 VDD.t29 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X167 VCO_C_0.INV_2_2.IN VCO_C_0.INV_2_0.OUT.t17 a_10161_4198.t49 VSS.t77 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X168 DFF_3_mag_0.INV_2_5.IN DFF_3_mag_0.INV_2_1.IN.t20 VDD.t337 VDD.t58 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X169 VDD DFF_3_mag_0.INV_2_5.IN.t24 DFF_3_mag_0.INV_2_5.OUT.t15 VDD.t169 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X170 VSS VCTRL2.t34 a_10161_4198.t16 VSS.t142 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X171 VSS DFF_3_mag_0.INV_2_1.IN.t21 DFF_3_mag_0.INV_2_5.IN.t15 VSS.t55 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X172 VDD VCO_C_0.OUTB.t32 DFF_3_mag_0.INV_2_0.OUT.t5 VDD.t317 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X173 VSS VCTRL2.t35 a_1424_1033.t43 VSS.t147 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X174 VDD.t226 VDD.t224 VDD.t226 VDD.t225 pfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X175 VSS VCTRL2.t36 a_10161_4198.t17 VSS.t150 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X176 DFF_3_mag_0.INV_2_0.OUT VCO_C_0.OUTB.t33 VDD.t346 VDD.t320 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X177 VSS.t316 VSS.t315 VSS.t316 VSS.t296 nfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X178 VCO_C_0.INV_2_0.OUT VCO_C_0.INV_2_0.IN.t42 VDD.t65 VDD.t64 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X179 VDD VCO_C_0.INV_2_2.IN.t43 VCO_C_0.INV_2_3.IN.t14 VDD.t29 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X180 VSS.t314 VSS.t312 VSS.t314 VSS.t313 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X181 DFF_3_mag_0.INV_2_4.OUT DFF_3_mag_0.INV_2_0.OUT.t21 DFF_3_mag_0.INV_2_3.IN.t6 VSS.t59 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X182 VCO_C_0.INV_2_4.IN VCO_C_0.INV_2_2.IN.t44 VDD.t276 VDD.t262 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X183 DFF_3_mag_0.INV_2_4.OUT OUT.t22 VSS.t87 VSS.t68 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X184 VSS VCTRL2.t37 a_1424_1033.t42 VSS.t153 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X185 VDD VCO_C_0.INV_2_1.IN.t18 VCO_C_0.OUTB.t3 VDD.t387 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X186 VDD VCO_C_0.INV_2_4.IN.t17 VCO_C_0.OUT.t3 VDD.t96 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X187 VSS VCTRL2.t38 a_1424_1033.t41 VSS.t147 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X188 DFF_3_mag_0.INV_2_4.OUT OUT.t23 VDD.t151 VDD.t150 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X189 VDD VCTRL.t8 VCO_C_0.INV_2_2.IN.t15 VDD.t330 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X190 VCO_C_0.OUT VCO_C_0.INV_2_4.IN.t18 VDD.t301 VDD.t154 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X191 VDD VCTRL.t9 VCO_C_0.INV_2_5.IN.t20 VDD.t245 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.84u
X192 OUTB OUT.t24 VDD.t152 VDD.t119 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X193 VDD VCO_C_0.INV_2_5.IN.t42 VCO_C_0.INV_2_0.IN.t24 VDD.t136 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X194 VCO_C_0.INV_2_3.IN VCTRL.t10 VDD.t368 VDD.t199 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.84u
X195 VDD VCO_C_0.INV_2_5.IN.t43 VCO_C_0.INV_2_5.OUT.t4 VDD.t139 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X196 VDD.t223 VDD.t222 VDD.t223 VDD.t208 pfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X197 VCO_C_0.INV_2_4.IN VCO_C_0.INV_2_2.IN.t45 VSS.t110 VSS.t109 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X198 VSS VCTRL2.t39 a_1424_1033.t40 VSS.t153 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X199 VCO_C_0.INV_2_5.OUT VCO_C_0.INV_2_5.IN.t44 VDD.t143 VDD.t142 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X200 DFF_3_mag_0.INV_2_5.OUT a_17597_1404.t8 DFF_3_mag_0.INV_2_1.IN.t13 VDD.t77 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X201 VDD VCO_C_0.INV_2_2.IN.t46 VCO_C_0.INV_2_3.IN.t13 VDD.t2 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X202 VCO_C_0.OUT VCO_C_0.INV_2_4.IN.t19 VDD.t302 VDD.t294 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X203 VDD VCO_C_0.INV_2_3.IN.t43 VCO_C_0.INV_2_1.IN.t3 VDD.t26 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X204 VDD.t221 VDD.t219 VDD.t221 VDD.t220 pfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X205 VDD.t218 VDD.t216 VDD.t218 VDD.t217 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X206 VCO_C_0.INV_2_5.IN VCO_C_0.INV_2_0.IN.t43 VDD.t67 VDD.t66 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X207 VCO_C_0.INV_2_5.IN VCO_C_0.OUTB.t35 a_1424_1033.t4 VSS.t35 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X208 VCO_C_0.INV_2_0.IN VCO_C_0.OUT.t15 a_1424_1033.t16 VSS.t35 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X209 VCO_C_0.INV_2_3.IN VCO_C_0.INV_2_2.IN.t47 VDD.t273 VDD.t0 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X210 VDD VCO_C_0.INV_2_3.IN.t44 VCO_C_0.INV_2_2.IN.t8 VDD.t23 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X211 VSS VCO_C_0.INV_2_4.IN.t20 VCO_C_0.OUT.t10 VSS.t119 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X212 VDD VCO_C_0.INV_2_3.IN.t45 VCO_C_0.INV_2_2.IN.t9 VDD.t2 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X213 VDD OUT.t25 DFF_3_mag_0.INV_2_4.OUT.t7 VDD.t156 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X214 VDD.t215 VDD.t213 VDD.t215 VDD.t214 pfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X215 VSS DFF_3_mag_0.INV_2_5.IN.t25 DFF_3_mag_0.INV_2_5.OUT.t4 VSS.t55 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X216 VCO_C_0.OUT VCO_C_0.INV_2_4.IN.t21 VSS.t64 VSS.t63 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X217 VDD VCO_C_0.INV_2_0.IN.t44 VCO_C_0.INV_2_5.IN.t11 VDD.t68 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X218 VCO_C_0.INV_2_5.IN VCO_C_0.INV_2_0.IN.t45 VDD.t72 VDD.t71 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X219 VDD OUT.t26 OUTB.t9 VDD.t113 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X220 VSS.t311 VSS.t310 VSS.t311 VSS.t293 nfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X221 OUTB a_17597_2884.t8 DFF_3_mag_0.INV_2_1.IN.t6 VDD.t77 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X222 DFF_3_mag_0.INV_2_4.OUT OUT.t27 VDD.t162 VDD.t161 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X223 VDD VCO_C_0.INV_2_0.IN.t46 VCO_C_0.INV_2_0.OUT.t2 VDD.t73 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X224 DFF_3_mag_0.INV_2_4.OUT a_20434_1083.t9 DFF_3_mag_0.INV_2_3.IN.t11 VDD.t53 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X225 VCO_C_0.INV_2_2.IN VCTRL.t11 VDD.t369 VDD.t330 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X226 VDD OUT.t28 DFF_3_mag_0.INV_2_4.OUT.t5 VDD.t163 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X227 VDD.t212 VDD.t210 VDD.t212 VDD.t211 pfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X228 VCO_C_0.INV_2_2.IN VCO_C_0.INV_2_3.IN.t46 VDD.t20 VDD.t0 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X229 VDD OUT.t29 OUTB.t8 VDD.t50 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X230 VDD VCO_C_0.INV_2_2.IN.t48 VCO_C_0.INV_2_3.IN.t12 VDD.t23 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X231 VSS VCO_C_0.OUTB.t36 DFF_3_mag_0.INV_2_0.OUT.t9 VSS.t131 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X232 VCO_C_0.INV_2_0.IN VCO_C_0.OUT.t17 a_1424_1033.t14 VSS.t103 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X233 VCO_C_0.INV_2_0.IN VCO_C_0.INV_2_5.IN.t45 VDD.t144 VDD.t71 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X234 VSS VCTRL2.t44 a_10161_4198.t3 VSS.t7 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X235 VSS VCO_C_0.INV_2_5.IN.t46 VCO_C_0.INV_2_5.OUT.t9 VSS.t49 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X236 VSS VCTRL2.t46 a_10161_4198.t5 VSS.t12 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X237 DFF_3_mag_0.INV_2_5.IN VCO_C_0.OUTB.t37 DFF_3_mag_0.INV_2_3.IN.t1 VSS.t134 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X238 VSS.t309 VSS.t307 VSS.t309 VSS.t308 nfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X239 VCO_C_0.INV_2_5.IN VCO_C_0.OUTB.t38 a_1424_1033.t3 VSS.t35 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X240 VCO_C_0.INV_2_0.IN VCTRL.t12 VDD.t370 VDD.t245 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X241 VSS.t306 VSS.t305 VSS.t306 VSS.t293 nfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X242 VDD DFF_3_mag_0.INV_2_1.IN.t22 DFF_3_mag_0.INV_2_5.IN.t8 VDD.t317 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X243 VSS.t304 VSS.t303 VSS.t304 VSS.t264 nfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X244 OUTB OUT.t30 VDD.t168 VDD.t48 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X245 VCO_C_0.INV_2_0.IN VCO_C_0.INV_2_5.IN.t47 VDD.t146 VDD.t145 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X246 VSS VCTRL2.t48 a_10161_4198.t7 VSS.t12 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X247 VDD VCO_C_0.INV_2_1.IN.t19 VCO_C_0.OUTB.t2 VDD.t387 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X248 VCO_C_0.INV_2_2.IN VCO_C_0.INV_2_3.IN.t47 VDD.t19 VDD.t18 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X249 VSS VCTRL2.t50 a_1424_1033.t38 VSS.t147 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X250 VCO_C_0.INV_2_5.IN VCO_C_0.OUTB.t40 a_1424_1033.t1 VSS.t103 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X251 VDD.t209 VDD.t207 VDD.t209 VDD.t208 pfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X252 VSS VCO_C_0.INV_2_3.IN.t48 VCO_C_0.INV_2_1.IN.t9 VSS.t375 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X253 VCO_C_0.INV_2_2.IN VCO_C_0.INV_2_0.OUT.t19 a_10161_4198.t47 VSS.t48 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X254 VDD VCO_C_0.OUTB.t42 a_17597_1404.t1 VDD.t77 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X255 VDD VCO_C_0.INV_2_1.IN.t20 VCO_C_0.OUTB.t1 VDD.t61 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X256 VCO_C_0.INV_2_3.IN VCO_C_0.INV_2_5.OUT.t18 a_10161_4198.t8 VSS.t48 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X257 VCO_C_0.INV_2_3.IN VCO_C_0.INV_2_2.IN.t49 VDD.t270 VDD.t18 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X258 VDD VCO_C_0.INV_2_5.IN.t48 VCO_C_0.INV_2_0.IN.t21 VDD.t108 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X259 VSS.t302 VSS.t301 VSS.t302 VSS.t78 nfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X260 DFF_3_mag_0.INV_2_1.IN DFF_3_mag_0.INV_2_0.OUT.t22 OUTB.t6 VSS.t70 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X261 VSS VCTRL2.t53 a_1424_1033.t35 VSS.t147 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X262 VCO_C_0.INV_2_0.IN VCO_C_0.INV_2_5.IN.t49 VDD.t149 VDD.t111 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X263 VSS.t300 VSS.t298 VSS.t300 VSS.t299 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X264 VCO_C_0.INV_2_4.IN VCO_C_0.INV_2_2.IN.t50 VDD.t269 VDD.t268 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X265 VSS VCO_C_0.INV_2_0.IN.t47 VCO_C_0.INV_2_0.OUT.t3 VSS.t52 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X266 VDD.t206 VDD.t204 VDD.t206 VDD.t205 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X267 VSS.t297 VSS.t295 VSS.t297 VSS.t296 nfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X268 VCO_C_0.INV_2_2.IN VCO_C_0.INV_2_3.IN.t49 VDD.t17 VDD.t16 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X269 DFF_3_mag_0.INV_2_5.IN DFF_3_mag_0.INV_2_1.IN.t23 VDD.t321 VDD.t320 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X270 VDD.t203 VDD.t201 VDD.t203 VDD.t202 pfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X271 VDD DFF_3_mag_0.INV_2_0.OUT.t23 a_20434_1083.t4 VDD.t53 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X272 VSS VCTRL2.t57 a_10161_4198.t41 VSS.t150 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X273 VCO_C_0.INV_2_0.IN VCO_C_0.OUT.t19 a_1424_1033.t12 VSS.t103 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X274 VDD VCO_C_0.INV_2_0.IN.t48 VCO_C_0.INV_2_5.IN.t24 VDD.t103 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X275 OUT DFF_3_mag_0.INV_2_3.IN.t21 VDD.t120 VDD.t119 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X276 DFF_3_mag_0.INV_2_4.OUT DFF_3_mag_0.INV_2_0.OUT.t24 DFF_3_mag_0.INV_2_3.IN.t4 VSS.t43 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X277 VDD VCO_C_0.OUTB.t44 DFF_3_mag_0.INV_2_0.OUT.t3 VDD.t180 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X278 VDD VCO_C_0.INV_2_0.IN.t49 VCO_C_0.INV_2_0.OUT.t8 VDD.t73 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X279 DFF_3_mag_0.INV_2_5.OUT DFF_3_mag_0.INV_2_5.IN.t26 VDD.t82 VDD.t81 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X280 VDD.t200 VDD.t198 VDD.t200 VDD.t199 pfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X281 VDD VCO_C_0.OUTB.t45 a_20434_3437.t1 VDD.t127 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X282 VCO_C_0.INV_2_3.IN VCO_C_0.INV_2_2.IN.t51 VDD.t267 VDD.t16 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X283 DFF_3_mag_0.INV_2_5.IN DFF_3_mag_0.INV_2_1.IN.t24 VSS.t39 VSS.t38 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X284 DFF_3_mag_0.INV_2_0.OUT VCO_C_0.OUTB.t46 VDD.t185 VDD.t58 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X285 VCO_C_0.OUT VCO_C_0.INV_2_4.IN.t22 VDD.t295 VDD.t294 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X286 DFF_3_mag_0.INV_2_5.OUT DFF_3_mag_0.INV_2_5.IN.t27 VDD.t83 VDD.t81 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X287 VCO_C_0.INV_2_2.IN VCTRL.t13 VDD.t371 VDD.t199 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X288 VSS.t294 VSS.t292 VSS.t294 VSS.t293 nfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X289 VSS.t291 VSS.t289 VSS.t291 VSS.t290 nfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X290 VDD VCTRL.t14 VCO_C_0.INV_2_5.IN.t19 VDD.t325 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X291 OUTB OUT.t31 VSS.t97 VSS.t96 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X292 VSS VCTRL2.t58 a_10161_4198.t25 VSS.t150 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X293 VSS VCO_C_0.INV_2_1.IN.t21 VCO_C_0.OUTB.t9 VSS.t122 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X294 VCO_C_0.INV_2_4.IN VCO_C_0.INV_2_2.IN.t52 VSS.t108 VSS.t107 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X295 VDD.t197 VDD.t195 VDD.t197 VDD.t196 pfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X296 VSS VCTRL2.t59 a_1424_1033.t31 VSS.t153 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X297 VCO_C_0.INV_2_3.IN VCO_C_0.INV_2_5.OUT.t20 a_10161_4198.t9 VSS.t48 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X298 VSS VCO_C_0.INV_2_1.IN.t22 VCO_C_0.OUTB.t8 VSS.t71 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X299 VDD VCO_C_0.INV_2_5.IN.t50 VCO_C_0.INV_2_5.OUT.t2 VDD.t355 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X300 DFF_3_mag_0.INV_2_4.OUT DFF_3_mag_0.INV_2_0.OUT.t26 DFF_3_mag_0.INV_2_3.IN.t5 VSS.t59 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X301 VDD VCO_C_0.INV_2_0.IN.t50 VCO_C_0.INV_2_5.IN.t25 VDD.t136 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X302 OUTB DFF_3_mag_0.INV_2_0.OUT.t27 DFF_3_mag_0.INV_2_1.IN.t8 VSS.t40 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X303 VSS.t288 VSS.t287 VSS.t288 VSS.t78 nfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X304 VSS VCTRL2.t60 a_1424_1033.t30 VSS.t185 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X305 VCO_C_0.INV_2_5.OUT VCO_C_0.INV_2_5.IN.t51 VDD.t374 VDD.t358 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X306 VDD DFF_3_mag_0.INV_2_3.IN.t22 OUT.t10 VDD.t113 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X307 OUT DFF_3_mag_0.INV_2_3.IN.t23 VSS.t20 VSS.t19 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X308 DFF_3_mag_0.INV_2_5.IN VCO_C_0.OUTB.t47 DFF_3_mag_0.INV_2_3.IN.t0 VSS.t362 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X309 VSS.t286 VSS.t285 VSS.t286 VSS.t78 nfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X310 OUT DFF_3_mag_0.INV_2_3.IN.t24 VDD.t49 VDD.t48 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X311 VSS VCTRL2.t61 a_1424_1033.t29 VSS.t185 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X312 VDD VCO_C_0.INV_2_0.IN.t51 VCO_C_0.INV_2_5.IN.t26 VDD.t68 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X313 VCO_C_0.INV_2_1.IN VCO_C_0.INV_2_3.IN.t50 VDD.t15 VDD.t13 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X314 VCO_C_0.OUT VCO_C_0.INV_2_4.IN.t23 VSS.t118 VSS.t117 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X315 VDD DFF_3_mag_0.INV_2_3.IN.t25 OUT.t2 VDD.t50 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X316 VDD VCO_C_0.INV_2_0.IN.t52 VCO_C_0.INV_2_0.OUT.t9 VDD.t311 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X317 VCO_C_0.INV_2_0.IN VCO_C_0.INV_2_5.IN.t52 VDD.t375 VDD.t66 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X318 VSS VCO_C_0.OUTB.t48 DFF_3_mag_0.INV_2_0.OUT.t8 VSS.t363 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X319 VCO_C_0.INV_2_1.IN VCO_C_0.INV_2_3.IN.t51 VDD.t14 VDD.t13 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X320 VDD VCO_C_0.INV_2_5.IN.t53 VCO_C_0.INV_2_0.IN.t18 VDD.t68 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X321 DFF_3_mag_0.INV_2_3.IN a_20434_3437.t8 DFF_3_mag_0.INV_2_5.IN.t19 VDD.t123 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X322 DFF_3_mag_0.INV_2_5.OUT DFF_3_mag_0.INV_2_5.IN.t28 VSS.t58 VSS.t38 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X323 DFF_3_mag_0.INV_2_3.IN DFF_3_mag_0.INV_2_0.OUT.t29 DFF_3_mag_0.INV_2_4.OUT.t19 VSS.t125 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X324 VSS VCTRL2.t65 a_10161_4198.t28 VSS.t7 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X325 VSS VCO_C_0.INV_2_5.IN.t54 VCO_C_0.INV_2_5.OUT.t8 VSS.t52 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X326 DFF_3_mag_0.INV_2_5.OUT a_17597_1404.t9 DFF_3_mag_0.INV_2_1.IN.t12 VDD.t78 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X327 VDD DFF_3_mag_0.INV_2_5.IN.t29 DFF_3_mag_0.INV_2_5.OUT.t8 VDD.t84 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X328 VDD.t194 VDD.t192 VDD.t194 VDD.t193 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X329 VSS.t284 VSS.t282 VSS.t284 VSS.t283 nfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X330 VSS.t281 VSS.t280 VSS.t281 VSS.t275 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X331 VSS DFF_3_mag_0.INV_2_3.IN.t26 OUT.t3 VSS.t21 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X332 DFF_3_mag_0.INV_2_1.IN DFF_3_mag_0.INV_2_0.OUT.t30 OUTB.t19 VSS.t46 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X333 VDD.t191 VDD.t189 VDD.t191 VDD.t190 pfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X334 VCO_C_0.INV_2_3.IN VCO_C_0.INV_2_2.IN.t53 VDD.t266 VDD.t8 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X335 VSS.t279 VSS.t277 VSS.t279 VSS.t278 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X336 VDD VCO_C_0.INV_2_3.IN.t52 VCO_C_0.INV_2_2.IN.t4 VDD.t10 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X337 VSS VCTRL2.t69 a_10161_4198.t42 VSS.t7 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X338 VSS DFF_3_mag_0.INV_2_3.IN.t27 OUT.t4 VSS.t24 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X339 VSS VCO_C_0.OUTB.t49 a_20434_3437.t4 VSS.t366 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X340 VSS.t276 VSS.t274 VSS.t276 VSS.t275 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X341 OUTB a_17597_2884.t9 DFF_3_mag_0.INV_2_1.IN.t7 VDD.t78 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X342 VDD VCTRL.t15 VCO_C_0.INV_2_5.IN.t18 VDD.t245 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X343 DFF_3_mag_0.INV_2_5.IN DFF_3_mag_0.INV_2_1.IN.t25 VDD.t59 VDD.t58 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X344 DFF_3_mag_0.INV_2_4.OUT OUT.t32 VSS.t98 VSS.t19 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X345 VSS.t273 VSS.t272 VSS.t273 VSS.t270 nfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X346 VCO_C_0.INV_2_2.IN VCO_C_0.INV_2_3.IN.t53 VDD.t9 VDD.t8 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X347 VDD VCTRL.t16 VCO_C_0.INV_2_3.IN VDD.t330 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X348 DFF_3_mag_0.INV_2_5.IN a_20434_3437.t9 DFF_3_mag_0.INV_2_3.IN.t7 VDD.t127 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X349 VCO_C_0.OUTB VCO_C_0.INV_2_1.IN.t23 VDD.t390 VDD.t385 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X350 VDD VCO_C_0.INV_2_2.IN.t54 VCO_C_0.INV_2_3.IN.t11 VDD.t10 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X351 VCO_C_0.INV_2_5.IN VCO_C_0.INV_2_0.IN.t53 VDD.t314 VDD.t145 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X352 VDD VCO_C_0.INV_2_5.IN.t55 VCO_C_0.INV_2_0.IN.t17 VDD.t108 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X353 VCO_C_0.INV_2_0.IN VCO_C_0.INV_2_5.IN.t56 VDD.t380 VDD.t111 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X354 VCO_C_0.INV_2_1.IN VCO_C_0.INV_2_3.IN.t54 VSS.t221 VSS.t220 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X355 VSS.t271 VSS.t269 VSS.t271 VSS.t270 nfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X356 VCO_C_0.INV_2_4.IN VCO_C_0.INV_2_2.IN.t55 VDD.t263 VDD.t262 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X357 VSS VCTRL2.t72 a_1424_1033.t24 VSS.t147 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X358 VDD DFF_3_mag_0.INV_2_0.OUT.t31 a_17597_2884.t5 VDD.t77 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X359 DFF_3_mag_0.INV_2_5.OUT DFF_3_mag_0.INV_2_5.IN.t30 VDD.t88 VDD.t87 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X360 VDD VCTRL.t17 VCO_C_0.INV_2_0.IN.t10 VDD.t325 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.84u
X361 VSS VCTRL2.t73 a_1424_1033.t23 VSS.t172 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X362 VDD VCO_C_0.INV_2_0.IN.t54 VCO_C_0.INV_2_5.IN.t28 VDD.t108 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X363 VDD DFF_3_mag_0.INV_2_1.IN.t26 DFF_3_mag_0.INV_2_5.IN.t5 VDD.t180 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X364 VDD VCO_C_0.INV_2_3.IN.t55 VCO_C_0.INV_2_1.IN.t0 VDD.t5 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X365 VCO_C_0.INV_2_5.IN VCO_C_0.INV_2_0.IN.t55 VDD.t339 VDD.t111 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X366 VSS VCTRL2.t74 a_10161_4198.t44 VSS.t142 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X367 VCO_C_0.INV_2_0.OUT VCO_C_0.INV_2_0.IN.t56 VSS.t130 VSS.t129 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X368 VSS VCTRL2.t75 a_1424_1033.t22 VSS.t185 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X369 VDD.t188 VDD.t186 VDD.t188 VDD.t187 pfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X370 VSS VCTRL2.t76 a_10161_4198.t38 VSS.t150 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X371 VDD VCO_C_0.OUTB.t51 DFF_3_mag_0.INV_2_0.OUT.t1 VDD.t317 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X372 VDD VCO_C_0.INV_2_0.IN.t57 VCO_C_0.INV_2_0.OUT.t11 VDD.t311 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X373 DFF_3_mag_0.INV_2_5.OUT DFF_3_mag_0.INV_2_5.IN.t31 VDD.t153 VDD.t87 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X374 VSS VCTRL2.t77 a_1424_1033.t21 VSS.t172 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X375 VDD VCO_C_0.INV_2_2.IN.t56 VCO_C_0.INV_2_4.IN.t1 VDD.t259 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X376 DFF_3_mag_0.INV_2_5.IN DFF_3_mag_0.INV_2_1.IN.t27 VSS.t374 VSS.t91 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X377 VSS OUT.t33 DFF_3_mag_0.INV_2_4.OUT.t13 VSS.t21 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X378 DFF_3_mag_0.INV_2_0.OUT VCO_C_0.OUTB.t52 VDD.t418 VDD.t320 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X379 VDD VCO_C_0.OUTB.t53 a_17597_1404.t0 VDD.t78 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X380 VCO_C_0.INV_2_2.IN VCTRL.t18 VDD.t335 VDD.t330 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.84u
X381 VCO_C_0.INV_2_5.IN VCTRL.t19 VDD.t336 VDD.t245 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X382 VSS VCTRL2.t78 a_10161_4198.t39 VSS.t150 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X383 VDD VCO_C_0.INV_2_2.IN.t57 VCO_C_0.INV_2_3.IN.t10 VDD.t29 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X384 VDD VCO_C_0.INV_2_3.IN.t56 VCO_C_0.INV_2_2.IN.t28 VDD.t2 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X385 VSS.t268 VSS.t266 VSS.t268 VSS.t267 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X386 VSS OUT.t34 DFF_3_mag_0.INV_2_4.OUT.t12 VSS.t24 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X387 VDD VCO_C_0.INV_2_2.IN.t58 VCO_C_0.INV_2_4.IN.t0 VDD.t254 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X388 DFF_3_mag_0.INV_2_4.OUT OUT.t35 VDD.t176 VDD.t150 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X389 VSS.t265 VSS.t263 VSS.t265 VSS.t264 nfet_03v3 ad=0 pd=0 as=0.22p ps=1.88u w=0.5u l=0.84u
X390 VSS VCTRL2.t79 a_1424_1033.t20 VSS.t185 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X391 VDD VCO_C_0.INV_2_5.IN.t57 VCO_C_0.INV_2_0.IN.t15 VDD.t103 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X392 VCO_C_0.INV_2_2.IN VCO_C_0.INV_2_0.OUT.t21 a_10161_4198.t45 VSS.t77 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X393 VDD VCO_C_0.INV_2_0.IN.t58 VCO_C_0.INV_2_5.IN.t30 VDD.t136 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X394 VDD VCO_C_0.INV_2_5.IN.t58 VCO_C_0.INV_2_5.OUT.t0 VDD.t139 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X395 VCO_C_0.INV_2_2.IN VCO_C_0.INV_2_3.IN.t57 VDD.t1 VDD.t0 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
R0 VCO_C_0.INV_2_0.OUT.n7 VCO_C_0.INV_2_0.OUT.t14 14.1829
R1 VCO_C_0.INV_2_0.OUT.n6 VCO_C_0.INV_2_0.OUT.t16 13.9657
R2 VCO_C_0.INV_2_0.OUT.n1 VCO_C_0.INV_2_0.OUT.t12 13.3574
R3 VCO_C_0.INV_2_0.OUT.n1 VCO_C_0.INV_2_0.OUT.t18 13.1401
R4 VCO_C_0.INV_2_0.OUT.n1 VCO_C_0.INV_2_0.OUT.t15 12.9025
R5 VCO_C_0.INV_2_0.OUT.n1 VCO_C_0.INV_2_0.OUT.t19 12.6187
R6 VCO_C_0.INV_2_0.OUT.n4 VCO_C_0.INV_2_0.OUT.t13 8.77788
R7 VCO_C_0.INV_2_0.OUT.n5 VCO_C_0.INV_2_0.OUT.t21 8.64752
R8 VCO_C_0.INV_2_0.OUT.n5 VCO_C_0.INV_2_0.OUT.t17 8.56062
R9 VCO_C_0.INV_2_0.OUT.n4 VCO_C_0.INV_2_0.OUT.t20 8.43026
R10 VCO_C_0.INV_2_0.OUT.n2 VCO_C_0.INV_2_0.OUT.n5 6.11825
R11 VCO_C_0.INV_2_0.OUT.n2 VCO_C_0.INV_2_0.OUT.n4 5.88354
R12 VCO_C_0.INV_2_0.OUT VCO_C_0.INV_2_0.OUT.n3 4.64372
R13 VCO_C_0.INV_2_0.OUT.n18 VCO_C_0.INV_2_0.OUT.t9 3.6405
R14 VCO_C_0.INV_2_0.OUT.n18 VCO_C_0.INV_2_0.OUT.n17 3.6405
R15 VCO_C_0.INV_2_0.OUT.n14 VCO_C_0.INV_2_0.OUT.t2 3.6405
R16 VCO_C_0.INV_2_0.OUT.n14 VCO_C_0.INV_2_0.OUT.n13 3.6405
R17 VCO_C_0.INV_2_0.OUT.n16 VCO_C_0.INV_2_0.OUT.t8 3.6405
R18 VCO_C_0.INV_2_0.OUT.n16 VCO_C_0.INV_2_0.OUT.n15 3.6405
R19 VCO_C_0.INV_2_0.OUT.n20 VCO_C_0.INV_2_0.OUT.t11 3.6405
R20 VCO_C_0.INV_2_0.OUT.n20 VCO_C_0.INV_2_0.OUT.n19 3.6405
R21 VCO_C_0.INV_2_0.OUT VCO_C_0.INV_2_0.OUT.n10 3.50463
R22 VCO_C_0.INV_2_0.OUT.n0 VCO_C_0.INV_2_0.OUT.n12 3.50463
R23 VCO_C_0.INV_2_0.OUT.n10 VCO_C_0.INV_2_0.OUT.t3 3.2765
R24 VCO_C_0.INV_2_0.OUT.n10 VCO_C_0.INV_2_0.OUT.n9 3.2765
R25 VCO_C_0.INV_2_0.OUT.n12 VCO_C_0.INV_2_0.OUT.t0 3.2765
R26 VCO_C_0.INV_2_0.OUT.n12 VCO_C_0.INV_2_0.OUT.n11 3.2765
R27 VCO_C_0.INV_2_0.OUT.n0 VCO_C_0.INV_2_0.OUT.n16 3.06224
R28 VCO_C_0.INV_2_0.OUT VCO_C_0.INV_2_0.OUT.n20 3.06224
R29 VCO_C_0.INV_2_0.OUT.n2 VCO_C_0.INV_2_0.OUT.n1 2.65077
R30 VCO_C_0.INV_2_0.OUT.n0 VCO_C_0.INV_2_0.OUT.n14 2.6005
R31 VCO_C_0.INV_2_0.OUT VCO_C_0.INV_2_0.OUT.n18 2.6005
R32 VCO_C_0.INV_2_0.OUT.n3 VCO_C_0.INV_2_0.OUT.n8 2.3804
R33 VCO_C_0.INV_2_0.OUT VCO_C_0.INV_2_0.OUT.n0 1.73202
R34 VCO_C_0.INV_2_0.OUT VCO_C_0.INV_2_0.OUT.n3 1.15983
R35 VCO_C_0.INV_2_0.OUT.n6 VCO_C_0.INV_2_0.OUT.n2 1.58291
R36 VCO_C_0.INV_2_0.OUT.n8 VCO_C_0.INV_2_0.OUT.n7 1.33917
R37 VCO_C_0.INV_2_0.OUT.n7 VCO_C_0.INV_2_0.OUT.n6 1.23958
R38 VCO_C_0.INV_2_2.IN.n71 VCO_C_0.INV_2_2.IN.n70 15.8172
R39 VCO_C_0.INV_2_2.IN.n72 VCO_C_0.INV_2_2.IN.n71 15.8172
R40 VCO_C_0.INV_2_2.IN.n73 VCO_C_0.INV_2_2.IN.n72 15.8172
R41 VCO_C_0.INV_2_2.IN.n71 VCO_C_0.INV_2_2.IN.t42 14.8925
R42 VCO_C_0.INV_2_2.IN.n72 VCO_C_0.INV_2_2.IN.t55 14.8925
R43 VCO_C_0.INV_2_2.IN.n69 VCO_C_0.INV_2_2.IN.n68 12.2457
R44 VCO_C_0.INV_2_2.IN.n68 VCO_C_0.INV_2_2.IN.n66 12.2457
R45 VCO_C_0.INV_2_2.IN.n66 VCO_C_0.INV_2_2.IN.n64 12.2457
R46 VCO_C_0.INV_2_2.IN.n74 VCO_C_0.INV_2_2.IN.t41 11.6285
R47 VCO_C_0.INV_2_2.IN.n19 VCO_C_0.INV_2_2.IN.t39 9.57577
R48 VCO_C_0.INV_2_2.IN.n22 VCO_C_0.INV_2_2.IN.t54 9.55796
R49 VCO_C_0.INV_2_2.IN.n64 VCO_C_0.INV_2_2.IN.t36 8.9065
R50 VCO_C_0.INV_2_2.IN.n66 VCO_C_0.INV_2_2.IN.t58 8.9065
R51 VCO_C_0.INV_2_2.IN.n68 VCO_C_0.INV_2_2.IN.t44 8.9065
R52 VCO_C_0.INV_2_2.IN.n69 VCO_C_0.INV_2_2.IN.t56 8.9065
R53 VCO_C_0.INV_2_2.IN.n70 VCO_C_0.INV_2_2.IN.t45 8.6145
R54 VCO_C_0.INV_2_2.IN.n71 VCO_C_0.INV_2_2.IN.t38 8.6145
R55 VCO_C_0.INV_2_2.IN.n72 VCO_C_0.INV_2_2.IN.t52 8.6145
R56 VCO_C_0.INV_2_2.IN.n73 VCO_C_0.INV_2_2.IN.t37 8.59715
R57 VCO_C_0.INV_2_2.IN.n61 VCO_C_0.INV_2_2.IN.n60 8.59228
R58 VCO_C_0.INV_2_2.IN.n19 VCO_C_0.INV_2_2.IN.t35 8.56851
R59 VCO_C_0.INV_2_2.IN.n20 VCO_C_0.INV_2_2.IN.t34 8.56851
R60 VCO_C_0.INV_2_2.IN.n21 VCO_C_0.INV_2_2.IN.t31 8.56851
R61 VCO_C_0.INV_2_2.IN.n5 VCO_C_0.INV_2_2.IN.t47 8.5214
R62 VCO_C_0.INV_2_2.IN.n1 VCO_C_0.INV_2_2.IN.t57 8.5214
R63 VCO_C_0.INV_2_2.IN.n2 VCO_C_0.INV_2_2.IN.t46 8.5214
R64 VCO_C_0.INV_2_2.IN.n7 VCO_C_0.INV_2_2.IN.t53 8.5214
R65 VCO_C_0.INV_2_2.IN.n24 VCO_C_0.INV_2_2.IN.t48 8.5112
R66 VCO_C_0.INV_2_2.IN.n23 VCO_C_0.INV_2_2.IN.t49 8.5112
R67 VCO_C_0.INV_2_2.IN.n22 VCO_C_0.INV_2_2.IN.t51 8.5112
R68 VCO_C_0.INV_2_2.IN.n1 VCO_C_0.INV_2_2.IN.t43 8.34992
R69 VCO_C_0.INV_2_2.IN.n64 VCO_C_0.INV_2_2.IN.t50 8.3225
R70 VCO_C_0.INV_2_2.IN.t41 VCO_C_0.INV_2_2.IN.n69 8.3225
R71 VCO_C_0.INV_2_2.IN.n55 VCO_C_0.INV_2_2.IN.n75 8.65114
R72 VCO_C_0.INV_2_2.IN.n7 VCO_C_0.INV_2_2.IN.t40 8.30779
R73 VCO_C_0.INV_2_2.IN.n2 VCO_C_0.INV_2_2.IN.t32 8.30779
R74 VCO_C_0.INV_2_2.IN.n5 VCO_C_0.INV_2_2.IN.t33 8.30779
R75 VCO_C_0.INV_2_2.IN.n54 VCO_C_0.INV_2_2.IN.n52 7.40037
R76 VCO_C_0.INV_2_2.IN.n4 VCO_C_0.INV_2_2.IN.t19 7.05758
R77 VCO_C_0.INV_2_2.IN.n3 VCO_C_0.INV_2_2.IN.n10 6.80072
R78 VCO_C_0.INV_2_2.IN.n61 VCO_C_0.INV_2_2.IN.n59 6.73941
R79 VCO_C_0.INV_2_2.IN VCO_C_0.INV_2_2.IN.t14 6.45366
R80 VCO_C_0.INV_2_2.IN.n17 VCO_C_0.INV_2_2.IN.t20 6.2092
R81 VCO_C_0.INV_2_2.IN.n14 VCO_C_0.INV_2_2.IN.n11 5.83551
R82 VCO_C_0.INV_2_2.IN.n46 VCO_C_0.INV_2_2.IN.t1 5.28839
R83 VCO_C_0.INV_2_2.IN.n36 VCO_C_0.INV_2_2.IN.t6 4.89657
R84 VCO_C_0.INV_2_2.IN.n32 VCO_C_0.INV_2_2.IN.n31 4.89653
R85 VCO_C_0.INV_2_2.IN.n54 VCO_C_0.INV_2_2.IN.n53 4.88218
R86 VCO_C_0.INV_2_2.IN.n63 VCO_C_0.INV_2_2.IN 4.87529
R87 VCO_C_0.INV_2_2.IN.n6 VCO_C_0.INV_2_2.IN.t13 4.6632
R88 VCO_C_0.INV_2_2.IN.n40 VCO_C_0.INV_2_2.IN.t4 4.63112
R89 VCO_C_0.INV_2_2.IN VCO_C_0.INV_2_2.IN.n74 4.223
R90 VCO_C_0.INV_2_2.IN.n33 VCO_C_0.INV_2_2.IN.n32 4.04562
R91 VCO_C_0.INV_2_2.IN.n47 VCO_C_0.INV_2_2.IN.n46 4.02915
R92 VCO_C_0.INV_2_2.IN.n49 VCO_C_0.INV_2_2.IN.n48 4.01867
R93 VCO_C_0.INV_2_2.IN.n62 VCO_C_0.INV_2_2.IN.n58 3.9838
R94 VCO_C_0.INV_2_2.IN.n0 VCO_C_0.INV_2_2.IN.n63 3.96161
R95 VCO_C_0.INV_2_2.IN.n49 VCO_C_0.INV_2_2.IN.n54 3.87403
R96 VCO_C_0.INV_2_2.IN.t58 VCO_C_0.INV_2_2.IN.n65 3.6505
R97 VCO_C_0.INV_2_2.IN.t44 VCO_C_0.INV_2_2.IN.n67 3.6505
R98 VCO_C_0.INV_2_2.IN.n58 VCO_C_0.INV_2_2.IN.t15 3.6405
R99 VCO_C_0.INV_2_2.IN.n58 VCO_C_0.INV_2_2.IN.n57 3.6405
R100 VCO_C_0.INV_2_2.IN.n38 VCO_C_0.INV_2_2.IN.t7 3.6405
R101 VCO_C_0.INV_2_2.IN.n38 VCO_C_0.INV_2_2.IN.n37 3.6405
R102 VCO_C_0.INV_2_2.IN.n29 VCO_C_0.INV_2_2.IN.t9 3.6405
R103 VCO_C_0.INV_2_2.IN.n29 VCO_C_0.INV_2_2.IN.n28 3.6405
R104 VCO_C_0.INV_2_2.IN.n43 VCO_C_0.INV_2_2.IN.t28 3.6405
R105 VCO_C_0.INV_2_2.IN.n43 VCO_C_0.INV_2_2.IN.n42 3.6405
R106 VCO_C_0.INV_2_2.IN.n51 VCO_C_0.INV_2_2.IN.t8 3.6405
R107 VCO_C_0.INV_2_2.IN.n51 VCO_C_0.INV_2_2.IN.n50 3.6405
R108 VCO_C_0.INV_2_2.IN.n13 VCO_C_0.INV_2_2.IN.t22 3.47629
R109 VCO_C_0.INV_2_2.IN.n16 VCO_C_0.INV_2_2.IN.t21 3.47629
R110 VCO_C_0.INV_2_2.IN.n9 VCO_C_0.INV_2_2.IN.t18 3.47617
R111 VCO_C_0.INV_2_2.IN.n14 VCO_C_0.INV_2_2.IN.n13 3.3987
R112 VCO_C_0.INV_2_2.IN.n74 VCO_C_0.INV_2_2.IN.n73 3.1807
R113 VCO_C_0.INV_2_2.IN.n35 VCO_C_0.INV_2_2.IN.n38 5.42442
R114 VCO_C_0.INV_2_2.IN.n45 VCO_C_0.INV_2_2.IN.n44 2.88562
R115 VCO_C_0.INV_2_2.IN.n9 VCO_C_0.INV_2_2.IN.n8 2.86157
R116 VCO_C_0.INV_2_2.IN.n16 VCO_C_0.INV_2_2.IN.n15 2.86147
R117 VCO_C_0.INV_2_2.IN.n13 VCO_C_0.INV_2_2.IN.n12 2.86147
R118 VCO_C_0.INV_2_2.IN.n4 VCO_C_0.INV_2_2.IN.n16 2.48336
R119 VCO_C_0.INV_2_2.IN.n3 VCO_C_0.INV_2_2.IN.n9 2.47781
R120 VCO_C_0.INV_2_2.IN.n0 VCO_C_0.INV_2_2.IN 2.35499
R121 VCO_C_0.INV_2_2.IN.n18 VCO_C_0.INV_2_2.IN 2.30073
R122 VCO_C_0.INV_2_2.IN.n6 VCO_C_0.INV_2_2.IN.n39 2.24532
R123 VCO_C_0.INV_2_2.IN.n39 VCO_C_0.INV_2_2.IN.n27 2.21522
R124 VCO_C_0.INV_2_2.IN.n35 VCO_C_0.INV_2_2.IN.n34 1.7262
R125 VCO_C_0.INV_2_2.IN.n27 VCO_C_0.INV_2_2.IN.n26 1.71923
R126 VCO_C_0.INV_2_2.IN.n44 VCO_C_0.INV_2_2.IN.n43 1.65851
R127 VCO_C_0.INV_2_2.IN.n25 VCO_C_0.INV_2_2.IN.n24 1.61187
R128 VCO_C_0.INV_2_2.IN.n25 VCO_C_0.INV_2_2.IN.n21 1.57365
R129 VCO_C_0.INV_2_2.IN VCO_C_0.INV_2_2.IN.n62 1.51605
R130 VCO_C_0.INV_2_2.IN.n41 VCO_C_0.INV_2_2.IN.n40 1.51564
R131 VCO_C_0.INV_2_2.IN VCO_C_0.INV_2_2.IN.n0 1.51518
R132 VCO_C_0.INV_2_2.IN.n26 VCO_C_0.INV_2_2.IN.n30 1.49487
R133 VCO_C_0.INV_2_2.IN.n34 VCO_C_0.INV_2_2.IN.n36 1.49463
R134 VCO_C_0.INV_2_2.IN.n48 VCO_C_0.INV_2_2.IN.n51 1.25753
R135 VCO_C_0.INV_2_2.IN.n30 VCO_C_0.INV_2_2.IN.n29 1.25657
R136 VCO_C_0.INV_2_2.IN.n3 VCO_C_0.INV_2_2.IN.n4 1.05601
R137 VCO_C_0.INV_2_2.IN.n18 VCO_C_0.INV_2_2.IN.n17 1.01067
R138 VCO_C_0.INV_2_2.IN.n23 VCO_C_0.INV_2_2.IN.n22 0.996664
R139 VCO_C_0.INV_2_2.IN.n1 VCO_C_0.INV_2_2.IN.n5 0.992966
R140 VCO_C_0.INV_2_2.IN.n4 VCO_C_0.INV_2_2.IN.n14 0.983286
R141 VCO_C_0.INV_2_2.IN.n2 VCO_C_0.INV_2_2.IN.n1 0.975705
R142 VCO_C_0.INV_2_2.IN.n56 VCO_C_0.INV_2_2.IN.n41 0.969569
R143 VCO_C_0.INV_2_2.IN.n63 VCO_C_0.INV_2_2.IN.n56 0.955885
R144 VCO_C_0.INV_2_2.IN.n20 VCO_C_0.INV_2_2.IN.n19 0.953514
R145 VCO_C_0.INV_2_2.IN.n17 VCO_C_0.INV_2_2.IN.n3 0.907492
R146 VCO_C_0.INV_2_2.IN.n47 VCO_C_0.INV_2_2.IN.n49 0.856289
R147 VCO_C_0.INV_2_2.IN.n45 VCO_C_0.INV_2_2.IN.n55 0.843096
R148 VCO_C_0.INV_2_2.IN.n27 VCO_C_0.INV_2_2.IN.n33 0.8015
R149 VCO_C_0.INV_2_2.IN.n62 VCO_C_0.INV_2_2.IN.n61 0.800717
R150 VCO_C_0.INV_2_2.IN.n40 VCO_C_0.INV_2_2.IN.n6 0.741058
R151 VCO_C_0.INV_2_2.IN.n41 VCO_C_0.INV_2_2.IN.n7 0.69855
R152 VCO_C_0.INV_2_2.IN.n56 VCO_C_0.INV_2_2.IN.n45 0.656716
R153 VCO_C_0.INV_2_2.IN.n0 VCO_C_0.INV_2_2.IN.n18 0.555846
R154 VCO_C_0.INV_2_2.IN.n55 VCO_C_0.INV_2_2.IN.n47 0.398395
R155 VCO_C_0.INV_2_2.IN.n33 VCO_C_0.INV_2_2.IN.n35 0.3875
R156 VCO_C_0.INV_2_2.IN.n21 VCO_C_0.INV_2_2.IN.n20 0.364199
R157 VCO_C_0.INV_2_2.IN.n7 VCO_C_0.INV_2_2.IN.n2 0.359267
R158 VCO_C_0.INV_2_2.IN.n24 VCO_C_0.INV_2_2.IN.n23 0.323514
R159 VCO_C_0.INV_2_2.IN.n5 VCO_C_0.INV_2_2.IN.n25 0.319815
R160 a_10161_4198.n66 a_10161_4198.n59 9.67588
R161 a_10161_4198.n24 a_10161_4198.n21 3.74722
R162 a_10161_4198.n0 a_10161_4198.n50 3.71799
R163 a_10161_4198.n3 a_10161_4198.n38 3.74413
R164 a_10161_4198.n2 a_10161_4198.n9 3.70973
R165 a_10161_4198.n77 a_10161_4198.t9 3.2765
R166 a_10161_4198.n77 a_10161_4198.n76 3.2765
R167 a_10161_4198.n79 a_10161_4198.t59 3.2765
R168 a_10161_4198.n79 a_10161_4198.n78 3.2765
R169 a_10161_4198.n85 a_10161_4198.t50 3.2765
R170 a_10161_4198.n85 a_10161_4198.n84 3.2765
R171 a_10161_4198.n68 a_10161_4198.t47 3.2765
R172 a_10161_4198.n68 a_10161_4198.n67 3.2765
R173 a_10161_4198.n61 a_10161_4198.t51 3.2765
R174 a_10161_4198.n61 a_10161_4198.n60 3.2765
R175 a_10161_4198.n63 a_10161_4198.t37 3.2765
R176 a_10161_4198.n63 a_10161_4198.n62 3.2765
R177 a_10161_4198.n81 a_10161_4198.t11 3.2765
R178 a_10161_4198.n81 a_10161_4198.n80 3.2765
R179 a_10161_4198.n70 a_10161_4198.t49 3.2765
R180 a_10161_4198.n70 a_10161_4198.n69 3.2765
R181 a_10161_4198.n72 a_10161_4198.t45 3.2765
R182 a_10161_4198.n72 a_10161_4198.n71 3.2765
R183 a_10161_4198.n17 a_10161_4198.t58 3.2765
R184 a_10161_4198.n17 a_10161_4198.n16 3.2765
R185 a_10161_4198.n27 a_10161_4198.t28 3.2765
R186 a_10161_4198.n27 a_10161_4198.n26 3.2765
R187 a_10161_4198.n19 a_10161_4198.t3 3.2765
R188 a_10161_4198.n19 a_10161_4198.n18 3.2765
R189 a_10161_4198.n52 a_10161_4198.t39 3.2765
R190 a_10161_4198.n52 a_10161_4198.n51 3.2765
R191 a_10161_4198.n48 a_10161_4198.t17 3.2765
R192 a_10161_4198.n48 a_10161_4198.n47 3.2765
R193 a_10161_4198.n55 a_10161_4198.t41 3.2765
R194 a_10161_4198.n55 a_10161_4198.n54 3.2765
R195 a_10161_4198.n46 a_10161_4198.t38 3.2765
R196 a_10161_4198.n46 a_10161_4198.n45 3.2765
R197 a_10161_4198.n32 a_10161_4198.t5 3.2765
R198 a_10161_4198.n32 a_10161_4198.n31 3.2765
R199 a_10161_4198.n34 a_10161_4198.t19 3.2765
R200 a_10161_4198.n34 a_10161_4198.n33 3.2765
R201 a_10161_4198.n14 a_10161_4198.t22 3.2765
R202 a_10161_4198.n14 a_10161_4198.n13 3.2765
R203 a_10161_4198.n5 a_10161_4198.t15 3.2765
R204 a_10161_4198.n5 a_10161_4198.n4 3.2765
R205 a_10161_4198.n7 a_10161_4198.t44 3.2765
R206 a_10161_4198.n7 a_10161_4198.n6 3.2765
R207 a_10161_4198.n11 a_10161_4198.t16 3.2765
R208 a_10161_4198.n11 a_10161_4198.n10 3.2765
R209 a_10161_4198.n9 a_10161_4198.t23 3.2765
R210 a_10161_4198.n9 a_10161_4198.n8 3.2765
R211 a_10161_4198.n36 a_10161_4198.t34 3.2765
R212 a_10161_4198.n36 a_10161_4198.n35 3.2765
R213 a_10161_4198.n41 a_10161_4198.t7 3.2765
R214 a_10161_4198.n41 a_10161_4198.n40 3.2765
R215 a_10161_4198.n38 a_10161_4198.t21 3.2765
R216 a_10161_4198.n38 a_10161_4198.n37 3.2765
R217 a_10161_4198.n50 a_10161_4198.t25 3.2765
R218 a_10161_4198.n50 a_10161_4198.n49 3.2765
R219 a_10161_4198.n23 a_10161_4198.t32 3.2765
R220 a_10161_4198.n23 a_10161_4198.n22 3.2765
R221 a_10161_4198.n21 a_10161_4198.t42 3.2765
R222 a_10161_4198.n21 a_10161_4198.n20 3.2765
R223 a_10161_4198.n93 a_10161_4198.t8 3.2765
R224 a_10161_4198.n94 a_10161_4198.n93 3.2765
R225 a_10161_4198.n15 a_10161_4198.n5 3.1505
R226 a_10161_4198.n12 a_10161_4198.n7 3.1505
R227 a_10161_4198.n42 a_10161_4198.n36 3.1505
R228 a_10161_4198.n44 a_10161_4198.n32 3.1505
R229 a_10161_4198.n57 a_10161_4198.n46 3.1505
R230 a_10161_4198.n53 a_10161_4198.n48 3.1505
R231 a_10161_4198.n25 a_10161_4198.n19 3.1505
R232 a_10161_4198.n29 a_10161_4198.n17 3.1505
R233 a_10161_4198.n73 a_10161_4198.n72 3.1505
R234 a_10161_4198.n74 a_10161_4198.n70 3.1505
R235 a_10161_4198.n82 a_10161_4198.n81 3.1505
R236 a_10161_4198.n64 a_10161_4198.n63 3.1505
R237 a_10161_4198.n65 a_10161_4198.n61 3.1505
R238 a_10161_4198.n91 a_10161_4198.n68 3.1505
R239 a_10161_4198.n86 a_10161_4198.n85 3.1505
R240 a_10161_4198.n88 a_10161_4198.n79 3.1505
R241 a_10161_4198.n89 a_10161_4198.n77 3.1505
R242 a_10161_4198.n93 a_10161_4198.n92 3.1505
R243 a_10161_4198.n3 a_10161_4198.n39 2.24571
R244 a_10161_4198.n24 a_10161_4198.n23 1.84747
R245 a_10161_4198.n3 a_10161_4198.n41 1.84743
R246 a_10161_4198.n2 a_10161_4198.n11 1.84737
R247 a_10161_4198.n1 a_10161_4198.n14 1.84737
R248 a_10161_4198.n43 a_10161_4198.n34 1.84737
R249 a_10161_4198.n28 a_10161_4198.n27 1.84737
R250 a_10161_4198.n56 a_10161_4198.n55 1.84732
R251 a_10161_4198.n0 a_10161_4198.n52 1.84618
R252 a_10161_4198.n90 a_10161_4198.n75 0.972891
R253 a_10161_4198.n87 a_10161_4198.n83 0.972891
R254 a_10161_4198.n58 a_10161_4198.n57 0.899822
R255 a_10161_4198.n30 a_10161_4198.n29 0.899822
R256 a_10161_4198.n74 a_10161_4198.n73 0.758798
R257 a_10161_4198.n89 a_10161_4198.n88 0.758798
R258 a_10161_4198.n92 a_10161_4198.n66 0.724996
R259 a_10161_4198.n65 a_10161_4198.n64 0.7205
R260 a_10161_4198.n92 a_10161_4198.n91 0.7205
R261 a_10161_4198.n53 a_10161_4198.n0 0.66786
R262 a_10161_4198.n66 a_10161_4198.n65 0.636952
R263 a_10161_4198.n12 a_10161_4198.n2 0.627536
R264 a_10161_4198.n57 a_10161_4198.n56 0.610652
R265 a_10161_4198.n44 a_10161_4198.n43 0.607482
R266 a_10161_4198.n15 a_10161_4198.n1 0.604163
R267 a_10161_4198.n29 a_10161_4198.n28 0.60198
R268 a_10161_4198.n28 a_10161_4198.n25 0.601834
R269 a_10161_4198.n25 a_10161_4198.n24 0.601076
R270 a_10161_4198.n1 a_10161_4198.n12 0.598753
R271 a_10161_4198.n43 a_10161_4198.n42 0.595434
R272 a_10161_4198.n42 a_10161_4198.n3 0.593116
R273 a_10161_4198.n56 a_10161_4198.n53 0.592154
R274 a_10161_4198.n83 a_10161_4198.n82 0.555819
R275 a_10161_4198.n87 a_10161_4198.n86 0.555819
R276 a_10161_4198.n91 a_10161_4198.n90 0.551989
R277 a_10161_4198.n59 a_10161_4198.n58 0.378745
R278 a_10161_4198.n75 a_10161_4198.n74 0.283904
R279 a_10161_4198.n90 a_10161_4198.n89 0.283904
R280 a_10161_4198.n88 a_10161_4198.n87 0.280074
R281 a_10161_4198.n59 a_10161_4198.n30 0.248582
R282 a_10161_4198.n30 a_10161_4198.n15 0.247022
R283 a_10161_4198.n58 a_10161_4198.n44 0.247022
R284 VSS.n2427 VSS.n2426 5.93814e+06
R285 VSS.n1220 VSS.n1218 6613.27
R286 VSS.n1191 VSS.t290 6602.99
R287 VSS.t343 VSS.t299 4969.11
R288 VSS.n1126 VSS.t355 4768.34
R289 VSS.n1509 VSS.n1508 3480.07
R290 VSS.n2426 VSS.n2425 3326.77
R291 VSS.n0 VSS.t217 2458.99
R292 VSS.n1120 VSS.t360 2371.62
R293 VSS.n1598 VSS.t343 2308.88
R294 VSS.t372 VSS.t366 1753.97
R295 VSS.n1955 VSS.n1954 1514.17
R296 VSS.n531 VSS.n530 953.981
R297 VSS.n95 VSS.n94 944.048
R298 VSS.n375 VSS.n374 929.726
R299 VSS.n1221 VSS.n1220 632.529
R300 VSS.n2026 VSS.n2025 594.688
R301 VSS.n2668 VSS.n2667 588.614
R302 VSS.n1220 VSS.n1219 506.783
R303 VSS.n2662 VSS.n2661 489.312
R304 VSS.n0 VSS.t372 421.296
R305 VSS.n2728 VSS.n2727 407.524
R306 VSS.n1315 VSS.n1314 218.591
R307 VSS.n109 VSS.t125 154.649
R308 VSS.n557 VSS.t34 137.732
R309 VSS.n2921 VSS.n2920 132.9
R310 VSS.n2027 VSS.n2026 129.446
R311 VSS.n1277 VSS.t52 127.856
R312 VSS.n1568 VSS.n1567 127.8
R313 VSS.n2705 VSS.n2704 116.502
R314 VSS.n129 VSS.n128 109.445
R315 VSS.n1383 VSS.n1382 107.07
R316 VSS.t220 VSS.t109 88.6679
R317 VSS.n1599 VSS.n1598 77.5641
R318 VSS.n2052 VSS.t63 75.4357
R319 VSS.n2706 VSS.n2705 71.3171
R320 VSS.n1304 VSS.t129 70.1147
R321 VSS.n339 VSS.t21 68.7194
R322 VSS.n385 VSS.t19 68.7194
R323 VSS.n475 VSS.t55 68.7194
R324 VSS.n525 VSS.t38 68.7194
R325 VSS.n3122 VSS.t134 67.9645
R326 VSS.n43 VSS.t59 64.2392
R327 VSS.n1287 VSS.t61 61.866
R328 VSS.n2934 VSS.t31 60.4094
R329 VSS.n1961 VSS.t375 57.9753
R330 VSS.n162 VSS.n161 57.5226
R331 VSS.n1510 VSS.n1509 55.7009
R332 VSS.n2034 VSS.t122 53.4338
R333 VSS.n2073 VSS.t119 53.4338
R334 VSS.n2174 VSS.t293 51.6521
R335 VSS.n2007 VSS.t111 51.1548
R336 VSS.n3043 VSS.n3042 50.289
R337 VSS.n2315 VSS.t283 49.6265
R338 VSS.n3070 VSS.t40 49.4366
R339 VSS.n2043 VSS.t71 47.1475
R340 VSS.n2082 VSS.t88 47.1475
R341 VSS.n1121 VSS.n1120 44.0982
R342 VSS.n2581 VSS.t104 41.5243
R343 VSS.n1865 VSS.t264 41.5243
R344 VSS.n2627 VSS.n2626 39.4988
R345 VSS.n2007 VSS.t136 37.5136
R346 VSS.n2606 VSS.t35 35.4477
R347 VSS.n1028 VSS.t10 34.0944
R348 VSS.n2640 VSS.n2639 32.4093
R349 VSS.n1215 VSS.n1214 31.7508
R350 VSS.n1099 VSS.t78 30.8689
R351 VSS.n1961 VSS.t114 30.6931
R352 VSS.n1620 VSS.t150 30.685
R353 VSS.n1608 VSS.t296 30.685
R354 VSS.n2513 VSS.t199 28.3582
R355 VSS.n1799 VSS.t185 26.3327
R356 VSS.n105 VSS.t43 26.1718
R357 VSS.n2955 VSS.n2954 26.0884
R358 VSS.n1662 VSS.t322 25.5709
R359 VSS.n2088 VSS.t66 25.1456
R360 VSS.n2940 VSS.t30 24.1641
R361 VSS.n1 VSS.n0 22.6552
R362 VSS.n698 VSS.t70 22.1615
R363 VSS.n3015 VSS.n3014 20.5962
R364 VSS.n96 VSS.n95 19.0342
R365 VSS.n1061 VSS.t3 18.7521
R366 VSS.n2554 VSS.t172 18.2305
R367 VSS.n2013 VSS.t220 17.0519
R368 VSS.n456 VSS.t27 16.9915
R369 VSS.n288 VSS.t79 16.0849
R370 VSS.n450 VSS.t362 16.0476
R371 VSS.n626 VSS.t363 16.0476
R372 VSS.n678 VSS.t28 16.0476
R373 VSS.n1653 VSS.t7 15.3427
R374 VSS.n2290 VSS.t147 15.1921
R375 VSS.n36 VSS.t81 15.1388
R376 VSS.n258 VSS.t96 14.1926
R377 VSS.n1040 VSS.t0 13.6381
R378 VSS.n1769 VSS.t267 13.1666
R379 VSS.n2589 VSS.t103 13.1666
R380 VSS.n2284 VSS.t140 13.1666
R381 VSS.n1257 VSS.n1256 12.9423
R382 VSS.n193 VSS.n192 11.5049
R383 VSS.n1202 VSS.t60 11.4659
R384 VSS.n1034 VSS.t142 10.2287
R385 VSS.n2547 VSS.t175 10.1283
R386 VSS.n1737 VSS.n1736 9.61182
R387 VSS.n1745 VSS.t310 9.55913
R388 VSS.n1089 VSS.t354 9.55885
R389 VSS.n980 VSS.t298 9.54136
R390 VSS.n1752 VSS.t357 9.54089
R391 VSS.n1751 VSS.t305 9.51568
R392 VSS.n998 VSS.t342 9.5154
R393 VSS.n1753 VSS.t333 9.5085
R394 VSS.n967 VSS.t289 9.50824
R395 VSS.n1088 VSS.t359 9.49457
R396 VSS.n782 VSS.t285 9.49428
R397 VSS.n781 VSS.t287 9.49428
R398 VSS.n780 VSS.t326 9.49428
R399 VSS.n812 VSS.t301 9.49428
R400 VSS.n1940 VSS.t328 9.49403
R401 VSS.n1941 VSS.t347 9.49403
R402 VSS.n2059 VSS.t312 9.49403
R403 VSS.n2098 VSS.t324 9.49403
R404 VSS.n1918 VSS.t292 9.49372
R405 VSS.n813 VSS.t349 9.45083
R406 VSS.n1756 VSS.t266 9.45057
R407 VSS.n996 VSS.t336 9.43205
R408 VSS.n1086 VSS.t295 9.43205
R409 VSS.n986 VSS.t317 9.43205
R410 VSS.n978 VSS.t352 9.43205
R411 VSS.n969 VSS.t315 9.43205
R412 VSS.n2223 VSS.t263 9.43205
R413 VSS.n1903 VSS.t319 9.43205
R414 VSS.n1887 VSS.t303 9.43205
R415 VSS.n1749 VSS.t338 9.43205
R416 VSS.n1880 VSS.t340 9.43205
R417 VSS.n770 VSS.t280 9.3886
R418 VSS.n732 VSS.t277 9.3886
R419 VSS.n2405 VSS.t269 9.3886
R420 VSS.n2398 VSS.t282 9.3886
R421 VSS.n724 VSS.t345 9.34514
R422 VSS.n886 VSS.t321 9.34514
R423 VSS.n865 VSS.t274 9.34514
R424 VSS.n2366 VSS.t331 9.34514
R425 VSS.n2332 VSS.t307 9.34514
R426 VSS.n2337 VSS.t272 9.34514
R427 VSS.n510 VSS.n508 9.13939
R428 VSS.n2006 VSS.n1990 9.13939
R429 VSS.n2008 VSS.n2006 9.13939
R430 VSS.n1969 VSS.n1952 9.13939
R431 VSS.n1971 VSS.n1969 9.13939
R432 VSS.n1288 VSS.n1286 9.13939
R433 VSS.n1286 VSS.n1284 9.13939
R434 VSS.n2042 VSS.n1946 9.13939
R435 VSS.n2044 VSS.n2042 9.13939
R436 VSS.n2081 VSS.n2064 9.13939
R437 VSS.n2083 VSS.n2081 9.13939
R438 VSS.n1296 VSS.n1295 9.13939
R439 VSS.n1298 VSS.n1296 9.13939
R440 VSS.n363 VSS.n361 9.13939
R441 VSS.n643 VSS.n641 8.16717
R442 VSS.n371 VSS.n369 7.58383
R443 VSS.n501 VSS.n499 7.48661
R444 VSS.n2156 VSS.t65 7.08994
R445 VSS.n1626 VSS.t15 6.81928
R446 VSS.n1982 VSS.t221 6.65541
R447 VSS.n1957 VSS.n1953 6.65541
R448 VSS.n1994 VSS.n1991 6.65541
R449 VSS.n2019 VSS.t110 6.65541
R450 VSS.n2069 VSS.n2065 6.65541
R451 VSS.n2094 VSS.t64 6.65541
R452 VSS.n2055 VSS.t67 6.65541
R453 VSS.n2030 VSS.n1947 6.65541
R454 VSS.n1271 VSS.n778 6.65541
R455 VSS.n1271 VSS.n779 6.65541
R456 VSS.n1312 VSS.t135 6.65541
R457 VSS.n1312 VSS.t130 6.65541
R458 VSS.n332 VSS.n325 6.65541
R459 VSS.n332 VSS.n326 6.65541
R460 VSS.n378 VSS.t20 6.65541
R461 VSS.n378 VSS.t98 6.65541
R462 VSS.n686 VSS.t29 6.65541
R463 VSS.n622 VSS.n616 6.65541
R464 VSS.n468 VSS.n461 6.65541
R465 VSS.n468 VSS.n462 6.65541
R466 VSS.n534 VSS.t39 6.65541
R467 VSS.n534 VSS.t58 6.65541
R468 VSS.n310 VSS.t80 6.65541
R469 VSS.n241 VSS.n40 6.65541
R470 VSS.n1087 VSS.t297 6.63905
R471 VSS.n2225 VSS.t265 6.6371
R472 VSS.n771 VSS.t281 6.63522
R473 VSS.n733 VSS.t279 6.63522
R474 VSS.n2399 VSS.t284 6.63522
R475 VSS.n2406 VSS.t271 6.63522
R476 VSS.n725 VSS.t346 6.63331
R477 VSS.n2333 VSS.t309 6.63331
R478 VSS.n885 VSS.t323 6.5165
R479 VSS.n2367 VSS.t332 6.5165
R480 VSS.n866 VSS.t276 6.50525
R481 VSS.n2338 VSS.t273 6.50525
R482 VSS.n821 VSS.t201 6.4265
R483 VSS.n819 VSS.t260 6.4265
R484 VSS.n814 VSS.t198 6.4265
R485 VSS.n988 VSS.t337 6.4265
R486 VSS.n981 VSS.t318 6.4265
R487 VSS.n968 VSS.t353 6.4265
R488 VSS.n970 VSS.t316 6.4265
R489 VSS.n729 VSS.n728 6.4265
R490 VSS.n860 VSS.n859 6.4265
R491 VSS.n862 VSS.n861 6.4265
R492 VSS.n2303 VSS.t242 6.4265
R493 VSS.n2334 VSS.t200 6.4265
R494 VSS.n2329 VSS.t233 6.4265
R495 VSS.n2227 VSS.n2226 6.4265
R496 VSS.n2220 VSS.t339 6.4265
R497 VSS.n1897 VSS.t304 6.4265
R498 VSS.n2201 VSS.n2200 6.4265
R499 VSS.n1746 VSS.t320 6.4265
R500 VSS.n2204 VSS.n2203 6.4265
R501 VSS.n1881 VSS.t341 6.4265
R502 VSS.n1105 VSS.t77 6.17418
R503 VSS.n77 VSS.n76 5.80511
R504 VSS.n555 VSS.n554 5.26318
R505 VSS.n1266 VSS.n1265 5.2005
R506 VSS.n369 VSS.n368 5.2005
R507 VSS.n691 VSS.n690 5.2005
R508 VSS.n693 VSS.n692 5.2005
R509 VSS.n695 VSS.n694 5.2005
R510 VSS.n706 VSS.n705 5.2005
R511 VSS.n705 VSS.n704 5.2005
R512 VSS.n703 VSS.n702 5.2005
R513 VSS.n702 VSS.n701 5.2005
R514 VSS.n679 VSS.n678 5.2005
R515 VSS.n643 VSS.n642 5.2005
R516 VSS.n665 VSS.n664 5.2005
R517 VSS.n576 VSS.n575 5.2005
R518 VSS.n575 VSS.n574 5.2005
R519 VSS.n579 VSS.n578 5.2005
R520 VSS.n578 VSS.n577 5.2005
R521 VSS.n583 VSS.n581 5.2005
R522 VSS.n583 VSS.n582 5.2005
R523 VSS.n568 VSS.n567 5.2005
R524 VSS.n558 VSS.n557 5.2005
R525 VSS.n501 VSS.n491 5.2005
R526 VSS.n501 VSS.n500 5.2005
R527 VSS.n59 VSS.n58 5.2005
R528 VSS.n48 VSS.n47 5.2005
R529 VSS.n47 VSS.n46 5.2005
R530 VSS.n51 VSS.n50 5.2005
R531 VSS.n50 VSS.n49 5.2005
R532 VSS.n71 VSS.n70 5.2005
R533 VSS.n275 VSS.n274 5.2005
R534 VSS.n251 VSS.n250 5.2005
R535 VSS.n263 VSS.n262 5.2005
R536 VSS.n262 VSS.n261 5.2005
R537 VSS.n426 VSS.n425 5.2005
R538 VSS.n293 VSS.n292 5.2005
R539 VSS.n292 VSS.n291 5.2005
R540 VSS.n2 VSS.n1 5.2005
R541 VSS.n4 VSS.n3 5.2005
R542 VSS.n618 VSS.n617 5.2005
R543 VSS.n296 VSS.n295 5.2005
R544 VSS.n295 VSS.n294 5.2005
R545 VSS.n711 VSS.n710 5.12343
R546 VSS.n817 VSS.t4 5.1234
R547 VSS.n1081 VSS.t259 5.12337
R548 VSS.n2229 VSS.n2199 5.12337
R549 VSS.n2301 VSS.t206 5.12332
R550 VSS.n2207 VSS.n2206 5.12328
R551 VSS.n2310 VSS.t234 5.12118
R552 VSS.n752 VSS.n751 5.12105
R553 VSS.n45 VSS.n42 4.88449
R554 VSS.n573 VSS.n570 4.88277
R555 VSS.n700 VSS.n697 4.88215
R556 VSS.n664 VSS.t131 4.72022
R557 VSS.n1264 VSS.n1263 4.5005
R558 VSS.n323 VSS.n322 4.5005
R559 VSS.n700 VSS.n699 4.5005
R560 VSS.n699 VSS.n698 4.5005
R561 VSS.n676 VSS.n675 4.5005
R562 VSS.n663 VSS.n662 4.5005
R563 VSS.n635 VSS.n634 4.5005
R564 VSS.n586 VSS.n585 4.5005
R565 VSS.n585 VSS.n584 4.5005
R566 VSS.n563 VSS.n562 4.5005
R567 VSS.n562 VSS.n561 4.5005
R568 VSS.n573 VSS.n572 4.5005
R569 VSS.n572 VSS.n571 4.5005
R570 VSS.n504 VSS.n497 4.5005
R571 VSS.n504 VSS.n503 4.5005
R572 VSS.n80 VSS.n79 4.5005
R573 VSS.n79 VSS.n78 4.5005
R574 VSS.n45 VSS.n44 4.5005
R575 VSS.n44 VSS.n43 4.5005
R576 VSS.n68 VSS.n67 4.5005
R577 VSS.n67 VSS.n66 4.5005
R578 VSS.n278 VSS.n277 4.5005
R579 VSS.n254 VSS.n253 4.5005
R580 VSS.n269 VSS.n268 4.5005
R581 VSS.n268 VSS.n267 4.5005
R582 VSS.n429 VSS.n428 4.5005
R583 VSS.n299 VSS.n298 4.5005
R584 VSS.n298 VSS.n297 4.5005
R585 VSS.n1297 VSS.t49 4.12487
R586 VSS.n2616 VSS.n2615 4.05161
R587 VSS.n2612 VSS.n2610 4.05161
R588 VSS.n2612 VSS.n2611 4.05161
R589 VSS.n2607 VSS.n2605 4.05161
R590 VSS.n2607 VSS.n2606 4.05161
R591 VSS.n2602 VSS.n2601 4.05161
R592 VSS.n2598 VSS.n2597 4.05161
R593 VSS.n2594 VSS.n2593 4.05161
R594 VSS.n2590 VSS.n2589 4.05161
R595 VSS.n2586 VSS.n2585 4.05161
R596 VSS.n2582 VSS.n2581 4.05161
R597 VSS.n360 VSS.t68 4.04279
R598 VSS.n398 VSS.t24 4.04279
R599 VSS.n487 VSS.t91 4.04279
R600 VSS.n512 VSS.t93 4.04279
R601 VSS.n302 VSS.n301 3.95365
R602 VSS.n3017 VSS.n3013 3.59971
R603 VSS.n3045 VSS.n3044 3.59911
R604 VSS.n1951 VSS.t36 3.41078
R605 VSS.n1989 VSS.t107 3.41078
R606 VSS.n3073 VSS.t46 3.40989
R607 VSS.n1950 VSS.n1949 3.37941
R608 VSS.n1988 VSS.n1987 3.37941
R609 VSS.n2062 VSS.n2061 3.37941
R610 VSS.n1944 VSS.n1943 3.37941
R611 VSS.n1293 VSS.n1290 3.37941
R612 VSS.n1293 VSS.n1292 3.37941
R613 VSS.n321 VSS.n318 3.37941
R614 VSS.n321 VSS.n320 3.37941
R615 VSS.n639 VSS.n638 3.37941
R616 VSS.n506 VSS.n493 3.37941
R617 VSS.n506 VSS.n495 3.37941
R618 VSS.n264 VSS.n11 3.37941
R619 VSS.n1088 VSS.t361 3.333
R620 VSS.n1918 VSS.t294 3.33271
R621 VSS.n980 VSS.t300 3.33057
R622 VSS.n1752 VSS.t358 3.33036
R623 VSS.n1940 VSS.t330 3.32608
R624 VSS.n1941 VSS.t348 3.32608
R625 VSS.n2059 VSS.t314 3.32608
R626 VSS.n2098 VSS.t325 3.32608
R627 VSS.n782 VSS.t286 3.32582
R628 VSS.n781 VSS.t288 3.32582
R629 VSS.n780 VSS.t327 3.32582
R630 VSS.n812 VSS.t302 3.32582
R631 VSS.n1756 VSS.t268 3.32512
R632 VSS.n813 VSS.t351 3.32486
R633 VSS.n1089 VSS.t356 3.31238
R634 VSS.n1745 VSS.t311 3.31209
R635 VSS.n967 VSS.t291 3.31186
R636 VSS.n1753 VSS.t335 3.3116
R637 VSS.n998 VSS.t344 3.31143
R638 VSS.n1751 VSS.t306 3.31114
R639 VSS.n932 VSS.t215 3.2765
R640 VSS.n932 VSS.n931 3.2765
R641 VSS.n935 VSS.t230 3.2765
R642 VSS.n935 VSS.n934 3.2765
R643 VSS.n938 VSS.t139 3.2765
R644 VSS.n938 VSS.n937 3.2765
R645 VSS.n837 VSS.t2 3.2765
R646 VSS.n837 VSS.n836 3.2765
R647 VSS.n840 VSS.t162 3.2765
R648 VSS.n840 VSS.n839 3.2765
R649 VSS.n834 VSS.t258 3.2765
R650 VSS.n834 VSS.n833 3.2765
R651 VSS.n830 VSS.t188 3.2765
R652 VSS.n830 VSS.n829 3.2765
R653 VSS.n826 VSS.t1 3.2765
R654 VSS.n826 VSS.n825 3.2765
R655 VSS.n928 VSS.t168 3.2765
R656 VSS.n928 VSS.n927 3.2765
R657 VSS.n925 VSS.t16 3.2765
R658 VSS.n925 VSS.n924 3.2765
R659 VSS.n843 VSS.t205 3.2765
R660 VSS.n843 VSS.n842 3.2765
R661 VSS.n847 VSS.t204 3.2765
R662 VSS.n847 VSS.n846 3.2765
R663 VSS.n851 VSS.t11 3.2765
R664 VSS.n851 VSS.n850 3.2765
R665 VSS.n854 VSS.t209 3.2765
R666 VSS.n854 VSS.n853 3.2765
R667 VSS.n857 VSS.t246 3.2765
R668 VSS.n857 VSS.n856 3.2765
R669 VSS.n1839 VSS.t243 3.2765
R670 VSS.n1839 VSS.n1838 3.2765
R671 VSS.n1841 VSS.t238 3.2765
R672 VSS.n1841 VSS.n1840 3.2765
R673 VSS.n2233 VSS.t176 3.2765
R674 VSS.n2233 VSS.n2232 3.2765
R675 VSS.n2237 VSS.t247 3.2765
R676 VSS.n2237 VSS.n2236 3.2765
R677 VSS.n2231 VSS.t239 3.2765
R678 VSS.n2231 VSS.n2230 3.2765
R679 VSS.n2254 VSS.t216 3.2765
R680 VSS.n2254 VSS.n2253 3.2765
R681 VSS.n1830 VSS.t165 3.2765
R682 VSS.n1830 VSS.n1829 3.2765
R683 VSS.n1828 VSS.t6 3.2765
R684 VSS.n1828 VSS.n1827 3.2765
R685 VSS.n1824 VSS.t189 3.2765
R686 VSS.n1824 VSS.n1823 3.2765
R687 VSS.n1826 VSS.t212 3.2765
R688 VSS.n1826 VSS.n1825 3.2765
R689 VSS.n2248 VSS.t184 3.2765
R690 VSS.n2248 VSS.n2247 3.2765
R691 VSS.n2346 VSS.t141 3.2765
R692 VSS.n2346 VSS.n2345 3.2765
R693 VSS.n2344 VSS.t237 3.2765
R694 VSS.n2344 VSS.n2343 3.2765
R695 VSS.n2342 VSS.t181 3.2765
R696 VSS.n2342 VSS.n2341 3.2765
R697 VSS.n2340 VSS.t169 3.2765
R698 VSS.n2340 VSS.n2339 3.2765
R699 VSS.n1949 VSS.t37 3.2765
R700 VSS.n1949 VSS.n1948 3.2765
R701 VSS.n1987 VSS.t108 3.2765
R702 VSS.n1987 VSS.n1986 3.2765
R703 VSS.n2061 VSS.t118 3.2765
R704 VSS.n2061 VSS.n2060 3.2765
R705 VSS.n1943 VSS.t257 3.2765
R706 VSS.n1943 VSS.n1942 3.2765
R707 VSS.n1292 VSS.t62 3.2765
R708 VSS.n1292 VSS.n1291 3.2765
R709 VSS.n1290 VSS.t74 3.2765
R710 VSS.n1290 VSS.n1289 3.2765
R711 VSS.n320 VSS.t87 3.2765
R712 VSS.n320 VSS.n319 3.2765
R713 VSS.n318 VSS.t69 3.2765
R714 VSS.n318 VSS.n317 3.2765
R715 VSS.n638 VSS.t371 3.2765
R716 VSS.n638 VSS.n637 3.2765
R717 VSS.n495 VSS.t92 3.2765
R718 VSS.n495 VSS.n494 3.2765
R719 VSS.n493 VSS.t374 3.2765
R720 VSS.n493 VSS.n492 3.2765
R721 VSS.n11 VSS.t97 3.2765
R722 VSS.n11 VSS.n10 3.2765
R723 VSS.n929 VSS.n928 3.1505
R724 VSS.n858 VSS.n857 3.1505
R725 VSS.n855 VSS.n854 3.1505
R726 VSS.n848 VSS.n847 3.1505
R727 VSS.n831 VSS.n830 3.1505
R728 VSS.n841 VSS.n840 3.1505
R729 VSS.n838 VSS.n837 3.1505
R730 VSS.n939 VSS.n938 3.1505
R731 VSS.n936 VSS.n935 3.1505
R732 VSS.n1834 VSS.n1826 3.1505
R733 VSS.n1835 VSS.n1824 3.1505
R734 VSS.n1831 VSS.n1830 3.1505
R735 VSS.n2351 VSS.n2340 3.1505
R736 VSS.n2350 VSS.n2342 3.1505
R737 VSS.n2347 VSS.n2346 3.1505
R738 VSS.n2238 VSS.n2237 3.1505
R739 VSS.n1842 VSS.n1841 3.1505
R740 VSS.n1843 VSS.n1839 3.1505
R741 VSS.n1945 VSS.t256 3.14363
R742 VSS.n2063 VSS.t117 3.14363
R743 VSS.n1261 VSS.n1260 3.07743
R744 VSS.n2620 VSS.n2619 3.03883
R745 VSS.n1165 VSS.n1164 2.83943
R746 VSS.n1169 VSS.n1168 2.83943
R747 VSS.n2118 VSS.n2117 2.83943
R748 VSS.n2122 VSS.n2121 2.83943
R749 VSS.n2125 VSS.n2124 2.83943
R750 VSS.n2128 VSS.n2127 2.83943
R751 VSS.n2132 VSS.n2131 2.83943
R752 VSS.n1957 VSS.n1956 2.64393
R753 VSS.n1994 VSS.n1993 2.64393
R754 VSS.n926 VSS.n925 2.6255
R755 VSS.n852 VSS.n851 2.6255
R756 VSS.n835 VSS.n834 2.6255
R757 VSS.n933 VSS.n932 2.6255
R758 VSS.n1833 VSS.n1828 2.6255
R759 VSS.n2349 VSS.n2344 2.6255
R760 VSS.n2239 VSS.n2231 2.6255
R761 VSS.n2234 VSS.n2233 2.6255
R762 VSS.n2266 VSS.n1744 2.61042
R763 VSS.n2293 VSS.n2280 2.61042
R764 VSS.n2325 VSS.n2298 2.61042
R765 VSS.n2490 VSS.n2489 2.60873
R766 VSS.n1689 VSS.n777 2.60818
R767 VSS.n434 VSS.n9 2.60616
R768 VSS.n20 VSS.n14 2.60562
R769 VSS.n331 VSS.n328 2.60491
R770 VSS.n377 VSS.n376 2.60491
R771 VSS.n467 VSS.n464 2.60491
R772 VSS.n533 VSS.n532 2.60491
R773 VSS.n2376 VSS.n2375 2.60246
R774 VSS.n2402 VSS.n2401 2.60244
R775 VSS.n2409 VSS.n2408 2.60244
R776 VSS.n880 VSS.n873 2.60148
R777 VSS.n736 VSS.n727 2.60147
R778 VSS.n1361 VSS.n1360 2.6005
R779 VSS.n1371 VSS.n1370 2.6005
R780 VSS.n1369 VSS.n1368 2.6005
R781 VSS.n1366 VSS.n1365 2.6005
R782 VSS.n1364 VSS.n1363 2.6005
R783 VSS.n1375 VSS.n1374 2.6005
R784 VSS.n1359 VSS.n1358 2.6005
R785 VSS.n1358 VSS.n1357 2.6005
R786 VSS.n1356 VSS.n1355 2.6005
R787 VSS.n1355 VSS.n1354 2.6005
R788 VSS.n1353 VSS.n1352 2.6005
R789 VSS.n1352 VSS.n1351 2.6005
R790 VSS.n1350 VSS.n1349 2.6005
R791 VSS.n1349 VSS.n1348 2.6005
R792 VSS.n1347 VSS.n1346 2.6005
R793 VSS.n1346 VSS.n1345 2.6005
R794 VSS.n1344 VSS.n1343 2.6005
R795 VSS.n1343 VSS.n1342 2.6005
R796 VSS.n1341 VSS.n1340 2.6005
R797 VSS.n1340 VSS.n1339 2.6005
R798 VSS.n1338 VSS.n1337 2.6005
R799 VSS.n1337 VSS.n1336 2.6005
R800 VSS.n1335 VSS.n1334 2.6005
R801 VSS.n1334 VSS.n1333 2.6005
R802 VSS.n1332 VSS.n1331 2.6005
R803 VSS.n1331 VSS.n1330 2.6005
R804 VSS.n1329 VSS.n1328 2.6005
R805 VSS.n1328 VSS.n1327 2.6005
R806 VSS.n1326 VSS.n1325 2.6005
R807 VSS.n1325 VSS.n1324 2.6005
R808 VSS.n1323 VSS.n1322 2.6005
R809 VSS.n1322 VSS.n1321 2.6005
R810 VSS.n1320 VSS.n1319 2.6005
R811 VSS.n1319 VSS.n1318 2.6005
R812 VSS.n2424 VSS.n2423 2.6005
R813 VSS.n2423 VSS.n2422 2.6005
R814 VSS.n2429 VSS.n2428 2.6005
R815 VSS.n2428 VSS.n2427 2.6005
R816 VSS.n2431 VSS.n2430 2.6005
R817 VSS.n2417 VSS.n2416 2.6005
R818 VSS.n2185 VSS.n2184 2.6005
R819 VSS.n2184 VSS.n2183 2.6005
R820 VSS.n2317 VSS.n2316 2.6005
R821 VSS.n2316 VSS.n2315 2.6005
R822 VSS.n2314 VSS.n2313 2.6005
R823 VSS.n2313 VSS.n2312 2.6005
R824 VSS.n2328 VSS.n2327 2.6005
R825 VSS.n2327 VSS.n2326 2.6005
R826 VSS.n2420 VSS.n2419 2.6005
R827 VSS.n1798 VSS.n1797 2.6005
R828 VSS.n2144 VSS.n2143 2.6005
R829 VSS.n2133 VSS.n2132 2.6005
R830 VSS.n2129 VSS.n2128 2.6005
R831 VSS.n2126 VSS.n2125 2.6005
R832 VSS.n2123 VSS.n2122 2.6005
R833 VSS.n2119 VSS.n2118 2.6005
R834 VSS.n2116 VSS.n2115 2.6005
R835 VSS.n2113 VSS.n2112 2.6005
R836 VSS.n2110 VSS.n2109 2.6005
R837 VSS.n2107 VSS.n2106 2.6005
R838 VSS.n2104 VSS.n2103 2.6005
R839 VSS.n2102 VSS.n2101 2.6005
R840 VSS.n2100 VSS.n2099 2.6005
R841 VSS.n1759 VSS.n1758 2.6005
R842 VSS.n1762 VSS.n1761 2.6005
R843 VSS.n2146 VSS.n2145 2.6005
R844 VSS.n1763 VSS.n1755 2.6005
R845 VSS.n1755 VSS.n1754 2.6005
R846 VSS.n1766 VSS.n1765 2.6005
R847 VSS.n1765 VSS.n1764 2.6005
R848 VSS.n1768 VSS.n1767 2.6005
R849 VSS.n1771 VSS.n1770 2.6005
R850 VSS.n1770 VSS.n1769 2.6005
R851 VSS.n1774 VSS.n1773 2.6005
R852 VSS.n1773 VSS.n1772 2.6005
R853 VSS.n1776 VSS.n1775 2.6005
R854 VSS.n1778 VSS.n1777 2.6005
R855 VSS.n1780 VSS.n1779 2.6005
R856 VSS.n1782 VSS.n1781 2.6005
R857 VSS.n1784 VSS.n1783 2.6005
R858 VSS.n1786 VSS.n1785 2.6005
R859 VSS.n1788 VSS.n1787 2.6005
R860 VSS.n1790 VSS.n1789 2.6005
R861 VSS.n1793 VSS.n1792 2.6005
R862 VSS.n1792 VSS.n1791 2.6005
R863 VSS.n1796 VSS.n1795 2.6005
R864 VSS.n1795 VSS.n1794 2.6005
R865 VSS.n2393 VSS.n2392 2.6005
R866 VSS.n2395 VSS.n2394 2.6005
R867 VSS.n2404 VSS.n2403 2.6005
R868 VSS.n2454 VSS.n2453 2.6005
R869 VSS.n2451 VSS.n2450 2.6005
R870 VSS.n2448 VSS.n2447 2.6005
R871 VSS.n2445 VSS.n2444 2.6005
R872 VSS.n2434 VSS.n2433 2.6005
R873 VSS.n2436 VSS.n2435 2.6005
R874 VSS.n2439 VSS.n2438 2.6005
R875 VSS.n2442 VSS.n2441 2.6005
R876 VSS.n2378 VSS.n2377 2.6005
R877 VSS.n2460 VSS.n2459 2.6005
R878 VSS.n2411 VSS.n2410 2.6005
R879 VSS.n2470 VSS.n2469 2.6005
R880 VSS.n2467 VSS.n2466 2.6005
R881 VSS.n2465 VSS.n2464 2.6005
R882 VSS.n2462 VSS.n2461 2.6005
R883 VSS.n2472 VSS.n2471 2.6005
R884 VSS.n2476 VSS.n2475 2.6005
R885 VSS.n2478 VSS.n2477 2.6005
R886 VSS.n2481 VSS.n2480 2.6005
R887 VSS.n2483 VSS.n2482 2.6005
R888 VSS.n2487 VSS.n2486 2.6005
R889 VSS.n2456 VSS.n2455 2.6005
R890 VSS.n2384 VSS.n2383 2.6005
R891 VSS.n2382 VSS.n2381 2.6005
R892 VSS.n2387 VSS.n2386 2.6005
R893 VSS.n2389 VSS.n2388 2.6005
R894 VSS.n1928 VSS.n1927 2.6005
R895 VSS.n1926 VSS.n1925 2.6005
R896 VSS.n1920 VSS.n1919 2.6005
R897 VSS.n1917 VSS.n1916 2.6005
R898 VSS.n1914 VSS.n1913 2.6005
R899 VSS.n1911 VSS.n1910 2.6005
R900 VSS.n1907 VSS.n1906 2.6005
R901 VSS.n1896 VSS.n1895 2.6005
R902 VSS.n1893 VSS.n1892 2.6005
R903 VSS.n1891 VSS.n1890 2.6005
R904 VSS.n1879 VSS.n1878 2.6005
R905 VSS.n1876 VSS.n1875 2.6005
R906 VSS.n1935 VSS.n1934 2.6005
R907 VSS.n1874 VSS.n1873 2.6005
R908 VSS.n1870 VSS.n1869 2.6005
R909 VSS.n1869 VSS.n1868 2.6005
R910 VSS.n1867 VSS.n1866 2.6005
R911 VSS.n1866 VSS.n1865 2.6005
R912 VSS.n1864 VSS.n1863 2.6005
R913 VSS.n1863 VSS.n1862 2.6005
R914 VSS.n1861 VSS.n1860 2.6005
R915 VSS.n1860 VSS.n1859 2.6005
R916 VSS.n1858 VSS.n1857 2.6005
R917 VSS.n1857 VSS.n1856 2.6005
R918 VSS.n1854 VSS.n1853 2.6005
R919 VSS.n1853 VSS.n1852 2.6005
R920 VSS.n1851 VSS.n1850 2.6005
R921 VSS.n1850 VSS.n1849 2.6005
R922 VSS.n1847 VSS.n1846 2.6005
R923 VSS.n1846 VSS.n1845 2.6005
R924 VSS.n1801 VSS.n1800 2.6005
R925 VSS.n1800 VSS.n1799 2.6005
R926 VSS.n1822 VSS.n1821 2.6005
R927 VSS.n1821 VSS.n1820 2.6005
R928 VSS.n1818 VSS.n1817 2.6005
R929 VSS.n1817 VSS.n1816 2.6005
R930 VSS.n1815 VSS.n1814 2.6005
R931 VSS.n1814 VSS.n1813 2.6005
R932 VSS.n1812 VSS.n1811 2.6005
R933 VSS.n1811 VSS.n1810 2.6005
R934 VSS.n1808 VSS.n1807 2.6005
R935 VSS.n1807 VSS.n1806 2.6005
R936 VSS.n1804 VSS.n1803 2.6005
R937 VSS.n1803 VSS.n1802 2.6005
R938 VSS.n2355 VSS.n2354 2.6005
R939 VSS.n2354 VSS.n2353 2.6005
R940 VSS.n2358 VSS.n2357 2.6005
R941 VSS.n2357 VSS.n2356 2.6005
R942 VSS.n2362 VSS.n2361 2.6005
R943 VSS.n2361 VSS.n2360 2.6005
R944 VSS.n2370 VSS.n2369 2.6005
R945 VSS.n2369 VSS.n2368 2.6005
R946 VSS.n2373 VSS.n2372 2.6005
R947 VSS.n2372 VSS.n2371 2.6005
R948 VSS.n2320 VSS.n2319 2.6005
R949 VSS.n2319 VSS.n2318 2.6005
R950 VSS.n2324 VSS.n2323 2.6005
R951 VSS.n2323 VSS.n2322 2.6005
R952 VSS.n2298 VSS.n2297 2.6005
R953 VSS.n2296 VSS.n2295 2.6005
R954 VSS.n2295 VSS.n2294 2.6005
R955 VSS.n2283 VSS.n2282 2.6005
R956 VSS.n2282 VSS.n2281 2.6005
R957 VSS.n2286 VSS.n2285 2.6005
R958 VSS.n2285 VSS.n2284 2.6005
R959 VSS.n2289 VSS.n2288 2.6005
R960 VSS.n2288 VSS.n2287 2.6005
R961 VSS.n2292 VSS.n2291 2.6005
R962 VSS.n2291 VSS.n2290 2.6005
R963 VSS.n2280 VSS.n2279 2.6005
R964 VSS.n2278 VSS.n2277 2.6005
R965 VSS.n2277 VSS.n2276 2.6005
R966 VSS.n2275 VSS.n2274 2.6005
R967 VSS.n2274 VSS.n2273 2.6005
R968 VSS.n2272 VSS.n2271 2.6005
R969 VSS.n2271 VSS.n2270 2.6005
R970 VSS.n2269 VSS.n2268 2.6005
R971 VSS.n2268 VSS.n2267 2.6005
R972 VSS.n1744 VSS.n1743 2.6005
R973 VSS.n2265 VSS.n2264 2.6005
R974 VSS.n2264 VSS.n2263 2.6005
R975 VSS.n2262 VSS.n2261 2.6005
R976 VSS.n2261 VSS.n2260 2.6005
R977 VSS.n2198 VSS.n2197 2.6005
R978 VSS.n2197 VSS.n2196 2.6005
R979 VSS.n2195 VSS.n2194 2.6005
R980 VSS.n2194 VSS.n2193 2.6005
R981 VSS.n2192 VSS.n2191 2.6005
R982 VSS.n2191 VSS.n2190 2.6005
R983 VSS.n2189 VSS.n2188 2.6005
R984 VSS.n2188 VSS.n2187 2.6005
R985 VSS.n1939 VSS.n1938 2.6005
R986 VSS.n1938 VSS.n1937 2.6005
R987 VSS.n2150 VSS.n2149 2.6005
R988 VSS.n2152 VSS.n2151 2.6005
R989 VSS.n2155 VSS.n2154 2.6005
R990 VSS.n2154 VSS.n2153 2.6005
R991 VSS.n2158 VSS.n2157 2.6005
R992 VSS.n2157 VSS.n2156 2.6005
R993 VSS.n2161 VSS.n2160 2.6005
R994 VSS.n2160 VSS.n2159 2.6005
R995 VSS.n2164 VSS.n2163 2.6005
R996 VSS.n2163 VSS.n2162 2.6005
R997 VSS.n2167 VSS.n2166 2.6005
R998 VSS.n2166 VSS.n2165 2.6005
R999 VSS.n2170 VSS.n2169 2.6005
R1000 VSS.n2169 VSS.n2168 2.6005
R1001 VSS.n2173 VSS.n2172 2.6005
R1002 VSS.n2172 VSS.n2171 2.6005
R1003 VSS.n2176 VSS.n2175 2.6005
R1004 VSS.n2175 VSS.n2174 2.6005
R1005 VSS.n2179 VSS.n2178 2.6005
R1006 VSS.n2178 VSS.n2177 2.6005
R1007 VSS.n2182 VSS.n2181 2.6005
R1008 VSS.n2181 VSS.n2180 2.6005
R1009 VSS.n2148 VSS.n2147 2.6005
R1010 VSS.n2493 VSS.n2492 2.6005
R1011 VSS.n2492 VSS.n2491 2.6005
R1012 VSS.n2496 VSS.n2495 2.6005
R1013 VSS.n2495 VSS.n2494 2.6005
R1014 VSS.n2499 VSS.n2498 2.6005
R1015 VSS.n2498 VSS.n2497 2.6005
R1016 VSS.n2503 VSS.n2502 2.6005
R1017 VSS.n2502 VSS.n2501 2.6005
R1018 VSS.n2506 VSS.n2505 2.6005
R1019 VSS.n2505 VSS.n2504 2.6005
R1020 VSS.n2509 VSS.n2508 2.6005
R1021 VSS.n2508 VSS.n2507 2.6005
R1022 VSS.n2512 VSS.n2511 2.6005
R1023 VSS.n2511 VSS.n2510 2.6005
R1024 VSS.n2515 VSS.n2514 2.6005
R1025 VSS.n2514 VSS.n2513 2.6005
R1026 VSS.n2518 VSS.n2517 2.6005
R1027 VSS.n2517 VSS.n2516 2.6005
R1028 VSS.n2521 VSS.n2520 2.6005
R1029 VSS.n2520 VSS.t153 2.6005
R1030 VSS.n2524 VSS.n2523 2.6005
R1031 VSS.n2523 VSS.n2522 2.6005
R1032 VSS.n2527 VSS.n2526 2.6005
R1033 VSS.n2526 VSS.n2525 2.6005
R1034 VSS.n2530 VSS.n2529 2.6005
R1035 VSS.n2529 VSS.n2528 2.6005
R1036 VSS.n2533 VSS.n2532 2.6005
R1037 VSS.n2532 VSS.n2531 2.6005
R1038 VSS.n2537 VSS.n2536 2.6005
R1039 VSS.n2536 VSS.n2535 2.6005
R1040 VSS.n2540 VSS.n2539 2.6005
R1041 VSS.n2539 VSS.n2538 2.6005
R1042 VSS.n2543 VSS.n2542 2.6005
R1043 VSS.n2542 VSS.n2541 2.6005
R1044 VSS.n2546 VSS.n2545 2.6005
R1045 VSS.n2545 VSS.n2544 2.6005
R1046 VSS.n2549 VSS.n2548 2.6005
R1047 VSS.n2548 VSS.n2547 2.6005
R1048 VSS.n2553 VSS.n2552 2.6005
R1049 VSS.n2552 VSS.n2551 2.6005
R1050 VSS.n2556 VSS.n2555 2.6005
R1051 VSS.n2555 VSS.n2554 2.6005
R1052 VSS.n2559 VSS.n2558 2.6005
R1053 VSS.n2558 VSS.n2557 2.6005
R1054 VSS.n2562 VSS.n2561 2.6005
R1055 VSS.n2561 VSS.n2560 2.6005
R1056 VSS.n2565 VSS.n2564 2.6005
R1057 VSS.n2564 VSS.n2563 2.6005
R1058 VSS.n2568 VSS.n2567 2.6005
R1059 VSS.n2567 VSS.n2566 2.6005
R1060 VSS.n2571 VSS.n2570 2.6005
R1061 VSS.n2570 VSS.n2569 2.6005
R1062 VSS.n2574 VSS.n2573 2.6005
R1063 VSS.n2573 VSS.n2572 2.6005
R1064 VSS.n2577 VSS.n2576 2.6005
R1065 VSS.n2576 VSS.n2575 2.6005
R1066 VSS.n2580 VSS.n2579 2.6005
R1067 VSS.n2579 VSS.n2578 2.6005
R1068 VSS.n2584 VSS.n2583 2.6005
R1069 VSS.n2583 VSS.n2582 2.6005
R1070 VSS.n2588 VSS.n2587 2.6005
R1071 VSS.n2587 VSS.n2586 2.6005
R1072 VSS.n2592 VSS.n2591 2.6005
R1073 VSS.n2591 VSS.n2590 2.6005
R1074 VSS.n2596 VSS.n2595 2.6005
R1075 VSS.n2595 VSS.n2594 2.6005
R1076 VSS.n2600 VSS.n2599 2.6005
R1077 VSS.n2599 VSS.n2598 2.6005
R1078 VSS.n2604 VSS.n2603 2.6005
R1079 VSS.n2603 VSS.n2602 2.6005
R1080 VSS.n2068 VSS.n2067 2.6005
R1081 VSS.n2067 VSS.n2066 2.6005
R1082 VSS.n2072 VSS.n2071 2.6005
R1083 VSS.n2071 VSS.n2070 2.6005
R1084 VSS.n2075 VSS.n2074 2.6005
R1085 VSS.n2074 VSS.n2073 2.6005
R1086 VSS.n2078 VSS.n2077 2.6005
R1087 VSS.n2077 VSS.n2076 2.6005
R1088 VSS.n2079 VSS.n2064 2.6005
R1089 VSS.n2064 VSS.n2063 2.6005
R1090 VSS.n2081 VSS 2.6005
R1091 VSS.n2081 VSS.n2080 2.6005
R1092 VSS.n2084 VSS.n2083 2.6005
R1093 VSS.n2083 VSS.n2082 2.6005
R1094 VSS.n2087 VSS.n2086 2.6005
R1095 VSS.n2086 VSS.n2085 2.6005
R1096 VSS.n2090 VSS.n2089 2.6005
R1097 VSS.n2089 VSS.n2088 2.6005
R1098 VSS.n2093 VSS.n2092 2.6005
R1099 VSS.n2092 VSS.n2091 2.6005
R1100 VSS.n2097 VSS.n2096 2.6005
R1101 VSS.n2096 VSS.n2095 2.6005
R1102 VSS.n2029 VSS.n2028 2.6005
R1103 VSS.n2028 VSS.n2027 2.6005
R1104 VSS.n2033 VSS.n2032 2.6005
R1105 VSS.n2032 VSS.n2031 2.6005
R1106 VSS.n2036 VSS.n2035 2.6005
R1107 VSS.n2035 VSS.n2034 2.6005
R1108 VSS.n2039 VSS.n2038 2.6005
R1109 VSS.n2038 VSS.n2037 2.6005
R1110 VSS.n2040 VSS.n1946 2.6005
R1111 VSS.n1946 VSS.n1945 2.6005
R1112 VSS.n2042 VSS 2.6005
R1113 VSS.n2042 VSS.n2041 2.6005
R1114 VSS.n2045 VSS.n2044 2.6005
R1115 VSS.n2044 VSS.n2043 2.6005
R1116 VSS.n2048 VSS.n2047 2.6005
R1117 VSS.n2047 VSS.n2046 2.6005
R1118 VSS.n2051 VSS.n2050 2.6005
R1119 VSS.n2050 VSS.n2049 2.6005
R1120 VSS.n2054 VSS.n2053 2.6005
R1121 VSS.n2053 VSS.n2052 2.6005
R1122 VSS.n2058 VSS.n2057 2.6005
R1123 VSS.n2057 VSS.n2056 2.6005
R1124 VSS.n1317 VSS.n1313 2.6005
R1125 VSS.n1275 VSS.n1272 2.6005
R1126 VSS.n1279 VSS.n1276 2.6005
R1127 VSS.n1283 VSS.n1281 2.6005
R1128 VSS.n1281 VSS.n1280 2.6005
R1129 VSS.n1294 VSS.n1288 2.6005
R1130 VSS.n1288 VSS.n1287 2.6005
R1131 VSS.n1286 VSS 2.6005
R1132 VSS.n1286 VSS.n1285 2.6005
R1133 VSS.n1303 VSS.n1301 2.6005
R1134 VSS.n1301 VSS.n1300 2.6005
R1135 VSS.n1307 VSS.n1305 2.6005
R1136 VSS.n1305 VSS.n1304 2.6005
R1137 VSS.n1311 VSS.n1309 2.6005
R1138 VSS.n1309 VSS.n1308 2.6005
R1139 VSS.n1269 VSS.n1262 2.6005
R1140 VSS.n1275 VSS.n1274 2.6005
R1141 VSS.n1274 VSS.n1273 2.6005
R1142 VSS.n1279 VSS.n1278 2.6005
R1143 VSS.n1278 VSS.n1277 2.6005
R1144 VSS.n1283 VSS.n1282 2.6005
R1145 VSS.n1295 VSS.n1294 2.6005
R1146 VSS.n1296 VSS 2.6005
R1147 VSS.n1299 VSS.n1298 2.6005
R1148 VSS.n1298 VSS.n1297 2.6005
R1149 VSS.n1303 VSS.n1302 2.6005
R1150 VSS.n1307 VSS.n1306 2.6005
R1151 VSS.n1311 VSS.n1310 2.6005
R1152 VSS.n1317 VSS.n1316 2.6005
R1153 VSS.n1316 VSS.n1315 2.6005
R1154 VSS.n1269 VSS.n1268 2.6005
R1155 VSS.n1268 VSS.n1267 2.6005
R1156 VSS.n1534 VSS.n1533 2.6005
R1157 VSS.n1533 VSS.n1532 2.6005
R1158 VSS.n1531 VSS.n1530 2.6005
R1159 VSS.n1530 VSS.n1529 2.6005
R1160 VSS.n1528 VSS.n1527 2.6005
R1161 VSS.n1527 VSS.n1526 2.6005
R1162 VSS.n1525 VSS.n1524 2.6005
R1163 VSS.n1524 VSS.n1523 2.6005
R1164 VSS.n1522 VSS.n1521 2.6005
R1165 VSS.n1521 VSS.n1520 2.6005
R1166 VSS.n1519 VSS.n1518 2.6005
R1167 VSS.n1518 VSS.n1517 2.6005
R1168 VSS.n1516 VSS.n1515 2.6005
R1169 VSS.n1515 VSS.n1514 2.6005
R1170 VSS.n1513 VSS.n1512 2.6005
R1171 VSS.n1507 VSS.n1506 2.6005
R1172 VSS.n1504 VSS.n1503 2.6005
R1173 VSS.n1501 VSS.n1500 2.6005
R1174 VSS.n1499 VSS.n1498 2.6005
R1175 VSS.n1496 VSS.n1495 2.6005
R1176 VSS.n1494 VSS.n1493 2.6005
R1177 VSS.n1491 VSS.n1490 2.6005
R1178 VSS.n1489 VSS.n1488 2.6005
R1179 VSS.n1487 VSS.n1486 2.6005
R1180 VSS.n1486 VSS.n1485 2.6005
R1181 VSS.n1484 VSS.n1483 2.6005
R1182 VSS.n1483 VSS.n1482 2.6005
R1183 VSS.n1481 VSS.n1480 2.6005
R1184 VSS.n1480 VSS.n1479 2.6005
R1185 VSS.n1478 VSS.n1477 2.6005
R1186 VSS.n1477 VSS.n1476 2.6005
R1187 VSS.n1475 VSS.n1474 2.6005
R1188 VSS.n1474 VSS.n1473 2.6005
R1189 VSS.n1472 VSS.n1471 2.6005
R1190 VSS.n1471 VSS.n1470 2.6005
R1191 VSS.n1469 VSS.n1468 2.6005
R1192 VSS.n1468 VSS.n1467 2.6005
R1193 VSS.n1466 VSS.n1465 2.6005
R1194 VSS.n1465 VSS.n1464 2.6005
R1195 VSS.n1463 VSS.n1462 2.6005
R1196 VSS.n1462 VSS.n1461 2.6005
R1197 VSS.n1460 VSS.n1459 2.6005
R1198 VSS.n1459 VSS.n1458 2.6005
R1199 VSS.n1457 VSS.n1456 2.6005
R1200 VSS.n1456 VSS.n1455 2.6005
R1201 VSS.n1454 VSS.n1453 2.6005
R1202 VSS.n1453 VSS.n1452 2.6005
R1203 VSS.n1451 VSS.n1450 2.6005
R1204 VSS.n1450 VSS.n1449 2.6005
R1205 VSS.n1448 VSS.n1447 2.6005
R1206 VSS.n1447 VSS.n1446 2.6005
R1207 VSS.n1445 VSS.n1444 2.6005
R1208 VSS.n1444 VSS.n1443 2.6005
R1209 VSS.n1442 VSS.n1441 2.6005
R1210 VSS.n1441 VSS.n1440 2.6005
R1211 VSS.n1439 VSS.n1438 2.6005
R1212 VSS.n1438 VSS.n1437 2.6005
R1213 VSS.n1436 VSS.n1435 2.6005
R1214 VSS.n1435 VSS.n1434 2.6005
R1215 VSS.n1433 VSS.n1432 2.6005
R1216 VSS.n1432 VSS.n1431 2.6005
R1217 VSS.n1430 VSS.n1429 2.6005
R1218 VSS.n1429 VSS.n1428 2.6005
R1219 VSS.n1427 VSS.n1426 2.6005
R1220 VSS.n1426 VSS.n1425 2.6005
R1221 VSS.n1424 VSS.n1423 2.6005
R1222 VSS.n1423 VSS.n1422 2.6005
R1223 VSS.n1421 VSS.n1420 2.6005
R1224 VSS.n1420 VSS.n1419 2.6005
R1225 VSS.n1418 VSS.n1417 2.6005
R1226 VSS.n1417 VSS.n1416 2.6005
R1227 VSS.n1415 VSS.n1414 2.6005
R1228 VSS.n1414 VSS.n1413 2.6005
R1229 VSS.n1412 VSS.n1411 2.6005
R1230 VSS.n1411 VSS.n1410 2.6005
R1231 VSS.n1409 VSS.n1408 2.6005
R1232 VSS.n1408 VSS.n1407 2.6005
R1233 VSS.n1406 VSS.n1405 2.6005
R1234 VSS.n1405 VSS.n1404 2.6005
R1235 VSS.n1403 VSS.n1402 2.6005
R1236 VSS.n1402 VSS.n1401 2.6005
R1237 VSS.n1400 VSS.n1399 2.6005
R1238 VSS.n1399 VSS.n1398 2.6005
R1239 VSS.n1397 VSS.n1396 2.6005
R1240 VSS.n1396 VSS.n1395 2.6005
R1241 VSS.n1394 VSS.n1393 2.6005
R1242 VSS.n1393 VSS.n1392 2.6005
R1243 VSS.n1391 VSS.n1390 2.6005
R1244 VSS.n1390 VSS.n1389 2.6005
R1245 VSS.n1388 VSS.n1387 2.6005
R1246 VSS.n1387 VSS.n1386 2.6005
R1247 VSS.n1385 VSS.n1384 2.6005
R1248 VSS.n1384 VSS.n1383 2.6005
R1249 VSS.n1381 VSS.n1380 2.6005
R1250 VSS.n1380 VSS.n1379 2.6005
R1251 VSS.n1378 VSS.n1377 2.6005
R1252 VSS.n1377 VSS.n1376 2.6005
R1253 VSS.n2609 VSS.n2608 2.6005
R1254 VSS.n2608 VSS.n2607 2.6005
R1255 VSS.n2614 VSS.n2613 2.6005
R1256 VSS.n2613 VSS.n2612 2.6005
R1257 VSS.n2618 VSS.n2617 2.6005
R1258 VSS.n2617 VSS.n2616 2.6005
R1259 VSS.n2622 VSS.n2621 2.6005
R1260 VSS.n2621 VSS.n2620 2.6005
R1261 VSS.n2625 VSS.n2624 2.6005
R1262 VSS.n2624 VSS.n2623 2.6005
R1263 VSS.n2629 VSS.n2628 2.6005
R1264 VSS.n2628 VSS.n2627 2.6005
R1265 VSS.n2632 VSS.n2631 2.6005
R1266 VSS.n2631 VSS.n2630 2.6005
R1267 VSS.n2635 VSS.n2634 2.6005
R1268 VSS.n2634 VSS.n2633 2.6005
R1269 VSS.n2638 VSS.n2637 2.6005
R1270 VSS.n2637 VSS.n2636 2.6005
R1271 VSS.n2642 VSS.n2641 2.6005
R1272 VSS.n2641 VSS.n2640 2.6005
R1273 VSS.n2645 VSS.n2644 2.6005
R1274 VSS.n2644 VSS.n2643 2.6005
R1275 VSS.n2648 VSS.n2647 2.6005
R1276 VSS.n2647 VSS.n2646 2.6005
R1277 VSS.n2651 VSS.n2650 2.6005
R1278 VSS.n2650 VSS.n2649 2.6005
R1279 VSS.n2654 VSS.n2653 2.6005
R1280 VSS.n2653 VSS.n2652 2.6005
R1281 VSS.n2657 VSS.n2656 2.6005
R1282 VSS.n2656 VSS.n2655 2.6005
R1283 VSS.n2660 VSS.n2659 2.6005
R1284 VSS.n2659 VSS.n2658 2.6005
R1285 VSS.n2664 VSS.n2663 2.6005
R1286 VSS.n2663 VSS.n2662 2.6005
R1287 VSS.n2666 VSS.n2665 2.6005
R1288 VSS.n2670 VSS.n2669 2.6005
R1289 VSS.n2669 VSS.n2668 2.6005
R1290 VSS.n2673 VSS.n2672 2.6005
R1291 VSS.n2672 VSS.n2671 2.6005
R1292 VSS.n2676 VSS.n2675 2.6005
R1293 VSS.n2675 VSS.n2674 2.6005
R1294 VSS.n2679 VSS.n2678 2.6005
R1295 VSS.n2678 VSS.n2677 2.6005
R1296 VSS.n2682 VSS.n2681 2.6005
R1297 VSS.n2681 VSS.n2680 2.6005
R1298 VSS.n2685 VSS.n2684 2.6005
R1299 VSS.n2684 VSS.n2683 2.6005
R1300 VSS.n2688 VSS.n2687 2.6005
R1301 VSS.n2687 VSS.n2686 2.6005
R1302 VSS.n2804 VSS.n2803 2.6005
R1303 VSS.n2803 VSS.n2802 2.6005
R1304 VSS.n2807 VSS.n2806 2.6005
R1305 VSS.n2806 VSS.n2805 2.6005
R1306 VSS.n2738 VSS.n2737 2.6005
R1307 VSS.n2737 VSS.n2736 2.6005
R1308 VSS.n2741 VSS.n2740 2.6005
R1309 VSS.n2740 VSS.n2739 2.6005
R1310 VSS.n2744 VSS.n2743 2.6005
R1311 VSS.n2743 VSS.n2742 2.6005
R1312 VSS.n2747 VSS.n2746 2.6005
R1313 VSS.n2746 VSS.n2745 2.6005
R1314 VSS.n2750 VSS.n2749 2.6005
R1315 VSS.n2749 VSS.n2748 2.6005
R1316 VSS.n2753 VSS.n2752 2.6005
R1317 VSS.n2752 VSS.n2751 2.6005
R1318 VSS.n2756 VSS.n2755 2.6005
R1319 VSS.n2755 VSS.n2754 2.6005
R1320 VSS.n2759 VSS.n2758 2.6005
R1321 VSS.n2758 VSS.n2757 2.6005
R1322 VSS.n2762 VSS.n2761 2.6005
R1323 VSS.n2761 VSS.n2760 2.6005
R1324 VSS.n2765 VSS.n2764 2.6005
R1325 VSS.n2764 VSS.n2763 2.6005
R1326 VSS.n2768 VSS.n2767 2.6005
R1327 VSS.n2767 VSS.n2766 2.6005
R1328 VSS.n2771 VSS.n2770 2.6005
R1329 VSS.n2770 VSS.n2769 2.6005
R1330 VSS.n2774 VSS.n2773 2.6005
R1331 VSS.n2773 VSS.n2772 2.6005
R1332 VSS.n2777 VSS.n2776 2.6005
R1333 VSS.n2776 VSS.n2775 2.6005
R1334 VSS.n2780 VSS.n2779 2.6005
R1335 VSS.n2779 VSS.n2778 2.6005
R1336 VSS.n2783 VSS.n2782 2.6005
R1337 VSS.n2782 VSS.n2781 2.6005
R1338 VSS.n2786 VSS.n2785 2.6005
R1339 VSS.n2785 VSS.n2784 2.6005
R1340 VSS.n2789 VSS.n2788 2.6005
R1341 VSS.n2788 VSS.n2787 2.6005
R1342 VSS.n2792 VSS.n2791 2.6005
R1343 VSS.n2791 VSS.n2790 2.6005
R1344 VSS.n2795 VSS.n2794 2.6005
R1345 VSS.n2794 VSS.n2793 2.6005
R1346 VSS.n2798 VSS.n2797 2.6005
R1347 VSS.n2797 VSS.n2796 2.6005
R1348 VSS.n2801 VSS.n2800 2.6005
R1349 VSS.n2800 VSS.n2799 2.6005
R1350 VSS.n2732 VSS.n2731 2.6005
R1351 VSS.n2735 VSS.n2734 2.6005
R1352 VSS.n2708 VSS.n2707 2.6005
R1353 VSS.n2707 VSS.n2706 2.6005
R1354 VSS.n2711 VSS.n2710 2.6005
R1355 VSS.n2710 VSS.n2709 2.6005
R1356 VSS.n2714 VSS.n2713 2.6005
R1357 VSS.n2713 VSS.n2712 2.6005
R1358 VSS.n2717 VSS.n2716 2.6005
R1359 VSS.n2716 VSS.n2715 2.6005
R1360 VSS.n2720 VSS.n2719 2.6005
R1361 VSS.n2719 VSS.n2718 2.6005
R1362 VSS.n2723 VSS.n2722 2.6005
R1363 VSS.n2722 VSS.n2721 2.6005
R1364 VSS.n2726 VSS.n2725 2.6005
R1365 VSS.n2725 VSS.n2724 2.6005
R1366 VSS.n2730 VSS.n2729 2.6005
R1367 VSS.n2729 VSS.n2728 2.6005
R1368 VSS.n2691 VSS.n2690 2.6005
R1369 VSS.n2693 VSS.n2692 2.6005
R1370 VSS.n2696 VSS.n2695 2.6005
R1371 VSS.n2699 VSS.n2698 2.6005
R1372 VSS.n2703 VSS.n2702 2.6005
R1373 VSS.n1985 VSS.n1984 2.6005
R1374 VSS.n1984 VSS.n1983 2.6005
R1375 VSS.n1960 VSS.n1959 2.6005
R1376 VSS.n1959 VSS.n1958 2.6005
R1377 VSS.n1963 VSS.n1962 2.6005
R1378 VSS.n1962 VSS.n1961 2.6005
R1379 VSS.n1966 VSS.n1965 2.6005
R1380 VSS.n1965 VSS.n1964 2.6005
R1381 VSS.n1967 VSS.n1952 2.6005
R1382 VSS.n1952 VSS.n1951 2.6005
R1383 VSS.n1969 VSS 2.6005
R1384 VSS.n1969 VSS.n1968 2.6005
R1385 VSS.n1972 VSS.n1971 2.6005
R1386 VSS.n1971 VSS.n1970 2.6005
R1387 VSS.n1975 VSS.n1974 2.6005
R1388 VSS.n1974 VSS.n1973 2.6005
R1389 VSS.n1978 VSS.n1977 2.6005
R1390 VSS.n1977 VSS.n1976 2.6005
R1391 VSS.n1981 VSS.n1980 2.6005
R1392 VSS.n1980 VSS.n1979 2.6005
R1393 VSS.n1956 VSS.n1955 2.6005
R1394 VSS.n1993 VSS.n1992 2.6005
R1395 VSS.n1997 VSS.n1996 2.6005
R1396 VSS.n1996 VSS.n1995 2.6005
R1397 VSS.n2000 VSS.n1999 2.6005
R1398 VSS.n1999 VSS.n1998 2.6005
R1399 VSS.n2003 VSS.n2002 2.6005
R1400 VSS.n2002 VSS.n2001 2.6005
R1401 VSS.n2004 VSS.n1990 2.6005
R1402 VSS.n1990 VSS.n1989 2.6005
R1403 VSS.n2006 VSS 2.6005
R1404 VSS.n2006 VSS.n2005 2.6005
R1405 VSS.n2009 VSS.n2008 2.6005
R1406 VSS.n2008 VSS.n2007 2.6005
R1407 VSS.n2012 VSS.n2011 2.6005
R1408 VSS.n2011 VSS.n2010 2.6005
R1409 VSS.n2015 VSS.n2014 2.6005
R1410 VSS.n2014 VSS.n2013 2.6005
R1411 VSS.n2018 VSS.n2017 2.6005
R1412 VSS.n2017 VSS.n2016 2.6005
R1413 VSS.n2022 VSS.n2021 2.6005
R1414 VSS.n2021 VSS.n2020 2.6005
R1415 VSS.n1255 VSS.n811 2.6005
R1416 VSS.n811 VSS.n810 2.6005
R1417 VSS.n805 VSS.n804 2.6005
R1418 VSS.n804 VSS.n803 2.6005
R1419 VSS.n802 VSS.n801 2.6005
R1420 VSS.n801 VSS.n800 2.6005
R1421 VSS.n798 VSS.n797 2.6005
R1422 VSS.n797 VSS.n796 2.6005
R1423 VSS.n795 VSS.n794 2.6005
R1424 VSS.n794 VSS.n793 2.6005
R1425 VSS.n792 VSS.n791 2.6005
R1426 VSS.n791 VSS.n790 2.6005
R1427 VSS.n788 VSS.n787 2.6005
R1428 VSS.n787 VSS.n786 2.6005
R1429 VSS.n785 VSS.n784 2.6005
R1430 VSS.n784 VSS.n783 2.6005
R1431 VSS.n1092 VSS.n1091 2.6005
R1432 VSS.n1091 VSS.n1090 2.6005
R1433 VSS.n1098 VSS.n1097 2.6005
R1434 VSS.n1094 VSS.n1093 2.6005
R1435 VSS.n808 VSS.n807 2.6005
R1436 VSS.n807 VSS.n806 2.6005
R1437 VSS.n1240 VSS.n1239 2.6005
R1438 VSS.n1239 VSS.n1238 2.6005
R1439 VSS.n1243 VSS.n1242 2.6005
R1440 VSS.n1242 VSS.n1241 2.6005
R1441 VSS.n1247 VSS.n1246 2.6005
R1442 VSS.n1246 VSS.n1245 2.6005
R1443 VSS.n1250 VSS.n1249 2.6005
R1444 VSS.n1249 VSS.n1248 2.6005
R1445 VSS.n1253 VSS.n1252 2.6005
R1446 VSS.n1252 VSS.n1251 2.6005
R1447 VSS.n1223 VSS.n1222 2.6005
R1448 VSS.n1222 VSS.n1221 2.6005
R1449 VSS.n1227 VSS.n1226 2.6005
R1450 VSS.n1229 VSS.n1228 2.6005
R1451 VSS.n1232 VSS.n1231 2.6005
R1452 VSS.n1235 VSS.n1234 2.6005
R1453 VSS.n1237 VSS.n1236 2.6005
R1454 VSS.n1259 VSS.n1258 2.6005
R1455 VSS.n1258 VSS.n1257 2.6005
R1456 VSS.n1571 VSS.n1570 2.6005
R1457 VSS.n1566 VSS.n1565 2.6005
R1458 VSS.n1564 VSS.n1563 2.6005
R1459 VSS.n1561 VSS.n1560 2.6005
R1460 VSS.n1559 VSS.n1558 2.6005
R1461 VSS.n1556 VSS.n1555 2.6005
R1462 VSS.n1554 VSS.n1553 2.6005
R1463 VSS.n1551 VSS.n1550 2.6005
R1464 VSS.n1549 VSS.n1548 2.6005
R1465 VSS.n1546 VSS.n1545 2.6005
R1466 VSS.n1544 VSS.n1543 2.6005
R1467 VSS.n1541 VSS.n1540 2.6005
R1468 VSS.n1539 VSS.n1538 2.6005
R1469 VSS.n1536 VSS.n1535 2.6005
R1470 VSS.n1123 VSS.n1122 2.6005
R1471 VSS.n1122 VSS.n1121 2.6005
R1472 VSS.n1119 VSS.n1118 2.6005
R1473 VSS.n1118 VSS.n1117 2.6005
R1474 VSS.n1116 VSS.n1115 2.6005
R1475 VSS.n1115 VSS.n1114 2.6005
R1476 VSS.n1113 VSS.n1112 2.6005
R1477 VSS.n1112 VSS.n1111 2.6005
R1478 VSS.n1110 VSS.n1109 2.6005
R1479 VSS.n1109 VSS.n1108 2.6005
R1480 VSS.n1107 VSS.n1106 2.6005
R1481 VSS.n1106 VSS.n1105 2.6005
R1482 VSS.n1104 VSS.n1103 2.6005
R1483 VSS.n1103 VSS.n1102 2.6005
R1484 VSS.n1101 VSS.n1100 2.6005
R1485 VSS.n1100 VSS.n1099 2.6005
R1486 VSS.n1195 VSS.n1194 2.6005
R1487 VSS.n1194 VSS.n1193 2.6005
R1488 VSS.n1198 VSS.n1197 2.6005
R1489 VSS.n1197 VSS.n1196 2.6005
R1490 VSS.n1201 VSS.n1200 2.6005
R1491 VSS.n1200 VSS.n1199 2.6005
R1492 VSS.n1204 VSS.n1203 2.6005
R1493 VSS.n1203 VSS.n1202 2.6005
R1494 VSS.n1207 VSS.n1206 2.6005
R1495 VSS.n1206 VSS.n1205 2.6005
R1496 VSS.n1210 VSS.n1209 2.6005
R1497 VSS.n1209 VSS.n1208 2.6005
R1498 VSS.n1213 VSS.n1212 2.6005
R1499 VSS.n1212 VSS.n1211 2.6005
R1500 VSS.n1217 VSS.n1216 2.6005
R1501 VSS.n1216 VSS.n1215 2.6005
R1502 VSS.n1592 VSS.n1591 2.6005
R1503 VSS.n1591 VSS.n1590 2.6005
R1504 VSS.n1589 VSS.n1588 2.6005
R1505 VSS.n1588 VSS.n1587 2.6005
R1506 VSS.n1586 VSS.n1585 2.6005
R1507 VSS.n1585 VSS.n1584 2.6005
R1508 VSS.n1583 VSS.n1582 2.6005
R1509 VSS.n1582 VSS.n1581 2.6005
R1510 VSS.n1580 VSS.n1579 2.6005
R1511 VSS.n1579 VSS.n1578 2.6005
R1512 VSS.n1577 VSS.n1576 2.6005
R1513 VSS.n1576 VSS.n1575 2.6005
R1514 VSS.n1574 VSS.n1573 2.6005
R1515 VSS.n1573 VSS.n1572 2.6005
R1516 VSS.n1129 VSS.n1128 2.6005
R1517 VSS.n1125 VSS.n1124 2.6005
R1518 VSS.n1192 VSS.n1191 2.6005
R1519 VSS.n1597 VSS.n1596 2.6005
R1520 VSS.n1594 VSS.n1593 2.6005
R1521 VSS.n377 VSS.n373 2.6005
R1522 VSS.n373 VSS.n372 2.6005
R1523 VSS.n335 VSS.n334 2.6005
R1524 VSS.n334 VSS.n333 2.6005
R1525 VSS.n341 VSS.n340 2.6005
R1526 VSS.n340 VSS.n339 2.6005
R1527 VSS.n347 VSS.n346 2.6005
R1528 VSS.n346 VSS.n345 2.6005
R1529 VSS.n361 VSS.n359 2.6005
R1530 VSS.n361 VSS.n360 2.6005
R1531 VSS VSS.n363 2.6005
R1532 VSS.n363 VSS.n362 2.6005
R1533 VSS.n403 VSS.n402 2.6005
R1534 VSS.n402 VSS.n401 2.6005
R1535 VSS.n396 VSS.n395 2.6005
R1536 VSS.n395 VSS.n394 2.6005
R1537 VSS.n390 VSS.n389 2.6005
R1538 VSS.n389 VSS.n388 2.6005
R1539 VSS.n384 VSS.n383 2.6005
R1540 VSS.n383 VSS.n382 2.6005
R1541 VSS.n328 VSS.n327 2.6005
R1542 VSS VSS.n371 2.6005
R1543 VSS.n371 VSS.n370 2.6005
R1544 VSS.n400 VSS.n399 2.6005
R1545 VSS.n399 VSS.n398 2.6005
R1546 VSS.n393 VSS.n392 2.6005
R1547 VSS.n392 VSS.n391 2.6005
R1548 VSS.n387 VSS.n386 2.6005
R1549 VSS.n386 VSS.n385 2.6005
R1550 VSS.n381 VSS.n380 2.6005
R1551 VSS.n380 VSS.n379 2.6005
R1552 VSS.n376 VSS.n375 2.6005
R1553 VSS.n331 VSS.n330 2.6005
R1554 VSS.n330 VSS.n329 2.6005
R1555 VSS.n338 VSS.n337 2.6005
R1556 VSS.n337 VSS.n336 2.6005
R1557 VSS.n344 VSS.n343 2.6005
R1558 VSS.n343 VSS.n342 2.6005
R1559 VSS.n350 VSS.n349 2.6005
R1560 VSS.n349 VSS.n348 2.6005
R1561 VSS.n367 VSS.n365 2.6005
R1562 VSS.n367 VSS.n366 2.6005
R1563 VSS.n879 VSS.n878 2.6005
R1564 VSS.n878 VSS.n877 2.6005
R1565 VSS.n876 VSS.n875 2.6005
R1566 VSS.n875 VSS.n874 2.6005
R1567 VSS.n911 VSS.n910 2.6005
R1568 VSS.n910 VSS.n909 2.6005
R1569 VSS.n907 VSS.n906 2.6005
R1570 VSS.n906 VSS.n905 2.6005
R1571 VSS.n904 VSS.n903 2.6005
R1572 VSS.n903 VSS.n902 2.6005
R1573 VSS.n901 VSS.n900 2.6005
R1574 VSS.n900 VSS.n899 2.6005
R1575 VSS.n891 VSS.n890 2.6005
R1576 VSS.n890 VSS.n889 2.6005
R1577 VSS.n897 VSS.n896 2.6005
R1578 VSS.n896 VSS.n895 2.6005
R1579 VSS.n894 VSS.n893 2.6005
R1580 VSS.n893 VSS.n892 2.6005
R1581 VSS.n824 VSS.n823 2.6005
R1582 VSS.n823 VSS.n822 2.6005
R1583 VSS.n919 VSS.n918 2.6005
R1584 VSS.n918 VSS.n917 2.6005
R1585 VSS.n923 VSS.n922 2.6005
R1586 VSS.n922 VSS.n921 2.6005
R1587 VSS.n943 VSS.n942 2.6005
R1588 VSS.n942 VSS.n941 2.6005
R1589 VSS.n947 VSS.n946 2.6005
R1590 VSS.n946 VSS.n945 2.6005
R1591 VSS.n950 VSS.n949 2.6005
R1592 VSS.n949 VSS.n948 2.6005
R1593 VSS.n954 VSS.n953 2.6005
R1594 VSS.n953 VSS.n952 2.6005
R1595 VSS.n957 VSS.n956 2.6005
R1596 VSS.n956 VSS.n955 2.6005
R1597 VSS.n960 VSS.n959 2.6005
R1598 VSS.n959 VSS.n958 2.6005
R1599 VSS.n963 VSS.n962 2.6005
R1600 VSS.n962 VSS.n961 2.6005
R1601 VSS.n966 VSS.n965 2.6005
R1602 VSS.n965 VSS.n964 2.6005
R1603 VSS.n1187 VSS.n1186 2.6005
R1604 VSS.n1184 VSS.n1183 2.6005
R1605 VSS.n1173 VSS.n1172 2.6005
R1606 VSS.n1170 VSS.n1169 2.6005
R1607 VSS.n1166 VSS.n1165 2.6005
R1608 VSS.n1162 VSS.n1161 2.6005
R1609 VSS.n1011 VSS.n1010 2.6005
R1610 VSS.n1010 VSS.n1009 2.6005
R1611 VSS.n1020 VSS.n1019 2.6005
R1612 VSS.n1019 VSS.n1018 2.6005
R1613 VSS.n1024 VSS.n1023 2.6005
R1614 VSS.n1023 VSS.n1022 2.6005
R1615 VSS.n1027 VSS.n1026 2.6005
R1616 VSS.n1026 VSS.n1025 2.6005
R1617 VSS.n1030 VSS.n1029 2.6005
R1618 VSS.n1029 VSS.n1028 2.6005
R1619 VSS.n1033 VSS.n1032 2.6005
R1620 VSS.n1032 VSS.n1031 2.6005
R1621 VSS.n1036 VSS.n1035 2.6005
R1622 VSS.n1035 VSS.n1034 2.6005
R1623 VSS.n1039 VSS.n1038 2.6005
R1624 VSS.n1038 VSS.n1037 2.6005
R1625 VSS.n1042 VSS.n1041 2.6005
R1626 VSS.n1041 VSS.n1040 2.6005
R1627 VSS.n1045 VSS.n1044 2.6005
R1628 VSS.n1044 VSS.n1043 2.6005
R1629 VSS.n1048 VSS.n1047 2.6005
R1630 VSS.n1047 VSS.n1046 2.6005
R1631 VSS.n1051 VSS.n1050 2.6005
R1632 VSS.n1050 VSS.n1049 2.6005
R1633 VSS.n1054 VSS.n1053 2.6005
R1634 VSS.n1053 VSS.n1052 2.6005
R1635 VSS.n1057 VSS.n1056 2.6005
R1636 VSS.n1056 VSS.n1055 2.6005
R1637 VSS.n1060 VSS.n1059 2.6005
R1638 VSS.n1059 VSS.n1058 2.6005
R1639 VSS.n1063 VSS.n1062 2.6005
R1640 VSS.n1062 VSS.n1061 2.6005
R1641 VSS.n1066 VSS.n1065 2.6005
R1642 VSS.n1065 VSS.n1064 2.6005
R1643 VSS.n1132 VSS.n1131 2.6005
R1644 VSS.n1131 VSS.n1130 2.6005
R1645 VSS.n1134 VSS.n1133 2.6005
R1646 VSS.n1138 VSS.n1137 2.6005
R1647 VSS.n1137 VSS.n1136 2.6005
R1648 VSS.n1069 VSS.n1068 2.6005
R1649 VSS.n1068 VSS.n1067 2.6005
R1650 VSS.n1072 VSS.n1071 2.6005
R1651 VSS.n1071 VSS.n1070 2.6005
R1652 VSS.n1075 VSS.n1074 2.6005
R1653 VSS.n1074 VSS.n1073 2.6005
R1654 VSS.n1078 VSS.n1077 2.6005
R1655 VSS.n1077 VSS.n1076 2.6005
R1656 VSS.n1014 VSS.n1013 2.6005
R1657 VSS.n1013 VSS.n1012 2.6005
R1658 VSS.n1017 VSS.n1016 2.6005
R1659 VSS.n1016 VSS.n1015 2.6005
R1660 VSS.n1148 VSS.n1147 2.6005
R1661 VSS.n1145 VSS.n1144 2.6005
R1662 VSS.n1143 VSS.n1142 2.6005
R1663 VSS.n1140 VSS.n1139 2.6005
R1664 VSS.n1152 VSS.n1151 2.6005
R1665 VSS.n1155 VSS.n1154 2.6005
R1666 VSS.n1008 VSS.n1007 2.6005
R1667 VSS.n1006 VSS.n1005 2.6005
R1668 VSS.n1003 VSS.n1002 2.6005
R1669 VSS.n1707 VSS.n1706 2.6005
R1670 VSS.n1704 VSS.n1703 2.6005
R1671 VSS.n1701 VSS.n1700 2.6005
R1672 VSS.n1698 VSS.n1697 2.6005
R1673 VSS.n1696 VSS.n1695 2.6005
R1674 VSS.n1694 VSS.n1693 2.6005
R1675 VSS.n1692 VSS.n1691 2.6005
R1676 VSS.n1710 VSS.n1709 2.6005
R1677 VSS.n1713 VSS.n1712 2.6005
R1678 VSS.n1715 VSS.n1714 2.6005
R1679 VSS.n1718 VSS.n1717 2.6005
R1680 VSS.n1720 VSS.n1719 2.6005
R1681 VSS.n1723 VSS.n1722 2.6005
R1682 VSS.n1725 VSS.n1724 2.6005
R1683 VSS.n748 VSS.n747 2.6005
R1684 VSS.n774 VSS.n773 2.6005
R1685 VSS.n735 VSS.n734 2.6005
R1686 VSS.n738 VSS.n737 2.6005
R1687 VSS.n741 VSS.n740 2.6005
R1688 VSS.n744 VSS.n743 2.6005
R1689 VSS.n870 VSS.n869 2.6005
R1690 VSS.n872 VSS.n871 2.6005
R1691 VSS.n1729 VSS.n1728 2.6005
R1692 VSS.n3028 VSS.n3027 2.6005
R1693 VSS.n3031 VSS.n3030 2.6005
R1694 VSS.n3034 VSS.n3033 2.6005
R1695 VSS.n3037 VSS.n3036 2.6005
R1696 VSS.n3039 VSS.n3038 2.6005
R1697 VSS.n1732 VSS.n1731 2.6005
R1698 VSS.n1159 VSS.n1158 2.6005
R1699 VSS.n1176 VSS.n1175 2.6005
R1700 VSS.n883 VSS.n882 2.6005
R1701 VSS.n1190 VSS.n1189 2.6005
R1702 VSS.n1688 VSS.n1687 2.6005
R1703 VSS.n1687 VSS.n1686 2.6005
R1704 VSS.n1685 VSS.n1684 2.6005
R1705 VSS.n1684 VSS.n1683 2.6005
R1706 VSS.n1682 VSS.n1681 2.6005
R1707 VSS.n1681 VSS.n1680 2.6005
R1708 VSS.n1679 VSS.n1678 2.6005
R1709 VSS.n1678 VSS.n1677 2.6005
R1710 VSS.n1676 VSS.n1675 2.6005
R1711 VSS.n1675 VSS.n1674 2.6005
R1712 VSS.n1673 VSS.n1672 2.6005
R1713 VSS.n1672 VSS.n1671 2.6005
R1714 VSS.n1670 VSS.n1669 2.6005
R1715 VSS.n1669 VSS.n1668 2.6005
R1716 VSS.n1667 VSS.n1666 2.6005
R1717 VSS.n1666 VSS.n1665 2.6005
R1718 VSS.n1664 VSS.n1663 2.6005
R1719 VSS.n1663 VSS.n1662 2.6005
R1720 VSS.n1661 VSS.n1660 2.6005
R1721 VSS.n1660 VSS.n1659 2.6005
R1722 VSS.n1658 VSS.n1657 2.6005
R1723 VSS.n1657 VSS.n1656 2.6005
R1724 VSS.n1655 VSS.n1654 2.6005
R1725 VSS.n1654 VSS.n1653 2.6005
R1726 VSS.n1652 VSS.n1651 2.6005
R1727 VSS.n1651 VSS.n1650 2.6005
R1728 VSS.n1649 VSS.n1648 2.6005
R1729 VSS.n1648 VSS.n1647 2.6005
R1730 VSS.n1646 VSS.n1645 2.6005
R1731 VSS.n1645 VSS.n1644 2.6005
R1732 VSS.n1643 VSS.n1642 2.6005
R1733 VSS.n1642 VSS.n1641 2.6005
R1734 VSS.n1640 VSS.n1639 2.6005
R1735 VSS.n1639 VSS.n1638 2.6005
R1736 VSS.n1637 VSS.n1636 2.6005
R1737 VSS.n1636 VSS.n1635 2.6005
R1738 VSS.n1634 VSS.n1633 2.6005
R1739 VSS.n1633 VSS.n1632 2.6005
R1740 VSS.n1631 VSS.n1630 2.6005
R1741 VSS.n1630 VSS.n1629 2.6005
R1742 VSS.n1628 VSS.n1627 2.6005
R1743 VSS.n1627 VSS.n1626 2.6005
R1744 VSS.n1625 VSS.n1624 2.6005
R1745 VSS.n1624 VSS.n1623 2.6005
R1746 VSS.n1622 VSS.n1621 2.6005
R1747 VSS.n1621 VSS.n1620 2.6005
R1748 VSS.n1619 VSS.n1618 2.6005
R1749 VSS.n1618 VSS.n1617 2.6005
R1750 VSS.n1616 VSS.n1615 2.6005
R1751 VSS.n1615 VSS.n1614 2.6005
R1752 VSS.n1613 VSS.n1612 2.6005
R1753 VSS.n1612 VSS.n1611 2.6005
R1754 VSS.n1610 VSS.n1609 2.6005
R1755 VSS.n1609 VSS.n1608 2.6005
R1756 VSS.n1607 VSS.n1606 2.6005
R1757 VSS.n1606 VSS.n1605 2.6005
R1758 VSS.n1604 VSS.n1603 2.6005
R1759 VSS.n1603 VSS.n1602 2.6005
R1760 VSS.n1601 VSS.n1600 2.6005
R1761 VSS.n1600 VSS.n1599 2.6005
R1762 VSS.n621 VSS.n620 2.6005
R1763 VSS.n620 VSS.n619 2.6005
R1764 VSS.n680 VSS.n677 2.6005
R1765 VSS.n644 VSS.n636 2.6005
R1766 VSS.n625 VSS.n624 2.6005
R1767 VSS.n624 VSS.n623 2.6005
R1768 VSS.n628 VSS.n627 2.6005
R1769 VSS.n627 VSS.n626 2.6005
R1770 VSS.n631 VSS.n630 2.6005
R1771 VSS.n630 VSS.n629 2.6005
R1772 VSS.n645 VSS.n644 2.6005
R1773 VSS.n641 VSS 2.6005
R1774 VSS.n641 VSS.n640 2.6005
R1775 VSS.n667 VSS.n666 2.6005
R1776 VSS.n671 VSS.n670 2.6005
R1777 VSS.n670 VSS.n669 2.6005
R1778 VSS.n681 VSS.n680 2.6005
R1779 VSS.n685 VSS.n684 2.6005
R1780 VSS.n684 VSS.n683 2.6005
R1781 VSS.n689 VSS.n688 2.6005
R1782 VSS.n688 VSS.n687 2.6005
R1783 VSS.n560 VSS.n559 2.6005
R1784 VSS.n2828 VSS.n2827 2.6005
R1785 VSS.n1738 VSS.n1737 2.6005
R1786 VSS.n1740 VSS.n1739 2.6005
R1787 VSS.n2841 VSS.n2840 2.6005
R1788 VSS.n2840 VSS.n2839 2.6005
R1789 VSS.n2844 VSS.n2843 2.6005
R1790 VSS.n2843 VSS.n2842 2.6005
R1791 VSS.n2847 VSS.n2846 2.6005
R1792 VSS.n2846 VSS.n2845 2.6005
R1793 VSS.n2850 VSS.n2849 2.6005
R1794 VSS.n2849 VSS.n2848 2.6005
R1795 VSS.n2853 VSS.n2852 2.6005
R1796 VSS.n2852 VSS.n2851 2.6005
R1797 VSS.n2857 VSS.n2856 2.6005
R1798 VSS.n2856 VSS.n2855 2.6005
R1799 VSS.n2860 VSS.n2859 2.6005
R1800 VSS.n2859 VSS.n2858 2.6005
R1801 VSS.n2863 VSS.n2862 2.6005
R1802 VSS.n2862 VSS.n2861 2.6005
R1803 VSS.n2866 VSS.n2865 2.6005
R1804 VSS.n2865 VSS.n2864 2.6005
R1805 VSS.n2869 VSS.n2868 2.6005
R1806 VSS.n2868 VSS.n2867 2.6005
R1807 VSS.n1735 VSS.n1734 2.6005
R1808 VSS.n1734 VSS.n1733 2.6005
R1809 VSS.n2873 VSS.n2872 2.6005
R1810 VSS.n2872 VSS.n2871 2.6005
R1811 VSS.n2876 VSS.n2875 2.6005
R1812 VSS.n2875 VSS.n2874 2.6005
R1813 VSS.n2879 VSS.n2878 2.6005
R1814 VSS.n2878 VSS.n2877 2.6005
R1815 VSS.n2882 VSS.n2881 2.6005
R1816 VSS.n2881 VSS.n2880 2.6005
R1817 VSS.n2885 VSS.n2884 2.6005
R1818 VSS.n2884 VSS.n2883 2.6005
R1819 VSS.n2837 VSS.n2836 2.6005
R1820 VSS.n2836 VSS.n2835 2.6005
R1821 VSS.n2834 VSS.n2833 2.6005
R1822 VSS.n2833 VSS.n2832 2.6005
R1823 VSS.n2831 VSS.n2830 2.6005
R1824 VSS.n2830 VSS.n2829 2.6005
R1825 VSS.n2810 VSS.n2809 2.6005
R1826 VSS.n2812 VSS.n2811 2.6005
R1827 VSS.n2815 VSS.n2814 2.6005
R1828 VSS.n2818 VSS.n2817 2.6005
R1829 VSS.n2822 VSS.n2821 2.6005
R1830 VSS.n2824 VSS.n2823 2.6005
R1831 VSS.n3021 VSS.n3020 2.6005
R1832 VSS.n533 VSS.n529 2.6005
R1833 VSS.n529 VSS.n528 2.6005
R1834 VSS.n471 VSS.n470 2.6005
R1835 VSS.n470 VSS.n469 2.6005
R1836 VSS.n477 VSS.n476 2.6005
R1837 VSS.n476 VSS.n475 2.6005
R1838 VSS.n483 VSS.n482 2.6005
R1839 VSS.n482 VSS.n481 2.6005
R1840 VSS.n489 VSS.n488 2.6005
R1841 VSS.n488 VSS.n487 2.6005
R1842 VSS.n508 VSS 2.6005
R1843 VSS.n508 VSS.n507 2.6005
R1844 VSS.n511 VSS.n510 2.6005
R1845 VSS.n510 VSS.n509 2.6005
R1846 VSS.n517 VSS.n516 2.6005
R1847 VSS.n516 VSS.n515 2.6005
R1848 VSS.n524 VSS.n523 2.6005
R1849 VSS.n523 VSS.n522 2.6005
R1850 VSS.n540 VSS.n539 2.6005
R1851 VSS.n539 VSS.n538 2.6005
R1852 VSS.n464 VSS.n463 2.6005
R1853 VSS.n505 VSS.n502 2.6005
R1854 VSS.n474 VSS.n473 2.6005
R1855 VSS.n473 VSS.n472 2.6005
R1856 VSS.n480 VSS.n479 2.6005
R1857 VSS.n479 VSS.n478 2.6005
R1858 VSS.n486 VSS.n485 2.6005
R1859 VSS.n485 VSS.n484 2.6005
R1860 VSS.n499 VSS.n498 2.6005
R1861 VSS VSS.n505 2.6005
R1862 VSS.n514 VSS.n513 2.6005
R1863 VSS.n513 VSS.n512 2.6005
R1864 VSS.n521 VSS.n520 2.6005
R1865 VSS.n520 VSS.n519 2.6005
R1866 VSS.n527 VSS.n526 2.6005
R1867 VSS.n526 VSS.n525 2.6005
R1868 VSS.n537 VSS.n536 2.6005
R1869 VSS.n536 VSS.n535 2.6005
R1870 VSS.n532 VSS.n531 2.6005
R1871 VSS.n467 VSS.n466 2.6005
R1872 VSS.n466 VSS.n465 2.6005
R1873 VSS.n75 VSS.n74 2.6005
R1874 VSS.n72 VSS.n69 2.6005
R1875 VSS.n73 VSS.n72 2.6005
R1876 VSS.n236 VSS.n235 2.6005
R1877 VSS.n167 VSS.n166 2.6005
R1878 VSS.n166 VSS.n165 2.6005
R1879 VSS.n170 VSS.n169 2.6005
R1880 VSS.n169 VSS.n168 2.6005
R1881 VSS.n173 VSS.n172 2.6005
R1882 VSS.n172 VSS.n171 2.6005
R1883 VSS.n176 VSS.n175 2.6005
R1884 VSS.n175 VSS.n174 2.6005
R1885 VSS.n179 VSS.n178 2.6005
R1886 VSS.n178 VSS.n177 2.6005
R1887 VSS.n182 VSS.n181 2.6005
R1888 VSS.n181 VSS.n180 2.6005
R1889 VSS.n185 VSS.n184 2.6005
R1890 VSS.n184 VSS.n183 2.6005
R1891 VSS.n188 VSS.n187 2.6005
R1892 VSS.n187 VSS.n186 2.6005
R1893 VSS.n191 VSS.n190 2.6005
R1894 VSS.n190 VSS.n189 2.6005
R1895 VSS.n195 VSS.n194 2.6005
R1896 VSS.n194 VSS.n193 2.6005
R1897 VSS.n198 VSS.n197 2.6005
R1898 VSS.n197 VSS.n196 2.6005
R1899 VSS.n201 VSS.n200 2.6005
R1900 VSS.n200 VSS.n199 2.6005
R1901 VSS.n204 VSS.n203 2.6005
R1902 VSS.n203 VSS.n202 2.6005
R1903 VSS.n207 VSS.n206 2.6005
R1904 VSS.n206 VSS.n205 2.6005
R1905 VSS.n210 VSS.n209 2.6005
R1906 VSS.n209 VSS.n208 2.6005
R1907 VSS.n213 VSS.n212 2.6005
R1908 VSS.n212 VSS.n211 2.6005
R1909 VSS.n216 VSS.n215 2.6005
R1910 VSS.n215 VSS.n214 2.6005
R1911 VSS.n219 VSS.n218 2.6005
R1912 VSS.n218 VSS.n217 2.6005
R1913 VSS.n222 VSS.n221 2.6005
R1914 VSS.n221 VSS.n220 2.6005
R1915 VSS.n225 VSS.n224 2.6005
R1916 VSS.n224 VSS.n223 2.6005
R1917 VSS.n228 VSS.n227 2.6005
R1918 VSS.n227 VSS.n226 2.6005
R1919 VSS.n231 VSS.n230 2.6005
R1920 VSS.n230 VSS.n229 2.6005
R1921 VSS.n234 VSS.n233 2.6005
R1922 VSS.n19 VSS.n18 2.6005
R1923 VSS.n17 VSS.n16 2.6005
R1924 VSS.n164 VSS.n163 2.6005
R1925 VSS.n163 VSS.n162 2.6005
R1926 VSS.n156 VSS.n155 2.6005
R1927 VSS.n154 VSS.n153 2.6005
R1928 VSS.n152 VSS.n151 2.6005
R1929 VSS.n151 VSS.n150 2.6005
R1930 VSS.n149 VSS.n148 2.6005
R1931 VSS.n148 VSS.n147 2.6005
R1932 VSS.n146 VSS.n145 2.6005
R1933 VSS.n145 VSS.n144 2.6005
R1934 VSS.n143 VSS.n142 2.6005
R1935 VSS.n142 VSS.n141 2.6005
R1936 VSS.n140 VSS.n139 2.6005
R1937 VSS.n139 VSS.n138 2.6005
R1938 VSS.n137 VSS.n136 2.6005
R1939 VSS.n136 VSS.n135 2.6005
R1940 VSS.n134 VSS.n133 2.6005
R1941 VSS.n133 VSS.n132 2.6005
R1942 VSS.n131 VSS.n130 2.6005
R1943 VSS.n130 VSS.n129 2.6005
R1944 VSS.n127 VSS.n126 2.6005
R1945 VSS.n126 VSS.n125 2.6005
R1946 VSS.n124 VSS.n123 2.6005
R1947 VSS.n123 VSS.n122 2.6005
R1948 VSS.n121 VSS.n120 2.6005
R1949 VSS.n120 VSS.n119 2.6005
R1950 VSS.n118 VSS.n117 2.6005
R1951 VSS.n117 VSS.n116 2.6005
R1952 VSS.n114 VSS.n113 2.6005
R1953 VSS.n113 VSS.n112 2.6005
R1954 VSS.n111 VSS.n110 2.6005
R1955 VSS.n110 VSS.n109 2.6005
R1956 VSS.n107 VSS.n106 2.6005
R1957 VSS.n106 VSS.n105 2.6005
R1958 VSS.n104 VSS.n103 2.6005
R1959 VSS.n103 VSS.n102 2.6005
R1960 VSS.n101 VSS.n100 2.6005
R1961 VSS.n100 VSS.n99 2.6005
R1962 VSS.n98 VSS.n97 2.6005
R1963 VSS.n97 VSS.n96 2.6005
R1964 VSS.n93 VSS.n92 2.6005
R1965 VSS.n92 VSS.n91 2.6005
R1966 VSS.n2898 VSS.n2897 2.6005
R1967 VSS.n2897 VSS.n2896 2.6005
R1968 VSS.n2901 VSS.n2900 2.6005
R1969 VSS.n2900 VSS.n2899 2.6005
R1970 VSS.n2904 VSS.n2903 2.6005
R1971 VSS.n2903 VSS.n2902 2.6005
R1972 VSS.n2907 VSS.n2906 2.6005
R1973 VSS.n2906 VSS.n2905 2.6005
R1974 VSS.n2910 VSS.n2909 2.6005
R1975 VSS.n2909 VSS.n2908 2.6005
R1976 VSS.n2913 VSS.n2912 2.6005
R1977 VSS.n2912 VSS.n2911 2.6005
R1978 VSS.n2916 VSS.n2915 2.6005
R1979 VSS.n2915 VSS.n2914 2.6005
R1980 VSS.n2919 VSS.n2918 2.6005
R1981 VSS.n2918 VSS.n2917 2.6005
R1982 VSS.n2923 VSS.n2922 2.6005
R1983 VSS.n2922 VSS.n2921 2.6005
R1984 VSS.n2926 VSS.n2925 2.6005
R1985 VSS.n2925 VSS.n2924 2.6005
R1986 VSS.n2929 VSS.n2928 2.6005
R1987 VSS.n2928 VSS.n2927 2.6005
R1988 VSS.n2933 VSS.n2932 2.6005
R1989 VSS.n2932 VSS.n2931 2.6005
R1990 VSS.n2936 VSS.n2935 2.6005
R1991 VSS.n2935 VSS.n2934 2.6005
R1992 VSS.n2939 VSS.n2938 2.6005
R1993 VSS.n2938 VSS.n2937 2.6005
R1994 VSS.n2942 VSS.n2941 2.6005
R1995 VSS.n2941 VSS.n2940 2.6005
R1996 VSS.n2945 VSS.n2944 2.6005
R1997 VSS.n2944 VSS.n2943 2.6005
R1998 VSS.n2947 VSS.n2946 2.6005
R1999 VSS.n2951 VSS.n2950 2.6005
R2000 VSS.n2953 VSS.n2952 2.6005
R2001 VSS.n160 VSS.n159 2.6005
R2002 VSS.n2957 VSS.n2956 2.6005
R2003 VSS.n2956 VSS.n2955 2.6005
R2004 VSS.n2959 VSS.n2958 2.6005
R2005 VSS.n2961 VSS.n2960 2.6005
R2006 VSS.n2895 VSS.n2894 2.6005
R2007 VSS.n2894 VSS.n2893 2.6005
R2008 VSS.n2980 VSS.n2979 2.6005
R2009 VSS.n2979 VSS.n2978 2.6005
R2010 VSS.n2995 VSS.n2994 2.6005
R2011 VSS.n2994 VSS.n2993 2.6005
R2012 VSS.n2999 VSS.n2998 2.6005
R2013 VSS.n2998 VSS.n2997 2.6005
R2014 VSS.n3011 VSS.n3010 2.6005
R2015 VSS.n3010 VSS.n3009 2.6005
R2016 VSS.n3008 VSS.n3007 2.6005
R2017 VSS.n3007 VSS.n3006 2.6005
R2018 VSS.n3005 VSS.n3004 2.6005
R2019 VSS.n3004 VSS.n3003 2.6005
R2020 VSS.n3002 VSS.n3001 2.6005
R2021 VSS.n3001 VSS.n3000 2.6005
R2022 VSS.n3016 VSS.n3015 2.6005
R2023 VSS.n2992 VSS.n2991 2.6005
R2024 VSS.n2991 VSS.n2990 2.6005
R2025 VSS.n2989 VSS.n2988 2.6005
R2026 VSS.n2988 VSS.n2987 2.6005
R2027 VSS.n2986 VSS.n2985 2.6005
R2028 VSS.n2985 VSS.n2984 2.6005
R2029 VSS.n2983 VSS.n2982 2.6005
R2030 VSS.n2982 VSS.n2981 2.6005
R2031 VSS.n2976 VSS.n2975 2.6005
R2032 VSS.n2975 VSS.n2974 2.6005
R2033 VSS.n2973 VSS.n2972 2.6005
R2034 VSS.n2972 VSS.n2971 2.6005
R2035 VSS.n2970 VSS.n2969 2.6005
R2036 VSS.n2969 VSS.n2968 2.6005
R2037 VSS.n2967 VSS.n2966 2.6005
R2038 VSS.n2966 VSS.n2965 2.6005
R2039 VSS.n23 VSS.n22 2.6005
R2040 VSS.n22 VSS.n21 2.6005
R2041 VSS.n26 VSS.n25 2.6005
R2042 VSS.n25 VSS.n24 2.6005
R2043 VSS.n29 VSS.n28 2.6005
R2044 VSS.n28 VSS.n27 2.6005
R2045 VSS.n38 VSS.n37 2.6005
R2046 VSS.n37 VSS.n36 2.6005
R2047 VSS.n35 VSS.n34 2.6005
R2048 VSS.n34 VSS.n33 2.6005
R2049 VSS.n32 VSS.n31 2.6005
R2050 VSS.n31 VSS.n30 2.6005
R2051 VSS.n7 VSS.n6 2.6005
R2052 VSS.n6 VSS.n5 2.6005
R2053 VSS.n9 VSS.n8 2.6005
R2054 VSS.n430 VSS.n427 2.6005
R2055 VSS.n279 VSS.n276 2.6005
R2056 VSS.n266 VSS.n265 2.6005
R2057 VSS.n255 VSS.n252 2.6005
R2058 VSS.n244 VSS.n243 2.6005
R2059 VSS.n243 VSS.n242 2.6005
R2060 VSS.n248 VSS.n247 2.6005
R2061 VSS.n247 VSS.n246 2.6005
R2062 VSS.n256 VSS.n255 2.6005
R2063 VSS.n260 VSS.n259 2.6005
R2064 VSS.n259 VSS.n258 2.6005
R2065 VSS.n266 VSS 2.6005
R2066 VSS.n272 VSS.n271 2.6005
R2067 VSS.n271 VSS.n270 2.6005
R2068 VSS.n280 VSS.n279 2.6005
R2069 VSS.n290 VSS.n289 2.6005
R2070 VSS.n289 VSS.n288 2.6005
R2071 VSS.n431 VSS.n430 2.6005
R2072 VSS.n308 VSS.n307 2.6005
R2073 VSS.n307 VSS.n306 2.6005
R2074 VSS.n240 VSS.n239 2.6005
R2075 VSS.n239 VSS.n238 2.6005
R2076 VSS.n437 VSS.n436 2.6005
R2077 VSS.n436 VSS.n435 2.6005
R2078 VSS.n440 VSS.n439 2.6005
R2079 VSS.n439 VSS.n438 2.6005
R2080 VSS.n443 VSS.n442 2.6005
R2081 VSS.n442 VSS.n441 2.6005
R2082 VSS.n446 VSS.n445 2.6005
R2083 VSS.n445 VSS.n444 2.6005
R2084 VSS.n449 VSS.n448 2.6005
R2085 VSS.n448 VSS.n447 2.6005
R2086 VSS.n452 VSS.n451 2.6005
R2087 VSS.n451 VSS.n450 2.6005
R2088 VSS.n455 VSS.n454 2.6005
R2089 VSS.n454 VSS.n453 2.6005
R2090 VSS.n458 VSS.n457 2.6005
R2091 VSS.n457 VSS.n456 2.6005
R2092 VSS.n3124 VSS.n3123 2.6005
R2093 VSS.n3123 VSS.n3122 2.6005
R2094 VSS.n3121 VSS.n3120 2.6005
R2095 VSS.n3120 VSS.n3119 2.6005
R2096 VSS.n3118 VSS.n3117 2.6005
R2097 VSS.n3117 VSS.n3116 2.6005
R2098 VSS.n3115 VSS.n3114 2.6005
R2099 VSS.n3114 VSS.n3113 2.6005
R2100 VSS.n3112 VSS.n3111 2.6005
R2101 VSS.n3111 VSS.n3110 2.6005
R2102 VSS.n3109 VSS.n3108 2.6005
R2103 VSS.n3108 VSS.n3107 2.6005
R2104 VSS.n3106 VSS.n3105 2.6005
R2105 VSS.n3105 VSS.n3104 2.6005
R2106 VSS.n3103 VSS.n3102 2.6005
R2107 VSS.n3102 VSS.n3101 2.6005
R2108 VSS.n3100 VSS.n3099 2.6005
R2109 VSS.n3099 VSS.n3098 2.6005
R2110 VSS.n3097 VSS.n3096 2.6005
R2111 VSS.n3096 VSS.n3095 2.6005
R2112 VSS.n3093 VSS.n3092 2.6005
R2113 VSS.n3092 VSS.n3091 2.6005
R2114 VSS.n3090 VSS.n3089 2.6005
R2115 VSS.n3089 VSS.n3088 2.6005
R2116 VSS.n3087 VSS.n3086 2.6005
R2117 VSS.n3086 VSS.n3085 2.6005
R2118 VSS.n3084 VSS.n3083 2.6005
R2119 VSS.n3083 VSS.n3082 2.6005
R2120 VSS.n3081 VSS.n3080 2.6005
R2121 VSS.n3080 VSS.n3079 2.6005
R2122 VSS.n3078 VSS.n3077 2.6005
R2123 VSS.n3077 VSS.n3076 2.6005
R2124 VSS.n3075 VSS.n3074 2.6005
R2125 VSS.n3074 VSS.n3073 2.6005
R2126 VSS.n3072 VSS.n3071 2.6005
R2127 VSS.n3071 VSS.n3070 2.6005
R2128 VSS.n3069 VSS.n3068 2.6005
R2129 VSS.n3068 VSS.n3067 2.6005
R2130 VSS.n3065 VSS.n3064 2.6005
R2131 VSS.n3064 VSS.n3063 2.6005
R2132 VSS.n3062 VSS.n3061 2.6005
R2133 VSS.n3061 VSS.n3060 2.6005
R2134 VSS.n3059 VSS.n3058 2.6005
R2135 VSS.n3058 VSS.n3057 2.6005
R2136 VSS.n3056 VSS.n3055 2.6005
R2137 VSS.n3055 VSS.n3054 2.6005
R2138 VSS.n3053 VSS.n3052 2.6005
R2139 VSS.n3052 VSS.n3051 2.6005
R2140 VSS.n3050 VSS.n3049 2.6005
R2141 VSS.n3049 VSS.n3048 2.6005
R2142 VSS.n709 VSS.n708 2.6005
R2143 VSS.n2888 VSS.n2887 2.6005
R2144 VSS.n2890 VSS.n2889 2.6005
R2145 VSS.n2892 VSS.n2891 2.6005
R2146 VSS.n2931 VSS.n2930 2.41686
R2147 VSS.n1700 VSS.n1699 2.29396
R2148 VSS.n1703 VSS.n1702 2.29396
R2149 VSS.n3036 VSS.n3035 2.29396
R2150 VSS.n3033 VSS.n3032 2.29396
R2151 VSS.n3030 VSS.n3029 2.29396
R2152 VSS.n2447 VSS.n2446 2.28399
R2153 VSS.n2450 VSS.n2449 2.28399
R2154 VSS.n2695 VSS.n2694 2.28399
R2155 VSS.n2698 VSS.n2697 2.28399
R2156 VSS.n2814 VSS.n2813 2.28399
R2157 VSS.n2817 VSS.n2816 2.28399
R2158 VSS.n763 VSS.n762 2.25676
R2159 VSS.n545 VSS.n541 2.25575
R2160 VSS.n305 VSS.n304 2.25285
R2161 VSS.n87 VSS.n86 2.2505
R2162 VSS.n405 VSS.n404 2.2505
R2163 VSS.n358 VSS.n357 2.2505
R2164 VSS.n648 VSS.n647 2.2505
R2165 VSS.n660 VSS.n659 2.2505
R2166 VSS.n56 VSS.n55 2.2505
R2167 VSS.n65 VSS.n64 2.2505
R2168 VSS.n423 VSS.n422 2.2505
R2169 VSS.n286 VSS.n285 2.2505
R2170 VSS.n303 VSS.n302 2.24654
R2171 VSS.n2256 VSS.n2255 2.24613
R2172 VSS.n2250 VSS.n2249 2.24465
R2173 VSS.n2246 VSS.n2241 2.24345
R2174 VSS.n2252 VSS.n2240 2.24345
R2175 VSS.n413 VSS.n412 2.12849
R2176 VSS.n585 VSS.n583 2.04928
R2177 VSS.n301 VSS.t373 2.02838
R2178 VSS.n42 VSS.t126 2.02837
R2179 VSS.t313 VSS.t329 2.02605
R2180 VSS.t267 VSS.t313 2.02605
R2181 VSS.n1816 VSS.t5 2.02605
R2182 VSS.n697 VSS.n696 2.0097
R2183 VSS.n570 VSS.n569 2.00969
R2184 VSS.n583 VSS.n568 1.96391
R2185 VSS VSS.n1317 1.9362
R2186 VSS.n3095 VSS.n3094 1.88839
R2187 VSS.n1097 VSS.n1096 1.87053
R2188 VSS.n827 VSS.n826 1.85822
R2189 VSS.n844 VSS.n843 1.85787
R2190 VSS.n2255 VSS.n2254 1.85765
R2191 VSS.n2249 VSS.n2248 1.85765
R2192 VSS.n2416 VSS.n2415 1.83785
R2193 VSS.n1183 VSS.n1182 1.83785
R2194 VSS.n1128 VSS.n1127 1.83757
R2195 VSS.n1005 VSS.n1004 1.83724
R2196 VSS.n727 VSS.n726 1.83716
R2197 VSS.n740 VSS.n739 1.83716
R2198 VSS.n747 VSS.n746 1.83716
R2199 VSS.n1154 VSS.n1153 1.83716
R2200 VSS.n1910 VSS.n1909 1.83716
R2201 VSS.n1916 VSS.n1915 1.83716
R2202 VSS.n1925 VSS.n1924 1.83716
R2203 VSS.n1934 VSS.n1933 1.83716
R2204 VSS.n2392 VSS.n2391 1.83716
R2205 VSS.n2401 VSS.n2400 1.83716
R2206 VSS.n2408 VSS.n2407 1.83716
R2207 VSS.n1002 VSS.n1001 1.83716
R2208 VSS.n869 VSS.n868 1.83716
R2209 VSS.n610 VSS.n609 1.82536
R2210 VSS.n570 VSS.t369 1.82525
R2211 VSS.n697 VSS.t47 1.82525
R2212 VSS.n417 VSS.n416 1.82479
R2213 VSS.n42 VSS.n41 1.80405
R2214 VSS.n301 VSS.n300 1.80404
R2215 VSS.n2962 VSS.n2959 1.8001
R2216 VSS.n2887 VSS.n2886 1.8001
R2217 VSS.n2950 VSS.n2949 1.79951
R2218 VSS.n159 VSS.n158 1.79951
R2219 VSS.n2962 VSS.n2961 1.79951
R2220 VSS.n3017 VSS.n3016 1.79951
R2221 VSS.n3045 VSS.n3041 1.79951
R2222 VSS.n559 VSS.n558 1.79318
R2223 VSS.n255 VSS.n251 1.7505
R2224 VSS.n882 VSS.n881 1.7444
R2225 VSS.n14 VSS.n13 1.70902
R2226 VSS.n1234 VSS.n1233 1.68127
R2227 VSS.n505 VSS.n501 1.65328
R2228 VSS.n72 VSS.n71 1.62245
R2229 VSS.t78 VSS.t350 1.61822
R2230 VSS.n1761 VSS.n1760 1.60209
R2231 VSS.n1158 VSS.n1157 1.60209
R2232 VSS.n1147 VSS.n1146 1.60199
R2233 VSS.n1172 VSS.n1171 1.60199
R2234 VSS.n2143 VSS.n2142 1.60199
R2235 VSS.n1741 VSS.n1738 1.59295
R2236 VSS.n1712 VSS.n1711 1.5924
R2237 VSS.n1717 VSS.n1716 1.5924
R2238 VSS.n1722 VSS.n1721 1.5924
R2239 VSS.n1728 VSS.n1727 1.5924
R2240 VSS.n1741 VSS.n1740 1.5924
R2241 VSS.n1368 VSS.n1367 1.58814
R2242 VSS.n1512 VSS.n1511 1.58814
R2243 VSS.n1503 VSS.n1502 1.58814
R2244 VSS.n1498 VSS.n1497 1.58814
R2245 VSS.n1493 VSS.n1492 1.58814
R2246 VSS.n2827 VSS.n2826 1.58814
R2247 VSS.n1570 VSS.n1569 1.58814
R2248 VSS.n1596 VSS.n1595 1.58814
R2249 VSS.n1363 VSS.n1362 1.58759
R2250 VSS.n1374 VSS.n1373 1.58759
R2251 VSS.n2734 VSS.n2733 1.58759
R2252 VSS.n2459 VSS.n2458 1.58747
R2253 VSS.n2464 VSS.n2463 1.58747
R2254 VSS.n2469 VSS.n2468 1.58747
R2255 VSS.n2475 VSS.n2474 1.58747
R2256 VSS.n2480 VSS.n2479 1.58747
R2257 VSS.n2486 VSS.n2485 1.58747
R2258 VSS.n1563 VSS.n1562 1.58747
R2259 VSS.n1558 VSS.n1557 1.58747
R2260 VSS.n1553 VSS.n1552 1.58747
R2261 VSS.n1548 VSS.n1547 1.58747
R2262 VSS.n1543 VSS.n1542 1.58747
R2263 VSS.n1538 VSS.n1537 1.58747
R2264 VSS.n80 VSS.n77 1.56241
R2265 VSS.n16 VSS.n15 1.55933
R2266 VSS.n233 VSS.n232 1.55922
R2267 VSS.n369 VSS.n367 1.55606
R2268 VSS.n589 VSS.n587 1.5005
R2269 VSS.n430 VSS.n426 1.45883
R2270 VSS.n1268 VSS.n1266 1.45883
R2271 VSS.n3025 VSS.n3023 1.45452
R2272 VSS.n3025 VSS.n3024 1.45452
R2273 VSS.n2258 VSS.n2257 1.43813
R2274 VSS.n680 VSS.n679 1.36161
R2275 VSS.n1691 VSS.n1690 1.33389
R2276 VSS.n1731 VSS.n1730 1.33389
R2277 VSS.n1706 VSS.n1705 1.33375
R2278 VSS.n3027 VSS.n3026 1.33375
R2279 VSS.n1226 VSS.n1225 1.33085
R2280 VSS.n2441 VSS.n2440 1.32883
R2281 VSS.n2702 VSS.n2701 1.32883
R2282 VSS.n2821 VSS.n2820 1.32883
R2283 VSS.n2809 VSS.n2808 1.32869
R2284 VSS.n2690 VSS.n2689 1.32869
R2285 VSS.n2433 VSS.n2432 1.32869
R2286 VSS.n2438 VSS.n2437 1.32869
R2287 VSS.n2453 VSS.n2452 1.32869
R2288 VSS.n1231 VSS.n1230 1.32419
R2289 VSS.n2217 VSS.n2216 1.28654
R2290 VSS.n721 VSS.n720 1.26956
R2291 VSS.n644 VSS.n635 1.26439
R2292 VSS.n666 VSS.n663 1.26439
R2293 VSS.n2114 VSS.n2058 1.22037
R2294 VSS.n2141 VSS.n2134 1.18179
R2295 VSS.n2141 VSS.n2135 1.18179
R2296 VSS.n2141 VSS.n2136 1.18179
R2297 VSS.n2141 VSS.n2137 1.18179
R2298 VSS.n2141 VSS.n2138 1.18179
R2299 VSS.n2141 VSS.n2139 1.18179
R2300 VSS.n2141 VSS.n2140 1.18179
R2301 VSS.n1181 VSS.n1179 1.18179
R2302 VSS.n279 VSS.n275 1.16717
R2303 VSS.n2108 VSS.n2097 1.15537
R2304 VSS.n406 VSS.n405 1.1255
R2305 VSS.n605 VSS.n553 1.09796
R2306 VSS.n606 VSS.n605 1.09475
R2307 VSS.n268 VSS.n266 1.06994
R2308 VSS.n279 VSS.n278 1.06994
R2309 VSS.n2827 VSS.n2825 1.03151
R2310 VSS.t293 VSS.t334 1.01328
R2311 VSS.t283 VSS.t270 1.01328
R2312 VSS.t270 VSS.t308 1.01328
R2313 VSS.n644 VSS.n643 0.972722
R2314 VSS.n666 VSS.n665 0.972722
R2315 VSS.n270 VSS.t84 0.946643
R2316 VSS.n636 VSS.t370 0.944444
R2317 VSS.n421 VSS.n420 0.931406
R2318 VSS.n615 VSS.n614 0.929276
R2319 VSS.n550 VSS.n549 0.928071
R2320 VSS.n353 VSS.n352 0.925894
R2321 VSS.n1708 VSS.n775 0.919029
R2322 VSS.n1726 VSS.n749 0.919029
R2323 VSS.n604 VSS.n598 0.897993
R2324 VSS.n2257 VSS.n2239 0.895896
R2325 VSS.n1587 VSS.t48 0.882454
R2326 VSS.n680 VSS.n676 0.8755
R2327 VSS.t322 VSS.t275 0.852847
R2328 VSS.t275 VSS.t278 0.852847
R2329 VSS.n822 VSS.t12 0.852847
R2330 VSS.n1181 VSS.n1178 0.852847
R2331 VSS.n2701 VSS.n2700 0.849401
R2332 VSS.n2820 VSS.n2819 0.849401
R2333 VSS.n1225 VSS.n1224 0.847764
R2334 VSS.n3026 VSS.n3025 0.845835
R2335 VSS.n608 VSS.n545 0.829906
R2336 VSS.n621 VSS.n618 0.79929
R2337 VSS.n430 VSS.n429 0.778278
R2338 VSS.n1268 VSS.n1264 0.778278
R2339 VSS.n605 VSS.n604 0.768418
R2340 VSS.n691 VSS.n689 0.726531
R2341 VSS.n367 VSS.n323 0.681056
R2342 VSS.n1181 VSS.n1180 0.66722
R2343 VSS.n2142 VSS.n2141 0.66701
R2344 VSS.n858 VSS.n855 0.642239
R2345 VSS.n841 VSS.n838 0.642239
R2346 VSS.n939 VSS.n936 0.642239
R2347 VSS.n1835 VSS.n1834 0.642239
R2348 VSS.n2351 VSS.n2350 0.642239
R2349 VSS.n1843 VSS.n1842 0.642239
R2350 VSS.n1080 VSS.n1079 0.611951
R2351 VSS.n2259 VSS.n2258 0.610998
R2352 VSS.n855 VSS.n852 0.597879
R2353 VSS.n2350 VSS.n2349 0.597879
R2354 VSS.n838 VSS.n835 0.596788
R2355 VSS.n1834 VSS.n1833 0.596788
R2356 VSS.n936 VSS.n933 0.595696
R2357 VSS.n930 VSS.n929 0.587994
R2358 VSS.n2238 VSS.n2235 0.587128
R2359 VSS.n832 VSS.n831 0.586903
R2360 VSS.n1832 VSS.n1831 0.586037
R2361 VSS.n849 VSS.n848 0.585812
R2362 VSS.n2348 VSS.n2347 0.584946
R2363 VSS.n505 VSS.n504 0.583833
R2364 VSS.n831 VSS.n828 0.574288
R2365 VSS.n848 VSS.n845 0.573197
R2366 VSS.n2321 VSS.n2311 0.557842
R2367 VSS.n929 VSS.n926 0.550283
R2368 VSS.n2239 VSS.n2238 0.550283
R2369 VSS.n755 VSS.n754 0.54076
R2370 VSS.n2257 VSS.n2256 0.54028
R2371 VSS.n1373 VSS.n1372 0.508005
R2372 VSS.n1511 VSS.n1510 0.508005
R2373 VSS.n1569 VSS.n1568 0.508005
R2374 VSS.n2485 VSS.n2484 0.507764
R2375 VSS.n1742 VSS.n1741 0.505601
R2376 VSS.n758 VSS.n757 0.502362
R2377 VSS.n2251 VSS.n2250 0.502362
R2378 VSS.n761 VSS.n760 0.497425
R2379 VSS.n2245 VSS.n2244 0.497402
R2380 VSS.n255 VSS.n254 0.486611
R2381 VSS.n308 VSS 0.449668
R2382 VSS.n13 VSS.n12 0.447284
R2383 VSS.n970 VSS.n969 0.435547
R2384 VSS.n1881 VSS.n1880 0.434956
R2385 VSS.n880 VSS.n879 0.427022
R2386 VSS.n2376 VSS.n2373 0.426043
R2387 VSS VSS.n305 0.405813
R2388 VSS.n2949 VSS.n2948 0.402035
R2389 VSS.n158 VSS.n157 0.402035
R2390 VSS.n3044 VSS.n3043 0.402035
R2391 VSS.n2963 VSS.n2962 0.402035
R2392 VSS.n3018 VSS.n3017 0.402035
R2393 VSS.n3046 VSS.n3045 0.402035
R2394 VSS.n1094 VSS.n1092 0.393137
R2395 VSS.n2148 VSS.n2146 0.393137
R2396 VSS.n2550 VSS.n2266 0.391771
R2397 VSS.n2534 VSS.n2293 0.391771
R2398 VSS.n2519 VSS.n2325 0.391771
R2399 VSS.n3021 VSS.n3018 0.390642
R2400 VSS.n1127 VSS.n1126 0.383302
R2401 VSS.n2415 VSS.n2414 0.383166
R2402 VSS.n1182 VSS.n1181 0.383166
R2403 VSS.n2414 VSS.n2413 0.382921
R2404 VSS.n2414 VSS.n2412 0.382921
R2405 VSS.n1932 VSS.n1930 0.382921
R2406 VSS.n1932 VSS.n1931 0.382921
R2407 VSS.n1933 VSS.n1932 0.382921
R2408 VSS.n746 VSS.n745 0.382921
R2409 VSS.n1141 VSS.n1089 0.376519
R2410 VSS.n1160 VSS.n998 0.376518
R2411 VSS.n1929 VSS.n1745 0.37489
R2412 VSS.n1908 VSS.n1751 0.374889
R2413 VSS.n951 VSS.n821 0.372135
R2414 VSS.n718 VSS.n717 0.371392
R2415 VSS.n2211 VSS.n2210 0.371022
R2416 VSS.n715 VSS.n714 0.370645
R2417 VSS.n2214 VSS.n2213 0.370645
R2418 VSS.n1096 VSS.n1095 0.366825
R2419 VSS.n2500 VSS.n2421 0.365076
R2420 VSS.n1192 VSS.n1190 0.358977
R2421 VSS.n1798 VSS.n1796 0.358977
R2422 VSS.n1177 VSS.n967 0.356537
R2423 VSS.n1877 VSS.n1753 0.354994
R2424 VSS.n1920 VSS.n1918 0.347591
R2425 VSS.n820 VSS.n819 0.341179
R2426 VSS.n2204 VSS.n2202 0.340476
R2427 VSS.n863 VSS.n862 0.338978
R2428 VSS.n2335 VSS.n2334 0.338978
R2429 VSS.n240 VSS.n237 0.327038
R2430 VSS.n2489 VSS.n2488 0.326081
R2431 VSS.n1894 VSS.n1752 0.321363
R2432 VSS.n1167 VSS.n980 0.320022
R2433 VSS.n2207 VSS.n2205 0.31827
R2434 VSS.n818 VSS.n817 0.318076
R2435 VSS.n1149 VSS.n1088 0.313628
R2436 VSS.n77 VSS.n75 0.302495
R2437 VSS.n777 VSS.n776 0.3005
R2438 VSS.n2105 VSS.n2098 0.292445
R2439 VSS.n984 VSS.n983 0.291512
R2440 VSS.n1254 VSS.n812 0.290903
R2441 VSS.n1757 VSS.n1756 0.289506
R2442 VSS.n2111 VSS.n2059 0.288772
R2443 VSS.n1244 VSS.n813 0.287963
R2444 VSS.n809 VSS.n780 0.287229
R2445 VSS.n2130 VSS.n1940 0.285098
R2446 VSS.n2120 VSS.n1941 0.285098
R2447 VSS.n789 VSS.n782 0.283556
R2448 VSS.n799 VSS.n781 0.283556
R2449 VSS.n3046 VSS 0.281962
R2450 VSS.n913 VSS.n912 0.2753
R2451 VSS.n2363 VSS.n2352 0.2753
R2452 VSS.n915 VSS.n914 0.2729
R2453 VSS.n940 VSS.n939 0.272046
R2454 VSS.n1844 VSS.n1843 0.27149
R2455 VSS.n912 VSS.n888 0.269479
R2456 VSS.n2364 VSS.n2363 0.269479
R2457 VSS.n1082 VSS.n1081 0.254764
R2458 VSS.n913 VSS.n858 0.250935
R2459 VSS.n915 VSS.n841 0.250935
R2460 VSS.n1836 VSS.n1835 0.250935
R2461 VSS.n2352 VSS.n2351 0.250935
R2462 VSS.n1186 VSS.n1185 0.2505
R2463 VSS.n1873 VSS.n1872 0.2505
R2464 VSS.n2229 VSS.n2228 0.249688
R2465 VSS.n815 VSS.n814 0.24562
R2466 VSS.n730 VSS.n729 0.241152
R2467 VSS.n2303 VSS.n2302 0.241152
R2468 VSS.n2219 VSS.n2218 0.239887
R2469 VSS.n2305 VSS.n2303 0.235283
R2470 VSS.n3066 VSS.n707 0.224214
R2471 VSS.n2330 VSS.n2329 0.217674
R2472 VSS.n1844 VSS.n1837 0.2141
R2473 VSS.n987 VSS.n981 0.213053
R2474 VSS.n997 VSS.n988 0.213053
R2475 VSS.n979 VSS.n968 0.213053
R2476 VSS.n2024 VSS.n2023 0.205045
R2477 VSS.n2228 VSS.n2227 0.201811
R2478 VSS.n2218 VSS.n2217 0.200222
R2479 VSS.n816 VSS.n815 0.199702
R2480 VSS.n115 VSS.n57 0.1985
R2481 VSS.n976 VSS.n975 0.196132
R2482 VSS.n245 VSS.n39 0.193921
R2483 VSS.n434 VSS.n433 0.193087
R2484 VSS.n3126 VSS.n3125 0.190786
R2485 VSS.n722 VSS.n721 0.189956
R2486 VSS.n108 VSS.n90 0.188079
R2487 VSS.n914 VSS.n913 0.1865
R2488 VSS.n54 VSS.n53 0.185092
R2489 VSS.n916 VSS.n915 0.1805
R2490 VSS.n1837 VSS.n1836 0.1805
R2491 VSS.n1132 VSS.n1129 0.174181
R2492 VSS.n2182 VSS.n2179 0.17414
R2493 VSS.n2302 VSS.n2301 0.172819
R2494 VSS.n994 VSS.n993 0.170926
R2495 VSS.n1748 VSS.n1747 0.165596
R2496 VSS.n3020 VSS.n3019 0.164562
R2497 VSS.n2202 VSS.n2201 0.163136
R2498 VSS.n2029 VSS.n2024 0.16275
R2499 VSS.n821 VSS.n820 0.162433
R2500 VSS.n693 VSS.n691 0.161214
R2501 VSS.n618 VSS.n4 0.161214
R2502 VSS.n2957 VSS.n2953 0.160198
R2503 VSS.n736 VSS.n733 0.157329
R2504 VSS.n2402 VSS.n2399 0.15648
R2505 VSS VSS.n693 0.155589
R2506 VSS.n2409 VSS.n2406 0.155512
R2507 VSS.n742 VSS.n725 0.153637
R2508 VSS.n2205 VSS.n2204 0.153513
R2509 VSS.n1083 VSS.n1082 0.152808
R2510 VSS.n819 VSS.n818 0.152738
R2511 VSS.n1137 VSS.n1135 0.152674
R2512 VSS.n293 VSS.n2 0.151571
R2513 VSS.n1240 VSS.n1237 0.150235
R2514 VSS.n1763 VSS.n1762 0.150235
R2515 VSS.n1195 VSS.n1192 0.148852
R2516 VSS.n1198 VSS.n1195 0.148852
R2517 VSS.n1201 VSS.n1198 0.148852
R2518 VSS.n1204 VSS.n1201 0.148852
R2519 VSS.n1207 VSS.n1204 0.148852
R2520 VSS.n1210 VSS.n1207 0.148852
R2521 VSS.n1213 VSS.n1210 0.148852
R2522 VSS.n1217 VSS.n1213 0.148852
R2523 VSS.n1223 VSS.n1217 0.148852
R2524 VSS.n1125 VSS.n1123 0.148852
R2525 VSS.n1123 VSS.n1119 0.148852
R2526 VSS.n1119 VSS.n1116 0.148852
R2527 VSS.n1116 VSS.n1113 0.148852
R2528 VSS.n1113 VSS.n1110 0.148852
R2529 VSS.n1110 VSS.n1107 0.148852
R2530 VSS.n1107 VSS.n1104 0.148852
R2531 VSS.n1104 VSS.n1101 0.148852
R2532 VSS.n1101 VSS.n1098 0.148852
R2533 VSS.n1098 VSS.n1094 0.148852
R2534 VSS.n2150 VSS.n2148 0.148852
R2535 VSS.n2152 VSS.n2150 0.148852
R2536 VSS.n2155 VSS.n2152 0.148852
R2537 VSS.n2158 VSS.n2155 0.148852
R2538 VSS.n2161 VSS.n2158 0.148852
R2539 VSS.n2164 VSS.n2161 0.148852
R2540 VSS.n2167 VSS.n2164 0.148852
R2541 VSS.n2170 VSS.n2167 0.148852
R2542 VSS.n2173 VSS.n2170 0.148852
R2543 VSS.n2176 VSS.n2173 0.148852
R2544 VSS.n1778 VSS.n1776 0.148852
R2545 VSS.n1780 VSS.n1778 0.148852
R2546 VSS.n1782 VSS.n1780 0.148852
R2547 VSS.n1784 VSS.n1782 0.148852
R2548 VSS.n1786 VSS.n1784 0.148852
R2549 VSS.n1788 VSS.n1786 0.148852
R2550 VSS.n1790 VSS.n1788 0.148852
R2551 VSS.n1793 VSS.n1790 0.148852
R2552 VSS.n1796 VSS.n1793 0.148852
R2553 VSS.n950 VSS.n947 0.147239
R2554 VSS.n748 VSS.n744 0.147239
R2555 VSS.n872 VSS.n870 0.147239
R2556 VSS.n907 VSS.n904 0.147239
R2557 VSS.n904 VSS.n901 0.147239
R2558 VSS.n879 VSS.n876 0.147239
R2559 VSS.n897 VSS.n894 0.147239
R2560 VSS.n894 VSS.n824 0.147239
R2561 VSS.n741 VSS.n738 0.147239
R2562 VSS.n1008 VSS.n1006 0.147239
R2563 VSS.n1006 VSS.n1003 0.147239
R2564 VSS.n2358 VSS.n2355 0.147239
R2565 VSS.n1818 VSS.n1815 0.147239
R2566 VSS.n1815 VSS.n1812 0.147239
R2567 VSS.n1854 VSS.n1851 0.147239
R2568 VSS.n2373 VSS.n2370 0.147239
R2569 VSS.n2384 VSS.n2382 0.147239
R2570 VSS.n2389 VSS.n2387 0.147239
R2571 VSS.n1014 VSS.n1011 0.144304
R2572 VSS.n2404 VSS.n2402 0.142348
R2573 VSS.n736 VSS.n735 0.14137
R2574 VSS.n1129 VSS.n1125 0.139951
R2575 VSS.n2179 VSS.n2176 0.139951
R2576 VSS.n2306 VSS.n2305 0.137463
R2577 VSS.n768 VSS.n767 0.136472
R2578 VSS.n580 VSS.n579 0.132286
R2579 VSS.n885 VSS.n884 0.131851
R2580 VSS.n411 VSS.n410 0.131587
R2581 VSS.n957 VSS.n954 0.130588
R2582 VSS.n866 VSS.n865 0.130302
R2583 VSS.n1861 VSS.n1858 0.130084
R2584 VSS.n2338 VSS.n2337 0.129374
R2585 VSS.n2336 VSS.n2335 0.125349
R2586 VSS.n657 VSS.n656 0.12483
R2587 VSS.n864 VSS.n863 0.124421
R2588 VSS.n2305 VSS.n2304 0.123458
R2589 VSS.n886 VSS.n885 0.122817
R2590 VSS.n1011 VSS.n1008 0.122783
R2591 VSS.n2331 VSS.n2330 0.122669
R2592 VSS.n769 VSS.n768 0.122609
R2593 VSS.n420 VSS.n419 0.1225
R2594 VSS.n2367 VSS.n2366 0.121959
R2595 VSS.n771 VSS.n770 0.121915
R2596 VSS.n733 VSS.n732 0.121915
R2597 VSS.n2399 VSS.n2398 0.121915
R2598 VSS.n2406 VSS.n2405 0.121915
R2599 VSS.n723 VSS.n722 0.121893
R2600 VSS.n863 VSS.n860 0.121804
R2601 VSS.n731 VSS.n730 0.121641
R2602 VSS.n923 VSS.n920 0.120826
R2603 VSS.n2378 VSS.n2376 0.120826
R2604 VSS.n1187 VSS.n1184 0.119969
R2605 VSS.n1145 VSS.n1143 0.119969
R2606 VSS.n1148 VSS.n1145 0.119969
R2607 VSS.n1155 VSS.n1152 0.119969
R2608 VSS.n788 VSS.n785 0.119969
R2609 VSS.n795 VSS.n792 0.119969
R2610 VSS.n798 VSS.n795 0.119969
R2611 VSS.n805 VSS.n802 0.119969
R2612 VSS.n808 VSS.n805 0.119969
R2613 VSS.n1259 VSS.n1255 0.119969
R2614 VSS.n1253 VSS.n1250 0.119969
R2615 VSS.n1250 VSS.n1247 0.119969
R2616 VSS.n1243 VSS.n1240 0.119969
R2617 VSS.n1762 VSS.n1759 0.119969
R2618 VSS.n2102 VSS.n2100 0.119969
R2619 VSS.n2104 VSS.n2102 0.119969
R2620 VSS.n2119 VSS.n2116 0.119969
R2621 VSS.n2126 VSS.n2123 0.119969
R2622 VSS.n2129 VSS.n2126 0.119969
R2623 VSS.n2144 VSS.n2133 0.119969
R2624 VSS.n2146 VSS.n2144 0.119969
R2625 VSS.n1917 VSS.n1914 0.119969
R2626 VSS.n1876 VSS.n1874 0.119969
R2627 VSS.n1928 VSS.n1926 0.119969
R2628 VSS.n883 VSS.n880 0.119848
R2629 VSS.n1819 VSS.n1801 0.119848
R2630 VSS.n651 VSS.n650 0.119263
R2631 VSS.n614 VSS.n613 0.119263
R2632 VSS.n1138 VSS.n1134 0.119173
R2633 VSS.n1027 VSS.n1024 0.118921
R2634 VSS.n1030 VSS.n1027 0.118921
R2635 VSS.n1033 VSS.n1030 0.118921
R2636 VSS.n1036 VSS.n1033 0.118921
R2637 VSS.n1039 VSS.n1036 0.118921
R2638 VSS.n1042 VSS.n1039 0.118921
R2639 VSS.n1045 VSS.n1042 0.118921
R2640 VSS.n1048 VSS.n1045 0.118921
R2641 VSS.n1054 VSS.n1051 0.118921
R2642 VSS.n1057 VSS.n1054 0.118921
R2643 VSS.n1060 VSS.n1057 0.118921
R2644 VSS.n1063 VSS.n1060 0.118921
R2645 VSS.n1066 VSS.n1063 0.118921
R2646 VSS.n2272 VSS.n2269 0.118921
R2647 VSS.n2275 VSS.n2272 0.118921
R2648 VSS.n2292 VSS.n2289 0.118921
R2649 VSS.n2289 VSS.n2286 0.118921
R2650 VSS.n2286 VSS.n2283 0.118921
R2651 VSS.n2265 VSS.n2262 0.118921
R2652 VSS.n865 VSS.n864 0.118335
R2653 VSS.n2337 VSS.n2336 0.118335
R2654 VSS.n1134 VSS.n1132 0.116783
R2655 VSS.n2325 VSS.n2324 0.116553
R2656 VSS.n2317 VSS.n2314 0.115403
R2657 VSS.n2186 VSS.n2185 0.115328
R2658 VSS.n1017 VSS.n1014 0.115214
R2659 VSS.n2185 VSS.n2182 0.113776
R2660 VSS.n1926 VSS.n1923 0.113597
R2661 VSS.n545 VSS.n544 0.113103
R2662 VSS.n1688 VSS.n1685 0.113
R2663 VSS.n2824 VSS.n2822 0.113
R2664 VSS.n772 VSS.n771 0.111845
R2665 VSS.n725 VSS.n724 0.111448
R2666 VSS.n2333 VSS.n2332 0.111448
R2667 VSS.n2951 VSS.n2947 0.111156
R2668 VSS.n2953 VSS.n2951 0.111156
R2669 VSS.n2947 VSS.n2945 0.11043
R2670 VSS.n26 VSS.n23 0.110256
R2671 VSS.n29 VSS.n26 0.110256
R2672 VSS.n38 VSS.n35 0.110256
R2673 VSS.n35 VSS.n32 0.110256
R2674 VSS.n32 VSS.n7 0.110256
R2675 VSS.n3011 VSS.n3008 0.110256
R2676 VSS.n3008 VSS.n3005 0.110256
R2677 VSS.n3005 VSS.n3002 0.110256
R2678 VSS.n3002 VSS.n2999 0.110256
R2679 VSS.n2992 VSS.n2989 0.110256
R2680 VSS.n2989 VSS.n2986 0.110256
R2681 VSS.n2986 VSS.n2983 0.110256
R2682 VSS.n2983 VSS.n2980 0.110256
R2683 VSS.n2976 VSS.n2973 0.110256
R2684 VSS.n2973 VSS.n2970 0.110256
R2685 VSS.n2970 VSS.n2967 0.110256
R2686 VSS.n160 VSS.n156 0.110256
R2687 VSS.n156 VSS.n154 0.110256
R2688 VSS.n154 VSS.n152 0.110256
R2689 VSS.n152 VSS.n149 0.110256
R2690 VSS.n149 VSS.n146 0.110256
R2691 VSS.n146 VSS.n143 0.110256
R2692 VSS.n143 VSS.n140 0.110256
R2693 VSS.n140 VSS.n137 0.110256
R2694 VSS.n137 VSS.n134 0.110256
R2695 VSS.n134 VSS.n131 0.110256
R2696 VSS.n131 VSS.n127 0.110256
R2697 VSS.n127 VSS.n124 0.110256
R2698 VSS.n124 VSS.n121 0.110256
R2699 VSS.n121 VSS.n118 0.110256
R2700 VSS.n114 VSS.n111 0.110256
R2701 VSS.n107 VSS.n104 0.110256
R2702 VSS.n104 VSS.n101 0.110256
R2703 VSS.n101 VSS.n98 0.110256
R2704 VSS.n98 VSS.n93 0.110256
R2705 VSS.n2901 VSS.n2898 0.110256
R2706 VSS.n2904 VSS.n2901 0.110256
R2707 VSS.n2907 VSS.n2904 0.110256
R2708 VSS.n2910 VSS.n2907 0.110256
R2709 VSS.n2913 VSS.n2910 0.110256
R2710 VSS.n2916 VSS.n2913 0.110256
R2711 VSS.n2919 VSS.n2916 0.110256
R2712 VSS.n2923 VSS.n2919 0.110256
R2713 VSS.n2926 VSS.n2923 0.110256
R2714 VSS.n2929 VSS.n2926 0.110256
R2715 VSS.n2933 VSS.n2929 0.110256
R2716 VSS.n2936 VSS.n2933 0.110256
R2717 VSS.n2939 VSS.n2936 0.110256
R2718 VSS.n2942 VSS.n2939 0.110256
R2719 VSS.n2945 VSS.n2942 0.110256
R2720 VSS.n19 VSS.n17 0.110256
R2721 VSS.n236 VSS.n234 0.110256
R2722 VSS.n234 VSS.n231 0.110256
R2723 VSS.n231 VSS.n228 0.110256
R2724 VSS.n228 VSS.n225 0.110256
R2725 VSS.n225 VSS.n222 0.110256
R2726 VSS.n222 VSS.n219 0.110256
R2727 VSS.n219 VSS.n216 0.110256
R2728 VSS.n216 VSS.n213 0.110256
R2729 VSS.n213 VSS.n210 0.110256
R2730 VSS.n210 VSS.n207 0.110256
R2731 VSS.n207 VSS.n204 0.110256
R2732 VSS.n204 VSS.n201 0.110256
R2733 VSS.n201 VSS.n198 0.110256
R2734 VSS.n198 VSS.n195 0.110256
R2735 VSS.n195 VSS.n191 0.110256
R2736 VSS.n191 VSS.n188 0.110256
R2737 VSS.n188 VSS.n185 0.110256
R2738 VSS.n185 VSS.n182 0.110256
R2739 VSS.n182 VSS.n179 0.110256
R2740 VSS.n179 VSS.n176 0.110256
R2741 VSS.n176 VSS.n173 0.110256
R2742 VSS.n173 VSS.n170 0.110256
R2743 VSS.n170 VSS.n167 0.110256
R2744 VSS.n167 VSS.n164 0.110256
R2745 VSS.n440 VSS.n437 0.110256
R2746 VSS.n443 VSS.n440 0.110256
R2747 VSS.n446 VSS.n443 0.110256
R2748 VSS.n449 VSS.n446 0.110256
R2749 VSS.n452 VSS.n449 0.110256
R2750 VSS.n455 VSS.n452 0.110256
R2751 VSS.n458 VSS.n455 0.110256
R2752 VSS.n3124 VSS.n3121 0.110256
R2753 VSS.n3121 VSS.n3118 0.110256
R2754 VSS.n3118 VSS.n3115 0.110256
R2755 VSS.n3115 VSS.n3112 0.110256
R2756 VSS.n3112 VSS.n3109 0.110256
R2757 VSS.n3109 VSS.n3106 0.110256
R2758 VSS.n3106 VSS.n3103 0.110256
R2759 VSS.n3103 VSS.n3100 0.110256
R2760 VSS.n3100 VSS.n3097 0.110256
R2761 VSS.n3097 VSS.n3093 0.110256
R2762 VSS.n3093 VSS.n3090 0.110256
R2763 VSS.n3090 VSS.n3087 0.110256
R2764 VSS.n3087 VSS.n3084 0.110256
R2765 VSS.n3084 VSS.n3081 0.110256
R2766 VSS.n3081 VSS.n3078 0.110256
R2767 VSS.n3078 VSS.n3075 0.110256
R2768 VSS.n3075 VSS.n3072 0.110256
R2769 VSS.n3072 VSS.n3069 0.110256
R2770 VSS.n3065 VSS.n3062 0.110256
R2771 VSS.n3062 VSS.n3059 0.110256
R2772 VSS.n3059 VSS.n3056 0.110256
R2773 VSS.n3056 VSS.n3053 0.110256
R2774 VSS.n3053 VSS.n3050 0.110256
R2775 VSS.n2888 VSS.n709 0.110256
R2776 VSS.n2890 VSS.n2888 0.110256
R2777 VSS.n2892 VSS.n2890 0.110256
R2778 VSS.n887 VSS.n886 0.109357
R2779 VSS.n2366 VSS.n2365 0.109357
R2780 VSS.n1505 VSS 0.109087
R2781 VSS.n2390 VSS.n2333 0.108345
R2782 VSS.n2398 VSS.n2397 0.10833
R2783 VSS.n770 VSS.n769 0.10833
R2784 VSS.n732 VSS.n731 0.10833
R2785 VSS.n1072 VSS.n1069 0.108109
R2786 VSS.n2192 VSS.n2189 0.108109
R2787 VSS.n39 VSS.n29 0.108061
R2788 VSS.n2964 VSS.n2957 0.108061
R2789 VSS.n2411 VSS.n2409 0.10713
R2790 VSS.n2293 VSS.n2278 0.107079
R2791 VSS.n60 VSS 0.107055
R2792 VSS.n2111 VSS.n2110 0.106429
R2793 VSS.n3012 VSS.n3011 0.105134
R2794 VSS.n1020 VSS.n1017 0.104711
R2795 VSS.n2320 VSS.n2317 0.104711
R2796 VSS.n870 VSS.n867 0.104196
R2797 VSS.n2385 VSS.n2384 0.104196
R2798 VSS.n1893 VSS.n1891 0.10383
R2799 VSS.n1173 VSS.n1170 0.103507
R2800 VSS.n1190 VSS.n1188 0.103243
R2801 VSS.n963 VSS.n960 0.103217
R2802 VSS.n1867 VSS.n1864 0.103217
R2803 VSS.n2114 VSS.n2113 0.102447
R2804 VSS.n1871 VSS.n1798 0.102447
R2805 VSS.n960 VSS.n957 0.102239
R2806 VSS.n966 VSS.n963 0.102239
R2807 VSS.n1870 VSS.n1867 0.102239
R2808 VSS.n1864 VSS.n1861 0.102239
R2809 VSS.n912 VSS.n911 0.0999444
R2810 VSS.n943 VSS.n940 0.0999444
R2811 VSS.n1808 VSS.n1805 0.0999444
R2812 VSS.n1847 VSS.n1844 0.0999444
R2813 VSS.n2363 VSS.n2362 0.0999444
R2814 VSS.n1689 VSS.n1688 0.0998293
R2815 VSS.n1162 VSS.n1160 0.0992611
R2816 VSS.n724 VSS.n723 0.0990345
R2817 VSS.n2332 VSS.n2331 0.0990345
R2818 VSS.n1000 VSS.n999 0.0986818
R2819 VSS.n1908 VSS.n1907 0.0984646
R2820 VSS.n1923 VSS.n1922 0.0978681
R2821 VSS.n1227 VSS.n1223 0.0974231
R2822 VSS.n1229 VSS.n1227 0.0974231
R2823 VSS.n1235 VSS.n1232 0.0974231
R2824 VSS.n1768 VSS.n1766 0.0974231
R2825 VSS.n1774 VSS.n1771 0.0974231
R2826 VSS.n1776 VSS.n1774 0.0974231
R2827 VSS.n2421 VSS.n2420 0.0973478
R2828 VSS.n1232 VSS.n1229 0.0964341
R2829 VSS.n1771 VSS.n1768 0.0964341
R2830 VSS.n2409 VSS.n2404 0.0963696
R2831 VSS.n802 VSS.n799 0.0952788
R2832 VSS.n2120 VSS.n2119 0.0952788
R2833 VSS.n2222 VSS.n2221 0.0945909
R2834 VSS.n2380 VSS.n2367 0.0945541
R2835 VSS.n1075 VSS.n1072 0.0942929
R2836 VSS.n2195 VSS.n2192 0.0941041
R2837 VSS.n1935 VSS.n1929 0.0928894
R2838 VSS.n2365 VSS.n2364 0.0922143
R2839 VSS.n1141 VSS.n1140 0.0920929
R2840 VSS.n888 VSS.n887 0.0913571
R2841 VSS.n89 VSS.n88 0.0907679
R2842 VSS.n867 VSS.n866 0.0905
R2843 VSS.n775 VSS.n774 0.0905
R2844 VSS.n1255 VSS.n1254 0.0905
R2845 VSS.n2107 VSS.n2105 0.0905
R2846 VSS.n2385 VSS.n2338 0.0905
R2847 VSS.n23 VSS.n20 0.0897683
R2848 VSS.n1871 VSS.n1870 0.0895217
R2849 VSS.n1879 VSS.n1877 0.0889071
R2850 VSS.n1188 VSS.n966 0.0885435
R2851 VSS.n1177 VSS.n1176 0.0881106
R2852 VSS.n1078 VSS.n1075 0.0873421
R2853 VSS.n2198 VSS.n2195 0.0873421
R2854 VSS.n352 VSS.n313 0.0862944
R2855 VSS.n355 VSS.n354 0.0862944
R2856 VSS.n2418 VSS.n2411 0.0856087
R2857 VSS.n2600 VSS.n2596 0.0854057
R2858 VSS.n2596 VSS.n2592 0.0854057
R2859 VSS.n2592 VSS.n2588 0.0854057
R2860 VSS.n2588 VSS.n2584 0.0854057
R2861 VSS.n2584 VSS.n2580 0.0854057
R2862 VSS.n2580 VSS.n2577 0.0854057
R2863 VSS.n2577 VSS.n2574 0.0854057
R2864 VSS.n2574 VSS.n2571 0.0854057
R2865 VSS.n2571 VSS.n2568 0.0854057
R2866 VSS.n2568 VSS.n2565 0.0854057
R2867 VSS.n2565 VSS.n2562 0.0854057
R2868 VSS.n2562 VSS.n2559 0.0854057
R2869 VSS.n2559 VSS.n2556 0.0854057
R2870 VSS.n2556 VSS.n2553 0.0854057
R2871 VSS.n2549 VSS.n2546 0.0854057
R2872 VSS.n2546 VSS.n2543 0.0854057
R2873 VSS.n2543 VSS.n2540 0.0854057
R2874 VSS.n2540 VSS.n2537 0.0854057
R2875 VSS.n2533 VSS.n2530 0.0854057
R2876 VSS.n2530 VSS.n2527 0.0854057
R2877 VSS.n2527 VSS.n2524 0.0854057
R2878 VSS.n2524 VSS.n2521 0.0854057
R2879 VSS.n2518 VSS.n2515 0.0854057
R2880 VSS.n2515 VSS.n2512 0.0854057
R2881 VSS.n2512 VSS.n2509 0.0854057
R2882 VSS.n2509 VSS.n2506 0.0854057
R2883 VSS.n2506 VSS.n2503 0.0854057
R2884 VSS.n2499 VSS.n2496 0.0854057
R2885 VSS.n2496 VSS.n2493 0.0854057
R2886 VSS.n752 VSS.n750 0.0846795
R2887 VSS.n2393 VSS.n2390 0.0846304
R2888 VSS.n2604 VSS.n2600 0.0843639
R2889 VSS.n1140 VSS.n1138 0.0841283
R2890 VSS.n789 VSS.n788 0.0841283
R2891 VSS.n2133 VSS.n2130 0.0841283
R2892 VSS.n1907 VSS.n1905 0.0838349
R2893 VSS.n2375 VSS.n2374 0.0838333
R2894 VSS.n1896 VSS.n1894 0.0837469
R2895 VSS.n1167 VSS.n1166 0.0832732
R2896 VSS.n1939 VSS.n1935 0.0832014
R2897 VSS.n2609 VSS.n2604 0.0830864
R2898 VSS.n1163 VSS.n1162 0.0830384
R2899 VSS.n1904 VSS.n1897 0.0828404
R2900 VSS.n1922 VSS.n1921 0.0828404
R2901 VSS.n1720 VSS.n1718 0.0828171
R2902 VSS.n1375 VSS.n1371 0.0828171
R2903 VSS.n1371 VSS.n1369 0.0828171
R2904 VSS.n1369 VSS.n1366 0.0828171
R2905 VSS.n1366 VSS.n1364 0.0828171
R2906 VSS.n1364 VSS.n1361 0.0828171
R2907 VSS.n1361 VSS.n1359 0.0828171
R2908 VSS.n1359 VSS.n1356 0.0828171
R2909 VSS.n1356 VSS.n1353 0.0828171
R2910 VSS.n1353 VSS.n1350 0.0828171
R2911 VSS.n1350 VSS.n1347 0.0828171
R2912 VSS.n1347 VSS.n1344 0.0828171
R2913 VSS.n1344 VSS.n1341 0.0828171
R2914 VSS.n1341 VSS.n1338 0.0828171
R2915 VSS.n1338 VSS.n1335 0.0828171
R2916 VSS.n1335 VSS.n1332 0.0828171
R2917 VSS.n1332 VSS.n1329 0.0828171
R2918 VSS.n1329 VSS.n1326 0.0828171
R2919 VSS.n1326 VSS.n1323 0.0828171
R2920 VSS.n1323 VSS.n1320 0.0828171
R2921 VSS.n2429 VSS.n2424 0.0828171
R2922 VSS.n2431 VSS.n2429 0.0828171
R2923 VSS.n2434 VSS.n2431 0.0828171
R2924 VSS.n2436 VSS.n2434 0.0828171
R2925 VSS.n2439 VSS.n2436 0.0828171
R2926 VSS.n2442 VSS.n2439 0.0828171
R2927 VSS.n2448 VSS.n2445 0.0828171
R2928 VSS.n2451 VSS.n2448 0.0828171
R2929 VSS.n2454 VSS.n2451 0.0828171
R2930 VSS.n2456 VSS.n2454 0.0828171
R2931 VSS.n2462 VSS.n2460 0.0828171
R2932 VSS.n2465 VSS.n2462 0.0828171
R2933 VSS.n2467 VSS.n2465 0.0828171
R2934 VSS.n2470 VSS.n2467 0.0828171
R2935 VSS.n2472 VSS.n2470 0.0828171
R2936 VSS.n2478 VSS.n2476 0.0828171
R2937 VSS.n2481 VSS.n2478 0.0828171
R2938 VSS.n2483 VSS.n2481 0.0828171
R2939 VSS.n2487 VSS.n2483 0.0828171
R2940 VSS.n1685 VSS.n1682 0.0828171
R2941 VSS.n1682 VSS.n1679 0.0828171
R2942 VSS.n1679 VSS.n1676 0.0828171
R2943 VSS.n1676 VSS.n1673 0.0828171
R2944 VSS.n1673 VSS.n1670 0.0828171
R2945 VSS.n1670 VSS.n1667 0.0828171
R2946 VSS.n1667 VSS.n1664 0.0828171
R2947 VSS.n1664 VSS.n1661 0.0828171
R2948 VSS.n1661 VSS.n1658 0.0828171
R2949 VSS.n1658 VSS.n1655 0.0828171
R2950 VSS.n1655 VSS.n1652 0.0828171
R2951 VSS.n1652 VSS.n1649 0.0828171
R2952 VSS.n1649 VSS.n1646 0.0828171
R2953 VSS.n1646 VSS.n1643 0.0828171
R2954 VSS.n1643 VSS.n1640 0.0828171
R2955 VSS.n1640 VSS.n1637 0.0828171
R2956 VSS.n1637 VSS.n1634 0.0828171
R2957 VSS.n1634 VSS.n1631 0.0828171
R2958 VSS.n1631 VSS.n1628 0.0828171
R2959 VSS.n1628 VSS.n1625 0.0828171
R2960 VSS.n1625 VSS.n1622 0.0828171
R2961 VSS.n1622 VSS.n1619 0.0828171
R2962 VSS.n1619 VSS.n1616 0.0828171
R2963 VSS.n1616 VSS.n1613 0.0828171
R2964 VSS.n1613 VSS.n1610 0.0828171
R2965 VSS.n1610 VSS.n1607 0.0828171
R2966 VSS.n1607 VSS.n1604 0.0828171
R2967 VSS.n1604 VSS.n1601 0.0828171
R2968 VSS.n1601 VSS.n1597 0.0828171
R2969 VSS.n1597 VSS.n1594 0.0828171
R2970 VSS.n1594 VSS.n1592 0.0828171
R2971 VSS.n1592 VSS.n1589 0.0828171
R2972 VSS.n1589 VSS.n1586 0.0828171
R2973 VSS.n1586 VSS.n1583 0.0828171
R2974 VSS.n1583 VSS.n1580 0.0828171
R2975 VSS.n1580 VSS.n1577 0.0828171
R2976 VSS.n1577 VSS.n1574 0.0828171
R2977 VSS.n1574 VSS.n1571 0.0828171
R2978 VSS.n1571 VSS.n1566 0.0828171
R2979 VSS.n1566 VSS.n1564 0.0828171
R2980 VSS.n1564 VSS.n1561 0.0828171
R2981 VSS.n1561 VSS.n1559 0.0828171
R2982 VSS.n1559 VSS.n1556 0.0828171
R2983 VSS.n1556 VSS.n1554 0.0828171
R2984 VSS.n1554 VSS.n1551 0.0828171
R2985 VSS.n1551 VSS.n1549 0.0828171
R2986 VSS.n1549 VSS.n1546 0.0828171
R2987 VSS.n1546 VSS.n1544 0.0828171
R2988 VSS.n1544 VSS.n1541 0.0828171
R2989 VSS.n1541 VSS.n1539 0.0828171
R2990 VSS.n1539 VSS.n1536 0.0828171
R2991 VSS.n1536 VSS.n1534 0.0828171
R2992 VSS.n1534 VSS.n1531 0.0828171
R2993 VSS.n1531 VSS.n1528 0.0828171
R2994 VSS.n1528 VSS.n1525 0.0828171
R2995 VSS.n1525 VSS.n1522 0.0828171
R2996 VSS.n1522 VSS.n1519 0.0828171
R2997 VSS.n1519 VSS.n1516 0.0828171
R2998 VSS.n1516 VSS.n1513 0.0828171
R2999 VSS.n1513 VSS.n1507 0.0828171
R3000 VSS.n1504 VSS.n1501 0.0828171
R3001 VSS.n1501 VSS.n1499 0.0828171
R3002 VSS.n1499 VSS.n1496 0.0828171
R3003 VSS.n1496 VSS.n1494 0.0828171
R3004 VSS.n1494 VSS.n1491 0.0828171
R3005 VSS.n1491 VSS.n1489 0.0828171
R3006 VSS.n1489 VSS.n1487 0.0828171
R3007 VSS.n1487 VSS.n1484 0.0828171
R3008 VSS.n1484 VSS.n1481 0.0828171
R3009 VSS.n1481 VSS.n1478 0.0828171
R3010 VSS.n1478 VSS.n1475 0.0828171
R3011 VSS.n1475 VSS.n1472 0.0828171
R3012 VSS.n1472 VSS.n1469 0.0828171
R3013 VSS.n1469 VSS.n1466 0.0828171
R3014 VSS.n1466 VSS.n1463 0.0828171
R3015 VSS.n1463 VSS.n1460 0.0828171
R3016 VSS.n1460 VSS.n1457 0.0828171
R3017 VSS.n1457 VSS.n1454 0.0828171
R3018 VSS.n1454 VSS.n1451 0.0828171
R3019 VSS.n1451 VSS.n1448 0.0828171
R3020 VSS.n1448 VSS.n1445 0.0828171
R3021 VSS.n1445 VSS.n1442 0.0828171
R3022 VSS.n1442 VSS.n1439 0.0828171
R3023 VSS.n1439 VSS.n1436 0.0828171
R3024 VSS.n1436 VSS.n1433 0.0828171
R3025 VSS.n1433 VSS.n1430 0.0828171
R3026 VSS.n1430 VSS.n1427 0.0828171
R3027 VSS.n1427 VSS.n1424 0.0828171
R3028 VSS.n1424 VSS.n1421 0.0828171
R3029 VSS.n1421 VSS.n1418 0.0828171
R3030 VSS.n1418 VSS.n1415 0.0828171
R3031 VSS.n1415 VSS.n1412 0.0828171
R3032 VSS.n1412 VSS.n1409 0.0828171
R3033 VSS.n1409 VSS.n1406 0.0828171
R3034 VSS.n1406 VSS.n1403 0.0828171
R3035 VSS.n1403 VSS.n1400 0.0828171
R3036 VSS.n1400 VSS.n1397 0.0828171
R3037 VSS.n1397 VSS.n1394 0.0828171
R3038 VSS.n1394 VSS.n1391 0.0828171
R3039 VSS.n1391 VSS.n1388 0.0828171
R3040 VSS.n1388 VSS.n1385 0.0828171
R3041 VSS.n1385 VSS.n1381 0.0828171
R3042 VSS.n1381 VSS.n1378 0.0828171
R3043 VSS.n1694 VSS.n1692 0.0828171
R3044 VSS.n1696 VSS.n1694 0.0828171
R3045 VSS.n1698 VSS.n1696 0.0828171
R3046 VSS.n1701 VSS.n1698 0.0828171
R3047 VSS.n1704 VSS.n1701 0.0828171
R3048 VSS.n1707 VSS.n1704 0.0828171
R3049 VSS.n1713 VSS.n1710 0.0828171
R3050 VSS.n1715 VSS.n1713 0.0828171
R3051 VSS.n1718 VSS.n1715 0.0828171
R3052 VSS.n1723 VSS.n1720 0.0828171
R3053 VSS.n1725 VSS.n1723 0.0828171
R3054 VSS.n1732 VSS.n1729 0.0828171
R3055 VSS.n3039 VSS.n3037 0.0828171
R3056 VSS.n3037 VSS.n3034 0.0828171
R3057 VSS.n3034 VSS.n3031 0.0828171
R3058 VSS.n3031 VSS.n3028 0.0828171
R3059 VSS.n2885 VSS.n2882 0.0828171
R3060 VSS.n2882 VSS.n2879 0.0828171
R3061 VSS.n2879 VSS.n2876 0.0828171
R3062 VSS.n2876 VSS.n2873 0.0828171
R3063 VSS.n2869 VSS.n2866 0.0828171
R3064 VSS.n2866 VSS.n2863 0.0828171
R3065 VSS.n2863 VSS.n2860 0.0828171
R3066 VSS.n2860 VSS.n2857 0.0828171
R3067 VSS.n2850 VSS.n2847 0.0828171
R3068 VSS.n2847 VSS.n2844 0.0828171
R3069 VSS.n2844 VSS.n2841 0.0828171
R3070 VSS.n2837 VSS.n2834 0.0828171
R3071 VSS.n2834 VSS.n2831 0.0828171
R3072 VSS.n2828 VSS.n2824 0.0828171
R3073 VSS.n2822 VSS.n2818 0.0828171
R3074 VSS.n2818 VSS.n2815 0.0828171
R3075 VSS.n2815 VSS.n2812 0.0828171
R3076 VSS.n2812 VSS.n2810 0.0828171
R3077 VSS.n2810 VSS.n2807 0.0828171
R3078 VSS.n2807 VSS.n2804 0.0828171
R3079 VSS.n2804 VSS.n2801 0.0828171
R3080 VSS.n2801 VSS.n2798 0.0828171
R3081 VSS.n2798 VSS.n2795 0.0828171
R3082 VSS.n2795 VSS.n2792 0.0828171
R3083 VSS.n2792 VSS.n2789 0.0828171
R3084 VSS.n2789 VSS.n2786 0.0828171
R3085 VSS.n2786 VSS.n2783 0.0828171
R3086 VSS.n2783 VSS.n2780 0.0828171
R3087 VSS.n2780 VSS.n2777 0.0828171
R3088 VSS.n2777 VSS.n2774 0.0828171
R3089 VSS.n2774 VSS.n2771 0.0828171
R3090 VSS.n2771 VSS.n2768 0.0828171
R3091 VSS.n2768 VSS.n2765 0.0828171
R3092 VSS.n2765 VSS.n2762 0.0828171
R3093 VSS.n2762 VSS.n2759 0.0828171
R3094 VSS.n2759 VSS.n2756 0.0828171
R3095 VSS.n2756 VSS.n2753 0.0828171
R3096 VSS.n2753 VSS.n2750 0.0828171
R3097 VSS.n2750 VSS.n2747 0.0828171
R3098 VSS.n2747 VSS.n2744 0.0828171
R3099 VSS.n2744 VSS.n2741 0.0828171
R3100 VSS.n2741 VSS.n2738 0.0828171
R3101 VSS.n2738 VSS.n2735 0.0828171
R3102 VSS.n2735 VSS.n2732 0.0828171
R3103 VSS.n2732 VSS.n2730 0.0828171
R3104 VSS.n2730 VSS.n2726 0.0828171
R3105 VSS.n2726 VSS.n2723 0.0828171
R3106 VSS.n2723 VSS.n2720 0.0828171
R3107 VSS.n2720 VSS.n2717 0.0828171
R3108 VSS.n2717 VSS.n2714 0.0828171
R3109 VSS.n2714 VSS.n2711 0.0828171
R3110 VSS.n2711 VSS.n2708 0.0828171
R3111 VSS.n2708 VSS.n2703 0.0828171
R3112 VSS.n2703 VSS.n2699 0.0828171
R3113 VSS.n2699 VSS.n2696 0.0828171
R3114 VSS.n2696 VSS.n2693 0.0828171
R3115 VSS.n2693 VSS.n2691 0.0828171
R3116 VSS.n2691 VSS.n2688 0.0828171
R3117 VSS.n2688 VSS.n2685 0.0828171
R3118 VSS.n2685 VSS.n2682 0.0828171
R3119 VSS.n2682 VSS.n2679 0.0828171
R3120 VSS.n2679 VSS.n2676 0.0828171
R3121 VSS.n2676 VSS.n2673 0.0828171
R3122 VSS.n2673 VSS.n2670 0.0828171
R3123 VSS.n2670 VSS.n2666 0.0828171
R3124 VSS.n2666 VSS.n2664 0.0828171
R3125 VSS.n2664 VSS.n2660 0.0828171
R3126 VSS.n2660 VSS.n2657 0.0828171
R3127 VSS.n2657 VSS.n2654 0.0828171
R3128 VSS.n2654 VSS.n2651 0.0828171
R3129 VSS.n2651 VSS.n2648 0.0828171
R3130 VSS.n2648 VSS.n2645 0.0828171
R3131 VSS.n2645 VSS.n2642 0.0828171
R3132 VSS.n2642 VSS.n2638 0.0828171
R3133 VSS.n2638 VSS.n2635 0.0828171
R3134 VSS.n2635 VSS.n2632 0.0828171
R3135 VSS.n2632 VSS.n2629 0.0828171
R3136 VSS.n2629 VSS.n2625 0.0828171
R3137 VSS.n2625 VSS.n2622 0.0828171
R3138 VSS.n2622 VSS.n2618 0.0828171
R3139 VSS.n2618 VSS.n2614 0.0828171
R3140 VSS.n2614 VSS.n2609 0.0828171
R3141 VSS.n2420 VSS.n2418 0.0826739
R3142 VSS.n1176 VSS.n1174 0.082242
R3143 VSS.n2841 VSS.n2838 0.0817195
R3144 VSS.n164 VSS.n160 0.0817195
R3145 VSS.n947 VSS.n944 0.0816957
R3146 VSS.n556 VSS.n555 0.0816607
R3147 VSS.n2024 VSS.n1985 0.0815383
R3148 VSS.n1889 VSS.n1879 0.0814455
R3149 VSS.n1507 VSS.n1505 0.0811707
R3150 VSS.n1914 VSS.n1912 0.0809425
R3151 VSS.n707 VSS.n695 0.0808571
R3152 VSS.n3126 VSS.n4 0.0808571
R3153 VSS.n1851 VSS.n1848 0.0807174
R3154 VSS VSS.n3040 0.0803113
R3155 VSS.n1079 VSS.n1078 0.0802368
R3156 VSS.n1156 VSS.n1155 0.080146
R3157 VSS.n597 VSS.n596 0.079766
R3158 VSS.n2259 VSS.n2198 0.0794474
R3159 VSS.n603 VSS.n602 0.0794283
R3160 VSS.n20 VSS.n19 0.0787927
R3161 VSS.n434 VSS.n7 0.0773293
R3162 VSS.n3125 VSS.n3124 0.0773293
R3163 VSS.n988 VSS.n987 0.0770957
R3164 VSS.n1750 VSS.n1746 0.0770957
R3165 VSS.n2269 VSS.n2266 0.077079
R3166 VSS.n1247 VSS.n1244 0.0769602
R3167 VSS.n2521 VSS.n2519 0.0769151
R3168 VSS.n1938 VSS.n1936 0.076587
R3169 VSS.n3040 VSS.n3039 0.0762317
R3170 VSS VSS.n3126 0.0760357
R3171 VSS.n1809 VSS.n1804 0.0758261
R3172 VSS.n608 VSS.n550 0.0752
R3173 VSS.n901 VSS.n898 0.0748478
R3174 VSS.n2490 VSS.n2487 0.0745854
R3175 VSS.n2278 VSS 0.0739211
R3176 VSS.n2382 VSS.n2380 0.0738696
R3177 VSS VSS.n1048 0.0731316
R3178 VSS.n566 VSS.n565 0.0728214
R3179 VSS.n1260 VSS.n809 0.0721814
R3180 VSS.n1152 VSS.n1150 0.071385
R3181 VSS.n316 VSS.n315 0.0713069
R3182 VSS.n2110 VSS.n2108 0.0705885
R3183 VSS.n707 VSS.n706 0.0704107
R3184 VSS.n56 VSS.n51 0.0704107
R3185 VSS.n59 VSS.n57 0.0704107
R3186 VSS.n237 VSS.n236 0.0700122
R3187 VSS.n3012 VSS.n2892 0.0700122
R3188 VSS.n2476 VSS.n2473 0.0696463
R3189 VSS.n1086 VSS.n1085 0.0687418
R3190 VSS.n2224 VSS.n2223 0.0687418
R3191 VSS.n2457 VSS.n2456 0.0685488
R3192 VSS.n2266 VSS.n2265 0.0676053
R3193 VSS.n979 VSS.n970 0.0675213
R3194 VSS.n1888 VSS.n1881 0.0675213
R3195 VSS.n2321 VSS.n2320 0.0673304
R3196 VSS.n1021 VSS.n1020 0.067297
R3197 VSS.n2967 VSS.n2964 0.0670854
R3198 VSS.n2189 VSS.n2186 0.0670217
R3199 VSS.n996 VSS.n995 0.0666326
R3200 VSS.n1903 VSS.n1902 0.0661354
R3201 VSS.n3047 VSS.n709 0.0656219
R3202 VSS.n2550 VSS.n2549 0.0655943
R3203 VSS.n2500 VSS.n2499 0.0655943
R3204 VSS.n978 VSS.n977 0.0649262
R3205 VSS.n1887 VSS.n1886 0.0644344
R3206 VSS.n991 VSS.n990 0.0640294
R3207 VSS.n1904 VSS.n1903 0.0636492
R3208 VSS.n997 VSS.n996 0.0636492
R3209 VSS.n1087 VSS.n1086 0.0633022
R3210 VSS.n2390 VSS.n2389 0.0631087
R3211 VSS.n979 VSS.n978 0.062959
R3212 VSS.n1888 VSS.n1887 0.062959
R3213 VSS.n2977 VSS.n2976 0.0626951
R3214 VSS.n1750 VSS.n1749 0.0622838
R3215 VSS.n987 VSS.n986 0.0622838
R3216 VSS.n738 VSS.n736 0.0621304
R3217 VSS.n2311 VSS.n2310 0.0618391
R3218 VSS.n1912 VSS.n1750 0.0616757
R3219 VSS.n600 VSS.n599 0.0616009
R3220 VSS.n592 VSS.n591 0.0616009
R3221 VSS.n1150 VSS.n1087 0.0613736
R3222 VSS.n898 VSS.n897 0.0611522
R3223 VSS.n3069 VSS.n3066 0.0605
R3224 VSS.n1855 VSS.n1854 0.0603902
R3225 VSS.n1812 VSS.n1809 0.0601739
R3226 VSS.n1963 VSS.n1960 0.0596608
R3227 VSS.n1966 VSS.n1963 0.0596608
R3228 VSS.n1967 VSS.n1966 0.0596608
R3229 VSS VSS.n1967 0.0596608
R3230 VSS.n1975 VSS.n1972 0.0596608
R3231 VSS.n1978 VSS.n1975 0.0596608
R3232 VSS.n1981 VSS.n1978 0.0596608
R3233 VSS.n2000 VSS.n1997 0.0596608
R3234 VSS.n2003 VSS.n2000 0.0596608
R3235 VSS.n2004 VSS.n2003 0.0596608
R3236 VSS VSS.n2004 0.0596608
R3237 VSS.n2012 VSS.n2009 0.0596608
R3238 VSS.n2015 VSS.n2012 0.0596608
R3239 VSS.n2018 VSS.n2015 0.0596608
R3240 VSS.n2075 VSS.n2072 0.0596608
R3241 VSS.n2078 VSS.n2075 0.0596608
R3242 VSS.n2079 VSS.n2078 0.0596608
R3243 VSS VSS.n2079 0.0596608
R3244 VSS.n2087 VSS.n2084 0.0596608
R3245 VSS.n2090 VSS.n2087 0.0596608
R3246 VSS.n2093 VSS.n2090 0.0596608
R3247 VSS.n2036 VSS.n2033 0.0596608
R3248 VSS.n2039 VSS.n2036 0.0596608
R3249 VSS.n2040 VSS.n2039 0.0596608
R3250 VSS VSS.n2040 0.0596608
R3251 VSS.n2048 VSS.n2045 0.0596608
R3252 VSS.n2051 VSS.n2048 0.0596608
R3253 VSS.n2054 VSS.n2051 0.0596608
R3254 VSS.n628 VSS.n625 0.0596608
R3255 VSS.n631 VSS.n628 0.0596608
R3256 VSS.n951 VSS.n950 0.0594119
R3257 VSS.n2996 VSS.n2992 0.0583049
R3258 VSS.n260 VSS.n257 0.0574719
R3259 VSS.n1003 VSS.n775 0.0572391
R3260 VSS.n1237 VSS.n1235 0.0568736
R3261 VSS.n1766 VSS.n1763 0.0568736
R3262 VSS.n2493 VSS.n2490 0.0559717
R3263 VSS.n118 VSS.n115 0.055378
R3264 VSS.n115 VSS.n114 0.055378
R3265 VSS.n111 VSS.n108 0.055378
R3266 VSS.n108 VSS.n107 0.055378
R3267 VSS.n1848 VSS.n1801 0.0552826
R3268 VSS.n1972 VSS.n1950 0.0552552
R3269 VSS.n2009 VSS.n1988 0.0552552
R3270 VSS.n2084 VSS.n2062 0.0552552
R3271 VSS.n2045 VSS.n1944 0.0552552
R3272 VSS.n919 VSS 0.0549444
R3273 VSS VSS.n1822 0.0543889
R3274 VSS.n944 VSS.n923 0.0543043
R3275 VSS.n272 VSS.n269 0.0536953
R3276 VSS VSS.n633 0.0533671
R3277 VSS.n671 VSS.n668 0.0533671
R3278 VSS.n1024 VSS.n1021 0.0530777
R3279 VSS.n2324 VSS.n2321 0.0530398
R3280 VSS.n263 VSS.n260 0.0521084
R3281 VSS.n273 VSS.n272 0.0521084
R3282 VSS.n2023 VSS.n2022 0.0513891
R3283 VSS.n2379 VSS.n2378 0.0513696
R3284 VSS.n685 VSS.n682 0.0508497
R3285 VSS.n1708 VSS.n1707 0.050439
R3286 VSS.n3066 VSS.n3065 0.0502561
R3287 VSS.n1729 VSS.n1726 0.0498902
R3288 VSS.n2838 VSS.n2837 0.0498902
R3289 VSS.n2108 VSS.n2107 0.0498805
R3290 VSS.n611 VSS.n610 0.0496753
R3291 VSS.n2537 VSS.n2534 0.0486132
R3292 VSS.n249 VSS.n248 0.0483322
R3293 VSS.n3022 VSS.n2885 0.0476951
R3294 VSS.n1902 VSS.n1899 0.0468235
R3295 VSS.n1051 VSS 0.0462895
R3296 VSS.n1837 VSS 0.0460556
R3297 VSS.n3050 VSS.n3047 0.0458659
R3298 VSS.n986 VSS.n985 0.0457432
R3299 VSS VSS.n916 0.0455
R3300 VSS VSS.n2275 0.0455
R3301 VSS.n2402 VSS.n2396 0.0455
R3302 VSS.n1749 VSS.n1748 0.0452568
R3303 VSS.n977 VSS.n972 0.04425
R3304 VSS.n1886 VSS.n1883 0.04425
R3305 VSS.n2069 VSS.n2068 0.0439266
R3306 VSS.n2030 VSS.n2029 0.0439266
R3307 VSS.n622 VSS.n621 0.0439266
R3308 VSS.n2387 VSS.n2385 0.0435435
R3309 VSS.n1244 VSS.n1243 0.0435088
R3310 VSS.n1759 VSS.n1757 0.0427124
R3311 VSS.n993 VSS.n992 0.0426277
R3312 VSS.n415 VSS.n407 0.0425561
R3313 VSS.n2445 VSS.n2443 0.0422073
R3314 VSS.n2443 VSS.n2442 0.0411098
R3315 VSS.n2222 VSS.n2220 0.0407128
R3316 VSS.n1159 VSS.n1156 0.040323
R3317 VSS.n433 VSS.n432 0.0401503
R3318 VSS.n1912 VSS.n1911 0.0395266
R3319 VSS.n742 VSS.n741 0.0386522
R3320 VSS.n437 VSS.n434 0.0385488
R3321 VSS.n2293 VSS.n2292 0.0376053
R3322 VSS.n2534 VSS.n2533 0.0372925
R3323 VSS.n2873 VSS.n2870 0.0367195
R3324 VSS.n2396 VSS.n2393 0.0366957
R3325 VSS.n792 VSS.n789 0.0363407
R3326 VSS.n2130 VSS.n2129 0.0363407
R3327 VSS.n309 VSS.n308 0.0357448
R3328 VSS.n767 VSS.n766 0.0352779
R3329 VSS.n2307 VSS.n2306 0.0352465
R3330 VSS.n1985 VSS.n1982 0.0351154
R3331 VSS.n2022 VSS.n2019 0.0351154
R3332 VSS.n2097 VSS.n2094 0.0351154
R3333 VSS.n2058 VSS.n2055 0.0351154
R3334 VSS.n672 VSS.n671 0.0351154
R3335 VSS.n689 VSS.n686 0.0351154
R3336 VSS.n241 VSS.n240 0.0351154
R3337 VSS.n1260 VSS.n1259 0.0347478
R3338 VSS.n290 VSS.n287 0.034486
R3339 VSS.n303 VSS.n299 0.0334464
R3340 VSS.n1726 VSS.n1725 0.0334268
R3341 VSS.n2857 VSS.n2854 0.0334268
R3342 VSS.n3125 VSS.n458 0.0334268
R3343 VSS.n1149 VSS.n1148 0.0331549
R3344 VSS.n1710 VSS.n1708 0.032878
R3345 VSS.n632 VSS.n631 0.0325979
R3346 VSS.n1184 VSS.n1177 0.0323584
R3347 VSS.n248 VSS.n245 0.0319685
R3348 VSS.n1279 VSS.n1275 0.0318333
R3349 VSS.n1283 VSS.n1279 0.0318333
R3350 VSS.n1294 VSS.n1283 0.0318333
R3351 VSS.n1299 VSS 0.0318333
R3352 VSS.n1303 VSS.n1299 0.0318333
R3353 VSS.n1307 VSS.n1303 0.0318333
R3354 VSS.n1311 VSS.n1307 0.0318333
R3355 VSS.n1877 VSS.n1876 0.0315619
R3356 VSS.n604 VSS.n603 0.0305726
R3357 VSS.n1254 VSS.n1253 0.029969
R3358 VSS.n2105 VSS.n2104 0.029969
R3359 VSS.n1294 VSS.n1293 0.0295
R3360 VSS.n613 VSS.n612 0.0292629
R3361 VSS.n639 VSS.n459 0.0288217
R3362 VSS.n576 VSS.n573 0.028625
R3363 VSS.n703 VSS.n700 0.028625
R3364 VSS.n48 VSS.n45 0.028625
R3365 VSS.n299 VSS.n296 0.028625
R3366 VSS.n1692 VSS.n1689 0.0284878
R3367 VSS.n543 VSS.n542 0.0284
R3368 VSS.n1143 VSS.n1141 0.0283761
R3369 VSS.n612 VSS.n611 0.0283351
R3370 VSS.n245 VSS.n244 0.0281923
R3371 VSS.n2325 VSS.n2296 0.0281316
R3372 VSS.n55 VSS.n54 0.028051
R3373 VSS.n1929 VSS.n1928 0.0275796
R3374 VSS.n544 VSS.n543 0.0275
R3375 VSS.n983 VSS.n982 0.0273085
R3376 VSS.n2220 VSS.n2219 0.0273085
R3377 VSS.n749 VSS.n748 0.026913
R3378 VSS.n762 VSS.n761 0.0265939
R3379 VSS.n406 VSS.n313 0.0265748
R3380 VSS.n2244 VSS.n2243 0.0261799
R3381 VSS.n602 VSS.n601 0.0260963
R3382 VSS.n760 VSS.n759 0.0259717
R3383 VSS.n2246 VSS.n2245 0.0259717
R3384 VSS.n407 VSS.n406 0.0257336
R3385 VSS.n405 VSS.n316 0.0257336
R3386 VSS.n341 VSS.n338 0.0256748
R3387 VSS.n347 VSS.n344 0.0256748
R3388 VSS.n393 VSS.n390 0.0256748
R3389 VSS.n387 VSS.n384 0.0256748
R3390 VSS.n477 VSS.n474 0.0256748
R3391 VSS.n483 VSS.n480 0.0256748
R3392 VSS.n489 VSS.n486 0.0256748
R3393 VSS.n517 VSS.n514 0.0256748
R3394 VSS.n524 VSS.n521 0.0256748
R3395 VSS.n601 VSS.n600 0.0252706
R3396 VSS.n598 VSS.n597 0.0252706
R3397 VSS.n799 VSS.n798 0.0251903
R3398 VSS.n2123 VSS.n2120 0.0251903
R3399 VSS.n1982 VSS.n1981 0.0250455
R3400 VSS.n2019 VSS.n2018 0.0250455
R3401 VSS.n2094 VSS.n2093 0.0250455
R3402 VSS.n2055 VSS.n2054 0.0250455
R3403 VSS.n400 VSS.n397 0.0250455
R3404 VSS.n686 VSS.n685 0.0250455
R3405 VSS.n244 VSS.n241 0.0250455
R3406 VSS.n2307 VSS.n2299 0.0247308
R3407 VSS.n491 VSS.n490 0.0247308
R3408 VSS.n412 VSS.n411 0.024574
R3409 VSS.n1378 VSS.n1375 0.0240976
R3410 VSS.n2831 VSS.n2828 0.0240976
R3411 VSS.n2421 VSS.n2328 0.0239783
R3412 VSS.n1317 VSS.n1312 0.0235
R3413 VSS.n2256 VSS.n2252 0.0234789
R3414 VSS.n954 VSS.n951 0.0232368
R3415 VSS.n756 VSS.n755 0.0230525
R3416 VSS.n2380 VSS.n2379 0.023
R3417 VSS.n1858 VSS.n1855 0.0227632
R3418 VSS.n714 VSS.n713 0.0220702
R3419 VSS.n1911 VSS.n1908 0.0220044
R3420 VSS.n73 VSS.n68 0.0217195
R3421 VSS.n563 VSS.n560 0.0213929
R3422 VSS.n717 VSS.n716 0.0213264
R3423 VSS.n2215 VSS.n2214 0.0213264
R3424 VSS.n2212 VSS.n2211 0.0213264
R3425 VSS.n766 VSS.n765 0.0212692
R3426 VSS.n1160 VSS.n1159 0.021208
R3427 VSS.n1085 VSS.n1000 0.0209545
R3428 VSS.n2224 VSS.n2222 0.0209545
R3429 VSS.n757 VSS.n756 0.0208774
R3430 VSS.n410 VSS.n409 0.0207174
R3431 VSS.n552 VSS.n551 0.0207174
R3432 VSS.n364 VSS 0.0206399
R3433 VSS.n1170 VSS.n1167 0.0204115
R3434 VSS.n590 VSS.n589 0.0203165
R3435 VSS.n2553 VSS.n2550 0.0203113
R3436 VSS.n2503 VSS.n2500 0.0203113
R3437 VSS.n1081 VSS.n1080 0.0200985
R3438 VSS.n884 VSS.n883 0.0200652
R3439 VSS.n409 VSS.n408 0.0200652
R3440 VSS.n553 VSS.n552 0.0200652
R3441 VSS.n2258 VSS.n2229 0.0200447
R3442 VSS.n2252 VSS.n2251 0.0200283
R3443 VSS.n652 VSS.n651 0.0199845
R3444 VSS.n720 VSS.n719 0.0198388
R3445 VSS.n2217 VSS.n2207 0.0198346
R3446 VSS.n587 VSS.n566 0.0197857
R3447 VSS.n1894 VSS.n1893 0.019615
R3448 VSS.n817 VSS.n816 0.0196091
R3449 VSS.n845 VSS.n844 0.0191251
R3450 VSS.n828 VSS.n827 0.0191251
R3451 VSS.n2209 VSS.n2208 0.019095
R3452 VSS.n884 VSS.n872 0.019087
R3453 VSS.n649 VSS.n648 0.0190567
R3454 VSS.n581 VSS.n580 0.0189821
R3455 VSS.n63 VSS.n62 0.0188673
R3456 VSS.n721 VSS.n711 0.0188391
R3457 VSS.n1833 VSS.n1832 0.0186836
R3458 VSS.n2349 VSS.n2348 0.0186836
R3459 VSS.n2235 VSS.n2234 0.0186836
R3460 VSS.n596 VSS.n595 0.0186651
R3461 VSS.n284 VSS.n283 0.0185
R3462 VSS.n609 VSS.n608 0.0185
R3463 VSS.n2210 VSS.n2209 0.0184602
R3464 VSS.n351 VSS.n350 0.0184371
R3465 VSS.n659 VSS.n658 0.0181289
R3466 VSS.n744 VSS.n742 0.0181087
R3467 VSS.n2301 VSS.n2300 0.0181073
R3468 VSS.n719 VSS.n718 0.0180867
R3469 VSS.n2116 VSS.n2114 0.0180221
R3470 VSS.n1874 VSS.n1871 0.0180221
R3471 VSS.n594 VSS.n593 0.0178394
R3472 VSS.n852 VSS.n849 0.0178182
R3473 VSS.n835 VSS.n832 0.0178182
R3474 VSS.n933 VSS.n930 0.0178182
R3475 VSS.n332 VSS.n331 0.0178077
R3476 VSS.n378 VSS.n377 0.0178077
R3477 VSS.n468 VSS.n467 0.0178077
R3478 VSS.n534 VSS.n533 0.0178077
R3479 VSS.n285 VSS.n282 0.0175
R3480 VSS.n541 VSS.n527 0.017493
R3481 VSS.n560 VSS.n556 0.017375
R3482 VSS.n565 VSS.n564 0.017375
R3483 VSS.n1188 VSS.n1187 0.0172257
R3484 VSS.n867 VSS.n749 0.0171304
R3485 VSS.n82 VSS.n81 0.0170306
R3486 VSS.n312 VSS.n311 0.0165
R3487 VSS.n1150 VSS.n1149 0.0164292
R3488 VSS.n656 VSS.n655 0.0162732
R3489 VSS.n1960 VSS.n1957 0.0162343
R3490 VSS.n1997 VSS.n1994 0.0162343
R3491 VSS.n2072 VSS.n2069 0.0162343
R3492 VSS.n2033 VSS.n2030 0.0162343
R3493 VSS.n625 VSS.n622 0.0162343
R3494 VSS.n1819 VSS.n1818 0.0161522
R3495 VSS.n86 VSS.n85 0.0161122
R3496 VSS.n2854 VSS.n2850 0.0158659
R3497 VSS.n2213 VSS.n2212 0.015852
R3498 VSS.n548 VSS.n547 0.0158
R3499 VSS.n404 VSS 0.0156049
R3500 VSS.n422 VSS.n312 0.0155
R3501 VSS.n2250 VSS.n2246 0.015398
R3502 VSS.n920 VSS.n824 0.0151739
R3503 VSS.n716 VSS.n715 0.0151082
R3504 VSS.n2216 VSS.n2215 0.0151082
R3505 VSS.n1923 VSS.n1917 0.0148363
R3506 VSS.n2310 VSS.n2309 0.0148234
R3507 VSS.n763 VSS.n752 0.0148073
R3508 VSS.n2460 VSS.n2457 0.0147683
R3509 VSS.n713 VSS.n712 0.0147345
R3510 VSS.n511 VSS.n460 0.0146608
R3511 VSS.n759 VSS.n758 0.014549
R3512 VSS.n65 VSS.n60 0.0144024
R3513 VSS.n586 VSS 0.0141607
R3514 VSS.n87 VSS.n80 0.0141607
R3515 VSS.n415 VSS.n414 0.0141607
R3516 VSS.n809 VSS.n808 0.0140398
R3517 VSS.n2113 VSS.n2111 0.0140398
R3518 VSS.n356 VSS.n355 0.0139579
R3519 VSS.n1271 VSS.n1270 0.0138333
R3520 VSS.n2473 VSS.n2472 0.0136707
R3521 VSS.n1275 VSS.n1271 0.0135
R3522 VSS.n655 VSS.n654 0.0134897
R3523 VSS.n647 VSS.n646 0.0130874
R3524 VSS.n414 VSS.n413 0.0126543
R3525 VSS.n2870 VSS.n2869 0.0125732
R3526 VSS.n285 VSS.n284 0.0125
R3527 VSS.n661 VSS.n660 0.012458
R3528 VSS.n85 VSS.n84 0.0124388
R3529 VSS.n994 VSS.n989 0.0124337
R3530 VSS.n1905 VSS.n1904 0.0124337
R3531 VSS.n1084 VSS.n1083 0.0123681
R3532 VSS.n976 VSS.n973 0.0123033
R3533 VSS.n1889 VSS.n1888 0.0123033
R3534 VSS.n357 VSS.n356 0.0122757
R3535 VSS.n547 VSS.n546 0.0122
R3536 VSS.n992 VSS.n991 0.0119894
R3537 VSS.n1163 VSS.n997 0.0119365
R3538 VSS.n1901 VSS.n1900 0.0119365
R3539 VSS.n2228 VSS.n2225 0.0118736
R3540 VSS.n256 VSS.n249 0.0118287
R3541 VSS.n1174 VSS.n979 0.0118115
R3542 VSS.n1885 VSS.n1884 0.0118115
R3543 VSS.n57 VSS.n56 0.01175
R3544 VSS.n53 VSS.n52 0.0115204
R3545 VSS.n975 VSS.n974 0.0113172
R3546 VSS.n1899 VSS.n1898 0.0113172
R3547 VSS.n286 VSS.n281 0.0111993
R3548 VSS.n579 VSS.n576 0.0109464
R3549 VSS.n88 VSS.n87 0.0109464
R3550 VSS.n706 VSS.n703 0.0109464
R3551 VSS.n658 VSS.n657 0.0107062
R3552 VSS.n404 VSS.n403 0.0105699
R3553 VSS.n674 VSS.n673 0.0105699
R3554 VSS.n433 VSS.n290 0.0105699
R3555 VSS.n416 VSS.n415 0.0101429
R3556 VSS.n51 VSS.n48 0.0101429
R3557 VSS.n296 VSS.n293 0.0101429
R3558 VSS.n90 VSS.n73 0.0100122
R3559 VSS.n1891 VSS.n1889 0.00997368
R3560 VSS.n432 VSS.n431 0.00994056
R3561 VSS.n424 VSS.n423 0.00994056
R3562 VSS.n650 VSS.n649 0.00977835
R3563 VSS.n659 VSS.n652 0.00977835
R3564 VSS.n64 VSS.n63 0.00968367
R3565 VSS.n315 VSS.n314 0.00965814
R3566 VSS.n607 VSS.n606 0.00958707
R3567 VSS.n1174 VSS.n1173 0.0095
R3568 VSS.n673 VSS.n672 0.00931119
R3569 VSS.n682 VSS.n681 0.00931119
R3570 VSS.n972 VSS.n971 0.00925
R3571 VSS.n1883 VSS.n1882 0.00925
R3572 VSS.n1166 VSS.n1163 0.00902632
R3573 VSS.n2519 VSS.n2518 0.00899057
R3574 VSS.n1312 VSS.n1311 0.00883333
R3575 VSS.n646 VSS.n645 0.00868182
R3576 VSS.n667 VSS.n661 0.00868182
R3577 VSS.n541 VSS.n540 0.00868182
R3578 VSS.n310 VSS.n309 0.00868182
R3579 VSS.n1905 VSS.n1896 0.00855263
R3580 VSS.n335 VSS.n332 0.00836713
R3581 VSS.n381 VSS.n378 0.00836713
R3582 VSS.n471 VSS.n468 0.00836713
R3583 VSS.n537 VSS.n534 0.00836713
R3584 VSS.n908 VSS.n907 0.00832609
R3585 VSS.n280 VSS.n273 0.00805245
R3586 VSS.n287 VSS.n286 0.00805245
R3587 VSS.n595 VSS.n594 0.00793119
R3588 VSS.n593 VSS.n592 0.00793119
R3589 VSS.n83 VSS.n82 0.00784694
R3590 VSS.n68 VSS.n65 0.00781707
R3591 VSS.n564 VSS.n563 0.00773214
R3592 VSS.n2262 VSS.n2259 0.00760526
R3593 VSS.n418 VSS.n417 0.00757142
R3594 VSS.n269 VSS 0.00742308
R3595 VSS.n281 VSS.n280 0.00742308
R3596 VSS.n608 VSS.n607 0.00735714
R3597 VSS.n2359 VSS.n2358 0.00734783
R3598 VSS.n3040 VSS.n1732 0.00708537
R3599 VSS.n2999 VSS.n2996 0.00708537
R3600 VSS.n1886 VSS.n1885 0.00689344
R3601 VSS.n1079 VSS.n1066 0.00681579
R3602 VSS.n647 VSS.n632 0.00679371
R3603 VSS.n645 VSS.n633 0.00679371
R3604 VSS.n660 VSS.n459 0.00679371
R3605 VSS.n668 VSS.n667 0.00679371
R3606 VSS.n419 VSS.n418 0.0065
R3607 VSS.n3022 VSS.n3021 0.0064434
R3608 VSS.n2870 VSS.n1735 0.0064434
R3609 VSS.n2854 VSS.n2853 0.0064434
R3610 VSS.n2838 VSS.n1742 0.0064434
R3611 VSS.n977 VSS.n976 0.00640164
R3612 VSS.n591 VSS.n590 0.00627982
R3613 VSS.n305 VSS.n303 0.00622751
R3614 VSS.n681 VSS.n674 0.00616434
R3615 VSS.n581 VSS 0.006125
R3616 VSS.n695 VSS 0.006125
R3617 VSS.n1902 VSS.n1901 0.00596961
R3618 VSS.n496 VSS.n460 0.00584965
R3619 VSS.n358 VSS.n351 0.00553496
R3620 VSS.n365 VSS.n364 0.00553496
R3621 VSS.n431 VSS.n424 0.00553496
R3622 VSS.n1270 VSS.n1269 0.0055
R3623 VSS.n995 VSS.n994 0.00547238
R3624 VSS.n774 VSS.n772 0.0053913
R3625 VSS.n587 VSS.n586 0.00532143
R3626 VSS VSS.n59 0.00532143
R3627 VSS VSS.n2 0.00532143
R3628 VSS.n764 VSS.n763 0.00511538
R3629 VSS.n2309 VSS.n2308 0.00511538
R3630 VSS.n86 VSS.n83 0.00509184
R3631 VSS VSS.n1950 0.00490559
R3632 VSS VSS.n1988 0.00490559
R3633 VSS VSS.n2062 0.00490559
R3634 VSS VSS.n1944 0.00490559
R3635 VSS.n338 VSS.n335 0.00490559
R3636 VSS.n344 VSS.n341 0.00490559
R3637 VSS.n350 VSS.n347 0.00490559
R3638 VSS.n403 VSS.n400 0.00490559
R3639 VSS.n396 VSS.n393 0.00490559
R3640 VSS.n390 VSS.n387 0.00490559
R3641 VSS.n384 VSS.n381 0.00490559
R3642 VSS VSS.n639 0.00490559
R3643 VSS.n474 VSS.n471 0.00490559
R3644 VSS.n480 VSS.n477 0.00490559
R3645 VSS.n486 VSS.n483 0.00490559
R3646 VSS.n490 VSS.n489 0.00490559
R3647 VSS.n514 VSS.n511 0.00490559
R3648 VSS.n527 VSS.n524 0.00490559
R3649 VSS.n540 VSS.n537 0.00490559
R3650 VSS VSS.n264 0.00490559
R3651 VSS.n90 VSS.n89 0.00489024
R3652 VSS.n357 VSS.n353 0.00456316
R3653 VSS.n654 VSS.n653 0.00446899
R3654 VSS.n497 VSS.n496 0.00427622
R3655 VSS.n521 VSS.n518 0.00427622
R3656 VSS.n985 VSS.n984 0.00414865
R3657 VSS.n422 VSS.n421 0.00396834
R3658 VSS.n2308 VSS.n2307 0.00396154
R3659 VSS.n1923 VSS.n1920 0.00371429
R3660 VSS.n257 VSS.n256 0.00364685
R3661 VSS.n264 VSS.n263 0.00364685
R3662 VSS.n3018 VSS.n3012 0.0034717
R3663 VSS.n2996 VSS.n2995 0.0034717
R3664 VSS.n2977 VSS.n2895 0.0034717
R3665 VSS.n2964 VSS.n2963 0.0034717
R3666 VSS.n3047 VSS.n3046 0.0034717
R3667 VSS.n1269 VSS.n1261 0.00316667
R3668 VSS.n549 VSS.n548 0.00313878
R3669 VSS.n1085 VSS.n1084 0.00297253
R3670 VSS.n2225 VSS.n2224 0.00297253
R3671 VSS.n589 VSS.n588 0.00287973
R3672 VSS.n648 VSS.n615 0.00283689
R3673 VSS.n1293 VSS 0.00283333
R3674 VSS.n766 VSS.n764 0.00280769
R3675 VSS.n359 VSS.n358 0.0027028
R3676 VSS.n359 VSS.n324 0.0027028
R3677 VSS.n365 VSS.n324 0.0027028
R3678 VSS VSS.n321 0.0027028
R3679 VSS VSS.n321 0.0027028
R3680 VSS VSS.n506 0.0027028
R3681 VSS.n506 VSS 0.0027028
R3682 VSS.n39 VSS.n38 0.00269512
R3683 VSS.n2980 VSS.n2977 0.00269512
R3684 VSS VSS.n497 0.00238811
R3685 VSS.n2243 VSS.n2242 0.00224148
R3686 VSS.n1809 VSS.n1808 0.00216667
R3687 VSS.n1822 VSS.n1819 0.00216667
R3688 VSS.n1848 VSS.n1847 0.00216667
R3689 VSS.n2362 VSS.n2359 0.00216667
R3690 VSS.n1505 VSS.n1504 0.00214634
R3691 VSS.n2396 VSS.n2395 0.00189535
R3692 VSS.n2418 VSS.n2417 0.00189535
R3693 VSS.n64 VSS.n61 0.00185388
R3694 VSS.n762 VSS.n753 0.0018278
R3695 VSS.n423 VSS.n310 0.00175874
R3696 VSS.n911 VSS.n908 0.00161111
R3697 VSS.n898 VSS.n891 0.00161111
R3698 VSS.n920 VSS.n919 0.00161111
R3699 VSS.n944 VSS.n943 0.00161111
R3700 VSS.n3028 VSS.n3022 0.00159756
R3701 VSS VSS.n491 0.00144406
R3702 VSS.n2186 VSS.n1939 0.00127586
R3703 VSS.n397 VSS.n396 0.00112937
R3704 VSS.n518 VSS.n517 0.00112937
R3705 VCO_C_0.INV_2_3.IN.n70 VCO_C_0.INV_2_3.IN.t51 23.6945
R3706 VCO_C_0.INV_2_3.IN.t35 VCO_C_0.INV_2_3.IN.n71 23.6945
R3707 VCO_C_0.INV_2_3.IN.n71 VCO_C_0.INV_2_3.IN.n70 18.8035
R3708 VCO_C_0.INV_2_3.IN.n68 VCO_C_0.INV_2_3.IN.n66 15.8172
R3709 VCO_C_0.INV_2_3.IN.n68 VCO_C_0.INV_2_3.IN.n67 15.8172
R3710 VCO_C_0.INV_2_3.IN.n67 VCO_C_0.INV_2_3.IN.n63 15.8172
R3711 VCO_C_0.INV_2_3.IN.n66 VCO_C_0.INV_2_3.IN.t50 14.8925
R3712 VCO_C_0.INV_2_3.IN.t38 VCO_C_0.INV_2_3.IN.n68 14.8925
R3713 VCO_C_0.INV_2_3.IN.n67 VCO_C_0.INV_2_3.IN.t32 14.8925
R3714 VCO_C_0.INV_2_3.IN.n72 VCO_C_0.INV_2_3.IN.n64 12.2457
R3715 VCO_C_0.INV_2_3.IN.n69 VCO_C_0.INV_2_3.IN.n64 12.2457
R3716 VCO_C_0.INV_2_3.IN.n69 VCO_C_0.INV_2_3.IN.n65 12.2457
R3717 VCO_C_0.INV_2_3.IN.n73 VCO_C_0.INV_2_3.IN.t43 11.6285
R3718 VCO_C_0.INV_2_3.IN.n15 VCO_C_0.INV_2_3.IN.t57 9.07401
R3719 VCO_C_0.INV_2_3.IN.n19 VCO_C_0.INV_2_3.IN.t56 8.94931
R3720 VCO_C_0.INV_2_3.IN.n13 VCO_C_0.INV_2_3.IN.t53 8.91612
R3721 VCO_C_0.INV_2_3.IN.n12 VCO_C_0.INV_2_3.IN.t45 8.91612
R3722 VCO_C_0.INV_2_3.IN.n9 VCO_C_0.INV_2_3.IN.t30 8.91612
R3723 VCO_C_0.INV_2_3.IN.n65 VCO_C_0.INV_2_3.IN.t51 8.9065
R3724 VCO_C_0.INV_2_3.IN.t55 VCO_C_0.INV_2_3.IN.n69 8.9065
R3725 VCO_C_0.INV_2_3.IN.t31 VCO_C_0.INV_2_3.IN.n64 8.9065
R3726 VCO_C_0.INV_2_3.IN.n72 VCO_C_0.INV_2_3.IN.t35 8.9065
R3727 VCO_C_0.INV_2_3.IN.n7 VCO_C_0.INV_2_3.IN.t33 8.88203
R3728 VCO_C_0.INV_2_3.IN.n17 VCO_C_0.INV_2_3.IN.t42 8.78079
R3729 VCO_C_0.INV_2_3.IN.n20 VCO_C_0.INV_2_3.IN.t39 8.78079
R3730 VCO_C_0.INV_2_3.IN.n16 VCO_C_0.INV_2_3.IN.t47 8.76459
R3731 VCO_C_0.INV_2_3.IN.n15 VCO_C_0.INV_2_3.IN.t44 8.76459
R3732 VCO_C_0.INV_2_3.IN.n51 VCO_C_0.INV_2_3.IN.n49 8.71932
R3733 VCO_C_0.INV_2_3.IN.n8 VCO_C_0.INV_2_3.IN.t34 8.71352
R3734 VCO_C_0.INV_2_3.IN.n11 VCO_C_0.INV_2_3.IN.t37 8.71352
R3735 VCO_C_0.INV_2_3.IN.n68 VCO_C_0.INV_2_3.IN.t41 8.6145
R3736 VCO_C_0.INV_2_3.IN.n66 VCO_C_0.INV_2_3.IN.t54 8.6145
R3737 VCO_C_0.INV_2_3.IN.n67 VCO_C_0.INV_2_3.IN.t36 8.6145
R3738 VCO_C_0.INV_2_3.IN.n63 VCO_C_0.INV_2_3.IN.t48 8.59715
R3739 VCO_C_0.INV_2_3.IN.n14 VCO_C_0.INV_2_3.IN.t40 8.50287
R3740 VCO_C_0.INV_2_3.IN.n0 VCO_C_0.INV_2_3.IN.t52 8.38543
R3741 VCO_C_0.INV_2_3.IN.t50 VCO_C_0.INV_2_3.IN.n65 8.3225
R3742 VCO_C_0.INV_2_3.IN.n69 VCO_C_0.INV_2_3.IN.t38 8.3225
R3743 VCO_C_0.INV_2_3.IN.t32 VCO_C_0.INV_2_3.IN.n64 8.3225
R3744 VCO_C_0.INV_2_3.IN.t43 VCO_C_0.INV_2_3.IN.n72 8.3225
R3745 VCO_C_0.INV_2_3.IN.n41 VCO_C_0.INV_2_3.IN.t10 8.51681
R3746 VCO_C_0.INV_2_3.IN.n18 VCO_C_0.INV_2_3.IN.t49 8.30117
R3747 VCO_C_0.INV_2_3.IN.n3 VCO_C_0.INV_2_3.IN.n2 8.23463
R3748 VCO_C_0.INV_2_3.IN.n7 VCO_C_0.INV_2_3.IN.t46 7.39905
R3749 VCO_C_0.INV_2_3.IN.n81 VCO_C_0.INV_2_3.IN.n80 6.43594
R3750 VCO_C_0.INV_2_3.IN.n60 VCO_C_0.INV_2_3.IN.n59 6.42178
R3751 VCO_C_0.INV_2_3.IN.n1 VCO_C_0.INV_2_3.IN.n82 6.3977
R3752 VCO_C_0.INV_2_3.IN.n6 VCO_C_0.INV_2_3.IN.n5 6.02773
R3753 VCO_C_0.INV_2_3.IN.n57 VCO_C_0.INV_2_3.IN.t21 5.83006
R3754 VCO_C_0.INV_2_3.IN.n45 VCO_C_0.INV_2_3.IN.n32 5.43818
R3755 VCO_C_0.INV_2_3.IN.n60 VCO_C_0.INV_2_3.IN.n54 5.23259
R3756 VCO_C_0.INV_2_3.IN.n43 VCO_C_0.INV_2_3.IN.n42 4.89653
R3757 VCO_C_0.INV_2_3.IN.n21 VCO_C_0.INV_2_3.IN.t15 4.89315
R3758 VCO_C_0.INV_2_3.IN.n51 VCO_C_0.INV_2_3.IN.n50 4.72831
R3759 VCO_C_0.INV_2_3.IN.n58 VCO_C_0.INV_2_3.IN.t23 4.70462
R3760 VCO_C_0.INV_2_3.IN.n59 VCO_C_0.INV_2_3.IN.t4 4.70337
R3761 VCO_C_0.INV_2_3.IN.n40 VCO_C_0.INV_2_3.IN.n36 4.55468
R3762 VCO_C_0.INV_2_3.IN VCO_C_0.INV_2_3.IN.n73 4.22145
R3763 VCO_C_0.INV_2_3.IN.n33 VCO_C_0.INV_2_3.IN.t14 4.04969
R3764 VCO_C_0.INV_2_3.IN.n40 VCO_C_0.INV_2_3.IN.n39 4.00854
R3765 VCO_C_0.INV_2_3.IN.n23 VCO_C_0.INV_2_3.IN.n22 4.00757
R3766 VCO_C_0.INV_2_3.IN.n4 VCO_C_0.INV_2_3.IN.t11 4.00481
R3767 VCO_C_0.INV_2_3.IN.n52 VCO_C_0.INV_2_3.IN.n48 3.90715
R3768 VCO_C_0.INV_2_3.IN.n75 VCO_C_0.INV_2_3.IN.n74 3.79925
R3769 VCO_C_0.INV_2_3.IN.n57 VCO_C_0.INV_2_3.IN.n56 3.77445
R3770 VCO_C_0.INV_2_3.IN.n26 VCO_C_0.INV_2_3.IN.n25 3.76954
R3771 VCO_C_0.INV_2_3.IN.n81 VCO_C_0.INV_2_3.IN.n79 3.76191
R3772 VCO_C_0.INV_2_3.IN.n79 VCO_C_0.INV_2_3.IN.t26 3.7183
R3773 VCO_C_0.INV_2_3.IN.n70 VCO_C_0.INV_2_3.IN.t55 3.6505
R3774 VCO_C_0.INV_2_3.IN.n71 VCO_C_0.INV_2_3.IN.t31 3.6505
R3775 VCO_C_0.INV_2_3.IN.n38 VCO_C_0.INV_2_3.IN.t16 3.6405
R3776 VCO_C_0.INV_2_3.IN.n38 VCO_C_0.INV_2_3.IN.n37 3.6405
R3777 VCO_C_0.INV_2_3.IN.n36 VCO_C_0.INV_2_3.IN.t13 3.6405
R3778 VCO_C_0.INV_2_3.IN.n36 VCO_C_0.INV_2_3.IN.n35 3.6405
R3779 VCO_C_0.INV_2_3.IN.n32 VCO_C_0.INV_2_3.IN.t12 3.6405
R3780 VCO_C_0.INV_2_3.IN.n32 VCO_C_0.INV_2_3.IN.n31 3.6405
R3781 VCO_C_0.INV_2_3.IN.n54 VCO_C_0.INV_2_3.IN.t24 3.47629
R3782 VCO_C_0.INV_2_3.IN.n56 VCO_C_0.INV_2_3.IN.t2 3.47627
R3783 VCO_C_0.INV_2_3.IN.n61 VCO_C_0.INV_2_3.IN.n60 3.3208
R3784 VCO_C_0.INV_2_3.IN.n26 VCO_C_0.INV_2_3.IN.t17 3.26269
R3785 VCO_C_0.INV_2_3.IN.n79 VCO_C_0.INV_2_3.IN.n78 3.25601
R3786 VCO_C_0.INV_2_3.IN.n73 VCO_C_0.INV_2_3.IN.n63 3.1807
R3787 VCO_C_0.INV_2_3.IN.n75 VCO_C_0.INV_2_3.IN.n62 3.14573
R3788 VCO_C_0.INV_2_3.IN.n58 VCO_C_0.INV_2_3.IN.n57 2.88663
R3789 VCO_C_0.INV_2_3.IN.n56 VCO_C_0.INV_2_3.IN.n55 2.86148
R3790 VCO_C_0.INV_2_3.IN.n54 VCO_C_0.INV_2_3.IN.n53 2.86147
R3791 VCO_C_0.INV_2_3.IN.n61 VCO_C_0.INV_2_3.IN.n52 2.83772
R3792 VCO_C_0.INV_2_3.IN.n28 VCO_C_0.INV_2_3.IN.n27 2.75932
R3793 VCO_C_0.INV_2_3.IN.n45 VCO_C_0.INV_2_3.IN.n3 2.62155
R3794 VCO_C_0.INV_2_3.IN.n74 VCO_C_0.INV_2_3.IN 2.36584
R3795 VCO_C_0.INV_2_3.IN.n76 VCO_C_0.INV_2_3.IN.n75 2.35159
R3796 VCO_C_0.INV_2_3.IN.n62 VCO_C_0.INV_2_3.IN 2.30603
R3797 VCO_C_0.INV_2_3.IN.n24 VCO_C_0.INV_2_3.IN.n23 2.2491
R3798 VCO_C_0.INV_2_3.IN.n34 VCO_C_0.INV_2_3.IN.n33 2.24586
R3799 VCO_C_0.INV_2_3.IN.n47 VCO_C_0.INV_2_3.IN.n46 2.03309
R3800 VCO_C_0.INV_2_3.IN.n74 VCO_C_0.INV_2_3.IN 1.93478
R3801 VCO_C_0.INV_2_3.IN.n27 VCO_C_0.INV_2_3.IN.n24 1.85135
R3802 VCO_C_0.INV_2_3.IN.n3 VCO_C_0.INV_2_3.IN.n44 1.79127
R3803 VCO_C_0.INV_2_3.IN.n41 VCO_C_0.INV_2_3.IN.n34 1.76701
R3804 VCO_C_0.INV_2_3.IN.n30 VCO_C_0.INV_2_3.IN.n4 1.50938
R3805 VCO_C_0.INV_2_3.IN.n27 VCO_C_0.INV_2_3.IN.n26 5.14667
R3806 VCO_C_0.INV_2_3.IN VCO_C_0.INV_2_3.IN.n1 3.15982
R3807 VCO_C_0.INV_2_3.IN.n3 VCO_C_0.INV_2_3.IN.n41 1.6295
R3808 VCO_C_0.INV_2_3.IN.n44 VCO_C_0.INV_2_3.IN.n43 1.495
R3809 VCO_C_0.INV_2_3.IN.n77 VCO_C_0.INV_2_3.IN.n76 1.47463
R3810 VCO_C_0.INV_2_3.IN.n39 VCO_C_0.INV_2_3.IN.n38 1.25653
R3811 VCO_C_0.INV_2_3.IN.n46 VCO_C_0.INV_2_3.IN.n45 1.22576
R3812 VCO_C_0.INV_2_3.IN.n29 VCO_C_0.INV_2_3.IN.n0 1.19023
R3813 VCO_C_0.INV_2_3.IN.n41 VCO_C_0.INV_2_3.IN.n40 1.1585
R3814 VCO_C_0.INV_2_3.IN.n28 VCO_C_0.INV_2_3.IN.n21 1.1379
R3815 VCO_C_0.INV_2_3.IN.n1 VCO_C_0.INV_2_3.IN.n77 0.931417
R3816 VCO_C_0.INV_2_3.IN.n1 VCO_C_0.INV_2_3.IN.n81 0.878898
R3817 VCO_C_0.INV_2_3.IN.n47 VCO_C_0.INV_2_3.IN.n30 0.836865
R3818 VCO_C_0.INV_2_3.IN.n18 VCO_C_0.INV_2_3.IN.n17 0.650226
R3819 VCO_C_0.INV_2_3.IN.n76 VCO_C_0.INV_2_3.IN.n47 0.597881
R3820 VCO_C_0.INV_2_3.IN.n62 VCO_C_0.INV_2_3.IN.n61 0.488268
R3821 VCO_C_0.INV_2_3.IN.n10 VCO_C_0.INV_2_3.IN.n9 0.487486
R3822 VCO_C_0.INV_2_3.IN.n52 VCO_C_0.INV_2_3.IN.n51 0.477758
R3823 VCO_C_0.INV_2_3.IN.n59 VCO_C_0.INV_2_3.IN.n58 0.472731
R3824 VCO_C_0.INV_2_3.IN.n0 VCO_C_0.INV_2_3.IN.n28 0.384538
R3825 VCO_C_0.INV_2_3.IN.n8 VCO_C_0.INV_2_3.IN.n7 0.345705
R3826 VCO_C_0.INV_2_3.IN.n20 VCO_C_0.INV_2_3.IN.n19 0.345705
R3827 VCO_C_0.INV_2_3.IN.n0 VCO_C_0.INV_2_3.IN.n20 0.34324
R3828 VCO_C_0.INV_2_3.IN.n13 VCO_C_0.INV_2_3.IN.n12 0.342007
R3829 VCO_C_0.INV_2_3.IN.n16 VCO_C_0.INV_2_3.IN.n15 0.342007
R3830 VCO_C_0.INV_2_3.IN.n12 VCO_C_0.INV_2_3.IN.n11 0.33461
R3831 VCO_C_0.INV_2_3.IN.n17 VCO_C_0.INV_2_3.IN.n16 0.325979
R3832 VCO_C_0.INV_2_3.IN.n19 VCO_C_0.INV_2_3.IN.n18 0.318582
R3833 VCO_C_0.INV_2_3.IN.n9 VCO_C_0.INV_2_3.IN.n8 0.312418
R3834 VCO_C_0.INV_2_3.IN.n14 VCO_C_0.INV_2_3.IN.n13 0.312418
R3835 VCO_C_0.INV_2_3.IN.n30 VCO_C_0.INV_2_3.IN.n29 0.216605
R3836 VCO_C_0.INV_2_3.IN.n10 VCO_C_0.INV_2_3.IN.n6 0.215773
R3837 VCO_C_0.INV_2_3.IN.n29 VCO_C_0.INV_2_3.IN.n14 0.198993
R3838 VCO_C_0.INV_2_3.IN.n11 VCO_C_0.INV_2_3.IN.n10 0.169404
R3839 VDD.n1087 VDD.n1086 102.362
R3840 VDD.n797 VDD.n796 102.362
R3841 VDD.n1481 VDD.t199 70.1759
R3842 VDD.n951 VDD.t245 70.1759
R3843 VDD.n1493 VDD.t250 67.252
R3844 VDD.n939 VDD.t214 67.252
R3845 VDD.n115 VDD.t77 60.7435
R3846 VDD.t132 VDD.n247 59.702
R3847 VDD.t76 VDD.n113 59.0509
R3848 VDD.n114 VDD.t76 52.7113
R3849 VDD.n248 VDD.t53 51.7418
R3850 VDD.t250 VDD.n1492 50.3542
R3851 VDD.t214 VDD.n938 49.9381
R3852 VDD.n248 VDD.t132 49.7517
R3853 VDD.t77 VDD.n114 49.6993
R3854 VDD.t245 VDD.n950 45.361
R3855 VDD.t199 VDD.n1480 45.361
R3856 VDD.n252 VDD.t123 43.7816
R3857 VDD.n247 VDD.t127 41.7915
R3858 VDD.n115 VDD.t56 41.6672
R3859 VDD.n1423 VDD.t26 39.6722
R3860 VDD.n1398 VDD.t387 39.6722
R3861 VDD.n1066 VDD.t259 39.6722
R3862 VDD.n1041 VDD.t96 39.6722
R3863 VDD.n1004 VDD.t101 39.6722
R3864 VDD.n479 VDD.t358 39.6722
R3865 VDD.n350 VDD.t156 39.6722
R3866 VDD.n1485 VDD.n1484 38.0122
R3867 VDD.n947 VDD.n946 38.0122
R3868 VDD.n16 VDD.t169 32.8322
R3869 VDD.n113 VDD.t78 24.6667
R3870 VDD.n667 VDD.t68 23.7307
R3871 VDD.n1007 VDD.n516 23.2342
R3872 VDD.n1417 VDD.t43 21.8883
R3873 VDD.n1392 VDD.t79 21.8883
R3874 VDD.n1060 VDD.t262 21.8883
R3875 VDD.n1024 VDD.t294 21.8883
R3876 VDD.n1014 VDD.t73 21.8883
R3877 VDD.n486 VDD.t355 21.8883
R3878 VDD.n363 VDD.t161 21.8883
R3879 VDD.n45 VDD.t87 21.8883
R3880 VDD.n1565 VDD.t18 21.6491
R3881 VDD.n1194 VDD.t205 21.2328
R3882 VDD.n1007 VDD.n1003 20.395
R3883 VDD.n317 VDD.t119 19.8363
R3884 VDD.n893 VDD.t111 17.4859
R3885 VDD.n1539 VDD.t2 17.0696
R3886 VDD.n1131 VDD.t8 14.5717
R3887 VDD.n702 VDD.t108 14.1554
R3888 VDD.n1408 VDD.t13 13.6804
R3889 VDD.n1383 VDD.t385 13.6804
R3890 VDD.n1051 VDD.t268 13.6804
R3891 VDD.n1031 VDD.t154 13.6804
R3892 VDD.n505 VDD.t311 13.6804
R3893 VDD.n496 VDD.t139 13.6804
R3894 VDD.n373 VDD.t150 13.6804
R3895 VDD.n36 VDD.t81 13.6804
R3896 VDD.n282 VDD.t50 10.9444
R3897 VDD.n1159 VDD.t29 9.99217
R3898 VDD.n1112 VDD.t202 9.99217
R3899 VDD.n720 VDD.t190 9.99217
R3900 VDD.n674 VDD.t66 9.57585
R3901 VDD.n413 VDD.t204 9.55982
R3902 VDD.n414 VDD.t242 9.55982
R3903 VDD.n415 VDD.t230 9.55982
R3904 VDD.n416 VDD.t232 9.55982
R3905 VDD.n579 VDD.t238 9.51591
R3906 VDD.n578 VDD.t207 9.51591
R3907 VDD.n577 VDD.t222 9.51591
R3908 VDD.n576 VDD.t195 9.51591
R3909 VDD.n1416 VDD.n1366 8.488
R3910 VDD.n1391 VDD.n1379 8.488
R3911 VDD.n1059 VDD.n453 8.488
R3912 VDD.n1017 VDD.n1013 8.488
R3913 VDD.n491 VDD.n489 8.488
R3914 VDD.n368 VDD.n366 8.488
R3915 VDD.n309 VDD.n285 8.488
R3916 VDD.n308 VDD.n306 8.488
R3917 VDD.n44 VDD.n32 8.488
R3918 VDD.n1418 VDD.n1416 8.2255
R3919 VDD.n1393 VDD.n1391 8.2255
R3920 VDD.n1061 VDD.n1059 8.2255
R3921 VDD.n1027 VDD.n1025 8.2255
R3922 VDD.n1017 VDD.n1015 8.2255
R3923 VDD.n489 VDD.n487 8.2255
R3924 VDD.n173 VDD.n171 8.2255
R3925 VDD.n366 VDD.n364 8.2255
R3926 VDD.n310 VDD.n309 8.2255
R3927 VDD.n308 VDD.n283 8.2255
R3928 VDD.n46 VDD.n44 8.2255
R3929 VDD.n856 VDD.t145 7.91057
R3930 VDD.n1571 VDD.t23 7.49426
R3931 VDD.n181 VDD.n179 7.1755
R3932 VDD.n1315 VDD.t368 6.94485
R3933 VDD.n729 VDD.n727 6.94485
R3934 VDD.n206 VDD.t317 6.84045
R3935 VDD.n151 VDD.t58 6.84045
R3936 VDD.n297 VDD.t113 6.84045
R3937 VDD.n1380 VDD.t390 6.70224
R3938 VDD.n1368 VDD.t15 6.70224
R3939 VDD.n1028 VDD.t301 6.70224
R3940 VDD.n467 VDD.n466 6.70224
R3941 VDD.n464 VDD.n462 6.70224
R3942 VDD.n455 VDD.t269 6.70224
R3943 VDD.n103 VDD.t423 6.70224
R3944 VDD.n74 VDD.n73 6.70224
R3945 VDD.n342 VDD.t151 6.70224
R3946 VDD.n288 VDD.n286 6.70224
R3947 VDD.n291 VDD.n290 6.70224
R3948 VDD.n33 VDD.t82 6.70224
R3949 VDD.n1002 VDD.t296 6.68489
R3950 VDD.n1432 VDD.n1430 6.68371
R3951 VDD.n1371 VDD.n1369 6.65503
R3952 VDD.n474 VDD.t359 6.65503
R3953 VDD.n458 VDD.n457 6.65503
R3954 VDD.n444 VDD.n443 6.65503
R3955 VDD.n105 VDD.t59 6.65503
R3956 VDD.n77 VDD.n75 6.65503
R3957 VDD.n345 VDD.n343 6.65503
R3958 VDD.n270 VDD.t401 6.65503
R3959 VDD.n2 VDD.n0 6.65503
R3960 VDD.n337 VDD.t120 6.64521
R3961 VDD.n1308 VDD.t219 6.43191
R3962 VDD.n1316 VDD.t240 6.43124
R3963 VDD.n1302 VDD.t201 6.4298
R3964 VDD.n742 VDD.t247 6.42961
R3965 VDD.n736 VDD.t235 6.37351
R3966 VDD.n1314 VDD.t192 6.37275
R3967 VDD.n730 VDD.t186 6.37256
R3968 VDD.n726 VDD.t189 6.37217
R3969 VDD.n818 VDD.t213 6.36486
R3970 VDD.n817 VDD.t244 6.36262
R3971 VDD.n517 VDD.t210 6.36128
R3972 VDD.n1358 VDD.t198 6.30795
R3973 VDD.n1357 VDD.t249 6.30193
R3974 VDD.n194 VDD.n193 6.3005
R3975 VDD.n95 VDD.n94 6.3005
R3976 VDD.n86 VDD.n85 6.3005
R3977 VDD.n378 VDD.n377 6.3005
R3978 VDD.n50 VDD.n49 6.3005
R3979 VDD.n49 VDD.n48 6.3005
R3980 VDD.n18 VDD.n17 6.3005
R3981 VDD.n17 VDD.n16 6.3005
R3982 VDD.n21 VDD.n20 6.3005
R3983 VDD.n53 VDD.n52 6.3005
R3984 VDD.n52 VDD.n51 6.3005
R3985 VDD.n432 VDD.t224 6.29942
R3986 VDD.n518 VDD.t227 6.29685
R3987 VDD.n337 VDD.t414 6.26273
R3988 VDD.n1432 VDD.n1431 6.24167
R3989 VDD.n1315 VDD.t335 6.2405
R3990 VDD.n1380 VDD.t386 6.2405
R3991 VDD.n1371 VDD.n1370 6.2405
R3992 VDD.n1368 VDD.t14 6.2405
R3993 VDD.n1028 VDD.t155 6.2405
R3994 VDD.n474 VDD.t374 6.2405
R3995 VDD.n467 VDD.n465 6.2405
R3996 VDD.n464 VDD.n463 6.2405
R3997 VDD.n729 VDD.n728 6.2405
R3998 VDD.n519 VDD.t229 6.2405
R3999 VDD.n1002 VDD.t102 6.2405
R4000 VDD.n458 VDD.n456 6.2405
R4001 VDD.n455 VDD.t282 6.2405
R4002 VDD.n444 VDD.n442 6.2405
R4003 VDD.n429 VDD.t218 6.2405
R4004 VDD.n103 VDD.t185 6.2405
R4005 VDD.n105 VDD.t337 6.2405
R4006 VDD.n77 VDD.n76 6.2405
R4007 VDD.n74 VDD.n72 6.2405
R4008 VDD.n345 VDD.n344 6.2405
R4009 VDD.n342 VDD.t176 6.2405
R4010 VDD.n291 VDD.n289 6.2405
R4011 VDD.n288 VDD.n287 6.2405
R4012 VDD.n270 VDD.t152 6.2405
R4013 VDD.n33 VDD.t83 6.2405
R4014 VDD.n2 VDD.n1 6.2405
R4015 VDD.n430 VDD.t216 6.23498
R4016 VDD.n122 VDD.n121 5.77744
R4017 VDD.n111 VDD.n110 5.77744
R4018 VDD.n242 VDD.t124 5.77744
R4019 VDD.n237 VDD.t179 5.77744
R4020 VDD.n1509 VDD.n1507 5.10682
R4021 VDD.n926 VDD.n924 5.10682
R4022 VDD.n112 VDD.t57 5.07264
R4023 VDD.n244 VDD.n243 5.07264
R4024 VDD.n239 VDD.n238 5.07264
R4025 VDD.n606 VDD.t196 4.99634
R4026 VDD.n127 VDD.t60 4.79075
R4027 VDD.n181 VDD.n180 4.5005
R4028 VDD.n191 VDD.n190 4.5005
R4029 VDD.n92 VDD.n91 4.5005
R4030 VDD.n91 VDD.n90 4.5005
R4031 VDD.n56 VDD.n55 4.5005
R4032 VDD.n55 VDD.n54 4.5005
R4033 VDD.n24 VDD.n23 4.5005
R4034 VDD.n23 VDD.n22 4.5005
R4035 VDD.n6 VDD.n5 4.5005
R4036 VDD.n1365 VDD.t5 4.10447
R4037 VDD.n1378 VDD.t61 4.10447
R4038 VDD.n452 VDD.t254 4.10447
R4039 VDD.n1037 VDD.t93 4.10447
R4040 VDD.n1012 VDD.t64 4.10447
R4041 VDD.n490 VDD.t142 4.10447
R4042 VDD.n367 VDD.t163 4.10447
R4043 VDD.n31 VDD.t84 4.10447
R4044 VDD.n419 VDD.t1 3.6405
R4045 VDD.n419 VDD.n418 3.6405
R4046 VDD.n1269 VDD.t266 3.6405
R4047 VDD.n1269 VDD.n1268 3.6405
R4048 VDD.n1272 VDD.t284 3.6405
R4049 VDD.n1272 VDD.n1271 3.6405
R4050 VDD.n1255 VDD.t20 3.6405
R4051 VDD.n1255 VDD.n1254 3.6405
R4052 VDD.n1558 VDD.t270 3.6405
R4053 VDD.n1558 VDD.n1557 3.6405
R4054 VDD.n1278 VDD.t267 3.6405
R4055 VDD.n1278 VDD.n1277 3.6405
R4056 VDD.n1281 VDD.t9 3.6405
R4057 VDD.n1281 VDD.n1280 3.6405
R4058 VDD.n1304 VDD.t369 3.6405
R4059 VDD.n1304 VDD.n1303 3.6405
R4060 VDD.n1306 VDD.t394 3.6405
R4061 VDD.n1306 VDD.n1305 3.6405
R4062 VDD.n1310 VDD.t395 3.6405
R4063 VDD.n1310 VDD.n1309 3.6405
R4064 VDD.n1312 VDD.t371 3.6405
R4065 VDD.n1312 VDD.n1311 3.6405
R4066 VDD.n1375 VDD.t89 3.6405
R4067 VDD.n1375 VDD.n1374 3.6405
R4068 VDD.n1373 VDD.t80 3.6405
R4069 VDD.n1373 VDD.n1372 3.6405
R4070 VDD.n1362 VDD.t45 3.6405
R4071 VDD.n1362 VDD.n1361 3.6405
R4072 VDD.n1360 VDD.t44 3.6405
R4073 VDD.n1360 VDD.n1359 3.6405
R4074 VDD.n1020 VDD.t302 3.6405
R4075 VDD.n1020 VDD.n1019 3.6405
R4076 VDD.n1022 VDD.t295 3.6405
R4077 VDD.n1022 VDD.n1021 3.6405
R4078 VDD.n469 VDD.t338 3.6405
R4079 VDD.n469 VDD.n468 3.6405
R4080 VDD.n471 VDD.t143 3.6405
R4081 VDD.n471 VDD.n470 3.6405
R4082 VDD.n515 VDD.t65 3.6405
R4083 VDD.n515 VDD.n514 3.6405
R4084 VDD.n513 VDD.t106 3.6405
R4085 VDD.n513 VDD.n512 3.6405
R4086 VDD.n740 VDD.t393 3.6405
R4087 VDD.n740 VDD.n739 3.6405
R4088 VDD.n738 VDD.t370 3.6405
R4089 VDD.n738 VDD.n737 3.6405
R4090 VDD.n734 VDD.t400 3.6405
R4091 VDD.n734 VDD.n733 3.6405
R4092 VDD.n732 VDD.t336 3.6405
R4093 VDD.n732 VDD.n731 3.6405
R4094 VDD.n573 VDD.t314 3.6405
R4095 VDD.n573 VDD.n572 3.6405
R4096 VDD.n559 VDD.t375 3.6405
R4097 VDD.n559 VDD.n558 3.6405
R4098 VDD.n543 VDD.t149 3.6405
R4099 VDD.n543 VDD.n542 3.6405
R4100 VDD.n530 VDD.t107 3.6405
R4101 VDD.n530 VDD.n529 3.6405
R4102 VDD.n523 VDD.t351 3.6405
R4103 VDD.n523 VDD.n522 3.6405
R4104 VDD.n526 VDD.t144 3.6405
R4105 VDD.n526 VDD.n525 3.6405
R4106 VDD.n538 VDD.t339 3.6405
R4107 VDD.n538 VDD.n537 3.6405
R4108 VDD.n535 VDD.t112 3.6405
R4109 VDD.n535 VDD.n534 3.6405
R4110 VDD.n551 VDD.t67 3.6405
R4111 VDD.n551 VDD.n550 3.6405
R4112 VDD.n554 VDD.t297 3.6405
R4113 VDD.n554 VDD.n553 3.6405
R4114 VDD.n569 VDD.t352 3.6405
R4115 VDD.n569 VDD.n568 3.6405
R4116 VDD.n566 VDD.t146 3.6405
R4117 VDD.n566 VDD.n565 3.6405
R4118 VDD.n562 VDD.t298 3.6405
R4119 VDD.n562 VDD.n561 3.6405
R4120 VDD.n832 VDD.t380 3.6405
R4121 VDD.n832 VDD.n831 3.6405
R4122 VDD.n828 VDD.t72 3.6405
R4123 VDD.n828 VDD.n827 3.6405
R4124 VDD.n546 VDD.t350 3.6405
R4125 VDD.n546 VDD.n545 3.6405
R4126 VDD.n447 VDD.t276 3.6405
R4127 VDD.n447 VDD.n446 3.6405
R4128 VDD.n449 VDD.t263 3.6405
R4129 VDD.n449 VDD.n448 3.6405
R4130 VDD.n1248 VDD.t273 3.6405
R4131 VDD.n1248 VDD.n1247 3.6405
R4132 VDD.n1251 VDD.t289 3.6405
R4133 VDD.n1251 VDD.n1250 3.6405
R4134 VDD.n1553 VDD.t40 3.6405
R4135 VDD.n1553 VDD.n1552 3.6405
R4136 VDD.n1550 VDD.t19 3.6405
R4137 VDD.n1550 VDD.n1549 3.6405
R4138 VDD.n1263 VDD.t17 3.6405
R4139 VDD.n1263 VDD.n1262 3.6405
R4140 VDD.n1266 VDD.t37 3.6405
R4141 VDD.n1266 VDD.n1265 3.6405
R4142 VDD.n426 VDD.t34 3.6405
R4143 VDD.n426 VDD.n425 3.6405
R4144 VDD.n422 VDD.t287 3.6405
R4145 VDD.n422 VDD.n421 3.6405
R4146 VDD.n1545 VDD.t288 3.6405
R4147 VDD.n1545 VDD.n1544 3.6405
R4148 VDD.n99 VDD.t418 3.6405
R4149 VDD.n99 VDD.n98 3.6405
R4150 VDD.n97 VDD.t346 3.6405
R4151 VDD.n97 VDD.n96 3.6405
R4152 VDD.n166 VDD.t321 3.6405
R4153 VDD.n166 VDD.n165 3.6405
R4154 VDD.n168 VDD.t322 3.6405
R4155 VDD.n168 VDD.n167 3.6405
R4156 VDD.n359 VDD.t162 3.6405
R4157 VDD.n359 VDD.n358 3.6405
R4158 VDD.n357 VDD.t404 3.6405
R4159 VDD.n357 VDD.n356 3.6405
R4160 VDD.n277 VDD.t49 3.6405
R4161 VDD.n277 VDD.n276 3.6405
R4162 VDD.n279 VDD.t116 3.6405
R4163 VDD.n279 VDD.n278 3.6405
R4164 VDD.n274 VDD.t405 3.6405
R4165 VDD.n274 VDD.n273 3.6405
R4166 VDD.n272 VDD.t168 3.6405
R4167 VDD.n272 VDD.n271 3.6405
R4168 VDD.n28 VDD.t88 3.6405
R4169 VDD.n28 VDD.n27 3.6405
R4170 VDD.n26 VDD.t153 3.6405
R4171 VDD.n26 VDD.n25 3.6405
R4172 VDD.n886 VDD.t136 3.33106
R4173 VDD.n411 VDD.n410 3.32815
R4174 VDD.n1307 VDD.n1306 3.30485
R4175 VDD.n1313 VDD.n1312 3.30485
R4176 VDD.n741 VDD.n738 3.30485
R4177 VDD.n735 VDD.n732 3.30485
R4178 VDD.n1106 VDD.n1104 3.28454
R4179 VDD.n579 VDD.t239 3.22394
R4180 VDD.n578 VDD.t209 3.22394
R4181 VDD.n577 VDD.t223 3.22394
R4182 VDD.n576 VDD.t197 3.22394
R4183 VDD.n413 VDD.t206 3.22347
R4184 VDD.n414 VDD.t243 3.22347
R4185 VDD.n415 VDD.t231 3.22347
R4186 VDD.n416 VDD.t234 3.22347
R4187 VDD.n1314 VDD.t194 3.21802
R4188 VDD.n730 VDD.t188 3.21788
R4189 VDD.n742 VDD.t248 3.21785
R4190 VDD.n1316 VDD.t241 3.21781
R4191 VDD.n726 VDD.t191 3.21767
R4192 VDD.n1302 VDD.t203 3.21766
R4193 VDD.n783 VDD.n782 3.21752
R4194 VDD.n1308 VDD.t221 3.21671
R4195 VDD.n736 VDD.t237 3.21657
R4196 VDD.n1358 VDD.t200 3.19864
R4197 VDD.n517 VDD.t212 3.19113
R4198 VDD.n432 VDD.t226 3.19113
R4199 VDD.n817 VDD.t246 3.18927
R4200 VDD.n1357 VDD.t251 3.1878
R4201 VDD.n818 VDD.t215 3.1878
R4202 VDD.n634 VDD.n575 3.16769
R4203 VDD.n1200 VDD.n417 3.16769
R4204 VDD.n116 VDD.n115 3.15287
R4205 VDD.n114 VDD 3.15287
R4206 VDD.n253 VDD.n252 3.15287
R4207 VDD.n249 VDD.n248 3.15287
R4208 VDD.n247 VDD.n246 3.15287
R4209 VDD.n929 VDD.n821 3.15151
R4210 VDD.n1595 VDD.n1594 3.1505
R4211 VDD.n1594 VDD.n1593 3.1505
R4212 VDD.n1501 VDD.n1356 3.1505
R4213 VDD.n1500 VDD.n1499 3.1505
R4214 VDD.n1495 VDD.n1494 3.1505
R4215 VDD.n1494 VDD.n1493 3.1505
R4216 VDD.n1490 VDD.n1489 3.1505
R4217 VDD.n1489 VDD.n1488 3.1505
R4218 VDD.n1487 VDD.n1486 3.1505
R4219 VDD.n1486 VDD.n1485 3.1505
R4220 VDD.n1483 VDD.n1482 3.1505
R4221 VDD.n1482 VDD.n1481 3.1505
R4222 VDD.n1478 VDD.n1477 3.1505
R4223 VDD.n1477 VDD.n1476 3.1505
R4224 VDD.n1475 VDD.n1474 3.1505
R4225 VDD.n1498 VDD.n1497 3.1505
R4226 VDD.n1497 VDD.n1496 3.1505
R4227 VDD.n1472 VDD.n1471 3.1505
R4228 VDD.n1389 VDD.n1379 3.1505
R4229 VDD.n1379 VDD.n1378 3.1505
R4230 VDD.n1388 VDD.n1387 3.1505
R4231 VDD.n1387 VDD.n1386 3.1505
R4232 VDD.n1385 VDD.n1384 3.1505
R4233 VDD.n1384 VDD.n1383 3.1505
R4234 VDD.n1382 VDD.n1381 3.1505
R4235 VDD.n1403 VDD.n1402 3.1505
R4236 VDD.n1400 VDD.n1399 3.1505
R4237 VDD.n1399 VDD.n1398 3.1505
R4238 VDD.n1397 VDD.n1396 3.1505
R4239 VDD.n1396 VDD.n1395 3.1505
R4240 VDD.n1394 VDD.n1393 3.1505
R4241 VDD.n1393 VDD.n1392 3.1505
R4242 VDD.n1391 VDD 3.1505
R4243 VDD.n1391 VDD.n1390 3.1505
R4244 VDD.n1407 VDD.n1367 3.1505
R4245 VDD.n1414 VDD.n1366 3.1505
R4246 VDD.n1366 VDD.n1365 3.1505
R4247 VDD.n1413 VDD.n1412 3.1505
R4248 VDD.n1412 VDD.n1411 3.1505
R4249 VDD.n1410 VDD.n1409 3.1505
R4250 VDD.n1409 VDD.n1408 3.1505
R4251 VDD.n1428 VDD.n1427 3.1505
R4252 VDD.n1425 VDD.n1424 3.1505
R4253 VDD.n1424 VDD.n1423 3.1505
R4254 VDD.n1422 VDD.n1421 3.1505
R4255 VDD.n1421 VDD.n1420 3.1505
R4256 VDD.n1419 VDD.n1418 3.1505
R4257 VDD.n1418 VDD.n1417 3.1505
R4258 VDD.n1416 VDD 3.1505
R4259 VDD.n1416 VDD.n1415 3.1505
R4260 VDD.n1469 VDD.n1468 3.1505
R4261 VDD.n1465 VDD.n1464 3.1505
R4262 VDD.n1462 VDD.n1461 3.1505
R4263 VDD.n1459 VDD.n1458 3.1505
R4264 VDD.n1456 VDD.n1455 3.1505
R4265 VDD.n1453 VDD.n1452 3.1505
R4266 VDD.n1450 VDD.n1449 3.1505
R4267 VDD.n1447 VDD.n1446 3.1505
R4268 VDD.n1444 VDD.n1443 3.1505
R4269 VDD.n1441 VDD.n1440 3.1505
R4270 VDD.n1438 VDD.n1437 3.1505
R4271 VDD.n1435 VDD.n1434 3.1505
R4272 VDD.n435 VDD.n434 3.1505
R4273 VDD.n438 VDD.n437 3.1505
R4274 VDD.n441 VDD.n440 3.1505
R4275 VDD.n1030 VDD.n1029 3.1505
R4276 VDD VDD.n1027 3.1505
R4277 VDD.n1027 VDD.n1026 3.1505
R4278 VDD.n1039 VDD.n1038 3.1505
R4279 VDD.n1038 VDD.n1037 3.1505
R4280 VDD.n1036 VDD.n1035 3.1505
R4281 VDD.n1035 VDD.n1034 3.1505
R4282 VDD.n1033 VDD.n1032 3.1505
R4283 VDD.n1032 VDD.n1031 3.1505
R4284 VDD.n489 VDD 3.1505
R4285 VDD.n489 VDD.n488 3.1505
R4286 VDD.n487 VDD.n485 3.1505
R4287 VDD.n487 VDD.n486 3.1505
R4288 VDD.n484 VDD.n483 3.1505
R4289 VDD.n483 VDD.n482 3.1505
R4290 VDD.n481 VDD.n480 3.1505
R4291 VDD.n480 VDD.n479 3.1505
R4292 VDD.n478 VDD.n477 3.1505
R4293 VDD.n500 VDD.n499 3.1505
R4294 VDD.n498 VDD.n497 3.1505
R4295 VDD.n497 VDD.n496 3.1505
R4296 VDD.n495 VDD.n494 3.1505
R4297 VDD.n494 VDD.n493 3.1505
R4298 VDD.n492 VDD.n491 3.1505
R4299 VDD.n491 VDD.n490 3.1505
R4300 VDD.n510 VDD.n509 3.1505
R4301 VDD.n509 VDD.n508 3.1505
R4302 VDD.n507 VDD.n506 3.1505
R4303 VDD.n506 VDD.n505 3.1505
R4304 VDD.n504 VDD.n503 3.1505
R4305 VDD.n633 VDD.n632 3.1505
R4306 VDD.n632 VDD.n631 3.1505
R4307 VDD.n630 VDD.n629 3.1505
R4308 VDD.n629 VDD.n628 3.1505
R4309 VDD.n627 VDD.n626 3.1505
R4310 VDD.n626 VDD.n625 3.1505
R4311 VDD.n623 VDD.n622 3.1505
R4312 VDD.n622 VDD.n621 3.1505
R4313 VDD.n620 VDD.n619 3.1505
R4314 VDD.n619 VDD.n618 3.1505
R4315 VDD.n617 VDD.n616 3.1505
R4316 VDD.n616 VDD.n615 3.1505
R4317 VDD.n614 VDD.n613 3.1505
R4318 VDD.n613 VDD.n612 3.1505
R4319 VDD.n610 VDD.n609 3.1505
R4320 VDD.n609 VDD.n608 3.1505
R4321 VDD.n605 VDD.n604 3.1505
R4322 VDD.n604 VDD.n603 3.1505
R4323 VDD.n602 VDD.n601 3.1505
R4324 VDD.n601 VDD.n600 3.1505
R4325 VDD.n598 VDD.n597 3.1505
R4326 VDD.n597 VDD.n596 3.1505
R4327 VDD.n595 VDD.n594 3.1505
R4328 VDD.n594 VDD.n593 3.1505
R4329 VDD.n592 VDD.n591 3.1505
R4330 VDD.n591 VDD.n590 3.1505
R4331 VDD.n589 VDD.n588 3.1505
R4332 VDD.n588 VDD.n587 3.1505
R4333 VDD.n585 VDD.n584 3.1505
R4334 VDD.n584 VDD.n583 3.1505
R4335 VDD.n582 VDD.n581 3.1505
R4336 VDD.n638 VDD.n637 3.1505
R4337 VDD.n641 VDD.n640 3.1505
R4338 VDD.n640 VDD.n639 3.1505
R4339 VDD.n644 VDD.n643 3.1505
R4340 VDD.n643 VDD.n642 3.1505
R4341 VDD.n647 VDD.n646 3.1505
R4342 VDD.n646 VDD.n645 3.1505
R4343 VDD.n650 VDD.n649 3.1505
R4344 VDD.n649 VDD.n648 3.1505
R4345 VDD.n653 VDD.n652 3.1505
R4346 VDD.n652 VDD.n651 3.1505
R4347 VDD.n656 VDD.n655 3.1505
R4348 VDD.n655 VDD.n654 3.1505
R4349 VDD.n660 VDD.n659 3.1505
R4350 VDD.n659 VDD.n658 3.1505
R4351 VDD.n663 VDD.n662 3.1505
R4352 VDD.n662 VDD.n661 3.1505
R4353 VDD.n666 VDD.n665 3.1505
R4354 VDD.n665 VDD.n664 3.1505
R4355 VDD.n669 VDD.n668 3.1505
R4356 VDD.n668 VDD.n667 3.1505
R4357 VDD.n673 VDD.n672 3.1505
R4358 VDD.n672 VDD.n671 3.1505
R4359 VDD.n676 VDD.n675 3.1505
R4360 VDD.n675 VDD.n674 3.1505
R4361 VDD.n679 VDD.n678 3.1505
R4362 VDD.n678 VDD.n677 3.1505
R4363 VDD.n682 VDD.n681 3.1505
R4364 VDD.n681 VDD.n680 3.1505
R4365 VDD.n685 VDD.n684 3.1505
R4366 VDD.n684 VDD.n683 3.1505
R4367 VDD.n688 VDD.n687 3.1505
R4368 VDD.n687 VDD.n686 3.1505
R4369 VDD.n691 VDD.n690 3.1505
R4370 VDD.n690 VDD.n689 3.1505
R4371 VDD.n695 VDD.n694 3.1505
R4372 VDD.n694 VDD.n693 3.1505
R4373 VDD.n698 VDD.n697 3.1505
R4374 VDD.n697 VDD.n696 3.1505
R4375 VDD.n701 VDD.n700 3.1505
R4376 VDD.n700 VDD.n699 3.1505
R4377 VDD.n704 VDD.n703 3.1505
R4378 VDD.n703 VDD.n702 3.1505
R4379 VDD.n708 VDD.n707 3.1505
R4380 VDD.n707 VDD.n706 3.1505
R4381 VDD.n710 VDD.n709 3.1505
R4382 VDD.n709 VDD.t71 3.1505
R4383 VDD.n713 VDD.n712 3.1505
R4384 VDD.n712 VDD.n711 3.1505
R4385 VDD.n716 VDD.n715 3.1505
R4386 VDD.n715 VDD.n714 3.1505
R4387 VDD.n719 VDD.n718 3.1505
R4388 VDD.n718 VDD.n717 3.1505
R4389 VDD.n722 VDD.n721 3.1505
R4390 VDD.n721 VDD.n720 3.1505
R4391 VDD.n725 VDD.n724 3.1505
R4392 VDD.n724 VDD.n723 3.1505
R4393 VDD.n962 VDD.n961 3.1505
R4394 VDD.n960 VDD.n959 3.1505
R4395 VDD.n957 VDD.n956 3.1505
R4396 VDD.n956 VDD.n955 3.1505
R4397 VDD.n953 VDD.n952 3.1505
R4398 VDD.n952 VDD.n951 3.1505
R4399 VDD.n949 VDD.n948 3.1505
R4400 VDD.n948 VDD.n947 3.1505
R4401 VDD.n945 VDD.n944 3.1505
R4402 VDD.n944 VDD.n943 3.1505
R4403 VDD.n941 VDD.n940 3.1505
R4404 VDD.n940 VDD.n939 3.1505
R4405 VDD.n937 VDD.n936 3.1505
R4406 VDD.n936 VDD.n935 3.1505
R4407 VDD.n931 VDD.n930 3.1505
R4408 VDD.n934 VDD.n933 3.1505
R4409 VDD.n839 VDD.n838 3.1505
R4410 VDD.n838 VDD.n837 3.1505
R4411 VDD.n836 VDD.n835 3.1505
R4412 VDD.n821 VDD.n820 3.1505
R4413 VDD.n927 VDD.n926 3.1505
R4414 VDD.n926 VDD.n925 3.1505
R4415 VDD.n923 VDD.n922 3.1505
R4416 VDD.n922 VDD.n921 3.1505
R4417 VDD.n920 VDD.n919 3.1505
R4418 VDD.n919 VDD.n918 3.1505
R4419 VDD.n917 VDD.n916 3.1505
R4420 VDD.n916 VDD.n915 3.1505
R4421 VDD.n914 VDD.n913 3.1505
R4422 VDD.n913 VDD.n912 3.1505
R4423 VDD.n911 VDD.n910 3.1505
R4424 VDD.n910 VDD.n909 3.1505
R4425 VDD.n908 VDD.n907 3.1505
R4426 VDD.n907 VDD.n906 3.1505
R4427 VDD.n904 VDD.n903 3.1505
R4428 VDD.n903 VDD.n902 3.1505
R4429 VDD.n901 VDD.n900 3.1505
R4430 VDD.n900 VDD.n899 3.1505
R4431 VDD.n898 VDD.n897 3.1505
R4432 VDD.n897 VDD.n896 3.1505
R4433 VDD.n895 VDD.n894 3.1505
R4434 VDD.n894 VDD.n893 3.1505
R4435 VDD.n891 VDD.n890 3.1505
R4436 VDD.n890 VDD.n889 3.1505
R4437 VDD.n888 VDD.n887 3.1505
R4438 VDD.n887 VDD.n886 3.1505
R4439 VDD.n885 VDD.n884 3.1505
R4440 VDD.n884 VDD.n883 3.1505
R4441 VDD.n882 VDD.n881 3.1505
R4442 VDD.n881 VDD.n880 3.1505
R4443 VDD.n879 VDD.n878 3.1505
R4444 VDD.n878 VDD.n877 3.1505
R4445 VDD.n876 VDD.n875 3.1505
R4446 VDD.n875 VDD.n874 3.1505
R4447 VDD.n873 VDD.n872 3.1505
R4448 VDD.n872 VDD.n871 3.1505
R4449 VDD.n867 VDD.n866 3.1505
R4450 VDD.n866 VDD.n865 3.1505
R4451 VDD.n864 VDD.n863 3.1505
R4452 VDD.n863 VDD.n862 3.1505
R4453 VDD.n861 VDD.n860 3.1505
R4454 VDD.n860 VDD.n859 3.1505
R4455 VDD.n858 VDD.n857 3.1505
R4456 VDD.n857 VDD.n856 3.1505
R4457 VDD.n854 VDD.n853 3.1505
R4458 VDD.n853 VDD.n852 3.1505
R4459 VDD.n851 VDD.n850 3.1505
R4460 VDD.n850 VDD.n849 3.1505
R4461 VDD.n848 VDD.n847 3.1505
R4462 VDD.n847 VDD.n846 3.1505
R4463 VDD.n845 VDD.n844 3.1505
R4464 VDD.n844 VDD.n843 3.1505
R4465 VDD.n842 VDD.n841 3.1505
R4466 VDD.n841 VDD.n840 3.1505
R4467 VDD.n826 VDD.n825 3.1505
R4468 VDD.n823 VDD.n822 3.1505
R4469 VDD.n746 VDD.n745 3.1505
R4470 VDD.n749 VDD.n748 3.1505
R4471 VDD.n751 VDD.n750 3.1505
R4472 VDD.n753 VDD.n752 3.1505
R4473 VDD.n757 VDD.n756 3.1505
R4474 VDD.n760 VDD.n759 3.1505
R4475 VDD.n763 VDD.n762 3.1505
R4476 VDD.n766 VDD.n765 3.1505
R4477 VDD.n769 VDD.n768 3.1505
R4478 VDD.n772 VDD.n771 3.1505
R4479 VDD.n776 VDD.n775 3.1505
R4480 VDD.n778 VDD.n777 3.1505
R4481 VDD.n784 VDD.n783 3.1505
R4482 VDD.n809 VDD.n808 3.1505
R4483 VDD.n806 VDD.n805 3.1505
R4484 VDD.n805 VDD.n804 3.1505
R4485 VDD.n802 VDD.n801 3.1505
R4486 VDD.n801 VDD.n800 3.1505
R4487 VDD.n799 VDD.n798 3.1505
R4488 VDD.n798 VDD.n797 3.1505
R4489 VDD.n795 VDD.n794 3.1505
R4490 VDD.n794 VDD.n793 3.1505
R4491 VDD.n791 VDD.n790 3.1505
R4492 VDD.n787 VDD.n786 3.1505
R4493 VDD.n811 VDD.n810 3.1505
R4494 VDD.n814 VDD.n813 3.1505
R4495 VDD.n816 VDD.n815 3.1505
R4496 VDD.n997 VDD.n996 3.1505
R4497 VDD.n994 VDD.n993 3.1505
R4498 VDD.n991 VDD.n990 3.1505
R4499 VDD.n988 VDD.n987 3.1505
R4500 VDD.n985 VDD.n984 3.1505
R4501 VDD.n982 VDD.n981 3.1505
R4502 VDD.n979 VDD.n978 3.1505
R4503 VDD.n976 VDD.n975 3.1505
R4504 VDD.n973 VDD.n972 3.1505
R4505 VDD.n970 VDD.n969 3.1505
R4506 VDD.n967 VDD.n966 3.1505
R4507 VDD.n965 VDD.n964 3.1505
R4508 VDD.n1001 VDD.n1000 3.1505
R4509 VDD.n1013 VDD.n511 3.1505
R4510 VDD.n1013 VDD.n1012 3.1505
R4511 VDD VDD.n1017 3.1505
R4512 VDD.n1017 VDD.n1016 3.1505
R4513 VDD.n1015 VDD.n1011 3.1505
R4514 VDD.n1015 VDD.n1014 3.1505
R4515 VDD.n1010 VDD.n1009 3.1505
R4516 VDD.n1009 VDD.n1008 3.1505
R4517 VDD.n1005 VDD.n1004 3.1505
R4518 VDD.n1025 VDD.n1024 3.1505
R4519 VDD.n460 VDD.n459 3.1505
R4520 VDD.n1046 VDD.n1045 3.1505
R4521 VDD.n1043 VDD.n1042 3.1505
R4522 VDD.n1042 VDD.n1041 3.1505
R4523 VDD.n1050 VDD.n454 3.1505
R4524 VDD.n1057 VDD.n453 3.1505
R4525 VDD.n453 VDD.n452 3.1505
R4526 VDD.n1056 VDD.n1055 3.1505
R4527 VDD.n1055 VDD.n1054 3.1505
R4528 VDD.n1053 VDD.n1052 3.1505
R4529 VDD.n1052 VDD.n1051 3.1505
R4530 VDD.n1071 VDD.n1070 3.1505
R4531 VDD.n1068 VDD.n1067 3.1505
R4532 VDD.n1067 VDD.n1066 3.1505
R4533 VDD.n1065 VDD.n1064 3.1505
R4534 VDD.n1064 VDD.n1063 3.1505
R4535 VDD.n1062 VDD.n1061 3.1505
R4536 VDD.n1061 VDD.n1060 3.1505
R4537 VDD.n1059 VDD 3.1505
R4538 VDD.n1059 VDD.n1058 3.1505
R4539 VDD.n1099 VDD.n1098 3.1505
R4540 VDD.n1096 VDD.n1095 3.1505
R4541 VDD.n1092 VDD.n1091 3.1505
R4542 VDD.n1091 VDD.n1090 3.1505
R4543 VDD.n1089 VDD.n1088 3.1505
R4544 VDD.n1088 VDD.n1087 3.1505
R4545 VDD.n1085 VDD.n1084 3.1505
R4546 VDD.n1084 VDD.n1083 3.1505
R4547 VDD.n1081 VDD.n1080 3.1505
R4548 VDD.n1080 VDD.n1079 3.1505
R4549 VDD.n1078 VDD.n1077 3.1505
R4550 VDD.n1075 VDD.n1074 3.1505
R4551 VDD.n1103 VDD.n1102 3.1505
R4552 VDD.n1101 VDD.n1100 3.1505
R4553 VDD.n1319 VDD.n1318 3.1505
R4554 VDD.n1322 VDD.n1321 3.1505
R4555 VDD.n1325 VDD.n1324 3.1505
R4556 VDD.n1328 VDD.n1327 3.1505
R4557 VDD.n1331 VDD.n1330 3.1505
R4558 VDD.n1334 VDD.n1333 3.1505
R4559 VDD.n1338 VDD.n1337 3.1505
R4560 VDD.n1340 VDD.n1339 3.1505
R4561 VDD.n1343 VDD.n1342 3.1505
R4562 VDD.n1346 VDD.n1345 3.1505
R4563 VDD.n1352 VDD.n1351 3.1505
R4564 VDD.n1354 VDD.n1353 3.1505
R4565 VDD.n1107 VDD.n1106 3.1505
R4566 VDD.n1505 VDD.n1504 3.1505
R4567 VDD.n1504 VDD.n1503 3.1505
R4568 VDD.n1513 VDD.n1512 3.1505
R4569 VDD.n1512 VDD.n1511 3.1505
R4570 VDD.n1510 VDD.n1509 3.1505
R4571 VDD.n1509 VDD.n1508 3.1505
R4572 VDD.n1528 VDD.n1527 3.1505
R4573 VDD.n1527 VDD.n1526 3.1505
R4574 VDD.n1525 VDD.n1524 3.1505
R4575 VDD.n1524 VDD.n1523 3.1505
R4576 VDD.n1522 VDD.n1521 3.1505
R4577 VDD.n1521 VDD.n1520 3.1505
R4578 VDD.n1519 VDD.n1518 3.1505
R4579 VDD.n1518 VDD.n1517 3.1505
R4580 VDD.n1516 VDD.n1515 3.1505
R4581 VDD.n1515 VDD.n1514 3.1505
R4582 VDD.n1589 VDD.n1588 3.1505
R4583 VDD.n1588 VDD.n1587 3.1505
R4584 VDD.n1586 VDD.n1585 3.1505
R4585 VDD.n1585 VDD.n1584 3.1505
R4586 VDD.n1583 VDD.n1582 3.1505
R4587 VDD.n1582 VDD.n1581 3.1505
R4588 VDD.n1580 VDD.n1579 3.1505
R4589 VDD.n1579 VDD.n1578 3.1505
R4590 VDD.n1577 VDD.n1576 3.1505
R4591 VDD.n1576 VDD.n1575 3.1505
R4592 VDD.n1573 VDD.n1572 3.1505
R4593 VDD.n1572 VDD.n1571 3.1505
R4594 VDD.n1570 VDD.n1569 3.1505
R4595 VDD.n1569 VDD.n1568 3.1505
R4596 VDD.n1567 VDD.n1566 3.1505
R4597 VDD.n1566 VDD.n1565 3.1505
R4598 VDD.n1564 VDD.n1563 3.1505
R4599 VDD.n1563 VDD.n1562 3.1505
R4600 VDD.n1260 VDD.n1259 3.1505
R4601 VDD.n1259 VDD.n1258 3.1505
R4602 VDD.n1286 VDD.n1285 3.1505
R4603 VDD.n1285 VDD.n1284 3.1505
R4604 VDD.n1289 VDD.n1288 3.1505
R4605 VDD.n1288 VDD.n1287 3.1505
R4606 VDD.n1292 VDD.n1291 3.1505
R4607 VDD.n1291 VDD.n1290 3.1505
R4608 VDD.n1295 VDD.n1294 3.1505
R4609 VDD.n1294 VDD.n1293 3.1505
R4610 VDD.n1298 VDD.n1297 3.1505
R4611 VDD.n1297 VDD.n1296 3.1505
R4612 VDD.n1301 VDD.n1300 3.1505
R4613 VDD.n1300 VDD.n1299 3.1505
R4614 VDD.n1541 VDD.n1540 3.1505
R4615 VDD.n1540 VDD.n1539 3.1505
R4616 VDD.n1538 VDD.n1537 3.1505
R4617 VDD.n1537 VDD.n1536 3.1505
R4618 VDD.n1535 VDD.n1534 3.1505
R4619 VDD.n1534 VDD.n1533 3.1505
R4620 VDD.n1532 VDD.n1531 3.1505
R4621 VDD.n1531 VDD.n1530 3.1505
R4622 VDD.n1592 VDD.n1591 3.1505
R4623 VDD.n1591 VDD.n1590 3.1505
R4624 VDD.n1199 VDD.n1198 3.1505
R4625 VDD.n1198 VDD.n1197 3.1505
R4626 VDD.n1196 VDD.n1195 3.1505
R4627 VDD.n1195 VDD.n1194 3.1505
R4628 VDD.n1193 VDD.n1192 3.1505
R4629 VDD.n1192 VDD.n1191 3.1505
R4630 VDD.n1190 VDD.n1189 3.1505
R4631 VDD.n1189 VDD.n1188 3.1505
R4632 VDD.n1187 VDD.n1186 3.1505
R4633 VDD.n1186 VDD.n1185 3.1505
R4634 VDD.n1184 VDD.n1183 3.1505
R4635 VDD.n1183 VDD.n1182 3.1505
R4636 VDD.n1181 VDD.n1180 3.1505
R4637 VDD.n1180 VDD.n1179 3.1505
R4638 VDD.n1177 VDD.n1176 3.1505
R4639 VDD.n1176 VDD.n1175 3.1505
R4640 VDD.n1174 VDD.n1173 3.1505
R4641 VDD.n1173 VDD.n1172 3.1505
R4642 VDD.n1171 VDD.n1170 3.1505
R4643 VDD.n1170 VDD.n1169 3.1505
R4644 VDD.n1168 VDD.n1167 3.1505
R4645 VDD.n1167 VDD.n1166 3.1505
R4646 VDD.n1164 VDD.n1163 3.1505
R4647 VDD.n1163 VDD.n1162 3.1505
R4648 VDD.n1161 VDD.n1160 3.1505
R4649 VDD.n1160 VDD.n1159 3.1505
R4650 VDD.n1158 VDD.n1157 3.1505
R4651 VDD.n1157 VDD.n1156 3.1505
R4652 VDD.n1155 VDD.n1154 3.1505
R4653 VDD.n1154 VDD.n1153 3.1505
R4654 VDD.n1152 VDD.n1151 3.1505
R4655 VDD.n1151 VDD.n1150 3.1505
R4656 VDD.n1149 VDD.n1148 3.1505
R4657 VDD.n1148 VDD.n1147 3.1505
R4658 VDD.n1146 VDD.n1145 3.1505
R4659 VDD.n1145 VDD.n1144 3.1505
R4660 VDD.n1142 VDD.n1141 3.1505
R4661 VDD.n1141 VDD.n1140 3.1505
R4662 VDD.n1139 VDD.n1138 3.1505
R4663 VDD.n1138 VDD.n1137 3.1505
R4664 VDD.n1136 VDD.n1135 3.1505
R4665 VDD.n1135 VDD.n1134 3.1505
R4666 VDD.n1133 VDD.n1132 3.1505
R4667 VDD.n1132 VDD.n1131 3.1505
R4668 VDD.n1129 VDD.n1128 3.1505
R4669 VDD.n1128 VDD.n1127 3.1505
R4670 VDD.n1126 VDD.n1125 3.1505
R4671 VDD.n1125 VDD.n1124 3.1505
R4672 VDD.n1123 VDD.n1122 3.1505
R4673 VDD.n1122 VDD.n1121 3.1505
R4674 VDD.n1120 VDD.n1119 3.1505
R4675 VDD.n1119 VDD.n1118 3.1505
R4676 VDD.n1117 VDD.n1116 3.1505
R4677 VDD.n1116 VDD.n1115 3.1505
R4678 VDD.n1114 VDD.n1113 3.1505
R4679 VDD.n1113 VDD.n1112 3.1505
R4680 VDD.n1111 VDD.n1110 3.1505
R4681 VDD.n1110 VDD.n1109 3.1505
R4682 VDD.n1203 VDD.n1202 3.1505
R4683 VDD.n1205 VDD.n1204 3.1505
R4684 VDD.n1207 VDD.n1206 3.1505
R4685 VDD.n1210 VDD.n1209 3.1505
R4686 VDD.n1212 VDD.n1211 3.1505
R4687 VDD.n1215 VDD.n1214 3.1505
R4688 VDD.n1217 VDD.n1216 3.1505
R4689 VDD.n1221 VDD.n1220 3.1505
R4690 VDD.n1223 VDD.n1222 3.1505
R4691 VDD.n1226 VDD.n1225 3.1505
R4692 VDD.n1229 VDD.n1228 3.1505
R4693 VDD.n1232 VDD.n1231 3.1505
R4694 VDD.n1234 VDD.n1233 3.1505
R4695 VDD.n1237 VDD.n1236 3.1505
R4696 VDD.n1240 VDD.n1239 3.1505
R4697 VDD.n1245 VDD.n1244 3.1505
R4698 VDD.n135 VDD.n104 3.1505
R4699 VDD.n171 VDD.n164 3.1505
R4700 VDD.n171 VDD.n170 3.1505
R4701 VDD.n162 VDD.n161 3.1505
R4702 VDD.n161 VDD.n160 3.1505
R4703 VDD.n156 VDD.n155 3.1505
R4704 VDD.n155 VDD.n154 3.1505
R4705 VDD.n149 VDD.n148 3.1505
R4706 VDD.n148 VDD.n147 3.1505
R4707 VDD.n163 VDD.n102 3.1505
R4708 VDD.n102 VDD.n101 3.1505
R4709 VDD.n159 VDD.n158 3.1505
R4710 VDD.n158 VDD.n157 3.1505
R4711 VDD.n153 VDD.n152 3.1505
R4712 VDD.n152 VDD.n151 3.1505
R4713 VDD VDD.n173 3.1505
R4714 VDD.n173 VDD.n172 3.1505
R4715 VDD.n179 VDD 3.1505
R4716 VDD.n179 VDD.n178 3.1505
R4717 VDD.n208 VDD.n207 3.1505
R4718 VDD.n207 VDD.n206 3.1505
R4719 VDD.n201 VDD.n200 3.1505
R4720 VDD.n200 VDD.n199 3.1505
R4721 VDD.n188 VDD.n187 3.1505
R4722 VDD.n187 VDD.n186 3.1505
R4723 VDD.n83 VDD.n82 3.1505
R4724 VDD.n82 VDD.n81 3.1505
R4725 VDD.n195 VDD.n192 3.1505
R4726 VDD.n196 VDD.n195 3.1505
R4727 VDD.n184 VDD.n183 3.1505
R4728 VDD.n183 VDD.n182 3.1505
R4729 VDD.n88 VDD.n87 3.1505
R4730 VDD.n79 VDD.n78 3.1505
R4731 VDD.n89 VDD.n88 3.1505
R4732 VDD.n205 VDD.n204 3.1505
R4733 VDD.n204 VDD.n203 3.1505
R4734 VDD.n349 VDD.n348 3.1505
R4735 VDD.n352 VDD.n351 3.1505
R4736 VDD.n351 VDD.n350 3.1505
R4737 VDD.n355 VDD.n354 3.1505
R4738 VDD.n354 VDD.n353 3.1505
R4739 VDD.n364 VDD.n362 3.1505
R4740 VDD.n364 VDD.n363 3.1505
R4741 VDD.n366 VDD 3.1505
R4742 VDD.n366 VDD.n365 3.1505
R4743 VDD.n369 VDD.n368 3.1505
R4744 VDD.n368 VDD.n367 3.1505
R4745 VDD.n372 VDD.n371 3.1505
R4746 VDD.n371 VDD.n370 3.1505
R4747 VDD.n375 VDD.n374 3.1505
R4748 VDD.n374 VDD.n373 3.1505
R4749 VDD.n381 VDD.n380 3.1505
R4750 VDD.n296 VDD.n295 3.1505
R4751 VDD.n295 VDD.n294 3.1505
R4752 VDD.n300 VDD.n298 3.1505
R4753 VDD.n298 VDD.n297 3.1505
R4754 VDD.n304 VDD.n301 3.1505
R4755 VDD.n296 VDD.n293 3.1505
R4756 VDD.n300 VDD.n299 3.1505
R4757 VDD.n304 VDD.n303 3.1505
R4758 VDD.n303 VDD.n302 3.1505
R4759 VDD.n305 VDD.n285 3.1505
R4760 VDD.n285 VDD.n284 3.1505
R4761 VDD VDD.n308 3.1505
R4762 VDD.n308 VDD.n307 3.1505
R4763 VDD.n311 VDD.n283 3.1505
R4764 VDD.n283 VDD.n282 3.1505
R4765 VDD.n315 VDD.n313 3.1505
R4766 VDD.n313 VDD.n312 3.1505
R4767 VDD.n319 VDD.n316 3.1505
R4768 VDD.n323 VDD.n321 3.1505
R4769 VDD.n321 VDD.n320 3.1505
R4770 VDD.n328 VDD.n325 3.1505
R4771 VDD.n309 VDD 3.1505
R4772 VDD.n311 VDD.n310 3.1505
R4773 VDD.n315 VDD.n314 3.1505
R4774 VDD.n319 VDD.n318 3.1505
R4775 VDD.n318 VDD.n317 3.1505
R4776 VDD.n323 VDD.n322 3.1505
R4777 VDD.n42 VDD.n32 3.1505
R4778 VDD.n32 VDD.n31 3.1505
R4779 VDD.n41 VDD.n40 3.1505
R4780 VDD.n40 VDD.n39 3.1505
R4781 VDD.n38 VDD.n37 3.1505
R4782 VDD.n37 VDD.n36 3.1505
R4783 VDD.n35 VDD.n34 3.1505
R4784 VDD.n8 VDD.n7 3.1505
R4785 VDD.n47 VDD.n46 3.1505
R4786 VDD.n46 VDD.n45 3.1505
R4787 VDD.n44 VDD 3.1505
R4788 VDD.n44 VDD.n43 3.1505
R4789 VDD.n9 VDD.n8 3.14819
R4790 VDD.n1376 VDD.n1373 3.06224
R4791 VDD.n1363 VDD.n1360 3.06224
R4792 VDD.n1023 VDD.n1022 3.06224
R4793 VDD.n472 VDD.n471 3.06224
R4794 VDD.n516 VDD.n513 3.06224
R4795 VDD.n450 VDD.n449 3.06224
R4796 VDD.n169 VDD.n168 3.06224
R4797 VDD.n100 VDD.n97 3.06224
R4798 VDD.n360 VDD.n357 3.06224
R4799 VDD.n275 VDD.n272 3.06224
R4800 VDD.n280 VDD.n279 3.06224
R4801 VDD.n29 VDD.n26 3.06224
R4802 VDD.n1182 VDD.t0 2.91474
R4803 VDD.n1296 VDD.t16 2.91474
R4804 VDD.n122 VDD.n120 2.87637
R4805 VDD.n111 VDD.n109 2.87637
R4806 VDD.n242 VDD.n241 2.87637
R4807 VDD.n237 VDD.n236 2.87637
R4808 VDD.n1559 VDD.n1558 2.6005
R4809 VDD.n1279 VDD.n1278 2.6005
R4810 VDD.n1282 VDD.n1281 2.6005
R4811 VDD.n1307 VDD.n1304 2.6005
R4812 VDD.n1313 VDD.n1310 2.6005
R4813 VDD.n1376 VDD.n1375 2.6005
R4814 VDD.n1363 VDD.n1362 2.6005
R4815 VDD.n1023 VDD.n1020 2.6005
R4816 VDD.n472 VDD.n469 2.6005
R4817 VDD.n516 VDD.n515 2.6005
R4818 VDD.n741 VDD.n740 2.6005
R4819 VDD.n735 VDD.n734 2.6005
R4820 VDD.n833 VDD.n832 2.6005
R4821 VDD.n829 VDD.n828 2.6005
R4822 VDD.n547 VDD.n546 2.6005
R4823 VDD.n563 VDD.n562 2.6005
R4824 VDD.n567 VDD.n566 2.6005
R4825 VDD.n570 VDD.n569 2.6005
R4826 VDD.n555 VDD.n554 2.6005
R4827 VDD.n552 VDD.n551 2.6005
R4828 VDD.n536 VDD.n535 2.6005
R4829 VDD.n539 VDD.n538 2.6005
R4830 VDD.n527 VDD.n526 2.6005
R4831 VDD.n524 VDD.n523 2.6005
R4832 VDD.n531 VDD.n530 2.6005
R4833 VDD.n544 VDD.n543 2.6005
R4834 VDD.n560 VDD.n559 2.6005
R4835 VDD.n574 VDD.n573 2.6005
R4836 VDD.n450 VDD.n447 2.6005
R4837 VDD.n1252 VDD.n1251 2.6005
R4838 VDD.n1249 VDD.n1248 2.6005
R4839 VDD.n1256 VDD.n1255 2.6005
R4840 VDD.n1551 VDD.n1550 2.6005
R4841 VDD.n1554 VDD.n1553 2.6005
R4842 VDD.n1267 VDD.n1266 2.6005
R4843 VDD.n1264 VDD.n1263 2.6005
R4844 VDD.n428 VDD.n426 2.6005
R4845 VDD.n1273 VDD.n1272 2.6005
R4846 VDD.n1270 VDD.n1269 2.6005
R4847 VDD.n424 VDD.n422 2.6005
R4848 VDD.n1546 VDD.n1545 2.6005
R4849 VDD.n420 VDD.n419 2.6005
R4850 VDD.n169 VDD.n166 2.6005
R4851 VDD.n100 VDD.n99 2.6005
R4852 VDD.n360 VDD.n359 2.6005
R4853 VDD.n275 VDD.n274 2.6005
R4854 VDD.n280 VDD.n277 2.6005
R4855 VDD.n29 VDD.n28 2.6005
R4856 VDD.n1437 VDD.n1436 2.59264
R4857 VDD.n1443 VDD.n1442 2.59264
R4858 VDD.n1449 VDD.n1448 2.59264
R4859 VDD.n1455 VDD.n1454 2.59264
R4860 VDD.n1461 VDD.n1460 2.59264
R4861 VDD.n437 VDD.n436 2.59264
R4862 VDD.n972 VDD.n971 2.59264
R4863 VDD.n978 VDD.n977 2.59264
R4864 VDD.n984 VDD.n983 2.59264
R4865 VDD.n990 VDD.n989 2.59264
R4866 VDD.n608 VDD.n607 2.58448
R4867 VDD.n1440 VDD.n1439 2.5167
R4868 VDD.n1446 VDD.n1445 2.5167
R4869 VDD.n1452 VDD.n1451 2.5167
R4870 VDD.n1458 VDD.n1457 2.5167
R4871 VDD.n434 VDD.n433 2.5167
R4872 VDD.n975 VDD.n974 2.5167
R4873 VDD.n981 VDD.n980 2.5167
R4874 VDD.n987 VDD.n986 2.5167
R4875 VDD.n993 VDD.n992 2.5167
R4876 VDD.n651 VDD.t103 2.49842
R4877 VDD.n607 VDD.n606 2.49842
R4878 VDD.n1464 VDD.n1463 2.47755
R4879 VDD.n969 VDD.n968 2.47755
R4880 VDD.n339 VDD.n338 2.31932
R4881 VDD.n128 VDD.n127 2.29638
R4882 VDD.n128 VDD.n125 2.29115
R4883 VDD.n134 VDD.n133 2.2804
R4884 VDD.n502 VDD.n501 2.25904
R4885 VDD.n143 VDD.n142 2.2505
R4886 VDD.n220 VDD.n210 2.2505
R4887 VDD.n334 VDD.n333 2.2505
R4888 VDD.n255 VDD.n254 2.2505
R4889 VDD.n120 VDD.t90 2.16717
R4890 VDD.n120 VDD.n119 2.16717
R4891 VDD.n109 VDD.t347 2.16717
R4892 VDD.n109 VDD.n108 2.16717
R4893 VDD.n241 VDD.t133 2.16717
R4894 VDD.n241 VDD.n240 2.16717
R4895 VDD.n236 VDD.t415 2.16717
R4896 VDD.n236 VDD.n235 2.16717
R4897 VDD.n186 VDD.t320 2.05248
R4898 VDD.n101 VDD.t180 2.05248
R4899 VDD.n284 VDD.t48 2.05248
R4900 VDD.n775 VDD.n774 2.04615
R4901 VDD.n637 VDD.n636 2.00555
R4902 VDD.n1324 VDD.n1323 1.94746
R4903 VDD.n768 VDD.n767 1.94734
R4904 VDD.n132 VDD.n128 1.94241
R4905 VDD.n1006 VDD.n1005 1.8985
R4906 VDD.n1356 VDD.n1355 1.87282
R4907 VDD.n933 VDD.n932 1.87228
R4908 VDD.n145 VDD.n144 1.85344
R4909 VDD.n146 VDD.n145 1.85344
R4910 VDD.n327 VDD.n326 1.85344
R4911 VDD.n328 VDD.n327 1.85344
R4912 VDD.n1337 VDD.n1336 1.83513
R4913 VDD.n756 VDD.n755 1.835
R4914 VDD.n1342 VDD.n1341 1.82925
R4915 VDD.n113 VDD 1.82452
R4916 VDD.n1025 VDD.n461 1.80965
R4917 VDD.n461 VDD.n460 1.80912
R4918 VDD.n195 VDD.n194 1.7505
R4919 VDD.n1351 VDD.n1350 1.69252
R4920 VDD.n1330 VDD.n1329 1.69252
R4921 VDD.n1106 VDD.n1105 1.69252
R4922 VDD.n762 VDD.n761 1.69238
R4923 VDD.n783 VDD.n781 1.69238
R4924 VDD.n1214 VDD.n1213 1.65963
R4925 VDD.n1220 VDD.n1219 1.65963
R4926 VDD.n1225 VDD.n1224 1.65963
R4927 VDD.n1231 VDD.n1230 1.65963
R4928 VDD.n1236 VDD.n1235 1.65963
R4929 VDD.n1244 VDD.n1243 1.65963
R4930 VDD.n23 VDD.n21 1.5755
R4931 VDD.n440 VDD.n439 1.54574
R4932 VDD.n813 VDD.n812 1.54559
R4933 VDD.n964 VDD.n963 1.52056
R4934 VDD.n1000 VDD.n999 1.52056
R4935 VDD.n1468 VDD.n1467 1.52041
R4936 VDD.n996 VDD.n995 1.52041
R4937 VDD.n61 VDD.n58 1.5005
R4938 VDD.n869 VDD.n834 1.49724
R4939 VDD.n1560 VDD.n1543 1.49724
R4940 VDD.n8 VDD.n4 1.488
R4941 VDD.n405 VDD.n401 1.42211
R4942 VDD.n392 VDD.n391 1.42018
R4943 VDD.n825 VDD.n824 1.3744
R4944 VDD.n745 VDD.n744 1.3744
R4945 VDD.n1202 VDD.n1201 1.36284
R4946 VDD.n1003 VDD.n1001 1.35142
R4947 VDD.t199 VDD.t225 1.24946
R4948 VDD.t245 VDD.t211 1.24946
R4949 VDD.n390 VDD.n385 1.2474
R4950 VDD.n412 VDD.n411 1.14837
R4951 VDD.n999 VDD.n998 1.08825
R4952 VDD.n1467 VDD.n1466 1.08806
R4953 VDD.n1275 VDD.n1274 1.06485
R4954 VDD.n183 VDD.n181 1.0505
R4955 VDD.n380 VDD.n378 1.0505
R4956 VDD.n869 VDD.n868 1.01789
R4957 VDD.n1543 VDD.n1283 1.01789
R4958 VDD.n1073 VDD.n1072 0.984049
R4959 VDD.n183 VDD.n95 0.963
R4960 VDD.n394 VDD.n392 0.950899
R4961 VDD.n1597 VDD.n1596 0.931466
R4962 VDD.n224 VDD.n223 0.927241
R4963 VDD.n409 VDD.n408 0.92659
R4964 VDD.n229 VDD.n221 0.904541
R4965 VDD.n340 VDD.n339 0.899617
R4966 VDD.n133 VDD.n132 0.898206
R4967 VDD.n394 VDD.n393 0.897926
R4968 VDD.n400 VDD.n255 0.897926
R4969 VDD.t202 VDD.t193 0.833139
R4970 VDD.t193 VDD.t220 0.833139
R4971 VDD.t187 VDD.t236 0.833139
R4972 VDD.t190 VDD.t187 0.833139
R4973 VDD.t196 VDD.t208 0.833139
R4974 VDD.n412 VDD 0.830218
R4975 VDD.n570 VDD.n567 0.802674
R4976 VDD.n555 VDD.n552 0.802674
R4977 VDD.n539 VDD.n536 0.802674
R4978 VDD.n527 VDD.n524 0.802674
R4979 VDD.n1252 VDD.n1249 0.802674
R4980 VDD.n1554 VDD.n1551 0.802674
R4981 VDD.n1267 VDD.n1264 0.802674
R4982 VDD.n1273 VDD.n1270 0.802674
R4983 VDD.n1470 VDD.n1433 0.795217
R4984 VDD.n401 VDD.n400 0.792748
R4985 VDD.n1242 VDD.n1241 0.746686
R4986 VDD.n1243 VDD.n1242 0.746686
R4987 VDD.n1350 VDD.n1349 0.730547
R4988 VDD.n781 VDD.n780 0.73031
R4989 VDD.n123 VDD.n122 0.7187
R4990 VDD.n1040 VDD.n461 0.674731
R4991 VDD.n780 VDD.n779 0.661938
R4992 VDD.n112 VDD.n111 0.6395
R4993 VDD.n244 VDD.n242 0.6395
R4994 VDD.n239 VDD.n237 0.6395
R4995 VDD.n88 VDD.n86 0.613
R4996 VDD.n965 VDD.n962 0.593699
R4997 VDD.n705 VDD.n531 0.581587
R4998 VDD.n692 VDD.n544 0.581587
R4999 VDD.n670 VDD.n560 0.581587
R5000 VDD.n657 VDD.n574 0.581587
R5001 VDD.n1130 VDD.n428 0.581587
R5002 VDD.n1143 VDD.n424 0.581587
R5003 VDD.n1178 VDD.n420 0.581587
R5004 VDD.n636 VDD.n635 0.573727
R5005 VDD.n1007 VDD.n1006 0.569476
R5006 VDD.n1349 VDD.n1348 0.553668
R5007 VDD.n401 VDD.n229 0.539532
R5008 VDD.n1344 VDD.n1307 0.536587
R5009 VDD.n1332 VDD.n1313 0.536587
R5010 VDD.n1320 VDD.n1315 0.536587
R5011 VDD.n747 VDD.n741 0.536587
R5012 VDD.n758 VDD.n735 0.536587
R5013 VDD.n770 VDD.n729 0.536587
R5014 VDD.n8 VDD.n6 0.5255
R5015 VDD.n814 VDD.n811 0.495796
R5016 VDD VDD.n100 0.485717
R5017 VDD VDD.n169 0.485717
R5018 VDD VDD.n1023 0.474784
R5019 VDD.n1560 VDD.n1559 0.467817
R5020 VDD.n1283 VDD.n1282 0.466777
R5021 VDD.n830 VDD.n829 0.466777
R5022 VDD.n391 VDD.n390 0.462817
R5023 VDD.n571 VDD.n570 0.440717
R5024 VDD.n1249 VDD.n1246 0.440717
R5025 VDD.n1543 VDD.n1279 0.430935
R5026 VDD.n834 VDD.n833 0.430935
R5027 VDD.n1257 VDD.n1256 0.430935
R5028 VDD.n567 VDD.n564 0.421152
R5029 VDD.n1253 VDD.n1252 0.421152
R5030 VDD.n1124 VDD.t10 0.41682
R5031 VDD.t330 VDD.t217 0.41682
R5032 VDD.t250 VDD.t330 0.41682
R5033 VDD.t205 VDD.t233 0.41682
R5034 VDD.t214 VDD.t325 0.41682
R5035 VDD.t325 VDD.t228 0.41682
R5036 VDD.n787 VDD.n785 0.405977
R5037 VDD.n1108 VDD.n1099 0.405977
R5038 VDD.n905 VDD.n830 0.394968
R5039 VDD.n870 VDD.n869 0.394968
R5040 VDD.n1561 VDD.n1560 0.394968
R5041 VDD.n531 VDD.n528 0.389848
R5042 VDD.n428 VDD.n427 0.389848
R5043 VDD.n1382 VDD.n1380 0.389323
R5044 VDD.n1030 VDD.n1028 0.389323
R5045 VDD.n35 VDD.n33 0.389323
R5046 VDD.n1406 VDD.n1368 0.376152
R5047 VDD.n501 VDD.n467 0.376152
R5048 VDD.n502 VDD.n464 0.376152
R5049 VDD.n1049 VDD.n455 0.376152
R5050 VDD.n137 VDD.n103 0.376152
R5051 VDD.n80 VDD.n74 0.376152
R5052 VDD.n383 VDD.n342 0.376152
R5053 VDD.n292 VDD.n288 0.376152
R5054 VDD.n292 VDD.n291 0.376152
R5055 VDD.n1377 VDD.n1376 0.374196
R5056 VDD.n1364 VDD.n1363 0.374196
R5057 VDD.n473 VDD.n472 0.374196
R5058 VDD.n451 VDD.n450 0.374196
R5059 VDD.n361 VDD.n360 0.374196
R5060 VDD.n281 VDD.n275 0.374196
R5061 VDD.n281 VDD.n280 0.374196
R5062 VDD.n30 VDD.n29 0.374196
R5063 VDD.n1040 VDD.n1018 0.372931
R5064 VDD.n1470 VDD.n1469 0.359918
R5065 VDD.n1574 VDD.n1257 0.358543
R5066 VDD.n892 VDD.n834 0.358543
R5067 VDD.n1543 VDD.n1542 0.358543
R5068 VDD.n4 VDD.n3 0.350287
R5069 VDD.n556 VDD.n555 0.327239
R5070 VDD.n1551 VDD.n1548 0.327239
R5071 VDD.n540 VDD.n539 0.323326
R5072 VDD.n528 VDD.n527 0.323326
R5073 VDD.n1264 VDD.n1261 0.323326
R5074 VDD.n1406 VDD.n1405 0.312794
R5075 VDD.n1279 VDD.n1276 0.311587
R5076 VDD.n1049 VDD.n1048 0.306039
R5077 VDD.n1238 VDD.n413 0.292144
R5078 VDD.n1227 VDD.n414 0.292144
R5079 VDD.n1218 VDD.n415 0.292144
R5080 VDD.n1559 VDD.n1556 0.292022
R5081 VDD.n548 VDD.n547 0.292022
R5082 VDD.n564 VDD.n563 0.292022
R5083 VDD.n536 VDD.n533 0.292022
R5084 VDD.n524 VDD.n521 0.292022
R5085 VDD.n1256 VDD.n1253 0.292022
R5086 VDD.n1275 VDD.n1267 0.292022
R5087 VDD.n1274 VDD.n1273 0.292022
R5088 VDD.n586 VDD.n579 0.291683
R5089 VDD.n599 VDD.n578 0.291683
R5090 VDD.n611 VDD.n577 0.291683
R5091 VDD.n1208 VDD.n416 0.288544
R5092 VDD.n624 VDD.n576 0.288083
R5093 VDD.n552 VDD.n549 0.278326
R5094 VDD.n1555 VDD.n1554 0.278326
R5095 VDD.n560 VDD.n557 0.272457
R5096 VDD.n574 VDD.n571 0.272457
R5097 VDD.n1547 VDD.n1546 0.272457
R5098 VDD.n544 VDD.n541 0.266587
R5099 VDD.n424 VDD.n423 0.266587
R5100 VDD.n773 VDD.n726 0.266523
R5101 VDD.n1317 VDD.n1316 0.26536
R5102 VDD.n743 VDD.n742 0.264528
R5103 VDD.n1347 VDD.n1302 0.263373
R5104 VDD.n195 VDD.n191 0.263
R5105 VDD.n764 VDD.n730 0.262011
R5106 VDD.n1326 VDD.n1314 0.260887
R5107 VDD.n754 VDD.n736 0.257984
R5108 VDD.n1335 VDD.n1308 0.257526
R5109 VDD.n954 VDD.n817 0.25389
R5110 VDD.n9 VDD.n2 0.253803
R5111 VDD.n1596 VDD.n1595 0.252505
R5112 VDD.n1075 VDD.n1073 0.248505
R5113 VDD.n942 VDD.n818 0.238241
R5114 VDD.n1479 VDD.n1358 0.238069
R5115 VDD.n1491 VDD.n1357 0.237294
R5116 VDD.n475 VDD.n474 0.237044
R5117 VDD.n445 VDD.n444 0.237044
R5118 VDD.n346 VDD.n345 0.237044
R5119 VDD.n79 VDD.n77 0.233429
R5120 VDD.n1405 VDD.n1371 0.229786
R5121 VDD.n1048 VDD.n458 0.229786
R5122 VDD.n134 VDD.n105 0.229786
R5123 VDD.n330 VDD.n270 0.229786
R5124 VDD.n1082 VDD.n432 0.221442
R5125 VDD.n803 VDD.n517 0.220495
R5126 VDD.n392 VDD.n340 0.217222
R5127 VDD.n638 VDD.n634 0.209826
R5128 VDD.n1200 VDD.n1199 0.209826
R5129 VDD.n581 VDD.n580 0.183919
R5130 VDD.n348 VDD.n347 0.182274
R5131 VDD.n1402 VDD.n1401 0.182033
R5132 VDD.n1427 VDD.n1426 0.182033
R5133 VDD.n477 VDD.n476 0.182033
R5134 VDD.n1045 VDD.n1044 0.182033
R5135 VDD.n1070 VDD.n1069 0.182033
R5136 VDD.n1097 VDD.n429 0.17667
R5137 VDD.n1500 VDD.n1498 0.176655
R5138 VDD.n937 VDD.n934 0.176655
R5139 VDD.n1433 VDD.n1429 0.174122
R5140 VDD.n725 VDD.n722 0.17241
R5141 VDD.n1114 VDD.n1111 0.17241
R5142 VDD.n927 VDD.n923 0.171399
R5143 VDD.n1513 VDD.n1510 0.171399
R5144 VDD.n769 VDD.n766 0.163357
R5145 VDD.n1325 VDD.n1322 0.163357
R5146 VDD.n923 VDD.n920 0.157434
R5147 VDD.n1516 VDD.n1513 0.15672
R5148 VDD.n644 VDD.n641 0.153197
R5149 VDD.n1196 VDD.n1193 0.153197
R5150 VDD.n839 VDD.n836 0.146319
R5151 VDD.n776 VDD.n773 0.146214
R5152 VDD.n641 VDD.n638 0.146118
R5153 VDD.n1199 VDD.n1196 0.146118
R5154 VDD.n1595 VDD.n1592 0.146022
R5155 VDD.n1505 VDD.n1501 0.143084
R5156 VDD.n772 VDD.n770 0.143
R5157 VDD.n1111 VDD.n1108 0.142944
R5158 VDD.n785 VDD.n725 0.142944
R5159 VDD.n520 VDD.n519 0.142202
R5160 VDD.n931 VDD.n929 0.142073
R5161 VDD.n1320 VDD.n1319 0.141929
R5162 VDD.n1501 VDD.n1500 0.141062
R5163 VDD.n934 VDD.n931 0.141062
R5164 VDD.n753 VDD.n751 0.140857
R5165 VDD.n1340 VDD.n1338 0.140857
R5166 VDD.n634 VDD.n633 0.14038
R5167 VDD.n1203 VDD.n1200 0.14038
R5168 VDD.n751 VDD.n749 0.139786
R5169 VDD.n778 VDD.n776 0.139786
R5170 VDD.n1103 VDD.n1101 0.139786
R5171 VDD.n1343 VDD.n1340 0.139786
R5172 VDD VDD.n123 0.139763
R5173 VDD.n1073 VDD.n441 0.139295
R5174 VDD.n441 VDD.n438 0.138211
R5175 VDD.n816 VDD.n814 0.138211
R5176 VDD.n757 VDD.n754 0.137643
R5177 VDD.n1335 VDD.n1334 0.137643
R5178 VDD.n722 VDD.n719 0.137017
R5179 VDD.n1117 VDD.n1114 0.136006
R5180 VDD.n438 VDD.n435 0.133873
R5181 VDD.n1438 VDD.n1435 0.133873
R5182 VDD.n1444 VDD.n1441 0.133873
R5183 VDD.n1450 VDD.n1447 0.133873
R5184 VDD.n1456 VDD.n1453 0.133873
R5185 VDD.n1462 VDD.n1459 0.133873
R5186 VDD.n1469 VDD.n1465 0.133873
R5187 VDD.n967 VDD.n965 0.133873
R5188 VDD.n973 VDD.n970 0.133873
R5189 VDD.n979 VDD.n976 0.133873
R5190 VDD.n985 VDD.n982 0.133873
R5191 VDD.n991 VDD.n988 0.133873
R5192 VDD.n997 VDD.n994 0.133873
R5193 VDD.n1498 VDD.n1495 0.133833
R5194 VDD.n1490 VDD.n1487 0.133833
R5195 VDD.n1487 VDD.n1483 0.133833
R5196 VDD.n1478 VDD.n1475 0.133833
R5197 VDD.n960 VDD.n957 0.133833
R5198 VDD.n953 VDD.n949 0.133833
R5199 VDD.n949 VDD.n945 0.133833
R5200 VDD.n941 VDD.n937 0.133833
R5201 VDD.n821 VDD.n819 0.133132
R5202 VDD VDD.n177 0.131587
R5203 VDD.n1093 VDD.n431 0.131498
R5204 VDD.n792 VDD.n520 0.13055
R5205 VDD.n1334 VDD.n1332 0.130143
R5206 VDD.n174 VDD 0.12963
R5207 VDD.n585 VDD.n582 0.129536
R5208 VDD.n592 VDD.n589 0.129536
R5209 VDD.n595 VDD.n592 0.129536
R5210 VDD.n598 VDD.n595 0.129536
R5211 VDD.n605 VDD.n602 0.129536
R5212 VDD.n610 VDD.n605 0.129536
R5213 VDD.n617 VDD.n614 0.129536
R5214 VDD.n620 VDD.n617 0.129536
R5215 VDD.n623 VDD.n620 0.129536
R5216 VDD.n630 VDD.n627 0.129536
R5217 VDD.n633 VDD.n630 0.129536
R5218 VDD.n1205 VDD.n1203 0.129536
R5219 VDD.n1207 VDD.n1205 0.129536
R5220 VDD.n1212 VDD.n1210 0.129536
R5221 VDD.n1215 VDD.n1212 0.129536
R5222 VDD.n1217 VDD.n1215 0.129536
R5223 VDD.n1223 VDD.n1221 0.129536
R5224 VDD.n1226 VDD.n1223 0.129536
R5225 VDD.n1232 VDD.n1229 0.129536
R5226 VDD.n1234 VDD.n1232 0.129536
R5227 VDD.n1237 VDD.n1234 0.129536
R5228 VDD.n1245 VDD.n1240 0.129536
R5229 VDD.n380 VDD.n379 0.129141
R5230 VDD.n758 VDD.n757 0.129071
R5231 VDD.n520 VDD.n518 0.128395
R5232 VDD.n431 VDD.n430 0.128395
R5233 VDD.n1441 VDD.n1438 0.127367
R5234 VDD.n1447 VDD.n1444 0.127367
R5235 VDD.n1453 VDD.n1450 0.127367
R5236 VDD.n1459 VDD.n1456 0.127367
R5237 VDD.n586 VDD.n585 0.127367
R5238 VDD.n976 VDD.n973 0.127367
R5239 VDD.n982 VDD.n979 0.127367
R5240 VDD.n988 VDD.n985 0.127367
R5241 VDD.n994 VDD.n991 0.127367
R5242 VDD.n1240 VDD.n1238 0.127367
R5243 VDD.n333 VDD.n332 0.126143
R5244 VDD.n1465 VDD.n1462 0.124114
R5245 VDD.n970 VDD.n967 0.124114
R5246 VDD.n811 VDD.n809 0.123227
R5247 VDD.n809 VDD.n806 0.123227
R5248 VDD.n802 VDD.n799 0.123227
R5249 VDD.n799 VDD.n795 0.123227
R5250 VDD.n1092 VDD.n1089 0.123227
R5251 VDD.n1089 VDD.n1085 0.123227
R5252 VDD.n1081 VDD.n1078 0.123227
R5253 VDD.n1078 VDD.n1075 0.123227
R5254 VDD.n611 VDD.n610 0.12303
R5255 VDD.n1221 VDD.n1218 0.12303
R5256 VDD.n803 VDD.n802 0.122205
R5257 VDD.n1085 VDD.n1082 0.122205
R5258 VDD.n719 VDD.n716 0.120837
R5259 VDD.n716 VDD.n713 0.120837
R5260 VDD.n713 VDD.n710 0.120837
R5261 VDD.n710 VDD.n708 0.120837
R5262 VDD.n704 VDD.n701 0.120837
R5263 VDD.n701 VDD.n698 0.120837
R5264 VDD.n698 VDD.n695 0.120837
R5265 VDD.n691 VDD.n688 0.120837
R5266 VDD.n688 VDD.n685 0.120837
R5267 VDD.n685 VDD.n682 0.120837
R5268 VDD.n682 VDD.n679 0.120837
R5269 VDD.n679 VDD.n676 0.120837
R5270 VDD.n676 VDD.n673 0.120837
R5271 VDD.n669 VDD.n666 0.120837
R5272 VDD.n666 VDD.n663 0.120837
R5273 VDD.n663 VDD.n660 0.120837
R5274 VDD.n656 VDD.n653 0.120837
R5275 VDD.n653 VDD.n650 0.120837
R5276 VDD.n650 VDD.n647 0.120837
R5277 VDD.n647 VDD.n644 0.120837
R5278 VDD.n1193 VDD.n1190 0.120837
R5279 VDD.n1190 VDD.n1187 0.120837
R5280 VDD.n1187 VDD.n1184 0.120837
R5281 VDD.n1184 VDD.n1181 0.120837
R5282 VDD.n1177 VDD.n1174 0.120837
R5283 VDD.n1174 VDD.n1171 0.120837
R5284 VDD.n1171 VDD.n1168 0.120837
R5285 VDD.n1164 VDD.n1161 0.120837
R5286 VDD.n1161 VDD.n1158 0.120837
R5287 VDD.n1158 VDD.n1155 0.120837
R5288 VDD.n1155 VDD.n1152 0.120837
R5289 VDD.n1152 VDD.n1149 0.120837
R5290 VDD.n1149 VDD.n1146 0.120837
R5291 VDD.n1142 VDD.n1139 0.120837
R5292 VDD.n1139 VDD.n1136 0.120837
R5293 VDD.n1136 VDD.n1133 0.120837
R5294 VDD.n1129 VDD.n1126 0.120837
R5295 VDD.n1126 VDD.n1123 0.120837
R5296 VDD.n1123 VDD.n1120 0.120837
R5297 VDD.n1120 VDD.n1117 0.120837
R5298 VDD.n1472 VDD.n1470 0.119037
R5299 VDD.n826 VDD.n823 0.117286
R5300 VDD.n763 VDD.n760 0.117286
R5301 VDD.n784 VDD.n778 0.117286
R5302 VDD.n1107 VDD.n1103 0.117286
R5303 VDD.n1331 VDD.n1328 0.117286
R5304 VDD.n1354 VDD.n1352 0.117286
R5305 VDD.n1096 VDD.n1093 0.113
R5306 VDD.n792 VDD.n791 0.111977
R5307 VDD.n1178 VDD.n1177 0.110725
R5308 VDD.n660 VDD.n657 0.109713
R5309 VDD.n928 VDD.n826 0.108714
R5310 VDD.n1346 VDD.n1344 0.107643
R5311 VDD.n1506 VDD.n1354 0.107643
R5312 VDD.n390 VDD.n389 0.106797
R5313 VDD.n747 VDD.n746 0.106571
R5314 VDD.n705 VDD.n704 0.103646
R5315 VDD.n1133 VDD.n1130 0.102635
R5316 VDD.n408 VDD.n407 0.101088
R5317 VDD.n842 VDD.n839 0.1005
R5318 VDD.n1592 VDD.n1589 0.1005
R5319 VDD.n1495 VDD.n1491 0.0971667
R5320 VDD.n942 VDD.n941 0.0971667
R5321 VDD.n1352 VDD.n1347 0.0947857
R5322 VDD.n1506 VDD.n1505 0.0945449
R5323 VDD.n1475 VDD.n1472 0.0938198
R5324 VDD.n962 VDD.n960 0.0938198
R5325 VDD.n929 VDD.n928 0.0935337
R5326 VDD.n117 VDD.n112 0.0893158
R5327 VDD.n245 VDD.n239 0.0893158
R5328 VDD.n245 VDD.n244 0.0893158
R5329 VDD.n1099 VDD.n1097 0.0884545
R5330 VDD.n1143 VDD.n1142 0.0874663
R5331 VDD.n788 VDD.n787 0.0874318
R5332 VDD.n695 VDD.n692 0.0864551
R5333 VDD.n1483 VDD.n1479 0.0860556
R5334 VDD.n954 VDD.n953 0.0860556
R5335 VDD.n920 VDD.n917 0.0855
R5336 VDD.n917 VDD.n914 0.0855
R5337 VDD.n914 VDD.n911 0.0855
R5338 VDD.n911 VDD.n908 0.0855
R5339 VDD.n904 VDD.n901 0.0855
R5340 VDD.n901 VDD.n898 0.0855
R5341 VDD.n898 VDD.n895 0.0855
R5342 VDD.n891 VDD.n888 0.0855
R5343 VDD.n888 VDD.n885 0.0855
R5344 VDD.n885 VDD.n882 0.0855
R5345 VDD.n879 VDD.n876 0.0855
R5346 VDD.n876 VDD.n873 0.0855
R5347 VDD.n867 VDD.n864 0.0855
R5348 VDD.n864 VDD.n861 0.0855
R5349 VDD.n861 VDD.n858 0.0855
R5350 VDD.n854 VDD.n851 0.0855
R5351 VDD.n851 VDD.n848 0.0855
R5352 VDD.n848 VDD.n845 0.0855
R5353 VDD.n845 VDD.n842 0.0855
R5354 VDD.n1528 VDD.n1525 0.0855
R5355 VDD.n1525 VDD.n1522 0.0855
R5356 VDD.n1522 VDD.n1519 0.0855
R5357 VDD.n1519 VDD.n1516 0.0855
R5358 VDD.n1589 VDD.n1586 0.0855
R5359 VDD.n1586 VDD.n1583 0.0855
R5360 VDD.n1583 VDD.n1580 0.0855
R5361 VDD.n1580 VDD.n1577 0.0855
R5362 VDD.n1573 VDD.n1570 0.0855
R5363 VDD.n1570 VDD.n1567 0.0855
R5364 VDD.n1567 VDD.n1564 0.0855
R5365 VDD.n1286 VDD.n1260 0.0855
R5366 VDD.n1289 VDD.n1286 0.0855
R5367 VDD.n1295 VDD.n1292 0.0855
R5368 VDD.n1298 VDD.n1295 0.0855
R5369 VDD.n1301 VDD.n1298 0.0855
R5370 VDD.n1541 VDD.n1538 0.0855
R5371 VDD.n1538 VDD.n1535 0.0855
R5372 VDD.n1535 VDD.n1532 0.0855
R5373 VDD.n627 VDD.n624 0.0850783
R5374 VDD.n1208 VDD.n1207 0.0850783
R5375 VDD.n1574 VDD.n1573 0.0847857
R5376 VDD.n858 VDD.n855 0.0840714
R5377 VDD.n116 VDD 0.0836933
R5378 VDD.n1001 VDD.n997 0.0818253
R5379 VDD.n670 VDD.n669 0.0803876
R5380 VDD.n1168 VDD.n1165 0.0793764
R5381 VDD.n231 VDD.n230 0.0790106
R5382 VDD.n246 VDD 0.0774922
R5383 VDD.n928 VDD.n927 0.0773539
R5384 VDD.n1510 VDD.n1506 0.0773539
R5385 VDD.n766 VDD.n764 0.0765714
R5386 VDD.n1326 VDD.n1325 0.0765714
R5387 VDD.n1474 VDD.n1473 0.074985
R5388 VDD.n959 VDD.n958 0.074985
R5389 VDD.n602 VDD.n599 0.0742349
R5390 VDD.n1227 VDD.n1226 0.0742349
R5391 VDD.n338 VDD.n337 0.07388
R5392 VDD.n1001 VDD.n816 0.0731506
R5393 VDD.n131 VDD.n130 0.0717174
R5394 VDD.n1388 VDD.n1385 0.0714756
R5395 VDD.n1413 VDD.n1410 0.0714756
R5396 VDD.n1036 VDD.n1033 0.0714756
R5397 VDD.n498 VDD.n495 0.0714756
R5398 VDD.n510 VDD.n507 0.0714756
R5399 VDD.n1011 VDD.n1010 0.0714756
R5400 VDD.n1056 VDD.n1053 0.0714756
R5401 VDD.n375 VDD.n372 0.0714756
R5402 VDD.n41 VDD.n38 0.0714756
R5403 VDD.n396 VDD.n395 0.0714615
R5404 VDD VDD.n1389 0.0713871
R5405 VDD VDD.n1414 0.0713871
R5406 VDD.n492 VDD 0.0713871
R5407 VDD VDD.n1057 0.0713871
R5408 VDD.n369 VDD 0.0713871
R5409 VDD VDD.n42 0.0713871
R5410 VDD.n1403 VDD.n1400 0.0709032
R5411 VDD.n1397 VDD.n1394 0.0709032
R5412 VDD.n1428 VDD.n1425 0.0709032
R5413 VDD.n1422 VDD.n1419 0.0709032
R5414 VDD.n485 VDD.n484 0.0709032
R5415 VDD.n481 VDD.n478 0.0709032
R5416 VDD.n1046 VDD.n1043 0.0709032
R5417 VDD.n1071 VDD.n1068 0.0709032
R5418 VDD.n1065 VDD.n1062 0.0709032
R5419 VDD.n352 VDD.n349 0.0709032
R5420 VDD.n362 VDD.n355 0.0709032
R5421 VDD.n50 VDD.n47 0.0701774
R5422 VDD.n1389 VDD.n1388 0.0692805
R5423 VDD.n1385 VDD.n1382 0.0692805
R5424 VDD.n1414 VDD.n1413 0.0692805
R5425 VDD.n1410 VDD.n1407 0.0692805
R5426 VDD.n1039 VDD.n1036 0.0692805
R5427 VDD.n1033 VDD.n1030 0.0692805
R5428 VDD.n500 VDD.n498 0.0692805
R5429 VDD.n495 VDD.n492 0.0692805
R5430 VDD.n507 VDD.n504 0.0692805
R5431 VDD.n511 VDD.n510 0.0692805
R5432 VDD VDD.n1011 0.0692805
R5433 VDD.n1057 VDD.n1056 0.0692805
R5434 VDD.n1053 VDD.n1050 0.0692805
R5435 VDD.n372 VDD.n369 0.0692805
R5436 VDD.n42 VDD.n41 0.0692805
R5437 VDD.n38 VDD.n35 0.0692805
R5438 VDD.n1404 VDD.n1403 0.0687258
R5439 VDD.n1400 VDD.n1397 0.0687258
R5440 VDD.n1429 VDD.n1428 0.0687258
R5441 VDD.n1425 VDD.n1422 0.0687258
R5442 VDD.n484 VDD.n481 0.0687258
R5443 VDD.n478 VDD.n475 0.0687258
R5444 VDD.n1047 VDD.n1046 0.0687258
R5445 VDD.n1068 VDD.n1065 0.0687258
R5446 VDD.n349 VDD.n346 0.0687258
R5447 VDD.n355 VDD.n352 0.0687258
R5448 VDD.n1542 VDD.n1541 0.0683571
R5449 VDD.n895 VDD.n892 0.0676429
R5450 VDD.n213 VDD.n212 0.0669486
R5451 VDD.n225 VDD.n224 0.0669486
R5452 VDD.n1504 VDD.n1502 0.0668158
R5453 VDD.n905 VDD.n904 0.0662143
R5454 VDD.n1532 VDD.n1529 0.0662143
R5455 VDD.n218 VDD.n217 0.0661075
R5456 VDD.n228 VDD.n227 0.0661075
R5457 VDD.n117 VDD.n116 0.0647857
R5458 VDD.n234 VDD.n233 0.0646489
R5459 VDD.n1394 VDD.n1377 0.0629194
R5460 VDD.n1419 VDD.n1364 0.0629194
R5461 VDD.n485 VDD.n473 0.0629194
R5462 VDD.n1062 VDD.n451 0.0629194
R5463 VDD.n362 VDD.n361 0.0629194
R5464 VDD.n47 VDD.n30 0.0629194
R5465 VDD.n246 VDD.n245 0.0606172
R5466 VDD.n1040 VDD.n1039 0.0605
R5467 VDD.n376 VDD.n375 0.0605
R5468 VDD.n399 VDD.n398 0.0584808
R5469 VDD.n599 VDD.n598 0.0558012
R5470 VDD.n1229 VDD.n1227 0.0558012
R5471 VDD.n1018 VDD 0.055378
R5472 VDD.n404 VDD.n403 0.0534412
R5473 VDD.n64 VDD.n63 0.0534412
R5474 VDD.n549 VDD.n548 0.0533261
R5475 VDD.n1556 VDD.n1555 0.0533261
R5476 VDD.n1108 VDD.n1107 0.053
R5477 VDD.n1010 VDD.n1007 0.0524512
R5478 VDD.n785 VDD.n784 0.0519286
R5479 VDD.n125 VDD.n107 0.0509
R5480 VDD.n251 VDD.n250 0.0504219
R5481 VDD.n1043 VDD.n1040 0.0498548
R5482 VDD.n870 VDD.n867 0.0497857
R5483 VDD.n1564 VDD.n1561 0.0497857
R5484 VDD.n882 VDD 0.0483571
R5485 VDD.n1479 VDD.n1478 0.0482778
R5486 VDD.n957 VDD.n954 0.0482778
R5487 VDD.n1292 VDD 0.0462143
R5488 VDD.n624 VDD.n623 0.0449578
R5489 VDD.n1210 VDD.n1208 0.0449578
R5490 VDD.n1165 VDD.n1164 0.0419607
R5491 VDD.n764 VDD.n763 0.0412143
R5492 VDD.n773 VDD.n772 0.0412143
R5493 VDD.n1319 VDD.n1317 0.0412143
R5494 VDD.n1328 VDD.n1326 0.0412143
R5495 VDD.n18 VDD.n15 0.0411452
R5496 VDD.n673 VDD.n670 0.0409494
R5497 VDD.n70 VDD.n69 0.0408043
R5498 VDD VDD.n1289 0.0397857
R5499 VDD.n1596 VDD.n1245 0.0395361
R5500 VDD VDD.n1597 0.0393983
R5501 VDD VDD.n879 0.0376429
R5502 VDD.n1072 VDD.n445 0.0375161
R5503 VDD.n1491 VDD.n1490 0.0371667
R5504 VDD.n945 VDD.n942 0.0371667
R5505 VDD.n1433 VDD.n1432 0.0369005
R5506 VDD.n254 VDD.n253 0.0367109
R5507 VDD.n791 VDD.n788 0.0362955
R5508 VDD.n873 VDD.n870 0.0362143
R5509 VDD.n1561 VDD.n1260 0.0362143
R5510 VDD.n304 VDD.n300 0.0359878
R5511 VDD VDD.n305 0.0359436
R5512 VDD.n315 VDD.n311 0.0357016
R5513 VDD.n323 VDD.n319 0.0357016
R5514 VDD.n1097 VDD.n1096 0.0352727
R5515 VDD.n300 VDD.n296 0.0348902
R5516 VDD.n305 VDD.n304 0.0348902
R5517 VDD.n692 VDD.n691 0.034882
R5518 VDD.n749 VDD.n747 0.0347857
R5519 VDD.n319 VDD.n315 0.0346129
R5520 VDD.n269 VDD.n268 0.0340503
R5521 VDD.n1146 VDD.n1143 0.0338708
R5522 VDD.n541 VDD.n540 0.0337609
R5523 VDD.n1344 VDD.n1343 0.0337143
R5524 VDD.n336 VDD.n335 0.0335178
R5525 VDD.n400 VDD.n399 0.0331389
R5526 VDD.n395 VDD.n394 0.0322736
R5527 VDD.n1072 VDD.n1071 0.0317097
R5528 VDD.n311 VDD.n281 0.0317097
R5529 VDD.n255 VDD.n234 0.0301809
R5530 VDD.n132 VDD.n131 0.0299176
R5531 VDD.n232 VDD.n231 0.0292234
R5532 VDD.n233 VDD.n232 0.0292234
R5533 VDD.n1095 VDD.n1094 0.0291956
R5534 VDD.n808 VDD.n807 0.0291956
R5535 VDD.n790 VDD.n789 0.0291956
R5536 VDD.n1077 VDD.n1076 0.0291956
R5537 VDD.n163 VDD.n162 0.0289211
R5538 VDD.n159 VDD.n156 0.0289211
R5539 VDD.n407 VDD.n406 0.0278529
R5540 VDD.n403 VDD.n402 0.0278529
R5541 VDD.n258 VDD.n257 0.0277596
R5542 VDD.n261 VDD.n260 0.0273269
R5543 VDD.n1003 VDD.n1002 0.0270909
R5544 VDD.n227 VDD.n226 0.0265748
R5545 VDD.n397 VDD.n396 0.0264615
R5546 VDD.n398 VDD.n397 0.0264615
R5547 VDD.n226 VDD.n225 0.0257336
R5548 VDD.n153 VDD.n150 0.0256417
R5549 VDD.n324 VDD.n323 0.0251774
R5550 VDD.n13 VDD.n12 0.0247707
R5551 VDD.n133 VDD.n106 0.0247609
R5552 VDD.n557 VDD.n556 0.0239783
R5553 VDD.n1548 VDD.n1547 0.0239783
R5554 VDD.n130 VDD.n129 0.0239783
R5555 VDD.n266 VDD.n262 0.0235488
R5556 VDD.n174 VDD.n164 0.0234555
R5557 VDD.n406 VDD.n405 0.0234412
R5558 VDD.n746 VDD.n743 0.023
R5559 VDD.n1322 VDD.n1320 0.023
R5560 VDD.n1347 VDD.n1346 0.023
R5561 VDD.n205 VDD.n202 0.0227267
R5562 VDD.n62 VDD.n61 0.0225588
R5563 VDD.n60 VDD.n59 0.0225588
R5564 VDD.n80 VDD.n79 0.0223623
R5565 VDD.n770 VDD.n769 0.0219286
R5566 VDD.n189 VDD.n188 0.0216336
R5567 VDD.n229 VDD.n228 0.0206869
R5568 VDD.n533 VDD.n532 0.0200652
R5569 VDD.n1276 VDD.n1275 0.0200652
R5570 VDD.n139 VDD.n138 0.0200652
R5571 VDD.n142 VDD.n141 0.0200652
R5572 VDD.n219 VDD.n218 0.0198458
R5573 VDD.n908 VDD.n905 0.0197857
R5574 VDD.n1529 VDD.n1528 0.0197857
R5575 VDD.n250 VDD.n249 0.0191328
R5576 VDD.n127 VDD.n126 0.0191207
R5577 VDD.n136 VDD.n135 0.019083
R5578 VDD.n391 VDD.n341 0.0190047
R5579 VDD.n1130 VDD.n1129 0.0187022
R5580 VDD.n58 VDD.n24 0.0186452
R5581 VDD.n57 VDD.n56 0.0186452
R5582 VDD.n892 VDD.n891 0.0183571
R5583 VDD.n708 VDD.n705 0.017691
R5584 VDD.n1542 VDD.n1301 0.0176429
R5585 VDD.n216 VDD.n215 0.0173224
R5586 VDD.n214 VDD.n213 0.0173224
R5587 VDD.n1018 VDD.n511 0.0165976
R5588 VDD.n56 VDD.n53 0.0164677
R5589 VDD.n340 VDD.n261 0.0160453
R5590 VDD.n334 VDD.n269 0.0159438
R5591 VDD.n335 VDD.n334 0.0159438
R5592 VDD.n339 VDD.n336 0.0159438
R5593 VDD.n410 VDD.n409 0.0157992
R5594 VDD.n389 VDD.n388 0.0156402
R5595 VDD.n66 VDD.n65 0.015009
R5596 VDD.n125 VDD.n124 0.0149
R5597 VDD.n123 VDD.n107 0.014
R5598 VDD.n1407 VDD.n1406 0.0136707
R5599 VDD.n501 VDD.n500 0.0136707
R5600 VDD.n504 VDD.n502 0.0136707
R5601 VDD.n1050 VDD.n1049 0.0136707
R5602 VDD.n24 VDD.n19 0.0135645
R5603 VDD.n257 VDD.n256 0.0130481
R5604 VDD.n259 VDD.n258 0.0130481
R5605 VDD.n260 VDD.n259 0.0130481
R5606 VDD.n71 VDD.n70 0.0122391
R5607 VDD.n209 VDD.n208 0.0121599
R5608 VDD.n15 VDD.n14 0.0121129
R5609 VDD.n65 VDD.n64 0.0119706
R5610 VDD.n118 VDD.n117 0.0118445
R5611 VDD.n795 VDD.n792 0.01175
R5612 VDD.n657 VDD.n656 0.0116236
R5613 VDD.n212 VDD.n211 0.0114346
R5614 VDD.n760 VDD.n758 0.0112143
R5615 VDD.n1093 VDD.n1092 0.0107273
R5616 VDD.n1181 VDD.n1178 0.0106124
R5617 VDD.n388 VDD.n387 0.0105935
R5618 VDD.n1332 VDD.n1331 0.0101429
R5619 VDD.n268 VDD.n267 0.0100858
R5620 VDD.n328 VDD.n324 0.00993548
R5621 VDD.n217 VDD.n216 0.00975234
R5622 VDD.n1040 VDD 0.00932353
R5623 VDD.n253 VDD.n251 0.00928906
R5624 VDD.n381 VDD.n376 0.00928049
R5625 VDD.n385 VDD.n384 0.00928049
R5626 VDD.n215 VDD.n214 0.00891121
R5627 VDD.n210 VDD.n92 0.00888057
R5628 VDD.n382 VDD.n381 0.00854878
R5629 VDD.n384 VDD.n383 0.00854878
R5630 VDD.n264 VDD.n263 0.00853674
R5631 VDD.n177 VDD.n176 0.00851619
R5632 VDD.n123 VDD.n118 0.00806303
R5633 VDD.n196 VDD.n189 0.00778745
R5634 VDD.n1405 VDD.n1404 0.00775806
R5635 VDD.n1048 VDD.n1047 0.00775806
R5636 VDD.n68 VDD.n67 0.00754348
R5637 VDD.n164 VDD.n163 0.00742308
R5638 VDD.n156 VDD.n153 0.00742308
R5639 VDD.n208 VDD.n205 0.00742308
R5640 VDD.n14 VDD.n13 0.00738437
R5641 VDD.n296 VDD.n292 0.00708537
R5642 VDD.n83 VDD.n80 0.0070587
R5643 VDD.n175 VDD.n93 0.0070587
R5644 VDD.n614 VDD.n611 0.00700602
R5645 VDD.n1218 VDD.n1217 0.00700602
R5646 VDD.n202 VDD.n201 0.00669433
R5647 VDD.n10 VDD.n9 0.00661998
R5648 VDD.n220 VDD.n219 0.00638785
R5649 VDD.n162 VDD.n159 0.00632996
R5650 VDD.n149 VDD.n146 0.00632996
R5651 VDD.n143 VDD.n137 0.00632996
R5652 VDD.n92 VDD.n89 0.00632996
R5653 VDD VDD.n1377 0.00630645
R5654 VDD VDD.n1364 0.00630645
R5655 VDD.n473 VDD 0.00630645
R5656 VDD VDD.n451 0.00630645
R5657 VDD.n361 VDD 0.00630645
R5658 VDD VDD.n30 0.00630645
R5659 VDD.n267 VDD.n266 0.00582544
R5660 VDD.n63 VDD.n62 0.00579412
R5661 VDD.n221 VDD.n220 0.00572908
R5662 VDD.n383 VDD.n382 0.00562195
R5663 VDD.n67 VDD.n66 0.00558696
R5664 VDD.n387 VDD.n386 0.00489628
R5665 VDD.n184 VDD.n93 0.00487247
R5666 VDD.n69 VDD.n68 0.00480435
R5667 VDD.n185 VDD.n184 0.0045081
R5668 VDD.n176 VDD.n175 0.0045081
R5669 VDD.n141 VDD.n140 0.00441304
R5670 VDD.n135 VDD.n134 0.00414372
R5671 VDD.n198 VDD.n197 0.00414372
R5672 VDD.n331 VDD.n330 0.00412903
R5673 VDD.n19 VDD.n18 0.00412903
R5674 VDD.n405 VDD.n404 0.00402941
R5675 VDD.n61 VDD.n60 0.00402941
R5676 VDD.n150 VDD.n149 0.00377935
R5677 VDD.n137 VDD.n136 0.00377935
R5678 VDD.n84 VDD.n83 0.00377935
R5679 VDD.n330 VDD.n329 0.00376613
R5680 VDD.n754 VDD.n753 0.00371429
R5681 VDD.n1338 VDD.n1335 0.00371429
R5682 VDD.n409 VDD.n71 0.00360796
R5683 VDD.n265 VDD.n264 0.00350186
R5684 VDD.n188 VDD.n185 0.00341498
R5685 VDD VDD.n281 0.00340323
R5686 VDD.n58 VDD.n57 0.00340323
R5687 VDD.n89 VDD.n84 0.00305061
R5688 VDD.n210 VDD.n209 0.00305061
R5689 VDD.n332 VDD.n331 0.00304032
R5690 VDD.n223 VDD.n222 0.00283401
R5691 VDD.n589 VDD.n586 0.00266867
R5692 VDD.n1238 VDD.n1237 0.00266867
R5693 VDD.n124 VDD 0.00254545
R5694 VDD.n14 VDD.n11 0.00254545
R5695 VDD.n177 VDD.n174 0.00245652
R5696 VDD.n142 VDD.n139 0.00206522
R5697 VDD.n855 VDD.n854 0.00192857
R5698 VDD.n201 VDD.n198 0.00159312
R5699 VDD.n197 VDD.n196 0.00159312
R5700 VDD.n806 VDD.n803 0.00152273
R5701 VDD.n1082 VDD.n1081 0.00152273
R5702 VDD VDD.n412 0.00151695
R5703 VDD.n146 VDD.n143 0.00122874
R5704 VDD.n53 VDD.n50 0.00122581
R5705 VDD.n1577 VDD.n1574 0.00121429
R5706 VDD.n266 VDD.n265 0.00103254
R5707 VDD.n11 VDD.n10 0.00101136
R5708 VDD.n329 VDD.n328 0.000862903
R5709 VDD.n249 VDD 0.000851563
R5710 VCTRL.n0 VCTRL.t0 27.5268
R5711 VCTRL.n13 VCTRL.t19 27.5268
R5712 VCTRL.n15 VCTRL.t6 25.3421
R5713 VCTRL.n3 VCTRL.t8 25.3421
R5714 VCTRL VCTRL.n12 9.02002
R5715 VCTRL.n17 VCTRL.t17 8.86359
R5716 VCTRL.n5 VCTRL.t18 8.86319
R5717 VCTRL.n20 VCTRL.t12 7.92693
R5718 VCTRL.n7 VCTRL.t7 7.92693
R5719 VCTRL.n4 VCTRL.t13 7.79605
R5720 VCTRL.n18 VCTRL.t4 7.79604
R5721 VCTRL.n1 VCTRL.t10 7.57548
R5722 VCTRL.n14 VCTRL.t9 7.54055
R5723 VCTRL.n2 VCTRL.t3 7.49426
R5724 VCTRL.n19 VCTRL.t14 7.49422
R5725 VCTRL.n8 VCTRL.t16 6.73304
R5726 VCTRL.n21 VCTRL.t1 6.73129
R5727 VCTRL.n1 VCTRL.n0 4.72106
R5728 VCTRL.n14 VCTRL.n13 4.72106
R5729 VCTRL.n6 VCTRL.n3 3.90288
R5730 VCTRL.n16 VCTRL.n15 3.90053
R5731 VCTRL.n11 VCTRL 2.50091
R5732 VCTRL.n24 VCTRL 2.46425
R5733 VCTRL.n12 VCTRL 2.32969
R5734 VCTRL.n15 VCTRL.t5 2.17312
R5735 VCTRL.n0 VCTRL.t2 2.17312
R5736 VCTRL.n3 VCTRL.t11 2.17312
R5737 VCTRL.n13 VCTRL.t15 2.17312
R5738 VCTRL.n25 VCTRL.n24 1.89901
R5739 VCTRL.n22 VCTRL.n21 1.89604
R5740 VCTRL.n9 VCTRL.n8 1.89145
R5741 VCTRL.n23 VCTRL.n22 1.5395
R5742 VCTRL.n10 VCTRL.n9 1.5395
R5743 VCTRL.n26 VCTRL.n25 1.4706
R5744 VCTRL.n7 VCTRL.n6 1.05913
R5745 VCTRL.n9 VCTRL.n2 0.957464
R5746 VCTRL.n22 VCTRL.n19 0.95718
R5747 VCTRL.n12 VCTRL.n11 0.798473
R5748 VCTRL.n5 VCTRL.n4 0.749817
R5749 VCTRL.n18 VCTRL.n17 0.749568
R5750 VCTRL.n19 VCTRL.n18 0.62372
R5751 VCTRL.n4 VCTRL.n2 0.622675
R5752 VCTRL.n17 VCTRL.n16 0.602194
R5753 VCTRL.n6 VCTRL.n5 0.602194
R5754 VCTRL VCTRL.n26 0.550625
R5755 VCTRL.n8 VCTRL.n7 0.453053
R5756 VCTRL.n21 VCTRL.n20 0.451554
R5757 VCTRL.n11 VCTRL.n10 0.43025
R5758 VCTRL.n24 VCTRL.n23 0.43025
R5759 VCTRL.n10 VCTRL.n1 0.266
R5760 VCTRL.n23 VCTRL.n14 0.266
R5761 VCTRL.n26 VCTRL 0.231324
R5762 VCTRL.n25 VCTRL 0.0563767
R5763 VCO_C_0.INV_2_1.IN.n23 VCO_C_0.INV_2_1.IN.t14 23.6945
R5764 VCO_C_0.INV_2_1.IN.t18 VCO_C_0.INV_2_1.IN.n24 23.6945
R5765 VCO_C_0.INV_2_1.IN.n24 VCO_C_0.INV_2_1.IN.n23 18.8035
R5766 VCO_C_0.INV_2_1.IN.n21 VCO_C_0.INV_2_1.IN.n19 15.8172
R5767 VCO_C_0.INV_2_1.IN.n21 VCO_C_0.INV_2_1.IN.n20 15.8172
R5768 VCO_C_0.INV_2_1.IN.n20 VCO_C_0.INV_2_1.IN.n16 15.8172
R5769 VCO_C_0.INV_2_1.IN.n19 VCO_C_0.INV_2_1.IN.t23 14.8925
R5770 VCO_C_0.INV_2_1.IN.t20 VCO_C_0.INV_2_1.IN.n21 14.8925
R5771 VCO_C_0.INV_2_1.IN.n20 VCO_C_0.INV_2_1.IN.t13 14.8925
R5772 VCO_C_0.INV_2_1.IN.n25 VCO_C_0.INV_2_1.IN.n17 12.2457
R5773 VCO_C_0.INV_2_1.IN.n22 VCO_C_0.INV_2_1.IN.n17 12.2457
R5774 VCO_C_0.INV_2_1.IN.n22 VCO_C_0.INV_2_1.IN.n18 12.2457
R5775 VCO_C_0.INV_2_1.IN.n26 VCO_C_0.INV_2_1.IN.t19 11.6285
R5776 VCO_C_0.INV_2_1.IN.n18 VCO_C_0.INV_2_1.IN.t14 8.9065
R5777 VCO_C_0.INV_2_1.IN.t15 VCO_C_0.INV_2_1.IN.n22 8.9065
R5778 VCO_C_0.INV_2_1.IN.t17 VCO_C_0.INV_2_1.IN.n17 8.9065
R5779 VCO_C_0.INV_2_1.IN.n25 VCO_C_0.INV_2_1.IN.t18 8.9065
R5780 VCO_C_0.INV_2_1.IN.n21 VCO_C_0.INV_2_1.IN.t22 8.6145
R5781 VCO_C_0.INV_2_1.IN.n19 VCO_C_0.INV_2_1.IN.t12 8.6145
R5782 VCO_C_0.INV_2_1.IN.n20 VCO_C_0.INV_2_1.IN.t16 8.6145
R5783 VCO_C_0.INV_2_1.IN.n16 VCO_C_0.INV_2_1.IN.t21 8.59715
R5784 VCO_C_0.INV_2_1.IN.t23 VCO_C_0.INV_2_1.IN.n18 8.3225
R5785 VCO_C_0.INV_2_1.IN.n22 VCO_C_0.INV_2_1.IN.t20 8.3225
R5786 VCO_C_0.INV_2_1.IN.t13 VCO_C_0.INV_2_1.IN.n17 8.3225
R5787 VCO_C_0.INV_2_1.IN.t19 VCO_C_0.INV_2_1.IN.n25 8.3225
R5788 VCO_C_0.INV_2_1.IN VCO_C_0.INV_2_1.IN.n26 4.223
R5789 VCO_C_0.INV_2_1.IN.n23 VCO_C_0.INV_2_1.IN.t15 3.6505
R5790 VCO_C_0.INV_2_1.IN.n24 VCO_C_0.INV_2_1.IN.t17 3.6505
R5791 VCO_C_0.INV_2_1.IN.n10 VCO_C_0.INV_2_1.IN.t3 3.6405
R5792 VCO_C_0.INV_2_1.IN.n10 VCO_C_0.INV_2_1.IN.n9 3.6405
R5793 VCO_C_0.INV_2_1.IN.n3 VCO_C_0.INV_2_1.IN.t4 3.6405
R5794 VCO_C_0.INV_2_1.IN.n3 VCO_C_0.INV_2_1.IN.n2 3.6405
R5795 VCO_C_0.INV_2_1.IN.n5 VCO_C_0.INV_2_1.IN.t0 3.6405
R5796 VCO_C_0.INV_2_1.IN.n5 VCO_C_0.INV_2_1.IN.n4 3.6405
R5797 VCO_C_0.INV_2_1.IN.n12 VCO_C_0.INV_2_1.IN.t5 3.6405
R5798 VCO_C_0.INV_2_1.IN.n12 VCO_C_0.INV_2_1.IN.n11 3.6405
R5799 VCO_C_0.INV_2_1.IN.n14 VCO_C_0.INV_2_1.IN.n8 3.50463
R5800 VCO_C_0.INV_2_1.IN.n15 VCO_C_0.INV_2_1.IN.n1 3.50463
R5801 VCO_C_0.INV_2_1.IN.n8 VCO_C_0.INV_2_1.IN.t9 3.2765
R5802 VCO_C_0.INV_2_1.IN.n8 VCO_C_0.INV_2_1.IN.n7 3.2765
R5803 VCO_C_0.INV_2_1.IN.n1 VCO_C_0.INV_2_1.IN.t10 3.2765
R5804 VCO_C_0.INV_2_1.IN.n1 VCO_C_0.INV_2_1.IN.n0 3.2765
R5805 VCO_C_0.INV_2_1.IN.n26 VCO_C_0.INV_2_1.IN.n16 3.1807
R5806 VCO_C_0.INV_2_1.IN.n6 VCO_C_0.INV_2_1.IN.n5 3.06224
R5807 VCO_C_0.INV_2_1.IN.n13 VCO_C_0.INV_2_1.IN.n12 3.06224
R5808 VCO_C_0.INV_2_1.IN.n6 VCO_C_0.INV_2_1.IN.n3 2.6005
R5809 VCO_C_0.INV_2_1.IN.n13 VCO_C_0.INV_2_1.IN.n10 2.6005
R5810 VCO_C_0.INV_2_1.IN.n15 VCO_C_0.INV_2_1.IN.n14 0.798761
R5811 VCO_C_0.INV_2_1.IN VCO_C_0.INV_2_1.IN.n15 0.562022
R5812 VCO_C_0.INV_2_1.IN.n15 VCO_C_0.INV_2_1.IN.n6 0.18637
R5813 VCO_C_0.INV_2_1.IN.n14 VCO_C_0.INV_2_1.IN.n13 0.18637
R5814 VCO_C_0.OUTB.n20 VCO_C_0.OUTB.t17 45.6363
R5815 VCO_C_0.OUTB.n26 VCO_C_0.OUTB.t47 45.6363
R5816 VCO_C_0.OUTB.n23 VCO_C_0.OUTB.t19 29.6446
R5817 VCO_C_0.OUTB.t53 VCO_C_0.OUTB.n24 29.6446
R5818 VCO_C_0.OUTB.n29 VCO_C_0.OUTB.t45 29.6446
R5819 VCO_C_0.OUTB.t43 VCO_C_0.OUTB.n30 29.6446
R5820 VCO_C_0.OUTB.n19 VCO_C_0.OUTB.t20 24.6117
R5821 VCO_C_0.OUTB.n28 VCO_C_0.OUTB.t28 24.6117
R5822 VCO_C_0.OUTB.n40 VCO_C_0.OUTB.t46 23.6945
R5823 VCO_C_0.OUTB.t32 VCO_C_0.OUTB.n41 23.6945
R5824 VCO_C_0.OUTB.n24 VCO_C_0.OUTB.n23 22.2047
R5825 VCO_C_0.OUTB.n30 VCO_C_0.OUTB.n29 22.2047
R5826 VCO_C_0.OUTB.t17 VCO_C_0.OUTB.t14 22.1925
R5827 VCO_C_0.OUTB.t47 VCO_C_0.OUTB.t13 22.1925
R5828 VCO_C_0.OUTB.n21 VCO_C_0.OUTB.n20 20.9314
R5829 VCO_C_0.OUTB.n27 VCO_C_0.OUTB.n26 20.9314
R5830 VCO_C_0.OUTB.n41 VCO_C_0.OUTB.n40 18.8035
R5831 VCO_C_0.OUTB VCO_C_0.OUTB.t43 18.5191
R5832 VCO_C_0.OUTB.n25 VCO_C_0.OUTB.t53 17.9055
R5833 VCO_C_0.OUTB.n38 VCO_C_0.OUTB.n36 15.8172
R5834 VCO_C_0.OUTB.n38 VCO_C_0.OUTB.n37 15.8172
R5835 VCO_C_0.OUTB.n37 VCO_C_0.OUTB.n33 15.8172
R5836 VCO_C_0.OUTB.n46 VCO_C_0.OUTB.t12 15.4917
R5837 VCO_C_0.OUTB.n48 VCO_C_0.OUTB.t38 15.3942
R5838 VCO_C_0.OUTB.n49 VCO_C_0.OUTB.t41 14.9265
R5839 VCO_C_0.OUTB.n36 VCO_C_0.OUTB.t24 14.8925
R5840 VCO_C_0.OUTB.t44 VCO_C_0.OUTB.n38 14.8925
R5841 VCO_C_0.OUTB.n37 VCO_C_0.OUTB.t33 14.8925
R5842 VCO_C_0.OUTB.n53 VCO_C_0.OUTB.t29 14.7749
R5843 VCO_C_0.OUTB.n47 VCO_C_0.OUTB.t39 13.6019
R5844 VCO_C_0.OUTB.n53 VCO_C_0.OUTB.t35 13.5312
R5845 VCO_C_0.OUTB.n51 VCO_C_0.OUTB.t22 13.4877
R5846 VCO_C_0.OUTB.n49 VCO_C_0.OUTB.t31 13.227
R5847 VCO_C_0.OUTB.n50 VCO_C_0.OUTB.t30 13.1835
R5848 VCO_C_0.OUTB.n42 VCO_C_0.OUTB.n34 12.2457
R5849 VCO_C_0.OUTB.n39 VCO_C_0.OUTB.n34 12.2457
R5850 VCO_C_0.OUTB.n39 VCO_C_0.OUTB.n35 12.2457
R5851 VCO_C_0.OUTB.n43 VCO_C_0.OUTB.t51 11.6285
R5852 VCO_C_0.OUTB.n45 VCO_C_0.OUTB.n2 9.0064
R5853 VCO_C_0.OUTB.n35 VCO_C_0.OUTB.t46 8.9065
R5854 VCO_C_0.OUTB.t23 VCO_C_0.OUTB.n39 8.9065
R5855 VCO_C_0.OUTB.t52 VCO_C_0.OUTB.n34 8.9065
R5856 VCO_C_0.OUTB.n42 VCO_C_0.OUTB.t32 8.9065
R5857 VCO_C_0.OUTB.n38 VCO_C_0.OUTB.t36 8.6145
R5858 VCO_C_0.OUTB.n36 VCO_C_0.OUTB.t16 8.6145
R5859 VCO_C_0.OUTB.n37 VCO_C_0.OUTB.t26 8.6145
R5860 VCO_C_0.OUTB.n33 VCO_C_0.OUTB.t48 8.59715
R5861 VCO_C_0.OUTB.t24 VCO_C_0.OUTB.n35 8.3225
R5862 VCO_C_0.OUTB.n39 VCO_C_0.OUTB.t44 8.3225
R5863 VCO_C_0.OUTB.t33 VCO_C_0.OUTB.n34 8.3225
R5864 VCO_C_0.OUTB.t51 VCO_C_0.OUTB.n42 8.3225
R5865 VCO_C_0.OUTB.n2 VCO_C_0.OUTB.n25 8.24338
R5866 VCO_C_0.OUTB.n46 VCO_C_0.OUTB.t40 8.1387
R5867 VCO_C_0.OUTB.n23 VCO_C_0.OUTB.t42 6.1325
R5868 VCO_C_0.OUTB.n24 VCO_C_0.OUTB.t34 6.1325
R5869 VCO_C_0.OUTB.n19 VCO_C_0.OUTB.t25 6.1325
R5870 VCO_C_0.OUTB.n20 VCO_C_0.OUTB.t27 6.1325
R5871 VCO_C_0.OUTB.n21 VCO_C_0.OUTB.t21 6.1325
R5872 VCO_C_0.OUTB.n28 VCO_C_0.OUTB.t49 6.1325
R5873 VCO_C_0.OUTB.n29 VCO_C_0.OUTB.t50 6.1325
R5874 VCO_C_0.OUTB.n30 VCO_C_0.OUTB.t18 6.1325
R5875 VCO_C_0.OUTB.n26 VCO_C_0.OUTB.t15 6.1325
R5876 VCO_C_0.OUTB.n27 VCO_C_0.OUTB.t37 6.1325
R5877 VCO_C_0.OUTB.n32 VCO_C_0.OUTB.n27 5.5044
R5878 VCO_C_0.OUTB.n22 VCO_C_0.OUTB.n21 5.38991
R5879 VCO_C_0.OUTB.n22 VCO_C_0.OUTB.n19 4.83094
R5880 VCO_C_0.OUTB.n31 VCO_C_0.OUTB.n28 4.83094
R5881 VCO_C_0.OUTB VCO_C_0.OUTB.n43 4.223
R5882 VCO_C_0.OUTB.n40 VCO_C_0.OUTB.t23 3.6505
R5883 VCO_C_0.OUTB.n41 VCO_C_0.OUTB.t52 3.6505
R5884 VCO_C_0.OUTB.n13 VCO_C_0.OUTB.t3 3.6405
R5885 VCO_C_0.OUTB.n13 VCO_C_0.OUTB.n12 3.6405
R5886 VCO_C_0.OUTB.n6 VCO_C_0.OUTB.t1 3.6405
R5887 VCO_C_0.OUTB.n6 VCO_C_0.OUTB.n5 3.6405
R5888 VCO_C_0.OUTB.n8 VCO_C_0.OUTB.t5 3.6405
R5889 VCO_C_0.OUTB.n8 VCO_C_0.OUTB.n7 3.6405
R5890 VCO_C_0.OUTB.n15 VCO_C_0.OUTB.t2 3.6405
R5891 VCO_C_0.OUTB.n15 VCO_C_0.OUTB.n14 3.6405
R5892 VCO_C_0.OUTB.n17 VCO_C_0.OUTB.n11 3.50463
R5893 VCO_C_0.OUTB.n18 VCO_C_0.OUTB.n4 3.50463
R5894 VCO_C_0.OUTB.n11 VCO_C_0.OUTB.t9 3.2765
R5895 VCO_C_0.OUTB.n11 VCO_C_0.OUTB.n10 3.2765
R5896 VCO_C_0.OUTB.n4 VCO_C_0.OUTB.t8 3.2765
R5897 VCO_C_0.OUTB.n4 VCO_C_0.OUTB.n3 3.2765
R5898 VCO_C_0.OUTB.n43 VCO_C_0.OUTB.n33 3.1807
R5899 VCO_C_0.OUTB.n9 VCO_C_0.OUTB.n8 3.06224
R5900 VCO_C_0.OUTB.n16 VCO_C_0.OUTB.n13 3.06224
R5901 VCO_C_0.OUTB.n2 VCO_C_0.OUTB.n44 2.82705
R5902 VCO_C_0.OUTB.n9 VCO_C_0.OUTB.n6 2.6005
R5903 VCO_C_0.OUTB.n16 VCO_C_0.OUTB.n15 2.6005
R5904 VCO_C_0.OUTB.n2 VCO_C_0.OUTB 2.36547
R5905 VCO_C_0.OUTB VCO_C_0.OUTB.n56 2.30807
R5906 VCO_C_0.OUTB.n0 VCO_C_0.OUTB.n1 1.10603
R5907 VCO_C_0.OUTB.n56 VCO_C_0.OUTB.n55 2.2505
R5908 VCO_C_0.OUTB.n52 VCO_C_0.OUTB.n48 1.5982
R5909 VCO_C_0.OUTB.n54 VCO_C_0.OUTB.n52 1.18336
R5910 VCO_C_0.OUTB.n55 VCO_C_0.OUTB.n54 0.977746
R5911 VCO_C_0.OUTB.n18 VCO_C_0.OUTB.n17 0.798761
R5912 VCO_C_0.OUTB.n45 VCO_C_0.OUTB.n0 0.66931
R5913 VCO_C_0.OUTB VCO_C_0.OUTB.n22 0.658318
R5914 VCO_C_0.OUTB.n31 VCO_C_0.OUTB 0.637045
R5915 VCO_C_0.OUTB.n25 VCO_C_0.OUTB 0.6125
R5916 VCO_C_0.OUTB VCO_C_0.OUTB.n18 0.562022
R5917 VCO_C_0.OUTB.n32 VCO_C_0.OUTB.n31 0.458758
R5918 VCO_C_0.OUTB.n47 VCO_C_0.OUTB.n46 0.381495
R5919 VCO_C_0.OUTB.n54 VCO_C_0.OUTB.n53 0.37501
R5920 VCO_C_0.OUTB.n48 VCO_C_0.OUTB.n47 0.355126
R5921 VCO_C_0.OUTB.n51 VCO_C_0.OUTB.n50 0.31227
R5922 VCO_C_0.OUTB.n50 VCO_C_0.OUTB.n49 0.298874
R5923 VCO_C_0.OUTB.n56 VCO_C_0.OUTB.n0 0.281082
R5924 VCO_C_0.OUTB.n44 VCO_C_0.OUTB.n32 0.238532
R5925 VCO_C_0.OUTB.n52 VCO_C_0.OUTB.n51 0.233052
R5926 VCO_C_0.OUTB.n18 VCO_C_0.OUTB.n9 0.18637
R5927 VCO_C_0.OUTB.n17 VCO_C_0.OUTB.n16 0.18637
R5928 VCO_C_0.OUTB VCO_C_0.OUTB.n1 0.203752
R5929 VCO_C_0.OUTB.n55 VCO_C_0.OUTB.n45 0.137564
R5930 VCO_C_0.OUTB.n44 VCO_C_0.OUTB 0.104622
R5931 VCO_C_0.OUTB.n1 VCO_C_0.OUTB 0.147946
R5932 VCO_C_0.INV_2_5.IN.n12 VCO_C_0.INV_2_5.IN.t43 23.6945
R5933 VCO_C_0.INV_2_5.IN.n13 VCO_C_0.INV_2_5.IN.t51 23.6945
R5934 VCO_C_0.INV_2_5.IN.n13 VCO_C_0.INV_2_5.IN.n12 18.8035
R5935 VCO_C_0.INV_2_5.IN.n10 VCO_C_0.INV_2_5.IN.n7 15.8172
R5936 VCO_C_0.INV_2_5.IN.n16 VCO_C_0.INV_2_5.IN.n15 15.8172
R5937 VCO_C_0.INV_2_5.IN.n15 VCO_C_0.INV_2_5.IN.n7 15.8172
R5938 VCO_C_0.INV_2_5.IN.t58 VCO_C_0.INV_2_5.IN.n10 14.8925
R5939 VCO_C_0.INV_2_5.IN.t44 VCO_C_0.INV_2_5.IN.n7 14.8925
R5940 VCO_C_0.INV_2_5.IN.n15 VCO_C_0.INV_2_5.IN.t50 14.8925
R5941 VCO_C_0.INV_2_5.IN.n14 VCO_C_0.INV_2_5.IN.n8 12.2457
R5942 VCO_C_0.INV_2_5.IN.n14 VCO_C_0.INV_2_5.IN.n9 12.2457
R5943 VCO_C_0.INV_2_5.IN.n11 VCO_C_0.INV_2_5.IN.n9 12.2457
R5944 VCO_C_0.INV_2_5.IN.n17 VCO_C_0.INV_2_5.IN.t39 11.6285
R5945 VCO_C_0.INV_2_5.IN.n62 VCO_C_0.INV_2_5.IN.t57 9.07373
R5946 VCO_C_0.INV_2_5.IN.n66 VCO_C_0.INV_2_5.IN.t49 8.94903
R5947 VCO_C_0.INV_2_5.IN.n72 VCO_C_0.INV_2_5.IN.t55 8.91906
R5948 VCO_C_0.INV_2_5.IN.n71 VCO_C_0.INV_2_5.IN.t56 8.91906
R5949 VCO_C_0.INV_2_5.IN.n70 VCO_C_0.INV_2_5.IN.t33 8.91906
R5950 VCO_C_0.INV_2_5.IN.t43 VCO_C_0.INV_2_5.IN.n11 8.9065
R5951 VCO_C_0.INV_2_5.IN.t31 VCO_C_0.INV_2_5.IN.n9 8.9065
R5952 VCO_C_0.INV_2_5.IN.n14 VCO_C_0.INV_2_5.IN.t38 8.9065
R5953 VCO_C_0.INV_2_5.IN.t51 VCO_C_0.INV_2_5.IN.n8 8.9065
R5954 VCO_C_0.INV_2_5.IN.n68 VCO_C_0.INV_2_5.IN.t47 8.88175
R5955 VCO_C_0.INV_2_5.IN.n64 VCO_C_0.INV_2_5.IN.t52 8.78051
R5956 VCO_C_0.INV_2_5.IN.n67 VCO_C_0.INV_2_5.IN.t48 8.78051
R5957 VCO_C_0.INV_2_5.IN.n63 VCO_C_0.INV_2_5.IN.t53 8.76753
R5958 VCO_C_0.INV_2_5.IN.n62 VCO_C_0.INV_2_5.IN.t36 8.76753
R5959 VCO_C_0.INV_2_5.IN.n30 VCO_C_0.INV_2_5.IN.t5 8.71893
R5960 VCO_C_0.INV_2_5.IN.n69 VCO_C_0.INV_2_5.IN.t40 8.71324
R5961 VCO_C_0.INV_2_5.IN.n2 VCO_C_0.INV_2_5.IN.t42 8.71324
R5962 VCO_C_0.INV_2_5.IN.n10 VCO_C_0.INV_2_5.IN.t54 8.6145
R5963 VCO_C_0.INV_2_5.IN.n7 VCO_C_0.INV_2_5.IN.t41 8.6145
R5964 VCO_C_0.INV_2_5.IN.n15 VCO_C_0.INV_2_5.IN.t46 8.6145
R5965 VCO_C_0.INV_2_5.IN.n16 VCO_C_0.INV_2_5.IN.t35 8.59715
R5966 VCO_C_0.INV_2_5.IN.n0 VCO_C_0.INV_2_5.IN.t34 8.50259
R5967 VCO_C_0.INV_2_5.IN.n4 VCO_C_0.INV_2_5.IN.t45 8.38837
R5968 VCO_C_0.INV_2_5.IN.n11 VCO_C_0.INV_2_5.IN.t58 8.3225
R5969 VCO_C_0.INV_2_5.IN.n9 VCO_C_0.INV_2_5.IN.t44 8.3225
R5970 VCO_C_0.INV_2_5.IN.t50 VCO_C_0.INV_2_5.IN.n14 8.3225
R5971 VCO_C_0.INV_2_5.IN.n8 VCO_C_0.INV_2_5.IN.t39 8.3225
R5972 VCO_C_0.INV_2_5.IN.n65 VCO_C_0.INV_2_5.IN.t32 8.30411
R5973 VCO_C_0.INV_2_5.IN.n6 VCO_C_0.INV_2_5.IN.t13 7.93952
R5974 VCO_C_0.INV_2_5.IN.n68 VCO_C_0.INV_2_5.IN.t37 7.40199
R5975 VCO_C_0.INV_2_5.IN.n81 VCO_C_0.INV_2_5.IN.t20 6.43598
R5976 VCO_C_0.INV_2_5.IN.n29 VCO_C_0.INV_2_5.IN.n26 6.42121
R5977 VCO_C_0.INV_2_5.IN.n5 VCO_C_0.INV_2_5.IN.t19 6.39767
R5978 VCO_C_0.INV_2_5.IN.n1 VCO_C_0.INV_2_5.IN.t30 6.02861
R5979 VCO_C_0.INV_2_5.IN.n24 VCO_C_0.INV_2_5.IN.n23 5.82997
R5980 VCO_C_0.INV_2_5.IN.n47 VCO_C_0.INV_2_5.IN.n46 5.30071
R5981 VCO_C_0.INV_2_5.IN.n29 VCO_C_0.INV_2_5.IN.n28 5.23266
R5982 VCO_C_0.INV_2_5.IN.n39 VCO_C_0.INV_2_5.IN.t24 4.89657
R5983 VCO_C_0.INV_2_5.IN.n60 VCO_C_0.INV_2_5.IN.n59 4.89332
R5984 VCO_C_0.INV_2_5.IN VCO_C_0.INV_2_5.IN.n82 4.88822
R5985 VCO_C_0.INV_2_5.IN.n30 VCO_C_0.INV_2_5.IN.t2 4.76585
R5986 VCO_C_0.INV_2_5.IN.n25 VCO_C_0.INV_2_5.IN.n20 4.70534
R5987 VCO_C_0.INV_2_5.IN.n26 VCO_C_0.INV_2_5.IN.n19 4.70317
R5988 VCO_C_0.INV_2_5.IN VCO_C_0.INV_2_5.IN.n17 4.60939
R5989 VCO_C_0.INV_2_5.IN.n61 VCO_C_0.INV_2_5.IN.n84 4.53389
R5990 VCO_C_0.INV_2_5.IN.n61 VCO_C_0.INV_2_5.IN.n83 4.10346
R5991 VCO_C_0.INV_2_5.IN.n42 VCO_C_0.INV_2_5.IN.n41 4.04842
R5992 VCO_C_0.INV_2_5.IN.n83 VCO_C_0.INV_2_5.IN.t25 4.00791
R5993 VCO_C_0.INV_2_5.IN.n74 VCO_C_0.INV_2_5.IN.n73 3.96274
R5994 VCO_C_0.INV_2_5.IN.n34 VCO_C_0.INV_2_5.IN.n18 3.95313
R5995 VCO_C_0.INV_2_5.IN.n31 VCO_C_0.INV_2_5.IN.t6 3.94347
R5996 VCO_C_0.INV_2_5.IN.n85 VCO_C_0.INV_2_5.IN.t11 3.80888
R5997 VCO_C_0.INV_2_5.IN.n24 VCO_C_0.INV_2_5.IN.n22 3.77407
R5998 VCO_C_0.INV_2_5.IN.n81 VCO_C_0.INV_2_5.IN.n80 3.75752
R5999 VCO_C_0.INV_2_5.IN.n18 VCO_C_0.INV_2_5.IN 3.73676
R6000 VCO_C_0.INV_2_5.IN.n80 VCO_C_0.INV_2_5.IN.n79 3.65963
R6001 VCO_C_0.INV_2_5.IN.n12 VCO_C_0.INV_2_5.IN.t31 3.6505
R6002 VCO_C_0.INV_2_5.IN.t38 VCO_C_0.INV_2_5.IN.n13 3.6505
R6003 VCO_C_0.INV_2_5.IN.n55 VCO_C_0.INV_2_5.IN.t28 3.6405
R6004 VCO_C_0.INV_2_5.IN.n55 VCO_C_0.INV_2_5.IN.n54 3.6405
R6005 VCO_C_0.INV_2_5.IN.n49 VCO_C_0.INV_2_5.IN.t15 3.6405
R6006 VCO_C_0.INV_2_5.IN.n49 VCO_C_0.INV_2_5.IN.n48 3.6405
R6007 VCO_C_0.INV_2_5.IN.n36 VCO_C_0.INV_2_5.IN.t26 3.6405
R6008 VCO_C_0.INV_2_5.IN.n36 VCO_C_0.INV_2_5.IN.n35 3.6405
R6009 VCO_C_0.INV_2_5.IN.n28 VCO_C_0.INV_2_5.IN.n27 3.47613
R6010 VCO_C_0.INV_2_5.IN.n22 VCO_C_0.INV_2_5.IN.n21 3.47611
R6011 VCO_C_0.INV_2_5.IN.n32 VCO_C_0.INV_2_5.IN.n29 3.3208
R6012 VCO_C_0.INV_2_5.IN.n80 VCO_C_0.INV_2_5.IN.t18 3.31772
R6013 VCO_C_0.INV_2_5.IN.n85 VCO_C_0.INV_2_5.IN.n86 3.21498
R6014 VCO_C_0.INV_2_5.IN.n17 VCO_C_0.INV_2_5.IN.n16 3.1807
R6015 VCO_C_0.INV_2_5.IN VCO_C_0.INV_2_5.IN.n5 3.15891
R6016 VCO_C_0.INV_2_5.IN.n34 VCO_C_0.INV_2_5.IN.n33 3.14573
R6017 VCO_C_0.INV_2_5.IN.n25 VCO_C_0.INV_2_5.IN.n24 2.88722
R6018 VCO_C_0.INV_2_5.IN.n22 VCO_C_0.INV_2_5.IN.t4 2.86261
R6019 VCO_C_0.INV_2_5.IN.n28 VCO_C_0.INV_2_5.IN.t3 2.8626
R6020 VCO_C_0.INV_2_5.IN.n32 VCO_C_0.INV_2_5.IN.n31 2.83609
R6021 VCO_C_0.INV_2_5.IN.n3 VCO_C_0.INV_2_5.IN.n61 2.75901
R6022 VCO_C_0.INV_2_5.IN.n57 VCO_C_0.INV_2_5.IN.n6 2.62313
R6023 VCO_C_0.INV_2_5.IN.n18 VCO_C_0.INV_2_5.IN 2.36584
R6024 VCO_C_0.INV_2_5.IN.n77 VCO_C_0.INV_2_5.IN.n34 2.35267
R6025 VCO_C_0.INV_2_5.IN.n33 VCO_C_0.INV_2_5.IN 2.30603
R6026 VCO_C_0.INV_2_5.IN.n43 VCO_C_0.INV_2_5.IN.n42 2.24883
R6027 VCO_C_0.INV_2_5.IN.n76 VCO_C_0.INV_2_5.IN.n58 2.03424
R6028 VCO_C_0.INV_2_5.IN.n57 VCO_C_0.INV_2_5.IN.n38 1.94273
R6029 VCO_C_0.INV_2_5.IN.n6 VCO_C_0.INV_2_5.IN.n40 1.78522
R6030 VCO_C_0.INV_2_5.IN.n52 VCO_C_0.INV_2_5.IN.n53 1.77736
R6031 VCO_C_0.INV_2_5.IN.n52 VCO_C_0.INV_2_5.IN.n51 1.77011
R6032 VCO_C_0.INV_2_5.IN.n44 VCO_C_0.INV_2_5.IN.n43 1.76105
R6033 VCO_C_0.INV_2_5.IN.n44 VCO_C_0.INV_2_5.IN.n45 1.71456
R6034 VCO_C_0.INV_2_5.IN.n56 VCO_C_0.INV_2_5.IN.n55 1.66033
R6035 VCO_C_0.INV_2_5.IN.n6 VCO_C_0.INV_2_5.IN.n44 1.5995
R6036 VCO_C_0.INV_2_5.IN.n75 VCO_C_0.INV_2_5.IN.n74 1.5089
R6037 VCO_C_0.INV_2_5.IN.n40 VCO_C_0.INV_2_5.IN.n39 1.495
R6038 VCO_C_0.INV_2_5.IN.n51 VCO_C_0.INV_2_5.IN.n50 1.49487
R6039 VCO_C_0.INV_2_5.IN.n38 VCO_C_0.INV_2_5.IN.n37 1.49487
R6040 VCO_C_0.INV_2_5.IN.n78 VCO_C_0.INV_2_5.IN.n77 1.47485
R6041 VCO_C_0.INV_2_5.IN.n37 VCO_C_0.INV_2_5.IN.n36 1.25757
R6042 VCO_C_0.INV_2_5.IN.n50 VCO_C_0.INV_2_5.IN.n49 1.25657
R6043 VCO_C_0.INV_2_5.IN.n58 VCO_C_0.INV_2_5.IN.n57 1.22576
R6044 VCO_C_0.INV_2_5.IN.n0 VCO_C_0.INV_2_5.IN.n4 1.19023
R6045 VCO_C_0.INV_2_5.IN.n44 VCO_C_0.INV_2_5.IN.n52 1.1585
R6046 VCO_C_0.INV_2_5.IN.n3 VCO_C_0.INV_2_5.IN.n60 1.1375
R6047 VCO_C_0.INV_2_5.IN.n45 VCO_C_0.INV_2_5.IN.n47 1.1242
R6048 VCO_C_0.INV_2_5.IN.n53 VCO_C_0.INV_2_5.IN.n56 1.12383
R6049 VCO_C_0.INV_2_5.IN.n84 VCO_C_0.INV_2_5.IN.n85 1.00902
R6050 VCO_C_0.INV_2_5.IN.n5 VCO_C_0.INV_2_5.IN.n78 0.932551
R6051 VCO_C_0.INV_2_5.IN.n5 VCO_C_0.INV_2_5.IN.n81 0.878175
R6052 VCO_C_0.INV_2_5.IN.n76 VCO_C_0.INV_2_5.IN.n75 0.836557
R6053 VCO_C_0.INV_2_5.IN.n65 VCO_C_0.INV_2_5.IN.n64 0.650226
R6054 VCO_C_0.INV_2_5.IN.n77 VCO_C_0.INV_2_5.IN.n76 0.596796
R6055 VCO_C_0.INV_2_5.IN.n33 VCO_C_0.INV_2_5.IN.n32 0.488268
R6056 VCO_C_0.INV_2_5.IN.n2 VCO_C_0.INV_2_5.IN.n70 0.486253
R6057 VCO_C_0.INV_2_5.IN.n31 VCO_C_0.INV_2_5.IN.n30 0.476518
R6058 VCO_C_0.INV_2_5.IN.n26 VCO_C_0.INV_2_5.IN.n25 0.471952
R6059 VCO_C_0.INV_2_5.IN.n75 VCO_C_0.INV_2_5.IN.n0 0.412247
R6060 VCO_C_0.INV_2_5.IN.n2 VCO_C_0.INV_2_5.IN.n1 0.387961
R6061 VCO_C_0.INV_2_5.IN.n4 VCO_C_0.INV_2_5.IN.n3 0.382089
R6062 VCO_C_0.INV_2_5.IN.n67 VCO_C_0.INV_2_5.IN.n66 0.345705
R6063 VCO_C_0.INV_2_5.IN.n69 VCO_C_0.INV_2_5.IN.n68 0.345705
R6064 VCO_C_0.INV_2_5.IN.n4 VCO_C_0.INV_2_5.IN.n67 0.34324
R6065 VCO_C_0.INV_2_5.IN.n63 VCO_C_0.INV_2_5.IN.n62 0.342007
R6066 VCO_C_0.INV_2_5.IN.n72 VCO_C_0.INV_2_5.IN.n71 0.342007
R6067 VCO_C_0.INV_2_5.IN.n71 VCO_C_0.INV_2_5.IN.n2 0.33461
R6068 VCO_C_0.INV_2_5.IN.n64 VCO_C_0.INV_2_5.IN.n63 0.325979
R6069 VCO_C_0.INV_2_5.IN.n66 VCO_C_0.INV_2_5.IN.n65 0.318582
R6070 VCO_C_0.INV_2_5.IN.n0 VCO_C_0.INV_2_5.IN.n72 0.312418
R6071 VCO_C_0.INV_2_5.IN.n70 VCO_C_0.INV_2_5.IN.n69 0.312418
R6072 VCO_C_0.INV_2_5.OUT.n2 VCO_C_0.INV_2_5.OUT.t14 15.4917
R6073 VCO_C_0.INV_2_5.OUT.n4 VCO_C_0.INV_2_5.OUT.t13 15.3942
R6074 VCO_C_0.INV_2_5.OUT.n5 VCO_C_0.INV_2_5.OUT.t20 14.904
R6075 VCO_C_0.INV_2_5.OUT.n9 VCO_C_0.INV_2_5.OUT.t18 14.7749
R6076 VCO_C_0.INV_2_5.OUT.n3 VCO_C_0.INV_2_5.OUT.t12 13.6019
R6077 VCO_C_0.INV_2_5.OUT.n9 VCO_C_0.INV_2_5.OUT.t16 13.5312
R6078 VCO_C_0.INV_2_5.OUT.n7 VCO_C_0.INV_2_5.OUT.t17 13.4877
R6079 VCO_C_0.INV_2_5.OUT.n5 VCO_C_0.INV_2_5.OUT.t21 13.227
R6080 VCO_C_0.INV_2_5.OUT.n6 VCO_C_0.INV_2_5.OUT.t15 13.1835
R6081 VCO_C_0.INV_2_5.OUT.n2 VCO_C_0.INV_2_5.OUT.t19 8.17943
R6082 VCO_C_0.INV_2_5.OUT VCO_C_0.INV_2_5.OUT.n0 4.7425
R6083 VCO_C_0.INV_2_5.OUT.n26 VCO_C_0.INV_2_5.OUT.t0 3.6405
R6084 VCO_C_0.INV_2_5.OUT.n26 VCO_C_0.INV_2_5.OUT.n25 3.6405
R6085 VCO_C_0.INV_2_5.OUT.n18 VCO_C_0.INV_2_5.OUT.t2 3.6405
R6086 VCO_C_0.INV_2_5.OUT.n18 VCO_C_0.INV_2_5.OUT.n17 3.6405
R6087 VCO_C_0.INV_2_5.OUT.n16 VCO_C_0.INV_2_5.OUT.t6 3.6405
R6088 VCO_C_0.INV_2_5.OUT.n16 VCO_C_0.INV_2_5.OUT.n15 3.6405
R6089 VCO_C_0.INV_2_5.OUT.n24 VCO_C_0.INV_2_5.OUT.t4 3.6405
R6090 VCO_C_0.INV_2_5.OUT.n24 VCO_C_0.INV_2_5.OUT.n23 3.6405
R6091 VCO_C_0.INV_2_5.OUT.n28 VCO_C_0.INV_2_5.OUT.n14 3.50463
R6092 VCO_C_0.INV_2_5.OUT.n22 VCO_C_0.INV_2_5.OUT.n21 3.50463
R6093 VCO_C_0.INV_2_5.OUT.n14 VCO_C_0.INV_2_5.OUT.t8 3.2765
R6094 VCO_C_0.INV_2_5.OUT.n14 VCO_C_0.INV_2_5.OUT.n13 3.2765
R6095 VCO_C_0.INV_2_5.OUT.n21 VCO_C_0.INV_2_5.OUT.t9 3.2765
R6096 VCO_C_0.INV_2_5.OUT.n21 VCO_C_0.INV_2_5.OUT.n20 3.2765
R6097 VCO_C_0.INV_2_5.OUT.n19 VCO_C_0.INV_2_5.OUT.n16 3.06224
R6098 VCO_C_0.INV_2_5.OUT.n27 VCO_C_0.INV_2_5.OUT.n24 3.06224
R6099 VCO_C_0.INV_2_5.OUT.n19 VCO_C_0.INV_2_5.OUT.n18 2.6005
R6100 VCO_C_0.INV_2_5.OUT.n27 VCO_C_0.INV_2_5.OUT.n26 2.6005
R6101 VCO_C_0.INV_2_5.OUT.n1 VCO_C_0.INV_2_5.OUT 2.28587
R6102 VCO_C_0.INV_2_5.OUT.n12 VCO_C_0.INV_2_5.OUT.n1 2.2505
R6103 VCO_C_0.INV_2_5.OUT.n8 VCO_C_0.INV_2_5.OUT.n4 1.5982
R6104 VCO_C_0.INV_2_5.OUT.n10 VCO_C_0.INV_2_5.OUT.n8 1.18336
R6105 VCO_C_0.INV_2_5.OUT.n11 VCO_C_0.INV_2_5.OUT.n10 0.961395
R6106 VCO_C_0.INV_2_5.OUT.n1 VCO_C_0.INV_2_5.OUT.n11 0.806561
R6107 VCO_C_0.INV_2_5.OUT.n28 VCO_C_0.INV_2_5.OUT.n22 0.798761
R6108 VCO_C_0.INV_2_5.OUT.n0 VCO_C_0.INV_2_5.OUT 0.65726
R6109 VCO_C_0.INV_2_5.OUT.n1 VCO_C_0.INV_2_5.OUT.n0 0.56461
R6110 VCO_C_0.INV_2_5.OUT VCO_C_0.INV_2_5.OUT.n28 0.539611
R6111 VCO_C_0.INV_2_5.OUT.n3 VCO_C_0.INV_2_5.OUT.n2 0.381495
R6112 VCO_C_0.INV_2_5.OUT.n10 VCO_C_0.INV_2_5.OUT.n9 0.37501
R6113 VCO_C_0.INV_2_5.OUT.n4 VCO_C_0.INV_2_5.OUT.n3 0.355126
R6114 VCO_C_0.INV_2_5.OUT.n7 VCO_C_0.INV_2_5.OUT.n6 0.31227
R6115 VCO_C_0.INV_2_5.OUT.n6 VCO_C_0.INV_2_5.OUT.n5 0.298874
R6116 VCO_C_0.INV_2_5.OUT.n8 VCO_C_0.INV_2_5.OUT.n7 0.233052
R6117 VCO_C_0.INV_2_5.OUT.n22 VCO_C_0.INV_2_5.OUT.n19 0.18637
R6118 VCO_C_0.INV_2_5.OUT.n28 VCO_C_0.INV_2_5.OUT.n27 0.18637
R6119 VCO_C_0.INV_2_5.OUT VCO_C_0.INV_2_5.OUT.n12 0.185454
R6120 a_17597_1404.n5 a_17597_1404.t9 29.2961
R6121 a_17597_1404.n6 a_17597_1404.n5 21.9292
R6122 a_17597_1404.n7 a_17597_1404.n6 18.1271
R6123 a_17597_1404.n7 a_17597_1404.t6 11.1695
R6124 a_17597_1404.n3 a_17597_1404.t5 10.2143
R6125 a_17597_1404.n5 a_17597_1404.t7 6.1325
R6126 a_17597_1404.n6 a_17597_1404.t8 6.1325
R6127 a_17597_1404.n3 a_17597_1404.n2 4.68517
R6128 a_17597_1404.n8 a_17597_1404.n7 4.6311
R6129 a_17597_1404.n9 a_17597_1404.n8 2.85093
R6130 a_17597_1404.n1 a_17597_1404.t0 2.16717
R6131 a_17597_1404.n1 a_17597_1404.n0 2.16717
R6132 a_17597_1404.n9 a_17597_1404.t1 2.16717
R6133 a_17597_1404.n10 a_17597_1404.n9 2.16717
R6134 a_17597_1404.n4 a_17597_1404.n3 1.58582
R6135 a_17597_1404.n4 a_17597_1404.n1 1.24371
R6136 a_17597_1404.n8 a_17597_1404.n4 0.971051
R6137 DFF_3_mag_0.INV_2_5.OUT.n3 DFF_3_mag_0.INV_2_5.OUT.n2 5.81586
R6138 DFF_3_mag_0.INV_2_5.OUT.n8 DFF_3_mag_0.INV_2_5.OUT.t1 5.10148
R6139 DFF_3_mag_0.INV_2_5.OUT.n5 DFF_3_mag_0.INV_2_5.OUT.t2 5.1005
R6140 DFF_3_mag_0.INV_2_5.OUT.n4 DFF_3_mag_0.INV_2_5.OUT.t19 5.08021
R6141 DFF_3_mag_0.INV_2_5.OUT.n8 DFF_3_mag_0.INV_2_5.OUT.n7 4.66166
R6142 DFF_3_mag_0.INV_2_5.OUT.n19 DFF_3_mag_0.INV_2_5.OUT.t15 3.6405
R6143 DFF_3_mag_0.INV_2_5.OUT.n19 DFF_3_mag_0.INV_2_5.OUT.n18 3.6405
R6144 DFF_3_mag_0.INV_2_5.OUT.n21 DFF_3_mag_0.INV_2_5.OUT.t11 3.6405
R6145 DFF_3_mag_0.INV_2_5.OUT.n21 DFF_3_mag_0.INV_2_5.OUT.n20 3.6405
R6146 DFF_3_mag_0.INV_2_5.OUT.n12 DFF_3_mag_0.INV_2_5.OUT.t13 3.6405
R6147 DFF_3_mag_0.INV_2_5.OUT.n12 DFF_3_mag_0.INV_2_5.OUT.n11 3.6405
R6148 DFF_3_mag_0.INV_2_5.OUT.n14 DFF_3_mag_0.INV_2_5.OUT.t8 3.6405
R6149 DFF_3_mag_0.INV_2_5.OUT.n14 DFF_3_mag_0.INV_2_5.OUT.n13 3.6405
R6150 DFF_3_mag_0.INV_2_5.OUT.n23 DFF_3_mag_0.INV_2_5.OUT.n17 3.50463
R6151 DFF_3_mag_0.INV_2_5.OUT.n24 DFF_3_mag_0.INV_2_5.OUT.n10 3.50463
R6152 DFF_3_mag_0.INV_2_5.OUT.n17 DFF_3_mag_0.INV_2_5.OUT.t4 3.2765
R6153 DFF_3_mag_0.INV_2_5.OUT.n17 DFF_3_mag_0.INV_2_5.OUT.n16 3.2765
R6154 DFF_3_mag_0.INV_2_5.OUT.n10 DFF_3_mag_0.INV_2_5.OUT.t14 3.2765
R6155 DFF_3_mag_0.INV_2_5.OUT.n10 DFF_3_mag_0.INV_2_5.OUT.n9 3.2765
R6156 DFF_3_mag_0.INV_2_5.OUT.n22 DFF_3_mag_0.INV_2_5.OUT.n21 3.06224
R6157 DFF_3_mag_0.INV_2_5.OUT.n15 DFF_3_mag_0.INV_2_5.OUT.n14 3.06224
R6158 DFF_3_mag_0.INV_2_5.OUT.n3 DFF_3_mag_0.INV_2_5.OUT.n1 2.85093
R6159 DFF_3_mag_0.INV_2_5.OUT.n22 DFF_3_mag_0.INV_2_5.OUT.n19 2.6005
R6160 DFF_3_mag_0.INV_2_5.OUT.n15 DFF_3_mag_0.INV_2_5.OUT.n12 2.6005
R6161 DFF_3_mag_0.INV_2_5.OUT.n1 DFF_3_mag_0.INV_2_5.OUT.t18 2.16717
R6162 DFF_3_mag_0.INV_2_5.OUT.n1 DFF_3_mag_0.INV_2_5.OUT.n0 2.16717
R6163 DFF_3_mag_0.INV_2_5.OUT.n7 DFF_3_mag_0.INV_2_5.OUT.t0 1.9505
R6164 DFF_3_mag_0.INV_2_5.OUT.n7 DFF_3_mag_0.INV_2_5.OUT.n6 1.9505
R6165 DFF_3_mag_0.INV_2_5.OUT.n24 DFF_3_mag_0.INV_2_5.OUT.n23 0.798761
R6166 DFF_3_mag_0.INV_2_5.OUT.n4 DFF_3_mag_0.INV_2_5.OUT.n3 0.644196
R6167 DFF_3_mag_0.INV_2_5.OUT DFF_3_mag_0.INV_2_5.OUT.n24 0.562022
R6168 DFF_3_mag_0.INV_2_5.OUT.n5 DFF_3_mag_0.INV_2_5.OUT.n4 0.447229
R6169 DFF_3_mag_0.INV_2_5.OUT DFF_3_mag_0.INV_2_5.OUT.n5 0.392597
R6170 DFF_3_mag_0.INV_2_5.OUT DFF_3_mag_0.INV_2_5.OUT.n8 0.308628
R6171 DFF_3_mag_0.INV_2_5.OUT.n23 DFF_3_mag_0.INV_2_5.OUT.n22 0.18637
R6172 DFF_3_mag_0.INV_2_5.OUT.n24 DFF_3_mag_0.INV_2_5.OUT.n15 0.18637
R6173 DFF_3_mag_0.INV_2_1.IN.n27 DFF_3_mag_0.INV_2_1.IN.t17 23.6945
R6174 DFF_3_mag_0.INV_2_1.IN.n28 DFF_3_mag_0.INV_2_1.IN.t20 23.6945
R6175 DFF_3_mag_0.INV_2_1.IN.n28 DFF_3_mag_0.INV_2_1.IN.n27 18.8035
R6176 DFF_3_mag_0.INV_2_1.IN.n25 DFF_3_mag_0.INV_2_1.IN.n22 15.8172
R6177 DFF_3_mag_0.INV_2_1.IN.n31 DFF_3_mag_0.INV_2_1.IN.n30 15.8172
R6178 DFF_3_mag_0.INV_2_1.IN.n30 DFF_3_mag_0.INV_2_1.IN.n22 15.8172
R6179 DFF_3_mag_0.INV_2_1.IN.t22 DFF_3_mag_0.INV_2_1.IN.n25 14.8925
R6180 DFF_3_mag_0.INV_2_1.IN.t16 DFF_3_mag_0.INV_2_1.IN.n22 14.8925
R6181 DFF_3_mag_0.INV_2_1.IN.n30 DFF_3_mag_0.INV_2_1.IN.t19 14.8925
R6182 DFF_3_mag_0.INV_2_1.IN.n29 DFF_3_mag_0.INV_2_1.IN.n23 12.2457
R6183 DFF_3_mag_0.INV_2_1.IN.n29 DFF_3_mag_0.INV_2_1.IN.n24 12.2457
R6184 DFF_3_mag_0.INV_2_1.IN.n26 DFF_3_mag_0.INV_2_1.IN.n24 12.2457
R6185 DFF_3_mag_0.INV_2_1.IN.n32 DFF_3_mag_0.INV_2_1.IN.t25 11.6285
R6186 DFF_3_mag_0.INV_2_1.IN.t17 DFF_3_mag_0.INV_2_1.IN.n26 8.9065
R6187 DFF_3_mag_0.INV_2_1.IN.t23 DFF_3_mag_0.INV_2_1.IN.n24 8.9065
R6188 DFF_3_mag_0.INV_2_1.IN.n29 DFF_3_mag_0.INV_2_1.IN.t26 8.9065
R6189 DFF_3_mag_0.INV_2_1.IN.t20 DFF_3_mag_0.INV_2_1.IN.n23 8.9065
R6190 DFF_3_mag_0.INV_2_1.IN.n25 DFF_3_mag_0.INV_2_1.IN.t21 8.6145
R6191 DFF_3_mag_0.INV_2_1.IN.n22 DFF_3_mag_0.INV_2_1.IN.t27 8.6145
R6192 DFF_3_mag_0.INV_2_1.IN.n30 DFF_3_mag_0.INV_2_1.IN.t18 8.6145
R6193 DFF_3_mag_0.INV_2_1.IN.n31 DFF_3_mag_0.INV_2_1.IN.t24 8.59715
R6194 DFF_3_mag_0.INV_2_1.IN.n26 DFF_3_mag_0.INV_2_1.IN.t22 8.3225
R6195 DFF_3_mag_0.INV_2_1.IN.n24 DFF_3_mag_0.INV_2_1.IN.t16 8.3225
R6196 DFF_3_mag_0.INV_2_1.IN.t19 DFF_3_mag_0.INV_2_1.IN.n29 8.3225
R6197 DFF_3_mag_0.INV_2_1.IN.n23 DFF_3_mag_0.INV_2_1.IN.t25 8.3225
R6198 DFF_3_mag_0.INV_2_1.IN.n33 DFF_3_mag_0.INV_2_1.IN 6.97731
R6199 DFF_3_mag_0.INV_2_1.IN.n0 DFF_3_mag_0.INV_2_1.IN.n18 6.74326
R6200 DFF_3_mag_0.INV_2_1.IN.n1 DFF_3_mag_0.INV_2_1.IN.n8 6.74326
R6201 DFF_3_mag_0.INV_2_1.IN.n0 DFF_3_mag_0.INV_2_1.IN.n19 5.1005
R6202 DFF_3_mag_0.INV_2_1.IN.n1 DFF_3_mag_0.INV_2_1.IN.n9 5.1005
R6203 DFF_3_mag_0.INV_2_1.IN DFF_3_mag_0.INV_2_1.IN.n32 4.21749
R6204 DFF_3_mag_0.INV_2_1.IN.n27 DFF_3_mag_0.INV_2_1.IN.t23 3.6505
R6205 DFF_3_mag_0.INV_2_1.IN.t26 DFF_3_mag_0.INV_2_1.IN.n28 3.6505
R6206 DFF_3_mag_0.INV_2_1.IN.n6 DFF_3_mag_0.INV_2_1.IN.n3 3.57508
R6207 DFF_3_mag_0.INV_2_1.IN.n16 DFF_3_mag_0.INV_2_1.IN.n15 3.5743
R6208 DFF_3_mag_0.INV_2_1.IN.n1 DFF_3_mag_0.INV_2_1.IN.t0 3.40075
R6209 DFF_3_mag_0.INV_2_1.IN.n0 DFF_3_mag_0.INV_2_1.IN.t8 3.40065
R6210 DFF_3_mag_0.INV_2_1.IN.n32 DFF_3_mag_0.INV_2_1.IN.n31 3.1807
R6211 DFF_3_mag_0.INV_2_1.IN.n20 DFF_3_mag_0.INV_2_1.IN.n17 3.00034
R6212 DFF_3_mag_0.INV_2_1.IN.n10 DFF_3_mag_0.INV_2_1.IN.n7 3.00032
R6213 DFF_3_mag_0.INV_2_1.IN DFF_3_mag_0.INV_2_1.IN.n21 2.58093
R6214 DFF_3_mag_0.INV_2_1.IN DFF_3_mag_0.INV_2_1.IN.n11 2.5808
R6215 DFF_3_mag_0.INV_2_1.IN.n13 DFF_3_mag_0.INV_2_1.IN.t6 2.16717
R6216 DFF_3_mag_0.INV_2_1.IN.n13 DFF_3_mag_0.INV_2_1.IN.n12 2.16717
R6217 DFF_3_mag_0.INV_2_1.IN.n15 DFF_3_mag_0.INV_2_1.IN.t7 2.16717
R6218 DFF_3_mag_0.INV_2_1.IN.n15 DFF_3_mag_0.INV_2_1.IN.n14 2.16717
R6219 DFF_3_mag_0.INV_2_1.IN.n3 DFF_3_mag_0.INV_2_1.IN.t12 2.16717
R6220 DFF_3_mag_0.INV_2_1.IN.n3 DFF_3_mag_0.INV_2_1.IN.n2 2.16717
R6221 DFF_3_mag_0.INV_2_1.IN.n5 DFF_3_mag_0.INV_2_1.IN.t13 2.16717
R6222 DFF_3_mag_0.INV_2_1.IN.n5 DFF_3_mag_0.INV_2_1.IN.n4 2.16717
R6223 DFF_3_mag_0.INV_2_1.IN.n11 DFF_3_mag_0.INV_2_1.IN.n10 1.8481
R6224 DFF_3_mag_0.INV_2_1.IN.n21 DFF_3_mag_0.INV_2_1.IN.n20 1.847
R6225 DFF_3_mag_0.INV_2_1.IN.n16 DFF_3_mag_0.INV_2_1.IN.n13 1.25225
R6226 DFF_3_mag_0.INV_2_1.IN.n6 DFF_3_mag_0.INV_2_1.IN.n5 1.25187
R6227 DFF_3_mag_0.INV_2_1.IN.n21 DFF_3_mag_0.INV_2_1.IN.n16 1.12594
R6228 DFF_3_mag_0.INV_2_1.IN.n11 DFF_3_mag_0.INV_2_1.IN.n6 1.12561
R6229 DFF_3_mag_0.INV_2_1.IN.n33 DFF_3_mag_0.INV_2_1.IN 0.812356
R6230 DFF_3_mag_0.INV_2_1.IN DFF_3_mag_0.INV_2_1.IN.n33 0.728851
R6231 DFF_3_mag_0.INV_2_1.IN.n20 DFF_3_mag_0.INV_2_1.IN.n0 0.559412
R6232 DFF_3_mag_0.INV_2_1.IN.n10 DFF_3_mag_0.INV_2_1.IN.n1 0.558374
R6233 VCTRL2.n65 VCTRL2.n63 10.0043
R6234 VCTRL2.n123 VCTRL2.n65 9.34779
R6235 VCTRL2.n115 VCTRL2.t45 8.213
R6236 VCTRL2.n83 VCTRL2.t42 8.213
R6237 VCTRL2.n52 VCTRL2.t59 8.16955
R6238 VCTRL2.n40 VCTRL2.t30 8.16955
R6239 VCTRL2.n88 VCTRL2.t11 8.16955
R6240 VCTRL2.n74 VCTRL2.t10 8.16955
R6241 VCTRL2.n79 VCTRL2.t36 8.16955
R6242 VCTRL2.n120 VCTRL2.t44 8.16955
R6243 VCTRL2.n30 VCTRL2.t19 8.1261
R6244 VCTRL2.n23 VCTRL2.t43 8.1261
R6245 VCTRL2.n36 VCTRL2.t13 8.1261
R6246 VCTRL2.n57 VCTRL2.t5 8.1261
R6247 VCTRL2.n101 VCTRL2.t0 8.1261
R6248 VCTRL2.n70 VCTRL2.t74 8.1261
R6249 VCTRL2.n17 VCTRL2.t72 8.08264
R6250 VCTRL2.n9 VCTRL2.t54 8.08264
R6251 VCTRL2.n106 VCTRL2.t4 7.51776
R6252 VCTRL2.n81 VCTRL2.t1 7.51776
R6253 VCTRL2.n49 VCTRL2.t24 7.47431
R6254 VCTRL2.n38 VCTRL2.t77 7.47431
R6255 VCTRL2.n118 VCTRL2.t3 7.47431
R6256 VCTRL2.n86 VCTRL2.t47 7.47431
R6257 VCTRL2.n72 VCTRL2.t46 7.47431
R6258 VCTRL2.n113 VCTRL2.t66 7.47431
R6259 VCTRL2.n76 VCTRL2.t76 7.47431
R6260 VCTRL2.n82 VCTRL2.t62 7.47431
R6261 VCTRL2.n28 VCTRL2.t61 7.43086
R6262 VCTRL2.n21 VCTRL2.t12 7.43086
R6263 VCTRL2.n51 VCTRL2.t39 7.43086
R6264 VCTRL2.n34 VCTRL2.t56 7.43086
R6265 VCTRL2.n55 VCTRL2.t52 7.43086
R6266 VCTRL2.n39 VCTRL2.t14 7.43086
R6267 VCTRL2.n87 VCTRL2.t27 7.43086
R6268 VCTRL2.n73 VCTRL2.t26 7.43086
R6269 VCTRL2.n96 VCTRL2.t40 7.43086
R6270 VCTRL2.n67 VCTRL2.t33 7.43086
R6271 VCTRL2.n77 VCTRL2.t57 7.43086
R6272 VCTRL2.n119 VCTRL2.t65 7.43086
R6273 VCTRL2.n29 VCTRL2.t79 7.3874
R6274 VCTRL2.n22 VCTRL2.t25 7.3874
R6275 VCTRL2.n12 VCTRL2.t38 7.3874
R6276 VCTRL2.n6 VCTRL2.t18 7.3874
R6277 VCTRL2.n35 VCTRL2.t71 7.3874
R6278 VCTRL2.n56 VCTRL2.t67 7.3874
R6279 VCTRL2.n97 VCTRL2.t20 7.3874
R6280 VCTRL2.n68 VCTRL2.t15 7.3874
R6281 VCTRL2.n16 VCTRL2.t53 7.34395
R6282 VCTRL2.n8 VCTRL2.t32 7.34395
R6283 VCTRL2.n18 VCTRL2.t50 7.3005
R6284 VCTRL2.n10 VCTRL2.t28 7.3005
R6285 VCTRL2.n37 VCTRL2.t68 7.25705
R6286 VCTRL2.n31 VCTRL2.t75 7.25705
R6287 VCTRL2.n24 VCTRL2.t21 7.25705
R6288 VCTRL2.t72 VCTRL2.n16 7.25705
R6289 VCTRL2.t54 VCTRL2.n8 7.25705
R6290 VCTRL2.n58 VCTRL2.t63 7.25705
R6291 VCTRL2.n102 VCTRL2.t23 7.25705
R6292 VCTRL2.n71 VCTRL2.t17 7.25705
R6293 VCTRL2.n41 VCTRL2.t8 7.2136
R6294 VCTRL2.t19 VCTRL2.n29 7.2136
R6295 VCTRL2.t43 VCTRL2.n22 7.2136
R6296 VCTRL2.t53 VCTRL2.n12 7.2136
R6297 VCTRL2.t32 VCTRL2.n6 7.2136
R6298 VCTRL2.n53 VCTRL2.t37 7.2136
R6299 VCTRL2.t13 VCTRL2.n35 7.2136
R6300 VCTRL2.t5 VCTRL2.n56 7.2136
R6301 VCTRL2.n89 VCTRL2.t31 7.2136
R6302 VCTRL2.n75 VCTRL2.t29 7.2136
R6303 VCTRL2.t0 VCTRL2.n97 7.2136
R6304 VCTRL2.t74 VCTRL2.n68 7.2136
R6305 VCTRL2.n80 VCTRL2.t58 7.2136
R6306 VCTRL2.n121 VCTRL2.t69 7.2136
R6307 VCTRL2.t79 VCTRL2.n28 7.17014
R6308 VCTRL2.t25 VCTRL2.n21 7.17014
R6309 VCTRL2.t59 VCTRL2.n51 7.17014
R6310 VCTRL2.t71 VCTRL2.n34 7.17014
R6311 VCTRL2.t67 VCTRL2.n55 7.17014
R6312 VCTRL2.t30 VCTRL2.n39 7.17014
R6313 VCTRL2.t11 VCTRL2.n87 7.17014
R6314 VCTRL2.t10 VCTRL2.n73 7.17014
R6315 VCTRL2.t20 VCTRL2.n96 7.17014
R6316 VCTRL2.t15 VCTRL2.n67 7.17014
R6317 VCTRL2.n116 VCTRL2.t70 7.17014
R6318 VCTRL2.t36 VCTRL2.n77 7.17014
R6319 VCTRL2.t44 VCTRL2.n119 7.17014
R6320 VCTRL2.n84 VCTRL2.t64 7.17014
R6321 VCTRL2.t39 VCTRL2.n49 7.12669
R6322 VCTRL2.t14 VCTRL2.n38 7.12669
R6323 VCTRL2.t27 VCTRL2.n86 7.12669
R6324 VCTRL2.t26 VCTRL2.n72 7.12669
R6325 VCTRL2.t45 VCTRL2.n113 7.12669
R6326 VCTRL2.t57 VCTRL2.n76 7.12669
R6327 VCTRL2.t65 VCTRL2.n118 7.12669
R6328 VCTRL2.t42 VCTRL2.n82 7.12669
R6329 VCTRL2.t66 VCTRL2.n106 7.08324
R6330 VCTRL2.n116 VCTRL2.t7 7.08324
R6331 VCTRL2.t62 VCTRL2.n81 7.08324
R6332 VCTRL2.n84 VCTRL2.t2 7.08324
R6333 VCTRL2.n53 VCTRL2.t22 7.03979
R6334 VCTRL2.n41 VCTRL2.t73 7.03979
R6335 VCTRL2.n89 VCTRL2.t49 7.03979
R6336 VCTRL2.n75 VCTRL2.t48 7.03979
R6337 VCTRL2.n80 VCTRL2.t78 7.03979
R6338 VCTRL2.n121 VCTRL2.t6 7.03979
R6339 VCTRL2.n37 VCTRL2.t55 6.99633
R6340 VCTRL2.n31 VCTRL2.t60 6.99633
R6341 VCTRL2.n24 VCTRL2.t9 6.99633
R6342 VCTRL2.n58 VCTRL2.t51 6.99633
R6343 VCTRL2.n102 VCTRL2.t41 6.99633
R6344 VCTRL2.n71 VCTRL2.t34 6.99633
R6345 VCTRL2.n18 VCTRL2.t35 6.95288
R6346 VCTRL2.n10 VCTRL2.t16 6.95288
R6347 VCTRL2.t35 VCTRL2.n17 6.51836
R6348 VCTRL2.t16 VCTRL2.n9 6.51836
R6349 VCTRL2.t55 VCTRL2.n36 6.4749
R6350 VCTRL2.t60 VCTRL2.n30 6.4749
R6351 VCTRL2.t9 VCTRL2.n23 6.4749
R6352 VCTRL2.t51 VCTRL2.n57 6.4749
R6353 VCTRL2.t41 VCTRL2.n101 6.4749
R6354 VCTRL2.t34 VCTRL2.n70 6.4749
R6355 VCTRL2.t22 VCTRL2.n52 6.43145
R6356 VCTRL2.t73 VCTRL2.n40 6.43145
R6357 VCTRL2.t49 VCTRL2.n88 6.43145
R6358 VCTRL2.t48 VCTRL2.n74 6.43145
R6359 VCTRL2.t78 VCTRL2.n79 6.43145
R6360 VCTRL2.t6 VCTRL2.n120 6.43145
R6361 VCTRL2.t7 VCTRL2.n115 6.388
R6362 VCTRL2.t2 VCTRL2.n83 6.388
R6363 VCTRL2.n85 VCTRL2.n84 4.03166
R6364 VCTRL2.n42 VCTRL2.n41 4.0306
R6365 VCTRL2.n59 VCTRL2.n58 3.63007
R6366 VCTRL2.n122 VCTRL2.n121 3.62933
R6367 VCTRL2.n43 VCTRL2.n31 3.62466
R6368 VCTRL2.n30 VCTRL2.n26 3.62466
R6369 VCTRL2.n49 VCTRL2.n48 3.62466
R6370 VCTRL2.n67 VCTRL2.n66 3.62466
R6371 VCTRL2.n96 VCTRL2.n95 3.62466
R6372 VCTRL2.n85 VCTRL2.n80 3.62466
R6373 VCTRL2.n91 VCTRL2.n75 3.62466
R6374 VCTRL2.n104 VCTRL2.n71 3.62466
R6375 VCTRL2.n28 VCTRL2.n27 3.62466
R6376 VCTRL2.n52 VCTRL2.n47 3.62466
R6377 VCTRL2.n54 VCTRL2.n53 3.62466
R6378 VCTRL2.n51 VCTRL2.n50 3.62466
R6379 VCTRL2.n101 VCTRL2.n100 3.62466
R6380 VCTRL2.n103 VCTRL2.n102 3.62466
R6381 VCTRL2.n70 VCTRL2.n69 3.62466
R6382 VCTRL2.n79 VCTRL2.n78 3.62466
R6383 VCTRL2.n42 VCTRL2.n37 3.62462
R6384 VCTRL2.n23 VCTRL2.n19 3.62462
R6385 VCTRL2.n44 VCTRL2.n24 3.62462
R6386 VCTRL2.n21 VCTRL2.n20 3.62462
R6387 VCTRL2.n45 VCTRL2.n18 3.62462
R6388 VCTRL2.n12 VCTRL2.n11 3.62462
R6389 VCTRL2.n16 VCTRL2.n15 3.62462
R6390 VCTRL2.n9 VCTRL2.n4 3.62462
R6391 VCTRL2.n46 VCTRL2.n10 3.62462
R6392 VCTRL2.n6 VCTRL2.n5 3.62462
R6393 VCTRL2.n8 VCTRL2.n7 3.62462
R6394 VCTRL2.n35 VCTRL2.n32 3.62462
R6395 VCTRL2.n34 VCTRL2.n33 3.62462
R6396 VCTRL2.n90 VCTRL2.n89 3.62462
R6397 VCTRL2.n106 VCTRL2.n105 3.62462
R6398 VCTRL2.n115 VCTRL2.n114 3.62462
R6399 VCTRL2.n117 VCTRL2.n116 3.62462
R6400 VCTRL2.n113 VCTRL2.n112 3.62462
R6401 VCTRL2.n62 VCTRL2.n61 2.2505
R6402 VCTRL2.n65 VCTRL2.n64 1.5049
R6403 VCTRL2 VCTRL2.n125 1.16594
R6404 VCTRL2 VCTRL2.n2 1.16341
R6405 VCTRL2.n62 VCTRL2.n59 1.05045
R6406 VCTRL2.n123 VCTRL2.n122 0.984409
R6407 VCTRL2.n60 VCTRL2 0.936261
R6408 VCTRL2.n0 VCTRL2 0.936261
R6409 VCTRL2.n64 VCTRL2 0.61117
R6410 VCTRL2.n59 VCTRL2.n54 0.442081
R6411 VCTRL2.n122 VCTRL2.n117 0.441056
R6412 VCTRL2.n109 VCTRL2.n108 0.404715
R6413 VCTRL2.n99 VCTRL2.n98 0.404715
R6414 VCTRL2.n91 VCTRL2.n90 0.404715
R6415 VCTRL2.n14 VCTRL2.n13 0.404539
R6416 VCTRL2.n44 VCTRL2.n43 0.404539
R6417 VCTRL2.n94 VCTRL2.n93 0.404539
R6418 VCTRL2.n103 VCTRL2.n91 0.401155
R6419 VCTRL2.n110 VCTRL2.n109 0.401155
R6420 VCTRL2.n100 VCTRL2.n99 0.401155
R6421 VCTRL2.n95 VCTRL2.n94 0.401155
R6422 VCTRL2.n15 VCTRL2.n14 0.400353
R6423 VCTRL2.n45 VCTRL2.n44 0.400353
R6424 VCTRL2.n104 VCTRL2.n103 0.398905
R6425 VCTRL2.n111 VCTRL2.n110 0.398484
R6426 VCTRL2.n112 VCTRL2.n111 0.398165
R6427 VCTRL2.n4 VCTRL2.n3 0.397928
R6428 VCTRL2.n117 VCTRL2.n104 0.397919
R6429 VCTRL2.n54 VCTRL2.n46 0.397919
R6430 VCTRL2.n46 VCTRL2.n45 0.397753
R6431 VCTRL2.n108 VCTRL2.n107 0.389969
R6432 VCTRL2.n43 VCTRL2.n42 0.389723
R6433 VCTRL2.n93 VCTRL2.n92 0.389723
R6434 VCTRL2.n26 VCTRL2.n25 0.389547
R6435 VCTRL2.n90 VCTRL2.n85 0.389547
R6436 VCTRL2.n64 VCTRL2 0.10046
R6437 VCTRL2.n63 VCTRL2.n2 0.0698976
R6438 VCTRL2.n125 VCTRL2.n124 0.0695909
R6439 VCTRL2.n61 VCTRL2 0.0362534
R6440 VCTRL2 VCTRL2.n1 0.0362534
R6441 VCTRL2.n63 VCTRL2.n62 0.0124277
R6442 VCTRL2.n124 VCTRL2.n123 0.00395428
R6443 VCTRL2.n61 VCTRL2.n60 0.00173288
R6444 VCTRL2.n1 VCTRL2.n0 0.00173288
R6445 VCO_C_0.INV_2_4.IN.n21 VCO_C_0.INV_2_4.IN.t15 23.6945
R6446 VCO_C_0.INV_2_4.IN.n22 VCO_C_0.INV_2_4.IN.t14 23.6945
R6447 VCO_C_0.INV_2_4.IN.n22 VCO_C_0.INV_2_4.IN.n21 18.8035
R6448 VCO_C_0.INV_2_4.IN.n19 VCO_C_0.INV_2_4.IN.n16 15.8172
R6449 VCO_C_0.INV_2_4.IN.n24 VCO_C_0.INV_2_4.IN.n16 15.8172
R6450 VCO_C_0.INV_2_4.IN.n25 VCO_C_0.INV_2_4.IN.n24 15.8172
R6451 VCO_C_0.INV_2_4.IN.t18 VCO_C_0.INV_2_4.IN.n19 14.8925
R6452 VCO_C_0.INV_2_4.IN.t13 VCO_C_0.INV_2_4.IN.n16 14.8925
R6453 VCO_C_0.INV_2_4.IN.n24 VCO_C_0.INV_2_4.IN.t22 14.8925
R6454 VCO_C_0.INV_2_4.IN.n23 VCO_C_0.INV_2_4.IN.n17 12.2457
R6455 VCO_C_0.INV_2_4.IN.n23 VCO_C_0.INV_2_4.IN.n18 12.2457
R6456 VCO_C_0.INV_2_4.IN.n20 VCO_C_0.INV_2_4.IN.n18 12.2457
R6457 VCO_C_0.INV_2_4.IN.n26 VCO_C_0.INV_2_4.IN.t17 11.6285
R6458 VCO_C_0.INV_2_4.IN.t15 VCO_C_0.INV_2_4.IN.n20 8.9065
R6459 VCO_C_0.INV_2_4.IN.t12 VCO_C_0.INV_2_4.IN.n18 8.9065
R6460 VCO_C_0.INV_2_4.IN.n23 VCO_C_0.INV_2_4.IN.t19 8.9065
R6461 VCO_C_0.INV_2_4.IN.t14 VCO_C_0.INV_2_4.IN.n17 8.9065
R6462 VCO_C_0.INV_2_4.IN.n19 VCO_C_0.INV_2_4.IN.t21 8.6145
R6463 VCO_C_0.INV_2_4.IN.n16 VCO_C_0.INV_2_4.IN.t16 8.6145
R6464 VCO_C_0.INV_2_4.IN.n24 VCO_C_0.INV_2_4.IN.t23 8.6145
R6465 VCO_C_0.INV_2_4.IN.n25 VCO_C_0.INV_2_4.IN.t20 8.59715
R6466 VCO_C_0.INV_2_4.IN.n20 VCO_C_0.INV_2_4.IN.t18 8.3225
R6467 VCO_C_0.INV_2_4.IN.n18 VCO_C_0.INV_2_4.IN.t13 8.3225
R6468 VCO_C_0.INV_2_4.IN.t22 VCO_C_0.INV_2_4.IN.n23 8.3225
R6469 VCO_C_0.INV_2_4.IN.n17 VCO_C_0.INV_2_4.IN.t17 8.3225
R6470 VCO_C_0.INV_2_4.IN VCO_C_0.INV_2_4.IN.n26 4.223
R6471 VCO_C_0.INV_2_4.IN.n21 VCO_C_0.INV_2_4.IN.t12 3.6505
R6472 VCO_C_0.INV_2_4.IN.t19 VCO_C_0.INV_2_4.IN.n22 3.6505
R6473 VCO_C_0.INV_2_4.IN.n13 VCO_C_0.INV_2_4.IN.t5 3.6405
R6474 VCO_C_0.INV_2_4.IN.n13 VCO_C_0.INV_2_4.IN.n12 3.6405
R6475 VCO_C_0.INV_2_4.IN.n5 VCO_C_0.INV_2_4.IN.t6 3.6405
R6476 VCO_C_0.INV_2_4.IN.n5 VCO_C_0.INV_2_4.IN.n4 3.6405
R6477 VCO_C_0.INV_2_4.IN.n3 VCO_C_0.INV_2_4.IN.t1 3.6405
R6478 VCO_C_0.INV_2_4.IN.n3 VCO_C_0.INV_2_4.IN.n2 3.6405
R6479 VCO_C_0.INV_2_4.IN.n11 VCO_C_0.INV_2_4.IN.t0 3.6405
R6480 VCO_C_0.INV_2_4.IN.n11 VCO_C_0.INV_2_4.IN.n10 3.6405
R6481 VCO_C_0.INV_2_4.IN.n15 VCO_C_0.INV_2_4.IN.n1 3.50463
R6482 VCO_C_0.INV_2_4.IN.n9 VCO_C_0.INV_2_4.IN.n8 3.50463
R6483 VCO_C_0.INV_2_4.IN.n1 VCO_C_0.INV_2_4.IN.t10 3.2765
R6484 VCO_C_0.INV_2_4.IN.n1 VCO_C_0.INV_2_4.IN.n0 3.2765
R6485 VCO_C_0.INV_2_4.IN.n8 VCO_C_0.INV_2_4.IN.t11 3.2765
R6486 VCO_C_0.INV_2_4.IN.n8 VCO_C_0.INV_2_4.IN.n7 3.2765
R6487 VCO_C_0.INV_2_4.IN.n26 VCO_C_0.INV_2_4.IN.n25 3.1807
R6488 VCO_C_0.INV_2_4.IN.n6 VCO_C_0.INV_2_4.IN.n3 3.06224
R6489 VCO_C_0.INV_2_4.IN.n14 VCO_C_0.INV_2_4.IN.n11 3.06224
R6490 VCO_C_0.INV_2_4.IN.n6 VCO_C_0.INV_2_4.IN.n5 2.6005
R6491 VCO_C_0.INV_2_4.IN.n14 VCO_C_0.INV_2_4.IN.n13 2.6005
R6492 VCO_C_0.INV_2_4.IN.n15 VCO_C_0.INV_2_4.IN.n9 0.798761
R6493 VCO_C_0.INV_2_4.IN VCO_C_0.INV_2_4.IN.n15 0.562022
R6494 VCO_C_0.INV_2_4.IN.n9 VCO_C_0.INV_2_4.IN.n6 0.18637
R6495 VCO_C_0.INV_2_4.IN.n15 VCO_C_0.INV_2_4.IN.n14 0.18637
R6496 VCO_C_0.OUT.n24 VCO_C_0.OUT.t15 14.1829
R6497 VCO_C_0.OUT.n23 VCO_C_0.OUT.t21 13.9657
R6498 VCO_C_0.OUT.n17 VCO_C_0.OUT.t17 13.3574
R6499 VCO_C_0.OUT.n16 VCO_C_0.OUT.t14 13.1401
R6500 VCO_C_0.OUT.n16 VCO_C_0.OUT.t16 12.9025
R6501 VCO_C_0.OUT.n18 VCO_C_0.OUT.t20 12.6187
R6502 VCO_C_0.OUT.n20 VCO_C_0.OUT.t13 8.77788
R6503 VCO_C_0.OUT.n19 VCO_C_0.OUT.t18 8.64752
R6504 VCO_C_0.OUT.n19 VCO_C_0.OUT.t12 8.56062
R6505 VCO_C_0.OUT.n20 VCO_C_0.OUT.t19 8.43026
R6506 VCO_C_0.OUT.n21 VCO_C_0.OUT.n19 6.11825
R6507 VCO_C_0.OUT.n21 VCO_C_0.OUT.n20 5.88354
R6508 VCO_C_0.OUT.n13 VCO_C_0.OUT.t6 3.6405
R6509 VCO_C_0.OUT.n13 VCO_C_0.OUT.n12 3.6405
R6510 VCO_C_0.OUT.n5 VCO_C_0.OUT.t3 3.6405
R6511 VCO_C_0.OUT.n5 VCO_C_0.OUT.n4 3.6405
R6512 VCO_C_0.OUT.n3 VCO_C_0.OUT.t5 3.6405
R6513 VCO_C_0.OUT.n3 VCO_C_0.OUT.n2 3.6405
R6514 VCO_C_0.OUT.n11 VCO_C_0.OUT.t7 3.6405
R6515 VCO_C_0.OUT.n11 VCO_C_0.OUT.n10 3.6405
R6516 VCO_C_0.OUT.n15 VCO_C_0.OUT.n1 3.50463
R6517 VCO_C_0.OUT.n9 VCO_C_0.OUT.n8 3.50463
R6518 VCO_C_0.OUT.n1 VCO_C_0.OUT.t11 3.2765
R6519 VCO_C_0.OUT.n1 VCO_C_0.OUT.n0 3.2765
R6520 VCO_C_0.OUT.n8 VCO_C_0.OUT.t10 3.2765
R6521 VCO_C_0.OUT.n8 VCO_C_0.OUT.n7 3.2765
R6522 VCO_C_0.OUT.n6 VCO_C_0.OUT.n3 3.06224
R6523 VCO_C_0.OUT.n14 VCO_C_0.OUT.n11 3.06224
R6524 VCO_C_0.OUT VCO_C_0.OUT.n24 2.91964
R6525 VCO_C_0.OUT.n6 VCO_C_0.OUT.n5 2.6005
R6526 VCO_C_0.OUT.n14 VCO_C_0.OUT.n13 2.6005
R6527 VCO_C_0.OUT.n23 VCO_C_0.OUT.n22 1.58291
R6528 VCO_C_0.OUT.n22 VCO_C_0.OUT.n18 1.47586
R6529 VCO_C_0.OUT.n24 VCO_C_0.OUT.n23 1.23958
R6530 VCO_C_0.OUT.n15 VCO_C_0.OUT.n9 0.798761
R6531 VCO_C_0.OUT VCO_C_0.OUT.n15 0.561439
R6532 VCO_C_0.OUT.n22 VCO_C_0.OUT.n21 0.448735
R6533 VCO_C_0.OUT.n18 VCO_C_0.OUT.n17 0.386992
R6534 VCO_C_0.OUT.n17 VCO_C_0.OUT.n16 0.340685
R6535 VCO_C_0.OUT.n9 VCO_C_0.OUT.n6 0.18637
R6536 VCO_C_0.OUT.n15 VCO_C_0.OUT.n14 0.18637
R6537 VCO_C_0.INV_2_0.IN.n9 VCO_C_0.INV_2_0.IN.n8 15.8172
R6538 VCO_C_0.INV_2_0.IN.n11 VCO_C_0.INV_2_0.IN.n10 15.8172
R6539 VCO_C_0.INV_2_0.IN.n10 VCO_C_0.INV_2_0.IN.n9 15.8172
R6540 VCO_C_0.INV_2_0.IN.n9 VCO_C_0.INV_2_0.IN.t37 14.8925
R6541 VCO_C_0.INV_2_0.IN.n10 VCO_C_0.INV_2_0.IN.t46 14.8925
R6542 VCO_C_0.INV_2_0.IN.n17 VCO_C_0.INV_2_0.IN.n16 12.2457
R6543 VCO_C_0.INV_2_0.IN.n16 VCO_C_0.INV_2_0.IN.n14 12.2457
R6544 VCO_C_0.INV_2_0.IN.n14 VCO_C_0.INV_2_0.IN.n12 12.2457
R6545 VCO_C_0.INV_2_0.IN.n18 VCO_C_0.INV_2_0.IN.t31 11.6285
R6546 VCO_C_0.INV_2_0.IN.n52 VCO_C_0.INV_2_0.IN.t38 9.5787
R6547 VCO_C_0.INV_2_0.IN.n49 VCO_C_0.INV_2_0.IN.t45 9.55768
R6548 VCO_C_0.INV_2_0.IN.n12 VCO_C_0.INV_2_0.IN.t57 8.9065
R6549 VCO_C_0.INV_2_0.IN.n14 VCO_C_0.INV_2_0.IN.t42 8.9065
R6550 VCO_C_0.INV_2_0.IN.n16 VCO_C_0.INV_2_0.IN.t49 8.9065
R6551 VCO_C_0.INV_2_0.IN.n17 VCO_C_0.INV_2_0.IN.t35 8.9065
R6552 VCO_C_0.INV_2_0.IN.n66 VCO_C_0.INV_2_0.IN.n62 8.86038
R6553 VCO_C_0.INV_2_0.IN.n9 VCO_C_0.INV_2_0.IN.t34 8.6145
R6554 VCO_C_0.INV_2_0.IN.n8 VCO_C_0.INV_2_0.IN.t47 8.6145
R6555 VCO_C_0.INV_2_0.IN.n10 VCO_C_0.INV_2_0.IN.t41 8.6145
R6556 VCO_C_0.INV_2_0.IN.n11 VCO_C_0.INV_2_0.IN.t56 8.59715
R6557 VCO_C_0.INV_2_0.IN.n52 VCO_C_0.INV_2_0.IN.t50 8.57144
R6558 VCO_C_0.INV_2_0.IN.n53 VCO_C_0.INV_2_0.IN.t44 8.57144
R6559 VCO_C_0.INV_2_0.IN.n54 VCO_C_0.INV_2_0.IN.t53 8.57144
R6560 VCO_C_0.INV_2_0.IN.n31 VCO_C_0.INV_2_0.IN.t10 8.54728
R6561 VCO_C_0.INV_2_0.IN.n5 VCO_C_0.INV_2_0.IN.t36 8.52112
R6562 VCO_C_0.INV_2_0.IN.n0 VCO_C_0.INV_2_0.IN.t32 8.52112
R6563 VCO_C_0.INV_2_0.IN.n2 VCO_C_0.INV_2_0.IN.t55 8.52112
R6564 VCO_C_0.INV_2_0.IN.n7 VCO_C_0.INV_2_0.IN.t54 8.52112
R6565 VCO_C_0.INV_2_0.IN.n51 VCO_C_0.INV_2_0.IN.t33 8.51092
R6566 VCO_C_0.INV_2_0.IN.n50 VCO_C_0.INV_2_0.IN.t51 8.51092
R6567 VCO_C_0.INV_2_0.IN.n49 VCO_C_0.INV_2_0.IN.t58 8.51092
R6568 VCO_C_0.INV_2_0.IN.n0 VCO_C_0.INV_2_0.IN.t43 8.35286
R6569 VCO_C_0.INV_2_0.IN.n12 VCO_C_0.INV_2_0.IN.t52 8.3225
R6570 VCO_C_0.INV_2_0.IN.t31 VCO_C_0.INV_2_0.IN.n17 8.3225
R6571 VCO_C_0.INV_2_0.IN.n7 VCO_C_0.INV_2_0.IN.t39 8.31073
R6572 VCO_C_0.INV_2_0.IN.n2 VCO_C_0.INV_2_0.IN.t40 8.31073
R6573 VCO_C_0.INV_2_0.IN.n5 VCO_C_0.INV_2_0.IN.t48 8.31073
R6574 VCO_C_0.INV_2_0.IN.n4 VCO_C_0.INV_2_0.IN.n22 7.05764
R6575 VCO_C_0.INV_2_0.IN.n3 VCO_C_0.INV_2_0.IN.t0 6.83153
R6576 VCO_C_0.INV_2_0.IN.n31 VCO_C_0.INV_2_0.IN.t14 6.78441
R6577 VCO_C_0.INV_2_0.IN VCO_C_0.INV_2_0.IN.n35 6.45366
R6578 VCO_C_0.INV_2_0.IN.n29 VCO_C_0.INV_2_0.IN.n28 6.20932
R6579 VCO_C_0.INV_2_0.IN.n21 VCO_C_0.INV_2_0.IN.t1 5.87174
R6580 VCO_C_0.INV_2_0.IN.n42 VCO_C_0.INV_2_0.IN.n41 5.28839
R6581 VCO_C_0.INV_2_0.IN.n68 VCO_C_0.INV_2_0.IN.n59 5.21368
R6582 VCO_C_0.INV_2_0.IN.n1 VCO_C_0.INV_2_0.IN.t15 4.92134
R6583 VCO_C_0.INV_2_0.IN.n60 VCO_C_0.INV_2_0.IN.t24 4.89657
R6584 VCO_C_0.INV_2_0.IN.n44 VCO_C_0.INV_2_0.IN.t26 4.89616
R6585 VCO_C_0.INV_2_0.IN.n73 VCO_C_0.INV_2_0.IN.n36 4.87698
R6586 VCO_C_0.INV_2_0.IN.n6 VCO_C_0.INV_2_0.IN.n57 4.63042
R6587 VCO_C_0.INV_2_0.IN.n70 VCO_C_0.INV_2_0.IN.n56 4.63037
R6588 VCO_C_0.INV_2_0.IN.n45 VCO_C_0.INV_2_0.IN.n1 4.22693
R6589 VCO_C_0.INV_2_0.IN VCO_C_0.INV_2_0.IN.n18 4.223
R6590 VCO_C_0.INV_2_0.IN.n46 VCO_C_0.INV_2_0.IN.n42 4.02972
R6591 VCO_C_0.INV_2_0.IN.n34 VCO_C_0.INV_2_0.IN.n33 4.0288
R6592 VCO_C_0.INV_2_0.IN.n74 VCO_C_0.INV_2_0.IN.n73 3.96222
R6593 VCO_C_0.INV_2_0.IN.t42 VCO_C_0.INV_2_0.IN.n13 3.6505
R6594 VCO_C_0.INV_2_0.IN.t49 VCO_C_0.INV_2_0.IN.n15 3.6505
R6595 VCO_C_0.INV_2_0.IN.n77 VCO_C_0.INV_2_0.IN.t18 3.6405
R6596 VCO_C_0.INV_2_0.IN.n77 VCO_C_0.INV_2_0.IN.n78 3.6405
R6597 VCO_C_0.INV_2_0.IN.n59 VCO_C_0.INV_2_0.IN.t17 3.6405
R6598 VCO_C_0.INV_2_0.IN.n59 VCO_C_0.INV_2_0.IN.n58 3.6405
R6599 VCO_C_0.INV_2_0.IN.n64 VCO_C_0.INV_2_0.IN.t25 3.6405
R6600 VCO_C_0.INV_2_0.IN.n64 VCO_C_0.INV_2_0.IN.n63 3.6405
R6601 VCO_C_0.INV_2_0.IN.n38 VCO_C_0.INV_2_0.IN.t21 3.6405
R6602 VCO_C_0.INV_2_0.IN.n38 VCO_C_0.INV_2_0.IN.n37 3.6405
R6603 VCO_C_0.INV_2_0.IN.n33 VCO_C_0.INV_2_0.IN.t13 3.6405
R6604 VCO_C_0.INV_2_0.IN.n33 VCO_C_0.INV_2_0.IN.n32 3.6405
R6605 VCO_C_0.INV_2_0.IN.n24 VCO_C_0.INV_2_0.IN.n23 3.47613
R6606 VCO_C_0.INV_2_0.IN.n20 VCO_C_0.INV_2_0.IN.n19 3.47609
R6607 VCO_C_0.INV_2_0.IN.n26 VCO_C_0.INV_2_0.IN.n25 3.47601
R6608 VCO_C_0.INV_2_0.IN.n21 VCO_C_0.INV_2_0.IN.n20 3.39857
R6609 VCO_C_0.INV_2_0.IN.n45 VCO_C_0.INV_2_0.IN.n76 3.27464
R6610 VCO_C_0.INV_2_0.IN.n18 VCO_C_0.INV_2_0.IN.n11 3.1807
R6611 VCO_C_0.INV_2_0.IN VCO_C_0.INV_2_0.IN.n75 3.16877
R6612 VCO_C_0.INV_2_0.IN.n26 VCO_C_0.INV_2_0.IN.t2 2.8627
R6613 VCO_C_0.INV_2_0.IN.n20 VCO_C_0.INV_2_0.IN.t3 2.86263
R6614 VCO_C_0.INV_2_0.IN.n24 VCO_C_0.INV_2_0.IN.t4 2.8626
R6615 VCO_C_0.INV_2_0.IN.n69 VCO_C_0.INV_2_0.IN.n68 2.60609
R6616 VCO_C_0.INV_2_0.IN.n4 VCO_C_0.INV_2_0.IN.n24 2.48343
R6617 VCO_C_0.INV_2_0.IN.n30 VCO_C_0.INV_2_0.IN 2.30073
R6618 VCO_C_0.INV_2_0.IN.n75 VCO_C_0.INV_2_0.IN 2.29178
R6619 VCO_C_0.INV_2_0.IN.n3 VCO_C_0.INV_2_0.IN.n27 2.24606
R6620 VCO_C_0.INV_2_0.IN.n6 VCO_C_0.INV_2_0.IN.n69 2.24505
R6621 VCO_C_0.INV_2_0.IN.n66 VCO_C_0.INV_2_0.IN.n65 3.77141
R6622 VCO_C_0.INV_2_0.IN.n67 VCO_C_0.INV_2_0.IN.n61 1.8072
R6623 VCO_C_0.INV_2_0.IN.n48 VCO_C_0.INV_2_0.IN.n40 1.76824
R6624 VCO_C_0.INV_2_0.IN.n65 VCO_C_0.INV_2_0.IN.n64 1.65829
R6625 VCO_C_0.INV_2_0.IN.n39 VCO_C_0.INV_2_0.IN.n38 1.65829
R6626 VCO_C_0.INV_2_0.IN.n55 VCO_C_0.INV_2_0.IN.n51 1.6131
R6627 VCO_C_0.INV_2_0.IN.n55 VCO_C_0.INV_2_0.IN.n54 1.57488
R6628 VCO_C_0.INV_2_0.IN.n44 VCO_C_0.INV_2_0.IN.n43 1.53436
R6629 VCO_C_0.INV_2_0.IN.n71 VCO_C_0.INV_2_0.IN.n70 1.51602
R6630 VCO_C_0.INV_2_0.IN.n47 VCO_C_0.INV_2_0.IN.t30 8.25008
R6631 VCO_C_0.INV_2_0.IN.n1 VCO_C_0.INV_2_0.IN.n44 2.52627
R6632 VCO_C_0.INV_2_0.IN.n61 VCO_C_0.INV_2_0.IN.n60 1.49487
R6633 VCO_C_0.INV_2_0.IN.n36 VCO_C_0.INV_2_0.IN.n34 1.32452
R6634 VCO_C_0.INV_2_0.IN.n76 VCO_C_0.INV_2_0.IN.n77 1.25757
R6635 VCO_C_0.INV_2_0.IN.n40 VCO_C_0.INV_2_0.IN.n39 1.12313
R6636 VCO_C_0.INV_2_0.IN.n3 VCO_C_0.INV_2_0.IN.n4 1.05601
R6637 VCO_C_0.INV_2_0.IN.n30 VCO_C_0.INV_2_0.IN.n29 1.01067
R6638 VCO_C_0.INV_2_0.IN.n50 VCO_C_0.INV_2_0.IN.n49 0.996664
R6639 VCO_C_0.INV_2_0.IN.n0 VCO_C_0.INV_2_0.IN.n5 0.992966
R6640 VCO_C_0.INV_2_0.IN.n4 VCO_C_0.INV_2_0.IN.n21 0.983287
R6641 VCO_C_0.INV_2_0.IN.n27 VCO_C_0.INV_2_0.IN.n26 0.982856
R6642 VCO_C_0.INV_2_0.IN.n2 VCO_C_0.INV_2_0.IN.n0 0.975705
R6643 VCO_C_0.INV_2_0.IN.n72 VCO_C_0.INV_2_0.IN.n71 0.968726
R6644 VCO_C_0.INV_2_0.IN.n73 VCO_C_0.INV_2_0.IN.n72 0.955885
R6645 VCO_C_0.INV_2_0.IN.n53 VCO_C_0.INV_2_0.IN.n52 0.953514
R6646 VCO_C_0.INV_2_0.IN.n29 VCO_C_0.INV_2_0.IN.n3 0.911933
R6647 VCO_C_0.INV_2_0.IN.n46 VCO_C_0.INV_2_0.IN.n45 0.856289
R6648 VCO_C_0.INV_2_0.IN.n48 VCO_C_0.INV_2_0.IN.n47 0.843442
R6649 VCO_C_0.INV_2_0.IN.n68 VCO_C_0.INV_2_0.IN.n67 0.8015
R6650 VCO_C_0.INV_2_0.IN.n70 VCO_C_0.INV_2_0.IN.n6 0.741046
R6651 VCO_C_0.INV_2_0.IN.n34 VCO_C_0.INV_2_0.IN.n31 0.710717
R6652 VCO_C_0.INV_2_0.IN.n71 VCO_C_0.INV_2_0.IN.n7 0.698938
R6653 VCO_C_0.INV_2_0.IN.n72 VCO_C_0.INV_2_0.IN.n48 0.656959
R6654 VCO_C_0.INV_2_0.IN.n47 VCO_C_0.INV_2_0.IN.n46 0.398395
R6655 VCO_C_0.INV_2_0.IN.n67 VCO_C_0.INV_2_0.IN.n66 0.3875
R6656 VCO_C_0.INV_2_0.IN.n54 VCO_C_0.INV_2_0.IN.n53 0.364199
R6657 VCO_C_0.INV_2_0.IN.n74 VCO_C_0.INV_2_0.IN.n30 0.362023
R6658 VCO_C_0.INV_2_0.IN.n7 VCO_C_0.INV_2_0.IN.n2 0.359267
R6659 VCO_C_0.INV_2_0.IN.n51 VCO_C_0.INV_2_0.IN.n50 0.323514
R6660 VCO_C_0.INV_2_0.IN.n5 VCO_C_0.INV_2_0.IN.n55 0.321048
R6661 VCO_C_0.INV_2_0.IN.n75 VCO_C_0.INV_2_0.IN.n74 0.271283
R6662 VCO_C_0.INV_2_0.IN.n36 VCO_C_0.INV_2_0.IN 0.147028
R6663 DFF_3_mag_0.INV_2_5.IN.n20 DFF_3_mag_0.INV_2_5.IN.t27 23.6945
R6664 DFF_3_mag_0.INV_2_5.IN.t20 DFF_3_mag_0.INV_2_5.IN.n21 23.6945
R6665 DFF_3_mag_0.INV_2_5.IN.n21 DFF_3_mag_0.INV_2_5.IN.n20 18.8035
R6666 DFF_3_mag_0.INV_2_5.IN.n18 DFF_3_mag_0.INV_2_5.IN.n16 15.8172
R6667 DFF_3_mag_0.INV_2_5.IN.n18 DFF_3_mag_0.INV_2_5.IN.n17 15.8172
R6668 DFF_3_mag_0.INV_2_5.IN.n17 DFF_3_mag_0.INV_2_5.IN.n13 15.8172
R6669 DFF_3_mag_0.INV_2_5.IN.n16 DFF_3_mag_0.INV_2_5.IN.t26 14.8925
R6670 DFF_3_mag_0.INV_2_5.IN.t22 DFF_3_mag_0.INV_2_5.IN.n18 14.8925
R6671 DFF_3_mag_0.INV_2_5.IN.n17 DFF_3_mag_0.INV_2_5.IN.t31 14.8925
R6672 DFF_3_mag_0.INV_2_5.IN.n22 DFF_3_mag_0.INV_2_5.IN.n14 12.2457
R6673 DFF_3_mag_0.INV_2_5.IN.n19 DFF_3_mag_0.INV_2_5.IN.n14 12.2457
R6674 DFF_3_mag_0.INV_2_5.IN.n19 DFF_3_mag_0.INV_2_5.IN.n15 12.2457
R6675 DFF_3_mag_0.INV_2_5.IN.n23 DFF_3_mag_0.INV_2_5.IN.t24 11.6285
R6676 DFF_3_mag_0.INV_2_5.IN.n15 DFF_3_mag_0.INV_2_5.IN.t27 8.9065
R6677 DFF_3_mag_0.INV_2_5.IN.t29 DFF_3_mag_0.INV_2_5.IN.n19 8.9065
R6678 DFF_3_mag_0.INV_2_5.IN.t30 DFF_3_mag_0.INV_2_5.IN.n14 8.9065
R6679 DFF_3_mag_0.INV_2_5.IN.n22 DFF_3_mag_0.INV_2_5.IN.t20 8.9065
R6680 DFF_3_mag_0.INV_2_5.IN.n18 DFF_3_mag_0.INV_2_5.IN.t23 8.6145
R6681 DFF_3_mag_0.INV_2_5.IN.n16 DFF_3_mag_0.INV_2_5.IN.t28 8.6145
R6682 DFF_3_mag_0.INV_2_5.IN.n17 DFF_3_mag_0.INV_2_5.IN.t21 8.6145
R6683 DFF_3_mag_0.INV_2_5.IN.n13 DFF_3_mag_0.INV_2_5.IN.t25 8.59715
R6684 DFF_3_mag_0.INV_2_5.IN.t26 DFF_3_mag_0.INV_2_5.IN.n15 8.3225
R6685 DFF_3_mag_0.INV_2_5.IN.n19 DFF_3_mag_0.INV_2_5.IN.t22 8.3225
R6686 DFF_3_mag_0.INV_2_5.IN.t31 DFF_3_mag_0.INV_2_5.IN.n14 8.3225
R6687 DFF_3_mag_0.INV_2_5.IN.t24 DFF_3_mag_0.INV_2_5.IN.n22 8.3225
R6688 DFF_3_mag_0.INV_2_5.IN.n24 DFF_3_mag_0.INV_2_5.IN.n12 5.24044
R6689 DFF_3_mag_0.INV_2_5.IN.n7 DFF_3_mag_0.INV_2_5.IN.n4 5.10151
R6690 DFF_3_mag_0.INV_2_5.IN.n9 DFF_3_mag_0.INV_2_5.IN.n3 5.10119
R6691 DFF_3_mag_0.INV_2_5.IN.n10 DFF_3_mag_0.INV_2_5.IN.n2 5.08021
R6692 DFF_3_mag_0.INV_2_5.IN.n7 DFF_3_mag_0.INV_2_5.IN.n6 4.66164
R6693 DFF_3_mag_0.INV_2_5.IN DFF_3_mag_0.INV_2_5.IN.n23 4.223
R6694 DFF_3_mag_0.INV_2_5.IN.n20 DFF_3_mag_0.INV_2_5.IN.t29 3.6505
R6695 DFF_3_mag_0.INV_2_5.IN.n21 DFF_3_mag_0.INV_2_5.IN.t30 3.6505
R6696 DFF_3_mag_0.INV_2_5.IN.n36 DFF_3_mag_0.INV_2_5.IN.t11 3.6405
R6697 DFF_3_mag_0.INV_2_5.IN.n36 DFF_3_mag_0.INV_2_5.IN.n35 3.6405
R6698 DFF_3_mag_0.INV_2_5.IN.n30 DFF_3_mag_0.INV_2_5.IN.t10 3.6405
R6699 DFF_3_mag_0.INV_2_5.IN.n30 DFF_3_mag_0.INV_2_5.IN.n29 3.6405
R6700 DFF_3_mag_0.INV_2_5.IN.n28 DFF_3_mag_0.INV_2_5.IN.t5 3.6405
R6701 DFF_3_mag_0.INV_2_5.IN.n28 DFF_3_mag_0.INV_2_5.IN.n27 3.6405
R6702 DFF_3_mag_0.INV_2_5.IN.n38 DFF_3_mag_0.INV_2_5.IN.t8 3.6405
R6703 DFF_3_mag_0.INV_2_5.IN.n38 DFF_3_mag_0.INV_2_5.IN.n37 3.6405
R6704 DFF_3_mag_0.INV_2_5.IN.n40 DFF_3_mag_0.INV_2_5.IN.n26 3.50463
R6705 DFF_3_mag_0.INV_2_5.IN.n34 DFF_3_mag_0.INV_2_5.IN.n33 3.50463
R6706 DFF_3_mag_0.INV_2_5.IN.n12 DFF_3_mag_0.INV_2_5.IN.t19 3.40711
R6707 DFF_3_mag_0.INV_2_5.IN.n26 DFF_3_mag_0.INV_2_5.IN.t15 3.2765
R6708 DFF_3_mag_0.INV_2_5.IN.n26 DFF_3_mag_0.INV_2_5.IN.n25 3.2765
R6709 DFF_3_mag_0.INV_2_5.IN.n33 DFF_3_mag_0.INV_2_5.IN.t16 3.2765
R6710 DFF_3_mag_0.INV_2_5.IN.n33 DFF_3_mag_0.INV_2_5.IN.n32 3.2765
R6711 DFF_3_mag_0.INV_2_5.IN.n23 DFF_3_mag_0.INV_2_5.IN.n13 3.1807
R6712 DFF_3_mag_0.INV_2_5.IN.n31 DFF_3_mag_0.INV_2_5.IN.n28 3.06224
R6713 DFF_3_mag_0.INV_2_5.IN.n39 DFF_3_mag_0.INV_2_5.IN.n36 3.06224
R6714 DFF_3_mag_0.INV_2_5.IN.n11 DFF_3_mag_0.INV_2_5.IN.n1 2.85093
R6715 DFF_3_mag_0.INV_2_5.IN.n31 DFF_3_mag_0.INV_2_5.IN.n30 2.6005
R6716 DFF_3_mag_0.INV_2_5.IN.n39 DFF_3_mag_0.INV_2_5.IN.n38 2.6005
R6717 DFF_3_mag_0.INV_2_5.IN.n8 DFF_3_mag_0.INV_2_5.IN 2.36593
R6718 DFF_3_mag_0.INV_2_5.IN.n1 DFF_3_mag_0.INV_2_5.IN.t17 2.16717
R6719 DFF_3_mag_0.INV_2_5.IN.n1 DFF_3_mag_0.INV_2_5.IN.n0 2.16717
R6720 DFF_3_mag_0.INV_2_5.IN.n24 DFF_3_mag_0.INV_2_5.IN 2.01183
R6721 DFF_3_mag_0.INV_2_5.IN.n6 DFF_3_mag_0.INV_2_5.IN.t3 1.9505
R6722 DFF_3_mag_0.INV_2_5.IN.n6 DFF_3_mag_0.INV_2_5.IN.n5 1.9505
R6723 DFF_3_mag_0.INV_2_5.IN.n12 DFF_3_mag_0.INV_2_5.IN.n11 1.0205
R6724 DFF_3_mag_0.INV_2_5.IN.n40 DFF_3_mag_0.INV_2_5.IN.n34 0.798761
R6725 DFF_3_mag_0.INV_2_5.IN.n11 DFF_3_mag_0.INV_2_5.IN.n10 0.644196
R6726 DFF_3_mag_0.INV_2_5.IN DFF_3_mag_0.INV_2_5.IN.n40 0.562022
R6727 DFF_3_mag_0.INV_2_5.IN.n10 DFF_3_mag_0.INV_2_5.IN.n9 0.450799
R6728 DFF_3_mag_0.INV_2_5.IN.n8 DFF_3_mag_0.INV_2_5.IN.n7 0.358456
R6729 DFF_3_mag_0.INV_2_5.IN DFF_3_mag_0.INV_2_5.IN.n24 0.278326
R6730 DFF_3_mag_0.INV_2_5.IN.n9 DFF_3_mag_0.INV_2_5.IN.n8 0.229792
R6731 DFF_3_mag_0.INV_2_5.IN.n34 DFF_3_mag_0.INV_2_5.IN.n31 0.18637
R6732 DFF_3_mag_0.INV_2_5.IN.n40 DFF_3_mag_0.INV_2_5.IN.n39 0.18637
R6733 OUT.n7 OUT.t26 23.6945
R6734 OUT.t24 OUT.n8 23.6945
R6735 OUT.n35 OUT.t35 23.6945
R6736 OUT.t13 OUT.n36 23.6945
R6737 OUT.n8 OUT.n7 18.8035
R6738 OUT.n36 OUT.n35 18.8035
R6739 OUT.n5 OUT.n3 15.8172
R6740 OUT.n4 OUT.n0 15.8172
R6741 OUT.n5 OUT.n4 15.8172
R6742 OUT.n33 OUT.n31 15.8172
R6743 OUT.n33 OUT.n32 15.8172
R6744 OUT.n32 OUT.n28 15.8172
R6745 OUT.n3 OUT.t17 14.8925
R6746 OUT.t30 OUT.n5 14.8925
R6747 OUT.n4 OUT.t18 14.8925
R6748 OUT.n31 OUT.t23 14.8925
R6749 OUT.t28 OUT.n33 14.8925
R6750 OUT.n32 OUT.t14 14.8925
R6751 OUT.n9 OUT.n1 12.2457
R6752 OUT.n6 OUT.n1 12.2457
R6753 OUT.n6 OUT.n2 12.2457
R6754 OUT.n37 OUT.n29 12.2457
R6755 OUT.n34 OUT.n29 12.2457
R6756 OUT.n34 OUT.n30 12.2457
R6757 OUT.n10 OUT.t12 11.6285
R6758 OUT.n38 OUT.t25 11.6285
R6759 OUT.n2 OUT.t26 8.9065
R6760 OUT.t15 OUT.n6 8.9065
R6761 OUT.t29 OUT.n1 8.9065
R6762 OUT.n9 OUT.t24 8.9065
R6763 OUT.n30 OUT.t35 8.9065
R6764 OUT.t16 OUT.n34 8.9065
R6765 OUT.t27 OUT.n29 8.9065
R6766 OUT.n37 OUT.t13 8.9065
R6767 OUT.n5 OUT.t31 8.6145
R6768 OUT.n3 OUT.t20 8.6145
R6769 OUT.n4 OUT.t21 8.6145
R6770 OUT.n33 OUT.t34 8.6145
R6771 OUT.n31 OUT.t32 8.6145
R6772 OUT.n32 OUT.t22 8.6145
R6773 OUT.n0 OUT.t19 8.59715
R6774 OUT.n28 OUT.t33 8.59715
R6775 OUT.t17 OUT.n2 8.3225
R6776 OUT.n6 OUT.t30 8.3225
R6777 OUT.t18 OUT.n1 8.3225
R6778 OUT.t12 OUT.n9 8.3225
R6779 OUT.t23 OUT.n30 8.3225
R6780 OUT.n34 OUT.t28 8.3225
R6781 OUT.t14 OUT.n29 8.3225
R6782 OUT.t25 OUT.n37 8.3225
R6783 OUT.n11 OUT 4.9636
R6784 OUT OUT.n10 4.223
R6785 OUT OUT.n38 4.223
R6786 OUT.n7 OUT.t15 3.6505
R6787 OUT.n8 OUT.t29 3.6505
R6788 OUT.n35 OUT.t16 3.6505
R6789 OUT.n36 OUT.t27 3.6505
R6790 OUT.n15 OUT.t10 3.6405
R6791 OUT.n15 OUT.n14 3.6405
R6792 OUT.n13 OUT.t5 3.6405
R6793 OUT.n13 OUT.n12 3.6405
R6794 OUT.n22 OUT.t2 3.6405
R6795 OUT.n22 OUT.n21 3.6405
R6796 OUT.n20 OUT.t7 3.6405
R6797 OUT.n20 OUT.n19 3.6405
R6798 OUT.n27 OUT.n18 3.50463
R6799 OUT.n26 OUT.n25 3.50463
R6800 OUT.n18 OUT.t3 3.2765
R6801 OUT.n18 OUT.n17 3.2765
R6802 OUT.n25 OUT.t4 3.2765
R6803 OUT.n25 OUT.n24 3.2765
R6804 OUT.n10 OUT.n0 3.1807
R6805 OUT.n38 OUT.n28 3.1807
R6806 OUT.n16 OUT.n13 3.06224
R6807 OUT.n23 OUT.n20 3.06224
R6808 OUT.n16 OUT.n15 2.6005
R6809 OUT.n23 OUT.n22 2.6005
R6810 OUT.n11 OUT 1.45743
R6811 OUT.n39 OUT 1.24006
R6812 OUT.n27 OUT.n26 0.798761
R6813 OUT.n40 OUT.n39 0.611422
R6814 OUT OUT.n27 0.562022
R6815 OUT.n39 OUT 0.247022
R6816 OUT.n40 OUT.n11 0.202264
R6817 OUT OUT.n40 0.19218
R6818 OUT.n27 OUT.n16 0.18637
R6819 OUT.n26 OUT.n23 0.18637
R6820 OUTB.n26 OUTB 6.6528
R6821 OUTB.n22 OUTB.n21 5.81586
R6822 OUTB.n18 OUTB.t6 5.10151
R6823 OUTB.n24 OUTB.t5 5.1005
R6824 OUTB.n23 OUTB.t0 5.08021
R6825 OUTB.n18 OUTB.n17 4.66164
R6826 OUTB.n3 OUTB.t12 3.6405
R6827 OUTB.n3 OUTB.n2 3.6405
R6828 OUTB.n5 OUTB.t9 3.6405
R6829 OUTB.n5 OUTB.n4 3.6405
R6830 OUTB.n10 OUTB.t11 3.6405
R6831 OUTB.n10 OUTB.n9 3.6405
R6832 OUTB.n12 OUTB.t8 3.6405
R6833 OUTB.n12 OUTB.n11 3.6405
R6834 OUTB.n15 OUTB.n1 3.50463
R6835 OUTB.n14 OUTB.n8 3.50463
R6836 OUTB.n1 OUTB.t17 3.2765
R6837 OUTB.n1 OUTB.n0 3.2765
R6838 OUTB.n8 OUTB.t16 3.2765
R6839 OUTB.n8 OUTB.n7 3.2765
R6840 OUTB.n6 OUTB.n5 3.06224
R6841 OUTB.n13 OUTB.n12 3.06224
R6842 OUTB.n22 OUTB.n20 2.85093
R6843 OUTB.n6 OUTB.n3 2.6005
R6844 OUTB.n13 OUTB.n10 2.6005
R6845 OUTB.n20 OUTB.t1 2.16717
R6846 OUTB.n20 OUTB.n19 2.16717
R6847 OUTB.n17 OUTB.t19 1.9505
R6848 OUTB.n17 OUTB.n16 1.9505
R6849 OUTB.n27 OUTB.n26 1.47848
R6850 OUTB.n26 OUTB 1.05814
R6851 OUTB.n15 OUTB.n14 0.798761
R6852 OUTB.n23 OUTB.n22 0.644196
R6853 OUTB OUTB.n15 0.562022
R6854 OUTB.n24 OUTB.n23 0.447229
R6855 OUTB.n25 OUTB.n18 0.308586
R6856 OUTB.n25 OUTB.n24 0.277162
R6857 OUTB.n15 OUTB.n6 0.18637
R6858 OUTB.n14 OUTB.n13 0.18637
R6859 OUTB.n27 OUTB 0.161224
R6860 OUTB OUTB.n25 0.115935
R6861 OUTB OUTB.n27 0.0483126
R6862 a_1424_1033.n86 a_1424_1033.n73 9.67588
R6863 a_1424_1033.n76 a_1424_1033.n75 3.74875
R6864 a_1424_1033.n3 a_1424_1033.n20 3.72928
R6865 a_1424_1033.n97 a_1424_1033.n95 3.71799
R6866 a_1424_1033.n1 a_1424_1033.n8 3.71559
R6867 a_1424_1033.n13 a_1424_1033.n12 3.71016
R6868 a_1424_1033.n26 a_1424_1033.t23 3.2765
R6869 a_1424_1033.n26 a_1424_1033.n25 3.2765
R6870 a_1424_1033.n28 a_1424_1033.t45 3.2765
R6871 a_1424_1033.n28 a_1424_1033.n27 3.2765
R6872 a_1424_1033.n93 a_1424_1033.t54 3.2765
R6873 a_1424_1033.n93 a_1424_1033.n92 3.2765
R6874 a_1424_1033.n30 a_1424_1033.t21 3.2765
R6875 a_1424_1033.n30 a_1424_1033.n29 3.2765
R6876 a_1424_1033.n54 a_1424_1033.t14 3.2765
R6877 a_1424_1033.n54 a_1424_1033.n53 3.2765
R6878 a_1424_1033.n51 a_1424_1033.t5 3.2765
R6879 a_1424_1033.n51 a_1424_1033.n50 3.2765
R6880 a_1424_1033.n47 a_1424_1033.t18 3.2765
R6881 a_1424_1033.n47 a_1424_1033.n46 3.2765
R6882 a_1424_1033.n44 a_1424_1033.t12 3.2765
R6883 a_1424_1033.n44 a_1424_1033.n43 3.2765
R6884 a_1424_1033.n40 a_1424_1033.t1 3.2765
R6885 a_1424_1033.n40 a_1424_1033.n39 3.2765
R6886 a_1424_1033.n71 a_1424_1033.t4 3.2765
R6887 a_1424_1033.n71 a_1424_1033.n70 3.2765
R6888 a_1424_1033.n68 a_1424_1033.t17 3.2765
R6889 a_1424_1033.n68 a_1424_1033.n67 3.2765
R6890 a_1424_1033.n64 a_1424_1033.t8 3.2765
R6891 a_1424_1033.n64 a_1424_1033.n63 3.2765
R6892 a_1424_1033.n61 a_1424_1033.t3 3.2765
R6893 a_1424_1033.n61 a_1424_1033.n60 3.2765
R6894 a_1424_1033.n57 a_1424_1033.t16 3.2765
R6895 a_1424_1033.n57 a_1424_1033.n56 3.2765
R6896 a_1424_1033.n83 a_1424_1033.t48 3.2765
R6897 a_1424_1033.n83 a_1424_1033.n82 3.2765
R6898 a_1424_1033.n90 a_1424_1033.t40 3.2765
R6899 a_1424_1033.n90 a_1424_1033.n89 3.2765
R6900 a_1424_1033.n17 a_1424_1033.t31 3.2765
R6901 a_1424_1033.n17 a_1424_1033.n16 3.2765
R6902 a_1424_1033.n15 a_1424_1033.t49 3.2765
R6903 a_1424_1033.n15 a_1424_1033.n14 3.2765
R6904 a_1424_1033.n10 a_1424_1033.t30 3.2765
R6905 a_1424_1033.n10 a_1424_1033.n9 3.2765
R6906 a_1424_1033.n8 a_1424_1033.t22 3.2765
R6907 a_1424_1033.n8 a_1424_1033.n7 3.2765
R6908 a_1424_1033.n32 a_1424_1033.t51 3.2765
R6909 a_1424_1033.n32 a_1424_1033.n31 3.2765
R6910 a_1424_1033.n35 a_1424_1033.t20 3.2765
R6911 a_1424_1033.n35 a_1424_1033.n34 3.2765
R6912 a_1424_1033.n78 a_1424_1033.t35 3.2765
R6913 a_1424_1033.n78 a_1424_1033.n77 3.2765
R6914 a_1424_1033.n75 a_1424_1033.t24 3.2765
R6915 a_1424_1033.n75 a_1424_1033.n74 3.2765
R6916 a_1424_1033.n22 a_1424_1033.t43 3.2765
R6917 a_1424_1033.n22 a_1424_1033.n21 3.2765
R6918 a_1424_1033.n12 a_1424_1033.t38 3.2765
R6919 a_1424_1033.n12 a_1424_1033.n11 3.2765
R6920 a_1424_1033.n80 a_1424_1033.t41 3.2765
R6921 a_1424_1033.n80 a_1424_1033.n79 3.2765
R6922 a_1424_1033.n37 a_1424_1033.t29 3.2765
R6923 a_1424_1033.n37 a_1424_1033.n36 3.2765
R6924 a_1424_1033.n20 a_1424_1033.t42 3.2765
R6925 a_1424_1033.n20 a_1424_1033.n19 3.2765
R6926 a_1424_1033.t58 a_1424_1033.n97 3.2765
R6927 a_1424_1033.n97 a_1424_1033.n96 3.2765
R6928 a_1424_1033.n58 a_1424_1033.n57 3.1505
R6929 a_1424_1033.n62 a_1424_1033.n61 3.1505
R6930 a_1424_1033.n65 a_1424_1033.n64 3.1505
R6931 a_1424_1033.n69 a_1424_1033.n68 3.1505
R6932 a_1424_1033.n72 a_1424_1033.n71 3.1505
R6933 a_1424_1033.n41 a_1424_1033.n40 3.1505
R6934 a_1424_1033.n45 a_1424_1033.n44 3.1505
R6935 a_1424_1033.n48 a_1424_1033.n47 3.1505
R6936 a_1424_1033.n52 a_1424_1033.n51 3.1505
R6937 a_1424_1033.n55 a_1424_1033.n54 3.1505
R6938 a_1424_1033.n81 a_1424_1033.n80 3.1505
R6939 a_1424_1033.n38 a_1424_1033.n37 3.1505
R6940 a_1424_1033.n33 a_1424_1033.n32 3.1505
R6941 a_1424_1033.n18 a_1424_1033.n17 3.1505
R6942 a_1424_1033.n84 a_1424_1033.n83 3.1505
R6943 a_1424_1033.n88 a_1424_1033.n30 3.1505
R6944 a_1424_1033.n94 a_1424_1033.n28 3.1505
R6945 a_1424_1033.n5 a_1424_1033.n22 4.10259
R6946 a_1424_1033.n5 a_1424_1033.n13 2.24345
R6947 a_1424_1033.n2 a_1424_1033.n1 2.24324
R6948 a_1424_1033.n4 a_1424_1033.n91 2.10504
R6949 a_1424_1033.n3 a_1424_1033.n15 1.8475
R6950 a_1424_1033.n4 a_1424_1033.n93 1.84743
R6951 a_1424_1033.n76 a_1424_1033.n78 1.84737
R6952 a_1424_1033.n91 a_1424_1033.n90 3.35151
R6953 a_1424_1033.n1 a_1424_1033.n10 1.87597
R6954 a_1424_1033.n0 a_1424_1033.n35 1.84728
R6955 a_1424_1033.n6 a_1424_1033.n26 1.84618
R6956 a_1424_1033.n6 a_1424_1033.n24 1.69983
R6957 a_1424_1033.n5 a_1424_1033.n3 1.48093
R6958 a_1424_1033.n85 a_1424_1033.n84 0.899822
R6959 a_1424_1033.n88 a_1424_1033.n87 0.899822
R6960 a_1424_1033.n65 a_1424_1033.n62 0.758798
R6961 a_1424_1033.n48 a_1424_1033.n45 0.758798
R6962 a_1424_1033.n73 a_1424_1033.n55 0.724996
R6963 a_1424_1033.n72 a_1424_1033.n69 0.7205
R6964 a_1424_1033.n55 a_1424_1033.n52 0.7205
R6965 a_1424_1033.n73 a_1424_1033.n72 0.636952
R6966 a_1424_1033.n6 a_1424_1033.n94 0.622339
R6967 a_1424_1033.n3 a_1424_1033.n18 0.618999
R6968 a_1424_1033.n4 a_1424_1033.n88 0.610699
R6969 a_1424_1033.n38 a_1424_1033.n0 0.607127
R6970 a_1424_1033.n81 a_1424_1033.n76 0.604163
R6971 a_1424_1033.n0 a_1424_1033.n33 0.59579
R6972 a_1424_1033.n94 a_1424_1033.n4 0.593116
R6973 a_1424_1033.n2 a_1424_1033.n23 0.566952
R6974 a_1424_1033.n59 a_1424_1033.n58 0.555819
R6975 a_1424_1033.n42 a_1424_1033.n41 0.555819
R6976 a_1424_1033.n69 a_1424_1033.n66 0.551989
R6977 a_1424_1033.n52 a_1424_1033.n49 0.551989
R6978 a_1424_1033.n87 a_1424_1033.n86 0.3917
R6979 a_1424_1033.n66 a_1424_1033.n65 0.283904
R6980 a_1424_1033.n49 a_1424_1033.n48 0.283904
R6981 a_1424_1033.n62 a_1424_1033.n59 0.280074
R6982 a_1424_1033.n45 a_1424_1033.n42 0.280074
R6983 a_1424_1033.n86 a_1424_1033.n85 0.2621
R6984 a_1424_1033.n85 a_1424_1033.n81 0.247022
R6985 a_1424_1033.n87 a_1424_1033.n38 0.247022
R6986 a_1424_1033.n95 a_1424_1033.n6 0.0460206
R6987 a_1424_1033.n24 a_1424_1033.n2 0.0425768
R6988 a_1424_1033.n23 a_1424_1033.n5 0.0408697
R6989 DFF_3_mag_0.INV_2_4.OUT.n18 DFF_3_mag_0.INV_2_4.OUT.t3 5.81586
R6990 DFF_3_mag_0.INV_2_4.OUT.n26 DFF_3_mag_0.INV_2_4.OUT.n23 5.10148
R6991 DFF_3_mag_0.INV_2_4.OUT.n22 DFF_3_mag_0.INV_2_4.OUT.n21 5.10116
R6992 DFF_3_mag_0.INV_2_4.OUT.n20 DFF_3_mag_0.INV_2_4.OUT.n19 5.08021
R6993 DFF_3_mag_0.INV_2_4.OUT.n26 DFF_3_mag_0.INV_2_4.OUT.n25 4.66166
R6994 DFF_3_mag_0.INV_2_4.OUT.n10 DFF_3_mag_0.INV_2_4.OUT.t7 3.6405
R6995 DFF_3_mag_0.INV_2_4.OUT.n10 DFF_3_mag_0.INV_2_4.OUT.n9 3.6405
R6996 DFF_3_mag_0.INV_2_4.OUT.n3 DFF_3_mag_0.INV_2_4.OUT.t5 3.6405
R6997 DFF_3_mag_0.INV_2_4.OUT.n3 DFF_3_mag_0.INV_2_4.OUT.n2 3.6405
R6998 DFF_3_mag_0.INV_2_4.OUT.n5 DFF_3_mag_0.INV_2_4.OUT.t9 3.6405
R6999 DFF_3_mag_0.INV_2_4.OUT.n5 DFF_3_mag_0.INV_2_4.OUT.n4 3.6405
R7000 DFF_3_mag_0.INV_2_4.OUT.n12 DFF_3_mag_0.INV_2_4.OUT.t11 3.6405
R7001 DFF_3_mag_0.INV_2_4.OUT.n12 DFF_3_mag_0.INV_2_4.OUT.n11 3.6405
R7002 DFF_3_mag_0.INV_2_4.OUT.n14 DFF_3_mag_0.INV_2_4.OUT.n8 3.50463
R7003 DFF_3_mag_0.INV_2_4.OUT.n15 DFF_3_mag_0.INV_2_4.OUT.n1 3.50463
R7004 DFF_3_mag_0.INV_2_4.OUT.n8 DFF_3_mag_0.INV_2_4.OUT.t13 3.2765
R7005 DFF_3_mag_0.INV_2_4.OUT.n8 DFF_3_mag_0.INV_2_4.OUT.n7 3.2765
R7006 DFF_3_mag_0.INV_2_4.OUT.n1 DFF_3_mag_0.INV_2_4.OUT.t12 3.2765
R7007 DFF_3_mag_0.INV_2_4.OUT.n1 DFF_3_mag_0.INV_2_4.OUT.n0 3.2765
R7008 DFF_3_mag_0.INV_2_4.OUT.n6 DFF_3_mag_0.INV_2_4.OUT.n5 3.06224
R7009 DFF_3_mag_0.INV_2_4.OUT.n13 DFF_3_mag_0.INV_2_4.OUT.n12 3.06224
R7010 DFF_3_mag_0.INV_2_4.OUT.n18 DFF_3_mag_0.INV_2_4.OUT.n17 2.85093
R7011 DFF_3_mag_0.INV_2_4.OUT.n6 DFF_3_mag_0.INV_2_4.OUT.n3 2.6005
R7012 DFF_3_mag_0.INV_2_4.OUT.n13 DFF_3_mag_0.INV_2_4.OUT.n10 2.6005
R7013 DFF_3_mag_0.INV_2_4.OUT DFF_3_mag_0.INV_2_4.OUT.n27 2.36593
R7014 DFF_3_mag_0.INV_2_4.OUT.n17 DFF_3_mag_0.INV_2_4.OUT.t17 2.16717
R7015 DFF_3_mag_0.INV_2_4.OUT.n17 DFF_3_mag_0.INV_2_4.OUT.n16 2.16717
R7016 DFF_3_mag_0.INV_2_4.OUT.n25 DFF_3_mag_0.INV_2_4.OUT.t19 1.9505
R7017 DFF_3_mag_0.INV_2_4.OUT.n25 DFF_3_mag_0.INV_2_4.OUT.n24 1.9505
R7018 DFF_3_mag_0.INV_2_4.OUT.n15 DFF_3_mag_0.INV_2_4.OUT.n14 0.798761
R7019 DFF_3_mag_0.INV_2_4.OUT.n20 DFF_3_mag_0.INV_2_4.OUT.n18 0.644196
R7020 DFF_3_mag_0.INV_2_4.OUT DFF_3_mag_0.INV_2_4.OUT.n15 0.562022
R7021 DFF_3_mag_0.INV_2_4.OUT.n22 DFF_3_mag_0.INV_2_4.OUT.n20 0.450839
R7022 DFF_3_mag_0.INV_2_4.OUT.n27 DFF_3_mag_0.INV_2_4.OUT.n26 0.358498
R7023 DFF_3_mag_0.INV_2_4.OUT.n27 DFF_3_mag_0.INV_2_4.OUT.n22 0.229792
R7024 DFF_3_mag_0.INV_2_4.OUT.n15 DFF_3_mag_0.INV_2_4.OUT.n6 0.18637
R7025 DFF_3_mag_0.INV_2_4.OUT.n14 DFF_3_mag_0.INV_2_4.OUT.n13 0.18637
R7026 DFF_3_mag_0.INV_2_3.IN.n7 DFF_3_mag_0.INV_2_3.IN.t17 23.6945
R7027 DFF_3_mag_0.INV_2_3.IN.n8 DFF_3_mag_0.INV_2_3.IN.t16 23.6945
R7028 DFF_3_mag_0.INV_2_3.IN.n8 DFF_3_mag_0.INV_2_3.IN.n7 18.8035
R7029 DFF_3_mag_0.INV_2_3.IN.n5 DFF_3_mag_0.INV_2_3.IN.n2 15.8172
R7030 DFF_3_mag_0.INV_2_3.IN.n11 DFF_3_mag_0.INV_2_3.IN.n10 15.8172
R7031 DFF_3_mag_0.INV_2_3.IN.n10 DFF_3_mag_0.INV_2_3.IN.n2 15.8172
R7032 DFF_3_mag_0.INV_2_3.IN.t22 DFF_3_mag_0.INV_2_3.IN.n5 14.8925
R7033 DFF_3_mag_0.INV_2_3.IN.t18 DFF_3_mag_0.INV_2_3.IN.n2 14.8925
R7034 DFF_3_mag_0.INV_2_3.IN.n10 DFF_3_mag_0.INV_2_3.IN.t25 14.8925
R7035 DFF_3_mag_0.INV_2_3.IN.n9 DFF_3_mag_0.INV_2_3.IN.n3 12.2457
R7036 DFF_3_mag_0.INV_2_3.IN.n9 DFF_3_mag_0.INV_2_3.IN.n4 12.2457
R7037 DFF_3_mag_0.INV_2_3.IN.n6 DFF_3_mag_0.INV_2_3.IN.n4 12.2457
R7038 DFF_3_mag_0.INV_2_3.IN.n12 DFF_3_mag_0.INV_2_3.IN.t21 11.6285
R7039 DFF_3_mag_0.INV_2_3.IN.t17 DFF_3_mag_0.INV_2_3.IN.n6 8.9065
R7040 DFF_3_mag_0.INV_2_3.IN.t24 DFF_3_mag_0.INV_2_3.IN.n4 8.9065
R7041 DFF_3_mag_0.INV_2_3.IN.n9 DFF_3_mag_0.INV_2_3.IN.t19 8.9065
R7042 DFF_3_mag_0.INV_2_3.IN.t16 DFF_3_mag_0.INV_2_3.IN.n3 8.9065
R7043 DFF_3_mag_0.INV_2_3.IN.n5 DFF_3_mag_0.INV_2_3.IN.t26 8.6145
R7044 DFF_3_mag_0.INV_2_3.IN.n2 DFF_3_mag_0.INV_2_3.IN.t20 8.6145
R7045 DFF_3_mag_0.INV_2_3.IN.n10 DFF_3_mag_0.INV_2_3.IN.t27 8.6145
R7046 DFF_3_mag_0.INV_2_3.IN.n11 DFF_3_mag_0.INV_2_3.IN.t23 8.59715
R7047 DFF_3_mag_0.INV_2_3.IN.n6 DFF_3_mag_0.INV_2_3.IN.t22 8.3225
R7048 DFF_3_mag_0.INV_2_3.IN.n4 DFF_3_mag_0.INV_2_3.IN.t18 8.3225
R7049 DFF_3_mag_0.INV_2_3.IN.t25 DFF_3_mag_0.INV_2_3.IN.n9 8.3225
R7050 DFF_3_mag_0.INV_2_3.IN.n3 DFF_3_mag_0.INV_2_3.IN.t21 8.3225
R7051 DFF_3_mag_0.INV_2_3.IN.n1 DFF_3_mag_0.INV_2_3.IN.t1 6.74388
R7052 DFF_3_mag_0.INV_2_3.IN.n0 DFF_3_mag_0.INV_2_3.IN.t4 6.74332
R7053 DFF_3_mag_0.INV_2_3.IN.n0 DFF_3_mag_0.INV_2_3.IN.t5 5.1005
R7054 DFF_3_mag_0.INV_2_3.IN.n1 DFF_3_mag_0.INV_2_3.IN.t0 5.1005
R7055 DFF_3_mag_0.INV_2_3.IN DFF_3_mag_0.INV_2_3.IN.n12 4.223
R7056 DFF_3_mag_0.INV_2_3.IN.n7 DFF_3_mag_0.INV_2_3.IN.t24 3.6505
R7057 DFF_3_mag_0.INV_2_3.IN.t19 DFF_3_mag_0.INV_2_3.IN.n8 3.6505
R7058 DFF_3_mag_0.INV_2_3.IN.n19 DFF_3_mag_0.INV_2_3.IN.n16 3.57508
R7059 DFF_3_mag_0.INV_2_3.IN.n28 DFF_3_mag_0.INV_2_3.IN.n27 3.5743
R7060 DFF_3_mag_0.INV_2_3.IN.n0 DFF_3_mag_0.INV_2_3.IN.n13 3.40011
R7061 DFF_3_mag_0.INV_2_3.IN.n1 DFF_3_mag_0.INV_2_3.IN.n22 3.40001
R7062 DFF_3_mag_0.INV_2_3.IN.n12 DFF_3_mag_0.INV_2_3.IN.n11 3.1807
R7063 DFF_3_mag_0.INV_2_3.IN.n14 DFF_3_mag_0.INV_2_3.IN.t6 3.00158
R7064 DFF_3_mag_0.INV_2_3.IN.n23 DFF_3_mag_0.INV_2_3.IN.t3 3.00077
R7065 DFF_3_mag_0.INV_2_3.IN DFF_3_mag_0.INV_2_3.IN.n20 2.58112
R7066 DFF_3_mag_0.INV_2_3.IN DFF_3_mag_0.INV_2_3.IN.n29 2.58112
R7067 DFF_3_mag_0.INV_2_3.IN.n18 DFF_3_mag_0.INV_2_3.IN.t9 2.16717
R7068 DFF_3_mag_0.INV_2_3.IN.n18 DFF_3_mag_0.INV_2_3.IN.n17 2.16717
R7069 DFF_3_mag_0.INV_2_3.IN.n16 DFF_3_mag_0.INV_2_3.IN.t11 2.16717
R7070 DFF_3_mag_0.INV_2_3.IN.n16 DFF_3_mag_0.INV_2_3.IN.n15 2.16717
R7071 DFF_3_mag_0.INV_2_3.IN.n25 DFF_3_mag_0.INV_2_3.IN.t7 2.16717
R7072 DFF_3_mag_0.INV_2_3.IN.n25 DFF_3_mag_0.INV_2_3.IN.n24 2.16717
R7073 DFF_3_mag_0.INV_2_3.IN.n27 DFF_3_mag_0.INV_2_3.IN.t14 2.16717
R7074 DFF_3_mag_0.INV_2_3.IN.n27 DFF_3_mag_0.INV_2_3.IN.n26 2.16717
R7075 DFF_3_mag_0.INV_2_3.IN.n20 DFF_3_mag_0.INV_2_3.IN.n14 1.84821
R7076 DFF_3_mag_0.INV_2_3.IN.n29 DFF_3_mag_0.INV_2_3.IN.n23 1.84769
R7077 DFF_3_mag_0.INV_2_3.IN.n19 DFF_3_mag_0.INV_2_3.IN.n18 1.25233
R7078 DFF_3_mag_0.INV_2_3.IN.n28 DFF_3_mag_0.INV_2_3.IN.n25 1.25225
R7079 DFF_3_mag_0.INV_2_3.IN.n29 DFF_3_mag_0.INV_2_3.IN.n28 1.12575
R7080 DFF_3_mag_0.INV_2_3.IN.n20 DFF_3_mag_0.INV_2_3.IN.n19 1.12554
R7081 DFF_3_mag_0.INV_2_3.IN DFF_3_mag_0.INV_2_3.IN.n21 0.784521
R7082 DFF_3_mag_0.INV_2_3.IN.n21 DFF_3_mag_0.INV_2_3.IN 0.689881
R7083 DFF_3_mag_0.INV_2_3.IN.n23 DFF_3_mag_0.INV_2_3.IN.n1 0.559952
R7084 DFF_3_mag_0.INV_2_3.IN.n14 DFF_3_mag_0.INV_2_3.IN.n0 0.558372
R7085 DFF_3_mag_0.INV_2_3.IN.n21 DFF_3_mag_0.INV_2_3.IN 0.25925
R7086 a_17597_2884.n5 a_17597_2884.t9 29.3691
R7087 a_17597_2884.n6 a_17597_2884.n5 21.9292
R7088 a_17597_2884.n7 a_17597_2884.n6 18.1271
R7089 a_17597_2884.n7 a_17597_2884.t6 11.2425
R7090 a_17597_2884.n3 a_17597_2884.t0 10.2135
R7091 a_17597_2884.n5 a_17597_2884.t7 6.1325
R7092 a_17597_2884.n6 a_17597_2884.t8 6.1325
R7093 a_17597_2884.n3 a_17597_2884.n2 4.68398
R7094 a_17597_2884.n8 a_17597_2884.n7 4.6302
R7095 a_17597_2884.n9 a_17597_2884.n8 2.85093
R7096 a_17597_2884.n1 a_17597_2884.t4 2.16717
R7097 a_17597_2884.n1 a_17597_2884.n0 2.16717
R7098 a_17597_2884.n9 a_17597_2884.t5 2.16717
R7099 a_17597_2884.n10 a_17597_2884.n9 2.16717
R7100 a_17597_2884.n4 a_17597_2884.n3 1.58582
R7101 a_17597_2884.n4 a_17597_2884.n1 1.24371
R7102 a_17597_2884.n8 a_17597_2884.n4 0.971051
R7103 a_20434_3437.n3 a_20434_3437.t8 29.3691
R7104 a_20434_3437.n4 a_20434_3437.n3 21.9292
R7105 a_20434_3437.n5 a_20434_3437.n4 18.1271
R7106 a_20434_3437.n5 a_20434_3437.t9 11.2425
R7107 a_20434_3437.n8 a_20434_3437.n7 10.1038
R7108 a_20434_3437.n3 a_20434_3437.t7 6.1325
R7109 a_20434_3437.n4 a_20434_3437.t6 6.1325
R7110 a_20434_3437.n8 a_20434_3437.t4 4.70149
R7111 a_20434_3437.n6 a_20434_3437.n5 4.6302
R7112 a_20434_3437.n6 a_20434_3437.n2 2.85093
R7113 a_20434_3437.n2 a_20434_3437.t1 2.16717
R7114 a_20434_3437.n2 a_20434_3437.n1 2.16717
R7115 a_20434_3437.t3 a_20434_3437.n10 2.16717
R7116 a_20434_3437.n10 a_20434_3437.n0 2.16717
R7117 a_20434_3437.n9 a_20434_3437.n8 1.58618
R7118 a_20434_3437.n10 a_20434_3437.n9 1.24388
R7119 a_20434_3437.n9 a_20434_3437.n6 0.97169
R7120 a_20434_1083.n2 a_20434_1083.t6 29.2961
R7121 a_20434_1083.n3 a_20434_1083.n2 21.9292
R7122 a_20434_1083.n4 a_20434_1083.n3 18.1271
R7123 a_20434_1083.n4 a_20434_1083.t7 11.1695
R7124 a_20434_1083.n2 a_20434_1083.t9 6.1325
R7125 a_20434_1083.n3 a_20434_1083.t8 6.1325
R7126 a_20434_1083.n7 a_20434_1083.n6 4.93252
R7127 a_20434_1083.n7 a_20434_1083.t0 4.70348
R7128 a_20434_1083.n5 a_20434_1083.n4 4.6311
R7129 a_20434_1083.n5 a_20434_1083.n1 2.85093
R7130 a_20434_1083.n1 a_20434_1083.t2 2.16717
R7131 a_20434_1083.n1 a_20434_1083.n0 2.16717
R7132 a_20434_1083.n9 a_20434_1083.t4 2.16717
R7133 a_20434_1083.n10 a_20434_1083.n9 2.16717
R7134 a_20434_1083.n8 a_20434_1083.n7 1.58583
R7135 a_20434_1083.n9 a_20434_1083.n8 1.24398
R7136 a_20434_1083.n8 a_20434_1083.n5 0.971047
R7137 DFF_3_mag_0.INV_2_0.OUT.n26 DFF_3_mag_0.INV_2_0.OUT.t22 45.6363
R7138 DFF_3_mag_0.INV_2_0.OUT.n22 DFF_3_mag_0.INV_2_0.OUT.t26 45.6363
R7139 DFF_3_mag_0.INV_2_0.OUT.n17 DFF_3_mag_0.INV_2_0.OUT.t19 29.6446
R7140 DFF_3_mag_0.INV_2_0.OUT.t14 DFF_3_mag_0.INV_2_0.OUT.n18 29.6446
R7141 DFF_3_mag_0.INV_2_0.OUT.n19 DFF_3_mag_0.INV_2_0.OUT.t15 29.6446
R7142 DFF_3_mag_0.INV_2_0.OUT.t13 DFF_3_mag_0.INV_2_0.OUT.n20 29.6446
R7143 DFF_3_mag_0.INV_2_0.OUT.n16 DFF_3_mag_0.INV_2_0.OUT.t16 24.6117
R7144 DFF_3_mag_0.INV_2_0.OUT.n21 DFF_3_mag_0.INV_2_0.OUT.t28 24.6117
R7145 DFF_3_mag_0.INV_2_0.OUT.n18 DFF_3_mag_0.INV_2_0.OUT.n17 22.2047
R7146 DFF_3_mag_0.INV_2_0.OUT.n20 DFF_3_mag_0.INV_2_0.OUT.n19 22.2047
R7147 DFF_3_mag_0.INV_2_0.OUT.t22 DFF_3_mag_0.INV_2_0.OUT.t12 22.1925
R7148 DFF_3_mag_0.INV_2_0.OUT.t26 DFF_3_mag_0.INV_2_0.OUT.t21 22.1925
R7149 DFF_3_mag_0.INV_2_0.OUT DFF_3_mag_0.INV_2_0.OUT.t14 21.8613
R7150 DFF_3_mag_0.INV_2_0.OUT.n27 DFF_3_mag_0.INV_2_0.OUT.n26 20.9314
R7151 DFF_3_mag_0.INV_2_0.OUT.n23 DFF_3_mag_0.INV_2_0.OUT.n22 20.9314
R7152 DFF_3_mag_0.INV_2_0.OUT.n25 DFF_3_mag_0.INV_2_0.OUT.t13 17.8613
R7153 DFF_3_mag_0.INV_2_0.OUT DFF_3_mag_0.INV_2_0.OUT.n28 10.8592
R7154 DFF_3_mag_0.INV_2_0.OUT DFF_3_mag_0.INV_2_0.OUT.n25 8.94379
R7155 DFF_3_mag_0.INV_2_0.OUT DFF_3_mag_0.INV_2_0.OUT.n16 8.87094
R7156 DFF_3_mag_0.INV_2_0.OUT.n26 DFF_3_mag_0.INV_2_0.OUT.t27 6.1325
R7157 DFF_3_mag_0.INV_2_0.OUT.n27 DFF_3_mag_0.INV_2_0.OUT.t30 6.1325
R7158 DFF_3_mag_0.INV_2_0.OUT.n17 DFF_3_mag_0.INV_2_0.OUT.t31 6.1325
R7159 DFF_3_mag_0.INV_2_0.OUT.n18 DFF_3_mag_0.INV_2_0.OUT.t25 6.1325
R7160 DFF_3_mag_0.INV_2_0.OUT.n16 DFF_3_mag_0.INV_2_0.OUT.t18 6.1325
R7161 DFF_3_mag_0.INV_2_0.OUT.n19 DFF_3_mag_0.INV_2_0.OUT.t20 6.1325
R7162 DFF_3_mag_0.INV_2_0.OUT.n20 DFF_3_mag_0.INV_2_0.OUT.t23 6.1325
R7163 DFF_3_mag_0.INV_2_0.OUT.n21 DFF_3_mag_0.INV_2_0.OUT.t17 6.1325
R7164 DFF_3_mag_0.INV_2_0.OUT.n22 DFF_3_mag_0.INV_2_0.OUT.t29 6.1325
R7165 DFF_3_mag_0.INV_2_0.OUT.n23 DFF_3_mag_0.INV_2_0.OUT.t24 6.1325
R7166 DFF_3_mag_0.INV_2_0.OUT.n24 DFF_3_mag_0.INV_2_0.OUT.n23 5.38991
R7167 DFF_3_mag_0.INV_2_0.OUT.n28 DFF_3_mag_0.INV_2_0.OUT.n27 5.12094
R7168 DFF_3_mag_0.INV_2_0.OUT.n24 DFF_3_mag_0.INV_2_0.OUT.n21 4.83094
R7169 DFF_3_mag_0.INV_2_0.OUT.n11 DFF_3_mag_0.INV_2_0.OUT.t3 3.6405
R7170 DFF_3_mag_0.INV_2_0.OUT.n11 DFF_3_mag_0.INV_2_0.OUT.n10 3.6405
R7171 DFF_3_mag_0.INV_2_0.OUT.n5 DFF_3_mag_0.INV_2_0.OUT.t1 3.6405
R7172 DFF_3_mag_0.INV_2_0.OUT.n5 DFF_3_mag_0.INV_2_0.OUT.n4 3.6405
R7173 DFF_3_mag_0.INV_2_0.OUT.n7 DFF_3_mag_0.INV_2_0.OUT.t5 3.6405
R7174 DFF_3_mag_0.INV_2_0.OUT.n7 DFF_3_mag_0.INV_2_0.OUT.n6 3.6405
R7175 DFF_3_mag_0.INV_2_0.OUT.n13 DFF_3_mag_0.INV_2_0.OUT.t7 3.6405
R7176 DFF_3_mag_0.INV_2_0.OUT.n13 DFF_3_mag_0.INV_2_0.OUT.n12 3.6405
R7177 DFF_3_mag_0.INV_2_0.OUT.n15 DFF_3_mag_0.INV_2_0.OUT.n1 3.50463
R7178 DFF_3_mag_0.INV_2_0.OUT.n9 DFF_3_mag_0.INV_2_0.OUT.n3 3.50463
R7179 DFF_3_mag_0.INV_2_0.OUT.n1 DFF_3_mag_0.INV_2_0.OUT.t9 3.2765
R7180 DFF_3_mag_0.INV_2_0.OUT.n1 DFF_3_mag_0.INV_2_0.OUT.n0 3.2765
R7181 DFF_3_mag_0.INV_2_0.OUT.n3 DFF_3_mag_0.INV_2_0.OUT.t8 3.2765
R7182 DFF_3_mag_0.INV_2_0.OUT.n3 DFF_3_mag_0.INV_2_0.OUT.n2 3.2765
R7183 DFF_3_mag_0.INV_2_0.OUT.n8 DFF_3_mag_0.INV_2_0.OUT.n7 3.06224
R7184 DFF_3_mag_0.INV_2_0.OUT.n14 DFF_3_mag_0.INV_2_0.OUT.n13 3.06224
R7185 DFF_3_mag_0.INV_2_0.OUT.n8 DFF_3_mag_0.INV_2_0.OUT.n5 2.6005
R7186 DFF_3_mag_0.INV_2_0.OUT.n14 DFF_3_mag_0.INV_2_0.OUT.n11 2.6005
R7187 DFF_3_mag_0.INV_2_0.OUT.n28 DFF_3_mag_0.INV_2_0.OUT 1.07267
R7188 DFF_3_mag_0.INV_2_0.OUT.n15 DFF_3_mag_0.INV_2_0.OUT.n9 0.798761
R7189 DFF_3_mag_0.INV_2_0.OUT DFF_3_mag_0.INV_2_0.OUT.n24 0.658318
R7190 DFF_3_mag_0.INV_2_0.OUT.n25 DFF_3_mag_0.INV_2_0.OUT 0.628846
R7191 DFF_3_mag_0.INV_2_0.OUT DFF_3_mag_0.INV_2_0.OUT.n15 0.562022
R7192 DFF_3_mag_0.INV_2_0.OUT.n9 DFF_3_mag_0.INV_2_0.OUT.n8 0.18637
R7193 DFF_3_mag_0.INV_2_0.OUT.n15 DFF_3_mag_0.INV_2_0.OUT.n14 0.18637
C0 VCO_C_0.INV_2_2.IN VCO_C_0.OUTB 0.0179f
C1 VCO_C_0.INV_2_0.IN m1_5752_3074# 0.103f
C2 VCO_C_0.OUTB DFF_3_mag_0.INV_2_0.OUT 0.703f
C3 DFF_3_mag_0.INV_2_0.OUT DFF_3_mag_0.INV_2_4.OUT 0.488f
C4 VCTRL VCO_C_0.OUTB 0.0222f
C5 VCO_C_0.INV_2_5.IN m1_5752_3074# 0.00112f
C6 VCO_C_0.INV_2_3.IN VCO_C_0.OUTB 0.348f
C7 VCO_C_0.INV_2_4.IN VCO_C_0.OUTB 0.00204f
C8 VCO_C_0.OUTB OUTB 0.725f
C9 DFF_3_mag_0.INV_2_3.IN DFF_3_mag_0.INV_2_5.IN 1.21f
C10 VDD VCO_C_0.INV_2_0.IN 14.8f
C11 DFF_3_mag_0.INV_2_5.IN DFF_3_mag_0.INV_2_5.OUT 0.381f
C12 VDD VCO_C_0.INV_2_1.IN 2.15f
C13 VCO_C_0.INV_2_0.IN VCTRL2 0.338f
C14 VDD VCO_C_0.INV_2_5.IN 12.4f
C15 VDD VCO_C_0.INV_2_0.OUT 0.893f
C16 VCO_C_0.INV_2_5.OUT VCO_C_0.INV_2_0.IN 3.46e-19
C17 VCO_C_0.INV_2_2.IN VCO_C_0.INV_2_1.IN 7.5e-19
C18 VCO_C_0.INV_2_5.IN VCTRL2 0.354f
C19 VCO_C_0.INV_2_0.IN VCTRL 1.57f
C20 VCO_C_0.INV_2_0.OUT VCTRL2 0.0273f
C21 VCO_C_0.INV_2_5.OUT VCO_C_0.INV_2_5.IN 0.391f
C22 VCTRL VCO_C_0.INV_2_1.IN 0.0107f
C23 VCO_C_0.INV_2_0.OUT VCO_C_0.INV_2_2.IN 1.2f
C24 DFF_3_mag_0.INV_2_1.IN DFF_3_mag_0.INV_2_5.OUT 1.21f
C25 VCO_C_0.INV_2_5.IN VCTRL 3.24f
C26 DFF_3_mag_0.INV_2_1.IN DFF_3_mag_0.INV_2_5.IN 0.403f
C27 OUT DFF_3_mag_0.INV_2_3.IN 0.577f
C28 VCO_C_0.INV_2_3.IN VCO_C_0.INV_2_1.IN 0.389f
C29 VCO_C_0.INV_2_5.OUT VCO_C_0.INV_2_0.OUT 1.64f
C30 VCO_C_0.INV_2_0.IN VCO_C_0.INV_2_4.IN 0.00756f
C31 VDD VCO_C_0.OUT 0.723f
C32 VCO_C_0.INV_2_0.OUT VCTRL 0.02f
C33 VDD DFF_3_mag_0.INV_2_3.IN 2.59f
C34 VCO_C_0.INV_2_4.IN VCO_C_0.INV_2_1.IN 0.0108f
C35 VCO_C_0.INV_2_0.OUT VCO_C_0.INV_2_3.IN 0.809f
C36 VCTRL2 VCO_C_0.OUT 0.0145f
C37 VCO_C_0.INV_2_5.IN VCO_C_0.INV_2_4.IN 0.00342f
C38 VCO_C_0.INV_2_2.IN VCO_C_0.OUT 9.22e-19
C39 OUT DFF_3_mag_0.INV_2_5.IN 0.0191f
C40 VDD DFF_3_mag_0.INV_2_5.OUT 0.958f
C41 VCTRL VCO_C_0.OUT 0.0471f
C42 VDD DFF_3_mag_0.INV_2_5.IN 2.87f
C43 DFF_3_mag_0.INV_2_0.OUT DFF_3_mag_0.INV_2_3.IN 0.39f
C44 VDD m1_9610_3407# 0.0434f
C45 VCO_C_0.INV_2_0.IN VCO_C_0.OUTB 0.915f
C46 VDD m1_5752_3074# 0.0163f
C47 VCO_C_0.INV_2_4.IN VCO_C_0.OUT 0.385f
C48 VCO_C_0.OUTB VCO_C_0.INV_2_1.IN 0.419f
C49 DFF_3_mag_0.INV_2_0.OUT DFF_3_mag_0.INV_2_5.OUT 0.00977f
C50 VCO_C_0.INV_2_5.IN VCO_C_0.OUTB 0.618f
C51 OUTB DFF_3_mag_0.INV_2_3.IN 0.0234f
C52 DFF_3_mag_0.INV_2_0.OUT DFF_3_mag_0.INV_2_5.IN 0.306f
C53 VCO_C_0.INV_2_2.IN m1_9610_3407# 0.106f
C54 VDD DFF_3_mag_0.INV_2_1.IN 2.74f
C55 VCTRL m1_9610_3407# 5.46e-20
C56 VCTRL m1_5752_3074# 0.0168f
C57 VCO_C_0.INV_2_3.IN m1_9610_3407# 0.00112f
C58 OUTB DFF_3_mag_0.INV_2_5.IN 0.00852f
C59 VCO_C_0.OUT VCO_C_0.OUTB 1.64f
C60 VDD OUT 4.42f
C61 DFF_3_mag_0.INV_2_0.OUT DFF_3_mag_0.INV_2_1.IN 0.546f
C62 VCO_C_0.OUTB DFF_3_mag_0.INV_2_3.IN 0.403f
C63 DFF_3_mag_0.INV_2_3.IN DFF_3_mag_0.INV_2_4.OUT 1.27f
C64 VDD VCTRL2 1.01f
C65 OUTB DFF_3_mag_0.INV_2_1.IN 1.27f
C66 DFF_3_mag_0.INV_2_0.OUT OUT 0.00102f
C67 VDD VCO_C_0.INV_2_2.IN 14.9f
C68 VCO_C_0.OUTB DFF_3_mag_0.INV_2_5.OUT 0.765f
C69 VCO_C_0.OUTB DFF_3_mag_0.INV_2_5.IN 0.652f
C70 DFF_3_mag_0.INV_2_5.IN DFF_3_mag_0.INV_2_4.OUT 7.97e-19
C71 VDD VCO_C_0.INV_2_5.OUT 0.795f
C72 VCO_C_0.INV_2_0.IN VCO_C_0.INV_2_1.IN 3.61e-20
C73 VDD DFF_3_mag_0.INV_2_0.OUT 3.8f
C74 VCO_C_0.INV_2_2.IN VCTRL2 0.108f
C75 VCO_C_0.INV_2_5.IN VCO_C_0.INV_2_0.IN 10.4f
C76 VDD VCTRL 9.76f
C77 VCO_C_0.INV_2_5.OUT VCTRL2 0.198f
C78 VDD VCO_C_0.INV_2_3.IN 12.6f
C79 VCO_C_0.INV_2_5.IN VCO_C_0.INV_2_1.IN 0.00409f
C80 VCO_C_0.INV_2_0.OUT VCO_C_0.INV_2_0.IN 0.388f
C81 OUTB OUT 0.5f
C82 VCO_C_0.INV_2_5.OUT VCO_C_0.INV_2_2.IN 0.915f
C83 VCTRL2 VCTRL 0.0235f
C84 VCO_C_0.INV_2_2.IN VCTRL 1.63f
C85 VDD VCO_C_0.INV_2_4.IN 2.16f
C86 VDD OUTB 0.781f
C87 VCO_C_0.INV_2_3.IN VCTRL2 0.0917f
C88 VCO_C_0.INV_2_0.OUT VCO_C_0.INV_2_5.IN 3.46e-19
C89 VCO_C_0.INV_2_5.OUT VCTRL 0.00912f
C90 VCO_C_0.INV_2_3.IN VCO_C_0.INV_2_2.IN 10.3f
C91 VCO_C_0.OUTB DFF_3_mag_0.INV_2_1.IN 0.624f
C92 VCO_C_0.INV_2_5.OUT VCO_C_0.INV_2_3.IN 0.674f
C93 VCO_C_0.INV_2_0.IN VCO_C_0.OUT 1.19f
C94 VCO_C_0.INV_2_2.IN VCO_C_0.INV_2_4.IN 0.4f
C95 VCO_C_0.INV_2_3.IN VCTRL 3.19f
C96 VCO_C_0.OUT VCO_C_0.INV_2_1.IN 5.91e-19
C97 DFF_3_mag_0.INV_2_0.OUT OUTB 0.493f
C98 VCTRL VCO_C_0.INV_2_4.IN 0.13f
C99 VCO_C_0.INV_2_5.IN VCO_C_0.OUT 0.791f
C100 VCO_C_0.OUTB OUT 0.00703f
C101 OUT DFF_3_mag_0.INV_2_4.OUT 0.382f
C102 VCO_C_0.INV_2_3.IN VCO_C_0.INV_2_4.IN 2.23e-19
C103 VDD VCO_C_0.OUTB 5.93f
C104 VDD DFF_3_mag_0.INV_2_4.OUT 0.921f
C105 VCTRL2 VCO_C_0.OUTB 0.00407f
C106 m1_9610_3407# VSS 0.196f $ **FLOATING
C107 m1_5752_3074# VSS 0.199f $ **FLOATING
C108 DFF_3_mag_0.INV_2_4.OUT VSS 1.68f
C109 DFF_3_mag_0.INV_2_5.OUT VSS 3.77f
C110 DFF_3_mag_0.INV_2_5.IN VSS 3.79f
C111 DFF_3_mag_0.INV_2_3.IN VSS 3.33f
C112 OUT VSS 6.2f
C113 DFF_3_mag_0.INV_2_1.IN VSS 4.03f
C114 OUTB VSS 6.02f
C115 DFF_3_mag_0.INV_2_0.OUT VSS 6.35f
C116 VCO_C_0.INV_2_1.IN VSS 1.97f
C117 VCO_C_0.OUTB VSS 20.9f
C118 VCO_C_0.OUT VSS 5f
C119 VCO_C_0.INV_2_4.IN VSS 1.95f
C120 VCTRL VSS 7.26f
C121 VCTRL2 VSS 45f
C122 VCO_C_0.INV_2_0.IN VSS 6.8f
C123 VCO_C_0.INV_2_5.IN VSS 9.1f
C124 VCO_C_0.INV_2_2.IN VSS 7.23f
C125 VCO_C_0.INV_2_3.IN VSS 8.85f
C126 VCO_C_0.INV_2_0.OUT VSS 5.46f
C127 VCO_C_0.INV_2_5.OUT VSS 6.52f
C128 VDD VSS 0.135p
C129 DFF_3_mag_0.INV_2_0.OUT.t9 VSS 0.00847f
C130 DFF_3_mag_0.INV_2_0.OUT.n0 VSS 0.00847f
C131 DFF_3_mag_0.INV_2_0.OUT.n1 VSS 0.019f
C132 DFF_3_mag_0.INV_2_0.OUT.t8 VSS 0.00847f
C133 DFF_3_mag_0.INV_2_0.OUT.n2 VSS 0.00847f
C134 DFF_3_mag_0.INV_2_0.OUT.n3 VSS 0.019f
C135 DFF_3_mag_0.INV_2_0.OUT.t1 VSS 0.00847f
C136 DFF_3_mag_0.INV_2_0.OUT.n4 VSS 0.00847f
C137 DFF_3_mag_0.INV_2_0.OUT.n5 VSS 0.0169f
C138 DFF_3_mag_0.INV_2_0.OUT.t5 VSS 0.00847f
C139 DFF_3_mag_0.INV_2_0.OUT.n6 VSS 0.00847f
C140 DFF_3_mag_0.INV_2_0.OUT.n7 VSS 0.0207f
C141 DFF_3_mag_0.INV_2_0.OUT.n8 VSS 0.0459f
C142 DFF_3_mag_0.INV_2_0.OUT.n9 VSS 0.0733f
C143 DFF_3_mag_0.INV_2_0.OUT.t3 VSS 0.00847f
C144 DFF_3_mag_0.INV_2_0.OUT.n10 VSS 0.00847f
C145 DFF_3_mag_0.INV_2_0.OUT.n11 VSS 0.0169f
C146 DFF_3_mag_0.INV_2_0.OUT.t7 VSS 0.00847f
C147 DFF_3_mag_0.INV_2_0.OUT.n12 VSS 0.00847f
C148 DFF_3_mag_0.INV_2_0.OUT.n13 VSS 0.0207f
C149 DFF_3_mag_0.INV_2_0.OUT.n14 VSS 0.0459f
C150 DFF_3_mag_0.INV_2_0.OUT.n15 VSS 0.0914f
C151 DFF_3_mag_0.INV_2_0.OUT.t18 VSS 0.0267f
C152 DFF_3_mag_0.INV_2_0.OUT.t16 VSS 0.0684f
C153 DFF_3_mag_0.INV_2_0.OUT.n16 VSS 0.124f
C154 DFF_3_mag_0.INV_2_0.OUT.t25 VSS 0.0267f
C155 DFF_3_mag_0.INV_2_0.OUT.t31 VSS 0.0267f
C156 DFF_3_mag_0.INV_2_0.OUT.t19 VSS 0.0665f
C157 DFF_3_mag_0.INV_2_0.OUT.n17 VSS 0.0765f
C158 DFF_3_mag_0.INV_2_0.OUT.n18 VSS 0.0765f
C159 DFF_3_mag_0.INV_2_0.OUT.t14 VSS 0.11f
C160 DFF_3_mag_0.INV_2_0.OUT.t23 VSS 0.0267f
C161 DFF_3_mag_0.INV_2_0.OUT.t20 VSS 0.0267f
C162 DFF_3_mag_0.INV_2_0.OUT.t15 VSS 0.0665f
C163 DFF_3_mag_0.INV_2_0.OUT.n19 VSS 0.0765f
C164 DFF_3_mag_0.INV_2_0.OUT.n20 VSS 0.0765f
C165 DFF_3_mag_0.INV_2_0.OUT.t13 VSS 0.0967f
C166 DFF_3_mag_0.INV_2_0.OUT.t17 VSS 0.0267f
C167 DFF_3_mag_0.INV_2_0.OUT.t28 VSS 0.0684f
C168 DFF_3_mag_0.INV_2_0.OUT.n21 VSS 0.0796f
C169 DFF_3_mag_0.INV_2_0.OUT.t24 VSS 0.0267f
C170 DFF_3_mag_0.INV_2_0.OUT.t29 VSS 0.0267f
C171 DFF_3_mag_0.INV_2_0.OUT.t21 VSS 0.0625f
C172 DFF_3_mag_0.INV_2_0.OUT.t26 VSS 0.119f
C173 DFF_3_mag_0.INV_2_0.OUT.n22 VSS 0.0883f
C174 DFF_3_mag_0.INV_2_0.OUT.n23 VSS 0.0645f
C175 DFF_3_mag_0.INV_2_0.OUT.n24 VSS 0.215f
C176 DFF_3_mag_0.INV_2_0.OUT.n25 VSS 0.422f
C177 DFF_3_mag_0.INV_2_0.OUT.t30 VSS 0.0267f
C178 DFF_3_mag_0.INV_2_0.OUT.t27 VSS 0.0267f
C179 DFF_3_mag_0.INV_2_0.OUT.t12 VSS 0.0625f
C180 DFF_3_mag_0.INV_2_0.OUT.t22 VSS 0.119f
C181 DFF_3_mag_0.INV_2_0.OUT.n26 VSS 0.0883f
C182 DFF_3_mag_0.INV_2_0.OUT.n27 VSS 0.0605f
C183 DFF_3_mag_0.INV_2_0.OUT.n28 VSS 0.113f
C184 DFF_3_mag_0.INV_2_3.IN.n0 VSS 0.182f
C185 DFF_3_mag_0.INV_2_3.IN.n1 VSS 0.182f
C186 DFF_3_mag_0.INV_2_3.IN.t21 VSS 0.0291f
C187 DFF_3_mag_0.INV_2_3.IN.t20 VSS 0.0138f
C188 DFF_3_mag_0.INV_2_3.IN.n2 VSS 0.0449f
C189 DFF_3_mag_0.INV_2_3.IN.n3 VSS 0.032f
C190 DFF_3_mag_0.INV_2_3.IN.t18 VSS 0.0338f
C191 DFF_3_mag_0.INV_2_3.IN.n4 VSS 0.0388f
C192 DFF_3_mag_0.INV_2_3.IN.t26 VSS 0.0138f
C193 DFF_3_mag_0.INV_2_3.IN.n5 VSS 0.0396f
C194 DFF_3_mag_0.INV_2_3.IN.t22 VSS 0.0338f
C195 DFF_3_mag_0.INV_2_3.IN.n6 VSS 0.032f
C196 DFF_3_mag_0.INV_2_3.IN.t17 VSS 0.0445f
C197 DFF_3_mag_0.INV_2_3.IN.t24 VSS 0.0183f
C198 DFF_3_mag_0.INV_2_3.IN.n7 VSS 0.0489f
C199 DFF_3_mag_0.INV_2_3.IN.t16 VSS 0.0445f
C200 DFF_3_mag_0.INV_2_3.IN.n8 VSS 0.0489f
C201 DFF_3_mag_0.INV_2_3.IN.t19 VSS 0.0183f
C202 DFF_3_mag_0.INV_2_3.IN.n9 VSS 0.0388f
C203 DFF_3_mag_0.INV_2_3.IN.t25 VSS 0.0338f
C204 DFF_3_mag_0.INV_2_3.IN.t27 VSS 0.0138f
C205 DFF_3_mag_0.INV_2_3.IN.n10 VSS 0.0449f
C206 DFF_3_mag_0.INV_2_3.IN.t23 VSS 0.0138f
C207 DFF_3_mag_0.INV_2_3.IN.n11 VSS 0.0227f
C208 DFF_3_mag_0.INV_2_3.IN.n12 VSS 0.0229f
C209 DFF_3_mag_0.INV_2_3.IN.t6 VSS 0.0171f
C210 DFF_3_mag_0.INV_2_3.IN.t4 VSS 0.0681f
C211 DFF_3_mag_0.INV_2_3.IN.n13 VSS 0.0188f
C212 DFF_3_mag_0.INV_2_3.IN.t5 VSS 0.023f
C213 DFF_3_mag_0.INV_2_3.IN.n14 VSS 0.0488f
C214 DFF_3_mag_0.INV_2_3.IN.t11 VSS 0.00929f
C215 DFF_3_mag_0.INV_2_3.IN.n15 VSS 0.00929f
C216 DFF_3_mag_0.INV_2_3.IN.n16 VSS 0.0291f
C217 DFF_3_mag_0.INV_2_3.IN.t9 VSS 0.00929f
C218 DFF_3_mag_0.INV_2_3.IN.n17 VSS 0.00929f
C219 DFF_3_mag_0.INV_2_3.IN.n18 VSS 0.0187f
C220 DFF_3_mag_0.INV_2_3.IN.n19 VSS 0.0943f
C221 DFF_3_mag_0.INV_2_3.IN.n20 VSS 0.165f
C222 DFF_3_mag_0.INV_2_3.IN.n21 VSS 0.181f
C223 DFF_3_mag_0.INV_2_3.IN.t1 VSS 0.0681f
C224 DFF_3_mag_0.INV_2_3.IN.n22 VSS 0.0188f
C225 DFF_3_mag_0.INV_2_3.IN.t0 VSS 0.023f
C226 DFF_3_mag_0.INV_2_3.IN.t3 VSS 0.0171f
C227 DFF_3_mag_0.INV_2_3.IN.n23 VSS 0.0487f
C228 DFF_3_mag_0.INV_2_3.IN.t7 VSS 0.00929f
C229 DFF_3_mag_0.INV_2_3.IN.n24 VSS 0.00929f
C230 DFF_3_mag_0.INV_2_3.IN.n25 VSS 0.0187f
C231 DFF_3_mag_0.INV_2_3.IN.t14 VSS 0.00929f
C232 DFF_3_mag_0.INV_2_3.IN.n26 VSS 0.00929f
C233 DFF_3_mag_0.INV_2_3.IN.n27 VSS 0.0291f
C234 DFF_3_mag_0.INV_2_3.IN.n28 VSS 0.0943f
C235 DFF_3_mag_0.INV_2_3.IN.n29 VSS 0.165f
C236 a_1424_1033.n0 VSS 0.0859f
C237 a_1424_1033.n1 VSS 0.113f
C238 a_1424_1033.n2 VSS 0.089f
C239 a_1424_1033.n3 VSS 0.15f
C240 a_1424_1033.n4 VSS 0.194f
C241 a_1424_1033.n5 VSS 0.173f
C242 a_1424_1033.n6 VSS 0.0692f
C243 a_1424_1033.t22 VSS 0.00968f
C244 a_1424_1033.n7 VSS 0.00968f
C245 a_1424_1033.n8 VSS 0.0244f
C246 a_1424_1033.t30 VSS 0.00968f
C247 a_1424_1033.n9 VSS 0.00968f
C248 a_1424_1033.n10 VSS 0.0194f
C249 a_1424_1033.t38 VSS 0.00968f
C250 a_1424_1033.n11 VSS 0.00968f
C251 a_1424_1033.n12 VSS 0.0243f
C252 a_1424_1033.n13 VSS 0.064f
C253 a_1424_1033.t49 VSS 0.00968f
C254 a_1424_1033.n14 VSS 0.00968f
C255 a_1424_1033.n15 VSS 0.0194f
C256 a_1424_1033.t31 VSS 0.00968f
C257 a_1424_1033.n16 VSS 0.00968f
C258 a_1424_1033.n17 VSS 0.0194f
C259 a_1424_1033.n18 VSS 0.0528f
C260 a_1424_1033.t42 VSS 0.00968f
C261 a_1424_1033.n19 VSS 0.00968f
C262 a_1424_1033.n20 VSS 0.0246f
C263 a_1424_1033.t43 VSS 0.00968f
C264 a_1424_1033.n21 VSS 0.00968f
C265 a_1424_1033.n22 VSS 0.0463f
C266 a_1424_1033.n23 VSS 0.08f
C267 a_1424_1033.n24 VSS 0.136f
C268 a_1424_1033.t23 VSS 0.00968f
C269 a_1424_1033.n25 VSS 0.00968f
C270 a_1424_1033.n26 VSS 0.0194f
C271 a_1424_1033.t45 VSS 0.00968f
C272 a_1424_1033.n27 VSS 0.00968f
C273 a_1424_1033.n28 VSS 0.0194f
C274 a_1424_1033.t21 VSS 0.00968f
C275 a_1424_1033.n29 VSS 0.00968f
C276 a_1424_1033.n30 VSS 0.0194f
C277 a_1424_1033.t51 VSS 0.00968f
C278 a_1424_1033.n31 VSS 0.00968f
C279 a_1424_1033.n32 VSS 0.0194f
C280 a_1424_1033.n33 VSS 0.053f
C281 a_1424_1033.t20 VSS 0.00968f
C282 a_1424_1033.n34 VSS 0.00968f
C283 a_1424_1033.n35 VSS 0.0194f
C284 a_1424_1033.t29 VSS 0.00968f
C285 a_1424_1033.n36 VSS 0.00968f
C286 a_1424_1033.n37 VSS 0.0194f
C287 a_1424_1033.n38 VSS 0.0363f
C288 a_1424_1033.t1 VSS 0.00968f
C289 a_1424_1033.n39 VSS 0.00968f
C290 a_1424_1033.n40 VSS 0.0194f
C291 a_1424_1033.n41 VSS 0.0953f
C292 a_1424_1033.n42 VSS 0.0807f
C293 a_1424_1033.t12 VSS 0.00968f
C294 a_1424_1033.n43 VSS 0.00968f
C295 a_1424_1033.n44 VSS 0.0194f
C296 a_1424_1033.n45 VSS 0.0474f
C297 a_1424_1033.t18 VSS 0.00968f
C298 a_1424_1033.n46 VSS 0.00968f
C299 a_1424_1033.n47 VSS 0.0194f
C300 a_1424_1033.n48 VSS 0.0476f
C301 a_1424_1033.n49 VSS 0.0807f
C302 a_1424_1033.t5 VSS 0.00968f
C303 a_1424_1033.n50 VSS 0.00968f
C304 a_1424_1033.n51 VSS 0.0194f
C305 a_1424_1033.n52 VSS 0.0581f
C306 a_1424_1033.t14 VSS 0.00968f
C307 a_1424_1033.n53 VSS 0.00968f
C308 a_1424_1033.n54 VSS 0.0194f
C309 a_1424_1033.n55 VSS 0.068f
C310 a_1424_1033.t16 VSS 0.00968f
C311 a_1424_1033.n56 VSS 0.00968f
C312 a_1424_1033.n57 VSS 0.0194f
C313 a_1424_1033.n58 VSS 0.0951f
C314 a_1424_1033.n59 VSS 0.0807f
C315 a_1424_1033.t3 VSS 0.00968f
C316 a_1424_1033.n60 VSS 0.00968f
C317 a_1424_1033.n61 VSS 0.0194f
C318 a_1424_1033.n62 VSS 0.0474f
C319 a_1424_1033.t8 VSS 0.00968f
C320 a_1424_1033.n63 VSS 0.00968f
C321 a_1424_1033.n64 VSS 0.0194f
C322 a_1424_1033.n65 VSS 0.0476f
C323 a_1424_1033.n66 VSS 0.0807f
C324 a_1424_1033.t17 VSS 0.00968f
C325 a_1424_1033.n67 VSS 0.00968f
C326 a_1424_1033.n68 VSS 0.0194f
C327 a_1424_1033.n69 VSS 0.0581f
C328 a_1424_1033.t4 VSS 0.00968f
C329 a_1424_1033.n70 VSS 0.00968f
C330 a_1424_1033.n71 VSS 0.0194f
C331 a_1424_1033.n72 VSS 0.064f
C332 a_1424_1033.n73 VSS 0.474f
C333 a_1424_1033.t24 VSS 0.00968f
C334 a_1424_1033.n74 VSS 0.00968f
C335 a_1424_1033.n75 VSS 0.028f
C336 a_1424_1033.n76 VSS 0.129f
C337 a_1424_1033.t35 VSS 0.00968f
C338 a_1424_1033.n77 VSS 0.00968f
C339 a_1424_1033.n78 VSS 0.0194f
C340 a_1424_1033.t41 VSS 0.00968f
C341 a_1424_1033.n79 VSS 0.00968f
C342 a_1424_1033.n80 VSS 0.0194f
C343 a_1424_1033.n81 VSS 0.0376f
C344 a_1424_1033.t48 VSS 0.00968f
C345 a_1424_1033.n82 VSS 0.00968f
C346 a_1424_1033.n83 VSS 0.0194f
C347 a_1424_1033.n84 VSS 0.105f
C348 a_1424_1033.n85 VSS 0.143f
C349 a_1424_1033.n86 VSS 0.451f
C350 a_1424_1033.n87 VSS 0.158f
C351 a_1424_1033.n88 VSS 0.105f
C352 a_1424_1033.t40 VSS 0.00968f
C353 a_1424_1033.n89 VSS 0.00968f
C354 a_1424_1033.n90 VSS 0.0763f
C355 a_1424_1033.n91 VSS 0.463f
C356 a_1424_1033.t54 VSS 0.00968f
C357 a_1424_1033.n92 VSS 0.00968f
C358 a_1424_1033.n93 VSS 0.0194f
C359 a_1424_1033.n94 VSS 0.0538f
C360 a_1424_1033.n95 VSS 0.0592f
C361 a_1424_1033.n96 VSS 0.00968f
C362 a_1424_1033.n97 VSS 0.0244f
C363 a_1424_1033.t58 VSS 0.00968f
C364 OUT.t19 VSS 0.0215f
C365 OUT.n0 VSS 0.0353f
C366 OUT.n1 VSS 0.0605f
C367 OUT.t29 VSS 0.0285f
C368 OUT.t26 VSS 0.0694f
C369 OUT.n2 VSS 0.0498f
C370 OUT.t20 VSS 0.0216f
C371 OUT.t17 VSS 0.0527f
C372 OUT.n3 VSS 0.0617f
C373 OUT.t31 VSS 0.0216f
C374 OUT.t21 VSS 0.0216f
C375 OUT.t18 VSS 0.0527f
C376 OUT.n4 VSS 0.07f
C377 OUT.n5 VSS 0.07f
C378 OUT.t30 VSS 0.0527f
C379 OUT.n6 VSS 0.0605f
C380 OUT.t15 VSS 0.0285f
C381 OUT.n7 VSS 0.0762f
C382 OUT.n8 VSS 0.0762f
C383 OUT.t24 VSS 0.0694f
C384 OUT.n9 VSS 0.0498f
C385 OUT.t12 VSS 0.0454f
C386 OUT.n10 VSS 0.0357f
C387 OUT.n11 VSS 0.639f
C388 OUT.t5 VSS 0.00862f
C389 OUT.n12 VSS 0.00862f
C390 OUT.n13 VSS 0.0211f
C391 OUT.t10 VSS 0.00862f
C392 OUT.n14 VSS 0.00862f
C393 OUT.n15 VSS 0.0172f
C394 OUT.n16 VSS 0.0468f
C395 OUT.t3 VSS 0.00862f
C396 OUT.n17 VSS 0.00862f
C397 OUT.n18 VSS 0.0194f
C398 OUT.t7 VSS 0.00862f
C399 OUT.n19 VSS 0.00862f
C400 OUT.n20 VSS 0.0211f
C401 OUT.t2 VSS 0.00862f
C402 OUT.n21 VSS 0.00862f
C403 OUT.n22 VSS 0.0172f
C404 OUT.n23 VSS 0.0468f
C405 OUT.t4 VSS 0.00862f
C406 OUT.n24 VSS 0.00862f
C407 OUT.n25 VSS 0.0194f
C408 OUT.n26 VSS 0.0747f
C409 OUT.n27 VSS 0.0931f
C410 OUT.t33 VSS 0.0215f
C411 OUT.n28 VSS 0.0353f
C412 OUT.n29 VSS 0.0605f
C413 OUT.t27 VSS 0.0285f
C414 OUT.t35 VSS 0.0694f
C415 OUT.n30 VSS 0.0498f
C416 OUT.t32 VSS 0.0216f
C417 OUT.t23 VSS 0.0527f
C418 OUT.n31 VSS 0.0617f
C419 OUT.t34 VSS 0.0216f
C420 OUT.t22 VSS 0.0216f
C421 OUT.t14 VSS 0.0527f
C422 OUT.n32 VSS 0.07f
C423 OUT.n33 VSS 0.07f
C424 OUT.t28 VSS 0.0527f
C425 OUT.n34 VSS 0.0605f
C426 OUT.t16 VSS 0.0285f
C427 OUT.n35 VSS 0.0762f
C428 OUT.n36 VSS 0.0762f
C429 OUT.t13 VSS 0.0694f
C430 OUT.n37 VSS 0.0498f
C431 OUT.t25 VSS 0.0454f
C432 OUT.n38 VSS 0.0357f
C433 OUT.n39 VSS 0.279f
C434 OUT.n40 VSS 0.0601f
C435 DFF_3_mag_0.INV_2_5.IN.t17 VSS 0.0143f
C436 DFF_3_mag_0.INV_2_5.IN.n0 VSS 0.0143f
C437 DFF_3_mag_0.INV_2_5.IN.n1 VSS 0.0304f
C438 DFF_3_mag_0.INV_2_5.IN.n2 VSS 0.0353f
C439 DFF_3_mag_0.INV_2_5.IN.n3 VSS 0.0352f
C440 DFF_3_mag_0.INV_2_5.IN.n4 VSS 0.0353f
C441 DFF_3_mag_0.INV_2_5.IN.t3 VSS 0.0143f
C442 DFF_3_mag_0.INV_2_5.IN.n5 VSS 0.0143f
C443 DFF_3_mag_0.INV_2_5.IN.n6 VSS 0.0537f
C444 DFF_3_mag_0.INV_2_5.IN.n7 VSS 0.145f
C445 DFF_3_mag_0.INV_2_5.IN.n8 VSS 0.0233f
C446 DFF_3_mag_0.INV_2_5.IN.n9 VSS 0.0407f
C447 DFF_3_mag_0.INV_2_5.IN.n10 VSS 0.099f
C448 DFF_3_mag_0.INV_2_5.IN.n11 VSS 0.0943f
C449 DFF_3_mag_0.INV_2_5.IN.t19 VSS 0.0266f
C450 DFF_3_mag_0.INV_2_5.IN.n12 VSS 0.191f
C451 DFF_3_mag_0.INV_2_5.IN.t25 VSS 0.0212f
C452 DFF_3_mag_0.INV_2_5.IN.n13 VSS 0.0347f
C453 DFF_3_mag_0.INV_2_5.IN.n14 VSS 0.0595f
C454 DFF_3_mag_0.INV_2_5.IN.t30 VSS 0.0281f
C455 DFF_3_mag_0.INV_2_5.IN.t27 VSS 0.0682f
C456 DFF_3_mag_0.INV_2_5.IN.n15 VSS 0.049f
C457 DFF_3_mag_0.INV_2_5.IN.t28 VSS 0.0212f
C458 DFF_3_mag_0.INV_2_5.IN.t26 VSS 0.0519f
C459 DFF_3_mag_0.INV_2_5.IN.n16 VSS 0.0607f
C460 DFF_3_mag_0.INV_2_5.IN.t23 VSS 0.0212f
C461 DFF_3_mag_0.INV_2_5.IN.t21 VSS 0.0212f
C462 DFF_3_mag_0.INV_2_5.IN.t31 VSS 0.0519f
C463 DFF_3_mag_0.INV_2_5.IN.n17 VSS 0.0688f
C464 DFF_3_mag_0.INV_2_5.IN.n18 VSS 0.0688f
C465 DFF_3_mag_0.INV_2_5.IN.t22 VSS 0.0519f
C466 DFF_3_mag_0.INV_2_5.IN.n19 VSS 0.0595f
C467 DFF_3_mag_0.INV_2_5.IN.t29 VSS 0.0281f
C468 DFF_3_mag_0.INV_2_5.IN.n20 VSS 0.075f
C469 DFF_3_mag_0.INV_2_5.IN.n21 VSS 0.075f
C470 DFF_3_mag_0.INV_2_5.IN.t20 VSS 0.0682f
C471 DFF_3_mag_0.INV_2_5.IN.n22 VSS 0.049f
C472 DFF_3_mag_0.INV_2_5.IN.t24 VSS 0.0447f
C473 DFF_3_mag_0.INV_2_5.IN.n23 VSS 0.0351f
C474 DFF_3_mag_0.INV_2_5.IN.n24 VSS 0.27f
C475 DFF_3_mag_0.INV_2_5.IN.t15 VSS 0.00848f
C476 DFF_3_mag_0.INV_2_5.IN.n25 VSS 0.00848f
C477 DFF_3_mag_0.INV_2_5.IN.n26 VSS 0.0191f
C478 DFF_3_mag_0.INV_2_5.IN.t5 VSS 0.00848f
C479 DFF_3_mag_0.INV_2_5.IN.n27 VSS 0.00848f
C480 DFF_3_mag_0.INV_2_5.IN.n28 VSS 0.0207f
C481 DFF_3_mag_0.INV_2_5.IN.t10 VSS 0.00848f
C482 DFF_3_mag_0.INV_2_5.IN.n29 VSS 0.00848f
C483 DFF_3_mag_0.INV_2_5.IN.n30 VSS 0.017f
C484 DFF_3_mag_0.INV_2_5.IN.n31 VSS 0.046f
C485 DFF_3_mag_0.INV_2_5.IN.t16 VSS 0.00848f
C486 DFF_3_mag_0.INV_2_5.IN.n32 VSS 0.00848f
C487 DFF_3_mag_0.INV_2_5.IN.n33 VSS 0.0191f
C488 DFF_3_mag_0.INV_2_5.IN.n34 VSS 0.0735f
C489 DFF_3_mag_0.INV_2_5.IN.t11 VSS 0.00848f
C490 DFF_3_mag_0.INV_2_5.IN.n35 VSS 0.00848f
C491 DFF_3_mag_0.INV_2_5.IN.n36 VSS 0.0207f
C492 DFF_3_mag_0.INV_2_5.IN.t8 VSS 0.00848f
C493 DFF_3_mag_0.INV_2_5.IN.n37 VSS 0.00848f
C494 DFF_3_mag_0.INV_2_5.IN.n38 VSS 0.017f
C495 DFF_3_mag_0.INV_2_5.IN.n39 VSS 0.046f
C496 DFF_3_mag_0.INV_2_5.IN.n40 VSS 0.0916f
C497 VCO_C_0.INV_2_0.IN.n0 VSS 0.631f
C498 VCO_C_0.INV_2_0.IN.n1 VSS 0.366f
C499 VCO_C_0.INV_2_0.IN.n2 VSS 0.501f
C500 VCO_C_0.INV_2_0.IN.n3 VSS 0.622f
C501 VCO_C_0.INV_2_0.IN.n4 VSS 0.586f
C502 VCO_C_0.INV_2_0.IN.n5 VSS 0.501f
C503 VCO_C_0.INV_2_0.IN.n6 VSS 0.118f
C504 VCO_C_0.INV_2_0.IN.n7 VSS 0.457f
C505 VCO_C_0.INV_2_0.IN.t47 VSS 0.0406f
C506 VCO_C_0.INV_2_0.IN.n8 VSS 0.116f
C507 VCO_C_0.INV_2_0.IN.t34 VSS 0.0406f
C508 VCO_C_0.INV_2_0.IN.t37 VSS 0.0992f
C509 VCO_C_0.INV_2_0.IN.n9 VSS 0.132f
C510 VCO_C_0.INV_2_0.IN.t41 VSS 0.0406f
C511 VCO_C_0.INV_2_0.IN.t46 VSS 0.0992f
C512 VCO_C_0.INV_2_0.IN.n10 VSS 0.132f
C513 VCO_C_0.INV_2_0.IN.t56 VSS 0.0405f
C514 VCO_C_0.INV_2_0.IN.n11 VSS 0.0664f
C515 VCO_C_0.INV_2_0.IN.t52 VSS 0.0992f
C516 VCO_C_0.INV_2_0.IN.t57 VSS 0.13f
C517 VCO_C_0.INV_2_0.IN.n12 VSS 0.0937f
C518 VCO_C_0.INV_2_0.IN.n13 VSS 0.143f
C519 VCO_C_0.INV_2_0.IN.t42 VSS 0.0537f
C520 VCO_C_0.INV_2_0.IN.n14 VSS 0.114f
C521 VCO_C_0.INV_2_0.IN.n15 VSS 0.143f
C522 VCO_C_0.INV_2_0.IN.t49 VSS 0.0537f
C523 VCO_C_0.INV_2_0.IN.n16 VSS 0.114f
C524 VCO_C_0.INV_2_0.IN.t35 VSS 0.13f
C525 VCO_C_0.INV_2_0.IN.n17 VSS 0.0937f
C526 VCO_C_0.INV_2_0.IN.t31 VSS 0.0855f
C527 VCO_C_0.INV_2_0.IN.n18 VSS 0.0672f
C528 VCO_C_0.INV_2_0.IN.n19 VSS 0.0176f
C529 VCO_C_0.INV_2_0.IN.t3 VSS 0.0149f
C530 VCO_C_0.INV_2_0.IN.n20 VSS 0.105f
C531 VCO_C_0.INV_2_0.IN.t1 VSS 0.0577f
C532 VCO_C_0.INV_2_0.IN.n21 VSS 0.525f
C533 VCO_C_0.INV_2_0.IN.n22 VSS 0.0926f
C534 VCO_C_0.INV_2_0.IN.n23 VSS 0.0176f
C535 VCO_C_0.INV_2_0.IN.t4 VSS 0.0149f
C536 VCO_C_0.INV_2_0.IN.n24 VSS 0.0586f
C537 VCO_C_0.INV_2_0.IN.t0 VSS 0.103f
C538 VCO_C_0.INV_2_0.IN.n25 VSS 0.0176f
C539 VCO_C_0.INV_2_0.IN.t2 VSS 0.0149f
C540 VCO_C_0.INV_2_0.IN.n26 VSS 0.0326f
C541 VCO_C_0.INV_2_0.IN.n27 VSS 0.0547f
C542 VCO_C_0.INV_2_0.IN.n28 VSS 0.0537f
C543 VCO_C_0.INV_2_0.IN.n29 VSS 0.453f
C544 VCO_C_0.INV_2_0.IN.n30 VSS 0.315f
C545 VCO_C_0.INV_2_0.IN.t10 VSS 0.093f
C546 VCO_C_0.INV_2_0.IN.t14 VSS 0.0385f
C547 VCO_C_0.INV_2_0.IN.n31 VSS 0.507f
C548 VCO_C_0.INV_2_0.IN.t13 VSS 0.0162f
C549 VCO_C_0.INV_2_0.IN.n32 VSS 0.0162f
C550 VCO_C_0.INV_2_0.IN.n33 VSS 0.0802f
C551 VCO_C_0.INV_2_0.IN.n34 VSS 0.349f
C552 VCO_C_0.INV_2_0.IN.n35 VSS 0.0345f
C553 VCO_C_0.INV_2_0.IN.n36 VSS 0.372f
C554 VCO_C_0.INV_2_0.IN.t21 VSS 0.0162f
C555 VCO_C_0.INV_2_0.IN.n37 VSS 0.0162f
C556 VCO_C_0.INV_2_0.IN.n38 VSS 0.0325f
C557 VCO_C_0.INV_2_0.IN.n39 VSS 0.0337f
C558 VCO_C_0.INV_2_0.IN.n40 VSS 0.0484f
C559 VCO_C_0.INV_2_0.IN.n41 VSS 0.0283f
C560 VCO_C_0.INV_2_0.IN.n42 VSS 0.0842f
C561 VCO_C_0.INV_2_0.IN.t26 VSS 0.0262f
C562 VCO_C_0.INV_2_0.IN.n43 VSS 0.0399f
C563 VCO_C_0.INV_2_0.IN.n44 VSS 0.29f
C564 VCO_C_0.INV_2_0.IN.t15 VSS 0.0254f
C565 VCO_C_0.INV_2_0.IN.n45 VSS 0.473f
C566 VCO_C_0.INV_2_0.IN.n46 VSS 0.249f
C567 VCO_C_0.INV_2_0.IN.t30 VSS 0.0666f
C568 VCO_C_0.INV_2_0.IN.n47 VSS 0.326f
C569 VCO_C_0.INV_2_0.IN.n48 VSS 0.3f
C570 VCO_C_0.INV_2_0.IN.t39 VSS 0.11f
C571 VCO_C_0.INV_2_0.IN.t54 VSS 0.113f
C572 VCO_C_0.INV_2_0.IN.t40 VSS 0.11f
C573 VCO_C_0.INV_2_0.IN.t55 VSS 0.113f
C574 VCO_C_0.INV_2_0.IN.t43 VSS 0.114f
C575 VCO_C_0.INV_2_0.IN.t32 VSS 0.11f
C576 VCO_C_0.INV_2_0.IN.t48 VSS 0.111f
C577 VCO_C_0.INV_2_0.IN.t36 VSS 0.11f
C578 VCO_C_0.INV_2_0.IN.t33 VSS 0.115f
C579 VCO_C_0.INV_2_0.IN.t51 VSS 0.115f
C580 VCO_C_0.INV_2_0.IN.t58 VSS 0.112f
C581 VCO_C_0.INV_2_0.IN.t45 VSS 0.15f
C582 VCO_C_0.INV_2_0.IN.n49 VSS 0.842f
C583 VCO_C_0.INV_2_0.IN.n50 VSS 0.387f
C584 VCO_C_0.INV_2_0.IN.n51 VSS 0.511f
C585 VCO_C_0.INV_2_0.IN.t53 VSS 0.11f
C586 VCO_C_0.INV_2_0.IN.t44 VSS 0.11f
C587 VCO_C_0.INV_2_0.IN.t50 VSS 0.111f
C588 VCO_C_0.INV_2_0.IN.t38 VSS 0.151f
C589 VCO_C_0.INV_2_0.IN.n52 VSS 0.82f
C590 VCO_C_0.INV_2_0.IN.n53 VSS 0.371f
C591 VCO_C_0.INV_2_0.IN.n54 VSS 0.496f
C592 VCO_C_0.INV_2_0.IN.n55 VSS 0.676f
C593 VCO_C_0.INV_2_0.IN.n56 VSS 0.0239f
C594 VCO_C_0.INV_2_0.IN.n57 VSS 0.0239f
C595 VCO_C_0.INV_2_0.IN.t17 VSS 0.0162f
C596 VCO_C_0.INV_2_0.IN.n58 VSS 0.0162f
C597 VCO_C_0.INV_2_0.IN.n59 VSS 0.0757f
C598 VCO_C_0.INV_2_0.IN.t24 VSS 0.0262f
C599 VCO_C_0.INV_2_0.IN.n60 VSS 0.0654f
C600 VCO_C_0.INV_2_0.IN.n61 VSS 0.0505f
C601 VCO_C_0.INV_2_0.IN.n62 VSS 0.0645f
C602 VCO_C_0.INV_2_0.IN.t25 VSS 0.0162f
C603 VCO_C_0.INV_2_0.IN.n63 VSS 0.0162f
C604 VCO_C_0.INV_2_0.IN.n64 VSS 0.0325f
C605 VCO_C_0.INV_2_0.IN.n65 VSS 0.177f
C606 VCO_C_0.INV_2_0.IN.n66 VSS 0.7f
C607 VCO_C_0.INV_2_0.IN.n67 VSS 0.24f
C608 VCO_C_0.INV_2_0.IN.n68 VSS 0.456f
C609 VCO_C_0.INV_2_0.IN.n69 VSS 0.112f
C610 VCO_C_0.INV_2_0.IN.n70 VSS 0.118f
C611 VCO_C_0.INV_2_0.IN.n71 VSS 0.177f
C612 VCO_C_0.INV_2_0.IN.n72 VSS 0.473f
C613 VCO_C_0.INV_2_0.IN.n73 VSS 2.22f
C614 VCO_C_0.INV_2_0.IN.n74 VSS 0.931f
C615 VCO_C_0.INV_2_0.IN.n75 VSS 0.66f
C616 VCO_C_0.INV_2_0.IN.n76 VSS 0.0631f
C617 VCO_C_0.INV_2_0.IN.n77 VSS 0.0326f
C618 VCO_C_0.INV_2_0.IN.n78 VSS 0.0162f
C619 VCO_C_0.INV_2_0.IN.t18 VSS 0.0162f
C620 VCO_C_0.INV_2_4.IN.t10 VSS 0.011f
C621 VCO_C_0.INV_2_4.IN.n0 VSS 0.011f
C622 VCO_C_0.INV_2_4.IN.n1 VSS 0.0248f
C623 VCO_C_0.INV_2_4.IN.t1 VSS 0.011f
C624 VCO_C_0.INV_2_4.IN.n2 VSS 0.011f
C625 VCO_C_0.INV_2_4.IN.n3 VSS 0.027f
C626 VCO_C_0.INV_2_4.IN.t6 VSS 0.011f
C627 VCO_C_0.INV_2_4.IN.n4 VSS 0.011f
C628 VCO_C_0.INV_2_4.IN.n5 VSS 0.0221f
C629 VCO_C_0.INV_2_4.IN.n6 VSS 0.0599f
C630 VCO_C_0.INV_2_4.IN.t11 VSS 0.011f
C631 VCO_C_0.INV_2_4.IN.n7 VSS 0.011f
C632 VCO_C_0.INV_2_4.IN.n8 VSS 0.0248f
C633 VCO_C_0.INV_2_4.IN.n9 VSS 0.0956f
C634 VCO_C_0.INV_2_4.IN.t0 VSS 0.011f
C635 VCO_C_0.INV_2_4.IN.n10 VSS 0.011f
C636 VCO_C_0.INV_2_4.IN.n11 VSS 0.027f
C637 VCO_C_0.INV_2_4.IN.t5 VSS 0.011f
C638 VCO_C_0.INV_2_4.IN.n12 VSS 0.011f
C639 VCO_C_0.INV_2_4.IN.n13 VSS 0.0221f
C640 VCO_C_0.INV_2_4.IN.n14 VSS 0.0599f
C641 VCO_C_0.INV_2_4.IN.n15 VSS 0.119f
C642 VCO_C_0.INV_2_4.IN.t17 VSS 0.0582f
C643 VCO_C_0.INV_2_4.IN.t16 VSS 0.0276f
C644 VCO_C_0.INV_2_4.IN.n16 VSS 0.0896f
C645 VCO_C_0.INV_2_4.IN.n17 VSS 0.0638f
C646 VCO_C_0.INV_2_4.IN.t13 VSS 0.0675f
C647 VCO_C_0.INV_2_4.IN.n18 VSS 0.0775f
C648 VCO_C_0.INV_2_4.IN.t14 VSS 0.0888f
C649 VCO_C_0.INV_2_4.IN.t21 VSS 0.0276f
C650 VCO_C_0.INV_2_4.IN.n19 VSS 0.079f
C651 VCO_C_0.INV_2_4.IN.t18 VSS 0.0675f
C652 VCO_C_0.INV_2_4.IN.n20 VSS 0.0638f
C653 VCO_C_0.INV_2_4.IN.t15 VSS 0.0888f
C654 VCO_C_0.INV_2_4.IN.t12 VSS 0.0365f
C655 VCO_C_0.INV_2_4.IN.n21 VSS 0.0976f
C656 VCO_C_0.INV_2_4.IN.n22 VSS 0.0976f
C657 VCO_C_0.INV_2_4.IN.t19 VSS 0.0365f
C658 VCO_C_0.INV_2_4.IN.n23 VSS 0.0775f
C659 VCO_C_0.INV_2_4.IN.t22 VSS 0.0675f
C660 VCO_C_0.INV_2_4.IN.t23 VSS 0.0276f
C661 VCO_C_0.INV_2_4.IN.n24 VSS 0.0896f
C662 VCO_C_0.INV_2_4.IN.t20 VSS 0.0276f
C663 VCO_C_0.INV_2_4.IN.n25 VSS 0.0452f
C664 VCO_C_0.INV_2_4.IN.n26 VSS 0.0457f
C665 VCTRL2.n0 VSS 0.0391f
C666 VCTRL2.n1 VSS 0.015f
C667 VCTRL2.n2 VSS 0.0646f
C668 VCTRL2.t28 VSS 0.023f
C669 VCTRL2.n3 VSS 0.0337f
C670 VCTRL2.n4 VSS 0.0336f
C671 VCTRL2.n5 VSS 0.0336f
C672 VCTRL2.t18 VSS 0.0232f
C673 VCTRL2.n6 VSS 0.0449f
C674 VCTRL2.t32 VSS 0.0427f
C675 VCTRL2.n7 VSS 0.0336f
C676 VCTRL2.n8 VSS 0.0449f
C677 VCTRL2.t54 VSS 0.045f
C678 VCTRL2.n9 VSS 0.0449f
C679 VCTRL2.t16 VSS 0.0395f
C680 VCTRL2.n10 VSS 0.0438f
C681 VCTRL2.t50 VSS 0.023f
C682 VCTRL2.n11 VSS 0.0337f
C683 VCTRL2.t38 VSS 0.0232f
C684 VCTRL2.n12 VSS 0.0449f
C685 VCTRL2.t53 VSS 0.0427f
C686 VCTRL2.n13 VSS 0.0335f
C687 VCTRL2.n14 VSS 0.0339f
C688 VCTRL2.n15 VSS 0.0337f
C689 VCTRL2.n16 VSS 0.0449f
C690 VCTRL2.t72 VSS 0.045f
C691 VCTRL2.n17 VSS 0.0449f
C692 VCTRL2.t35 VSS 0.0395f
C693 VCTRL2.n18 VSS 0.0438f
C694 VCTRL2.t21 VSS 0.0228f
C695 VCTRL2.n19 VSS 0.0339f
C696 VCTRL2.n20 VSS 0.0339f
C697 VCTRL2.t12 VSS 0.0233f
C698 VCTRL2.n21 VSS 0.0449f
C699 VCTRL2.t25 VSS 0.0427f
C700 VCTRL2.n22 VSS 0.0449f
C701 VCTRL2.t43 VSS 0.045f
C702 VCTRL2.n23 VSS 0.0449f
C703 VCTRL2.t9 VSS 0.0395f
C704 VCTRL2.n24 VSS 0.0438f
C705 VCTRL2.t75 VSS 0.0228f
C706 VCTRL2.n25 VSS 0.0567f
C707 VCTRL2.n26 VSS 0.0335f
C708 VCTRL2.n27 VSS 0.0335f
C709 VCTRL2.t61 VSS 0.0233f
C710 VCTRL2.n28 VSS 0.0449f
C711 VCTRL2.t79 VSS 0.0427f
C712 VCTRL2.n29 VSS 0.0449f
C713 VCTRL2.t19 VSS 0.045f
C714 VCTRL2.n30 VSS 0.0449f
C715 VCTRL2.t60 VSS 0.0395f
C716 VCTRL2.n31 VSS 0.0438f
C717 VCTRL2.t68 VSS 0.0228f
C718 VCTRL2.n32 VSS 0.0567f
C719 VCTRL2.n33 VSS 0.0567f
C720 VCTRL2.t56 VSS 0.0233f
C721 VCTRL2.n34 VSS 0.0449f
C722 VCTRL2.t71 VSS 0.0427f
C723 VCTRL2.n35 VSS 0.0449f
C724 VCTRL2.t13 VSS 0.045f
C725 VCTRL2.n36 VSS 0.0449f
C726 VCTRL2.t55 VSS 0.0395f
C727 VCTRL2.n37 VSS 0.0438f
C728 VCTRL2.t8 VSS 0.0227f
C729 VCTRL2.t77 VSS 0.0235f
C730 VCTRL2.n38 VSS 0.0474f
C731 VCTRL2.t14 VSS 0.0427f
C732 VCTRL2.n39 VSS 0.0474f
C733 VCTRL2.t30 VSS 0.045f
C734 VCTRL2.n40 VSS 0.0474f
C735 VCTRL2.t73 VSS 0.0395f
C736 VCTRL2.n41 VSS 0.0464f
C737 VCTRL2.n42 VSS 0.0567f
C738 VCTRL2.n43 VSS 0.0335f
C739 VCTRL2.n44 VSS 0.0339f
C740 VCTRL2.n45 VSS 0.0337f
C741 VCTRL2.n46 VSS 0.0336f
C742 VCTRL2.t37 VSS 0.0227f
C743 VCTRL2.n47 VSS 0.0587f
C744 VCTRL2.n48 VSS 0.0587f
C745 VCTRL2.t24 VSS 0.0235f
C746 VCTRL2.n49 VSS 0.0449f
C747 VCTRL2.t39 VSS 0.0427f
C748 VCTRL2.n50 VSS 0.0587f
C749 VCTRL2.n51 VSS 0.0449f
C750 VCTRL2.t59 VSS 0.045f
C751 VCTRL2.n52 VSS 0.0449f
C752 VCTRL2.t22 VSS 0.0395f
C753 VCTRL2.n53 VSS 0.0438f
C754 VCTRL2.n54 VSS 0.0347f
C755 VCTRL2.t63 VSS 0.0228f
C756 VCTRL2.t52 VSS 0.0233f
C757 VCTRL2.n55 VSS 0.0478f
C758 VCTRL2.t67 VSS 0.0427f
C759 VCTRL2.n56 VSS 0.0478f
C760 VCTRL2.t5 VSS 0.045f
C761 VCTRL2.n57 VSS 0.0478f
C762 VCTRL2.t51 VSS 0.0395f
C763 VCTRL2.n58 VSS 0.0438f
C764 VCTRL2.n59 VSS 0.0544f
C765 VCTRL2.n60 VSS 0.0391f
C766 VCTRL2.n61 VSS 0.015f
C767 VCTRL2.n62 VSS 0.0313f
C768 VCTRL2.n63 VSS 0.931f
C769 VCTRL2.n64 VSS 0.148f
C770 VCTRL2.n65 VSS 1.88f
C771 VCTRL2.t33 VSS 0.0233f
C772 VCTRL2.n66 VSS 0.0336f
C773 VCTRL2.n67 VSS 0.0449f
C774 VCTRL2.t15 VSS 0.0427f
C775 VCTRL2.n68 VSS 0.0449f
C776 VCTRL2.t74 VSS 0.045f
C777 VCTRL2.n69 VSS 0.0336f
C778 VCTRL2.n70 VSS 0.0449f
C779 VCTRL2.t34 VSS 0.0395f
C780 VCTRL2.t17 VSS 0.0228f
C781 VCTRL2.n71 VSS 0.0438f
C782 VCTRL2.t46 VSS 0.0235f
C783 VCTRL2.n72 VSS 0.0449f
C784 VCTRL2.t26 VSS 0.0427f
C785 VCTRL2.n73 VSS 0.0449f
C786 VCTRL2.t10 VSS 0.045f
C787 VCTRL2.n74 VSS 0.0449f
C788 VCTRL2.t48 VSS 0.0395f
C789 VCTRL2.t29 VSS 0.0227f
C790 VCTRL2.n75 VSS 0.0438f
C791 VCTRL2.t76 VSS 0.0235f
C792 VCTRL2.n76 VSS 0.0449f
C793 VCTRL2.t57 VSS 0.0427f
C794 VCTRL2.n77 VSS 0.0449f
C795 VCTRL2.t36 VSS 0.045f
C796 VCTRL2.n78 VSS 0.0567f
C797 VCTRL2.n79 VSS 0.0449f
C798 VCTRL2.t78 VSS 0.0395f
C799 VCTRL2.t58 VSS 0.0227f
C800 VCTRL2.n80 VSS 0.0438f
C801 VCTRL2.t1 VSS 0.0236f
C802 VCTRL2.n81 VSS 0.0474f
C803 VCTRL2.t62 VSS 0.0427f
C804 VCTRL2.n82 VSS 0.0474f
C805 VCTRL2.t42 VSS 0.045f
C806 VCTRL2.n83 VSS 0.0474f
C807 VCTRL2.t2 VSS 0.0395f
C808 VCTRL2.t64 VSS 0.0226f
C809 VCTRL2.n84 VSS 0.0464f
C810 VCTRL2.n85 VSS 0.0567f
C811 VCTRL2.t47 VSS 0.0235f
C812 VCTRL2.n86 VSS 0.0449f
C813 VCTRL2.t27 VSS 0.0427f
C814 VCTRL2.n87 VSS 0.0449f
C815 VCTRL2.t11 VSS 0.045f
C816 VCTRL2.n88 VSS 0.0449f
C817 VCTRL2.t49 VSS 0.0395f
C818 VCTRL2.t31 VSS 0.0227f
C819 VCTRL2.n89 VSS 0.0438f
C820 VCTRL2.n90 VSS 0.0336f
C821 VCTRL2.n91 VSS 0.0338f
C822 VCTRL2.t40 VSS 0.0233f
C823 VCTRL2.n92 VSS 0.0567f
C824 VCTRL2.n93 VSS 0.0336f
C825 VCTRL2.n94 VSS 0.0338f
C826 VCTRL2.n95 VSS 0.0337f
C827 VCTRL2.n96 VSS 0.0449f
C828 VCTRL2.t20 VSS 0.0427f
C829 VCTRL2.n97 VSS 0.0449f
C830 VCTRL2.t0 VSS 0.045f
C831 VCTRL2.n98 VSS 0.0336f
C832 VCTRL2.n99 VSS 0.0338f
C833 VCTRL2.n100 VSS 0.0337f
C834 VCTRL2.n101 VSS 0.0449f
C835 VCTRL2.t41 VSS 0.0395f
C836 VCTRL2.t23 VSS 0.0228f
C837 VCTRL2.n102 VSS 0.0438f
C838 VCTRL2.n103 VSS 0.0337f
C839 VCTRL2.n104 VSS 0.0336f
C840 VCTRL2.t4 VSS 0.0236f
C841 VCTRL2.n105 VSS 0.0588f
C842 VCTRL2.n106 VSS 0.0449f
C843 VCTRL2.t66 VSS 0.0427f
C844 VCTRL2.n107 VSS 0.0567f
C845 VCTRL2.n108 VSS 0.0336f
C846 VCTRL2.n109 VSS 0.0338f
C847 VCTRL2.n110 VSS 0.0337f
C848 VCTRL2.n111 VSS 0.0336f
C849 VCTRL2.n112 VSS 0.0588f
C850 VCTRL2.n113 VSS 0.0449f
C851 VCTRL2.t45 VSS 0.045f
C852 VCTRL2.n114 VSS 0.0588f
C853 VCTRL2.n115 VSS 0.0449f
C854 VCTRL2.t7 VSS 0.0395f
C855 VCTRL2.t70 VSS 0.0226f
C856 VCTRL2.n116 VSS 0.0438f
C857 VCTRL2.n117 VSS 0.0347f
C858 VCTRL2.t3 VSS 0.0235f
C859 VCTRL2.n118 VSS 0.0478f
C860 VCTRL2.t65 VSS 0.0427f
C861 VCTRL2.n119 VSS 0.0478f
C862 VCTRL2.t44 VSS 0.045f
C863 VCTRL2.n120 VSS 0.0478f
C864 VCTRL2.t6 VSS 0.0395f
C865 VCTRL2.t69 VSS 0.0227f
C866 VCTRL2.n121 VSS 0.0438f
C867 VCTRL2.n122 VSS 0.0531f
C868 VCTRL2.n123 VSS 0.902f
C869 VCTRL2.n124 VSS 0.00725f
C870 VCTRL2.n125 VSS 0.0635f
C871 DFF_3_mag_0.INV_2_1.IN.n0 VSS 0.175f
C872 DFF_3_mag_0.INV_2_1.IN.n1 VSS 0.175f
C873 DFF_3_mag_0.INV_2_1.IN.t12 VSS 0.00891f
C874 DFF_3_mag_0.INV_2_1.IN.n2 VSS 0.00891f
C875 DFF_3_mag_0.INV_2_1.IN.n3 VSS 0.0279f
C876 DFF_3_mag_0.INV_2_1.IN.t13 VSS 0.00891f
C877 DFF_3_mag_0.INV_2_1.IN.n4 VSS 0.00891f
C878 DFF_3_mag_0.INV_2_1.IN.n5 VSS 0.0179f
C879 DFF_3_mag_0.INV_2_1.IN.n6 VSS 0.0904f
C880 DFF_3_mag_0.INV_2_1.IN.n7 VSS 0.0164f
C881 DFF_3_mag_0.INV_2_1.IN.t0 VSS 0.018f
C882 DFF_3_mag_0.INV_2_1.IN.n8 VSS 0.0652f
C883 DFF_3_mag_0.INV_2_1.IN.n9 VSS 0.022f
C884 DFF_3_mag_0.INV_2_1.IN.n10 VSS 0.0467f
C885 DFF_3_mag_0.INV_2_1.IN.n11 VSS 0.158f
C886 DFF_3_mag_0.INV_2_1.IN.t6 VSS 0.00891f
C887 DFF_3_mag_0.INV_2_1.IN.n12 VSS 0.00891f
C888 DFF_3_mag_0.INV_2_1.IN.n13 VSS 0.0179f
C889 DFF_3_mag_0.INV_2_1.IN.t7 VSS 0.00891f
C890 DFF_3_mag_0.INV_2_1.IN.n14 VSS 0.00891f
C891 DFF_3_mag_0.INV_2_1.IN.n15 VSS 0.0279f
C892 DFF_3_mag_0.INV_2_1.IN.n16 VSS 0.0904f
C893 DFF_3_mag_0.INV_2_1.IN.n17 VSS 0.0164f
C894 DFF_3_mag_0.INV_2_1.IN.t8 VSS 0.018f
C895 DFF_3_mag_0.INV_2_1.IN.n18 VSS 0.0652f
C896 DFF_3_mag_0.INV_2_1.IN.n19 VSS 0.022f
C897 DFF_3_mag_0.INV_2_1.IN.n20 VSS 0.0467f
C898 DFF_3_mag_0.INV_2_1.IN.n21 VSS 0.158f
C899 DFF_3_mag_0.INV_2_1.IN.t25 VSS 0.0279f
C900 DFF_3_mag_0.INV_2_1.IN.t27 VSS 0.0133f
C901 DFF_3_mag_0.INV_2_1.IN.n22 VSS 0.043f
C902 DFF_3_mag_0.INV_2_1.IN.n23 VSS 0.0306f
C903 DFF_3_mag_0.INV_2_1.IN.t16 VSS 0.0324f
C904 DFF_3_mag_0.INV_2_1.IN.n24 VSS 0.0372f
C905 DFF_3_mag_0.INV_2_1.IN.t21 VSS 0.0133f
C906 DFF_3_mag_0.INV_2_1.IN.n25 VSS 0.0379f
C907 DFF_3_mag_0.INV_2_1.IN.t22 VSS 0.0324f
C908 DFF_3_mag_0.INV_2_1.IN.n26 VSS 0.0306f
C909 DFF_3_mag_0.INV_2_1.IN.t17 VSS 0.0426f
C910 DFF_3_mag_0.INV_2_1.IN.t23 VSS 0.0175f
C911 DFF_3_mag_0.INV_2_1.IN.n27 VSS 0.0469f
C912 DFF_3_mag_0.INV_2_1.IN.t20 VSS 0.0426f
C913 DFF_3_mag_0.INV_2_1.IN.n28 VSS 0.0469f
C914 DFF_3_mag_0.INV_2_1.IN.t26 VSS 0.0175f
C915 DFF_3_mag_0.INV_2_1.IN.n29 VSS 0.0372f
C916 DFF_3_mag_0.INV_2_1.IN.t19 VSS 0.0324f
C917 DFF_3_mag_0.INV_2_1.IN.t18 VSS 0.0133f
C918 DFF_3_mag_0.INV_2_1.IN.n30 VSS 0.043f
C919 DFF_3_mag_0.INV_2_1.IN.t24 VSS 0.0132f
C920 DFF_3_mag_0.INV_2_1.IN.n31 VSS 0.0217f
C921 DFF_3_mag_0.INV_2_1.IN.n32 VSS 0.0219f
C922 DFF_3_mag_0.INV_2_1.IN.n33 VSS 0.271f
C923 VCO_C_0.INV_2_5.IN.n0 VSS 0.562f
C924 VCO_C_0.INV_2_5.IN.n1 VSS 0.144f
C925 VCO_C_0.INV_2_5.IN.n2 VSS 0.4f
C926 VCO_C_0.INV_2_5.IN.n3 VSS 0.286f
C927 VCO_C_0.INV_2_5.IN.n4 VSS 0.557f
C928 VCO_C_0.INV_2_5.IN.n5 VSS 0.674f
C929 VCO_C_0.INV_2_5.IN.n6 VSS 0.835f
C930 VCO_C_0.INV_2_5.IN.t39 VSS 0.0904f
C931 VCO_C_0.INV_2_5.IN.t41 VSS 0.0429f
C932 VCO_C_0.INV_2_5.IN.n7 VSS 0.139f
C933 VCO_C_0.INV_2_5.IN.n8 VSS 0.0991f
C934 VCO_C_0.INV_2_5.IN.t44 VSS 0.105f
C935 VCO_C_0.INV_2_5.IN.n9 VSS 0.12f
C936 VCO_C_0.INV_2_5.IN.t54 VSS 0.0429f
C937 VCO_C_0.INV_2_5.IN.n10 VSS 0.123f
C938 VCO_C_0.INV_2_5.IN.t58 VSS 0.105f
C939 VCO_C_0.INV_2_5.IN.n11 VSS 0.0991f
C940 VCO_C_0.INV_2_5.IN.t43 VSS 0.138f
C941 VCO_C_0.INV_2_5.IN.t31 VSS 0.0568f
C942 VCO_C_0.INV_2_5.IN.n12 VSS 0.152f
C943 VCO_C_0.INV_2_5.IN.t51 VSS 0.138f
C944 VCO_C_0.INV_2_5.IN.n13 VSS 0.152f
C945 VCO_C_0.INV_2_5.IN.t38 VSS 0.0568f
C946 VCO_C_0.INV_2_5.IN.n14 VSS 0.12f
C947 VCO_C_0.INV_2_5.IN.t50 VSS 0.105f
C948 VCO_C_0.INV_2_5.IN.t46 VSS 0.0429f
C949 VCO_C_0.INV_2_5.IN.n15 VSS 0.139f
C950 VCO_C_0.INV_2_5.IN.t35 VSS 0.0428f
C951 VCO_C_0.INV_2_5.IN.n16 VSS 0.0703f
C952 VCO_C_0.INV_2_5.IN.n17 VSS 0.0776f
C953 VCO_C_0.INV_2_5.IN.n18 VSS 1.02f
C954 VCO_C_0.INV_2_5.IN.n19 VSS 0.0296f
C955 VCO_C_0.INV_2_5.IN.n20 VSS 0.0296f
C956 VCO_C_0.INV_2_5.IN.n21 VSS 0.0186f
C957 VCO_C_0.INV_2_5.IN.t4 VSS 0.0158f
C958 VCO_C_0.INV_2_5.IN.n22 VSS 0.14f
C959 VCO_C_0.INV_2_5.IN.n23 VSS 0.0449f
C960 VCO_C_0.INV_2_5.IN.n24 VSS 0.739f
C961 VCO_C_0.INV_2_5.IN.n25 VSS 0.303f
C962 VCO_C_0.INV_2_5.IN.n26 VSS 0.42f
C963 VCO_C_0.INV_2_5.IN.n27 VSS 0.0186f
C964 VCO_C_0.INV_2_5.IN.t3 VSS 0.0158f
C965 VCO_C_0.INV_2_5.IN.n28 VSS 0.162f
C966 VCO_C_0.INV_2_5.IN.n29 VSS 0.757f
C967 VCO_C_0.INV_2_5.IN.t5 VSS 0.205f
C968 VCO_C_0.INV_2_5.IN.t2 VSS 0.029f
C969 VCO_C_0.INV_2_5.IN.n30 VSS 0.683f
C970 VCO_C_0.INV_2_5.IN.t6 VSS 0.0265f
C971 VCO_C_0.INV_2_5.IN.n31 VSS 0.251f
C972 VCO_C_0.INV_2_5.IN.n32 VSS 0.405f
C973 VCO_C_0.INV_2_5.IN.n33 VSS 0.479f
C974 VCO_C_0.INV_2_5.IN.n34 VSS 0.905f
C975 VCO_C_0.INV_2_5.IN.t26 VSS 0.0172f
C976 VCO_C_0.INV_2_5.IN.n35 VSS 0.0172f
C977 VCO_C_0.INV_2_5.IN.n36 VSS 0.0345f
C978 VCO_C_0.INV_2_5.IN.n37 VSS 0.0387f
C979 VCO_C_0.INV_2_5.IN.n38 VSS 0.0602f
C980 VCO_C_0.INV_2_5.IN.t24 VSS 0.0277f
C981 VCO_C_0.INV_2_5.IN.n39 VSS 0.0692f
C982 VCO_C_0.INV_2_5.IN.n40 VSS 0.0523f
C983 VCO_C_0.INV_2_5.IN.n41 VSS 0.0243f
C984 VCO_C_0.INV_2_5.IN.n42 VSS 0.0726f
C985 VCO_C_0.INV_2_5.IN.n43 VSS 0.0515f
C986 VCO_C_0.INV_2_5.IN.n44 VSS 0.528f
C987 VCO_C_0.INV_2_5.IN.n45 VSS 0.049f
C988 VCO_C_0.INV_2_5.IN.n46 VSS 0.0301f
C989 VCO_C_0.INV_2_5.IN.n47 VSS 0.0815f
C990 VCO_C_0.INV_2_5.IN.t15 VSS 0.0172f
C991 VCO_C_0.INV_2_5.IN.n48 VSS 0.0172f
C992 VCO_C_0.INV_2_5.IN.n49 VSS 0.0345f
C993 VCO_C_0.INV_2_5.IN.n50 VSS 0.0387f
C994 VCO_C_0.INV_2_5.IN.n51 VSS 0.0515f
C995 VCO_C_0.INV_2_5.IN.n52 VSS 0.35f
C996 VCO_C_0.INV_2_5.IN.n53 VSS 0.0529f
C997 VCO_C_0.INV_2_5.IN.t28 VSS 0.0172f
C998 VCO_C_0.INV_2_5.IN.n54 VSS 0.0172f
C999 VCO_C_0.INV_2_5.IN.n55 VSS 0.0346f
C1000 VCO_C_0.INV_2_5.IN.n56 VSS 0.0509f
C1001 VCO_C_0.INV_2_5.IN.t13 VSS 0.0699f
C1002 VCO_C_0.INV_2_5.IN.n57 VSS 0.58f
C1003 VCO_C_0.INV_2_5.IN.n58 VSS 0.491f
C1004 VCO_C_0.INV_2_5.IN.n59 VSS 0.0277f
C1005 VCO_C_0.INV_2_5.IN.n60 VSS 0.278f
C1006 VCO_C_0.INV_2_5.IN.n61 VSS 0.82f
C1007 VCO_C_0.INV_2_5.IN.t45 VSS 0.117f
C1008 VCO_C_0.INV_2_5.IN.t48 VSS 0.122f
C1009 VCO_C_0.INV_2_5.IN.t49 VSS 0.122f
C1010 VCO_C_0.INV_2_5.IN.t32 VSS 0.116f
C1011 VCO_C_0.INV_2_5.IN.t52 VSS 0.12f
C1012 VCO_C_0.INV_2_5.IN.t53 VSS 0.125f
C1013 VCO_C_0.INV_2_5.IN.t36 VSS 0.125f
C1014 VCO_C_0.INV_2_5.IN.t57 VSS 0.129f
C1015 VCO_C_0.INV_2_5.IN.n62 VSS 0.512f
C1016 VCO_C_0.INV_2_5.IN.n63 VSS 0.269f
C1017 VCO_C_0.INV_2_5.IN.n64 VSS 0.329f
C1018 VCO_C_0.INV_2_5.IN.n65 VSS 0.322f
C1019 VCO_C_0.INV_2_5.IN.n66 VSS 0.269f
C1020 VCO_C_0.INV_2_5.IN.n67 VSS 0.275f
C1021 VCO_C_0.INV_2_5.IN.t34 VSS 0.118f
C1022 VCO_C_0.INV_2_5.IN.t55 VSS 0.123f
C1023 VCO_C_0.INV_2_5.IN.t56 VSS 0.123f
C1024 VCO_C_0.INV_2_5.IN.t42 VSS 0.119f
C1025 VCO_C_0.INV_2_5.IN.t33 VSS 0.123f
C1026 VCO_C_0.INV_2_5.IN.t40 VSS 0.123f
C1027 VCO_C_0.INV_2_5.IN.t47 VSS 0.123f
C1028 VCO_C_0.INV_2_5.IN.t37 VSS 0.142f
C1029 VCO_C_0.INV_2_5.IN.n68 VSS 0.495f
C1030 VCO_C_0.INV_2_5.IN.n69 VSS 0.263f
C1031 VCO_C_0.INV_2_5.IN.n70 VSS 0.297f
C1032 VCO_C_0.INV_2_5.IN.t30 VSS 0.0407f
C1033 VCO_C_0.INV_2_5.IN.n71 VSS 0.275f
C1034 VCO_C_0.INV_2_5.IN.n72 VSS 0.271f
C1035 VCO_C_0.INV_2_5.IN.n73 VSS 0.0243f
C1036 VCO_C_0.INV_2_5.IN.n74 VSS 0.28f
C1037 VCO_C_0.INV_2_5.IN.n75 VSS 0.0734f
C1038 VCO_C_0.INV_2_5.IN.n76 VSS 0.436f
C1039 VCO_C_0.INV_2_5.IN.n77 VSS 0.506f
C1040 VCO_C_0.INV_2_5.IN.n78 VSS 0.351f
C1041 VCO_C_0.INV_2_5.IN.n79 VSS 0.0177f
C1042 VCO_C_0.INV_2_5.IN.t18 VSS 0.0164f
C1043 VCO_C_0.INV_2_5.IN.n80 VSS 0.139f
C1044 VCO_C_0.INV_2_5.IN.t20 VSS 0.0413f
C1045 VCO_C_0.INV_2_5.IN.n81 VSS 0.579f
C1046 VCO_C_0.INV_2_5.IN.t19 VSS 0.0409f
C1047 VCO_C_0.INV_2_5.IN.n82 VSS 0.0276f
C1048 VCO_C_0.INV_2_5.IN.n83 VSS 0.0978f
C1049 VCO_C_0.INV_2_5.IN.t25 VSS 0.0243f
C1050 VCO_C_0.INV_2_5.IN.n84 VSS 0.143f
C1051 VCO_C_0.INV_2_5.IN.n85 VSS 0.0345f
C1052 VCO_C_0.INV_2_5.IN.n86 VSS 0.0159f
C1053 VCO_C_0.INV_2_5.IN.t11 VSS 0.0184f
C1054 VCO_C_0.OUTB.n0 VSS 0.0359f
C1055 VCO_C_0.OUTB.n1 VSS 0.0163f
C1056 VCO_C_0.OUTB.n2 VSS 2.18f
C1057 VCO_C_0.OUTB.t8 VSS 0.00227f
C1058 VCO_C_0.OUTB.n3 VSS 0.00227f
C1059 VCO_C_0.OUTB.n4 VSS 0.00509f
C1060 VCO_C_0.OUTB.t1 VSS 0.00227f
C1061 VCO_C_0.OUTB.n5 VSS 0.00227f
C1062 VCO_C_0.OUTB.n6 VSS 0.00453f
C1063 VCO_C_0.OUTB.t5 VSS 0.00227f
C1064 VCO_C_0.OUTB.n7 VSS 0.00227f
C1065 VCO_C_0.OUTB.n8 VSS 0.00553f
C1066 VCO_C_0.OUTB.n9 VSS 0.0123f
C1067 VCO_C_0.OUTB.t9 VSS 0.00227f
C1068 VCO_C_0.OUTB.n10 VSS 0.00227f
C1069 VCO_C_0.OUTB.n11 VSS 0.00509f
C1070 VCO_C_0.OUTB.t3 VSS 0.00227f
C1071 VCO_C_0.OUTB.n12 VSS 0.00227f
C1072 VCO_C_0.OUTB.n13 VSS 0.00553f
C1073 VCO_C_0.OUTB.t2 VSS 0.00227f
C1074 VCO_C_0.OUTB.n14 VSS 0.00227f
C1075 VCO_C_0.OUTB.n15 VSS 0.00453f
C1076 VCO_C_0.OUTB.n16 VSS 0.0123f
C1077 VCO_C_0.OUTB.n17 VSS 0.0196f
C1078 VCO_C_0.OUTB.n18 VSS 0.0244f
C1079 VCO_C_0.OUTB.t25 VSS 0.00714f
C1080 VCO_C_0.OUTB.t20 VSS 0.0183f
C1081 VCO_C_0.OUTB.n19 VSS 0.0213f
C1082 VCO_C_0.OUTB.t21 VSS 0.00714f
C1083 VCO_C_0.OUTB.t27 VSS 0.00714f
C1084 VCO_C_0.OUTB.t14 VSS 0.0167f
C1085 VCO_C_0.OUTB.t17 VSS 0.0319f
C1086 VCO_C_0.OUTB.n20 VSS 0.0236f
C1087 VCO_C_0.OUTB.n21 VSS 0.0173f
C1088 VCO_C_0.OUTB.n22 VSS 0.0576f
C1089 VCO_C_0.OUTB.t34 VSS 0.00714f
C1090 VCO_C_0.OUTB.t42 VSS 0.00714f
C1091 VCO_C_0.OUTB.t19 VSS 0.0178f
C1092 VCO_C_0.OUTB.n23 VSS 0.0205f
C1093 VCO_C_0.OUTB.n24 VSS 0.0205f
C1094 VCO_C_0.OUTB.t53 VSS 0.0259f
C1095 VCO_C_0.OUTB.n25 VSS 0.111f
C1096 VCO_C_0.OUTB.t37 VSS 0.00714f
C1097 VCO_C_0.OUTB.t15 VSS 0.00714f
C1098 VCO_C_0.OUTB.t13 VSS 0.0167f
C1099 VCO_C_0.OUTB.t47 VSS 0.0319f
C1100 VCO_C_0.OUTB.n26 VSS 0.0236f
C1101 VCO_C_0.OUTB.n27 VSS 0.0178f
C1102 VCO_C_0.OUTB.t49 VSS 0.00714f
C1103 VCO_C_0.OUTB.t28 VSS 0.0183f
C1104 VCO_C_0.OUTB.n28 VSS 0.0213f
C1105 VCO_C_0.OUTB.t18 VSS 0.00714f
C1106 VCO_C_0.OUTB.t50 VSS 0.00714f
C1107 VCO_C_0.OUTB.t45 VSS 0.0178f
C1108 VCO_C_0.OUTB.n29 VSS 0.0205f
C1109 VCO_C_0.OUTB.n30 VSS 0.0205f
C1110 VCO_C_0.OUTB.t43 VSS 0.0269f
C1111 VCO_C_0.OUTB.n31 VSS 0.036f
C1112 VCO_C_0.OUTB.n32 VSS 0.0339f
C1113 VCO_C_0.OUTB.t48 VSS 0.00566f
C1114 VCO_C_0.OUTB.n33 VSS 0.00928f
C1115 VCO_C_0.OUTB.n34 VSS 0.0159f
C1116 VCO_C_0.OUTB.t52 VSS 0.00749f
C1117 VCO_C_0.OUTB.t46 VSS 0.0182f
C1118 VCO_C_0.OUTB.n35 VSS 0.0131f
C1119 VCO_C_0.OUTB.t16 VSS 0.00566f
C1120 VCO_C_0.OUTB.t24 VSS 0.0139f
C1121 VCO_C_0.OUTB.n36 VSS 0.0162f
C1122 VCO_C_0.OUTB.t36 VSS 0.00566f
C1123 VCO_C_0.OUTB.t26 VSS 0.00566f
C1124 VCO_C_0.OUTB.t33 VSS 0.0139f
C1125 VCO_C_0.OUTB.n37 VSS 0.0184f
C1126 VCO_C_0.OUTB.n38 VSS 0.0184f
C1127 VCO_C_0.OUTB.t44 VSS 0.0139f
C1128 VCO_C_0.OUTB.n39 VSS 0.0159f
C1129 VCO_C_0.OUTB.t23 VSS 0.00749f
C1130 VCO_C_0.OUTB.n40 VSS 0.02f
C1131 VCO_C_0.OUTB.n41 VSS 0.02f
C1132 VCO_C_0.OUTB.t32 VSS 0.0182f
C1133 VCO_C_0.OUTB.n42 VSS 0.0131f
C1134 VCO_C_0.OUTB.t51 VSS 0.0119f
C1135 VCO_C_0.OUTB.n43 VSS 0.00938f
C1136 VCO_C_0.OUTB.n44 VSS 0.016f
C1137 VCO_C_0.OUTB.n45 VSS 1.48f
C1138 VCO_C_0.OUTB.t38 VSS 0.0277f
C1139 VCO_C_0.OUTB.t39 VSS 0.0251f
C1140 VCO_C_0.OUTB.t40 VSS 0.0304f
C1141 VCO_C_0.OUTB.t12 VSS 0.0286f
C1142 VCO_C_0.OUTB.n46 VSS 0.0681f
C1143 VCO_C_0.OUTB.n47 VSS 0.0394f
C1144 VCO_C_0.OUTB.n48 VSS 0.0605f
C1145 VCO_C_0.OUTB.t22 VSS 0.0246f
C1146 VCO_C_0.OUTB.t30 VSS 0.0247f
C1147 VCO_C_0.OUTB.t31 VSS 0.0241f
C1148 VCO_C_0.OUTB.t41 VSS 0.0285f
C1149 VCO_C_0.OUTB.n49 VSS 0.0847f
C1150 VCO_C_0.OUTB.n50 VSS 0.0465f
C1151 VCO_C_0.OUTB.n51 VSS 0.045f
C1152 VCO_C_0.OUTB.n52 VSS 0.0555f
C1153 VCO_C_0.OUTB.t35 VSS 0.0244f
C1154 VCO_C_0.OUTB.t29 VSS 0.028f
C1155 VCO_C_0.OUTB.n53 VSS 0.0919f
C1156 VCO_C_0.OUTB.n54 VSS 0.0387f
C1157 VCO_C_0.OUTB.n55 VSS 0.0255f
C1158 VCO_C_0.OUTB.n56 VSS 0.00893f
C1159 VCO_C_0.INV_2_1.IN.t10 VSS 0.0111f
C1160 VCO_C_0.INV_2_1.IN.n0 VSS 0.0111f
C1161 VCO_C_0.INV_2_1.IN.n1 VSS 0.0249f
C1162 VCO_C_0.INV_2_1.IN.t4 VSS 0.0111f
C1163 VCO_C_0.INV_2_1.IN.n2 VSS 0.0111f
C1164 VCO_C_0.INV_2_1.IN.n3 VSS 0.0221f
C1165 VCO_C_0.INV_2_1.IN.t0 VSS 0.0111f
C1166 VCO_C_0.INV_2_1.IN.n4 VSS 0.0111f
C1167 VCO_C_0.INV_2_1.IN.n5 VSS 0.027f
C1168 VCO_C_0.INV_2_1.IN.n6 VSS 0.0599f
C1169 VCO_C_0.INV_2_1.IN.t9 VSS 0.0111f
C1170 VCO_C_0.INV_2_1.IN.n7 VSS 0.0111f
C1171 VCO_C_0.INV_2_1.IN.n8 VSS 0.0249f
C1172 VCO_C_0.INV_2_1.IN.t3 VSS 0.0111f
C1173 VCO_C_0.INV_2_1.IN.n9 VSS 0.0111f
C1174 VCO_C_0.INV_2_1.IN.n10 VSS 0.0221f
C1175 VCO_C_0.INV_2_1.IN.t5 VSS 0.0111f
C1176 VCO_C_0.INV_2_1.IN.n11 VSS 0.0111f
C1177 VCO_C_0.INV_2_1.IN.n12 VSS 0.027f
C1178 VCO_C_0.INV_2_1.IN.n13 VSS 0.0599f
C1179 VCO_C_0.INV_2_1.IN.n14 VSS 0.0958f
C1180 VCO_C_0.INV_2_1.IN.n15 VSS 0.119f
C1181 VCO_C_0.INV_2_1.IN.t21 VSS 0.0276f
C1182 VCO_C_0.INV_2_1.IN.n16 VSS 0.0453f
C1183 VCO_C_0.INV_2_1.IN.n17 VSS 0.0776f
C1184 VCO_C_0.INV_2_1.IN.t17 VSS 0.0366f
C1185 VCO_C_0.INV_2_1.IN.t14 VSS 0.0889f
C1186 VCO_C_0.INV_2_1.IN.n18 VSS 0.0639f
C1187 VCO_C_0.INV_2_1.IN.t12 VSS 0.0276f
C1188 VCO_C_0.INV_2_1.IN.t23 VSS 0.0676f
C1189 VCO_C_0.INV_2_1.IN.n19 VSS 0.0791f
C1190 VCO_C_0.INV_2_1.IN.t22 VSS 0.0276f
C1191 VCO_C_0.INV_2_1.IN.t16 VSS 0.0276f
C1192 VCO_C_0.INV_2_1.IN.t13 VSS 0.0676f
C1193 VCO_C_0.INV_2_1.IN.n20 VSS 0.0897f
C1194 VCO_C_0.INV_2_1.IN.n21 VSS 0.0897f
C1195 VCO_C_0.INV_2_1.IN.t20 VSS 0.0676f
C1196 VCO_C_0.INV_2_1.IN.n22 VSS 0.0776f
C1197 VCO_C_0.INV_2_1.IN.t15 VSS 0.0366f
C1198 VCO_C_0.INV_2_1.IN.n23 VSS 0.0977f
C1199 VCO_C_0.INV_2_1.IN.n24 VSS 0.0977f
C1200 VCO_C_0.INV_2_1.IN.t18 VSS 0.0889f
C1201 VCO_C_0.INV_2_1.IN.n25 VSS 0.0639f
C1202 VCO_C_0.INV_2_1.IN.t19 VSS 0.0582f
C1203 VCO_C_0.INV_2_1.IN.n26 VSS 0.0458f
C1204 VCTRL.t10 VSS 0.104f
C1205 VCTRL.t2 VSS 0.0317f
C1206 VCTRL.t0 VSS 0.166f
C1207 VCTRL.n0 VSS 0.235f
C1208 VCTRL.n1 VSS 0.655f
C1209 VCTRL.t3 VSS 0.0962f
C1210 VCTRL.n2 VSS 0.133f
C1211 VCTRL.t11 VSS 0.0317f
C1212 VCTRL.t8 VSS 0.165f
C1213 VCTRL.n3 VSS 0.164f
C1214 VCTRL.t13 VSS 0.106f
C1215 VCTRL.n4 VSS 0.147f
C1216 VCTRL.t18 VSS 0.121f
C1217 VCTRL.n5 VSS 0.495f
C1218 VCTRL.n6 VSS 0.515f
C1219 VCTRL.t7 VSS 0.1f
C1220 VCTRL.n7 VSS 0.255f
C1221 VCTRL.t16 VSS 0.0891f
C1222 VCTRL.n8 VSS 0.283f
C1223 VCTRL.n9 VSS 0.718f
C1224 VCTRL.n10 VSS 0.416f
C1225 VCTRL.n11 VSS 0.411f
C1226 VCTRL.n12 VSS 2.02f
C1227 VCTRL.t9 VSS 0.104f
C1228 VCTRL.t15 VSS 0.0317f
C1229 VCTRL.t19 VSS 0.166f
C1230 VCTRL.n13 VSS 0.235f
C1231 VCTRL.n14 VSS 0.655f
C1232 VCTRL.t5 VSS 0.0317f
C1233 VCTRL.t6 VSS 0.165f
C1234 VCTRL.n15 VSS 0.164f
C1235 VCTRL.n16 VSS 0.515f
C1236 VCTRL.t17 VSS 0.121f
C1237 VCTRL.n17 VSS 0.495f
C1238 VCTRL.t4 VSS 0.106f
C1239 VCTRL.n18 VSS 0.148f
C1240 VCTRL.t14 VSS 0.0962f
C1241 VCTRL.n19 VSS 0.133f
C1242 VCTRL.t1 VSS 0.0891f
C1243 VCTRL.t12 VSS 0.1f
C1244 VCTRL.n20 VSS 0.255f
C1245 VCTRL.n21 VSS 0.283f
C1246 VCTRL.n22 VSS 0.718f
C1247 VCTRL.n23 VSS 0.416f
C1248 VCTRL.n24 VSS 0.618f
C1249 VCTRL.n25 VSS 0.499f
C1250 VCTRL.n26 VSS 0.518f
C1251 VDD.n0 VSS 0.00913f
C1252 VDD.n1 VSS 0.00808f
C1253 VDD.n2 VSS 0.0518f
C1254 VDD.n3 VSS 0.0869f
C1255 VDD.n4 VSS 0.00527f
C1256 VDD.n5 VSS 0.0387f
C1257 VDD.n6 VSS 0.00516f
C1258 VDD.n7 VSS 0.0242f
C1259 VDD.n8 VSS 0.00129f
C1260 VDD.n9 VSS 0.0203f
C1261 VDD.n10 VSS 0.0816f
C1262 VDD.n11 VSS 6.86e-19
C1263 VDD.n12 VSS 0.0573f
C1264 VDD.n13 VSS 0.00611f
C1265 VDD.n14 VSS 0.00528f
C1266 VDD.n15 VSS 0.00696f
C1267 VDD.t169 VSS 0.049f
C1268 VDD.n16 VSS 0.0165f
C1269 VDD.n17 VSS 0.00511f
C1270 VDD.n18 VSS 0.00589f
C1271 VDD.n19 VSS 0.00222f
C1272 VDD.n20 VSS 0.0131f
C1273 VDD.n21 VSS 0.00129f
C1274 VDD.n22 VSS 0.041f
C1275 VDD.n23 VSS 0.00404f
C1276 VDD.n24 VSS 0.00415f
C1277 VDD.t153 VSS 0.00405f
C1278 VDD.n25 VSS 0.00405f
C1279 VDD.n26 VSS 0.0099f
C1280 VDD.t88 VSS 0.00405f
C1281 VDD.n27 VSS 0.00405f
C1282 VDD.n28 VSS 0.0081f
C1283 VDD.n29 VSS 0.0254f
C1284 VDD.n30 VSS 0.0159f
C1285 VDD.t84 VSS 0.0552f
C1286 VDD.n31 VSS 0.0552f
C1287 VDD.n32 VSS 0.0107f
C1288 VDD.t82 VSS 0.00929f
C1289 VDD.t83 VSS 0.00808f
C1290 VDD.n33 VSS 0.0384f
C1291 VDD.n34 VSS 0.214f
C1292 VDD.n35 VSS 0.0416f
C1293 VDD.t81 VSS 0.0591f
C1294 VDD.n36 VSS 0.0609f
C1295 VDD.n37 VSS 0.0107f
C1296 VDD.n38 VSS 0.0183f
C1297 VDD.n39 VSS 0.109f
C1298 VDD.n40 VSS 0.0107f
C1299 VDD.n41 VSS 0.0183f
C1300 VDD.n42 VSS 0.0183f
C1301 VDD.n43 VSS 0.107f
C1302 VDD.n44 VSS 0.0107f
C1303 VDD.t87 VSS 0.0547f
C1304 VDD.n45 VSS 0.0627f
C1305 VDD.n46 VSS 0.0107f
C1306 VDD.n47 VSS 0.0176f
C1307 VDD.n48 VSS 0.0461f
C1308 VDD.n49 VSS 0.00544f
C1309 VDD.n50 VSS 0.00937f
C1310 VDD.n51 VSS 0.0131f
C1311 VDD.n52 VSS 0.00129f
C1312 VDD.n53 VSS 0.00222f
C1313 VDD.n54 VSS 0.0433f
C1314 VDD.n55 VSS 0.00426f
C1315 VDD.n56 VSS 0.00454f
C1316 VDD.n57 VSS 0.0028f
C1317 VDD.n58 VSS 0.0028f
C1318 VDD.n59 VSS 0.00504f
C1319 VDD.n60 VSS 0.0023f
C1320 VDD.n61 VSS 0.0023f
C1321 VDD.n62 VSS 0.00246f
C1322 VDD.n63 VSS 0.00525f
C1323 VDD.n64 VSS 0.0058f
C1324 VDD.n65 VSS 0.00234f
C1325 VDD.n66 VSS 0.00392f
C1326 VDD.n67 VSS 0.00556f
C1327 VDD.n68 VSS 0.0052f
C1328 VDD.n69 VSS 0.0208f
C1329 VDD.n70 VSS 0.0238f
C1330 VDD.n71 VSS 0.0113f
C1331 VDD.n72 VSS 0.00808f
C1332 VDD.n73 VSS 0.00929f
C1333 VDD.n74 VSS 0.0373f
C1334 VDD.n75 VSS 0.00913f
C1335 VDD.n76 VSS 0.00808f
C1336 VDD.n77 VSS 0.0508f
C1337 VDD.n78 VSS 0.226f
C1338 VDD.n79 VSS 0.0441f
C1339 VDD.n80 VSS 0.0219f
C1340 VDD.n81 VSS 0.112f
C1341 VDD.n82 VSS 0.0121f
C1342 VDD.n83 VSS 0.0052f
C1343 VDD.n84 VSS 0.00308f
C1344 VDD.n85 VSS 0.0182f
C1345 VDD.n86 VSS 0.00527f
C1346 VDD.n87 VSS 0.0262f
C1347 VDD.n88 VSS 0.00129f
C1348 VDD.n89 VSS 0.00443f
C1349 VDD.n90 VSS 0.0775f
C1350 VDD.n91 VSS 0.00544f
C1351 VDD.n92 VSS 0.00753f
C1352 VDD.n93 VSS 0.00577f
C1353 VDD.n94 VSS 0.0182f
C1354 VDD.n95 VSS 0.00432f
C1355 VDD.t346 VSS 0.00405f
C1356 VDD.n96 VSS 0.00405f
C1357 VDD.n97 VSS 0.0099f
C1358 VDD.t418 VSS 0.00405f
C1359 VDD.n98 VSS 0.00405f
C1360 VDD.n99 VSS 0.0081f
C1361 VDD.n100 VSS 0.0275f
C1362 VDD.t180 VSS 0.0216f
C1363 VDD.n101 VSS 0.0923f
C1364 VDD.n102 VSS 0.0107f
C1365 VDD.t423 VSS 0.00929f
C1366 VDD.t185 VSS 0.00808f
C1367 VDD.n103 VSS 0.0373f
C1368 VDD.n104 VSS 0.227f
C1369 VDD.t337 VSS 0.00808f
C1370 VDD.t59 VSS 0.00913f
C1371 VDD.n105 VSS 0.0503f
C1372 VDD.n106 VSS 0.0109f
C1373 VDD.n107 VSS 0.0138f
C1374 VDD.t347 VSS 0.00681f
C1375 VDD.n108 VSS 0.00681f
C1376 VDD.n109 VSS 0.0147f
C1377 VDD.n110 VSS 0.0218f
C1378 VDD.n111 VSS 0.0796f
C1379 VDD.t57 VSS 0.0168f
C1380 VDD.n112 VSS 0.0435f
C1381 VDD.t78 VSS 0.34f
C1382 VDD.n113 VSS 0.355f
C1383 VDD.t76 VSS 0.349f
C1384 VDD.n114 VSS 0.331f
C1385 VDD.t77 VSS 0.341f
C1386 VDD.t56 VSS 0.337f
C1387 VDD.n115 VSS 0.331f
C1388 VDD.n116 VSS 0.0863f
C1389 VDD.n117 VSS 0.0415f
C1390 VDD.n118 VSS 0.524f
C1391 VDD.t90 VSS 0.00681f
C1392 VDD.n119 VSS 0.00681f
C1393 VDD.n120 VSS 0.0147f
C1394 VDD.n121 VSS 0.0218f
C1395 VDD.n122 VSS 0.0819f
C1396 VDD.n123 VSS 0.0601f
C1397 VDD.n124 VSS 0.0055f
C1398 VDD.n125 VSS 0.00618f
C1399 VDD.t60 VSS 0.0157f
C1400 VDD.n126 VSS 0.0209f
C1401 VDD.n127 VSS 0.0156f
C1402 VDD.n128 VSS 0.235f
C1403 VDD.n129 VSS 0.0139f
C1404 VDD.n130 VSS 0.0108f
C1405 VDD.n131 VSS 0.0119f
C1406 VDD.n132 VSS 0.184f
C1407 VDD.n133 VSS 0.0123f
C1408 VDD.n134 VSS 0.0427f
C1409 VDD.n135 VSS 0.0117f
C1410 VDD.n136 VSS 0.0115f
C1411 VDD.n137 VSS 0.0117f
C1412 VDD.n138 VSS 0.00873f
C1413 VDD.n139 VSS 0.00242f
C1414 VDD.n140 VSS 0.0086f
C1415 VDD.n141 VSS 0.00269f
C1416 VDD.n142 VSS 0.00242f
C1417 VDD.n143 VSS 0.00346f
C1418 VDD.n144 VSS 0.12f
C1419 VDD.n145 VSS 0.0121f
C1420 VDD.n146 VSS 0.00346f
C1421 VDD.n147 VSS 0.0957f
C1422 VDD.n148 VSS 0.0107f
C1423 VDD.n149 VSS 0.00481f
C1424 VDD.n150 VSS 0.015f
C1425 VDD.t58 VSS 0.0889f
C1426 VDD.n151 VSS 0.033f
C1427 VDD.n152 VSS 0.0107f
C1428 VDD.n153 VSS 0.0169f
C1429 VDD.n154 VSS 0.11f
C1430 VDD.n155 VSS 0.0107f
C1431 VDD.n156 VSS 0.0187f
C1432 VDD.n157 VSS 0.107f
C1433 VDD.n158 VSS 0.0107f
C1434 VDD.n159 VSS 0.0181f
C1435 VDD.n160 VSS 0.107f
C1436 VDD.n161 VSS 0.0107f
C1437 VDD.n162 VSS 0.0181f
C1438 VDD.n163 VSS 0.0187f
C1439 VDD.n164 VSS 0.0158f
C1440 VDD.t321 VSS 0.00405f
C1441 VDD.n165 VSS 0.00405f
C1442 VDD.n166 VSS 0.0081f
C1443 VDD.t322 VSS 0.00405f
C1444 VDD.n167 VSS 0.00405f
C1445 VDD.n168 VSS 0.0099f
C1446 VDD.n169 VSS 0.0275f
C1447 VDD.n170 VSS 0.107f
C1448 VDD.n171 VSS 0.0107f
C1449 VDD.n172 VSS 0.0934f
C1450 VDD.n173 VSS 0.0107f
C1451 VDD.n174 VSS 0.0145f
C1452 VDD.n175 VSS 0.00558f
C1453 VDD.n176 VSS 0.00636f
C1454 VDD.n177 VSS 0.00667f
C1455 VDD.n178 VSS 0.107f
C1456 VDD.n179 VSS 0.01f
C1457 VDD.n180 VSS 0.0889f
C1458 VDD.n181 VSS 0.00527f
C1459 VDD.n182 VSS 0.0262f
C1460 VDD.n183 VSS 0.00129f
C1461 VDD.n184 VSS 0.00443f
C1462 VDD.n185 VSS 0.00366f
C1463 VDD.t320 VSS 0.00911f
C1464 VDD.n186 VSS 0.0695f
C1465 VDD.n187 VSS 0.0107f
C1466 VDD.n188 VSS 0.0127f
C1467 VDD.n189 VSS 0.015f
C1468 VDD.n190 VSS 0.0182f
C1469 VDD.n191 VSS 0.00527f
C1470 VDD.n192 VSS 0.0262f
C1471 VDD.n193 VSS 0.0889f
C1472 VDD.n194 VSS 0.00482f
C1473 VDD.n195 VSS 0.00129f
C1474 VDD.n196 VSS 0.00443f
C1475 VDD.n197 VSS 0.0025f
C1476 VDD.n198 VSS 0.0025f
C1477 VDD.n199 VSS 0.104f
C1478 VDD.n200 VSS 0.0107f
C1479 VDD.n201 VSS 0.00385f
C1480 VDD.n202 VSS 0.015f
C1481 VDD.n203 VSS 0.11f
C1482 VDD.n204 VSS 0.00965f
C1483 VDD.n205 VSS 0.0154f
C1484 VDD.t317 VSS 0.0706f
C1485 VDD.n206 VSS 0.033f
C1486 VDD.n207 VSS 0.0107f
C1487 VDD.n208 VSS 0.00981f
C1488 VDD.n209 VSS 0.0075f
C1489 VDD.n210 VSS 0.00577f
C1490 VDD.n211 VSS 0.00258f
C1491 VDD.n212 VSS 0.00767f
C1492 VDD.n213 VSS 0.00825f
C1493 VDD.n214 VSS 0.0025f
C1494 VDD.n215 VSS 0.0025f
C1495 VDD.n216 VSS 0.00258f
C1496 VDD.n217 VSS 0.00742f
C1497 VDD.n218 VSS 0.00842f
C1498 VDD.n219 VSS 0.0025f
C1499 VDD.n220 VSS 0.0025f
C1500 VDD.n221 VSS 0.00517f
C1501 VDD.n222 VSS 0.00242f
C1502 VDD.n223 VSS 0.00653f
C1503 VDD.n224 VSS 0.0186f
C1504 VDD.n225 VSS 0.00909f
C1505 VDD.n226 VSS 0.00508f
C1506 VDD.n227 VSS 0.00909f
C1507 VDD.n228 VSS 0.0085f
C1508 VDD.n229 VSS 0.0503f
C1509 VDD.n230 VSS 0.0082f
C1510 VDD.n231 VSS 0.0082f
C1511 VDD.n232 VSS 0.00439f
C1512 VDD.n233 VSS 0.0071f
C1513 VDD.n234 VSS 0.00718f
C1514 VDD.t127 VSS 0.341f
C1515 VDD.t415 VSS 0.00681f
C1516 VDD.n235 VSS 0.00681f
C1517 VDD.n236 VSS 0.0147f
C1518 VDD.t179 VSS 0.0218f
C1519 VDD.n237 VSS 0.0796f
C1520 VDD.n238 VSS 0.0168f
C1521 VDD.n239 VSS 0.0435f
C1522 VDD.t133 VSS 0.00681f
C1523 VDD.n240 VSS 0.00681f
C1524 VDD.n241 VSS 0.0147f
C1525 VDD.t124 VSS 0.0218f
C1526 VDD.n242 VSS 0.0796f
C1527 VDD.n243 VSS 0.0168f
C1528 VDD.n244 VSS 0.0435f
C1529 VDD.n245 VSS 0.618f
C1530 VDD.n246 VSS 0.0918f
C1531 VDD.n247 VSS 0.333f
C1532 VDD.t132 VSS 0.345f
C1533 VDD.t53 VSS 0.345f
C1534 VDD.n248 VSS 0.333f
C1535 VDD.n249 VSS 0.0247f
C1536 VDD.n250 VSS 0.0389f
C1537 VDD.n251 VSS 0.0333f
C1538 VDD.t123 VSS 0.342f
C1539 VDD.n252 VSS 0.333f
C1540 VDD.n253 VSS 0.0395f
C1541 VDD.n254 VSS 0.629f
C1542 VDD.n255 VSS 0.0109f
C1543 VDD.n256 VSS 0.0174f
C1544 VDD.n257 VSS 0.0149f
C1545 VDD.n258 VSS 0.0149f
C1546 VDD.n259 VSS 0.0094f
C1547 VDD.n260 VSS 0.0147f
C1548 VDD.n261 VSS 0.0166f
C1549 VDD.n262 VSS 0.00351f
C1550 VDD.n263 VSS 0.00884f
C1551 VDD.n265 VSS 0.00237f
C1552 VDD.n266 VSS 0.00279f
C1553 VDD.n267 VSS 0.00369f
C1554 VDD.n268 VSS 0.0107f
C1555 VDD.n269 VSS 0.0121f
C1556 VDD.t401 VSS 0.00913f
C1557 VDD.t152 VSS 0.00808f
C1558 VDD.n270 VSS 0.0503f
C1559 VDD.t168 VSS 0.00405f
C1560 VDD.n271 VSS 0.00405f
C1561 VDD.n272 VSS 0.0099f
C1562 VDD.t405 VSS 0.00405f
C1563 VDD.n273 VSS 0.00405f
C1564 VDD.n274 VSS 0.0081f
C1565 VDD.n275 VSS 0.0254f
C1566 VDD.t49 VSS 0.00405f
C1567 VDD.n276 VSS 0.00405f
C1568 VDD.n277 VSS 0.0081f
C1569 VDD.t116 VSS 0.00405f
C1570 VDD.n278 VSS 0.00405f
C1571 VDD.n279 VSS 0.0099f
C1572 VDD.n280 VSS 0.0254f
C1573 VDD.n281 VSS 0.0319f
C1574 VDD.t50 VSS 0.11f
C1575 VDD.n282 VSS 0.125f
C1576 VDD.n283 VSS 0.0107f
C1577 VDD.t48 VSS 0.11f
C1578 VDD.n284 VSS 0.11f
C1579 VDD.n285 VSS 0.0107f
C1580 VDD.n286 VSS 0.00929f
C1581 VDD.n287 VSS 0.00808f
C1582 VDD.n288 VSS 0.0373f
C1583 VDD.n289 VSS 0.00808f
C1584 VDD.n290 VSS 0.00929f
C1585 VDD.n291 VSS 0.0373f
C1586 VDD.n292 VSS 0.064f
C1587 VDD.n293 VSS 0.0121f
C1588 VDD.n294 VSS 0.415f
C1589 VDD.n295 VSS 0.0121f
C1590 VDD.n296 VSS 0.0215f
C1591 VDD.t113 VSS 0.107f
C1592 VDD.n297 VSS 0.122f
C1593 VDD.n298 VSS 0.0107f
C1594 VDD.n299 VSS 0.0107f
C1595 VDD.n300 VSS 0.0366f
C1596 VDD.n301 VSS 0.0107f
C1597 VDD.n302 VSS 0.218f
C1598 VDD.n303 VSS 0.0107f
C1599 VDD.n304 VSS 0.0366f
C1600 VDD.n305 VSS 0.0366f
C1601 VDD.n306 VSS 0.0107f
C1602 VDD.n307 VSS 0.214f
C1603 VDD.n308 VSS 0.0107f
C1604 VDD.n309 VSS 0.0107f
C1605 VDD.n310 VSS 0.0107f
C1606 VDD.n311 VSS 0.0354f
C1607 VDD.n312 VSS 0.199f
C1608 VDD.n313 VSS 0.0107f
C1609 VDD.n314 VSS 0.0107f
C1610 VDD.n315 VSS 0.0369f
C1611 VDD.n316 VSS 0.0107f
C1612 VDD.t119 VSS 0.11f
C1613 VDD.n317 VSS 0.14f
C1614 VDD.n318 VSS 0.0107f
C1615 VDD.n319 VSS 0.0369f
C1616 VDD.n320 VSS 0.185f
C1617 VDD.n321 VSS 0.0107f
C1618 VDD.n322 VSS 0.0107f
C1619 VDD.n323 VSS 0.0319f
C1620 VDD.n324 VSS 0.0182f
C1621 VDD.n325 VSS 0.00931f
C1622 VDD.n326 VSS 0.248f
C1623 VDD.n327 VSS 0.00931f
C1624 VDD.n328 VSS 0.00522f
C1625 VDD.n329 VSS 0.00193f
C1626 VDD.n330 VSS 0.0128f
C1627 VDD.n331 VSS 0.0122f
C1628 VDD.n332 VSS 0.0283f
C1629 VDD.n333 VSS 0.0158f
C1630 VDD.n334 VSS 0.00764f
C1631 VDD.n335 VSS 0.012f
C1632 VDD.n336 VSS 0.012f
C1633 VDD.t120 VSS 0.0091f
C1634 VDD.t414 VSS 0.00812f
C1635 VDD.n337 VSS 0.0498f
C1636 VDD.n338 VSS 0.0379f
C1637 VDD.n339 VSS 0.019f
C1638 VDD.n340 VSS 0.0333f
C1639 VDD.n341 VSS 0.0147f
C1640 VDD.t151 VSS 0.00929f
C1641 VDD.t176 VSS 0.00808f
C1642 VDD.n342 VSS 0.0373f
C1643 VDD.n343 VSS 0.00913f
C1644 VDD.n344 VSS 0.00808f
C1645 VDD.n345 VSS 0.0509f
C1646 VDD.n346 VSS 0.122f
C1647 VDD.n347 VSS 0.131f
C1648 VDD.n348 VSS 0.0107f
C1649 VDD.n349 VSS 0.0185f
C1650 VDD.t156 VSS 0.0581f
C1651 VDD.n350 VSS 0.0701f
C1652 VDD.n351 VSS 0.0107f
C1653 VDD.n352 VSS 0.0185f
C1654 VDD.n353 VSS 0.0997f
C1655 VDD.n354 VSS 0.0107f
C1656 VDD.n355 VSS 0.0185f
C1657 VDD.t404 VSS 0.00405f
C1658 VDD.n356 VSS 0.00405f
C1659 VDD.n357 VSS 0.0099f
C1660 VDD.t162 VSS 0.00405f
C1661 VDD.n358 VSS 0.00405f
C1662 VDD.n359 VSS 0.0081f
C1663 VDD.n360 VSS 0.0254f
C1664 VDD.n361 VSS 0.0159f
C1665 VDD.n362 VSS 0.0177f
C1666 VDD.t161 VSS 0.0552f
C1667 VDD.n363 VSS 0.0627f
C1668 VDD.n364 VSS 0.0107f
C1669 VDD.n365 VSS 0.107f
C1670 VDD.n366 VSS 0.0107f
C1671 VDD.t163 VSS 0.0552f
C1672 VDD.n367 VSS 0.0552f
C1673 VDD.n368 VSS 0.0107f
C1674 VDD.n369 VSS 0.0183f
C1675 VDD.n370 VSS 0.109f
C1676 VDD.n371 VSS 0.0107f
C1677 VDD.n372 VSS 0.0183f
C1678 VDD.t150 VSS 0.0467f
C1679 VDD.n373 VSS 0.0609f
C1680 VDD.n374 VSS 0.01f
C1681 VDD.n375 VSS 0.0172f
C1682 VDD.n376 VSS 0.00901f
C1683 VDD.n377 VSS 0.0545f
C1684 VDD.n378 VSS 0.00527f
C1685 VDD.n379 VSS 0.147f
C1686 VDD.n380 VSS 0.00129f
C1687 VDD.n381 VSS 0.0022f
C1688 VDD.n382 VSS 0.0204f
C1689 VDD.n383 VSS 0.00861f
C1690 VDD.n384 VSS 0.0022f
C1691 VDD.n385 VSS 0.0543f
C1692 VDD.n386 VSS 0.00696f
C1693 VDD.n387 VSS 0.0025f
C1694 VDD.n388 VSS 0.0025f
C1695 VDD.n389 VSS 0.0144f
C1696 VDD.n390 VSS 0.0485f
C1697 VDD.n391 VSS 0.149f
C1698 VDD.n392 VSS 0.201f
C1699 VDD.n393 VSS 0.0102f
C1700 VDD.n394 VSS 0.0752f
C1701 VDD.n395 VSS 0.00998f
C1702 VDD.n396 VSS 0.00908f
C1703 VDD.n397 VSS 0.00486f
C1704 VDD.n398 VSS 0.00786f
C1705 VDD.n399 VSS 0.00884f
C1706 VDD.n400 VSS 0.0636f
C1707 VDD.n401 VSS 0.213f
C1708 VDD.n402 VSS 0.0101f
C1709 VDD.n403 VSS 0.00723f
C1710 VDD.n404 VSS 0.00509f
C1711 VDD.n405 VSS 0.109f
C1712 VDD.n406 VSS 0.00453f
C1713 VDD.n407 VSS 0.0115f
C1714 VDD.n408 VSS 0.0241f
C1715 VDD.n409 VSS 0.0025f
C1716 VDD.n410 VSS 0.769f
C1717 VDD.n411 VSS 1.23f
C1718 VDD.n412 VSS 0.24f
C1719 VDD.t204 VSS 0.0311f
C1720 VDD.t206 VSS 0.0177f
C1721 VDD.n413 VSS 0.0826f
C1722 VDD.t242 VSS 0.0311f
C1723 VDD.t243 VSS 0.0177f
C1724 VDD.n414 VSS 0.0826f
C1725 VDD.t230 VSS 0.0311f
C1726 VDD.t231 VSS 0.0177f
C1727 VDD.n415 VSS 0.0825f
C1728 VDD.t232 VSS 0.0311f
C1729 VDD.t234 VSS 0.0177f
C1730 VDD.n416 VSS 0.0824f
C1731 VDD.n417 VSS 0.289f
C1732 VDD.t1 VSS 0.00405f
C1733 VDD.n418 VSS 0.00405f
C1734 VDD.n419 VSS 0.0081f
C1735 VDD.n420 VSS 0.0156f
C1736 VDD.t287 VSS 0.00405f
C1737 VDD.n421 VSS 0.00405f
C1738 VDD.n422 VSS 0.0081f
C1739 VDD.n423 VSS 0.0372f
C1740 VDD.n424 VSS 0.0155f
C1741 VDD.t34 VSS 0.00405f
C1742 VDD.n425 VSS 0.00405f
C1743 VDD.n426 VSS 0.0081f
C1744 VDD.n427 VSS 0.0342f
C1745 VDD.n428 VSS 0.0178f
C1746 VDD.t218 VSS 0.017f
C1747 VDD.n429 VSS 0.0143f
C1748 VDD.t216 VSS 0.0323f
C1749 VDD.n430 VSS 0.0611f
C1750 VDD.n431 VSS 0.0196f
C1751 VDD.t224 VSS 0.0329f
C1752 VDD.t226 VSS 0.0172f
C1753 VDD.n432 VSS 0.0826f
C1754 VDD.n434 VSS 0.0165f
C1755 VDD.n435 VSS 0.0155f
C1756 VDD.n437 VSS 0.0171f
C1757 VDD.n438 VSS 0.0162f
C1758 VDD.n440 VSS 0.0401f
C1759 VDD.n441 VSS 0.0165f
C1760 VDD.n442 VSS 0.00808f
C1761 VDD.n443 VSS 0.00913f
C1762 VDD.n444 VSS 0.0509f
C1763 VDD.n445 VSS 0.118f
C1764 VDD.t276 VSS 0.00405f
C1765 VDD.n446 VSS 0.00405f
C1766 VDD.n447 VSS 0.0081f
C1767 VDD.t263 VSS 0.00405f
C1768 VDD.n448 VSS 0.00405f
C1769 VDD.n449 VSS 0.0099f
C1770 VDD.n450 VSS 0.0254f
C1771 VDD.n451 VSS 0.0159f
C1772 VDD.t254 VSS 0.0552f
C1773 VDD.n452 VSS 0.0552f
C1774 VDD.n453 VSS 0.0107f
C1775 VDD.n454 VSS 0.214f
C1776 VDD.t282 VSS 0.00808f
C1777 VDD.t269 VSS 0.00929f
C1778 VDD.n455 VSS 0.0373f
C1779 VDD.n456 VSS 0.00808f
C1780 VDD.n457 VSS 0.00913f
C1781 VDD.n458 VSS 0.0503f
C1782 VDD.n459 VSS 0.0997f
C1783 VDD.n460 VSS 0.0107f
C1784 VDD.n461 VSS 6.19e-20
C1785 VDD.n462 VSS 0.00929f
C1786 VDD.n463 VSS 0.00808f
C1787 VDD.n464 VSS 0.0373f
C1788 VDD.n465 VSS 0.00808f
C1789 VDD.n466 VSS 0.00929f
C1790 VDD.n467 VSS 0.0373f
C1791 VDD.t338 VSS 0.00405f
C1792 VDD.n468 VSS 0.00405f
C1793 VDD.n469 VSS 0.0081f
C1794 VDD.t143 VSS 0.00405f
C1795 VDD.n470 VSS 0.00405f
C1796 VDD.n471 VSS 0.0099f
C1797 VDD.n472 VSS 0.0254f
C1798 VDD.n473 VSS 0.0159f
C1799 VDD.t374 VSS 0.00808f
C1800 VDD.t359 VSS 0.00913f
C1801 VDD.n474 VSS 0.0509f
C1802 VDD.n475 VSS 0.122f
C1803 VDD.n476 VSS 0.131f
C1804 VDD.n477 VSS 0.0107f
C1805 VDD.n478 VSS 0.0185f
C1806 VDD.t358 VSS 0.0581f
C1807 VDD.n479 VSS 0.0701f
C1808 VDD.n480 VSS 0.0107f
C1809 VDD.n481 VSS 0.0185f
C1810 VDD.n482 VSS 0.0997f
C1811 VDD.n483 VSS 0.0107f
C1812 VDD.n484 VSS 0.0185f
C1813 VDD.n485 VSS 0.0177f
C1814 VDD.t355 VSS 0.0552f
C1815 VDD.n486 VSS 0.0627f
C1816 VDD.n487 VSS 0.0107f
C1817 VDD.n488 VSS 0.107f
C1818 VDD.n489 VSS 0.0107f
C1819 VDD.t142 VSS 0.0552f
C1820 VDD.n490 VSS 0.0552f
C1821 VDD.n491 VSS 0.0107f
C1822 VDD.n492 VSS 0.0183f
C1823 VDD.n493 VSS 0.109f
C1824 VDD.n494 VSS 0.0107f
C1825 VDD.n495 VSS 0.0183f
C1826 VDD.t139 VSS 0.0591f
C1827 VDD.n496 VSS 0.0609f
C1828 VDD.n497 VSS 0.0107f
C1829 VDD.n498 VSS 0.0183f
C1830 VDD.n499 VSS 0.214f
C1831 VDD.n500 VSS 0.0107f
C1832 VDD.n501 VSS 0.289f
C1833 VDD.n502 VSS 0.289f
C1834 VDD.n503 VSS 0.214f
C1835 VDD.n504 VSS 0.0107f
C1836 VDD.t311 VSS 0.0591f
C1837 VDD.n505 VSS 0.0609f
C1838 VDD.n506 VSS 0.0107f
C1839 VDD.n507 VSS 0.0183f
C1840 VDD.n508 VSS 0.109f
C1841 VDD.n509 VSS 0.0107f
C1842 VDD.n510 VSS 0.0183f
C1843 VDD.n511 VSS 0.0111f
C1844 VDD.t106 VSS 0.00405f
C1845 VDD.n512 VSS 0.00405f
C1846 VDD.n513 VSS 0.0099f
C1847 VDD.t65 VSS 0.00405f
C1848 VDD.n514 VSS 0.00405f
C1849 VDD.n515 VSS 0.0081f
C1850 VDD.n516 VSS 0.0324f
C1851 VDD.t212 VSS 0.0172f
C1852 VDD.t210 VSS 0.0329f
C1853 VDD.n517 VSS 0.0826f
C1854 VDD.t227 VSS 0.0322f
C1855 VDD.n518 VSS 0.0613f
C1856 VDD.t229 VSS 0.017f
C1857 VDD.n519 VSS 0.0142f
C1858 VDD.n520 VSS 0.0195f
C1859 VDD.n521 VSS 0.0342f
C1860 VDD.t351 VSS 0.00405f
C1861 VDD.n522 VSS 0.00405f
C1862 VDD.n523 VSS 0.0081f
C1863 VDD.n524 VSS 0.02f
C1864 VDD.t144 VSS 0.00405f
C1865 VDD.n525 VSS 0.00405f
C1866 VDD.n526 VSS 0.0081f
C1867 VDD.n527 VSS 0.0206f
C1868 VDD.n528 VSS 0.0342f
C1869 VDD.t107 VSS 0.00405f
C1870 VDD.n529 VSS 0.00405f
C1871 VDD.n530 VSS 0.0081f
C1872 VDD.n531 VSS 0.0178f
C1873 VDD.n532 VSS 0.0378f
C1874 VDD.n533 VSS 0.0268f
C1875 VDD.t112 VSS 0.00405f
C1876 VDD.n534 VSS 0.00405f
C1877 VDD.n535 VSS 0.0081f
C1878 VDD.n536 VSS 0.02f
C1879 VDD.t339 VSS 0.00405f
C1880 VDD.n537 VSS 0.00405f
C1881 VDD.n538 VSS 0.0081f
C1882 VDD.n539 VSS 0.0206f
C1883 VDD.n540 VSS 0.0277f
C1884 VDD.n541 VSS 0.0372f
C1885 VDD.t149 VSS 0.00405f
C1886 VDD.n542 VSS 0.00405f
C1887 VDD.n543 VSS 0.0081f
C1888 VDD.n544 VSS 0.0155f
C1889 VDD.t350 VSS 0.00405f
C1890 VDD.n545 VSS 0.00405f
C1891 VDD.n546 VSS 0.0081f
C1892 VDD.n547 VSS 0.0141f
C1893 VDD.n548 VSS 0.0275f
C1894 VDD.n549 VSS 0.0386f
C1895 VDD.t67 VSS 0.00405f
C1896 VDD.n550 VSS 0.00405f
C1897 VDD.n551 VSS 0.0081f
C1898 VDD.n552 VSS 0.0198f
C1899 VDD.t297 VSS 0.00405f
C1900 VDD.n553 VSS 0.00405f
C1901 VDD.n554 VSS 0.0081f
C1902 VDD.n555 VSS 0.0207f
C1903 VDD.n556 VSS 0.0388f
C1904 VDD.n557 VSS 0.0266f
C1905 VDD.t375 VSS 0.00405f
C1906 VDD.n558 VSS 0.00405f
C1907 VDD.n559 VSS 0.0081f
C1908 VDD.n560 VSS 0.0156f
C1909 VDD.t298 VSS 0.00405f
C1910 VDD.n561 VSS 0.00405f
C1911 VDD.n562 VSS 0.0081f
C1912 VDD.n563 VSS 0.0132f
C1913 VDD.n564 VSS 0.0342f
C1914 VDD.t146 VSS 0.00405f
C1915 VDD.n565 VSS 0.00405f
C1916 VDD.n566 VSS 0.0081f
C1917 VDD.n567 VSS 0.0224f
C1918 VDD.t352 VSS 0.00405f
C1919 VDD.n568 VSS 0.00405f
C1920 VDD.n569 VSS 0.0081f
C1921 VDD.n570 VSS 0.0228f
C1922 VDD.n571 VSS 0.0342f
C1923 VDD.t314 VSS 0.00405f
C1924 VDD.n572 VSS 0.00405f
C1925 VDD.n573 VSS 0.0081f
C1926 VDD.n574 VSS 0.0156f
C1927 VDD.n575 VSS 0.0337f
C1928 VDD.t197 VSS 0.0177f
C1929 VDD.t195 VSS 0.0311f
C1930 VDD.n576 VSS 0.0825f
C1931 VDD.t223 VSS 0.0177f
C1932 VDD.t222 VSS 0.0311f
C1933 VDD.n577 VSS 0.0825f
C1934 VDD.t209 VSS 0.0177f
C1935 VDD.t207 VSS 0.0311f
C1936 VDD.n578 VSS 0.0826f
C1937 VDD.t239 VSS 0.0177f
C1938 VDD.t238 VSS 0.0311f
C1939 VDD.n579 VSS 0.0826f
C1940 VDD.n580 VSS 0.0688f
C1941 VDD.n581 VSS 0.0376f
C1942 VDD.n582 VSS 0.0304f
C1943 VDD.n583 VSS 0.0724f
C1944 VDD.n584 VSS 0.0198f
C1945 VDD.n585 VSS 0.0153f
C1946 VDD.n586 VSS 0.0208f
C1947 VDD.n587 VSS 0.0718f
C1948 VDD.n588 VSS 0.0198f
C1949 VDD.n589 VSS 0.00782f
C1950 VDD.n590 VSS 0.0443f
C1951 VDD.n591 VSS 0.0198f
C1952 VDD.n592 VSS 0.0154f
C1953 VDD.n593 VSS 0.0633f
C1954 VDD.n594 VSS 0.0198f
C1955 VDD.n595 VSS 0.0154f
C1956 VDD.n596 VSS 0.0718f
C1957 VDD.n597 VSS 0.0198f
C1958 VDD.n598 VSS 0.011f
C1959 VDD.n599 VSS 0.0208f
C1960 VDD.n600 VSS 0.0603f
C1961 VDD.n601 VSS 0.0198f
C1962 VDD.n602 VSS 0.0121f
C1963 VDD.n603 VSS 0.047f
C1964 VDD.n604 VSS 0.0198f
C1965 VDD.n605 VSS 0.0154f
C1966 VDD.t208 VSS 0.205f
C1967 VDD.t196 VSS 0.0621f
C1968 VDD.n606 VSS 0.0382f
C1969 VDD.n607 VSS 0.0471f
C1970 VDD.n608 VSS 0.0362f
C1971 VDD.n609 VSS 0.0198f
C1972 VDD.n610 VSS 0.015f
C1973 VDD.n611 VSS 0.0208f
C1974 VDD.n612 VSS 0.0718f
C1975 VDD.n613 VSS 0.0198f
C1976 VDD.n614 VSS 0.00808f
C1977 VDD.n615 VSS 0.041f
C1978 VDD.n616 VSS 0.0198f
C1979 VDD.n617 VSS 0.0154f
C1980 VDD.n618 VSS 0.0666f
C1981 VDD.n619 VSS 0.0198f
C1982 VDD.n620 VSS 0.0154f
C1983 VDD.n621 VSS 0.0718f
C1984 VDD.n622 VSS 0.0198f
C1985 VDD.n623 VSS 0.0103f
C1986 VDD.n624 VSS 0.0209f
C1987 VDD.n625 VSS 0.057f
C1988 VDD.n626 VSS 0.0198f
C1989 VDD.n627 VSS 0.0127f
C1990 VDD.n628 VSS 0.0507f
C1991 VDD.n629 VSS 0.0198f
C1992 VDD.n630 VSS 0.0154f
C1993 VDD.n631 VSS 0.088f
C1994 VDD.n632 VSS 0.0243f
C1995 VDD.n633 VSS 0.016f
C1996 VDD.n634 VSS 0.0307f
C1997 VDD.n635 VSS 0.165f
C1998 VDD.n637 VSS 0.0219f
C1999 VDD.n638 VSS 0.0243f
C2000 VDD.n639 VSS 0.131f
C2001 VDD.n640 VSS 0.0211f
C2002 VDD.n641 VSS 0.0205f
C2003 VDD.n642 VSS 0.262f
C2004 VDD.n643 VSS 0.0194f
C2005 VDD.n644 VSS 0.0187f
C2006 VDD.n645 VSS 0.223f
C2007 VDD.n646 VSS 0.0171f
C2008 VDD.n647 VSS 0.0165f
C2009 VDD.n648 VSS 0.223f
C2010 VDD.n649 VSS 0.0171f
C2011 VDD.n650 VSS 0.0165f
C2012 VDD.t103 VSS 0.206f
C2013 VDD.n651 VSS 0.0281f
C2014 VDD.n652 VSS 0.0171f
C2015 VDD.n653 VSS 0.0165f
C2016 VDD.n654 VSS 0.223f
C2017 VDD.n655 VSS 0.0171f
C2018 VDD.n656 VSS 0.00901f
C2019 VDD.n657 VSS 0.0189f
C2020 VDD.n658 VSS 0.223f
C2021 VDD.n659 VSS 0.0171f
C2022 VDD.n660 VSS 0.0157f
C2023 VDD.n661 VSS 0.187f
C2024 VDD.n662 VSS 0.0171f
C2025 VDD.n663 VSS 0.0165f
C2026 VDD.n664 VSS 0.223f
C2027 VDD.n665 VSS 0.0171f
C2028 VDD.n666 VSS 0.0165f
C2029 VDD.t68 VSS 0.206f
C2030 VDD.n667 VSS 0.124f
C2031 VDD.n668 VSS 0.0171f
C2032 VDD.n669 VSS 0.0137f
C2033 VDD.n670 VSS 0.0189f
C2034 VDD.n671 VSS 0.223f
C2035 VDD.n672 VSS 0.0171f
C2036 VDD.n673 VSS 0.011f
C2037 VDD.t66 VSS 0.206f
C2038 VDD.n674 VSS 0.0599f
C2039 VDD.n675 VSS 0.0171f
C2040 VDD.n676 VSS 0.0165f
C2041 VDD.n677 VSS 0.223f
C2042 VDD.n678 VSS 0.0171f
C2043 VDD.n679 VSS 0.0165f
C2044 VDD.n680 VSS 0.223f
C2045 VDD.n681 VSS 0.0171f
C2046 VDD.n682 VSS 0.0165f
C2047 VDD.n683 VSS 0.223f
C2048 VDD.n684 VSS 0.0171f
C2049 VDD.n685 VSS 0.0165f
C2050 VDD.n686 VSS 0.223f
C2051 VDD.n687 VSS 0.0171f
C2052 VDD.n688 VSS 0.0165f
C2053 VDD.n689 VSS 0.208f
C2054 VDD.n690 VSS 0.0171f
C2055 VDD.n691 VSS 0.0106f
C2056 VDD.n692 VSS 0.0189f
C2057 VDD.n693 VSS 0.223f
C2058 VDD.n694 VSS 0.0171f
C2059 VDD.n695 VSS 0.0141f
C2060 VDD.n696 VSS 0.144f
C2061 VDD.n697 VSS 0.0171f
C2062 VDD.n698 VSS 0.0165f
C2063 VDD.n699 VSS 0.223f
C2064 VDD.n700 VSS 0.0171f
C2065 VDD.n701 VSS 0.0165f
C2066 VDD.t108 VSS 0.206f
C2067 VDD.n702 VSS 0.0805f
C2068 VDD.n703 VSS 0.0171f
C2069 VDD.n704 VSS 0.0153f
C2070 VDD.n705 VSS 0.0189f
C2071 VDD.n706 VSS 0.223f
C2072 VDD.n707 VSS 0.0171f
C2073 VDD.n708 VSS 0.00943f
C2074 VDD.t71 VSS 0.223f
C2075 VDD.n709 VSS 0.0171f
C2076 VDD.n710 VSS 0.0165f
C2077 VDD.n711 VSS 0.223f
C2078 VDD.n712 VSS 0.0171f
C2079 VDD.n713 VSS 0.0165f
C2080 VDD.n714 VSS 0.223f
C2081 VDD.n715 VSS 0.0171f
C2082 VDD.n716 VSS 0.0165f
C2083 VDD.n717 VSS 0.223f
C2084 VDD.n718 VSS 0.0182f
C2085 VDD.n719 VSS 0.0176f
C2086 VDD.t236 VSS 0.0917f
C2087 VDD.t187 VSS 0.00749f
C2088 VDD.t190 VSS 0.0487f
C2089 VDD.n720 VSS 0.281f
C2090 VDD.n721 VSS 0.0219f
C2091 VDD.n722 VSS 0.0211f
C2092 VDD.n723 VSS 0.316f
C2093 VDD.n724 VSS 0.0228f
C2094 VDD.n725 VSS 0.022f
C2095 VDD.t191 VSS 0.0177f
C2096 VDD.t189 VSS 0.0338f
C2097 VDD.n726 VSS 0.0796f
C2098 VDD.n727 VSS 0.0103f
C2099 VDD.n728 VSS 0.00808f
C2100 VDD.n729 VSS 0.0481f
C2101 VDD.t188 VSS 0.0177f
C2102 VDD.t186 VSS 0.0574f
C2103 VDD.n730 VSS 0.0798f
C2104 VDD.t336 VSS 0.00405f
C2105 VDD.n731 VSS 0.00405f
C2106 VDD.n732 VSS 0.0116f
C2107 VDD.t400 VSS 0.00405f
C2108 VDD.n733 VSS 0.00405f
C2109 VDD.n734 VSS 0.0081f
C2110 VDD.n735 VSS 0.0356f
C2111 VDD.t237 VSS 0.0177f
C2112 VDD.t235 VSS 0.0338f
C2113 VDD.n736 VSS 0.0796f
C2114 VDD.t370 VSS 0.00405f
C2115 VDD.n737 VSS 0.00405f
C2116 VDD.n738 VSS 0.0116f
C2117 VDD.t393 VSS 0.00405f
C2118 VDD.n739 VSS 0.00405f
C2119 VDD.n740 VSS 0.0081f
C2120 VDD.n741 VSS 0.0356f
C2121 VDD.t248 VSS 0.0177f
C2122 VDD.t247 VSS 0.0338f
C2123 VDD.n742 VSS 0.0805f
C2124 VDD.n743 VSS 0.0214f
C2125 VDD.n745 VSS 0.0176f
C2126 VDD.n746 VSS 0.00785f
C2127 VDD.n747 VSS 0.0184f
C2128 VDD.n748 VSS 0.0191f
C2129 VDD.n749 VSS 0.0106f
C2130 VDD.n750 VSS 0.0191f
C2131 VDD.n751 VSS 0.0171f
C2132 VDD.n752 VSS 0.0192f
C2133 VDD.n753 VSS 0.00877f
C2134 VDD.n754 VSS 0.0229f
C2135 VDD.n756 VSS 0.0191f
C2136 VDD.n757 VSS 0.0162f
C2137 VDD.n758 VSS 0.0183f
C2138 VDD.n759 VSS 0.0175f
C2139 VDD.n760 VSS 0.00779f
C2140 VDD.n762 VSS 0.016f
C2141 VDD.n763 VSS 0.00962f
C2142 VDD.n764 VSS 0.0215f
C2143 VDD.n765 VSS 0.0191f
C2144 VDD.n766 VSS 0.0146f
C2145 VDD.n768 VSS 0.0223f
C2146 VDD.n769 VSS 0.0113f
C2147 VDD.n770 VSS 0.0198f
C2148 VDD.n771 VSS 0.024f
C2149 VDD.n772 VSS 0.0112f
C2150 VDD.n773 VSS 0.0256f
C2151 VDD.n775 VSS 0.0223f
C2152 VDD.n776 VSS 0.0174f
C2153 VDD.n777 VSS 0.0175f
C2154 VDD.n778 VSS 0.0156f
C2155 VDD.n780 VSS 0.316f
C2156 VDD.n782 VSS 0.0513f
C2157 VDD.n783 VSS 0.0115f
C2158 VDD.n784 VSS 0.0103f
C2159 VDD.n785 VSS 0.0505f
C2160 VDD.n786 VSS 0.0932f
C2161 VDD.n787 VSS 0.0347f
C2162 VDD.n788 VSS 0.0119f
C2163 VDD.n789 VSS 0.0239f
C2164 VDD.n790 VSS 0.0165f
C2165 VDD.n791 VSS 0.00987f
C2166 VDD.n792 VSS 0.0137f
C2167 VDD.n793 VSS 0.0225f
C2168 VDD.n794 VSS 0.0165f
C2169 VDD.n795 VSS 0.00898f
C2170 VDD.n796 VSS 0.0139f
C2171 VDD.n797 VSS 0.0132f
C2172 VDD.n798 VSS 0.0165f
C2173 VDD.n799 VSS 0.0165f
C2174 VDD.n800 VSS 0.0237f
C2175 VDD.n801 VSS 0.0165f
C2176 VDD.n802 VSS 0.0164f
C2177 VDD.n803 VSS 0.0218f
C2178 VDD.n804 VSS 0.0238f
C2179 VDD.n805 VSS 0.0165f
C2180 VDD.n806 VSS 0.0083f
C2181 VDD.n807 VSS 0.0238f
C2182 VDD.n808 VSS 0.0165f
C2183 VDD.n809 VSS 0.0165f
C2184 VDD.n810 VSS 0.073f
C2185 VDD.n811 VSS 0.0438f
C2186 VDD.n813 VSS 0.0401f
C2187 VDD.n814 VSS 0.0378f
C2188 VDD.n815 VSS 0.0171f
C2189 VDD.n816 VSS 0.0125f
C2190 VDD.t246 VSS 0.0172f
C2191 VDD.t244 VSS 0.0329f
C2192 VDD.n817 VSS 0.0839f
C2193 VDD.t215 VSS 0.0172f
C2194 VDD.t213 VSS 0.032f
C2195 VDD.n818 VSS 0.0834f
C2196 VDD.n819 VSS 0.0169f
C2197 VDD.n820 VSS 0.588f
C2198 VDD.n821 VSS 0.00696f
C2199 VDD.n822 VSS 0.016f
C2200 VDD.n823 VSS 0.0129f
C2201 VDD.n825 VSS 0.0152f
C2202 VDD.n826 VSS 0.0137f
C2203 VDD.t72 VSS 0.00405f
C2204 VDD.n827 VSS 0.00405f
C2205 VDD.n828 VSS 0.0081f
C2206 VDD.n829 VSS 0.0166f
C2207 VDD.n830 VSS 0.0351f
C2208 VDD.t380 VSS 0.00405f
C2209 VDD.n831 VSS 0.00405f
C2210 VDD.n832 VSS 0.0081f
C2211 VDD.n833 VSS 0.0136f
C2212 VDD.n834 VSS 0.0605f
C2213 VDD.n835 VSS 0.152f
C2214 VDD.n836 VSS 0.0312f
C2215 VDD.n837 VSS 0.283f
C2216 VDD.n838 VSS 0.0221f
C2217 VDD.n839 VSS 0.0278f
C2218 VDD.n840 VSS 0.223f
C2219 VDD.n841 VSS 0.0192f
C2220 VDD.n842 VSS 0.0254f
C2221 VDD.n843 VSS 0.223f
C2222 VDD.n844 VSS 0.0176f
C2223 VDD.n845 VSS 0.0234f
C2224 VDD.n846 VSS 0.211f
C2225 VDD.n847 VSS 0.0176f
C2226 VDD.n848 VSS 0.0234f
C2227 VDD.n849 VSS 0.223f
C2228 VDD.n850 VSS 0.0176f
C2229 VDD.n851 VSS 0.0234f
C2230 VDD.n852 VSS 0.223f
C2231 VDD.n853 VSS 0.0176f
C2232 VDD.n854 VSS 0.0119f
C2233 VDD.n855 VSS 0.0182f
C2234 VDD.t145 VSS 0.206f
C2235 VDD.n856 VSS 0.0524f
C2236 VDD.n857 VSS 0.0176f
C2237 VDD.n858 VSS 0.0232f
C2238 VDD.n859 VSS 0.223f
C2239 VDD.n860 VSS 0.0176f
C2240 VDD.n861 VSS 0.0234f
C2241 VDD.n862 VSS 0.116f
C2242 VDD.n863 VSS 0.0176f
C2243 VDD.n864 VSS 0.0234f
C2244 VDD.n865 VSS 0.223f
C2245 VDD.n866 VSS 0.0176f
C2246 VDD.n867 VSS 0.0185f
C2247 VDD.n868 VSS 0.0347f
C2248 VDD.n869 VSS 0.0625f
C2249 VDD.n870 VSS 0.0192f
C2250 VDD.n871 VSS 0.18f
C2251 VDD.n872 VSS 0.0176f
C2252 VDD.n873 VSS 0.0166f
C2253 VDD.n874 VSS 0.223f
C2254 VDD.n875 VSS 0.0176f
C2255 VDD.n876 VSS 0.0234f
C2256 VDD.n877 VSS 0.223f
C2257 VDD.n878 VSS 0.0176f
C2258 VDD.n879 VSS 0.0168f
C2259 VDD.n880 VSS 0.223f
C2260 VDD.n881 VSS 0.0176f
C2261 VDD.n882 VSS 0.0183f
C2262 VDD.n883 VSS 0.223f
C2263 VDD.n884 VSS 0.0176f
C2264 VDD.n885 VSS 0.0234f
C2265 VDD.t136 VSS 0.206f
C2266 VDD.n886 VSS 0.0318f
C2267 VDD.n887 VSS 0.0176f
C2268 VDD.n888 VSS 0.0234f
C2269 VDD.n889 VSS 0.223f
C2270 VDD.n890 VSS 0.0176f
C2271 VDD.n891 VSS 0.0141f
C2272 VDD.n892 VSS 0.0182f
C2273 VDD.t111 VSS 0.206f
C2274 VDD.n893 VSS 0.0954f
C2275 VDD.n894 VSS 0.0176f
C2276 VDD.n895 VSS 0.0209f
C2277 VDD.n896 VSS 0.223f
C2278 VDD.n897 VSS 0.0176f
C2279 VDD.n898 VSS 0.0234f
C2280 VDD.n899 VSS 0.159f
C2281 VDD.n900 VSS 0.0176f
C2282 VDD.n901 VSS 0.0234f
C2283 VDD.n902 VSS 0.223f
C2284 VDD.n903 VSS 0.0176f
C2285 VDD.n904 VSS 0.0207f
C2286 VDD.n905 VSS 0.0192f
C2287 VDD.n906 VSS 0.223f
C2288 VDD.n907 VSS 0.0176f
C2289 VDD.n908 VSS 0.0143f
C2290 VDD.n909 VSS 0.223f
C2291 VDD.n910 VSS 0.0176f
C2292 VDD.n911 VSS 0.0234f
C2293 VDD.n912 VSS 0.223f
C2294 VDD.n913 VSS 0.0176f
C2295 VDD.n914 VSS 0.0234f
C2296 VDD.n915 VSS 0.223f
C2297 VDD.n916 VSS 0.0176f
C2298 VDD.n917 VSS 0.0234f
C2299 VDD.n918 VSS 0.253f
C2300 VDD.n919 VSS 0.0237f
C2301 VDD.n920 VSS 0.0323f
C2302 VDD.n921 VSS 0.266f
C2303 VDD.n922 VSS 0.0274f
C2304 VDD.n923 VSS 0.0279f
C2305 VDD.n924 VSS 0.0196f
C2306 VDD.n925 VSS 0.283f
C2307 VDD.n926 VSS 0.0182f
C2308 VDD.n927 VSS 0.017f
C2309 VDD.n928 VSS 0.0183f
C2310 VDD.n929 VSS 0.0223f
C2311 VDD.n930 VSS 0.0204f
C2312 VDD.n931 VSS 0.0193f
C2313 VDD.n932 VSS 0.0859f
C2314 VDD.n933 VSS 0.0257f
C2315 VDD.n934 VSS 0.0241f
C2316 VDD.n935 VSS 0.0598f
C2317 VDD.n936 VSS 0.0226f
C2318 VDD.n937 VSS 0.0208f
C2319 VDD.n938 VSS 0.674f
C2320 VDD.t228 VSS 0.417f
C2321 VDD.t325 VSS 0.00374f
C2322 VDD.t214 VSS 0.259f
C2323 VDD.n939 VSS 0.0381f
C2324 VDD.n940 VSS 0.0165f
C2325 VDD.n941 VSS 0.0131f
C2326 VDD.n942 VSS 0.0223f
C2327 VDD.n943 VSS 0.0605f
C2328 VDD.n944 VSS 0.0165f
C2329 VDD.n945 VSS 0.00966f
C2330 VDD.n946 VSS 0.0322f
C2331 VDD.n947 VSS 0.029f
C2332 VDD.n948 VSS 0.0165f
C2333 VDD.n949 VSS 0.0151f
C2334 VDD.t211 VSS 0.726f
C2335 VDD.t245 VSS 0.486f
C2336 VDD.n951 VSS 0.0384f
C2337 VDD.n952 VSS 0.0165f
C2338 VDD.n953 VSS 0.0124f
C2339 VDD.n954 VSS 0.021f
C2340 VDD.n955 VSS 0.0645f
C2341 VDD.n956 VSS 0.0165f
C2342 VDD.n957 VSS 0.0103f
C2343 VDD.n958 VSS 0.0641f
C2344 VDD.n959 VSS 0.0165f
C2345 VDD.n960 VSS 0.0129f
C2346 VDD.n961 VSS 0.122f
C2347 VDD.n962 VSS 0.045f
C2348 VDD.n964 VSS 0.0428f
C2349 VDD.n965 VSS 0.0426f
C2350 VDD.n966 VSS 0.0163f
C2351 VDD.n967 VSS 0.0153f
C2352 VDD.n969 VSS 0.0163f
C2353 VDD.n970 VSS 0.0153f
C2354 VDD.n972 VSS 0.0165f
C2355 VDD.n973 VSS 0.0155f
C2356 VDD.n975 VSS 0.0165f
C2357 VDD.n976 VSS 0.0155f
C2358 VDD.n978 VSS 0.0165f
C2359 VDD.n979 VSS 0.0155f
C2360 VDD.n981 VSS 0.0165f
C2361 VDD.n982 VSS 0.0155f
C2362 VDD.n984 VSS 0.0165f
C2363 VDD.n985 VSS 0.0155f
C2364 VDD.n987 VSS 0.0165f
C2365 VDD.n988 VSS 0.0155f
C2366 VDD.n990 VSS 0.0165f
C2367 VDD.n991 VSS 0.0155f
C2368 VDD.n993 VSS 0.0165f
C2369 VDD.n994 VSS 0.0155f
C2370 VDD.n996 VSS 0.0165f
C2371 VDD.n997 VSS 0.0128f
C2372 VDD.n998 VSS 1f
C2373 VDD.n1000 VSS 0.0165f
C2374 VDD.n1001 VSS 0.128f
C2375 VDD.t296 VSS 0.00923f
C2376 VDD.t102 VSS 0.00808f
C2377 VDD.n1002 VSS 0.0383f
C2378 VDD.n1003 VSS 0.134f
C2379 VDD.t101 VSS 0.0605f
C2380 VDD.n1004 VSS 0.0701f
C2381 VDD.n1005 VSS 0.0108f
C2382 VDD.n1006 VSS 0.148f
C2383 VDD.n1007 VSS 0.144f
C2384 VDD.n1008 VSS 0.0997f
C2385 VDD.n1009 VSS 0.0107f
C2386 VDD.n1010 VSS 0.0161f
C2387 VDD.n1011 VSS 0.0183f
C2388 VDD.t64 VSS 0.0552f
C2389 VDD.n1012 VSS 0.0552f
C2390 VDD.n1013 VSS 0.0107f
C2391 VDD.t73 VSS 0.0552f
C2392 VDD.n1014 VSS 0.0627f
C2393 VDD.n1015 VSS 0.0107f
C2394 VDD.n1016 VSS 0.107f
C2395 VDD.n1017 VSS 0.0107f
C2396 VDD.n1018 VSS 0.115f
C2397 VDD.t302 VSS 0.00405f
C2398 VDD.n1019 VSS 0.00405f
C2399 VDD.n1020 VSS 0.0081f
C2400 VDD.t295 VSS 0.00405f
C2401 VDD.n1021 VSS 0.00405f
C2402 VDD.n1022 VSS 0.0099f
C2403 VDD.n1023 VSS 0.0273f
C2404 VDD.t294 VSS 0.0552f
C2405 VDD.n1024 VSS 0.0627f
C2406 VDD.n1025 VSS 0.0107f
C2407 VDD.n1026 VSS 0.107f
C2408 VDD.n1027 VSS 0.0107f
C2409 VDD.t155 VSS 0.00808f
C2410 VDD.t301 VSS 0.00929f
C2411 VDD.n1028 VSS 0.0384f
C2412 VDD.n1029 VSS 0.214f
C2413 VDD.n1030 VSS 0.0416f
C2414 VDD.t154 VSS 0.0591f
C2415 VDD.n1031 VSS 0.0609f
C2416 VDD.n1032 VSS 0.0107f
C2417 VDD.n1033 VSS 0.0183f
C2418 VDD.n1034 VSS 0.109f
C2419 VDD.n1035 VSS 0.0107f
C2420 VDD.n1036 VSS 0.0183f
C2421 VDD.t93 VSS 0.0552f
C2422 VDD.n1037 VSS 0.0552f
C2423 VDD.n1038 VSS 0.0107f
C2424 VDD.n1039 VSS 0.0169f
C2425 VDD.n1040 VSS 0.143f
C2426 VDD.t96 VSS 0.0581f
C2427 VDD.n1041 VSS 0.0701f
C2428 VDD.n1042 VSS 0.0107f
C2429 VDD.n1043 VSS 0.0159f
C2430 VDD.n1044 VSS 0.131f
C2431 VDD.n1045 VSS 0.0107f
C2432 VDD.n1046 VSS 0.0185f
C2433 VDD.n1047 VSS 0.102f
C2434 VDD.n1048 VSS 0.0331f
C2435 VDD.n1049 VSS 0.0365f
C2436 VDD.n1050 VSS 0.0107f
C2437 VDD.t268 VSS 0.0591f
C2438 VDD.n1051 VSS 0.0609f
C2439 VDD.n1052 VSS 0.0107f
C2440 VDD.n1053 VSS 0.0183f
C2441 VDD.n1054 VSS 0.109f
C2442 VDD.n1055 VSS 0.0107f
C2443 VDD.n1056 VSS 0.0183f
C2444 VDD.n1057 VSS 0.0183f
C2445 VDD.n1058 VSS 0.107f
C2446 VDD.n1059 VSS 0.0107f
C2447 VDD.t262 VSS 0.0552f
C2448 VDD.n1060 VSS 0.0627f
C2449 VDD.n1061 VSS 0.0107f
C2450 VDD.n1062 VSS 0.0177f
C2451 VDD.n1063 VSS 0.0997f
C2452 VDD.n1064 VSS 0.0107f
C2453 VDD.n1065 VSS 0.0185f
C2454 VDD.t259 VSS 0.0581f
C2455 VDD.n1066 VSS 0.0701f
C2456 VDD.n1067 VSS 0.0107f
C2457 VDD.n1068 VSS 0.0185f
C2458 VDD.n1069 VSS 0.131f
C2459 VDD.n1070 VSS 0.0107f
C2460 VDD.n1071 VSS 0.0135f
C2461 VDD.n1072 VSS 0.103f
C2462 VDD.n1073 VSS 0.117f
C2463 VDD.n1074 VSS 0.073f
C2464 VDD.n1075 VSS 0.0289f
C2465 VDD.n1076 VSS 0.0238f
C2466 VDD.n1077 VSS 0.0165f
C2467 VDD.n1078 VSS 0.0165f
C2468 VDD.n1079 VSS 0.0238f
C2469 VDD.n1080 VSS 0.0165f
C2470 VDD.n1081 VSS 0.0083f
C2471 VDD.n1082 VSS 0.0218f
C2472 VDD.n1083 VSS 0.0237f
C2473 VDD.n1084 VSS 0.0165f
C2474 VDD.n1085 VSS 0.0164f
C2475 VDD.n1086 VSS 0.0139f
C2476 VDD.n1087 VSS 0.0132f
C2477 VDD.n1088 VSS 0.0165f
C2478 VDD.n1089 VSS 0.0165f
C2479 VDD.n1090 VSS 0.0225f
C2480 VDD.n1091 VSS 0.0165f
C2481 VDD.n1092 VSS 0.00891f
C2482 VDD.n1093 VSS 0.0138f
C2483 VDD.n1094 VSS 0.0239f
C2484 VDD.n1095 VSS 0.0165f
C2485 VDD.n1096 VSS 0.00987f
C2486 VDD.n1097 VSS 0.0119f
C2487 VDD.n1098 VSS 0.0932f
C2488 VDD.n1099 VSS 0.0348f
C2489 VDD.n1100 VSS 0.0223f
C2490 VDD.n1101 VSS 0.0174f
C2491 VDD.n1102 VSS 0.0175f
C2492 VDD.n1103 VSS 0.0156f
C2493 VDD.n1104 VSS 0.0514f
C2494 VDD.n1106 VSS 0.0116f
C2495 VDD.n1107 VSS 0.0103f
C2496 VDD.n1108 VSS 0.0506f
C2497 VDD.n1109 VSS 0.316f
C2498 VDD.n1110 VSS 0.0228f
C2499 VDD.n1111 VSS 0.022f
C2500 VDD.t220 VSS 0.0917f
C2501 VDD.t193 VSS 0.00749f
C2502 VDD.t202 VSS 0.0487f
C2503 VDD.n1112 VSS 0.279f
C2504 VDD.n1113 VSS 0.0218f
C2505 VDD.n1114 VSS 0.0211f
C2506 VDD.n1115 VSS 0.223f
C2507 VDD.n1116 VSS 0.0181f
C2508 VDD.n1117 VSS 0.0175f
C2509 VDD.n1118 VSS 0.223f
C2510 VDD.n1119 VSS 0.0171f
C2511 VDD.n1120 VSS 0.0165f
C2512 VDD.n1121 VSS 0.223f
C2513 VDD.n1122 VSS 0.0171f
C2514 VDD.n1123 VSS 0.0165f
C2515 VDD.t10 VSS 0.206f
C2516 VDD.n1124 VSS 0.0187f
C2517 VDD.n1125 VSS 0.0171f
C2518 VDD.n1126 VSS 0.0165f
C2519 VDD.n1127 VSS 0.223f
C2520 VDD.n1128 VSS 0.0171f
C2521 VDD.n1129 VSS 0.0095f
C2522 VDD.n1130 VSS 0.0189f
C2523 VDD.t8 VSS 0.206f
C2524 VDD.n1131 VSS 0.0823f
C2525 VDD.n1132 VSS 0.0171f
C2526 VDD.n1133 VSS 0.0153f
C2527 VDD.n1134 VSS 0.223f
C2528 VDD.n1135 VSS 0.0171f
C2529 VDD.n1136 VSS 0.0165f
C2530 VDD.n1137 VSS 0.146f
C2531 VDD.n1138 VSS 0.0171f
C2532 VDD.n1139 VSS 0.0165f
C2533 VDD.n1140 VSS 0.223f
C2534 VDD.n1141 VSS 0.0171f
C2535 VDD.n1142 VSS 0.0142f
C2536 VDD.n1143 VSS 0.0189f
C2537 VDD.n1144 VSS 0.21f
C2538 VDD.n1145 VSS 0.0171f
C2539 VDD.n1146 VSS 0.0105f
C2540 VDD.n1147 VSS 0.223f
C2541 VDD.n1148 VSS 0.0171f
C2542 VDD.n1149 VSS 0.0165f
C2543 VDD.n1150 VSS 0.223f
C2544 VDD.n1151 VSS 0.0171f
C2545 VDD.n1152 VSS 0.0165f
C2546 VDD.n1153 VSS 0.223f
C2547 VDD.n1154 VSS 0.0171f
C2548 VDD.n1155 VSS 0.0165f
C2549 VDD.n1156 VSS 0.223f
C2550 VDD.n1157 VSS 0.0171f
C2551 VDD.n1158 VSS 0.0165f
C2552 VDD.t29 VSS 0.206f
C2553 VDD.n1159 VSS 0.0618f
C2554 VDD.n1160 VSS 0.0171f
C2555 VDD.n1161 VSS 0.0165f
C2556 VDD.n1162 VSS 0.223f
C2557 VDD.n1163 VSS 0.0171f
C2558 VDD.n1164 VSS 0.0111f
C2559 VDD.n1165 VSS 0.0189f
C2560 VDD.n1166 VSS 0.125f
C2561 VDD.n1167 VSS 0.0171f
C2562 VDD.n1168 VSS 0.0137f
C2563 VDD.n1169 VSS 0.223f
C2564 VDD.n1170 VSS 0.0171f
C2565 VDD.n1171 VSS 0.0165f
C2566 VDD.n1172 VSS 0.189f
C2567 VDD.n1173 VSS 0.0171f
C2568 VDD.n1174 VSS 0.0165f
C2569 VDD.n1175 VSS 0.223f
C2570 VDD.n1176 VSS 0.0171f
C2571 VDD.n1177 VSS 0.0158f
C2572 VDD.n1178 VSS 0.0189f
C2573 VDD.n1179 VSS 0.223f
C2574 VDD.n1180 VSS 0.0171f
C2575 VDD.n1181 VSS 0.00894f
C2576 VDD.t0 VSS 0.206f
C2577 VDD.n1182 VSS 0.0299f
C2578 VDD.n1183 VSS 0.0171f
C2579 VDD.n1184 VSS 0.0165f
C2580 VDD.n1185 VSS 0.223f
C2581 VDD.n1186 VSS 0.0171f
C2582 VDD.n1187 VSS 0.0165f
C2583 VDD.n1188 VSS 0.223f
C2584 VDD.n1189 VSS 0.0171f
C2585 VDD.n1190 VSS 0.0165f
C2586 VDD.n1191 VSS 0.262f
C2587 VDD.n1192 VSS 0.0194f
C2588 VDD.n1193 VSS 0.0187f
C2589 VDD.t233 VSS 0.245f
C2590 VDD.t205 VSS 0.0281f
C2591 VDD.n1194 VSS 0.133f
C2592 VDD.n1195 VSS 0.0211f
C2593 VDD.n1196 VSS 0.0205f
C2594 VDD.n1197 VSS 0.399f
C2595 VDD.n1198 VSS 0.0219f
C2596 VDD.n1199 VSS 0.0243f
C2597 VDD.n1200 VSS 0.0308f
C2598 VDD.n1202 VSS 0.0243f
C2599 VDD.n1203 VSS 0.016f
C2600 VDD.n1204 VSS 0.0198f
C2601 VDD.n1205 VSS 0.0154f
C2602 VDD.n1206 VSS 0.0198f
C2603 VDD.n1207 VSS 0.0127f
C2604 VDD.n1208 VSS 0.0209f
C2605 VDD.n1209 VSS 0.0198f
C2606 VDD.n1210 VSS 0.0103f
C2607 VDD.n1211 VSS 0.0198f
C2608 VDD.n1212 VSS 0.0154f
C2609 VDD.n1214 VSS 0.0198f
C2610 VDD.n1215 VSS 0.0154f
C2611 VDD.n1216 VSS 0.0198f
C2612 VDD.n1217 VSS 0.00808f
C2613 VDD.n1218 VSS 0.0209f
C2614 VDD.n1220 VSS 0.0198f
C2615 VDD.n1221 VSS 0.015f
C2616 VDD.n1222 VSS 0.0198f
C2617 VDD.n1223 VSS 0.0154f
C2618 VDD.n1225 VSS 0.0198f
C2619 VDD.n1226 VSS 0.0121f
C2620 VDD.n1227 VSS 0.0209f
C2621 VDD.n1228 VSS 0.0198f
C2622 VDD.n1229 VSS 0.011f
C2623 VDD.n1231 VSS 0.0198f
C2624 VDD.n1232 VSS 0.0154f
C2625 VDD.n1233 VSS 0.0198f
C2626 VDD.n1234 VSS 0.0154f
C2627 VDD.n1236 VSS 0.0198f
C2628 VDD.n1237 VSS 0.00782f
C2629 VDD.n1238 VSS 0.0209f
C2630 VDD.n1239 VSS 0.0198f
C2631 VDD.n1240 VSS 0.0153f
C2632 VDD.n1242 VSS 0.533f
C2633 VDD.n1244 VSS 0.0376f
C2634 VDD.n1245 VSS 0.01f
C2635 VDD.n1246 VSS 0.0342f
C2636 VDD.t273 VSS 0.00405f
C2637 VDD.n1247 VSS 0.00405f
C2638 VDD.n1248 VSS 0.0081f
C2639 VDD.n1249 VSS 0.0228f
C2640 VDD.t289 VSS 0.00405f
C2641 VDD.n1250 VSS 0.00405f
C2642 VDD.n1251 VSS 0.0081f
C2643 VDD.n1252 VSS 0.0224f
C2644 VDD.n1253 VSS 0.0342f
C2645 VDD.t20 VSS 0.00405f
C2646 VDD.n1254 VSS 0.00405f
C2647 VDD.n1255 VSS 0.0081f
C2648 VDD.n1256 VSS 0.0132f
C2649 VDD.n1257 VSS 0.0347f
C2650 VDD.n1258 VSS 0.178f
C2651 VDD.n1259 VSS 0.0176f
C2652 VDD.n1260 VSS 0.0166f
C2653 VDD.n1261 VSS 0.0277f
C2654 VDD.t17 VSS 0.00405f
C2655 VDD.n1262 VSS 0.00405f
C2656 VDD.n1263 VSS 0.0081f
C2657 VDD.n1264 VSS 0.0206f
C2658 VDD.t37 VSS 0.00405f
C2659 VDD.n1265 VSS 0.00405f
C2660 VDD.n1266 VSS 0.0081f
C2661 VDD.n1267 VSS 0.02f
C2662 VDD.t266 VSS 0.00405f
C2663 VDD.n1268 VSS 0.00405f
C2664 VDD.n1269 VSS 0.0081f
C2665 VDD.n1270 VSS 0.0206f
C2666 VDD.t284 VSS 0.00405f
C2667 VDD.n1271 VSS 0.00405f
C2668 VDD.n1272 VSS 0.0081f
C2669 VDD.n1273 VSS 0.02f
C2670 VDD.n1274 VSS 0.0342f
C2671 VDD.n1275 VSS 0.0268f
C2672 VDD.n1276 VSS 0.0378f
C2673 VDD.t267 VSS 0.00405f
C2674 VDD.n1277 VSS 0.00405f
C2675 VDD.n1278 VSS 0.0081f
C2676 VDD.n1279 VSS 0.0136f
C2677 VDD.t9 VSS 0.00405f
C2678 VDD.n1280 VSS 0.00405f
C2679 VDD.n1281 VSS 0.0081f
C2680 VDD.n1282 VSS 0.0166f
C2681 VDD.n1283 VSS 0.0351f
C2682 VDD.n1284 VSS 0.223f
C2683 VDD.n1285 VSS 0.0176f
C2684 VDD.n1286 VSS 0.0234f
C2685 VDD.n1287 VSS 0.223f
C2686 VDD.n1288 VSS 0.0176f
C2687 VDD.n1289 VSS 0.0171f
C2688 VDD.n1290 VSS 0.223f
C2689 VDD.n1291 VSS 0.0176f
C2690 VDD.n1292 VSS 0.018f
C2691 VDD.n1293 VSS 0.223f
C2692 VDD.n1294 VSS 0.0176f
C2693 VDD.n1295 VSS 0.0234f
C2694 VDD.t16 VSS 0.206f
C2695 VDD.n1296 VSS 0.0299f
C2696 VDD.n1297 VSS 0.0176f
C2697 VDD.n1298 VSS 0.0234f
C2698 VDD.n1299 VSS 0.223f
C2699 VDD.n1300 VSS 0.0176f
C2700 VDD.n1301 VSS 0.014f
C2701 VDD.t201 VSS 0.0338f
C2702 VDD.t203 VSS 0.0177f
C2703 VDD.n1302 VSS 0.0805f
C2704 VDD.t369 VSS 0.00405f
C2705 VDD.n1303 VSS 0.00405f
C2706 VDD.n1304 VSS 0.0081f
C2707 VDD.t394 VSS 0.00405f
C2708 VDD.n1305 VSS 0.00405f
C2709 VDD.n1306 VSS 0.0116f
C2710 VDD.n1307 VSS 0.0356f
C2711 VDD.t219 VSS 0.0338f
C2712 VDD.t221 VSS 0.0177f
C2713 VDD.n1308 VSS 0.0797f
C2714 VDD.t395 VSS 0.00405f
C2715 VDD.n1309 VSS 0.00405f
C2716 VDD.n1310 VSS 0.0081f
C2717 VDD.t371 VSS 0.00405f
C2718 VDD.n1311 VSS 0.00405f
C2719 VDD.n1312 VSS 0.0116f
C2720 VDD.n1313 VSS 0.0356f
C2721 VDD.t192 VSS 0.0574f
C2722 VDD.t194 VSS 0.0177f
C2723 VDD.n1314 VSS 0.0798f
C2724 VDD.t335 VSS 0.00808f
C2725 VDD.t368 VSS 0.0103f
C2726 VDD.n1315 VSS 0.0481f
C2727 VDD.t240 VSS 0.0338f
C2728 VDD.t241 VSS 0.0177f
C2729 VDD.n1316 VSS 0.0797f
C2730 VDD.n1317 VSS 0.0256f
C2731 VDD.n1318 VSS 0.024f
C2732 VDD.n1319 VSS 0.0111f
C2733 VDD.n1320 VSS 0.0198f
C2734 VDD.n1321 VSS 0.0223f
C2735 VDD.n1322 VSS 0.0113f
C2736 VDD.n1324 VSS 0.0191f
C2737 VDD.n1325 VSS 0.0146f
C2738 VDD.n1326 VSS 0.0215f
C2739 VDD.n1327 VSS 0.016f
C2740 VDD.n1328 VSS 0.00962f
C2741 VDD.n1330 VSS 0.0175f
C2742 VDD.n1331 VSS 0.00772f
C2743 VDD.n1332 VSS 0.0183f
C2744 VDD.n1333 VSS 0.0191f
C2745 VDD.n1334 VSS 0.0163f
C2746 VDD.n1335 VSS 0.0229f
C2747 VDD.n1337 VSS 0.0192f
C2748 VDD.n1338 VSS 0.00877f
C2749 VDD.n1339 VSS 0.0191f
C2750 VDD.n1340 VSS 0.0171f
C2751 VDD.n1342 VSS 0.0191f
C2752 VDD.n1343 VSS 0.0105f
C2753 VDD.n1344 VSS 0.0184f
C2754 VDD.n1345 VSS 0.0176f
C2755 VDD.n1346 VSS 0.00792f
C2756 VDD.n1347 VSS 0.0214f
C2757 VDD.n1349 VSS 0.316f
C2758 VDD.n1351 VSS 0.016f
C2759 VDD.n1352 VSS 0.0129f
C2760 VDD.n1353 VSS 0.0152f
C2761 VDD.n1354 VSS 0.0137f
C2762 VDD.n1355 VSS 0.0859f
C2763 VDD.n1356 VSS 0.0204f
C2764 VDD.t249 VSS 0.032f
C2765 VDD.t251 VSS 0.0172f
C2766 VDD.n1357 VSS 0.0834f
C2767 VDD.t198 VSS 0.033f
C2768 VDD.t200 VSS 0.0173f
C2769 VDD.n1358 VSS 0.0832f
C2770 VDD.t44 VSS 0.00405f
C2771 VDD.n1359 VSS 0.00405f
C2772 VDD.n1360 VSS 0.0099f
C2773 VDD.t45 VSS 0.00405f
C2774 VDD.n1361 VSS 0.00405f
C2775 VDD.n1362 VSS 0.0081f
C2776 VDD.n1363 VSS 0.0254f
C2777 VDD.n1364 VSS 0.0159f
C2778 VDD.t5 VSS 0.0552f
C2779 VDD.n1365 VSS 0.0552f
C2780 VDD.n1366 VSS 0.0107f
C2781 VDD.n1367 VSS 0.214f
C2782 VDD.t15 VSS 0.00929f
C2783 VDD.t14 VSS 0.00808f
C2784 VDD.n1368 VSS 0.0373f
C2785 VDD.n1369 VSS 0.00913f
C2786 VDD.n1370 VSS 0.00808f
C2787 VDD.n1371 VSS 0.0503f
C2788 VDD.t80 VSS 0.00405f
C2789 VDD.n1372 VSS 0.00405f
C2790 VDD.n1373 VSS 0.0099f
C2791 VDD.t89 VSS 0.00405f
C2792 VDD.n1374 VSS 0.00405f
C2793 VDD.n1375 VSS 0.0081f
C2794 VDD.n1376 VSS 0.0254f
C2795 VDD.n1377 VSS 0.0159f
C2796 VDD.t61 VSS 0.0552f
C2797 VDD.n1378 VSS 0.0552f
C2798 VDD.n1379 VSS 0.0107f
C2799 VDD.t390 VSS 0.00929f
C2800 VDD.t386 VSS 0.00808f
C2801 VDD.n1380 VSS 0.0384f
C2802 VDD.n1381 VSS 0.214f
C2803 VDD.n1382 VSS 0.0416f
C2804 VDD.t385 VSS 0.0591f
C2805 VDD.n1383 VSS 0.0609f
C2806 VDD.n1384 VSS 0.0107f
C2807 VDD.n1385 VSS 0.0183f
C2808 VDD.n1386 VSS 0.109f
C2809 VDD.n1387 VSS 0.0107f
C2810 VDD.n1388 VSS 0.0183f
C2811 VDD.n1389 VSS 0.0183f
C2812 VDD.n1390 VSS 0.107f
C2813 VDD.n1391 VSS 0.0107f
C2814 VDD.t79 VSS 0.0552f
C2815 VDD.n1392 VSS 0.0627f
C2816 VDD.n1393 VSS 0.0107f
C2817 VDD.n1394 VSS 0.0177f
C2818 VDD.n1395 VSS 0.0997f
C2819 VDD.n1396 VSS 0.0107f
C2820 VDD.n1397 VSS 0.0185f
C2821 VDD.t387 VSS 0.0581f
C2822 VDD.n1398 VSS 0.0701f
C2823 VDD.n1399 VSS 0.0107f
C2824 VDD.n1400 VSS 0.0185f
C2825 VDD.n1401 VSS 0.131f
C2826 VDD.n1402 VSS 0.0107f
C2827 VDD.n1403 VSS 0.0185f
C2828 VDD.n1404 VSS 0.102f
C2829 VDD.n1405 VSS 0.0311f
C2830 VDD.n1406 VSS 0.0351f
C2831 VDD.n1407 VSS 0.0107f
C2832 VDD.t13 VSS 0.0591f
C2833 VDD.n1408 VSS 0.0609f
C2834 VDD.n1409 VSS 0.0107f
C2835 VDD.n1410 VSS 0.0183f
C2836 VDD.n1411 VSS 0.109f
C2837 VDD.n1412 VSS 0.0107f
C2838 VDD.n1413 VSS 0.0183f
C2839 VDD.n1414 VSS 0.0183f
C2840 VDD.n1415 VSS 0.107f
C2841 VDD.n1416 VSS 0.0107f
C2842 VDD.t43 VSS 0.0552f
C2843 VDD.n1417 VSS 0.0627f
C2844 VDD.n1418 VSS 0.0107f
C2845 VDD.n1419 VSS 0.0177f
C2846 VDD.n1420 VSS 0.0997f
C2847 VDD.n1421 VSS 0.0107f
C2848 VDD.n1422 VSS 0.0185f
C2849 VDD.t26 VSS 0.0581f
C2850 VDD.n1423 VSS 0.0701f
C2851 VDD.n1424 VSS 0.0107f
C2852 VDD.n1425 VSS 0.0185f
C2853 VDD.n1426 VSS 0.131f
C2854 VDD.n1427 VSS 0.0107f
C2855 VDD.n1428 VSS 0.0185f
C2856 VDD.n1429 VSS 0.119f
C2857 VDD.n1430 VSS 0.00922f
C2858 VDD.n1431 VSS 0.00808f
C2859 VDD.n1432 VSS 0.0369f
C2860 VDD.n1433 VSS 0.0888f
C2861 VDD.n1434 VSS 0.0165f
C2862 VDD.n1435 VSS 0.0155f
C2863 VDD.n1437 VSS 0.0165f
C2864 VDD.n1438 VSS 0.0155f
C2865 VDD.n1440 VSS 0.0165f
C2866 VDD.n1441 VSS 0.0155f
C2867 VDD.n1443 VSS 0.0165f
C2868 VDD.n1444 VSS 0.0155f
C2869 VDD.n1446 VSS 0.0165f
C2870 VDD.n1447 VSS 0.0155f
C2871 VDD.n1449 VSS 0.0165f
C2872 VDD.n1450 VSS 0.0155f
C2873 VDD.n1452 VSS 0.0165f
C2874 VDD.n1453 VSS 0.0155f
C2875 VDD.n1455 VSS 0.0165f
C2876 VDD.n1456 VSS 0.0155f
C2877 VDD.n1458 VSS 0.0165f
C2878 VDD.n1459 VSS 0.0155f
C2879 VDD.n1461 VSS 0.0163f
C2880 VDD.n1462 VSS 0.0153f
C2881 VDD.n1464 VSS 0.0163f
C2882 VDD.n1465 VSS 0.0153f
C2883 VDD.n1466 VSS 0.999f
C2884 VDD.n1468 VSS 0.0428f
C2885 VDD.n1469 VSS 0.029f
C2886 VDD.n1470 VSS 0.112f
C2887 VDD.n1471 VSS 0.122f
C2888 VDD.n1472 VSS 0.0173f
C2889 VDD.n1473 VSS 0.0641f
C2890 VDD.n1474 VSS 0.0165f
C2891 VDD.n1475 VSS 0.0129f
C2892 VDD.n1476 VSS 0.0645f
C2893 VDD.n1477 VSS 0.0165f
C2894 VDD.n1478 VSS 0.0103f
C2895 VDD.n1479 VSS 0.0215f
C2896 VDD.t225 VSS 0.728f
C2897 VDD.t199 VSS 0.484f
C2898 VDD.n1481 VSS 0.0384f
C2899 VDD.n1482 VSS 0.0165f
C2900 VDD.n1483 VSS 0.0124f
C2901 VDD.n1484 VSS 0.0322f
C2902 VDD.n1485 VSS 0.029f
C2903 VDD.n1486 VSS 0.0165f
C2904 VDD.n1487 VSS 0.0151f
C2905 VDD.n1488 VSS 0.0605f
C2906 VDD.n1489 VSS 0.0165f
C2907 VDD.n1490 VSS 0.00966f
C2908 VDD.n1491 VSS 0.0223f
C2909 VDD.t217 VSS 0.417f
C2910 VDD.t330 VSS 0.00374f
C2911 VDD.n1492 VSS 0.674f
C2912 VDD.t250 VSS 0.261f
C2913 VDD.n1493 VSS 0.0381f
C2914 VDD.n1494 VSS 0.0165f
C2915 VDD.n1495 VSS 0.0131f
C2916 VDD.n1496 VSS 0.0598f
C2917 VDD.n1497 VSS 0.0225f
C2918 VDD.n1498 VSS 0.0207f
C2919 VDD.n1499 VSS 0.0257f
C2920 VDD.n1500 VSS 0.0241f
C2921 VDD.n1501 VSS 0.0194f
C2922 VDD.n1502 VSS 0.0169f
C2923 VDD.n1503 VSS 0.588f
C2924 VDD.n1504 VSS 0.00688f
C2925 VDD.n1505 VSS 0.0223f
C2926 VDD.n1506 VSS 0.0183f
C2927 VDD.n1507 VSS 0.0196f
C2928 VDD.n1508 VSS 0.283f
C2929 VDD.n1509 VSS 0.0182f
C2930 VDD.n1510 VSS 0.017f
C2931 VDD.n1511 VSS 0.266f
C2932 VDD.n1512 VSS 0.0273f
C2933 VDD.n1513 VSS 0.0278f
C2934 VDD.n1514 VSS 0.251f
C2935 VDD.n1515 VSS 0.0236f
C2936 VDD.n1516 VSS 0.0322f
C2937 VDD.n1517 VSS 0.223f
C2938 VDD.n1518 VSS 0.0176f
C2939 VDD.n1519 VSS 0.0234f
C2940 VDD.n1520 VSS 0.223f
C2941 VDD.n1521 VSS 0.0176f
C2942 VDD.n1522 VSS 0.0234f
C2943 VDD.n1523 VSS 0.223f
C2944 VDD.n1524 VSS 0.0176f
C2945 VDD.n1525 VSS 0.0234f
C2946 VDD.n1526 VSS 0.221f
C2947 VDD.n1527 VSS 0.0176f
C2948 VDD.n1528 VSS 0.0143f
C2949 VDD.n1529 VSS 0.0192f
C2950 VDD.n1530 VSS 0.223f
C2951 VDD.n1531 VSS 0.0176f
C2952 VDD.n1532 VSS 0.0207f
C2953 VDD.n1533 VSS 0.157f
C2954 VDD.n1534 VSS 0.0176f
C2955 VDD.n1535 VSS 0.0234f
C2956 VDD.n1536 VSS 0.223f
C2957 VDD.n1537 VSS 0.0176f
C2958 VDD.n1538 VSS 0.0234f
C2959 VDD.t2 VSS 0.206f
C2960 VDD.n1539 VSS 0.0936f
C2961 VDD.n1540 VSS 0.0176f
C2962 VDD.n1541 VSS 0.021f
C2963 VDD.n1542 VSS 0.0182f
C2964 VDD.n1543 VSS 0.0605f
C2965 VDD.t288 VSS 0.00405f
C2966 VDD.n1544 VSS 0.00405f
C2967 VDD.n1545 VSS 0.0081f
C2968 VDD.n1546 VSS 0.0156f
C2969 VDD.n1547 VSS 0.0266f
C2970 VDD.n1548 VSS 0.0388f
C2971 VDD.t19 VSS 0.00405f
C2972 VDD.n1549 VSS 0.00405f
C2973 VDD.n1550 VSS 0.0081f
C2974 VDD.n1551 VSS 0.0207f
C2975 VDD.t40 VSS 0.00405f
C2976 VDD.n1552 VSS 0.00405f
C2977 VDD.n1553 VSS 0.0081f
C2978 VDD.n1554 VSS 0.0198f
C2979 VDD.n1555 VSS 0.0386f
C2980 VDD.n1556 VSS 0.0275f
C2981 VDD.t270 VSS 0.00405f
C2982 VDD.n1557 VSS 0.00405f
C2983 VDD.n1558 VSS 0.0081f
C2984 VDD.n1559 VSS 0.0141f
C2985 VDD.n1560 VSS 0.0625f
C2986 VDD.n1561 VSS 0.0192f
C2987 VDD.n1562 VSS 0.223f
C2988 VDD.n1563 VSS 0.0176f
C2989 VDD.n1564 VSS 0.0185f
C2990 VDD.t18 VSS 0.206f
C2991 VDD.n1565 VSS 0.114f
C2992 VDD.n1566 VSS 0.0176f
C2993 VDD.n1567 VSS 0.0234f
C2994 VDD.n1568 VSS 0.223f
C2995 VDD.n1569 VSS 0.0176f
C2996 VDD.n1570 VSS 0.0234f
C2997 VDD.t23 VSS 0.206f
C2998 VDD.n1571 VSS 0.0505f
C2999 VDD.n1572 VSS 0.0176f
C3000 VDD.n1573 VSS 0.0233f
C3001 VDD.n1574 VSS 0.0182f
C3002 VDD.n1575 VSS 0.223f
C3003 VDD.n1576 VSS 0.0176f
C3004 VDD.n1577 VSS 0.0118f
C3005 VDD.n1578 VSS 0.223f
C3006 VDD.n1579 VSS 0.0176f
C3007 VDD.n1580 VSS 0.0234f
C3008 VDD.n1581 VSS 0.21f
C3009 VDD.n1582 VSS 0.0176f
C3010 VDD.n1583 VSS 0.0234f
C3011 VDD.n1584 VSS 0.223f
C3012 VDD.n1585 VSS 0.0176f
C3013 VDD.n1586 VSS 0.0234f
C3014 VDD.n1587 VSS 0.223f
C3015 VDD.n1588 VSS 0.0192f
C3016 VDD.n1589 VSS 0.0254f
C3017 VDD.n1590 VSS 0.283f
C3018 VDD.n1591 VSS 0.0221f
C3019 VDD.n1592 VSS 0.0279f
C3020 VDD.n1593 VSS 0.159f
C3021 VDD.n1594 VSS 0.0349f
C3022 VDD.n1595 VSS 0.0294f
C3023 VDD.n1596 VSS 0.0434f
C3024 VDD.n1597 VSS 0.083f
C3025 VCO_C_0.INV_2_3.IN.n0 VSS 0.561f
C3026 VCO_C_0.INV_2_3.IN.n1 VSS 0.678f
C3027 VCO_C_0.INV_2_3.IN.n2 VSS 0.0733f
C3028 VCO_C_0.INV_2_3.IN.n3 VSS 0.828f
C3029 VCO_C_0.INV_2_3.IN.t11 VSS 0.0244f
C3030 VCO_C_0.INV_2_3.IN.n4 VSS 0.282f
C3031 VCO_C_0.INV_2_3.IN.t40 VSS 0.118f
C3032 VCO_C_0.INV_2_3.IN.t53 VSS 0.124f
C3033 VCO_C_0.INV_2_3.IN.t45 VSS 0.124f
C3034 VCO_C_0.INV_2_3.IN.t37 VSS 0.12f
C3035 VCO_C_0.INV_2_3.IN.n5 VSS 0.041f
C3036 VCO_C_0.INV_2_3.IN.n6 VSS 0.145f
C3037 VCO_C_0.INV_2_3.IN.t30 VSS 0.123f
C3038 VCO_C_0.INV_2_3.IN.t34 VSS 0.124f
C3039 VCO_C_0.INV_2_3.IN.t33 VSS 0.124f
C3040 VCO_C_0.INV_2_3.IN.t46 VSS 0.143f
C3041 VCO_C_0.INV_2_3.IN.n7 VSS 0.499f
C3042 VCO_C_0.INV_2_3.IN.n8 VSS 0.265f
C3043 VCO_C_0.INV_2_3.IN.n9 VSS 0.3f
C3044 VCO_C_0.INV_2_3.IN.n10 VSS 0.172f
C3045 VCO_C_0.INV_2_3.IN.n11 VSS 0.231f
C3046 VCO_C_0.INV_2_3.IN.n12 VSS 0.277f
C3047 VCO_C_0.INV_2_3.IN.n13 VSS 0.272f
C3048 VCO_C_0.INV_2_3.IN.n14 VSS 0.233f
C3049 VCO_C_0.INV_2_3.IN.t52 VSS 0.118f
C3050 VCO_C_0.INV_2_3.IN.t39 VSS 0.123f
C3051 VCO_C_0.INV_2_3.IN.t56 VSS 0.123f
C3052 VCO_C_0.INV_2_3.IN.t49 VSS 0.117f
C3053 VCO_C_0.INV_2_3.IN.t42 VSS 0.121f
C3054 VCO_C_0.INV_2_3.IN.t47 VSS 0.126f
C3055 VCO_C_0.INV_2_3.IN.t44 VSS 0.126f
C3056 VCO_C_0.INV_2_3.IN.t57 VSS 0.13f
C3057 VCO_C_0.INV_2_3.IN.n15 VSS 0.515f
C3058 VCO_C_0.INV_2_3.IN.n16 VSS 0.271f
C3059 VCO_C_0.INV_2_3.IN.n17 VSS 0.331f
C3060 VCO_C_0.INV_2_3.IN.n18 VSS 0.324f
C3061 VCO_C_0.INV_2_3.IN.n19 VSS 0.27f
C3062 VCO_C_0.INV_2_3.IN.n20 VSS 0.277f
C3063 VCO_C_0.INV_2_3.IN.t15 VSS 0.0278f
C3064 VCO_C_0.INV_2_3.IN.n21 VSS 0.28f
C3065 VCO_C_0.INV_2_3.IN.n22 VSS 0.0245f
C3066 VCO_C_0.INV_2_3.IN.n23 VSS 0.0731f
C3067 VCO_C_0.INV_2_3.IN.n24 VSS 0.0563f
C3068 VCO_C_0.INV_2_3.IN.n25 VSS 0.0183f
C3069 VCO_C_0.INV_2_3.IN.t17 VSS 0.0161f
C3070 VCO_C_0.INV_2_3.IN.n26 VSS 0.155f
C3071 VCO_C_0.INV_2_3.IN.n27 VSS 0.818f
C3072 VCO_C_0.INV_2_3.IN.n28 VSS 0.288f
C3073 VCO_C_0.INV_2_3.IN.n29 VSS 0.334f
C3074 VCO_C_0.INV_2_3.IN.n30 VSS 0.0736f
C3075 VCO_C_0.INV_2_3.IN.t12 VSS 0.0173f
C3076 VCO_C_0.INV_2_3.IN.n31 VSS 0.0173f
C3077 VCO_C_0.INV_2_3.IN.n32 VSS 0.0862f
C3078 VCO_C_0.INV_2_3.IN.t14 VSS 0.0245f
C3079 VCO_C_0.INV_2_3.IN.n33 VSS 0.073f
C3080 VCO_C_0.INV_2_3.IN.n34 VSS 0.0517f
C3081 VCO_C_0.INV_2_3.IN.t13 VSS 0.0173f
C3082 VCO_C_0.INV_2_3.IN.n35 VSS 0.0173f
C3083 VCO_C_0.INV_2_3.IN.n36 VSS 0.0881f
C3084 VCO_C_0.INV_2_3.IN.t16 VSS 0.0173f
C3085 VCO_C_0.INV_2_3.IN.n37 VSS 0.0173f
C3086 VCO_C_0.INV_2_3.IN.n38 VSS 0.0347f
C3087 VCO_C_0.INV_2_3.IN.n39 VSS 0.0617f
C3088 VCO_C_0.INV_2_3.IN.n40 VSS 0.433f
C3089 VCO_C_0.INV_2_3.IN.n41 VSS 0.622f
C3090 VCO_C_0.INV_2_3.IN.n42 VSS 0.0279f
C3091 VCO_C_0.INV_2_3.IN.n43 VSS 0.0697f
C3092 VCO_C_0.INV_2_3.IN.n44 VSS 0.0509f
C3093 VCO_C_0.INV_2_3.IN.n45 VSS 0.632f
C3094 VCO_C_0.INV_2_3.IN.n46 VSS 0.494f
C3095 VCO_C_0.INV_2_3.IN.n47 VSS 0.439f
C3096 VCO_C_0.INV_2_3.IN.n48 VSS 0.0267f
C3097 VCO_C_0.INV_2_3.IN.n49 VSS 0.207f
C3098 VCO_C_0.INV_2_3.IN.n50 VSS 0.0291f
C3099 VCO_C_0.INV_2_3.IN.n51 VSS 0.688f
C3100 VCO_C_0.INV_2_3.IN.n52 VSS 0.252f
C3101 VCO_C_0.INV_2_3.IN.n53 VSS 0.0159f
C3102 VCO_C_0.INV_2_3.IN.t24 VSS 0.0187f
C3103 VCO_C_0.INV_2_3.IN.n54 VSS 0.163f
C3104 VCO_C_0.INV_2_3.IN.t21 VSS 0.0452f
C3105 VCO_C_0.INV_2_3.IN.n55 VSS 0.0159f
C3106 VCO_C_0.INV_2_3.IN.t2 VSS 0.0187f
C3107 VCO_C_0.INV_2_3.IN.n56 VSS 0.141f
C3108 VCO_C_0.INV_2_3.IN.n57 VSS 0.744f
C3109 VCO_C_0.INV_2_3.IN.t23 VSS 0.0298f
C3110 VCO_C_0.INV_2_3.IN.n58 VSS 0.305f
C3111 VCO_C_0.INV_2_3.IN.t4 VSS 0.0298f
C3112 VCO_C_0.INV_2_3.IN.n59 VSS 0.422f
C3113 VCO_C_0.INV_2_3.IN.n60 VSS 0.761f
C3114 VCO_C_0.INV_2_3.IN.n61 VSS 0.408f
C3115 VCO_C_0.INV_2_3.IN.n62 VSS 0.482f
C3116 VCO_C_0.INV_2_3.IN.t48 VSS 0.0431f
C3117 VCO_C_0.INV_2_3.IN.n63 VSS 0.0707f
C3118 VCO_C_0.INV_2_3.IN.n64 VSS 0.121f
C3119 VCO_C_0.INV_2_3.IN.t31 VSS 0.0571f
C3120 VCO_C_0.INV_2_3.IN.t51 VSS 0.139f
C3121 VCO_C_0.INV_2_3.IN.n65 VSS 0.0998f
C3122 VCO_C_0.INV_2_3.IN.t54 VSS 0.0432f
C3123 VCO_C_0.INV_2_3.IN.t50 VSS 0.106f
C3124 VCO_C_0.INV_2_3.IN.n66 VSS 0.124f
C3125 VCO_C_0.INV_2_3.IN.t41 VSS 0.0432f
C3126 VCO_C_0.INV_2_3.IN.t36 VSS 0.0432f
C3127 VCO_C_0.INV_2_3.IN.t32 VSS 0.106f
C3128 VCO_C_0.INV_2_3.IN.n67 VSS 0.14f
C3129 VCO_C_0.INV_2_3.IN.n68 VSS 0.14f
C3130 VCO_C_0.INV_2_3.IN.t38 VSS 0.106f
C3131 VCO_C_0.INV_2_3.IN.n69 VSS 0.121f
C3132 VCO_C_0.INV_2_3.IN.t55 VSS 0.0571f
C3133 VCO_C_0.INV_2_3.IN.n70 VSS 0.153f
C3134 VCO_C_0.INV_2_3.IN.n71 VSS 0.153f
C3135 VCO_C_0.INV_2_3.IN.t35 VSS 0.139f
C3136 VCO_C_0.INV_2_3.IN.n72 VSS 0.0998f
C3137 VCO_C_0.INV_2_3.IN.t43 VSS 0.091f
C3138 VCO_C_0.INV_2_3.IN.n73 VSS 0.0715f
C3139 VCO_C_0.INV_2_3.IN.n74 VSS 0.891f
C3140 VCO_C_0.INV_2_3.IN.n75 VSS 0.898f
C3141 VCO_C_0.INV_2_3.IN.n76 VSS 0.51f
C3142 VCO_C_0.INV_2_3.IN.n77 VSS 0.353f
C3143 VCO_C_0.INV_2_3.IN.t26 VSS 0.0181f
C3144 VCO_C_0.INV_2_3.IN.n78 VSS 0.0163f
C3145 VCO_C_0.INV_2_3.IN.n79 VSS 0.139f
C3146 VCO_C_0.INV_2_3.IN.n80 VSS 0.0416f
C3147 VCO_C_0.INV_2_3.IN.n81 VSS 0.583f
C3148 VCO_C_0.INV_2_3.IN.n82 VSS 0.0412f
C3149 VCO_C_0.INV_2_3.IN.t10 VSS 0.0712f
C3150 a_10161_4198.n0 VSS 0.144f
C3151 a_10161_4198.n1 VSS 0.0962f
C3152 a_10161_4198.n2 VSS 0.127f
C3153 a_10161_4198.n3 VSS 0.289f
C3154 a_10161_4198.t8 VSS 0.0108f
C3155 a_10161_4198.t15 VSS 0.0108f
C3156 a_10161_4198.n4 VSS 0.0108f
C3157 a_10161_4198.n5 VSS 0.0217f
C3158 a_10161_4198.t44 VSS 0.0108f
C3159 a_10161_4198.n6 VSS 0.0108f
C3160 a_10161_4198.n7 VSS 0.0217f
C3161 a_10161_4198.t23 VSS 0.0108f
C3162 a_10161_4198.n8 VSS 0.0108f
C3163 a_10161_4198.n9 VSS 0.0273f
C3164 a_10161_4198.t16 VSS 0.0108f
C3165 a_10161_4198.n10 VSS 0.0108f
C3166 a_10161_4198.n11 VSS 0.0217f
C3167 a_10161_4198.n12 VSS 0.0581f
C3168 a_10161_4198.t22 VSS 0.0108f
C3169 a_10161_4198.n13 VSS 0.0108f
C3170 a_10161_4198.n14 VSS 0.0217f
C3171 a_10161_4198.n15 VSS 0.042f
C3172 a_10161_4198.t58 VSS 0.0108f
C3173 a_10161_4198.n16 VSS 0.0108f
C3174 a_10161_4198.n17 VSS 0.0217f
C3175 a_10161_4198.t3 VSS 0.0108f
C3176 a_10161_4198.n18 VSS 0.0108f
C3177 a_10161_4198.n19 VSS 0.0217f
C3178 a_10161_4198.t42 VSS 0.0108f
C3179 a_10161_4198.n20 VSS 0.0108f
C3180 a_10161_4198.n21 VSS 0.0295f
C3181 a_10161_4198.t32 VSS 0.0108f
C3182 a_10161_4198.n22 VSS 0.0108f
C3183 a_10161_4198.n23 VSS 0.0217f
C3184 a_10161_4198.n24 VSS 0.424f
C3185 a_10161_4198.n25 VSS 0.0707f
C3186 a_10161_4198.t28 VSS 0.0108f
C3187 a_10161_4198.n26 VSS 0.0108f
C3188 a_10161_4198.n27 VSS 0.0217f
C3189 a_10161_4198.n28 VSS 0.392f
C3190 a_10161_4198.n29 VSS 0.118f
C3191 a_10161_4198.n30 VSS 0.159f
C3192 a_10161_4198.t5 VSS 0.0108f
C3193 a_10161_4198.n31 VSS 0.0108f
C3194 a_10161_4198.n32 VSS 0.0217f
C3195 a_10161_4198.t19 VSS 0.0108f
C3196 a_10161_4198.n33 VSS 0.0108f
C3197 a_10161_4198.n34 VSS 0.0217f
C3198 a_10161_4198.t34 VSS 0.0108f
C3199 a_10161_4198.n35 VSS 0.0108f
C3200 a_10161_4198.n36 VSS 0.0217f
C3201 a_10161_4198.t21 VSS 0.0108f
C3202 a_10161_4198.n37 VSS 0.0108f
C3203 a_10161_4198.n38 VSS 0.0292f
C3204 a_10161_4198.n39 VSS 0.0876f
C3205 a_10161_4198.t7 VSS 0.0108f
C3206 a_10161_4198.n40 VSS 0.0108f
C3207 a_10161_4198.n41 VSS 0.0217f
C3208 a_10161_4198.n42 VSS 0.0593f
C3209 a_10161_4198.n43 VSS 0.0939f
C3210 a_10161_4198.n44 VSS 0.043f
C3211 a_10161_4198.t38 VSS 0.0108f
C3212 a_10161_4198.n45 VSS 0.0108f
C3213 a_10161_4198.n46 VSS 0.0217f
C3214 a_10161_4198.t17 VSS 0.0108f
C3215 a_10161_4198.n47 VSS 0.0108f
C3216 a_10161_4198.n48 VSS 0.0217f
C3217 a_10161_4198.t25 VSS 0.0108f
C3218 a_10161_4198.n49 VSS 0.0108f
C3219 a_10161_4198.n50 VSS 0.0273f
C3220 a_10161_4198.t39 VSS 0.0108f
C3221 a_10161_4198.n51 VSS 0.0108f
C3222 a_10161_4198.n52 VSS 0.0217f
C3223 a_10161_4198.n53 VSS 0.0602f
C3224 a_10161_4198.t41 VSS 0.0108f
C3225 a_10161_4198.n54 VSS 0.0108f
C3226 a_10161_4198.n55 VSS 0.0217f
C3227 a_10161_4198.n56 VSS 0.386f
C3228 a_10161_4198.n57 VSS 0.128f
C3229 a_10161_4198.n58 VSS 0.175f
C3230 a_10161_4198.n59 VSS 0.525f
C3231 a_10161_4198.t51 VSS 0.0108f
C3232 a_10161_4198.n60 VSS 0.0108f
C3233 a_10161_4198.n61 VSS 0.0217f
C3234 a_10161_4198.t37 VSS 0.0108f
C3235 a_10161_4198.n62 VSS 0.0108f
C3236 a_10161_4198.n63 VSS 0.0217f
C3237 a_10161_4198.n64 VSS 0.065f
C3238 a_10161_4198.n65 VSS 0.0716f
C3239 a_10161_4198.n66 VSS 0.53f
C3240 a_10161_4198.t47 VSS 0.0108f
C3241 a_10161_4198.n67 VSS 0.0108f
C3242 a_10161_4198.n68 VSS 0.0217f
C3243 a_10161_4198.t49 VSS 0.0108f
C3244 a_10161_4198.n69 VSS 0.0108f
C3245 a_10161_4198.n70 VSS 0.0217f
C3246 a_10161_4198.t45 VSS 0.0108f
C3247 a_10161_4198.n71 VSS 0.0108f
C3248 a_10161_4198.n72 VSS 0.0217f
C3249 a_10161_4198.n73 VSS 0.0531f
C3250 a_10161_4198.n74 VSS 0.0533f
C3251 a_10161_4198.n75 VSS 0.0904f
C3252 a_10161_4198.t9 VSS 0.0108f
C3253 a_10161_4198.n76 VSS 0.0108f
C3254 a_10161_4198.n77 VSS 0.0217f
C3255 a_10161_4198.t59 VSS 0.0108f
C3256 a_10161_4198.n78 VSS 0.0108f
C3257 a_10161_4198.n79 VSS 0.0217f
C3258 a_10161_4198.t11 VSS 0.0108f
C3259 a_10161_4198.n80 VSS 0.0108f
C3260 a_10161_4198.n81 VSS 0.0217f
C3261 a_10161_4198.n82 VSS 0.106f
C3262 a_10161_4198.n83 VSS 0.0904f
C3263 a_10161_4198.t50 VSS 0.0108f
C3264 a_10161_4198.n84 VSS 0.0108f
C3265 a_10161_4198.n85 VSS 0.0217f
C3266 a_10161_4198.n86 VSS 0.107f
C3267 a_10161_4198.n87 VSS 0.0904f
C3268 a_10161_4198.n88 VSS 0.0531f
C3269 a_10161_4198.n89 VSS 0.0533f
C3270 a_10161_4198.n90 VSS 0.0904f
C3271 a_10161_4198.n91 VSS 0.065f
C3272 a_10161_4198.n92 VSS 0.0762f
C3273 a_10161_4198.n93 VSS 0.0217f
C3274 a_10161_4198.n94 VSS 0.0108f
C3275 VCO_C_0.INV_2_2.IN.n0 VSS 1.78f
C3276 VCO_C_0.INV_2_2.IN.n1 VSS 0.624f
C3277 VCO_C_0.INV_2_2.IN.n2 VSS 0.495f
C3278 VCO_C_0.INV_2_2.IN.n3 VSS 0.636f
C3279 VCO_C_0.INV_2_2.IN.n4 VSS 0.579f
C3280 VCO_C_0.INV_2_2.IN.n5 VSS 0.495f
C3281 VCO_C_0.INV_2_2.IN.n6 VSS 0.117f
C3282 VCO_C_0.INV_2_2.IN.n7 VSS 0.451f
C3283 VCO_C_0.INV_2_2.IN.t20 VSS 0.0531f
C3284 VCO_C_0.INV_2_2.IN.n8 VSS 0.0147f
C3285 VCO_C_0.INV_2_2.IN.t18 VSS 0.0174f
C3286 VCO_C_0.INV_2_2.IN.n9 VSS 0.0648f
C3287 VCO_C_0.INV_2_2.IN.n10 VSS 0.102f
C3288 VCO_C_0.INV_2_2.IN.t19 VSS 0.0915f
C3289 VCO_C_0.INV_2_2.IN.n11 VSS 0.0572f
C3290 VCO_C_0.INV_2_2.IN.n12 VSS 0.0147f
C3291 VCO_C_0.INV_2_2.IN.t22 VSS 0.0174f
C3292 VCO_C_0.INV_2_2.IN.n13 VSS 0.104f
C3293 VCO_C_0.INV_2_2.IN.n14 VSS 0.519f
C3294 VCO_C_0.INV_2_2.IN.n15 VSS 0.0147f
C3295 VCO_C_0.INV_2_2.IN.t21 VSS 0.0174f
C3296 VCO_C_0.INV_2_2.IN.n16 VSS 0.0579f
C3297 VCO_C_0.INV_2_2.IN.n17 VSS 0.447f
C3298 VCO_C_0.INV_2_2.IN.n18 VSS 0.312f
C3299 VCO_C_0.INV_2_2.IN.t40 VSS 0.108f
C3300 VCO_C_0.INV_2_2.IN.t53 VSS 0.111f
C3301 VCO_C_0.INV_2_2.IN.t32 VSS 0.108f
C3302 VCO_C_0.INV_2_2.IN.t46 VSS 0.111f
C3303 VCO_C_0.INV_2_2.IN.t43 VSS 0.113f
C3304 VCO_C_0.INV_2_2.IN.t57 VSS 0.109f
C3305 VCO_C_0.INV_2_2.IN.t33 VSS 0.109f
C3306 VCO_C_0.INV_2_2.IN.t47 VSS 0.109f
C3307 VCO_C_0.INV_2_2.IN.t31 VSS 0.109f
C3308 VCO_C_0.INV_2_2.IN.t34 VSS 0.109f
C3309 VCO_C_0.INV_2_2.IN.t35 VSS 0.11f
C3310 VCO_C_0.INV_2_2.IN.t39 VSS 0.149f
C3311 VCO_C_0.INV_2_2.IN.n19 VSS 0.811f
C3312 VCO_C_0.INV_2_2.IN.n20 VSS 0.367f
C3313 VCO_C_0.INV_2_2.IN.n21 VSS 0.49f
C3314 VCO_C_0.INV_2_2.IN.t48 VSS 0.114f
C3315 VCO_C_0.INV_2_2.IN.t49 VSS 0.114f
C3316 VCO_C_0.INV_2_2.IN.t51 VSS 0.111f
C3317 VCO_C_0.INV_2_2.IN.t54 VSS 0.148f
C3318 VCO_C_0.INV_2_2.IN.n22 VSS 0.832f
C3319 VCO_C_0.INV_2_2.IN.n23 VSS 0.383f
C3320 VCO_C_0.INV_2_2.IN.n24 VSS 0.505f
C3321 VCO_C_0.INV_2_2.IN.n25 VSS 0.668f
C3322 VCO_C_0.INV_2_2.IN.t4 VSS 0.0236f
C3323 VCO_C_0.INV_2_2.IN.n26 VSS 0.0461f
C3324 VCO_C_0.INV_2_2.IN.n27 VSS 0.398f
C3325 VCO_C_0.INV_2_2.IN.t9 VSS 0.016f
C3326 VCO_C_0.INV_2_2.IN.n28 VSS 0.016f
C3327 VCO_C_0.INV_2_2.IN.n29 VSS 0.0322f
C3328 VCO_C_0.INV_2_2.IN.n30 VSS 0.0361f
C3329 VCO_C_0.INV_2_2.IN.n31 VSS 0.0259f
C3330 VCO_C_0.INV_2_2.IN.n32 VSS 0.0869f
C3331 VCO_C_0.INV_2_2.IN.n33 VSS 0.265f
C3332 VCO_C_0.INV_2_2.IN.n34 VSS 0.0461f
C3333 VCO_C_0.INV_2_2.IN.n35 VSS 0.672f
C3334 VCO_C_0.INV_2_2.IN.t6 VSS 0.0259f
C3335 VCO_C_0.INV_2_2.IN.n36 VSS 0.0647f
C3336 VCO_C_0.INV_2_2.IN.t7 VSS 0.016f
C3337 VCO_C_0.INV_2_2.IN.n37 VSS 0.016f
C3338 VCO_C_0.INV_2_2.IN.n38 VSS 0.154f
C3339 VCO_C_0.INV_2_2.IN.n39 VSS 0.123f
C3340 VCO_C_0.INV_2_2.IN.t13 VSS 0.0237f
C3341 VCO_C_0.INV_2_2.IN.n40 VSS 0.116f
C3342 VCO_C_0.INV_2_2.IN.n41 VSS 0.175f
C3343 VCO_C_0.INV_2_2.IN.t28 VSS 0.016f
C3344 VCO_C_0.INV_2_2.IN.n42 VSS 0.016f
C3345 VCO_C_0.INV_2_2.IN.n43 VSS 0.0321f
C3346 VCO_C_0.INV_2_2.IN.n44 VSS 0.0626f
C3347 VCO_C_0.INV_2_2.IN.n45 VSS 0.315f
C3348 VCO_C_0.INV_2_2.IN.t1 VSS 0.0279f
C3349 VCO_C_0.INV_2_2.IN.n46 VSS 0.0832f
C3350 VCO_C_0.INV_2_2.IN.n47 VSS 0.246f
C3351 VCO_C_0.INV_2_2.IN.n48 VSS 0.0574f
C3352 VCO_C_0.INV_2_2.IN.n49 VSS 0.47f
C3353 VCO_C_0.INV_2_2.IN.t8 VSS 0.016f
C3354 VCO_C_0.INV_2_2.IN.n50 VSS 0.016f
C3355 VCO_C_0.INV_2_2.IN.n51 VSS 0.0322f
C3356 VCO_C_0.INV_2_2.IN.n52 VSS 0.136f
C3357 VCO_C_0.INV_2_2.IN.n53 VSS 0.025f
C3358 VCO_C_0.INV_2_2.IN.n54 VSS 0.58f
C3359 VCO_C_0.INV_2_2.IN.n55 VSS 0.319f
C3360 VCO_C_0.INV_2_2.IN.n56 VSS 0.468f
C3361 VCO_C_0.INV_2_2.IN.t14 VSS 0.034f
C3362 VCO_C_0.INV_2_2.IN.t15 VSS 0.016f
C3363 VCO_C_0.INV_2_2.IN.n57 VSS 0.016f
C3364 VCO_C_0.INV_2_2.IN.n58 VSS 0.0772f
C3365 VCO_C_0.INV_2_2.IN.n59 VSS 0.0373f
C3366 VCO_C_0.INV_2_2.IN.n60 VSS 0.0938f
C3367 VCO_C_0.INV_2_2.IN.n61 VSS 0.5f
C3368 VCO_C_0.INV_2_2.IN.n62 VSS 0.344f
C3369 VCO_C_0.INV_2_2.IN.n63 VSS 2.19f
C3370 VCO_C_0.INV_2_2.IN.t36 VSS 0.129f
C3371 VCO_C_0.INV_2_2.IN.t50 VSS 0.0981f
C3372 VCO_C_0.INV_2_2.IN.n64 VSS 0.0927f
C3373 VCO_C_0.INV_2_2.IN.n65 VSS 0.142f
C3374 VCO_C_0.INV_2_2.IN.t58 VSS 0.053f
C3375 VCO_C_0.INV_2_2.IN.n66 VSS 0.113f
C3376 VCO_C_0.INV_2_2.IN.n67 VSS 0.142f
C3377 VCO_C_0.INV_2_2.IN.t44 VSS 0.053f
C3378 VCO_C_0.INV_2_2.IN.n68 VSS 0.113f
C3379 VCO_C_0.INV_2_2.IN.t56 VSS 0.129f
C3380 VCO_C_0.INV_2_2.IN.n69 VSS 0.0927f
C3381 VCO_C_0.INV_2_2.IN.t41 VSS 0.0845f
C3382 VCO_C_0.INV_2_2.IN.t45 VSS 0.0401f
C3383 VCO_C_0.INV_2_2.IN.n70 VSS 0.115f
C3384 VCO_C_0.INV_2_2.IN.t42 VSS 0.0981f
C3385 VCO_C_0.INV_2_2.IN.t38 VSS 0.0401f
C3386 VCO_C_0.INV_2_2.IN.n71 VSS 0.13f
C3387 VCO_C_0.INV_2_2.IN.t55 VSS 0.0981f
C3388 VCO_C_0.INV_2_2.IN.t52 VSS 0.0401f
C3389 VCO_C_0.INV_2_2.IN.n72 VSS 0.13f
C3390 VCO_C_0.INV_2_2.IN.t37 VSS 0.04f
C3391 VCO_C_0.INV_2_2.IN.n73 VSS 0.0657f
C3392 VCO_C_0.INV_2_2.IN.n74 VSS 0.0664f
C3393 VCO_C_0.INV_2_2.IN.n75 VSS 0.0697f
.ends

