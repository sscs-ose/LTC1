magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2558 -2501 2558 2501
<< psubdiff >>
rect -558 479 558 501
rect -558 433 -536 479
rect -490 433 -422 479
rect -376 433 -308 479
rect -262 433 -194 479
rect -148 433 -80 479
rect -34 433 34 479
rect 80 433 148 479
rect 194 433 262 479
rect 308 433 376 479
rect 422 433 490 479
rect 536 433 558 479
rect -558 365 558 433
rect -558 319 -536 365
rect -490 319 -422 365
rect -376 319 -308 365
rect -262 319 -194 365
rect -148 319 -80 365
rect -34 319 34 365
rect 80 319 148 365
rect 194 319 262 365
rect 308 319 376 365
rect 422 319 490 365
rect 536 319 558 365
rect -558 251 558 319
rect -558 205 -536 251
rect -490 205 -422 251
rect -376 205 -308 251
rect -262 205 -194 251
rect -148 205 -80 251
rect -34 205 34 251
rect 80 205 148 251
rect 194 205 262 251
rect 308 205 376 251
rect 422 205 490 251
rect 536 205 558 251
rect -558 137 558 205
rect -558 91 -536 137
rect -490 91 -422 137
rect -376 91 -308 137
rect -262 91 -194 137
rect -148 91 -80 137
rect -34 91 34 137
rect 80 91 148 137
rect 194 91 262 137
rect 308 91 376 137
rect 422 91 490 137
rect 536 91 558 137
rect -558 23 558 91
rect -558 -23 -536 23
rect -490 -23 -422 23
rect -376 -23 -308 23
rect -262 -23 -194 23
rect -148 -23 -80 23
rect -34 -23 34 23
rect 80 -23 148 23
rect 194 -23 262 23
rect 308 -23 376 23
rect 422 -23 490 23
rect 536 -23 558 23
rect -558 -91 558 -23
rect -558 -137 -536 -91
rect -490 -137 -422 -91
rect -376 -137 -308 -91
rect -262 -137 -194 -91
rect -148 -137 -80 -91
rect -34 -137 34 -91
rect 80 -137 148 -91
rect 194 -137 262 -91
rect 308 -137 376 -91
rect 422 -137 490 -91
rect 536 -137 558 -91
rect -558 -205 558 -137
rect -558 -251 -536 -205
rect -490 -251 -422 -205
rect -376 -251 -308 -205
rect -262 -251 -194 -205
rect -148 -251 -80 -205
rect -34 -251 34 -205
rect 80 -251 148 -205
rect 194 -251 262 -205
rect 308 -251 376 -205
rect 422 -251 490 -205
rect 536 -251 558 -205
rect -558 -319 558 -251
rect -558 -365 -536 -319
rect -490 -365 -422 -319
rect -376 -365 -308 -319
rect -262 -365 -194 -319
rect -148 -365 -80 -319
rect -34 -365 34 -319
rect 80 -365 148 -319
rect 194 -365 262 -319
rect 308 -365 376 -319
rect 422 -365 490 -319
rect 536 -365 558 -319
rect -558 -433 558 -365
rect -558 -479 -536 -433
rect -490 -479 -422 -433
rect -376 -479 -308 -433
rect -262 -479 -194 -433
rect -148 -479 -80 -433
rect -34 -479 34 -433
rect 80 -479 148 -433
rect 194 -479 262 -433
rect 308 -479 376 -433
rect 422 -479 490 -433
rect 536 -479 558 -433
rect -558 -501 558 -479
<< psubdiffcont >>
rect -536 433 -490 479
rect -422 433 -376 479
rect -308 433 -262 479
rect -194 433 -148 479
rect -80 433 -34 479
rect 34 433 80 479
rect 148 433 194 479
rect 262 433 308 479
rect 376 433 422 479
rect 490 433 536 479
rect -536 319 -490 365
rect -422 319 -376 365
rect -308 319 -262 365
rect -194 319 -148 365
rect -80 319 -34 365
rect 34 319 80 365
rect 148 319 194 365
rect 262 319 308 365
rect 376 319 422 365
rect 490 319 536 365
rect -536 205 -490 251
rect -422 205 -376 251
rect -308 205 -262 251
rect -194 205 -148 251
rect -80 205 -34 251
rect 34 205 80 251
rect 148 205 194 251
rect 262 205 308 251
rect 376 205 422 251
rect 490 205 536 251
rect -536 91 -490 137
rect -422 91 -376 137
rect -308 91 -262 137
rect -194 91 -148 137
rect -80 91 -34 137
rect 34 91 80 137
rect 148 91 194 137
rect 262 91 308 137
rect 376 91 422 137
rect 490 91 536 137
rect -536 -23 -490 23
rect -422 -23 -376 23
rect -308 -23 -262 23
rect -194 -23 -148 23
rect -80 -23 -34 23
rect 34 -23 80 23
rect 148 -23 194 23
rect 262 -23 308 23
rect 376 -23 422 23
rect 490 -23 536 23
rect -536 -137 -490 -91
rect -422 -137 -376 -91
rect -308 -137 -262 -91
rect -194 -137 -148 -91
rect -80 -137 -34 -91
rect 34 -137 80 -91
rect 148 -137 194 -91
rect 262 -137 308 -91
rect 376 -137 422 -91
rect 490 -137 536 -91
rect -536 -251 -490 -205
rect -422 -251 -376 -205
rect -308 -251 -262 -205
rect -194 -251 -148 -205
rect -80 -251 -34 -205
rect 34 -251 80 -205
rect 148 -251 194 -205
rect 262 -251 308 -205
rect 376 -251 422 -205
rect 490 -251 536 -205
rect -536 -365 -490 -319
rect -422 -365 -376 -319
rect -308 -365 -262 -319
rect -194 -365 -148 -319
rect -80 -365 -34 -319
rect 34 -365 80 -319
rect 148 -365 194 -319
rect 262 -365 308 -319
rect 376 -365 422 -319
rect 490 -365 536 -319
rect -536 -479 -490 -433
rect -422 -479 -376 -433
rect -308 -479 -262 -433
rect -194 -479 -148 -433
rect -80 -479 -34 -433
rect 34 -479 80 -433
rect 148 -479 194 -433
rect 262 -479 308 -433
rect 376 -479 422 -433
rect 490 -479 536 -433
<< metal1 >>
rect -547 479 547 490
rect -547 433 -536 479
rect -490 433 -422 479
rect -376 433 -308 479
rect -262 433 -194 479
rect -148 433 -80 479
rect -34 433 34 479
rect 80 433 148 479
rect 194 433 262 479
rect 308 433 376 479
rect 422 433 490 479
rect 536 433 547 479
rect -547 365 547 433
rect -547 319 -536 365
rect -490 319 -422 365
rect -376 319 -308 365
rect -262 319 -194 365
rect -148 319 -80 365
rect -34 319 34 365
rect 80 319 148 365
rect 194 319 262 365
rect 308 319 376 365
rect 422 319 490 365
rect 536 319 547 365
rect -547 251 547 319
rect -547 205 -536 251
rect -490 205 -422 251
rect -376 205 -308 251
rect -262 205 -194 251
rect -148 205 -80 251
rect -34 205 34 251
rect 80 205 148 251
rect 194 205 262 251
rect 308 205 376 251
rect 422 205 490 251
rect 536 205 547 251
rect -547 137 547 205
rect -547 91 -536 137
rect -490 91 -422 137
rect -376 91 -308 137
rect -262 91 -194 137
rect -148 91 -80 137
rect -34 91 34 137
rect 80 91 148 137
rect 194 91 262 137
rect 308 91 376 137
rect 422 91 490 137
rect 536 91 547 137
rect -547 23 547 91
rect -547 -23 -536 23
rect -490 -23 -422 23
rect -376 -23 -308 23
rect -262 -23 -194 23
rect -148 -23 -80 23
rect -34 -23 34 23
rect 80 -23 148 23
rect 194 -23 262 23
rect 308 -23 376 23
rect 422 -23 490 23
rect 536 -23 547 23
rect -547 -91 547 -23
rect -547 -137 -536 -91
rect -490 -137 -422 -91
rect -376 -137 -308 -91
rect -262 -137 -194 -91
rect -148 -137 -80 -91
rect -34 -137 34 -91
rect 80 -137 148 -91
rect 194 -137 262 -91
rect 308 -137 376 -91
rect 422 -137 490 -91
rect 536 -137 547 -91
rect -547 -205 547 -137
rect -547 -251 -536 -205
rect -490 -251 -422 -205
rect -376 -251 -308 -205
rect -262 -251 -194 -205
rect -148 -251 -80 -205
rect -34 -251 34 -205
rect 80 -251 148 -205
rect 194 -251 262 -205
rect 308 -251 376 -205
rect 422 -251 490 -205
rect 536 -251 547 -205
rect -547 -319 547 -251
rect -547 -365 -536 -319
rect -490 -365 -422 -319
rect -376 -365 -308 -319
rect -262 -365 -194 -319
rect -148 -365 -80 -319
rect -34 -365 34 -319
rect 80 -365 148 -319
rect 194 -365 262 -319
rect 308 -365 376 -319
rect 422 -365 490 -319
rect 536 -365 547 -319
rect -547 -433 547 -365
rect -547 -479 -536 -433
rect -490 -479 -422 -433
rect -376 -479 -308 -433
rect -262 -479 -194 -433
rect -148 -479 -80 -433
rect -34 -479 34 -433
rect 80 -479 148 -433
rect 194 -479 262 -433
rect 308 -479 376 -433
rect 422 -479 490 -433
rect 536 -479 547 -433
rect -547 -490 547 -479
<< end >>
