magic
tech gf180mcuC
magscale 1 10
timestamp 1699896181
<< nwell >>
rect -260 1850 2668 2179
rect -260 -60 -60 1850
rect 1721 1802 1751 1850
rect 1499 -60 2059 68
rect 2468 -60 2668 1850
rect -260 -260 2668 -60
<< nsubdiff >>
rect -210 2107 2618 2124
rect -210 2061 -193 2107
rect -147 2061 -95 2107
rect -48 2061 4 2107
rect 50 2061 102 2107
rect 148 2061 200 2107
rect 246 2061 298 2107
rect 344 2061 396 2107
rect 442 2061 494 2107
rect 540 2061 592 2107
rect 638 2061 690 2107
rect 736 2061 788 2107
rect 834 2061 886 2107
rect 932 2061 984 2107
rect 1030 2061 1082 2107
rect 1128 2061 1180 2107
rect 1226 2061 1278 2107
rect 1324 2061 1376 2107
rect 1422 2061 1474 2107
rect 1520 2061 1572 2107
rect 1618 2061 1670 2107
rect 1716 2061 1768 2107
rect 1814 2061 1866 2107
rect 1912 2061 1964 2107
rect 2010 2061 2062 2107
rect 2108 2061 2160 2107
rect 2206 2061 2258 2107
rect 2304 2061 2356 2107
rect 2402 2061 2454 2107
rect 2500 2061 2555 2107
rect 2601 2061 2618 2107
rect -210 2044 2618 2061
rect -210 2009 -130 2044
rect -210 1963 -193 2009
rect -147 1963 -130 2009
rect -210 1911 -130 1963
rect -210 1865 -193 1911
rect -147 1865 -130 1911
rect -210 1813 -130 1865
rect -210 1767 -193 1813
rect -147 1767 -130 1813
rect -210 1715 -130 1767
rect -210 1669 -193 1715
rect -147 1669 -130 1715
rect -210 1617 -130 1669
rect -210 1571 -193 1617
rect -147 1571 -130 1617
rect -210 1519 -130 1571
rect -210 1473 -193 1519
rect -147 1473 -130 1519
rect -210 1421 -130 1473
rect -210 1375 -193 1421
rect -147 1375 -130 1421
rect -210 1323 -130 1375
rect -210 1277 -193 1323
rect -147 1277 -130 1323
rect -210 1225 -130 1277
rect -210 1179 -193 1225
rect -147 1179 -130 1225
rect -210 1127 -130 1179
rect -210 1081 -193 1127
rect -147 1081 -130 1127
rect -210 1029 -130 1081
rect -210 983 -193 1029
rect -147 983 -130 1029
rect -210 931 -130 983
rect -210 885 -193 931
rect -147 885 -130 931
rect -210 833 -130 885
rect -210 787 -193 833
rect -147 787 -130 833
rect -210 735 -130 787
rect -210 689 -193 735
rect -147 689 -130 735
rect -210 637 -130 689
rect -210 591 -193 637
rect -147 591 -130 637
rect -210 539 -130 591
rect -210 493 -193 539
rect -147 493 -130 539
rect -210 441 -130 493
rect -210 395 -193 441
rect -147 395 -130 441
rect -210 343 -130 395
rect -210 297 -193 343
rect -147 297 -130 343
rect -210 245 -130 297
rect -210 199 -193 245
rect -147 199 -130 245
rect -210 147 -130 199
rect -210 101 -193 147
rect -147 101 -130 147
rect -210 49 -130 101
rect -210 3 -193 49
rect -147 3 -130 49
rect -210 -49 -130 3
rect -210 -95 -193 -49
rect -147 -95 -130 -49
rect -210 -130 -130 -95
rect 2538 2009 2618 2044
rect 2538 1963 2555 2009
rect 2601 1963 2618 2009
rect 2538 1911 2618 1963
rect 2538 1865 2555 1911
rect 2601 1865 2618 1911
rect 2538 1813 2618 1865
rect 2538 1767 2555 1813
rect 2601 1767 2618 1813
rect 2538 1715 2618 1767
rect 2538 1669 2555 1715
rect 2601 1669 2618 1715
rect 2538 1617 2618 1669
rect 2538 1571 2555 1617
rect 2601 1571 2618 1617
rect 2538 1519 2618 1571
rect 2538 1473 2555 1519
rect 2601 1473 2618 1519
rect 2538 1421 2618 1473
rect 2538 1375 2555 1421
rect 2601 1375 2618 1421
rect 2538 1323 2618 1375
rect 2538 1277 2555 1323
rect 2601 1277 2618 1323
rect 2538 1225 2618 1277
rect 2538 1179 2555 1225
rect 2601 1179 2618 1225
rect 2538 1127 2618 1179
rect 2538 1081 2555 1127
rect 2601 1081 2618 1127
rect 2538 1029 2618 1081
rect 2538 983 2555 1029
rect 2601 983 2618 1029
rect 2538 931 2618 983
rect 2538 885 2555 931
rect 2601 885 2618 931
rect 2538 833 2618 885
rect 2538 787 2555 833
rect 2601 787 2618 833
rect 2538 735 2618 787
rect 2538 689 2555 735
rect 2601 689 2618 735
rect 2538 637 2618 689
rect 2538 591 2555 637
rect 2601 591 2618 637
rect 2538 539 2618 591
rect 2538 493 2555 539
rect 2601 493 2618 539
rect 2538 441 2618 493
rect 2538 395 2555 441
rect 2601 395 2618 441
rect 2538 343 2618 395
rect 2538 297 2555 343
rect 2601 297 2618 343
rect 2538 245 2618 297
rect 2538 199 2555 245
rect 2601 199 2618 245
rect 2538 147 2618 199
rect 2538 101 2555 147
rect 2601 101 2618 147
rect 2538 49 2618 101
rect 2538 3 2555 49
rect 2601 3 2618 49
rect 2538 -49 2618 3
rect 2538 -95 2555 -49
rect 2601 -95 2618 -49
rect 2538 -130 2618 -95
rect -210 -147 2618 -130
rect -210 -193 -193 -147
rect -147 -193 -95 -147
rect -49 -193 3 -147
rect 49 -193 101 -147
rect 147 -193 199 -147
rect 245 -193 297 -147
rect 343 -193 395 -147
rect 441 -193 493 -147
rect 539 -193 591 -147
rect 637 -193 689 -147
rect 735 -193 787 -147
rect 833 -193 885 -147
rect 931 -193 983 -147
rect 1029 -193 1081 -147
rect 1127 -193 1179 -147
rect 1225 -193 1277 -147
rect 1323 -193 1375 -147
rect 1421 -193 1473 -147
rect 1519 -193 1571 -147
rect 1617 -193 1669 -147
rect 1715 -193 1767 -147
rect 1813 -193 1865 -147
rect 1911 -193 1963 -147
rect 2009 -193 2061 -147
rect 2107 -193 2159 -147
rect 2205 -193 2257 -147
rect 2303 -193 2355 -147
rect 2401 -193 2453 -147
rect 2499 -193 2551 -147
rect 2601 -193 2618 -147
rect -210 -210 2618 -193
<< nsubdiffcont >>
rect -193 2061 -147 2107
rect -95 2061 -48 2107
rect 4 2061 50 2107
rect 102 2061 148 2107
rect 200 2061 246 2107
rect 298 2061 344 2107
rect 396 2061 442 2107
rect 494 2061 540 2107
rect 592 2061 638 2107
rect 690 2061 736 2107
rect 788 2061 834 2107
rect 886 2061 932 2107
rect 984 2061 1030 2107
rect 1082 2061 1128 2107
rect 1180 2061 1226 2107
rect 1278 2061 1324 2107
rect 1376 2061 1422 2107
rect 1474 2061 1520 2107
rect 1572 2061 1618 2107
rect 1670 2061 1716 2107
rect 1768 2061 1814 2107
rect 1866 2061 1912 2107
rect 1964 2061 2010 2107
rect 2062 2061 2108 2107
rect 2160 2061 2206 2107
rect 2258 2061 2304 2107
rect 2356 2061 2402 2107
rect 2454 2061 2500 2107
rect 2555 2061 2601 2107
rect -193 1963 -147 2009
rect -193 1865 -147 1911
rect -193 1767 -147 1813
rect -193 1669 -147 1715
rect -193 1571 -147 1617
rect -193 1473 -147 1519
rect -193 1375 -147 1421
rect -193 1277 -147 1323
rect -193 1179 -147 1225
rect -193 1081 -147 1127
rect -193 983 -147 1029
rect -193 885 -147 931
rect -193 787 -147 833
rect -193 689 -147 735
rect -193 591 -147 637
rect -193 493 -147 539
rect -193 395 -147 441
rect -193 297 -147 343
rect -193 199 -147 245
rect -193 101 -147 147
rect -193 3 -147 49
rect -193 -95 -147 -49
rect 2555 1963 2601 2009
rect 2555 1865 2601 1911
rect 2555 1767 2601 1813
rect 2555 1669 2601 1715
rect 2555 1571 2601 1617
rect 2555 1473 2601 1519
rect 2555 1375 2601 1421
rect 2555 1277 2601 1323
rect 2555 1179 2601 1225
rect 2555 1081 2601 1127
rect 2555 983 2601 1029
rect 2555 885 2601 931
rect 2555 787 2601 833
rect 2555 689 2601 735
rect 2555 591 2601 637
rect 2555 493 2601 539
rect 2555 395 2601 441
rect 2555 297 2601 343
rect 2555 199 2601 245
rect 2555 101 2601 147
rect 2555 3 2601 49
rect 2555 -95 2601 -49
rect -193 -193 -147 -147
rect -95 -193 -49 -147
rect 3 -193 49 -147
rect 101 -193 147 -147
rect 199 -193 245 -147
rect 297 -193 343 -147
rect 395 -193 441 -147
rect 493 -193 539 -147
rect 591 -193 637 -147
rect 689 -193 735 -147
rect 787 -193 833 -147
rect 885 -193 931 -147
rect 983 -193 1029 -147
rect 1081 -193 1127 -147
rect 1179 -193 1225 -147
rect 1277 -193 1323 -147
rect 1375 -193 1421 -147
rect 1473 -193 1519 -147
rect 1571 -193 1617 -147
rect 1669 -193 1715 -147
rect 1767 -193 1813 -147
rect 1865 -193 1911 -147
rect 1963 -193 2009 -147
rect 2061 -193 2107 -147
rect 2159 -193 2205 -147
rect 2257 -193 2303 -147
rect 2355 -193 2401 -147
rect 2453 -193 2499 -147
rect 2551 -193 2601 -147
<< metal1 >>
rect -210 2107 2618 2124
rect -210 2061 -193 2107
rect -147 2061 -95 2107
rect -48 2061 4 2107
rect 50 2061 102 2107
rect 148 2061 200 2107
rect 246 2061 298 2107
rect 344 2061 396 2107
rect 442 2061 494 2107
rect 540 2061 592 2107
rect 638 2061 690 2107
rect 736 2061 788 2107
rect 834 2061 886 2107
rect 932 2061 984 2107
rect 1030 2061 1082 2107
rect 1128 2061 1180 2107
rect 1226 2061 1278 2107
rect 1324 2061 1376 2107
rect 1422 2061 1474 2107
rect 1520 2061 1572 2107
rect 1618 2061 1670 2107
rect 1716 2061 1768 2107
rect 1814 2061 1866 2107
rect 1912 2061 1964 2107
rect 2010 2061 2062 2107
rect 2108 2061 2160 2107
rect 2206 2061 2258 2107
rect 2304 2061 2356 2107
rect 2402 2061 2454 2107
rect 2500 2061 2555 2107
rect 2601 2061 2618 2107
rect -210 2044 2618 2061
rect -210 2009 -130 2044
rect -210 1963 -193 2009
rect -147 1963 -130 2009
rect -210 1911 -130 1963
rect -210 1865 -193 1911
rect -147 1865 -130 1911
rect -210 1813 -130 1865
rect -210 1767 -193 1813
rect -147 1767 -130 1813
rect -210 1715 -130 1767
rect -210 1669 -193 1715
rect -147 1669 -130 1715
rect 127 1671 321 2044
rect 408 1670 602 2044
rect 975 1964 1721 1965
rect 966 1804 1721 1964
rect -210 1617 -130 1669
rect -210 1571 -193 1617
rect -147 1571 -130 1617
rect -210 1519 -130 1571
rect -210 1473 -193 1519
rect -147 1473 -130 1519
rect -210 1421 -130 1473
rect 687 1464 881 1716
rect 966 1668 1162 1804
rect -210 1375 -193 1421
rect -147 1375 -130 1421
rect -210 1323 -130 1375
rect -210 1277 -193 1323
rect -147 1277 -130 1323
rect -210 1225 -130 1277
rect 143 1270 881 1464
rect 1247 1587 1443 1723
rect 1525 1668 1721 1804
rect 1806 1722 2002 1723
rect 1806 1676 2003 1722
rect 1806 1587 2002 1676
rect 2088 1668 2282 2044
rect 2538 2009 2618 2044
rect 2538 1963 2555 2009
rect 2601 1963 2618 2009
rect 2538 1911 2618 1963
rect 2538 1865 2555 1911
rect 2601 1865 2618 1911
rect 2538 1813 2618 1865
rect 2538 1767 2555 1813
rect 2601 1767 2618 1813
rect 2538 1715 2618 1767
rect 2538 1669 2555 1715
rect 2601 1669 2618 1715
rect 1247 1427 2002 1587
rect 1256 1426 2002 1427
rect 2538 1617 2618 1669
rect 2538 1571 2555 1617
rect 2601 1571 2618 1617
rect 2538 1519 2618 1571
rect 2538 1473 2555 1519
rect 2601 1473 2618 1519
rect 2538 1421 2618 1473
rect 2538 1375 2555 1421
rect 2601 1375 2618 1421
rect 2538 1323 2618 1375
rect 2538 1277 2555 1323
rect 2601 1277 2618 1323
rect -210 1179 -193 1225
rect -147 1179 -130 1225
rect -210 1127 -130 1179
rect -210 1081 -193 1127
rect -147 1081 -130 1127
rect -210 1029 -130 1081
rect -210 983 -193 1029
rect -147 983 -130 1029
rect -210 931 -130 983
rect -210 885 -193 931
rect -147 885 -130 931
rect -210 833 -130 885
rect -210 787 -193 833
rect -147 787 -130 833
rect -210 735 -130 787
rect -210 689 -193 735
rect -147 689 -130 735
rect -210 637 -130 689
rect -210 591 -193 637
rect -147 591 -130 637
rect -210 539 -130 591
rect -210 493 -193 539
rect -147 493 -130 539
rect -210 441 -130 493
rect -210 395 -193 441
rect -147 395 -130 441
rect 2538 1225 2618 1277
rect 2538 1179 2555 1225
rect 2601 1179 2618 1225
rect 2538 1127 2618 1179
rect 2538 1081 2555 1127
rect 2601 1081 2618 1127
rect 2538 1029 2618 1081
rect 2538 983 2555 1029
rect 2601 983 2618 1029
rect 2538 931 2618 983
rect 2538 885 2555 931
rect 2601 885 2618 931
rect 2538 833 2618 885
rect 2538 787 2555 833
rect 2601 787 2618 833
rect 2538 735 2618 787
rect 2538 689 2555 735
rect 2601 689 2618 735
rect 2538 637 2618 689
rect 2538 591 2555 637
rect 2601 591 2618 637
rect 2538 539 2618 591
rect 2538 493 2555 539
rect 2601 493 2618 539
rect 2538 441 2618 493
rect 698 432 1444 433
rect -210 343 -130 395
rect -210 297 -193 343
rect -147 297 -130 343
rect -210 245 -130 297
rect -210 199 -193 245
rect -147 199 -130 245
rect -210 147 -130 199
rect 689 272 1444 432
rect -210 101 -193 147
rect -147 101 -130 147
rect -210 49 -130 101
rect -210 3 -193 49
rect -147 3 -130 49
rect -210 -49 -130 3
rect -210 -95 -193 -49
rect -147 -95 -130 -49
rect -210 -130 -130 -95
rect 126 -130 320 187
rect 406 77 603 185
rect 689 136 885 272
rect 967 77 1164 186
rect 1248 183 1444 272
rect 2538 395 2555 441
rect 2601 395 2618 441
rect 2538 343 2618 395
rect 2538 297 2555 343
rect 2601 297 2618 343
rect 2538 245 2618 297
rect 1248 137 1445 183
rect 1248 136 1444 137
rect 406 -84 1164 77
rect 1525 68 2003 228
rect 2538 199 2555 245
rect 2601 199 2618 245
rect 2084 -130 2278 185
rect 2538 147 2618 199
rect 2538 101 2555 147
rect 2601 101 2618 147
rect 2538 49 2618 101
rect 2538 3 2555 49
rect 2601 3 2618 49
rect 2538 -49 2618 3
rect 2538 -95 2555 -49
rect 2601 -95 2618 -49
rect 2538 -130 2618 -95
rect -210 -147 2618 -130
rect -210 -193 -193 -147
rect -147 -193 -95 -147
rect -49 -193 3 -147
rect 49 -193 101 -147
rect 147 -193 199 -147
rect 245 -193 297 -147
rect 343 -193 395 -147
rect 441 -193 493 -147
rect 539 -193 591 -147
rect 637 -193 689 -147
rect 735 -193 787 -147
rect 833 -193 885 -147
rect 931 -193 983 -147
rect 1029 -193 1081 -147
rect 1127 -193 1179 -147
rect 1225 -193 1277 -147
rect 1323 -193 1375 -147
rect 1421 -193 1473 -147
rect 1519 -193 1571 -147
rect 1617 -193 1669 -147
rect 1715 -193 1767 -147
rect 1813 -193 1865 -147
rect 1911 -193 1963 -147
rect 2009 -193 2061 -147
rect 2107 -193 2159 -147
rect 2205 -193 2257 -147
rect 2303 -193 2355 -147
rect 2401 -193 2453 -147
rect 2499 -193 2551 -147
rect 2601 -193 2618 -147
rect -210 -210 2618 -193
use ppolyf_u_PVCJS8  ppolyf_u_PVCJS8_0
timestamp 1699895628
transform 1 0 1204 0 1 926
box -1264 -986 1264 986
<< labels >>
flabel metal1 493 1958 493 1958 0 FreeSans 1600 0 0 0 VDD
port 0 nsew
flabel metal1 312 1363 312 1363 0 FreeSans 1600 0 0 0 VSS
port 1 nsew
flabel metal1 1779 108 1779 108 0 FreeSans 800 0 0 0 VCM_1.6
port 3 nsew
<< end >>
