magic
tech gf180mcuC
magscale 1 10
timestamp 1693455138
<< mimcap >>
rect -20427 20100 -427 20180
rect -20427 260 -20347 20100
rect -507 260 -427 20100
rect -20427 180 -427 260
rect 187 20100 20187 20180
rect 187 260 267 20100
rect 20107 260 20187 20100
rect 187 180 20187 260
rect -20427 -260 -427 -180
rect -20427 -20100 -20347 -260
rect -507 -20100 -427 -260
rect -20427 -20180 -427 -20100
rect 187 -260 20187 -180
rect 187 -20100 267 -260
rect 20107 -20100 20187 -260
rect 187 -20180 20187 -20100
<< mimcapcontact >>
rect -20347 260 -507 20100
rect 267 260 20107 20100
rect -20347 -20100 -507 -260
rect 267 -20100 20107 -260
<< metal4 >>
rect -20547 20233 -67 20300
rect -20547 20180 -217 20233
rect -20547 180 -20427 20180
rect -427 180 -217 20180
rect -20547 127 -217 180
rect -129 127 -67 20233
rect -20547 60 -67 127
rect 67 20233 20547 20300
rect 67 20180 20397 20233
rect 67 180 187 20180
rect 20187 180 20397 20180
rect 67 127 20397 180
rect 20485 127 20547 20233
rect 67 60 20547 127
rect -20547 -127 -67 -60
rect -20547 -180 -217 -127
rect -20547 -20180 -20427 -180
rect -427 -20180 -217 -180
rect -20547 -20233 -217 -20180
rect -129 -20233 -67 -127
rect -20547 -20300 -67 -20233
rect 67 -127 20547 -60
rect 67 -180 20397 -127
rect 67 -20180 187 -180
rect 20187 -20180 20397 -180
rect 67 -20233 20397 -20180
rect 20485 -20233 20547 -127
rect 67 -20300 20547 -20233
<< via4 >>
rect -217 127 -129 20233
rect 20397 127 20485 20233
rect -217 -20233 -129 -127
rect 20397 -20233 20485 -127
<< metal5 >>
rect -217 20233 -129 20243
rect 20397 20233 20485 20243
rect -217 117 -129 127
rect 20397 117 20485 127
rect -217 -127 -129 -117
rect 20397 -127 20485 -117
rect -217 -20243 -129 -20233
rect 20397 -20243 20485 -20233
<< properties >>
string FIXED_BBOX 67 60 20307 20300
string gencell mim_2p0fF
string library gf180mcu
string parameters w 100.0 l 100.0 val 258.0k carea 25.00 cperi 20.00 nx 2 ny 2 dummy 0 square 0 lmin 5.00 wmin 5.00 lmax 100.0 wmax 100.0 dc 0 bconnect 0 tconnect 0
<< end >>
