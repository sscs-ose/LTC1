magic
tech gf180mcuC
magscale 1 10
timestamp 1691670594
<< nwell >>
rect -64 794 1692 1032
rect 804 340 1688 794
<< pwell >>
rect 864 0 1624 236
<< nmos >>
rect 976 68 1032 168
rect 1136 68 1192 168
rect 1296 68 1352 168
rect 1456 68 1512 168
<< pmos >>
rect 978 470 1034 670
rect 1138 470 1194 670
rect 1298 470 1354 670
rect 1458 470 1514 670
<< ndiff >>
rect 888 155 976 168
rect 888 81 901 155
rect 947 81 976 155
rect 888 68 976 81
rect 1032 155 1136 168
rect 1032 81 1061 155
rect 1107 81 1136 155
rect 1032 68 1136 81
rect 1192 155 1296 168
rect 1192 81 1221 155
rect 1267 81 1296 155
rect 1192 68 1296 81
rect 1352 155 1456 168
rect 1352 81 1381 155
rect 1427 81 1456 155
rect 1352 68 1456 81
rect 1512 155 1600 168
rect 1512 81 1541 155
rect 1587 81 1600 155
rect 1512 68 1600 81
<< pdiff >>
rect 890 657 978 670
rect 890 483 903 657
rect 949 483 978 657
rect 890 470 978 483
rect 1034 657 1138 670
rect 1034 483 1063 657
rect 1109 483 1138 657
rect 1034 470 1138 483
rect 1194 657 1298 670
rect 1194 483 1223 657
rect 1269 483 1298 657
rect 1194 470 1298 483
rect 1354 657 1458 670
rect 1354 483 1383 657
rect 1429 483 1458 657
rect 1354 470 1458 483
rect 1514 657 1602 670
rect 1514 483 1543 657
rect 1589 483 1602 657
rect 1514 470 1602 483
<< ndiffc >>
rect 901 81 947 155
rect 1061 81 1107 155
rect 1221 81 1267 155
rect 1381 81 1427 155
rect 1541 81 1587 155
<< pdiffc >>
rect 903 483 949 657
rect 1063 483 1109 657
rect 1223 483 1269 657
rect 1383 483 1429 657
rect 1543 483 1589 657
<< psubdiff >>
rect 622 -55 929 -27
rect 622 -141 706 -55
rect 813 -141 929 -55
rect 622 -159 929 -141
<< nsubdiff >>
rect 656 957 973 996
rect 656 871 734 957
rect 879 871 973 957
rect 656 830 973 871
<< psubdiffcont >>
rect 706 -141 813 -55
<< nsubdiffcont >>
rect 734 871 879 957
<< polysilicon >>
rect 978 670 1034 714
rect 1138 670 1194 714
rect 1298 670 1354 714
rect 1458 670 1514 714
rect 978 428 1034 470
rect 110 341 169 428
rect 12 325 169 341
rect 12 242 29 325
rect 115 322 169 325
rect 271 322 330 427
rect 432 322 491 426
rect 590 322 649 428
rect 974 426 1034 428
rect 1138 427 1194 470
rect 974 341 1033 426
rect 876 325 1033 341
rect 115 270 654 322
rect 115 242 169 270
rect 12 227 169 242
rect 110 210 169 227
rect 271 209 330 270
rect 432 208 491 270
rect 590 210 649 270
rect 876 242 893 325
rect 979 322 1033 325
rect 1135 322 1194 427
rect 1298 426 1354 470
rect 1458 428 1514 470
rect 1454 426 1514 428
rect 1296 322 1355 426
rect 1454 322 1513 426
rect 979 270 1518 322
rect 979 242 1033 270
rect 876 227 1033 242
rect 974 210 1033 227
rect 976 168 1032 210
rect 1135 209 1194 270
rect 1136 168 1192 209
rect 1296 208 1355 270
rect 1454 210 1513 270
rect 1296 168 1352 208
rect 1456 168 1512 210
rect 976 24 1032 68
rect 1136 24 1192 68
rect 1296 24 1352 68
rect 1456 24 1512 68
<< polycontact >>
rect 29 242 115 325
rect 893 242 979 325
<< metal1 >>
rect -64 957 1692 1032
rect -64 871 734 957
rect 879 871 1692 957
rect -64 794 1692 871
rect 30 474 90 794
rect 12 325 140 330
rect 12 322 29 325
rect -63 256 29 322
rect 12 242 29 256
rect 115 242 140 325
rect 12 237 140 242
rect 190 321 250 677
rect 350 478 410 794
rect 507 321 567 681
rect 669 476 729 794
rect 894 657 954 794
rect 894 483 903 657
rect 949 483 954 657
rect 894 474 954 483
rect 1054 657 1114 677
rect 1054 483 1063 657
rect 1109 483 1114 657
rect 903 472 949 474
rect 876 325 1004 330
rect 876 321 893 325
rect 190 269 893 321
rect 30 3 86 171
rect 190 66 250 269
rect 350 3 406 166
rect 507 70 567 269
rect 876 242 893 269
rect 979 242 1004 325
rect 876 237 1004 242
rect 1054 321 1114 483
rect 1214 657 1274 794
rect 1214 483 1223 657
rect 1269 483 1274 657
rect 1214 478 1274 483
rect 1371 657 1431 681
rect 1371 483 1383 657
rect 1429 483 1431 657
rect 1223 472 1269 478
rect 1371 321 1431 483
rect 1533 657 1593 794
rect 1533 483 1543 657
rect 1589 483 1593 657
rect 1533 476 1593 483
rect 1543 472 1589 476
rect 1054 269 1651 321
rect 669 3 725 169
rect 894 155 950 171
rect 894 81 901 155
rect 947 81 950 155
rect 894 3 950 81
rect 1054 155 1114 269
rect 1054 81 1061 155
rect 1107 81 1114 155
rect 1054 66 1114 81
rect 1214 155 1270 166
rect 1214 81 1221 155
rect 1267 81 1270 155
rect 1214 3 1270 81
rect 1371 155 1431 269
rect 1371 81 1381 155
rect 1427 81 1431 155
rect 1371 70 1431 81
rect 1533 155 1589 169
rect 1533 81 1541 155
rect 1587 81 1589 155
rect 1533 3 1589 81
rect -56 -55 1693 3
rect -56 -141 706 -55
rect 813 -141 1693 -55
rect -56 -176 1693 -141
use nmos_3p3_5GGST2  nmos_3p3_5GGST2_0
timestamp 1691575691
transform 1 0 380 0 1 118
box -380 -118 380 118
use pmos_3p3_MWXUAR  pmos_3p3_MWXUAR_0
timestamp 1691575691
transform 1 0 382 0 1 570
box -442 -230 442 230
<< labels >>
flabel nsubdiffcont 810 910 810 910 0 FreeSans 320 0 0 0 VDD
port 0 nsew
flabel psubdiffcont 750 -100 750 -100 0 FreeSans 320 0 0 0 VSS
port 1 nsew
flabel metal1 1610 290 1610 290 0 FreeSans 320 0 0 0 OUT
port 2 nsew
flabel metal1 -40 290 -40 290 0 FreeSans 320 0 0 0 IN
port 3 nsew
<< end >>
