magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -2867 -1019 1019 1019
<< metal3 >>
rect -1867 14 19 19
rect -1867 -14 -1862 14
rect -1834 -14 -1796 14
rect -1768 -14 -1730 14
rect -1702 -14 -1664 14
rect -1636 -14 -1598 14
rect -1570 -14 -1532 14
rect -1504 -14 -1466 14
rect -1438 -14 -1400 14
rect -1372 -14 -1334 14
rect -1306 -14 -1268 14
rect -1240 -14 -1202 14
rect -1174 -14 -1136 14
rect -1108 -14 -1070 14
rect -1042 -14 -1004 14
rect -976 -14 -938 14
rect -910 -14 -872 14
rect -844 -14 -806 14
rect -778 -14 -740 14
rect -712 -14 -674 14
rect -646 -14 -608 14
rect -580 -14 -542 14
rect -514 -14 -476 14
rect -448 -14 -410 14
rect -382 -14 -344 14
rect -316 -14 -278 14
rect -250 -14 -212 14
rect -184 -14 -146 14
rect -118 -14 -80 14
rect -52 -14 -14 14
rect 14 -14 19 14
rect -1867 -19 19 -14
<< via3 >>
rect -1862 -14 -1834 14
rect -1796 -14 -1768 14
rect -1730 -14 -1702 14
rect -1664 -14 -1636 14
rect -1598 -14 -1570 14
rect -1532 -14 -1504 14
rect -1466 -14 -1438 14
rect -1400 -14 -1372 14
rect -1334 -14 -1306 14
rect -1268 -14 -1240 14
rect -1202 -14 -1174 14
rect -1136 -14 -1108 14
rect -1070 -14 -1042 14
rect -1004 -14 -976 14
rect -938 -14 -910 14
rect -872 -14 -844 14
rect -806 -14 -778 14
rect -740 -14 -712 14
rect -674 -14 -646 14
rect -608 -14 -580 14
rect -542 -14 -514 14
rect -476 -14 -448 14
rect -410 -14 -382 14
rect -344 -14 -316 14
rect -278 -14 -250 14
rect -212 -14 -184 14
rect -146 -14 -118 14
rect -80 -14 -52 14
rect -14 -14 14 14
<< metal4 >>
rect -1867 14 19 19
rect -1867 -14 -1862 14
rect -1834 -14 -1796 14
rect -1768 -14 -1730 14
rect -1702 -14 -1664 14
rect -1636 -14 -1598 14
rect -1570 -14 -1532 14
rect -1504 -14 -1466 14
rect -1438 -14 -1400 14
rect -1372 -14 -1334 14
rect -1306 -14 -1268 14
rect -1240 -14 -1202 14
rect -1174 -14 -1136 14
rect -1108 -14 -1070 14
rect -1042 -14 -1004 14
rect -976 -14 -938 14
rect -910 -14 -872 14
rect -844 -14 -806 14
rect -778 -14 -740 14
rect -712 -14 -674 14
rect -646 -14 -608 14
rect -580 -14 -542 14
rect -514 -14 -476 14
rect -448 -14 -410 14
rect -382 -14 -344 14
rect -316 -14 -278 14
rect -250 -14 -212 14
rect -184 -14 -146 14
rect -118 -14 -80 14
rect -52 -14 -14 14
rect 14 -14 19 14
rect -1867 -19 19 -14
<< end >>
