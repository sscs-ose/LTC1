magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2128 -4760 2128 4760
<< nwell >>
rect -128 -2760 128 2760
<< nsubdiff >>
rect -45 2655 45 2677
rect -45 -2655 -23 2655
rect 23 -2655 45 2655
rect -45 -2677 45 -2655
<< nsubdiffcont >>
rect -23 -2655 23 2655
<< metal1 >>
rect -34 2655 34 2666
rect -34 -2655 -23 2655
rect 23 -2655 34 2655
rect -34 -2666 34 -2655
<< end >>
