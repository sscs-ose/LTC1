magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -4883 -1748 4883 1748
<< metal4 >>
rect -3880 740 3880 745
rect -3880 712 -3875 740
rect -3847 712 -3809 740
rect -3781 712 -3743 740
rect -3715 712 -3677 740
rect -3649 712 -3611 740
rect -3583 712 -3545 740
rect -3517 712 -3479 740
rect -3451 712 -3413 740
rect -3385 712 -3347 740
rect -3319 712 -3281 740
rect -3253 712 -3215 740
rect -3187 712 -3149 740
rect -3121 712 -3083 740
rect -3055 712 -3017 740
rect -2989 712 -2951 740
rect -2923 712 -2885 740
rect -2857 712 -2819 740
rect -2791 712 -2753 740
rect -2725 712 -2687 740
rect -2659 712 -2621 740
rect -2593 712 -2555 740
rect -2527 712 -2489 740
rect -2461 712 -2423 740
rect -2395 712 -2357 740
rect -2329 712 -2291 740
rect -2263 712 -2225 740
rect -2197 712 -2159 740
rect -2131 712 -2093 740
rect -2065 712 -2027 740
rect -1999 712 -1961 740
rect -1933 712 -1895 740
rect -1867 712 -1829 740
rect -1801 712 -1763 740
rect -1735 712 -1697 740
rect -1669 712 -1631 740
rect -1603 712 -1565 740
rect -1537 712 -1499 740
rect -1471 712 -1433 740
rect -1405 712 -1367 740
rect -1339 712 -1301 740
rect -1273 712 -1235 740
rect -1207 712 -1169 740
rect -1141 712 -1103 740
rect -1075 712 -1037 740
rect -1009 712 -971 740
rect -943 712 -905 740
rect -877 712 -839 740
rect -811 712 -773 740
rect -745 712 -707 740
rect -679 712 -641 740
rect -613 712 -575 740
rect -547 712 -509 740
rect -481 712 -443 740
rect -415 712 -377 740
rect -349 712 -311 740
rect -283 712 -245 740
rect -217 712 -179 740
rect -151 712 -113 740
rect -85 712 -47 740
rect -19 712 19 740
rect 47 712 85 740
rect 113 712 151 740
rect 179 712 217 740
rect 245 712 283 740
rect 311 712 349 740
rect 377 712 415 740
rect 443 712 481 740
rect 509 712 547 740
rect 575 712 613 740
rect 641 712 679 740
rect 707 712 745 740
rect 773 712 811 740
rect 839 712 877 740
rect 905 712 943 740
rect 971 712 1009 740
rect 1037 712 1075 740
rect 1103 712 1141 740
rect 1169 712 1207 740
rect 1235 712 1273 740
rect 1301 712 1339 740
rect 1367 712 1405 740
rect 1433 712 1471 740
rect 1499 712 1537 740
rect 1565 712 1603 740
rect 1631 712 1669 740
rect 1697 712 1735 740
rect 1763 712 1801 740
rect 1829 712 1867 740
rect 1895 712 1933 740
rect 1961 712 1999 740
rect 2027 712 2065 740
rect 2093 712 2131 740
rect 2159 712 2197 740
rect 2225 712 2263 740
rect 2291 712 2329 740
rect 2357 712 2395 740
rect 2423 712 2461 740
rect 2489 712 2527 740
rect 2555 712 2593 740
rect 2621 712 2659 740
rect 2687 712 2725 740
rect 2753 712 2791 740
rect 2819 712 2857 740
rect 2885 712 2923 740
rect 2951 712 2989 740
rect 3017 712 3055 740
rect 3083 712 3121 740
rect 3149 712 3187 740
rect 3215 712 3253 740
rect 3281 712 3319 740
rect 3347 712 3385 740
rect 3413 712 3451 740
rect 3479 712 3517 740
rect 3545 712 3583 740
rect 3611 712 3649 740
rect 3677 712 3715 740
rect 3743 712 3781 740
rect 3809 712 3847 740
rect 3875 712 3880 740
rect -3880 674 3880 712
rect -3880 646 -3875 674
rect -3847 646 -3809 674
rect -3781 646 -3743 674
rect -3715 646 -3677 674
rect -3649 646 -3611 674
rect -3583 646 -3545 674
rect -3517 646 -3479 674
rect -3451 646 -3413 674
rect -3385 646 -3347 674
rect -3319 646 -3281 674
rect -3253 646 -3215 674
rect -3187 646 -3149 674
rect -3121 646 -3083 674
rect -3055 646 -3017 674
rect -2989 646 -2951 674
rect -2923 646 -2885 674
rect -2857 646 -2819 674
rect -2791 646 -2753 674
rect -2725 646 -2687 674
rect -2659 646 -2621 674
rect -2593 646 -2555 674
rect -2527 646 -2489 674
rect -2461 646 -2423 674
rect -2395 646 -2357 674
rect -2329 646 -2291 674
rect -2263 646 -2225 674
rect -2197 646 -2159 674
rect -2131 646 -2093 674
rect -2065 646 -2027 674
rect -1999 646 -1961 674
rect -1933 646 -1895 674
rect -1867 646 -1829 674
rect -1801 646 -1763 674
rect -1735 646 -1697 674
rect -1669 646 -1631 674
rect -1603 646 -1565 674
rect -1537 646 -1499 674
rect -1471 646 -1433 674
rect -1405 646 -1367 674
rect -1339 646 -1301 674
rect -1273 646 -1235 674
rect -1207 646 -1169 674
rect -1141 646 -1103 674
rect -1075 646 -1037 674
rect -1009 646 -971 674
rect -943 646 -905 674
rect -877 646 -839 674
rect -811 646 -773 674
rect -745 646 -707 674
rect -679 646 -641 674
rect -613 646 -575 674
rect -547 646 -509 674
rect -481 646 -443 674
rect -415 646 -377 674
rect -349 646 -311 674
rect -283 646 -245 674
rect -217 646 -179 674
rect -151 646 -113 674
rect -85 646 -47 674
rect -19 646 19 674
rect 47 646 85 674
rect 113 646 151 674
rect 179 646 217 674
rect 245 646 283 674
rect 311 646 349 674
rect 377 646 415 674
rect 443 646 481 674
rect 509 646 547 674
rect 575 646 613 674
rect 641 646 679 674
rect 707 646 745 674
rect 773 646 811 674
rect 839 646 877 674
rect 905 646 943 674
rect 971 646 1009 674
rect 1037 646 1075 674
rect 1103 646 1141 674
rect 1169 646 1207 674
rect 1235 646 1273 674
rect 1301 646 1339 674
rect 1367 646 1405 674
rect 1433 646 1471 674
rect 1499 646 1537 674
rect 1565 646 1603 674
rect 1631 646 1669 674
rect 1697 646 1735 674
rect 1763 646 1801 674
rect 1829 646 1867 674
rect 1895 646 1933 674
rect 1961 646 1999 674
rect 2027 646 2065 674
rect 2093 646 2131 674
rect 2159 646 2197 674
rect 2225 646 2263 674
rect 2291 646 2329 674
rect 2357 646 2395 674
rect 2423 646 2461 674
rect 2489 646 2527 674
rect 2555 646 2593 674
rect 2621 646 2659 674
rect 2687 646 2725 674
rect 2753 646 2791 674
rect 2819 646 2857 674
rect 2885 646 2923 674
rect 2951 646 2989 674
rect 3017 646 3055 674
rect 3083 646 3121 674
rect 3149 646 3187 674
rect 3215 646 3253 674
rect 3281 646 3319 674
rect 3347 646 3385 674
rect 3413 646 3451 674
rect 3479 646 3517 674
rect 3545 646 3583 674
rect 3611 646 3649 674
rect 3677 646 3715 674
rect 3743 646 3781 674
rect 3809 646 3847 674
rect 3875 646 3880 674
rect -3880 608 3880 646
rect -3880 580 -3875 608
rect -3847 580 -3809 608
rect -3781 580 -3743 608
rect -3715 580 -3677 608
rect -3649 580 -3611 608
rect -3583 580 -3545 608
rect -3517 580 -3479 608
rect -3451 580 -3413 608
rect -3385 580 -3347 608
rect -3319 580 -3281 608
rect -3253 580 -3215 608
rect -3187 580 -3149 608
rect -3121 580 -3083 608
rect -3055 580 -3017 608
rect -2989 580 -2951 608
rect -2923 580 -2885 608
rect -2857 580 -2819 608
rect -2791 580 -2753 608
rect -2725 580 -2687 608
rect -2659 580 -2621 608
rect -2593 580 -2555 608
rect -2527 580 -2489 608
rect -2461 580 -2423 608
rect -2395 580 -2357 608
rect -2329 580 -2291 608
rect -2263 580 -2225 608
rect -2197 580 -2159 608
rect -2131 580 -2093 608
rect -2065 580 -2027 608
rect -1999 580 -1961 608
rect -1933 580 -1895 608
rect -1867 580 -1829 608
rect -1801 580 -1763 608
rect -1735 580 -1697 608
rect -1669 580 -1631 608
rect -1603 580 -1565 608
rect -1537 580 -1499 608
rect -1471 580 -1433 608
rect -1405 580 -1367 608
rect -1339 580 -1301 608
rect -1273 580 -1235 608
rect -1207 580 -1169 608
rect -1141 580 -1103 608
rect -1075 580 -1037 608
rect -1009 580 -971 608
rect -943 580 -905 608
rect -877 580 -839 608
rect -811 580 -773 608
rect -745 580 -707 608
rect -679 580 -641 608
rect -613 580 -575 608
rect -547 580 -509 608
rect -481 580 -443 608
rect -415 580 -377 608
rect -349 580 -311 608
rect -283 580 -245 608
rect -217 580 -179 608
rect -151 580 -113 608
rect -85 580 -47 608
rect -19 580 19 608
rect 47 580 85 608
rect 113 580 151 608
rect 179 580 217 608
rect 245 580 283 608
rect 311 580 349 608
rect 377 580 415 608
rect 443 580 481 608
rect 509 580 547 608
rect 575 580 613 608
rect 641 580 679 608
rect 707 580 745 608
rect 773 580 811 608
rect 839 580 877 608
rect 905 580 943 608
rect 971 580 1009 608
rect 1037 580 1075 608
rect 1103 580 1141 608
rect 1169 580 1207 608
rect 1235 580 1273 608
rect 1301 580 1339 608
rect 1367 580 1405 608
rect 1433 580 1471 608
rect 1499 580 1537 608
rect 1565 580 1603 608
rect 1631 580 1669 608
rect 1697 580 1735 608
rect 1763 580 1801 608
rect 1829 580 1867 608
rect 1895 580 1933 608
rect 1961 580 1999 608
rect 2027 580 2065 608
rect 2093 580 2131 608
rect 2159 580 2197 608
rect 2225 580 2263 608
rect 2291 580 2329 608
rect 2357 580 2395 608
rect 2423 580 2461 608
rect 2489 580 2527 608
rect 2555 580 2593 608
rect 2621 580 2659 608
rect 2687 580 2725 608
rect 2753 580 2791 608
rect 2819 580 2857 608
rect 2885 580 2923 608
rect 2951 580 2989 608
rect 3017 580 3055 608
rect 3083 580 3121 608
rect 3149 580 3187 608
rect 3215 580 3253 608
rect 3281 580 3319 608
rect 3347 580 3385 608
rect 3413 580 3451 608
rect 3479 580 3517 608
rect 3545 580 3583 608
rect 3611 580 3649 608
rect 3677 580 3715 608
rect 3743 580 3781 608
rect 3809 580 3847 608
rect 3875 580 3880 608
rect -3880 542 3880 580
rect -3880 514 -3875 542
rect -3847 514 -3809 542
rect -3781 514 -3743 542
rect -3715 514 -3677 542
rect -3649 514 -3611 542
rect -3583 514 -3545 542
rect -3517 514 -3479 542
rect -3451 514 -3413 542
rect -3385 514 -3347 542
rect -3319 514 -3281 542
rect -3253 514 -3215 542
rect -3187 514 -3149 542
rect -3121 514 -3083 542
rect -3055 514 -3017 542
rect -2989 514 -2951 542
rect -2923 514 -2885 542
rect -2857 514 -2819 542
rect -2791 514 -2753 542
rect -2725 514 -2687 542
rect -2659 514 -2621 542
rect -2593 514 -2555 542
rect -2527 514 -2489 542
rect -2461 514 -2423 542
rect -2395 514 -2357 542
rect -2329 514 -2291 542
rect -2263 514 -2225 542
rect -2197 514 -2159 542
rect -2131 514 -2093 542
rect -2065 514 -2027 542
rect -1999 514 -1961 542
rect -1933 514 -1895 542
rect -1867 514 -1829 542
rect -1801 514 -1763 542
rect -1735 514 -1697 542
rect -1669 514 -1631 542
rect -1603 514 -1565 542
rect -1537 514 -1499 542
rect -1471 514 -1433 542
rect -1405 514 -1367 542
rect -1339 514 -1301 542
rect -1273 514 -1235 542
rect -1207 514 -1169 542
rect -1141 514 -1103 542
rect -1075 514 -1037 542
rect -1009 514 -971 542
rect -943 514 -905 542
rect -877 514 -839 542
rect -811 514 -773 542
rect -745 514 -707 542
rect -679 514 -641 542
rect -613 514 -575 542
rect -547 514 -509 542
rect -481 514 -443 542
rect -415 514 -377 542
rect -349 514 -311 542
rect -283 514 -245 542
rect -217 514 -179 542
rect -151 514 -113 542
rect -85 514 -47 542
rect -19 514 19 542
rect 47 514 85 542
rect 113 514 151 542
rect 179 514 217 542
rect 245 514 283 542
rect 311 514 349 542
rect 377 514 415 542
rect 443 514 481 542
rect 509 514 547 542
rect 575 514 613 542
rect 641 514 679 542
rect 707 514 745 542
rect 773 514 811 542
rect 839 514 877 542
rect 905 514 943 542
rect 971 514 1009 542
rect 1037 514 1075 542
rect 1103 514 1141 542
rect 1169 514 1207 542
rect 1235 514 1273 542
rect 1301 514 1339 542
rect 1367 514 1405 542
rect 1433 514 1471 542
rect 1499 514 1537 542
rect 1565 514 1603 542
rect 1631 514 1669 542
rect 1697 514 1735 542
rect 1763 514 1801 542
rect 1829 514 1867 542
rect 1895 514 1933 542
rect 1961 514 1999 542
rect 2027 514 2065 542
rect 2093 514 2131 542
rect 2159 514 2197 542
rect 2225 514 2263 542
rect 2291 514 2329 542
rect 2357 514 2395 542
rect 2423 514 2461 542
rect 2489 514 2527 542
rect 2555 514 2593 542
rect 2621 514 2659 542
rect 2687 514 2725 542
rect 2753 514 2791 542
rect 2819 514 2857 542
rect 2885 514 2923 542
rect 2951 514 2989 542
rect 3017 514 3055 542
rect 3083 514 3121 542
rect 3149 514 3187 542
rect 3215 514 3253 542
rect 3281 514 3319 542
rect 3347 514 3385 542
rect 3413 514 3451 542
rect 3479 514 3517 542
rect 3545 514 3583 542
rect 3611 514 3649 542
rect 3677 514 3715 542
rect 3743 514 3781 542
rect 3809 514 3847 542
rect 3875 514 3880 542
rect -3880 476 3880 514
rect -3880 448 -3875 476
rect -3847 448 -3809 476
rect -3781 448 -3743 476
rect -3715 448 -3677 476
rect -3649 448 -3611 476
rect -3583 448 -3545 476
rect -3517 448 -3479 476
rect -3451 448 -3413 476
rect -3385 448 -3347 476
rect -3319 448 -3281 476
rect -3253 448 -3215 476
rect -3187 448 -3149 476
rect -3121 448 -3083 476
rect -3055 448 -3017 476
rect -2989 448 -2951 476
rect -2923 448 -2885 476
rect -2857 448 -2819 476
rect -2791 448 -2753 476
rect -2725 448 -2687 476
rect -2659 448 -2621 476
rect -2593 448 -2555 476
rect -2527 448 -2489 476
rect -2461 448 -2423 476
rect -2395 448 -2357 476
rect -2329 448 -2291 476
rect -2263 448 -2225 476
rect -2197 448 -2159 476
rect -2131 448 -2093 476
rect -2065 448 -2027 476
rect -1999 448 -1961 476
rect -1933 448 -1895 476
rect -1867 448 -1829 476
rect -1801 448 -1763 476
rect -1735 448 -1697 476
rect -1669 448 -1631 476
rect -1603 448 -1565 476
rect -1537 448 -1499 476
rect -1471 448 -1433 476
rect -1405 448 -1367 476
rect -1339 448 -1301 476
rect -1273 448 -1235 476
rect -1207 448 -1169 476
rect -1141 448 -1103 476
rect -1075 448 -1037 476
rect -1009 448 -971 476
rect -943 448 -905 476
rect -877 448 -839 476
rect -811 448 -773 476
rect -745 448 -707 476
rect -679 448 -641 476
rect -613 448 -575 476
rect -547 448 -509 476
rect -481 448 -443 476
rect -415 448 -377 476
rect -349 448 -311 476
rect -283 448 -245 476
rect -217 448 -179 476
rect -151 448 -113 476
rect -85 448 -47 476
rect -19 448 19 476
rect 47 448 85 476
rect 113 448 151 476
rect 179 448 217 476
rect 245 448 283 476
rect 311 448 349 476
rect 377 448 415 476
rect 443 448 481 476
rect 509 448 547 476
rect 575 448 613 476
rect 641 448 679 476
rect 707 448 745 476
rect 773 448 811 476
rect 839 448 877 476
rect 905 448 943 476
rect 971 448 1009 476
rect 1037 448 1075 476
rect 1103 448 1141 476
rect 1169 448 1207 476
rect 1235 448 1273 476
rect 1301 448 1339 476
rect 1367 448 1405 476
rect 1433 448 1471 476
rect 1499 448 1537 476
rect 1565 448 1603 476
rect 1631 448 1669 476
rect 1697 448 1735 476
rect 1763 448 1801 476
rect 1829 448 1867 476
rect 1895 448 1933 476
rect 1961 448 1999 476
rect 2027 448 2065 476
rect 2093 448 2131 476
rect 2159 448 2197 476
rect 2225 448 2263 476
rect 2291 448 2329 476
rect 2357 448 2395 476
rect 2423 448 2461 476
rect 2489 448 2527 476
rect 2555 448 2593 476
rect 2621 448 2659 476
rect 2687 448 2725 476
rect 2753 448 2791 476
rect 2819 448 2857 476
rect 2885 448 2923 476
rect 2951 448 2989 476
rect 3017 448 3055 476
rect 3083 448 3121 476
rect 3149 448 3187 476
rect 3215 448 3253 476
rect 3281 448 3319 476
rect 3347 448 3385 476
rect 3413 448 3451 476
rect 3479 448 3517 476
rect 3545 448 3583 476
rect 3611 448 3649 476
rect 3677 448 3715 476
rect 3743 448 3781 476
rect 3809 448 3847 476
rect 3875 448 3880 476
rect -3880 410 3880 448
rect -3880 382 -3875 410
rect -3847 382 -3809 410
rect -3781 382 -3743 410
rect -3715 382 -3677 410
rect -3649 382 -3611 410
rect -3583 382 -3545 410
rect -3517 382 -3479 410
rect -3451 382 -3413 410
rect -3385 382 -3347 410
rect -3319 382 -3281 410
rect -3253 382 -3215 410
rect -3187 382 -3149 410
rect -3121 382 -3083 410
rect -3055 382 -3017 410
rect -2989 382 -2951 410
rect -2923 382 -2885 410
rect -2857 382 -2819 410
rect -2791 382 -2753 410
rect -2725 382 -2687 410
rect -2659 382 -2621 410
rect -2593 382 -2555 410
rect -2527 382 -2489 410
rect -2461 382 -2423 410
rect -2395 382 -2357 410
rect -2329 382 -2291 410
rect -2263 382 -2225 410
rect -2197 382 -2159 410
rect -2131 382 -2093 410
rect -2065 382 -2027 410
rect -1999 382 -1961 410
rect -1933 382 -1895 410
rect -1867 382 -1829 410
rect -1801 382 -1763 410
rect -1735 382 -1697 410
rect -1669 382 -1631 410
rect -1603 382 -1565 410
rect -1537 382 -1499 410
rect -1471 382 -1433 410
rect -1405 382 -1367 410
rect -1339 382 -1301 410
rect -1273 382 -1235 410
rect -1207 382 -1169 410
rect -1141 382 -1103 410
rect -1075 382 -1037 410
rect -1009 382 -971 410
rect -943 382 -905 410
rect -877 382 -839 410
rect -811 382 -773 410
rect -745 382 -707 410
rect -679 382 -641 410
rect -613 382 -575 410
rect -547 382 -509 410
rect -481 382 -443 410
rect -415 382 -377 410
rect -349 382 -311 410
rect -283 382 -245 410
rect -217 382 -179 410
rect -151 382 -113 410
rect -85 382 -47 410
rect -19 382 19 410
rect 47 382 85 410
rect 113 382 151 410
rect 179 382 217 410
rect 245 382 283 410
rect 311 382 349 410
rect 377 382 415 410
rect 443 382 481 410
rect 509 382 547 410
rect 575 382 613 410
rect 641 382 679 410
rect 707 382 745 410
rect 773 382 811 410
rect 839 382 877 410
rect 905 382 943 410
rect 971 382 1009 410
rect 1037 382 1075 410
rect 1103 382 1141 410
rect 1169 382 1207 410
rect 1235 382 1273 410
rect 1301 382 1339 410
rect 1367 382 1405 410
rect 1433 382 1471 410
rect 1499 382 1537 410
rect 1565 382 1603 410
rect 1631 382 1669 410
rect 1697 382 1735 410
rect 1763 382 1801 410
rect 1829 382 1867 410
rect 1895 382 1933 410
rect 1961 382 1999 410
rect 2027 382 2065 410
rect 2093 382 2131 410
rect 2159 382 2197 410
rect 2225 382 2263 410
rect 2291 382 2329 410
rect 2357 382 2395 410
rect 2423 382 2461 410
rect 2489 382 2527 410
rect 2555 382 2593 410
rect 2621 382 2659 410
rect 2687 382 2725 410
rect 2753 382 2791 410
rect 2819 382 2857 410
rect 2885 382 2923 410
rect 2951 382 2989 410
rect 3017 382 3055 410
rect 3083 382 3121 410
rect 3149 382 3187 410
rect 3215 382 3253 410
rect 3281 382 3319 410
rect 3347 382 3385 410
rect 3413 382 3451 410
rect 3479 382 3517 410
rect 3545 382 3583 410
rect 3611 382 3649 410
rect 3677 382 3715 410
rect 3743 382 3781 410
rect 3809 382 3847 410
rect 3875 382 3880 410
rect -3880 344 3880 382
rect -3880 316 -3875 344
rect -3847 316 -3809 344
rect -3781 316 -3743 344
rect -3715 316 -3677 344
rect -3649 316 -3611 344
rect -3583 316 -3545 344
rect -3517 316 -3479 344
rect -3451 316 -3413 344
rect -3385 316 -3347 344
rect -3319 316 -3281 344
rect -3253 316 -3215 344
rect -3187 316 -3149 344
rect -3121 316 -3083 344
rect -3055 316 -3017 344
rect -2989 316 -2951 344
rect -2923 316 -2885 344
rect -2857 316 -2819 344
rect -2791 316 -2753 344
rect -2725 316 -2687 344
rect -2659 316 -2621 344
rect -2593 316 -2555 344
rect -2527 316 -2489 344
rect -2461 316 -2423 344
rect -2395 316 -2357 344
rect -2329 316 -2291 344
rect -2263 316 -2225 344
rect -2197 316 -2159 344
rect -2131 316 -2093 344
rect -2065 316 -2027 344
rect -1999 316 -1961 344
rect -1933 316 -1895 344
rect -1867 316 -1829 344
rect -1801 316 -1763 344
rect -1735 316 -1697 344
rect -1669 316 -1631 344
rect -1603 316 -1565 344
rect -1537 316 -1499 344
rect -1471 316 -1433 344
rect -1405 316 -1367 344
rect -1339 316 -1301 344
rect -1273 316 -1235 344
rect -1207 316 -1169 344
rect -1141 316 -1103 344
rect -1075 316 -1037 344
rect -1009 316 -971 344
rect -943 316 -905 344
rect -877 316 -839 344
rect -811 316 -773 344
rect -745 316 -707 344
rect -679 316 -641 344
rect -613 316 -575 344
rect -547 316 -509 344
rect -481 316 -443 344
rect -415 316 -377 344
rect -349 316 -311 344
rect -283 316 -245 344
rect -217 316 -179 344
rect -151 316 -113 344
rect -85 316 -47 344
rect -19 316 19 344
rect 47 316 85 344
rect 113 316 151 344
rect 179 316 217 344
rect 245 316 283 344
rect 311 316 349 344
rect 377 316 415 344
rect 443 316 481 344
rect 509 316 547 344
rect 575 316 613 344
rect 641 316 679 344
rect 707 316 745 344
rect 773 316 811 344
rect 839 316 877 344
rect 905 316 943 344
rect 971 316 1009 344
rect 1037 316 1075 344
rect 1103 316 1141 344
rect 1169 316 1207 344
rect 1235 316 1273 344
rect 1301 316 1339 344
rect 1367 316 1405 344
rect 1433 316 1471 344
rect 1499 316 1537 344
rect 1565 316 1603 344
rect 1631 316 1669 344
rect 1697 316 1735 344
rect 1763 316 1801 344
rect 1829 316 1867 344
rect 1895 316 1933 344
rect 1961 316 1999 344
rect 2027 316 2065 344
rect 2093 316 2131 344
rect 2159 316 2197 344
rect 2225 316 2263 344
rect 2291 316 2329 344
rect 2357 316 2395 344
rect 2423 316 2461 344
rect 2489 316 2527 344
rect 2555 316 2593 344
rect 2621 316 2659 344
rect 2687 316 2725 344
rect 2753 316 2791 344
rect 2819 316 2857 344
rect 2885 316 2923 344
rect 2951 316 2989 344
rect 3017 316 3055 344
rect 3083 316 3121 344
rect 3149 316 3187 344
rect 3215 316 3253 344
rect 3281 316 3319 344
rect 3347 316 3385 344
rect 3413 316 3451 344
rect 3479 316 3517 344
rect 3545 316 3583 344
rect 3611 316 3649 344
rect 3677 316 3715 344
rect 3743 316 3781 344
rect 3809 316 3847 344
rect 3875 316 3880 344
rect -3880 278 3880 316
rect -3880 250 -3875 278
rect -3847 250 -3809 278
rect -3781 250 -3743 278
rect -3715 250 -3677 278
rect -3649 250 -3611 278
rect -3583 250 -3545 278
rect -3517 250 -3479 278
rect -3451 250 -3413 278
rect -3385 250 -3347 278
rect -3319 250 -3281 278
rect -3253 250 -3215 278
rect -3187 250 -3149 278
rect -3121 250 -3083 278
rect -3055 250 -3017 278
rect -2989 250 -2951 278
rect -2923 250 -2885 278
rect -2857 250 -2819 278
rect -2791 250 -2753 278
rect -2725 250 -2687 278
rect -2659 250 -2621 278
rect -2593 250 -2555 278
rect -2527 250 -2489 278
rect -2461 250 -2423 278
rect -2395 250 -2357 278
rect -2329 250 -2291 278
rect -2263 250 -2225 278
rect -2197 250 -2159 278
rect -2131 250 -2093 278
rect -2065 250 -2027 278
rect -1999 250 -1961 278
rect -1933 250 -1895 278
rect -1867 250 -1829 278
rect -1801 250 -1763 278
rect -1735 250 -1697 278
rect -1669 250 -1631 278
rect -1603 250 -1565 278
rect -1537 250 -1499 278
rect -1471 250 -1433 278
rect -1405 250 -1367 278
rect -1339 250 -1301 278
rect -1273 250 -1235 278
rect -1207 250 -1169 278
rect -1141 250 -1103 278
rect -1075 250 -1037 278
rect -1009 250 -971 278
rect -943 250 -905 278
rect -877 250 -839 278
rect -811 250 -773 278
rect -745 250 -707 278
rect -679 250 -641 278
rect -613 250 -575 278
rect -547 250 -509 278
rect -481 250 -443 278
rect -415 250 -377 278
rect -349 250 -311 278
rect -283 250 -245 278
rect -217 250 -179 278
rect -151 250 -113 278
rect -85 250 -47 278
rect -19 250 19 278
rect 47 250 85 278
rect 113 250 151 278
rect 179 250 217 278
rect 245 250 283 278
rect 311 250 349 278
rect 377 250 415 278
rect 443 250 481 278
rect 509 250 547 278
rect 575 250 613 278
rect 641 250 679 278
rect 707 250 745 278
rect 773 250 811 278
rect 839 250 877 278
rect 905 250 943 278
rect 971 250 1009 278
rect 1037 250 1075 278
rect 1103 250 1141 278
rect 1169 250 1207 278
rect 1235 250 1273 278
rect 1301 250 1339 278
rect 1367 250 1405 278
rect 1433 250 1471 278
rect 1499 250 1537 278
rect 1565 250 1603 278
rect 1631 250 1669 278
rect 1697 250 1735 278
rect 1763 250 1801 278
rect 1829 250 1867 278
rect 1895 250 1933 278
rect 1961 250 1999 278
rect 2027 250 2065 278
rect 2093 250 2131 278
rect 2159 250 2197 278
rect 2225 250 2263 278
rect 2291 250 2329 278
rect 2357 250 2395 278
rect 2423 250 2461 278
rect 2489 250 2527 278
rect 2555 250 2593 278
rect 2621 250 2659 278
rect 2687 250 2725 278
rect 2753 250 2791 278
rect 2819 250 2857 278
rect 2885 250 2923 278
rect 2951 250 2989 278
rect 3017 250 3055 278
rect 3083 250 3121 278
rect 3149 250 3187 278
rect 3215 250 3253 278
rect 3281 250 3319 278
rect 3347 250 3385 278
rect 3413 250 3451 278
rect 3479 250 3517 278
rect 3545 250 3583 278
rect 3611 250 3649 278
rect 3677 250 3715 278
rect 3743 250 3781 278
rect 3809 250 3847 278
rect 3875 250 3880 278
rect -3880 212 3880 250
rect -3880 184 -3875 212
rect -3847 184 -3809 212
rect -3781 184 -3743 212
rect -3715 184 -3677 212
rect -3649 184 -3611 212
rect -3583 184 -3545 212
rect -3517 184 -3479 212
rect -3451 184 -3413 212
rect -3385 184 -3347 212
rect -3319 184 -3281 212
rect -3253 184 -3215 212
rect -3187 184 -3149 212
rect -3121 184 -3083 212
rect -3055 184 -3017 212
rect -2989 184 -2951 212
rect -2923 184 -2885 212
rect -2857 184 -2819 212
rect -2791 184 -2753 212
rect -2725 184 -2687 212
rect -2659 184 -2621 212
rect -2593 184 -2555 212
rect -2527 184 -2489 212
rect -2461 184 -2423 212
rect -2395 184 -2357 212
rect -2329 184 -2291 212
rect -2263 184 -2225 212
rect -2197 184 -2159 212
rect -2131 184 -2093 212
rect -2065 184 -2027 212
rect -1999 184 -1961 212
rect -1933 184 -1895 212
rect -1867 184 -1829 212
rect -1801 184 -1763 212
rect -1735 184 -1697 212
rect -1669 184 -1631 212
rect -1603 184 -1565 212
rect -1537 184 -1499 212
rect -1471 184 -1433 212
rect -1405 184 -1367 212
rect -1339 184 -1301 212
rect -1273 184 -1235 212
rect -1207 184 -1169 212
rect -1141 184 -1103 212
rect -1075 184 -1037 212
rect -1009 184 -971 212
rect -943 184 -905 212
rect -877 184 -839 212
rect -811 184 -773 212
rect -745 184 -707 212
rect -679 184 -641 212
rect -613 184 -575 212
rect -547 184 -509 212
rect -481 184 -443 212
rect -415 184 -377 212
rect -349 184 -311 212
rect -283 184 -245 212
rect -217 184 -179 212
rect -151 184 -113 212
rect -85 184 -47 212
rect -19 184 19 212
rect 47 184 85 212
rect 113 184 151 212
rect 179 184 217 212
rect 245 184 283 212
rect 311 184 349 212
rect 377 184 415 212
rect 443 184 481 212
rect 509 184 547 212
rect 575 184 613 212
rect 641 184 679 212
rect 707 184 745 212
rect 773 184 811 212
rect 839 184 877 212
rect 905 184 943 212
rect 971 184 1009 212
rect 1037 184 1075 212
rect 1103 184 1141 212
rect 1169 184 1207 212
rect 1235 184 1273 212
rect 1301 184 1339 212
rect 1367 184 1405 212
rect 1433 184 1471 212
rect 1499 184 1537 212
rect 1565 184 1603 212
rect 1631 184 1669 212
rect 1697 184 1735 212
rect 1763 184 1801 212
rect 1829 184 1867 212
rect 1895 184 1933 212
rect 1961 184 1999 212
rect 2027 184 2065 212
rect 2093 184 2131 212
rect 2159 184 2197 212
rect 2225 184 2263 212
rect 2291 184 2329 212
rect 2357 184 2395 212
rect 2423 184 2461 212
rect 2489 184 2527 212
rect 2555 184 2593 212
rect 2621 184 2659 212
rect 2687 184 2725 212
rect 2753 184 2791 212
rect 2819 184 2857 212
rect 2885 184 2923 212
rect 2951 184 2989 212
rect 3017 184 3055 212
rect 3083 184 3121 212
rect 3149 184 3187 212
rect 3215 184 3253 212
rect 3281 184 3319 212
rect 3347 184 3385 212
rect 3413 184 3451 212
rect 3479 184 3517 212
rect 3545 184 3583 212
rect 3611 184 3649 212
rect 3677 184 3715 212
rect 3743 184 3781 212
rect 3809 184 3847 212
rect 3875 184 3880 212
rect -3880 146 3880 184
rect -3880 118 -3875 146
rect -3847 118 -3809 146
rect -3781 118 -3743 146
rect -3715 118 -3677 146
rect -3649 118 -3611 146
rect -3583 118 -3545 146
rect -3517 118 -3479 146
rect -3451 118 -3413 146
rect -3385 118 -3347 146
rect -3319 118 -3281 146
rect -3253 118 -3215 146
rect -3187 118 -3149 146
rect -3121 118 -3083 146
rect -3055 118 -3017 146
rect -2989 118 -2951 146
rect -2923 118 -2885 146
rect -2857 118 -2819 146
rect -2791 118 -2753 146
rect -2725 118 -2687 146
rect -2659 118 -2621 146
rect -2593 118 -2555 146
rect -2527 118 -2489 146
rect -2461 118 -2423 146
rect -2395 118 -2357 146
rect -2329 118 -2291 146
rect -2263 118 -2225 146
rect -2197 118 -2159 146
rect -2131 118 -2093 146
rect -2065 118 -2027 146
rect -1999 118 -1961 146
rect -1933 118 -1895 146
rect -1867 118 -1829 146
rect -1801 118 -1763 146
rect -1735 118 -1697 146
rect -1669 118 -1631 146
rect -1603 118 -1565 146
rect -1537 118 -1499 146
rect -1471 118 -1433 146
rect -1405 118 -1367 146
rect -1339 118 -1301 146
rect -1273 118 -1235 146
rect -1207 118 -1169 146
rect -1141 118 -1103 146
rect -1075 118 -1037 146
rect -1009 118 -971 146
rect -943 118 -905 146
rect -877 118 -839 146
rect -811 118 -773 146
rect -745 118 -707 146
rect -679 118 -641 146
rect -613 118 -575 146
rect -547 118 -509 146
rect -481 118 -443 146
rect -415 118 -377 146
rect -349 118 -311 146
rect -283 118 -245 146
rect -217 118 -179 146
rect -151 118 -113 146
rect -85 118 -47 146
rect -19 118 19 146
rect 47 118 85 146
rect 113 118 151 146
rect 179 118 217 146
rect 245 118 283 146
rect 311 118 349 146
rect 377 118 415 146
rect 443 118 481 146
rect 509 118 547 146
rect 575 118 613 146
rect 641 118 679 146
rect 707 118 745 146
rect 773 118 811 146
rect 839 118 877 146
rect 905 118 943 146
rect 971 118 1009 146
rect 1037 118 1075 146
rect 1103 118 1141 146
rect 1169 118 1207 146
rect 1235 118 1273 146
rect 1301 118 1339 146
rect 1367 118 1405 146
rect 1433 118 1471 146
rect 1499 118 1537 146
rect 1565 118 1603 146
rect 1631 118 1669 146
rect 1697 118 1735 146
rect 1763 118 1801 146
rect 1829 118 1867 146
rect 1895 118 1933 146
rect 1961 118 1999 146
rect 2027 118 2065 146
rect 2093 118 2131 146
rect 2159 118 2197 146
rect 2225 118 2263 146
rect 2291 118 2329 146
rect 2357 118 2395 146
rect 2423 118 2461 146
rect 2489 118 2527 146
rect 2555 118 2593 146
rect 2621 118 2659 146
rect 2687 118 2725 146
rect 2753 118 2791 146
rect 2819 118 2857 146
rect 2885 118 2923 146
rect 2951 118 2989 146
rect 3017 118 3055 146
rect 3083 118 3121 146
rect 3149 118 3187 146
rect 3215 118 3253 146
rect 3281 118 3319 146
rect 3347 118 3385 146
rect 3413 118 3451 146
rect 3479 118 3517 146
rect 3545 118 3583 146
rect 3611 118 3649 146
rect 3677 118 3715 146
rect 3743 118 3781 146
rect 3809 118 3847 146
rect 3875 118 3880 146
rect -3880 80 3880 118
rect -3880 52 -3875 80
rect -3847 52 -3809 80
rect -3781 52 -3743 80
rect -3715 52 -3677 80
rect -3649 52 -3611 80
rect -3583 52 -3545 80
rect -3517 52 -3479 80
rect -3451 52 -3413 80
rect -3385 52 -3347 80
rect -3319 52 -3281 80
rect -3253 52 -3215 80
rect -3187 52 -3149 80
rect -3121 52 -3083 80
rect -3055 52 -3017 80
rect -2989 52 -2951 80
rect -2923 52 -2885 80
rect -2857 52 -2819 80
rect -2791 52 -2753 80
rect -2725 52 -2687 80
rect -2659 52 -2621 80
rect -2593 52 -2555 80
rect -2527 52 -2489 80
rect -2461 52 -2423 80
rect -2395 52 -2357 80
rect -2329 52 -2291 80
rect -2263 52 -2225 80
rect -2197 52 -2159 80
rect -2131 52 -2093 80
rect -2065 52 -2027 80
rect -1999 52 -1961 80
rect -1933 52 -1895 80
rect -1867 52 -1829 80
rect -1801 52 -1763 80
rect -1735 52 -1697 80
rect -1669 52 -1631 80
rect -1603 52 -1565 80
rect -1537 52 -1499 80
rect -1471 52 -1433 80
rect -1405 52 -1367 80
rect -1339 52 -1301 80
rect -1273 52 -1235 80
rect -1207 52 -1169 80
rect -1141 52 -1103 80
rect -1075 52 -1037 80
rect -1009 52 -971 80
rect -943 52 -905 80
rect -877 52 -839 80
rect -811 52 -773 80
rect -745 52 -707 80
rect -679 52 -641 80
rect -613 52 -575 80
rect -547 52 -509 80
rect -481 52 -443 80
rect -415 52 -377 80
rect -349 52 -311 80
rect -283 52 -245 80
rect -217 52 -179 80
rect -151 52 -113 80
rect -85 52 -47 80
rect -19 52 19 80
rect 47 52 85 80
rect 113 52 151 80
rect 179 52 217 80
rect 245 52 283 80
rect 311 52 349 80
rect 377 52 415 80
rect 443 52 481 80
rect 509 52 547 80
rect 575 52 613 80
rect 641 52 679 80
rect 707 52 745 80
rect 773 52 811 80
rect 839 52 877 80
rect 905 52 943 80
rect 971 52 1009 80
rect 1037 52 1075 80
rect 1103 52 1141 80
rect 1169 52 1207 80
rect 1235 52 1273 80
rect 1301 52 1339 80
rect 1367 52 1405 80
rect 1433 52 1471 80
rect 1499 52 1537 80
rect 1565 52 1603 80
rect 1631 52 1669 80
rect 1697 52 1735 80
rect 1763 52 1801 80
rect 1829 52 1867 80
rect 1895 52 1933 80
rect 1961 52 1999 80
rect 2027 52 2065 80
rect 2093 52 2131 80
rect 2159 52 2197 80
rect 2225 52 2263 80
rect 2291 52 2329 80
rect 2357 52 2395 80
rect 2423 52 2461 80
rect 2489 52 2527 80
rect 2555 52 2593 80
rect 2621 52 2659 80
rect 2687 52 2725 80
rect 2753 52 2791 80
rect 2819 52 2857 80
rect 2885 52 2923 80
rect 2951 52 2989 80
rect 3017 52 3055 80
rect 3083 52 3121 80
rect 3149 52 3187 80
rect 3215 52 3253 80
rect 3281 52 3319 80
rect 3347 52 3385 80
rect 3413 52 3451 80
rect 3479 52 3517 80
rect 3545 52 3583 80
rect 3611 52 3649 80
rect 3677 52 3715 80
rect 3743 52 3781 80
rect 3809 52 3847 80
rect 3875 52 3880 80
rect -3880 14 3880 52
rect -3880 -14 -3875 14
rect -3847 -14 -3809 14
rect -3781 -14 -3743 14
rect -3715 -14 -3677 14
rect -3649 -14 -3611 14
rect -3583 -14 -3545 14
rect -3517 -14 -3479 14
rect -3451 -14 -3413 14
rect -3385 -14 -3347 14
rect -3319 -14 -3281 14
rect -3253 -14 -3215 14
rect -3187 -14 -3149 14
rect -3121 -14 -3083 14
rect -3055 -14 -3017 14
rect -2989 -14 -2951 14
rect -2923 -14 -2885 14
rect -2857 -14 -2819 14
rect -2791 -14 -2753 14
rect -2725 -14 -2687 14
rect -2659 -14 -2621 14
rect -2593 -14 -2555 14
rect -2527 -14 -2489 14
rect -2461 -14 -2423 14
rect -2395 -14 -2357 14
rect -2329 -14 -2291 14
rect -2263 -14 -2225 14
rect -2197 -14 -2159 14
rect -2131 -14 -2093 14
rect -2065 -14 -2027 14
rect -1999 -14 -1961 14
rect -1933 -14 -1895 14
rect -1867 -14 -1829 14
rect -1801 -14 -1763 14
rect -1735 -14 -1697 14
rect -1669 -14 -1631 14
rect -1603 -14 -1565 14
rect -1537 -14 -1499 14
rect -1471 -14 -1433 14
rect -1405 -14 -1367 14
rect -1339 -14 -1301 14
rect -1273 -14 -1235 14
rect -1207 -14 -1169 14
rect -1141 -14 -1103 14
rect -1075 -14 -1037 14
rect -1009 -14 -971 14
rect -943 -14 -905 14
rect -877 -14 -839 14
rect -811 -14 -773 14
rect -745 -14 -707 14
rect -679 -14 -641 14
rect -613 -14 -575 14
rect -547 -14 -509 14
rect -481 -14 -443 14
rect -415 -14 -377 14
rect -349 -14 -311 14
rect -283 -14 -245 14
rect -217 -14 -179 14
rect -151 -14 -113 14
rect -85 -14 -47 14
rect -19 -14 19 14
rect 47 -14 85 14
rect 113 -14 151 14
rect 179 -14 217 14
rect 245 -14 283 14
rect 311 -14 349 14
rect 377 -14 415 14
rect 443 -14 481 14
rect 509 -14 547 14
rect 575 -14 613 14
rect 641 -14 679 14
rect 707 -14 745 14
rect 773 -14 811 14
rect 839 -14 877 14
rect 905 -14 943 14
rect 971 -14 1009 14
rect 1037 -14 1075 14
rect 1103 -14 1141 14
rect 1169 -14 1207 14
rect 1235 -14 1273 14
rect 1301 -14 1339 14
rect 1367 -14 1405 14
rect 1433 -14 1471 14
rect 1499 -14 1537 14
rect 1565 -14 1603 14
rect 1631 -14 1669 14
rect 1697 -14 1735 14
rect 1763 -14 1801 14
rect 1829 -14 1867 14
rect 1895 -14 1933 14
rect 1961 -14 1999 14
rect 2027 -14 2065 14
rect 2093 -14 2131 14
rect 2159 -14 2197 14
rect 2225 -14 2263 14
rect 2291 -14 2329 14
rect 2357 -14 2395 14
rect 2423 -14 2461 14
rect 2489 -14 2527 14
rect 2555 -14 2593 14
rect 2621 -14 2659 14
rect 2687 -14 2725 14
rect 2753 -14 2791 14
rect 2819 -14 2857 14
rect 2885 -14 2923 14
rect 2951 -14 2989 14
rect 3017 -14 3055 14
rect 3083 -14 3121 14
rect 3149 -14 3187 14
rect 3215 -14 3253 14
rect 3281 -14 3319 14
rect 3347 -14 3385 14
rect 3413 -14 3451 14
rect 3479 -14 3517 14
rect 3545 -14 3583 14
rect 3611 -14 3649 14
rect 3677 -14 3715 14
rect 3743 -14 3781 14
rect 3809 -14 3847 14
rect 3875 -14 3880 14
rect -3880 -52 3880 -14
rect -3880 -80 -3875 -52
rect -3847 -80 -3809 -52
rect -3781 -80 -3743 -52
rect -3715 -80 -3677 -52
rect -3649 -80 -3611 -52
rect -3583 -80 -3545 -52
rect -3517 -80 -3479 -52
rect -3451 -80 -3413 -52
rect -3385 -80 -3347 -52
rect -3319 -80 -3281 -52
rect -3253 -80 -3215 -52
rect -3187 -80 -3149 -52
rect -3121 -80 -3083 -52
rect -3055 -80 -3017 -52
rect -2989 -80 -2951 -52
rect -2923 -80 -2885 -52
rect -2857 -80 -2819 -52
rect -2791 -80 -2753 -52
rect -2725 -80 -2687 -52
rect -2659 -80 -2621 -52
rect -2593 -80 -2555 -52
rect -2527 -80 -2489 -52
rect -2461 -80 -2423 -52
rect -2395 -80 -2357 -52
rect -2329 -80 -2291 -52
rect -2263 -80 -2225 -52
rect -2197 -80 -2159 -52
rect -2131 -80 -2093 -52
rect -2065 -80 -2027 -52
rect -1999 -80 -1961 -52
rect -1933 -80 -1895 -52
rect -1867 -80 -1829 -52
rect -1801 -80 -1763 -52
rect -1735 -80 -1697 -52
rect -1669 -80 -1631 -52
rect -1603 -80 -1565 -52
rect -1537 -80 -1499 -52
rect -1471 -80 -1433 -52
rect -1405 -80 -1367 -52
rect -1339 -80 -1301 -52
rect -1273 -80 -1235 -52
rect -1207 -80 -1169 -52
rect -1141 -80 -1103 -52
rect -1075 -80 -1037 -52
rect -1009 -80 -971 -52
rect -943 -80 -905 -52
rect -877 -80 -839 -52
rect -811 -80 -773 -52
rect -745 -80 -707 -52
rect -679 -80 -641 -52
rect -613 -80 -575 -52
rect -547 -80 -509 -52
rect -481 -80 -443 -52
rect -415 -80 -377 -52
rect -349 -80 -311 -52
rect -283 -80 -245 -52
rect -217 -80 -179 -52
rect -151 -80 -113 -52
rect -85 -80 -47 -52
rect -19 -80 19 -52
rect 47 -80 85 -52
rect 113 -80 151 -52
rect 179 -80 217 -52
rect 245 -80 283 -52
rect 311 -80 349 -52
rect 377 -80 415 -52
rect 443 -80 481 -52
rect 509 -80 547 -52
rect 575 -80 613 -52
rect 641 -80 679 -52
rect 707 -80 745 -52
rect 773 -80 811 -52
rect 839 -80 877 -52
rect 905 -80 943 -52
rect 971 -80 1009 -52
rect 1037 -80 1075 -52
rect 1103 -80 1141 -52
rect 1169 -80 1207 -52
rect 1235 -80 1273 -52
rect 1301 -80 1339 -52
rect 1367 -80 1405 -52
rect 1433 -80 1471 -52
rect 1499 -80 1537 -52
rect 1565 -80 1603 -52
rect 1631 -80 1669 -52
rect 1697 -80 1735 -52
rect 1763 -80 1801 -52
rect 1829 -80 1867 -52
rect 1895 -80 1933 -52
rect 1961 -80 1999 -52
rect 2027 -80 2065 -52
rect 2093 -80 2131 -52
rect 2159 -80 2197 -52
rect 2225 -80 2263 -52
rect 2291 -80 2329 -52
rect 2357 -80 2395 -52
rect 2423 -80 2461 -52
rect 2489 -80 2527 -52
rect 2555 -80 2593 -52
rect 2621 -80 2659 -52
rect 2687 -80 2725 -52
rect 2753 -80 2791 -52
rect 2819 -80 2857 -52
rect 2885 -80 2923 -52
rect 2951 -80 2989 -52
rect 3017 -80 3055 -52
rect 3083 -80 3121 -52
rect 3149 -80 3187 -52
rect 3215 -80 3253 -52
rect 3281 -80 3319 -52
rect 3347 -80 3385 -52
rect 3413 -80 3451 -52
rect 3479 -80 3517 -52
rect 3545 -80 3583 -52
rect 3611 -80 3649 -52
rect 3677 -80 3715 -52
rect 3743 -80 3781 -52
rect 3809 -80 3847 -52
rect 3875 -80 3880 -52
rect -3880 -118 3880 -80
rect -3880 -146 -3875 -118
rect -3847 -146 -3809 -118
rect -3781 -146 -3743 -118
rect -3715 -146 -3677 -118
rect -3649 -146 -3611 -118
rect -3583 -146 -3545 -118
rect -3517 -146 -3479 -118
rect -3451 -146 -3413 -118
rect -3385 -146 -3347 -118
rect -3319 -146 -3281 -118
rect -3253 -146 -3215 -118
rect -3187 -146 -3149 -118
rect -3121 -146 -3083 -118
rect -3055 -146 -3017 -118
rect -2989 -146 -2951 -118
rect -2923 -146 -2885 -118
rect -2857 -146 -2819 -118
rect -2791 -146 -2753 -118
rect -2725 -146 -2687 -118
rect -2659 -146 -2621 -118
rect -2593 -146 -2555 -118
rect -2527 -146 -2489 -118
rect -2461 -146 -2423 -118
rect -2395 -146 -2357 -118
rect -2329 -146 -2291 -118
rect -2263 -146 -2225 -118
rect -2197 -146 -2159 -118
rect -2131 -146 -2093 -118
rect -2065 -146 -2027 -118
rect -1999 -146 -1961 -118
rect -1933 -146 -1895 -118
rect -1867 -146 -1829 -118
rect -1801 -146 -1763 -118
rect -1735 -146 -1697 -118
rect -1669 -146 -1631 -118
rect -1603 -146 -1565 -118
rect -1537 -146 -1499 -118
rect -1471 -146 -1433 -118
rect -1405 -146 -1367 -118
rect -1339 -146 -1301 -118
rect -1273 -146 -1235 -118
rect -1207 -146 -1169 -118
rect -1141 -146 -1103 -118
rect -1075 -146 -1037 -118
rect -1009 -146 -971 -118
rect -943 -146 -905 -118
rect -877 -146 -839 -118
rect -811 -146 -773 -118
rect -745 -146 -707 -118
rect -679 -146 -641 -118
rect -613 -146 -575 -118
rect -547 -146 -509 -118
rect -481 -146 -443 -118
rect -415 -146 -377 -118
rect -349 -146 -311 -118
rect -283 -146 -245 -118
rect -217 -146 -179 -118
rect -151 -146 -113 -118
rect -85 -146 -47 -118
rect -19 -146 19 -118
rect 47 -146 85 -118
rect 113 -146 151 -118
rect 179 -146 217 -118
rect 245 -146 283 -118
rect 311 -146 349 -118
rect 377 -146 415 -118
rect 443 -146 481 -118
rect 509 -146 547 -118
rect 575 -146 613 -118
rect 641 -146 679 -118
rect 707 -146 745 -118
rect 773 -146 811 -118
rect 839 -146 877 -118
rect 905 -146 943 -118
rect 971 -146 1009 -118
rect 1037 -146 1075 -118
rect 1103 -146 1141 -118
rect 1169 -146 1207 -118
rect 1235 -146 1273 -118
rect 1301 -146 1339 -118
rect 1367 -146 1405 -118
rect 1433 -146 1471 -118
rect 1499 -146 1537 -118
rect 1565 -146 1603 -118
rect 1631 -146 1669 -118
rect 1697 -146 1735 -118
rect 1763 -146 1801 -118
rect 1829 -146 1867 -118
rect 1895 -146 1933 -118
rect 1961 -146 1999 -118
rect 2027 -146 2065 -118
rect 2093 -146 2131 -118
rect 2159 -146 2197 -118
rect 2225 -146 2263 -118
rect 2291 -146 2329 -118
rect 2357 -146 2395 -118
rect 2423 -146 2461 -118
rect 2489 -146 2527 -118
rect 2555 -146 2593 -118
rect 2621 -146 2659 -118
rect 2687 -146 2725 -118
rect 2753 -146 2791 -118
rect 2819 -146 2857 -118
rect 2885 -146 2923 -118
rect 2951 -146 2989 -118
rect 3017 -146 3055 -118
rect 3083 -146 3121 -118
rect 3149 -146 3187 -118
rect 3215 -146 3253 -118
rect 3281 -146 3319 -118
rect 3347 -146 3385 -118
rect 3413 -146 3451 -118
rect 3479 -146 3517 -118
rect 3545 -146 3583 -118
rect 3611 -146 3649 -118
rect 3677 -146 3715 -118
rect 3743 -146 3781 -118
rect 3809 -146 3847 -118
rect 3875 -146 3880 -118
rect -3880 -184 3880 -146
rect -3880 -212 -3875 -184
rect -3847 -212 -3809 -184
rect -3781 -212 -3743 -184
rect -3715 -212 -3677 -184
rect -3649 -212 -3611 -184
rect -3583 -212 -3545 -184
rect -3517 -212 -3479 -184
rect -3451 -212 -3413 -184
rect -3385 -212 -3347 -184
rect -3319 -212 -3281 -184
rect -3253 -212 -3215 -184
rect -3187 -212 -3149 -184
rect -3121 -212 -3083 -184
rect -3055 -212 -3017 -184
rect -2989 -212 -2951 -184
rect -2923 -212 -2885 -184
rect -2857 -212 -2819 -184
rect -2791 -212 -2753 -184
rect -2725 -212 -2687 -184
rect -2659 -212 -2621 -184
rect -2593 -212 -2555 -184
rect -2527 -212 -2489 -184
rect -2461 -212 -2423 -184
rect -2395 -212 -2357 -184
rect -2329 -212 -2291 -184
rect -2263 -212 -2225 -184
rect -2197 -212 -2159 -184
rect -2131 -212 -2093 -184
rect -2065 -212 -2027 -184
rect -1999 -212 -1961 -184
rect -1933 -212 -1895 -184
rect -1867 -212 -1829 -184
rect -1801 -212 -1763 -184
rect -1735 -212 -1697 -184
rect -1669 -212 -1631 -184
rect -1603 -212 -1565 -184
rect -1537 -212 -1499 -184
rect -1471 -212 -1433 -184
rect -1405 -212 -1367 -184
rect -1339 -212 -1301 -184
rect -1273 -212 -1235 -184
rect -1207 -212 -1169 -184
rect -1141 -212 -1103 -184
rect -1075 -212 -1037 -184
rect -1009 -212 -971 -184
rect -943 -212 -905 -184
rect -877 -212 -839 -184
rect -811 -212 -773 -184
rect -745 -212 -707 -184
rect -679 -212 -641 -184
rect -613 -212 -575 -184
rect -547 -212 -509 -184
rect -481 -212 -443 -184
rect -415 -212 -377 -184
rect -349 -212 -311 -184
rect -283 -212 -245 -184
rect -217 -212 -179 -184
rect -151 -212 -113 -184
rect -85 -212 -47 -184
rect -19 -212 19 -184
rect 47 -212 85 -184
rect 113 -212 151 -184
rect 179 -212 217 -184
rect 245 -212 283 -184
rect 311 -212 349 -184
rect 377 -212 415 -184
rect 443 -212 481 -184
rect 509 -212 547 -184
rect 575 -212 613 -184
rect 641 -212 679 -184
rect 707 -212 745 -184
rect 773 -212 811 -184
rect 839 -212 877 -184
rect 905 -212 943 -184
rect 971 -212 1009 -184
rect 1037 -212 1075 -184
rect 1103 -212 1141 -184
rect 1169 -212 1207 -184
rect 1235 -212 1273 -184
rect 1301 -212 1339 -184
rect 1367 -212 1405 -184
rect 1433 -212 1471 -184
rect 1499 -212 1537 -184
rect 1565 -212 1603 -184
rect 1631 -212 1669 -184
rect 1697 -212 1735 -184
rect 1763 -212 1801 -184
rect 1829 -212 1867 -184
rect 1895 -212 1933 -184
rect 1961 -212 1999 -184
rect 2027 -212 2065 -184
rect 2093 -212 2131 -184
rect 2159 -212 2197 -184
rect 2225 -212 2263 -184
rect 2291 -212 2329 -184
rect 2357 -212 2395 -184
rect 2423 -212 2461 -184
rect 2489 -212 2527 -184
rect 2555 -212 2593 -184
rect 2621 -212 2659 -184
rect 2687 -212 2725 -184
rect 2753 -212 2791 -184
rect 2819 -212 2857 -184
rect 2885 -212 2923 -184
rect 2951 -212 2989 -184
rect 3017 -212 3055 -184
rect 3083 -212 3121 -184
rect 3149 -212 3187 -184
rect 3215 -212 3253 -184
rect 3281 -212 3319 -184
rect 3347 -212 3385 -184
rect 3413 -212 3451 -184
rect 3479 -212 3517 -184
rect 3545 -212 3583 -184
rect 3611 -212 3649 -184
rect 3677 -212 3715 -184
rect 3743 -212 3781 -184
rect 3809 -212 3847 -184
rect 3875 -212 3880 -184
rect -3880 -250 3880 -212
rect -3880 -278 -3875 -250
rect -3847 -278 -3809 -250
rect -3781 -278 -3743 -250
rect -3715 -278 -3677 -250
rect -3649 -278 -3611 -250
rect -3583 -278 -3545 -250
rect -3517 -278 -3479 -250
rect -3451 -278 -3413 -250
rect -3385 -278 -3347 -250
rect -3319 -278 -3281 -250
rect -3253 -278 -3215 -250
rect -3187 -278 -3149 -250
rect -3121 -278 -3083 -250
rect -3055 -278 -3017 -250
rect -2989 -278 -2951 -250
rect -2923 -278 -2885 -250
rect -2857 -278 -2819 -250
rect -2791 -278 -2753 -250
rect -2725 -278 -2687 -250
rect -2659 -278 -2621 -250
rect -2593 -278 -2555 -250
rect -2527 -278 -2489 -250
rect -2461 -278 -2423 -250
rect -2395 -278 -2357 -250
rect -2329 -278 -2291 -250
rect -2263 -278 -2225 -250
rect -2197 -278 -2159 -250
rect -2131 -278 -2093 -250
rect -2065 -278 -2027 -250
rect -1999 -278 -1961 -250
rect -1933 -278 -1895 -250
rect -1867 -278 -1829 -250
rect -1801 -278 -1763 -250
rect -1735 -278 -1697 -250
rect -1669 -278 -1631 -250
rect -1603 -278 -1565 -250
rect -1537 -278 -1499 -250
rect -1471 -278 -1433 -250
rect -1405 -278 -1367 -250
rect -1339 -278 -1301 -250
rect -1273 -278 -1235 -250
rect -1207 -278 -1169 -250
rect -1141 -278 -1103 -250
rect -1075 -278 -1037 -250
rect -1009 -278 -971 -250
rect -943 -278 -905 -250
rect -877 -278 -839 -250
rect -811 -278 -773 -250
rect -745 -278 -707 -250
rect -679 -278 -641 -250
rect -613 -278 -575 -250
rect -547 -278 -509 -250
rect -481 -278 -443 -250
rect -415 -278 -377 -250
rect -349 -278 -311 -250
rect -283 -278 -245 -250
rect -217 -278 -179 -250
rect -151 -278 -113 -250
rect -85 -278 -47 -250
rect -19 -278 19 -250
rect 47 -278 85 -250
rect 113 -278 151 -250
rect 179 -278 217 -250
rect 245 -278 283 -250
rect 311 -278 349 -250
rect 377 -278 415 -250
rect 443 -278 481 -250
rect 509 -278 547 -250
rect 575 -278 613 -250
rect 641 -278 679 -250
rect 707 -278 745 -250
rect 773 -278 811 -250
rect 839 -278 877 -250
rect 905 -278 943 -250
rect 971 -278 1009 -250
rect 1037 -278 1075 -250
rect 1103 -278 1141 -250
rect 1169 -278 1207 -250
rect 1235 -278 1273 -250
rect 1301 -278 1339 -250
rect 1367 -278 1405 -250
rect 1433 -278 1471 -250
rect 1499 -278 1537 -250
rect 1565 -278 1603 -250
rect 1631 -278 1669 -250
rect 1697 -278 1735 -250
rect 1763 -278 1801 -250
rect 1829 -278 1867 -250
rect 1895 -278 1933 -250
rect 1961 -278 1999 -250
rect 2027 -278 2065 -250
rect 2093 -278 2131 -250
rect 2159 -278 2197 -250
rect 2225 -278 2263 -250
rect 2291 -278 2329 -250
rect 2357 -278 2395 -250
rect 2423 -278 2461 -250
rect 2489 -278 2527 -250
rect 2555 -278 2593 -250
rect 2621 -278 2659 -250
rect 2687 -278 2725 -250
rect 2753 -278 2791 -250
rect 2819 -278 2857 -250
rect 2885 -278 2923 -250
rect 2951 -278 2989 -250
rect 3017 -278 3055 -250
rect 3083 -278 3121 -250
rect 3149 -278 3187 -250
rect 3215 -278 3253 -250
rect 3281 -278 3319 -250
rect 3347 -278 3385 -250
rect 3413 -278 3451 -250
rect 3479 -278 3517 -250
rect 3545 -278 3583 -250
rect 3611 -278 3649 -250
rect 3677 -278 3715 -250
rect 3743 -278 3781 -250
rect 3809 -278 3847 -250
rect 3875 -278 3880 -250
rect -3880 -316 3880 -278
rect -3880 -344 -3875 -316
rect -3847 -344 -3809 -316
rect -3781 -344 -3743 -316
rect -3715 -344 -3677 -316
rect -3649 -344 -3611 -316
rect -3583 -344 -3545 -316
rect -3517 -344 -3479 -316
rect -3451 -344 -3413 -316
rect -3385 -344 -3347 -316
rect -3319 -344 -3281 -316
rect -3253 -344 -3215 -316
rect -3187 -344 -3149 -316
rect -3121 -344 -3083 -316
rect -3055 -344 -3017 -316
rect -2989 -344 -2951 -316
rect -2923 -344 -2885 -316
rect -2857 -344 -2819 -316
rect -2791 -344 -2753 -316
rect -2725 -344 -2687 -316
rect -2659 -344 -2621 -316
rect -2593 -344 -2555 -316
rect -2527 -344 -2489 -316
rect -2461 -344 -2423 -316
rect -2395 -344 -2357 -316
rect -2329 -344 -2291 -316
rect -2263 -344 -2225 -316
rect -2197 -344 -2159 -316
rect -2131 -344 -2093 -316
rect -2065 -344 -2027 -316
rect -1999 -344 -1961 -316
rect -1933 -344 -1895 -316
rect -1867 -344 -1829 -316
rect -1801 -344 -1763 -316
rect -1735 -344 -1697 -316
rect -1669 -344 -1631 -316
rect -1603 -344 -1565 -316
rect -1537 -344 -1499 -316
rect -1471 -344 -1433 -316
rect -1405 -344 -1367 -316
rect -1339 -344 -1301 -316
rect -1273 -344 -1235 -316
rect -1207 -344 -1169 -316
rect -1141 -344 -1103 -316
rect -1075 -344 -1037 -316
rect -1009 -344 -971 -316
rect -943 -344 -905 -316
rect -877 -344 -839 -316
rect -811 -344 -773 -316
rect -745 -344 -707 -316
rect -679 -344 -641 -316
rect -613 -344 -575 -316
rect -547 -344 -509 -316
rect -481 -344 -443 -316
rect -415 -344 -377 -316
rect -349 -344 -311 -316
rect -283 -344 -245 -316
rect -217 -344 -179 -316
rect -151 -344 -113 -316
rect -85 -344 -47 -316
rect -19 -344 19 -316
rect 47 -344 85 -316
rect 113 -344 151 -316
rect 179 -344 217 -316
rect 245 -344 283 -316
rect 311 -344 349 -316
rect 377 -344 415 -316
rect 443 -344 481 -316
rect 509 -344 547 -316
rect 575 -344 613 -316
rect 641 -344 679 -316
rect 707 -344 745 -316
rect 773 -344 811 -316
rect 839 -344 877 -316
rect 905 -344 943 -316
rect 971 -344 1009 -316
rect 1037 -344 1075 -316
rect 1103 -344 1141 -316
rect 1169 -344 1207 -316
rect 1235 -344 1273 -316
rect 1301 -344 1339 -316
rect 1367 -344 1405 -316
rect 1433 -344 1471 -316
rect 1499 -344 1537 -316
rect 1565 -344 1603 -316
rect 1631 -344 1669 -316
rect 1697 -344 1735 -316
rect 1763 -344 1801 -316
rect 1829 -344 1867 -316
rect 1895 -344 1933 -316
rect 1961 -344 1999 -316
rect 2027 -344 2065 -316
rect 2093 -344 2131 -316
rect 2159 -344 2197 -316
rect 2225 -344 2263 -316
rect 2291 -344 2329 -316
rect 2357 -344 2395 -316
rect 2423 -344 2461 -316
rect 2489 -344 2527 -316
rect 2555 -344 2593 -316
rect 2621 -344 2659 -316
rect 2687 -344 2725 -316
rect 2753 -344 2791 -316
rect 2819 -344 2857 -316
rect 2885 -344 2923 -316
rect 2951 -344 2989 -316
rect 3017 -344 3055 -316
rect 3083 -344 3121 -316
rect 3149 -344 3187 -316
rect 3215 -344 3253 -316
rect 3281 -344 3319 -316
rect 3347 -344 3385 -316
rect 3413 -344 3451 -316
rect 3479 -344 3517 -316
rect 3545 -344 3583 -316
rect 3611 -344 3649 -316
rect 3677 -344 3715 -316
rect 3743 -344 3781 -316
rect 3809 -344 3847 -316
rect 3875 -344 3880 -316
rect -3880 -382 3880 -344
rect -3880 -410 -3875 -382
rect -3847 -410 -3809 -382
rect -3781 -410 -3743 -382
rect -3715 -410 -3677 -382
rect -3649 -410 -3611 -382
rect -3583 -410 -3545 -382
rect -3517 -410 -3479 -382
rect -3451 -410 -3413 -382
rect -3385 -410 -3347 -382
rect -3319 -410 -3281 -382
rect -3253 -410 -3215 -382
rect -3187 -410 -3149 -382
rect -3121 -410 -3083 -382
rect -3055 -410 -3017 -382
rect -2989 -410 -2951 -382
rect -2923 -410 -2885 -382
rect -2857 -410 -2819 -382
rect -2791 -410 -2753 -382
rect -2725 -410 -2687 -382
rect -2659 -410 -2621 -382
rect -2593 -410 -2555 -382
rect -2527 -410 -2489 -382
rect -2461 -410 -2423 -382
rect -2395 -410 -2357 -382
rect -2329 -410 -2291 -382
rect -2263 -410 -2225 -382
rect -2197 -410 -2159 -382
rect -2131 -410 -2093 -382
rect -2065 -410 -2027 -382
rect -1999 -410 -1961 -382
rect -1933 -410 -1895 -382
rect -1867 -410 -1829 -382
rect -1801 -410 -1763 -382
rect -1735 -410 -1697 -382
rect -1669 -410 -1631 -382
rect -1603 -410 -1565 -382
rect -1537 -410 -1499 -382
rect -1471 -410 -1433 -382
rect -1405 -410 -1367 -382
rect -1339 -410 -1301 -382
rect -1273 -410 -1235 -382
rect -1207 -410 -1169 -382
rect -1141 -410 -1103 -382
rect -1075 -410 -1037 -382
rect -1009 -410 -971 -382
rect -943 -410 -905 -382
rect -877 -410 -839 -382
rect -811 -410 -773 -382
rect -745 -410 -707 -382
rect -679 -410 -641 -382
rect -613 -410 -575 -382
rect -547 -410 -509 -382
rect -481 -410 -443 -382
rect -415 -410 -377 -382
rect -349 -410 -311 -382
rect -283 -410 -245 -382
rect -217 -410 -179 -382
rect -151 -410 -113 -382
rect -85 -410 -47 -382
rect -19 -410 19 -382
rect 47 -410 85 -382
rect 113 -410 151 -382
rect 179 -410 217 -382
rect 245 -410 283 -382
rect 311 -410 349 -382
rect 377 -410 415 -382
rect 443 -410 481 -382
rect 509 -410 547 -382
rect 575 -410 613 -382
rect 641 -410 679 -382
rect 707 -410 745 -382
rect 773 -410 811 -382
rect 839 -410 877 -382
rect 905 -410 943 -382
rect 971 -410 1009 -382
rect 1037 -410 1075 -382
rect 1103 -410 1141 -382
rect 1169 -410 1207 -382
rect 1235 -410 1273 -382
rect 1301 -410 1339 -382
rect 1367 -410 1405 -382
rect 1433 -410 1471 -382
rect 1499 -410 1537 -382
rect 1565 -410 1603 -382
rect 1631 -410 1669 -382
rect 1697 -410 1735 -382
rect 1763 -410 1801 -382
rect 1829 -410 1867 -382
rect 1895 -410 1933 -382
rect 1961 -410 1999 -382
rect 2027 -410 2065 -382
rect 2093 -410 2131 -382
rect 2159 -410 2197 -382
rect 2225 -410 2263 -382
rect 2291 -410 2329 -382
rect 2357 -410 2395 -382
rect 2423 -410 2461 -382
rect 2489 -410 2527 -382
rect 2555 -410 2593 -382
rect 2621 -410 2659 -382
rect 2687 -410 2725 -382
rect 2753 -410 2791 -382
rect 2819 -410 2857 -382
rect 2885 -410 2923 -382
rect 2951 -410 2989 -382
rect 3017 -410 3055 -382
rect 3083 -410 3121 -382
rect 3149 -410 3187 -382
rect 3215 -410 3253 -382
rect 3281 -410 3319 -382
rect 3347 -410 3385 -382
rect 3413 -410 3451 -382
rect 3479 -410 3517 -382
rect 3545 -410 3583 -382
rect 3611 -410 3649 -382
rect 3677 -410 3715 -382
rect 3743 -410 3781 -382
rect 3809 -410 3847 -382
rect 3875 -410 3880 -382
rect -3880 -448 3880 -410
rect -3880 -476 -3875 -448
rect -3847 -476 -3809 -448
rect -3781 -476 -3743 -448
rect -3715 -476 -3677 -448
rect -3649 -476 -3611 -448
rect -3583 -476 -3545 -448
rect -3517 -476 -3479 -448
rect -3451 -476 -3413 -448
rect -3385 -476 -3347 -448
rect -3319 -476 -3281 -448
rect -3253 -476 -3215 -448
rect -3187 -476 -3149 -448
rect -3121 -476 -3083 -448
rect -3055 -476 -3017 -448
rect -2989 -476 -2951 -448
rect -2923 -476 -2885 -448
rect -2857 -476 -2819 -448
rect -2791 -476 -2753 -448
rect -2725 -476 -2687 -448
rect -2659 -476 -2621 -448
rect -2593 -476 -2555 -448
rect -2527 -476 -2489 -448
rect -2461 -476 -2423 -448
rect -2395 -476 -2357 -448
rect -2329 -476 -2291 -448
rect -2263 -476 -2225 -448
rect -2197 -476 -2159 -448
rect -2131 -476 -2093 -448
rect -2065 -476 -2027 -448
rect -1999 -476 -1961 -448
rect -1933 -476 -1895 -448
rect -1867 -476 -1829 -448
rect -1801 -476 -1763 -448
rect -1735 -476 -1697 -448
rect -1669 -476 -1631 -448
rect -1603 -476 -1565 -448
rect -1537 -476 -1499 -448
rect -1471 -476 -1433 -448
rect -1405 -476 -1367 -448
rect -1339 -476 -1301 -448
rect -1273 -476 -1235 -448
rect -1207 -476 -1169 -448
rect -1141 -476 -1103 -448
rect -1075 -476 -1037 -448
rect -1009 -476 -971 -448
rect -943 -476 -905 -448
rect -877 -476 -839 -448
rect -811 -476 -773 -448
rect -745 -476 -707 -448
rect -679 -476 -641 -448
rect -613 -476 -575 -448
rect -547 -476 -509 -448
rect -481 -476 -443 -448
rect -415 -476 -377 -448
rect -349 -476 -311 -448
rect -283 -476 -245 -448
rect -217 -476 -179 -448
rect -151 -476 -113 -448
rect -85 -476 -47 -448
rect -19 -476 19 -448
rect 47 -476 85 -448
rect 113 -476 151 -448
rect 179 -476 217 -448
rect 245 -476 283 -448
rect 311 -476 349 -448
rect 377 -476 415 -448
rect 443 -476 481 -448
rect 509 -476 547 -448
rect 575 -476 613 -448
rect 641 -476 679 -448
rect 707 -476 745 -448
rect 773 -476 811 -448
rect 839 -476 877 -448
rect 905 -476 943 -448
rect 971 -476 1009 -448
rect 1037 -476 1075 -448
rect 1103 -476 1141 -448
rect 1169 -476 1207 -448
rect 1235 -476 1273 -448
rect 1301 -476 1339 -448
rect 1367 -476 1405 -448
rect 1433 -476 1471 -448
rect 1499 -476 1537 -448
rect 1565 -476 1603 -448
rect 1631 -476 1669 -448
rect 1697 -476 1735 -448
rect 1763 -476 1801 -448
rect 1829 -476 1867 -448
rect 1895 -476 1933 -448
rect 1961 -476 1999 -448
rect 2027 -476 2065 -448
rect 2093 -476 2131 -448
rect 2159 -476 2197 -448
rect 2225 -476 2263 -448
rect 2291 -476 2329 -448
rect 2357 -476 2395 -448
rect 2423 -476 2461 -448
rect 2489 -476 2527 -448
rect 2555 -476 2593 -448
rect 2621 -476 2659 -448
rect 2687 -476 2725 -448
rect 2753 -476 2791 -448
rect 2819 -476 2857 -448
rect 2885 -476 2923 -448
rect 2951 -476 2989 -448
rect 3017 -476 3055 -448
rect 3083 -476 3121 -448
rect 3149 -476 3187 -448
rect 3215 -476 3253 -448
rect 3281 -476 3319 -448
rect 3347 -476 3385 -448
rect 3413 -476 3451 -448
rect 3479 -476 3517 -448
rect 3545 -476 3583 -448
rect 3611 -476 3649 -448
rect 3677 -476 3715 -448
rect 3743 -476 3781 -448
rect 3809 -476 3847 -448
rect 3875 -476 3880 -448
rect -3880 -514 3880 -476
rect -3880 -542 -3875 -514
rect -3847 -542 -3809 -514
rect -3781 -542 -3743 -514
rect -3715 -542 -3677 -514
rect -3649 -542 -3611 -514
rect -3583 -542 -3545 -514
rect -3517 -542 -3479 -514
rect -3451 -542 -3413 -514
rect -3385 -542 -3347 -514
rect -3319 -542 -3281 -514
rect -3253 -542 -3215 -514
rect -3187 -542 -3149 -514
rect -3121 -542 -3083 -514
rect -3055 -542 -3017 -514
rect -2989 -542 -2951 -514
rect -2923 -542 -2885 -514
rect -2857 -542 -2819 -514
rect -2791 -542 -2753 -514
rect -2725 -542 -2687 -514
rect -2659 -542 -2621 -514
rect -2593 -542 -2555 -514
rect -2527 -542 -2489 -514
rect -2461 -542 -2423 -514
rect -2395 -542 -2357 -514
rect -2329 -542 -2291 -514
rect -2263 -542 -2225 -514
rect -2197 -542 -2159 -514
rect -2131 -542 -2093 -514
rect -2065 -542 -2027 -514
rect -1999 -542 -1961 -514
rect -1933 -542 -1895 -514
rect -1867 -542 -1829 -514
rect -1801 -542 -1763 -514
rect -1735 -542 -1697 -514
rect -1669 -542 -1631 -514
rect -1603 -542 -1565 -514
rect -1537 -542 -1499 -514
rect -1471 -542 -1433 -514
rect -1405 -542 -1367 -514
rect -1339 -542 -1301 -514
rect -1273 -542 -1235 -514
rect -1207 -542 -1169 -514
rect -1141 -542 -1103 -514
rect -1075 -542 -1037 -514
rect -1009 -542 -971 -514
rect -943 -542 -905 -514
rect -877 -542 -839 -514
rect -811 -542 -773 -514
rect -745 -542 -707 -514
rect -679 -542 -641 -514
rect -613 -542 -575 -514
rect -547 -542 -509 -514
rect -481 -542 -443 -514
rect -415 -542 -377 -514
rect -349 -542 -311 -514
rect -283 -542 -245 -514
rect -217 -542 -179 -514
rect -151 -542 -113 -514
rect -85 -542 -47 -514
rect -19 -542 19 -514
rect 47 -542 85 -514
rect 113 -542 151 -514
rect 179 -542 217 -514
rect 245 -542 283 -514
rect 311 -542 349 -514
rect 377 -542 415 -514
rect 443 -542 481 -514
rect 509 -542 547 -514
rect 575 -542 613 -514
rect 641 -542 679 -514
rect 707 -542 745 -514
rect 773 -542 811 -514
rect 839 -542 877 -514
rect 905 -542 943 -514
rect 971 -542 1009 -514
rect 1037 -542 1075 -514
rect 1103 -542 1141 -514
rect 1169 -542 1207 -514
rect 1235 -542 1273 -514
rect 1301 -542 1339 -514
rect 1367 -542 1405 -514
rect 1433 -542 1471 -514
rect 1499 -542 1537 -514
rect 1565 -542 1603 -514
rect 1631 -542 1669 -514
rect 1697 -542 1735 -514
rect 1763 -542 1801 -514
rect 1829 -542 1867 -514
rect 1895 -542 1933 -514
rect 1961 -542 1999 -514
rect 2027 -542 2065 -514
rect 2093 -542 2131 -514
rect 2159 -542 2197 -514
rect 2225 -542 2263 -514
rect 2291 -542 2329 -514
rect 2357 -542 2395 -514
rect 2423 -542 2461 -514
rect 2489 -542 2527 -514
rect 2555 -542 2593 -514
rect 2621 -542 2659 -514
rect 2687 -542 2725 -514
rect 2753 -542 2791 -514
rect 2819 -542 2857 -514
rect 2885 -542 2923 -514
rect 2951 -542 2989 -514
rect 3017 -542 3055 -514
rect 3083 -542 3121 -514
rect 3149 -542 3187 -514
rect 3215 -542 3253 -514
rect 3281 -542 3319 -514
rect 3347 -542 3385 -514
rect 3413 -542 3451 -514
rect 3479 -542 3517 -514
rect 3545 -542 3583 -514
rect 3611 -542 3649 -514
rect 3677 -542 3715 -514
rect 3743 -542 3781 -514
rect 3809 -542 3847 -514
rect 3875 -542 3880 -514
rect -3880 -580 3880 -542
rect -3880 -608 -3875 -580
rect -3847 -608 -3809 -580
rect -3781 -608 -3743 -580
rect -3715 -608 -3677 -580
rect -3649 -608 -3611 -580
rect -3583 -608 -3545 -580
rect -3517 -608 -3479 -580
rect -3451 -608 -3413 -580
rect -3385 -608 -3347 -580
rect -3319 -608 -3281 -580
rect -3253 -608 -3215 -580
rect -3187 -608 -3149 -580
rect -3121 -608 -3083 -580
rect -3055 -608 -3017 -580
rect -2989 -608 -2951 -580
rect -2923 -608 -2885 -580
rect -2857 -608 -2819 -580
rect -2791 -608 -2753 -580
rect -2725 -608 -2687 -580
rect -2659 -608 -2621 -580
rect -2593 -608 -2555 -580
rect -2527 -608 -2489 -580
rect -2461 -608 -2423 -580
rect -2395 -608 -2357 -580
rect -2329 -608 -2291 -580
rect -2263 -608 -2225 -580
rect -2197 -608 -2159 -580
rect -2131 -608 -2093 -580
rect -2065 -608 -2027 -580
rect -1999 -608 -1961 -580
rect -1933 -608 -1895 -580
rect -1867 -608 -1829 -580
rect -1801 -608 -1763 -580
rect -1735 -608 -1697 -580
rect -1669 -608 -1631 -580
rect -1603 -608 -1565 -580
rect -1537 -608 -1499 -580
rect -1471 -608 -1433 -580
rect -1405 -608 -1367 -580
rect -1339 -608 -1301 -580
rect -1273 -608 -1235 -580
rect -1207 -608 -1169 -580
rect -1141 -608 -1103 -580
rect -1075 -608 -1037 -580
rect -1009 -608 -971 -580
rect -943 -608 -905 -580
rect -877 -608 -839 -580
rect -811 -608 -773 -580
rect -745 -608 -707 -580
rect -679 -608 -641 -580
rect -613 -608 -575 -580
rect -547 -608 -509 -580
rect -481 -608 -443 -580
rect -415 -608 -377 -580
rect -349 -608 -311 -580
rect -283 -608 -245 -580
rect -217 -608 -179 -580
rect -151 -608 -113 -580
rect -85 -608 -47 -580
rect -19 -608 19 -580
rect 47 -608 85 -580
rect 113 -608 151 -580
rect 179 -608 217 -580
rect 245 -608 283 -580
rect 311 -608 349 -580
rect 377 -608 415 -580
rect 443 -608 481 -580
rect 509 -608 547 -580
rect 575 -608 613 -580
rect 641 -608 679 -580
rect 707 -608 745 -580
rect 773 -608 811 -580
rect 839 -608 877 -580
rect 905 -608 943 -580
rect 971 -608 1009 -580
rect 1037 -608 1075 -580
rect 1103 -608 1141 -580
rect 1169 -608 1207 -580
rect 1235 -608 1273 -580
rect 1301 -608 1339 -580
rect 1367 -608 1405 -580
rect 1433 -608 1471 -580
rect 1499 -608 1537 -580
rect 1565 -608 1603 -580
rect 1631 -608 1669 -580
rect 1697 -608 1735 -580
rect 1763 -608 1801 -580
rect 1829 -608 1867 -580
rect 1895 -608 1933 -580
rect 1961 -608 1999 -580
rect 2027 -608 2065 -580
rect 2093 -608 2131 -580
rect 2159 -608 2197 -580
rect 2225 -608 2263 -580
rect 2291 -608 2329 -580
rect 2357 -608 2395 -580
rect 2423 -608 2461 -580
rect 2489 -608 2527 -580
rect 2555 -608 2593 -580
rect 2621 -608 2659 -580
rect 2687 -608 2725 -580
rect 2753 -608 2791 -580
rect 2819 -608 2857 -580
rect 2885 -608 2923 -580
rect 2951 -608 2989 -580
rect 3017 -608 3055 -580
rect 3083 -608 3121 -580
rect 3149 -608 3187 -580
rect 3215 -608 3253 -580
rect 3281 -608 3319 -580
rect 3347 -608 3385 -580
rect 3413 -608 3451 -580
rect 3479 -608 3517 -580
rect 3545 -608 3583 -580
rect 3611 -608 3649 -580
rect 3677 -608 3715 -580
rect 3743 -608 3781 -580
rect 3809 -608 3847 -580
rect 3875 -608 3880 -580
rect -3880 -646 3880 -608
rect -3880 -674 -3875 -646
rect -3847 -674 -3809 -646
rect -3781 -674 -3743 -646
rect -3715 -674 -3677 -646
rect -3649 -674 -3611 -646
rect -3583 -674 -3545 -646
rect -3517 -674 -3479 -646
rect -3451 -674 -3413 -646
rect -3385 -674 -3347 -646
rect -3319 -674 -3281 -646
rect -3253 -674 -3215 -646
rect -3187 -674 -3149 -646
rect -3121 -674 -3083 -646
rect -3055 -674 -3017 -646
rect -2989 -674 -2951 -646
rect -2923 -674 -2885 -646
rect -2857 -674 -2819 -646
rect -2791 -674 -2753 -646
rect -2725 -674 -2687 -646
rect -2659 -674 -2621 -646
rect -2593 -674 -2555 -646
rect -2527 -674 -2489 -646
rect -2461 -674 -2423 -646
rect -2395 -674 -2357 -646
rect -2329 -674 -2291 -646
rect -2263 -674 -2225 -646
rect -2197 -674 -2159 -646
rect -2131 -674 -2093 -646
rect -2065 -674 -2027 -646
rect -1999 -674 -1961 -646
rect -1933 -674 -1895 -646
rect -1867 -674 -1829 -646
rect -1801 -674 -1763 -646
rect -1735 -674 -1697 -646
rect -1669 -674 -1631 -646
rect -1603 -674 -1565 -646
rect -1537 -674 -1499 -646
rect -1471 -674 -1433 -646
rect -1405 -674 -1367 -646
rect -1339 -674 -1301 -646
rect -1273 -674 -1235 -646
rect -1207 -674 -1169 -646
rect -1141 -674 -1103 -646
rect -1075 -674 -1037 -646
rect -1009 -674 -971 -646
rect -943 -674 -905 -646
rect -877 -674 -839 -646
rect -811 -674 -773 -646
rect -745 -674 -707 -646
rect -679 -674 -641 -646
rect -613 -674 -575 -646
rect -547 -674 -509 -646
rect -481 -674 -443 -646
rect -415 -674 -377 -646
rect -349 -674 -311 -646
rect -283 -674 -245 -646
rect -217 -674 -179 -646
rect -151 -674 -113 -646
rect -85 -674 -47 -646
rect -19 -674 19 -646
rect 47 -674 85 -646
rect 113 -674 151 -646
rect 179 -674 217 -646
rect 245 -674 283 -646
rect 311 -674 349 -646
rect 377 -674 415 -646
rect 443 -674 481 -646
rect 509 -674 547 -646
rect 575 -674 613 -646
rect 641 -674 679 -646
rect 707 -674 745 -646
rect 773 -674 811 -646
rect 839 -674 877 -646
rect 905 -674 943 -646
rect 971 -674 1009 -646
rect 1037 -674 1075 -646
rect 1103 -674 1141 -646
rect 1169 -674 1207 -646
rect 1235 -674 1273 -646
rect 1301 -674 1339 -646
rect 1367 -674 1405 -646
rect 1433 -674 1471 -646
rect 1499 -674 1537 -646
rect 1565 -674 1603 -646
rect 1631 -674 1669 -646
rect 1697 -674 1735 -646
rect 1763 -674 1801 -646
rect 1829 -674 1867 -646
rect 1895 -674 1933 -646
rect 1961 -674 1999 -646
rect 2027 -674 2065 -646
rect 2093 -674 2131 -646
rect 2159 -674 2197 -646
rect 2225 -674 2263 -646
rect 2291 -674 2329 -646
rect 2357 -674 2395 -646
rect 2423 -674 2461 -646
rect 2489 -674 2527 -646
rect 2555 -674 2593 -646
rect 2621 -674 2659 -646
rect 2687 -674 2725 -646
rect 2753 -674 2791 -646
rect 2819 -674 2857 -646
rect 2885 -674 2923 -646
rect 2951 -674 2989 -646
rect 3017 -674 3055 -646
rect 3083 -674 3121 -646
rect 3149 -674 3187 -646
rect 3215 -674 3253 -646
rect 3281 -674 3319 -646
rect 3347 -674 3385 -646
rect 3413 -674 3451 -646
rect 3479 -674 3517 -646
rect 3545 -674 3583 -646
rect 3611 -674 3649 -646
rect 3677 -674 3715 -646
rect 3743 -674 3781 -646
rect 3809 -674 3847 -646
rect 3875 -674 3880 -646
rect -3880 -712 3880 -674
rect -3880 -740 -3875 -712
rect -3847 -740 -3809 -712
rect -3781 -740 -3743 -712
rect -3715 -740 -3677 -712
rect -3649 -740 -3611 -712
rect -3583 -740 -3545 -712
rect -3517 -740 -3479 -712
rect -3451 -740 -3413 -712
rect -3385 -740 -3347 -712
rect -3319 -740 -3281 -712
rect -3253 -740 -3215 -712
rect -3187 -740 -3149 -712
rect -3121 -740 -3083 -712
rect -3055 -740 -3017 -712
rect -2989 -740 -2951 -712
rect -2923 -740 -2885 -712
rect -2857 -740 -2819 -712
rect -2791 -740 -2753 -712
rect -2725 -740 -2687 -712
rect -2659 -740 -2621 -712
rect -2593 -740 -2555 -712
rect -2527 -740 -2489 -712
rect -2461 -740 -2423 -712
rect -2395 -740 -2357 -712
rect -2329 -740 -2291 -712
rect -2263 -740 -2225 -712
rect -2197 -740 -2159 -712
rect -2131 -740 -2093 -712
rect -2065 -740 -2027 -712
rect -1999 -740 -1961 -712
rect -1933 -740 -1895 -712
rect -1867 -740 -1829 -712
rect -1801 -740 -1763 -712
rect -1735 -740 -1697 -712
rect -1669 -740 -1631 -712
rect -1603 -740 -1565 -712
rect -1537 -740 -1499 -712
rect -1471 -740 -1433 -712
rect -1405 -740 -1367 -712
rect -1339 -740 -1301 -712
rect -1273 -740 -1235 -712
rect -1207 -740 -1169 -712
rect -1141 -740 -1103 -712
rect -1075 -740 -1037 -712
rect -1009 -740 -971 -712
rect -943 -740 -905 -712
rect -877 -740 -839 -712
rect -811 -740 -773 -712
rect -745 -740 -707 -712
rect -679 -740 -641 -712
rect -613 -740 -575 -712
rect -547 -740 -509 -712
rect -481 -740 -443 -712
rect -415 -740 -377 -712
rect -349 -740 -311 -712
rect -283 -740 -245 -712
rect -217 -740 -179 -712
rect -151 -740 -113 -712
rect -85 -740 -47 -712
rect -19 -740 19 -712
rect 47 -740 85 -712
rect 113 -740 151 -712
rect 179 -740 217 -712
rect 245 -740 283 -712
rect 311 -740 349 -712
rect 377 -740 415 -712
rect 443 -740 481 -712
rect 509 -740 547 -712
rect 575 -740 613 -712
rect 641 -740 679 -712
rect 707 -740 745 -712
rect 773 -740 811 -712
rect 839 -740 877 -712
rect 905 -740 943 -712
rect 971 -740 1009 -712
rect 1037 -740 1075 -712
rect 1103 -740 1141 -712
rect 1169 -740 1207 -712
rect 1235 -740 1273 -712
rect 1301 -740 1339 -712
rect 1367 -740 1405 -712
rect 1433 -740 1471 -712
rect 1499 -740 1537 -712
rect 1565 -740 1603 -712
rect 1631 -740 1669 -712
rect 1697 -740 1735 -712
rect 1763 -740 1801 -712
rect 1829 -740 1867 -712
rect 1895 -740 1933 -712
rect 1961 -740 1999 -712
rect 2027 -740 2065 -712
rect 2093 -740 2131 -712
rect 2159 -740 2197 -712
rect 2225 -740 2263 -712
rect 2291 -740 2329 -712
rect 2357 -740 2395 -712
rect 2423 -740 2461 -712
rect 2489 -740 2527 -712
rect 2555 -740 2593 -712
rect 2621 -740 2659 -712
rect 2687 -740 2725 -712
rect 2753 -740 2791 -712
rect 2819 -740 2857 -712
rect 2885 -740 2923 -712
rect 2951 -740 2989 -712
rect 3017 -740 3055 -712
rect 3083 -740 3121 -712
rect 3149 -740 3187 -712
rect 3215 -740 3253 -712
rect 3281 -740 3319 -712
rect 3347 -740 3385 -712
rect 3413 -740 3451 -712
rect 3479 -740 3517 -712
rect 3545 -740 3583 -712
rect 3611 -740 3649 -712
rect 3677 -740 3715 -712
rect 3743 -740 3781 -712
rect 3809 -740 3847 -712
rect 3875 -740 3880 -712
rect -3880 -745 3880 -740
<< via4 >>
rect -3875 712 -3847 740
rect -3809 712 -3781 740
rect -3743 712 -3715 740
rect -3677 712 -3649 740
rect -3611 712 -3583 740
rect -3545 712 -3517 740
rect -3479 712 -3451 740
rect -3413 712 -3385 740
rect -3347 712 -3319 740
rect -3281 712 -3253 740
rect -3215 712 -3187 740
rect -3149 712 -3121 740
rect -3083 712 -3055 740
rect -3017 712 -2989 740
rect -2951 712 -2923 740
rect -2885 712 -2857 740
rect -2819 712 -2791 740
rect -2753 712 -2725 740
rect -2687 712 -2659 740
rect -2621 712 -2593 740
rect -2555 712 -2527 740
rect -2489 712 -2461 740
rect -2423 712 -2395 740
rect -2357 712 -2329 740
rect -2291 712 -2263 740
rect -2225 712 -2197 740
rect -2159 712 -2131 740
rect -2093 712 -2065 740
rect -2027 712 -1999 740
rect -1961 712 -1933 740
rect -1895 712 -1867 740
rect -1829 712 -1801 740
rect -1763 712 -1735 740
rect -1697 712 -1669 740
rect -1631 712 -1603 740
rect -1565 712 -1537 740
rect -1499 712 -1471 740
rect -1433 712 -1405 740
rect -1367 712 -1339 740
rect -1301 712 -1273 740
rect -1235 712 -1207 740
rect -1169 712 -1141 740
rect -1103 712 -1075 740
rect -1037 712 -1009 740
rect -971 712 -943 740
rect -905 712 -877 740
rect -839 712 -811 740
rect -773 712 -745 740
rect -707 712 -679 740
rect -641 712 -613 740
rect -575 712 -547 740
rect -509 712 -481 740
rect -443 712 -415 740
rect -377 712 -349 740
rect -311 712 -283 740
rect -245 712 -217 740
rect -179 712 -151 740
rect -113 712 -85 740
rect -47 712 -19 740
rect 19 712 47 740
rect 85 712 113 740
rect 151 712 179 740
rect 217 712 245 740
rect 283 712 311 740
rect 349 712 377 740
rect 415 712 443 740
rect 481 712 509 740
rect 547 712 575 740
rect 613 712 641 740
rect 679 712 707 740
rect 745 712 773 740
rect 811 712 839 740
rect 877 712 905 740
rect 943 712 971 740
rect 1009 712 1037 740
rect 1075 712 1103 740
rect 1141 712 1169 740
rect 1207 712 1235 740
rect 1273 712 1301 740
rect 1339 712 1367 740
rect 1405 712 1433 740
rect 1471 712 1499 740
rect 1537 712 1565 740
rect 1603 712 1631 740
rect 1669 712 1697 740
rect 1735 712 1763 740
rect 1801 712 1829 740
rect 1867 712 1895 740
rect 1933 712 1961 740
rect 1999 712 2027 740
rect 2065 712 2093 740
rect 2131 712 2159 740
rect 2197 712 2225 740
rect 2263 712 2291 740
rect 2329 712 2357 740
rect 2395 712 2423 740
rect 2461 712 2489 740
rect 2527 712 2555 740
rect 2593 712 2621 740
rect 2659 712 2687 740
rect 2725 712 2753 740
rect 2791 712 2819 740
rect 2857 712 2885 740
rect 2923 712 2951 740
rect 2989 712 3017 740
rect 3055 712 3083 740
rect 3121 712 3149 740
rect 3187 712 3215 740
rect 3253 712 3281 740
rect 3319 712 3347 740
rect 3385 712 3413 740
rect 3451 712 3479 740
rect 3517 712 3545 740
rect 3583 712 3611 740
rect 3649 712 3677 740
rect 3715 712 3743 740
rect 3781 712 3809 740
rect 3847 712 3875 740
rect -3875 646 -3847 674
rect -3809 646 -3781 674
rect -3743 646 -3715 674
rect -3677 646 -3649 674
rect -3611 646 -3583 674
rect -3545 646 -3517 674
rect -3479 646 -3451 674
rect -3413 646 -3385 674
rect -3347 646 -3319 674
rect -3281 646 -3253 674
rect -3215 646 -3187 674
rect -3149 646 -3121 674
rect -3083 646 -3055 674
rect -3017 646 -2989 674
rect -2951 646 -2923 674
rect -2885 646 -2857 674
rect -2819 646 -2791 674
rect -2753 646 -2725 674
rect -2687 646 -2659 674
rect -2621 646 -2593 674
rect -2555 646 -2527 674
rect -2489 646 -2461 674
rect -2423 646 -2395 674
rect -2357 646 -2329 674
rect -2291 646 -2263 674
rect -2225 646 -2197 674
rect -2159 646 -2131 674
rect -2093 646 -2065 674
rect -2027 646 -1999 674
rect -1961 646 -1933 674
rect -1895 646 -1867 674
rect -1829 646 -1801 674
rect -1763 646 -1735 674
rect -1697 646 -1669 674
rect -1631 646 -1603 674
rect -1565 646 -1537 674
rect -1499 646 -1471 674
rect -1433 646 -1405 674
rect -1367 646 -1339 674
rect -1301 646 -1273 674
rect -1235 646 -1207 674
rect -1169 646 -1141 674
rect -1103 646 -1075 674
rect -1037 646 -1009 674
rect -971 646 -943 674
rect -905 646 -877 674
rect -839 646 -811 674
rect -773 646 -745 674
rect -707 646 -679 674
rect -641 646 -613 674
rect -575 646 -547 674
rect -509 646 -481 674
rect -443 646 -415 674
rect -377 646 -349 674
rect -311 646 -283 674
rect -245 646 -217 674
rect -179 646 -151 674
rect -113 646 -85 674
rect -47 646 -19 674
rect 19 646 47 674
rect 85 646 113 674
rect 151 646 179 674
rect 217 646 245 674
rect 283 646 311 674
rect 349 646 377 674
rect 415 646 443 674
rect 481 646 509 674
rect 547 646 575 674
rect 613 646 641 674
rect 679 646 707 674
rect 745 646 773 674
rect 811 646 839 674
rect 877 646 905 674
rect 943 646 971 674
rect 1009 646 1037 674
rect 1075 646 1103 674
rect 1141 646 1169 674
rect 1207 646 1235 674
rect 1273 646 1301 674
rect 1339 646 1367 674
rect 1405 646 1433 674
rect 1471 646 1499 674
rect 1537 646 1565 674
rect 1603 646 1631 674
rect 1669 646 1697 674
rect 1735 646 1763 674
rect 1801 646 1829 674
rect 1867 646 1895 674
rect 1933 646 1961 674
rect 1999 646 2027 674
rect 2065 646 2093 674
rect 2131 646 2159 674
rect 2197 646 2225 674
rect 2263 646 2291 674
rect 2329 646 2357 674
rect 2395 646 2423 674
rect 2461 646 2489 674
rect 2527 646 2555 674
rect 2593 646 2621 674
rect 2659 646 2687 674
rect 2725 646 2753 674
rect 2791 646 2819 674
rect 2857 646 2885 674
rect 2923 646 2951 674
rect 2989 646 3017 674
rect 3055 646 3083 674
rect 3121 646 3149 674
rect 3187 646 3215 674
rect 3253 646 3281 674
rect 3319 646 3347 674
rect 3385 646 3413 674
rect 3451 646 3479 674
rect 3517 646 3545 674
rect 3583 646 3611 674
rect 3649 646 3677 674
rect 3715 646 3743 674
rect 3781 646 3809 674
rect 3847 646 3875 674
rect -3875 580 -3847 608
rect -3809 580 -3781 608
rect -3743 580 -3715 608
rect -3677 580 -3649 608
rect -3611 580 -3583 608
rect -3545 580 -3517 608
rect -3479 580 -3451 608
rect -3413 580 -3385 608
rect -3347 580 -3319 608
rect -3281 580 -3253 608
rect -3215 580 -3187 608
rect -3149 580 -3121 608
rect -3083 580 -3055 608
rect -3017 580 -2989 608
rect -2951 580 -2923 608
rect -2885 580 -2857 608
rect -2819 580 -2791 608
rect -2753 580 -2725 608
rect -2687 580 -2659 608
rect -2621 580 -2593 608
rect -2555 580 -2527 608
rect -2489 580 -2461 608
rect -2423 580 -2395 608
rect -2357 580 -2329 608
rect -2291 580 -2263 608
rect -2225 580 -2197 608
rect -2159 580 -2131 608
rect -2093 580 -2065 608
rect -2027 580 -1999 608
rect -1961 580 -1933 608
rect -1895 580 -1867 608
rect -1829 580 -1801 608
rect -1763 580 -1735 608
rect -1697 580 -1669 608
rect -1631 580 -1603 608
rect -1565 580 -1537 608
rect -1499 580 -1471 608
rect -1433 580 -1405 608
rect -1367 580 -1339 608
rect -1301 580 -1273 608
rect -1235 580 -1207 608
rect -1169 580 -1141 608
rect -1103 580 -1075 608
rect -1037 580 -1009 608
rect -971 580 -943 608
rect -905 580 -877 608
rect -839 580 -811 608
rect -773 580 -745 608
rect -707 580 -679 608
rect -641 580 -613 608
rect -575 580 -547 608
rect -509 580 -481 608
rect -443 580 -415 608
rect -377 580 -349 608
rect -311 580 -283 608
rect -245 580 -217 608
rect -179 580 -151 608
rect -113 580 -85 608
rect -47 580 -19 608
rect 19 580 47 608
rect 85 580 113 608
rect 151 580 179 608
rect 217 580 245 608
rect 283 580 311 608
rect 349 580 377 608
rect 415 580 443 608
rect 481 580 509 608
rect 547 580 575 608
rect 613 580 641 608
rect 679 580 707 608
rect 745 580 773 608
rect 811 580 839 608
rect 877 580 905 608
rect 943 580 971 608
rect 1009 580 1037 608
rect 1075 580 1103 608
rect 1141 580 1169 608
rect 1207 580 1235 608
rect 1273 580 1301 608
rect 1339 580 1367 608
rect 1405 580 1433 608
rect 1471 580 1499 608
rect 1537 580 1565 608
rect 1603 580 1631 608
rect 1669 580 1697 608
rect 1735 580 1763 608
rect 1801 580 1829 608
rect 1867 580 1895 608
rect 1933 580 1961 608
rect 1999 580 2027 608
rect 2065 580 2093 608
rect 2131 580 2159 608
rect 2197 580 2225 608
rect 2263 580 2291 608
rect 2329 580 2357 608
rect 2395 580 2423 608
rect 2461 580 2489 608
rect 2527 580 2555 608
rect 2593 580 2621 608
rect 2659 580 2687 608
rect 2725 580 2753 608
rect 2791 580 2819 608
rect 2857 580 2885 608
rect 2923 580 2951 608
rect 2989 580 3017 608
rect 3055 580 3083 608
rect 3121 580 3149 608
rect 3187 580 3215 608
rect 3253 580 3281 608
rect 3319 580 3347 608
rect 3385 580 3413 608
rect 3451 580 3479 608
rect 3517 580 3545 608
rect 3583 580 3611 608
rect 3649 580 3677 608
rect 3715 580 3743 608
rect 3781 580 3809 608
rect 3847 580 3875 608
rect -3875 514 -3847 542
rect -3809 514 -3781 542
rect -3743 514 -3715 542
rect -3677 514 -3649 542
rect -3611 514 -3583 542
rect -3545 514 -3517 542
rect -3479 514 -3451 542
rect -3413 514 -3385 542
rect -3347 514 -3319 542
rect -3281 514 -3253 542
rect -3215 514 -3187 542
rect -3149 514 -3121 542
rect -3083 514 -3055 542
rect -3017 514 -2989 542
rect -2951 514 -2923 542
rect -2885 514 -2857 542
rect -2819 514 -2791 542
rect -2753 514 -2725 542
rect -2687 514 -2659 542
rect -2621 514 -2593 542
rect -2555 514 -2527 542
rect -2489 514 -2461 542
rect -2423 514 -2395 542
rect -2357 514 -2329 542
rect -2291 514 -2263 542
rect -2225 514 -2197 542
rect -2159 514 -2131 542
rect -2093 514 -2065 542
rect -2027 514 -1999 542
rect -1961 514 -1933 542
rect -1895 514 -1867 542
rect -1829 514 -1801 542
rect -1763 514 -1735 542
rect -1697 514 -1669 542
rect -1631 514 -1603 542
rect -1565 514 -1537 542
rect -1499 514 -1471 542
rect -1433 514 -1405 542
rect -1367 514 -1339 542
rect -1301 514 -1273 542
rect -1235 514 -1207 542
rect -1169 514 -1141 542
rect -1103 514 -1075 542
rect -1037 514 -1009 542
rect -971 514 -943 542
rect -905 514 -877 542
rect -839 514 -811 542
rect -773 514 -745 542
rect -707 514 -679 542
rect -641 514 -613 542
rect -575 514 -547 542
rect -509 514 -481 542
rect -443 514 -415 542
rect -377 514 -349 542
rect -311 514 -283 542
rect -245 514 -217 542
rect -179 514 -151 542
rect -113 514 -85 542
rect -47 514 -19 542
rect 19 514 47 542
rect 85 514 113 542
rect 151 514 179 542
rect 217 514 245 542
rect 283 514 311 542
rect 349 514 377 542
rect 415 514 443 542
rect 481 514 509 542
rect 547 514 575 542
rect 613 514 641 542
rect 679 514 707 542
rect 745 514 773 542
rect 811 514 839 542
rect 877 514 905 542
rect 943 514 971 542
rect 1009 514 1037 542
rect 1075 514 1103 542
rect 1141 514 1169 542
rect 1207 514 1235 542
rect 1273 514 1301 542
rect 1339 514 1367 542
rect 1405 514 1433 542
rect 1471 514 1499 542
rect 1537 514 1565 542
rect 1603 514 1631 542
rect 1669 514 1697 542
rect 1735 514 1763 542
rect 1801 514 1829 542
rect 1867 514 1895 542
rect 1933 514 1961 542
rect 1999 514 2027 542
rect 2065 514 2093 542
rect 2131 514 2159 542
rect 2197 514 2225 542
rect 2263 514 2291 542
rect 2329 514 2357 542
rect 2395 514 2423 542
rect 2461 514 2489 542
rect 2527 514 2555 542
rect 2593 514 2621 542
rect 2659 514 2687 542
rect 2725 514 2753 542
rect 2791 514 2819 542
rect 2857 514 2885 542
rect 2923 514 2951 542
rect 2989 514 3017 542
rect 3055 514 3083 542
rect 3121 514 3149 542
rect 3187 514 3215 542
rect 3253 514 3281 542
rect 3319 514 3347 542
rect 3385 514 3413 542
rect 3451 514 3479 542
rect 3517 514 3545 542
rect 3583 514 3611 542
rect 3649 514 3677 542
rect 3715 514 3743 542
rect 3781 514 3809 542
rect 3847 514 3875 542
rect -3875 448 -3847 476
rect -3809 448 -3781 476
rect -3743 448 -3715 476
rect -3677 448 -3649 476
rect -3611 448 -3583 476
rect -3545 448 -3517 476
rect -3479 448 -3451 476
rect -3413 448 -3385 476
rect -3347 448 -3319 476
rect -3281 448 -3253 476
rect -3215 448 -3187 476
rect -3149 448 -3121 476
rect -3083 448 -3055 476
rect -3017 448 -2989 476
rect -2951 448 -2923 476
rect -2885 448 -2857 476
rect -2819 448 -2791 476
rect -2753 448 -2725 476
rect -2687 448 -2659 476
rect -2621 448 -2593 476
rect -2555 448 -2527 476
rect -2489 448 -2461 476
rect -2423 448 -2395 476
rect -2357 448 -2329 476
rect -2291 448 -2263 476
rect -2225 448 -2197 476
rect -2159 448 -2131 476
rect -2093 448 -2065 476
rect -2027 448 -1999 476
rect -1961 448 -1933 476
rect -1895 448 -1867 476
rect -1829 448 -1801 476
rect -1763 448 -1735 476
rect -1697 448 -1669 476
rect -1631 448 -1603 476
rect -1565 448 -1537 476
rect -1499 448 -1471 476
rect -1433 448 -1405 476
rect -1367 448 -1339 476
rect -1301 448 -1273 476
rect -1235 448 -1207 476
rect -1169 448 -1141 476
rect -1103 448 -1075 476
rect -1037 448 -1009 476
rect -971 448 -943 476
rect -905 448 -877 476
rect -839 448 -811 476
rect -773 448 -745 476
rect -707 448 -679 476
rect -641 448 -613 476
rect -575 448 -547 476
rect -509 448 -481 476
rect -443 448 -415 476
rect -377 448 -349 476
rect -311 448 -283 476
rect -245 448 -217 476
rect -179 448 -151 476
rect -113 448 -85 476
rect -47 448 -19 476
rect 19 448 47 476
rect 85 448 113 476
rect 151 448 179 476
rect 217 448 245 476
rect 283 448 311 476
rect 349 448 377 476
rect 415 448 443 476
rect 481 448 509 476
rect 547 448 575 476
rect 613 448 641 476
rect 679 448 707 476
rect 745 448 773 476
rect 811 448 839 476
rect 877 448 905 476
rect 943 448 971 476
rect 1009 448 1037 476
rect 1075 448 1103 476
rect 1141 448 1169 476
rect 1207 448 1235 476
rect 1273 448 1301 476
rect 1339 448 1367 476
rect 1405 448 1433 476
rect 1471 448 1499 476
rect 1537 448 1565 476
rect 1603 448 1631 476
rect 1669 448 1697 476
rect 1735 448 1763 476
rect 1801 448 1829 476
rect 1867 448 1895 476
rect 1933 448 1961 476
rect 1999 448 2027 476
rect 2065 448 2093 476
rect 2131 448 2159 476
rect 2197 448 2225 476
rect 2263 448 2291 476
rect 2329 448 2357 476
rect 2395 448 2423 476
rect 2461 448 2489 476
rect 2527 448 2555 476
rect 2593 448 2621 476
rect 2659 448 2687 476
rect 2725 448 2753 476
rect 2791 448 2819 476
rect 2857 448 2885 476
rect 2923 448 2951 476
rect 2989 448 3017 476
rect 3055 448 3083 476
rect 3121 448 3149 476
rect 3187 448 3215 476
rect 3253 448 3281 476
rect 3319 448 3347 476
rect 3385 448 3413 476
rect 3451 448 3479 476
rect 3517 448 3545 476
rect 3583 448 3611 476
rect 3649 448 3677 476
rect 3715 448 3743 476
rect 3781 448 3809 476
rect 3847 448 3875 476
rect -3875 382 -3847 410
rect -3809 382 -3781 410
rect -3743 382 -3715 410
rect -3677 382 -3649 410
rect -3611 382 -3583 410
rect -3545 382 -3517 410
rect -3479 382 -3451 410
rect -3413 382 -3385 410
rect -3347 382 -3319 410
rect -3281 382 -3253 410
rect -3215 382 -3187 410
rect -3149 382 -3121 410
rect -3083 382 -3055 410
rect -3017 382 -2989 410
rect -2951 382 -2923 410
rect -2885 382 -2857 410
rect -2819 382 -2791 410
rect -2753 382 -2725 410
rect -2687 382 -2659 410
rect -2621 382 -2593 410
rect -2555 382 -2527 410
rect -2489 382 -2461 410
rect -2423 382 -2395 410
rect -2357 382 -2329 410
rect -2291 382 -2263 410
rect -2225 382 -2197 410
rect -2159 382 -2131 410
rect -2093 382 -2065 410
rect -2027 382 -1999 410
rect -1961 382 -1933 410
rect -1895 382 -1867 410
rect -1829 382 -1801 410
rect -1763 382 -1735 410
rect -1697 382 -1669 410
rect -1631 382 -1603 410
rect -1565 382 -1537 410
rect -1499 382 -1471 410
rect -1433 382 -1405 410
rect -1367 382 -1339 410
rect -1301 382 -1273 410
rect -1235 382 -1207 410
rect -1169 382 -1141 410
rect -1103 382 -1075 410
rect -1037 382 -1009 410
rect -971 382 -943 410
rect -905 382 -877 410
rect -839 382 -811 410
rect -773 382 -745 410
rect -707 382 -679 410
rect -641 382 -613 410
rect -575 382 -547 410
rect -509 382 -481 410
rect -443 382 -415 410
rect -377 382 -349 410
rect -311 382 -283 410
rect -245 382 -217 410
rect -179 382 -151 410
rect -113 382 -85 410
rect -47 382 -19 410
rect 19 382 47 410
rect 85 382 113 410
rect 151 382 179 410
rect 217 382 245 410
rect 283 382 311 410
rect 349 382 377 410
rect 415 382 443 410
rect 481 382 509 410
rect 547 382 575 410
rect 613 382 641 410
rect 679 382 707 410
rect 745 382 773 410
rect 811 382 839 410
rect 877 382 905 410
rect 943 382 971 410
rect 1009 382 1037 410
rect 1075 382 1103 410
rect 1141 382 1169 410
rect 1207 382 1235 410
rect 1273 382 1301 410
rect 1339 382 1367 410
rect 1405 382 1433 410
rect 1471 382 1499 410
rect 1537 382 1565 410
rect 1603 382 1631 410
rect 1669 382 1697 410
rect 1735 382 1763 410
rect 1801 382 1829 410
rect 1867 382 1895 410
rect 1933 382 1961 410
rect 1999 382 2027 410
rect 2065 382 2093 410
rect 2131 382 2159 410
rect 2197 382 2225 410
rect 2263 382 2291 410
rect 2329 382 2357 410
rect 2395 382 2423 410
rect 2461 382 2489 410
rect 2527 382 2555 410
rect 2593 382 2621 410
rect 2659 382 2687 410
rect 2725 382 2753 410
rect 2791 382 2819 410
rect 2857 382 2885 410
rect 2923 382 2951 410
rect 2989 382 3017 410
rect 3055 382 3083 410
rect 3121 382 3149 410
rect 3187 382 3215 410
rect 3253 382 3281 410
rect 3319 382 3347 410
rect 3385 382 3413 410
rect 3451 382 3479 410
rect 3517 382 3545 410
rect 3583 382 3611 410
rect 3649 382 3677 410
rect 3715 382 3743 410
rect 3781 382 3809 410
rect 3847 382 3875 410
rect -3875 316 -3847 344
rect -3809 316 -3781 344
rect -3743 316 -3715 344
rect -3677 316 -3649 344
rect -3611 316 -3583 344
rect -3545 316 -3517 344
rect -3479 316 -3451 344
rect -3413 316 -3385 344
rect -3347 316 -3319 344
rect -3281 316 -3253 344
rect -3215 316 -3187 344
rect -3149 316 -3121 344
rect -3083 316 -3055 344
rect -3017 316 -2989 344
rect -2951 316 -2923 344
rect -2885 316 -2857 344
rect -2819 316 -2791 344
rect -2753 316 -2725 344
rect -2687 316 -2659 344
rect -2621 316 -2593 344
rect -2555 316 -2527 344
rect -2489 316 -2461 344
rect -2423 316 -2395 344
rect -2357 316 -2329 344
rect -2291 316 -2263 344
rect -2225 316 -2197 344
rect -2159 316 -2131 344
rect -2093 316 -2065 344
rect -2027 316 -1999 344
rect -1961 316 -1933 344
rect -1895 316 -1867 344
rect -1829 316 -1801 344
rect -1763 316 -1735 344
rect -1697 316 -1669 344
rect -1631 316 -1603 344
rect -1565 316 -1537 344
rect -1499 316 -1471 344
rect -1433 316 -1405 344
rect -1367 316 -1339 344
rect -1301 316 -1273 344
rect -1235 316 -1207 344
rect -1169 316 -1141 344
rect -1103 316 -1075 344
rect -1037 316 -1009 344
rect -971 316 -943 344
rect -905 316 -877 344
rect -839 316 -811 344
rect -773 316 -745 344
rect -707 316 -679 344
rect -641 316 -613 344
rect -575 316 -547 344
rect -509 316 -481 344
rect -443 316 -415 344
rect -377 316 -349 344
rect -311 316 -283 344
rect -245 316 -217 344
rect -179 316 -151 344
rect -113 316 -85 344
rect -47 316 -19 344
rect 19 316 47 344
rect 85 316 113 344
rect 151 316 179 344
rect 217 316 245 344
rect 283 316 311 344
rect 349 316 377 344
rect 415 316 443 344
rect 481 316 509 344
rect 547 316 575 344
rect 613 316 641 344
rect 679 316 707 344
rect 745 316 773 344
rect 811 316 839 344
rect 877 316 905 344
rect 943 316 971 344
rect 1009 316 1037 344
rect 1075 316 1103 344
rect 1141 316 1169 344
rect 1207 316 1235 344
rect 1273 316 1301 344
rect 1339 316 1367 344
rect 1405 316 1433 344
rect 1471 316 1499 344
rect 1537 316 1565 344
rect 1603 316 1631 344
rect 1669 316 1697 344
rect 1735 316 1763 344
rect 1801 316 1829 344
rect 1867 316 1895 344
rect 1933 316 1961 344
rect 1999 316 2027 344
rect 2065 316 2093 344
rect 2131 316 2159 344
rect 2197 316 2225 344
rect 2263 316 2291 344
rect 2329 316 2357 344
rect 2395 316 2423 344
rect 2461 316 2489 344
rect 2527 316 2555 344
rect 2593 316 2621 344
rect 2659 316 2687 344
rect 2725 316 2753 344
rect 2791 316 2819 344
rect 2857 316 2885 344
rect 2923 316 2951 344
rect 2989 316 3017 344
rect 3055 316 3083 344
rect 3121 316 3149 344
rect 3187 316 3215 344
rect 3253 316 3281 344
rect 3319 316 3347 344
rect 3385 316 3413 344
rect 3451 316 3479 344
rect 3517 316 3545 344
rect 3583 316 3611 344
rect 3649 316 3677 344
rect 3715 316 3743 344
rect 3781 316 3809 344
rect 3847 316 3875 344
rect -3875 250 -3847 278
rect -3809 250 -3781 278
rect -3743 250 -3715 278
rect -3677 250 -3649 278
rect -3611 250 -3583 278
rect -3545 250 -3517 278
rect -3479 250 -3451 278
rect -3413 250 -3385 278
rect -3347 250 -3319 278
rect -3281 250 -3253 278
rect -3215 250 -3187 278
rect -3149 250 -3121 278
rect -3083 250 -3055 278
rect -3017 250 -2989 278
rect -2951 250 -2923 278
rect -2885 250 -2857 278
rect -2819 250 -2791 278
rect -2753 250 -2725 278
rect -2687 250 -2659 278
rect -2621 250 -2593 278
rect -2555 250 -2527 278
rect -2489 250 -2461 278
rect -2423 250 -2395 278
rect -2357 250 -2329 278
rect -2291 250 -2263 278
rect -2225 250 -2197 278
rect -2159 250 -2131 278
rect -2093 250 -2065 278
rect -2027 250 -1999 278
rect -1961 250 -1933 278
rect -1895 250 -1867 278
rect -1829 250 -1801 278
rect -1763 250 -1735 278
rect -1697 250 -1669 278
rect -1631 250 -1603 278
rect -1565 250 -1537 278
rect -1499 250 -1471 278
rect -1433 250 -1405 278
rect -1367 250 -1339 278
rect -1301 250 -1273 278
rect -1235 250 -1207 278
rect -1169 250 -1141 278
rect -1103 250 -1075 278
rect -1037 250 -1009 278
rect -971 250 -943 278
rect -905 250 -877 278
rect -839 250 -811 278
rect -773 250 -745 278
rect -707 250 -679 278
rect -641 250 -613 278
rect -575 250 -547 278
rect -509 250 -481 278
rect -443 250 -415 278
rect -377 250 -349 278
rect -311 250 -283 278
rect -245 250 -217 278
rect -179 250 -151 278
rect -113 250 -85 278
rect -47 250 -19 278
rect 19 250 47 278
rect 85 250 113 278
rect 151 250 179 278
rect 217 250 245 278
rect 283 250 311 278
rect 349 250 377 278
rect 415 250 443 278
rect 481 250 509 278
rect 547 250 575 278
rect 613 250 641 278
rect 679 250 707 278
rect 745 250 773 278
rect 811 250 839 278
rect 877 250 905 278
rect 943 250 971 278
rect 1009 250 1037 278
rect 1075 250 1103 278
rect 1141 250 1169 278
rect 1207 250 1235 278
rect 1273 250 1301 278
rect 1339 250 1367 278
rect 1405 250 1433 278
rect 1471 250 1499 278
rect 1537 250 1565 278
rect 1603 250 1631 278
rect 1669 250 1697 278
rect 1735 250 1763 278
rect 1801 250 1829 278
rect 1867 250 1895 278
rect 1933 250 1961 278
rect 1999 250 2027 278
rect 2065 250 2093 278
rect 2131 250 2159 278
rect 2197 250 2225 278
rect 2263 250 2291 278
rect 2329 250 2357 278
rect 2395 250 2423 278
rect 2461 250 2489 278
rect 2527 250 2555 278
rect 2593 250 2621 278
rect 2659 250 2687 278
rect 2725 250 2753 278
rect 2791 250 2819 278
rect 2857 250 2885 278
rect 2923 250 2951 278
rect 2989 250 3017 278
rect 3055 250 3083 278
rect 3121 250 3149 278
rect 3187 250 3215 278
rect 3253 250 3281 278
rect 3319 250 3347 278
rect 3385 250 3413 278
rect 3451 250 3479 278
rect 3517 250 3545 278
rect 3583 250 3611 278
rect 3649 250 3677 278
rect 3715 250 3743 278
rect 3781 250 3809 278
rect 3847 250 3875 278
rect -3875 184 -3847 212
rect -3809 184 -3781 212
rect -3743 184 -3715 212
rect -3677 184 -3649 212
rect -3611 184 -3583 212
rect -3545 184 -3517 212
rect -3479 184 -3451 212
rect -3413 184 -3385 212
rect -3347 184 -3319 212
rect -3281 184 -3253 212
rect -3215 184 -3187 212
rect -3149 184 -3121 212
rect -3083 184 -3055 212
rect -3017 184 -2989 212
rect -2951 184 -2923 212
rect -2885 184 -2857 212
rect -2819 184 -2791 212
rect -2753 184 -2725 212
rect -2687 184 -2659 212
rect -2621 184 -2593 212
rect -2555 184 -2527 212
rect -2489 184 -2461 212
rect -2423 184 -2395 212
rect -2357 184 -2329 212
rect -2291 184 -2263 212
rect -2225 184 -2197 212
rect -2159 184 -2131 212
rect -2093 184 -2065 212
rect -2027 184 -1999 212
rect -1961 184 -1933 212
rect -1895 184 -1867 212
rect -1829 184 -1801 212
rect -1763 184 -1735 212
rect -1697 184 -1669 212
rect -1631 184 -1603 212
rect -1565 184 -1537 212
rect -1499 184 -1471 212
rect -1433 184 -1405 212
rect -1367 184 -1339 212
rect -1301 184 -1273 212
rect -1235 184 -1207 212
rect -1169 184 -1141 212
rect -1103 184 -1075 212
rect -1037 184 -1009 212
rect -971 184 -943 212
rect -905 184 -877 212
rect -839 184 -811 212
rect -773 184 -745 212
rect -707 184 -679 212
rect -641 184 -613 212
rect -575 184 -547 212
rect -509 184 -481 212
rect -443 184 -415 212
rect -377 184 -349 212
rect -311 184 -283 212
rect -245 184 -217 212
rect -179 184 -151 212
rect -113 184 -85 212
rect -47 184 -19 212
rect 19 184 47 212
rect 85 184 113 212
rect 151 184 179 212
rect 217 184 245 212
rect 283 184 311 212
rect 349 184 377 212
rect 415 184 443 212
rect 481 184 509 212
rect 547 184 575 212
rect 613 184 641 212
rect 679 184 707 212
rect 745 184 773 212
rect 811 184 839 212
rect 877 184 905 212
rect 943 184 971 212
rect 1009 184 1037 212
rect 1075 184 1103 212
rect 1141 184 1169 212
rect 1207 184 1235 212
rect 1273 184 1301 212
rect 1339 184 1367 212
rect 1405 184 1433 212
rect 1471 184 1499 212
rect 1537 184 1565 212
rect 1603 184 1631 212
rect 1669 184 1697 212
rect 1735 184 1763 212
rect 1801 184 1829 212
rect 1867 184 1895 212
rect 1933 184 1961 212
rect 1999 184 2027 212
rect 2065 184 2093 212
rect 2131 184 2159 212
rect 2197 184 2225 212
rect 2263 184 2291 212
rect 2329 184 2357 212
rect 2395 184 2423 212
rect 2461 184 2489 212
rect 2527 184 2555 212
rect 2593 184 2621 212
rect 2659 184 2687 212
rect 2725 184 2753 212
rect 2791 184 2819 212
rect 2857 184 2885 212
rect 2923 184 2951 212
rect 2989 184 3017 212
rect 3055 184 3083 212
rect 3121 184 3149 212
rect 3187 184 3215 212
rect 3253 184 3281 212
rect 3319 184 3347 212
rect 3385 184 3413 212
rect 3451 184 3479 212
rect 3517 184 3545 212
rect 3583 184 3611 212
rect 3649 184 3677 212
rect 3715 184 3743 212
rect 3781 184 3809 212
rect 3847 184 3875 212
rect -3875 118 -3847 146
rect -3809 118 -3781 146
rect -3743 118 -3715 146
rect -3677 118 -3649 146
rect -3611 118 -3583 146
rect -3545 118 -3517 146
rect -3479 118 -3451 146
rect -3413 118 -3385 146
rect -3347 118 -3319 146
rect -3281 118 -3253 146
rect -3215 118 -3187 146
rect -3149 118 -3121 146
rect -3083 118 -3055 146
rect -3017 118 -2989 146
rect -2951 118 -2923 146
rect -2885 118 -2857 146
rect -2819 118 -2791 146
rect -2753 118 -2725 146
rect -2687 118 -2659 146
rect -2621 118 -2593 146
rect -2555 118 -2527 146
rect -2489 118 -2461 146
rect -2423 118 -2395 146
rect -2357 118 -2329 146
rect -2291 118 -2263 146
rect -2225 118 -2197 146
rect -2159 118 -2131 146
rect -2093 118 -2065 146
rect -2027 118 -1999 146
rect -1961 118 -1933 146
rect -1895 118 -1867 146
rect -1829 118 -1801 146
rect -1763 118 -1735 146
rect -1697 118 -1669 146
rect -1631 118 -1603 146
rect -1565 118 -1537 146
rect -1499 118 -1471 146
rect -1433 118 -1405 146
rect -1367 118 -1339 146
rect -1301 118 -1273 146
rect -1235 118 -1207 146
rect -1169 118 -1141 146
rect -1103 118 -1075 146
rect -1037 118 -1009 146
rect -971 118 -943 146
rect -905 118 -877 146
rect -839 118 -811 146
rect -773 118 -745 146
rect -707 118 -679 146
rect -641 118 -613 146
rect -575 118 -547 146
rect -509 118 -481 146
rect -443 118 -415 146
rect -377 118 -349 146
rect -311 118 -283 146
rect -245 118 -217 146
rect -179 118 -151 146
rect -113 118 -85 146
rect -47 118 -19 146
rect 19 118 47 146
rect 85 118 113 146
rect 151 118 179 146
rect 217 118 245 146
rect 283 118 311 146
rect 349 118 377 146
rect 415 118 443 146
rect 481 118 509 146
rect 547 118 575 146
rect 613 118 641 146
rect 679 118 707 146
rect 745 118 773 146
rect 811 118 839 146
rect 877 118 905 146
rect 943 118 971 146
rect 1009 118 1037 146
rect 1075 118 1103 146
rect 1141 118 1169 146
rect 1207 118 1235 146
rect 1273 118 1301 146
rect 1339 118 1367 146
rect 1405 118 1433 146
rect 1471 118 1499 146
rect 1537 118 1565 146
rect 1603 118 1631 146
rect 1669 118 1697 146
rect 1735 118 1763 146
rect 1801 118 1829 146
rect 1867 118 1895 146
rect 1933 118 1961 146
rect 1999 118 2027 146
rect 2065 118 2093 146
rect 2131 118 2159 146
rect 2197 118 2225 146
rect 2263 118 2291 146
rect 2329 118 2357 146
rect 2395 118 2423 146
rect 2461 118 2489 146
rect 2527 118 2555 146
rect 2593 118 2621 146
rect 2659 118 2687 146
rect 2725 118 2753 146
rect 2791 118 2819 146
rect 2857 118 2885 146
rect 2923 118 2951 146
rect 2989 118 3017 146
rect 3055 118 3083 146
rect 3121 118 3149 146
rect 3187 118 3215 146
rect 3253 118 3281 146
rect 3319 118 3347 146
rect 3385 118 3413 146
rect 3451 118 3479 146
rect 3517 118 3545 146
rect 3583 118 3611 146
rect 3649 118 3677 146
rect 3715 118 3743 146
rect 3781 118 3809 146
rect 3847 118 3875 146
rect -3875 52 -3847 80
rect -3809 52 -3781 80
rect -3743 52 -3715 80
rect -3677 52 -3649 80
rect -3611 52 -3583 80
rect -3545 52 -3517 80
rect -3479 52 -3451 80
rect -3413 52 -3385 80
rect -3347 52 -3319 80
rect -3281 52 -3253 80
rect -3215 52 -3187 80
rect -3149 52 -3121 80
rect -3083 52 -3055 80
rect -3017 52 -2989 80
rect -2951 52 -2923 80
rect -2885 52 -2857 80
rect -2819 52 -2791 80
rect -2753 52 -2725 80
rect -2687 52 -2659 80
rect -2621 52 -2593 80
rect -2555 52 -2527 80
rect -2489 52 -2461 80
rect -2423 52 -2395 80
rect -2357 52 -2329 80
rect -2291 52 -2263 80
rect -2225 52 -2197 80
rect -2159 52 -2131 80
rect -2093 52 -2065 80
rect -2027 52 -1999 80
rect -1961 52 -1933 80
rect -1895 52 -1867 80
rect -1829 52 -1801 80
rect -1763 52 -1735 80
rect -1697 52 -1669 80
rect -1631 52 -1603 80
rect -1565 52 -1537 80
rect -1499 52 -1471 80
rect -1433 52 -1405 80
rect -1367 52 -1339 80
rect -1301 52 -1273 80
rect -1235 52 -1207 80
rect -1169 52 -1141 80
rect -1103 52 -1075 80
rect -1037 52 -1009 80
rect -971 52 -943 80
rect -905 52 -877 80
rect -839 52 -811 80
rect -773 52 -745 80
rect -707 52 -679 80
rect -641 52 -613 80
rect -575 52 -547 80
rect -509 52 -481 80
rect -443 52 -415 80
rect -377 52 -349 80
rect -311 52 -283 80
rect -245 52 -217 80
rect -179 52 -151 80
rect -113 52 -85 80
rect -47 52 -19 80
rect 19 52 47 80
rect 85 52 113 80
rect 151 52 179 80
rect 217 52 245 80
rect 283 52 311 80
rect 349 52 377 80
rect 415 52 443 80
rect 481 52 509 80
rect 547 52 575 80
rect 613 52 641 80
rect 679 52 707 80
rect 745 52 773 80
rect 811 52 839 80
rect 877 52 905 80
rect 943 52 971 80
rect 1009 52 1037 80
rect 1075 52 1103 80
rect 1141 52 1169 80
rect 1207 52 1235 80
rect 1273 52 1301 80
rect 1339 52 1367 80
rect 1405 52 1433 80
rect 1471 52 1499 80
rect 1537 52 1565 80
rect 1603 52 1631 80
rect 1669 52 1697 80
rect 1735 52 1763 80
rect 1801 52 1829 80
rect 1867 52 1895 80
rect 1933 52 1961 80
rect 1999 52 2027 80
rect 2065 52 2093 80
rect 2131 52 2159 80
rect 2197 52 2225 80
rect 2263 52 2291 80
rect 2329 52 2357 80
rect 2395 52 2423 80
rect 2461 52 2489 80
rect 2527 52 2555 80
rect 2593 52 2621 80
rect 2659 52 2687 80
rect 2725 52 2753 80
rect 2791 52 2819 80
rect 2857 52 2885 80
rect 2923 52 2951 80
rect 2989 52 3017 80
rect 3055 52 3083 80
rect 3121 52 3149 80
rect 3187 52 3215 80
rect 3253 52 3281 80
rect 3319 52 3347 80
rect 3385 52 3413 80
rect 3451 52 3479 80
rect 3517 52 3545 80
rect 3583 52 3611 80
rect 3649 52 3677 80
rect 3715 52 3743 80
rect 3781 52 3809 80
rect 3847 52 3875 80
rect -3875 -14 -3847 14
rect -3809 -14 -3781 14
rect -3743 -14 -3715 14
rect -3677 -14 -3649 14
rect -3611 -14 -3583 14
rect -3545 -14 -3517 14
rect -3479 -14 -3451 14
rect -3413 -14 -3385 14
rect -3347 -14 -3319 14
rect -3281 -14 -3253 14
rect -3215 -14 -3187 14
rect -3149 -14 -3121 14
rect -3083 -14 -3055 14
rect -3017 -14 -2989 14
rect -2951 -14 -2923 14
rect -2885 -14 -2857 14
rect -2819 -14 -2791 14
rect -2753 -14 -2725 14
rect -2687 -14 -2659 14
rect -2621 -14 -2593 14
rect -2555 -14 -2527 14
rect -2489 -14 -2461 14
rect -2423 -14 -2395 14
rect -2357 -14 -2329 14
rect -2291 -14 -2263 14
rect -2225 -14 -2197 14
rect -2159 -14 -2131 14
rect -2093 -14 -2065 14
rect -2027 -14 -1999 14
rect -1961 -14 -1933 14
rect -1895 -14 -1867 14
rect -1829 -14 -1801 14
rect -1763 -14 -1735 14
rect -1697 -14 -1669 14
rect -1631 -14 -1603 14
rect -1565 -14 -1537 14
rect -1499 -14 -1471 14
rect -1433 -14 -1405 14
rect -1367 -14 -1339 14
rect -1301 -14 -1273 14
rect -1235 -14 -1207 14
rect -1169 -14 -1141 14
rect -1103 -14 -1075 14
rect -1037 -14 -1009 14
rect -971 -14 -943 14
rect -905 -14 -877 14
rect -839 -14 -811 14
rect -773 -14 -745 14
rect -707 -14 -679 14
rect -641 -14 -613 14
rect -575 -14 -547 14
rect -509 -14 -481 14
rect -443 -14 -415 14
rect -377 -14 -349 14
rect -311 -14 -283 14
rect -245 -14 -217 14
rect -179 -14 -151 14
rect -113 -14 -85 14
rect -47 -14 -19 14
rect 19 -14 47 14
rect 85 -14 113 14
rect 151 -14 179 14
rect 217 -14 245 14
rect 283 -14 311 14
rect 349 -14 377 14
rect 415 -14 443 14
rect 481 -14 509 14
rect 547 -14 575 14
rect 613 -14 641 14
rect 679 -14 707 14
rect 745 -14 773 14
rect 811 -14 839 14
rect 877 -14 905 14
rect 943 -14 971 14
rect 1009 -14 1037 14
rect 1075 -14 1103 14
rect 1141 -14 1169 14
rect 1207 -14 1235 14
rect 1273 -14 1301 14
rect 1339 -14 1367 14
rect 1405 -14 1433 14
rect 1471 -14 1499 14
rect 1537 -14 1565 14
rect 1603 -14 1631 14
rect 1669 -14 1697 14
rect 1735 -14 1763 14
rect 1801 -14 1829 14
rect 1867 -14 1895 14
rect 1933 -14 1961 14
rect 1999 -14 2027 14
rect 2065 -14 2093 14
rect 2131 -14 2159 14
rect 2197 -14 2225 14
rect 2263 -14 2291 14
rect 2329 -14 2357 14
rect 2395 -14 2423 14
rect 2461 -14 2489 14
rect 2527 -14 2555 14
rect 2593 -14 2621 14
rect 2659 -14 2687 14
rect 2725 -14 2753 14
rect 2791 -14 2819 14
rect 2857 -14 2885 14
rect 2923 -14 2951 14
rect 2989 -14 3017 14
rect 3055 -14 3083 14
rect 3121 -14 3149 14
rect 3187 -14 3215 14
rect 3253 -14 3281 14
rect 3319 -14 3347 14
rect 3385 -14 3413 14
rect 3451 -14 3479 14
rect 3517 -14 3545 14
rect 3583 -14 3611 14
rect 3649 -14 3677 14
rect 3715 -14 3743 14
rect 3781 -14 3809 14
rect 3847 -14 3875 14
rect -3875 -80 -3847 -52
rect -3809 -80 -3781 -52
rect -3743 -80 -3715 -52
rect -3677 -80 -3649 -52
rect -3611 -80 -3583 -52
rect -3545 -80 -3517 -52
rect -3479 -80 -3451 -52
rect -3413 -80 -3385 -52
rect -3347 -80 -3319 -52
rect -3281 -80 -3253 -52
rect -3215 -80 -3187 -52
rect -3149 -80 -3121 -52
rect -3083 -80 -3055 -52
rect -3017 -80 -2989 -52
rect -2951 -80 -2923 -52
rect -2885 -80 -2857 -52
rect -2819 -80 -2791 -52
rect -2753 -80 -2725 -52
rect -2687 -80 -2659 -52
rect -2621 -80 -2593 -52
rect -2555 -80 -2527 -52
rect -2489 -80 -2461 -52
rect -2423 -80 -2395 -52
rect -2357 -80 -2329 -52
rect -2291 -80 -2263 -52
rect -2225 -80 -2197 -52
rect -2159 -80 -2131 -52
rect -2093 -80 -2065 -52
rect -2027 -80 -1999 -52
rect -1961 -80 -1933 -52
rect -1895 -80 -1867 -52
rect -1829 -80 -1801 -52
rect -1763 -80 -1735 -52
rect -1697 -80 -1669 -52
rect -1631 -80 -1603 -52
rect -1565 -80 -1537 -52
rect -1499 -80 -1471 -52
rect -1433 -80 -1405 -52
rect -1367 -80 -1339 -52
rect -1301 -80 -1273 -52
rect -1235 -80 -1207 -52
rect -1169 -80 -1141 -52
rect -1103 -80 -1075 -52
rect -1037 -80 -1009 -52
rect -971 -80 -943 -52
rect -905 -80 -877 -52
rect -839 -80 -811 -52
rect -773 -80 -745 -52
rect -707 -80 -679 -52
rect -641 -80 -613 -52
rect -575 -80 -547 -52
rect -509 -80 -481 -52
rect -443 -80 -415 -52
rect -377 -80 -349 -52
rect -311 -80 -283 -52
rect -245 -80 -217 -52
rect -179 -80 -151 -52
rect -113 -80 -85 -52
rect -47 -80 -19 -52
rect 19 -80 47 -52
rect 85 -80 113 -52
rect 151 -80 179 -52
rect 217 -80 245 -52
rect 283 -80 311 -52
rect 349 -80 377 -52
rect 415 -80 443 -52
rect 481 -80 509 -52
rect 547 -80 575 -52
rect 613 -80 641 -52
rect 679 -80 707 -52
rect 745 -80 773 -52
rect 811 -80 839 -52
rect 877 -80 905 -52
rect 943 -80 971 -52
rect 1009 -80 1037 -52
rect 1075 -80 1103 -52
rect 1141 -80 1169 -52
rect 1207 -80 1235 -52
rect 1273 -80 1301 -52
rect 1339 -80 1367 -52
rect 1405 -80 1433 -52
rect 1471 -80 1499 -52
rect 1537 -80 1565 -52
rect 1603 -80 1631 -52
rect 1669 -80 1697 -52
rect 1735 -80 1763 -52
rect 1801 -80 1829 -52
rect 1867 -80 1895 -52
rect 1933 -80 1961 -52
rect 1999 -80 2027 -52
rect 2065 -80 2093 -52
rect 2131 -80 2159 -52
rect 2197 -80 2225 -52
rect 2263 -80 2291 -52
rect 2329 -80 2357 -52
rect 2395 -80 2423 -52
rect 2461 -80 2489 -52
rect 2527 -80 2555 -52
rect 2593 -80 2621 -52
rect 2659 -80 2687 -52
rect 2725 -80 2753 -52
rect 2791 -80 2819 -52
rect 2857 -80 2885 -52
rect 2923 -80 2951 -52
rect 2989 -80 3017 -52
rect 3055 -80 3083 -52
rect 3121 -80 3149 -52
rect 3187 -80 3215 -52
rect 3253 -80 3281 -52
rect 3319 -80 3347 -52
rect 3385 -80 3413 -52
rect 3451 -80 3479 -52
rect 3517 -80 3545 -52
rect 3583 -80 3611 -52
rect 3649 -80 3677 -52
rect 3715 -80 3743 -52
rect 3781 -80 3809 -52
rect 3847 -80 3875 -52
rect -3875 -146 -3847 -118
rect -3809 -146 -3781 -118
rect -3743 -146 -3715 -118
rect -3677 -146 -3649 -118
rect -3611 -146 -3583 -118
rect -3545 -146 -3517 -118
rect -3479 -146 -3451 -118
rect -3413 -146 -3385 -118
rect -3347 -146 -3319 -118
rect -3281 -146 -3253 -118
rect -3215 -146 -3187 -118
rect -3149 -146 -3121 -118
rect -3083 -146 -3055 -118
rect -3017 -146 -2989 -118
rect -2951 -146 -2923 -118
rect -2885 -146 -2857 -118
rect -2819 -146 -2791 -118
rect -2753 -146 -2725 -118
rect -2687 -146 -2659 -118
rect -2621 -146 -2593 -118
rect -2555 -146 -2527 -118
rect -2489 -146 -2461 -118
rect -2423 -146 -2395 -118
rect -2357 -146 -2329 -118
rect -2291 -146 -2263 -118
rect -2225 -146 -2197 -118
rect -2159 -146 -2131 -118
rect -2093 -146 -2065 -118
rect -2027 -146 -1999 -118
rect -1961 -146 -1933 -118
rect -1895 -146 -1867 -118
rect -1829 -146 -1801 -118
rect -1763 -146 -1735 -118
rect -1697 -146 -1669 -118
rect -1631 -146 -1603 -118
rect -1565 -146 -1537 -118
rect -1499 -146 -1471 -118
rect -1433 -146 -1405 -118
rect -1367 -146 -1339 -118
rect -1301 -146 -1273 -118
rect -1235 -146 -1207 -118
rect -1169 -146 -1141 -118
rect -1103 -146 -1075 -118
rect -1037 -146 -1009 -118
rect -971 -146 -943 -118
rect -905 -146 -877 -118
rect -839 -146 -811 -118
rect -773 -146 -745 -118
rect -707 -146 -679 -118
rect -641 -146 -613 -118
rect -575 -146 -547 -118
rect -509 -146 -481 -118
rect -443 -146 -415 -118
rect -377 -146 -349 -118
rect -311 -146 -283 -118
rect -245 -146 -217 -118
rect -179 -146 -151 -118
rect -113 -146 -85 -118
rect -47 -146 -19 -118
rect 19 -146 47 -118
rect 85 -146 113 -118
rect 151 -146 179 -118
rect 217 -146 245 -118
rect 283 -146 311 -118
rect 349 -146 377 -118
rect 415 -146 443 -118
rect 481 -146 509 -118
rect 547 -146 575 -118
rect 613 -146 641 -118
rect 679 -146 707 -118
rect 745 -146 773 -118
rect 811 -146 839 -118
rect 877 -146 905 -118
rect 943 -146 971 -118
rect 1009 -146 1037 -118
rect 1075 -146 1103 -118
rect 1141 -146 1169 -118
rect 1207 -146 1235 -118
rect 1273 -146 1301 -118
rect 1339 -146 1367 -118
rect 1405 -146 1433 -118
rect 1471 -146 1499 -118
rect 1537 -146 1565 -118
rect 1603 -146 1631 -118
rect 1669 -146 1697 -118
rect 1735 -146 1763 -118
rect 1801 -146 1829 -118
rect 1867 -146 1895 -118
rect 1933 -146 1961 -118
rect 1999 -146 2027 -118
rect 2065 -146 2093 -118
rect 2131 -146 2159 -118
rect 2197 -146 2225 -118
rect 2263 -146 2291 -118
rect 2329 -146 2357 -118
rect 2395 -146 2423 -118
rect 2461 -146 2489 -118
rect 2527 -146 2555 -118
rect 2593 -146 2621 -118
rect 2659 -146 2687 -118
rect 2725 -146 2753 -118
rect 2791 -146 2819 -118
rect 2857 -146 2885 -118
rect 2923 -146 2951 -118
rect 2989 -146 3017 -118
rect 3055 -146 3083 -118
rect 3121 -146 3149 -118
rect 3187 -146 3215 -118
rect 3253 -146 3281 -118
rect 3319 -146 3347 -118
rect 3385 -146 3413 -118
rect 3451 -146 3479 -118
rect 3517 -146 3545 -118
rect 3583 -146 3611 -118
rect 3649 -146 3677 -118
rect 3715 -146 3743 -118
rect 3781 -146 3809 -118
rect 3847 -146 3875 -118
rect -3875 -212 -3847 -184
rect -3809 -212 -3781 -184
rect -3743 -212 -3715 -184
rect -3677 -212 -3649 -184
rect -3611 -212 -3583 -184
rect -3545 -212 -3517 -184
rect -3479 -212 -3451 -184
rect -3413 -212 -3385 -184
rect -3347 -212 -3319 -184
rect -3281 -212 -3253 -184
rect -3215 -212 -3187 -184
rect -3149 -212 -3121 -184
rect -3083 -212 -3055 -184
rect -3017 -212 -2989 -184
rect -2951 -212 -2923 -184
rect -2885 -212 -2857 -184
rect -2819 -212 -2791 -184
rect -2753 -212 -2725 -184
rect -2687 -212 -2659 -184
rect -2621 -212 -2593 -184
rect -2555 -212 -2527 -184
rect -2489 -212 -2461 -184
rect -2423 -212 -2395 -184
rect -2357 -212 -2329 -184
rect -2291 -212 -2263 -184
rect -2225 -212 -2197 -184
rect -2159 -212 -2131 -184
rect -2093 -212 -2065 -184
rect -2027 -212 -1999 -184
rect -1961 -212 -1933 -184
rect -1895 -212 -1867 -184
rect -1829 -212 -1801 -184
rect -1763 -212 -1735 -184
rect -1697 -212 -1669 -184
rect -1631 -212 -1603 -184
rect -1565 -212 -1537 -184
rect -1499 -212 -1471 -184
rect -1433 -212 -1405 -184
rect -1367 -212 -1339 -184
rect -1301 -212 -1273 -184
rect -1235 -212 -1207 -184
rect -1169 -212 -1141 -184
rect -1103 -212 -1075 -184
rect -1037 -212 -1009 -184
rect -971 -212 -943 -184
rect -905 -212 -877 -184
rect -839 -212 -811 -184
rect -773 -212 -745 -184
rect -707 -212 -679 -184
rect -641 -212 -613 -184
rect -575 -212 -547 -184
rect -509 -212 -481 -184
rect -443 -212 -415 -184
rect -377 -212 -349 -184
rect -311 -212 -283 -184
rect -245 -212 -217 -184
rect -179 -212 -151 -184
rect -113 -212 -85 -184
rect -47 -212 -19 -184
rect 19 -212 47 -184
rect 85 -212 113 -184
rect 151 -212 179 -184
rect 217 -212 245 -184
rect 283 -212 311 -184
rect 349 -212 377 -184
rect 415 -212 443 -184
rect 481 -212 509 -184
rect 547 -212 575 -184
rect 613 -212 641 -184
rect 679 -212 707 -184
rect 745 -212 773 -184
rect 811 -212 839 -184
rect 877 -212 905 -184
rect 943 -212 971 -184
rect 1009 -212 1037 -184
rect 1075 -212 1103 -184
rect 1141 -212 1169 -184
rect 1207 -212 1235 -184
rect 1273 -212 1301 -184
rect 1339 -212 1367 -184
rect 1405 -212 1433 -184
rect 1471 -212 1499 -184
rect 1537 -212 1565 -184
rect 1603 -212 1631 -184
rect 1669 -212 1697 -184
rect 1735 -212 1763 -184
rect 1801 -212 1829 -184
rect 1867 -212 1895 -184
rect 1933 -212 1961 -184
rect 1999 -212 2027 -184
rect 2065 -212 2093 -184
rect 2131 -212 2159 -184
rect 2197 -212 2225 -184
rect 2263 -212 2291 -184
rect 2329 -212 2357 -184
rect 2395 -212 2423 -184
rect 2461 -212 2489 -184
rect 2527 -212 2555 -184
rect 2593 -212 2621 -184
rect 2659 -212 2687 -184
rect 2725 -212 2753 -184
rect 2791 -212 2819 -184
rect 2857 -212 2885 -184
rect 2923 -212 2951 -184
rect 2989 -212 3017 -184
rect 3055 -212 3083 -184
rect 3121 -212 3149 -184
rect 3187 -212 3215 -184
rect 3253 -212 3281 -184
rect 3319 -212 3347 -184
rect 3385 -212 3413 -184
rect 3451 -212 3479 -184
rect 3517 -212 3545 -184
rect 3583 -212 3611 -184
rect 3649 -212 3677 -184
rect 3715 -212 3743 -184
rect 3781 -212 3809 -184
rect 3847 -212 3875 -184
rect -3875 -278 -3847 -250
rect -3809 -278 -3781 -250
rect -3743 -278 -3715 -250
rect -3677 -278 -3649 -250
rect -3611 -278 -3583 -250
rect -3545 -278 -3517 -250
rect -3479 -278 -3451 -250
rect -3413 -278 -3385 -250
rect -3347 -278 -3319 -250
rect -3281 -278 -3253 -250
rect -3215 -278 -3187 -250
rect -3149 -278 -3121 -250
rect -3083 -278 -3055 -250
rect -3017 -278 -2989 -250
rect -2951 -278 -2923 -250
rect -2885 -278 -2857 -250
rect -2819 -278 -2791 -250
rect -2753 -278 -2725 -250
rect -2687 -278 -2659 -250
rect -2621 -278 -2593 -250
rect -2555 -278 -2527 -250
rect -2489 -278 -2461 -250
rect -2423 -278 -2395 -250
rect -2357 -278 -2329 -250
rect -2291 -278 -2263 -250
rect -2225 -278 -2197 -250
rect -2159 -278 -2131 -250
rect -2093 -278 -2065 -250
rect -2027 -278 -1999 -250
rect -1961 -278 -1933 -250
rect -1895 -278 -1867 -250
rect -1829 -278 -1801 -250
rect -1763 -278 -1735 -250
rect -1697 -278 -1669 -250
rect -1631 -278 -1603 -250
rect -1565 -278 -1537 -250
rect -1499 -278 -1471 -250
rect -1433 -278 -1405 -250
rect -1367 -278 -1339 -250
rect -1301 -278 -1273 -250
rect -1235 -278 -1207 -250
rect -1169 -278 -1141 -250
rect -1103 -278 -1075 -250
rect -1037 -278 -1009 -250
rect -971 -278 -943 -250
rect -905 -278 -877 -250
rect -839 -278 -811 -250
rect -773 -278 -745 -250
rect -707 -278 -679 -250
rect -641 -278 -613 -250
rect -575 -278 -547 -250
rect -509 -278 -481 -250
rect -443 -278 -415 -250
rect -377 -278 -349 -250
rect -311 -278 -283 -250
rect -245 -278 -217 -250
rect -179 -278 -151 -250
rect -113 -278 -85 -250
rect -47 -278 -19 -250
rect 19 -278 47 -250
rect 85 -278 113 -250
rect 151 -278 179 -250
rect 217 -278 245 -250
rect 283 -278 311 -250
rect 349 -278 377 -250
rect 415 -278 443 -250
rect 481 -278 509 -250
rect 547 -278 575 -250
rect 613 -278 641 -250
rect 679 -278 707 -250
rect 745 -278 773 -250
rect 811 -278 839 -250
rect 877 -278 905 -250
rect 943 -278 971 -250
rect 1009 -278 1037 -250
rect 1075 -278 1103 -250
rect 1141 -278 1169 -250
rect 1207 -278 1235 -250
rect 1273 -278 1301 -250
rect 1339 -278 1367 -250
rect 1405 -278 1433 -250
rect 1471 -278 1499 -250
rect 1537 -278 1565 -250
rect 1603 -278 1631 -250
rect 1669 -278 1697 -250
rect 1735 -278 1763 -250
rect 1801 -278 1829 -250
rect 1867 -278 1895 -250
rect 1933 -278 1961 -250
rect 1999 -278 2027 -250
rect 2065 -278 2093 -250
rect 2131 -278 2159 -250
rect 2197 -278 2225 -250
rect 2263 -278 2291 -250
rect 2329 -278 2357 -250
rect 2395 -278 2423 -250
rect 2461 -278 2489 -250
rect 2527 -278 2555 -250
rect 2593 -278 2621 -250
rect 2659 -278 2687 -250
rect 2725 -278 2753 -250
rect 2791 -278 2819 -250
rect 2857 -278 2885 -250
rect 2923 -278 2951 -250
rect 2989 -278 3017 -250
rect 3055 -278 3083 -250
rect 3121 -278 3149 -250
rect 3187 -278 3215 -250
rect 3253 -278 3281 -250
rect 3319 -278 3347 -250
rect 3385 -278 3413 -250
rect 3451 -278 3479 -250
rect 3517 -278 3545 -250
rect 3583 -278 3611 -250
rect 3649 -278 3677 -250
rect 3715 -278 3743 -250
rect 3781 -278 3809 -250
rect 3847 -278 3875 -250
rect -3875 -344 -3847 -316
rect -3809 -344 -3781 -316
rect -3743 -344 -3715 -316
rect -3677 -344 -3649 -316
rect -3611 -344 -3583 -316
rect -3545 -344 -3517 -316
rect -3479 -344 -3451 -316
rect -3413 -344 -3385 -316
rect -3347 -344 -3319 -316
rect -3281 -344 -3253 -316
rect -3215 -344 -3187 -316
rect -3149 -344 -3121 -316
rect -3083 -344 -3055 -316
rect -3017 -344 -2989 -316
rect -2951 -344 -2923 -316
rect -2885 -344 -2857 -316
rect -2819 -344 -2791 -316
rect -2753 -344 -2725 -316
rect -2687 -344 -2659 -316
rect -2621 -344 -2593 -316
rect -2555 -344 -2527 -316
rect -2489 -344 -2461 -316
rect -2423 -344 -2395 -316
rect -2357 -344 -2329 -316
rect -2291 -344 -2263 -316
rect -2225 -344 -2197 -316
rect -2159 -344 -2131 -316
rect -2093 -344 -2065 -316
rect -2027 -344 -1999 -316
rect -1961 -344 -1933 -316
rect -1895 -344 -1867 -316
rect -1829 -344 -1801 -316
rect -1763 -344 -1735 -316
rect -1697 -344 -1669 -316
rect -1631 -344 -1603 -316
rect -1565 -344 -1537 -316
rect -1499 -344 -1471 -316
rect -1433 -344 -1405 -316
rect -1367 -344 -1339 -316
rect -1301 -344 -1273 -316
rect -1235 -344 -1207 -316
rect -1169 -344 -1141 -316
rect -1103 -344 -1075 -316
rect -1037 -344 -1009 -316
rect -971 -344 -943 -316
rect -905 -344 -877 -316
rect -839 -344 -811 -316
rect -773 -344 -745 -316
rect -707 -344 -679 -316
rect -641 -344 -613 -316
rect -575 -344 -547 -316
rect -509 -344 -481 -316
rect -443 -344 -415 -316
rect -377 -344 -349 -316
rect -311 -344 -283 -316
rect -245 -344 -217 -316
rect -179 -344 -151 -316
rect -113 -344 -85 -316
rect -47 -344 -19 -316
rect 19 -344 47 -316
rect 85 -344 113 -316
rect 151 -344 179 -316
rect 217 -344 245 -316
rect 283 -344 311 -316
rect 349 -344 377 -316
rect 415 -344 443 -316
rect 481 -344 509 -316
rect 547 -344 575 -316
rect 613 -344 641 -316
rect 679 -344 707 -316
rect 745 -344 773 -316
rect 811 -344 839 -316
rect 877 -344 905 -316
rect 943 -344 971 -316
rect 1009 -344 1037 -316
rect 1075 -344 1103 -316
rect 1141 -344 1169 -316
rect 1207 -344 1235 -316
rect 1273 -344 1301 -316
rect 1339 -344 1367 -316
rect 1405 -344 1433 -316
rect 1471 -344 1499 -316
rect 1537 -344 1565 -316
rect 1603 -344 1631 -316
rect 1669 -344 1697 -316
rect 1735 -344 1763 -316
rect 1801 -344 1829 -316
rect 1867 -344 1895 -316
rect 1933 -344 1961 -316
rect 1999 -344 2027 -316
rect 2065 -344 2093 -316
rect 2131 -344 2159 -316
rect 2197 -344 2225 -316
rect 2263 -344 2291 -316
rect 2329 -344 2357 -316
rect 2395 -344 2423 -316
rect 2461 -344 2489 -316
rect 2527 -344 2555 -316
rect 2593 -344 2621 -316
rect 2659 -344 2687 -316
rect 2725 -344 2753 -316
rect 2791 -344 2819 -316
rect 2857 -344 2885 -316
rect 2923 -344 2951 -316
rect 2989 -344 3017 -316
rect 3055 -344 3083 -316
rect 3121 -344 3149 -316
rect 3187 -344 3215 -316
rect 3253 -344 3281 -316
rect 3319 -344 3347 -316
rect 3385 -344 3413 -316
rect 3451 -344 3479 -316
rect 3517 -344 3545 -316
rect 3583 -344 3611 -316
rect 3649 -344 3677 -316
rect 3715 -344 3743 -316
rect 3781 -344 3809 -316
rect 3847 -344 3875 -316
rect -3875 -410 -3847 -382
rect -3809 -410 -3781 -382
rect -3743 -410 -3715 -382
rect -3677 -410 -3649 -382
rect -3611 -410 -3583 -382
rect -3545 -410 -3517 -382
rect -3479 -410 -3451 -382
rect -3413 -410 -3385 -382
rect -3347 -410 -3319 -382
rect -3281 -410 -3253 -382
rect -3215 -410 -3187 -382
rect -3149 -410 -3121 -382
rect -3083 -410 -3055 -382
rect -3017 -410 -2989 -382
rect -2951 -410 -2923 -382
rect -2885 -410 -2857 -382
rect -2819 -410 -2791 -382
rect -2753 -410 -2725 -382
rect -2687 -410 -2659 -382
rect -2621 -410 -2593 -382
rect -2555 -410 -2527 -382
rect -2489 -410 -2461 -382
rect -2423 -410 -2395 -382
rect -2357 -410 -2329 -382
rect -2291 -410 -2263 -382
rect -2225 -410 -2197 -382
rect -2159 -410 -2131 -382
rect -2093 -410 -2065 -382
rect -2027 -410 -1999 -382
rect -1961 -410 -1933 -382
rect -1895 -410 -1867 -382
rect -1829 -410 -1801 -382
rect -1763 -410 -1735 -382
rect -1697 -410 -1669 -382
rect -1631 -410 -1603 -382
rect -1565 -410 -1537 -382
rect -1499 -410 -1471 -382
rect -1433 -410 -1405 -382
rect -1367 -410 -1339 -382
rect -1301 -410 -1273 -382
rect -1235 -410 -1207 -382
rect -1169 -410 -1141 -382
rect -1103 -410 -1075 -382
rect -1037 -410 -1009 -382
rect -971 -410 -943 -382
rect -905 -410 -877 -382
rect -839 -410 -811 -382
rect -773 -410 -745 -382
rect -707 -410 -679 -382
rect -641 -410 -613 -382
rect -575 -410 -547 -382
rect -509 -410 -481 -382
rect -443 -410 -415 -382
rect -377 -410 -349 -382
rect -311 -410 -283 -382
rect -245 -410 -217 -382
rect -179 -410 -151 -382
rect -113 -410 -85 -382
rect -47 -410 -19 -382
rect 19 -410 47 -382
rect 85 -410 113 -382
rect 151 -410 179 -382
rect 217 -410 245 -382
rect 283 -410 311 -382
rect 349 -410 377 -382
rect 415 -410 443 -382
rect 481 -410 509 -382
rect 547 -410 575 -382
rect 613 -410 641 -382
rect 679 -410 707 -382
rect 745 -410 773 -382
rect 811 -410 839 -382
rect 877 -410 905 -382
rect 943 -410 971 -382
rect 1009 -410 1037 -382
rect 1075 -410 1103 -382
rect 1141 -410 1169 -382
rect 1207 -410 1235 -382
rect 1273 -410 1301 -382
rect 1339 -410 1367 -382
rect 1405 -410 1433 -382
rect 1471 -410 1499 -382
rect 1537 -410 1565 -382
rect 1603 -410 1631 -382
rect 1669 -410 1697 -382
rect 1735 -410 1763 -382
rect 1801 -410 1829 -382
rect 1867 -410 1895 -382
rect 1933 -410 1961 -382
rect 1999 -410 2027 -382
rect 2065 -410 2093 -382
rect 2131 -410 2159 -382
rect 2197 -410 2225 -382
rect 2263 -410 2291 -382
rect 2329 -410 2357 -382
rect 2395 -410 2423 -382
rect 2461 -410 2489 -382
rect 2527 -410 2555 -382
rect 2593 -410 2621 -382
rect 2659 -410 2687 -382
rect 2725 -410 2753 -382
rect 2791 -410 2819 -382
rect 2857 -410 2885 -382
rect 2923 -410 2951 -382
rect 2989 -410 3017 -382
rect 3055 -410 3083 -382
rect 3121 -410 3149 -382
rect 3187 -410 3215 -382
rect 3253 -410 3281 -382
rect 3319 -410 3347 -382
rect 3385 -410 3413 -382
rect 3451 -410 3479 -382
rect 3517 -410 3545 -382
rect 3583 -410 3611 -382
rect 3649 -410 3677 -382
rect 3715 -410 3743 -382
rect 3781 -410 3809 -382
rect 3847 -410 3875 -382
rect -3875 -476 -3847 -448
rect -3809 -476 -3781 -448
rect -3743 -476 -3715 -448
rect -3677 -476 -3649 -448
rect -3611 -476 -3583 -448
rect -3545 -476 -3517 -448
rect -3479 -476 -3451 -448
rect -3413 -476 -3385 -448
rect -3347 -476 -3319 -448
rect -3281 -476 -3253 -448
rect -3215 -476 -3187 -448
rect -3149 -476 -3121 -448
rect -3083 -476 -3055 -448
rect -3017 -476 -2989 -448
rect -2951 -476 -2923 -448
rect -2885 -476 -2857 -448
rect -2819 -476 -2791 -448
rect -2753 -476 -2725 -448
rect -2687 -476 -2659 -448
rect -2621 -476 -2593 -448
rect -2555 -476 -2527 -448
rect -2489 -476 -2461 -448
rect -2423 -476 -2395 -448
rect -2357 -476 -2329 -448
rect -2291 -476 -2263 -448
rect -2225 -476 -2197 -448
rect -2159 -476 -2131 -448
rect -2093 -476 -2065 -448
rect -2027 -476 -1999 -448
rect -1961 -476 -1933 -448
rect -1895 -476 -1867 -448
rect -1829 -476 -1801 -448
rect -1763 -476 -1735 -448
rect -1697 -476 -1669 -448
rect -1631 -476 -1603 -448
rect -1565 -476 -1537 -448
rect -1499 -476 -1471 -448
rect -1433 -476 -1405 -448
rect -1367 -476 -1339 -448
rect -1301 -476 -1273 -448
rect -1235 -476 -1207 -448
rect -1169 -476 -1141 -448
rect -1103 -476 -1075 -448
rect -1037 -476 -1009 -448
rect -971 -476 -943 -448
rect -905 -476 -877 -448
rect -839 -476 -811 -448
rect -773 -476 -745 -448
rect -707 -476 -679 -448
rect -641 -476 -613 -448
rect -575 -476 -547 -448
rect -509 -476 -481 -448
rect -443 -476 -415 -448
rect -377 -476 -349 -448
rect -311 -476 -283 -448
rect -245 -476 -217 -448
rect -179 -476 -151 -448
rect -113 -476 -85 -448
rect -47 -476 -19 -448
rect 19 -476 47 -448
rect 85 -476 113 -448
rect 151 -476 179 -448
rect 217 -476 245 -448
rect 283 -476 311 -448
rect 349 -476 377 -448
rect 415 -476 443 -448
rect 481 -476 509 -448
rect 547 -476 575 -448
rect 613 -476 641 -448
rect 679 -476 707 -448
rect 745 -476 773 -448
rect 811 -476 839 -448
rect 877 -476 905 -448
rect 943 -476 971 -448
rect 1009 -476 1037 -448
rect 1075 -476 1103 -448
rect 1141 -476 1169 -448
rect 1207 -476 1235 -448
rect 1273 -476 1301 -448
rect 1339 -476 1367 -448
rect 1405 -476 1433 -448
rect 1471 -476 1499 -448
rect 1537 -476 1565 -448
rect 1603 -476 1631 -448
rect 1669 -476 1697 -448
rect 1735 -476 1763 -448
rect 1801 -476 1829 -448
rect 1867 -476 1895 -448
rect 1933 -476 1961 -448
rect 1999 -476 2027 -448
rect 2065 -476 2093 -448
rect 2131 -476 2159 -448
rect 2197 -476 2225 -448
rect 2263 -476 2291 -448
rect 2329 -476 2357 -448
rect 2395 -476 2423 -448
rect 2461 -476 2489 -448
rect 2527 -476 2555 -448
rect 2593 -476 2621 -448
rect 2659 -476 2687 -448
rect 2725 -476 2753 -448
rect 2791 -476 2819 -448
rect 2857 -476 2885 -448
rect 2923 -476 2951 -448
rect 2989 -476 3017 -448
rect 3055 -476 3083 -448
rect 3121 -476 3149 -448
rect 3187 -476 3215 -448
rect 3253 -476 3281 -448
rect 3319 -476 3347 -448
rect 3385 -476 3413 -448
rect 3451 -476 3479 -448
rect 3517 -476 3545 -448
rect 3583 -476 3611 -448
rect 3649 -476 3677 -448
rect 3715 -476 3743 -448
rect 3781 -476 3809 -448
rect 3847 -476 3875 -448
rect -3875 -542 -3847 -514
rect -3809 -542 -3781 -514
rect -3743 -542 -3715 -514
rect -3677 -542 -3649 -514
rect -3611 -542 -3583 -514
rect -3545 -542 -3517 -514
rect -3479 -542 -3451 -514
rect -3413 -542 -3385 -514
rect -3347 -542 -3319 -514
rect -3281 -542 -3253 -514
rect -3215 -542 -3187 -514
rect -3149 -542 -3121 -514
rect -3083 -542 -3055 -514
rect -3017 -542 -2989 -514
rect -2951 -542 -2923 -514
rect -2885 -542 -2857 -514
rect -2819 -542 -2791 -514
rect -2753 -542 -2725 -514
rect -2687 -542 -2659 -514
rect -2621 -542 -2593 -514
rect -2555 -542 -2527 -514
rect -2489 -542 -2461 -514
rect -2423 -542 -2395 -514
rect -2357 -542 -2329 -514
rect -2291 -542 -2263 -514
rect -2225 -542 -2197 -514
rect -2159 -542 -2131 -514
rect -2093 -542 -2065 -514
rect -2027 -542 -1999 -514
rect -1961 -542 -1933 -514
rect -1895 -542 -1867 -514
rect -1829 -542 -1801 -514
rect -1763 -542 -1735 -514
rect -1697 -542 -1669 -514
rect -1631 -542 -1603 -514
rect -1565 -542 -1537 -514
rect -1499 -542 -1471 -514
rect -1433 -542 -1405 -514
rect -1367 -542 -1339 -514
rect -1301 -542 -1273 -514
rect -1235 -542 -1207 -514
rect -1169 -542 -1141 -514
rect -1103 -542 -1075 -514
rect -1037 -542 -1009 -514
rect -971 -542 -943 -514
rect -905 -542 -877 -514
rect -839 -542 -811 -514
rect -773 -542 -745 -514
rect -707 -542 -679 -514
rect -641 -542 -613 -514
rect -575 -542 -547 -514
rect -509 -542 -481 -514
rect -443 -542 -415 -514
rect -377 -542 -349 -514
rect -311 -542 -283 -514
rect -245 -542 -217 -514
rect -179 -542 -151 -514
rect -113 -542 -85 -514
rect -47 -542 -19 -514
rect 19 -542 47 -514
rect 85 -542 113 -514
rect 151 -542 179 -514
rect 217 -542 245 -514
rect 283 -542 311 -514
rect 349 -542 377 -514
rect 415 -542 443 -514
rect 481 -542 509 -514
rect 547 -542 575 -514
rect 613 -542 641 -514
rect 679 -542 707 -514
rect 745 -542 773 -514
rect 811 -542 839 -514
rect 877 -542 905 -514
rect 943 -542 971 -514
rect 1009 -542 1037 -514
rect 1075 -542 1103 -514
rect 1141 -542 1169 -514
rect 1207 -542 1235 -514
rect 1273 -542 1301 -514
rect 1339 -542 1367 -514
rect 1405 -542 1433 -514
rect 1471 -542 1499 -514
rect 1537 -542 1565 -514
rect 1603 -542 1631 -514
rect 1669 -542 1697 -514
rect 1735 -542 1763 -514
rect 1801 -542 1829 -514
rect 1867 -542 1895 -514
rect 1933 -542 1961 -514
rect 1999 -542 2027 -514
rect 2065 -542 2093 -514
rect 2131 -542 2159 -514
rect 2197 -542 2225 -514
rect 2263 -542 2291 -514
rect 2329 -542 2357 -514
rect 2395 -542 2423 -514
rect 2461 -542 2489 -514
rect 2527 -542 2555 -514
rect 2593 -542 2621 -514
rect 2659 -542 2687 -514
rect 2725 -542 2753 -514
rect 2791 -542 2819 -514
rect 2857 -542 2885 -514
rect 2923 -542 2951 -514
rect 2989 -542 3017 -514
rect 3055 -542 3083 -514
rect 3121 -542 3149 -514
rect 3187 -542 3215 -514
rect 3253 -542 3281 -514
rect 3319 -542 3347 -514
rect 3385 -542 3413 -514
rect 3451 -542 3479 -514
rect 3517 -542 3545 -514
rect 3583 -542 3611 -514
rect 3649 -542 3677 -514
rect 3715 -542 3743 -514
rect 3781 -542 3809 -514
rect 3847 -542 3875 -514
rect -3875 -608 -3847 -580
rect -3809 -608 -3781 -580
rect -3743 -608 -3715 -580
rect -3677 -608 -3649 -580
rect -3611 -608 -3583 -580
rect -3545 -608 -3517 -580
rect -3479 -608 -3451 -580
rect -3413 -608 -3385 -580
rect -3347 -608 -3319 -580
rect -3281 -608 -3253 -580
rect -3215 -608 -3187 -580
rect -3149 -608 -3121 -580
rect -3083 -608 -3055 -580
rect -3017 -608 -2989 -580
rect -2951 -608 -2923 -580
rect -2885 -608 -2857 -580
rect -2819 -608 -2791 -580
rect -2753 -608 -2725 -580
rect -2687 -608 -2659 -580
rect -2621 -608 -2593 -580
rect -2555 -608 -2527 -580
rect -2489 -608 -2461 -580
rect -2423 -608 -2395 -580
rect -2357 -608 -2329 -580
rect -2291 -608 -2263 -580
rect -2225 -608 -2197 -580
rect -2159 -608 -2131 -580
rect -2093 -608 -2065 -580
rect -2027 -608 -1999 -580
rect -1961 -608 -1933 -580
rect -1895 -608 -1867 -580
rect -1829 -608 -1801 -580
rect -1763 -608 -1735 -580
rect -1697 -608 -1669 -580
rect -1631 -608 -1603 -580
rect -1565 -608 -1537 -580
rect -1499 -608 -1471 -580
rect -1433 -608 -1405 -580
rect -1367 -608 -1339 -580
rect -1301 -608 -1273 -580
rect -1235 -608 -1207 -580
rect -1169 -608 -1141 -580
rect -1103 -608 -1075 -580
rect -1037 -608 -1009 -580
rect -971 -608 -943 -580
rect -905 -608 -877 -580
rect -839 -608 -811 -580
rect -773 -608 -745 -580
rect -707 -608 -679 -580
rect -641 -608 -613 -580
rect -575 -608 -547 -580
rect -509 -608 -481 -580
rect -443 -608 -415 -580
rect -377 -608 -349 -580
rect -311 -608 -283 -580
rect -245 -608 -217 -580
rect -179 -608 -151 -580
rect -113 -608 -85 -580
rect -47 -608 -19 -580
rect 19 -608 47 -580
rect 85 -608 113 -580
rect 151 -608 179 -580
rect 217 -608 245 -580
rect 283 -608 311 -580
rect 349 -608 377 -580
rect 415 -608 443 -580
rect 481 -608 509 -580
rect 547 -608 575 -580
rect 613 -608 641 -580
rect 679 -608 707 -580
rect 745 -608 773 -580
rect 811 -608 839 -580
rect 877 -608 905 -580
rect 943 -608 971 -580
rect 1009 -608 1037 -580
rect 1075 -608 1103 -580
rect 1141 -608 1169 -580
rect 1207 -608 1235 -580
rect 1273 -608 1301 -580
rect 1339 -608 1367 -580
rect 1405 -608 1433 -580
rect 1471 -608 1499 -580
rect 1537 -608 1565 -580
rect 1603 -608 1631 -580
rect 1669 -608 1697 -580
rect 1735 -608 1763 -580
rect 1801 -608 1829 -580
rect 1867 -608 1895 -580
rect 1933 -608 1961 -580
rect 1999 -608 2027 -580
rect 2065 -608 2093 -580
rect 2131 -608 2159 -580
rect 2197 -608 2225 -580
rect 2263 -608 2291 -580
rect 2329 -608 2357 -580
rect 2395 -608 2423 -580
rect 2461 -608 2489 -580
rect 2527 -608 2555 -580
rect 2593 -608 2621 -580
rect 2659 -608 2687 -580
rect 2725 -608 2753 -580
rect 2791 -608 2819 -580
rect 2857 -608 2885 -580
rect 2923 -608 2951 -580
rect 2989 -608 3017 -580
rect 3055 -608 3083 -580
rect 3121 -608 3149 -580
rect 3187 -608 3215 -580
rect 3253 -608 3281 -580
rect 3319 -608 3347 -580
rect 3385 -608 3413 -580
rect 3451 -608 3479 -580
rect 3517 -608 3545 -580
rect 3583 -608 3611 -580
rect 3649 -608 3677 -580
rect 3715 -608 3743 -580
rect 3781 -608 3809 -580
rect 3847 -608 3875 -580
rect -3875 -674 -3847 -646
rect -3809 -674 -3781 -646
rect -3743 -674 -3715 -646
rect -3677 -674 -3649 -646
rect -3611 -674 -3583 -646
rect -3545 -674 -3517 -646
rect -3479 -674 -3451 -646
rect -3413 -674 -3385 -646
rect -3347 -674 -3319 -646
rect -3281 -674 -3253 -646
rect -3215 -674 -3187 -646
rect -3149 -674 -3121 -646
rect -3083 -674 -3055 -646
rect -3017 -674 -2989 -646
rect -2951 -674 -2923 -646
rect -2885 -674 -2857 -646
rect -2819 -674 -2791 -646
rect -2753 -674 -2725 -646
rect -2687 -674 -2659 -646
rect -2621 -674 -2593 -646
rect -2555 -674 -2527 -646
rect -2489 -674 -2461 -646
rect -2423 -674 -2395 -646
rect -2357 -674 -2329 -646
rect -2291 -674 -2263 -646
rect -2225 -674 -2197 -646
rect -2159 -674 -2131 -646
rect -2093 -674 -2065 -646
rect -2027 -674 -1999 -646
rect -1961 -674 -1933 -646
rect -1895 -674 -1867 -646
rect -1829 -674 -1801 -646
rect -1763 -674 -1735 -646
rect -1697 -674 -1669 -646
rect -1631 -674 -1603 -646
rect -1565 -674 -1537 -646
rect -1499 -674 -1471 -646
rect -1433 -674 -1405 -646
rect -1367 -674 -1339 -646
rect -1301 -674 -1273 -646
rect -1235 -674 -1207 -646
rect -1169 -674 -1141 -646
rect -1103 -674 -1075 -646
rect -1037 -674 -1009 -646
rect -971 -674 -943 -646
rect -905 -674 -877 -646
rect -839 -674 -811 -646
rect -773 -674 -745 -646
rect -707 -674 -679 -646
rect -641 -674 -613 -646
rect -575 -674 -547 -646
rect -509 -674 -481 -646
rect -443 -674 -415 -646
rect -377 -674 -349 -646
rect -311 -674 -283 -646
rect -245 -674 -217 -646
rect -179 -674 -151 -646
rect -113 -674 -85 -646
rect -47 -674 -19 -646
rect 19 -674 47 -646
rect 85 -674 113 -646
rect 151 -674 179 -646
rect 217 -674 245 -646
rect 283 -674 311 -646
rect 349 -674 377 -646
rect 415 -674 443 -646
rect 481 -674 509 -646
rect 547 -674 575 -646
rect 613 -674 641 -646
rect 679 -674 707 -646
rect 745 -674 773 -646
rect 811 -674 839 -646
rect 877 -674 905 -646
rect 943 -674 971 -646
rect 1009 -674 1037 -646
rect 1075 -674 1103 -646
rect 1141 -674 1169 -646
rect 1207 -674 1235 -646
rect 1273 -674 1301 -646
rect 1339 -674 1367 -646
rect 1405 -674 1433 -646
rect 1471 -674 1499 -646
rect 1537 -674 1565 -646
rect 1603 -674 1631 -646
rect 1669 -674 1697 -646
rect 1735 -674 1763 -646
rect 1801 -674 1829 -646
rect 1867 -674 1895 -646
rect 1933 -674 1961 -646
rect 1999 -674 2027 -646
rect 2065 -674 2093 -646
rect 2131 -674 2159 -646
rect 2197 -674 2225 -646
rect 2263 -674 2291 -646
rect 2329 -674 2357 -646
rect 2395 -674 2423 -646
rect 2461 -674 2489 -646
rect 2527 -674 2555 -646
rect 2593 -674 2621 -646
rect 2659 -674 2687 -646
rect 2725 -674 2753 -646
rect 2791 -674 2819 -646
rect 2857 -674 2885 -646
rect 2923 -674 2951 -646
rect 2989 -674 3017 -646
rect 3055 -674 3083 -646
rect 3121 -674 3149 -646
rect 3187 -674 3215 -646
rect 3253 -674 3281 -646
rect 3319 -674 3347 -646
rect 3385 -674 3413 -646
rect 3451 -674 3479 -646
rect 3517 -674 3545 -646
rect 3583 -674 3611 -646
rect 3649 -674 3677 -646
rect 3715 -674 3743 -646
rect 3781 -674 3809 -646
rect 3847 -674 3875 -646
rect -3875 -740 -3847 -712
rect -3809 -740 -3781 -712
rect -3743 -740 -3715 -712
rect -3677 -740 -3649 -712
rect -3611 -740 -3583 -712
rect -3545 -740 -3517 -712
rect -3479 -740 -3451 -712
rect -3413 -740 -3385 -712
rect -3347 -740 -3319 -712
rect -3281 -740 -3253 -712
rect -3215 -740 -3187 -712
rect -3149 -740 -3121 -712
rect -3083 -740 -3055 -712
rect -3017 -740 -2989 -712
rect -2951 -740 -2923 -712
rect -2885 -740 -2857 -712
rect -2819 -740 -2791 -712
rect -2753 -740 -2725 -712
rect -2687 -740 -2659 -712
rect -2621 -740 -2593 -712
rect -2555 -740 -2527 -712
rect -2489 -740 -2461 -712
rect -2423 -740 -2395 -712
rect -2357 -740 -2329 -712
rect -2291 -740 -2263 -712
rect -2225 -740 -2197 -712
rect -2159 -740 -2131 -712
rect -2093 -740 -2065 -712
rect -2027 -740 -1999 -712
rect -1961 -740 -1933 -712
rect -1895 -740 -1867 -712
rect -1829 -740 -1801 -712
rect -1763 -740 -1735 -712
rect -1697 -740 -1669 -712
rect -1631 -740 -1603 -712
rect -1565 -740 -1537 -712
rect -1499 -740 -1471 -712
rect -1433 -740 -1405 -712
rect -1367 -740 -1339 -712
rect -1301 -740 -1273 -712
rect -1235 -740 -1207 -712
rect -1169 -740 -1141 -712
rect -1103 -740 -1075 -712
rect -1037 -740 -1009 -712
rect -971 -740 -943 -712
rect -905 -740 -877 -712
rect -839 -740 -811 -712
rect -773 -740 -745 -712
rect -707 -740 -679 -712
rect -641 -740 -613 -712
rect -575 -740 -547 -712
rect -509 -740 -481 -712
rect -443 -740 -415 -712
rect -377 -740 -349 -712
rect -311 -740 -283 -712
rect -245 -740 -217 -712
rect -179 -740 -151 -712
rect -113 -740 -85 -712
rect -47 -740 -19 -712
rect 19 -740 47 -712
rect 85 -740 113 -712
rect 151 -740 179 -712
rect 217 -740 245 -712
rect 283 -740 311 -712
rect 349 -740 377 -712
rect 415 -740 443 -712
rect 481 -740 509 -712
rect 547 -740 575 -712
rect 613 -740 641 -712
rect 679 -740 707 -712
rect 745 -740 773 -712
rect 811 -740 839 -712
rect 877 -740 905 -712
rect 943 -740 971 -712
rect 1009 -740 1037 -712
rect 1075 -740 1103 -712
rect 1141 -740 1169 -712
rect 1207 -740 1235 -712
rect 1273 -740 1301 -712
rect 1339 -740 1367 -712
rect 1405 -740 1433 -712
rect 1471 -740 1499 -712
rect 1537 -740 1565 -712
rect 1603 -740 1631 -712
rect 1669 -740 1697 -712
rect 1735 -740 1763 -712
rect 1801 -740 1829 -712
rect 1867 -740 1895 -712
rect 1933 -740 1961 -712
rect 1999 -740 2027 -712
rect 2065 -740 2093 -712
rect 2131 -740 2159 -712
rect 2197 -740 2225 -712
rect 2263 -740 2291 -712
rect 2329 -740 2357 -712
rect 2395 -740 2423 -712
rect 2461 -740 2489 -712
rect 2527 -740 2555 -712
rect 2593 -740 2621 -712
rect 2659 -740 2687 -712
rect 2725 -740 2753 -712
rect 2791 -740 2819 -712
rect 2857 -740 2885 -712
rect 2923 -740 2951 -712
rect 2989 -740 3017 -712
rect 3055 -740 3083 -712
rect 3121 -740 3149 -712
rect 3187 -740 3215 -712
rect 3253 -740 3281 -712
rect 3319 -740 3347 -712
rect 3385 -740 3413 -712
rect 3451 -740 3479 -712
rect 3517 -740 3545 -712
rect 3583 -740 3611 -712
rect 3649 -740 3677 -712
rect 3715 -740 3743 -712
rect 3781 -740 3809 -712
rect 3847 -740 3875 -712
<< metal5 >>
rect -3883 740 3883 748
rect -3883 712 -3875 740
rect -3847 712 -3809 740
rect -3781 712 -3743 740
rect -3715 712 -3677 740
rect -3649 712 -3611 740
rect -3583 712 -3545 740
rect -3517 712 -3479 740
rect -3451 712 -3413 740
rect -3385 712 -3347 740
rect -3319 712 -3281 740
rect -3253 712 -3215 740
rect -3187 712 -3149 740
rect -3121 712 -3083 740
rect -3055 712 -3017 740
rect -2989 712 -2951 740
rect -2923 712 -2885 740
rect -2857 712 -2819 740
rect -2791 712 -2753 740
rect -2725 712 -2687 740
rect -2659 712 -2621 740
rect -2593 712 -2555 740
rect -2527 712 -2489 740
rect -2461 712 -2423 740
rect -2395 712 -2357 740
rect -2329 712 -2291 740
rect -2263 712 -2225 740
rect -2197 712 -2159 740
rect -2131 712 -2093 740
rect -2065 712 -2027 740
rect -1999 712 -1961 740
rect -1933 712 -1895 740
rect -1867 712 -1829 740
rect -1801 712 -1763 740
rect -1735 712 -1697 740
rect -1669 712 -1631 740
rect -1603 712 -1565 740
rect -1537 712 -1499 740
rect -1471 712 -1433 740
rect -1405 712 -1367 740
rect -1339 712 -1301 740
rect -1273 712 -1235 740
rect -1207 712 -1169 740
rect -1141 712 -1103 740
rect -1075 712 -1037 740
rect -1009 712 -971 740
rect -943 712 -905 740
rect -877 712 -839 740
rect -811 712 -773 740
rect -745 712 -707 740
rect -679 712 -641 740
rect -613 712 -575 740
rect -547 712 -509 740
rect -481 712 -443 740
rect -415 712 -377 740
rect -349 712 -311 740
rect -283 712 -245 740
rect -217 712 -179 740
rect -151 712 -113 740
rect -85 712 -47 740
rect -19 712 19 740
rect 47 712 85 740
rect 113 712 151 740
rect 179 712 217 740
rect 245 712 283 740
rect 311 712 349 740
rect 377 712 415 740
rect 443 712 481 740
rect 509 712 547 740
rect 575 712 613 740
rect 641 712 679 740
rect 707 712 745 740
rect 773 712 811 740
rect 839 712 877 740
rect 905 712 943 740
rect 971 712 1009 740
rect 1037 712 1075 740
rect 1103 712 1141 740
rect 1169 712 1207 740
rect 1235 712 1273 740
rect 1301 712 1339 740
rect 1367 712 1405 740
rect 1433 712 1471 740
rect 1499 712 1537 740
rect 1565 712 1603 740
rect 1631 712 1669 740
rect 1697 712 1735 740
rect 1763 712 1801 740
rect 1829 712 1867 740
rect 1895 712 1933 740
rect 1961 712 1999 740
rect 2027 712 2065 740
rect 2093 712 2131 740
rect 2159 712 2197 740
rect 2225 712 2263 740
rect 2291 712 2329 740
rect 2357 712 2395 740
rect 2423 712 2461 740
rect 2489 712 2527 740
rect 2555 712 2593 740
rect 2621 712 2659 740
rect 2687 712 2725 740
rect 2753 712 2791 740
rect 2819 712 2857 740
rect 2885 712 2923 740
rect 2951 712 2989 740
rect 3017 712 3055 740
rect 3083 712 3121 740
rect 3149 712 3187 740
rect 3215 712 3253 740
rect 3281 712 3319 740
rect 3347 712 3385 740
rect 3413 712 3451 740
rect 3479 712 3517 740
rect 3545 712 3583 740
rect 3611 712 3649 740
rect 3677 712 3715 740
rect 3743 712 3781 740
rect 3809 712 3847 740
rect 3875 712 3883 740
rect -3883 674 3883 712
rect -3883 646 -3875 674
rect -3847 646 -3809 674
rect -3781 646 -3743 674
rect -3715 646 -3677 674
rect -3649 646 -3611 674
rect -3583 646 -3545 674
rect -3517 646 -3479 674
rect -3451 646 -3413 674
rect -3385 646 -3347 674
rect -3319 646 -3281 674
rect -3253 646 -3215 674
rect -3187 646 -3149 674
rect -3121 646 -3083 674
rect -3055 646 -3017 674
rect -2989 646 -2951 674
rect -2923 646 -2885 674
rect -2857 646 -2819 674
rect -2791 646 -2753 674
rect -2725 646 -2687 674
rect -2659 646 -2621 674
rect -2593 646 -2555 674
rect -2527 646 -2489 674
rect -2461 646 -2423 674
rect -2395 646 -2357 674
rect -2329 646 -2291 674
rect -2263 646 -2225 674
rect -2197 646 -2159 674
rect -2131 646 -2093 674
rect -2065 646 -2027 674
rect -1999 646 -1961 674
rect -1933 646 -1895 674
rect -1867 646 -1829 674
rect -1801 646 -1763 674
rect -1735 646 -1697 674
rect -1669 646 -1631 674
rect -1603 646 -1565 674
rect -1537 646 -1499 674
rect -1471 646 -1433 674
rect -1405 646 -1367 674
rect -1339 646 -1301 674
rect -1273 646 -1235 674
rect -1207 646 -1169 674
rect -1141 646 -1103 674
rect -1075 646 -1037 674
rect -1009 646 -971 674
rect -943 646 -905 674
rect -877 646 -839 674
rect -811 646 -773 674
rect -745 646 -707 674
rect -679 646 -641 674
rect -613 646 -575 674
rect -547 646 -509 674
rect -481 646 -443 674
rect -415 646 -377 674
rect -349 646 -311 674
rect -283 646 -245 674
rect -217 646 -179 674
rect -151 646 -113 674
rect -85 646 -47 674
rect -19 646 19 674
rect 47 646 85 674
rect 113 646 151 674
rect 179 646 217 674
rect 245 646 283 674
rect 311 646 349 674
rect 377 646 415 674
rect 443 646 481 674
rect 509 646 547 674
rect 575 646 613 674
rect 641 646 679 674
rect 707 646 745 674
rect 773 646 811 674
rect 839 646 877 674
rect 905 646 943 674
rect 971 646 1009 674
rect 1037 646 1075 674
rect 1103 646 1141 674
rect 1169 646 1207 674
rect 1235 646 1273 674
rect 1301 646 1339 674
rect 1367 646 1405 674
rect 1433 646 1471 674
rect 1499 646 1537 674
rect 1565 646 1603 674
rect 1631 646 1669 674
rect 1697 646 1735 674
rect 1763 646 1801 674
rect 1829 646 1867 674
rect 1895 646 1933 674
rect 1961 646 1999 674
rect 2027 646 2065 674
rect 2093 646 2131 674
rect 2159 646 2197 674
rect 2225 646 2263 674
rect 2291 646 2329 674
rect 2357 646 2395 674
rect 2423 646 2461 674
rect 2489 646 2527 674
rect 2555 646 2593 674
rect 2621 646 2659 674
rect 2687 646 2725 674
rect 2753 646 2791 674
rect 2819 646 2857 674
rect 2885 646 2923 674
rect 2951 646 2989 674
rect 3017 646 3055 674
rect 3083 646 3121 674
rect 3149 646 3187 674
rect 3215 646 3253 674
rect 3281 646 3319 674
rect 3347 646 3385 674
rect 3413 646 3451 674
rect 3479 646 3517 674
rect 3545 646 3583 674
rect 3611 646 3649 674
rect 3677 646 3715 674
rect 3743 646 3781 674
rect 3809 646 3847 674
rect 3875 646 3883 674
rect -3883 608 3883 646
rect -3883 580 -3875 608
rect -3847 580 -3809 608
rect -3781 580 -3743 608
rect -3715 580 -3677 608
rect -3649 580 -3611 608
rect -3583 580 -3545 608
rect -3517 580 -3479 608
rect -3451 580 -3413 608
rect -3385 580 -3347 608
rect -3319 580 -3281 608
rect -3253 580 -3215 608
rect -3187 580 -3149 608
rect -3121 580 -3083 608
rect -3055 580 -3017 608
rect -2989 580 -2951 608
rect -2923 580 -2885 608
rect -2857 580 -2819 608
rect -2791 580 -2753 608
rect -2725 580 -2687 608
rect -2659 580 -2621 608
rect -2593 580 -2555 608
rect -2527 580 -2489 608
rect -2461 580 -2423 608
rect -2395 580 -2357 608
rect -2329 580 -2291 608
rect -2263 580 -2225 608
rect -2197 580 -2159 608
rect -2131 580 -2093 608
rect -2065 580 -2027 608
rect -1999 580 -1961 608
rect -1933 580 -1895 608
rect -1867 580 -1829 608
rect -1801 580 -1763 608
rect -1735 580 -1697 608
rect -1669 580 -1631 608
rect -1603 580 -1565 608
rect -1537 580 -1499 608
rect -1471 580 -1433 608
rect -1405 580 -1367 608
rect -1339 580 -1301 608
rect -1273 580 -1235 608
rect -1207 580 -1169 608
rect -1141 580 -1103 608
rect -1075 580 -1037 608
rect -1009 580 -971 608
rect -943 580 -905 608
rect -877 580 -839 608
rect -811 580 -773 608
rect -745 580 -707 608
rect -679 580 -641 608
rect -613 580 -575 608
rect -547 580 -509 608
rect -481 580 -443 608
rect -415 580 -377 608
rect -349 580 -311 608
rect -283 580 -245 608
rect -217 580 -179 608
rect -151 580 -113 608
rect -85 580 -47 608
rect -19 580 19 608
rect 47 580 85 608
rect 113 580 151 608
rect 179 580 217 608
rect 245 580 283 608
rect 311 580 349 608
rect 377 580 415 608
rect 443 580 481 608
rect 509 580 547 608
rect 575 580 613 608
rect 641 580 679 608
rect 707 580 745 608
rect 773 580 811 608
rect 839 580 877 608
rect 905 580 943 608
rect 971 580 1009 608
rect 1037 580 1075 608
rect 1103 580 1141 608
rect 1169 580 1207 608
rect 1235 580 1273 608
rect 1301 580 1339 608
rect 1367 580 1405 608
rect 1433 580 1471 608
rect 1499 580 1537 608
rect 1565 580 1603 608
rect 1631 580 1669 608
rect 1697 580 1735 608
rect 1763 580 1801 608
rect 1829 580 1867 608
rect 1895 580 1933 608
rect 1961 580 1999 608
rect 2027 580 2065 608
rect 2093 580 2131 608
rect 2159 580 2197 608
rect 2225 580 2263 608
rect 2291 580 2329 608
rect 2357 580 2395 608
rect 2423 580 2461 608
rect 2489 580 2527 608
rect 2555 580 2593 608
rect 2621 580 2659 608
rect 2687 580 2725 608
rect 2753 580 2791 608
rect 2819 580 2857 608
rect 2885 580 2923 608
rect 2951 580 2989 608
rect 3017 580 3055 608
rect 3083 580 3121 608
rect 3149 580 3187 608
rect 3215 580 3253 608
rect 3281 580 3319 608
rect 3347 580 3385 608
rect 3413 580 3451 608
rect 3479 580 3517 608
rect 3545 580 3583 608
rect 3611 580 3649 608
rect 3677 580 3715 608
rect 3743 580 3781 608
rect 3809 580 3847 608
rect 3875 580 3883 608
rect -3883 542 3883 580
rect -3883 514 -3875 542
rect -3847 514 -3809 542
rect -3781 514 -3743 542
rect -3715 514 -3677 542
rect -3649 514 -3611 542
rect -3583 514 -3545 542
rect -3517 514 -3479 542
rect -3451 514 -3413 542
rect -3385 514 -3347 542
rect -3319 514 -3281 542
rect -3253 514 -3215 542
rect -3187 514 -3149 542
rect -3121 514 -3083 542
rect -3055 514 -3017 542
rect -2989 514 -2951 542
rect -2923 514 -2885 542
rect -2857 514 -2819 542
rect -2791 514 -2753 542
rect -2725 514 -2687 542
rect -2659 514 -2621 542
rect -2593 514 -2555 542
rect -2527 514 -2489 542
rect -2461 514 -2423 542
rect -2395 514 -2357 542
rect -2329 514 -2291 542
rect -2263 514 -2225 542
rect -2197 514 -2159 542
rect -2131 514 -2093 542
rect -2065 514 -2027 542
rect -1999 514 -1961 542
rect -1933 514 -1895 542
rect -1867 514 -1829 542
rect -1801 514 -1763 542
rect -1735 514 -1697 542
rect -1669 514 -1631 542
rect -1603 514 -1565 542
rect -1537 514 -1499 542
rect -1471 514 -1433 542
rect -1405 514 -1367 542
rect -1339 514 -1301 542
rect -1273 514 -1235 542
rect -1207 514 -1169 542
rect -1141 514 -1103 542
rect -1075 514 -1037 542
rect -1009 514 -971 542
rect -943 514 -905 542
rect -877 514 -839 542
rect -811 514 -773 542
rect -745 514 -707 542
rect -679 514 -641 542
rect -613 514 -575 542
rect -547 514 -509 542
rect -481 514 -443 542
rect -415 514 -377 542
rect -349 514 -311 542
rect -283 514 -245 542
rect -217 514 -179 542
rect -151 514 -113 542
rect -85 514 -47 542
rect -19 514 19 542
rect 47 514 85 542
rect 113 514 151 542
rect 179 514 217 542
rect 245 514 283 542
rect 311 514 349 542
rect 377 514 415 542
rect 443 514 481 542
rect 509 514 547 542
rect 575 514 613 542
rect 641 514 679 542
rect 707 514 745 542
rect 773 514 811 542
rect 839 514 877 542
rect 905 514 943 542
rect 971 514 1009 542
rect 1037 514 1075 542
rect 1103 514 1141 542
rect 1169 514 1207 542
rect 1235 514 1273 542
rect 1301 514 1339 542
rect 1367 514 1405 542
rect 1433 514 1471 542
rect 1499 514 1537 542
rect 1565 514 1603 542
rect 1631 514 1669 542
rect 1697 514 1735 542
rect 1763 514 1801 542
rect 1829 514 1867 542
rect 1895 514 1933 542
rect 1961 514 1999 542
rect 2027 514 2065 542
rect 2093 514 2131 542
rect 2159 514 2197 542
rect 2225 514 2263 542
rect 2291 514 2329 542
rect 2357 514 2395 542
rect 2423 514 2461 542
rect 2489 514 2527 542
rect 2555 514 2593 542
rect 2621 514 2659 542
rect 2687 514 2725 542
rect 2753 514 2791 542
rect 2819 514 2857 542
rect 2885 514 2923 542
rect 2951 514 2989 542
rect 3017 514 3055 542
rect 3083 514 3121 542
rect 3149 514 3187 542
rect 3215 514 3253 542
rect 3281 514 3319 542
rect 3347 514 3385 542
rect 3413 514 3451 542
rect 3479 514 3517 542
rect 3545 514 3583 542
rect 3611 514 3649 542
rect 3677 514 3715 542
rect 3743 514 3781 542
rect 3809 514 3847 542
rect 3875 514 3883 542
rect -3883 476 3883 514
rect -3883 448 -3875 476
rect -3847 448 -3809 476
rect -3781 448 -3743 476
rect -3715 448 -3677 476
rect -3649 448 -3611 476
rect -3583 448 -3545 476
rect -3517 448 -3479 476
rect -3451 448 -3413 476
rect -3385 448 -3347 476
rect -3319 448 -3281 476
rect -3253 448 -3215 476
rect -3187 448 -3149 476
rect -3121 448 -3083 476
rect -3055 448 -3017 476
rect -2989 448 -2951 476
rect -2923 448 -2885 476
rect -2857 448 -2819 476
rect -2791 448 -2753 476
rect -2725 448 -2687 476
rect -2659 448 -2621 476
rect -2593 448 -2555 476
rect -2527 448 -2489 476
rect -2461 448 -2423 476
rect -2395 448 -2357 476
rect -2329 448 -2291 476
rect -2263 448 -2225 476
rect -2197 448 -2159 476
rect -2131 448 -2093 476
rect -2065 448 -2027 476
rect -1999 448 -1961 476
rect -1933 448 -1895 476
rect -1867 448 -1829 476
rect -1801 448 -1763 476
rect -1735 448 -1697 476
rect -1669 448 -1631 476
rect -1603 448 -1565 476
rect -1537 448 -1499 476
rect -1471 448 -1433 476
rect -1405 448 -1367 476
rect -1339 448 -1301 476
rect -1273 448 -1235 476
rect -1207 448 -1169 476
rect -1141 448 -1103 476
rect -1075 448 -1037 476
rect -1009 448 -971 476
rect -943 448 -905 476
rect -877 448 -839 476
rect -811 448 -773 476
rect -745 448 -707 476
rect -679 448 -641 476
rect -613 448 -575 476
rect -547 448 -509 476
rect -481 448 -443 476
rect -415 448 -377 476
rect -349 448 -311 476
rect -283 448 -245 476
rect -217 448 -179 476
rect -151 448 -113 476
rect -85 448 -47 476
rect -19 448 19 476
rect 47 448 85 476
rect 113 448 151 476
rect 179 448 217 476
rect 245 448 283 476
rect 311 448 349 476
rect 377 448 415 476
rect 443 448 481 476
rect 509 448 547 476
rect 575 448 613 476
rect 641 448 679 476
rect 707 448 745 476
rect 773 448 811 476
rect 839 448 877 476
rect 905 448 943 476
rect 971 448 1009 476
rect 1037 448 1075 476
rect 1103 448 1141 476
rect 1169 448 1207 476
rect 1235 448 1273 476
rect 1301 448 1339 476
rect 1367 448 1405 476
rect 1433 448 1471 476
rect 1499 448 1537 476
rect 1565 448 1603 476
rect 1631 448 1669 476
rect 1697 448 1735 476
rect 1763 448 1801 476
rect 1829 448 1867 476
rect 1895 448 1933 476
rect 1961 448 1999 476
rect 2027 448 2065 476
rect 2093 448 2131 476
rect 2159 448 2197 476
rect 2225 448 2263 476
rect 2291 448 2329 476
rect 2357 448 2395 476
rect 2423 448 2461 476
rect 2489 448 2527 476
rect 2555 448 2593 476
rect 2621 448 2659 476
rect 2687 448 2725 476
rect 2753 448 2791 476
rect 2819 448 2857 476
rect 2885 448 2923 476
rect 2951 448 2989 476
rect 3017 448 3055 476
rect 3083 448 3121 476
rect 3149 448 3187 476
rect 3215 448 3253 476
rect 3281 448 3319 476
rect 3347 448 3385 476
rect 3413 448 3451 476
rect 3479 448 3517 476
rect 3545 448 3583 476
rect 3611 448 3649 476
rect 3677 448 3715 476
rect 3743 448 3781 476
rect 3809 448 3847 476
rect 3875 448 3883 476
rect -3883 410 3883 448
rect -3883 382 -3875 410
rect -3847 382 -3809 410
rect -3781 382 -3743 410
rect -3715 382 -3677 410
rect -3649 382 -3611 410
rect -3583 382 -3545 410
rect -3517 382 -3479 410
rect -3451 382 -3413 410
rect -3385 382 -3347 410
rect -3319 382 -3281 410
rect -3253 382 -3215 410
rect -3187 382 -3149 410
rect -3121 382 -3083 410
rect -3055 382 -3017 410
rect -2989 382 -2951 410
rect -2923 382 -2885 410
rect -2857 382 -2819 410
rect -2791 382 -2753 410
rect -2725 382 -2687 410
rect -2659 382 -2621 410
rect -2593 382 -2555 410
rect -2527 382 -2489 410
rect -2461 382 -2423 410
rect -2395 382 -2357 410
rect -2329 382 -2291 410
rect -2263 382 -2225 410
rect -2197 382 -2159 410
rect -2131 382 -2093 410
rect -2065 382 -2027 410
rect -1999 382 -1961 410
rect -1933 382 -1895 410
rect -1867 382 -1829 410
rect -1801 382 -1763 410
rect -1735 382 -1697 410
rect -1669 382 -1631 410
rect -1603 382 -1565 410
rect -1537 382 -1499 410
rect -1471 382 -1433 410
rect -1405 382 -1367 410
rect -1339 382 -1301 410
rect -1273 382 -1235 410
rect -1207 382 -1169 410
rect -1141 382 -1103 410
rect -1075 382 -1037 410
rect -1009 382 -971 410
rect -943 382 -905 410
rect -877 382 -839 410
rect -811 382 -773 410
rect -745 382 -707 410
rect -679 382 -641 410
rect -613 382 -575 410
rect -547 382 -509 410
rect -481 382 -443 410
rect -415 382 -377 410
rect -349 382 -311 410
rect -283 382 -245 410
rect -217 382 -179 410
rect -151 382 -113 410
rect -85 382 -47 410
rect -19 382 19 410
rect 47 382 85 410
rect 113 382 151 410
rect 179 382 217 410
rect 245 382 283 410
rect 311 382 349 410
rect 377 382 415 410
rect 443 382 481 410
rect 509 382 547 410
rect 575 382 613 410
rect 641 382 679 410
rect 707 382 745 410
rect 773 382 811 410
rect 839 382 877 410
rect 905 382 943 410
rect 971 382 1009 410
rect 1037 382 1075 410
rect 1103 382 1141 410
rect 1169 382 1207 410
rect 1235 382 1273 410
rect 1301 382 1339 410
rect 1367 382 1405 410
rect 1433 382 1471 410
rect 1499 382 1537 410
rect 1565 382 1603 410
rect 1631 382 1669 410
rect 1697 382 1735 410
rect 1763 382 1801 410
rect 1829 382 1867 410
rect 1895 382 1933 410
rect 1961 382 1999 410
rect 2027 382 2065 410
rect 2093 382 2131 410
rect 2159 382 2197 410
rect 2225 382 2263 410
rect 2291 382 2329 410
rect 2357 382 2395 410
rect 2423 382 2461 410
rect 2489 382 2527 410
rect 2555 382 2593 410
rect 2621 382 2659 410
rect 2687 382 2725 410
rect 2753 382 2791 410
rect 2819 382 2857 410
rect 2885 382 2923 410
rect 2951 382 2989 410
rect 3017 382 3055 410
rect 3083 382 3121 410
rect 3149 382 3187 410
rect 3215 382 3253 410
rect 3281 382 3319 410
rect 3347 382 3385 410
rect 3413 382 3451 410
rect 3479 382 3517 410
rect 3545 382 3583 410
rect 3611 382 3649 410
rect 3677 382 3715 410
rect 3743 382 3781 410
rect 3809 382 3847 410
rect 3875 382 3883 410
rect -3883 344 3883 382
rect -3883 316 -3875 344
rect -3847 316 -3809 344
rect -3781 316 -3743 344
rect -3715 316 -3677 344
rect -3649 316 -3611 344
rect -3583 316 -3545 344
rect -3517 316 -3479 344
rect -3451 316 -3413 344
rect -3385 316 -3347 344
rect -3319 316 -3281 344
rect -3253 316 -3215 344
rect -3187 316 -3149 344
rect -3121 316 -3083 344
rect -3055 316 -3017 344
rect -2989 316 -2951 344
rect -2923 316 -2885 344
rect -2857 316 -2819 344
rect -2791 316 -2753 344
rect -2725 316 -2687 344
rect -2659 316 -2621 344
rect -2593 316 -2555 344
rect -2527 316 -2489 344
rect -2461 316 -2423 344
rect -2395 316 -2357 344
rect -2329 316 -2291 344
rect -2263 316 -2225 344
rect -2197 316 -2159 344
rect -2131 316 -2093 344
rect -2065 316 -2027 344
rect -1999 316 -1961 344
rect -1933 316 -1895 344
rect -1867 316 -1829 344
rect -1801 316 -1763 344
rect -1735 316 -1697 344
rect -1669 316 -1631 344
rect -1603 316 -1565 344
rect -1537 316 -1499 344
rect -1471 316 -1433 344
rect -1405 316 -1367 344
rect -1339 316 -1301 344
rect -1273 316 -1235 344
rect -1207 316 -1169 344
rect -1141 316 -1103 344
rect -1075 316 -1037 344
rect -1009 316 -971 344
rect -943 316 -905 344
rect -877 316 -839 344
rect -811 316 -773 344
rect -745 316 -707 344
rect -679 316 -641 344
rect -613 316 -575 344
rect -547 316 -509 344
rect -481 316 -443 344
rect -415 316 -377 344
rect -349 316 -311 344
rect -283 316 -245 344
rect -217 316 -179 344
rect -151 316 -113 344
rect -85 316 -47 344
rect -19 316 19 344
rect 47 316 85 344
rect 113 316 151 344
rect 179 316 217 344
rect 245 316 283 344
rect 311 316 349 344
rect 377 316 415 344
rect 443 316 481 344
rect 509 316 547 344
rect 575 316 613 344
rect 641 316 679 344
rect 707 316 745 344
rect 773 316 811 344
rect 839 316 877 344
rect 905 316 943 344
rect 971 316 1009 344
rect 1037 316 1075 344
rect 1103 316 1141 344
rect 1169 316 1207 344
rect 1235 316 1273 344
rect 1301 316 1339 344
rect 1367 316 1405 344
rect 1433 316 1471 344
rect 1499 316 1537 344
rect 1565 316 1603 344
rect 1631 316 1669 344
rect 1697 316 1735 344
rect 1763 316 1801 344
rect 1829 316 1867 344
rect 1895 316 1933 344
rect 1961 316 1999 344
rect 2027 316 2065 344
rect 2093 316 2131 344
rect 2159 316 2197 344
rect 2225 316 2263 344
rect 2291 316 2329 344
rect 2357 316 2395 344
rect 2423 316 2461 344
rect 2489 316 2527 344
rect 2555 316 2593 344
rect 2621 316 2659 344
rect 2687 316 2725 344
rect 2753 316 2791 344
rect 2819 316 2857 344
rect 2885 316 2923 344
rect 2951 316 2989 344
rect 3017 316 3055 344
rect 3083 316 3121 344
rect 3149 316 3187 344
rect 3215 316 3253 344
rect 3281 316 3319 344
rect 3347 316 3385 344
rect 3413 316 3451 344
rect 3479 316 3517 344
rect 3545 316 3583 344
rect 3611 316 3649 344
rect 3677 316 3715 344
rect 3743 316 3781 344
rect 3809 316 3847 344
rect 3875 316 3883 344
rect -3883 278 3883 316
rect -3883 250 -3875 278
rect -3847 250 -3809 278
rect -3781 250 -3743 278
rect -3715 250 -3677 278
rect -3649 250 -3611 278
rect -3583 250 -3545 278
rect -3517 250 -3479 278
rect -3451 250 -3413 278
rect -3385 250 -3347 278
rect -3319 250 -3281 278
rect -3253 250 -3215 278
rect -3187 250 -3149 278
rect -3121 250 -3083 278
rect -3055 250 -3017 278
rect -2989 250 -2951 278
rect -2923 250 -2885 278
rect -2857 250 -2819 278
rect -2791 250 -2753 278
rect -2725 250 -2687 278
rect -2659 250 -2621 278
rect -2593 250 -2555 278
rect -2527 250 -2489 278
rect -2461 250 -2423 278
rect -2395 250 -2357 278
rect -2329 250 -2291 278
rect -2263 250 -2225 278
rect -2197 250 -2159 278
rect -2131 250 -2093 278
rect -2065 250 -2027 278
rect -1999 250 -1961 278
rect -1933 250 -1895 278
rect -1867 250 -1829 278
rect -1801 250 -1763 278
rect -1735 250 -1697 278
rect -1669 250 -1631 278
rect -1603 250 -1565 278
rect -1537 250 -1499 278
rect -1471 250 -1433 278
rect -1405 250 -1367 278
rect -1339 250 -1301 278
rect -1273 250 -1235 278
rect -1207 250 -1169 278
rect -1141 250 -1103 278
rect -1075 250 -1037 278
rect -1009 250 -971 278
rect -943 250 -905 278
rect -877 250 -839 278
rect -811 250 -773 278
rect -745 250 -707 278
rect -679 250 -641 278
rect -613 250 -575 278
rect -547 250 -509 278
rect -481 250 -443 278
rect -415 250 -377 278
rect -349 250 -311 278
rect -283 250 -245 278
rect -217 250 -179 278
rect -151 250 -113 278
rect -85 250 -47 278
rect -19 250 19 278
rect 47 250 85 278
rect 113 250 151 278
rect 179 250 217 278
rect 245 250 283 278
rect 311 250 349 278
rect 377 250 415 278
rect 443 250 481 278
rect 509 250 547 278
rect 575 250 613 278
rect 641 250 679 278
rect 707 250 745 278
rect 773 250 811 278
rect 839 250 877 278
rect 905 250 943 278
rect 971 250 1009 278
rect 1037 250 1075 278
rect 1103 250 1141 278
rect 1169 250 1207 278
rect 1235 250 1273 278
rect 1301 250 1339 278
rect 1367 250 1405 278
rect 1433 250 1471 278
rect 1499 250 1537 278
rect 1565 250 1603 278
rect 1631 250 1669 278
rect 1697 250 1735 278
rect 1763 250 1801 278
rect 1829 250 1867 278
rect 1895 250 1933 278
rect 1961 250 1999 278
rect 2027 250 2065 278
rect 2093 250 2131 278
rect 2159 250 2197 278
rect 2225 250 2263 278
rect 2291 250 2329 278
rect 2357 250 2395 278
rect 2423 250 2461 278
rect 2489 250 2527 278
rect 2555 250 2593 278
rect 2621 250 2659 278
rect 2687 250 2725 278
rect 2753 250 2791 278
rect 2819 250 2857 278
rect 2885 250 2923 278
rect 2951 250 2989 278
rect 3017 250 3055 278
rect 3083 250 3121 278
rect 3149 250 3187 278
rect 3215 250 3253 278
rect 3281 250 3319 278
rect 3347 250 3385 278
rect 3413 250 3451 278
rect 3479 250 3517 278
rect 3545 250 3583 278
rect 3611 250 3649 278
rect 3677 250 3715 278
rect 3743 250 3781 278
rect 3809 250 3847 278
rect 3875 250 3883 278
rect -3883 212 3883 250
rect -3883 184 -3875 212
rect -3847 184 -3809 212
rect -3781 184 -3743 212
rect -3715 184 -3677 212
rect -3649 184 -3611 212
rect -3583 184 -3545 212
rect -3517 184 -3479 212
rect -3451 184 -3413 212
rect -3385 184 -3347 212
rect -3319 184 -3281 212
rect -3253 184 -3215 212
rect -3187 184 -3149 212
rect -3121 184 -3083 212
rect -3055 184 -3017 212
rect -2989 184 -2951 212
rect -2923 184 -2885 212
rect -2857 184 -2819 212
rect -2791 184 -2753 212
rect -2725 184 -2687 212
rect -2659 184 -2621 212
rect -2593 184 -2555 212
rect -2527 184 -2489 212
rect -2461 184 -2423 212
rect -2395 184 -2357 212
rect -2329 184 -2291 212
rect -2263 184 -2225 212
rect -2197 184 -2159 212
rect -2131 184 -2093 212
rect -2065 184 -2027 212
rect -1999 184 -1961 212
rect -1933 184 -1895 212
rect -1867 184 -1829 212
rect -1801 184 -1763 212
rect -1735 184 -1697 212
rect -1669 184 -1631 212
rect -1603 184 -1565 212
rect -1537 184 -1499 212
rect -1471 184 -1433 212
rect -1405 184 -1367 212
rect -1339 184 -1301 212
rect -1273 184 -1235 212
rect -1207 184 -1169 212
rect -1141 184 -1103 212
rect -1075 184 -1037 212
rect -1009 184 -971 212
rect -943 184 -905 212
rect -877 184 -839 212
rect -811 184 -773 212
rect -745 184 -707 212
rect -679 184 -641 212
rect -613 184 -575 212
rect -547 184 -509 212
rect -481 184 -443 212
rect -415 184 -377 212
rect -349 184 -311 212
rect -283 184 -245 212
rect -217 184 -179 212
rect -151 184 -113 212
rect -85 184 -47 212
rect -19 184 19 212
rect 47 184 85 212
rect 113 184 151 212
rect 179 184 217 212
rect 245 184 283 212
rect 311 184 349 212
rect 377 184 415 212
rect 443 184 481 212
rect 509 184 547 212
rect 575 184 613 212
rect 641 184 679 212
rect 707 184 745 212
rect 773 184 811 212
rect 839 184 877 212
rect 905 184 943 212
rect 971 184 1009 212
rect 1037 184 1075 212
rect 1103 184 1141 212
rect 1169 184 1207 212
rect 1235 184 1273 212
rect 1301 184 1339 212
rect 1367 184 1405 212
rect 1433 184 1471 212
rect 1499 184 1537 212
rect 1565 184 1603 212
rect 1631 184 1669 212
rect 1697 184 1735 212
rect 1763 184 1801 212
rect 1829 184 1867 212
rect 1895 184 1933 212
rect 1961 184 1999 212
rect 2027 184 2065 212
rect 2093 184 2131 212
rect 2159 184 2197 212
rect 2225 184 2263 212
rect 2291 184 2329 212
rect 2357 184 2395 212
rect 2423 184 2461 212
rect 2489 184 2527 212
rect 2555 184 2593 212
rect 2621 184 2659 212
rect 2687 184 2725 212
rect 2753 184 2791 212
rect 2819 184 2857 212
rect 2885 184 2923 212
rect 2951 184 2989 212
rect 3017 184 3055 212
rect 3083 184 3121 212
rect 3149 184 3187 212
rect 3215 184 3253 212
rect 3281 184 3319 212
rect 3347 184 3385 212
rect 3413 184 3451 212
rect 3479 184 3517 212
rect 3545 184 3583 212
rect 3611 184 3649 212
rect 3677 184 3715 212
rect 3743 184 3781 212
rect 3809 184 3847 212
rect 3875 184 3883 212
rect -3883 146 3883 184
rect -3883 118 -3875 146
rect -3847 118 -3809 146
rect -3781 118 -3743 146
rect -3715 118 -3677 146
rect -3649 118 -3611 146
rect -3583 118 -3545 146
rect -3517 118 -3479 146
rect -3451 118 -3413 146
rect -3385 118 -3347 146
rect -3319 118 -3281 146
rect -3253 118 -3215 146
rect -3187 118 -3149 146
rect -3121 118 -3083 146
rect -3055 118 -3017 146
rect -2989 118 -2951 146
rect -2923 118 -2885 146
rect -2857 118 -2819 146
rect -2791 118 -2753 146
rect -2725 118 -2687 146
rect -2659 118 -2621 146
rect -2593 118 -2555 146
rect -2527 118 -2489 146
rect -2461 118 -2423 146
rect -2395 118 -2357 146
rect -2329 118 -2291 146
rect -2263 118 -2225 146
rect -2197 118 -2159 146
rect -2131 118 -2093 146
rect -2065 118 -2027 146
rect -1999 118 -1961 146
rect -1933 118 -1895 146
rect -1867 118 -1829 146
rect -1801 118 -1763 146
rect -1735 118 -1697 146
rect -1669 118 -1631 146
rect -1603 118 -1565 146
rect -1537 118 -1499 146
rect -1471 118 -1433 146
rect -1405 118 -1367 146
rect -1339 118 -1301 146
rect -1273 118 -1235 146
rect -1207 118 -1169 146
rect -1141 118 -1103 146
rect -1075 118 -1037 146
rect -1009 118 -971 146
rect -943 118 -905 146
rect -877 118 -839 146
rect -811 118 -773 146
rect -745 118 -707 146
rect -679 118 -641 146
rect -613 118 -575 146
rect -547 118 -509 146
rect -481 118 -443 146
rect -415 118 -377 146
rect -349 118 -311 146
rect -283 118 -245 146
rect -217 118 -179 146
rect -151 118 -113 146
rect -85 118 -47 146
rect -19 118 19 146
rect 47 118 85 146
rect 113 118 151 146
rect 179 118 217 146
rect 245 118 283 146
rect 311 118 349 146
rect 377 118 415 146
rect 443 118 481 146
rect 509 118 547 146
rect 575 118 613 146
rect 641 118 679 146
rect 707 118 745 146
rect 773 118 811 146
rect 839 118 877 146
rect 905 118 943 146
rect 971 118 1009 146
rect 1037 118 1075 146
rect 1103 118 1141 146
rect 1169 118 1207 146
rect 1235 118 1273 146
rect 1301 118 1339 146
rect 1367 118 1405 146
rect 1433 118 1471 146
rect 1499 118 1537 146
rect 1565 118 1603 146
rect 1631 118 1669 146
rect 1697 118 1735 146
rect 1763 118 1801 146
rect 1829 118 1867 146
rect 1895 118 1933 146
rect 1961 118 1999 146
rect 2027 118 2065 146
rect 2093 118 2131 146
rect 2159 118 2197 146
rect 2225 118 2263 146
rect 2291 118 2329 146
rect 2357 118 2395 146
rect 2423 118 2461 146
rect 2489 118 2527 146
rect 2555 118 2593 146
rect 2621 118 2659 146
rect 2687 118 2725 146
rect 2753 118 2791 146
rect 2819 118 2857 146
rect 2885 118 2923 146
rect 2951 118 2989 146
rect 3017 118 3055 146
rect 3083 118 3121 146
rect 3149 118 3187 146
rect 3215 118 3253 146
rect 3281 118 3319 146
rect 3347 118 3385 146
rect 3413 118 3451 146
rect 3479 118 3517 146
rect 3545 118 3583 146
rect 3611 118 3649 146
rect 3677 118 3715 146
rect 3743 118 3781 146
rect 3809 118 3847 146
rect 3875 118 3883 146
rect -3883 80 3883 118
rect -3883 52 -3875 80
rect -3847 52 -3809 80
rect -3781 52 -3743 80
rect -3715 52 -3677 80
rect -3649 52 -3611 80
rect -3583 52 -3545 80
rect -3517 52 -3479 80
rect -3451 52 -3413 80
rect -3385 52 -3347 80
rect -3319 52 -3281 80
rect -3253 52 -3215 80
rect -3187 52 -3149 80
rect -3121 52 -3083 80
rect -3055 52 -3017 80
rect -2989 52 -2951 80
rect -2923 52 -2885 80
rect -2857 52 -2819 80
rect -2791 52 -2753 80
rect -2725 52 -2687 80
rect -2659 52 -2621 80
rect -2593 52 -2555 80
rect -2527 52 -2489 80
rect -2461 52 -2423 80
rect -2395 52 -2357 80
rect -2329 52 -2291 80
rect -2263 52 -2225 80
rect -2197 52 -2159 80
rect -2131 52 -2093 80
rect -2065 52 -2027 80
rect -1999 52 -1961 80
rect -1933 52 -1895 80
rect -1867 52 -1829 80
rect -1801 52 -1763 80
rect -1735 52 -1697 80
rect -1669 52 -1631 80
rect -1603 52 -1565 80
rect -1537 52 -1499 80
rect -1471 52 -1433 80
rect -1405 52 -1367 80
rect -1339 52 -1301 80
rect -1273 52 -1235 80
rect -1207 52 -1169 80
rect -1141 52 -1103 80
rect -1075 52 -1037 80
rect -1009 52 -971 80
rect -943 52 -905 80
rect -877 52 -839 80
rect -811 52 -773 80
rect -745 52 -707 80
rect -679 52 -641 80
rect -613 52 -575 80
rect -547 52 -509 80
rect -481 52 -443 80
rect -415 52 -377 80
rect -349 52 -311 80
rect -283 52 -245 80
rect -217 52 -179 80
rect -151 52 -113 80
rect -85 52 -47 80
rect -19 52 19 80
rect 47 52 85 80
rect 113 52 151 80
rect 179 52 217 80
rect 245 52 283 80
rect 311 52 349 80
rect 377 52 415 80
rect 443 52 481 80
rect 509 52 547 80
rect 575 52 613 80
rect 641 52 679 80
rect 707 52 745 80
rect 773 52 811 80
rect 839 52 877 80
rect 905 52 943 80
rect 971 52 1009 80
rect 1037 52 1075 80
rect 1103 52 1141 80
rect 1169 52 1207 80
rect 1235 52 1273 80
rect 1301 52 1339 80
rect 1367 52 1405 80
rect 1433 52 1471 80
rect 1499 52 1537 80
rect 1565 52 1603 80
rect 1631 52 1669 80
rect 1697 52 1735 80
rect 1763 52 1801 80
rect 1829 52 1867 80
rect 1895 52 1933 80
rect 1961 52 1999 80
rect 2027 52 2065 80
rect 2093 52 2131 80
rect 2159 52 2197 80
rect 2225 52 2263 80
rect 2291 52 2329 80
rect 2357 52 2395 80
rect 2423 52 2461 80
rect 2489 52 2527 80
rect 2555 52 2593 80
rect 2621 52 2659 80
rect 2687 52 2725 80
rect 2753 52 2791 80
rect 2819 52 2857 80
rect 2885 52 2923 80
rect 2951 52 2989 80
rect 3017 52 3055 80
rect 3083 52 3121 80
rect 3149 52 3187 80
rect 3215 52 3253 80
rect 3281 52 3319 80
rect 3347 52 3385 80
rect 3413 52 3451 80
rect 3479 52 3517 80
rect 3545 52 3583 80
rect 3611 52 3649 80
rect 3677 52 3715 80
rect 3743 52 3781 80
rect 3809 52 3847 80
rect 3875 52 3883 80
rect -3883 14 3883 52
rect -3883 -14 -3875 14
rect -3847 -14 -3809 14
rect -3781 -14 -3743 14
rect -3715 -14 -3677 14
rect -3649 -14 -3611 14
rect -3583 -14 -3545 14
rect -3517 -14 -3479 14
rect -3451 -14 -3413 14
rect -3385 -14 -3347 14
rect -3319 -14 -3281 14
rect -3253 -14 -3215 14
rect -3187 -14 -3149 14
rect -3121 -14 -3083 14
rect -3055 -14 -3017 14
rect -2989 -14 -2951 14
rect -2923 -14 -2885 14
rect -2857 -14 -2819 14
rect -2791 -14 -2753 14
rect -2725 -14 -2687 14
rect -2659 -14 -2621 14
rect -2593 -14 -2555 14
rect -2527 -14 -2489 14
rect -2461 -14 -2423 14
rect -2395 -14 -2357 14
rect -2329 -14 -2291 14
rect -2263 -14 -2225 14
rect -2197 -14 -2159 14
rect -2131 -14 -2093 14
rect -2065 -14 -2027 14
rect -1999 -14 -1961 14
rect -1933 -14 -1895 14
rect -1867 -14 -1829 14
rect -1801 -14 -1763 14
rect -1735 -14 -1697 14
rect -1669 -14 -1631 14
rect -1603 -14 -1565 14
rect -1537 -14 -1499 14
rect -1471 -14 -1433 14
rect -1405 -14 -1367 14
rect -1339 -14 -1301 14
rect -1273 -14 -1235 14
rect -1207 -14 -1169 14
rect -1141 -14 -1103 14
rect -1075 -14 -1037 14
rect -1009 -14 -971 14
rect -943 -14 -905 14
rect -877 -14 -839 14
rect -811 -14 -773 14
rect -745 -14 -707 14
rect -679 -14 -641 14
rect -613 -14 -575 14
rect -547 -14 -509 14
rect -481 -14 -443 14
rect -415 -14 -377 14
rect -349 -14 -311 14
rect -283 -14 -245 14
rect -217 -14 -179 14
rect -151 -14 -113 14
rect -85 -14 -47 14
rect -19 -14 19 14
rect 47 -14 85 14
rect 113 -14 151 14
rect 179 -14 217 14
rect 245 -14 283 14
rect 311 -14 349 14
rect 377 -14 415 14
rect 443 -14 481 14
rect 509 -14 547 14
rect 575 -14 613 14
rect 641 -14 679 14
rect 707 -14 745 14
rect 773 -14 811 14
rect 839 -14 877 14
rect 905 -14 943 14
rect 971 -14 1009 14
rect 1037 -14 1075 14
rect 1103 -14 1141 14
rect 1169 -14 1207 14
rect 1235 -14 1273 14
rect 1301 -14 1339 14
rect 1367 -14 1405 14
rect 1433 -14 1471 14
rect 1499 -14 1537 14
rect 1565 -14 1603 14
rect 1631 -14 1669 14
rect 1697 -14 1735 14
rect 1763 -14 1801 14
rect 1829 -14 1867 14
rect 1895 -14 1933 14
rect 1961 -14 1999 14
rect 2027 -14 2065 14
rect 2093 -14 2131 14
rect 2159 -14 2197 14
rect 2225 -14 2263 14
rect 2291 -14 2329 14
rect 2357 -14 2395 14
rect 2423 -14 2461 14
rect 2489 -14 2527 14
rect 2555 -14 2593 14
rect 2621 -14 2659 14
rect 2687 -14 2725 14
rect 2753 -14 2791 14
rect 2819 -14 2857 14
rect 2885 -14 2923 14
rect 2951 -14 2989 14
rect 3017 -14 3055 14
rect 3083 -14 3121 14
rect 3149 -14 3187 14
rect 3215 -14 3253 14
rect 3281 -14 3319 14
rect 3347 -14 3385 14
rect 3413 -14 3451 14
rect 3479 -14 3517 14
rect 3545 -14 3583 14
rect 3611 -14 3649 14
rect 3677 -14 3715 14
rect 3743 -14 3781 14
rect 3809 -14 3847 14
rect 3875 -14 3883 14
rect -3883 -52 3883 -14
rect -3883 -80 -3875 -52
rect -3847 -80 -3809 -52
rect -3781 -80 -3743 -52
rect -3715 -80 -3677 -52
rect -3649 -80 -3611 -52
rect -3583 -80 -3545 -52
rect -3517 -80 -3479 -52
rect -3451 -80 -3413 -52
rect -3385 -80 -3347 -52
rect -3319 -80 -3281 -52
rect -3253 -80 -3215 -52
rect -3187 -80 -3149 -52
rect -3121 -80 -3083 -52
rect -3055 -80 -3017 -52
rect -2989 -80 -2951 -52
rect -2923 -80 -2885 -52
rect -2857 -80 -2819 -52
rect -2791 -80 -2753 -52
rect -2725 -80 -2687 -52
rect -2659 -80 -2621 -52
rect -2593 -80 -2555 -52
rect -2527 -80 -2489 -52
rect -2461 -80 -2423 -52
rect -2395 -80 -2357 -52
rect -2329 -80 -2291 -52
rect -2263 -80 -2225 -52
rect -2197 -80 -2159 -52
rect -2131 -80 -2093 -52
rect -2065 -80 -2027 -52
rect -1999 -80 -1961 -52
rect -1933 -80 -1895 -52
rect -1867 -80 -1829 -52
rect -1801 -80 -1763 -52
rect -1735 -80 -1697 -52
rect -1669 -80 -1631 -52
rect -1603 -80 -1565 -52
rect -1537 -80 -1499 -52
rect -1471 -80 -1433 -52
rect -1405 -80 -1367 -52
rect -1339 -80 -1301 -52
rect -1273 -80 -1235 -52
rect -1207 -80 -1169 -52
rect -1141 -80 -1103 -52
rect -1075 -80 -1037 -52
rect -1009 -80 -971 -52
rect -943 -80 -905 -52
rect -877 -80 -839 -52
rect -811 -80 -773 -52
rect -745 -80 -707 -52
rect -679 -80 -641 -52
rect -613 -80 -575 -52
rect -547 -80 -509 -52
rect -481 -80 -443 -52
rect -415 -80 -377 -52
rect -349 -80 -311 -52
rect -283 -80 -245 -52
rect -217 -80 -179 -52
rect -151 -80 -113 -52
rect -85 -80 -47 -52
rect -19 -80 19 -52
rect 47 -80 85 -52
rect 113 -80 151 -52
rect 179 -80 217 -52
rect 245 -80 283 -52
rect 311 -80 349 -52
rect 377 -80 415 -52
rect 443 -80 481 -52
rect 509 -80 547 -52
rect 575 -80 613 -52
rect 641 -80 679 -52
rect 707 -80 745 -52
rect 773 -80 811 -52
rect 839 -80 877 -52
rect 905 -80 943 -52
rect 971 -80 1009 -52
rect 1037 -80 1075 -52
rect 1103 -80 1141 -52
rect 1169 -80 1207 -52
rect 1235 -80 1273 -52
rect 1301 -80 1339 -52
rect 1367 -80 1405 -52
rect 1433 -80 1471 -52
rect 1499 -80 1537 -52
rect 1565 -80 1603 -52
rect 1631 -80 1669 -52
rect 1697 -80 1735 -52
rect 1763 -80 1801 -52
rect 1829 -80 1867 -52
rect 1895 -80 1933 -52
rect 1961 -80 1999 -52
rect 2027 -80 2065 -52
rect 2093 -80 2131 -52
rect 2159 -80 2197 -52
rect 2225 -80 2263 -52
rect 2291 -80 2329 -52
rect 2357 -80 2395 -52
rect 2423 -80 2461 -52
rect 2489 -80 2527 -52
rect 2555 -80 2593 -52
rect 2621 -80 2659 -52
rect 2687 -80 2725 -52
rect 2753 -80 2791 -52
rect 2819 -80 2857 -52
rect 2885 -80 2923 -52
rect 2951 -80 2989 -52
rect 3017 -80 3055 -52
rect 3083 -80 3121 -52
rect 3149 -80 3187 -52
rect 3215 -80 3253 -52
rect 3281 -80 3319 -52
rect 3347 -80 3385 -52
rect 3413 -80 3451 -52
rect 3479 -80 3517 -52
rect 3545 -80 3583 -52
rect 3611 -80 3649 -52
rect 3677 -80 3715 -52
rect 3743 -80 3781 -52
rect 3809 -80 3847 -52
rect 3875 -80 3883 -52
rect -3883 -118 3883 -80
rect -3883 -146 -3875 -118
rect -3847 -146 -3809 -118
rect -3781 -146 -3743 -118
rect -3715 -146 -3677 -118
rect -3649 -146 -3611 -118
rect -3583 -146 -3545 -118
rect -3517 -146 -3479 -118
rect -3451 -146 -3413 -118
rect -3385 -146 -3347 -118
rect -3319 -146 -3281 -118
rect -3253 -146 -3215 -118
rect -3187 -146 -3149 -118
rect -3121 -146 -3083 -118
rect -3055 -146 -3017 -118
rect -2989 -146 -2951 -118
rect -2923 -146 -2885 -118
rect -2857 -146 -2819 -118
rect -2791 -146 -2753 -118
rect -2725 -146 -2687 -118
rect -2659 -146 -2621 -118
rect -2593 -146 -2555 -118
rect -2527 -146 -2489 -118
rect -2461 -146 -2423 -118
rect -2395 -146 -2357 -118
rect -2329 -146 -2291 -118
rect -2263 -146 -2225 -118
rect -2197 -146 -2159 -118
rect -2131 -146 -2093 -118
rect -2065 -146 -2027 -118
rect -1999 -146 -1961 -118
rect -1933 -146 -1895 -118
rect -1867 -146 -1829 -118
rect -1801 -146 -1763 -118
rect -1735 -146 -1697 -118
rect -1669 -146 -1631 -118
rect -1603 -146 -1565 -118
rect -1537 -146 -1499 -118
rect -1471 -146 -1433 -118
rect -1405 -146 -1367 -118
rect -1339 -146 -1301 -118
rect -1273 -146 -1235 -118
rect -1207 -146 -1169 -118
rect -1141 -146 -1103 -118
rect -1075 -146 -1037 -118
rect -1009 -146 -971 -118
rect -943 -146 -905 -118
rect -877 -146 -839 -118
rect -811 -146 -773 -118
rect -745 -146 -707 -118
rect -679 -146 -641 -118
rect -613 -146 -575 -118
rect -547 -146 -509 -118
rect -481 -146 -443 -118
rect -415 -146 -377 -118
rect -349 -146 -311 -118
rect -283 -146 -245 -118
rect -217 -146 -179 -118
rect -151 -146 -113 -118
rect -85 -146 -47 -118
rect -19 -146 19 -118
rect 47 -146 85 -118
rect 113 -146 151 -118
rect 179 -146 217 -118
rect 245 -146 283 -118
rect 311 -146 349 -118
rect 377 -146 415 -118
rect 443 -146 481 -118
rect 509 -146 547 -118
rect 575 -146 613 -118
rect 641 -146 679 -118
rect 707 -146 745 -118
rect 773 -146 811 -118
rect 839 -146 877 -118
rect 905 -146 943 -118
rect 971 -146 1009 -118
rect 1037 -146 1075 -118
rect 1103 -146 1141 -118
rect 1169 -146 1207 -118
rect 1235 -146 1273 -118
rect 1301 -146 1339 -118
rect 1367 -146 1405 -118
rect 1433 -146 1471 -118
rect 1499 -146 1537 -118
rect 1565 -146 1603 -118
rect 1631 -146 1669 -118
rect 1697 -146 1735 -118
rect 1763 -146 1801 -118
rect 1829 -146 1867 -118
rect 1895 -146 1933 -118
rect 1961 -146 1999 -118
rect 2027 -146 2065 -118
rect 2093 -146 2131 -118
rect 2159 -146 2197 -118
rect 2225 -146 2263 -118
rect 2291 -146 2329 -118
rect 2357 -146 2395 -118
rect 2423 -146 2461 -118
rect 2489 -146 2527 -118
rect 2555 -146 2593 -118
rect 2621 -146 2659 -118
rect 2687 -146 2725 -118
rect 2753 -146 2791 -118
rect 2819 -146 2857 -118
rect 2885 -146 2923 -118
rect 2951 -146 2989 -118
rect 3017 -146 3055 -118
rect 3083 -146 3121 -118
rect 3149 -146 3187 -118
rect 3215 -146 3253 -118
rect 3281 -146 3319 -118
rect 3347 -146 3385 -118
rect 3413 -146 3451 -118
rect 3479 -146 3517 -118
rect 3545 -146 3583 -118
rect 3611 -146 3649 -118
rect 3677 -146 3715 -118
rect 3743 -146 3781 -118
rect 3809 -146 3847 -118
rect 3875 -146 3883 -118
rect -3883 -184 3883 -146
rect -3883 -212 -3875 -184
rect -3847 -212 -3809 -184
rect -3781 -212 -3743 -184
rect -3715 -212 -3677 -184
rect -3649 -212 -3611 -184
rect -3583 -212 -3545 -184
rect -3517 -212 -3479 -184
rect -3451 -212 -3413 -184
rect -3385 -212 -3347 -184
rect -3319 -212 -3281 -184
rect -3253 -212 -3215 -184
rect -3187 -212 -3149 -184
rect -3121 -212 -3083 -184
rect -3055 -212 -3017 -184
rect -2989 -212 -2951 -184
rect -2923 -212 -2885 -184
rect -2857 -212 -2819 -184
rect -2791 -212 -2753 -184
rect -2725 -212 -2687 -184
rect -2659 -212 -2621 -184
rect -2593 -212 -2555 -184
rect -2527 -212 -2489 -184
rect -2461 -212 -2423 -184
rect -2395 -212 -2357 -184
rect -2329 -212 -2291 -184
rect -2263 -212 -2225 -184
rect -2197 -212 -2159 -184
rect -2131 -212 -2093 -184
rect -2065 -212 -2027 -184
rect -1999 -212 -1961 -184
rect -1933 -212 -1895 -184
rect -1867 -212 -1829 -184
rect -1801 -212 -1763 -184
rect -1735 -212 -1697 -184
rect -1669 -212 -1631 -184
rect -1603 -212 -1565 -184
rect -1537 -212 -1499 -184
rect -1471 -212 -1433 -184
rect -1405 -212 -1367 -184
rect -1339 -212 -1301 -184
rect -1273 -212 -1235 -184
rect -1207 -212 -1169 -184
rect -1141 -212 -1103 -184
rect -1075 -212 -1037 -184
rect -1009 -212 -971 -184
rect -943 -212 -905 -184
rect -877 -212 -839 -184
rect -811 -212 -773 -184
rect -745 -212 -707 -184
rect -679 -212 -641 -184
rect -613 -212 -575 -184
rect -547 -212 -509 -184
rect -481 -212 -443 -184
rect -415 -212 -377 -184
rect -349 -212 -311 -184
rect -283 -212 -245 -184
rect -217 -212 -179 -184
rect -151 -212 -113 -184
rect -85 -212 -47 -184
rect -19 -212 19 -184
rect 47 -212 85 -184
rect 113 -212 151 -184
rect 179 -212 217 -184
rect 245 -212 283 -184
rect 311 -212 349 -184
rect 377 -212 415 -184
rect 443 -212 481 -184
rect 509 -212 547 -184
rect 575 -212 613 -184
rect 641 -212 679 -184
rect 707 -212 745 -184
rect 773 -212 811 -184
rect 839 -212 877 -184
rect 905 -212 943 -184
rect 971 -212 1009 -184
rect 1037 -212 1075 -184
rect 1103 -212 1141 -184
rect 1169 -212 1207 -184
rect 1235 -212 1273 -184
rect 1301 -212 1339 -184
rect 1367 -212 1405 -184
rect 1433 -212 1471 -184
rect 1499 -212 1537 -184
rect 1565 -212 1603 -184
rect 1631 -212 1669 -184
rect 1697 -212 1735 -184
rect 1763 -212 1801 -184
rect 1829 -212 1867 -184
rect 1895 -212 1933 -184
rect 1961 -212 1999 -184
rect 2027 -212 2065 -184
rect 2093 -212 2131 -184
rect 2159 -212 2197 -184
rect 2225 -212 2263 -184
rect 2291 -212 2329 -184
rect 2357 -212 2395 -184
rect 2423 -212 2461 -184
rect 2489 -212 2527 -184
rect 2555 -212 2593 -184
rect 2621 -212 2659 -184
rect 2687 -212 2725 -184
rect 2753 -212 2791 -184
rect 2819 -212 2857 -184
rect 2885 -212 2923 -184
rect 2951 -212 2989 -184
rect 3017 -212 3055 -184
rect 3083 -212 3121 -184
rect 3149 -212 3187 -184
rect 3215 -212 3253 -184
rect 3281 -212 3319 -184
rect 3347 -212 3385 -184
rect 3413 -212 3451 -184
rect 3479 -212 3517 -184
rect 3545 -212 3583 -184
rect 3611 -212 3649 -184
rect 3677 -212 3715 -184
rect 3743 -212 3781 -184
rect 3809 -212 3847 -184
rect 3875 -212 3883 -184
rect -3883 -250 3883 -212
rect -3883 -278 -3875 -250
rect -3847 -278 -3809 -250
rect -3781 -278 -3743 -250
rect -3715 -278 -3677 -250
rect -3649 -278 -3611 -250
rect -3583 -278 -3545 -250
rect -3517 -278 -3479 -250
rect -3451 -278 -3413 -250
rect -3385 -278 -3347 -250
rect -3319 -278 -3281 -250
rect -3253 -278 -3215 -250
rect -3187 -278 -3149 -250
rect -3121 -278 -3083 -250
rect -3055 -278 -3017 -250
rect -2989 -278 -2951 -250
rect -2923 -278 -2885 -250
rect -2857 -278 -2819 -250
rect -2791 -278 -2753 -250
rect -2725 -278 -2687 -250
rect -2659 -278 -2621 -250
rect -2593 -278 -2555 -250
rect -2527 -278 -2489 -250
rect -2461 -278 -2423 -250
rect -2395 -278 -2357 -250
rect -2329 -278 -2291 -250
rect -2263 -278 -2225 -250
rect -2197 -278 -2159 -250
rect -2131 -278 -2093 -250
rect -2065 -278 -2027 -250
rect -1999 -278 -1961 -250
rect -1933 -278 -1895 -250
rect -1867 -278 -1829 -250
rect -1801 -278 -1763 -250
rect -1735 -278 -1697 -250
rect -1669 -278 -1631 -250
rect -1603 -278 -1565 -250
rect -1537 -278 -1499 -250
rect -1471 -278 -1433 -250
rect -1405 -278 -1367 -250
rect -1339 -278 -1301 -250
rect -1273 -278 -1235 -250
rect -1207 -278 -1169 -250
rect -1141 -278 -1103 -250
rect -1075 -278 -1037 -250
rect -1009 -278 -971 -250
rect -943 -278 -905 -250
rect -877 -278 -839 -250
rect -811 -278 -773 -250
rect -745 -278 -707 -250
rect -679 -278 -641 -250
rect -613 -278 -575 -250
rect -547 -278 -509 -250
rect -481 -278 -443 -250
rect -415 -278 -377 -250
rect -349 -278 -311 -250
rect -283 -278 -245 -250
rect -217 -278 -179 -250
rect -151 -278 -113 -250
rect -85 -278 -47 -250
rect -19 -278 19 -250
rect 47 -278 85 -250
rect 113 -278 151 -250
rect 179 -278 217 -250
rect 245 -278 283 -250
rect 311 -278 349 -250
rect 377 -278 415 -250
rect 443 -278 481 -250
rect 509 -278 547 -250
rect 575 -278 613 -250
rect 641 -278 679 -250
rect 707 -278 745 -250
rect 773 -278 811 -250
rect 839 -278 877 -250
rect 905 -278 943 -250
rect 971 -278 1009 -250
rect 1037 -278 1075 -250
rect 1103 -278 1141 -250
rect 1169 -278 1207 -250
rect 1235 -278 1273 -250
rect 1301 -278 1339 -250
rect 1367 -278 1405 -250
rect 1433 -278 1471 -250
rect 1499 -278 1537 -250
rect 1565 -278 1603 -250
rect 1631 -278 1669 -250
rect 1697 -278 1735 -250
rect 1763 -278 1801 -250
rect 1829 -278 1867 -250
rect 1895 -278 1933 -250
rect 1961 -278 1999 -250
rect 2027 -278 2065 -250
rect 2093 -278 2131 -250
rect 2159 -278 2197 -250
rect 2225 -278 2263 -250
rect 2291 -278 2329 -250
rect 2357 -278 2395 -250
rect 2423 -278 2461 -250
rect 2489 -278 2527 -250
rect 2555 -278 2593 -250
rect 2621 -278 2659 -250
rect 2687 -278 2725 -250
rect 2753 -278 2791 -250
rect 2819 -278 2857 -250
rect 2885 -278 2923 -250
rect 2951 -278 2989 -250
rect 3017 -278 3055 -250
rect 3083 -278 3121 -250
rect 3149 -278 3187 -250
rect 3215 -278 3253 -250
rect 3281 -278 3319 -250
rect 3347 -278 3385 -250
rect 3413 -278 3451 -250
rect 3479 -278 3517 -250
rect 3545 -278 3583 -250
rect 3611 -278 3649 -250
rect 3677 -278 3715 -250
rect 3743 -278 3781 -250
rect 3809 -278 3847 -250
rect 3875 -278 3883 -250
rect -3883 -316 3883 -278
rect -3883 -344 -3875 -316
rect -3847 -344 -3809 -316
rect -3781 -344 -3743 -316
rect -3715 -344 -3677 -316
rect -3649 -344 -3611 -316
rect -3583 -344 -3545 -316
rect -3517 -344 -3479 -316
rect -3451 -344 -3413 -316
rect -3385 -344 -3347 -316
rect -3319 -344 -3281 -316
rect -3253 -344 -3215 -316
rect -3187 -344 -3149 -316
rect -3121 -344 -3083 -316
rect -3055 -344 -3017 -316
rect -2989 -344 -2951 -316
rect -2923 -344 -2885 -316
rect -2857 -344 -2819 -316
rect -2791 -344 -2753 -316
rect -2725 -344 -2687 -316
rect -2659 -344 -2621 -316
rect -2593 -344 -2555 -316
rect -2527 -344 -2489 -316
rect -2461 -344 -2423 -316
rect -2395 -344 -2357 -316
rect -2329 -344 -2291 -316
rect -2263 -344 -2225 -316
rect -2197 -344 -2159 -316
rect -2131 -344 -2093 -316
rect -2065 -344 -2027 -316
rect -1999 -344 -1961 -316
rect -1933 -344 -1895 -316
rect -1867 -344 -1829 -316
rect -1801 -344 -1763 -316
rect -1735 -344 -1697 -316
rect -1669 -344 -1631 -316
rect -1603 -344 -1565 -316
rect -1537 -344 -1499 -316
rect -1471 -344 -1433 -316
rect -1405 -344 -1367 -316
rect -1339 -344 -1301 -316
rect -1273 -344 -1235 -316
rect -1207 -344 -1169 -316
rect -1141 -344 -1103 -316
rect -1075 -344 -1037 -316
rect -1009 -344 -971 -316
rect -943 -344 -905 -316
rect -877 -344 -839 -316
rect -811 -344 -773 -316
rect -745 -344 -707 -316
rect -679 -344 -641 -316
rect -613 -344 -575 -316
rect -547 -344 -509 -316
rect -481 -344 -443 -316
rect -415 -344 -377 -316
rect -349 -344 -311 -316
rect -283 -344 -245 -316
rect -217 -344 -179 -316
rect -151 -344 -113 -316
rect -85 -344 -47 -316
rect -19 -344 19 -316
rect 47 -344 85 -316
rect 113 -344 151 -316
rect 179 -344 217 -316
rect 245 -344 283 -316
rect 311 -344 349 -316
rect 377 -344 415 -316
rect 443 -344 481 -316
rect 509 -344 547 -316
rect 575 -344 613 -316
rect 641 -344 679 -316
rect 707 -344 745 -316
rect 773 -344 811 -316
rect 839 -344 877 -316
rect 905 -344 943 -316
rect 971 -344 1009 -316
rect 1037 -344 1075 -316
rect 1103 -344 1141 -316
rect 1169 -344 1207 -316
rect 1235 -344 1273 -316
rect 1301 -344 1339 -316
rect 1367 -344 1405 -316
rect 1433 -344 1471 -316
rect 1499 -344 1537 -316
rect 1565 -344 1603 -316
rect 1631 -344 1669 -316
rect 1697 -344 1735 -316
rect 1763 -344 1801 -316
rect 1829 -344 1867 -316
rect 1895 -344 1933 -316
rect 1961 -344 1999 -316
rect 2027 -344 2065 -316
rect 2093 -344 2131 -316
rect 2159 -344 2197 -316
rect 2225 -344 2263 -316
rect 2291 -344 2329 -316
rect 2357 -344 2395 -316
rect 2423 -344 2461 -316
rect 2489 -344 2527 -316
rect 2555 -344 2593 -316
rect 2621 -344 2659 -316
rect 2687 -344 2725 -316
rect 2753 -344 2791 -316
rect 2819 -344 2857 -316
rect 2885 -344 2923 -316
rect 2951 -344 2989 -316
rect 3017 -344 3055 -316
rect 3083 -344 3121 -316
rect 3149 -344 3187 -316
rect 3215 -344 3253 -316
rect 3281 -344 3319 -316
rect 3347 -344 3385 -316
rect 3413 -344 3451 -316
rect 3479 -344 3517 -316
rect 3545 -344 3583 -316
rect 3611 -344 3649 -316
rect 3677 -344 3715 -316
rect 3743 -344 3781 -316
rect 3809 -344 3847 -316
rect 3875 -344 3883 -316
rect -3883 -382 3883 -344
rect -3883 -410 -3875 -382
rect -3847 -410 -3809 -382
rect -3781 -410 -3743 -382
rect -3715 -410 -3677 -382
rect -3649 -410 -3611 -382
rect -3583 -410 -3545 -382
rect -3517 -410 -3479 -382
rect -3451 -410 -3413 -382
rect -3385 -410 -3347 -382
rect -3319 -410 -3281 -382
rect -3253 -410 -3215 -382
rect -3187 -410 -3149 -382
rect -3121 -410 -3083 -382
rect -3055 -410 -3017 -382
rect -2989 -410 -2951 -382
rect -2923 -410 -2885 -382
rect -2857 -410 -2819 -382
rect -2791 -410 -2753 -382
rect -2725 -410 -2687 -382
rect -2659 -410 -2621 -382
rect -2593 -410 -2555 -382
rect -2527 -410 -2489 -382
rect -2461 -410 -2423 -382
rect -2395 -410 -2357 -382
rect -2329 -410 -2291 -382
rect -2263 -410 -2225 -382
rect -2197 -410 -2159 -382
rect -2131 -410 -2093 -382
rect -2065 -410 -2027 -382
rect -1999 -410 -1961 -382
rect -1933 -410 -1895 -382
rect -1867 -410 -1829 -382
rect -1801 -410 -1763 -382
rect -1735 -410 -1697 -382
rect -1669 -410 -1631 -382
rect -1603 -410 -1565 -382
rect -1537 -410 -1499 -382
rect -1471 -410 -1433 -382
rect -1405 -410 -1367 -382
rect -1339 -410 -1301 -382
rect -1273 -410 -1235 -382
rect -1207 -410 -1169 -382
rect -1141 -410 -1103 -382
rect -1075 -410 -1037 -382
rect -1009 -410 -971 -382
rect -943 -410 -905 -382
rect -877 -410 -839 -382
rect -811 -410 -773 -382
rect -745 -410 -707 -382
rect -679 -410 -641 -382
rect -613 -410 -575 -382
rect -547 -410 -509 -382
rect -481 -410 -443 -382
rect -415 -410 -377 -382
rect -349 -410 -311 -382
rect -283 -410 -245 -382
rect -217 -410 -179 -382
rect -151 -410 -113 -382
rect -85 -410 -47 -382
rect -19 -410 19 -382
rect 47 -410 85 -382
rect 113 -410 151 -382
rect 179 -410 217 -382
rect 245 -410 283 -382
rect 311 -410 349 -382
rect 377 -410 415 -382
rect 443 -410 481 -382
rect 509 -410 547 -382
rect 575 -410 613 -382
rect 641 -410 679 -382
rect 707 -410 745 -382
rect 773 -410 811 -382
rect 839 -410 877 -382
rect 905 -410 943 -382
rect 971 -410 1009 -382
rect 1037 -410 1075 -382
rect 1103 -410 1141 -382
rect 1169 -410 1207 -382
rect 1235 -410 1273 -382
rect 1301 -410 1339 -382
rect 1367 -410 1405 -382
rect 1433 -410 1471 -382
rect 1499 -410 1537 -382
rect 1565 -410 1603 -382
rect 1631 -410 1669 -382
rect 1697 -410 1735 -382
rect 1763 -410 1801 -382
rect 1829 -410 1867 -382
rect 1895 -410 1933 -382
rect 1961 -410 1999 -382
rect 2027 -410 2065 -382
rect 2093 -410 2131 -382
rect 2159 -410 2197 -382
rect 2225 -410 2263 -382
rect 2291 -410 2329 -382
rect 2357 -410 2395 -382
rect 2423 -410 2461 -382
rect 2489 -410 2527 -382
rect 2555 -410 2593 -382
rect 2621 -410 2659 -382
rect 2687 -410 2725 -382
rect 2753 -410 2791 -382
rect 2819 -410 2857 -382
rect 2885 -410 2923 -382
rect 2951 -410 2989 -382
rect 3017 -410 3055 -382
rect 3083 -410 3121 -382
rect 3149 -410 3187 -382
rect 3215 -410 3253 -382
rect 3281 -410 3319 -382
rect 3347 -410 3385 -382
rect 3413 -410 3451 -382
rect 3479 -410 3517 -382
rect 3545 -410 3583 -382
rect 3611 -410 3649 -382
rect 3677 -410 3715 -382
rect 3743 -410 3781 -382
rect 3809 -410 3847 -382
rect 3875 -410 3883 -382
rect -3883 -448 3883 -410
rect -3883 -476 -3875 -448
rect -3847 -476 -3809 -448
rect -3781 -476 -3743 -448
rect -3715 -476 -3677 -448
rect -3649 -476 -3611 -448
rect -3583 -476 -3545 -448
rect -3517 -476 -3479 -448
rect -3451 -476 -3413 -448
rect -3385 -476 -3347 -448
rect -3319 -476 -3281 -448
rect -3253 -476 -3215 -448
rect -3187 -476 -3149 -448
rect -3121 -476 -3083 -448
rect -3055 -476 -3017 -448
rect -2989 -476 -2951 -448
rect -2923 -476 -2885 -448
rect -2857 -476 -2819 -448
rect -2791 -476 -2753 -448
rect -2725 -476 -2687 -448
rect -2659 -476 -2621 -448
rect -2593 -476 -2555 -448
rect -2527 -476 -2489 -448
rect -2461 -476 -2423 -448
rect -2395 -476 -2357 -448
rect -2329 -476 -2291 -448
rect -2263 -476 -2225 -448
rect -2197 -476 -2159 -448
rect -2131 -476 -2093 -448
rect -2065 -476 -2027 -448
rect -1999 -476 -1961 -448
rect -1933 -476 -1895 -448
rect -1867 -476 -1829 -448
rect -1801 -476 -1763 -448
rect -1735 -476 -1697 -448
rect -1669 -476 -1631 -448
rect -1603 -476 -1565 -448
rect -1537 -476 -1499 -448
rect -1471 -476 -1433 -448
rect -1405 -476 -1367 -448
rect -1339 -476 -1301 -448
rect -1273 -476 -1235 -448
rect -1207 -476 -1169 -448
rect -1141 -476 -1103 -448
rect -1075 -476 -1037 -448
rect -1009 -476 -971 -448
rect -943 -476 -905 -448
rect -877 -476 -839 -448
rect -811 -476 -773 -448
rect -745 -476 -707 -448
rect -679 -476 -641 -448
rect -613 -476 -575 -448
rect -547 -476 -509 -448
rect -481 -476 -443 -448
rect -415 -476 -377 -448
rect -349 -476 -311 -448
rect -283 -476 -245 -448
rect -217 -476 -179 -448
rect -151 -476 -113 -448
rect -85 -476 -47 -448
rect -19 -476 19 -448
rect 47 -476 85 -448
rect 113 -476 151 -448
rect 179 -476 217 -448
rect 245 -476 283 -448
rect 311 -476 349 -448
rect 377 -476 415 -448
rect 443 -476 481 -448
rect 509 -476 547 -448
rect 575 -476 613 -448
rect 641 -476 679 -448
rect 707 -476 745 -448
rect 773 -476 811 -448
rect 839 -476 877 -448
rect 905 -476 943 -448
rect 971 -476 1009 -448
rect 1037 -476 1075 -448
rect 1103 -476 1141 -448
rect 1169 -476 1207 -448
rect 1235 -476 1273 -448
rect 1301 -476 1339 -448
rect 1367 -476 1405 -448
rect 1433 -476 1471 -448
rect 1499 -476 1537 -448
rect 1565 -476 1603 -448
rect 1631 -476 1669 -448
rect 1697 -476 1735 -448
rect 1763 -476 1801 -448
rect 1829 -476 1867 -448
rect 1895 -476 1933 -448
rect 1961 -476 1999 -448
rect 2027 -476 2065 -448
rect 2093 -476 2131 -448
rect 2159 -476 2197 -448
rect 2225 -476 2263 -448
rect 2291 -476 2329 -448
rect 2357 -476 2395 -448
rect 2423 -476 2461 -448
rect 2489 -476 2527 -448
rect 2555 -476 2593 -448
rect 2621 -476 2659 -448
rect 2687 -476 2725 -448
rect 2753 -476 2791 -448
rect 2819 -476 2857 -448
rect 2885 -476 2923 -448
rect 2951 -476 2989 -448
rect 3017 -476 3055 -448
rect 3083 -476 3121 -448
rect 3149 -476 3187 -448
rect 3215 -476 3253 -448
rect 3281 -476 3319 -448
rect 3347 -476 3385 -448
rect 3413 -476 3451 -448
rect 3479 -476 3517 -448
rect 3545 -476 3583 -448
rect 3611 -476 3649 -448
rect 3677 -476 3715 -448
rect 3743 -476 3781 -448
rect 3809 -476 3847 -448
rect 3875 -476 3883 -448
rect -3883 -514 3883 -476
rect -3883 -542 -3875 -514
rect -3847 -542 -3809 -514
rect -3781 -542 -3743 -514
rect -3715 -542 -3677 -514
rect -3649 -542 -3611 -514
rect -3583 -542 -3545 -514
rect -3517 -542 -3479 -514
rect -3451 -542 -3413 -514
rect -3385 -542 -3347 -514
rect -3319 -542 -3281 -514
rect -3253 -542 -3215 -514
rect -3187 -542 -3149 -514
rect -3121 -542 -3083 -514
rect -3055 -542 -3017 -514
rect -2989 -542 -2951 -514
rect -2923 -542 -2885 -514
rect -2857 -542 -2819 -514
rect -2791 -542 -2753 -514
rect -2725 -542 -2687 -514
rect -2659 -542 -2621 -514
rect -2593 -542 -2555 -514
rect -2527 -542 -2489 -514
rect -2461 -542 -2423 -514
rect -2395 -542 -2357 -514
rect -2329 -542 -2291 -514
rect -2263 -542 -2225 -514
rect -2197 -542 -2159 -514
rect -2131 -542 -2093 -514
rect -2065 -542 -2027 -514
rect -1999 -542 -1961 -514
rect -1933 -542 -1895 -514
rect -1867 -542 -1829 -514
rect -1801 -542 -1763 -514
rect -1735 -542 -1697 -514
rect -1669 -542 -1631 -514
rect -1603 -542 -1565 -514
rect -1537 -542 -1499 -514
rect -1471 -542 -1433 -514
rect -1405 -542 -1367 -514
rect -1339 -542 -1301 -514
rect -1273 -542 -1235 -514
rect -1207 -542 -1169 -514
rect -1141 -542 -1103 -514
rect -1075 -542 -1037 -514
rect -1009 -542 -971 -514
rect -943 -542 -905 -514
rect -877 -542 -839 -514
rect -811 -542 -773 -514
rect -745 -542 -707 -514
rect -679 -542 -641 -514
rect -613 -542 -575 -514
rect -547 -542 -509 -514
rect -481 -542 -443 -514
rect -415 -542 -377 -514
rect -349 -542 -311 -514
rect -283 -542 -245 -514
rect -217 -542 -179 -514
rect -151 -542 -113 -514
rect -85 -542 -47 -514
rect -19 -542 19 -514
rect 47 -542 85 -514
rect 113 -542 151 -514
rect 179 -542 217 -514
rect 245 -542 283 -514
rect 311 -542 349 -514
rect 377 -542 415 -514
rect 443 -542 481 -514
rect 509 -542 547 -514
rect 575 -542 613 -514
rect 641 -542 679 -514
rect 707 -542 745 -514
rect 773 -542 811 -514
rect 839 -542 877 -514
rect 905 -542 943 -514
rect 971 -542 1009 -514
rect 1037 -542 1075 -514
rect 1103 -542 1141 -514
rect 1169 -542 1207 -514
rect 1235 -542 1273 -514
rect 1301 -542 1339 -514
rect 1367 -542 1405 -514
rect 1433 -542 1471 -514
rect 1499 -542 1537 -514
rect 1565 -542 1603 -514
rect 1631 -542 1669 -514
rect 1697 -542 1735 -514
rect 1763 -542 1801 -514
rect 1829 -542 1867 -514
rect 1895 -542 1933 -514
rect 1961 -542 1999 -514
rect 2027 -542 2065 -514
rect 2093 -542 2131 -514
rect 2159 -542 2197 -514
rect 2225 -542 2263 -514
rect 2291 -542 2329 -514
rect 2357 -542 2395 -514
rect 2423 -542 2461 -514
rect 2489 -542 2527 -514
rect 2555 -542 2593 -514
rect 2621 -542 2659 -514
rect 2687 -542 2725 -514
rect 2753 -542 2791 -514
rect 2819 -542 2857 -514
rect 2885 -542 2923 -514
rect 2951 -542 2989 -514
rect 3017 -542 3055 -514
rect 3083 -542 3121 -514
rect 3149 -542 3187 -514
rect 3215 -542 3253 -514
rect 3281 -542 3319 -514
rect 3347 -542 3385 -514
rect 3413 -542 3451 -514
rect 3479 -542 3517 -514
rect 3545 -542 3583 -514
rect 3611 -542 3649 -514
rect 3677 -542 3715 -514
rect 3743 -542 3781 -514
rect 3809 -542 3847 -514
rect 3875 -542 3883 -514
rect -3883 -580 3883 -542
rect -3883 -608 -3875 -580
rect -3847 -608 -3809 -580
rect -3781 -608 -3743 -580
rect -3715 -608 -3677 -580
rect -3649 -608 -3611 -580
rect -3583 -608 -3545 -580
rect -3517 -608 -3479 -580
rect -3451 -608 -3413 -580
rect -3385 -608 -3347 -580
rect -3319 -608 -3281 -580
rect -3253 -608 -3215 -580
rect -3187 -608 -3149 -580
rect -3121 -608 -3083 -580
rect -3055 -608 -3017 -580
rect -2989 -608 -2951 -580
rect -2923 -608 -2885 -580
rect -2857 -608 -2819 -580
rect -2791 -608 -2753 -580
rect -2725 -608 -2687 -580
rect -2659 -608 -2621 -580
rect -2593 -608 -2555 -580
rect -2527 -608 -2489 -580
rect -2461 -608 -2423 -580
rect -2395 -608 -2357 -580
rect -2329 -608 -2291 -580
rect -2263 -608 -2225 -580
rect -2197 -608 -2159 -580
rect -2131 -608 -2093 -580
rect -2065 -608 -2027 -580
rect -1999 -608 -1961 -580
rect -1933 -608 -1895 -580
rect -1867 -608 -1829 -580
rect -1801 -608 -1763 -580
rect -1735 -608 -1697 -580
rect -1669 -608 -1631 -580
rect -1603 -608 -1565 -580
rect -1537 -608 -1499 -580
rect -1471 -608 -1433 -580
rect -1405 -608 -1367 -580
rect -1339 -608 -1301 -580
rect -1273 -608 -1235 -580
rect -1207 -608 -1169 -580
rect -1141 -608 -1103 -580
rect -1075 -608 -1037 -580
rect -1009 -608 -971 -580
rect -943 -608 -905 -580
rect -877 -608 -839 -580
rect -811 -608 -773 -580
rect -745 -608 -707 -580
rect -679 -608 -641 -580
rect -613 -608 -575 -580
rect -547 -608 -509 -580
rect -481 -608 -443 -580
rect -415 -608 -377 -580
rect -349 -608 -311 -580
rect -283 -608 -245 -580
rect -217 -608 -179 -580
rect -151 -608 -113 -580
rect -85 -608 -47 -580
rect -19 -608 19 -580
rect 47 -608 85 -580
rect 113 -608 151 -580
rect 179 -608 217 -580
rect 245 -608 283 -580
rect 311 -608 349 -580
rect 377 -608 415 -580
rect 443 -608 481 -580
rect 509 -608 547 -580
rect 575 -608 613 -580
rect 641 -608 679 -580
rect 707 -608 745 -580
rect 773 -608 811 -580
rect 839 -608 877 -580
rect 905 -608 943 -580
rect 971 -608 1009 -580
rect 1037 -608 1075 -580
rect 1103 -608 1141 -580
rect 1169 -608 1207 -580
rect 1235 -608 1273 -580
rect 1301 -608 1339 -580
rect 1367 -608 1405 -580
rect 1433 -608 1471 -580
rect 1499 -608 1537 -580
rect 1565 -608 1603 -580
rect 1631 -608 1669 -580
rect 1697 -608 1735 -580
rect 1763 -608 1801 -580
rect 1829 -608 1867 -580
rect 1895 -608 1933 -580
rect 1961 -608 1999 -580
rect 2027 -608 2065 -580
rect 2093 -608 2131 -580
rect 2159 -608 2197 -580
rect 2225 -608 2263 -580
rect 2291 -608 2329 -580
rect 2357 -608 2395 -580
rect 2423 -608 2461 -580
rect 2489 -608 2527 -580
rect 2555 -608 2593 -580
rect 2621 -608 2659 -580
rect 2687 -608 2725 -580
rect 2753 -608 2791 -580
rect 2819 -608 2857 -580
rect 2885 -608 2923 -580
rect 2951 -608 2989 -580
rect 3017 -608 3055 -580
rect 3083 -608 3121 -580
rect 3149 -608 3187 -580
rect 3215 -608 3253 -580
rect 3281 -608 3319 -580
rect 3347 -608 3385 -580
rect 3413 -608 3451 -580
rect 3479 -608 3517 -580
rect 3545 -608 3583 -580
rect 3611 -608 3649 -580
rect 3677 -608 3715 -580
rect 3743 -608 3781 -580
rect 3809 -608 3847 -580
rect 3875 -608 3883 -580
rect -3883 -646 3883 -608
rect -3883 -674 -3875 -646
rect -3847 -674 -3809 -646
rect -3781 -674 -3743 -646
rect -3715 -674 -3677 -646
rect -3649 -674 -3611 -646
rect -3583 -674 -3545 -646
rect -3517 -674 -3479 -646
rect -3451 -674 -3413 -646
rect -3385 -674 -3347 -646
rect -3319 -674 -3281 -646
rect -3253 -674 -3215 -646
rect -3187 -674 -3149 -646
rect -3121 -674 -3083 -646
rect -3055 -674 -3017 -646
rect -2989 -674 -2951 -646
rect -2923 -674 -2885 -646
rect -2857 -674 -2819 -646
rect -2791 -674 -2753 -646
rect -2725 -674 -2687 -646
rect -2659 -674 -2621 -646
rect -2593 -674 -2555 -646
rect -2527 -674 -2489 -646
rect -2461 -674 -2423 -646
rect -2395 -674 -2357 -646
rect -2329 -674 -2291 -646
rect -2263 -674 -2225 -646
rect -2197 -674 -2159 -646
rect -2131 -674 -2093 -646
rect -2065 -674 -2027 -646
rect -1999 -674 -1961 -646
rect -1933 -674 -1895 -646
rect -1867 -674 -1829 -646
rect -1801 -674 -1763 -646
rect -1735 -674 -1697 -646
rect -1669 -674 -1631 -646
rect -1603 -674 -1565 -646
rect -1537 -674 -1499 -646
rect -1471 -674 -1433 -646
rect -1405 -674 -1367 -646
rect -1339 -674 -1301 -646
rect -1273 -674 -1235 -646
rect -1207 -674 -1169 -646
rect -1141 -674 -1103 -646
rect -1075 -674 -1037 -646
rect -1009 -674 -971 -646
rect -943 -674 -905 -646
rect -877 -674 -839 -646
rect -811 -674 -773 -646
rect -745 -674 -707 -646
rect -679 -674 -641 -646
rect -613 -674 -575 -646
rect -547 -674 -509 -646
rect -481 -674 -443 -646
rect -415 -674 -377 -646
rect -349 -674 -311 -646
rect -283 -674 -245 -646
rect -217 -674 -179 -646
rect -151 -674 -113 -646
rect -85 -674 -47 -646
rect -19 -674 19 -646
rect 47 -674 85 -646
rect 113 -674 151 -646
rect 179 -674 217 -646
rect 245 -674 283 -646
rect 311 -674 349 -646
rect 377 -674 415 -646
rect 443 -674 481 -646
rect 509 -674 547 -646
rect 575 -674 613 -646
rect 641 -674 679 -646
rect 707 -674 745 -646
rect 773 -674 811 -646
rect 839 -674 877 -646
rect 905 -674 943 -646
rect 971 -674 1009 -646
rect 1037 -674 1075 -646
rect 1103 -674 1141 -646
rect 1169 -674 1207 -646
rect 1235 -674 1273 -646
rect 1301 -674 1339 -646
rect 1367 -674 1405 -646
rect 1433 -674 1471 -646
rect 1499 -674 1537 -646
rect 1565 -674 1603 -646
rect 1631 -674 1669 -646
rect 1697 -674 1735 -646
rect 1763 -674 1801 -646
rect 1829 -674 1867 -646
rect 1895 -674 1933 -646
rect 1961 -674 1999 -646
rect 2027 -674 2065 -646
rect 2093 -674 2131 -646
rect 2159 -674 2197 -646
rect 2225 -674 2263 -646
rect 2291 -674 2329 -646
rect 2357 -674 2395 -646
rect 2423 -674 2461 -646
rect 2489 -674 2527 -646
rect 2555 -674 2593 -646
rect 2621 -674 2659 -646
rect 2687 -674 2725 -646
rect 2753 -674 2791 -646
rect 2819 -674 2857 -646
rect 2885 -674 2923 -646
rect 2951 -674 2989 -646
rect 3017 -674 3055 -646
rect 3083 -674 3121 -646
rect 3149 -674 3187 -646
rect 3215 -674 3253 -646
rect 3281 -674 3319 -646
rect 3347 -674 3385 -646
rect 3413 -674 3451 -646
rect 3479 -674 3517 -646
rect 3545 -674 3583 -646
rect 3611 -674 3649 -646
rect 3677 -674 3715 -646
rect 3743 -674 3781 -646
rect 3809 -674 3847 -646
rect 3875 -674 3883 -646
rect -3883 -712 3883 -674
rect -3883 -740 -3875 -712
rect -3847 -740 -3809 -712
rect -3781 -740 -3743 -712
rect -3715 -740 -3677 -712
rect -3649 -740 -3611 -712
rect -3583 -740 -3545 -712
rect -3517 -740 -3479 -712
rect -3451 -740 -3413 -712
rect -3385 -740 -3347 -712
rect -3319 -740 -3281 -712
rect -3253 -740 -3215 -712
rect -3187 -740 -3149 -712
rect -3121 -740 -3083 -712
rect -3055 -740 -3017 -712
rect -2989 -740 -2951 -712
rect -2923 -740 -2885 -712
rect -2857 -740 -2819 -712
rect -2791 -740 -2753 -712
rect -2725 -740 -2687 -712
rect -2659 -740 -2621 -712
rect -2593 -740 -2555 -712
rect -2527 -740 -2489 -712
rect -2461 -740 -2423 -712
rect -2395 -740 -2357 -712
rect -2329 -740 -2291 -712
rect -2263 -740 -2225 -712
rect -2197 -740 -2159 -712
rect -2131 -740 -2093 -712
rect -2065 -740 -2027 -712
rect -1999 -740 -1961 -712
rect -1933 -740 -1895 -712
rect -1867 -740 -1829 -712
rect -1801 -740 -1763 -712
rect -1735 -740 -1697 -712
rect -1669 -740 -1631 -712
rect -1603 -740 -1565 -712
rect -1537 -740 -1499 -712
rect -1471 -740 -1433 -712
rect -1405 -740 -1367 -712
rect -1339 -740 -1301 -712
rect -1273 -740 -1235 -712
rect -1207 -740 -1169 -712
rect -1141 -740 -1103 -712
rect -1075 -740 -1037 -712
rect -1009 -740 -971 -712
rect -943 -740 -905 -712
rect -877 -740 -839 -712
rect -811 -740 -773 -712
rect -745 -740 -707 -712
rect -679 -740 -641 -712
rect -613 -740 -575 -712
rect -547 -740 -509 -712
rect -481 -740 -443 -712
rect -415 -740 -377 -712
rect -349 -740 -311 -712
rect -283 -740 -245 -712
rect -217 -740 -179 -712
rect -151 -740 -113 -712
rect -85 -740 -47 -712
rect -19 -740 19 -712
rect 47 -740 85 -712
rect 113 -740 151 -712
rect 179 -740 217 -712
rect 245 -740 283 -712
rect 311 -740 349 -712
rect 377 -740 415 -712
rect 443 -740 481 -712
rect 509 -740 547 -712
rect 575 -740 613 -712
rect 641 -740 679 -712
rect 707 -740 745 -712
rect 773 -740 811 -712
rect 839 -740 877 -712
rect 905 -740 943 -712
rect 971 -740 1009 -712
rect 1037 -740 1075 -712
rect 1103 -740 1141 -712
rect 1169 -740 1207 -712
rect 1235 -740 1273 -712
rect 1301 -740 1339 -712
rect 1367 -740 1405 -712
rect 1433 -740 1471 -712
rect 1499 -740 1537 -712
rect 1565 -740 1603 -712
rect 1631 -740 1669 -712
rect 1697 -740 1735 -712
rect 1763 -740 1801 -712
rect 1829 -740 1867 -712
rect 1895 -740 1933 -712
rect 1961 -740 1999 -712
rect 2027 -740 2065 -712
rect 2093 -740 2131 -712
rect 2159 -740 2197 -712
rect 2225 -740 2263 -712
rect 2291 -740 2329 -712
rect 2357 -740 2395 -712
rect 2423 -740 2461 -712
rect 2489 -740 2527 -712
rect 2555 -740 2593 -712
rect 2621 -740 2659 -712
rect 2687 -740 2725 -712
rect 2753 -740 2791 -712
rect 2819 -740 2857 -712
rect 2885 -740 2923 -712
rect 2951 -740 2989 -712
rect 3017 -740 3055 -712
rect 3083 -740 3121 -712
rect 3149 -740 3187 -712
rect 3215 -740 3253 -712
rect 3281 -740 3319 -712
rect 3347 -740 3385 -712
rect 3413 -740 3451 -712
rect 3479 -740 3517 -712
rect 3545 -740 3583 -712
rect 3611 -740 3649 -712
rect 3677 -740 3715 -712
rect 3743 -740 3781 -712
rect 3809 -740 3847 -712
rect 3875 -740 3883 -712
rect -3883 -748 3883 -740
<< end >>
