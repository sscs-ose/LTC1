magic
tech gf180mcuC
magscale 1 10
timestamp 1714126980
<< error_p >>
rect -371 -48 -325 48
rect -197 -48 -151 48
rect -23 -48 23 48
rect 151 -48 197 48
rect 325 -48 371 48
<< nwell >>
rect -470 -180 470 180
<< pmos >>
rect -296 -50 -226 50
rect -122 -50 -52 50
rect 52 -50 122 50
rect 226 -50 296 50
<< pdiff >>
rect -384 37 -296 50
rect -384 -37 -371 37
rect -325 -37 -296 37
rect -384 -50 -296 -37
rect -226 37 -122 50
rect -226 -37 -197 37
rect -151 -37 -122 37
rect -226 -50 -122 -37
rect -52 37 52 50
rect -52 -37 -23 37
rect 23 -37 52 37
rect -52 -50 52 -37
rect 122 37 226 50
rect 122 -37 151 37
rect 197 -37 226 37
rect 122 -50 226 -37
rect 296 37 384 50
rect 296 -37 325 37
rect 371 -37 384 37
rect 296 -50 384 -37
<< pdiffc >>
rect -371 -37 -325 37
rect -197 -37 -151 37
rect -23 -37 23 37
rect 151 -37 197 37
rect 325 -37 371 37
<< polysilicon >>
rect -296 50 -226 94
rect -122 50 -52 94
rect 52 50 122 94
rect 226 50 296 94
rect -296 -94 -226 -50
rect -122 -94 -52 -50
rect 52 -94 122 -50
rect 226 -94 296 -50
<< metal1 >>
rect -371 37 -325 48
rect -371 -48 -325 -37
rect -197 37 -151 48
rect -197 -48 -151 -37
rect -23 37 23 48
rect -23 -48 23 -37
rect 151 37 197 48
rect 151 -48 197 -37
rect 325 37 371 48
rect 325 -48 371 -37
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 0.5 l 0.35 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
