magic
tech gf180mcuC
magscale 1 10
timestamp 1699986627
<< metal1 >>
rect 3663 19860 128522 20014
rect 3663 19845 113574 19860
rect 3663 19789 24715 19845
rect 24771 19789 24825 19845
rect 24881 19789 24935 19845
rect 24991 19789 25045 19845
rect 25101 19789 25155 19845
rect 25211 19789 25265 19845
rect 25321 19789 25375 19845
rect 25431 19804 113574 19845
rect 113630 19804 113684 19860
rect 113740 19804 113794 19860
rect 113850 19804 113904 19860
rect 113960 19804 114014 19860
rect 114070 19804 114124 19860
rect 114180 19804 114234 19860
rect 114290 19804 128522 19860
rect 25431 19789 128522 19804
rect 3663 19750 128522 19789
rect 3663 19735 113574 19750
rect 3663 19679 24715 19735
rect 24771 19679 24825 19735
rect 24881 19679 24935 19735
rect 24991 19679 25045 19735
rect 25101 19679 25155 19735
rect 25211 19679 25265 19735
rect 25321 19679 25375 19735
rect 25431 19694 113574 19735
rect 113630 19694 113684 19750
rect 113740 19694 113794 19750
rect 113850 19694 113904 19750
rect 113960 19694 114014 19750
rect 114070 19694 114124 19750
rect 114180 19694 114234 19750
rect 114290 19694 128522 19750
rect 25431 19679 128522 19694
rect 3663 19640 128522 19679
rect 3663 19625 113574 19640
rect 3663 19569 24715 19625
rect 24771 19569 24825 19625
rect 24881 19569 24935 19625
rect 24991 19569 25045 19625
rect 25101 19569 25155 19625
rect 25211 19569 25265 19625
rect 25321 19569 25375 19625
rect 25431 19584 113574 19625
rect 113630 19584 113684 19640
rect 113740 19584 113794 19640
rect 113850 19584 113904 19640
rect 113960 19584 114014 19640
rect 114070 19584 114124 19640
rect 114180 19584 114234 19640
rect 114290 19584 128522 19640
rect 25431 19569 128522 19584
rect 3663 19530 128522 19569
rect 3663 19515 113574 19530
rect 3663 19459 24715 19515
rect 24771 19459 24825 19515
rect 24881 19459 24935 19515
rect 24991 19459 25045 19515
rect 25101 19459 25155 19515
rect 25211 19459 25265 19515
rect 25321 19459 25375 19515
rect 25431 19474 113574 19515
rect 113630 19474 113684 19530
rect 113740 19474 113794 19530
rect 113850 19474 113904 19530
rect 113960 19474 114014 19530
rect 114070 19474 114124 19530
rect 114180 19474 114234 19530
rect 114290 19474 128522 19530
rect 25431 19459 128522 19474
rect 3663 19420 128522 19459
rect 3663 19405 113574 19420
rect 3663 19349 24715 19405
rect 24771 19349 24825 19405
rect 24881 19349 24935 19405
rect 24991 19349 25045 19405
rect 25101 19349 25155 19405
rect 25211 19349 25265 19405
rect 25321 19349 25375 19405
rect 25431 19364 113574 19405
rect 113630 19364 113684 19420
rect 113740 19364 113794 19420
rect 113850 19364 113904 19420
rect 113960 19364 114014 19420
rect 114070 19364 114124 19420
rect 114180 19364 114234 19420
rect 114290 19364 128522 19420
rect 25431 19349 128522 19364
rect 3663 19310 128522 19349
rect 3663 19295 113574 19310
rect 3663 19239 24715 19295
rect 24771 19239 24825 19295
rect 24881 19239 24935 19295
rect 24991 19239 25045 19295
rect 25101 19239 25155 19295
rect 25211 19239 25265 19295
rect 25321 19239 25375 19295
rect 25431 19254 113574 19295
rect 113630 19254 113684 19310
rect 113740 19254 113794 19310
rect 113850 19254 113904 19310
rect 113960 19254 114014 19310
rect 114070 19254 114124 19310
rect 114180 19254 114234 19310
rect 114290 19254 128522 19310
rect 25431 19239 128522 19254
rect 3663 19114 128522 19239
rect 7038 15257 8653 19114
rect 9433 18785 25861 18786
rect 26830 18785 114552 18786
rect 115597 18785 128522 18786
rect 9433 18616 128522 18785
rect 9433 18560 25931 18616
rect 25987 18560 26041 18616
rect 26097 18560 26151 18616
rect 26207 18560 26261 18616
rect 26317 18560 26371 18616
rect 26427 18560 26481 18616
rect 26537 18560 26591 18616
rect 26647 18575 128522 18616
rect 26647 18560 114647 18575
rect 9433 18519 114647 18560
rect 114703 18519 114757 18575
rect 114813 18519 114867 18575
rect 114923 18519 114977 18575
rect 115033 18519 115087 18575
rect 115143 18519 115197 18575
rect 115253 18519 115307 18575
rect 115363 18519 128522 18575
rect 9433 18506 128522 18519
rect 9433 18450 25931 18506
rect 25987 18450 26041 18506
rect 26097 18450 26151 18506
rect 26207 18450 26261 18506
rect 26317 18450 26371 18506
rect 26427 18450 26481 18506
rect 26537 18450 26591 18506
rect 26647 18465 128522 18506
rect 26647 18450 114647 18465
rect 9433 18409 114647 18450
rect 114703 18409 114757 18465
rect 114813 18409 114867 18465
rect 114923 18409 114977 18465
rect 115033 18409 115087 18465
rect 115143 18409 115197 18465
rect 115253 18409 115307 18465
rect 115363 18409 128522 18465
rect 9433 18396 128522 18409
rect 9433 18340 25931 18396
rect 25987 18340 26041 18396
rect 26097 18340 26151 18396
rect 26207 18340 26261 18396
rect 26317 18340 26371 18396
rect 26427 18340 26481 18396
rect 26537 18340 26591 18396
rect 26647 18355 128522 18396
rect 26647 18340 114647 18355
rect 9433 18299 114647 18340
rect 114703 18299 114757 18355
rect 114813 18299 114867 18355
rect 114923 18299 114977 18355
rect 115033 18299 115087 18355
rect 115143 18299 115197 18355
rect 115253 18299 115307 18355
rect 115363 18299 128522 18355
rect 9433 18286 128522 18299
rect 9433 18230 25931 18286
rect 25987 18230 26041 18286
rect 26097 18230 26151 18286
rect 26207 18230 26261 18286
rect 26317 18230 26371 18286
rect 26427 18230 26481 18286
rect 26537 18230 26591 18286
rect 26647 18245 128522 18286
rect 26647 18230 114647 18245
rect 9433 18189 114647 18230
rect 114703 18189 114757 18245
rect 114813 18189 114867 18245
rect 114923 18189 114977 18245
rect 115033 18189 115087 18245
rect 115143 18189 115197 18245
rect 115253 18189 115307 18245
rect 115363 18189 128522 18245
rect 9433 18176 128522 18189
rect 9433 18120 25931 18176
rect 25987 18120 26041 18176
rect 26097 18120 26151 18176
rect 26207 18120 26261 18176
rect 26317 18120 26371 18176
rect 26427 18120 26481 18176
rect 26537 18120 26591 18176
rect 26647 18135 128522 18176
rect 26647 18120 114647 18135
rect 9433 18079 114647 18120
rect 114703 18079 114757 18135
rect 114813 18079 114867 18135
rect 114923 18079 114977 18135
rect 115033 18079 115087 18135
rect 115143 18079 115197 18135
rect 115253 18079 115307 18135
rect 115363 18079 128522 18135
rect 9433 18066 128522 18079
rect 9433 18010 25931 18066
rect 25987 18010 26041 18066
rect 26097 18010 26151 18066
rect 26207 18010 26261 18066
rect 26317 18010 26371 18066
rect 26427 18010 26481 18066
rect 26537 18010 26591 18066
rect 26647 18025 128522 18066
rect 26647 18010 114647 18025
rect 9433 17969 114647 18010
rect 114703 17969 114757 18025
rect 114813 17969 114867 18025
rect 114923 17969 114977 18025
rect 115033 17969 115087 18025
rect 115143 17969 115197 18025
rect 115253 17969 115307 18025
rect 115363 17969 128522 18025
rect 9433 17886 128522 17969
rect 55786 15424 56696 17886
rect 59193 15346 60103 17886
rect 62184 15476 63094 17886
rect 65305 15398 66215 17886
rect 67905 15476 68815 17886
rect 71338 15372 72248 17886
rect 73653 15294 74563 17886
rect 113495 13098 114290 13134
rect 113495 13042 113535 13098
rect 113591 13042 113645 13098
rect 113701 13042 113755 13098
rect 113811 13042 113865 13098
rect 113921 13042 113975 13098
rect 114031 13042 114085 13098
rect 114141 13042 114195 13098
rect 114251 13042 114290 13098
rect 113495 12988 114290 13042
rect 113495 12932 113535 12988
rect 113591 12932 113645 12988
rect 113701 12932 113755 12988
rect 113811 12932 113865 12988
rect 113921 12932 113975 12988
rect 114031 12932 114085 12988
rect 114141 12932 114195 12988
rect 114251 12968 114290 12988
rect 114251 12932 129059 12968
rect 113495 12878 129059 12932
rect 113495 12822 113535 12878
rect 113591 12822 113645 12878
rect 113701 12822 113755 12878
rect 113811 12822 113865 12878
rect 113921 12822 113975 12878
rect 114031 12822 114085 12878
rect 114141 12822 114195 12878
rect 114251 12822 129059 12878
rect 113495 12768 129059 12822
rect 113495 12712 113535 12768
rect 113591 12712 113645 12768
rect 113701 12712 113755 12768
rect 113811 12712 113865 12768
rect 113921 12712 113975 12768
rect 114031 12712 114085 12768
rect 114141 12712 114195 12768
rect 114251 12712 129059 12768
rect 113495 12658 129059 12712
rect 113495 12602 113535 12658
rect 113591 12602 113645 12658
rect 113701 12602 113755 12658
rect 113811 12602 113865 12658
rect 113921 12602 113975 12658
rect 114031 12602 114085 12658
rect 114141 12602 114195 12658
rect 114251 12602 129059 12658
rect 113495 12548 129059 12602
rect 113495 12492 113535 12548
rect 113591 12492 113645 12548
rect 113701 12492 113755 12548
rect 113811 12492 113865 12548
rect 113921 12492 113975 12548
rect 114031 12492 114085 12548
rect 114141 12492 114195 12548
rect 114251 12511 129059 12548
rect 114251 12492 114290 12511
rect 113495 12452 114290 12492
rect 3200 3035 3627 11341
rect 129229 10872 131180 11421
rect 129237 10561 131188 10567
rect 129237 10385 131196 10561
rect 129237 10018 131188 10385
rect 116760 9949 116770 10005
rect 116826 9949 116836 10005
rect 129233 8972 131184 9347
rect 129233 8796 131196 8972
rect 129224 8466 131175 8641
rect 116723 8430 116888 8438
rect 116723 8374 116770 8430
rect 116826 8374 116888 8430
rect 116723 8320 116888 8374
rect 116723 8264 116770 8320
rect 116826 8264 116888 8320
rect 116723 8210 116888 8264
rect 116723 8154 116770 8210
rect 116826 8154 116888 8210
rect 116723 8100 116888 8154
rect 116723 8044 116770 8100
rect 116826 8044 116888 8100
rect 129224 8290 131185 8466
rect 129224 8092 131175 8290
rect 116723 7990 116888 8044
rect 116723 7934 116770 7990
rect 116826 7934 116888 7990
rect 116723 7880 116888 7934
rect 116723 7824 116770 7880
rect 116826 7824 116888 7880
rect 129237 7832 130481 7872
rect 129237 7830 130252 7832
rect 116723 7787 116888 7824
rect 129233 7774 129243 7830
rect 129299 7774 129353 7830
rect 129409 7776 130252 7830
rect 130308 7776 130362 7832
rect 130418 7776 130481 7832
rect 129409 7774 130481 7776
rect 129237 7740 130481 7774
rect 46392 6309 46957 6314
rect 43879 6293 44495 6294
rect 43879 6250 44498 6293
rect 43879 6194 43928 6250
rect 43984 6194 44038 6250
rect 44094 6194 44148 6250
rect 44204 6194 44258 6250
rect 44314 6194 44368 6250
rect 44424 6194 44498 6250
rect 43879 6140 44498 6194
rect 43879 6084 43928 6140
rect 43984 6084 44038 6140
rect 44094 6084 44148 6140
rect 44204 6084 44258 6140
rect 44314 6084 44368 6140
rect 44424 6084 44498 6140
rect 43879 6030 44498 6084
rect 43879 5974 43928 6030
rect 43984 5974 44038 6030
rect 44094 5974 44148 6030
rect 44204 5974 44258 6030
rect 44314 5974 44368 6030
rect 44424 5998 44498 6030
rect 46392 6253 46418 6309
rect 46474 6253 46528 6309
rect 46584 6253 46638 6309
rect 46694 6253 46748 6309
rect 46804 6253 46858 6309
rect 46914 6290 46957 6309
rect 46914 6253 46958 6290
rect 46392 6199 46958 6253
rect 46392 6143 46638 6199
rect 46694 6143 46748 6199
rect 46804 6143 46858 6199
rect 46914 6143 46958 6199
rect 46392 6089 46958 6143
rect 46392 6033 46638 6089
rect 46694 6033 46748 6089
rect 46804 6033 46858 6089
rect 46914 6033 46958 6089
rect 44424 5974 44495 5998
rect 46392 5996 46958 6033
rect 43879 5958 44495 5974
rect -1632 2948 3627 3035
rect -1632 2892 -808 2948
rect -752 2892 -698 2948
rect -642 2892 -588 2948
rect -532 2892 -478 2948
rect -422 2892 -368 2948
rect -312 2892 -258 2948
rect -202 2892 -148 2948
rect -92 2892 3627 2948
rect -1632 2838 3627 2892
rect -1632 2782 -808 2838
rect -752 2782 -698 2838
rect -642 2782 -588 2838
rect -532 2782 -478 2838
rect -422 2782 -368 2838
rect -312 2782 -258 2838
rect -202 2782 -148 2838
rect -92 2782 3627 2838
rect 10737 3443 12429 3485
rect 10737 3387 10800 3443
rect 10856 3387 10910 3443
rect 10966 3387 11020 3443
rect 11076 3387 11130 3443
rect 11186 3387 11240 3443
rect 11296 3387 11350 3443
rect 11406 3387 11460 3443
rect 11516 3387 11624 3443
rect 11680 3387 11734 3443
rect 11790 3387 11844 3443
rect 11900 3387 11954 3443
rect 12010 3387 12064 3443
rect 12120 3387 12174 3443
rect 12230 3387 12284 3443
rect 12340 3387 12429 3443
rect 10737 3333 12429 3387
rect 10737 3277 10800 3333
rect 10856 3277 10910 3333
rect 10966 3277 11020 3333
rect 11076 3277 11130 3333
rect 11186 3277 11240 3333
rect 11296 3277 11350 3333
rect 11406 3277 11460 3333
rect 11516 3277 11624 3333
rect 11680 3277 11734 3333
rect 11790 3277 11844 3333
rect 11900 3277 11954 3333
rect 12010 3277 12064 3333
rect 12120 3277 12174 3333
rect 12230 3277 12284 3333
rect 12340 3277 12429 3333
rect 10737 3223 12429 3277
rect 10737 3167 10800 3223
rect 10856 3167 10910 3223
rect 10966 3167 11020 3223
rect 11076 3167 11130 3223
rect 11186 3167 11240 3223
rect 11296 3167 11350 3223
rect 11406 3167 11460 3223
rect 11516 3167 11624 3223
rect 11680 3167 11734 3223
rect 11790 3167 11844 3223
rect 11900 3167 11954 3223
rect 12010 3167 12064 3223
rect 12120 3167 12174 3223
rect 12230 3167 12284 3223
rect 12340 3167 12429 3223
rect 10737 3113 12429 3167
rect 10737 3057 10800 3113
rect 10856 3057 10910 3113
rect 10966 3057 11020 3113
rect 11076 3057 11130 3113
rect 11186 3057 11240 3113
rect 11296 3057 11350 3113
rect 11406 3057 11460 3113
rect 11516 3057 11624 3113
rect 11680 3057 11734 3113
rect 11790 3057 11844 3113
rect 11900 3057 11954 3113
rect 12010 3057 12064 3113
rect 12120 3057 12174 3113
rect 12230 3057 12284 3113
rect 12340 3057 12429 3113
rect 10737 3003 12429 3057
rect 10737 2947 10800 3003
rect 10856 2947 10910 3003
rect 10966 2947 11020 3003
rect 11076 2947 11130 3003
rect 11186 2947 11240 3003
rect 11296 2947 11350 3003
rect 11406 2947 11460 3003
rect 11516 2947 11624 3003
rect 11680 2947 11734 3003
rect 11790 2947 11844 3003
rect 11900 2947 11954 3003
rect 12010 2947 12064 3003
rect 12120 2947 12174 3003
rect 12230 2947 12284 3003
rect 12340 2947 12429 3003
rect 10737 2893 12429 2947
rect 10737 2837 10800 2893
rect 10856 2837 10910 2893
rect 10966 2837 11020 2893
rect 11076 2837 11130 2893
rect 11186 2837 11240 2893
rect 11296 2837 11350 2893
rect 11406 2837 11460 2893
rect 11516 2837 11624 2893
rect 11680 2837 11734 2893
rect 11790 2837 11844 2893
rect 11900 2837 11954 2893
rect 12010 2837 12064 2893
rect 12120 2837 12174 2893
rect 12230 2837 12284 2893
rect 12340 2837 12429 2893
rect 10737 2795 12429 2837
rect -1632 2728 3627 2782
rect -1632 2672 -808 2728
rect -752 2672 -698 2728
rect -642 2672 -588 2728
rect -532 2672 -478 2728
rect -422 2672 -368 2728
rect -312 2672 -258 2728
rect -202 2672 -148 2728
rect -92 2672 3627 2728
rect -1632 2637 3627 2672
rect -1632 2618 3111 2637
rect -1632 2562 -808 2618
rect -752 2562 -698 2618
rect -642 2562 -588 2618
rect -532 2562 -478 2618
rect -422 2562 -368 2618
rect -312 2562 -258 2618
rect -202 2562 -148 2618
rect -92 2581 3111 2618
rect 3167 2581 3221 2637
rect 3277 2581 3331 2637
rect 3387 2581 3441 2637
rect 3497 2581 3627 2637
rect -92 2562 3627 2581
rect -1632 2527 3627 2562
rect -1632 2508 3111 2527
rect -1632 2452 -808 2508
rect -752 2452 -698 2508
rect -642 2452 -588 2508
rect -532 2452 -478 2508
rect -422 2452 -368 2508
rect -312 2452 -258 2508
rect -202 2452 -148 2508
rect -92 2471 3111 2508
rect 3167 2471 3221 2527
rect 3277 2471 3331 2527
rect 3387 2471 3441 2527
rect 3497 2471 3627 2527
rect -92 2452 3627 2471
rect -1632 2417 3627 2452
rect -1632 2398 3111 2417
rect -1632 2342 -808 2398
rect -752 2342 -698 2398
rect -642 2342 -588 2398
rect -532 2342 -478 2398
rect -422 2342 -368 2398
rect -312 2342 -258 2398
rect -202 2342 -148 2398
rect -92 2361 3111 2398
rect 3167 2361 3221 2417
rect 3277 2361 3331 2417
rect 3387 2361 3441 2417
rect 3497 2361 3627 2417
rect -92 2342 3627 2361
rect -1632 2307 3627 2342
rect -1632 2282 3111 2307
rect 3089 2251 3111 2282
rect 3167 2251 3221 2307
rect 3277 2251 3331 2307
rect 3387 2251 3441 2307
rect 3497 2251 3627 2307
rect 3089 2226 3627 2251
rect 6286 1204 7074 1217
rect 22871 1204 23661 1220
rect 28340 1204 29128 1206
rect 43885 1204 44489 5958
rect 6286 1192 23661 1204
rect 6286 1186 22896 1192
rect 6286 1130 6315 1186
rect 6371 1130 6425 1186
rect 6481 1130 6535 1186
rect 6591 1130 6645 1186
rect 6701 1130 6755 1186
rect 6811 1130 6865 1186
rect 6921 1130 6975 1186
rect 7031 1136 22896 1186
rect 22952 1136 23006 1192
rect 23062 1136 23116 1192
rect 23172 1136 23226 1192
rect 23282 1136 23336 1192
rect 23392 1136 23446 1192
rect 23502 1136 23556 1192
rect 23612 1136 23661 1192
rect 7031 1130 23661 1136
rect 6286 1082 23661 1130
rect 6286 1076 22896 1082
rect 6286 1020 6315 1076
rect 6371 1020 6425 1076
rect 6481 1020 6535 1076
rect 6591 1020 6645 1076
rect 6701 1020 6755 1076
rect 6811 1020 6865 1076
rect 6921 1020 6975 1076
rect 7031 1026 22896 1076
rect 22952 1026 23006 1082
rect 23062 1026 23116 1082
rect 23172 1026 23226 1082
rect 23282 1026 23336 1082
rect 23392 1026 23446 1082
rect 23502 1026 23556 1082
rect 23612 1026 23661 1082
rect 7031 1020 23661 1026
rect 6286 972 23661 1020
rect 6286 966 22896 972
rect 6286 910 6315 966
rect 6371 910 6425 966
rect 6481 910 6535 966
rect 6591 910 6645 966
rect 6701 910 6755 966
rect 6811 910 6865 966
rect 6921 910 6975 966
rect 7031 916 22896 966
rect 22952 916 23006 972
rect 23062 916 23116 972
rect 23172 916 23226 972
rect 23282 916 23336 972
rect 23392 916 23446 972
rect 23502 916 23556 972
rect 23612 916 23661 972
rect 7031 910 23661 916
rect 6286 862 23661 910
rect 6286 856 22896 862
rect 6286 800 6315 856
rect 6371 800 6425 856
rect 6481 800 6535 856
rect 6591 800 6645 856
rect 6701 800 6755 856
rect 6811 800 6865 856
rect 6921 800 6975 856
rect 7031 806 22896 856
rect 22952 806 23006 862
rect 23062 806 23116 862
rect 23172 806 23226 862
rect 23282 806 23336 862
rect 23392 806 23446 862
rect 23502 806 23556 862
rect 23612 806 23661 862
rect 7031 800 23661 806
rect 6286 752 23661 800
rect 6286 746 22896 752
rect 6286 690 6315 746
rect 6371 690 6425 746
rect 6481 690 6535 746
rect 6591 690 6645 746
rect 6701 690 6755 746
rect 6811 690 6865 746
rect 6921 690 6975 746
rect 7031 696 22896 746
rect 22952 696 23006 752
rect 23062 696 23116 752
rect 23172 696 23226 752
rect 23282 696 23336 752
rect 23392 696 23446 752
rect 23502 696 23556 752
rect 23612 696 23661 752
rect 7031 690 23661 696
rect 6286 642 23661 690
rect 6286 636 22896 642
rect 6286 580 6315 636
rect 6371 580 6425 636
rect 6481 580 6535 636
rect 6591 580 6645 636
rect 6701 580 6755 636
rect 6811 580 6865 636
rect 6921 580 6975 636
rect 7031 586 22896 636
rect 22952 586 23006 642
rect 23062 586 23116 642
rect 23172 586 23226 642
rect 23282 586 23336 642
rect 23392 586 23446 642
rect 23502 586 23556 642
rect 23612 586 23661 642
rect 7031 580 23661 586
rect 6286 560 23661 580
rect 28331 1188 44529 1204
rect 28331 1132 28369 1188
rect 28425 1132 28479 1188
rect 28535 1132 28589 1188
rect 28645 1132 28699 1188
rect 28755 1132 28809 1188
rect 28865 1132 28919 1188
rect 28975 1132 29029 1188
rect 29085 1132 44529 1188
rect 28331 1078 44529 1132
rect 28331 1022 28369 1078
rect 28425 1022 28479 1078
rect 28535 1022 28589 1078
rect 28645 1022 28699 1078
rect 28755 1022 28809 1078
rect 28865 1022 28919 1078
rect 28975 1022 29029 1078
rect 29085 1022 44529 1078
rect 28331 968 44529 1022
rect 28331 912 28369 968
rect 28425 912 28479 968
rect 28535 912 28589 968
rect 28645 912 28699 968
rect 28755 912 28809 968
rect 28865 912 28919 968
rect 28975 912 29029 968
rect 29085 912 44529 968
rect 28331 858 44529 912
rect 28331 802 28369 858
rect 28425 802 28479 858
rect 28535 802 28589 858
rect 28645 802 28699 858
rect 28755 802 28809 858
rect 28865 802 28919 858
rect 28975 802 29029 858
rect 29085 802 44529 858
rect 28331 748 44529 802
rect 28331 692 28369 748
rect 28425 692 28479 748
rect 28535 692 28589 748
rect 28645 692 28699 748
rect 28755 692 28809 748
rect 28865 692 28919 748
rect 28975 692 29029 748
rect 29085 692 44529 748
rect 28331 638 44529 692
rect 28331 582 28369 638
rect 28425 582 28479 638
rect 28535 582 28589 638
rect 28645 582 28699 638
rect 28755 582 28809 638
rect 28865 582 28919 638
rect 28975 582 29029 638
rect 29085 582 44529 638
rect 28331 560 44529 582
rect 22871 559 23661 560
rect 43885 500 44489 560
rect 7578 377 9499 391
rect 45101 377 45681 2391
rect 46368 377 46948 2418
rect 47594 377 48174 2431
rect 48564 377 49144 2431
rect 62378 377 62961 2038
rect 63802 377 64385 2051
rect 64982 377 65565 2078
rect 67070 377 67653 2038
rect 70285 377 70868 2038
rect 72048 377 72631 1997
rect 73269 377 73852 2065
rect 74543 377 75126 2024
rect 97978 377 98736 7500
rect 99825 377 100583 7610
rect 101479 377 102237 7527
rect 103491 377 104249 7569
rect 104952 377 105710 7624
rect 116723 6920 116888 6928
rect 116723 6864 116770 6920
rect 116826 6864 116888 6920
rect 116723 6810 116888 6864
rect 107171 6784 116351 6808
rect 107171 6728 107204 6784
rect 107260 6728 107314 6784
rect 107370 6728 107424 6784
rect 107480 6728 107534 6784
rect 107590 6728 107644 6784
rect 107700 6728 107754 6784
rect 107810 6728 107864 6784
rect 107920 6728 116351 6784
rect 107171 6674 116351 6728
rect 107171 6618 107204 6674
rect 107260 6618 107314 6674
rect 107370 6618 107424 6674
rect 107480 6618 107534 6674
rect 107590 6618 107644 6674
rect 107700 6618 107754 6674
rect 107810 6618 107864 6674
rect 107920 6618 116351 6674
rect 107171 6564 116351 6618
rect 107171 6508 107204 6564
rect 107260 6508 107314 6564
rect 107370 6508 107424 6564
rect 107480 6508 107534 6564
rect 107590 6508 107644 6564
rect 107700 6508 107754 6564
rect 107810 6508 107864 6564
rect 107920 6508 116351 6564
rect 107171 6454 116351 6508
rect 107171 6398 107204 6454
rect 107260 6398 107314 6454
rect 107370 6398 107424 6454
rect 107480 6398 107534 6454
rect 107590 6398 107644 6454
rect 107700 6398 107754 6454
rect 107810 6398 107864 6454
rect 107920 6398 116351 6454
rect 107171 6344 116351 6398
rect 107171 6288 107204 6344
rect 107260 6288 107314 6344
rect 107370 6288 107424 6344
rect 107480 6288 107534 6344
rect 107590 6288 107644 6344
rect 107700 6288 107754 6344
rect 107810 6288 107864 6344
rect 107920 6288 116351 6344
rect 107171 6234 116351 6288
rect 116723 6754 116770 6810
rect 116826 6754 116888 6810
rect 116723 6700 116888 6754
rect 116723 6644 116770 6700
rect 116826 6644 116888 6700
rect 116723 6590 116888 6644
rect 116723 6534 116770 6590
rect 116826 6534 116888 6590
rect 116723 6480 116888 6534
rect 116723 6424 116770 6480
rect 116826 6424 116888 6480
rect 116723 6370 116888 6424
rect 116723 6314 116770 6370
rect 116826 6314 116888 6370
rect 116723 6277 116888 6314
rect 107171 6178 107204 6234
rect 107260 6178 107314 6234
rect 107370 6178 107424 6234
rect 107480 6178 107534 6234
rect 107590 6178 107644 6234
rect 107700 6178 107754 6234
rect 107810 6178 107864 6234
rect 107920 6178 116351 6234
rect 129256 6230 131207 6779
rect 107171 6124 116351 6178
rect 107171 6068 107204 6124
rect 107260 6068 107314 6124
rect 107370 6068 107424 6124
rect 107480 6068 107534 6124
rect 107590 6068 107644 6124
rect 107700 6068 107754 6124
rect 107810 6068 107864 6124
rect 107920 6068 116351 6124
rect 107171 6014 116351 6068
rect 107171 5958 107204 6014
rect 107260 5958 107314 6014
rect 107370 5958 107424 6014
rect 107480 5958 107534 6014
rect 107590 5958 107644 6014
rect 107700 5958 107754 6014
rect 107810 5958 107864 6014
rect 107920 5958 116351 6014
rect 107171 5938 116351 5958
rect 129240 5567 131191 6116
rect 116723 5500 116888 5508
rect 116723 5444 116770 5500
rect 116826 5444 116888 5500
rect 116723 5390 116888 5444
rect 116723 5334 116770 5390
rect 116826 5334 116888 5390
rect 116723 5280 116888 5334
rect 116723 5224 116770 5280
rect 116826 5224 116888 5280
rect 129242 5338 130828 5366
rect 129242 5333 130585 5338
rect 129242 5277 129259 5333
rect 129315 5277 129369 5333
rect 129425 5282 130585 5333
rect 130641 5282 130695 5338
rect 130751 5282 130828 5338
rect 129425 5277 130828 5282
rect 129242 5241 130828 5277
rect 116723 5170 116888 5224
rect 116723 5114 116770 5170
rect 116826 5114 116888 5170
rect 116723 5060 116888 5114
rect 116723 5004 116770 5060
rect 116826 5004 116888 5060
rect 116723 4950 116888 5004
rect 116723 4894 116770 4950
rect 116826 4894 116888 4950
rect 116723 4857 116888 4894
rect 129297 4091 131248 4640
rect 129180 3267 131131 3816
rect 117172 377 117438 2225
rect 117919 377 118185 2233
rect 119423 377 119689 2267
rect 120425 377 120691 2233
rect 121361 377 121627 2247
rect 122056 377 122322 2233
rect 122931 377 123197 2240
rect 123834 377 124100 2272
rect 124539 377 124805 2272
rect 125597 377 125868 2258
rect 126502 377 126773 2246
rect 127325 377 127596 2211
rect 128348 377 128619 2246
rect 5980 214 128736 377
rect 5980 159 29849 214
rect 5980 103 24709 159
rect 24765 103 24819 159
rect 24875 103 24929 159
rect 24985 103 25039 159
rect 25095 103 25149 159
rect 25205 103 25259 159
rect 25315 103 25369 159
rect 25425 158 29849 159
rect 29905 158 29959 214
rect 30015 158 30069 214
rect 30125 158 30179 214
rect 30235 158 30289 214
rect 30345 158 30399 214
rect 30455 158 30509 214
rect 30565 211 128736 214
rect 30565 158 113565 211
rect 25425 155 113565 158
rect 113621 155 113675 211
rect 113731 155 113785 211
rect 113841 155 113895 211
rect 113951 155 114005 211
rect 114061 155 114115 211
rect 114171 155 114225 211
rect 114281 155 128736 211
rect 25425 118 128736 155
rect 25425 114 89511 118
rect 25425 108 74565 114
rect 25425 104 71847 108
rect 25425 103 29849 104
rect 5980 49 29849 103
rect 5980 -7 24709 49
rect 24765 -7 24819 49
rect 24875 -7 24929 49
rect 24985 -7 25039 49
rect 25095 -7 25149 49
rect 25205 -7 25259 49
rect 25315 -7 25369 49
rect 25425 48 29849 49
rect 29905 48 29959 104
rect 30015 48 30069 104
rect 30125 48 30179 104
rect 30235 48 30289 104
rect 30345 48 30399 104
rect 30455 48 30509 104
rect 30565 103 71847 104
rect 30565 48 69220 103
rect 25425 47 69220 48
rect 69276 47 69330 103
rect 69386 47 69440 103
rect 69496 47 69550 103
rect 69606 47 69660 103
rect 69716 47 69770 103
rect 69826 47 69880 103
rect 69936 52 71847 103
rect 71903 52 71957 108
rect 72013 52 72067 108
rect 72123 52 72177 108
rect 72233 52 72287 108
rect 72343 52 72397 108
rect 72453 52 72507 108
rect 72563 58 74565 108
rect 74621 58 74675 114
rect 74731 58 74785 114
rect 74841 58 74895 114
rect 74951 58 75005 114
rect 75061 58 75115 114
rect 75171 58 75225 114
rect 75281 109 89511 114
rect 75281 100 80687 109
rect 75281 58 77637 100
rect 72563 52 77637 58
rect 69936 47 77637 52
rect 25425 44 77637 47
rect 77693 44 77747 100
rect 77803 44 77857 100
rect 77913 44 77967 100
rect 78023 44 78077 100
rect 78133 44 78187 100
rect 78243 44 78297 100
rect 78353 53 80687 100
rect 80743 53 80797 109
rect 80853 53 80907 109
rect 80963 53 81017 109
rect 81073 53 81127 109
rect 81183 53 81237 109
rect 81293 53 81347 109
rect 81403 53 83528 109
rect 83584 53 83638 109
rect 83694 53 83748 109
rect 83804 53 83858 109
rect 83914 53 83968 109
rect 84024 53 84078 109
rect 84134 53 84188 109
rect 84244 106 89511 109
rect 84244 53 86316 106
rect 78353 50 86316 53
rect 86372 50 86426 106
rect 86482 50 86536 106
rect 86592 50 86646 106
rect 86702 50 86756 106
rect 86812 50 86866 106
rect 86922 50 86976 106
rect 87032 62 89511 106
rect 89567 62 89621 118
rect 89677 62 89731 118
rect 89787 62 89841 118
rect 89897 62 89951 118
rect 90007 62 90061 118
rect 90117 62 90171 118
rect 90227 110 128736 118
rect 90227 107 95994 110
rect 90227 62 92852 107
rect 87032 51 92852 62
rect 92908 51 92962 107
rect 93018 51 93072 107
rect 93128 51 93182 107
rect 93238 51 93292 107
rect 93348 51 93402 107
rect 93458 51 93512 107
rect 93568 54 95994 107
rect 96050 54 96104 110
rect 96160 54 96214 110
rect 96270 54 96324 110
rect 96380 54 96434 110
rect 96490 54 96544 110
rect 96600 54 96654 110
rect 96710 108 128736 110
rect 96710 54 99280 108
rect 93568 52 99280 54
rect 99336 52 99390 108
rect 99446 52 99500 108
rect 99556 52 99610 108
rect 99666 52 99720 108
rect 99776 52 99830 108
rect 99886 52 99940 108
rect 99996 101 128736 108
rect 99996 52 113565 101
rect 93568 51 113565 52
rect 87032 50 113565 51
rect 78353 45 113565 50
rect 113621 45 113675 101
rect 113731 45 113785 101
rect 113841 45 113895 101
rect 113951 45 114005 101
rect 114061 45 114115 101
rect 114171 45 114225 101
rect 114281 45 128736 101
rect 78353 44 128736 45
rect 25425 8 128736 44
rect 25425 4 89511 8
rect 25425 -2 74565 4
rect 25425 -6 71847 -2
rect 25425 -7 29849 -6
rect 5980 -61 29849 -7
rect 5980 -117 24709 -61
rect 24765 -117 24819 -61
rect 24875 -117 24929 -61
rect 24985 -117 25039 -61
rect 25095 -117 25149 -61
rect 25205 -117 25259 -61
rect 25315 -117 25369 -61
rect 25425 -62 29849 -61
rect 29905 -62 29959 -6
rect 30015 -62 30069 -6
rect 30125 -62 30179 -6
rect 30235 -62 30289 -6
rect 30345 -62 30399 -6
rect 30455 -62 30509 -6
rect 30565 -7 71847 -6
rect 30565 -62 69220 -7
rect 25425 -63 69220 -62
rect 69276 -63 69330 -7
rect 69386 -63 69440 -7
rect 69496 -63 69550 -7
rect 69606 -63 69660 -7
rect 69716 -63 69770 -7
rect 69826 -63 69880 -7
rect 69936 -58 71847 -7
rect 71903 -58 71957 -2
rect 72013 -58 72067 -2
rect 72123 -58 72177 -2
rect 72233 -58 72287 -2
rect 72343 -58 72397 -2
rect 72453 -58 72507 -2
rect 72563 -52 74565 -2
rect 74621 -52 74675 4
rect 74731 -52 74785 4
rect 74841 -52 74895 4
rect 74951 -52 75005 4
rect 75061 -52 75115 4
rect 75171 -52 75225 4
rect 75281 -1 89511 4
rect 75281 -10 80687 -1
rect 75281 -52 77637 -10
rect 72563 -58 77637 -52
rect 69936 -63 77637 -58
rect 25425 -66 77637 -63
rect 77693 -66 77747 -10
rect 77803 -66 77857 -10
rect 77913 -66 77967 -10
rect 78023 -66 78077 -10
rect 78133 -66 78187 -10
rect 78243 -66 78297 -10
rect 78353 -57 80687 -10
rect 80743 -57 80797 -1
rect 80853 -57 80907 -1
rect 80963 -57 81017 -1
rect 81073 -57 81127 -1
rect 81183 -57 81237 -1
rect 81293 -57 81347 -1
rect 81403 -57 83528 -1
rect 83584 -57 83638 -1
rect 83694 -57 83748 -1
rect 83804 -57 83858 -1
rect 83914 -57 83968 -1
rect 84024 -57 84078 -1
rect 84134 -57 84188 -1
rect 84244 -4 89511 -1
rect 84244 -57 86316 -4
rect 78353 -60 86316 -57
rect 86372 -60 86426 -4
rect 86482 -60 86536 -4
rect 86592 -60 86646 -4
rect 86702 -60 86756 -4
rect 86812 -60 86866 -4
rect 86922 -60 86976 -4
rect 87032 -48 89511 -4
rect 89567 -48 89621 8
rect 89677 -48 89731 8
rect 89787 -48 89841 8
rect 89897 -48 89951 8
rect 90007 -48 90061 8
rect 90117 -48 90171 8
rect 90227 0 128736 8
rect 90227 -3 95994 0
rect 90227 -48 92852 -3
rect 87032 -59 92852 -48
rect 92908 -59 92962 -3
rect 93018 -59 93072 -3
rect 93128 -59 93182 -3
rect 93238 -59 93292 -3
rect 93348 -59 93402 -3
rect 93458 -59 93512 -3
rect 93568 -56 95994 -3
rect 96050 -56 96104 0
rect 96160 -56 96214 0
rect 96270 -56 96324 0
rect 96380 -56 96434 0
rect 96490 -56 96544 0
rect 96600 -56 96654 0
rect 96710 -2 128736 0
rect 96710 -56 99280 -2
rect 93568 -58 99280 -56
rect 99336 -58 99390 -2
rect 99446 -58 99500 -2
rect 99556 -58 99610 -2
rect 99666 -58 99720 -2
rect 99776 -58 99830 -2
rect 99886 -58 99940 -2
rect 99996 -9 128736 -2
rect 99996 -58 113565 -9
rect 93568 -59 113565 -58
rect 87032 -60 113565 -59
rect 78353 -65 113565 -60
rect 113621 -65 113675 -9
rect 113731 -65 113785 -9
rect 113841 -65 113895 -9
rect 113951 -65 114005 -9
rect 114061 -65 114115 -9
rect 114171 -65 114225 -9
rect 114281 -65 128736 -9
rect 78353 -66 128736 -65
rect 25425 -102 128736 -66
rect 25425 -106 89511 -102
rect 25425 -112 74565 -106
rect 25425 -116 71847 -112
rect 25425 -117 29849 -116
rect 5980 -171 29849 -117
rect 5980 -227 24709 -171
rect 24765 -227 24819 -171
rect 24875 -227 24929 -171
rect 24985 -227 25039 -171
rect 25095 -227 25149 -171
rect 25205 -227 25259 -171
rect 25315 -227 25369 -171
rect 25425 -172 29849 -171
rect 29905 -172 29959 -116
rect 30015 -172 30069 -116
rect 30125 -172 30179 -116
rect 30235 -172 30289 -116
rect 30345 -172 30399 -116
rect 30455 -172 30509 -116
rect 30565 -117 71847 -116
rect 30565 -172 69220 -117
rect 25425 -173 69220 -172
rect 69276 -173 69330 -117
rect 69386 -173 69440 -117
rect 69496 -173 69550 -117
rect 69606 -173 69660 -117
rect 69716 -173 69770 -117
rect 69826 -173 69880 -117
rect 69936 -168 71847 -117
rect 71903 -168 71957 -112
rect 72013 -168 72067 -112
rect 72123 -168 72177 -112
rect 72233 -168 72287 -112
rect 72343 -168 72397 -112
rect 72453 -168 72507 -112
rect 72563 -162 74565 -112
rect 74621 -162 74675 -106
rect 74731 -162 74785 -106
rect 74841 -162 74895 -106
rect 74951 -162 75005 -106
rect 75061 -162 75115 -106
rect 75171 -162 75225 -106
rect 75281 -111 89511 -106
rect 75281 -120 80687 -111
rect 75281 -162 77637 -120
rect 72563 -168 77637 -162
rect 69936 -173 77637 -168
rect 25425 -176 77637 -173
rect 77693 -176 77747 -120
rect 77803 -176 77857 -120
rect 77913 -176 77967 -120
rect 78023 -176 78077 -120
rect 78133 -176 78187 -120
rect 78243 -176 78297 -120
rect 78353 -167 80687 -120
rect 80743 -167 80797 -111
rect 80853 -167 80907 -111
rect 80963 -167 81017 -111
rect 81073 -167 81127 -111
rect 81183 -167 81237 -111
rect 81293 -167 81347 -111
rect 81403 -167 83528 -111
rect 83584 -167 83638 -111
rect 83694 -167 83748 -111
rect 83804 -167 83858 -111
rect 83914 -167 83968 -111
rect 84024 -167 84078 -111
rect 84134 -167 84188 -111
rect 84244 -114 89511 -111
rect 84244 -167 86316 -114
rect 78353 -170 86316 -167
rect 86372 -170 86426 -114
rect 86482 -170 86536 -114
rect 86592 -170 86646 -114
rect 86702 -170 86756 -114
rect 86812 -170 86866 -114
rect 86922 -170 86976 -114
rect 87032 -158 89511 -114
rect 89567 -158 89621 -102
rect 89677 -158 89731 -102
rect 89787 -158 89841 -102
rect 89897 -158 89951 -102
rect 90007 -158 90061 -102
rect 90117 -158 90171 -102
rect 90227 -110 128736 -102
rect 90227 -113 95994 -110
rect 90227 -158 92852 -113
rect 87032 -169 92852 -158
rect 92908 -169 92962 -113
rect 93018 -169 93072 -113
rect 93128 -169 93182 -113
rect 93238 -169 93292 -113
rect 93348 -169 93402 -113
rect 93458 -169 93512 -113
rect 93568 -166 95994 -113
rect 96050 -166 96104 -110
rect 96160 -166 96214 -110
rect 96270 -166 96324 -110
rect 96380 -166 96434 -110
rect 96490 -166 96544 -110
rect 96600 -166 96654 -110
rect 96710 -112 128736 -110
rect 96710 -166 99280 -112
rect 93568 -168 99280 -166
rect 99336 -168 99390 -112
rect 99446 -168 99500 -112
rect 99556 -168 99610 -112
rect 99666 -168 99720 -112
rect 99776 -168 99830 -112
rect 99886 -168 99940 -112
rect 99996 -119 128736 -112
rect 99996 -168 113565 -119
rect 93568 -169 113565 -168
rect 87032 -170 113565 -169
rect 78353 -175 113565 -170
rect 113621 -175 113675 -119
rect 113731 -175 113785 -119
rect 113841 -175 113895 -119
rect 113951 -175 114005 -119
rect 114061 -175 114115 -119
rect 114171 -175 114225 -119
rect 114281 -175 128736 -119
rect 78353 -176 128736 -175
rect 25425 -212 128736 -176
rect 25425 -216 89511 -212
rect 25425 -222 74565 -216
rect 25425 -226 71847 -222
rect 25425 -227 29849 -226
rect 5980 -281 29849 -227
rect 5980 -337 24709 -281
rect 24765 -337 24819 -281
rect 24875 -337 24929 -281
rect 24985 -337 25039 -281
rect 25095 -337 25149 -281
rect 25205 -337 25259 -281
rect 25315 -337 25369 -281
rect 25425 -282 29849 -281
rect 29905 -282 29959 -226
rect 30015 -282 30069 -226
rect 30125 -282 30179 -226
rect 30235 -282 30289 -226
rect 30345 -282 30399 -226
rect 30455 -282 30509 -226
rect 30565 -227 71847 -226
rect 30565 -282 69220 -227
rect 25425 -283 69220 -282
rect 69276 -283 69330 -227
rect 69386 -283 69440 -227
rect 69496 -283 69550 -227
rect 69606 -283 69660 -227
rect 69716 -283 69770 -227
rect 69826 -283 69880 -227
rect 69936 -278 71847 -227
rect 71903 -278 71957 -222
rect 72013 -278 72067 -222
rect 72123 -278 72177 -222
rect 72233 -278 72287 -222
rect 72343 -278 72397 -222
rect 72453 -278 72507 -222
rect 72563 -272 74565 -222
rect 74621 -272 74675 -216
rect 74731 -272 74785 -216
rect 74841 -272 74895 -216
rect 74951 -272 75005 -216
rect 75061 -272 75115 -216
rect 75171 -272 75225 -216
rect 75281 -221 89511 -216
rect 75281 -230 80687 -221
rect 75281 -272 77637 -230
rect 72563 -278 77637 -272
rect 69936 -283 77637 -278
rect 25425 -286 77637 -283
rect 77693 -286 77747 -230
rect 77803 -286 77857 -230
rect 77913 -286 77967 -230
rect 78023 -286 78077 -230
rect 78133 -286 78187 -230
rect 78243 -286 78297 -230
rect 78353 -277 80687 -230
rect 80743 -277 80797 -221
rect 80853 -277 80907 -221
rect 80963 -277 81017 -221
rect 81073 -277 81127 -221
rect 81183 -277 81237 -221
rect 81293 -277 81347 -221
rect 81403 -277 83528 -221
rect 83584 -277 83638 -221
rect 83694 -277 83748 -221
rect 83804 -277 83858 -221
rect 83914 -277 83968 -221
rect 84024 -277 84078 -221
rect 84134 -277 84188 -221
rect 84244 -224 89511 -221
rect 84244 -277 86316 -224
rect 78353 -280 86316 -277
rect 86372 -280 86426 -224
rect 86482 -280 86536 -224
rect 86592 -280 86646 -224
rect 86702 -280 86756 -224
rect 86812 -280 86866 -224
rect 86922 -280 86976 -224
rect 87032 -268 89511 -224
rect 89567 -268 89621 -212
rect 89677 -268 89731 -212
rect 89787 -268 89841 -212
rect 89897 -268 89951 -212
rect 90007 -268 90061 -212
rect 90117 -268 90171 -212
rect 90227 -220 128736 -212
rect 90227 -223 95994 -220
rect 90227 -268 92852 -223
rect 87032 -279 92852 -268
rect 92908 -279 92962 -223
rect 93018 -279 93072 -223
rect 93128 -279 93182 -223
rect 93238 -279 93292 -223
rect 93348 -279 93402 -223
rect 93458 -279 93512 -223
rect 93568 -276 95994 -223
rect 96050 -276 96104 -220
rect 96160 -276 96214 -220
rect 96270 -276 96324 -220
rect 96380 -276 96434 -220
rect 96490 -276 96544 -220
rect 96600 -276 96654 -220
rect 96710 -222 128736 -220
rect 96710 -276 99280 -222
rect 93568 -278 99280 -276
rect 99336 -278 99390 -222
rect 99446 -278 99500 -222
rect 99556 -278 99610 -222
rect 99666 -278 99720 -222
rect 99776 -278 99830 -222
rect 99886 -278 99940 -222
rect 99996 -229 128736 -222
rect 99996 -278 113565 -229
rect 93568 -279 113565 -278
rect 87032 -280 113565 -279
rect 78353 -285 113565 -280
rect 113621 -285 113675 -229
rect 113731 -285 113785 -229
rect 113841 -285 113895 -229
rect 113951 -285 114005 -229
rect 114061 -285 114115 -229
rect 114171 -285 114225 -229
rect 114281 -285 128736 -229
rect 78353 -286 128736 -285
rect 25425 -322 128736 -286
rect 25425 -326 89511 -322
rect 25425 -332 74565 -326
rect 25425 -336 71847 -332
rect 25425 -337 29849 -336
rect 5980 -391 29849 -337
rect 5980 -447 24709 -391
rect 24765 -447 24819 -391
rect 24875 -447 24929 -391
rect 24985 -447 25039 -391
rect 25095 -447 25149 -391
rect 25205 -447 25259 -391
rect 25315 -447 25369 -391
rect 25425 -392 29849 -391
rect 29905 -392 29959 -336
rect 30015 -392 30069 -336
rect 30125 -392 30179 -336
rect 30235 -392 30289 -336
rect 30345 -392 30399 -336
rect 30455 -392 30509 -336
rect 30565 -337 71847 -336
rect 30565 -392 69220 -337
rect 25425 -393 69220 -392
rect 69276 -393 69330 -337
rect 69386 -393 69440 -337
rect 69496 -393 69550 -337
rect 69606 -393 69660 -337
rect 69716 -393 69770 -337
rect 69826 -393 69880 -337
rect 69936 -388 71847 -337
rect 71903 -388 71957 -332
rect 72013 -388 72067 -332
rect 72123 -388 72177 -332
rect 72233 -388 72287 -332
rect 72343 -388 72397 -332
rect 72453 -388 72507 -332
rect 72563 -382 74565 -332
rect 74621 -382 74675 -326
rect 74731 -382 74785 -326
rect 74841 -382 74895 -326
rect 74951 -382 75005 -326
rect 75061 -382 75115 -326
rect 75171 -382 75225 -326
rect 75281 -331 89511 -326
rect 75281 -340 80687 -331
rect 75281 -382 77637 -340
rect 72563 -388 77637 -382
rect 69936 -393 77637 -388
rect 25425 -396 77637 -393
rect 77693 -396 77747 -340
rect 77803 -396 77857 -340
rect 77913 -396 77967 -340
rect 78023 -396 78077 -340
rect 78133 -396 78187 -340
rect 78243 -396 78297 -340
rect 78353 -387 80687 -340
rect 80743 -387 80797 -331
rect 80853 -387 80907 -331
rect 80963 -387 81017 -331
rect 81073 -387 81127 -331
rect 81183 -387 81237 -331
rect 81293 -387 81347 -331
rect 81403 -387 83528 -331
rect 83584 -387 83638 -331
rect 83694 -387 83748 -331
rect 83804 -387 83858 -331
rect 83914 -387 83968 -331
rect 84024 -387 84078 -331
rect 84134 -387 84188 -331
rect 84244 -334 89511 -331
rect 84244 -387 86316 -334
rect 78353 -390 86316 -387
rect 86372 -390 86426 -334
rect 86482 -390 86536 -334
rect 86592 -390 86646 -334
rect 86702 -390 86756 -334
rect 86812 -390 86866 -334
rect 86922 -390 86976 -334
rect 87032 -378 89511 -334
rect 89567 -378 89621 -322
rect 89677 -378 89731 -322
rect 89787 -378 89841 -322
rect 89897 -378 89951 -322
rect 90007 -378 90061 -322
rect 90117 -378 90171 -322
rect 90227 -330 128736 -322
rect 90227 -333 95994 -330
rect 90227 -378 92852 -333
rect 87032 -389 92852 -378
rect 92908 -389 92962 -333
rect 93018 -389 93072 -333
rect 93128 -389 93182 -333
rect 93238 -389 93292 -333
rect 93348 -389 93402 -333
rect 93458 -389 93512 -333
rect 93568 -386 95994 -333
rect 96050 -386 96104 -330
rect 96160 -386 96214 -330
rect 96270 -386 96324 -330
rect 96380 -386 96434 -330
rect 96490 -386 96544 -330
rect 96600 -386 96654 -330
rect 96710 -332 128736 -330
rect 96710 -386 99280 -332
rect 93568 -388 99280 -386
rect 99336 -388 99390 -332
rect 99446 -388 99500 -332
rect 99556 -388 99610 -332
rect 99666 -388 99720 -332
rect 99776 -388 99830 -332
rect 99886 -388 99940 -332
rect 99996 -339 128736 -332
rect 99996 -388 113565 -339
rect 93568 -389 113565 -388
rect 87032 -390 113565 -389
rect 78353 -395 113565 -390
rect 113621 -395 113675 -339
rect 113731 -395 113785 -339
rect 113841 -395 113895 -339
rect 113951 -395 114005 -339
rect 114061 -395 114115 -339
rect 114171 -395 114225 -339
rect 114281 -395 128736 -339
rect 78353 -396 128736 -395
rect 25425 -432 128736 -396
rect 25425 -436 89511 -432
rect 25425 -442 74565 -436
rect 25425 -447 71847 -442
rect 5980 -503 69220 -447
rect 69276 -503 69330 -447
rect 69386 -503 69440 -447
rect 69496 -503 69550 -447
rect 69606 -503 69660 -447
rect 69716 -503 69770 -447
rect 69826 -503 69880 -447
rect 69936 -498 71847 -447
rect 71903 -498 71957 -442
rect 72013 -498 72067 -442
rect 72123 -498 72177 -442
rect 72233 -498 72287 -442
rect 72343 -498 72397 -442
rect 72453 -498 72507 -442
rect 72563 -492 74565 -442
rect 74621 -492 74675 -436
rect 74731 -492 74785 -436
rect 74841 -492 74895 -436
rect 74951 -492 75005 -436
rect 75061 -492 75115 -436
rect 75171 -492 75225 -436
rect 75281 -441 89511 -436
rect 75281 -450 80687 -441
rect 75281 -492 77637 -450
rect 72563 -498 77637 -492
rect 69936 -503 77637 -498
rect 5980 -506 77637 -503
rect 77693 -506 77747 -450
rect 77803 -506 77857 -450
rect 77913 -506 77967 -450
rect 78023 -506 78077 -450
rect 78133 -506 78187 -450
rect 78243 -506 78297 -450
rect 78353 -497 80687 -450
rect 80743 -497 80797 -441
rect 80853 -497 80907 -441
rect 80963 -497 81017 -441
rect 81073 -497 81127 -441
rect 81183 -497 81237 -441
rect 81293 -497 81347 -441
rect 81403 -497 83528 -441
rect 83584 -497 83638 -441
rect 83694 -497 83748 -441
rect 83804 -497 83858 -441
rect 83914 -497 83968 -441
rect 84024 -497 84078 -441
rect 84134 -497 84188 -441
rect 84244 -444 89511 -441
rect 84244 -497 86316 -444
rect 78353 -500 86316 -497
rect 86372 -500 86426 -444
rect 86482 -500 86536 -444
rect 86592 -500 86646 -444
rect 86702 -500 86756 -444
rect 86812 -500 86866 -444
rect 86922 -500 86976 -444
rect 87032 -488 89511 -444
rect 89567 -488 89621 -432
rect 89677 -488 89731 -432
rect 89787 -488 89841 -432
rect 89897 -488 89951 -432
rect 90007 -488 90061 -432
rect 90117 -488 90171 -432
rect 90227 -440 128736 -432
rect 90227 -443 95994 -440
rect 90227 -488 92852 -443
rect 87032 -499 92852 -488
rect 92908 -499 92962 -443
rect 93018 -499 93072 -443
rect 93128 -499 93182 -443
rect 93238 -499 93292 -443
rect 93348 -499 93402 -443
rect 93458 -499 93512 -443
rect 93568 -496 95994 -443
rect 96050 -496 96104 -440
rect 96160 -496 96214 -440
rect 96270 -496 96324 -440
rect 96380 -496 96434 -440
rect 96490 -496 96544 -440
rect 96600 -496 96654 -440
rect 96710 -442 128736 -440
rect 96710 -496 99280 -442
rect 93568 -498 99280 -496
rect 99336 -498 99390 -442
rect 99446 -498 99500 -442
rect 99556 -498 99610 -442
rect 99666 -498 99720 -442
rect 99776 -498 99830 -442
rect 99886 -498 99940 -442
rect 99996 -498 128736 -442
rect 93568 -499 128736 -498
rect 87032 -500 128736 -499
rect 78353 -506 128736 -500
rect 5980 -523 128736 -506
rect 5522 -1584 5951 -1568
rect 5522 -1640 5544 -1584
rect 5600 -1640 5654 -1584
rect 5710 -1640 5764 -1584
rect 5820 -1640 5874 -1584
rect 5930 -1640 5951 -1584
rect 5522 -1694 5951 -1640
rect 5522 -1750 5544 -1694
rect 5600 -1750 5654 -1694
rect 5710 -1750 5764 -1694
rect 5820 -1750 5874 -1694
rect 5930 -1750 5951 -1694
rect 5522 -1804 5951 -1750
rect 5522 -1860 5544 -1804
rect 5600 -1860 5654 -1804
rect 5710 -1860 5764 -1804
rect 5820 -1860 5874 -1804
rect 5930 -1860 5951 -1804
rect 5522 -1914 5951 -1860
rect 5522 -1970 5544 -1914
rect 5600 -1970 5654 -1914
rect 5710 -1970 5764 -1914
rect 5820 -1970 5874 -1914
rect 5930 -1970 5951 -1914
rect 5522 -2013 5949 -1970
rect -1821 -2181 5949 -2013
rect -1821 -2237 138 -2181
rect 194 -2237 248 -2181
rect 304 -2237 358 -2181
rect 414 -2237 468 -2181
rect 524 -2237 578 -2181
rect 634 -2237 688 -2181
rect 744 -2237 798 -2181
rect 854 -2237 5949 -2181
rect -1821 -2291 5949 -2237
rect -1821 -2347 138 -2291
rect 194 -2347 248 -2291
rect 304 -2347 358 -2291
rect 414 -2347 468 -2291
rect 524 -2347 578 -2291
rect 634 -2347 688 -2291
rect 744 -2347 798 -2291
rect 854 -2347 5949 -2291
rect -1821 -2401 5949 -2347
rect -1821 -2457 138 -2401
rect 194 -2457 248 -2401
rect 304 -2457 358 -2401
rect 414 -2457 468 -2401
rect 524 -2457 578 -2401
rect 634 -2457 688 -2401
rect 744 -2457 798 -2401
rect 854 -2440 5949 -2401
rect 854 -2457 2839 -2440
rect -1821 -2511 2839 -2457
rect -1821 -2567 138 -2511
rect 194 -2567 248 -2511
rect 304 -2567 358 -2511
rect 414 -2567 468 -2511
rect 524 -2567 578 -2511
rect 634 -2567 688 -2511
rect 744 -2567 798 -2511
rect 854 -2567 2839 -2511
rect -1821 -2621 2839 -2567
rect -1821 -2677 138 -2621
rect 194 -2677 248 -2621
rect 304 -2677 358 -2621
rect 414 -2677 468 -2621
rect 524 -2677 578 -2621
rect 634 -2677 688 -2621
rect 744 -2677 798 -2621
rect 854 -2677 2839 -2621
rect -1821 -2731 2839 -2677
rect -1821 -2787 138 -2731
rect 194 -2787 248 -2731
rect 304 -2787 358 -2731
rect 414 -2787 468 -2731
rect 524 -2787 578 -2731
rect 634 -2787 688 -2731
rect 744 -2787 798 -2731
rect 854 -2787 2839 -2731
rect -1821 -2846 2839 -2787
rect 2412 -7045 2839 -2846
rect 7578 -2912 9780 -523
rect 77608 -526 78396 -523
rect 123834 -528 124100 -523
rect 124539 -528 124805 -523
rect 10763 -1128 128737 -973
rect 10763 -1184 10881 -1128
rect 10937 -1184 10991 -1128
rect 11047 -1184 11101 -1128
rect 11157 -1184 11211 -1128
rect 11267 -1184 11321 -1128
rect 11377 -1184 11431 -1128
rect 11487 -1184 11541 -1128
rect 11597 -1184 11670 -1128
rect 11726 -1184 11780 -1128
rect 11836 -1184 11890 -1128
rect 11946 -1184 12000 -1128
rect 12056 -1184 12110 -1128
rect 12166 -1184 12220 -1128
rect 12276 -1184 12330 -1128
rect 12386 -1146 128737 -1128
rect 12386 -1184 25927 -1146
rect 10763 -1202 25927 -1184
rect 25983 -1202 26037 -1146
rect 26093 -1202 26147 -1146
rect 26203 -1202 26257 -1146
rect 26313 -1202 26367 -1146
rect 26423 -1202 26477 -1146
rect 26533 -1202 26587 -1146
rect 26643 -1199 128737 -1146
rect 26643 -1202 114635 -1199
rect 10763 -1238 114635 -1202
rect 10763 -1294 10881 -1238
rect 10937 -1294 10991 -1238
rect 11047 -1294 11101 -1238
rect 11157 -1294 11211 -1238
rect 11267 -1294 11321 -1238
rect 11377 -1294 11431 -1238
rect 11487 -1294 11541 -1238
rect 11597 -1294 11670 -1238
rect 11726 -1294 11780 -1238
rect 11836 -1294 11890 -1238
rect 11946 -1294 12000 -1238
rect 12056 -1294 12110 -1238
rect 12166 -1294 12220 -1238
rect 12276 -1294 12330 -1238
rect 12386 -1255 114635 -1238
rect 114691 -1255 114745 -1199
rect 114801 -1255 114855 -1199
rect 114911 -1255 114965 -1199
rect 115021 -1255 115075 -1199
rect 115131 -1255 115185 -1199
rect 115241 -1255 115295 -1199
rect 115351 -1255 128737 -1199
rect 12386 -1256 128737 -1255
rect 12386 -1294 25927 -1256
rect 10763 -1312 25927 -1294
rect 25983 -1312 26037 -1256
rect 26093 -1312 26147 -1256
rect 26203 -1312 26257 -1256
rect 26313 -1312 26367 -1256
rect 26423 -1312 26477 -1256
rect 26533 -1312 26587 -1256
rect 26643 -1309 128737 -1256
rect 26643 -1312 114635 -1309
rect 10763 -1348 114635 -1312
rect 10763 -1404 10881 -1348
rect 10937 -1404 10991 -1348
rect 11047 -1404 11101 -1348
rect 11157 -1404 11211 -1348
rect 11267 -1404 11321 -1348
rect 11377 -1404 11431 -1348
rect 11487 -1404 11541 -1348
rect 11597 -1404 11670 -1348
rect 11726 -1404 11780 -1348
rect 11836 -1404 11890 -1348
rect 11946 -1404 12000 -1348
rect 12056 -1404 12110 -1348
rect 12166 -1404 12220 -1348
rect 12276 -1404 12330 -1348
rect 12386 -1365 114635 -1348
rect 114691 -1365 114745 -1309
rect 114801 -1365 114855 -1309
rect 114911 -1365 114965 -1309
rect 115021 -1365 115075 -1309
rect 115131 -1365 115185 -1309
rect 115241 -1365 115295 -1309
rect 115351 -1365 128737 -1309
rect 12386 -1366 128737 -1365
rect 12386 -1404 25927 -1366
rect 10763 -1422 25927 -1404
rect 25983 -1422 26037 -1366
rect 26093 -1422 26147 -1366
rect 26203 -1422 26257 -1366
rect 26313 -1422 26367 -1366
rect 26423 -1422 26477 -1366
rect 26533 -1422 26587 -1366
rect 26643 -1419 128737 -1366
rect 26643 -1422 114635 -1419
rect 10763 -1458 114635 -1422
rect 10763 -1514 10881 -1458
rect 10937 -1514 10991 -1458
rect 11047 -1514 11101 -1458
rect 11157 -1514 11211 -1458
rect 11267 -1514 11321 -1458
rect 11377 -1514 11431 -1458
rect 11487 -1514 11541 -1458
rect 11597 -1514 11670 -1458
rect 11726 -1514 11780 -1458
rect 11836 -1514 11890 -1458
rect 11946 -1514 12000 -1458
rect 12056 -1514 12110 -1458
rect 12166 -1514 12220 -1458
rect 12276 -1514 12330 -1458
rect 12386 -1475 114635 -1458
rect 114691 -1475 114745 -1419
rect 114801 -1475 114855 -1419
rect 114911 -1475 114965 -1419
rect 115021 -1475 115075 -1419
rect 115131 -1475 115185 -1419
rect 115241 -1475 115295 -1419
rect 115351 -1475 128737 -1419
rect 12386 -1476 128737 -1475
rect 12386 -1514 25927 -1476
rect 10763 -1532 25927 -1514
rect 25983 -1532 26037 -1476
rect 26093 -1532 26147 -1476
rect 26203 -1532 26257 -1476
rect 26313 -1532 26367 -1476
rect 26423 -1532 26477 -1476
rect 26533 -1532 26587 -1476
rect 26643 -1529 128737 -1476
rect 26643 -1532 114635 -1529
rect 10763 -1568 114635 -1532
rect 10763 -1624 10881 -1568
rect 10937 -1624 10991 -1568
rect 11047 -1624 11101 -1568
rect 11157 -1624 11211 -1568
rect 11267 -1624 11321 -1568
rect 11377 -1624 11431 -1568
rect 11487 -1624 11541 -1568
rect 11597 -1624 11670 -1568
rect 11726 -1624 11780 -1568
rect 11836 -1624 11890 -1568
rect 11946 -1624 12000 -1568
rect 12056 -1624 12110 -1568
rect 12166 -1624 12220 -1568
rect 12276 -1624 12330 -1568
rect 12386 -1585 114635 -1568
rect 114691 -1585 114745 -1529
rect 114801 -1585 114855 -1529
rect 114911 -1585 114965 -1529
rect 115021 -1585 115075 -1529
rect 115131 -1585 115185 -1529
rect 115241 -1585 115295 -1529
rect 115351 -1585 128737 -1529
rect 12386 -1586 128737 -1585
rect 12386 -1624 25927 -1586
rect 10763 -1642 25927 -1624
rect 25983 -1642 26037 -1586
rect 26093 -1642 26147 -1586
rect 26203 -1642 26257 -1586
rect 26313 -1642 26367 -1586
rect 26423 -1642 26477 -1586
rect 26533 -1642 26587 -1586
rect 26643 -1639 128737 -1586
rect 26643 -1642 114635 -1639
rect 10763 -1678 114635 -1642
rect 10763 -1734 10881 -1678
rect 10937 -1734 10991 -1678
rect 11047 -1734 11101 -1678
rect 11157 -1734 11211 -1678
rect 11267 -1734 11321 -1678
rect 11377 -1734 11431 -1678
rect 11487 -1734 11541 -1678
rect 11597 -1734 11670 -1678
rect 11726 -1734 11780 -1678
rect 11836 -1734 11890 -1678
rect 11946 -1734 12000 -1678
rect 12056 -1734 12110 -1678
rect 12166 -1734 12220 -1678
rect 12276 -1734 12330 -1678
rect 12386 -1695 114635 -1678
rect 114691 -1695 114745 -1639
rect 114801 -1695 114855 -1639
rect 114911 -1695 114965 -1639
rect 115021 -1695 115075 -1639
rect 115131 -1695 115185 -1639
rect 115241 -1695 115295 -1639
rect 115351 -1695 128737 -1639
rect 12386 -1696 128737 -1695
rect 12386 -1734 25927 -1696
rect 10763 -1752 25927 -1734
rect 25983 -1752 26037 -1696
rect 26093 -1752 26147 -1696
rect 26203 -1752 26257 -1696
rect 26313 -1752 26367 -1696
rect 26423 -1752 26477 -1696
rect 26533 -1752 26587 -1696
rect 26643 -1749 128737 -1696
rect 26643 -1752 114635 -1749
rect 10763 -1805 114635 -1752
rect 114691 -1805 114745 -1749
rect 114801 -1805 114855 -1749
rect 114911 -1805 114965 -1749
rect 115021 -1805 115075 -1749
rect 115131 -1805 115185 -1749
rect 115241 -1805 115295 -1749
rect 115351 -1805 128737 -1749
rect 10763 -1873 128737 -1805
rect 29765 -2220 30664 -2127
rect 29765 -2276 29884 -2220
rect 29940 -2276 29994 -2220
rect 30050 -2276 30104 -2220
rect 30160 -2276 30214 -2220
rect 30270 -2276 30324 -2220
rect 30380 -2276 30434 -2220
rect 30490 -2276 30544 -2220
rect 30600 -2276 30664 -2220
rect 29765 -2312 30664 -2276
rect 29858 -2314 30630 -2312
rect 43577 -3315 44477 -1873
rect 47339 -3376 48239 -1873
rect 50279 -3193 51179 -1873
rect 53483 -3298 54383 -1873
rect 56765 -3376 57665 -1873
rect 59180 -3271 60080 -1873
rect 61307 -3376 62207 -1873
rect 63408 -3219 64308 -1873
rect 113520 -2289 114315 -2253
rect 113520 -2345 113560 -2289
rect 113616 -2345 113670 -2289
rect 113726 -2345 113780 -2289
rect 113836 -2345 113890 -2289
rect 113946 -2345 114000 -2289
rect 114056 -2345 114110 -2289
rect 114166 -2345 114220 -2289
rect 114276 -2324 114315 -2289
rect 114276 -2345 128946 -2324
rect 113520 -2399 128946 -2345
rect 113520 -2455 113560 -2399
rect 113616 -2455 113670 -2399
rect 113726 -2455 113780 -2399
rect 113836 -2455 113890 -2399
rect 113946 -2455 114000 -2399
rect 114056 -2455 114110 -2399
rect 114166 -2455 114220 -2399
rect 114276 -2455 128946 -2399
rect 113520 -2509 128946 -2455
rect 113520 -2565 113560 -2509
rect 113616 -2565 113670 -2509
rect 113726 -2565 113780 -2509
rect 113836 -2565 113890 -2509
rect 113946 -2565 114000 -2509
rect 114056 -2565 114110 -2509
rect 114166 -2565 114220 -2509
rect 114276 -2565 128946 -2509
rect 113520 -2619 128946 -2565
rect 113520 -2675 113560 -2619
rect 113616 -2675 113670 -2619
rect 113726 -2675 113780 -2619
rect 113836 -2675 113890 -2619
rect 113946 -2675 114000 -2619
rect 114056 -2675 114110 -2619
rect 114166 -2675 114220 -2619
rect 114276 -2675 128946 -2619
rect 113520 -2729 128946 -2675
rect 113520 -2785 113560 -2729
rect 113616 -2785 113670 -2729
rect 113726 -2785 113780 -2729
rect 113836 -2785 113890 -2729
rect 113946 -2785 114000 -2729
rect 114056 -2785 114110 -2729
rect 114166 -2785 114220 -2729
rect 114276 -2785 128946 -2729
rect 113520 -2803 128946 -2785
rect 113520 -2839 114315 -2803
rect 113520 -2895 113560 -2839
rect 113616 -2895 113670 -2839
rect 113726 -2895 113780 -2839
rect 113836 -2895 113890 -2839
rect 113946 -2895 114000 -2839
rect 114056 -2895 114110 -2839
rect 114166 -2895 114220 -2839
rect 114276 -2895 114315 -2839
rect 113520 -2935 114315 -2895
rect 69221 -3325 70009 -3307
rect 69221 -3381 69250 -3325
rect 69306 -3381 69360 -3325
rect 69416 -3381 69470 -3325
rect 69526 -3381 69580 -3325
rect 69636 -3381 69690 -3325
rect 69746 -3381 69800 -3325
rect 69856 -3381 69910 -3325
rect 69966 -3381 70009 -3325
rect 89492 -3329 90280 -3311
rect 80670 -3356 81458 -3338
rect 69221 -3435 70009 -3381
rect 69221 -3491 69250 -3435
rect 69306 -3491 69360 -3435
rect 69416 -3491 69470 -3435
rect 69526 -3491 69580 -3435
rect 69636 -3491 69690 -3435
rect 69746 -3491 69800 -3435
rect 69856 -3491 69910 -3435
rect 69966 -3491 70009 -3435
rect 69221 -3545 70009 -3491
rect 69221 -3601 69250 -3545
rect 69306 -3601 69360 -3545
rect 69416 -3601 69470 -3545
rect 69526 -3601 69580 -3545
rect 69636 -3601 69690 -3545
rect 69746 -3601 69800 -3545
rect 69856 -3601 69910 -3545
rect 69966 -3601 70009 -3545
rect 69221 -3655 70009 -3601
rect 69221 -3711 69250 -3655
rect 69306 -3711 69360 -3655
rect 69416 -3711 69470 -3655
rect 69526 -3711 69580 -3655
rect 69636 -3711 69690 -3655
rect 69746 -3711 69800 -3655
rect 69856 -3711 69910 -3655
rect 69966 -3711 70009 -3655
rect 69221 -3765 70009 -3711
rect 69221 -3821 69250 -3765
rect 69306 -3821 69360 -3765
rect 69416 -3821 69470 -3765
rect 69526 -3821 69580 -3765
rect 69636 -3821 69690 -3765
rect 69746 -3821 69800 -3765
rect 69856 -3821 69910 -3765
rect 69966 -3821 70009 -3765
rect 69221 -3875 70009 -3821
rect 69221 -3931 69250 -3875
rect 69306 -3931 69360 -3875
rect 69416 -3931 69470 -3875
rect 69526 -3931 69580 -3875
rect 69636 -3931 69690 -3875
rect 69746 -3931 69800 -3875
rect 69856 -3931 69910 -3875
rect 69966 -3931 70009 -3875
rect 69221 -3951 70009 -3931
rect 71834 -3388 72622 -3370
rect 71834 -3444 71863 -3388
rect 71919 -3444 71973 -3388
rect 72029 -3444 72083 -3388
rect 72139 -3444 72193 -3388
rect 72249 -3444 72303 -3388
rect 72359 -3444 72413 -3388
rect 72469 -3444 72523 -3388
rect 72579 -3444 72622 -3388
rect 77616 -3384 78404 -3366
rect 71834 -3498 72622 -3444
rect 71834 -3554 71863 -3498
rect 71919 -3554 71973 -3498
rect 72029 -3554 72083 -3498
rect 72139 -3554 72193 -3498
rect 72249 -3554 72303 -3498
rect 72359 -3554 72413 -3498
rect 72469 -3554 72523 -3498
rect 72579 -3554 72622 -3498
rect 71834 -3608 72622 -3554
rect 71834 -3664 71863 -3608
rect 71919 -3664 71973 -3608
rect 72029 -3664 72083 -3608
rect 72139 -3664 72193 -3608
rect 72249 -3664 72303 -3608
rect 72359 -3664 72413 -3608
rect 72469 -3664 72523 -3608
rect 72579 -3664 72622 -3608
rect 71834 -3718 72622 -3664
rect 71834 -3774 71863 -3718
rect 71919 -3774 71973 -3718
rect 72029 -3774 72083 -3718
rect 72139 -3774 72193 -3718
rect 72249 -3774 72303 -3718
rect 72359 -3774 72413 -3718
rect 72469 -3774 72523 -3718
rect 72579 -3774 72622 -3718
rect 71834 -3828 72622 -3774
rect 71834 -3884 71863 -3828
rect 71919 -3884 71973 -3828
rect 72029 -3884 72083 -3828
rect 72139 -3884 72193 -3828
rect 72249 -3884 72303 -3828
rect 72359 -3884 72413 -3828
rect 72469 -3884 72523 -3828
rect 72579 -3884 72622 -3828
rect 71834 -3938 72622 -3884
rect 71834 -3994 71863 -3938
rect 71919 -3994 71973 -3938
rect 72029 -3994 72083 -3938
rect 72139 -3994 72193 -3938
rect 72249 -3994 72303 -3938
rect 72359 -3994 72413 -3938
rect 72469 -3994 72523 -3938
rect 72579 -3994 72622 -3938
rect 71834 -4014 72622 -3994
rect 74548 -3410 75336 -3392
rect 74548 -3466 74577 -3410
rect 74633 -3466 74687 -3410
rect 74743 -3466 74797 -3410
rect 74853 -3466 74907 -3410
rect 74963 -3466 75017 -3410
rect 75073 -3466 75127 -3410
rect 75183 -3466 75237 -3410
rect 75293 -3466 75336 -3410
rect 74548 -3520 75336 -3466
rect 74548 -3576 74577 -3520
rect 74633 -3576 74687 -3520
rect 74743 -3576 74797 -3520
rect 74853 -3576 74907 -3520
rect 74963 -3576 75017 -3520
rect 75073 -3576 75127 -3520
rect 75183 -3576 75237 -3520
rect 75293 -3576 75336 -3520
rect 74548 -3630 75336 -3576
rect 74548 -3686 74577 -3630
rect 74633 -3686 74687 -3630
rect 74743 -3686 74797 -3630
rect 74853 -3686 74907 -3630
rect 74963 -3686 75017 -3630
rect 75073 -3686 75127 -3630
rect 75183 -3686 75237 -3630
rect 75293 -3686 75336 -3630
rect 74548 -3740 75336 -3686
rect 74548 -3796 74577 -3740
rect 74633 -3796 74687 -3740
rect 74743 -3796 74797 -3740
rect 74853 -3796 74907 -3740
rect 74963 -3796 75017 -3740
rect 75073 -3796 75127 -3740
rect 75183 -3796 75237 -3740
rect 75293 -3796 75336 -3740
rect 74548 -3850 75336 -3796
rect 74548 -3906 74577 -3850
rect 74633 -3906 74687 -3850
rect 74743 -3906 74797 -3850
rect 74853 -3906 74907 -3850
rect 74963 -3906 75017 -3850
rect 75073 -3906 75127 -3850
rect 75183 -3906 75237 -3850
rect 75293 -3906 75336 -3850
rect 74548 -3960 75336 -3906
rect 74548 -4016 74577 -3960
rect 74633 -4016 74687 -3960
rect 74743 -4016 74797 -3960
rect 74853 -4016 74907 -3960
rect 74963 -4016 75017 -3960
rect 75073 -4016 75127 -3960
rect 75183 -4016 75237 -3960
rect 75293 -4016 75336 -3960
rect 77616 -3440 77645 -3384
rect 77701 -3440 77755 -3384
rect 77811 -3440 77865 -3384
rect 77921 -3440 77975 -3384
rect 78031 -3440 78085 -3384
rect 78141 -3440 78195 -3384
rect 78251 -3440 78305 -3384
rect 78361 -3440 78404 -3384
rect 77616 -3494 78404 -3440
rect 77616 -3550 77645 -3494
rect 77701 -3550 77755 -3494
rect 77811 -3550 77865 -3494
rect 77921 -3550 77975 -3494
rect 78031 -3550 78085 -3494
rect 78141 -3550 78195 -3494
rect 78251 -3550 78305 -3494
rect 78361 -3550 78404 -3494
rect 77616 -3604 78404 -3550
rect 77616 -3660 77645 -3604
rect 77701 -3660 77755 -3604
rect 77811 -3660 77865 -3604
rect 77921 -3660 77975 -3604
rect 78031 -3660 78085 -3604
rect 78141 -3660 78195 -3604
rect 78251 -3660 78305 -3604
rect 78361 -3660 78404 -3604
rect 77616 -3714 78404 -3660
rect 77616 -3770 77645 -3714
rect 77701 -3770 77755 -3714
rect 77811 -3770 77865 -3714
rect 77921 -3770 77975 -3714
rect 78031 -3770 78085 -3714
rect 78141 -3770 78195 -3714
rect 78251 -3770 78305 -3714
rect 78361 -3770 78404 -3714
rect 77616 -3824 78404 -3770
rect 77616 -3880 77645 -3824
rect 77701 -3880 77755 -3824
rect 77811 -3880 77865 -3824
rect 77921 -3880 77975 -3824
rect 78031 -3880 78085 -3824
rect 78141 -3880 78195 -3824
rect 78251 -3880 78305 -3824
rect 78361 -3880 78404 -3824
rect 77616 -3934 78404 -3880
rect 77616 -3990 77645 -3934
rect 77701 -3990 77755 -3934
rect 77811 -3990 77865 -3934
rect 77921 -3990 77975 -3934
rect 78031 -3990 78085 -3934
rect 78141 -3990 78195 -3934
rect 78251 -3990 78305 -3934
rect 78361 -3990 78404 -3934
rect 80670 -3412 80699 -3356
rect 80755 -3412 80809 -3356
rect 80865 -3412 80919 -3356
rect 80975 -3412 81029 -3356
rect 81085 -3412 81139 -3356
rect 81195 -3412 81249 -3356
rect 81305 -3412 81359 -3356
rect 81415 -3412 81458 -3356
rect 80670 -3466 81458 -3412
rect 80670 -3522 80699 -3466
rect 80755 -3522 80809 -3466
rect 80865 -3522 80919 -3466
rect 80975 -3522 81029 -3466
rect 81085 -3522 81139 -3466
rect 81195 -3522 81249 -3466
rect 81305 -3522 81359 -3466
rect 81415 -3522 81458 -3466
rect 80670 -3576 81458 -3522
rect 80670 -3632 80699 -3576
rect 80755 -3632 80809 -3576
rect 80865 -3632 80919 -3576
rect 80975 -3632 81029 -3576
rect 81085 -3632 81139 -3576
rect 81195 -3632 81249 -3576
rect 81305 -3632 81359 -3576
rect 81415 -3632 81458 -3576
rect 80670 -3686 81458 -3632
rect 80670 -3742 80699 -3686
rect 80755 -3742 80809 -3686
rect 80865 -3742 80919 -3686
rect 80975 -3742 81029 -3686
rect 81085 -3742 81139 -3686
rect 81195 -3742 81249 -3686
rect 81305 -3742 81359 -3686
rect 81415 -3742 81458 -3686
rect 80670 -3796 81458 -3742
rect 80670 -3852 80699 -3796
rect 80755 -3852 80809 -3796
rect 80865 -3852 80919 -3796
rect 80975 -3852 81029 -3796
rect 81085 -3852 81139 -3796
rect 81195 -3852 81249 -3796
rect 81305 -3852 81359 -3796
rect 81415 -3852 81458 -3796
rect 80670 -3906 81458 -3852
rect 80670 -3962 80699 -3906
rect 80755 -3962 80809 -3906
rect 80865 -3962 80919 -3906
rect 80975 -3962 81029 -3906
rect 81085 -3962 81139 -3906
rect 81195 -3962 81249 -3906
rect 81305 -3962 81359 -3906
rect 81415 -3962 81458 -3906
rect 80670 -3982 81458 -3962
rect 83523 -3352 84311 -3334
rect 83523 -3408 83552 -3352
rect 83608 -3408 83662 -3352
rect 83718 -3408 83772 -3352
rect 83828 -3408 83882 -3352
rect 83938 -3408 83992 -3352
rect 84048 -3408 84102 -3352
rect 84158 -3408 84212 -3352
rect 84268 -3408 84311 -3352
rect 83523 -3462 84311 -3408
rect 83523 -3518 83552 -3462
rect 83608 -3518 83662 -3462
rect 83718 -3518 83772 -3462
rect 83828 -3518 83882 -3462
rect 83938 -3518 83992 -3462
rect 84048 -3518 84102 -3462
rect 84158 -3518 84212 -3462
rect 84268 -3518 84311 -3462
rect 83523 -3572 84311 -3518
rect 83523 -3628 83552 -3572
rect 83608 -3628 83662 -3572
rect 83718 -3628 83772 -3572
rect 83828 -3628 83882 -3572
rect 83938 -3628 83992 -3572
rect 84048 -3628 84102 -3572
rect 84158 -3628 84212 -3572
rect 84268 -3628 84311 -3572
rect 83523 -3682 84311 -3628
rect 83523 -3738 83552 -3682
rect 83608 -3738 83662 -3682
rect 83718 -3738 83772 -3682
rect 83828 -3738 83882 -3682
rect 83938 -3738 83992 -3682
rect 84048 -3738 84102 -3682
rect 84158 -3738 84212 -3682
rect 84268 -3738 84311 -3682
rect 83523 -3792 84311 -3738
rect 83523 -3848 83552 -3792
rect 83608 -3848 83662 -3792
rect 83718 -3848 83772 -3792
rect 83828 -3848 83882 -3792
rect 83938 -3848 83992 -3792
rect 84048 -3848 84102 -3792
rect 84158 -3848 84212 -3792
rect 84268 -3848 84311 -3792
rect 83523 -3902 84311 -3848
rect 86310 -3376 87098 -3358
rect 86310 -3432 86339 -3376
rect 86395 -3432 86449 -3376
rect 86505 -3432 86559 -3376
rect 86615 -3432 86669 -3376
rect 86725 -3432 86779 -3376
rect 86835 -3432 86889 -3376
rect 86945 -3432 86999 -3376
rect 87055 -3432 87098 -3376
rect 86310 -3486 87098 -3432
rect 86310 -3542 86339 -3486
rect 86395 -3542 86449 -3486
rect 86505 -3542 86559 -3486
rect 86615 -3542 86669 -3486
rect 86725 -3542 86779 -3486
rect 86835 -3542 86889 -3486
rect 86945 -3542 86999 -3486
rect 87055 -3542 87098 -3486
rect 86310 -3596 87098 -3542
rect 86310 -3652 86339 -3596
rect 86395 -3652 86449 -3596
rect 86505 -3652 86559 -3596
rect 86615 -3652 86669 -3596
rect 86725 -3652 86779 -3596
rect 86835 -3652 86889 -3596
rect 86945 -3652 86999 -3596
rect 87055 -3652 87098 -3596
rect 86310 -3706 87098 -3652
rect 86310 -3762 86339 -3706
rect 86395 -3762 86449 -3706
rect 86505 -3762 86559 -3706
rect 86615 -3762 86669 -3706
rect 86725 -3762 86779 -3706
rect 86835 -3762 86889 -3706
rect 86945 -3762 86999 -3706
rect 87055 -3762 87098 -3706
rect 86310 -3816 87098 -3762
rect 86310 -3872 86339 -3816
rect 86395 -3872 86449 -3816
rect 86505 -3872 86559 -3816
rect 86615 -3872 86669 -3816
rect 86725 -3872 86779 -3816
rect 86835 -3872 86889 -3816
rect 86945 -3872 86999 -3816
rect 87055 -3872 87098 -3816
rect 86310 -3877 87098 -3872
rect 83523 -3958 83552 -3902
rect 83608 -3958 83662 -3902
rect 83718 -3958 83772 -3902
rect 83828 -3958 83882 -3902
rect 83938 -3958 83992 -3902
rect 84048 -3958 84102 -3902
rect 84158 -3958 84212 -3902
rect 84268 -3958 84311 -3902
rect 83523 -3978 84311 -3958
rect 86256 -3926 87098 -3877
rect 86256 -3982 86339 -3926
rect 86395 -3982 86449 -3926
rect 86505 -3982 86559 -3926
rect 86615 -3982 86669 -3926
rect 86725 -3982 86779 -3926
rect 86835 -3982 86889 -3926
rect 86945 -3982 86999 -3926
rect 87055 -3982 87098 -3926
rect 89492 -3385 89521 -3329
rect 89577 -3385 89631 -3329
rect 89687 -3385 89741 -3329
rect 89797 -3385 89851 -3329
rect 89907 -3385 89961 -3329
rect 90017 -3385 90071 -3329
rect 90127 -3385 90181 -3329
rect 90237 -3385 90280 -3329
rect 89492 -3439 90280 -3385
rect 89492 -3495 89521 -3439
rect 89577 -3495 89631 -3439
rect 89687 -3495 89741 -3439
rect 89797 -3495 89851 -3439
rect 89907 -3495 89961 -3439
rect 90017 -3495 90071 -3439
rect 90127 -3495 90181 -3439
rect 90237 -3495 90280 -3439
rect 89492 -3549 90280 -3495
rect 89492 -3605 89521 -3549
rect 89577 -3605 89631 -3549
rect 89687 -3605 89741 -3549
rect 89797 -3605 89851 -3549
rect 89907 -3605 89961 -3549
rect 90017 -3605 90071 -3549
rect 90127 -3605 90181 -3549
rect 90237 -3605 90280 -3549
rect 89492 -3659 90280 -3605
rect 89492 -3715 89521 -3659
rect 89577 -3715 89631 -3659
rect 89687 -3715 89741 -3659
rect 89797 -3715 89851 -3659
rect 89907 -3715 89961 -3659
rect 90017 -3715 90071 -3659
rect 90127 -3715 90181 -3659
rect 90237 -3715 90280 -3659
rect 89492 -3769 90280 -3715
rect 89492 -3825 89521 -3769
rect 89577 -3825 89631 -3769
rect 89687 -3825 89741 -3769
rect 89797 -3825 89851 -3769
rect 89907 -3825 89961 -3769
rect 90017 -3825 90071 -3769
rect 90127 -3825 90181 -3769
rect 90237 -3825 90280 -3769
rect 89492 -3879 90280 -3825
rect 89492 -3935 89521 -3879
rect 89577 -3935 89631 -3879
rect 89687 -3935 89741 -3879
rect 89797 -3935 89851 -3879
rect 89907 -3935 89961 -3879
rect 90017 -3935 90071 -3879
rect 90127 -3935 90181 -3879
rect 90237 -3935 90280 -3879
rect 89492 -3955 90280 -3935
rect 92836 -3354 93624 -3336
rect 92836 -3410 92865 -3354
rect 92921 -3410 92975 -3354
rect 93031 -3410 93085 -3354
rect 93141 -3410 93195 -3354
rect 93251 -3410 93305 -3354
rect 93361 -3410 93415 -3354
rect 93471 -3410 93525 -3354
rect 93581 -3410 93624 -3354
rect 92836 -3464 93624 -3410
rect 92836 -3520 92865 -3464
rect 92921 -3520 92975 -3464
rect 93031 -3520 93085 -3464
rect 93141 -3520 93195 -3464
rect 93251 -3520 93305 -3464
rect 93361 -3520 93415 -3464
rect 93471 -3520 93525 -3464
rect 93581 -3520 93624 -3464
rect 92836 -3574 93624 -3520
rect 92836 -3630 92865 -3574
rect 92921 -3630 92975 -3574
rect 93031 -3630 93085 -3574
rect 93141 -3630 93195 -3574
rect 93251 -3630 93305 -3574
rect 93361 -3630 93415 -3574
rect 93471 -3630 93525 -3574
rect 93581 -3630 93624 -3574
rect 92836 -3684 93624 -3630
rect 92836 -3740 92865 -3684
rect 92921 -3740 92975 -3684
rect 93031 -3740 93085 -3684
rect 93141 -3740 93195 -3684
rect 93251 -3740 93305 -3684
rect 93361 -3740 93415 -3684
rect 93471 -3740 93525 -3684
rect 93581 -3740 93624 -3684
rect 92836 -3794 93624 -3740
rect 92836 -3850 92865 -3794
rect 92921 -3850 92975 -3794
rect 93031 -3850 93085 -3794
rect 93141 -3850 93195 -3794
rect 93251 -3850 93305 -3794
rect 93361 -3850 93415 -3794
rect 93471 -3850 93525 -3794
rect 93581 -3850 93624 -3794
rect 92836 -3904 93624 -3850
rect 95969 -3384 96757 -3366
rect 95969 -3440 95998 -3384
rect 96054 -3440 96108 -3384
rect 96164 -3440 96218 -3384
rect 96274 -3440 96328 -3384
rect 96384 -3440 96438 -3384
rect 96494 -3440 96548 -3384
rect 96604 -3440 96658 -3384
rect 96714 -3440 96757 -3384
rect 95969 -3494 96757 -3440
rect 95969 -3550 95998 -3494
rect 96054 -3550 96108 -3494
rect 96164 -3550 96218 -3494
rect 96274 -3550 96328 -3494
rect 96384 -3550 96438 -3494
rect 96494 -3550 96548 -3494
rect 96604 -3550 96658 -3494
rect 96714 -3550 96757 -3494
rect 95969 -3604 96757 -3550
rect 95969 -3660 95998 -3604
rect 96054 -3660 96108 -3604
rect 96164 -3660 96218 -3604
rect 96274 -3660 96328 -3604
rect 96384 -3660 96438 -3604
rect 96494 -3660 96548 -3604
rect 96604 -3660 96658 -3604
rect 96714 -3660 96757 -3604
rect 95969 -3714 96757 -3660
rect 95969 -3770 95998 -3714
rect 96054 -3770 96108 -3714
rect 96164 -3770 96218 -3714
rect 96274 -3770 96328 -3714
rect 96384 -3770 96438 -3714
rect 96494 -3770 96548 -3714
rect 96604 -3770 96658 -3714
rect 96714 -3770 96757 -3714
rect 95969 -3824 96757 -3770
rect 95969 -3854 95998 -3824
rect 92836 -3960 92865 -3904
rect 92921 -3960 92975 -3904
rect 93031 -3960 93085 -3904
rect 93141 -3960 93195 -3904
rect 93251 -3960 93305 -3904
rect 93361 -3960 93415 -3904
rect 93471 -3960 93525 -3904
rect 93581 -3960 93624 -3904
rect 92836 -3980 93624 -3960
rect 95924 -3880 95998 -3854
rect 96054 -3880 96108 -3824
rect 96164 -3880 96218 -3824
rect 96274 -3880 96328 -3824
rect 96384 -3880 96438 -3824
rect 96494 -3880 96548 -3824
rect 96604 -3880 96658 -3824
rect 96714 -3880 96757 -3824
rect 95924 -3934 96757 -3880
rect 95924 -3980 95998 -3934
rect 77616 -4010 78404 -3990
rect 86256 -4002 87098 -3982
rect 95925 -3990 95998 -3980
rect 96054 -3990 96108 -3934
rect 96164 -3990 96218 -3934
rect 96274 -3990 96328 -3934
rect 96384 -3990 96438 -3934
rect 96494 -3990 96548 -3934
rect 96604 -3990 96658 -3934
rect 96714 -3990 96757 -3934
rect 86256 -4003 86336 -4002
rect 95925 -4010 96757 -3990
rect 99247 -3418 100035 -3400
rect 99247 -3474 99276 -3418
rect 99332 -3474 99386 -3418
rect 99442 -3474 99496 -3418
rect 99552 -3474 99606 -3418
rect 99662 -3474 99716 -3418
rect 99772 -3474 99826 -3418
rect 99882 -3474 99936 -3418
rect 99992 -3474 100035 -3418
rect 99247 -3528 100035 -3474
rect 99247 -3584 99276 -3528
rect 99332 -3584 99386 -3528
rect 99442 -3584 99496 -3528
rect 99552 -3584 99606 -3528
rect 99662 -3584 99716 -3528
rect 99772 -3584 99826 -3528
rect 99882 -3584 99936 -3528
rect 99992 -3584 100035 -3528
rect 99247 -3638 100035 -3584
rect 99247 -3694 99276 -3638
rect 99332 -3694 99386 -3638
rect 99442 -3694 99496 -3638
rect 99552 -3694 99606 -3638
rect 99662 -3694 99716 -3638
rect 99772 -3694 99826 -3638
rect 99882 -3694 99936 -3638
rect 99992 -3694 100035 -3638
rect 99247 -3748 100035 -3694
rect 99247 -3804 99276 -3748
rect 99332 -3804 99386 -3748
rect 99442 -3804 99496 -3748
rect 99552 -3804 99606 -3748
rect 99662 -3804 99716 -3748
rect 99772 -3804 99826 -3748
rect 99882 -3804 99936 -3748
rect 99992 -3804 100035 -3748
rect 99247 -3858 100035 -3804
rect 99247 -3914 99276 -3858
rect 99332 -3914 99386 -3858
rect 99442 -3914 99496 -3858
rect 99552 -3914 99606 -3858
rect 99662 -3914 99716 -3858
rect 99772 -3914 99826 -3858
rect 99882 -3914 99936 -3858
rect 99992 -3914 100035 -3858
rect 99247 -3968 100035 -3914
rect 74548 -4036 75336 -4016
rect 99247 -4024 99276 -3968
rect 99332 -4024 99386 -3968
rect 99442 -4024 99496 -3968
rect 99552 -4024 99606 -3968
rect 99662 -4024 99716 -3968
rect 99772 -4024 99826 -3968
rect 99882 -4024 99936 -3968
rect 99992 -4024 100035 -3968
rect 99247 -4044 100035 -4024
rect 30146 -4151 30811 -4126
rect 30146 -4207 30166 -4151
rect 30222 -4207 30276 -4151
rect 30332 -4207 30386 -4151
rect 30442 -4207 30496 -4151
rect 30552 -4207 30606 -4151
rect 30662 -4207 30716 -4151
rect 30772 -4207 30811 -4151
rect 30146 -4261 30811 -4207
rect 30146 -4317 30166 -4261
rect 30222 -4317 30276 -4261
rect 30332 -4317 30386 -4261
rect 30442 -4317 30496 -4261
rect 30552 -4317 30606 -4261
rect 30662 -4317 30716 -4261
rect 30772 -4317 30811 -4261
rect 30146 -4376 30811 -4317
rect 129124 -4373 131075 -3824
rect 31187 -4612 31622 -4590
rect 31187 -4668 31209 -4612
rect 31265 -4668 31319 -4612
rect 31375 -4668 31429 -4612
rect 31485 -4668 31539 -4612
rect 31595 -4668 31622 -4612
rect 31187 -4687 31622 -4668
rect 116615 -5220 116780 -5212
rect 116615 -5276 116662 -5220
rect 116718 -5276 116780 -5220
rect 129129 -5223 131080 -4674
rect 116615 -5330 116780 -5276
rect 116615 -5386 116662 -5330
rect 116718 -5386 116780 -5330
rect 116615 -5440 116780 -5386
rect 116615 -5496 116662 -5440
rect 116718 -5496 116780 -5440
rect 116615 -5550 116780 -5496
rect 116615 -5606 116662 -5550
rect 116718 -5606 116780 -5550
rect 116615 -5660 116780 -5606
rect 116615 -5716 116662 -5660
rect 116718 -5716 116780 -5660
rect 116615 -5770 116780 -5716
rect 116615 -5826 116662 -5770
rect 116718 -5826 116780 -5770
rect 116615 -5863 116780 -5826
rect 129129 -6278 131080 -5981
rect 129128 -6454 131080 -6278
rect 129129 -6530 131080 -6454
rect 116619 -6615 116784 -6607
rect 116619 -6671 116666 -6615
rect 116722 -6671 116784 -6615
rect 116619 -6725 116784 -6671
rect 116619 -6781 116666 -6725
rect 116722 -6781 116784 -6725
rect 116619 -6835 116784 -6781
rect 116619 -6891 116666 -6835
rect 116722 -6891 116784 -6835
rect 116619 -6945 116784 -6891
rect 116619 -7001 116666 -6945
rect 116722 -7001 116784 -6945
rect 2412 -7220 3204 -7045
rect 116619 -7055 116784 -7001
rect 116619 -7111 116666 -7055
rect 116722 -7111 116784 -7055
rect 116619 -7165 116784 -7111
rect 116619 -7221 116666 -7165
rect 116722 -7221 116784 -7165
rect 116619 -7258 116784 -7221
rect 129124 -7239 131075 -6690
rect 109049 -7895 116267 -7875
rect 109049 -7951 109078 -7895
rect 109134 -7951 109188 -7895
rect 109244 -7951 109298 -7895
rect 109354 -7951 109408 -7895
rect 109464 -7951 109518 -7895
rect 109574 -7951 109628 -7895
rect 109684 -7951 109738 -7895
rect 109794 -7951 116267 -7895
rect 109049 -8005 116267 -7951
rect 109049 -8061 109078 -8005
rect 109134 -8061 109188 -8005
rect 109244 -8061 109298 -8005
rect 109354 -8061 109408 -8005
rect 109464 -8061 109518 -8005
rect 109574 -8061 109628 -8005
rect 109684 -8061 109738 -8005
rect 109794 -8061 116267 -8005
rect 109049 -8115 116267 -8061
rect 109049 -8171 109078 -8115
rect 109134 -8171 109188 -8115
rect 109244 -8171 109298 -8115
rect 109354 -8171 109408 -8115
rect 109464 -8171 109518 -8115
rect 109574 -8171 109628 -8115
rect 109684 -8171 109738 -8115
rect 109794 -8171 116267 -8115
rect 109049 -8225 116267 -8171
rect 109049 -8281 109078 -8225
rect 109134 -8281 109188 -8225
rect 109244 -8281 109298 -8225
rect 109354 -8281 109408 -8225
rect 109464 -8281 109518 -8225
rect 109574 -8281 109628 -8225
rect 109684 -8281 109738 -8225
rect 109794 -8281 116267 -8225
rect 109049 -8335 116267 -8281
rect 109049 -8391 109078 -8335
rect 109134 -8391 109188 -8335
rect 109244 -8391 109298 -8335
rect 109354 -8391 109408 -8335
rect 109464 -8391 109518 -8335
rect 109574 -8391 109628 -8335
rect 109684 -8391 109738 -8335
rect 109794 -8391 116267 -8335
rect 109049 -8445 116267 -8391
rect 109049 -8501 109078 -8445
rect 109134 -8501 109188 -8445
rect 109244 -8501 109298 -8445
rect 109354 -8501 109408 -8445
rect 109464 -8501 109518 -8445
rect 109574 -8501 109628 -8445
rect 109684 -8501 109738 -8445
rect 109794 -8501 116267 -8445
rect 109049 -8555 116267 -8501
rect 109049 -8611 109078 -8555
rect 109134 -8611 109188 -8555
rect 109244 -8611 109298 -8555
rect 109354 -8611 109408 -8555
rect 109464 -8611 109518 -8555
rect 109574 -8611 109628 -8555
rect 109684 -8611 109738 -8555
rect 109794 -8611 116267 -8555
rect 109049 -8665 116267 -8611
rect 109049 -8721 109078 -8665
rect 109134 -8721 109188 -8665
rect 109244 -8721 109298 -8665
rect 109354 -8721 109408 -8665
rect 109464 -8721 109518 -8665
rect 109574 -8721 109628 -8665
rect 109684 -8721 109738 -8665
rect 109794 -8721 116267 -8665
rect 109049 -8741 116267 -8721
rect 116617 -8446 116782 -8438
rect 116617 -8502 116664 -8446
rect 116720 -8502 116782 -8446
rect 116617 -8556 116782 -8502
rect 116617 -8612 116664 -8556
rect 116720 -8612 116782 -8556
rect 116617 -8666 116782 -8612
rect 116617 -8722 116664 -8666
rect 116720 -8722 116782 -8666
rect 116617 -8776 116782 -8722
rect 116617 -8832 116664 -8776
rect 116720 -8832 116782 -8776
rect 116617 -8886 116782 -8832
rect 116617 -8942 116664 -8886
rect 116720 -8942 116782 -8886
rect 116617 -8996 116782 -8942
rect 116617 -9052 116664 -8996
rect 116720 -9052 116782 -8996
rect 129151 -9038 131102 -8489
rect 116617 -9089 116782 -9052
rect 129133 -9735 131084 -9186
rect 116618 -9764 116783 -9756
rect 116618 -9820 116665 -9764
rect 116721 -9820 116783 -9764
rect 116618 -9874 116783 -9820
rect 116618 -9930 116665 -9874
rect 116721 -9930 116783 -9874
rect 116618 -9984 116783 -9930
rect 116618 -10040 116665 -9984
rect 116721 -10040 116783 -9984
rect 116618 -10094 116783 -10040
rect 116618 -10150 116665 -10094
rect 116721 -10150 116783 -10094
rect 116618 -10204 116783 -10150
rect 116618 -10260 116665 -10204
rect 116721 -10260 116783 -10204
rect 116618 -10314 116783 -10260
rect 116618 -10370 116665 -10314
rect 116721 -10370 116783 -10314
rect 116618 -10407 116783 -10370
rect 129189 -11215 131140 -10666
rect 129075 -11992 131026 -11443
rect 119087 -13006 126960 -12972
rect 113504 -13207 126960 -13006
rect 113504 -13263 113550 -13207
rect 113606 -13263 113660 -13207
rect 113716 -13263 113770 -13207
rect 113826 -13263 113880 -13207
rect 113936 -13263 113990 -13207
rect 114046 -13263 114100 -13207
rect 114156 -13263 114210 -13207
rect 114266 -13263 126960 -13207
rect 113504 -13317 126960 -13263
rect 113504 -13373 113550 -13317
rect 113606 -13373 113660 -13317
rect 113716 -13373 113770 -13317
rect 113826 -13373 113880 -13317
rect 113936 -13373 113990 -13317
rect 114046 -13373 114100 -13317
rect 114156 -13373 114210 -13317
rect 114266 -13373 126960 -13317
rect 113504 -13427 126960 -13373
rect 113504 -13483 113550 -13427
rect 113606 -13483 113660 -13427
rect 113716 -13483 113770 -13427
rect 113826 -13483 113880 -13427
rect 113936 -13483 113990 -13427
rect 114046 -13483 114100 -13427
rect 114156 -13483 114210 -13427
rect 114266 -13483 126960 -13427
rect 113504 -13537 126960 -13483
rect 29479 -13656 30536 -13568
rect 29479 -13664 30193 -13656
rect 29479 -13720 29533 -13664
rect 29589 -13720 29643 -13664
rect 29699 -13720 29753 -13664
rect 29809 -13720 29863 -13664
rect 29919 -13720 29973 -13664
rect 30029 -13720 30083 -13664
rect 30139 -13712 30193 -13664
rect 30249 -13712 30303 -13656
rect 30359 -13712 30413 -13656
rect 30469 -13712 30536 -13656
rect 30139 -13720 30536 -13712
rect 29479 -13766 30536 -13720
rect 29479 -13774 30193 -13766
rect 29479 -13830 29533 -13774
rect 29589 -13830 29643 -13774
rect 29699 -13830 29753 -13774
rect 29809 -13830 29863 -13774
rect 29919 -13830 29973 -13774
rect 30029 -13830 30083 -13774
rect 30139 -13822 30193 -13774
rect 30249 -13822 30303 -13766
rect 30359 -13822 30413 -13766
rect 30469 -13822 30536 -13766
rect 30139 -13830 30536 -13822
rect 29479 -13897 30536 -13830
rect 113504 -13593 113550 -13537
rect 113606 -13593 113660 -13537
rect 113716 -13593 113770 -13537
rect 113826 -13593 113880 -13537
rect 113936 -13593 113990 -13537
rect 114046 -13593 114100 -13537
rect 114156 -13593 114210 -13537
rect 114266 -13593 126960 -13537
rect 113504 -13647 126960 -13593
rect 113504 -13703 113550 -13647
rect 113606 -13703 113660 -13647
rect 113716 -13703 113770 -13647
rect 113826 -13703 113880 -13647
rect 113936 -13703 113990 -13647
rect 114046 -13703 114100 -13647
rect 114156 -13703 114210 -13647
rect 114266 -13703 126960 -13647
rect 113504 -13757 126960 -13703
rect 113504 -13813 113550 -13757
rect 113606 -13813 113660 -13757
rect 113716 -13813 113770 -13757
rect 113826 -13813 113880 -13757
rect 113936 -13813 113990 -13757
rect 114046 -13813 114100 -13757
rect 114156 -13813 114210 -13757
rect 114266 -13813 126960 -13757
rect 113504 -13872 126960 -13813
rect 29799 -14469 30669 -14407
rect 29799 -14525 29852 -14469
rect 29908 -14525 29962 -14469
rect 30018 -14525 30072 -14469
rect 30128 -14525 30249 -14469
rect 30305 -14525 30359 -14469
rect 30415 -14525 30469 -14469
rect 30525 -14525 30669 -14469
rect 29799 -14579 30669 -14525
rect 29799 -14635 29852 -14579
rect 29908 -14635 29962 -14579
rect 30018 -14635 30072 -14579
rect 30128 -14635 30249 -14579
rect 30305 -14635 30359 -14579
rect 30415 -14635 30469 -14579
rect 30525 -14635 30669 -14579
rect 29799 -14722 30669 -14635
rect 10211 -15052 11790 -15012
rect 10211 -15108 10245 -15052
rect 10301 -15108 10355 -15052
rect 10411 -15108 10465 -15052
rect 10521 -15108 10575 -15052
rect 10631 -15108 10685 -15052
rect 10741 -15108 10795 -15052
rect 10851 -15108 10905 -15052
rect 10961 -15108 11034 -15052
rect 11090 -15108 11144 -15052
rect 11200 -15108 11254 -15052
rect 11310 -15108 11364 -15052
rect 11420 -15108 11474 -15052
rect 11530 -15108 11584 -15052
rect 11640 -15108 11694 -15052
rect 11750 -15108 11790 -15052
rect 10211 -15162 11790 -15108
rect 10211 -15218 10245 -15162
rect 10301 -15218 10355 -15162
rect 10411 -15218 10465 -15162
rect 10521 -15218 10575 -15162
rect 10631 -15218 10685 -15162
rect 10741 -15218 10795 -15162
rect 10851 -15218 10905 -15162
rect 10961 -15218 11034 -15162
rect 11090 -15218 11144 -15162
rect 11200 -15218 11254 -15162
rect 11310 -15218 11364 -15162
rect 11420 -15218 11474 -15162
rect 11530 -15218 11584 -15162
rect 11640 -15218 11694 -15162
rect 11750 -15218 11790 -15162
rect 10211 -15272 11790 -15218
rect 10211 -15328 10245 -15272
rect 10301 -15328 10355 -15272
rect 10411 -15328 10465 -15272
rect 10521 -15328 10575 -15272
rect 10631 -15328 10685 -15272
rect 10741 -15328 10795 -15272
rect 10851 -15328 10905 -15272
rect 10961 -15328 11034 -15272
rect 11090 -15328 11144 -15272
rect 11200 -15328 11254 -15272
rect 11310 -15328 11364 -15272
rect 11420 -15328 11474 -15272
rect 11530 -15328 11584 -15272
rect 11640 -15328 11694 -15272
rect 11750 -15328 11790 -15272
rect 10211 -15382 11790 -15328
rect 10211 -15438 10245 -15382
rect 10301 -15438 10355 -15382
rect 10411 -15438 10465 -15382
rect 10521 -15438 10575 -15382
rect 10631 -15438 10685 -15382
rect 10741 -15438 10795 -15382
rect 10851 -15438 10905 -15382
rect 10961 -15438 11034 -15382
rect 11090 -15438 11144 -15382
rect 11200 -15438 11254 -15382
rect 11310 -15438 11364 -15382
rect 11420 -15438 11474 -15382
rect 11530 -15438 11584 -15382
rect 11640 -15438 11694 -15382
rect 11750 -15438 11790 -15382
rect 10211 -15492 11790 -15438
rect 10211 -15548 10245 -15492
rect 10301 -15548 10355 -15492
rect 10411 -15548 10465 -15492
rect 10521 -15548 10575 -15492
rect 10631 -15548 10685 -15492
rect 10741 -15548 10795 -15492
rect 10851 -15548 10905 -15492
rect 10961 -15548 11034 -15492
rect 11090 -15548 11144 -15492
rect 11200 -15548 11254 -15492
rect 11310 -15548 11364 -15492
rect 11420 -15548 11474 -15492
rect 11530 -15548 11584 -15492
rect 11640 -15548 11694 -15492
rect 11750 -15548 11790 -15492
rect 10211 -15602 11790 -15548
rect 10211 -15658 10245 -15602
rect 10301 -15658 10355 -15602
rect 10411 -15658 10465 -15602
rect 10521 -15658 10575 -15602
rect 10631 -15658 10685 -15602
rect 10741 -15658 10795 -15602
rect 10851 -15658 10905 -15602
rect 10961 -15658 11034 -15602
rect 11090 -15658 11144 -15602
rect 11200 -15658 11254 -15602
rect 11310 -15658 11364 -15602
rect 11420 -15658 11474 -15602
rect 11530 -15658 11584 -15602
rect 11640 -15658 11694 -15602
rect 11750 -15658 11790 -15602
rect 10211 -15730 11790 -15658
rect 31290 -15618 31736 -15591
rect 31290 -15674 31310 -15618
rect 31366 -15674 31420 -15618
rect 31476 -15674 31530 -15618
rect 31586 -15674 31640 -15618
rect 31696 -15674 31736 -15618
rect 31290 -15728 31736 -15674
rect 31290 -15784 31310 -15728
rect 31366 -15784 31420 -15728
rect 31476 -15784 31530 -15728
rect 31586 -15784 31640 -15728
rect 31696 -15784 31736 -15728
rect 31290 -15817 31736 -15784
rect 29756 -19802 30209 -19778
rect 29756 -19858 29779 -19802
rect 29835 -19858 29889 -19802
rect 29945 -19858 29999 -19802
rect 30055 -19858 30109 -19802
rect 30165 -19858 30209 -19802
rect 29756 -19879 30209 -19858
rect 30310 -19809 30763 -19785
rect 30310 -19865 30333 -19809
rect 30389 -19865 30443 -19809
rect 30499 -19865 30553 -19809
rect 30609 -19865 30663 -19809
rect 30719 -19865 30763 -19809
rect 30310 -19886 30763 -19865
rect 30864 -19800 31317 -19776
rect 30864 -19856 30887 -19800
rect 30943 -19856 30997 -19800
rect 31053 -19856 31107 -19800
rect 31163 -19856 31217 -19800
rect 31273 -19856 31317 -19800
rect 30864 -19877 31317 -19856
rect 31404 -19816 31857 -19792
rect 31404 -19872 31427 -19816
rect 31483 -19872 31537 -19816
rect 31593 -19872 31647 -19816
rect 31703 -19872 31757 -19816
rect 31813 -19872 31857 -19816
rect 31404 -19893 31857 -19872
rect 25859 -21422 26715 -21402
rect 25859 -21478 25916 -21422
rect 25972 -21478 26026 -21422
rect 26082 -21478 26136 -21422
rect 26192 -21478 26246 -21422
rect 26302 -21478 26356 -21422
rect 26412 -21478 26466 -21422
rect 26522 -21478 26576 -21422
rect 26632 -21435 26715 -21422
rect 26632 -21478 32404 -21435
rect 25859 -21532 32404 -21478
rect 25859 -21588 25916 -21532
rect 25972 -21588 26026 -21532
rect 26082 -21588 26136 -21532
rect 26192 -21588 26246 -21532
rect 26302 -21588 26356 -21532
rect 26412 -21588 26466 -21532
rect 26522 -21588 26576 -21532
rect 26632 -21588 32404 -21532
rect 25859 -21642 32404 -21588
rect 25859 -21698 25916 -21642
rect 25972 -21698 26026 -21642
rect 26082 -21698 26136 -21642
rect 26192 -21698 26246 -21642
rect 26302 -21698 26356 -21642
rect 26412 -21698 26466 -21642
rect 26522 -21698 26576 -21642
rect 26632 -21698 32404 -21642
rect 25859 -21770 32404 -21698
rect 14282 -23938 25532 -23937
rect 14282 -23994 24635 -23938
rect 24691 -23994 24745 -23938
rect 24801 -23994 24855 -23938
rect 24911 -23994 24965 -23938
rect 25021 -23994 25075 -23938
rect 25131 -23994 25185 -23938
rect 25241 -23994 25295 -23938
rect 25351 -23994 25405 -23938
rect 25461 -23994 25532 -23938
rect 14282 -24048 25532 -23994
rect 14282 -24104 24635 -24048
rect 24691 -24104 24745 -24048
rect 24801 -24104 24855 -24048
rect 24911 -24104 24965 -24048
rect 25021 -24104 25075 -24048
rect 25131 -24104 25185 -24048
rect 25241 -24104 25295 -24048
rect 25351 -24104 25405 -24048
rect 25461 -24104 25532 -24048
rect 14282 -24158 25532 -24104
rect 14282 -24214 24635 -24158
rect 24691 -24214 24745 -24158
rect 24801 -24214 24855 -24158
rect 24911 -24214 24965 -24158
rect 25021 -24214 25075 -24158
rect 25131 -24214 25185 -24158
rect 25241 -24214 25295 -24158
rect 25351 -24214 25405 -24158
rect 25461 -24214 25532 -24158
rect 14282 -24268 25532 -24214
rect 14282 -24324 24635 -24268
rect 24691 -24324 24745 -24268
rect 24801 -24324 24855 -24268
rect 24911 -24324 24965 -24268
rect 25021 -24324 25075 -24268
rect 25131 -24324 25185 -24268
rect 25241 -24324 25295 -24268
rect 25351 -24324 25405 -24268
rect 25461 -24324 25532 -24268
rect 14282 -24378 25532 -24324
rect 14282 -24434 24635 -24378
rect 24691 -24434 24745 -24378
rect 24801 -24434 24855 -24378
rect 24911 -24434 24965 -24378
rect 25021 -24434 25075 -24378
rect 25131 -24434 25185 -24378
rect 25241 -24434 25295 -24378
rect 25351 -24434 25405 -24378
rect 25461 -24434 25532 -24378
rect 14282 -24488 25532 -24434
rect 14282 -24544 24635 -24488
rect 24691 -24544 24745 -24488
rect 24801 -24544 24855 -24488
rect 24911 -24544 24965 -24488
rect 25021 -24544 25075 -24488
rect 25131 -24544 25185 -24488
rect 25241 -24544 25295 -24488
rect 25351 -24544 25405 -24488
rect 25461 -24544 25532 -24488
rect 39287 -28947 40068 -26510
rect 41809 -27308 42183 -27305
rect 39287 -29003 39307 -28947
rect 39363 -29003 39417 -28947
rect 39473 -29003 39527 -28947
rect 39583 -29003 39637 -28947
rect 39693 -29003 39747 -28947
rect 39803 -29003 39857 -28947
rect 39913 -29003 39967 -28947
rect 40023 -29003 40068 -28947
rect 39287 -29057 40068 -29003
rect 39287 -29113 39307 -29057
rect 39363 -29113 39417 -29057
rect 39473 -29113 39527 -29057
rect 39583 -29113 39637 -29057
rect 39693 -29113 39747 -29057
rect 39803 -29113 39857 -29057
rect 39913 -29113 39967 -29057
rect 40023 -29113 40068 -29057
rect 39287 -29167 40068 -29113
rect 39287 -29223 39307 -29167
rect 39363 -29223 39417 -29167
rect 39473 -29223 39527 -29167
rect 39583 -29223 39637 -29167
rect 39693 -29223 39747 -29167
rect 39803 -29223 39857 -29167
rect 39913 -29223 39967 -29167
rect 40023 -29223 40068 -29167
rect 39287 -29277 40068 -29223
rect 39287 -29333 39307 -29277
rect 39363 -29333 39417 -29277
rect 39473 -29333 39527 -29277
rect 39583 -29333 39637 -29277
rect 39693 -29333 39747 -29277
rect 39803 -29333 39857 -29277
rect 39913 -29333 39967 -29277
rect 40023 -29333 40068 -29277
rect 39287 -29387 40068 -29333
rect 39287 -29443 39307 -29387
rect 39363 -29443 39417 -29387
rect 39473 -29443 39527 -29387
rect 39583 -29443 39637 -29387
rect 39693 -29443 39747 -29387
rect 39803 -29443 39857 -29387
rect 39913 -29443 39967 -29387
rect 40023 -29443 40068 -29387
rect 39287 -29497 40068 -29443
rect 39287 -29553 39307 -29497
rect 39363 -29553 39417 -29497
rect 39473 -29553 39527 -29497
rect 39583 -29553 39637 -29497
rect 39693 -29553 39747 -29497
rect 39803 -29553 39857 -29497
rect 39913 -29553 39967 -29497
rect 40023 -29553 40068 -29497
rect 10215 -29666 24123 -29577
rect 10214 -29695 24123 -29666
rect 10214 -29751 10249 -29695
rect 10305 -29751 10359 -29695
rect 10415 -29751 10469 -29695
rect 10525 -29751 10579 -29695
rect 10635 -29751 10689 -29695
rect 10745 -29751 10799 -29695
rect 10855 -29751 10909 -29695
rect 10965 -29751 11038 -29695
rect 11094 -29751 11148 -29695
rect 11204 -29751 11258 -29695
rect 11314 -29751 11368 -29695
rect 11424 -29751 11478 -29695
rect 11534 -29751 11588 -29695
rect 11644 -29751 11698 -29695
rect 11754 -29751 24123 -29695
rect 10214 -29805 24123 -29751
rect 10214 -29861 10249 -29805
rect 10305 -29861 10359 -29805
rect 10415 -29861 10469 -29805
rect 10525 -29861 10579 -29805
rect 10635 -29861 10689 -29805
rect 10745 -29861 10799 -29805
rect 10855 -29861 10909 -29805
rect 10965 -29861 11038 -29805
rect 11094 -29861 11148 -29805
rect 11204 -29861 11258 -29805
rect 11314 -29861 11368 -29805
rect 11424 -29861 11478 -29805
rect 11534 -29861 11588 -29805
rect 11644 -29861 11698 -29805
rect 11754 -29861 24123 -29805
rect 39287 -29607 40068 -29553
rect 39287 -29663 39307 -29607
rect 39363 -29663 39417 -29607
rect 39473 -29663 39527 -29607
rect 39583 -29663 39637 -29607
rect 39693 -29663 39747 -29607
rect 39803 -29663 39857 -29607
rect 39913 -29663 39967 -29607
rect 40023 -29663 40068 -29607
rect 39287 -29717 40068 -29663
rect 39287 -29773 39307 -29717
rect 39363 -29773 39417 -29717
rect 39473 -29773 39527 -29717
rect 39583 -29773 39637 -29717
rect 39693 -29773 39747 -29717
rect 39803 -29773 39857 -29717
rect 39913 -29773 39967 -29717
rect 40023 -29773 40068 -29717
rect 39287 -29832 40068 -29773
rect 10214 -29915 24123 -29861
rect 10214 -29971 10249 -29915
rect 10305 -29971 10359 -29915
rect 10415 -29971 10469 -29915
rect 10525 -29971 10579 -29915
rect 10635 -29971 10689 -29915
rect 10745 -29971 10799 -29915
rect 10855 -29971 10909 -29915
rect 10965 -29971 11038 -29915
rect 11094 -29971 11148 -29915
rect 11204 -29971 11258 -29915
rect 11314 -29971 11368 -29915
rect 11424 -29971 11478 -29915
rect 11534 -29971 11588 -29915
rect 11644 -29971 11698 -29915
rect 11754 -29971 24123 -29915
rect 10214 -30025 24123 -29971
rect 10214 -30081 10249 -30025
rect 10305 -30081 10359 -30025
rect 10415 -30081 10469 -30025
rect 10525 -30081 10579 -30025
rect 10635 -30081 10689 -30025
rect 10745 -30081 10799 -30025
rect 10855 -30081 10909 -30025
rect 10965 -30081 11038 -30025
rect 11094 -30081 11148 -30025
rect 11204 -30081 11258 -30025
rect 11314 -30081 11368 -30025
rect 11424 -30081 11478 -30025
rect 11534 -30081 11588 -30025
rect 11644 -30081 11698 -30025
rect 11754 -30081 24123 -30025
rect 10214 -30105 24123 -30081
rect 10214 -30194 24122 -30105
rect 41815 -30387 42183 -27308
rect 43208 -30387 43576 -27294
rect 45124 -30387 45492 -27261
rect 46707 -30387 47075 -27272
rect 48200 -30387 48568 -27305
rect 49593 -30387 49961 -27261
rect 50707 -30387 51075 -27261
rect 51454 -30387 51822 -27261
rect 54502 -30387 55314 -23109
rect 56577 -27796 57328 -26578
rect 56571 -27818 57329 -27796
rect 56571 -27874 56591 -27818
rect 56647 -27874 56701 -27818
rect 56757 -27874 56811 -27818
rect 56867 -27874 56921 -27818
rect 56977 -27874 57031 -27818
rect 57087 -27874 57141 -27818
rect 57197 -27874 57251 -27818
rect 57307 -27874 57329 -27818
rect 56571 -27928 57329 -27874
rect 56571 -27984 56591 -27928
rect 56647 -27984 56701 -27928
rect 56757 -27984 56811 -27928
rect 56867 -27984 56921 -27928
rect 56977 -27984 57031 -27928
rect 57087 -27984 57141 -27928
rect 57197 -27984 57251 -27928
rect 57307 -27984 57329 -27928
rect 56571 -28038 57329 -27984
rect 56571 -28094 56591 -28038
rect 56647 -28094 56701 -28038
rect 56757 -28094 56811 -28038
rect 56867 -28094 56921 -28038
rect 56977 -28094 57031 -28038
rect 57087 -28094 57141 -28038
rect 57197 -28094 57251 -28038
rect 57307 -28094 57329 -28038
rect 56571 -28148 57329 -28094
rect 56571 -28204 56591 -28148
rect 56647 -28204 56701 -28148
rect 56757 -28204 56811 -28148
rect 56867 -28204 56921 -28148
rect 56977 -28204 57031 -28148
rect 57087 -28204 57141 -28148
rect 57197 -28204 57251 -28148
rect 57307 -28204 57329 -28148
rect 56571 -28258 57329 -28204
rect 56571 -28314 56591 -28258
rect 56647 -28314 56701 -28258
rect 56757 -28314 56811 -28258
rect 56867 -28314 56921 -28258
rect 56977 -28314 57031 -28258
rect 57087 -28314 57141 -28258
rect 57197 -28314 57251 -28258
rect 57307 -28314 57329 -28258
rect 56571 -28368 57329 -28314
rect 56571 -28424 56591 -28368
rect 56647 -28424 56701 -28368
rect 56757 -28424 56811 -28368
rect 56867 -28424 56921 -28368
rect 56977 -28424 57031 -28368
rect 57087 -28424 57141 -28368
rect 57197 -28424 57251 -28368
rect 57307 -28424 57329 -28368
rect 56571 -28478 57329 -28424
rect 56571 -28534 56591 -28478
rect 56647 -28534 56701 -28478
rect 56757 -28534 56811 -28478
rect 56867 -28534 56921 -28478
rect 56977 -28534 57031 -28478
rect 57087 -28534 57141 -28478
rect 57197 -28534 57251 -28478
rect 57307 -28534 57329 -28478
rect 56571 -28588 57329 -28534
rect 56571 -28644 56591 -28588
rect 56647 -28644 56701 -28588
rect 56757 -28644 56811 -28588
rect 56867 -28644 56921 -28588
rect 56977 -28644 57031 -28588
rect 57087 -28644 57141 -28588
rect 57197 -28644 57251 -28588
rect 57307 -28644 57329 -28588
rect 56571 -28703 57329 -28644
rect 58734 -30387 59125 -27331
rect 59948 -30387 60339 -27331
rect 61345 -30387 61736 -27331
rect 62742 -30387 63133 -27304
rect 64021 -30387 64412 -27318
rect 65183 -30387 65574 -27318
rect 66488 -30387 66879 -27344
rect 67481 -30387 67872 -27304
rect 68447 -30387 68838 -27331
rect 4105 -30448 128964 -30387
rect 4105 -30497 113577 -30448
rect 4105 -30553 24746 -30497
rect 24802 -30553 24856 -30497
rect 24912 -30553 24966 -30497
rect 25022 -30553 25076 -30497
rect 25132 -30553 25186 -30497
rect 25242 -30553 25296 -30497
rect 25352 -30553 25406 -30497
rect 25462 -30504 113577 -30497
rect 113633 -30504 113687 -30448
rect 113743 -30504 113797 -30448
rect 113853 -30504 113907 -30448
rect 113963 -30504 114017 -30448
rect 114073 -30504 114127 -30448
rect 114183 -30504 114237 -30448
rect 114293 -30504 128964 -30448
rect 25462 -30553 128964 -30504
rect 4105 -30558 128964 -30553
rect 4105 -30607 113577 -30558
rect 4105 -30663 24746 -30607
rect 24802 -30663 24856 -30607
rect 24912 -30663 24966 -30607
rect 25022 -30663 25076 -30607
rect 25132 -30663 25186 -30607
rect 25242 -30663 25296 -30607
rect 25352 -30663 25406 -30607
rect 25462 -30614 113577 -30607
rect 113633 -30614 113687 -30558
rect 113743 -30614 113797 -30558
rect 113853 -30614 113907 -30558
rect 113963 -30614 114017 -30558
rect 114073 -30614 114127 -30558
rect 114183 -30614 114237 -30558
rect 114293 -30614 128964 -30558
rect 25462 -30663 128964 -30614
rect 4105 -30668 128964 -30663
rect 4105 -30717 113577 -30668
rect 4105 -30773 24746 -30717
rect 24802 -30773 24856 -30717
rect 24912 -30773 24966 -30717
rect 25022 -30773 25076 -30717
rect 25132 -30773 25186 -30717
rect 25242 -30773 25296 -30717
rect 25352 -30773 25406 -30717
rect 25462 -30724 113577 -30717
rect 113633 -30724 113687 -30668
rect 113743 -30724 113797 -30668
rect 113853 -30724 113907 -30668
rect 113963 -30724 114017 -30668
rect 114073 -30724 114127 -30668
rect 114183 -30724 114237 -30668
rect 114293 -30724 128964 -30668
rect 25462 -30773 128964 -30724
rect 4105 -30778 128964 -30773
rect 4105 -30827 113577 -30778
rect 4105 -30883 24746 -30827
rect 24802 -30883 24856 -30827
rect 24912 -30883 24966 -30827
rect 25022 -30883 25076 -30827
rect 25132 -30883 25186 -30827
rect 25242 -30883 25296 -30827
rect 25352 -30883 25406 -30827
rect 25462 -30834 113577 -30827
rect 113633 -30834 113687 -30778
rect 113743 -30834 113797 -30778
rect 113853 -30834 113907 -30778
rect 113963 -30834 114017 -30778
rect 114073 -30834 114127 -30778
rect 114183 -30834 114237 -30778
rect 114293 -30834 128964 -30778
rect 25462 -30883 128964 -30834
rect 4105 -30888 128964 -30883
rect 4105 -30937 113577 -30888
rect 4105 -30993 24746 -30937
rect 24802 -30993 24856 -30937
rect 24912 -30993 24966 -30937
rect 25022 -30993 25076 -30937
rect 25132 -30993 25186 -30937
rect 25242 -30993 25296 -30937
rect 25352 -30993 25406 -30937
rect 25462 -30944 113577 -30937
rect 113633 -30944 113687 -30888
rect 113743 -30944 113797 -30888
rect 113853 -30944 113907 -30888
rect 113963 -30944 114017 -30888
rect 114073 -30944 114127 -30888
rect 114183 -30944 114237 -30888
rect 114293 -30944 128964 -30888
rect 25462 -30993 128964 -30944
rect 4105 -30998 128964 -30993
rect 4105 -31047 113577 -30998
rect 4105 -31103 24746 -31047
rect 24802 -31103 24856 -31047
rect 24912 -31103 24966 -31047
rect 25022 -31103 25076 -31047
rect 25132 -31103 25186 -31047
rect 25242 -31103 25296 -31047
rect 25352 -31103 25406 -31047
rect 25462 -31054 113577 -31047
rect 113633 -31054 113687 -30998
rect 113743 -31054 113797 -30998
rect 113853 -31054 113907 -30998
rect 113963 -31054 114017 -30998
rect 114073 -31054 114127 -30998
rect 114183 -31054 114237 -30998
rect 114293 -31054 128964 -30998
rect 25462 -31103 128964 -31054
rect 4105 -31287 128964 -31103
rect 3997 -31614 128856 -31467
rect 3997 -31670 25910 -31614
rect 25966 -31670 26020 -31614
rect 26076 -31670 26130 -31614
rect 26186 -31670 26240 -31614
rect 26296 -31670 26350 -31614
rect 26406 -31670 26460 -31614
rect 26516 -31670 26570 -31614
rect 26626 -31659 128856 -31614
rect 26626 -31670 114633 -31659
rect 3997 -31672 114633 -31670
rect 3997 -31728 10247 -31672
rect 10303 -31728 10357 -31672
rect 10413 -31728 10467 -31672
rect 10523 -31728 10577 -31672
rect 10633 -31728 10687 -31672
rect 10743 -31728 10797 -31672
rect 10853 -31728 10907 -31672
rect 10963 -31728 11036 -31672
rect 11092 -31728 11146 -31672
rect 11202 -31728 11256 -31672
rect 11312 -31728 11366 -31672
rect 11422 -31728 11476 -31672
rect 11532 -31728 11586 -31672
rect 11642 -31728 11696 -31672
rect 11752 -31715 114633 -31672
rect 114689 -31715 114743 -31659
rect 114799 -31715 114853 -31659
rect 114909 -31715 114963 -31659
rect 115019 -31715 115073 -31659
rect 115129 -31715 115183 -31659
rect 115239 -31715 115293 -31659
rect 115349 -31715 128856 -31659
rect 11752 -31724 128856 -31715
rect 11752 -31728 25910 -31724
rect 3997 -31780 25910 -31728
rect 25966 -31780 26020 -31724
rect 26076 -31780 26130 -31724
rect 26186 -31780 26240 -31724
rect 26296 -31780 26350 -31724
rect 26406 -31780 26460 -31724
rect 26516 -31780 26570 -31724
rect 26626 -31769 128856 -31724
rect 26626 -31780 114633 -31769
rect 3997 -31782 114633 -31780
rect 3997 -31838 10247 -31782
rect 10303 -31838 10357 -31782
rect 10413 -31838 10467 -31782
rect 10523 -31838 10577 -31782
rect 10633 -31838 10687 -31782
rect 10743 -31838 10797 -31782
rect 10853 -31838 10907 -31782
rect 10963 -31838 11036 -31782
rect 11092 -31838 11146 -31782
rect 11202 -31838 11256 -31782
rect 11312 -31838 11366 -31782
rect 11422 -31838 11476 -31782
rect 11532 -31838 11586 -31782
rect 11642 -31838 11696 -31782
rect 11752 -31825 114633 -31782
rect 114689 -31825 114743 -31769
rect 114799 -31825 114853 -31769
rect 114909 -31825 114963 -31769
rect 115019 -31825 115073 -31769
rect 115129 -31825 115183 -31769
rect 115239 -31825 115293 -31769
rect 115349 -31825 128856 -31769
rect 11752 -31834 128856 -31825
rect 11752 -31838 25910 -31834
rect 3997 -31890 25910 -31838
rect 25966 -31890 26020 -31834
rect 26076 -31890 26130 -31834
rect 26186 -31890 26240 -31834
rect 26296 -31890 26350 -31834
rect 26406 -31890 26460 -31834
rect 26516 -31890 26570 -31834
rect 26626 -31879 128856 -31834
rect 26626 -31890 114633 -31879
rect 3997 -31892 114633 -31890
rect 3997 -31948 10247 -31892
rect 10303 -31948 10357 -31892
rect 10413 -31948 10467 -31892
rect 10523 -31948 10577 -31892
rect 10633 -31948 10687 -31892
rect 10743 -31948 10797 -31892
rect 10853 -31948 10907 -31892
rect 10963 -31948 11036 -31892
rect 11092 -31948 11146 -31892
rect 11202 -31948 11256 -31892
rect 11312 -31948 11366 -31892
rect 11422 -31948 11476 -31892
rect 11532 -31948 11586 -31892
rect 11642 -31948 11696 -31892
rect 11752 -31935 114633 -31892
rect 114689 -31935 114743 -31879
rect 114799 -31935 114853 -31879
rect 114909 -31935 114963 -31879
rect 115019 -31935 115073 -31879
rect 115129 -31935 115183 -31879
rect 115239 -31935 115293 -31879
rect 115349 -31935 128856 -31879
rect 11752 -31944 128856 -31935
rect 11752 -31948 25910 -31944
rect 3997 -32000 25910 -31948
rect 25966 -32000 26020 -31944
rect 26076 -32000 26130 -31944
rect 26186 -32000 26240 -31944
rect 26296 -32000 26350 -31944
rect 26406 -32000 26460 -31944
rect 26516 -32000 26570 -31944
rect 26626 -31989 128856 -31944
rect 26626 -32000 114633 -31989
rect 3997 -32002 114633 -32000
rect 3997 -32058 10247 -32002
rect 10303 -32058 10357 -32002
rect 10413 -32058 10467 -32002
rect 10523 -32058 10577 -32002
rect 10633 -32058 10687 -32002
rect 10743 -32058 10797 -32002
rect 10853 -32058 10907 -32002
rect 10963 -32058 11036 -32002
rect 11092 -32058 11146 -32002
rect 11202 -32058 11256 -32002
rect 11312 -32058 11366 -32002
rect 11422 -32058 11476 -32002
rect 11532 -32058 11586 -32002
rect 11642 -32058 11696 -32002
rect 11752 -32045 114633 -32002
rect 114689 -32045 114743 -31989
rect 114799 -32045 114853 -31989
rect 114909 -32045 114963 -31989
rect 115019 -32045 115073 -31989
rect 115129 -32045 115183 -31989
rect 115239 -32045 115293 -31989
rect 115349 -32045 128856 -31989
rect 11752 -32054 128856 -32045
rect 11752 -32058 25910 -32054
rect 3997 -32110 25910 -32058
rect 25966 -32110 26020 -32054
rect 26076 -32110 26130 -32054
rect 26186 -32110 26240 -32054
rect 26296 -32110 26350 -32054
rect 26406 -32110 26460 -32054
rect 26516 -32110 26570 -32054
rect 26626 -32099 128856 -32054
rect 26626 -32110 114633 -32099
rect 3997 -32112 114633 -32110
rect 3997 -32168 10247 -32112
rect 10303 -32168 10357 -32112
rect 10413 -32168 10467 -32112
rect 10523 -32168 10577 -32112
rect 10633 -32168 10687 -32112
rect 10743 -32168 10797 -32112
rect 10853 -32168 10907 -32112
rect 10963 -32168 11036 -32112
rect 11092 -32168 11146 -32112
rect 11202 -32168 11256 -32112
rect 11312 -32168 11366 -32112
rect 11422 -32168 11476 -32112
rect 11532 -32168 11586 -32112
rect 11642 -32168 11696 -32112
rect 11752 -32155 114633 -32112
rect 114689 -32155 114743 -32099
rect 114799 -32155 114853 -32099
rect 114909 -32155 114963 -32099
rect 115019 -32155 115073 -32099
rect 115129 -32155 115183 -32099
rect 115239 -32155 115293 -32099
rect 115349 -32155 128856 -32099
rect 11752 -32164 128856 -32155
rect 11752 -32168 25910 -32164
rect 3997 -32220 25910 -32168
rect 25966 -32220 26020 -32164
rect 26076 -32220 26130 -32164
rect 26186 -32220 26240 -32164
rect 26296 -32220 26350 -32164
rect 26406 -32220 26460 -32164
rect 26516 -32220 26570 -32164
rect 26626 -32209 128856 -32164
rect 26626 -32220 114633 -32209
rect 3997 -32222 114633 -32220
rect 3997 -32278 10247 -32222
rect 10303 -32278 10357 -32222
rect 10413 -32278 10467 -32222
rect 10523 -32278 10577 -32222
rect 10633 -32278 10687 -32222
rect 10743 -32278 10797 -32222
rect 10853 -32278 10907 -32222
rect 10963 -32278 11036 -32222
rect 11092 -32278 11146 -32222
rect 11202 -32278 11256 -32222
rect 11312 -32278 11366 -32222
rect 11422 -32278 11476 -32222
rect 11532 -32278 11586 -32222
rect 11642 -32278 11696 -32222
rect 11752 -32265 114633 -32222
rect 114689 -32265 114743 -32209
rect 114799 -32265 114853 -32209
rect 114909 -32265 114963 -32209
rect 115019 -32265 115073 -32209
rect 115129 -32265 115183 -32209
rect 115239 -32265 115293 -32209
rect 115349 -32265 128856 -32209
rect 11752 -32278 128856 -32265
rect 3997 -32367 128856 -32278
<< via1 >>
rect 24715 19789 24771 19845
rect 24825 19789 24881 19845
rect 24935 19789 24991 19845
rect 25045 19789 25101 19845
rect 25155 19789 25211 19845
rect 25265 19789 25321 19845
rect 25375 19789 25431 19845
rect 113574 19804 113630 19860
rect 113684 19804 113740 19860
rect 113794 19804 113850 19860
rect 113904 19804 113960 19860
rect 114014 19804 114070 19860
rect 114124 19804 114180 19860
rect 114234 19804 114290 19860
rect 24715 19679 24771 19735
rect 24825 19679 24881 19735
rect 24935 19679 24991 19735
rect 25045 19679 25101 19735
rect 25155 19679 25211 19735
rect 25265 19679 25321 19735
rect 25375 19679 25431 19735
rect 113574 19694 113630 19750
rect 113684 19694 113740 19750
rect 113794 19694 113850 19750
rect 113904 19694 113960 19750
rect 114014 19694 114070 19750
rect 114124 19694 114180 19750
rect 114234 19694 114290 19750
rect 24715 19569 24771 19625
rect 24825 19569 24881 19625
rect 24935 19569 24991 19625
rect 25045 19569 25101 19625
rect 25155 19569 25211 19625
rect 25265 19569 25321 19625
rect 25375 19569 25431 19625
rect 113574 19584 113630 19640
rect 113684 19584 113740 19640
rect 113794 19584 113850 19640
rect 113904 19584 113960 19640
rect 114014 19584 114070 19640
rect 114124 19584 114180 19640
rect 114234 19584 114290 19640
rect 24715 19459 24771 19515
rect 24825 19459 24881 19515
rect 24935 19459 24991 19515
rect 25045 19459 25101 19515
rect 25155 19459 25211 19515
rect 25265 19459 25321 19515
rect 25375 19459 25431 19515
rect 113574 19474 113630 19530
rect 113684 19474 113740 19530
rect 113794 19474 113850 19530
rect 113904 19474 113960 19530
rect 114014 19474 114070 19530
rect 114124 19474 114180 19530
rect 114234 19474 114290 19530
rect 24715 19349 24771 19405
rect 24825 19349 24881 19405
rect 24935 19349 24991 19405
rect 25045 19349 25101 19405
rect 25155 19349 25211 19405
rect 25265 19349 25321 19405
rect 25375 19349 25431 19405
rect 113574 19364 113630 19420
rect 113684 19364 113740 19420
rect 113794 19364 113850 19420
rect 113904 19364 113960 19420
rect 114014 19364 114070 19420
rect 114124 19364 114180 19420
rect 114234 19364 114290 19420
rect 24715 19239 24771 19295
rect 24825 19239 24881 19295
rect 24935 19239 24991 19295
rect 25045 19239 25101 19295
rect 25155 19239 25211 19295
rect 25265 19239 25321 19295
rect 25375 19239 25431 19295
rect 113574 19254 113630 19310
rect 113684 19254 113740 19310
rect 113794 19254 113850 19310
rect 113904 19254 113960 19310
rect 114014 19254 114070 19310
rect 114124 19254 114180 19310
rect 114234 19254 114290 19310
rect 25931 18560 25987 18616
rect 26041 18560 26097 18616
rect 26151 18560 26207 18616
rect 26261 18560 26317 18616
rect 26371 18560 26427 18616
rect 26481 18560 26537 18616
rect 26591 18560 26647 18616
rect 114647 18519 114703 18575
rect 114757 18519 114813 18575
rect 114867 18519 114923 18575
rect 114977 18519 115033 18575
rect 115087 18519 115143 18575
rect 115197 18519 115253 18575
rect 115307 18519 115363 18575
rect 25931 18450 25987 18506
rect 26041 18450 26097 18506
rect 26151 18450 26207 18506
rect 26261 18450 26317 18506
rect 26371 18450 26427 18506
rect 26481 18450 26537 18506
rect 26591 18450 26647 18506
rect 114647 18409 114703 18465
rect 114757 18409 114813 18465
rect 114867 18409 114923 18465
rect 114977 18409 115033 18465
rect 115087 18409 115143 18465
rect 115197 18409 115253 18465
rect 115307 18409 115363 18465
rect 25931 18340 25987 18396
rect 26041 18340 26097 18396
rect 26151 18340 26207 18396
rect 26261 18340 26317 18396
rect 26371 18340 26427 18396
rect 26481 18340 26537 18396
rect 26591 18340 26647 18396
rect 114647 18299 114703 18355
rect 114757 18299 114813 18355
rect 114867 18299 114923 18355
rect 114977 18299 115033 18355
rect 115087 18299 115143 18355
rect 115197 18299 115253 18355
rect 115307 18299 115363 18355
rect 25931 18230 25987 18286
rect 26041 18230 26097 18286
rect 26151 18230 26207 18286
rect 26261 18230 26317 18286
rect 26371 18230 26427 18286
rect 26481 18230 26537 18286
rect 26591 18230 26647 18286
rect 114647 18189 114703 18245
rect 114757 18189 114813 18245
rect 114867 18189 114923 18245
rect 114977 18189 115033 18245
rect 115087 18189 115143 18245
rect 115197 18189 115253 18245
rect 115307 18189 115363 18245
rect 25931 18120 25987 18176
rect 26041 18120 26097 18176
rect 26151 18120 26207 18176
rect 26261 18120 26317 18176
rect 26371 18120 26427 18176
rect 26481 18120 26537 18176
rect 26591 18120 26647 18176
rect 114647 18079 114703 18135
rect 114757 18079 114813 18135
rect 114867 18079 114923 18135
rect 114977 18079 115033 18135
rect 115087 18079 115143 18135
rect 115197 18079 115253 18135
rect 115307 18079 115363 18135
rect 25931 18010 25987 18066
rect 26041 18010 26097 18066
rect 26151 18010 26207 18066
rect 26261 18010 26317 18066
rect 26371 18010 26427 18066
rect 26481 18010 26537 18066
rect 26591 18010 26647 18066
rect 114647 17969 114703 18025
rect 114757 17969 114813 18025
rect 114867 17969 114923 18025
rect 114977 17969 115033 18025
rect 115087 17969 115143 18025
rect 115197 17969 115253 18025
rect 115307 17969 115363 18025
rect 113535 13042 113591 13098
rect 113645 13042 113701 13098
rect 113755 13042 113811 13098
rect 113865 13042 113921 13098
rect 113975 13042 114031 13098
rect 114085 13042 114141 13098
rect 114195 13042 114251 13098
rect 113535 12932 113591 12988
rect 113645 12932 113701 12988
rect 113755 12932 113811 12988
rect 113865 12932 113921 12988
rect 113975 12932 114031 12988
rect 114085 12932 114141 12988
rect 114195 12932 114251 12988
rect 113535 12822 113591 12878
rect 113645 12822 113701 12878
rect 113755 12822 113811 12878
rect 113865 12822 113921 12878
rect 113975 12822 114031 12878
rect 114085 12822 114141 12878
rect 114195 12822 114251 12878
rect 113535 12712 113591 12768
rect 113645 12712 113701 12768
rect 113755 12712 113811 12768
rect 113865 12712 113921 12768
rect 113975 12712 114031 12768
rect 114085 12712 114141 12768
rect 114195 12712 114251 12768
rect 113535 12602 113591 12658
rect 113645 12602 113701 12658
rect 113755 12602 113811 12658
rect 113865 12602 113921 12658
rect 113975 12602 114031 12658
rect 114085 12602 114141 12658
rect 114195 12602 114251 12658
rect 113535 12492 113591 12548
rect 113645 12492 113701 12548
rect 113755 12492 113811 12548
rect 113865 12492 113921 12548
rect 113975 12492 114031 12548
rect 114085 12492 114141 12548
rect 114195 12492 114251 12548
rect 116770 9949 116826 10005
rect 116770 9839 116826 9895
rect 116770 9729 116826 9785
rect 116770 9619 116826 9675
rect 116770 9509 116826 9565
rect 116770 9399 116826 9455
rect 116770 8374 116826 8430
rect 116770 8264 116826 8320
rect 116770 8154 116826 8210
rect 116770 8044 116826 8100
rect 116770 7934 116826 7990
rect 116770 7824 116826 7880
rect 129243 7774 129299 7830
rect 129353 7774 129409 7830
rect 130252 7776 130308 7832
rect 130362 7776 130418 7832
rect 43928 6194 43984 6250
rect 44038 6194 44094 6250
rect 44148 6194 44204 6250
rect 44258 6194 44314 6250
rect 44368 6194 44424 6250
rect 43928 6084 43984 6140
rect 44038 6084 44094 6140
rect 44148 6084 44204 6140
rect 44258 6084 44314 6140
rect 44368 6084 44424 6140
rect 43928 5974 43984 6030
rect 44038 5974 44094 6030
rect 44148 5974 44204 6030
rect 44258 5974 44314 6030
rect 44368 5974 44424 6030
rect 46418 6253 46474 6309
rect 46528 6253 46584 6309
rect 46638 6253 46694 6309
rect 46748 6253 46804 6309
rect 46858 6253 46914 6309
rect 46638 6143 46694 6199
rect 46748 6143 46804 6199
rect 46858 6143 46914 6199
rect 46638 6033 46694 6089
rect 46748 6033 46804 6089
rect 46858 6033 46914 6089
rect -808 2892 -752 2948
rect -698 2892 -642 2948
rect -588 2892 -532 2948
rect -478 2892 -422 2948
rect -368 2892 -312 2948
rect -258 2892 -202 2948
rect -148 2892 -92 2948
rect -808 2782 -752 2838
rect -698 2782 -642 2838
rect -588 2782 -532 2838
rect -478 2782 -422 2838
rect -368 2782 -312 2838
rect -258 2782 -202 2838
rect -148 2782 -92 2838
rect 10800 3387 10856 3443
rect 10910 3387 10966 3443
rect 11020 3387 11076 3443
rect 11130 3387 11186 3443
rect 11240 3387 11296 3443
rect 11350 3387 11406 3443
rect 11460 3387 11516 3443
rect 11624 3387 11680 3443
rect 11734 3387 11790 3443
rect 11844 3387 11900 3443
rect 11954 3387 12010 3443
rect 12064 3387 12120 3443
rect 12174 3387 12230 3443
rect 12284 3387 12340 3443
rect 10800 3277 10856 3333
rect 10910 3277 10966 3333
rect 11020 3277 11076 3333
rect 11130 3277 11186 3333
rect 11240 3277 11296 3333
rect 11350 3277 11406 3333
rect 11460 3277 11516 3333
rect 11624 3277 11680 3333
rect 11734 3277 11790 3333
rect 11844 3277 11900 3333
rect 11954 3277 12010 3333
rect 12064 3277 12120 3333
rect 12174 3277 12230 3333
rect 12284 3277 12340 3333
rect 10800 3167 10856 3223
rect 10910 3167 10966 3223
rect 11020 3167 11076 3223
rect 11130 3167 11186 3223
rect 11240 3167 11296 3223
rect 11350 3167 11406 3223
rect 11460 3167 11516 3223
rect 11624 3167 11680 3223
rect 11734 3167 11790 3223
rect 11844 3167 11900 3223
rect 11954 3167 12010 3223
rect 12064 3167 12120 3223
rect 12174 3167 12230 3223
rect 12284 3167 12340 3223
rect 10800 3057 10856 3113
rect 10910 3057 10966 3113
rect 11020 3057 11076 3113
rect 11130 3057 11186 3113
rect 11240 3057 11296 3113
rect 11350 3057 11406 3113
rect 11460 3057 11516 3113
rect 11624 3057 11680 3113
rect 11734 3057 11790 3113
rect 11844 3057 11900 3113
rect 11954 3057 12010 3113
rect 12064 3057 12120 3113
rect 12174 3057 12230 3113
rect 12284 3057 12340 3113
rect 10800 2947 10856 3003
rect 10910 2947 10966 3003
rect 11020 2947 11076 3003
rect 11130 2947 11186 3003
rect 11240 2947 11296 3003
rect 11350 2947 11406 3003
rect 11460 2947 11516 3003
rect 11624 2947 11680 3003
rect 11734 2947 11790 3003
rect 11844 2947 11900 3003
rect 11954 2947 12010 3003
rect 12064 2947 12120 3003
rect 12174 2947 12230 3003
rect 12284 2947 12340 3003
rect 10800 2837 10856 2893
rect 10910 2837 10966 2893
rect 11020 2837 11076 2893
rect 11130 2837 11186 2893
rect 11240 2837 11296 2893
rect 11350 2837 11406 2893
rect 11460 2837 11516 2893
rect 11624 2837 11680 2893
rect 11734 2837 11790 2893
rect 11844 2837 11900 2893
rect 11954 2837 12010 2893
rect 12064 2837 12120 2893
rect 12174 2837 12230 2893
rect 12284 2837 12340 2893
rect -808 2672 -752 2728
rect -698 2672 -642 2728
rect -588 2672 -532 2728
rect -478 2672 -422 2728
rect -368 2672 -312 2728
rect -258 2672 -202 2728
rect -148 2672 -92 2728
rect -808 2562 -752 2618
rect -698 2562 -642 2618
rect -588 2562 -532 2618
rect -478 2562 -422 2618
rect -368 2562 -312 2618
rect -258 2562 -202 2618
rect -148 2562 -92 2618
rect 3111 2581 3167 2637
rect 3221 2581 3277 2637
rect 3331 2581 3387 2637
rect 3441 2581 3497 2637
rect -808 2452 -752 2508
rect -698 2452 -642 2508
rect -588 2452 -532 2508
rect -478 2452 -422 2508
rect -368 2452 -312 2508
rect -258 2452 -202 2508
rect -148 2452 -92 2508
rect 3111 2471 3167 2527
rect 3221 2471 3277 2527
rect 3331 2471 3387 2527
rect 3441 2471 3497 2527
rect -808 2342 -752 2398
rect -698 2342 -642 2398
rect -588 2342 -532 2398
rect -478 2342 -422 2398
rect -368 2342 -312 2398
rect -258 2342 -202 2398
rect -148 2342 -92 2398
rect 3111 2361 3167 2417
rect 3221 2361 3277 2417
rect 3331 2361 3387 2417
rect 3441 2361 3497 2417
rect 3111 2251 3167 2307
rect 3221 2251 3277 2307
rect 3331 2251 3387 2307
rect 3441 2251 3497 2307
rect 6315 1130 6371 1186
rect 6425 1130 6481 1186
rect 6535 1130 6591 1186
rect 6645 1130 6701 1186
rect 6755 1130 6811 1186
rect 6865 1130 6921 1186
rect 6975 1130 7031 1186
rect 22896 1136 22952 1192
rect 23006 1136 23062 1192
rect 23116 1136 23172 1192
rect 23226 1136 23282 1192
rect 23336 1136 23392 1192
rect 23446 1136 23502 1192
rect 23556 1136 23612 1192
rect 6315 1020 6371 1076
rect 6425 1020 6481 1076
rect 6535 1020 6591 1076
rect 6645 1020 6701 1076
rect 6755 1020 6811 1076
rect 6865 1020 6921 1076
rect 6975 1020 7031 1076
rect 22896 1026 22952 1082
rect 23006 1026 23062 1082
rect 23116 1026 23172 1082
rect 23226 1026 23282 1082
rect 23336 1026 23392 1082
rect 23446 1026 23502 1082
rect 23556 1026 23612 1082
rect 6315 910 6371 966
rect 6425 910 6481 966
rect 6535 910 6591 966
rect 6645 910 6701 966
rect 6755 910 6811 966
rect 6865 910 6921 966
rect 6975 910 7031 966
rect 22896 916 22952 972
rect 23006 916 23062 972
rect 23116 916 23172 972
rect 23226 916 23282 972
rect 23336 916 23392 972
rect 23446 916 23502 972
rect 23556 916 23612 972
rect 6315 800 6371 856
rect 6425 800 6481 856
rect 6535 800 6591 856
rect 6645 800 6701 856
rect 6755 800 6811 856
rect 6865 800 6921 856
rect 6975 800 7031 856
rect 22896 806 22952 862
rect 23006 806 23062 862
rect 23116 806 23172 862
rect 23226 806 23282 862
rect 23336 806 23392 862
rect 23446 806 23502 862
rect 23556 806 23612 862
rect 6315 690 6371 746
rect 6425 690 6481 746
rect 6535 690 6591 746
rect 6645 690 6701 746
rect 6755 690 6811 746
rect 6865 690 6921 746
rect 6975 690 7031 746
rect 22896 696 22952 752
rect 23006 696 23062 752
rect 23116 696 23172 752
rect 23226 696 23282 752
rect 23336 696 23392 752
rect 23446 696 23502 752
rect 23556 696 23612 752
rect 6315 580 6371 636
rect 6425 580 6481 636
rect 6535 580 6591 636
rect 6645 580 6701 636
rect 6755 580 6811 636
rect 6865 580 6921 636
rect 6975 580 7031 636
rect 22896 586 22952 642
rect 23006 586 23062 642
rect 23116 586 23172 642
rect 23226 586 23282 642
rect 23336 586 23392 642
rect 23446 586 23502 642
rect 23556 586 23612 642
rect 28369 1132 28425 1188
rect 28479 1132 28535 1188
rect 28589 1132 28645 1188
rect 28699 1132 28755 1188
rect 28809 1132 28865 1188
rect 28919 1132 28975 1188
rect 29029 1132 29085 1188
rect 28369 1022 28425 1078
rect 28479 1022 28535 1078
rect 28589 1022 28645 1078
rect 28699 1022 28755 1078
rect 28809 1022 28865 1078
rect 28919 1022 28975 1078
rect 29029 1022 29085 1078
rect 28369 912 28425 968
rect 28479 912 28535 968
rect 28589 912 28645 968
rect 28699 912 28755 968
rect 28809 912 28865 968
rect 28919 912 28975 968
rect 29029 912 29085 968
rect 28369 802 28425 858
rect 28479 802 28535 858
rect 28589 802 28645 858
rect 28699 802 28755 858
rect 28809 802 28865 858
rect 28919 802 28975 858
rect 29029 802 29085 858
rect 28369 692 28425 748
rect 28479 692 28535 748
rect 28589 692 28645 748
rect 28699 692 28755 748
rect 28809 692 28865 748
rect 28919 692 28975 748
rect 29029 692 29085 748
rect 28369 582 28425 638
rect 28479 582 28535 638
rect 28589 582 28645 638
rect 28699 582 28755 638
rect 28809 582 28865 638
rect 28919 582 28975 638
rect 29029 582 29085 638
rect 116770 6864 116826 6920
rect 107204 6728 107260 6784
rect 107314 6728 107370 6784
rect 107424 6728 107480 6784
rect 107534 6728 107590 6784
rect 107644 6728 107700 6784
rect 107754 6728 107810 6784
rect 107864 6728 107920 6784
rect 107204 6618 107260 6674
rect 107314 6618 107370 6674
rect 107424 6618 107480 6674
rect 107534 6618 107590 6674
rect 107644 6618 107700 6674
rect 107754 6618 107810 6674
rect 107864 6618 107920 6674
rect 107204 6508 107260 6564
rect 107314 6508 107370 6564
rect 107424 6508 107480 6564
rect 107534 6508 107590 6564
rect 107644 6508 107700 6564
rect 107754 6508 107810 6564
rect 107864 6508 107920 6564
rect 107204 6398 107260 6454
rect 107314 6398 107370 6454
rect 107424 6398 107480 6454
rect 107534 6398 107590 6454
rect 107644 6398 107700 6454
rect 107754 6398 107810 6454
rect 107864 6398 107920 6454
rect 107204 6288 107260 6344
rect 107314 6288 107370 6344
rect 107424 6288 107480 6344
rect 107534 6288 107590 6344
rect 107644 6288 107700 6344
rect 107754 6288 107810 6344
rect 107864 6288 107920 6344
rect 116770 6754 116826 6810
rect 116770 6644 116826 6700
rect 116770 6534 116826 6590
rect 116770 6424 116826 6480
rect 116770 6314 116826 6370
rect 107204 6178 107260 6234
rect 107314 6178 107370 6234
rect 107424 6178 107480 6234
rect 107534 6178 107590 6234
rect 107644 6178 107700 6234
rect 107754 6178 107810 6234
rect 107864 6178 107920 6234
rect 107204 6068 107260 6124
rect 107314 6068 107370 6124
rect 107424 6068 107480 6124
rect 107534 6068 107590 6124
rect 107644 6068 107700 6124
rect 107754 6068 107810 6124
rect 107864 6068 107920 6124
rect 107204 5958 107260 6014
rect 107314 5958 107370 6014
rect 107424 5958 107480 6014
rect 107534 5958 107590 6014
rect 107644 5958 107700 6014
rect 107754 5958 107810 6014
rect 107864 5958 107920 6014
rect 116770 5444 116826 5500
rect 116770 5334 116826 5390
rect 116770 5224 116826 5280
rect 129259 5277 129315 5333
rect 129369 5277 129425 5333
rect 130585 5282 130641 5338
rect 130695 5282 130751 5338
rect 116770 5114 116826 5170
rect 116770 5004 116826 5060
rect 116770 4894 116826 4950
rect 24709 103 24765 159
rect 24819 103 24875 159
rect 24929 103 24985 159
rect 25039 103 25095 159
rect 25149 103 25205 159
rect 25259 103 25315 159
rect 25369 103 25425 159
rect 29849 158 29905 214
rect 29959 158 30015 214
rect 30069 158 30125 214
rect 30179 158 30235 214
rect 30289 158 30345 214
rect 30399 158 30455 214
rect 30509 158 30565 214
rect 113565 155 113621 211
rect 113675 155 113731 211
rect 113785 155 113841 211
rect 113895 155 113951 211
rect 114005 155 114061 211
rect 114115 155 114171 211
rect 114225 155 114281 211
rect 24709 -7 24765 49
rect 24819 -7 24875 49
rect 24929 -7 24985 49
rect 25039 -7 25095 49
rect 25149 -7 25205 49
rect 25259 -7 25315 49
rect 25369 -7 25425 49
rect 29849 48 29905 104
rect 29959 48 30015 104
rect 30069 48 30125 104
rect 30179 48 30235 104
rect 30289 48 30345 104
rect 30399 48 30455 104
rect 30509 48 30565 104
rect 69220 47 69276 103
rect 69330 47 69386 103
rect 69440 47 69496 103
rect 69550 47 69606 103
rect 69660 47 69716 103
rect 69770 47 69826 103
rect 69880 47 69936 103
rect 71847 52 71903 108
rect 71957 52 72013 108
rect 72067 52 72123 108
rect 72177 52 72233 108
rect 72287 52 72343 108
rect 72397 52 72453 108
rect 72507 52 72563 108
rect 74565 58 74621 114
rect 74675 58 74731 114
rect 74785 58 74841 114
rect 74895 58 74951 114
rect 75005 58 75061 114
rect 75115 58 75171 114
rect 75225 58 75281 114
rect 77637 44 77693 100
rect 77747 44 77803 100
rect 77857 44 77913 100
rect 77967 44 78023 100
rect 78077 44 78133 100
rect 78187 44 78243 100
rect 78297 44 78353 100
rect 80687 53 80743 109
rect 80797 53 80853 109
rect 80907 53 80963 109
rect 81017 53 81073 109
rect 81127 53 81183 109
rect 81237 53 81293 109
rect 81347 53 81403 109
rect 83528 53 83584 109
rect 83638 53 83694 109
rect 83748 53 83804 109
rect 83858 53 83914 109
rect 83968 53 84024 109
rect 84078 53 84134 109
rect 84188 53 84244 109
rect 86316 50 86372 106
rect 86426 50 86482 106
rect 86536 50 86592 106
rect 86646 50 86702 106
rect 86756 50 86812 106
rect 86866 50 86922 106
rect 86976 50 87032 106
rect 89511 62 89567 118
rect 89621 62 89677 118
rect 89731 62 89787 118
rect 89841 62 89897 118
rect 89951 62 90007 118
rect 90061 62 90117 118
rect 90171 62 90227 118
rect 92852 51 92908 107
rect 92962 51 93018 107
rect 93072 51 93128 107
rect 93182 51 93238 107
rect 93292 51 93348 107
rect 93402 51 93458 107
rect 93512 51 93568 107
rect 95994 54 96050 110
rect 96104 54 96160 110
rect 96214 54 96270 110
rect 96324 54 96380 110
rect 96434 54 96490 110
rect 96544 54 96600 110
rect 96654 54 96710 110
rect 99280 52 99336 108
rect 99390 52 99446 108
rect 99500 52 99556 108
rect 99610 52 99666 108
rect 99720 52 99776 108
rect 99830 52 99886 108
rect 99940 52 99996 108
rect 113565 45 113621 101
rect 113675 45 113731 101
rect 113785 45 113841 101
rect 113895 45 113951 101
rect 114005 45 114061 101
rect 114115 45 114171 101
rect 114225 45 114281 101
rect 24709 -117 24765 -61
rect 24819 -117 24875 -61
rect 24929 -117 24985 -61
rect 25039 -117 25095 -61
rect 25149 -117 25205 -61
rect 25259 -117 25315 -61
rect 25369 -117 25425 -61
rect 29849 -62 29905 -6
rect 29959 -62 30015 -6
rect 30069 -62 30125 -6
rect 30179 -62 30235 -6
rect 30289 -62 30345 -6
rect 30399 -62 30455 -6
rect 30509 -62 30565 -6
rect 69220 -63 69276 -7
rect 69330 -63 69386 -7
rect 69440 -63 69496 -7
rect 69550 -63 69606 -7
rect 69660 -63 69716 -7
rect 69770 -63 69826 -7
rect 69880 -63 69936 -7
rect 71847 -58 71903 -2
rect 71957 -58 72013 -2
rect 72067 -58 72123 -2
rect 72177 -58 72233 -2
rect 72287 -58 72343 -2
rect 72397 -58 72453 -2
rect 72507 -58 72563 -2
rect 74565 -52 74621 4
rect 74675 -52 74731 4
rect 74785 -52 74841 4
rect 74895 -52 74951 4
rect 75005 -52 75061 4
rect 75115 -52 75171 4
rect 75225 -52 75281 4
rect 77637 -66 77693 -10
rect 77747 -66 77803 -10
rect 77857 -66 77913 -10
rect 77967 -66 78023 -10
rect 78077 -66 78133 -10
rect 78187 -66 78243 -10
rect 78297 -66 78353 -10
rect 80687 -57 80743 -1
rect 80797 -57 80853 -1
rect 80907 -57 80963 -1
rect 81017 -57 81073 -1
rect 81127 -57 81183 -1
rect 81237 -57 81293 -1
rect 81347 -57 81403 -1
rect 83528 -57 83584 -1
rect 83638 -57 83694 -1
rect 83748 -57 83804 -1
rect 83858 -57 83914 -1
rect 83968 -57 84024 -1
rect 84078 -57 84134 -1
rect 84188 -57 84244 -1
rect 86316 -60 86372 -4
rect 86426 -60 86482 -4
rect 86536 -60 86592 -4
rect 86646 -60 86702 -4
rect 86756 -60 86812 -4
rect 86866 -60 86922 -4
rect 86976 -60 87032 -4
rect 89511 -48 89567 8
rect 89621 -48 89677 8
rect 89731 -48 89787 8
rect 89841 -48 89897 8
rect 89951 -48 90007 8
rect 90061 -48 90117 8
rect 90171 -48 90227 8
rect 92852 -59 92908 -3
rect 92962 -59 93018 -3
rect 93072 -59 93128 -3
rect 93182 -59 93238 -3
rect 93292 -59 93348 -3
rect 93402 -59 93458 -3
rect 93512 -59 93568 -3
rect 95994 -56 96050 0
rect 96104 -56 96160 0
rect 96214 -56 96270 0
rect 96324 -56 96380 0
rect 96434 -56 96490 0
rect 96544 -56 96600 0
rect 96654 -56 96710 0
rect 99280 -58 99336 -2
rect 99390 -58 99446 -2
rect 99500 -58 99556 -2
rect 99610 -58 99666 -2
rect 99720 -58 99776 -2
rect 99830 -58 99886 -2
rect 99940 -58 99996 -2
rect 113565 -65 113621 -9
rect 113675 -65 113731 -9
rect 113785 -65 113841 -9
rect 113895 -65 113951 -9
rect 114005 -65 114061 -9
rect 114115 -65 114171 -9
rect 114225 -65 114281 -9
rect 24709 -227 24765 -171
rect 24819 -227 24875 -171
rect 24929 -227 24985 -171
rect 25039 -227 25095 -171
rect 25149 -227 25205 -171
rect 25259 -227 25315 -171
rect 25369 -227 25425 -171
rect 29849 -172 29905 -116
rect 29959 -172 30015 -116
rect 30069 -172 30125 -116
rect 30179 -172 30235 -116
rect 30289 -172 30345 -116
rect 30399 -172 30455 -116
rect 30509 -172 30565 -116
rect 69220 -173 69276 -117
rect 69330 -173 69386 -117
rect 69440 -173 69496 -117
rect 69550 -173 69606 -117
rect 69660 -173 69716 -117
rect 69770 -173 69826 -117
rect 69880 -173 69936 -117
rect 71847 -168 71903 -112
rect 71957 -168 72013 -112
rect 72067 -168 72123 -112
rect 72177 -168 72233 -112
rect 72287 -168 72343 -112
rect 72397 -168 72453 -112
rect 72507 -168 72563 -112
rect 74565 -162 74621 -106
rect 74675 -162 74731 -106
rect 74785 -162 74841 -106
rect 74895 -162 74951 -106
rect 75005 -162 75061 -106
rect 75115 -162 75171 -106
rect 75225 -162 75281 -106
rect 77637 -176 77693 -120
rect 77747 -176 77803 -120
rect 77857 -176 77913 -120
rect 77967 -176 78023 -120
rect 78077 -176 78133 -120
rect 78187 -176 78243 -120
rect 78297 -176 78353 -120
rect 80687 -167 80743 -111
rect 80797 -167 80853 -111
rect 80907 -167 80963 -111
rect 81017 -167 81073 -111
rect 81127 -167 81183 -111
rect 81237 -167 81293 -111
rect 81347 -167 81403 -111
rect 83528 -167 83584 -111
rect 83638 -167 83694 -111
rect 83748 -167 83804 -111
rect 83858 -167 83914 -111
rect 83968 -167 84024 -111
rect 84078 -167 84134 -111
rect 84188 -167 84244 -111
rect 86316 -170 86372 -114
rect 86426 -170 86482 -114
rect 86536 -170 86592 -114
rect 86646 -170 86702 -114
rect 86756 -170 86812 -114
rect 86866 -170 86922 -114
rect 86976 -170 87032 -114
rect 89511 -158 89567 -102
rect 89621 -158 89677 -102
rect 89731 -158 89787 -102
rect 89841 -158 89897 -102
rect 89951 -158 90007 -102
rect 90061 -158 90117 -102
rect 90171 -158 90227 -102
rect 92852 -169 92908 -113
rect 92962 -169 93018 -113
rect 93072 -169 93128 -113
rect 93182 -169 93238 -113
rect 93292 -169 93348 -113
rect 93402 -169 93458 -113
rect 93512 -169 93568 -113
rect 95994 -166 96050 -110
rect 96104 -166 96160 -110
rect 96214 -166 96270 -110
rect 96324 -166 96380 -110
rect 96434 -166 96490 -110
rect 96544 -166 96600 -110
rect 96654 -166 96710 -110
rect 99280 -168 99336 -112
rect 99390 -168 99446 -112
rect 99500 -168 99556 -112
rect 99610 -168 99666 -112
rect 99720 -168 99776 -112
rect 99830 -168 99886 -112
rect 99940 -168 99996 -112
rect 113565 -175 113621 -119
rect 113675 -175 113731 -119
rect 113785 -175 113841 -119
rect 113895 -175 113951 -119
rect 114005 -175 114061 -119
rect 114115 -175 114171 -119
rect 114225 -175 114281 -119
rect 24709 -337 24765 -281
rect 24819 -337 24875 -281
rect 24929 -337 24985 -281
rect 25039 -337 25095 -281
rect 25149 -337 25205 -281
rect 25259 -337 25315 -281
rect 25369 -337 25425 -281
rect 29849 -282 29905 -226
rect 29959 -282 30015 -226
rect 30069 -282 30125 -226
rect 30179 -282 30235 -226
rect 30289 -282 30345 -226
rect 30399 -282 30455 -226
rect 30509 -282 30565 -226
rect 69220 -283 69276 -227
rect 69330 -283 69386 -227
rect 69440 -283 69496 -227
rect 69550 -283 69606 -227
rect 69660 -283 69716 -227
rect 69770 -283 69826 -227
rect 69880 -283 69936 -227
rect 71847 -278 71903 -222
rect 71957 -278 72013 -222
rect 72067 -278 72123 -222
rect 72177 -278 72233 -222
rect 72287 -278 72343 -222
rect 72397 -278 72453 -222
rect 72507 -278 72563 -222
rect 74565 -272 74621 -216
rect 74675 -272 74731 -216
rect 74785 -272 74841 -216
rect 74895 -272 74951 -216
rect 75005 -272 75061 -216
rect 75115 -272 75171 -216
rect 75225 -272 75281 -216
rect 77637 -286 77693 -230
rect 77747 -286 77803 -230
rect 77857 -286 77913 -230
rect 77967 -286 78023 -230
rect 78077 -286 78133 -230
rect 78187 -286 78243 -230
rect 78297 -286 78353 -230
rect 80687 -277 80743 -221
rect 80797 -277 80853 -221
rect 80907 -277 80963 -221
rect 81017 -277 81073 -221
rect 81127 -277 81183 -221
rect 81237 -277 81293 -221
rect 81347 -277 81403 -221
rect 83528 -277 83584 -221
rect 83638 -277 83694 -221
rect 83748 -277 83804 -221
rect 83858 -277 83914 -221
rect 83968 -277 84024 -221
rect 84078 -277 84134 -221
rect 84188 -277 84244 -221
rect 86316 -280 86372 -224
rect 86426 -280 86482 -224
rect 86536 -280 86592 -224
rect 86646 -280 86702 -224
rect 86756 -280 86812 -224
rect 86866 -280 86922 -224
rect 86976 -280 87032 -224
rect 89511 -268 89567 -212
rect 89621 -268 89677 -212
rect 89731 -268 89787 -212
rect 89841 -268 89897 -212
rect 89951 -268 90007 -212
rect 90061 -268 90117 -212
rect 90171 -268 90227 -212
rect 92852 -279 92908 -223
rect 92962 -279 93018 -223
rect 93072 -279 93128 -223
rect 93182 -279 93238 -223
rect 93292 -279 93348 -223
rect 93402 -279 93458 -223
rect 93512 -279 93568 -223
rect 95994 -276 96050 -220
rect 96104 -276 96160 -220
rect 96214 -276 96270 -220
rect 96324 -276 96380 -220
rect 96434 -276 96490 -220
rect 96544 -276 96600 -220
rect 96654 -276 96710 -220
rect 99280 -278 99336 -222
rect 99390 -278 99446 -222
rect 99500 -278 99556 -222
rect 99610 -278 99666 -222
rect 99720 -278 99776 -222
rect 99830 -278 99886 -222
rect 99940 -278 99996 -222
rect 113565 -285 113621 -229
rect 113675 -285 113731 -229
rect 113785 -285 113841 -229
rect 113895 -285 113951 -229
rect 114005 -285 114061 -229
rect 114115 -285 114171 -229
rect 114225 -285 114281 -229
rect 24709 -447 24765 -391
rect 24819 -447 24875 -391
rect 24929 -447 24985 -391
rect 25039 -447 25095 -391
rect 25149 -447 25205 -391
rect 25259 -447 25315 -391
rect 25369 -447 25425 -391
rect 29849 -392 29905 -336
rect 29959 -392 30015 -336
rect 30069 -392 30125 -336
rect 30179 -392 30235 -336
rect 30289 -392 30345 -336
rect 30399 -392 30455 -336
rect 30509 -392 30565 -336
rect 69220 -393 69276 -337
rect 69330 -393 69386 -337
rect 69440 -393 69496 -337
rect 69550 -393 69606 -337
rect 69660 -393 69716 -337
rect 69770 -393 69826 -337
rect 69880 -393 69936 -337
rect 71847 -388 71903 -332
rect 71957 -388 72013 -332
rect 72067 -388 72123 -332
rect 72177 -388 72233 -332
rect 72287 -388 72343 -332
rect 72397 -388 72453 -332
rect 72507 -388 72563 -332
rect 74565 -382 74621 -326
rect 74675 -382 74731 -326
rect 74785 -382 74841 -326
rect 74895 -382 74951 -326
rect 75005 -382 75061 -326
rect 75115 -382 75171 -326
rect 75225 -382 75281 -326
rect 77637 -396 77693 -340
rect 77747 -396 77803 -340
rect 77857 -396 77913 -340
rect 77967 -396 78023 -340
rect 78077 -396 78133 -340
rect 78187 -396 78243 -340
rect 78297 -396 78353 -340
rect 80687 -387 80743 -331
rect 80797 -387 80853 -331
rect 80907 -387 80963 -331
rect 81017 -387 81073 -331
rect 81127 -387 81183 -331
rect 81237 -387 81293 -331
rect 81347 -387 81403 -331
rect 83528 -387 83584 -331
rect 83638 -387 83694 -331
rect 83748 -387 83804 -331
rect 83858 -387 83914 -331
rect 83968 -387 84024 -331
rect 84078 -387 84134 -331
rect 84188 -387 84244 -331
rect 86316 -390 86372 -334
rect 86426 -390 86482 -334
rect 86536 -390 86592 -334
rect 86646 -390 86702 -334
rect 86756 -390 86812 -334
rect 86866 -390 86922 -334
rect 86976 -390 87032 -334
rect 89511 -378 89567 -322
rect 89621 -378 89677 -322
rect 89731 -378 89787 -322
rect 89841 -378 89897 -322
rect 89951 -378 90007 -322
rect 90061 -378 90117 -322
rect 90171 -378 90227 -322
rect 92852 -389 92908 -333
rect 92962 -389 93018 -333
rect 93072 -389 93128 -333
rect 93182 -389 93238 -333
rect 93292 -389 93348 -333
rect 93402 -389 93458 -333
rect 93512 -389 93568 -333
rect 95994 -386 96050 -330
rect 96104 -386 96160 -330
rect 96214 -386 96270 -330
rect 96324 -386 96380 -330
rect 96434 -386 96490 -330
rect 96544 -386 96600 -330
rect 96654 -386 96710 -330
rect 99280 -388 99336 -332
rect 99390 -388 99446 -332
rect 99500 -388 99556 -332
rect 99610 -388 99666 -332
rect 99720 -388 99776 -332
rect 99830 -388 99886 -332
rect 99940 -388 99996 -332
rect 113565 -395 113621 -339
rect 113675 -395 113731 -339
rect 113785 -395 113841 -339
rect 113895 -395 113951 -339
rect 114005 -395 114061 -339
rect 114115 -395 114171 -339
rect 114225 -395 114281 -339
rect 69220 -503 69276 -447
rect 69330 -503 69386 -447
rect 69440 -503 69496 -447
rect 69550 -503 69606 -447
rect 69660 -503 69716 -447
rect 69770 -503 69826 -447
rect 69880 -503 69936 -447
rect 71847 -498 71903 -442
rect 71957 -498 72013 -442
rect 72067 -498 72123 -442
rect 72177 -498 72233 -442
rect 72287 -498 72343 -442
rect 72397 -498 72453 -442
rect 72507 -498 72563 -442
rect 74565 -492 74621 -436
rect 74675 -492 74731 -436
rect 74785 -492 74841 -436
rect 74895 -492 74951 -436
rect 75005 -492 75061 -436
rect 75115 -492 75171 -436
rect 75225 -492 75281 -436
rect 77637 -506 77693 -450
rect 77747 -506 77803 -450
rect 77857 -506 77913 -450
rect 77967 -506 78023 -450
rect 78077 -506 78133 -450
rect 78187 -506 78243 -450
rect 78297 -506 78353 -450
rect 80687 -497 80743 -441
rect 80797 -497 80853 -441
rect 80907 -497 80963 -441
rect 81017 -497 81073 -441
rect 81127 -497 81183 -441
rect 81237 -497 81293 -441
rect 81347 -497 81403 -441
rect 83528 -497 83584 -441
rect 83638 -497 83694 -441
rect 83748 -497 83804 -441
rect 83858 -497 83914 -441
rect 83968 -497 84024 -441
rect 84078 -497 84134 -441
rect 84188 -497 84244 -441
rect 86316 -500 86372 -444
rect 86426 -500 86482 -444
rect 86536 -500 86592 -444
rect 86646 -500 86702 -444
rect 86756 -500 86812 -444
rect 86866 -500 86922 -444
rect 86976 -500 87032 -444
rect 89511 -488 89567 -432
rect 89621 -488 89677 -432
rect 89731 -488 89787 -432
rect 89841 -488 89897 -432
rect 89951 -488 90007 -432
rect 90061 -488 90117 -432
rect 90171 -488 90227 -432
rect 92852 -499 92908 -443
rect 92962 -499 93018 -443
rect 93072 -499 93128 -443
rect 93182 -499 93238 -443
rect 93292 -499 93348 -443
rect 93402 -499 93458 -443
rect 93512 -499 93568 -443
rect 95994 -496 96050 -440
rect 96104 -496 96160 -440
rect 96214 -496 96270 -440
rect 96324 -496 96380 -440
rect 96434 -496 96490 -440
rect 96544 -496 96600 -440
rect 96654 -496 96710 -440
rect 99280 -498 99336 -442
rect 99390 -498 99446 -442
rect 99500 -498 99556 -442
rect 99610 -498 99666 -442
rect 99720 -498 99776 -442
rect 99830 -498 99886 -442
rect 99940 -498 99996 -442
rect 5544 -1640 5600 -1584
rect 5654 -1640 5710 -1584
rect 5764 -1640 5820 -1584
rect 5874 -1640 5930 -1584
rect 5544 -1750 5600 -1694
rect 5654 -1750 5710 -1694
rect 5764 -1750 5820 -1694
rect 5874 -1750 5930 -1694
rect 5544 -1860 5600 -1804
rect 5654 -1860 5710 -1804
rect 5764 -1860 5820 -1804
rect 5874 -1860 5930 -1804
rect 5544 -1970 5600 -1914
rect 5654 -1970 5710 -1914
rect 5764 -1970 5820 -1914
rect 5874 -1970 5930 -1914
rect 138 -2237 194 -2181
rect 248 -2237 304 -2181
rect 358 -2237 414 -2181
rect 468 -2237 524 -2181
rect 578 -2237 634 -2181
rect 688 -2237 744 -2181
rect 798 -2237 854 -2181
rect 138 -2347 194 -2291
rect 248 -2347 304 -2291
rect 358 -2347 414 -2291
rect 468 -2347 524 -2291
rect 578 -2347 634 -2291
rect 688 -2347 744 -2291
rect 798 -2347 854 -2291
rect 138 -2457 194 -2401
rect 248 -2457 304 -2401
rect 358 -2457 414 -2401
rect 468 -2457 524 -2401
rect 578 -2457 634 -2401
rect 688 -2457 744 -2401
rect 798 -2457 854 -2401
rect 138 -2567 194 -2511
rect 248 -2567 304 -2511
rect 358 -2567 414 -2511
rect 468 -2567 524 -2511
rect 578 -2567 634 -2511
rect 688 -2567 744 -2511
rect 798 -2567 854 -2511
rect 138 -2677 194 -2621
rect 248 -2677 304 -2621
rect 358 -2677 414 -2621
rect 468 -2677 524 -2621
rect 578 -2677 634 -2621
rect 688 -2677 744 -2621
rect 798 -2677 854 -2621
rect 138 -2787 194 -2731
rect 248 -2787 304 -2731
rect 358 -2787 414 -2731
rect 468 -2787 524 -2731
rect 578 -2787 634 -2731
rect 688 -2787 744 -2731
rect 798 -2787 854 -2731
rect 10881 -1184 10937 -1128
rect 10991 -1184 11047 -1128
rect 11101 -1184 11157 -1128
rect 11211 -1184 11267 -1128
rect 11321 -1184 11377 -1128
rect 11431 -1184 11487 -1128
rect 11541 -1184 11597 -1128
rect 11670 -1184 11726 -1128
rect 11780 -1184 11836 -1128
rect 11890 -1184 11946 -1128
rect 12000 -1184 12056 -1128
rect 12110 -1184 12166 -1128
rect 12220 -1184 12276 -1128
rect 12330 -1184 12386 -1128
rect 25927 -1202 25983 -1146
rect 26037 -1202 26093 -1146
rect 26147 -1202 26203 -1146
rect 26257 -1202 26313 -1146
rect 26367 -1202 26423 -1146
rect 26477 -1202 26533 -1146
rect 26587 -1202 26643 -1146
rect 10881 -1294 10937 -1238
rect 10991 -1294 11047 -1238
rect 11101 -1294 11157 -1238
rect 11211 -1294 11267 -1238
rect 11321 -1294 11377 -1238
rect 11431 -1294 11487 -1238
rect 11541 -1294 11597 -1238
rect 11670 -1294 11726 -1238
rect 11780 -1294 11836 -1238
rect 11890 -1294 11946 -1238
rect 12000 -1294 12056 -1238
rect 12110 -1294 12166 -1238
rect 12220 -1294 12276 -1238
rect 12330 -1294 12386 -1238
rect 114635 -1255 114691 -1199
rect 114745 -1255 114801 -1199
rect 114855 -1255 114911 -1199
rect 114965 -1255 115021 -1199
rect 115075 -1255 115131 -1199
rect 115185 -1255 115241 -1199
rect 115295 -1255 115351 -1199
rect 25927 -1312 25983 -1256
rect 26037 -1312 26093 -1256
rect 26147 -1312 26203 -1256
rect 26257 -1312 26313 -1256
rect 26367 -1312 26423 -1256
rect 26477 -1312 26533 -1256
rect 26587 -1312 26643 -1256
rect 10881 -1404 10937 -1348
rect 10991 -1404 11047 -1348
rect 11101 -1404 11157 -1348
rect 11211 -1404 11267 -1348
rect 11321 -1404 11377 -1348
rect 11431 -1404 11487 -1348
rect 11541 -1404 11597 -1348
rect 11670 -1404 11726 -1348
rect 11780 -1404 11836 -1348
rect 11890 -1404 11946 -1348
rect 12000 -1404 12056 -1348
rect 12110 -1404 12166 -1348
rect 12220 -1404 12276 -1348
rect 12330 -1404 12386 -1348
rect 114635 -1365 114691 -1309
rect 114745 -1365 114801 -1309
rect 114855 -1365 114911 -1309
rect 114965 -1365 115021 -1309
rect 115075 -1365 115131 -1309
rect 115185 -1365 115241 -1309
rect 115295 -1365 115351 -1309
rect 25927 -1422 25983 -1366
rect 26037 -1422 26093 -1366
rect 26147 -1422 26203 -1366
rect 26257 -1422 26313 -1366
rect 26367 -1422 26423 -1366
rect 26477 -1422 26533 -1366
rect 26587 -1422 26643 -1366
rect 10881 -1514 10937 -1458
rect 10991 -1514 11047 -1458
rect 11101 -1514 11157 -1458
rect 11211 -1514 11267 -1458
rect 11321 -1514 11377 -1458
rect 11431 -1514 11487 -1458
rect 11541 -1514 11597 -1458
rect 11670 -1514 11726 -1458
rect 11780 -1514 11836 -1458
rect 11890 -1514 11946 -1458
rect 12000 -1514 12056 -1458
rect 12110 -1514 12166 -1458
rect 12220 -1514 12276 -1458
rect 12330 -1514 12386 -1458
rect 114635 -1475 114691 -1419
rect 114745 -1475 114801 -1419
rect 114855 -1475 114911 -1419
rect 114965 -1475 115021 -1419
rect 115075 -1475 115131 -1419
rect 115185 -1475 115241 -1419
rect 115295 -1475 115351 -1419
rect 25927 -1532 25983 -1476
rect 26037 -1532 26093 -1476
rect 26147 -1532 26203 -1476
rect 26257 -1532 26313 -1476
rect 26367 -1532 26423 -1476
rect 26477 -1532 26533 -1476
rect 26587 -1532 26643 -1476
rect 10881 -1624 10937 -1568
rect 10991 -1624 11047 -1568
rect 11101 -1624 11157 -1568
rect 11211 -1624 11267 -1568
rect 11321 -1624 11377 -1568
rect 11431 -1624 11487 -1568
rect 11541 -1624 11597 -1568
rect 11670 -1624 11726 -1568
rect 11780 -1624 11836 -1568
rect 11890 -1624 11946 -1568
rect 12000 -1624 12056 -1568
rect 12110 -1624 12166 -1568
rect 12220 -1624 12276 -1568
rect 12330 -1624 12386 -1568
rect 114635 -1585 114691 -1529
rect 114745 -1585 114801 -1529
rect 114855 -1585 114911 -1529
rect 114965 -1585 115021 -1529
rect 115075 -1585 115131 -1529
rect 115185 -1585 115241 -1529
rect 115295 -1585 115351 -1529
rect 25927 -1642 25983 -1586
rect 26037 -1642 26093 -1586
rect 26147 -1642 26203 -1586
rect 26257 -1642 26313 -1586
rect 26367 -1642 26423 -1586
rect 26477 -1642 26533 -1586
rect 26587 -1642 26643 -1586
rect 10881 -1734 10937 -1678
rect 10991 -1734 11047 -1678
rect 11101 -1734 11157 -1678
rect 11211 -1734 11267 -1678
rect 11321 -1734 11377 -1678
rect 11431 -1734 11487 -1678
rect 11541 -1734 11597 -1678
rect 11670 -1734 11726 -1678
rect 11780 -1734 11836 -1678
rect 11890 -1734 11946 -1678
rect 12000 -1734 12056 -1678
rect 12110 -1734 12166 -1678
rect 12220 -1734 12276 -1678
rect 12330 -1734 12386 -1678
rect 114635 -1695 114691 -1639
rect 114745 -1695 114801 -1639
rect 114855 -1695 114911 -1639
rect 114965 -1695 115021 -1639
rect 115075 -1695 115131 -1639
rect 115185 -1695 115241 -1639
rect 115295 -1695 115351 -1639
rect 25927 -1752 25983 -1696
rect 26037 -1752 26093 -1696
rect 26147 -1752 26203 -1696
rect 26257 -1752 26313 -1696
rect 26367 -1752 26423 -1696
rect 26477 -1752 26533 -1696
rect 26587 -1752 26643 -1696
rect 114635 -1805 114691 -1749
rect 114745 -1805 114801 -1749
rect 114855 -1805 114911 -1749
rect 114965 -1805 115021 -1749
rect 115075 -1805 115131 -1749
rect 115185 -1805 115241 -1749
rect 115295 -1805 115351 -1749
rect 29884 -2276 29940 -2220
rect 29994 -2276 30050 -2220
rect 30104 -2276 30160 -2220
rect 30214 -2276 30270 -2220
rect 30324 -2276 30380 -2220
rect 30434 -2276 30490 -2220
rect 30544 -2276 30600 -2220
rect 113560 -2345 113616 -2289
rect 113670 -2345 113726 -2289
rect 113780 -2345 113836 -2289
rect 113890 -2345 113946 -2289
rect 114000 -2345 114056 -2289
rect 114110 -2345 114166 -2289
rect 114220 -2345 114276 -2289
rect 113560 -2455 113616 -2399
rect 113670 -2455 113726 -2399
rect 113780 -2455 113836 -2399
rect 113890 -2455 113946 -2399
rect 114000 -2455 114056 -2399
rect 114110 -2455 114166 -2399
rect 114220 -2455 114276 -2399
rect 113560 -2565 113616 -2509
rect 113670 -2565 113726 -2509
rect 113780 -2565 113836 -2509
rect 113890 -2565 113946 -2509
rect 114000 -2565 114056 -2509
rect 114110 -2565 114166 -2509
rect 114220 -2565 114276 -2509
rect 113560 -2675 113616 -2619
rect 113670 -2675 113726 -2619
rect 113780 -2675 113836 -2619
rect 113890 -2675 113946 -2619
rect 114000 -2675 114056 -2619
rect 114110 -2675 114166 -2619
rect 114220 -2675 114276 -2619
rect 113560 -2785 113616 -2729
rect 113670 -2785 113726 -2729
rect 113780 -2785 113836 -2729
rect 113890 -2785 113946 -2729
rect 114000 -2785 114056 -2729
rect 114110 -2785 114166 -2729
rect 114220 -2785 114276 -2729
rect 113560 -2895 113616 -2839
rect 113670 -2895 113726 -2839
rect 113780 -2895 113836 -2839
rect 113890 -2895 113946 -2839
rect 114000 -2895 114056 -2839
rect 114110 -2895 114166 -2839
rect 114220 -2895 114276 -2839
rect 69250 -3381 69306 -3325
rect 69360 -3381 69416 -3325
rect 69470 -3381 69526 -3325
rect 69580 -3381 69636 -3325
rect 69690 -3381 69746 -3325
rect 69800 -3381 69856 -3325
rect 69910 -3381 69966 -3325
rect 69250 -3491 69306 -3435
rect 69360 -3491 69416 -3435
rect 69470 -3491 69526 -3435
rect 69580 -3491 69636 -3435
rect 69690 -3491 69746 -3435
rect 69800 -3491 69856 -3435
rect 69910 -3491 69966 -3435
rect 69250 -3601 69306 -3545
rect 69360 -3601 69416 -3545
rect 69470 -3601 69526 -3545
rect 69580 -3601 69636 -3545
rect 69690 -3601 69746 -3545
rect 69800 -3601 69856 -3545
rect 69910 -3601 69966 -3545
rect 69250 -3711 69306 -3655
rect 69360 -3711 69416 -3655
rect 69470 -3711 69526 -3655
rect 69580 -3711 69636 -3655
rect 69690 -3711 69746 -3655
rect 69800 -3711 69856 -3655
rect 69910 -3711 69966 -3655
rect 69250 -3821 69306 -3765
rect 69360 -3821 69416 -3765
rect 69470 -3821 69526 -3765
rect 69580 -3821 69636 -3765
rect 69690 -3821 69746 -3765
rect 69800 -3821 69856 -3765
rect 69910 -3821 69966 -3765
rect 69250 -3931 69306 -3875
rect 69360 -3931 69416 -3875
rect 69470 -3931 69526 -3875
rect 69580 -3931 69636 -3875
rect 69690 -3931 69746 -3875
rect 69800 -3931 69856 -3875
rect 69910 -3931 69966 -3875
rect 71863 -3444 71919 -3388
rect 71973 -3444 72029 -3388
rect 72083 -3444 72139 -3388
rect 72193 -3444 72249 -3388
rect 72303 -3444 72359 -3388
rect 72413 -3444 72469 -3388
rect 72523 -3444 72579 -3388
rect 71863 -3554 71919 -3498
rect 71973 -3554 72029 -3498
rect 72083 -3554 72139 -3498
rect 72193 -3554 72249 -3498
rect 72303 -3554 72359 -3498
rect 72413 -3554 72469 -3498
rect 72523 -3554 72579 -3498
rect 71863 -3664 71919 -3608
rect 71973 -3664 72029 -3608
rect 72083 -3664 72139 -3608
rect 72193 -3664 72249 -3608
rect 72303 -3664 72359 -3608
rect 72413 -3664 72469 -3608
rect 72523 -3664 72579 -3608
rect 71863 -3774 71919 -3718
rect 71973 -3774 72029 -3718
rect 72083 -3774 72139 -3718
rect 72193 -3774 72249 -3718
rect 72303 -3774 72359 -3718
rect 72413 -3774 72469 -3718
rect 72523 -3774 72579 -3718
rect 71863 -3884 71919 -3828
rect 71973 -3884 72029 -3828
rect 72083 -3884 72139 -3828
rect 72193 -3884 72249 -3828
rect 72303 -3884 72359 -3828
rect 72413 -3884 72469 -3828
rect 72523 -3884 72579 -3828
rect 71863 -3994 71919 -3938
rect 71973 -3994 72029 -3938
rect 72083 -3994 72139 -3938
rect 72193 -3994 72249 -3938
rect 72303 -3994 72359 -3938
rect 72413 -3994 72469 -3938
rect 72523 -3994 72579 -3938
rect 74577 -3466 74633 -3410
rect 74687 -3466 74743 -3410
rect 74797 -3466 74853 -3410
rect 74907 -3466 74963 -3410
rect 75017 -3466 75073 -3410
rect 75127 -3466 75183 -3410
rect 75237 -3466 75293 -3410
rect 74577 -3576 74633 -3520
rect 74687 -3576 74743 -3520
rect 74797 -3576 74853 -3520
rect 74907 -3576 74963 -3520
rect 75017 -3576 75073 -3520
rect 75127 -3576 75183 -3520
rect 75237 -3576 75293 -3520
rect 74577 -3686 74633 -3630
rect 74687 -3686 74743 -3630
rect 74797 -3686 74853 -3630
rect 74907 -3686 74963 -3630
rect 75017 -3686 75073 -3630
rect 75127 -3686 75183 -3630
rect 75237 -3686 75293 -3630
rect 74577 -3796 74633 -3740
rect 74687 -3796 74743 -3740
rect 74797 -3796 74853 -3740
rect 74907 -3796 74963 -3740
rect 75017 -3796 75073 -3740
rect 75127 -3796 75183 -3740
rect 75237 -3796 75293 -3740
rect 74577 -3906 74633 -3850
rect 74687 -3906 74743 -3850
rect 74797 -3906 74853 -3850
rect 74907 -3906 74963 -3850
rect 75017 -3906 75073 -3850
rect 75127 -3906 75183 -3850
rect 75237 -3906 75293 -3850
rect 74577 -4016 74633 -3960
rect 74687 -4016 74743 -3960
rect 74797 -4016 74853 -3960
rect 74907 -4016 74963 -3960
rect 75017 -4016 75073 -3960
rect 75127 -4016 75183 -3960
rect 75237 -4016 75293 -3960
rect 77645 -3440 77701 -3384
rect 77755 -3440 77811 -3384
rect 77865 -3440 77921 -3384
rect 77975 -3440 78031 -3384
rect 78085 -3440 78141 -3384
rect 78195 -3440 78251 -3384
rect 78305 -3440 78361 -3384
rect 77645 -3550 77701 -3494
rect 77755 -3550 77811 -3494
rect 77865 -3550 77921 -3494
rect 77975 -3550 78031 -3494
rect 78085 -3550 78141 -3494
rect 78195 -3550 78251 -3494
rect 78305 -3550 78361 -3494
rect 77645 -3660 77701 -3604
rect 77755 -3660 77811 -3604
rect 77865 -3660 77921 -3604
rect 77975 -3660 78031 -3604
rect 78085 -3660 78141 -3604
rect 78195 -3660 78251 -3604
rect 78305 -3660 78361 -3604
rect 77645 -3770 77701 -3714
rect 77755 -3770 77811 -3714
rect 77865 -3770 77921 -3714
rect 77975 -3770 78031 -3714
rect 78085 -3770 78141 -3714
rect 78195 -3770 78251 -3714
rect 78305 -3770 78361 -3714
rect 77645 -3880 77701 -3824
rect 77755 -3880 77811 -3824
rect 77865 -3880 77921 -3824
rect 77975 -3880 78031 -3824
rect 78085 -3880 78141 -3824
rect 78195 -3880 78251 -3824
rect 78305 -3880 78361 -3824
rect 77645 -3990 77701 -3934
rect 77755 -3990 77811 -3934
rect 77865 -3990 77921 -3934
rect 77975 -3990 78031 -3934
rect 78085 -3990 78141 -3934
rect 78195 -3990 78251 -3934
rect 78305 -3990 78361 -3934
rect 80699 -3412 80755 -3356
rect 80809 -3412 80865 -3356
rect 80919 -3412 80975 -3356
rect 81029 -3412 81085 -3356
rect 81139 -3412 81195 -3356
rect 81249 -3412 81305 -3356
rect 81359 -3412 81415 -3356
rect 80699 -3522 80755 -3466
rect 80809 -3522 80865 -3466
rect 80919 -3522 80975 -3466
rect 81029 -3522 81085 -3466
rect 81139 -3522 81195 -3466
rect 81249 -3522 81305 -3466
rect 81359 -3522 81415 -3466
rect 80699 -3632 80755 -3576
rect 80809 -3632 80865 -3576
rect 80919 -3632 80975 -3576
rect 81029 -3632 81085 -3576
rect 81139 -3632 81195 -3576
rect 81249 -3632 81305 -3576
rect 81359 -3632 81415 -3576
rect 80699 -3742 80755 -3686
rect 80809 -3742 80865 -3686
rect 80919 -3742 80975 -3686
rect 81029 -3742 81085 -3686
rect 81139 -3742 81195 -3686
rect 81249 -3742 81305 -3686
rect 81359 -3742 81415 -3686
rect 80699 -3852 80755 -3796
rect 80809 -3852 80865 -3796
rect 80919 -3852 80975 -3796
rect 81029 -3852 81085 -3796
rect 81139 -3852 81195 -3796
rect 81249 -3852 81305 -3796
rect 81359 -3852 81415 -3796
rect 80699 -3962 80755 -3906
rect 80809 -3962 80865 -3906
rect 80919 -3962 80975 -3906
rect 81029 -3962 81085 -3906
rect 81139 -3962 81195 -3906
rect 81249 -3962 81305 -3906
rect 81359 -3962 81415 -3906
rect 83552 -3408 83608 -3352
rect 83662 -3408 83718 -3352
rect 83772 -3408 83828 -3352
rect 83882 -3408 83938 -3352
rect 83992 -3408 84048 -3352
rect 84102 -3408 84158 -3352
rect 84212 -3408 84268 -3352
rect 83552 -3518 83608 -3462
rect 83662 -3518 83718 -3462
rect 83772 -3518 83828 -3462
rect 83882 -3518 83938 -3462
rect 83992 -3518 84048 -3462
rect 84102 -3518 84158 -3462
rect 84212 -3518 84268 -3462
rect 83552 -3628 83608 -3572
rect 83662 -3628 83718 -3572
rect 83772 -3628 83828 -3572
rect 83882 -3628 83938 -3572
rect 83992 -3628 84048 -3572
rect 84102 -3628 84158 -3572
rect 84212 -3628 84268 -3572
rect 83552 -3738 83608 -3682
rect 83662 -3738 83718 -3682
rect 83772 -3738 83828 -3682
rect 83882 -3738 83938 -3682
rect 83992 -3738 84048 -3682
rect 84102 -3738 84158 -3682
rect 84212 -3738 84268 -3682
rect 83552 -3848 83608 -3792
rect 83662 -3848 83718 -3792
rect 83772 -3848 83828 -3792
rect 83882 -3848 83938 -3792
rect 83992 -3848 84048 -3792
rect 84102 -3848 84158 -3792
rect 84212 -3848 84268 -3792
rect 86339 -3432 86395 -3376
rect 86449 -3432 86505 -3376
rect 86559 -3432 86615 -3376
rect 86669 -3432 86725 -3376
rect 86779 -3432 86835 -3376
rect 86889 -3432 86945 -3376
rect 86999 -3432 87055 -3376
rect 86339 -3542 86395 -3486
rect 86449 -3542 86505 -3486
rect 86559 -3542 86615 -3486
rect 86669 -3542 86725 -3486
rect 86779 -3542 86835 -3486
rect 86889 -3542 86945 -3486
rect 86999 -3542 87055 -3486
rect 86339 -3652 86395 -3596
rect 86449 -3652 86505 -3596
rect 86559 -3652 86615 -3596
rect 86669 -3652 86725 -3596
rect 86779 -3652 86835 -3596
rect 86889 -3652 86945 -3596
rect 86999 -3652 87055 -3596
rect 86339 -3762 86395 -3706
rect 86449 -3762 86505 -3706
rect 86559 -3762 86615 -3706
rect 86669 -3762 86725 -3706
rect 86779 -3762 86835 -3706
rect 86889 -3762 86945 -3706
rect 86999 -3762 87055 -3706
rect 86339 -3872 86395 -3816
rect 86449 -3872 86505 -3816
rect 86559 -3872 86615 -3816
rect 86669 -3872 86725 -3816
rect 86779 -3872 86835 -3816
rect 86889 -3872 86945 -3816
rect 86999 -3872 87055 -3816
rect 83552 -3958 83608 -3902
rect 83662 -3958 83718 -3902
rect 83772 -3958 83828 -3902
rect 83882 -3958 83938 -3902
rect 83992 -3958 84048 -3902
rect 84102 -3958 84158 -3902
rect 84212 -3958 84268 -3902
rect 86339 -3982 86395 -3926
rect 86449 -3982 86505 -3926
rect 86559 -3982 86615 -3926
rect 86669 -3982 86725 -3926
rect 86779 -3982 86835 -3926
rect 86889 -3982 86945 -3926
rect 86999 -3982 87055 -3926
rect 89521 -3385 89577 -3329
rect 89631 -3385 89687 -3329
rect 89741 -3385 89797 -3329
rect 89851 -3385 89907 -3329
rect 89961 -3385 90017 -3329
rect 90071 -3385 90127 -3329
rect 90181 -3385 90237 -3329
rect 89521 -3495 89577 -3439
rect 89631 -3495 89687 -3439
rect 89741 -3495 89797 -3439
rect 89851 -3495 89907 -3439
rect 89961 -3495 90017 -3439
rect 90071 -3495 90127 -3439
rect 90181 -3495 90237 -3439
rect 89521 -3605 89577 -3549
rect 89631 -3605 89687 -3549
rect 89741 -3605 89797 -3549
rect 89851 -3605 89907 -3549
rect 89961 -3605 90017 -3549
rect 90071 -3605 90127 -3549
rect 90181 -3605 90237 -3549
rect 89521 -3715 89577 -3659
rect 89631 -3715 89687 -3659
rect 89741 -3715 89797 -3659
rect 89851 -3715 89907 -3659
rect 89961 -3715 90017 -3659
rect 90071 -3715 90127 -3659
rect 90181 -3715 90237 -3659
rect 89521 -3825 89577 -3769
rect 89631 -3825 89687 -3769
rect 89741 -3825 89797 -3769
rect 89851 -3825 89907 -3769
rect 89961 -3825 90017 -3769
rect 90071 -3825 90127 -3769
rect 90181 -3825 90237 -3769
rect 89521 -3935 89577 -3879
rect 89631 -3935 89687 -3879
rect 89741 -3935 89797 -3879
rect 89851 -3935 89907 -3879
rect 89961 -3935 90017 -3879
rect 90071 -3935 90127 -3879
rect 90181 -3935 90237 -3879
rect 92865 -3410 92921 -3354
rect 92975 -3410 93031 -3354
rect 93085 -3410 93141 -3354
rect 93195 -3410 93251 -3354
rect 93305 -3410 93361 -3354
rect 93415 -3410 93471 -3354
rect 93525 -3410 93581 -3354
rect 92865 -3520 92921 -3464
rect 92975 -3520 93031 -3464
rect 93085 -3520 93141 -3464
rect 93195 -3520 93251 -3464
rect 93305 -3520 93361 -3464
rect 93415 -3520 93471 -3464
rect 93525 -3520 93581 -3464
rect 92865 -3630 92921 -3574
rect 92975 -3630 93031 -3574
rect 93085 -3630 93141 -3574
rect 93195 -3630 93251 -3574
rect 93305 -3630 93361 -3574
rect 93415 -3630 93471 -3574
rect 93525 -3630 93581 -3574
rect 92865 -3740 92921 -3684
rect 92975 -3740 93031 -3684
rect 93085 -3740 93141 -3684
rect 93195 -3740 93251 -3684
rect 93305 -3740 93361 -3684
rect 93415 -3740 93471 -3684
rect 93525 -3740 93581 -3684
rect 92865 -3850 92921 -3794
rect 92975 -3850 93031 -3794
rect 93085 -3850 93141 -3794
rect 93195 -3850 93251 -3794
rect 93305 -3850 93361 -3794
rect 93415 -3850 93471 -3794
rect 93525 -3850 93581 -3794
rect 95998 -3440 96054 -3384
rect 96108 -3440 96164 -3384
rect 96218 -3440 96274 -3384
rect 96328 -3440 96384 -3384
rect 96438 -3440 96494 -3384
rect 96548 -3440 96604 -3384
rect 96658 -3440 96714 -3384
rect 95998 -3550 96054 -3494
rect 96108 -3550 96164 -3494
rect 96218 -3550 96274 -3494
rect 96328 -3550 96384 -3494
rect 96438 -3550 96494 -3494
rect 96548 -3550 96604 -3494
rect 96658 -3550 96714 -3494
rect 95998 -3660 96054 -3604
rect 96108 -3660 96164 -3604
rect 96218 -3660 96274 -3604
rect 96328 -3660 96384 -3604
rect 96438 -3660 96494 -3604
rect 96548 -3660 96604 -3604
rect 96658 -3660 96714 -3604
rect 95998 -3770 96054 -3714
rect 96108 -3770 96164 -3714
rect 96218 -3770 96274 -3714
rect 96328 -3770 96384 -3714
rect 96438 -3770 96494 -3714
rect 96548 -3770 96604 -3714
rect 96658 -3770 96714 -3714
rect 92865 -3960 92921 -3904
rect 92975 -3960 93031 -3904
rect 93085 -3960 93141 -3904
rect 93195 -3960 93251 -3904
rect 93305 -3960 93361 -3904
rect 93415 -3960 93471 -3904
rect 93525 -3960 93581 -3904
rect 95998 -3880 96054 -3824
rect 96108 -3880 96164 -3824
rect 96218 -3880 96274 -3824
rect 96328 -3880 96384 -3824
rect 96438 -3880 96494 -3824
rect 96548 -3880 96604 -3824
rect 96658 -3880 96714 -3824
rect 95998 -3990 96054 -3934
rect 96108 -3990 96164 -3934
rect 96218 -3990 96274 -3934
rect 96328 -3990 96384 -3934
rect 96438 -3990 96494 -3934
rect 96548 -3990 96604 -3934
rect 96658 -3990 96714 -3934
rect 99276 -3474 99332 -3418
rect 99386 -3474 99442 -3418
rect 99496 -3474 99552 -3418
rect 99606 -3474 99662 -3418
rect 99716 -3474 99772 -3418
rect 99826 -3474 99882 -3418
rect 99936 -3474 99992 -3418
rect 99276 -3584 99332 -3528
rect 99386 -3584 99442 -3528
rect 99496 -3584 99552 -3528
rect 99606 -3584 99662 -3528
rect 99716 -3584 99772 -3528
rect 99826 -3584 99882 -3528
rect 99936 -3584 99992 -3528
rect 99276 -3694 99332 -3638
rect 99386 -3694 99442 -3638
rect 99496 -3694 99552 -3638
rect 99606 -3694 99662 -3638
rect 99716 -3694 99772 -3638
rect 99826 -3694 99882 -3638
rect 99936 -3694 99992 -3638
rect 99276 -3804 99332 -3748
rect 99386 -3804 99442 -3748
rect 99496 -3804 99552 -3748
rect 99606 -3804 99662 -3748
rect 99716 -3804 99772 -3748
rect 99826 -3804 99882 -3748
rect 99936 -3804 99992 -3748
rect 99276 -3914 99332 -3858
rect 99386 -3914 99442 -3858
rect 99496 -3914 99552 -3858
rect 99606 -3914 99662 -3858
rect 99716 -3914 99772 -3858
rect 99826 -3914 99882 -3858
rect 99936 -3914 99992 -3858
rect 99276 -4024 99332 -3968
rect 99386 -4024 99442 -3968
rect 99496 -4024 99552 -3968
rect 99606 -4024 99662 -3968
rect 99716 -4024 99772 -3968
rect 99826 -4024 99882 -3968
rect 99936 -4024 99992 -3968
rect 30166 -4207 30222 -4151
rect 30276 -4207 30332 -4151
rect 30386 -4207 30442 -4151
rect 30496 -4207 30552 -4151
rect 30606 -4207 30662 -4151
rect 30716 -4207 30772 -4151
rect 30166 -4317 30222 -4261
rect 30276 -4317 30332 -4261
rect 30386 -4317 30442 -4261
rect 30496 -4317 30552 -4261
rect 30606 -4317 30662 -4261
rect 30716 -4317 30772 -4261
rect 31209 -4668 31265 -4612
rect 31319 -4668 31375 -4612
rect 31429 -4668 31485 -4612
rect 31539 -4668 31595 -4612
rect 116662 -5276 116718 -5220
rect 116662 -5386 116718 -5330
rect 116662 -5496 116718 -5440
rect 116662 -5606 116718 -5550
rect 116662 -5716 116718 -5660
rect 116662 -5826 116718 -5770
rect 116666 -6671 116722 -6615
rect 116666 -6781 116722 -6725
rect 116666 -6891 116722 -6835
rect 116666 -7001 116722 -6945
rect 116666 -7111 116722 -7055
rect 116666 -7221 116722 -7165
rect 109078 -7951 109134 -7895
rect 109188 -7951 109244 -7895
rect 109298 -7951 109354 -7895
rect 109408 -7951 109464 -7895
rect 109518 -7951 109574 -7895
rect 109628 -7951 109684 -7895
rect 109738 -7951 109794 -7895
rect 109078 -8061 109134 -8005
rect 109188 -8061 109244 -8005
rect 109298 -8061 109354 -8005
rect 109408 -8061 109464 -8005
rect 109518 -8061 109574 -8005
rect 109628 -8061 109684 -8005
rect 109738 -8061 109794 -8005
rect 109078 -8171 109134 -8115
rect 109188 -8171 109244 -8115
rect 109298 -8171 109354 -8115
rect 109408 -8171 109464 -8115
rect 109518 -8171 109574 -8115
rect 109628 -8171 109684 -8115
rect 109738 -8171 109794 -8115
rect 109078 -8281 109134 -8225
rect 109188 -8281 109244 -8225
rect 109298 -8281 109354 -8225
rect 109408 -8281 109464 -8225
rect 109518 -8281 109574 -8225
rect 109628 -8281 109684 -8225
rect 109738 -8281 109794 -8225
rect 109078 -8391 109134 -8335
rect 109188 -8391 109244 -8335
rect 109298 -8391 109354 -8335
rect 109408 -8391 109464 -8335
rect 109518 -8391 109574 -8335
rect 109628 -8391 109684 -8335
rect 109738 -8391 109794 -8335
rect 109078 -8501 109134 -8445
rect 109188 -8501 109244 -8445
rect 109298 -8501 109354 -8445
rect 109408 -8501 109464 -8445
rect 109518 -8501 109574 -8445
rect 109628 -8501 109684 -8445
rect 109738 -8501 109794 -8445
rect 109078 -8611 109134 -8555
rect 109188 -8611 109244 -8555
rect 109298 -8611 109354 -8555
rect 109408 -8611 109464 -8555
rect 109518 -8611 109574 -8555
rect 109628 -8611 109684 -8555
rect 109738 -8611 109794 -8555
rect 109078 -8721 109134 -8665
rect 109188 -8721 109244 -8665
rect 109298 -8721 109354 -8665
rect 109408 -8721 109464 -8665
rect 109518 -8721 109574 -8665
rect 109628 -8721 109684 -8665
rect 109738 -8721 109794 -8665
rect 116664 -8502 116720 -8446
rect 116664 -8612 116720 -8556
rect 116664 -8722 116720 -8666
rect 116664 -8832 116720 -8776
rect 116664 -8942 116720 -8886
rect 116664 -9052 116720 -8996
rect 116665 -9820 116721 -9764
rect 116665 -9930 116721 -9874
rect 116665 -10040 116721 -9984
rect 116665 -10150 116721 -10094
rect 116665 -10260 116721 -10204
rect 116665 -10370 116721 -10314
rect 113550 -13263 113606 -13207
rect 113660 -13263 113716 -13207
rect 113770 -13263 113826 -13207
rect 113880 -13263 113936 -13207
rect 113990 -13263 114046 -13207
rect 114100 -13263 114156 -13207
rect 114210 -13263 114266 -13207
rect 113550 -13373 113606 -13317
rect 113660 -13373 113716 -13317
rect 113770 -13373 113826 -13317
rect 113880 -13373 113936 -13317
rect 113990 -13373 114046 -13317
rect 114100 -13373 114156 -13317
rect 114210 -13373 114266 -13317
rect 113550 -13483 113606 -13427
rect 113660 -13483 113716 -13427
rect 113770 -13483 113826 -13427
rect 113880 -13483 113936 -13427
rect 113990 -13483 114046 -13427
rect 114100 -13483 114156 -13427
rect 114210 -13483 114266 -13427
rect 29533 -13720 29589 -13664
rect 29643 -13720 29699 -13664
rect 29753 -13720 29809 -13664
rect 29863 -13720 29919 -13664
rect 29973 -13720 30029 -13664
rect 30083 -13720 30139 -13664
rect 30193 -13712 30249 -13656
rect 30303 -13712 30359 -13656
rect 30413 -13712 30469 -13656
rect 29533 -13830 29589 -13774
rect 29643 -13830 29699 -13774
rect 29753 -13830 29809 -13774
rect 29863 -13830 29919 -13774
rect 29973 -13830 30029 -13774
rect 30083 -13830 30139 -13774
rect 30193 -13822 30249 -13766
rect 30303 -13822 30359 -13766
rect 30413 -13822 30469 -13766
rect 113550 -13593 113606 -13537
rect 113660 -13593 113716 -13537
rect 113770 -13593 113826 -13537
rect 113880 -13593 113936 -13537
rect 113990 -13593 114046 -13537
rect 114100 -13593 114156 -13537
rect 114210 -13593 114266 -13537
rect 113550 -13703 113606 -13647
rect 113660 -13703 113716 -13647
rect 113770 -13703 113826 -13647
rect 113880 -13703 113936 -13647
rect 113990 -13703 114046 -13647
rect 114100 -13703 114156 -13647
rect 114210 -13703 114266 -13647
rect 113550 -13813 113606 -13757
rect 113660 -13813 113716 -13757
rect 113770 -13813 113826 -13757
rect 113880 -13813 113936 -13757
rect 113990 -13813 114046 -13757
rect 114100 -13813 114156 -13757
rect 114210 -13813 114266 -13757
rect 29852 -14525 29908 -14469
rect 29962 -14525 30018 -14469
rect 30072 -14525 30128 -14469
rect 30249 -14525 30305 -14469
rect 30359 -14525 30415 -14469
rect 30469 -14525 30525 -14469
rect 29852 -14635 29908 -14579
rect 29962 -14635 30018 -14579
rect 30072 -14635 30128 -14579
rect 30249 -14635 30305 -14579
rect 30359 -14635 30415 -14579
rect 30469 -14635 30525 -14579
rect 10245 -15108 10301 -15052
rect 10355 -15108 10411 -15052
rect 10465 -15108 10521 -15052
rect 10575 -15108 10631 -15052
rect 10685 -15108 10741 -15052
rect 10795 -15108 10851 -15052
rect 10905 -15108 10961 -15052
rect 11034 -15108 11090 -15052
rect 11144 -15108 11200 -15052
rect 11254 -15108 11310 -15052
rect 11364 -15108 11420 -15052
rect 11474 -15108 11530 -15052
rect 11584 -15108 11640 -15052
rect 11694 -15108 11750 -15052
rect 10245 -15218 10301 -15162
rect 10355 -15218 10411 -15162
rect 10465 -15218 10521 -15162
rect 10575 -15218 10631 -15162
rect 10685 -15218 10741 -15162
rect 10795 -15218 10851 -15162
rect 10905 -15218 10961 -15162
rect 11034 -15218 11090 -15162
rect 11144 -15218 11200 -15162
rect 11254 -15218 11310 -15162
rect 11364 -15218 11420 -15162
rect 11474 -15218 11530 -15162
rect 11584 -15218 11640 -15162
rect 11694 -15218 11750 -15162
rect 10245 -15328 10301 -15272
rect 10355 -15328 10411 -15272
rect 10465 -15328 10521 -15272
rect 10575 -15328 10631 -15272
rect 10685 -15328 10741 -15272
rect 10795 -15328 10851 -15272
rect 10905 -15328 10961 -15272
rect 11034 -15328 11090 -15272
rect 11144 -15328 11200 -15272
rect 11254 -15328 11310 -15272
rect 11364 -15328 11420 -15272
rect 11474 -15328 11530 -15272
rect 11584 -15328 11640 -15272
rect 11694 -15328 11750 -15272
rect 10245 -15438 10301 -15382
rect 10355 -15438 10411 -15382
rect 10465 -15438 10521 -15382
rect 10575 -15438 10631 -15382
rect 10685 -15438 10741 -15382
rect 10795 -15438 10851 -15382
rect 10905 -15438 10961 -15382
rect 11034 -15438 11090 -15382
rect 11144 -15438 11200 -15382
rect 11254 -15438 11310 -15382
rect 11364 -15438 11420 -15382
rect 11474 -15438 11530 -15382
rect 11584 -15438 11640 -15382
rect 11694 -15438 11750 -15382
rect 10245 -15548 10301 -15492
rect 10355 -15548 10411 -15492
rect 10465 -15548 10521 -15492
rect 10575 -15548 10631 -15492
rect 10685 -15548 10741 -15492
rect 10795 -15548 10851 -15492
rect 10905 -15548 10961 -15492
rect 11034 -15548 11090 -15492
rect 11144 -15548 11200 -15492
rect 11254 -15548 11310 -15492
rect 11364 -15548 11420 -15492
rect 11474 -15548 11530 -15492
rect 11584 -15548 11640 -15492
rect 11694 -15548 11750 -15492
rect 10245 -15658 10301 -15602
rect 10355 -15658 10411 -15602
rect 10465 -15658 10521 -15602
rect 10575 -15658 10631 -15602
rect 10685 -15658 10741 -15602
rect 10795 -15658 10851 -15602
rect 10905 -15658 10961 -15602
rect 11034 -15658 11090 -15602
rect 11144 -15658 11200 -15602
rect 11254 -15658 11310 -15602
rect 11364 -15658 11420 -15602
rect 11474 -15658 11530 -15602
rect 11584 -15658 11640 -15602
rect 11694 -15658 11750 -15602
rect 31310 -15674 31366 -15618
rect 31420 -15674 31476 -15618
rect 31530 -15674 31586 -15618
rect 31640 -15674 31696 -15618
rect 31310 -15784 31366 -15728
rect 31420 -15784 31476 -15728
rect 31530 -15784 31586 -15728
rect 31640 -15784 31696 -15728
rect 29779 -19858 29835 -19802
rect 29889 -19858 29945 -19802
rect 29999 -19858 30055 -19802
rect 30109 -19858 30165 -19802
rect 30333 -19865 30389 -19809
rect 30443 -19865 30499 -19809
rect 30553 -19865 30609 -19809
rect 30663 -19865 30719 -19809
rect 30887 -19856 30943 -19800
rect 30997 -19856 31053 -19800
rect 31107 -19856 31163 -19800
rect 31217 -19856 31273 -19800
rect 31427 -19872 31483 -19816
rect 31537 -19872 31593 -19816
rect 31647 -19872 31703 -19816
rect 31757 -19872 31813 -19816
rect 25916 -21478 25972 -21422
rect 26026 -21478 26082 -21422
rect 26136 -21478 26192 -21422
rect 26246 -21478 26302 -21422
rect 26356 -21478 26412 -21422
rect 26466 -21478 26522 -21422
rect 26576 -21478 26632 -21422
rect 25916 -21588 25972 -21532
rect 26026 -21588 26082 -21532
rect 26136 -21588 26192 -21532
rect 26246 -21588 26302 -21532
rect 26356 -21588 26412 -21532
rect 26466 -21588 26522 -21532
rect 26576 -21588 26632 -21532
rect 25916 -21698 25972 -21642
rect 26026 -21698 26082 -21642
rect 26136 -21698 26192 -21642
rect 26246 -21698 26302 -21642
rect 26356 -21698 26412 -21642
rect 26466 -21698 26522 -21642
rect 26576 -21698 26632 -21642
rect 24635 -23994 24691 -23938
rect 24745 -23994 24801 -23938
rect 24855 -23994 24911 -23938
rect 24965 -23994 25021 -23938
rect 25075 -23994 25131 -23938
rect 25185 -23994 25241 -23938
rect 25295 -23994 25351 -23938
rect 25405 -23994 25461 -23938
rect 24635 -24104 24691 -24048
rect 24745 -24104 24801 -24048
rect 24855 -24104 24911 -24048
rect 24965 -24104 25021 -24048
rect 25075 -24104 25131 -24048
rect 25185 -24104 25241 -24048
rect 25295 -24104 25351 -24048
rect 25405 -24104 25461 -24048
rect 24635 -24214 24691 -24158
rect 24745 -24214 24801 -24158
rect 24855 -24214 24911 -24158
rect 24965 -24214 25021 -24158
rect 25075 -24214 25131 -24158
rect 25185 -24214 25241 -24158
rect 25295 -24214 25351 -24158
rect 25405 -24214 25461 -24158
rect 24635 -24324 24691 -24268
rect 24745 -24324 24801 -24268
rect 24855 -24324 24911 -24268
rect 24965 -24324 25021 -24268
rect 25075 -24324 25131 -24268
rect 25185 -24324 25241 -24268
rect 25295 -24324 25351 -24268
rect 25405 -24324 25461 -24268
rect 24635 -24434 24691 -24378
rect 24745 -24434 24801 -24378
rect 24855 -24434 24911 -24378
rect 24965 -24434 25021 -24378
rect 25075 -24434 25131 -24378
rect 25185 -24434 25241 -24378
rect 25295 -24434 25351 -24378
rect 25405 -24434 25461 -24378
rect 24635 -24544 24691 -24488
rect 24745 -24544 24801 -24488
rect 24855 -24544 24911 -24488
rect 24965 -24544 25021 -24488
rect 25075 -24544 25131 -24488
rect 25185 -24544 25241 -24488
rect 25295 -24544 25351 -24488
rect 25405 -24544 25461 -24488
rect 39307 -29003 39363 -28947
rect 39417 -29003 39473 -28947
rect 39527 -29003 39583 -28947
rect 39637 -29003 39693 -28947
rect 39747 -29003 39803 -28947
rect 39857 -29003 39913 -28947
rect 39967 -29003 40023 -28947
rect 39307 -29113 39363 -29057
rect 39417 -29113 39473 -29057
rect 39527 -29113 39583 -29057
rect 39637 -29113 39693 -29057
rect 39747 -29113 39803 -29057
rect 39857 -29113 39913 -29057
rect 39967 -29113 40023 -29057
rect 39307 -29223 39363 -29167
rect 39417 -29223 39473 -29167
rect 39527 -29223 39583 -29167
rect 39637 -29223 39693 -29167
rect 39747 -29223 39803 -29167
rect 39857 -29223 39913 -29167
rect 39967 -29223 40023 -29167
rect 39307 -29333 39363 -29277
rect 39417 -29333 39473 -29277
rect 39527 -29333 39583 -29277
rect 39637 -29333 39693 -29277
rect 39747 -29333 39803 -29277
rect 39857 -29333 39913 -29277
rect 39967 -29333 40023 -29277
rect 39307 -29443 39363 -29387
rect 39417 -29443 39473 -29387
rect 39527 -29443 39583 -29387
rect 39637 -29443 39693 -29387
rect 39747 -29443 39803 -29387
rect 39857 -29443 39913 -29387
rect 39967 -29443 40023 -29387
rect 39307 -29553 39363 -29497
rect 39417 -29553 39473 -29497
rect 39527 -29553 39583 -29497
rect 39637 -29553 39693 -29497
rect 39747 -29553 39803 -29497
rect 39857 -29553 39913 -29497
rect 39967 -29553 40023 -29497
rect 10249 -29751 10305 -29695
rect 10359 -29751 10415 -29695
rect 10469 -29751 10525 -29695
rect 10579 -29751 10635 -29695
rect 10689 -29751 10745 -29695
rect 10799 -29751 10855 -29695
rect 10909 -29751 10965 -29695
rect 11038 -29751 11094 -29695
rect 11148 -29751 11204 -29695
rect 11258 -29751 11314 -29695
rect 11368 -29751 11424 -29695
rect 11478 -29751 11534 -29695
rect 11588 -29751 11644 -29695
rect 11698 -29751 11754 -29695
rect 10249 -29861 10305 -29805
rect 10359 -29861 10415 -29805
rect 10469 -29861 10525 -29805
rect 10579 -29861 10635 -29805
rect 10689 -29861 10745 -29805
rect 10799 -29861 10855 -29805
rect 10909 -29861 10965 -29805
rect 11038 -29861 11094 -29805
rect 11148 -29861 11204 -29805
rect 11258 -29861 11314 -29805
rect 11368 -29861 11424 -29805
rect 11478 -29861 11534 -29805
rect 11588 -29861 11644 -29805
rect 11698 -29861 11754 -29805
rect 39307 -29663 39363 -29607
rect 39417 -29663 39473 -29607
rect 39527 -29663 39583 -29607
rect 39637 -29663 39693 -29607
rect 39747 -29663 39803 -29607
rect 39857 -29663 39913 -29607
rect 39967 -29663 40023 -29607
rect 39307 -29773 39363 -29717
rect 39417 -29773 39473 -29717
rect 39527 -29773 39583 -29717
rect 39637 -29773 39693 -29717
rect 39747 -29773 39803 -29717
rect 39857 -29773 39913 -29717
rect 39967 -29773 40023 -29717
rect 10249 -29971 10305 -29915
rect 10359 -29971 10415 -29915
rect 10469 -29971 10525 -29915
rect 10579 -29971 10635 -29915
rect 10689 -29971 10745 -29915
rect 10799 -29971 10855 -29915
rect 10909 -29971 10965 -29915
rect 11038 -29971 11094 -29915
rect 11148 -29971 11204 -29915
rect 11258 -29971 11314 -29915
rect 11368 -29971 11424 -29915
rect 11478 -29971 11534 -29915
rect 11588 -29971 11644 -29915
rect 11698 -29971 11754 -29915
rect 10249 -30081 10305 -30025
rect 10359 -30081 10415 -30025
rect 10469 -30081 10525 -30025
rect 10579 -30081 10635 -30025
rect 10689 -30081 10745 -30025
rect 10799 -30081 10855 -30025
rect 10909 -30081 10965 -30025
rect 11038 -30081 11094 -30025
rect 11148 -30081 11204 -30025
rect 11258 -30081 11314 -30025
rect 11368 -30081 11424 -30025
rect 11478 -30081 11534 -30025
rect 11588 -30081 11644 -30025
rect 11698 -30081 11754 -30025
rect 56591 -27874 56647 -27818
rect 56701 -27874 56757 -27818
rect 56811 -27874 56867 -27818
rect 56921 -27874 56977 -27818
rect 57031 -27874 57087 -27818
rect 57141 -27874 57197 -27818
rect 57251 -27874 57307 -27818
rect 56591 -27984 56647 -27928
rect 56701 -27984 56757 -27928
rect 56811 -27984 56867 -27928
rect 56921 -27984 56977 -27928
rect 57031 -27984 57087 -27928
rect 57141 -27984 57197 -27928
rect 57251 -27984 57307 -27928
rect 56591 -28094 56647 -28038
rect 56701 -28094 56757 -28038
rect 56811 -28094 56867 -28038
rect 56921 -28094 56977 -28038
rect 57031 -28094 57087 -28038
rect 57141 -28094 57197 -28038
rect 57251 -28094 57307 -28038
rect 56591 -28204 56647 -28148
rect 56701 -28204 56757 -28148
rect 56811 -28204 56867 -28148
rect 56921 -28204 56977 -28148
rect 57031 -28204 57087 -28148
rect 57141 -28204 57197 -28148
rect 57251 -28204 57307 -28148
rect 56591 -28314 56647 -28258
rect 56701 -28314 56757 -28258
rect 56811 -28314 56867 -28258
rect 56921 -28314 56977 -28258
rect 57031 -28314 57087 -28258
rect 57141 -28314 57197 -28258
rect 57251 -28314 57307 -28258
rect 56591 -28424 56647 -28368
rect 56701 -28424 56757 -28368
rect 56811 -28424 56867 -28368
rect 56921 -28424 56977 -28368
rect 57031 -28424 57087 -28368
rect 57141 -28424 57197 -28368
rect 57251 -28424 57307 -28368
rect 56591 -28534 56647 -28478
rect 56701 -28534 56757 -28478
rect 56811 -28534 56867 -28478
rect 56921 -28534 56977 -28478
rect 57031 -28534 57087 -28478
rect 57141 -28534 57197 -28478
rect 57251 -28534 57307 -28478
rect 56591 -28644 56647 -28588
rect 56701 -28644 56757 -28588
rect 56811 -28644 56867 -28588
rect 56921 -28644 56977 -28588
rect 57031 -28644 57087 -28588
rect 57141 -28644 57197 -28588
rect 57251 -28644 57307 -28588
rect 24746 -30553 24802 -30497
rect 24856 -30553 24912 -30497
rect 24966 -30553 25022 -30497
rect 25076 -30553 25132 -30497
rect 25186 -30553 25242 -30497
rect 25296 -30553 25352 -30497
rect 25406 -30553 25462 -30497
rect 113577 -30504 113633 -30448
rect 113687 -30504 113743 -30448
rect 113797 -30504 113853 -30448
rect 113907 -30504 113963 -30448
rect 114017 -30504 114073 -30448
rect 114127 -30504 114183 -30448
rect 114237 -30504 114293 -30448
rect 24746 -30663 24802 -30607
rect 24856 -30663 24912 -30607
rect 24966 -30663 25022 -30607
rect 25076 -30663 25132 -30607
rect 25186 -30663 25242 -30607
rect 25296 -30663 25352 -30607
rect 25406 -30663 25462 -30607
rect 113577 -30614 113633 -30558
rect 113687 -30614 113743 -30558
rect 113797 -30614 113853 -30558
rect 113907 -30614 113963 -30558
rect 114017 -30614 114073 -30558
rect 114127 -30614 114183 -30558
rect 114237 -30614 114293 -30558
rect 24746 -30773 24802 -30717
rect 24856 -30773 24912 -30717
rect 24966 -30773 25022 -30717
rect 25076 -30773 25132 -30717
rect 25186 -30773 25242 -30717
rect 25296 -30773 25352 -30717
rect 25406 -30773 25462 -30717
rect 113577 -30724 113633 -30668
rect 113687 -30724 113743 -30668
rect 113797 -30724 113853 -30668
rect 113907 -30724 113963 -30668
rect 114017 -30724 114073 -30668
rect 114127 -30724 114183 -30668
rect 114237 -30724 114293 -30668
rect 24746 -30883 24802 -30827
rect 24856 -30883 24912 -30827
rect 24966 -30883 25022 -30827
rect 25076 -30883 25132 -30827
rect 25186 -30883 25242 -30827
rect 25296 -30883 25352 -30827
rect 25406 -30883 25462 -30827
rect 113577 -30834 113633 -30778
rect 113687 -30834 113743 -30778
rect 113797 -30834 113853 -30778
rect 113907 -30834 113963 -30778
rect 114017 -30834 114073 -30778
rect 114127 -30834 114183 -30778
rect 114237 -30834 114293 -30778
rect 24746 -30993 24802 -30937
rect 24856 -30993 24912 -30937
rect 24966 -30993 25022 -30937
rect 25076 -30993 25132 -30937
rect 25186 -30993 25242 -30937
rect 25296 -30993 25352 -30937
rect 25406 -30993 25462 -30937
rect 113577 -30944 113633 -30888
rect 113687 -30944 113743 -30888
rect 113797 -30944 113853 -30888
rect 113907 -30944 113963 -30888
rect 114017 -30944 114073 -30888
rect 114127 -30944 114183 -30888
rect 114237 -30944 114293 -30888
rect 24746 -31103 24802 -31047
rect 24856 -31103 24912 -31047
rect 24966 -31103 25022 -31047
rect 25076 -31103 25132 -31047
rect 25186 -31103 25242 -31047
rect 25296 -31103 25352 -31047
rect 25406 -31103 25462 -31047
rect 113577 -31054 113633 -30998
rect 113687 -31054 113743 -30998
rect 113797 -31054 113853 -30998
rect 113907 -31054 113963 -30998
rect 114017 -31054 114073 -30998
rect 114127 -31054 114183 -30998
rect 114237 -31054 114293 -30998
rect 25910 -31670 25966 -31614
rect 26020 -31670 26076 -31614
rect 26130 -31670 26186 -31614
rect 26240 -31670 26296 -31614
rect 26350 -31670 26406 -31614
rect 26460 -31670 26516 -31614
rect 26570 -31670 26626 -31614
rect 10247 -31728 10303 -31672
rect 10357 -31728 10413 -31672
rect 10467 -31728 10523 -31672
rect 10577 -31728 10633 -31672
rect 10687 -31728 10743 -31672
rect 10797 -31728 10853 -31672
rect 10907 -31728 10963 -31672
rect 11036 -31728 11092 -31672
rect 11146 -31728 11202 -31672
rect 11256 -31728 11312 -31672
rect 11366 -31728 11422 -31672
rect 11476 -31728 11532 -31672
rect 11586 -31728 11642 -31672
rect 11696 -31728 11752 -31672
rect 114633 -31715 114689 -31659
rect 114743 -31715 114799 -31659
rect 114853 -31715 114909 -31659
rect 114963 -31715 115019 -31659
rect 115073 -31715 115129 -31659
rect 115183 -31715 115239 -31659
rect 115293 -31715 115349 -31659
rect 25910 -31780 25966 -31724
rect 26020 -31780 26076 -31724
rect 26130 -31780 26186 -31724
rect 26240 -31780 26296 -31724
rect 26350 -31780 26406 -31724
rect 26460 -31780 26516 -31724
rect 26570 -31780 26626 -31724
rect 10247 -31838 10303 -31782
rect 10357 -31838 10413 -31782
rect 10467 -31838 10523 -31782
rect 10577 -31838 10633 -31782
rect 10687 -31838 10743 -31782
rect 10797 -31838 10853 -31782
rect 10907 -31838 10963 -31782
rect 11036 -31838 11092 -31782
rect 11146 -31838 11202 -31782
rect 11256 -31838 11312 -31782
rect 11366 -31838 11422 -31782
rect 11476 -31838 11532 -31782
rect 11586 -31838 11642 -31782
rect 11696 -31838 11752 -31782
rect 114633 -31825 114689 -31769
rect 114743 -31825 114799 -31769
rect 114853 -31825 114909 -31769
rect 114963 -31825 115019 -31769
rect 115073 -31825 115129 -31769
rect 115183 -31825 115239 -31769
rect 115293 -31825 115349 -31769
rect 25910 -31890 25966 -31834
rect 26020 -31890 26076 -31834
rect 26130 -31890 26186 -31834
rect 26240 -31890 26296 -31834
rect 26350 -31890 26406 -31834
rect 26460 -31890 26516 -31834
rect 26570 -31890 26626 -31834
rect 10247 -31948 10303 -31892
rect 10357 -31948 10413 -31892
rect 10467 -31948 10523 -31892
rect 10577 -31948 10633 -31892
rect 10687 -31948 10743 -31892
rect 10797 -31948 10853 -31892
rect 10907 -31948 10963 -31892
rect 11036 -31948 11092 -31892
rect 11146 -31948 11202 -31892
rect 11256 -31948 11312 -31892
rect 11366 -31948 11422 -31892
rect 11476 -31948 11532 -31892
rect 11586 -31948 11642 -31892
rect 11696 -31948 11752 -31892
rect 114633 -31935 114689 -31879
rect 114743 -31935 114799 -31879
rect 114853 -31935 114909 -31879
rect 114963 -31935 115019 -31879
rect 115073 -31935 115129 -31879
rect 115183 -31935 115239 -31879
rect 115293 -31935 115349 -31879
rect 25910 -32000 25966 -31944
rect 26020 -32000 26076 -31944
rect 26130 -32000 26186 -31944
rect 26240 -32000 26296 -31944
rect 26350 -32000 26406 -31944
rect 26460 -32000 26516 -31944
rect 26570 -32000 26626 -31944
rect 10247 -32058 10303 -32002
rect 10357 -32058 10413 -32002
rect 10467 -32058 10523 -32002
rect 10577 -32058 10633 -32002
rect 10687 -32058 10743 -32002
rect 10797 -32058 10853 -32002
rect 10907 -32058 10963 -32002
rect 11036 -32058 11092 -32002
rect 11146 -32058 11202 -32002
rect 11256 -32058 11312 -32002
rect 11366 -32058 11422 -32002
rect 11476 -32058 11532 -32002
rect 11586 -32058 11642 -32002
rect 11696 -32058 11752 -32002
rect 114633 -32045 114689 -31989
rect 114743 -32045 114799 -31989
rect 114853 -32045 114909 -31989
rect 114963 -32045 115019 -31989
rect 115073 -32045 115129 -31989
rect 115183 -32045 115239 -31989
rect 115293 -32045 115349 -31989
rect 25910 -32110 25966 -32054
rect 26020 -32110 26076 -32054
rect 26130 -32110 26186 -32054
rect 26240 -32110 26296 -32054
rect 26350 -32110 26406 -32054
rect 26460 -32110 26516 -32054
rect 26570 -32110 26626 -32054
rect 10247 -32168 10303 -32112
rect 10357 -32168 10413 -32112
rect 10467 -32168 10523 -32112
rect 10577 -32168 10633 -32112
rect 10687 -32168 10743 -32112
rect 10797 -32168 10853 -32112
rect 10907 -32168 10963 -32112
rect 11036 -32168 11092 -32112
rect 11146 -32168 11202 -32112
rect 11256 -32168 11312 -32112
rect 11366 -32168 11422 -32112
rect 11476 -32168 11532 -32112
rect 11586 -32168 11642 -32112
rect 11696 -32168 11752 -32112
rect 114633 -32155 114689 -32099
rect 114743 -32155 114799 -32099
rect 114853 -32155 114909 -32099
rect 114963 -32155 115019 -32099
rect 115073 -32155 115129 -32099
rect 115183 -32155 115239 -32099
rect 115293 -32155 115349 -32099
rect 25910 -32220 25966 -32164
rect 26020 -32220 26076 -32164
rect 26130 -32220 26186 -32164
rect 26240 -32220 26296 -32164
rect 26350 -32220 26406 -32164
rect 26460 -32220 26516 -32164
rect 26570 -32220 26626 -32164
rect 10247 -32278 10303 -32222
rect 10357 -32278 10413 -32222
rect 10467 -32278 10523 -32222
rect 10577 -32278 10633 -32222
rect 10687 -32278 10743 -32222
rect 10797 -32278 10853 -32222
rect 10907 -32278 10963 -32222
rect 11036 -32278 11092 -32222
rect 11146 -32278 11202 -32222
rect 11256 -32278 11312 -32222
rect 11366 -32278 11422 -32222
rect 11476 -32278 11532 -32222
rect 11586 -32278 11642 -32222
rect 11696 -32278 11752 -32222
rect 114633 -32265 114689 -32209
rect 114743 -32265 114799 -32209
rect 114853 -32265 114909 -32209
rect 114963 -32265 115019 -32209
rect 115073 -32265 115129 -32209
rect 115183 -32265 115239 -32209
rect 115293 -32265 115349 -32209
<< metal2 >>
rect 24632 19845 25532 19894
rect 24632 19789 24715 19845
rect 24771 19789 24825 19845
rect 24881 19789 24935 19845
rect 24991 19789 25045 19845
rect 25101 19789 25155 19845
rect 25211 19789 25265 19845
rect 25321 19789 25375 19845
rect 25431 19789 25532 19845
rect 24632 19735 25532 19789
rect 24632 19679 24715 19735
rect 24771 19679 24825 19735
rect 24881 19679 24935 19735
rect 24991 19679 25045 19735
rect 25101 19679 25155 19735
rect 25211 19679 25265 19735
rect 25321 19679 25375 19735
rect 25431 19679 25532 19735
rect 24632 19625 25532 19679
rect 24632 19569 24715 19625
rect 24771 19569 24825 19625
rect 24881 19569 24935 19625
rect 24991 19569 25045 19625
rect 25101 19569 25155 19625
rect 25211 19569 25265 19625
rect 25321 19569 25375 19625
rect 25431 19569 25532 19625
rect 24632 19515 25532 19569
rect 24632 19459 24715 19515
rect 24771 19459 24825 19515
rect 24881 19459 24935 19515
rect 24991 19459 25045 19515
rect 25101 19459 25155 19515
rect 25211 19459 25265 19515
rect 25321 19459 25375 19515
rect 25431 19459 25532 19515
rect 24632 19405 25532 19459
rect 24632 19349 24715 19405
rect 24771 19349 24825 19405
rect 24881 19349 24935 19405
rect 24991 19349 25045 19405
rect 25101 19349 25155 19405
rect 25211 19349 25265 19405
rect 25321 19349 25375 19405
rect 25431 19349 25532 19405
rect 24632 19295 25532 19349
rect 24632 19239 24715 19295
rect 24771 19239 24825 19295
rect 24881 19239 24935 19295
rect 24991 19239 25045 19295
rect 25101 19239 25155 19295
rect 25211 19239 25265 19295
rect 25321 19239 25375 19295
rect 25431 19239 25532 19295
rect 1185 15616 6043 16549
rect -836 2983 -82 3015
rect -836 2948 -67 2983
rect -836 2892 -808 2948
rect -752 2892 -698 2948
rect -642 2892 -588 2948
rect -532 2892 -478 2948
rect -422 2892 -368 2948
rect -312 2892 -258 2948
rect -202 2892 -148 2948
rect -92 2892 -67 2948
rect -836 2838 -67 2892
rect -836 2782 -808 2838
rect -752 2782 -698 2838
rect -642 2782 -588 2838
rect -532 2782 -478 2838
rect -422 2782 -368 2838
rect -312 2782 -258 2838
rect -202 2782 -148 2838
rect -92 2782 -67 2838
rect -836 2728 -67 2782
rect -836 2672 -808 2728
rect -752 2672 -698 2728
rect -642 2672 -588 2728
rect -532 2672 -478 2728
rect -422 2672 -368 2728
rect -312 2672 -258 2728
rect -202 2672 -148 2728
rect -92 2672 -67 2728
rect -836 2618 -67 2672
rect -836 2562 -808 2618
rect -752 2562 -698 2618
rect -642 2562 -588 2618
rect -532 2562 -478 2618
rect -422 2562 -368 2618
rect -312 2562 -258 2618
rect -202 2562 -148 2618
rect -92 2562 -67 2618
rect -836 2508 -67 2562
rect -836 2452 -808 2508
rect -752 2452 -698 2508
rect -642 2452 -588 2508
rect -532 2452 -478 2508
rect -422 2452 -368 2508
rect -312 2452 -258 2508
rect -202 2452 -148 2508
rect -92 2452 -67 2508
rect -836 2398 -67 2452
rect -836 2342 -808 2398
rect -752 2342 -698 2398
rect -642 2342 -588 2398
rect -532 2342 -478 2398
rect -422 2342 -368 2398
rect -312 2342 -258 2398
rect -202 2342 -148 2398
rect -92 2342 -67 2398
rect -836 2298 -67 2342
rect -836 -16384 -82 2298
rect 97 -2146 851 -2049
rect 97 -2181 879 -2146
rect 97 -2237 138 -2181
rect 194 -2237 248 -2181
rect 304 -2237 358 -2181
rect 414 -2237 468 -2181
rect 524 -2237 578 -2181
rect 634 -2237 688 -2181
rect 744 -2237 798 -2181
rect 854 -2237 879 -2181
rect 97 -2291 879 -2237
rect 97 -2347 138 -2291
rect 194 -2347 248 -2291
rect 304 -2347 358 -2291
rect 414 -2347 468 -2291
rect 524 -2347 578 -2291
rect 634 -2347 688 -2291
rect 744 -2347 798 -2291
rect 854 -2347 879 -2291
rect 97 -2401 879 -2347
rect 97 -2457 138 -2401
rect 194 -2457 248 -2401
rect 304 -2457 358 -2401
rect 414 -2457 468 -2401
rect 524 -2457 578 -2401
rect 634 -2457 688 -2401
rect 744 -2457 798 -2401
rect 854 -2457 879 -2401
rect 97 -2511 879 -2457
rect 97 -2567 138 -2511
rect 194 -2567 248 -2511
rect 304 -2567 358 -2511
rect 414 -2567 468 -2511
rect 524 -2567 578 -2511
rect 634 -2567 688 -2511
rect 744 -2567 798 -2511
rect 854 -2567 879 -2511
rect 97 -2621 879 -2567
rect 97 -2677 138 -2621
rect 194 -2677 248 -2621
rect 304 -2677 358 -2621
rect 414 -2677 468 -2621
rect 524 -2677 578 -2621
rect 634 -2677 688 -2621
rect 744 -2677 798 -2621
rect 854 -2677 879 -2621
rect 97 -2731 879 -2677
rect 97 -2787 138 -2731
rect 194 -2787 248 -2731
rect 304 -2787 358 -2731
rect 414 -2787 468 -2731
rect 524 -2787 578 -2731
rect 634 -2787 688 -2731
rect 744 -2787 798 -2731
rect 854 -2787 879 -2731
rect 97 -2831 879 -2787
rect -836 -16413 -78 -16384
rect -836 -16469 -814 -16413
rect -758 -16469 -704 -16413
rect -648 -16469 -594 -16413
rect -538 -16469 -484 -16413
rect -428 -16469 -374 -16413
rect -318 -16469 -264 -16413
rect -208 -16469 -154 -16413
rect -98 -16469 -78 -16413
rect -836 -16523 -78 -16469
rect -836 -16579 -814 -16523
rect -758 -16579 -704 -16523
rect -648 -16579 -594 -16523
rect -538 -16579 -484 -16523
rect -428 -16579 -374 -16523
rect -318 -16579 -264 -16523
rect -208 -16579 -154 -16523
rect -98 -16579 -78 -16523
rect -836 -16633 -78 -16579
rect -836 -16689 -814 -16633
rect -758 -16689 -704 -16633
rect -648 -16689 -594 -16633
rect -538 -16689 -484 -16633
rect -428 -16689 -374 -16633
rect -318 -16689 -264 -16633
rect -208 -16689 -154 -16633
rect -98 -16689 -78 -16633
rect -836 -16743 -78 -16689
rect -836 -16799 -814 -16743
rect -758 -16799 -704 -16743
rect -648 -16799 -594 -16743
rect -538 -16799 -484 -16743
rect -428 -16799 -374 -16743
rect -318 -16799 -264 -16743
rect -208 -16799 -154 -16743
rect -98 -16799 -78 -16743
rect -836 -16853 -78 -16799
rect -836 -16909 -814 -16853
rect -758 -16909 -704 -16853
rect -648 -16909 -594 -16853
rect -538 -16909 -484 -16853
rect -428 -16909 -374 -16853
rect -318 -16909 -264 -16853
rect -208 -16909 -154 -16853
rect -98 -16909 -78 -16853
rect -836 -16963 -78 -16909
rect -836 -17019 -814 -16963
rect -758 -17019 -704 -16963
rect -648 -17019 -594 -16963
rect -538 -17019 -484 -16963
rect -428 -17019 -374 -16963
rect -318 -17019 -264 -16963
rect -208 -17019 -154 -16963
rect -98 -17019 -78 -16963
rect -836 -17073 -78 -17019
rect -836 -17129 -814 -17073
rect -758 -17129 -704 -17073
rect -648 -17129 -594 -17073
rect -538 -17129 -484 -17073
rect -428 -17129 -374 -17073
rect -318 -17129 -264 -17073
rect -208 -17129 -154 -17073
rect -98 -17129 -78 -17073
rect -836 -17143 -78 -17129
rect -836 -17324 -82 -17143
rect 97 -17316 851 -2831
rect 97 -17327 861 -17316
rect 106 -17348 861 -17327
rect 106 -17404 121 -17348
rect 177 -17404 231 -17348
rect 287 -17404 341 -17348
rect 397 -17404 451 -17348
rect 507 -17404 561 -17348
rect 617 -17404 671 -17348
rect 727 -17404 781 -17348
rect 837 -17404 861 -17348
rect 106 -17458 861 -17404
rect 106 -17514 121 -17458
rect 177 -17514 231 -17458
rect 287 -17514 341 -17458
rect 397 -17514 451 -17458
rect 507 -17514 561 -17458
rect 617 -17514 671 -17458
rect 727 -17514 781 -17458
rect 837 -17514 861 -17458
rect 106 -17568 861 -17514
rect 106 -17624 121 -17568
rect 177 -17624 231 -17568
rect 287 -17624 341 -17568
rect 397 -17624 451 -17568
rect 507 -17624 561 -17568
rect 617 -17624 671 -17568
rect 727 -17624 781 -17568
rect 837 -17624 861 -17568
rect 106 -17678 861 -17624
rect 106 -17734 121 -17678
rect 177 -17734 231 -17678
rect 287 -17734 341 -17678
rect 397 -17734 451 -17678
rect 507 -17734 561 -17678
rect 617 -17734 671 -17678
rect 727 -17734 781 -17678
rect 837 -17734 861 -17678
rect 106 -17788 861 -17734
rect 106 -17844 121 -17788
rect 177 -17844 231 -17788
rect 287 -17844 341 -17788
rect 397 -17844 451 -17788
rect 507 -17844 561 -17788
rect 617 -17844 671 -17788
rect 727 -17844 781 -17788
rect 837 -17844 861 -17788
rect 106 -17898 861 -17844
rect 106 -17954 121 -17898
rect 177 -17954 231 -17898
rect 287 -17954 341 -17898
rect 397 -17954 451 -17898
rect 507 -17954 561 -17898
rect 617 -17954 671 -17898
rect 727 -17954 781 -17898
rect 837 -17954 861 -17898
rect 106 -18008 861 -17954
rect 106 -18064 121 -18008
rect 177 -18064 231 -18008
rect 287 -18064 341 -18008
rect 397 -18064 451 -18008
rect 507 -18064 561 -18008
rect 617 -18064 671 -18008
rect 727 -18064 781 -18008
rect 837 -18064 861 -18008
rect 106 -18076 861 -18064
rect 106 -18082 851 -18076
rect 1185 -18281 2118 15616
rect 4860 15377 6040 15616
rect 10753 3485 12429 3491
rect 10737 3443 12429 3485
rect 10737 3387 10800 3443
rect 10856 3387 10910 3443
rect 10966 3387 11020 3443
rect 11076 3387 11130 3443
rect 11186 3387 11240 3443
rect 11296 3387 11350 3443
rect 11406 3387 11460 3443
rect 11516 3387 11624 3443
rect 11680 3387 11734 3443
rect 11790 3387 11844 3443
rect 11900 3387 11954 3443
rect 12010 3387 12064 3443
rect 12120 3387 12174 3443
rect 12230 3387 12284 3443
rect 12340 3387 12429 3443
rect 10737 3333 12429 3387
rect 10737 3277 10800 3333
rect 10856 3277 10910 3333
rect 10966 3277 11020 3333
rect 11076 3277 11130 3333
rect 11186 3277 11240 3333
rect 11296 3277 11350 3333
rect 11406 3277 11460 3333
rect 11516 3277 11624 3333
rect 11680 3277 11734 3333
rect 11790 3277 11844 3333
rect 11900 3277 11954 3333
rect 12010 3277 12064 3333
rect 12120 3277 12174 3333
rect 12230 3277 12284 3333
rect 12340 3277 12429 3333
rect 10737 3223 12429 3277
rect 10737 3167 10800 3223
rect 10856 3167 10910 3223
rect 10966 3167 11020 3223
rect 11076 3167 11130 3223
rect 11186 3167 11240 3223
rect 11296 3167 11350 3223
rect 11406 3167 11460 3223
rect 11516 3167 11624 3223
rect 11680 3167 11734 3223
rect 11790 3167 11844 3223
rect 11900 3167 11954 3223
rect 12010 3167 12064 3223
rect 12120 3167 12174 3223
rect 12230 3167 12284 3223
rect 12340 3167 12429 3223
rect 10737 3113 12429 3167
rect 10737 3057 10800 3113
rect 10856 3057 10910 3113
rect 10966 3057 11020 3113
rect 11076 3057 11130 3113
rect 11186 3057 11240 3113
rect 11296 3057 11350 3113
rect 11406 3057 11460 3113
rect 11516 3057 11624 3113
rect 11680 3057 11734 3113
rect 11790 3057 11844 3113
rect 11900 3057 11954 3113
rect 12010 3057 12064 3113
rect 12120 3057 12174 3113
rect 12230 3057 12284 3113
rect 12340 3057 12429 3113
rect 10737 3003 12429 3057
rect 10737 2947 10800 3003
rect 10856 2947 10910 3003
rect 10966 2947 11020 3003
rect 11076 2947 11130 3003
rect 11186 2947 11240 3003
rect 11296 2947 11350 3003
rect 11406 2947 11460 3003
rect 11516 2947 11624 3003
rect 11680 2947 11734 3003
rect 11790 2947 11844 3003
rect 11900 2947 11954 3003
rect 12010 2947 12064 3003
rect 12120 2947 12174 3003
rect 12230 2947 12284 3003
rect 12340 2947 12429 3003
rect 10737 2893 12429 2947
rect 10737 2837 10800 2893
rect 10856 2837 10910 2893
rect 10966 2837 11020 2893
rect 11076 2837 11130 2893
rect 11186 2837 11240 2893
rect 11296 2837 11350 2893
rect 11406 2837 11460 2893
rect 11516 2837 11624 2893
rect 11680 2837 11734 2893
rect 11790 2837 11844 2893
rect 11900 2837 11954 2893
rect 12010 2837 12064 2893
rect 12120 2837 12174 2893
rect 12230 2837 12284 2893
rect 12340 2837 12429 2893
rect 10737 2795 12429 2837
rect 3089 2637 3518 2653
rect 3089 2581 3111 2637
rect 3167 2581 3221 2637
rect 3277 2581 3331 2637
rect 3387 2581 3441 2637
rect 3497 2581 3518 2637
rect 3089 2527 3518 2581
rect 3089 2471 3111 2527
rect 3167 2471 3221 2527
rect 3277 2471 3331 2527
rect 3387 2471 3441 2527
rect 3497 2471 3518 2527
rect 3089 2417 3518 2471
rect 3089 2361 3111 2417
rect 3167 2361 3221 2417
rect 3277 2361 3331 2417
rect 3387 2361 3441 2417
rect 3497 2361 3518 2417
rect 3089 2307 3518 2361
rect 3089 2251 3111 2307
rect 3167 2251 3221 2307
rect 3277 2251 3331 2307
rect 3387 2251 3441 2307
rect 3497 2251 3518 2307
rect 3089 2226 3518 2251
rect 3089 37 3316 2226
rect 6286 1186 7074 1217
rect 6286 1130 6315 1186
rect 6371 1130 6425 1186
rect 6481 1130 6535 1186
rect 6591 1130 6645 1186
rect 6701 1130 6755 1186
rect 6811 1130 6865 1186
rect 6921 1130 6975 1186
rect 7031 1130 7074 1186
rect 6286 1076 7074 1130
rect 6286 1020 6315 1076
rect 6371 1020 6425 1076
rect 6481 1020 6535 1076
rect 6591 1020 6645 1076
rect 6701 1020 6755 1076
rect 6811 1020 6865 1076
rect 6921 1020 6975 1076
rect 7031 1020 7074 1076
rect 6286 966 7074 1020
rect 6286 910 6315 966
rect 6371 910 6425 966
rect 6481 910 6535 966
rect 6591 910 6645 966
rect 6701 910 6755 966
rect 6811 910 6865 966
rect 6921 910 6975 966
rect 7031 910 7074 966
rect 6286 856 7074 910
rect 6286 800 6315 856
rect 6371 800 6425 856
rect 6481 800 6535 856
rect 6591 800 6645 856
rect 6701 800 6755 856
rect 6811 800 6865 856
rect 6921 800 6975 856
rect 7031 800 7074 856
rect 6286 746 7074 800
rect 6286 690 6315 746
rect 6371 690 6425 746
rect 6481 690 6535 746
rect 6591 690 6645 746
rect 6701 690 6755 746
rect 6811 690 6865 746
rect 6921 690 6975 746
rect 7031 690 7074 746
rect 6286 636 7074 690
rect 6286 580 6315 636
rect 6371 580 6425 636
rect 6481 580 6535 636
rect 6591 580 6645 636
rect 6701 580 6755 636
rect 6811 580 6865 636
rect 6921 580 6975 636
rect 7031 580 7074 636
rect 6286 560 7074 580
rect 4298 -658 4354 -648
rect 4298 -724 4354 -714
rect 4298 -768 4354 -758
rect 4298 -834 4354 -824
rect 5628 -1568 5855 525
rect 5522 -1584 5951 -1568
rect 5522 -1640 5544 -1584
rect 5600 -1640 5654 -1584
rect 5710 -1640 5764 -1584
rect 5820 -1640 5874 -1584
rect 5930 -1640 5951 -1584
rect 5522 -1694 5951 -1640
rect 5522 -1750 5544 -1694
rect 5600 -1750 5654 -1694
rect 5710 -1750 5764 -1694
rect 5820 -1750 5874 -1694
rect 5930 -1750 5951 -1694
rect 5522 -1804 5951 -1750
rect 5522 -1860 5544 -1804
rect 5600 -1860 5654 -1804
rect 5710 -1860 5764 -1804
rect 5820 -1860 5874 -1804
rect 5930 -1860 5951 -1804
rect 5522 -1914 5951 -1860
rect 5522 -1970 5544 -1914
rect 5600 -1970 5654 -1914
rect 5710 -1970 5764 -1914
rect 5820 -1970 5874 -1914
rect 5930 -1970 5951 -1914
rect 5522 -1995 5951 -1970
rect 6287 -2554 7055 560
rect 10753 -1128 12429 2795
rect 22871 1204 23661 1220
rect 10753 -1184 10881 -1128
rect 10937 -1184 10991 -1128
rect 11047 -1184 11101 -1128
rect 11157 -1184 11211 -1128
rect 11267 -1184 11321 -1128
rect 11377 -1184 11431 -1128
rect 11487 -1184 11541 -1128
rect 11597 -1184 11670 -1128
rect 11726 -1184 11780 -1128
rect 11836 -1184 11890 -1128
rect 11946 -1184 12000 -1128
rect 12056 -1184 12110 -1128
rect 12166 -1184 12220 -1128
rect 12276 -1184 12330 -1128
rect 12386 -1184 12429 -1128
rect 10753 -1238 12429 -1184
rect 10753 -1294 10881 -1238
rect 10937 -1294 10991 -1238
rect 11047 -1294 11101 -1238
rect 11157 -1294 11211 -1238
rect 11267 -1294 11321 -1238
rect 11377 -1294 11431 -1238
rect 11487 -1294 11541 -1238
rect 11597 -1294 11670 -1238
rect 11726 -1294 11780 -1238
rect 11836 -1294 11890 -1238
rect 11946 -1294 12000 -1238
rect 12056 -1294 12110 -1238
rect 12166 -1294 12220 -1238
rect 12276 -1294 12330 -1238
rect 12386 -1294 12429 -1238
rect 10753 -1348 12429 -1294
rect 10753 -1404 10881 -1348
rect 10937 -1404 10991 -1348
rect 11047 -1404 11101 -1348
rect 11157 -1404 11211 -1348
rect 11267 -1404 11321 -1348
rect 11377 -1404 11431 -1348
rect 11487 -1404 11541 -1348
rect 11597 -1404 11670 -1348
rect 11726 -1404 11780 -1348
rect 11836 -1404 11890 -1348
rect 11946 -1404 12000 -1348
rect 12056 -1404 12110 -1348
rect 12166 -1404 12220 -1348
rect 12276 -1404 12330 -1348
rect 12386 -1404 12429 -1348
rect 10753 -1458 12429 -1404
rect 10753 -1514 10881 -1458
rect 10937 -1514 10991 -1458
rect 11047 -1514 11101 -1458
rect 11157 -1514 11211 -1458
rect 11267 -1514 11321 -1458
rect 11377 -1514 11431 -1458
rect 11487 -1514 11541 -1458
rect 11597 -1514 11670 -1458
rect 11726 -1514 11780 -1458
rect 11836 -1514 11890 -1458
rect 11946 -1514 12000 -1458
rect 12056 -1514 12110 -1458
rect 12166 -1514 12220 -1458
rect 12276 -1514 12330 -1458
rect 12386 -1514 12429 -1458
rect 10753 -1568 12429 -1514
rect 10753 -1624 10881 -1568
rect 10937 -1624 10991 -1568
rect 11047 -1624 11101 -1568
rect 11157 -1624 11211 -1568
rect 11267 -1624 11321 -1568
rect 11377 -1624 11431 -1568
rect 11487 -1624 11541 -1568
rect 11597 -1624 11670 -1568
rect 11726 -1624 11780 -1568
rect 11836 -1624 11890 -1568
rect 11946 -1624 12000 -1568
rect 12056 -1624 12110 -1568
rect 12166 -1624 12220 -1568
rect 12276 -1624 12330 -1568
rect 12386 -1624 12429 -1568
rect 10753 -1678 12429 -1624
rect 10753 -1734 10881 -1678
rect 10937 -1734 10991 -1678
rect 11047 -1734 11101 -1678
rect 11157 -1734 11211 -1678
rect 11267 -1734 11321 -1678
rect 11377 -1734 11431 -1678
rect 11487 -1734 11541 -1678
rect 11597 -1734 11670 -1678
rect 11726 -1734 11780 -1678
rect 11836 -1734 11890 -1678
rect 11946 -1734 12000 -1678
rect 12056 -1734 12110 -1678
rect 12166 -1734 12220 -1678
rect 12276 -1734 12330 -1678
rect 12386 -1734 12429 -1678
rect 10753 -1870 12429 -1734
rect 22870 1192 23661 1204
rect 22870 1136 22896 1192
rect 22952 1136 23006 1192
rect 23062 1136 23116 1192
rect 23172 1136 23226 1192
rect 23282 1136 23336 1192
rect 23392 1136 23446 1192
rect 23502 1136 23556 1192
rect 23612 1136 23661 1192
rect 22870 1082 23661 1136
rect 22870 1026 22896 1082
rect 22952 1026 23006 1082
rect 23062 1026 23116 1082
rect 23172 1026 23226 1082
rect 23282 1026 23336 1082
rect 23392 1026 23446 1082
rect 23502 1026 23556 1082
rect 23612 1026 23661 1082
rect 22870 972 23661 1026
rect 22870 916 22896 972
rect 22952 916 23006 972
rect 23062 916 23116 972
rect 23172 916 23226 972
rect 23282 916 23336 972
rect 23392 916 23446 972
rect 23502 916 23556 972
rect 23612 916 23661 972
rect 22870 862 23661 916
rect 22870 806 22896 862
rect 22952 806 23006 862
rect 23062 806 23116 862
rect 23172 806 23226 862
rect 23282 806 23336 862
rect 23392 806 23446 862
rect 23502 806 23556 862
rect 23612 806 23661 862
rect 22870 752 23661 806
rect 22870 696 22896 752
rect 22952 696 23006 752
rect 23062 696 23116 752
rect 23172 696 23226 752
rect 23282 696 23336 752
rect 23392 696 23446 752
rect 23502 696 23556 752
rect 23612 696 23661 752
rect 22870 642 23661 696
rect 22870 586 22896 642
rect 22952 586 23006 642
rect 23062 586 23116 642
rect 23172 586 23226 642
rect 23282 586 23336 642
rect 23392 586 23446 642
rect 23502 586 23556 642
rect 23612 586 23661 642
rect 22870 559 23661 586
rect 4762 -2967 7055 -2554
rect 6287 -3034 7055 -2967
rect 6287 -3055 6685 -3034
rect 6486 -3198 6685 -3055
rect 10213 -15012 11793 -14930
rect 10211 -15052 11793 -15012
rect 10211 -15108 10245 -15052
rect 10301 -15108 10355 -15052
rect 10411 -15108 10465 -15052
rect 10521 -15108 10575 -15052
rect 10631 -15108 10685 -15052
rect 10741 -15108 10795 -15052
rect 10851 -15108 10905 -15052
rect 10961 -15108 11034 -15052
rect 11090 -15108 11144 -15052
rect 11200 -15108 11254 -15052
rect 11310 -15108 11364 -15052
rect 11420 -15108 11474 -15052
rect 11530 -15108 11584 -15052
rect 11640 -15108 11694 -15052
rect 11750 -15108 11793 -15052
rect 10211 -15162 11793 -15108
rect 10211 -15218 10245 -15162
rect 10301 -15218 10355 -15162
rect 10411 -15218 10465 -15162
rect 10521 -15218 10575 -15162
rect 10631 -15218 10685 -15162
rect 10741 -15218 10795 -15162
rect 10851 -15218 10905 -15162
rect 10961 -15218 11034 -15162
rect 11090 -15218 11144 -15162
rect 11200 -15218 11254 -15162
rect 11310 -15218 11364 -15162
rect 11420 -15218 11474 -15162
rect 11530 -15218 11584 -15162
rect 11640 -15218 11694 -15162
rect 11750 -15218 11793 -15162
rect 10211 -15272 11793 -15218
rect 10211 -15328 10245 -15272
rect 10301 -15328 10355 -15272
rect 10411 -15328 10465 -15272
rect 10521 -15328 10575 -15272
rect 10631 -15328 10685 -15272
rect 10741 -15328 10795 -15272
rect 10851 -15328 10905 -15272
rect 10961 -15328 11034 -15272
rect 11090 -15328 11144 -15272
rect 11200 -15328 11254 -15272
rect 11310 -15328 11364 -15272
rect 11420 -15328 11474 -15272
rect 11530 -15328 11584 -15272
rect 11640 -15328 11694 -15272
rect 11750 -15328 11793 -15272
rect 10211 -15382 11793 -15328
rect 10211 -15438 10245 -15382
rect 10301 -15438 10355 -15382
rect 10411 -15438 10465 -15382
rect 10521 -15438 10575 -15382
rect 10631 -15438 10685 -15382
rect 10741 -15438 10795 -15382
rect 10851 -15438 10905 -15382
rect 10961 -15438 11034 -15382
rect 11090 -15438 11144 -15382
rect 11200 -15438 11254 -15382
rect 11310 -15438 11364 -15382
rect 11420 -15438 11474 -15382
rect 11530 -15438 11584 -15382
rect 11640 -15438 11694 -15382
rect 11750 -15438 11793 -15382
rect 10211 -15492 11793 -15438
rect 10211 -15548 10245 -15492
rect 10301 -15548 10355 -15492
rect 10411 -15548 10465 -15492
rect 10521 -15548 10575 -15492
rect 10631 -15548 10685 -15492
rect 10741 -15548 10795 -15492
rect 10851 -15548 10905 -15492
rect 10961 -15548 11034 -15492
rect 11090 -15548 11144 -15492
rect 11200 -15548 11254 -15492
rect 11310 -15548 11364 -15492
rect 11420 -15548 11474 -15492
rect 11530 -15548 11584 -15492
rect 11640 -15548 11694 -15492
rect 11750 -15548 11793 -15492
rect 10211 -15602 11793 -15548
rect 10211 -15658 10245 -15602
rect 10301 -15658 10355 -15602
rect 10411 -15658 10465 -15602
rect 10521 -15658 10575 -15602
rect 10631 -15658 10685 -15602
rect 10741 -15658 10795 -15602
rect 10851 -15658 10905 -15602
rect 10961 -15658 11034 -15602
rect 11090 -15658 11144 -15602
rect 11200 -15658 11254 -15602
rect 11310 -15658 11364 -15602
rect 11420 -15658 11474 -15602
rect 11530 -15658 11584 -15602
rect 11640 -15658 11694 -15602
rect 11750 -15658 11793 -15602
rect 10211 -15687 11793 -15658
rect 1185 -18337 1236 -18281
rect 1292 -18337 1346 -18281
rect 1402 -18337 1456 -18281
rect 1512 -18337 1566 -18281
rect 1622 -18337 1676 -18281
rect 1732 -18337 1786 -18281
rect 1842 -18337 1896 -18281
rect 1952 -18337 2118 -18281
rect 1185 -18391 2118 -18337
rect 1185 -18447 1236 -18391
rect 1292 -18447 1346 -18391
rect 1402 -18447 1456 -18391
rect 1512 -18447 1566 -18391
rect 1622 -18447 1676 -18391
rect 1732 -18447 1786 -18391
rect 1842 -18447 1896 -18391
rect 1952 -18447 2118 -18391
rect 1185 -18501 2118 -18447
rect 1185 -18557 1236 -18501
rect 1292 -18557 1346 -18501
rect 1402 -18557 1456 -18501
rect 1512 -18557 1566 -18501
rect 1622 -18557 1676 -18501
rect 1732 -18557 1786 -18501
rect 1842 -18557 1896 -18501
rect 1952 -18557 2118 -18501
rect 1185 -18611 2118 -18557
rect 1185 -18667 1236 -18611
rect 1292 -18667 1346 -18611
rect 1402 -18667 1456 -18611
rect 1512 -18667 1566 -18611
rect 1622 -18667 1676 -18611
rect 1732 -18667 1786 -18611
rect 1842 -18667 1896 -18611
rect 1952 -18667 2118 -18611
rect 1185 -18721 2118 -18667
rect 1185 -18777 1236 -18721
rect 1292 -18777 1346 -18721
rect 1402 -18777 1456 -18721
rect 1512 -18777 1566 -18721
rect 1622 -18777 1676 -18721
rect 1732 -18777 1786 -18721
rect 1842 -18777 1896 -18721
rect 1952 -18777 2118 -18721
rect 1185 -18831 2118 -18777
rect 1185 -18887 1236 -18831
rect 1292 -18887 1346 -18831
rect 1402 -18887 1456 -18831
rect 1512 -18887 1566 -18831
rect 1622 -18887 1676 -18831
rect 1732 -18887 1786 -18831
rect 1842 -18887 1896 -18831
rect 1952 -18887 2118 -18831
rect 1185 -18941 2118 -18887
rect 1185 -18997 1236 -18941
rect 1292 -18997 1346 -18941
rect 1402 -18997 1456 -18941
rect 1512 -18997 1566 -18941
rect 1622 -18997 1676 -18941
rect 1732 -18997 1786 -18941
rect 1842 -18997 1896 -18941
rect 1952 -18997 2118 -18941
rect 1185 -19026 2118 -18997
rect 1189 -19028 2107 -19026
rect 10213 -29695 11793 -15687
rect 21736 -16439 22477 -16409
rect 21736 -16495 21746 -16439
rect 21802 -16495 21856 -16439
rect 21912 -16495 21966 -16439
rect 22022 -16495 22076 -16439
rect 22132 -16495 22186 -16439
rect 22242 -16495 22296 -16439
rect 22352 -16495 22406 -16439
rect 22462 -16495 22477 -16439
rect 21736 -16549 22477 -16495
rect 21736 -16605 21746 -16549
rect 21802 -16605 21856 -16549
rect 21912 -16605 21966 -16549
rect 22022 -16605 22076 -16549
rect 22132 -16605 22186 -16549
rect 22242 -16605 22296 -16549
rect 22352 -16605 22406 -16549
rect 22462 -16605 22477 -16549
rect 21736 -16659 22477 -16605
rect 21736 -16715 21746 -16659
rect 21802 -16715 21856 -16659
rect 21912 -16715 21966 -16659
rect 22022 -16715 22076 -16659
rect 22132 -16715 22186 -16659
rect 22242 -16715 22296 -16659
rect 22352 -16715 22406 -16659
rect 22462 -16715 22477 -16659
rect 21736 -16769 22477 -16715
rect 21736 -16825 21746 -16769
rect 21802 -16825 21856 -16769
rect 21912 -16825 21966 -16769
rect 22022 -16825 22076 -16769
rect 22132 -16825 22186 -16769
rect 22242 -16825 22296 -16769
rect 22352 -16825 22406 -16769
rect 22462 -16825 22477 -16769
rect 21736 -16879 22477 -16825
rect 21736 -16935 21746 -16879
rect 21802 -16935 21856 -16879
rect 21912 -16935 21966 -16879
rect 22022 -16935 22076 -16879
rect 22132 -16935 22186 -16879
rect 22242 -16935 22296 -16879
rect 22352 -16935 22406 -16879
rect 22462 -16935 22477 -16879
rect 21736 -16989 22477 -16935
rect 21736 -17045 21746 -16989
rect 21802 -17045 21856 -16989
rect 21912 -17045 21966 -16989
rect 22022 -17045 22076 -16989
rect 22132 -17045 22186 -16989
rect 22242 -17045 22296 -16989
rect 22352 -17045 22406 -16989
rect 22462 -17045 22477 -16989
rect 21736 -17099 22477 -17045
rect 21736 -17155 21746 -17099
rect 21802 -17155 21856 -17099
rect 21912 -17155 21966 -17099
rect 22022 -17155 22076 -17099
rect 22132 -17155 22186 -17099
rect 22242 -17155 22296 -17099
rect 22352 -17155 22406 -17099
rect 22462 -17155 22477 -17099
rect 15714 -17358 16453 -17330
rect 15714 -17414 15724 -17358
rect 15780 -17414 15834 -17358
rect 15890 -17414 15944 -17358
rect 16000 -17414 16054 -17358
rect 16110 -17414 16164 -17358
rect 16220 -17414 16274 -17358
rect 16330 -17414 16384 -17358
rect 16440 -17414 16453 -17358
rect 15714 -17468 16453 -17414
rect 15714 -17524 15724 -17468
rect 15780 -17524 15834 -17468
rect 15890 -17524 15944 -17468
rect 16000 -17524 16054 -17468
rect 16110 -17524 16164 -17468
rect 16220 -17524 16274 -17468
rect 16330 -17524 16384 -17468
rect 16440 -17524 16453 -17468
rect 15714 -17578 16453 -17524
rect 15714 -17634 15724 -17578
rect 15780 -17634 15834 -17578
rect 15890 -17634 15944 -17578
rect 16000 -17634 16054 -17578
rect 16110 -17634 16164 -17578
rect 16220 -17634 16274 -17578
rect 16330 -17634 16384 -17578
rect 16440 -17634 16453 -17578
rect 15714 -17688 16453 -17634
rect 15714 -17744 15724 -17688
rect 15780 -17744 15834 -17688
rect 15890 -17744 15944 -17688
rect 16000 -17744 16054 -17688
rect 16110 -17744 16164 -17688
rect 16220 -17744 16274 -17688
rect 16330 -17744 16384 -17688
rect 16440 -17744 16453 -17688
rect 15714 -17798 16453 -17744
rect 15714 -17854 15724 -17798
rect 15780 -17854 15834 -17798
rect 15890 -17854 15944 -17798
rect 16000 -17854 16054 -17798
rect 16110 -17854 16164 -17798
rect 16220 -17854 16274 -17798
rect 16330 -17854 16384 -17798
rect 16440 -17854 16453 -17798
rect 15714 -17908 16453 -17854
rect 15714 -17964 15724 -17908
rect 15780 -17964 15834 -17908
rect 15890 -17964 15944 -17908
rect 16000 -17964 16054 -17908
rect 16110 -17964 16164 -17908
rect 16220 -17964 16274 -17908
rect 16330 -17964 16384 -17908
rect 16440 -17964 16453 -17908
rect 15714 -18018 16453 -17964
rect 15714 -18074 15724 -18018
rect 15780 -18074 15834 -18018
rect 15890 -18074 15944 -18018
rect 16000 -18074 16054 -18018
rect 16110 -18074 16164 -18018
rect 16220 -18074 16274 -18018
rect 16330 -18074 16384 -18018
rect 16440 -18074 16453 -18018
rect 15714 -18094 16453 -18074
rect 13160 -19871 13901 -19827
rect 13160 -19927 13167 -19871
rect 13223 -19927 13277 -19871
rect 13333 -19927 13387 -19871
rect 13443 -19927 13497 -19871
rect 13553 -19927 13607 -19871
rect 13663 -19927 13717 -19871
rect 13773 -19927 13827 -19871
rect 13883 -19927 13901 -19871
rect 13160 -19981 13901 -19927
rect 13160 -20037 13167 -19981
rect 13223 -20037 13277 -19981
rect 13333 -20037 13387 -19981
rect 13443 -20037 13497 -19981
rect 13553 -20037 13607 -19981
rect 13663 -20037 13717 -19981
rect 13773 -20037 13827 -19981
rect 13883 -20037 13901 -19981
rect 13160 -20091 13901 -20037
rect 13160 -20147 13167 -20091
rect 13223 -20147 13277 -20091
rect 13333 -20147 13387 -20091
rect 13443 -20147 13497 -20091
rect 13553 -20147 13607 -20091
rect 13663 -20147 13717 -20091
rect 13773 -20147 13827 -20091
rect 13883 -20147 13901 -20091
rect 13160 -20201 13901 -20147
rect 13160 -20257 13167 -20201
rect 13223 -20257 13277 -20201
rect 13333 -20257 13387 -20201
rect 13443 -20257 13497 -20201
rect 13553 -20257 13607 -20201
rect 13663 -20257 13717 -20201
rect 13773 -20257 13827 -20201
rect 13883 -20257 13901 -20201
rect 13160 -20311 13901 -20257
rect 13160 -20367 13167 -20311
rect 13223 -20367 13277 -20311
rect 13333 -20367 13387 -20311
rect 13443 -20367 13497 -20311
rect 13553 -20367 13607 -20311
rect 13663 -20367 13717 -20311
rect 13773 -20367 13827 -20311
rect 13883 -20367 13901 -20311
rect 13160 -20421 13901 -20367
rect 13160 -20477 13167 -20421
rect 13223 -20477 13277 -20421
rect 13333 -20477 13387 -20421
rect 13443 -20477 13497 -20421
rect 13553 -20477 13607 -20421
rect 13663 -20477 13717 -20421
rect 13773 -20477 13827 -20421
rect 13883 -20477 13901 -20421
rect 13160 -20531 13901 -20477
rect 13160 -20587 13167 -20531
rect 13223 -20587 13277 -20531
rect 13333 -20587 13387 -20531
rect 13443 -20587 13497 -20531
rect 13553 -20587 13607 -20531
rect 13663 -20587 13717 -20531
rect 13773 -20587 13827 -20531
rect 13883 -20587 13901 -20531
rect 12266 -20757 13007 -20751
rect 12266 -20813 12283 -20757
rect 12339 -20813 12393 -20757
rect 12449 -20813 12503 -20757
rect 12559 -20813 12613 -20757
rect 12669 -20813 12723 -20757
rect 12779 -20813 12833 -20757
rect 12889 -20813 12943 -20757
rect 12999 -20813 13007 -20757
rect 12266 -20867 13007 -20813
rect 12266 -20923 12283 -20867
rect 12339 -20923 12393 -20867
rect 12449 -20923 12503 -20867
rect 12559 -20923 12613 -20867
rect 12669 -20923 12723 -20867
rect 12779 -20923 12833 -20867
rect 12889 -20923 12943 -20867
rect 12999 -20923 13007 -20867
rect 12266 -20977 13007 -20923
rect 12266 -21033 12283 -20977
rect 12339 -21033 12393 -20977
rect 12449 -21033 12503 -20977
rect 12559 -21033 12613 -20977
rect 12669 -21033 12723 -20977
rect 12779 -21033 12833 -20977
rect 12889 -21033 12943 -20977
rect 12999 -21033 13007 -20977
rect 12266 -21087 13007 -21033
rect 12266 -21143 12283 -21087
rect 12339 -21143 12393 -21087
rect 12449 -21143 12503 -21087
rect 12559 -21143 12613 -21087
rect 12669 -21143 12723 -21087
rect 12779 -21143 12833 -21087
rect 12889 -21143 12943 -21087
rect 12999 -21143 13007 -21087
rect 12266 -21197 13007 -21143
rect 12266 -21253 12283 -21197
rect 12339 -21253 12393 -21197
rect 12449 -21253 12503 -21197
rect 12559 -21253 12613 -21197
rect 12669 -21253 12723 -21197
rect 12779 -21253 12833 -21197
rect 12889 -21253 12943 -21197
rect 12999 -21253 13007 -21197
rect 12266 -21307 13007 -21253
rect 12266 -21363 12283 -21307
rect 12339 -21363 12393 -21307
rect 12449 -21363 12503 -21307
rect 12559 -21363 12613 -21307
rect 12669 -21363 12723 -21307
rect 12779 -21363 12833 -21307
rect 12889 -21363 12943 -21307
rect 12999 -21363 13007 -21307
rect 12266 -21417 13007 -21363
rect 12266 -21473 12283 -21417
rect 12339 -21473 12393 -21417
rect 12449 -21473 12503 -21417
rect 12559 -21473 12613 -21417
rect 12669 -21473 12723 -21417
rect 12779 -21473 12833 -21417
rect 12889 -21473 12943 -21417
rect 12999 -21473 13007 -21417
rect 12266 -28681 13007 -21473
rect 13160 -28255 13901 -20587
rect 15714 -24689 16455 -18094
rect 19487 -19860 20228 -19839
rect 19485 -19872 20228 -19860
rect 19485 -19928 19494 -19872
rect 19550 -19928 19604 -19872
rect 19660 -19928 19714 -19872
rect 19770 -19928 19824 -19872
rect 19880 -19928 19934 -19872
rect 19990 -19928 20044 -19872
rect 20100 -19928 20154 -19872
rect 20210 -19928 20228 -19872
rect 19485 -19982 20228 -19928
rect 19485 -20038 19494 -19982
rect 19550 -20038 19604 -19982
rect 19660 -20038 19714 -19982
rect 19770 -20038 19824 -19982
rect 19880 -20038 19934 -19982
rect 19990 -20038 20044 -19982
rect 20100 -20038 20154 -19982
rect 20210 -20038 20228 -19982
rect 19485 -20092 20228 -20038
rect 19485 -20148 19494 -20092
rect 19550 -20148 19604 -20092
rect 19660 -20148 19714 -20092
rect 19770 -20148 19824 -20092
rect 19880 -20148 19934 -20092
rect 19990 -20148 20044 -20092
rect 20100 -20148 20154 -20092
rect 20210 -20148 20228 -20092
rect 19485 -20202 20228 -20148
rect 19485 -20258 19494 -20202
rect 19550 -20258 19604 -20202
rect 19660 -20258 19714 -20202
rect 19770 -20258 19824 -20202
rect 19880 -20258 19934 -20202
rect 19990 -20258 20044 -20202
rect 20100 -20258 20154 -20202
rect 20210 -20258 20228 -20202
rect 19485 -20312 20228 -20258
rect 19485 -20368 19494 -20312
rect 19550 -20368 19604 -20312
rect 19660 -20368 19714 -20312
rect 19770 -20368 19824 -20312
rect 19880 -20368 19934 -20312
rect 19990 -20368 20044 -20312
rect 20100 -20368 20154 -20312
rect 20210 -20368 20228 -20312
rect 19485 -20422 20228 -20368
rect 19485 -20478 19494 -20422
rect 19550 -20478 19604 -20422
rect 19660 -20478 19714 -20422
rect 19770 -20478 19824 -20422
rect 19880 -20478 19934 -20422
rect 19990 -20478 20044 -20422
rect 20100 -20478 20154 -20422
rect 20210 -20478 20228 -20422
rect 19485 -20532 20228 -20478
rect 19485 -20588 19494 -20532
rect 19550 -20588 19604 -20532
rect 19660 -20588 19714 -20532
rect 19770 -20588 19824 -20532
rect 19880 -20588 19934 -20532
rect 19990 -20588 20044 -20532
rect 20100 -20588 20154 -20532
rect 20210 -20588 20228 -20532
rect 19485 -20593 20228 -20588
rect 18592 -20725 19333 -20719
rect 18591 -20752 19333 -20725
rect 18591 -20808 18599 -20752
rect 18655 -20808 18709 -20752
rect 18765 -20808 18819 -20752
rect 18875 -20808 18929 -20752
rect 18985 -20808 19039 -20752
rect 19095 -20808 19149 -20752
rect 19205 -20808 19259 -20752
rect 19315 -20808 19333 -20752
rect 18591 -20862 19333 -20808
rect 18591 -20918 18599 -20862
rect 18655 -20918 18709 -20862
rect 18765 -20918 18819 -20862
rect 18875 -20918 18929 -20862
rect 18985 -20918 19039 -20862
rect 19095 -20918 19149 -20862
rect 19205 -20918 19259 -20862
rect 19315 -20918 19333 -20862
rect 18591 -20972 19333 -20918
rect 18591 -21028 18599 -20972
rect 18655 -21028 18709 -20972
rect 18765 -21028 18819 -20972
rect 18875 -21028 18929 -20972
rect 18985 -21028 19039 -20972
rect 19095 -21028 19149 -20972
rect 19205 -21028 19259 -20972
rect 19315 -21028 19333 -20972
rect 18591 -21082 19333 -21028
rect 18591 -21138 18599 -21082
rect 18655 -21138 18709 -21082
rect 18765 -21138 18819 -21082
rect 18875 -21138 18929 -21082
rect 18985 -21138 19039 -21082
rect 19095 -21138 19149 -21082
rect 19205 -21138 19259 -21082
rect 19315 -21138 19333 -21082
rect 18591 -21192 19333 -21138
rect 18591 -21248 18599 -21192
rect 18655 -21248 18709 -21192
rect 18765 -21248 18819 -21192
rect 18875 -21248 18929 -21192
rect 18985 -21248 19039 -21192
rect 19095 -21248 19149 -21192
rect 19205 -21248 19259 -21192
rect 19315 -21248 19333 -21192
rect 18591 -21302 19333 -21248
rect 18591 -21358 18599 -21302
rect 18655 -21358 18709 -21302
rect 18765 -21358 18819 -21302
rect 18875 -21358 18929 -21302
rect 18985 -21358 19039 -21302
rect 19095 -21358 19149 -21302
rect 19205 -21358 19259 -21302
rect 19315 -21358 19333 -21302
rect 18591 -21412 19333 -21358
rect 18591 -21468 18599 -21412
rect 18655 -21468 18709 -21412
rect 18765 -21468 18819 -21412
rect 18875 -21468 18929 -21412
rect 18985 -21468 19039 -21412
rect 19095 -21468 19149 -21412
rect 19205 -21468 19259 -21412
rect 19315 -21468 19333 -21412
rect 18591 -21473 19333 -21468
rect 13159 -28608 14611 -28255
rect 18591 -28676 19332 -21473
rect 19485 -28171 20226 -20593
rect 21736 -24703 22477 -17155
rect 22870 -17431 23656 559
rect 24632 159 25532 19239
rect 113495 19860 114395 20024
rect 113495 19804 113574 19860
rect 113630 19804 113684 19860
rect 113740 19804 113794 19860
rect 113850 19804 113904 19860
rect 113960 19804 114014 19860
rect 114070 19804 114124 19860
rect 114180 19804 114234 19860
rect 114290 19804 114395 19860
rect 113495 19750 114395 19804
rect 113495 19694 113574 19750
rect 113630 19694 113684 19750
rect 113740 19694 113794 19750
rect 113850 19694 113904 19750
rect 113960 19694 114014 19750
rect 114070 19694 114124 19750
rect 114180 19694 114234 19750
rect 114290 19694 114395 19750
rect 113495 19640 114395 19694
rect 113495 19584 113574 19640
rect 113630 19584 113684 19640
rect 113740 19584 113794 19640
rect 113850 19584 113904 19640
rect 113960 19584 114014 19640
rect 114070 19584 114124 19640
rect 114180 19584 114234 19640
rect 114290 19584 114395 19640
rect 113495 19530 114395 19584
rect 113495 19474 113574 19530
rect 113630 19474 113684 19530
rect 113740 19474 113794 19530
rect 113850 19474 113904 19530
rect 113960 19474 114014 19530
rect 114070 19474 114124 19530
rect 114180 19474 114234 19530
rect 114290 19474 114395 19530
rect 113495 19420 114395 19474
rect 113495 19364 113574 19420
rect 113630 19364 113684 19420
rect 113740 19364 113794 19420
rect 113850 19364 113904 19420
rect 113960 19364 114014 19420
rect 114070 19364 114124 19420
rect 114180 19364 114234 19420
rect 114290 19364 114395 19420
rect 113495 19310 114395 19364
rect 113495 19254 113574 19310
rect 113630 19254 113684 19310
rect 113740 19254 113794 19310
rect 113850 19254 113904 19310
rect 113960 19254 114014 19310
rect 114070 19254 114124 19310
rect 114180 19254 114234 19310
rect 114290 19254 114395 19310
rect 24632 103 24709 159
rect 24765 103 24819 159
rect 24875 103 24929 159
rect 24985 103 25039 159
rect 25095 103 25149 159
rect 25205 103 25259 159
rect 25315 103 25369 159
rect 25425 103 25532 159
rect 24632 49 25532 103
rect 24632 -7 24709 49
rect 24765 -7 24819 49
rect 24875 -7 24929 49
rect 24985 -7 25039 49
rect 25095 -7 25149 49
rect 25205 -7 25259 49
rect 25315 -7 25369 49
rect 25425 -7 25532 49
rect 24632 -61 25532 -7
rect 24632 -117 24709 -61
rect 24765 -117 24819 -61
rect 24875 -117 24929 -61
rect 24985 -117 25039 -61
rect 25095 -117 25149 -61
rect 25205 -117 25259 -61
rect 25315 -117 25369 -61
rect 25425 -117 25532 -61
rect 24632 -171 25532 -117
rect 24632 -227 24709 -171
rect 24765 -227 24819 -171
rect 24875 -227 24929 -171
rect 24985 -227 25039 -171
rect 25095 -227 25149 -171
rect 25205 -227 25259 -171
rect 25315 -227 25369 -171
rect 25425 -227 25532 -171
rect 24632 -281 25532 -227
rect 24632 -337 24709 -281
rect 24765 -337 24819 -281
rect 24875 -337 24929 -281
rect 24985 -337 25039 -281
rect 25095 -337 25149 -281
rect 25205 -337 25259 -281
rect 25315 -337 25369 -281
rect 25425 -337 25532 -281
rect 24632 -391 25532 -337
rect 24632 -447 24709 -391
rect 24765 -447 24819 -391
rect 24875 -447 24929 -391
rect 24985 -447 25039 -391
rect 25095 -447 25149 -391
rect 25205 -447 25259 -391
rect 25315 -447 25369 -391
rect 25425 -447 25532 -391
rect 24632 -13596 25532 -447
rect 24632 -13652 24679 -13596
rect 24735 -13652 24789 -13596
rect 24845 -13652 24899 -13596
rect 24955 -13652 25009 -13596
rect 25065 -13652 25119 -13596
rect 25175 -13652 25229 -13596
rect 25285 -13652 25339 -13596
rect 25395 -13652 25532 -13596
rect 24632 -13706 25532 -13652
rect 24632 -13762 24679 -13706
rect 24735 -13762 24789 -13706
rect 24845 -13762 24899 -13706
rect 24955 -13762 25009 -13706
rect 25065 -13762 25119 -13706
rect 25175 -13762 25229 -13706
rect 25285 -13762 25339 -13706
rect 25395 -13762 25532 -13706
rect 24632 -13816 25532 -13762
rect 24632 -13872 24679 -13816
rect 24735 -13872 24789 -13816
rect 24845 -13872 24899 -13816
rect 24955 -13872 25009 -13816
rect 25065 -13872 25119 -13816
rect 25175 -13872 25229 -13816
rect 25285 -13872 25339 -13816
rect 25395 -13872 25532 -13816
rect 22870 -17450 23798 -17431
rect 22870 -17454 23387 -17450
rect 22870 -17510 22902 -17454
rect 22958 -17510 23012 -17454
rect 23068 -17510 23122 -17454
rect 23178 -17510 23232 -17454
rect 23288 -17506 23387 -17454
rect 23443 -17506 23497 -17450
rect 23553 -17506 23607 -17450
rect 23663 -17506 23717 -17450
rect 23773 -17506 23798 -17450
rect 23288 -17510 23798 -17506
rect 22870 -17560 23798 -17510
rect 22870 -17564 23387 -17560
rect 22870 -17620 22902 -17564
rect 22958 -17620 23012 -17564
rect 23068 -17620 23122 -17564
rect 23178 -17620 23232 -17564
rect 23288 -17616 23387 -17564
rect 23443 -17616 23497 -17560
rect 23553 -17616 23607 -17560
rect 23663 -17616 23717 -17560
rect 23773 -17616 23798 -17560
rect 23288 -17620 23798 -17616
rect 22870 -17670 23798 -17620
rect 22870 -17674 23387 -17670
rect 22870 -17730 22902 -17674
rect 22958 -17730 23012 -17674
rect 23068 -17730 23122 -17674
rect 23178 -17730 23232 -17674
rect 23288 -17726 23387 -17674
rect 23443 -17726 23497 -17670
rect 23553 -17726 23607 -17670
rect 23663 -17726 23717 -17670
rect 23773 -17726 23798 -17670
rect 23288 -17730 23798 -17726
rect 22870 -17780 23798 -17730
rect 22870 -17784 23387 -17780
rect 22870 -17840 22902 -17784
rect 22958 -17840 23012 -17784
rect 23068 -17840 23122 -17784
rect 23178 -17840 23232 -17784
rect 23288 -17836 23387 -17784
rect 23443 -17836 23497 -17780
rect 23553 -17836 23607 -17780
rect 23663 -17836 23717 -17780
rect 23773 -17836 23798 -17780
rect 23288 -17840 23798 -17836
rect 22870 -17877 23798 -17840
rect 22870 -17878 23656 -17877
rect 23189 -17879 23656 -17878
rect 24632 -23938 25532 -13872
rect 25861 18616 26761 18785
rect 25861 18560 25931 18616
rect 25987 18560 26041 18616
rect 26097 18560 26151 18616
rect 26207 18560 26261 18616
rect 26317 18560 26371 18616
rect 26427 18560 26481 18616
rect 26537 18560 26591 18616
rect 26647 18560 26761 18616
rect 25861 18506 26761 18560
rect 25861 18450 25931 18506
rect 25987 18450 26041 18506
rect 26097 18450 26151 18506
rect 26207 18450 26261 18506
rect 26317 18450 26371 18506
rect 26427 18450 26481 18506
rect 26537 18450 26591 18506
rect 26647 18450 26761 18506
rect 25861 18396 26761 18450
rect 25861 18340 25931 18396
rect 25987 18340 26041 18396
rect 26097 18340 26151 18396
rect 26207 18340 26261 18396
rect 26317 18340 26371 18396
rect 26427 18340 26481 18396
rect 26537 18340 26591 18396
rect 26647 18340 26761 18396
rect 25861 18286 26761 18340
rect 25861 18230 25931 18286
rect 25987 18230 26041 18286
rect 26097 18230 26151 18286
rect 26207 18230 26261 18286
rect 26317 18230 26371 18286
rect 26427 18230 26481 18286
rect 26537 18230 26591 18286
rect 26647 18230 26761 18286
rect 25861 18176 26761 18230
rect 25861 18120 25931 18176
rect 25987 18120 26041 18176
rect 26097 18120 26151 18176
rect 26207 18120 26261 18176
rect 26317 18120 26371 18176
rect 26427 18120 26481 18176
rect 26537 18120 26591 18176
rect 26647 18120 26761 18176
rect 25861 18066 26761 18120
rect 25861 18010 25931 18066
rect 25987 18010 26041 18066
rect 26097 18010 26151 18066
rect 26207 18010 26261 18066
rect 26317 18010 26371 18066
rect 26427 18010 26481 18066
rect 26537 18010 26591 18066
rect 26647 18010 26761 18066
rect 25861 -1146 26761 18010
rect 112010 17222 112992 17430
rect 112010 17166 112156 17222
rect 112212 17166 112266 17222
rect 112322 17166 112376 17222
rect 112432 17166 112486 17222
rect 112542 17166 112596 17222
rect 112652 17166 112706 17222
rect 112762 17166 112816 17222
rect 112872 17166 112992 17222
rect 112010 17112 112992 17166
rect 112010 17056 112156 17112
rect 112212 17056 112266 17112
rect 112322 17056 112376 17112
rect 112432 17056 112486 17112
rect 112542 17056 112596 17112
rect 112652 17056 112706 17112
rect 112762 17056 112816 17112
rect 112872 17056 112992 17112
rect 112010 17002 112992 17056
rect 112010 16946 112156 17002
rect 112212 16946 112266 17002
rect 112322 16946 112376 17002
rect 112432 16946 112486 17002
rect 112542 16946 112596 17002
rect 112652 16946 112706 17002
rect 112762 16946 112816 17002
rect 112872 16946 112992 17002
rect 112010 16892 112992 16946
rect 112010 16836 112156 16892
rect 112212 16836 112266 16892
rect 112322 16836 112376 16892
rect 112432 16836 112486 16892
rect 112542 16836 112596 16892
rect 112652 16836 112706 16892
rect 112762 16836 112816 16892
rect 112872 16836 112992 16892
rect 112010 16782 112992 16836
rect 112010 16726 112156 16782
rect 112212 16726 112266 16782
rect 112322 16726 112376 16782
rect 112432 16726 112486 16782
rect 112542 16726 112596 16782
rect 112652 16726 112706 16782
rect 112762 16726 112816 16782
rect 112872 16726 112992 16782
rect 112010 16672 112992 16726
rect 112010 16616 112156 16672
rect 112212 16616 112266 16672
rect 112322 16616 112376 16672
rect 112432 16616 112486 16672
rect 112542 16616 112596 16672
rect 112652 16616 112706 16672
rect 112762 16616 112816 16672
rect 112872 16616 112992 16672
rect 112010 16562 112992 16616
rect 112010 16506 112156 16562
rect 112212 16506 112266 16562
rect 112322 16506 112376 16562
rect 112432 16506 112486 16562
rect 112542 16506 112596 16562
rect 112652 16506 112706 16562
rect 112762 16506 112816 16562
rect 112872 16506 112992 16562
rect 27299 10665 27726 10700
rect 27299 10609 27330 10665
rect 27386 10609 27440 10665
rect 27496 10609 27550 10665
rect 27606 10609 27660 10665
rect 27716 10609 27726 10665
rect 27299 10555 27726 10609
rect 27299 10499 27330 10555
rect 27386 10499 27440 10555
rect 27496 10499 27550 10555
rect 27606 10499 27660 10555
rect 27716 10499 27726 10555
rect 27299 10445 27726 10499
rect 27299 10389 27330 10445
rect 27386 10389 27440 10445
rect 27496 10389 27550 10445
rect 27606 10389 27660 10445
rect 27716 10389 27726 10445
rect 27299 10335 27726 10389
rect 27299 10279 27330 10335
rect 27386 10279 27440 10335
rect 27496 10279 27550 10335
rect 27606 10279 27660 10335
rect 27716 10279 27726 10335
rect 27299 10225 27726 10279
rect 27299 10169 27330 10225
rect 27386 10169 27440 10225
rect 27496 10169 27550 10225
rect 27606 10169 27660 10225
rect 27716 10169 27726 10225
rect 27299 10115 27726 10169
rect 27299 10059 27330 10115
rect 27386 10059 27440 10115
rect 27496 10059 27550 10115
rect 27606 10059 27660 10115
rect 27716 10059 27726 10115
rect 27299 10005 27726 10059
rect 27299 9949 27330 10005
rect 27386 9949 27440 10005
rect 27496 9949 27550 10005
rect 27606 9949 27660 10005
rect 27716 9949 27726 10005
rect 27299 9895 27726 9949
rect 27299 9839 27330 9895
rect 27386 9839 27440 9895
rect 27496 9839 27550 9895
rect 27606 9839 27660 9895
rect 27716 9839 27726 9895
rect 27299 9773 27726 9839
rect 25861 -1202 25927 -1146
rect 25983 -1202 26037 -1146
rect 26093 -1202 26147 -1146
rect 26203 -1202 26257 -1146
rect 26313 -1202 26367 -1146
rect 26423 -1202 26477 -1146
rect 26533 -1202 26587 -1146
rect 26643 -1202 26761 -1146
rect 25861 -1256 26761 -1202
rect 25861 -1312 25927 -1256
rect 25983 -1312 26037 -1256
rect 26093 -1312 26147 -1256
rect 26203 -1312 26257 -1256
rect 26313 -1312 26367 -1256
rect 26423 -1312 26477 -1256
rect 26533 -1312 26587 -1256
rect 26643 -1312 26761 -1256
rect 25861 -1366 26761 -1312
rect 25861 -1422 25927 -1366
rect 25983 -1422 26037 -1366
rect 26093 -1422 26147 -1366
rect 26203 -1422 26257 -1366
rect 26313 -1422 26367 -1366
rect 26423 -1422 26477 -1366
rect 26533 -1422 26587 -1366
rect 26643 -1422 26761 -1366
rect 25861 -1476 26761 -1422
rect 25861 -1532 25927 -1476
rect 25983 -1532 26037 -1476
rect 26093 -1532 26147 -1476
rect 26203 -1532 26257 -1476
rect 26313 -1532 26367 -1476
rect 26423 -1532 26477 -1476
rect 26533 -1532 26587 -1476
rect 26643 -1532 26761 -1476
rect 25861 -1586 26761 -1532
rect 25861 -1642 25927 -1586
rect 25983 -1642 26037 -1586
rect 26093 -1642 26147 -1586
rect 26203 -1642 26257 -1586
rect 26313 -1642 26367 -1586
rect 26423 -1642 26477 -1586
rect 26533 -1642 26587 -1586
rect 26643 -1642 26761 -1586
rect 25861 -1696 26761 -1642
rect 25861 -1752 25927 -1696
rect 25983 -1752 26037 -1696
rect 26093 -1752 26147 -1696
rect 26203 -1752 26257 -1696
rect 26313 -1752 26367 -1696
rect 26423 -1752 26477 -1696
rect 26533 -1752 26587 -1696
rect 26643 -1752 26761 -1696
rect 25861 -4107 26761 -1752
rect 25861 -4146 26762 -4107
rect 25861 -4147 26470 -4146
rect 25861 -4203 25883 -4147
rect 25939 -4203 25993 -4147
rect 26049 -4203 26103 -4147
rect 26159 -4203 26213 -4147
rect 26269 -4203 26323 -4147
rect 26379 -4202 26470 -4147
rect 26526 -4202 26580 -4146
rect 26636 -4202 26690 -4146
rect 26746 -4202 26762 -4146
rect 26379 -4203 26762 -4202
rect 25861 -4256 26762 -4203
rect 25861 -4257 26470 -4256
rect 25861 -4313 25883 -4257
rect 25939 -4313 25993 -4257
rect 26049 -4313 26103 -4257
rect 26159 -4313 26213 -4257
rect 26269 -4313 26323 -4257
rect 26379 -4312 26470 -4257
rect 26526 -4312 26580 -4256
rect 26636 -4312 26690 -4256
rect 26746 -4312 26762 -4256
rect 26379 -4313 26762 -4312
rect 25861 -4351 26762 -4313
rect 25861 -14420 26761 -4351
rect 25861 -14476 25904 -14420
rect 25960 -14476 26014 -14420
rect 26070 -14476 26124 -14420
rect 26180 -14476 26234 -14420
rect 26290 -14476 26344 -14420
rect 26400 -14476 26454 -14420
rect 26510 -14476 26564 -14420
rect 26620 -14476 26761 -14420
rect 25861 -14530 26761 -14476
rect 25861 -14586 25904 -14530
rect 25960 -14586 26014 -14530
rect 26070 -14586 26124 -14530
rect 26180 -14586 26234 -14530
rect 26290 -14586 26344 -14530
rect 26400 -14586 26454 -14530
rect 26510 -14586 26564 -14530
rect 26620 -14586 26761 -14530
rect 25861 -14640 26761 -14586
rect 25861 -14696 25904 -14640
rect 25960 -14696 26014 -14640
rect 26070 -14696 26124 -14640
rect 26180 -14696 26234 -14640
rect 26290 -14696 26344 -14640
rect 26400 -14696 26454 -14640
rect 26510 -14696 26564 -14640
rect 26620 -14696 26761 -14640
rect 25861 -21402 26761 -14696
rect 25859 -21422 26761 -21402
rect 25859 -21478 25916 -21422
rect 25972 -21478 26026 -21422
rect 26082 -21478 26136 -21422
rect 26192 -21478 26246 -21422
rect 26302 -21478 26356 -21422
rect 26412 -21478 26466 -21422
rect 26522 -21478 26576 -21422
rect 26632 -21478 26761 -21422
rect 25859 -21532 26761 -21478
rect 25859 -21588 25916 -21532
rect 25972 -21588 26026 -21532
rect 26082 -21588 26136 -21532
rect 26192 -21588 26246 -21532
rect 26302 -21588 26356 -21532
rect 26412 -21588 26466 -21532
rect 26522 -21588 26576 -21532
rect 26632 -21588 26761 -21532
rect 25859 -21642 26761 -21588
rect 25859 -21698 25916 -21642
rect 25972 -21698 26026 -21642
rect 26082 -21698 26136 -21642
rect 26192 -21698 26246 -21642
rect 26302 -21698 26356 -21642
rect 26412 -21698 26466 -21642
rect 26522 -21698 26576 -21642
rect 26632 -21698 26761 -21642
rect 25859 -21770 26761 -21698
rect 24632 -23994 24635 -23938
rect 24691 -23994 24745 -23938
rect 24801 -23994 24855 -23938
rect 24911 -23994 24965 -23938
rect 25021 -23994 25075 -23938
rect 25131 -23994 25185 -23938
rect 25241 -23994 25295 -23938
rect 25351 -23994 25405 -23938
rect 25461 -23994 25532 -23938
rect 24632 -24048 25532 -23994
rect 24632 -24104 24635 -24048
rect 24691 -24104 24745 -24048
rect 24801 -24104 24855 -24048
rect 24911 -24104 24965 -24048
rect 25021 -24104 25075 -24048
rect 25131 -24104 25185 -24048
rect 25241 -24104 25295 -24048
rect 25351 -24104 25405 -24048
rect 25461 -24104 25532 -24048
rect 24632 -24158 25532 -24104
rect 24632 -24214 24635 -24158
rect 24691 -24214 24745 -24158
rect 24801 -24214 24855 -24158
rect 24911 -24214 24965 -24158
rect 25021 -24214 25075 -24158
rect 25131 -24214 25185 -24158
rect 25241 -24214 25295 -24158
rect 25351 -24214 25405 -24158
rect 25461 -24214 25532 -24158
rect 24632 -24268 25532 -24214
rect 24632 -24324 24635 -24268
rect 24691 -24324 24745 -24268
rect 24801 -24324 24855 -24268
rect 24911 -24324 24965 -24268
rect 25021 -24324 25075 -24268
rect 25131 -24324 25185 -24268
rect 25241 -24324 25295 -24268
rect 25351 -24324 25405 -24268
rect 25461 -24324 25532 -24268
rect 24632 -24378 25532 -24324
rect 24632 -24434 24635 -24378
rect 24691 -24434 24745 -24378
rect 24801 -24434 24855 -24378
rect 24911 -24434 24965 -24378
rect 25021 -24434 25075 -24378
rect 25131 -24434 25185 -24378
rect 25241 -24434 25295 -24378
rect 25351 -24434 25405 -24378
rect 25461 -24434 25532 -24378
rect 24632 -24488 25532 -24434
rect 24632 -24544 24635 -24488
rect 24691 -24544 24745 -24488
rect 24801 -24544 24855 -24488
rect 24911 -24544 24965 -24488
rect 25021 -24544 25075 -24488
rect 25131 -24544 25185 -24488
rect 25241 -24544 25295 -24488
rect 25351 -24544 25405 -24488
rect 25461 -24544 25532 -24488
rect 19485 -28529 20758 -28171
rect 12261 -29090 14643 -28681
rect 18591 -28889 20708 -28676
rect 18592 -29022 20708 -28889
rect 10213 -29751 10249 -29695
rect 10305 -29751 10359 -29695
rect 10415 -29751 10469 -29695
rect 10525 -29751 10579 -29695
rect 10635 -29751 10689 -29695
rect 10745 -29751 10799 -29695
rect 10855 -29751 10909 -29695
rect 10965 -29751 11038 -29695
rect 11094 -29751 11148 -29695
rect 11204 -29751 11258 -29695
rect 11314 -29751 11368 -29695
rect 11424 -29751 11478 -29695
rect 11534 -29751 11588 -29695
rect 11644 -29751 11698 -29695
rect 11754 -29751 11793 -29695
rect 10213 -29805 11793 -29751
rect 10213 -29861 10249 -29805
rect 10305 -29861 10359 -29805
rect 10415 -29861 10469 -29805
rect 10525 -29861 10579 -29805
rect 10635 -29861 10689 -29805
rect 10745 -29861 10799 -29805
rect 10855 -29861 10909 -29805
rect 10965 -29861 11038 -29805
rect 11094 -29861 11148 -29805
rect 11204 -29861 11258 -29805
rect 11314 -29861 11368 -29805
rect 11424 -29861 11478 -29805
rect 11534 -29861 11588 -29805
rect 11644 -29861 11698 -29805
rect 11754 -29861 11793 -29805
rect 10213 -29915 11793 -29861
rect 10213 -29971 10249 -29915
rect 10305 -29971 10359 -29915
rect 10415 -29971 10469 -29915
rect 10525 -29971 10579 -29915
rect 10635 -29971 10689 -29915
rect 10745 -29971 10799 -29915
rect 10855 -29971 10909 -29915
rect 10965 -29971 11038 -29915
rect 11094 -29971 11148 -29915
rect 11204 -29971 11258 -29915
rect 11314 -29971 11368 -29915
rect 11424 -29971 11478 -29915
rect 11534 -29971 11588 -29915
rect 11644 -29971 11698 -29915
rect 11754 -29971 11793 -29915
rect 10213 -30025 11793 -29971
rect 10213 -30081 10249 -30025
rect 10305 -30081 10359 -30025
rect 10415 -30081 10469 -30025
rect 10525 -30081 10579 -30025
rect 10635 -30081 10689 -30025
rect 10745 -30081 10799 -30025
rect 10855 -30081 10909 -30025
rect 10965 -30081 11038 -30025
rect 11094 -30081 11148 -30025
rect 11204 -30081 11258 -30025
rect 11314 -30081 11368 -30025
rect 11424 -30081 11478 -30025
rect 11534 -30081 11588 -30025
rect 11644 -30081 11698 -30025
rect 11754 -30081 11793 -30025
rect 10213 -31672 11793 -30081
rect 24632 -30497 25532 -24544
rect 24632 -30553 24746 -30497
rect 24802 -30553 24856 -30497
rect 24912 -30553 24966 -30497
rect 25022 -30553 25076 -30497
rect 25132 -30553 25186 -30497
rect 25242 -30553 25296 -30497
rect 25352 -30553 25406 -30497
rect 25462 -30553 25532 -30497
rect 24632 -30607 25532 -30553
rect 24632 -30663 24746 -30607
rect 24802 -30663 24856 -30607
rect 24912 -30663 24966 -30607
rect 25022 -30663 25076 -30607
rect 25132 -30663 25186 -30607
rect 25242 -30663 25296 -30607
rect 25352 -30663 25406 -30607
rect 25462 -30663 25532 -30607
rect 24632 -30717 25532 -30663
rect 24632 -30773 24746 -30717
rect 24802 -30773 24856 -30717
rect 24912 -30773 24966 -30717
rect 25022 -30773 25076 -30717
rect 25132 -30773 25186 -30717
rect 25242 -30773 25296 -30717
rect 25352 -30773 25406 -30717
rect 25462 -30773 25532 -30717
rect 24632 -30827 25532 -30773
rect 24632 -30883 24746 -30827
rect 24802 -30883 24856 -30827
rect 24912 -30883 24966 -30827
rect 25022 -30883 25076 -30827
rect 25132 -30883 25186 -30827
rect 25242 -30883 25296 -30827
rect 25352 -30883 25406 -30827
rect 25462 -30883 25532 -30827
rect 24632 -30937 25532 -30883
rect 24632 -30993 24746 -30937
rect 24802 -30993 24856 -30937
rect 24912 -30993 24966 -30937
rect 25022 -30993 25076 -30937
rect 25132 -30993 25186 -30937
rect 25242 -30993 25296 -30937
rect 25352 -30993 25406 -30937
rect 25462 -30993 25532 -30937
rect 24632 -31047 25532 -30993
rect 24632 -31103 24746 -31047
rect 24802 -31103 24856 -31047
rect 24912 -31103 24966 -31047
rect 25022 -31103 25076 -31047
rect 25132 -31103 25186 -31047
rect 25242 -31103 25296 -31047
rect 25352 -31103 25406 -31047
rect 25462 -31103 25532 -31047
rect 24632 -31293 25532 -31103
rect 10213 -31728 10247 -31672
rect 10303 -31728 10357 -31672
rect 10413 -31728 10467 -31672
rect 10523 -31728 10577 -31672
rect 10633 -31728 10687 -31672
rect 10743 -31728 10797 -31672
rect 10853 -31728 10907 -31672
rect 10963 -31728 11036 -31672
rect 11092 -31728 11146 -31672
rect 11202 -31728 11256 -31672
rect 11312 -31728 11366 -31672
rect 11422 -31728 11476 -31672
rect 11532 -31728 11586 -31672
rect 11642 -31728 11696 -31672
rect 11752 -31728 11793 -31672
rect 10213 -31782 11793 -31728
rect 10213 -31838 10247 -31782
rect 10303 -31838 10357 -31782
rect 10413 -31838 10467 -31782
rect 10523 -31838 10577 -31782
rect 10633 -31838 10687 -31782
rect 10743 -31838 10797 -31782
rect 10853 -31838 10907 -31782
rect 10963 -31838 11036 -31782
rect 11092 -31838 11146 -31782
rect 11202 -31838 11256 -31782
rect 11312 -31838 11366 -31782
rect 11422 -31838 11476 -31782
rect 11532 -31838 11586 -31782
rect 11642 -31838 11696 -31782
rect 11752 -31838 11793 -31782
rect 10213 -31892 11793 -31838
rect 10213 -31948 10247 -31892
rect 10303 -31948 10357 -31892
rect 10413 -31948 10467 -31892
rect 10523 -31948 10577 -31892
rect 10633 -31948 10687 -31892
rect 10743 -31948 10797 -31892
rect 10853 -31948 10907 -31892
rect 10963 -31948 11036 -31892
rect 11092 -31948 11146 -31892
rect 11202 -31948 11256 -31892
rect 11312 -31948 11366 -31892
rect 11422 -31948 11476 -31892
rect 11532 -31948 11586 -31892
rect 11642 -31948 11696 -31892
rect 11752 -31948 11793 -31892
rect 10213 -32002 11793 -31948
rect 10213 -32058 10247 -32002
rect 10303 -32058 10357 -32002
rect 10413 -32058 10467 -32002
rect 10523 -32058 10577 -32002
rect 10633 -32058 10687 -32002
rect 10743 -32058 10797 -32002
rect 10853 -32058 10907 -32002
rect 10963 -32058 11036 -32002
rect 11092 -32058 11146 -32002
rect 11202 -32058 11256 -32002
rect 11312 -32058 11366 -32002
rect 11422 -32058 11476 -32002
rect 11532 -32058 11586 -32002
rect 11642 -32058 11696 -32002
rect 11752 -32058 11793 -32002
rect 10213 -32112 11793 -32058
rect 10213 -32168 10247 -32112
rect 10303 -32168 10357 -32112
rect 10413 -32168 10467 -32112
rect 10523 -32168 10577 -32112
rect 10633 -32168 10687 -32112
rect 10743 -32168 10797 -32112
rect 10853 -32168 10907 -32112
rect 10963 -32168 11036 -32112
rect 11092 -32168 11146 -32112
rect 11202 -32168 11256 -32112
rect 11312 -32168 11366 -32112
rect 11422 -32168 11476 -32112
rect 11532 -32168 11586 -32112
rect 11642 -32168 11696 -32112
rect 11752 -32168 11793 -32112
rect 10213 -32222 11793 -32168
rect 10213 -32278 10247 -32222
rect 10303 -32278 10357 -32222
rect 10413 -32278 10467 -32222
rect 10523 -32278 10577 -32222
rect 10633 -32278 10687 -32222
rect 10743 -32278 10797 -32222
rect 10853 -32278 10907 -32222
rect 10963 -32278 11036 -32222
rect 11092 -32278 11146 -32222
rect 11202 -32278 11256 -32222
rect 11312 -32278 11366 -32222
rect 11422 -32278 11476 -32222
rect 11532 -32278 11586 -32222
rect 11642 -32278 11696 -32222
rect 11752 -32278 11793 -32222
rect 10213 -32361 11793 -32278
rect 25861 -31614 26761 -21770
rect 27246 -7685 27775 6908
rect 107175 6784 107963 6804
rect 107175 6728 107204 6784
rect 107260 6728 107314 6784
rect 107370 6728 107424 6784
rect 107480 6728 107534 6784
rect 107590 6728 107644 6784
rect 107700 6728 107754 6784
rect 107810 6728 107864 6784
rect 107920 6728 107963 6784
rect 107175 6674 107963 6728
rect 107175 6618 107204 6674
rect 107260 6618 107314 6674
rect 107370 6618 107424 6674
rect 107480 6618 107534 6674
rect 107590 6618 107644 6674
rect 107700 6618 107754 6674
rect 107810 6618 107864 6674
rect 107920 6618 107963 6674
rect 107175 6564 107963 6618
rect 107175 6508 107204 6564
rect 107260 6508 107314 6564
rect 107370 6508 107424 6564
rect 107480 6508 107534 6564
rect 107590 6508 107644 6564
rect 107700 6508 107754 6564
rect 107810 6508 107864 6564
rect 107920 6508 107963 6564
rect 107175 6454 107963 6508
rect 107175 6398 107204 6454
rect 107260 6398 107314 6454
rect 107370 6398 107424 6454
rect 107480 6398 107534 6454
rect 107590 6398 107644 6454
rect 107700 6398 107754 6454
rect 107810 6398 107864 6454
rect 107920 6398 107963 6454
rect 107175 6344 107963 6398
rect 46858 6314 46914 6319
rect 46392 6309 46957 6314
rect 43879 6293 44495 6294
rect 43879 6250 44498 6293
rect 43879 6194 43928 6250
rect 43984 6194 44038 6250
rect 44094 6194 44148 6250
rect 44204 6194 44258 6250
rect 44314 6194 44368 6250
rect 44424 6194 44498 6250
rect 30985 6145 31774 6185
rect 30985 6135 31776 6145
rect 30985 6079 31032 6135
rect 31088 6079 31142 6135
rect 31198 6079 31252 6135
rect 31308 6079 31362 6135
rect 31418 6079 31472 6135
rect 31528 6079 31582 6135
rect 31638 6079 31692 6135
rect 31748 6079 31776 6135
rect 30985 6025 31776 6079
rect 30985 5969 31032 6025
rect 31088 5969 31142 6025
rect 31198 5969 31252 6025
rect 31308 5969 31362 6025
rect 31418 5969 31472 6025
rect 31528 5969 31582 6025
rect 31638 5969 31692 6025
rect 31748 5969 31776 6025
rect 30985 5915 31776 5969
rect 43879 6140 44498 6194
rect 43879 6084 43928 6140
rect 43984 6084 44038 6140
rect 44094 6084 44148 6140
rect 44204 6084 44258 6140
rect 44314 6084 44368 6140
rect 44424 6084 44498 6140
rect 43879 6030 44498 6084
rect 43879 5974 43928 6030
rect 43984 5974 44038 6030
rect 44094 5974 44148 6030
rect 44204 5974 44258 6030
rect 44314 5974 44368 6030
rect 44424 5998 44498 6030
rect 46392 6253 46418 6309
rect 46474 6253 46528 6309
rect 46584 6253 46638 6309
rect 46694 6253 46748 6309
rect 46804 6253 46858 6309
rect 46914 6290 46957 6309
rect 46914 6253 46958 6290
rect 46392 6199 46958 6253
rect 46392 6198 46638 6199
rect 46392 6197 46530 6198
rect 46392 6141 46421 6197
rect 46477 6142 46530 6197
rect 46586 6143 46638 6198
rect 46694 6143 46748 6199
rect 46804 6143 46858 6199
rect 46914 6143 46958 6199
rect 46586 6142 46958 6143
rect 46477 6141 46958 6142
rect 46392 6092 46958 6141
rect 46392 6091 46527 6092
rect 46392 6035 46421 6091
rect 46477 6036 46527 6091
rect 46583 6089 46958 6092
rect 46583 6036 46638 6089
rect 46477 6035 46638 6036
rect 46392 6033 46638 6035
rect 46694 6033 46748 6089
rect 46804 6033 46858 6089
rect 46914 6033 46958 6089
rect 44424 5974 44495 5998
rect 46392 5996 46958 6033
rect 107175 6288 107204 6344
rect 107260 6288 107314 6344
rect 107370 6288 107424 6344
rect 107480 6288 107534 6344
rect 107590 6288 107644 6344
rect 107700 6288 107754 6344
rect 107810 6288 107864 6344
rect 107920 6288 107963 6344
rect 107175 6234 107963 6288
rect 107175 6178 107204 6234
rect 107260 6178 107314 6234
rect 107370 6178 107424 6234
rect 107480 6178 107534 6234
rect 107590 6178 107644 6234
rect 107700 6178 107754 6234
rect 107810 6178 107864 6234
rect 107920 6178 107963 6234
rect 107175 6124 107963 6178
rect 107175 6068 107204 6124
rect 107260 6068 107314 6124
rect 107370 6068 107424 6124
rect 107480 6068 107534 6124
rect 107590 6068 107644 6124
rect 107700 6068 107754 6124
rect 107810 6068 107864 6124
rect 107920 6068 107963 6124
rect 107175 6014 107963 6068
rect 43879 5958 44495 5974
rect 107175 5958 107204 6014
rect 107260 5958 107314 6014
rect 107370 5958 107424 6014
rect 107480 5958 107534 6014
rect 107590 5958 107644 6014
rect 107700 5958 107754 6014
rect 107810 5958 107864 6014
rect 107920 5958 107963 6014
rect 30985 5859 31032 5915
rect 31088 5859 31142 5915
rect 31198 5859 31252 5915
rect 31308 5859 31362 5915
rect 31418 5859 31472 5915
rect 31528 5859 31582 5915
rect 31638 5859 31692 5915
rect 31748 5859 31776 5915
rect 30985 5805 31776 5859
rect 30985 5749 31032 5805
rect 31088 5749 31142 5805
rect 31198 5749 31252 5805
rect 31308 5749 31362 5805
rect 31418 5749 31472 5805
rect 31528 5749 31582 5805
rect 31638 5749 31692 5805
rect 31748 5749 31776 5805
rect 30985 5695 31776 5749
rect 30985 5639 31032 5695
rect 31088 5639 31142 5695
rect 31198 5639 31252 5695
rect 31308 5639 31362 5695
rect 31418 5639 31472 5695
rect 31528 5639 31582 5695
rect 31638 5639 31692 5695
rect 31748 5639 31776 5695
rect 30985 5585 31776 5639
rect 30985 5529 31032 5585
rect 31088 5529 31142 5585
rect 31198 5529 31252 5585
rect 31308 5529 31362 5585
rect 31418 5529 31472 5585
rect 31528 5529 31582 5585
rect 31638 5529 31692 5585
rect 31748 5529 31776 5585
rect 30985 5475 31776 5529
rect 30985 5419 31032 5475
rect 31088 5419 31142 5475
rect 31198 5419 31252 5475
rect 31308 5419 31362 5475
rect 31418 5419 31472 5475
rect 31528 5419 31582 5475
rect 31638 5419 31692 5475
rect 31748 5419 31776 5475
rect 30985 5382 31776 5419
rect 28340 1188 29128 1206
rect 28340 1132 28369 1188
rect 28425 1132 28479 1188
rect 28535 1132 28589 1188
rect 28645 1132 28699 1188
rect 28755 1132 28809 1188
rect 28865 1132 28919 1188
rect 28975 1132 29029 1188
rect 29085 1132 29128 1188
rect 28340 1078 29128 1132
rect 28340 1022 28369 1078
rect 28425 1022 28479 1078
rect 28535 1022 28589 1078
rect 28645 1022 28699 1078
rect 28755 1022 28809 1078
rect 28865 1022 28919 1078
rect 28975 1022 29029 1078
rect 29085 1022 29128 1078
rect 28340 968 29128 1022
rect 28340 912 28369 968
rect 28425 912 28479 968
rect 28535 912 28589 968
rect 28645 912 28699 968
rect 28755 912 28809 968
rect 28865 912 28919 968
rect 28975 912 29029 968
rect 29085 912 29128 968
rect 28340 858 29128 912
rect 28340 802 28369 858
rect 28425 802 28479 858
rect 28535 802 28589 858
rect 28645 802 28699 858
rect 28755 802 28809 858
rect 28865 802 28919 858
rect 28975 802 29029 858
rect 29085 802 29128 858
rect 28340 748 29128 802
rect 28340 692 28369 748
rect 28425 692 28479 748
rect 28535 692 28589 748
rect 28645 692 28699 748
rect 28755 692 28809 748
rect 28865 692 28919 748
rect 28975 692 29029 748
rect 29085 692 29128 748
rect 28340 638 29128 692
rect 28340 582 28369 638
rect 28425 582 28479 638
rect 28535 582 28589 638
rect 28645 582 28699 638
rect 28755 582 28809 638
rect 28865 582 28919 638
rect 28975 582 29029 638
rect 29085 582 29128 638
rect 28340 -82 29128 582
rect 28339 -195 29128 -82
rect 29761 214 30663 374
rect 29761 158 29849 214
rect 29905 158 29959 214
rect 30015 158 30069 214
rect 30125 158 30179 214
rect 30235 158 30289 214
rect 30345 158 30399 214
rect 30455 158 30509 214
rect 30565 158 30663 214
rect 29761 104 30663 158
rect 29761 48 29849 104
rect 29905 48 29959 104
rect 30015 48 30069 104
rect 30125 48 30179 104
rect 30235 48 30289 104
rect 30345 48 30399 104
rect 30455 48 30509 104
rect 30565 48 30663 104
rect 29761 -6 30663 48
rect 29761 -62 29849 -6
rect 29905 -62 29959 -6
rect 30015 -62 30069 -6
rect 30125 -62 30179 -6
rect 30235 -62 30289 -6
rect 30345 -62 30399 -6
rect 30455 -62 30509 -6
rect 30565 -62 30663 -6
rect 29761 -116 30663 -62
rect 29761 -172 29849 -116
rect 29905 -172 29959 -116
rect 30015 -172 30069 -116
rect 30125 -172 30179 -116
rect 30235 -172 30289 -116
rect 30345 -172 30399 -116
rect 30455 -172 30509 -116
rect 30565 -172 30663 -116
rect 28339 -745 29127 -195
rect 27246 -7741 27262 -7685
rect 27318 -7741 27372 -7685
rect 27428 -7741 27482 -7685
rect 27538 -7741 27592 -7685
rect 27648 -7741 27702 -7685
rect 27758 -7741 27775 -7685
rect 27246 -7795 27775 -7741
rect 27246 -7851 27262 -7795
rect 27318 -7851 27372 -7795
rect 27428 -7851 27482 -7795
rect 27538 -7851 27592 -7795
rect 27648 -7851 27702 -7795
rect 27758 -7851 27775 -7795
rect 27246 -7905 27775 -7851
rect 27246 -7961 27262 -7905
rect 27318 -7961 27372 -7905
rect 27428 -7961 27482 -7905
rect 27538 -7961 27592 -7905
rect 27648 -7961 27702 -7905
rect 27758 -7961 27775 -7905
rect 27246 -8015 27775 -7961
rect 27246 -8071 27262 -8015
rect 27318 -8071 27372 -8015
rect 27428 -8071 27482 -8015
rect 27538 -8071 27592 -8015
rect 27648 -8071 27702 -8015
rect 27758 -8071 27775 -8015
rect 27246 -22685 27775 -8071
rect 28340 -16521 29127 -745
rect 29761 -226 30663 -172
rect 29761 -282 29849 -226
rect 29905 -282 29959 -226
rect 30015 -282 30069 -226
rect 30125 -282 30179 -226
rect 30235 -282 30289 -226
rect 30345 -282 30399 -226
rect 30455 -282 30509 -226
rect 30565 -282 30663 -226
rect 29761 -336 30663 -282
rect 29761 -392 29849 -336
rect 29905 -392 29959 -336
rect 30015 -392 30069 -336
rect 30125 -392 30179 -336
rect 30235 -392 30289 -336
rect 30345 -392 30399 -336
rect 30455 -392 30509 -336
rect 30565 -392 30663 -336
rect 29761 -2220 30663 -392
rect 29761 -2276 29884 -2220
rect 29940 -2276 29994 -2220
rect 30050 -2276 30104 -2220
rect 30160 -2276 30214 -2220
rect 30270 -2276 30324 -2220
rect 30380 -2276 30434 -2220
rect 30490 -2276 30544 -2220
rect 30600 -2276 30663 -2220
rect 29761 -2311 30663 -2276
rect 29858 -2314 30630 -2311
rect 30146 -4151 30811 -4126
rect 30146 -4207 30166 -4151
rect 30222 -4207 30276 -4151
rect 30332 -4207 30386 -4151
rect 30442 -4207 30496 -4151
rect 30552 -4207 30606 -4151
rect 30662 -4207 30716 -4151
rect 30772 -4207 30811 -4151
rect 30146 -4261 30811 -4207
rect 30146 -4317 30166 -4261
rect 30222 -4317 30276 -4261
rect 30332 -4317 30386 -4261
rect 30442 -4317 30496 -4261
rect 30552 -4317 30606 -4261
rect 30662 -4317 30716 -4261
rect 30772 -4317 30811 -4261
rect 30146 -4376 30811 -4317
rect 30989 -4612 31776 5382
rect 69191 118 69979 121
rect 71818 118 72606 126
rect 69184 103 70023 118
rect 69184 47 69220 103
rect 69276 47 69330 103
rect 69386 47 69440 103
rect 69496 47 69550 103
rect 69606 47 69660 103
rect 69716 47 69770 103
rect 69826 47 69880 103
rect 69936 47 70023 103
rect 69184 -7 70023 47
rect 69184 -63 69220 -7
rect 69276 -63 69330 -7
rect 69386 -63 69440 -7
rect 69496 -63 69550 -7
rect 69606 -63 69660 -7
rect 69716 -63 69770 -7
rect 69826 -63 69880 -7
rect 69936 -63 70023 -7
rect 69184 -117 70023 -63
rect 69184 -173 69220 -117
rect 69276 -173 69330 -117
rect 69386 -173 69440 -117
rect 69496 -173 69550 -117
rect 69606 -173 69660 -117
rect 69716 -173 69770 -117
rect 69826 -173 69880 -117
rect 69936 -173 70023 -117
rect 69184 -227 70023 -173
rect 69184 -283 69220 -227
rect 69276 -283 69330 -227
rect 69386 -283 69440 -227
rect 69496 -283 69550 -227
rect 69606 -283 69660 -227
rect 69716 -283 69770 -227
rect 69826 -283 69880 -227
rect 69936 -283 70023 -227
rect 69184 -337 70023 -283
rect 69184 -393 69220 -337
rect 69276 -393 69330 -337
rect 69386 -393 69440 -337
rect 69496 -393 69550 -337
rect 69606 -393 69660 -337
rect 69716 -393 69770 -337
rect 69826 -393 69880 -337
rect 69936 -393 70023 -337
rect 69184 -447 70023 -393
rect 69184 -503 69220 -447
rect 69276 -503 69330 -447
rect 69386 -503 69440 -447
rect 69496 -503 69550 -447
rect 69606 -503 69660 -447
rect 69716 -503 69770 -447
rect 69826 -503 69880 -447
rect 69936 -503 70023 -447
rect 69184 -3325 70023 -503
rect 69184 -3381 69250 -3325
rect 69306 -3381 69360 -3325
rect 69416 -3381 69470 -3325
rect 69526 -3381 69580 -3325
rect 69636 -3381 69690 -3325
rect 69746 -3381 69800 -3325
rect 69856 -3381 69910 -3325
rect 69966 -3381 70023 -3325
rect 69184 -3435 70023 -3381
rect 69184 -3491 69250 -3435
rect 69306 -3491 69360 -3435
rect 69416 -3491 69470 -3435
rect 69526 -3491 69580 -3435
rect 69636 -3491 69690 -3435
rect 69746 -3491 69800 -3435
rect 69856 -3491 69910 -3435
rect 69966 -3491 70023 -3435
rect 69184 -3545 70023 -3491
rect 69184 -3601 69250 -3545
rect 69306 -3601 69360 -3545
rect 69416 -3601 69470 -3545
rect 69526 -3601 69580 -3545
rect 69636 -3601 69690 -3545
rect 69746 -3601 69800 -3545
rect 69856 -3601 69910 -3545
rect 69966 -3601 70023 -3545
rect 69184 -3655 70023 -3601
rect 69184 -3711 69250 -3655
rect 69306 -3711 69360 -3655
rect 69416 -3711 69470 -3655
rect 69526 -3711 69580 -3655
rect 69636 -3711 69690 -3655
rect 69746 -3711 69800 -3655
rect 69856 -3711 69910 -3655
rect 69966 -3711 70023 -3655
rect 69184 -3765 70023 -3711
rect 69184 -3821 69250 -3765
rect 69306 -3821 69360 -3765
rect 69416 -3821 69470 -3765
rect 69526 -3821 69580 -3765
rect 69636 -3821 69690 -3765
rect 69746 -3821 69800 -3765
rect 69856 -3821 69910 -3765
rect 69966 -3821 70023 -3765
rect 69184 -3875 70023 -3821
rect 69184 -3931 69250 -3875
rect 69306 -3931 69360 -3875
rect 69416 -3931 69470 -3875
rect 69526 -3931 69580 -3875
rect 69636 -3931 69690 -3875
rect 69746 -3931 69800 -3875
rect 69856 -3931 69910 -3875
rect 69966 -3931 70023 -3875
rect 69184 -3956 70023 -3931
rect 71812 108 72651 118
rect 71812 52 71847 108
rect 71903 52 71957 108
rect 72013 52 72067 108
rect 72123 52 72177 108
rect 72233 52 72287 108
rect 72343 52 72397 108
rect 72453 52 72507 108
rect 72563 52 72651 108
rect 74536 114 75324 132
rect 74536 88 74565 114
rect 71812 -2 72651 52
rect 71812 -58 71847 -2
rect 71903 -58 71957 -2
rect 72013 -58 72067 -2
rect 72123 -58 72177 -2
rect 72233 -58 72287 -2
rect 72343 -58 72397 -2
rect 72453 -58 72507 -2
rect 72563 -58 72651 -2
rect 71812 -112 72651 -58
rect 71812 -168 71847 -112
rect 71903 -168 71957 -112
rect 72013 -168 72067 -112
rect 72123 -168 72177 -112
rect 72233 -168 72287 -112
rect 72343 -168 72397 -112
rect 72453 -168 72507 -112
rect 72563 -168 72651 -112
rect 71812 -222 72651 -168
rect 71812 -278 71847 -222
rect 71903 -278 71957 -222
rect 72013 -278 72067 -222
rect 72123 -278 72177 -222
rect 72233 -278 72287 -222
rect 72343 -278 72397 -222
rect 72453 -278 72507 -222
rect 72563 -278 72651 -222
rect 71812 -332 72651 -278
rect 71812 -388 71847 -332
rect 71903 -388 71957 -332
rect 72013 -388 72067 -332
rect 72123 -388 72177 -332
rect 72233 -388 72287 -332
rect 72343 -388 72397 -332
rect 72453 -388 72507 -332
rect 72563 -388 72651 -332
rect 71812 -442 72651 -388
rect 71812 -498 71847 -442
rect 71903 -498 71957 -442
rect 72013 -498 72067 -442
rect 72123 -498 72177 -442
rect 72233 -498 72287 -442
rect 72343 -498 72397 -442
rect 72453 -498 72507 -442
rect 72563 -498 72651 -442
rect 71812 -3388 72651 -498
rect 71812 -3444 71863 -3388
rect 71919 -3444 71973 -3388
rect 72029 -3444 72083 -3388
rect 72139 -3444 72193 -3388
rect 72249 -3444 72303 -3388
rect 72359 -3444 72413 -3388
rect 72469 -3444 72523 -3388
rect 72579 -3444 72651 -3388
rect 71812 -3498 72651 -3444
rect 71812 -3554 71863 -3498
rect 71919 -3554 71973 -3498
rect 72029 -3554 72083 -3498
rect 72139 -3554 72193 -3498
rect 72249 -3554 72303 -3498
rect 72359 -3554 72413 -3498
rect 72469 -3554 72523 -3498
rect 72579 -3554 72651 -3498
rect 71812 -3608 72651 -3554
rect 71812 -3664 71863 -3608
rect 71919 -3664 71973 -3608
rect 72029 -3664 72083 -3608
rect 72139 -3664 72193 -3608
rect 72249 -3664 72303 -3608
rect 72359 -3664 72413 -3608
rect 72469 -3664 72523 -3608
rect 72579 -3664 72651 -3608
rect 71812 -3718 72651 -3664
rect 71812 -3774 71863 -3718
rect 71919 -3774 71973 -3718
rect 72029 -3774 72083 -3718
rect 72139 -3774 72193 -3718
rect 72249 -3774 72303 -3718
rect 72359 -3774 72413 -3718
rect 72469 -3774 72523 -3718
rect 72579 -3774 72651 -3718
rect 71812 -3828 72651 -3774
rect 71812 -3884 71863 -3828
rect 71919 -3884 71973 -3828
rect 72029 -3884 72083 -3828
rect 72139 -3884 72193 -3828
rect 72249 -3884 72303 -3828
rect 72359 -3884 72413 -3828
rect 72469 -3884 72523 -3828
rect 72579 -3884 72651 -3828
rect 71812 -3938 72651 -3884
rect 71812 -3994 71863 -3938
rect 71919 -3994 71973 -3938
rect 72029 -3994 72083 -3938
rect 72139 -3994 72193 -3938
rect 72249 -3994 72303 -3938
rect 72359 -3994 72413 -3938
rect 72469 -3994 72523 -3938
rect 72579 -3994 72651 -3938
rect 71812 -4039 72651 -3994
rect 74527 58 74565 88
rect 74621 58 74675 114
rect 74731 58 74785 114
rect 74841 58 74895 114
rect 74951 58 75005 114
rect 75061 58 75115 114
rect 75171 58 75225 114
rect 75281 88 75324 114
rect 77608 102 78396 118
rect 80658 116 81446 127
rect 80642 109 81481 116
rect 77599 100 78438 102
rect 75281 58 75366 88
rect 74527 4 75366 58
rect 74527 -52 74565 4
rect 74621 -52 74675 4
rect 74731 -52 74785 4
rect 74841 -52 74895 4
rect 74951 -52 75005 4
rect 75061 -52 75115 4
rect 75171 -52 75225 4
rect 75281 -52 75366 4
rect 74527 -106 75366 -52
rect 74527 -162 74565 -106
rect 74621 -162 74675 -106
rect 74731 -162 74785 -106
rect 74841 -162 74895 -106
rect 74951 -162 75005 -106
rect 75061 -162 75115 -106
rect 75171 -162 75225 -106
rect 75281 -162 75366 -106
rect 74527 -216 75366 -162
rect 74527 -272 74565 -216
rect 74621 -272 74675 -216
rect 74731 -272 74785 -216
rect 74841 -272 74895 -216
rect 74951 -272 75005 -216
rect 75061 -272 75115 -216
rect 75171 -272 75225 -216
rect 75281 -272 75366 -216
rect 74527 -326 75366 -272
rect 74527 -382 74565 -326
rect 74621 -382 74675 -326
rect 74731 -382 74785 -326
rect 74841 -382 74895 -326
rect 74951 -382 75005 -326
rect 75061 -382 75115 -326
rect 75171 -382 75225 -326
rect 75281 -382 75366 -326
rect 74527 -436 75366 -382
rect 74527 -492 74565 -436
rect 74621 -492 74675 -436
rect 74731 -492 74785 -436
rect 74841 -492 74895 -436
rect 74951 -492 75005 -436
rect 75061 -492 75115 -436
rect 75171 -492 75225 -436
rect 75281 -492 75366 -436
rect 74527 -3410 75366 -492
rect 74527 -3466 74577 -3410
rect 74633 -3466 74687 -3410
rect 74743 -3466 74797 -3410
rect 74853 -3466 74907 -3410
rect 74963 -3466 75017 -3410
rect 75073 -3466 75127 -3410
rect 75183 -3466 75237 -3410
rect 75293 -3466 75366 -3410
rect 74527 -3520 75366 -3466
rect 74527 -3576 74577 -3520
rect 74633 -3576 74687 -3520
rect 74743 -3576 74797 -3520
rect 74853 -3576 74907 -3520
rect 74963 -3576 75017 -3520
rect 75073 -3576 75127 -3520
rect 75183 -3576 75237 -3520
rect 75293 -3576 75366 -3520
rect 74527 -3630 75366 -3576
rect 74527 -3686 74577 -3630
rect 74633 -3686 74687 -3630
rect 74743 -3686 74797 -3630
rect 74853 -3686 74907 -3630
rect 74963 -3686 75017 -3630
rect 75073 -3686 75127 -3630
rect 75183 -3686 75237 -3630
rect 75293 -3686 75366 -3630
rect 74527 -3740 75366 -3686
rect 74527 -3796 74577 -3740
rect 74633 -3796 74687 -3740
rect 74743 -3796 74797 -3740
rect 74853 -3796 74907 -3740
rect 74963 -3796 75017 -3740
rect 75073 -3796 75127 -3740
rect 75183 -3796 75237 -3740
rect 75293 -3796 75366 -3740
rect 74527 -3850 75366 -3796
rect 74527 -3906 74577 -3850
rect 74633 -3906 74687 -3850
rect 74743 -3906 74797 -3850
rect 74853 -3906 74907 -3850
rect 74963 -3906 75017 -3850
rect 75073 -3906 75127 -3850
rect 75183 -3906 75237 -3850
rect 75293 -3906 75366 -3850
rect 74527 -3960 75366 -3906
rect 74527 -4016 74577 -3960
rect 74633 -4016 74687 -3960
rect 74743 -4016 74797 -3960
rect 74853 -4016 74907 -3960
rect 74963 -4016 75017 -3960
rect 75073 -4016 75127 -3960
rect 75183 -4016 75237 -3960
rect 75293 -4016 75366 -3960
rect 74527 -4057 75366 -4016
rect 77599 44 77637 100
rect 77693 44 77747 100
rect 77803 44 77857 100
rect 77913 44 77967 100
rect 78023 44 78077 100
rect 78133 44 78187 100
rect 78243 44 78297 100
rect 78353 44 78438 100
rect 77599 -10 78438 44
rect 77599 -66 77637 -10
rect 77693 -66 77747 -10
rect 77803 -66 77857 -10
rect 77913 -66 77967 -10
rect 78023 -66 78077 -10
rect 78133 -66 78187 -10
rect 78243 -66 78297 -10
rect 78353 -66 78438 -10
rect 77599 -120 78438 -66
rect 77599 -176 77637 -120
rect 77693 -176 77747 -120
rect 77803 -176 77857 -120
rect 77913 -176 77967 -120
rect 78023 -176 78077 -120
rect 78133 -176 78187 -120
rect 78243 -176 78297 -120
rect 78353 -176 78438 -120
rect 77599 -230 78438 -176
rect 77599 -286 77637 -230
rect 77693 -286 77747 -230
rect 77803 -286 77857 -230
rect 77913 -286 77967 -230
rect 78023 -286 78077 -230
rect 78133 -286 78187 -230
rect 78243 -286 78297 -230
rect 78353 -286 78438 -230
rect 77599 -340 78438 -286
rect 77599 -396 77637 -340
rect 77693 -396 77747 -340
rect 77803 -396 77857 -340
rect 77913 -396 77967 -340
rect 78023 -396 78077 -340
rect 78133 -396 78187 -340
rect 78243 -396 78297 -340
rect 78353 -396 78438 -340
rect 77599 -450 78438 -396
rect 77599 -506 77637 -450
rect 77693 -506 77747 -450
rect 77803 -506 77857 -450
rect 77913 -506 77967 -450
rect 78023 -506 78077 -450
rect 78133 -506 78187 -450
rect 78243 -506 78297 -450
rect 78353 -506 78438 -450
rect 77599 -3384 78438 -506
rect 77599 -3440 77645 -3384
rect 77701 -3440 77755 -3384
rect 77811 -3440 77865 -3384
rect 77921 -3440 77975 -3384
rect 78031 -3440 78085 -3384
rect 78141 -3440 78195 -3384
rect 78251 -3440 78305 -3384
rect 78361 -3440 78438 -3384
rect 77599 -3494 78438 -3440
rect 77599 -3550 77645 -3494
rect 77701 -3550 77755 -3494
rect 77811 -3550 77865 -3494
rect 77921 -3550 77975 -3494
rect 78031 -3550 78085 -3494
rect 78141 -3550 78195 -3494
rect 78251 -3550 78305 -3494
rect 78361 -3550 78438 -3494
rect 77599 -3604 78438 -3550
rect 77599 -3660 77645 -3604
rect 77701 -3660 77755 -3604
rect 77811 -3660 77865 -3604
rect 77921 -3660 77975 -3604
rect 78031 -3660 78085 -3604
rect 78141 -3660 78195 -3604
rect 78251 -3660 78305 -3604
rect 78361 -3660 78438 -3604
rect 77599 -3714 78438 -3660
rect 77599 -3770 77645 -3714
rect 77701 -3770 77755 -3714
rect 77811 -3770 77865 -3714
rect 77921 -3770 77975 -3714
rect 78031 -3770 78085 -3714
rect 78141 -3770 78195 -3714
rect 78251 -3770 78305 -3714
rect 78361 -3770 78438 -3714
rect 77599 -3824 78438 -3770
rect 77599 -3880 77645 -3824
rect 77701 -3880 77755 -3824
rect 77811 -3880 77865 -3824
rect 77921 -3880 77975 -3824
rect 78031 -3880 78085 -3824
rect 78141 -3880 78195 -3824
rect 78251 -3880 78305 -3824
rect 78361 -3880 78438 -3824
rect 77599 -3934 78438 -3880
rect 77599 -3990 77645 -3934
rect 77701 -3990 77755 -3934
rect 77811 -3990 77865 -3934
rect 77921 -3990 77975 -3934
rect 78031 -3990 78085 -3934
rect 78141 -3990 78195 -3934
rect 78251 -3990 78305 -3934
rect 78361 -3990 78438 -3934
rect 77599 -4021 78438 -3990
rect 80642 53 80687 109
rect 80743 53 80797 109
rect 80853 53 80907 109
rect 80963 53 81017 109
rect 81073 53 81127 109
rect 81183 53 81237 109
rect 81293 53 81347 109
rect 81403 53 81481 109
rect 83499 109 84287 127
rect 83499 102 83528 109
rect 80642 -1 81481 53
rect 80642 -57 80687 -1
rect 80743 -57 80797 -1
rect 80853 -57 80907 -1
rect 80963 -57 81017 -1
rect 81073 -57 81127 -1
rect 81183 -57 81237 -1
rect 81293 -57 81347 -1
rect 81403 -57 81481 -1
rect 80642 -111 81481 -57
rect 80642 -167 80687 -111
rect 80743 -167 80797 -111
rect 80853 -167 80907 -111
rect 80963 -167 81017 -111
rect 81073 -167 81127 -111
rect 81183 -167 81237 -111
rect 81293 -167 81347 -111
rect 81403 -167 81481 -111
rect 80642 -221 81481 -167
rect 80642 -277 80687 -221
rect 80743 -277 80797 -221
rect 80853 -277 80907 -221
rect 80963 -277 81017 -221
rect 81073 -277 81127 -221
rect 81183 -277 81237 -221
rect 81293 -277 81347 -221
rect 81403 -277 81481 -221
rect 80642 -331 81481 -277
rect 80642 -387 80687 -331
rect 80743 -387 80797 -331
rect 80853 -387 80907 -331
rect 80963 -387 81017 -331
rect 81073 -387 81127 -331
rect 81183 -387 81237 -331
rect 81293 -387 81347 -331
rect 81403 -387 81481 -331
rect 80642 -441 81481 -387
rect 80642 -497 80687 -441
rect 80743 -497 80797 -441
rect 80853 -497 80907 -441
rect 80963 -497 81017 -441
rect 81073 -497 81127 -441
rect 81183 -497 81237 -441
rect 81293 -497 81347 -441
rect 81403 -497 81481 -441
rect 80642 -3356 81481 -497
rect 80642 -3412 80699 -3356
rect 80755 -3412 80809 -3356
rect 80865 -3412 80919 -3356
rect 80975 -3412 81029 -3356
rect 81085 -3412 81139 -3356
rect 81195 -3412 81249 -3356
rect 81305 -3412 81359 -3356
rect 81415 -3412 81481 -3356
rect 80642 -3466 81481 -3412
rect 80642 -3522 80699 -3466
rect 80755 -3522 80809 -3466
rect 80865 -3522 80919 -3466
rect 80975 -3522 81029 -3466
rect 81085 -3522 81139 -3466
rect 81195 -3522 81249 -3466
rect 81305 -3522 81359 -3466
rect 81415 -3522 81481 -3466
rect 80642 -3576 81481 -3522
rect 80642 -3632 80699 -3576
rect 80755 -3632 80809 -3576
rect 80865 -3632 80919 -3576
rect 80975 -3632 81029 -3576
rect 81085 -3632 81139 -3576
rect 81195 -3632 81249 -3576
rect 81305 -3632 81359 -3576
rect 81415 -3632 81481 -3576
rect 80642 -3686 81481 -3632
rect 80642 -3742 80699 -3686
rect 80755 -3742 80809 -3686
rect 80865 -3742 80919 -3686
rect 80975 -3742 81029 -3686
rect 81085 -3742 81139 -3686
rect 81195 -3742 81249 -3686
rect 81305 -3742 81359 -3686
rect 81415 -3742 81481 -3686
rect 80642 -3796 81481 -3742
rect 80642 -3852 80699 -3796
rect 80755 -3852 80809 -3796
rect 80865 -3852 80919 -3796
rect 80975 -3852 81029 -3796
rect 81085 -3852 81139 -3796
rect 81195 -3852 81249 -3796
rect 81305 -3852 81359 -3796
rect 81415 -3852 81481 -3796
rect 80642 -3906 81481 -3852
rect 80642 -3962 80699 -3906
rect 80755 -3962 80809 -3906
rect 80865 -3962 80919 -3906
rect 80975 -3962 81029 -3906
rect 81085 -3962 81139 -3906
rect 81195 -3962 81249 -3906
rect 81305 -3962 81359 -3906
rect 81415 -3962 81481 -3906
rect 80642 -3993 81481 -3962
rect 83489 53 83528 102
rect 83584 53 83638 109
rect 83694 53 83748 109
rect 83804 53 83858 109
rect 83914 53 83968 109
rect 84024 53 84078 109
rect 84134 53 84188 109
rect 84244 102 84287 109
rect 86280 106 87119 130
rect 84244 53 84328 102
rect 83489 -1 84328 53
rect 83489 -57 83528 -1
rect 83584 -57 83638 -1
rect 83694 -57 83748 -1
rect 83804 -57 83858 -1
rect 83914 -57 83968 -1
rect 84024 -57 84078 -1
rect 84134 -57 84188 -1
rect 84244 -57 84328 -1
rect 83489 -111 84328 -57
rect 83489 -167 83528 -111
rect 83584 -167 83638 -111
rect 83694 -167 83748 -111
rect 83804 -167 83858 -111
rect 83914 -167 83968 -111
rect 84024 -167 84078 -111
rect 84134 -167 84188 -111
rect 84244 -167 84328 -111
rect 83489 -221 84328 -167
rect 83489 -277 83528 -221
rect 83584 -277 83638 -221
rect 83694 -277 83748 -221
rect 83804 -277 83858 -221
rect 83914 -277 83968 -221
rect 84024 -277 84078 -221
rect 84134 -277 84188 -221
rect 84244 -277 84328 -221
rect 83489 -331 84328 -277
rect 83489 -387 83528 -331
rect 83584 -387 83638 -331
rect 83694 -387 83748 -331
rect 83804 -387 83858 -331
rect 83914 -387 83968 -331
rect 84024 -387 84078 -331
rect 84134 -387 84188 -331
rect 84244 -387 84328 -331
rect 83489 -441 84328 -387
rect 83489 -497 83528 -441
rect 83584 -497 83638 -441
rect 83694 -497 83748 -441
rect 83804 -497 83858 -441
rect 83914 -497 83968 -441
rect 84024 -497 84078 -441
rect 84134 -497 84188 -441
rect 84244 -497 84328 -441
rect 83489 -3352 84328 -497
rect 83489 -3408 83552 -3352
rect 83608 -3408 83662 -3352
rect 83718 -3408 83772 -3352
rect 83828 -3408 83882 -3352
rect 83938 -3408 83992 -3352
rect 84048 -3408 84102 -3352
rect 84158 -3408 84212 -3352
rect 84268 -3408 84328 -3352
rect 83489 -3462 84328 -3408
rect 83489 -3518 83552 -3462
rect 83608 -3518 83662 -3462
rect 83718 -3518 83772 -3462
rect 83828 -3518 83882 -3462
rect 83938 -3518 83992 -3462
rect 84048 -3518 84102 -3462
rect 84158 -3518 84212 -3462
rect 84268 -3518 84328 -3462
rect 83489 -3572 84328 -3518
rect 83489 -3628 83552 -3572
rect 83608 -3628 83662 -3572
rect 83718 -3628 83772 -3572
rect 83828 -3628 83882 -3572
rect 83938 -3628 83992 -3572
rect 84048 -3628 84102 -3572
rect 84158 -3628 84212 -3572
rect 84268 -3628 84328 -3572
rect 83489 -3682 84328 -3628
rect 83489 -3738 83552 -3682
rect 83608 -3738 83662 -3682
rect 83718 -3738 83772 -3682
rect 83828 -3738 83882 -3682
rect 83938 -3738 83992 -3682
rect 84048 -3738 84102 -3682
rect 84158 -3738 84212 -3682
rect 84268 -3738 84328 -3682
rect 83489 -3792 84328 -3738
rect 83489 -3848 83552 -3792
rect 83608 -3848 83662 -3792
rect 83718 -3848 83772 -3792
rect 83828 -3848 83882 -3792
rect 83938 -3848 83992 -3792
rect 84048 -3848 84102 -3792
rect 84158 -3848 84212 -3792
rect 84268 -3848 84328 -3792
rect 83489 -3902 84328 -3848
rect 83489 -3958 83552 -3902
rect 83608 -3958 83662 -3902
rect 83718 -3958 83772 -3902
rect 83828 -3958 83882 -3902
rect 83938 -3958 83992 -3902
rect 84048 -3958 84102 -3902
rect 84158 -3958 84212 -3902
rect 84268 -3958 84328 -3902
rect 83489 -3993 84328 -3958
rect 86280 50 86316 106
rect 86372 50 86426 106
rect 86482 50 86536 106
rect 86592 50 86646 106
rect 86702 50 86756 106
rect 86812 50 86866 106
rect 86922 50 86976 106
rect 87032 50 87119 106
rect 86280 -4 87119 50
rect 86280 -60 86316 -4
rect 86372 -60 86426 -4
rect 86482 -60 86536 -4
rect 86592 -60 86646 -4
rect 86702 -60 86756 -4
rect 86812 -60 86866 -4
rect 86922 -60 86976 -4
rect 87032 -60 87119 -4
rect 86280 -114 87119 -60
rect 86280 -170 86316 -114
rect 86372 -170 86426 -114
rect 86482 -170 86536 -114
rect 86592 -170 86646 -114
rect 86702 -170 86756 -114
rect 86812 -170 86866 -114
rect 86922 -170 86976 -114
rect 87032 -170 87119 -114
rect 86280 -224 87119 -170
rect 86280 -280 86316 -224
rect 86372 -280 86426 -224
rect 86482 -280 86536 -224
rect 86592 -280 86646 -224
rect 86702 -280 86756 -224
rect 86812 -280 86866 -224
rect 86922 -280 86976 -224
rect 87032 -280 87119 -224
rect 86280 -334 87119 -280
rect 86280 -390 86316 -334
rect 86372 -390 86426 -334
rect 86482 -390 86536 -334
rect 86592 -390 86646 -334
rect 86702 -390 86756 -334
rect 86812 -390 86866 -334
rect 86922 -390 86976 -334
rect 87032 -390 87119 -334
rect 86280 -444 87119 -390
rect 86280 -500 86316 -444
rect 86372 -500 86426 -444
rect 86482 -500 86536 -444
rect 86592 -500 86646 -444
rect 86702 -500 86756 -444
rect 86812 -500 86866 -444
rect 86922 -500 86976 -444
rect 87032 -500 87119 -444
rect 86280 -3376 87119 -500
rect 86280 -3432 86339 -3376
rect 86395 -3432 86449 -3376
rect 86505 -3432 86559 -3376
rect 86615 -3432 86669 -3376
rect 86725 -3432 86779 -3376
rect 86835 -3432 86889 -3376
rect 86945 -3432 86999 -3376
rect 87055 -3432 87119 -3376
rect 86280 -3486 87119 -3432
rect 86280 -3542 86339 -3486
rect 86395 -3542 86449 -3486
rect 86505 -3542 86559 -3486
rect 86615 -3542 86669 -3486
rect 86725 -3542 86779 -3486
rect 86835 -3542 86889 -3486
rect 86945 -3542 86999 -3486
rect 87055 -3542 87119 -3486
rect 86280 -3596 87119 -3542
rect 86280 -3652 86339 -3596
rect 86395 -3652 86449 -3596
rect 86505 -3652 86559 -3596
rect 86615 -3652 86669 -3596
rect 86725 -3652 86779 -3596
rect 86835 -3652 86889 -3596
rect 86945 -3652 86999 -3596
rect 87055 -3652 87119 -3596
rect 86280 -3706 87119 -3652
rect 86280 -3762 86339 -3706
rect 86395 -3762 86449 -3706
rect 86505 -3762 86559 -3706
rect 86615 -3762 86669 -3706
rect 86725 -3762 86779 -3706
rect 86835 -3762 86889 -3706
rect 86945 -3762 86999 -3706
rect 87055 -3762 87119 -3706
rect 86280 -3816 87119 -3762
rect 86280 -3872 86339 -3816
rect 86395 -3872 86449 -3816
rect 86505 -3872 86559 -3816
rect 86615 -3872 86669 -3816
rect 86725 -3872 86779 -3816
rect 86835 -3872 86889 -3816
rect 86945 -3872 86999 -3816
rect 87055 -3872 87119 -3816
rect 86280 -3926 87119 -3872
rect 86280 -3982 86339 -3926
rect 86395 -3982 86449 -3926
rect 86505 -3982 86559 -3926
rect 86615 -3982 86669 -3926
rect 86725 -3982 86779 -3926
rect 86835 -3982 86889 -3926
rect 86945 -3982 86999 -3926
rect 87055 -3982 87119 -3926
rect 89463 118 90302 186
rect 89463 62 89511 118
rect 89567 62 89621 118
rect 89677 62 89731 118
rect 89787 62 89841 118
rect 89897 62 89951 118
rect 90007 62 90061 118
rect 90117 62 90171 118
rect 90227 62 90302 118
rect 89463 8 90302 62
rect 89463 -48 89511 8
rect 89567 -48 89621 8
rect 89677 -48 89731 8
rect 89787 -48 89841 8
rect 89897 -48 89951 8
rect 90007 -48 90061 8
rect 90117 -48 90171 8
rect 90227 -48 90302 8
rect 89463 -102 90302 -48
rect 89463 -158 89511 -102
rect 89567 -158 89621 -102
rect 89677 -158 89731 -102
rect 89787 -158 89841 -102
rect 89897 -158 89951 -102
rect 90007 -158 90061 -102
rect 90117 -158 90171 -102
rect 90227 -158 90302 -102
rect 89463 -212 90302 -158
rect 89463 -268 89511 -212
rect 89567 -268 89621 -212
rect 89677 -268 89731 -212
rect 89787 -268 89841 -212
rect 89897 -268 89951 -212
rect 90007 -268 90061 -212
rect 90117 -268 90171 -212
rect 90227 -268 90302 -212
rect 89463 -322 90302 -268
rect 89463 -378 89511 -322
rect 89567 -378 89621 -322
rect 89677 -378 89731 -322
rect 89787 -378 89841 -322
rect 89897 -378 89951 -322
rect 90007 -378 90061 -322
rect 90117 -378 90171 -322
rect 90227 -378 90302 -322
rect 89463 -432 90302 -378
rect 89463 -488 89511 -432
rect 89567 -488 89621 -432
rect 89677 -488 89731 -432
rect 89787 -488 89841 -432
rect 89897 -488 89951 -432
rect 90007 -488 90061 -432
rect 90117 -488 90171 -432
rect 90227 -488 90302 -432
rect 89463 -3329 90302 -488
rect 89463 -3385 89521 -3329
rect 89577 -3385 89631 -3329
rect 89687 -3385 89741 -3329
rect 89797 -3385 89851 -3329
rect 89907 -3385 89961 -3329
rect 90017 -3385 90071 -3329
rect 90127 -3385 90181 -3329
rect 90237 -3385 90302 -3329
rect 89463 -3439 90302 -3385
rect 89463 -3495 89521 -3439
rect 89577 -3495 89631 -3439
rect 89687 -3495 89741 -3439
rect 89797 -3495 89851 -3439
rect 89907 -3495 89961 -3439
rect 90017 -3495 90071 -3439
rect 90127 -3495 90181 -3439
rect 90237 -3495 90302 -3439
rect 89463 -3549 90302 -3495
rect 89463 -3605 89521 -3549
rect 89577 -3605 89631 -3549
rect 89687 -3605 89741 -3549
rect 89797 -3605 89851 -3549
rect 89907 -3605 89961 -3549
rect 90017 -3605 90071 -3549
rect 90127 -3605 90181 -3549
rect 90237 -3605 90302 -3549
rect 89463 -3659 90302 -3605
rect 89463 -3715 89521 -3659
rect 89577 -3715 89631 -3659
rect 89687 -3715 89741 -3659
rect 89797 -3715 89851 -3659
rect 89907 -3715 89961 -3659
rect 90017 -3715 90071 -3659
rect 90127 -3715 90181 -3659
rect 90237 -3715 90302 -3659
rect 89463 -3769 90302 -3715
rect 89463 -3825 89521 -3769
rect 89577 -3825 89631 -3769
rect 89687 -3825 89741 -3769
rect 89797 -3825 89851 -3769
rect 89907 -3825 89961 -3769
rect 90017 -3825 90071 -3769
rect 90127 -3825 90181 -3769
rect 90237 -3825 90302 -3769
rect 89463 -3879 90302 -3825
rect 89463 -3935 89521 -3879
rect 89577 -3935 89631 -3879
rect 89687 -3935 89741 -3879
rect 89797 -3935 89851 -3879
rect 89907 -3935 89961 -3879
rect 90017 -3935 90071 -3879
rect 90127 -3935 90181 -3879
rect 90237 -3935 90302 -3879
rect 89463 -3975 90302 -3935
rect 92815 107 93654 130
rect 92815 51 92852 107
rect 92908 51 92962 107
rect 93018 51 93072 107
rect 93128 51 93182 107
rect 93238 51 93292 107
rect 93348 51 93402 107
rect 93458 51 93512 107
rect 93568 51 93654 107
rect 92815 -3 93654 51
rect 92815 -59 92852 -3
rect 92908 -59 92962 -3
rect 93018 -59 93072 -3
rect 93128 -59 93182 -3
rect 93238 -59 93292 -3
rect 93348 -59 93402 -3
rect 93458 -59 93512 -3
rect 93568 -59 93654 -3
rect 92815 -113 93654 -59
rect 92815 -169 92852 -113
rect 92908 -169 92962 -113
rect 93018 -169 93072 -113
rect 93128 -169 93182 -113
rect 93238 -169 93292 -113
rect 93348 -169 93402 -113
rect 93458 -169 93512 -113
rect 93568 -169 93654 -113
rect 92815 -223 93654 -169
rect 92815 -279 92852 -223
rect 92908 -279 92962 -223
rect 93018 -279 93072 -223
rect 93128 -279 93182 -223
rect 93238 -279 93292 -223
rect 93348 -279 93402 -223
rect 93458 -279 93512 -223
rect 93568 -279 93654 -223
rect 92815 -333 93654 -279
rect 92815 -389 92852 -333
rect 92908 -389 92962 -333
rect 93018 -389 93072 -333
rect 93128 -389 93182 -333
rect 93238 -389 93292 -333
rect 93348 -389 93402 -333
rect 93458 -389 93512 -333
rect 93568 -389 93654 -333
rect 92815 -443 93654 -389
rect 92815 -499 92852 -443
rect 92908 -499 92962 -443
rect 93018 -499 93072 -443
rect 93128 -499 93182 -443
rect 93238 -499 93292 -443
rect 93348 -499 93402 -443
rect 93458 -499 93512 -443
rect 93568 -499 93654 -443
rect 92815 -3354 93654 -499
rect 92815 -3410 92865 -3354
rect 92921 -3410 92975 -3354
rect 93031 -3410 93085 -3354
rect 93141 -3410 93195 -3354
rect 93251 -3410 93305 -3354
rect 93361 -3410 93415 -3354
rect 93471 -3410 93525 -3354
rect 93581 -3410 93654 -3354
rect 92815 -3464 93654 -3410
rect 92815 -3520 92865 -3464
rect 92921 -3520 92975 -3464
rect 93031 -3520 93085 -3464
rect 93141 -3520 93195 -3464
rect 93251 -3520 93305 -3464
rect 93361 -3520 93415 -3464
rect 93471 -3520 93525 -3464
rect 93581 -3520 93654 -3464
rect 92815 -3574 93654 -3520
rect 92815 -3630 92865 -3574
rect 92921 -3630 92975 -3574
rect 93031 -3630 93085 -3574
rect 93141 -3630 93195 -3574
rect 93251 -3630 93305 -3574
rect 93361 -3630 93415 -3574
rect 93471 -3630 93525 -3574
rect 93581 -3630 93654 -3574
rect 92815 -3684 93654 -3630
rect 92815 -3740 92865 -3684
rect 92921 -3740 92975 -3684
rect 93031 -3740 93085 -3684
rect 93141 -3740 93195 -3684
rect 93251 -3740 93305 -3684
rect 93361 -3740 93415 -3684
rect 93471 -3740 93525 -3684
rect 93581 -3740 93654 -3684
rect 92815 -3794 93654 -3740
rect 92815 -3850 92865 -3794
rect 92921 -3850 92975 -3794
rect 93031 -3850 93085 -3794
rect 93141 -3850 93195 -3794
rect 93251 -3850 93305 -3794
rect 93361 -3850 93415 -3794
rect 93471 -3850 93525 -3794
rect 93581 -3850 93654 -3794
rect 92815 -3904 93654 -3850
rect 92815 -3960 92865 -3904
rect 92921 -3960 92975 -3904
rect 93031 -3960 93085 -3904
rect 93141 -3960 93195 -3904
rect 93251 -3960 93305 -3904
rect 93361 -3960 93415 -3904
rect 93471 -3960 93525 -3904
rect 93581 -3960 93654 -3904
rect 86280 -4002 87119 -3982
rect 92815 -4011 93654 -3960
rect 95956 110 96795 144
rect 95956 54 95994 110
rect 96050 54 96104 110
rect 96160 54 96214 110
rect 96270 54 96324 110
rect 96380 54 96434 110
rect 96490 54 96544 110
rect 96600 54 96654 110
rect 96710 54 96795 110
rect 95956 0 96795 54
rect 95956 -56 95994 0
rect 96050 -56 96104 0
rect 96160 -56 96214 0
rect 96270 -56 96324 0
rect 96380 -56 96434 0
rect 96490 -56 96544 0
rect 96600 -56 96654 0
rect 96710 -56 96795 0
rect 95956 -110 96795 -56
rect 95956 -166 95994 -110
rect 96050 -166 96104 -110
rect 96160 -166 96214 -110
rect 96270 -166 96324 -110
rect 96380 -166 96434 -110
rect 96490 -166 96544 -110
rect 96600 -166 96654 -110
rect 96710 -166 96795 -110
rect 95956 -220 96795 -166
rect 95956 -276 95994 -220
rect 96050 -276 96104 -220
rect 96160 -276 96214 -220
rect 96270 -276 96324 -220
rect 96380 -276 96434 -220
rect 96490 -276 96544 -220
rect 96600 -276 96654 -220
rect 96710 -276 96795 -220
rect 95956 -330 96795 -276
rect 95956 -386 95994 -330
rect 96050 -386 96104 -330
rect 96160 -386 96214 -330
rect 96270 -386 96324 -330
rect 96380 -386 96434 -330
rect 96490 -386 96544 -330
rect 96600 -386 96654 -330
rect 96710 -386 96795 -330
rect 95956 -440 96795 -386
rect 95956 -496 95994 -440
rect 96050 -496 96104 -440
rect 96160 -496 96214 -440
rect 96270 -496 96324 -440
rect 96380 -496 96434 -440
rect 96490 -496 96544 -440
rect 96600 -496 96654 -440
rect 96710 -496 96795 -440
rect 95956 -3384 96795 -496
rect 95956 -3440 95998 -3384
rect 96054 -3440 96108 -3384
rect 96164 -3440 96218 -3384
rect 96274 -3440 96328 -3384
rect 96384 -3440 96438 -3384
rect 96494 -3440 96548 -3384
rect 96604 -3440 96658 -3384
rect 96714 -3440 96795 -3384
rect 95956 -3494 96795 -3440
rect 95956 -3550 95998 -3494
rect 96054 -3550 96108 -3494
rect 96164 -3550 96218 -3494
rect 96274 -3550 96328 -3494
rect 96384 -3550 96438 -3494
rect 96494 -3550 96548 -3494
rect 96604 -3550 96658 -3494
rect 96714 -3550 96795 -3494
rect 95956 -3604 96795 -3550
rect 95956 -3660 95998 -3604
rect 96054 -3660 96108 -3604
rect 96164 -3660 96218 -3604
rect 96274 -3660 96328 -3604
rect 96384 -3660 96438 -3604
rect 96494 -3660 96548 -3604
rect 96604 -3660 96658 -3604
rect 96714 -3660 96795 -3604
rect 95956 -3714 96795 -3660
rect 95956 -3770 95998 -3714
rect 96054 -3770 96108 -3714
rect 96164 -3770 96218 -3714
rect 96274 -3770 96328 -3714
rect 96384 -3770 96438 -3714
rect 96494 -3770 96548 -3714
rect 96604 -3770 96658 -3714
rect 96714 -3770 96795 -3714
rect 95956 -3824 96795 -3770
rect 95956 -3880 95998 -3824
rect 96054 -3880 96108 -3824
rect 96164 -3880 96218 -3824
rect 96274 -3880 96328 -3824
rect 96384 -3880 96438 -3824
rect 96494 -3880 96548 -3824
rect 96604 -3880 96658 -3824
rect 96714 -3880 96795 -3824
rect 95956 -3934 96795 -3880
rect 95956 -3990 95998 -3934
rect 96054 -3990 96108 -3934
rect 96164 -3990 96218 -3934
rect 96274 -3990 96328 -3934
rect 96384 -3990 96438 -3934
rect 96494 -3990 96548 -3934
rect 96604 -3990 96658 -3934
rect 96714 -3990 96795 -3934
rect 95956 -4039 96795 -3990
rect 99238 108 100077 144
rect 99238 52 99280 108
rect 99336 52 99390 108
rect 99446 52 99500 108
rect 99556 52 99610 108
rect 99666 52 99720 108
rect 99776 52 99830 108
rect 99886 52 99940 108
rect 99996 52 100077 108
rect 99238 -2 100077 52
rect 99238 -58 99280 -2
rect 99336 -58 99390 -2
rect 99446 -58 99500 -2
rect 99556 -58 99610 -2
rect 99666 -58 99720 -2
rect 99776 -58 99830 -2
rect 99886 -58 99940 -2
rect 99996 -58 100077 -2
rect 99238 -112 100077 -58
rect 99238 -168 99280 -112
rect 99336 -168 99390 -112
rect 99446 -168 99500 -112
rect 99556 -168 99610 -112
rect 99666 -168 99720 -112
rect 99776 -168 99830 -112
rect 99886 -168 99940 -112
rect 99996 -168 100077 -112
rect 99238 -222 100077 -168
rect 99238 -278 99280 -222
rect 99336 -278 99390 -222
rect 99446 -278 99500 -222
rect 99556 -278 99610 -222
rect 99666 -278 99720 -222
rect 99776 -278 99830 -222
rect 99886 -278 99940 -222
rect 99996 -278 100077 -222
rect 99238 -332 100077 -278
rect 99238 -388 99280 -332
rect 99336 -388 99390 -332
rect 99446 -388 99500 -332
rect 99556 -388 99610 -332
rect 99666 -388 99720 -332
rect 99776 -388 99830 -332
rect 99886 -388 99940 -332
rect 99996 -388 100077 -332
rect 99238 -442 100077 -388
rect 99238 -498 99280 -442
rect 99336 -498 99390 -442
rect 99446 -498 99500 -442
rect 99556 -498 99610 -442
rect 99666 -498 99720 -442
rect 99776 -498 99830 -442
rect 99886 -498 99940 -442
rect 99996 -498 100077 -442
rect 99238 -3418 100077 -498
rect 99238 -3474 99276 -3418
rect 99332 -3474 99386 -3418
rect 99442 -3474 99496 -3418
rect 99552 -3474 99606 -3418
rect 99662 -3474 99716 -3418
rect 99772 -3474 99826 -3418
rect 99882 -3474 99936 -3418
rect 99992 -3474 100077 -3418
rect 99238 -3528 100077 -3474
rect 99238 -3584 99276 -3528
rect 99332 -3584 99386 -3528
rect 99442 -3584 99496 -3528
rect 99552 -3584 99606 -3528
rect 99662 -3584 99716 -3528
rect 99772 -3584 99826 -3528
rect 99882 -3584 99936 -3528
rect 99992 -3584 100077 -3528
rect 99238 -3638 100077 -3584
rect 99238 -3694 99276 -3638
rect 99332 -3694 99386 -3638
rect 99442 -3694 99496 -3638
rect 99552 -3694 99606 -3638
rect 99662 -3694 99716 -3638
rect 99772 -3694 99826 -3638
rect 99882 -3694 99936 -3638
rect 99992 -3694 100077 -3638
rect 99238 -3748 100077 -3694
rect 99238 -3804 99276 -3748
rect 99332 -3804 99386 -3748
rect 99442 -3804 99496 -3748
rect 99552 -3804 99606 -3748
rect 99662 -3804 99716 -3748
rect 99772 -3804 99826 -3748
rect 99882 -3804 99936 -3748
rect 99992 -3804 100077 -3748
rect 99238 -3858 100077 -3804
rect 99238 -3914 99276 -3858
rect 99332 -3914 99386 -3858
rect 99442 -3914 99496 -3858
rect 99552 -3914 99606 -3858
rect 99662 -3914 99716 -3858
rect 99772 -3914 99826 -3858
rect 99882 -3914 99936 -3858
rect 99992 -3914 100077 -3858
rect 99238 -3968 100077 -3914
rect 99238 -4024 99276 -3968
rect 99332 -4024 99386 -3968
rect 99442 -4024 99496 -3968
rect 99552 -4024 99606 -3968
rect 99662 -4024 99716 -3968
rect 99772 -4024 99826 -3968
rect 99882 -4024 99936 -3968
rect 99992 -4024 100077 -3968
rect 99238 -4057 100077 -4024
rect 107175 -2423 107963 5958
rect 110597 1746 111385 1796
rect 110597 1723 110643 1746
rect 110594 1690 110643 1723
rect 110699 1690 110753 1746
rect 110809 1690 110863 1746
rect 110919 1690 110973 1746
rect 111029 1690 111083 1746
rect 111139 1690 111193 1746
rect 111249 1690 111303 1746
rect 111359 1723 111385 1746
rect 111359 1690 111580 1723
rect 110594 1636 111580 1690
rect 110594 1580 110643 1636
rect 110699 1580 110753 1636
rect 110809 1580 110863 1636
rect 110919 1580 110973 1636
rect 111029 1580 111083 1636
rect 111139 1580 111193 1636
rect 111249 1580 111303 1636
rect 111359 1580 111580 1636
rect 110594 1526 111580 1580
rect 110594 1470 110643 1526
rect 110699 1470 110753 1526
rect 110809 1470 110863 1526
rect 110919 1470 110973 1526
rect 111029 1470 111083 1526
rect 111139 1470 111193 1526
rect 111249 1470 111303 1526
rect 111359 1470 111580 1526
rect 110594 1416 111580 1470
rect 110594 1360 110643 1416
rect 110699 1360 110753 1416
rect 110809 1360 110863 1416
rect 110919 1360 110973 1416
rect 111029 1360 111083 1416
rect 111139 1360 111193 1416
rect 111249 1360 111303 1416
rect 111359 1360 111580 1416
rect 110594 1306 111580 1360
rect 110594 1250 110643 1306
rect 110699 1250 110753 1306
rect 110809 1250 110863 1306
rect 110919 1250 110973 1306
rect 111029 1250 111083 1306
rect 111139 1250 111193 1306
rect 111249 1250 111303 1306
rect 111359 1250 111580 1306
rect 110594 1196 111580 1250
rect 110594 1140 110643 1196
rect 110699 1140 110753 1196
rect 110809 1140 110863 1196
rect 110919 1140 110973 1196
rect 111029 1140 111083 1196
rect 111139 1140 111193 1196
rect 111249 1140 111303 1196
rect 111359 1140 111580 1196
rect 110594 1086 111580 1140
rect 110594 1030 110643 1086
rect 110699 1030 110753 1086
rect 110809 1030 110863 1086
rect 110919 1030 110973 1086
rect 111029 1030 111083 1086
rect 111139 1030 111193 1086
rect 111249 1030 111303 1086
rect 111359 1030 111580 1086
rect 107175 -2479 107221 -2423
rect 107277 -2479 107331 -2423
rect 107387 -2479 107441 -2423
rect 107497 -2479 107551 -2423
rect 107607 -2479 107661 -2423
rect 107717 -2479 107771 -2423
rect 107827 -2479 107881 -2423
rect 107937 -2479 107963 -2423
rect 107175 -2533 107963 -2479
rect 107175 -2589 107221 -2533
rect 107277 -2589 107331 -2533
rect 107387 -2589 107441 -2533
rect 107497 -2589 107551 -2533
rect 107607 -2589 107661 -2533
rect 107717 -2589 107771 -2533
rect 107827 -2589 107881 -2533
rect 107937 -2589 107963 -2533
rect 107175 -2643 107963 -2589
rect 107175 -2699 107221 -2643
rect 107277 -2699 107331 -2643
rect 107387 -2699 107441 -2643
rect 107497 -2699 107551 -2643
rect 107607 -2699 107661 -2643
rect 107717 -2699 107771 -2643
rect 107827 -2699 107881 -2643
rect 107937 -2699 107963 -2643
rect 107175 -2753 107963 -2699
rect 107175 -2809 107221 -2753
rect 107277 -2809 107331 -2753
rect 107387 -2809 107441 -2753
rect 107497 -2809 107551 -2753
rect 107607 -2809 107661 -2753
rect 107717 -2809 107771 -2753
rect 107827 -2809 107881 -2753
rect 107937 -2809 107963 -2753
rect 107175 -2863 107963 -2809
rect 107175 -2919 107221 -2863
rect 107277 -2919 107331 -2863
rect 107387 -2919 107441 -2863
rect 107497 -2919 107551 -2863
rect 107607 -2919 107661 -2863
rect 107717 -2919 107771 -2863
rect 107827 -2919 107881 -2863
rect 107937 -2919 107963 -2863
rect 107175 -2973 107963 -2919
rect 107175 -3029 107221 -2973
rect 107277 -3029 107331 -2973
rect 107387 -3029 107441 -2973
rect 107497 -3029 107551 -2973
rect 107607 -3029 107661 -2973
rect 107717 -3029 107771 -2973
rect 107827 -3029 107881 -2973
rect 107937 -3029 107963 -2973
rect 107175 -3083 107963 -3029
rect 107175 -3139 107221 -3083
rect 107277 -3139 107331 -3083
rect 107387 -3139 107441 -3083
rect 107497 -3139 107551 -3083
rect 107607 -3139 107661 -3083
rect 107717 -3139 107771 -3083
rect 107827 -3139 107881 -3083
rect 107937 -3139 107963 -3083
rect 30989 -4668 31209 -4612
rect 31265 -4668 31319 -4612
rect 31375 -4668 31429 -4612
rect 31485 -4668 31539 -4612
rect 31595 -4668 31776 -4612
rect 30989 -4738 31776 -4668
rect 31244 -11628 31777 -11619
rect 31244 -11684 31255 -11628
rect 31311 -11684 31365 -11628
rect 31421 -11684 31475 -11628
rect 31531 -11684 31585 -11628
rect 31641 -11684 31695 -11628
rect 31751 -11684 31777 -11628
rect 31244 -11738 31777 -11684
rect 31244 -11794 31255 -11738
rect 31311 -11794 31365 -11738
rect 31421 -11794 31475 -11738
rect 31531 -11794 31585 -11738
rect 31641 -11794 31695 -11738
rect 31751 -11794 31777 -11738
rect 31244 -11848 31777 -11794
rect 31244 -11904 31255 -11848
rect 31311 -11904 31365 -11848
rect 31421 -11904 31475 -11848
rect 31531 -11904 31585 -11848
rect 31641 -11904 31695 -11848
rect 31751 -11904 31777 -11848
rect 31244 -11958 31777 -11904
rect 31244 -12014 31255 -11958
rect 31311 -12014 31365 -11958
rect 31421 -12014 31475 -11958
rect 31531 -12014 31585 -11958
rect 31641 -12014 31695 -11958
rect 31751 -12014 31777 -11958
rect 31244 -12068 31777 -12014
rect 31244 -12124 31255 -12068
rect 31311 -12124 31365 -12068
rect 31421 -12124 31475 -12068
rect 31531 -12124 31585 -12068
rect 31641 -12124 31695 -12068
rect 31751 -12124 31777 -12068
rect 31244 -12161 31777 -12124
rect 29479 -13656 30536 -13568
rect 29479 -13664 30193 -13656
rect 29479 -13720 29533 -13664
rect 29589 -13720 29643 -13664
rect 29699 -13720 29753 -13664
rect 29809 -13720 29863 -13664
rect 29919 -13720 29973 -13664
rect 30029 -13720 30083 -13664
rect 30139 -13712 30193 -13664
rect 30249 -13712 30303 -13656
rect 30359 -13712 30413 -13656
rect 30469 -13712 30536 -13656
rect 30139 -13720 30536 -13712
rect 29479 -13766 30536 -13720
rect 29479 -13774 30193 -13766
rect 29479 -13830 29533 -13774
rect 29589 -13830 29643 -13774
rect 29699 -13830 29753 -13774
rect 29809 -13830 29863 -13774
rect 29919 -13830 29973 -13774
rect 30029 -13830 30083 -13774
rect 30139 -13822 30193 -13774
rect 30249 -13822 30303 -13766
rect 30359 -13822 30413 -13766
rect 30469 -13822 30536 -13766
rect 30139 -13830 30536 -13822
rect 29479 -13897 30536 -13830
rect 29799 -14469 30669 -14407
rect 29799 -14525 29852 -14469
rect 29908 -14525 29962 -14469
rect 30018 -14525 30072 -14469
rect 30128 -14525 30249 -14469
rect 30305 -14525 30359 -14469
rect 30415 -14525 30469 -14469
rect 30525 -14525 30669 -14469
rect 29799 -14579 30669 -14525
rect 29799 -14635 29852 -14579
rect 29908 -14635 29962 -14579
rect 30018 -14635 30072 -14579
rect 30128 -14635 30249 -14579
rect 30305 -14635 30359 -14579
rect 30415 -14635 30469 -14579
rect 30525 -14635 30669 -14579
rect 29799 -14722 30669 -14635
rect 31244 -15618 31776 -12161
rect 34037 -12382 34633 -12318
rect 34037 -12438 34121 -12382
rect 34177 -12438 34231 -12382
rect 34287 -12438 34341 -12382
rect 34397 -12438 34451 -12382
rect 34507 -12438 34633 -12382
rect 34037 -12492 34633 -12438
rect 34037 -12548 34121 -12492
rect 34177 -12548 34231 -12492
rect 34287 -12548 34341 -12492
rect 34397 -12548 34451 -12492
rect 34507 -12548 34633 -12492
rect 34037 -12602 34633 -12548
rect 34037 -12658 34121 -12602
rect 34177 -12658 34231 -12602
rect 34287 -12658 34341 -12602
rect 34397 -12658 34451 -12602
rect 34507 -12658 34633 -12602
rect 34037 -12712 34633 -12658
rect 34037 -12768 34121 -12712
rect 34177 -12768 34231 -12712
rect 34287 -12768 34341 -12712
rect 34397 -12768 34451 -12712
rect 34507 -12768 34633 -12712
rect 34037 -12827 34633 -12768
rect 36010 -12387 36795 -12344
rect 36010 -12443 36056 -12387
rect 36112 -12443 36166 -12387
rect 36222 -12443 36276 -12387
rect 36332 -12443 36386 -12387
rect 36442 -12443 36496 -12387
rect 36552 -12443 36606 -12387
rect 36662 -12443 36716 -12387
rect 36772 -12443 36795 -12387
rect 36010 -12497 36795 -12443
rect 36010 -12553 36056 -12497
rect 36112 -12553 36166 -12497
rect 36222 -12553 36276 -12497
rect 36332 -12553 36386 -12497
rect 36442 -12553 36496 -12497
rect 36552 -12553 36606 -12497
rect 36662 -12553 36716 -12497
rect 36772 -12553 36795 -12497
rect 36010 -12607 36795 -12553
rect 36010 -12663 36056 -12607
rect 36112 -12663 36166 -12607
rect 36222 -12663 36276 -12607
rect 36332 -12663 36386 -12607
rect 36442 -12663 36496 -12607
rect 36552 -12663 36606 -12607
rect 36662 -12663 36716 -12607
rect 36772 -12663 36795 -12607
rect 36010 -12717 36795 -12663
rect 36010 -12773 36056 -12717
rect 36112 -12773 36166 -12717
rect 36222 -12773 36276 -12717
rect 36332 -12773 36386 -12717
rect 36442 -12773 36496 -12717
rect 36552 -12773 36606 -12717
rect 36662 -12773 36716 -12717
rect 36772 -12773 36795 -12717
rect 36010 -12810 36795 -12773
rect 31244 -15674 31310 -15618
rect 31366 -15674 31420 -15618
rect 31476 -15674 31530 -15618
rect 31586 -15674 31640 -15618
rect 31696 -15674 31776 -15618
rect 31244 -15728 31776 -15674
rect 31244 -15784 31310 -15728
rect 31366 -15784 31420 -15728
rect 31476 -15784 31530 -15728
rect 31586 -15784 31640 -15728
rect 31696 -15784 31776 -15728
rect 31244 -15823 31776 -15784
rect 30854 -16519 31321 -16462
rect 28340 -16525 29304 -16521
rect 28338 -16558 29304 -16525
rect 28338 -16562 28873 -16558
rect 28338 -16618 28388 -16562
rect 28444 -16618 28498 -16562
rect 28554 -16618 28608 -16562
rect 28664 -16618 28718 -16562
rect 28774 -16614 28873 -16562
rect 28929 -16614 28983 -16558
rect 29039 -16614 29093 -16558
rect 29149 -16614 29203 -16558
rect 29259 -16614 29304 -16558
rect 28774 -16618 29304 -16614
rect 28338 -16668 29304 -16618
rect 28338 -16672 28873 -16668
rect 28338 -16728 28388 -16672
rect 28444 -16728 28498 -16672
rect 28554 -16728 28608 -16672
rect 28664 -16728 28718 -16672
rect 28774 -16724 28873 -16672
rect 28929 -16724 28983 -16668
rect 29039 -16724 29093 -16668
rect 29149 -16724 29203 -16668
rect 29259 -16724 29304 -16668
rect 28774 -16728 29304 -16724
rect 28338 -16778 29304 -16728
rect 28338 -16782 28873 -16778
rect 28338 -16838 28388 -16782
rect 28444 -16838 28498 -16782
rect 28554 -16838 28608 -16782
rect 28664 -16838 28718 -16782
rect 28774 -16834 28873 -16782
rect 28929 -16834 28983 -16778
rect 29039 -16834 29093 -16778
rect 29149 -16834 29203 -16778
rect 29259 -16834 29304 -16778
rect 28774 -16838 29304 -16834
rect 28338 -16888 29304 -16838
rect 28338 -16892 28873 -16888
rect 28338 -16948 28388 -16892
rect 28444 -16948 28498 -16892
rect 28554 -16948 28608 -16892
rect 28664 -16948 28718 -16892
rect 28774 -16944 28873 -16892
rect 28929 -16944 28983 -16888
rect 29039 -16944 29093 -16888
rect 29149 -16944 29203 -16888
rect 29259 -16944 29304 -16888
rect 28774 -16948 29304 -16944
rect 28338 -17014 29304 -16948
rect 30844 -16556 31325 -16519
rect 30844 -16612 30894 -16556
rect 30950 -16612 31004 -16556
rect 31060 -16612 31114 -16556
rect 31170 -16612 31224 -16556
rect 31280 -16612 31325 -16556
rect 30844 -16666 31325 -16612
rect 30844 -16722 30894 -16666
rect 30950 -16722 31004 -16666
rect 31060 -16722 31114 -16666
rect 31170 -16722 31224 -16666
rect 31280 -16722 31325 -16666
rect 30844 -16776 31325 -16722
rect 30844 -16832 30894 -16776
rect 30950 -16832 31004 -16776
rect 31060 -16832 31114 -16776
rect 31170 -16832 31224 -16776
rect 31280 -16832 31325 -16776
rect 30844 -16886 31325 -16832
rect 30844 -16942 30894 -16886
rect 30950 -16942 31004 -16886
rect 31060 -16942 31114 -16886
rect 31170 -16942 31224 -16886
rect 31280 -16942 31325 -16886
rect 30844 -17012 31325 -16942
rect 28338 -17018 29127 -17014
rect 28340 -17019 29127 -17018
rect 30162 -17411 30769 -17390
rect 30162 -17456 30771 -17411
rect 30162 -17512 30249 -17456
rect 30305 -17512 30359 -17456
rect 30415 -17512 30469 -17456
rect 30525 -17512 30579 -17456
rect 30635 -17512 30771 -17456
rect 30162 -17566 30771 -17512
rect 30162 -17622 30249 -17566
rect 30305 -17622 30359 -17566
rect 30415 -17622 30469 -17566
rect 30525 -17622 30579 -17566
rect 30635 -17622 30771 -17566
rect 30162 -17676 30771 -17622
rect 30162 -17732 30249 -17676
rect 30305 -17732 30359 -17676
rect 30415 -17732 30469 -17676
rect 30525 -17732 30579 -17676
rect 30635 -17732 30771 -17676
rect 30162 -17786 30771 -17732
rect 30162 -17842 30249 -17786
rect 30305 -17842 30359 -17786
rect 30415 -17842 30469 -17786
rect 30525 -17842 30579 -17786
rect 30635 -17842 30771 -17786
rect 30162 -17957 30771 -17842
rect 29741 -18335 30208 -18277
rect 29741 -18391 29788 -18335
rect 29844 -18391 29898 -18335
rect 29954 -18391 30008 -18335
rect 30064 -18391 30118 -18335
rect 30174 -18391 30208 -18335
rect 29741 -18445 30208 -18391
rect 29741 -18501 29788 -18445
rect 29844 -18501 29898 -18445
rect 29954 -18501 30008 -18445
rect 30064 -18501 30118 -18445
rect 30174 -18501 30208 -18445
rect 29741 -18573 30208 -18501
rect 29741 -18629 29782 -18573
rect 29838 -18629 29892 -18573
rect 29948 -18629 30002 -18573
rect 30058 -18629 30112 -18573
rect 30168 -18629 30208 -18573
rect 29741 -18683 30208 -18629
rect 29741 -18739 29782 -18683
rect 29838 -18739 29892 -18683
rect 29948 -18739 30002 -18683
rect 30058 -18739 30112 -18683
rect 30168 -18739 30208 -18683
rect 29741 -18793 30208 -18739
rect 29741 -18849 29782 -18793
rect 29838 -18849 29892 -18793
rect 29948 -18849 30002 -18793
rect 30058 -18849 30112 -18793
rect 30168 -18849 30208 -18793
rect 29741 -18903 30208 -18849
rect 29741 -18959 29782 -18903
rect 29838 -18959 29892 -18903
rect 29948 -18959 30002 -18903
rect 30058 -18959 30112 -18903
rect 30168 -18959 30208 -18903
rect 29741 -19778 30208 -18959
rect 29741 -19802 30209 -19778
rect 28768 -19951 29207 -19837
rect 29741 -19858 29779 -19802
rect 29835 -19858 29889 -19802
rect 29945 -19858 29999 -19802
rect 30055 -19858 30109 -19802
rect 30165 -19858 30209 -19802
rect 29741 -19879 30209 -19858
rect 30304 -19809 30771 -17957
rect 30304 -19865 30333 -19809
rect 30389 -19865 30443 -19809
rect 30499 -19865 30553 -19809
rect 30609 -19865 30663 -19809
rect 30719 -19865 30771 -19809
rect 29741 -19888 30208 -19879
rect 30304 -19895 30771 -19865
rect 30854 -19800 31321 -17012
rect 31430 -18619 31941 -18617
rect 31386 -18673 31942 -18619
rect 31386 -18729 31488 -18673
rect 31544 -18729 31598 -18673
rect 31654 -18729 31708 -18673
rect 31764 -18729 31818 -18673
rect 31874 -18729 31942 -18673
rect 31386 -18783 31942 -18729
rect 31386 -18839 31488 -18783
rect 31544 -18839 31598 -18783
rect 31654 -18839 31708 -18783
rect 31764 -18839 31818 -18783
rect 31874 -18839 31942 -18783
rect 31386 -18893 31942 -18839
rect 31386 -18949 31488 -18893
rect 31544 -18949 31598 -18893
rect 31654 -18949 31708 -18893
rect 31764 -18949 31818 -18893
rect 31874 -18949 31942 -18893
rect 31386 -19003 31942 -18949
rect 31386 -19059 31488 -19003
rect 31544 -19059 31598 -19003
rect 31654 -19059 31708 -19003
rect 31764 -19059 31818 -19003
rect 31874 -19059 31942 -19003
rect 31386 -19176 31942 -19059
rect 34040 -18725 34623 -12827
rect 107175 -16271 107963 -3139
rect 109049 -1002 109837 -951
rect 109049 -1058 109095 -1002
rect 109151 -1058 109205 -1002
rect 109261 -1058 109315 -1002
rect 109371 -1058 109425 -1002
rect 109481 -1058 109535 -1002
rect 109591 -1058 109645 -1002
rect 109701 -1058 109755 -1002
rect 109811 -1058 109837 -1002
rect 109049 -1112 109837 -1058
rect 109049 -1168 109095 -1112
rect 109151 -1168 109205 -1112
rect 109261 -1168 109315 -1112
rect 109371 -1168 109425 -1112
rect 109481 -1168 109535 -1112
rect 109591 -1168 109645 -1112
rect 109701 -1168 109755 -1112
rect 109811 -1168 109837 -1112
rect 109049 -1222 109837 -1168
rect 109049 -1278 109095 -1222
rect 109151 -1278 109205 -1222
rect 109261 -1278 109315 -1222
rect 109371 -1278 109425 -1222
rect 109481 -1278 109535 -1222
rect 109591 -1278 109645 -1222
rect 109701 -1278 109755 -1222
rect 109811 -1278 109837 -1222
rect 109049 -1332 109837 -1278
rect 109049 -1388 109095 -1332
rect 109151 -1388 109205 -1332
rect 109261 -1388 109315 -1332
rect 109371 -1388 109425 -1332
rect 109481 -1388 109535 -1332
rect 109591 -1388 109645 -1332
rect 109701 -1388 109755 -1332
rect 109811 -1388 109837 -1332
rect 109049 -1442 109837 -1388
rect 109049 -1498 109095 -1442
rect 109151 -1498 109205 -1442
rect 109261 -1498 109315 -1442
rect 109371 -1498 109425 -1442
rect 109481 -1498 109535 -1442
rect 109591 -1498 109645 -1442
rect 109701 -1498 109755 -1442
rect 109811 -1498 109837 -1442
rect 109049 -1552 109837 -1498
rect 109049 -1608 109095 -1552
rect 109151 -1608 109205 -1552
rect 109261 -1608 109315 -1552
rect 109371 -1608 109425 -1552
rect 109481 -1608 109535 -1552
rect 109591 -1608 109645 -1552
rect 109701 -1608 109755 -1552
rect 109811 -1608 109837 -1552
rect 109049 -1662 109837 -1608
rect 109049 -1718 109095 -1662
rect 109151 -1718 109205 -1662
rect 109261 -1718 109315 -1662
rect 109371 -1718 109425 -1662
rect 109481 -1718 109535 -1662
rect 109591 -1718 109645 -1662
rect 109701 -1718 109755 -1662
rect 109811 -1718 109837 -1662
rect 109049 -7895 109837 -1718
rect 109049 -7951 109078 -7895
rect 109134 -7951 109188 -7895
rect 109244 -7951 109298 -7895
rect 109354 -7951 109408 -7895
rect 109464 -7951 109518 -7895
rect 109574 -7951 109628 -7895
rect 109684 -7951 109738 -7895
rect 109794 -7951 109837 -7895
rect 109049 -8005 109837 -7951
rect 109049 -8061 109078 -8005
rect 109134 -8061 109188 -8005
rect 109244 -8061 109298 -8005
rect 109354 -8061 109408 -8005
rect 109464 -8061 109518 -8005
rect 109574 -8061 109628 -8005
rect 109684 -8061 109738 -8005
rect 109794 -8061 109837 -8005
rect 109049 -8115 109837 -8061
rect 109049 -8171 109078 -8115
rect 109134 -8171 109188 -8115
rect 109244 -8171 109298 -8115
rect 109354 -8171 109408 -8115
rect 109464 -8171 109518 -8115
rect 109574 -8171 109628 -8115
rect 109684 -8171 109738 -8115
rect 109794 -8171 109837 -8115
rect 109049 -8225 109837 -8171
rect 109049 -8281 109078 -8225
rect 109134 -8281 109188 -8225
rect 109244 -8281 109298 -8225
rect 109354 -8281 109408 -8225
rect 109464 -8281 109518 -8225
rect 109574 -8281 109628 -8225
rect 109684 -8281 109738 -8225
rect 109794 -8281 109837 -8225
rect 109049 -8335 109837 -8281
rect 109049 -8391 109078 -8335
rect 109134 -8391 109188 -8335
rect 109244 -8391 109298 -8335
rect 109354 -8391 109408 -8335
rect 109464 -8391 109518 -8335
rect 109574 -8391 109628 -8335
rect 109684 -8391 109738 -8335
rect 109794 -8391 109837 -8335
rect 109049 -8445 109837 -8391
rect 109049 -8501 109078 -8445
rect 109134 -8501 109188 -8445
rect 109244 -8501 109298 -8445
rect 109354 -8501 109408 -8445
rect 109464 -8501 109518 -8445
rect 109574 -8501 109628 -8445
rect 109684 -8501 109738 -8445
rect 109794 -8501 109837 -8445
rect 109049 -8555 109837 -8501
rect 109049 -8611 109078 -8555
rect 109134 -8611 109188 -8555
rect 109244 -8611 109298 -8555
rect 109354 -8611 109408 -8555
rect 109464 -8611 109518 -8555
rect 109574 -8611 109628 -8555
rect 109684 -8611 109738 -8555
rect 109794 -8611 109837 -8555
rect 109049 -8665 109837 -8611
rect 109049 -8721 109078 -8665
rect 109134 -8721 109188 -8665
rect 109244 -8721 109298 -8665
rect 109354 -8721 109408 -8665
rect 109464 -8721 109518 -8665
rect 109574 -8721 109628 -8665
rect 109684 -8721 109738 -8665
rect 109794 -8721 109837 -8665
rect 109049 -14902 109837 -8721
rect 109049 -14958 109096 -14902
rect 109152 -14958 109206 -14902
rect 109262 -14958 109316 -14902
rect 109372 -14958 109426 -14902
rect 109482 -14958 109536 -14902
rect 109592 -14958 109646 -14902
rect 109702 -14958 109756 -14902
rect 109812 -14958 109837 -14902
rect 109049 -15012 109837 -14958
rect 109049 -15068 109096 -15012
rect 109152 -15068 109206 -15012
rect 109262 -15068 109316 -15012
rect 109372 -15068 109426 -15012
rect 109482 -15068 109536 -15012
rect 109592 -15068 109646 -15012
rect 109702 -15068 109756 -15012
rect 109812 -15068 109837 -15012
rect 109049 -15122 109837 -15068
rect 109049 -15178 109096 -15122
rect 109152 -15178 109206 -15122
rect 109262 -15178 109316 -15122
rect 109372 -15178 109426 -15122
rect 109482 -15178 109536 -15122
rect 109592 -15178 109646 -15122
rect 109702 -15178 109756 -15122
rect 109812 -15178 109837 -15122
rect 109049 -15232 109837 -15178
rect 109049 -15288 109096 -15232
rect 109152 -15288 109206 -15232
rect 109262 -15288 109316 -15232
rect 109372 -15288 109426 -15232
rect 109482 -15288 109536 -15232
rect 109592 -15288 109646 -15232
rect 109702 -15288 109756 -15232
rect 109812 -15288 109837 -15232
rect 109049 -15342 109837 -15288
rect 109049 -15398 109096 -15342
rect 109152 -15398 109206 -15342
rect 109262 -15398 109316 -15342
rect 109372 -15398 109426 -15342
rect 109482 -15398 109536 -15342
rect 109592 -15398 109646 -15342
rect 109702 -15398 109756 -15342
rect 109812 -15398 109837 -15342
rect 109049 -15452 109837 -15398
rect 109049 -15508 109096 -15452
rect 109152 -15508 109206 -15452
rect 109262 -15508 109316 -15452
rect 109372 -15508 109426 -15452
rect 109482 -15508 109536 -15452
rect 109592 -15508 109646 -15452
rect 109702 -15508 109756 -15452
rect 109812 -15508 109837 -15452
rect 109049 -15562 109837 -15508
rect 109049 -15618 109096 -15562
rect 109152 -15618 109206 -15562
rect 109262 -15618 109316 -15562
rect 109372 -15618 109426 -15562
rect 109482 -15618 109536 -15562
rect 109592 -15618 109646 -15562
rect 109702 -15618 109756 -15562
rect 109812 -15618 109837 -15562
rect 109049 -15656 109837 -15618
rect 107175 -16327 107210 -16271
rect 107266 -16327 107320 -16271
rect 107376 -16327 107430 -16271
rect 107486 -16327 107540 -16271
rect 107596 -16327 107650 -16271
rect 107706 -16327 107760 -16271
rect 107816 -16327 107870 -16271
rect 107926 -16327 107963 -16271
rect 107175 -16381 107963 -16327
rect 107175 -16437 107210 -16381
rect 107266 -16437 107320 -16381
rect 107376 -16437 107430 -16381
rect 107486 -16437 107540 -16381
rect 107596 -16437 107650 -16381
rect 107706 -16437 107760 -16381
rect 107816 -16437 107870 -16381
rect 107926 -16437 107963 -16381
rect 107175 -16491 107963 -16437
rect 107175 -16547 107210 -16491
rect 107266 -16547 107320 -16491
rect 107376 -16547 107430 -16491
rect 107486 -16547 107540 -16491
rect 107596 -16547 107650 -16491
rect 107706 -16547 107760 -16491
rect 107816 -16547 107870 -16491
rect 107926 -16547 107963 -16491
rect 107175 -16601 107963 -16547
rect 107175 -16657 107210 -16601
rect 107266 -16657 107320 -16601
rect 107376 -16657 107430 -16601
rect 107486 -16657 107540 -16601
rect 107596 -16657 107650 -16601
rect 107706 -16657 107760 -16601
rect 107816 -16657 107870 -16601
rect 107926 -16657 107963 -16601
rect 107175 -16711 107963 -16657
rect 107175 -16767 107210 -16711
rect 107266 -16767 107320 -16711
rect 107376 -16767 107430 -16711
rect 107486 -16767 107540 -16711
rect 107596 -16767 107650 -16711
rect 107706 -16767 107760 -16711
rect 107816 -16767 107870 -16711
rect 107926 -16767 107963 -16711
rect 107175 -16821 107963 -16767
rect 107175 -16877 107210 -16821
rect 107266 -16877 107320 -16821
rect 107376 -16877 107430 -16821
rect 107486 -16877 107540 -16821
rect 107596 -16877 107650 -16821
rect 107706 -16877 107760 -16821
rect 107816 -16877 107870 -16821
rect 107926 -16877 107963 -16821
rect 107175 -16931 107963 -16877
rect 107175 -16987 107210 -16931
rect 107266 -16987 107320 -16931
rect 107376 -16987 107430 -16931
rect 107486 -16987 107540 -16931
rect 107596 -16987 107650 -16931
rect 107706 -16987 107760 -16931
rect 107816 -16987 107870 -16931
rect 107926 -16987 107963 -16931
rect 107175 -17023 107963 -16987
rect 34040 -18781 34132 -18725
rect 34188 -18781 34242 -18725
rect 34298 -18781 34352 -18725
rect 34408 -18781 34462 -18725
rect 34518 -18781 34623 -18725
rect 34040 -18835 34623 -18781
rect 34040 -18891 34132 -18835
rect 34188 -18891 34242 -18835
rect 34298 -18891 34352 -18835
rect 34408 -18891 34462 -18835
rect 34518 -18891 34623 -18835
rect 34040 -18945 34623 -18891
rect 34040 -19001 34132 -18945
rect 34188 -19001 34242 -18945
rect 34298 -19001 34352 -18945
rect 34408 -19001 34462 -18945
rect 34518 -19001 34623 -18945
rect 34040 -19055 34623 -19001
rect 34040 -19111 34132 -19055
rect 34188 -19111 34242 -19055
rect 34298 -19111 34352 -19055
rect 34408 -19111 34462 -19055
rect 34518 -19111 34623 -19055
rect 34040 -19173 34623 -19111
rect 94333 -18639 94715 -18638
rect 94333 -18675 94768 -18639
rect 94333 -18731 94359 -18675
rect 94415 -18731 94469 -18675
rect 94525 -18731 94579 -18675
rect 94635 -18731 94689 -18675
rect 94745 -18731 94768 -18675
rect 94333 -18785 94768 -18731
rect 94333 -18841 94359 -18785
rect 94415 -18841 94469 -18785
rect 94525 -18841 94579 -18785
rect 94635 -18841 94689 -18785
rect 94745 -18841 94768 -18785
rect 94333 -18895 94768 -18841
rect 94333 -18951 94359 -18895
rect 94415 -18951 94469 -18895
rect 94525 -18951 94579 -18895
rect 94635 -18951 94689 -18895
rect 94745 -18951 94768 -18895
rect 94333 -19005 94768 -18951
rect 94333 -19061 94359 -19005
rect 94415 -19061 94469 -19005
rect 94525 -19061 94579 -19005
rect 94635 -19061 94689 -19005
rect 94745 -19061 94768 -19005
rect 94333 -19115 94768 -19061
rect 94333 -19171 94359 -19115
rect 94415 -19171 94469 -19115
rect 94525 -19171 94579 -19115
rect 94635 -19171 94689 -19115
rect 94745 -19171 94768 -19115
rect 30854 -19856 30887 -19800
rect 30943 -19856 30997 -19800
rect 31053 -19856 31107 -19800
rect 31163 -19856 31217 -19800
rect 31273 -19856 31321 -19800
rect 30854 -19882 31321 -19856
rect 31391 -19816 31888 -19176
rect 94333 -19225 94768 -19171
rect 94333 -19281 94359 -19225
rect 94415 -19281 94469 -19225
rect 94525 -19281 94579 -19225
rect 94635 -19281 94689 -19225
rect 94745 -19281 94768 -19225
rect 94333 -19335 94768 -19281
rect 94333 -19391 94359 -19335
rect 94415 -19391 94469 -19335
rect 94525 -19391 94579 -19335
rect 94635 -19391 94689 -19335
rect 94745 -19391 94768 -19335
rect 94333 -19432 94768 -19391
rect 31391 -19872 31427 -19816
rect 31483 -19872 31537 -19816
rect 31593 -19872 31647 -19816
rect 31703 -19872 31757 -19816
rect 31813 -19872 31888 -19816
rect 31391 -19908 31888 -19872
rect 28768 -20007 28803 -19951
rect 28859 -20007 28913 -19951
rect 28969 -20007 29023 -19951
rect 29079 -20007 29133 -19951
rect 29189 -20007 29207 -19951
rect 28768 -20061 29207 -20007
rect 28768 -20117 28803 -20061
rect 28859 -20117 28913 -20061
rect 28969 -20117 29023 -20061
rect 29079 -20117 29133 -20061
rect 29189 -20117 29207 -20061
rect 28768 -20189 29207 -20117
rect 28768 -20245 28797 -20189
rect 28853 -20245 28907 -20189
rect 28963 -20245 29017 -20189
rect 29073 -20245 29127 -20189
rect 29183 -20245 29207 -20189
rect 28768 -20299 29207 -20245
rect 28768 -20355 28797 -20299
rect 28853 -20355 28907 -20299
rect 28963 -20355 29017 -20299
rect 29073 -20355 29127 -20299
rect 29183 -20355 29207 -20299
rect 28768 -20409 29207 -20355
rect 28768 -20465 28797 -20409
rect 28853 -20465 28907 -20409
rect 28963 -20465 29017 -20409
rect 29073 -20465 29127 -20409
rect 29183 -20465 29207 -20409
rect 28768 -20519 29207 -20465
rect 28768 -20575 28797 -20519
rect 28853 -20575 28907 -20519
rect 28963 -20575 29017 -20519
rect 29073 -20575 29127 -20519
rect 29183 -20575 29207 -20519
rect 28768 -20592 29207 -20575
rect 28837 -20718 29216 -20717
rect 28770 -20805 29216 -20718
rect 28770 -20861 28796 -20805
rect 28852 -20861 28906 -20805
rect 28962 -20861 29016 -20805
rect 29072 -20861 29126 -20805
rect 29182 -20861 29216 -20805
rect 93813 -20845 93869 -19564
rect 94077 -19869 94133 -19523
rect 94075 -19873 94510 -19869
rect 94074 -19905 94510 -19873
rect 94074 -19961 94101 -19905
rect 94157 -19961 94211 -19905
rect 94267 -19961 94321 -19905
rect 94377 -19961 94431 -19905
rect 94487 -19961 94510 -19905
rect 94074 -20015 94510 -19961
rect 94074 -20071 94101 -20015
rect 94157 -20071 94211 -20015
rect 94267 -20071 94321 -20015
rect 94377 -20071 94431 -20015
rect 94487 -20071 94510 -20015
rect 94074 -20125 94510 -20071
rect 94074 -20181 94101 -20125
rect 94157 -20181 94211 -20125
rect 94267 -20181 94321 -20125
rect 94377 -20181 94431 -20125
rect 94487 -20181 94510 -20125
rect 94074 -20235 94510 -20181
rect 94074 -20291 94101 -20235
rect 94157 -20291 94211 -20235
rect 94267 -20291 94321 -20235
rect 94377 -20291 94431 -20235
rect 94487 -20291 94510 -20235
rect 94074 -20345 94510 -20291
rect 94074 -20401 94101 -20345
rect 94157 -20401 94211 -20345
rect 94267 -20401 94321 -20345
rect 94377 -20401 94431 -20345
rect 94487 -20401 94510 -20345
rect 94074 -20455 94510 -20401
rect 94074 -20511 94101 -20455
rect 94157 -20511 94211 -20455
rect 94267 -20511 94321 -20455
rect 94377 -20511 94431 -20455
rect 94487 -20511 94510 -20455
rect 94074 -20565 94510 -20511
rect 94074 -20621 94101 -20565
rect 94157 -20621 94211 -20565
rect 94267 -20621 94321 -20565
rect 94377 -20621 94431 -20565
rect 94487 -20621 94510 -20565
rect 94074 -20661 94510 -20621
rect 94075 -20662 94510 -20661
rect 28770 -20915 29216 -20861
rect 28770 -20971 28796 -20915
rect 28852 -20971 28906 -20915
rect 28962 -20971 29016 -20915
rect 29072 -20971 29126 -20915
rect 29182 -20971 29216 -20915
rect 28770 -21043 29216 -20971
rect 28770 -21099 28790 -21043
rect 28846 -21099 28900 -21043
rect 28956 -21099 29010 -21043
rect 29066 -21099 29120 -21043
rect 29176 -21099 29216 -21043
rect 28770 -21153 29216 -21099
rect 28770 -21209 28790 -21153
rect 28846 -21209 28900 -21153
rect 28956 -21209 29010 -21153
rect 29066 -21209 29120 -21153
rect 29176 -21209 29216 -21153
rect 28770 -21263 29216 -21209
rect 28770 -21319 28790 -21263
rect 28846 -21319 28900 -21263
rect 28956 -21319 29010 -21263
rect 29066 -21319 29120 -21263
rect 29176 -21319 29216 -21263
rect 28770 -21373 29216 -21319
rect 28770 -21429 28790 -21373
rect 28846 -21429 28900 -21373
rect 28956 -21429 29010 -21373
rect 29066 -21429 29120 -21373
rect 29176 -21429 29216 -21373
rect 28770 -21473 29216 -21429
rect 93809 -20846 94191 -20845
rect 93809 -20882 94245 -20846
rect 93809 -20938 93836 -20882
rect 93892 -20938 93946 -20882
rect 94002 -20938 94056 -20882
rect 94112 -20938 94166 -20882
rect 94222 -20938 94245 -20882
rect 93809 -20992 94245 -20938
rect 93809 -21048 93836 -20992
rect 93892 -21048 93946 -20992
rect 94002 -21048 94056 -20992
rect 94112 -21048 94166 -20992
rect 94222 -21048 94245 -20992
rect 93809 -21102 94245 -21048
rect 93809 -21158 93836 -21102
rect 93892 -21158 93946 -21102
rect 94002 -21158 94056 -21102
rect 94112 -21158 94166 -21102
rect 94222 -21158 94245 -21102
rect 93809 -21212 94245 -21158
rect 93809 -21268 93836 -21212
rect 93892 -21268 93946 -21212
rect 94002 -21268 94056 -21212
rect 94112 -21268 94166 -21212
rect 94222 -21268 94245 -21212
rect 93809 -21322 94245 -21268
rect 93809 -21378 93836 -21322
rect 93892 -21378 93946 -21322
rect 94002 -21378 94056 -21322
rect 94112 -21378 94166 -21322
rect 94222 -21378 94245 -21322
rect 93809 -21432 94245 -21378
rect 93809 -21488 93836 -21432
rect 93892 -21488 93946 -21432
rect 94002 -21488 94056 -21432
rect 94112 -21488 94166 -21432
rect 94222 -21488 94245 -21432
rect 93809 -21542 94245 -21488
rect 93809 -21598 93836 -21542
rect 93892 -21598 93946 -21542
rect 94002 -21598 94056 -21542
rect 94112 -21598 94166 -21542
rect 94222 -21598 94245 -21542
rect 93809 -21633 94245 -21598
rect 93810 -21639 94245 -21633
rect 27246 -22741 27330 -22685
rect 27386 -22741 27440 -22685
rect 27496 -22741 27550 -22685
rect 27606 -22741 27660 -22685
rect 27716 -22741 27775 -22685
rect 27246 -22795 27775 -22741
rect 27246 -22851 27330 -22795
rect 27386 -22851 27440 -22795
rect 27496 -22851 27550 -22795
rect 27606 -22851 27660 -22795
rect 27716 -22851 27775 -22795
rect 27246 -22923 27775 -22851
rect 27246 -22979 27324 -22923
rect 27380 -22979 27434 -22923
rect 27490 -22979 27544 -22923
rect 27600 -22979 27654 -22923
rect 27710 -22979 27775 -22923
rect 27246 -23033 27775 -22979
rect 27246 -23089 27324 -23033
rect 27380 -23089 27434 -23033
rect 27490 -23089 27544 -23033
rect 27600 -23089 27654 -23033
rect 27710 -23089 27775 -23033
rect 27246 -23143 27775 -23089
rect 27246 -23199 27324 -23143
rect 27380 -23199 27434 -23143
rect 27490 -23199 27544 -23143
rect 27600 -23199 27654 -23143
rect 27710 -23199 27775 -23143
rect 27246 -23253 27775 -23199
rect 27246 -23309 27324 -23253
rect 27380 -23309 27434 -23253
rect 27490 -23309 27544 -23253
rect 27600 -23309 27654 -23253
rect 27710 -23309 27775 -23253
rect 27246 -23412 27775 -23309
rect 56571 -27818 57329 -27796
rect 56571 -27874 56591 -27818
rect 56647 -27874 56701 -27818
rect 56757 -27874 56811 -27818
rect 56867 -27874 56921 -27818
rect 56977 -27874 57031 -27818
rect 57087 -27874 57141 -27818
rect 57197 -27874 57251 -27818
rect 57307 -27874 57329 -27818
rect 56571 -27928 57329 -27874
rect 56571 -27984 56591 -27928
rect 56647 -27984 56701 -27928
rect 56757 -27984 56811 -27928
rect 56867 -27984 56921 -27928
rect 56977 -27984 57031 -27928
rect 57087 -27984 57141 -27928
rect 57197 -27984 57251 -27928
rect 57307 -27984 57329 -27928
rect 56571 -28038 57329 -27984
rect 56571 -28094 56591 -28038
rect 56647 -28094 56701 -28038
rect 56757 -28094 56811 -28038
rect 56867 -28094 56921 -28038
rect 56977 -28094 57031 -28038
rect 57087 -28094 57141 -28038
rect 57197 -28094 57251 -28038
rect 57307 -28094 57329 -28038
rect 56571 -28148 57329 -28094
rect 56571 -28204 56591 -28148
rect 56647 -28204 56701 -28148
rect 56757 -28204 56811 -28148
rect 56867 -28204 56921 -28148
rect 56977 -28204 57031 -28148
rect 57087 -28204 57141 -28148
rect 57197 -28204 57251 -28148
rect 57307 -28204 57329 -28148
rect 56571 -28258 57329 -28204
rect 56571 -28314 56591 -28258
rect 56647 -28314 56701 -28258
rect 56757 -28314 56811 -28258
rect 56867 -28314 56921 -28258
rect 56977 -28314 57031 -28258
rect 57087 -28314 57141 -28258
rect 57197 -28314 57251 -28258
rect 57307 -28314 57329 -28258
rect 56571 -28368 57329 -28314
rect 56571 -28424 56591 -28368
rect 56647 -28424 56701 -28368
rect 56757 -28424 56811 -28368
rect 56867 -28424 56921 -28368
rect 56977 -28424 57031 -28368
rect 57087 -28424 57141 -28368
rect 57197 -28424 57251 -28368
rect 57307 -28424 57329 -28368
rect 56571 -28478 57329 -28424
rect 56571 -28534 56591 -28478
rect 56647 -28534 56701 -28478
rect 56757 -28534 56811 -28478
rect 56867 -28534 56921 -28478
rect 56977 -28534 57031 -28478
rect 57087 -28534 57141 -28478
rect 57197 -28534 57251 -28478
rect 57307 -28534 57329 -28478
rect 56571 -28588 57329 -28534
rect 56571 -28644 56591 -28588
rect 56647 -28644 56701 -28588
rect 56757 -28644 56811 -28588
rect 56867 -28644 56921 -28588
rect 56977 -28644 57031 -28588
rect 57087 -28644 57141 -28588
rect 57197 -28644 57251 -28588
rect 57307 -28644 57329 -28588
rect 56571 -28703 57329 -28644
rect 39287 -28947 40045 -28925
rect 39287 -29003 39307 -28947
rect 39363 -29003 39417 -28947
rect 39473 -29003 39527 -28947
rect 39583 -29003 39637 -28947
rect 39693 -29003 39747 -28947
rect 39803 -29003 39857 -28947
rect 39913 -29003 39967 -28947
rect 40023 -29003 40045 -28947
rect 39287 -29057 40045 -29003
rect 39287 -29113 39307 -29057
rect 39363 -29113 39417 -29057
rect 39473 -29113 39527 -29057
rect 39583 -29113 39637 -29057
rect 39693 -29113 39747 -29057
rect 39803 -29113 39857 -29057
rect 39913 -29113 39967 -29057
rect 40023 -29113 40045 -29057
rect 39287 -29167 40045 -29113
rect 39287 -29223 39307 -29167
rect 39363 -29223 39417 -29167
rect 39473 -29223 39527 -29167
rect 39583 -29223 39637 -29167
rect 39693 -29223 39747 -29167
rect 39803 -29223 39857 -29167
rect 39913 -29223 39967 -29167
rect 40023 -29223 40045 -29167
rect 39287 -29277 40045 -29223
rect 39287 -29333 39307 -29277
rect 39363 -29333 39417 -29277
rect 39473 -29333 39527 -29277
rect 39583 -29333 39637 -29277
rect 39693 -29333 39747 -29277
rect 39803 -29333 39857 -29277
rect 39913 -29333 39967 -29277
rect 40023 -29333 40045 -29277
rect 39287 -29387 40045 -29333
rect 39287 -29443 39307 -29387
rect 39363 -29443 39417 -29387
rect 39473 -29443 39527 -29387
rect 39583 -29443 39637 -29387
rect 39693 -29443 39747 -29387
rect 39803 -29443 39857 -29387
rect 39913 -29443 39967 -29387
rect 40023 -29443 40045 -29387
rect 39287 -29497 40045 -29443
rect 39287 -29553 39307 -29497
rect 39363 -29553 39417 -29497
rect 39473 -29553 39527 -29497
rect 39583 -29553 39637 -29497
rect 39693 -29553 39747 -29497
rect 39803 -29553 39857 -29497
rect 39913 -29553 39967 -29497
rect 40023 -29553 40045 -29497
rect 39287 -29607 40045 -29553
rect 39287 -29663 39307 -29607
rect 39363 -29663 39417 -29607
rect 39473 -29663 39527 -29607
rect 39583 -29663 39637 -29607
rect 39693 -29663 39747 -29607
rect 39803 -29663 39857 -29607
rect 39913 -29663 39967 -29607
rect 40023 -29663 40045 -29607
rect 39287 -29717 40045 -29663
rect 39287 -29773 39307 -29717
rect 39363 -29773 39417 -29717
rect 39473 -29773 39527 -29717
rect 39583 -29773 39637 -29717
rect 39693 -29773 39747 -29717
rect 39803 -29773 39857 -29717
rect 39913 -29773 39967 -29717
rect 40023 -29773 40045 -29717
rect 39287 -29832 40045 -29773
rect 110594 -29024 111580 1030
rect 112010 -27858 112992 16506
rect 112010 -27914 112129 -27858
rect 112185 -27914 112239 -27858
rect 112295 -27914 112349 -27858
rect 112405 -27914 112459 -27858
rect 112515 -27914 112569 -27858
rect 112625 -27914 112679 -27858
rect 112735 -27914 112789 -27858
rect 112845 -27914 112992 -27858
rect 112010 -27968 112992 -27914
rect 112010 -28024 112129 -27968
rect 112185 -28024 112239 -27968
rect 112295 -28024 112349 -27968
rect 112405 -28024 112459 -27968
rect 112515 -28024 112569 -27968
rect 112625 -28024 112679 -27968
rect 112735 -28024 112789 -27968
rect 112845 -28024 112992 -27968
rect 112010 -28078 112992 -28024
rect 112010 -28134 112129 -28078
rect 112185 -28134 112239 -28078
rect 112295 -28134 112349 -28078
rect 112405 -28134 112459 -28078
rect 112515 -28134 112569 -28078
rect 112625 -28134 112679 -28078
rect 112735 -28134 112789 -28078
rect 112845 -28134 112992 -28078
rect 112010 -28188 112992 -28134
rect 112010 -28244 112129 -28188
rect 112185 -28244 112239 -28188
rect 112295 -28244 112349 -28188
rect 112405 -28244 112459 -28188
rect 112515 -28244 112569 -28188
rect 112625 -28244 112679 -28188
rect 112735 -28244 112789 -28188
rect 112845 -28244 112992 -28188
rect 112010 -28298 112992 -28244
rect 112010 -28354 112129 -28298
rect 112185 -28354 112239 -28298
rect 112295 -28354 112349 -28298
rect 112405 -28354 112459 -28298
rect 112515 -28354 112569 -28298
rect 112625 -28354 112679 -28298
rect 112735 -28354 112789 -28298
rect 112845 -28354 112992 -28298
rect 112010 -28408 112992 -28354
rect 112010 -28464 112129 -28408
rect 112185 -28464 112239 -28408
rect 112295 -28464 112349 -28408
rect 112405 -28464 112459 -28408
rect 112515 -28464 112569 -28408
rect 112625 -28464 112679 -28408
rect 112735 -28464 112789 -28408
rect 112845 -28464 112992 -28408
rect 112010 -28518 112992 -28464
rect 112010 -28574 112129 -28518
rect 112185 -28574 112239 -28518
rect 112295 -28574 112349 -28518
rect 112405 -28574 112459 -28518
rect 112515 -28574 112569 -28518
rect 112625 -28574 112679 -28518
rect 112735 -28574 112789 -28518
rect 112845 -28574 112992 -28518
rect 112010 -28703 112992 -28574
rect 113495 13098 114395 19254
rect 113495 13042 113535 13098
rect 113591 13042 113645 13098
rect 113701 13042 113755 13098
rect 113811 13042 113865 13098
rect 113921 13042 113975 13098
rect 114031 13042 114085 13098
rect 114141 13042 114195 13098
rect 114251 13042 114395 13098
rect 113495 12988 114395 13042
rect 113495 12932 113535 12988
rect 113591 12932 113645 12988
rect 113701 12932 113755 12988
rect 113811 12932 113865 12988
rect 113921 12932 113975 12988
rect 114031 12932 114085 12988
rect 114141 12932 114195 12988
rect 114251 12932 114395 12988
rect 113495 12878 114395 12932
rect 113495 12822 113535 12878
rect 113591 12822 113645 12878
rect 113701 12822 113755 12878
rect 113811 12822 113865 12878
rect 113921 12822 113975 12878
rect 114031 12822 114085 12878
rect 114141 12822 114195 12878
rect 114251 12822 114395 12878
rect 113495 12768 114395 12822
rect 113495 12712 113535 12768
rect 113591 12712 113645 12768
rect 113701 12712 113755 12768
rect 113811 12712 113865 12768
rect 113921 12712 113975 12768
rect 114031 12712 114085 12768
rect 114141 12712 114195 12768
rect 114251 12712 114395 12768
rect 113495 12658 114395 12712
rect 113495 12602 113535 12658
rect 113591 12602 113645 12658
rect 113701 12602 113755 12658
rect 113811 12602 113865 12658
rect 113921 12602 113975 12658
rect 114031 12602 114085 12658
rect 114141 12602 114195 12658
rect 114251 12602 114395 12658
rect 113495 12548 114395 12602
rect 113495 12492 113535 12548
rect 113591 12492 113645 12548
rect 113701 12492 113755 12548
rect 113811 12492 113865 12548
rect 113921 12492 113975 12548
rect 114031 12492 114085 12548
rect 114141 12492 114195 12548
rect 114251 12492 114395 12548
rect 113495 211 114395 12492
rect 113495 155 113565 211
rect 113621 155 113675 211
rect 113731 155 113785 211
rect 113841 155 113895 211
rect 113951 155 114005 211
rect 114061 155 114115 211
rect 114171 155 114225 211
rect 114281 155 114395 211
rect 113495 101 114395 155
rect 113495 45 113565 101
rect 113621 45 113675 101
rect 113731 45 113785 101
rect 113841 45 113895 101
rect 113951 45 114005 101
rect 114061 45 114115 101
rect 114171 45 114225 101
rect 114281 45 114395 101
rect 113495 -9 114395 45
rect 113495 -65 113565 -9
rect 113621 -65 113675 -9
rect 113731 -65 113785 -9
rect 113841 -65 113895 -9
rect 113951 -65 114005 -9
rect 114061 -65 114115 -9
rect 114171 -65 114225 -9
rect 114281 -65 114395 -9
rect 113495 -119 114395 -65
rect 113495 -175 113565 -119
rect 113621 -175 113675 -119
rect 113731 -175 113785 -119
rect 113841 -175 113895 -119
rect 113951 -175 114005 -119
rect 114061 -175 114115 -119
rect 114171 -175 114225 -119
rect 114281 -175 114395 -119
rect 113495 -229 114395 -175
rect 113495 -285 113565 -229
rect 113621 -285 113675 -229
rect 113731 -285 113785 -229
rect 113841 -285 113895 -229
rect 113951 -285 114005 -229
rect 114061 -285 114115 -229
rect 114171 -285 114225 -229
rect 114281 -285 114395 -229
rect 113495 -339 114395 -285
rect 113495 -395 113565 -339
rect 113621 -395 113675 -339
rect 113731 -395 113785 -339
rect 113841 -395 113895 -339
rect 113951 -395 114005 -339
rect 114061 -395 114115 -339
rect 114171 -395 114225 -339
rect 114281 -395 114395 -339
rect 113495 -2289 114395 -395
rect 113495 -2345 113560 -2289
rect 113616 -2345 113670 -2289
rect 113726 -2345 113780 -2289
rect 113836 -2345 113890 -2289
rect 113946 -2345 114000 -2289
rect 114056 -2345 114110 -2289
rect 114166 -2345 114220 -2289
rect 114276 -2345 114395 -2289
rect 113495 -2399 114395 -2345
rect 113495 -2455 113560 -2399
rect 113616 -2455 113670 -2399
rect 113726 -2455 113780 -2399
rect 113836 -2455 113890 -2399
rect 113946 -2455 114000 -2399
rect 114056 -2455 114110 -2399
rect 114166 -2455 114220 -2399
rect 114276 -2455 114395 -2399
rect 113495 -2509 114395 -2455
rect 113495 -2565 113560 -2509
rect 113616 -2565 113670 -2509
rect 113726 -2565 113780 -2509
rect 113836 -2565 113890 -2509
rect 113946 -2565 114000 -2509
rect 114056 -2565 114110 -2509
rect 114166 -2565 114220 -2509
rect 114276 -2565 114395 -2509
rect 113495 -2619 114395 -2565
rect 113495 -2675 113560 -2619
rect 113616 -2675 113670 -2619
rect 113726 -2675 113780 -2619
rect 113836 -2675 113890 -2619
rect 113946 -2675 114000 -2619
rect 114056 -2675 114110 -2619
rect 114166 -2675 114220 -2619
rect 114276 -2675 114395 -2619
rect 113495 -2729 114395 -2675
rect 113495 -2785 113560 -2729
rect 113616 -2785 113670 -2729
rect 113726 -2785 113780 -2729
rect 113836 -2785 113890 -2729
rect 113946 -2785 114000 -2729
rect 114056 -2785 114110 -2729
rect 114166 -2785 114220 -2729
rect 114276 -2785 114395 -2729
rect 113495 -2839 114395 -2785
rect 113495 -2895 113560 -2839
rect 113616 -2895 113670 -2839
rect 113726 -2895 113780 -2839
rect 113836 -2895 113890 -2839
rect 113946 -2895 114000 -2839
rect 114056 -2895 114110 -2839
rect 114166 -2895 114220 -2839
rect 114276 -2895 114395 -2839
rect 113495 -13207 114395 -2895
rect 113495 -13263 113550 -13207
rect 113606 -13263 113660 -13207
rect 113716 -13263 113770 -13207
rect 113826 -13263 113880 -13207
rect 113936 -13263 113990 -13207
rect 114046 -13263 114100 -13207
rect 114156 -13263 114210 -13207
rect 114266 -13263 114395 -13207
rect 113495 -13317 114395 -13263
rect 113495 -13373 113550 -13317
rect 113606 -13373 113660 -13317
rect 113716 -13373 113770 -13317
rect 113826 -13373 113880 -13317
rect 113936 -13373 113990 -13317
rect 114046 -13373 114100 -13317
rect 114156 -13373 114210 -13317
rect 114266 -13373 114395 -13317
rect 113495 -13427 114395 -13373
rect 113495 -13483 113550 -13427
rect 113606 -13483 113660 -13427
rect 113716 -13483 113770 -13427
rect 113826 -13483 113880 -13427
rect 113936 -13483 113990 -13427
rect 114046 -13483 114100 -13427
rect 114156 -13483 114210 -13427
rect 114266 -13483 114395 -13427
rect 113495 -13537 114395 -13483
rect 113495 -13593 113550 -13537
rect 113606 -13593 113660 -13537
rect 113716 -13593 113770 -13537
rect 113826 -13593 113880 -13537
rect 113936 -13593 113990 -13537
rect 114046 -13593 114100 -13537
rect 114156 -13593 114210 -13537
rect 114266 -13593 114395 -13537
rect 113495 -13647 114395 -13593
rect 113495 -13703 113550 -13647
rect 113606 -13703 113660 -13647
rect 113716 -13703 113770 -13647
rect 113826 -13703 113880 -13647
rect 113936 -13703 113990 -13647
rect 114046 -13703 114100 -13647
rect 114156 -13703 114210 -13647
rect 114266 -13703 114395 -13647
rect 113495 -13757 114395 -13703
rect 113495 -13813 113550 -13757
rect 113606 -13813 113660 -13757
rect 113716 -13813 113770 -13757
rect 113826 -13813 113880 -13757
rect 113936 -13813 113990 -13757
rect 114046 -13813 114100 -13757
rect 114156 -13813 114210 -13757
rect 114266 -13813 114395 -13757
rect 110594 -29080 110768 -29024
rect 110824 -29080 110878 -29024
rect 110934 -29080 110988 -29024
rect 111044 -29080 111098 -29024
rect 111154 -29080 111208 -29024
rect 111264 -29080 111318 -29024
rect 111374 -29080 111428 -29024
rect 111484 -29080 111580 -29024
rect 110594 -29134 111580 -29080
rect 110594 -29190 110768 -29134
rect 110824 -29190 110878 -29134
rect 110934 -29190 110988 -29134
rect 111044 -29190 111098 -29134
rect 111154 -29190 111208 -29134
rect 111264 -29190 111318 -29134
rect 111374 -29190 111428 -29134
rect 111484 -29190 111580 -29134
rect 110594 -29244 111580 -29190
rect 110594 -29300 110768 -29244
rect 110824 -29300 110878 -29244
rect 110934 -29300 110988 -29244
rect 111044 -29300 111098 -29244
rect 111154 -29300 111208 -29244
rect 111264 -29300 111318 -29244
rect 111374 -29300 111428 -29244
rect 111484 -29300 111580 -29244
rect 110594 -29354 111580 -29300
rect 110594 -29410 110768 -29354
rect 110824 -29410 110878 -29354
rect 110934 -29410 110988 -29354
rect 111044 -29410 111098 -29354
rect 111154 -29410 111208 -29354
rect 111264 -29410 111318 -29354
rect 111374 -29410 111428 -29354
rect 111484 -29410 111580 -29354
rect 110594 -29464 111580 -29410
rect 110594 -29520 110768 -29464
rect 110824 -29520 110878 -29464
rect 110934 -29520 110988 -29464
rect 111044 -29520 111098 -29464
rect 111154 -29520 111208 -29464
rect 111264 -29520 111318 -29464
rect 111374 -29520 111428 -29464
rect 111484 -29520 111580 -29464
rect 110594 -29574 111580 -29520
rect 110594 -29630 110768 -29574
rect 110824 -29630 110878 -29574
rect 110934 -29630 110988 -29574
rect 111044 -29630 111098 -29574
rect 111154 -29630 111208 -29574
rect 111264 -29630 111318 -29574
rect 111374 -29630 111428 -29574
rect 111484 -29630 111580 -29574
rect 110594 -29684 111580 -29630
rect 110594 -29740 110768 -29684
rect 110824 -29740 110878 -29684
rect 110934 -29740 110988 -29684
rect 111044 -29740 111098 -29684
rect 111154 -29740 111208 -29684
rect 111264 -29740 111318 -29684
rect 111374 -29740 111428 -29684
rect 111484 -29740 111580 -29684
rect 110594 -29825 111580 -29740
rect 113495 -30448 114395 -13813
rect 113495 -30504 113577 -30448
rect 113633 -30504 113687 -30448
rect 113743 -30504 113797 -30448
rect 113853 -30504 113907 -30448
rect 113963 -30504 114017 -30448
rect 114073 -30504 114127 -30448
rect 114183 -30504 114237 -30448
rect 114293 -30504 114395 -30448
rect 113495 -30558 114395 -30504
rect 113495 -30614 113577 -30558
rect 113633 -30614 113687 -30558
rect 113743 -30614 113797 -30558
rect 113853 -30614 113907 -30558
rect 113963 -30614 114017 -30558
rect 114073 -30614 114127 -30558
rect 114183 -30614 114237 -30558
rect 114293 -30614 114395 -30558
rect 113495 -30668 114395 -30614
rect 113495 -30724 113577 -30668
rect 113633 -30724 113687 -30668
rect 113743 -30724 113797 -30668
rect 113853 -30724 113907 -30668
rect 113963 -30724 114017 -30668
rect 114073 -30724 114127 -30668
rect 114183 -30724 114237 -30668
rect 114293 -30724 114395 -30668
rect 113495 -30778 114395 -30724
rect 113495 -30834 113577 -30778
rect 113633 -30834 113687 -30778
rect 113743 -30834 113797 -30778
rect 113853 -30834 113907 -30778
rect 113963 -30834 114017 -30778
rect 114073 -30834 114127 -30778
rect 114183 -30834 114237 -30778
rect 114293 -30834 114395 -30778
rect 113495 -30888 114395 -30834
rect 113495 -30944 113577 -30888
rect 113633 -30944 113687 -30888
rect 113743 -30944 113797 -30888
rect 113853 -30944 113907 -30888
rect 113963 -30944 114017 -30888
rect 114073 -30944 114127 -30888
rect 114183 -30944 114237 -30888
rect 114293 -30944 114395 -30888
rect 113495 -30998 114395 -30944
rect 113495 -31054 113577 -30998
rect 113633 -31054 113687 -30998
rect 113743 -31054 113797 -30998
rect 113853 -31054 113907 -30998
rect 113963 -31054 114017 -30998
rect 114073 -31054 114127 -30998
rect 114183 -31054 114237 -30998
rect 114293 -31054 114395 -30998
rect 113495 -31285 114395 -31054
rect 114563 18575 115463 18785
rect 114563 18519 114647 18575
rect 114703 18519 114757 18575
rect 114813 18519 114867 18575
rect 114923 18519 114977 18575
rect 115033 18519 115087 18575
rect 115143 18519 115197 18575
rect 115253 18519 115307 18575
rect 115363 18519 115463 18575
rect 114563 18465 115463 18519
rect 114563 18409 114647 18465
rect 114703 18409 114757 18465
rect 114813 18409 114867 18465
rect 114923 18409 114977 18465
rect 115033 18409 115087 18465
rect 115143 18409 115197 18465
rect 115253 18409 115307 18465
rect 115363 18409 115463 18465
rect 114563 18355 115463 18409
rect 114563 18299 114647 18355
rect 114703 18299 114757 18355
rect 114813 18299 114867 18355
rect 114923 18299 114977 18355
rect 115033 18299 115087 18355
rect 115143 18299 115197 18355
rect 115253 18299 115307 18355
rect 115363 18299 115463 18355
rect 114563 18245 115463 18299
rect 114563 18189 114647 18245
rect 114703 18189 114757 18245
rect 114813 18189 114867 18245
rect 114923 18189 114977 18245
rect 115033 18189 115087 18245
rect 115143 18189 115197 18245
rect 115253 18189 115307 18245
rect 115363 18189 115463 18245
rect 114563 18135 115463 18189
rect 114563 18079 114647 18135
rect 114703 18079 114757 18135
rect 114813 18079 114867 18135
rect 114923 18079 114977 18135
rect 115033 18079 115087 18135
rect 115143 18079 115197 18135
rect 115253 18079 115307 18135
rect 115363 18079 115463 18135
rect 114563 18025 115463 18079
rect 114563 17969 114647 18025
rect 114703 17969 114757 18025
rect 114813 17969 114867 18025
rect 114923 17969 114977 18025
rect 115033 17969 115087 18025
rect 115143 17969 115197 18025
rect 115253 17969 115307 18025
rect 115363 17969 115463 18025
rect 114563 10013 115463 17969
rect 116770 10013 116826 10015
rect 114563 10005 116888 10013
rect 114563 9949 116770 10005
rect 116826 9949 116888 10005
rect 114563 9895 116888 9949
rect 114563 9839 116770 9895
rect 116826 9839 116888 9895
rect 114563 9785 116888 9839
rect 114563 9729 116770 9785
rect 116826 9729 116888 9785
rect 114563 9675 116888 9729
rect 114563 9619 116770 9675
rect 116826 9619 116888 9675
rect 114563 9565 116888 9619
rect 114563 9509 116770 9565
rect 116826 9509 116888 9565
rect 114563 9455 116888 9509
rect 114563 9399 116770 9455
rect 116826 9399 116888 9455
rect 114563 9362 116888 9399
rect 114563 8395 115463 9362
rect 116188 8701 116402 9214
rect 116723 8430 116888 8438
rect 116723 8395 116770 8430
rect 114563 8374 116770 8395
rect 116826 8395 116888 8430
rect 116826 8374 116889 8395
rect 114563 8320 116889 8374
rect 114563 8264 116770 8320
rect 116826 8264 116889 8320
rect 114563 8210 116889 8264
rect 129873 8213 130140 8214
rect 114563 8154 116770 8210
rect 116826 8154 116889 8210
rect 129301 8157 130140 8213
rect 114563 8100 116889 8154
rect 114563 8044 116770 8100
rect 116826 8044 116889 8100
rect 114563 7990 116889 8044
rect 114563 7934 116770 7990
rect 116826 7934 116889 7990
rect 114563 7880 116889 7934
rect 114563 7824 116770 7880
rect 116826 7824 116889 7880
rect 114563 7787 116889 7824
rect 129237 7830 129427 7872
rect 114563 6885 115463 7787
rect 129237 7774 129243 7830
rect 129299 7774 129353 7830
rect 129409 7774 129427 7830
rect 129237 7740 129427 7774
rect 116723 6920 116888 6928
rect 116723 6885 116770 6920
rect 114563 6864 116770 6885
rect 116826 6864 116888 6920
rect 114563 6810 116888 6864
rect 114563 6754 116770 6810
rect 116826 6754 116888 6810
rect 114563 6700 116888 6754
rect 114563 6644 116770 6700
rect 116826 6644 116888 6700
rect 114563 6590 116888 6644
rect 114563 6534 116770 6590
rect 116826 6534 116888 6590
rect 114563 6480 116888 6534
rect 114563 6424 116770 6480
rect 116826 6424 116888 6480
rect 114563 6370 116888 6424
rect 114563 6314 116770 6370
rect 116826 6314 116888 6370
rect 114563 6277 116888 6314
rect 114563 5465 115463 6277
rect 116723 5500 116888 5508
rect 116723 5465 116770 5500
rect 114563 5444 116770 5465
rect 116826 5465 116888 5500
rect 116826 5444 116899 5465
rect 114563 5390 116899 5444
rect 114563 5334 116770 5390
rect 116826 5334 116899 5390
rect 114563 5280 116899 5334
rect 114563 5224 116770 5280
rect 116826 5224 116899 5280
rect 129242 5333 129478 5366
rect 129242 5277 129259 5333
rect 129315 5277 129369 5333
rect 129425 5277 129478 5333
rect 129242 5241 129478 5277
rect 114563 5170 116899 5224
rect 114563 5114 116770 5170
rect 116826 5114 116899 5170
rect 114563 5060 116899 5114
rect 114563 5004 116770 5060
rect 116826 5004 116899 5060
rect 114563 4950 116899 5004
rect 114563 4894 116770 4950
rect 116826 4894 116899 4950
rect 114563 4857 116899 4894
rect 114563 -1199 115463 4857
rect 128977 3904 129779 4024
rect 114563 -1255 114635 -1199
rect 114691 -1255 114745 -1199
rect 114801 -1255 114855 -1199
rect 114911 -1255 114965 -1199
rect 115021 -1255 115075 -1199
rect 115131 -1255 115185 -1199
rect 115241 -1255 115295 -1199
rect 115351 -1255 115463 -1199
rect 114563 -1309 115463 -1255
rect 114563 -1365 114635 -1309
rect 114691 -1365 114745 -1309
rect 114801 -1365 114855 -1309
rect 114911 -1365 114965 -1309
rect 115021 -1365 115075 -1309
rect 115131 -1365 115185 -1309
rect 115241 -1365 115295 -1309
rect 115351 -1365 115463 -1309
rect 114563 -1419 115463 -1365
rect 114563 -1475 114635 -1419
rect 114691 -1475 114745 -1419
rect 114801 -1475 114855 -1419
rect 114911 -1475 114965 -1419
rect 115021 -1475 115075 -1419
rect 115131 -1475 115185 -1419
rect 115241 -1475 115295 -1419
rect 115351 -1475 115463 -1419
rect 114563 -1529 115463 -1475
rect 114563 -1585 114635 -1529
rect 114691 -1585 114745 -1529
rect 114801 -1585 114855 -1529
rect 114911 -1585 114965 -1529
rect 115021 -1585 115075 -1529
rect 115131 -1585 115185 -1529
rect 115241 -1585 115295 -1529
rect 115351 -1585 115463 -1529
rect 114563 -1639 115463 -1585
rect 114563 -1695 114635 -1639
rect 114691 -1695 114745 -1639
rect 114801 -1695 114855 -1639
rect 114911 -1695 114965 -1639
rect 115021 -1695 115075 -1639
rect 115131 -1695 115185 -1639
rect 115241 -1695 115295 -1639
rect 115351 -1695 115463 -1639
rect 114563 -1749 115463 -1695
rect 114563 -1805 114635 -1749
rect 114691 -1805 114745 -1749
rect 114801 -1805 114855 -1749
rect 114911 -1805 114965 -1749
rect 115021 -1805 115075 -1749
rect 115131 -1805 115185 -1749
rect 115241 -1805 115295 -1749
rect 115351 -1805 115463 -1749
rect 114563 -5214 115463 -1805
rect 129549 1018 129779 3904
rect 129549 962 129566 1018
rect 129622 962 129676 1018
rect 129732 962 129779 1018
rect 129549 908 129779 962
rect 129549 852 129566 908
rect 129622 852 129676 908
rect 129732 852 129779 908
rect 129549 798 129779 852
rect 129549 742 129566 798
rect 129622 742 129676 798
rect 129732 742 129779 798
rect 129549 688 129779 742
rect 129549 632 129566 688
rect 129622 632 129676 688
rect 129732 632 129779 688
rect 129549 578 129779 632
rect 129549 522 129566 578
rect 129622 522 129676 578
rect 129732 522 129779 578
rect 129549 468 129779 522
rect 129549 412 129566 468
rect 129622 412 129676 468
rect 129732 412 129779 468
rect 129549 -4433 129779 412
rect 129043 -4553 129779 -4433
rect 129873 1703 130140 8157
rect 129873 1647 129891 1703
rect 129947 1647 130001 1703
rect 130057 1647 130140 1703
rect 129873 1593 130140 1647
rect 129873 1537 129891 1593
rect 129947 1537 130001 1593
rect 130057 1537 130140 1593
rect 129873 1483 130140 1537
rect 129873 1427 129891 1483
rect 129947 1427 130001 1483
rect 130057 1427 130140 1483
rect 129873 1373 130140 1427
rect 129873 1317 129891 1373
rect 129947 1317 130001 1373
rect 130057 1317 130140 1373
rect 129873 1263 130140 1317
rect 129873 1207 129891 1263
rect 129947 1207 130001 1263
rect 130057 1207 130140 1263
rect 129873 1153 130140 1207
rect 129873 1097 129891 1153
rect 129947 1097 130001 1153
rect 130057 1097 130140 1153
rect 116615 -5214 116780 -5212
rect 114563 -5220 116780 -5214
rect 114563 -5276 116662 -5220
rect 116718 -5276 116780 -5220
rect 114563 -5330 116780 -5276
rect 114563 -5386 116662 -5330
rect 116718 -5386 116780 -5330
rect 114563 -5440 116780 -5386
rect 114563 -5496 116662 -5440
rect 116718 -5496 116780 -5440
rect 114563 -5550 116780 -5496
rect 114563 -5606 116662 -5550
rect 116718 -5606 116780 -5550
rect 114563 -5660 116780 -5606
rect 114563 -5716 116662 -5660
rect 116718 -5716 116780 -5660
rect 114563 -5770 116780 -5716
rect 114563 -5826 116662 -5770
rect 116718 -5826 116780 -5770
rect 114563 -5862 116780 -5826
rect 114563 -6604 115463 -5862
rect 116615 -5863 116780 -5862
rect 114563 -6607 116781 -6604
rect 114563 -6615 116784 -6607
rect 114563 -6671 116666 -6615
rect 116722 -6671 116784 -6615
rect 114563 -6725 116784 -6671
rect 114563 -6781 116666 -6725
rect 116722 -6781 116784 -6725
rect 114563 -6835 116784 -6781
rect 114563 -6891 116666 -6835
rect 116722 -6891 116784 -6835
rect 114563 -6945 116784 -6891
rect 114563 -7001 116666 -6945
rect 116722 -7001 116784 -6945
rect 114563 -7055 116784 -7001
rect 129873 -7036 130140 1097
rect 130214 7832 130481 7872
rect 130214 7776 130252 7832
rect 130308 7776 130362 7832
rect 130418 7776 130481 7832
rect 130214 2376 130481 7776
rect 130214 2320 130234 2376
rect 130290 2320 130344 2376
rect 130400 2320 130481 2376
rect 130214 2266 130481 2320
rect 130214 2210 130234 2266
rect 130290 2210 130344 2266
rect 130400 2210 130481 2266
rect 130214 2156 130481 2210
rect 130214 2100 130234 2156
rect 130290 2100 130344 2156
rect 130400 2100 130481 2156
rect 130214 2046 130481 2100
rect 130214 1990 130234 2046
rect 130290 1990 130344 2046
rect 130400 1990 130481 2046
rect 130214 1936 130481 1990
rect 130214 1880 130234 1936
rect 130290 1880 130344 1936
rect 130400 1880 130481 1936
rect 130214 1826 130481 1880
rect 130214 1770 130234 1826
rect 130290 1770 130344 1826
rect 130400 1770 130481 1826
rect 114563 -7111 116666 -7055
rect 116722 -7111 116784 -7055
rect 129169 -7092 130143 -7036
rect 114563 -7165 116784 -7111
rect 114563 -7221 116666 -7165
rect 116722 -7221 116784 -7165
rect 114563 -7252 116784 -7221
rect 114563 -8438 115463 -7252
rect 116619 -7258 116784 -7252
rect 130214 -7420 130481 1770
rect 129151 -7476 130481 -7420
rect 130214 -7477 130481 -7476
rect 130559 5338 130826 5366
rect 130559 5282 130585 5338
rect 130641 5282 130695 5338
rect 130751 5282 130826 5338
rect 130559 3119 130826 5282
rect 130559 3063 130581 3119
rect 130637 3063 130691 3119
rect 130747 3063 130826 3119
rect 130559 3009 130826 3063
rect 130559 2953 130581 3009
rect 130637 2953 130691 3009
rect 130747 2953 130826 3009
rect 130559 2899 130826 2953
rect 130559 2843 130581 2899
rect 130637 2843 130691 2899
rect 130747 2843 130826 2899
rect 130559 2789 130826 2843
rect 130559 2733 130581 2789
rect 130637 2733 130691 2789
rect 130747 2733 130826 2789
rect 130559 2679 130826 2733
rect 130559 2623 130581 2679
rect 130637 2623 130691 2679
rect 130747 2623 130826 2679
rect 130559 2569 130826 2623
rect 130559 2513 130581 2569
rect 130637 2513 130691 2569
rect 130747 2513 130826 2569
rect 114563 -8446 116782 -8438
rect 114563 -8502 116664 -8446
rect 116720 -8502 116782 -8446
rect 114563 -8556 116782 -8502
rect 114563 -8612 116664 -8556
rect 116720 -8612 116782 -8556
rect 114563 -8666 116782 -8612
rect 114563 -8722 116664 -8666
rect 116720 -8722 116782 -8666
rect 114563 -8776 116782 -8722
rect 114563 -8832 116664 -8776
rect 116720 -8832 116782 -8776
rect 114563 -8886 116782 -8832
rect 114563 -8942 116664 -8886
rect 116720 -8942 116782 -8886
rect 114563 -8996 116782 -8942
rect 114563 -9052 116664 -8996
rect 116720 -9052 116782 -8996
rect 114563 -9086 116782 -9052
rect 114563 -9757 115463 -9086
rect 116617 -9089 116782 -9086
rect 116618 -9757 116783 -9756
rect 114563 -9764 116785 -9757
rect 114563 -9820 116665 -9764
rect 116721 -9820 116785 -9764
rect 114563 -9874 116785 -9820
rect 114563 -9930 116665 -9874
rect 116721 -9930 116785 -9874
rect 130559 -9914 130826 2513
rect 114563 -9984 116785 -9930
rect 129100 -9973 130826 -9914
rect 129100 -9974 130753 -9973
rect 114563 -10040 116665 -9984
rect 116721 -10040 116785 -9984
rect 114563 -10094 116785 -10040
rect 114563 -10150 116665 -10094
rect 116721 -10150 116785 -10094
rect 114563 -10204 116785 -10150
rect 114563 -10260 116665 -10204
rect 116721 -10260 116785 -10204
rect 114563 -10314 116785 -10260
rect 114563 -10370 116665 -10314
rect 116721 -10370 116785 -10314
rect 114563 -10405 116785 -10370
rect 25861 -31670 25910 -31614
rect 25966 -31670 26020 -31614
rect 26076 -31670 26130 -31614
rect 26186 -31670 26240 -31614
rect 26296 -31670 26350 -31614
rect 26406 -31670 26460 -31614
rect 26516 -31670 26570 -31614
rect 26626 -31670 26761 -31614
rect 25861 -31724 26761 -31670
rect 25861 -31780 25910 -31724
rect 25966 -31780 26020 -31724
rect 26076 -31780 26130 -31724
rect 26186 -31780 26240 -31724
rect 26296 -31780 26350 -31724
rect 26406 -31780 26460 -31724
rect 26516 -31780 26570 -31724
rect 26626 -31780 26761 -31724
rect 25861 -31834 26761 -31780
rect 25861 -31890 25910 -31834
rect 25966 -31890 26020 -31834
rect 26076 -31890 26130 -31834
rect 26186 -31890 26240 -31834
rect 26296 -31890 26350 -31834
rect 26406 -31890 26460 -31834
rect 26516 -31890 26570 -31834
rect 26626 -31890 26761 -31834
rect 25861 -31944 26761 -31890
rect 25861 -32000 25910 -31944
rect 25966 -32000 26020 -31944
rect 26076 -32000 26130 -31944
rect 26186 -32000 26240 -31944
rect 26296 -32000 26350 -31944
rect 26406 -32000 26460 -31944
rect 26516 -32000 26570 -31944
rect 26626 -32000 26761 -31944
rect 25861 -32054 26761 -32000
rect 25861 -32110 25910 -32054
rect 25966 -32110 26020 -32054
rect 26076 -32110 26130 -32054
rect 26186 -32110 26240 -32054
rect 26296 -32110 26350 -32054
rect 26406 -32110 26460 -32054
rect 26516 -32110 26570 -32054
rect 26626 -32110 26761 -32054
rect 25861 -32164 26761 -32110
rect 25861 -32220 25910 -32164
rect 25966 -32220 26020 -32164
rect 26076 -32220 26130 -32164
rect 26186 -32220 26240 -32164
rect 26296 -32220 26350 -32164
rect 26406 -32220 26460 -32164
rect 26516 -32220 26570 -32164
rect 26626 -32220 26761 -32164
rect 25861 -32362 26761 -32220
rect 114563 -31659 115463 -10405
rect 116618 -10407 116783 -10405
rect 114563 -31715 114633 -31659
rect 114689 -31715 114743 -31659
rect 114799 -31715 114853 -31659
rect 114909 -31715 114963 -31659
rect 115019 -31715 115073 -31659
rect 115129 -31715 115183 -31659
rect 115239 -31715 115293 -31659
rect 115349 -31715 115463 -31659
rect 114563 -31769 115463 -31715
rect 114563 -31825 114633 -31769
rect 114689 -31825 114743 -31769
rect 114799 -31825 114853 -31769
rect 114909 -31825 114963 -31769
rect 115019 -31825 115073 -31769
rect 115129 -31825 115183 -31769
rect 115239 -31825 115293 -31769
rect 115349 -31825 115463 -31769
rect 114563 -31879 115463 -31825
rect 114563 -31935 114633 -31879
rect 114689 -31935 114743 -31879
rect 114799 -31935 114853 -31879
rect 114909 -31935 114963 -31879
rect 115019 -31935 115073 -31879
rect 115129 -31935 115183 -31879
rect 115239 -31935 115293 -31879
rect 115349 -31935 115463 -31879
rect 114563 -31989 115463 -31935
rect 114563 -32045 114633 -31989
rect 114689 -32045 114743 -31989
rect 114799 -32045 114853 -31989
rect 114909 -32045 114963 -31989
rect 115019 -32045 115073 -31989
rect 115129 -32045 115183 -31989
rect 115239 -32045 115293 -31989
rect 115349 -32045 115463 -31989
rect 114563 -32099 115463 -32045
rect 114563 -32155 114633 -32099
rect 114689 -32155 114743 -32099
rect 114799 -32155 114853 -32099
rect 114909 -32155 114963 -32099
rect 115019 -32155 115073 -32099
rect 115129 -32155 115183 -32099
rect 115239 -32155 115293 -32099
rect 115349 -32155 115463 -32099
rect 114563 -32209 115463 -32155
rect 114563 -32265 114633 -32209
rect 114689 -32265 114743 -32209
rect 114799 -32265 114853 -32209
rect 114909 -32265 114963 -32209
rect 115019 -32265 115073 -32209
rect 115129 -32265 115183 -32209
rect 115239 -32265 115293 -32209
rect 115349 -32265 115463 -32209
rect 114563 -32350 115463 -32265
<< via2 >>
rect -814 -16469 -758 -16413
rect -704 -16469 -648 -16413
rect -594 -16469 -538 -16413
rect -484 -16469 -428 -16413
rect -374 -16469 -318 -16413
rect -264 -16469 -208 -16413
rect -154 -16469 -98 -16413
rect -814 -16579 -758 -16523
rect -704 -16579 -648 -16523
rect -594 -16579 -538 -16523
rect -484 -16579 -428 -16523
rect -374 -16579 -318 -16523
rect -264 -16579 -208 -16523
rect -154 -16579 -98 -16523
rect -814 -16689 -758 -16633
rect -704 -16689 -648 -16633
rect -594 -16689 -538 -16633
rect -484 -16689 -428 -16633
rect -374 -16689 -318 -16633
rect -264 -16689 -208 -16633
rect -154 -16689 -98 -16633
rect -814 -16799 -758 -16743
rect -704 -16799 -648 -16743
rect -594 -16799 -538 -16743
rect -484 -16799 -428 -16743
rect -374 -16799 -318 -16743
rect -264 -16799 -208 -16743
rect -154 -16799 -98 -16743
rect -814 -16909 -758 -16853
rect -704 -16909 -648 -16853
rect -594 -16909 -538 -16853
rect -484 -16909 -428 -16853
rect -374 -16909 -318 -16853
rect -264 -16909 -208 -16853
rect -154 -16909 -98 -16853
rect -814 -17019 -758 -16963
rect -704 -17019 -648 -16963
rect -594 -17019 -538 -16963
rect -484 -17019 -428 -16963
rect -374 -17019 -318 -16963
rect -264 -17019 -208 -16963
rect -154 -17019 -98 -16963
rect -814 -17129 -758 -17073
rect -704 -17129 -648 -17073
rect -594 -17129 -538 -17073
rect -484 -17129 -428 -17073
rect -374 -17129 -318 -17073
rect -264 -17129 -208 -17073
rect -154 -17129 -98 -17073
rect 121 -17404 177 -17348
rect 231 -17404 287 -17348
rect 341 -17404 397 -17348
rect 451 -17404 507 -17348
rect 561 -17404 617 -17348
rect 671 -17404 727 -17348
rect 781 -17404 837 -17348
rect 121 -17514 177 -17458
rect 231 -17514 287 -17458
rect 341 -17514 397 -17458
rect 451 -17514 507 -17458
rect 561 -17514 617 -17458
rect 671 -17514 727 -17458
rect 781 -17514 837 -17458
rect 121 -17624 177 -17568
rect 231 -17624 287 -17568
rect 341 -17624 397 -17568
rect 451 -17624 507 -17568
rect 561 -17624 617 -17568
rect 671 -17624 727 -17568
rect 781 -17624 837 -17568
rect 121 -17734 177 -17678
rect 231 -17734 287 -17678
rect 341 -17734 397 -17678
rect 451 -17734 507 -17678
rect 561 -17734 617 -17678
rect 671 -17734 727 -17678
rect 781 -17734 837 -17678
rect 121 -17844 177 -17788
rect 231 -17844 287 -17788
rect 341 -17844 397 -17788
rect 451 -17844 507 -17788
rect 561 -17844 617 -17788
rect 671 -17844 727 -17788
rect 781 -17844 837 -17788
rect 121 -17954 177 -17898
rect 231 -17954 287 -17898
rect 341 -17954 397 -17898
rect 451 -17954 507 -17898
rect 561 -17954 617 -17898
rect 671 -17954 727 -17898
rect 781 -17954 837 -17898
rect 121 -18064 177 -18008
rect 231 -18064 287 -18008
rect 341 -18064 397 -18008
rect 451 -18064 507 -18008
rect 561 -18064 617 -18008
rect 671 -18064 727 -18008
rect 781 -18064 837 -18008
rect 4298 -714 4354 -658
rect 4408 -714 4464 -658
rect 4518 -714 4574 -658
rect 4628 -714 4684 -658
rect 4298 -824 4354 -768
rect 4408 -824 4464 -768
rect 4518 -824 4574 -768
rect 4628 -824 4684 -768
rect 10881 -1514 10937 -1458
rect 10991 -1514 11047 -1458
rect 11101 -1514 11157 -1458
rect 11211 -1514 11267 -1458
rect 11321 -1514 11377 -1458
rect 11431 -1514 11487 -1458
rect 11541 -1514 11597 -1458
rect 11670 -1514 11726 -1458
rect 11780 -1514 11836 -1458
rect 11890 -1514 11946 -1458
rect 12000 -1514 12056 -1458
rect 12110 -1514 12166 -1458
rect 12220 -1514 12276 -1458
rect 12330 -1514 12386 -1458
rect 10881 -1624 10937 -1568
rect 10991 -1624 11047 -1568
rect 11101 -1624 11157 -1568
rect 11211 -1624 11267 -1568
rect 11321 -1624 11377 -1568
rect 11431 -1624 11487 -1568
rect 11541 -1624 11597 -1568
rect 11670 -1624 11726 -1568
rect 11780 -1624 11836 -1568
rect 11890 -1624 11946 -1568
rect 12000 -1624 12056 -1568
rect 12110 -1624 12166 -1568
rect 12220 -1624 12276 -1568
rect 12330 -1624 12386 -1568
rect 10881 -1734 10937 -1678
rect 10991 -1734 11047 -1678
rect 11101 -1734 11157 -1678
rect 11211 -1734 11267 -1678
rect 11321 -1734 11377 -1678
rect 11431 -1734 11487 -1678
rect 11541 -1734 11597 -1678
rect 11670 -1734 11726 -1678
rect 11780 -1734 11836 -1678
rect 11890 -1734 11946 -1678
rect 12000 -1734 12056 -1678
rect 12110 -1734 12166 -1678
rect 12220 -1734 12276 -1678
rect 12330 -1734 12386 -1678
rect 1236 -18337 1292 -18281
rect 1346 -18337 1402 -18281
rect 1456 -18337 1512 -18281
rect 1566 -18337 1622 -18281
rect 1676 -18337 1732 -18281
rect 1786 -18337 1842 -18281
rect 1896 -18337 1952 -18281
rect 1236 -18447 1292 -18391
rect 1346 -18447 1402 -18391
rect 1456 -18447 1512 -18391
rect 1566 -18447 1622 -18391
rect 1676 -18447 1732 -18391
rect 1786 -18447 1842 -18391
rect 1896 -18447 1952 -18391
rect 1236 -18557 1292 -18501
rect 1346 -18557 1402 -18501
rect 1456 -18557 1512 -18501
rect 1566 -18557 1622 -18501
rect 1676 -18557 1732 -18501
rect 1786 -18557 1842 -18501
rect 1896 -18557 1952 -18501
rect 1236 -18667 1292 -18611
rect 1346 -18667 1402 -18611
rect 1456 -18667 1512 -18611
rect 1566 -18667 1622 -18611
rect 1676 -18667 1732 -18611
rect 1786 -18667 1842 -18611
rect 1896 -18667 1952 -18611
rect 1236 -18777 1292 -18721
rect 1346 -18777 1402 -18721
rect 1456 -18777 1512 -18721
rect 1566 -18777 1622 -18721
rect 1676 -18777 1732 -18721
rect 1786 -18777 1842 -18721
rect 1896 -18777 1952 -18721
rect 1236 -18887 1292 -18831
rect 1346 -18887 1402 -18831
rect 1456 -18887 1512 -18831
rect 1566 -18887 1622 -18831
rect 1676 -18887 1732 -18831
rect 1786 -18887 1842 -18831
rect 1896 -18887 1952 -18831
rect 1236 -18997 1292 -18941
rect 1346 -18997 1402 -18941
rect 1456 -18997 1512 -18941
rect 1566 -18997 1622 -18941
rect 1676 -18997 1732 -18941
rect 1786 -18997 1842 -18941
rect 1896 -18997 1952 -18941
rect 21746 -16495 21802 -16439
rect 21856 -16495 21912 -16439
rect 21966 -16495 22022 -16439
rect 22076 -16495 22132 -16439
rect 22186 -16495 22242 -16439
rect 22296 -16495 22352 -16439
rect 22406 -16495 22462 -16439
rect 21746 -16605 21802 -16549
rect 21856 -16605 21912 -16549
rect 21966 -16605 22022 -16549
rect 22076 -16605 22132 -16549
rect 22186 -16605 22242 -16549
rect 22296 -16605 22352 -16549
rect 22406 -16605 22462 -16549
rect 21746 -16715 21802 -16659
rect 21856 -16715 21912 -16659
rect 21966 -16715 22022 -16659
rect 22076 -16715 22132 -16659
rect 22186 -16715 22242 -16659
rect 22296 -16715 22352 -16659
rect 22406 -16715 22462 -16659
rect 21746 -16825 21802 -16769
rect 21856 -16825 21912 -16769
rect 21966 -16825 22022 -16769
rect 22076 -16825 22132 -16769
rect 22186 -16825 22242 -16769
rect 22296 -16825 22352 -16769
rect 22406 -16825 22462 -16769
rect 21746 -16935 21802 -16879
rect 21856 -16935 21912 -16879
rect 21966 -16935 22022 -16879
rect 22076 -16935 22132 -16879
rect 22186 -16935 22242 -16879
rect 22296 -16935 22352 -16879
rect 22406 -16935 22462 -16879
rect 21746 -17045 21802 -16989
rect 21856 -17045 21912 -16989
rect 21966 -17045 22022 -16989
rect 22076 -17045 22132 -16989
rect 22186 -17045 22242 -16989
rect 22296 -17045 22352 -16989
rect 22406 -17045 22462 -16989
rect 21746 -17155 21802 -17099
rect 21856 -17155 21912 -17099
rect 21966 -17155 22022 -17099
rect 22076 -17155 22132 -17099
rect 22186 -17155 22242 -17099
rect 22296 -17155 22352 -17099
rect 22406 -17155 22462 -17099
rect 15724 -17414 15780 -17358
rect 15834 -17414 15890 -17358
rect 15944 -17414 16000 -17358
rect 16054 -17414 16110 -17358
rect 16164 -17414 16220 -17358
rect 16274 -17414 16330 -17358
rect 16384 -17414 16440 -17358
rect 15724 -17524 15780 -17468
rect 15834 -17524 15890 -17468
rect 15944 -17524 16000 -17468
rect 16054 -17524 16110 -17468
rect 16164 -17524 16220 -17468
rect 16274 -17524 16330 -17468
rect 16384 -17524 16440 -17468
rect 15724 -17634 15780 -17578
rect 15834 -17634 15890 -17578
rect 15944 -17634 16000 -17578
rect 16054 -17634 16110 -17578
rect 16164 -17634 16220 -17578
rect 16274 -17634 16330 -17578
rect 16384 -17634 16440 -17578
rect 15724 -17744 15780 -17688
rect 15834 -17744 15890 -17688
rect 15944 -17744 16000 -17688
rect 16054 -17744 16110 -17688
rect 16164 -17744 16220 -17688
rect 16274 -17744 16330 -17688
rect 16384 -17744 16440 -17688
rect 15724 -17854 15780 -17798
rect 15834 -17854 15890 -17798
rect 15944 -17854 16000 -17798
rect 16054 -17854 16110 -17798
rect 16164 -17854 16220 -17798
rect 16274 -17854 16330 -17798
rect 16384 -17854 16440 -17798
rect 15724 -17964 15780 -17908
rect 15834 -17964 15890 -17908
rect 15944 -17964 16000 -17908
rect 16054 -17964 16110 -17908
rect 16164 -17964 16220 -17908
rect 16274 -17964 16330 -17908
rect 16384 -17964 16440 -17908
rect 15724 -18074 15780 -18018
rect 15834 -18074 15890 -18018
rect 15944 -18074 16000 -18018
rect 16054 -18074 16110 -18018
rect 16164 -18074 16220 -18018
rect 16274 -18074 16330 -18018
rect 16384 -18074 16440 -18018
rect 13167 -19927 13223 -19871
rect 13277 -19927 13333 -19871
rect 13387 -19927 13443 -19871
rect 13497 -19927 13553 -19871
rect 13607 -19927 13663 -19871
rect 13717 -19927 13773 -19871
rect 13827 -19927 13883 -19871
rect 13167 -20037 13223 -19981
rect 13277 -20037 13333 -19981
rect 13387 -20037 13443 -19981
rect 13497 -20037 13553 -19981
rect 13607 -20037 13663 -19981
rect 13717 -20037 13773 -19981
rect 13827 -20037 13883 -19981
rect 13167 -20147 13223 -20091
rect 13277 -20147 13333 -20091
rect 13387 -20147 13443 -20091
rect 13497 -20147 13553 -20091
rect 13607 -20147 13663 -20091
rect 13717 -20147 13773 -20091
rect 13827 -20147 13883 -20091
rect 13167 -20257 13223 -20201
rect 13277 -20257 13333 -20201
rect 13387 -20257 13443 -20201
rect 13497 -20257 13553 -20201
rect 13607 -20257 13663 -20201
rect 13717 -20257 13773 -20201
rect 13827 -20257 13883 -20201
rect 13167 -20367 13223 -20311
rect 13277 -20367 13333 -20311
rect 13387 -20367 13443 -20311
rect 13497 -20367 13553 -20311
rect 13607 -20367 13663 -20311
rect 13717 -20367 13773 -20311
rect 13827 -20367 13883 -20311
rect 13167 -20477 13223 -20421
rect 13277 -20477 13333 -20421
rect 13387 -20477 13443 -20421
rect 13497 -20477 13553 -20421
rect 13607 -20477 13663 -20421
rect 13717 -20477 13773 -20421
rect 13827 -20477 13883 -20421
rect 13167 -20587 13223 -20531
rect 13277 -20587 13333 -20531
rect 13387 -20587 13443 -20531
rect 13497 -20587 13553 -20531
rect 13607 -20587 13663 -20531
rect 13717 -20587 13773 -20531
rect 13827 -20587 13883 -20531
rect 12283 -20813 12339 -20757
rect 12393 -20813 12449 -20757
rect 12503 -20813 12559 -20757
rect 12613 -20813 12669 -20757
rect 12723 -20813 12779 -20757
rect 12833 -20813 12889 -20757
rect 12943 -20813 12999 -20757
rect 12283 -20923 12339 -20867
rect 12393 -20923 12449 -20867
rect 12503 -20923 12559 -20867
rect 12613 -20923 12669 -20867
rect 12723 -20923 12779 -20867
rect 12833 -20923 12889 -20867
rect 12943 -20923 12999 -20867
rect 12283 -21033 12339 -20977
rect 12393 -21033 12449 -20977
rect 12503 -21033 12559 -20977
rect 12613 -21033 12669 -20977
rect 12723 -21033 12779 -20977
rect 12833 -21033 12889 -20977
rect 12943 -21033 12999 -20977
rect 12283 -21143 12339 -21087
rect 12393 -21143 12449 -21087
rect 12503 -21143 12559 -21087
rect 12613 -21143 12669 -21087
rect 12723 -21143 12779 -21087
rect 12833 -21143 12889 -21087
rect 12943 -21143 12999 -21087
rect 12283 -21253 12339 -21197
rect 12393 -21253 12449 -21197
rect 12503 -21253 12559 -21197
rect 12613 -21253 12669 -21197
rect 12723 -21253 12779 -21197
rect 12833 -21253 12889 -21197
rect 12943 -21253 12999 -21197
rect 12283 -21363 12339 -21307
rect 12393 -21363 12449 -21307
rect 12503 -21363 12559 -21307
rect 12613 -21363 12669 -21307
rect 12723 -21363 12779 -21307
rect 12833 -21363 12889 -21307
rect 12943 -21363 12999 -21307
rect 12283 -21473 12339 -21417
rect 12393 -21473 12449 -21417
rect 12503 -21473 12559 -21417
rect 12613 -21473 12669 -21417
rect 12723 -21473 12779 -21417
rect 12833 -21473 12889 -21417
rect 12943 -21473 12999 -21417
rect 19494 -19928 19550 -19872
rect 19604 -19928 19660 -19872
rect 19714 -19928 19770 -19872
rect 19824 -19928 19880 -19872
rect 19934 -19928 19990 -19872
rect 20044 -19928 20100 -19872
rect 20154 -19928 20210 -19872
rect 19494 -20038 19550 -19982
rect 19604 -20038 19660 -19982
rect 19714 -20038 19770 -19982
rect 19824 -20038 19880 -19982
rect 19934 -20038 19990 -19982
rect 20044 -20038 20100 -19982
rect 20154 -20038 20210 -19982
rect 19494 -20148 19550 -20092
rect 19604 -20148 19660 -20092
rect 19714 -20148 19770 -20092
rect 19824 -20148 19880 -20092
rect 19934 -20148 19990 -20092
rect 20044 -20148 20100 -20092
rect 20154 -20148 20210 -20092
rect 19494 -20258 19550 -20202
rect 19604 -20258 19660 -20202
rect 19714 -20258 19770 -20202
rect 19824 -20258 19880 -20202
rect 19934 -20258 19990 -20202
rect 20044 -20258 20100 -20202
rect 20154 -20258 20210 -20202
rect 19494 -20368 19550 -20312
rect 19604 -20368 19660 -20312
rect 19714 -20368 19770 -20312
rect 19824 -20368 19880 -20312
rect 19934 -20368 19990 -20312
rect 20044 -20368 20100 -20312
rect 20154 -20368 20210 -20312
rect 19494 -20478 19550 -20422
rect 19604 -20478 19660 -20422
rect 19714 -20478 19770 -20422
rect 19824 -20478 19880 -20422
rect 19934 -20478 19990 -20422
rect 20044 -20478 20100 -20422
rect 20154 -20478 20210 -20422
rect 19494 -20588 19550 -20532
rect 19604 -20588 19660 -20532
rect 19714 -20588 19770 -20532
rect 19824 -20588 19880 -20532
rect 19934 -20588 19990 -20532
rect 20044 -20588 20100 -20532
rect 20154 -20588 20210 -20532
rect 18599 -20808 18655 -20752
rect 18709 -20808 18765 -20752
rect 18819 -20808 18875 -20752
rect 18929 -20808 18985 -20752
rect 19039 -20808 19095 -20752
rect 19149 -20808 19205 -20752
rect 19259 -20808 19315 -20752
rect 18599 -20918 18655 -20862
rect 18709 -20918 18765 -20862
rect 18819 -20918 18875 -20862
rect 18929 -20918 18985 -20862
rect 19039 -20918 19095 -20862
rect 19149 -20918 19205 -20862
rect 19259 -20918 19315 -20862
rect 18599 -21028 18655 -20972
rect 18709 -21028 18765 -20972
rect 18819 -21028 18875 -20972
rect 18929 -21028 18985 -20972
rect 19039 -21028 19095 -20972
rect 19149 -21028 19205 -20972
rect 19259 -21028 19315 -20972
rect 18599 -21138 18655 -21082
rect 18709 -21138 18765 -21082
rect 18819 -21138 18875 -21082
rect 18929 -21138 18985 -21082
rect 19039 -21138 19095 -21082
rect 19149 -21138 19205 -21082
rect 19259 -21138 19315 -21082
rect 18599 -21248 18655 -21192
rect 18709 -21248 18765 -21192
rect 18819 -21248 18875 -21192
rect 18929 -21248 18985 -21192
rect 19039 -21248 19095 -21192
rect 19149 -21248 19205 -21192
rect 19259 -21248 19315 -21192
rect 18599 -21358 18655 -21302
rect 18709 -21358 18765 -21302
rect 18819 -21358 18875 -21302
rect 18929 -21358 18985 -21302
rect 19039 -21358 19095 -21302
rect 19149 -21358 19205 -21302
rect 19259 -21358 19315 -21302
rect 18599 -21468 18655 -21412
rect 18709 -21468 18765 -21412
rect 18819 -21468 18875 -21412
rect 18929 -21468 18985 -21412
rect 19039 -21468 19095 -21412
rect 19149 -21468 19205 -21412
rect 19259 -21468 19315 -21412
rect 24679 -13652 24735 -13596
rect 24789 -13652 24845 -13596
rect 24899 -13652 24955 -13596
rect 25009 -13652 25065 -13596
rect 25119 -13652 25175 -13596
rect 25229 -13652 25285 -13596
rect 25339 -13652 25395 -13596
rect 24679 -13762 24735 -13706
rect 24789 -13762 24845 -13706
rect 24899 -13762 24955 -13706
rect 25009 -13762 25065 -13706
rect 25119 -13762 25175 -13706
rect 25229 -13762 25285 -13706
rect 25339 -13762 25395 -13706
rect 24679 -13872 24735 -13816
rect 24789 -13872 24845 -13816
rect 24899 -13872 24955 -13816
rect 25009 -13872 25065 -13816
rect 25119 -13872 25175 -13816
rect 25229 -13872 25285 -13816
rect 25339 -13872 25395 -13816
rect 22902 -17510 22958 -17454
rect 23012 -17510 23068 -17454
rect 23122 -17510 23178 -17454
rect 23232 -17510 23288 -17454
rect 23387 -17506 23443 -17450
rect 23497 -17506 23553 -17450
rect 23607 -17506 23663 -17450
rect 23717 -17506 23773 -17450
rect 22902 -17620 22958 -17564
rect 23012 -17620 23068 -17564
rect 23122 -17620 23178 -17564
rect 23232 -17620 23288 -17564
rect 23387 -17616 23443 -17560
rect 23497 -17616 23553 -17560
rect 23607 -17616 23663 -17560
rect 23717 -17616 23773 -17560
rect 22902 -17730 22958 -17674
rect 23012 -17730 23068 -17674
rect 23122 -17730 23178 -17674
rect 23232 -17730 23288 -17674
rect 23387 -17726 23443 -17670
rect 23497 -17726 23553 -17670
rect 23607 -17726 23663 -17670
rect 23717 -17726 23773 -17670
rect 22902 -17840 22958 -17784
rect 23012 -17840 23068 -17784
rect 23122 -17840 23178 -17784
rect 23232 -17840 23288 -17784
rect 23387 -17836 23443 -17780
rect 23497 -17836 23553 -17780
rect 23607 -17836 23663 -17780
rect 23717 -17836 23773 -17780
rect 112156 17166 112212 17222
rect 112266 17166 112322 17222
rect 112376 17166 112432 17222
rect 112486 17166 112542 17222
rect 112596 17166 112652 17222
rect 112706 17166 112762 17222
rect 112816 17166 112872 17222
rect 112156 17056 112212 17112
rect 112266 17056 112322 17112
rect 112376 17056 112432 17112
rect 112486 17056 112542 17112
rect 112596 17056 112652 17112
rect 112706 17056 112762 17112
rect 112816 17056 112872 17112
rect 112156 16946 112212 17002
rect 112266 16946 112322 17002
rect 112376 16946 112432 17002
rect 112486 16946 112542 17002
rect 112596 16946 112652 17002
rect 112706 16946 112762 17002
rect 112816 16946 112872 17002
rect 112156 16836 112212 16892
rect 112266 16836 112322 16892
rect 112376 16836 112432 16892
rect 112486 16836 112542 16892
rect 112596 16836 112652 16892
rect 112706 16836 112762 16892
rect 112816 16836 112872 16892
rect 112156 16726 112212 16782
rect 112266 16726 112322 16782
rect 112376 16726 112432 16782
rect 112486 16726 112542 16782
rect 112596 16726 112652 16782
rect 112706 16726 112762 16782
rect 112816 16726 112872 16782
rect 112156 16616 112212 16672
rect 112266 16616 112322 16672
rect 112376 16616 112432 16672
rect 112486 16616 112542 16672
rect 112596 16616 112652 16672
rect 112706 16616 112762 16672
rect 112816 16616 112872 16672
rect 112156 16506 112212 16562
rect 112266 16506 112322 16562
rect 112376 16506 112432 16562
rect 112486 16506 112542 16562
rect 112596 16506 112652 16562
rect 112706 16506 112762 16562
rect 112816 16506 112872 16562
rect 27330 10609 27386 10665
rect 27440 10609 27496 10665
rect 27550 10609 27606 10665
rect 27660 10609 27716 10665
rect 27330 10499 27386 10555
rect 27440 10499 27496 10555
rect 27550 10499 27606 10555
rect 27660 10499 27716 10555
rect 27330 10389 27386 10445
rect 27440 10389 27496 10445
rect 27550 10389 27606 10445
rect 27660 10389 27716 10445
rect 27330 10279 27386 10335
rect 27440 10279 27496 10335
rect 27550 10279 27606 10335
rect 27660 10279 27716 10335
rect 27330 10169 27386 10225
rect 27440 10169 27496 10225
rect 27550 10169 27606 10225
rect 27660 10169 27716 10225
rect 27330 10059 27386 10115
rect 27440 10059 27496 10115
rect 27550 10059 27606 10115
rect 27660 10059 27716 10115
rect 27330 9949 27386 10005
rect 27440 9949 27496 10005
rect 27550 9949 27606 10005
rect 27660 9949 27716 10005
rect 27330 9839 27386 9895
rect 27440 9839 27496 9895
rect 27550 9839 27606 9895
rect 27660 9839 27716 9895
rect 25883 -4203 25939 -4147
rect 25993 -4203 26049 -4147
rect 26103 -4203 26159 -4147
rect 26213 -4203 26269 -4147
rect 26323 -4203 26379 -4147
rect 26470 -4202 26526 -4146
rect 26580 -4202 26636 -4146
rect 26690 -4202 26746 -4146
rect 25883 -4313 25939 -4257
rect 25993 -4313 26049 -4257
rect 26103 -4313 26159 -4257
rect 26213 -4313 26269 -4257
rect 26323 -4313 26379 -4257
rect 26470 -4312 26526 -4256
rect 26580 -4312 26636 -4256
rect 26690 -4312 26746 -4256
rect 25904 -14476 25960 -14420
rect 26014 -14476 26070 -14420
rect 26124 -14476 26180 -14420
rect 26234 -14476 26290 -14420
rect 26344 -14476 26400 -14420
rect 26454 -14476 26510 -14420
rect 26564 -14476 26620 -14420
rect 25904 -14586 25960 -14530
rect 26014 -14586 26070 -14530
rect 26124 -14586 26180 -14530
rect 26234 -14586 26290 -14530
rect 26344 -14586 26400 -14530
rect 26454 -14586 26510 -14530
rect 26564 -14586 26620 -14530
rect 25904 -14696 25960 -14640
rect 26014 -14696 26070 -14640
rect 26124 -14696 26180 -14640
rect 26234 -14696 26290 -14640
rect 26344 -14696 26400 -14640
rect 26454 -14696 26510 -14640
rect 26564 -14696 26620 -14640
rect 43928 6194 43984 6250
rect 44038 6194 44094 6250
rect 44148 6194 44204 6250
rect 44258 6194 44314 6250
rect 44368 6194 44424 6250
rect 31032 6079 31088 6135
rect 31142 6079 31198 6135
rect 31252 6079 31308 6135
rect 31362 6079 31418 6135
rect 31472 6079 31528 6135
rect 31582 6079 31638 6135
rect 31692 6079 31748 6135
rect 31032 5969 31088 6025
rect 31142 5969 31198 6025
rect 31252 5969 31308 6025
rect 31362 5969 31418 6025
rect 31472 5969 31528 6025
rect 31582 5969 31638 6025
rect 31692 5969 31748 6025
rect 43928 6084 43984 6140
rect 44038 6084 44094 6140
rect 44148 6084 44204 6140
rect 44258 6084 44314 6140
rect 44368 6084 44424 6140
rect 43928 5974 43984 6030
rect 44038 5974 44094 6030
rect 44148 5974 44204 6030
rect 44258 5974 44314 6030
rect 44368 5974 44424 6030
rect 46418 6253 46474 6309
rect 46528 6253 46584 6309
rect 46638 6253 46694 6309
rect 46748 6253 46804 6309
rect 46858 6253 46914 6309
rect 46421 6141 46477 6197
rect 46530 6142 46586 6198
rect 46638 6143 46694 6199
rect 46748 6143 46804 6199
rect 46858 6143 46914 6199
rect 46421 6035 46477 6091
rect 46527 6036 46583 6092
rect 46638 6033 46694 6089
rect 46748 6033 46804 6089
rect 46858 6033 46914 6089
rect 31032 5859 31088 5915
rect 31142 5859 31198 5915
rect 31252 5859 31308 5915
rect 31362 5859 31418 5915
rect 31472 5859 31528 5915
rect 31582 5859 31638 5915
rect 31692 5859 31748 5915
rect 31032 5749 31088 5805
rect 31142 5749 31198 5805
rect 31252 5749 31308 5805
rect 31362 5749 31418 5805
rect 31472 5749 31528 5805
rect 31582 5749 31638 5805
rect 31692 5749 31748 5805
rect 31032 5639 31088 5695
rect 31142 5639 31198 5695
rect 31252 5639 31308 5695
rect 31362 5639 31418 5695
rect 31472 5639 31528 5695
rect 31582 5639 31638 5695
rect 31692 5639 31748 5695
rect 31032 5529 31088 5585
rect 31142 5529 31198 5585
rect 31252 5529 31308 5585
rect 31362 5529 31418 5585
rect 31472 5529 31528 5585
rect 31582 5529 31638 5585
rect 31692 5529 31748 5585
rect 31032 5419 31088 5475
rect 31142 5419 31198 5475
rect 31252 5419 31308 5475
rect 31362 5419 31418 5475
rect 31472 5419 31528 5475
rect 31582 5419 31638 5475
rect 31692 5419 31748 5475
rect 27262 -7741 27318 -7685
rect 27372 -7741 27428 -7685
rect 27482 -7741 27538 -7685
rect 27592 -7741 27648 -7685
rect 27702 -7741 27758 -7685
rect 27262 -7851 27318 -7795
rect 27372 -7851 27428 -7795
rect 27482 -7851 27538 -7795
rect 27592 -7851 27648 -7795
rect 27702 -7851 27758 -7795
rect 27262 -7961 27318 -7905
rect 27372 -7961 27428 -7905
rect 27482 -7961 27538 -7905
rect 27592 -7961 27648 -7905
rect 27702 -7961 27758 -7905
rect 27262 -8071 27318 -8015
rect 27372 -8071 27428 -8015
rect 27482 -8071 27538 -8015
rect 27592 -8071 27648 -8015
rect 27702 -8071 27758 -8015
rect 30166 -4207 30222 -4151
rect 30276 -4207 30332 -4151
rect 30386 -4207 30442 -4151
rect 30496 -4207 30552 -4151
rect 30606 -4207 30662 -4151
rect 30716 -4207 30772 -4151
rect 30166 -4317 30222 -4261
rect 30276 -4317 30332 -4261
rect 30386 -4317 30442 -4261
rect 30496 -4317 30552 -4261
rect 30606 -4317 30662 -4261
rect 30716 -4317 30772 -4261
rect 110643 1690 110699 1746
rect 110753 1690 110809 1746
rect 110863 1690 110919 1746
rect 110973 1690 111029 1746
rect 111083 1690 111139 1746
rect 111193 1690 111249 1746
rect 111303 1690 111359 1746
rect 110643 1580 110699 1636
rect 110753 1580 110809 1636
rect 110863 1580 110919 1636
rect 110973 1580 111029 1636
rect 111083 1580 111139 1636
rect 111193 1580 111249 1636
rect 111303 1580 111359 1636
rect 110643 1470 110699 1526
rect 110753 1470 110809 1526
rect 110863 1470 110919 1526
rect 110973 1470 111029 1526
rect 111083 1470 111139 1526
rect 111193 1470 111249 1526
rect 111303 1470 111359 1526
rect 110643 1360 110699 1416
rect 110753 1360 110809 1416
rect 110863 1360 110919 1416
rect 110973 1360 111029 1416
rect 111083 1360 111139 1416
rect 111193 1360 111249 1416
rect 111303 1360 111359 1416
rect 110643 1250 110699 1306
rect 110753 1250 110809 1306
rect 110863 1250 110919 1306
rect 110973 1250 111029 1306
rect 111083 1250 111139 1306
rect 111193 1250 111249 1306
rect 111303 1250 111359 1306
rect 110643 1140 110699 1196
rect 110753 1140 110809 1196
rect 110863 1140 110919 1196
rect 110973 1140 111029 1196
rect 111083 1140 111139 1196
rect 111193 1140 111249 1196
rect 111303 1140 111359 1196
rect 110643 1030 110699 1086
rect 110753 1030 110809 1086
rect 110863 1030 110919 1086
rect 110973 1030 111029 1086
rect 111083 1030 111139 1086
rect 111193 1030 111249 1086
rect 111303 1030 111359 1086
rect 107221 -2479 107277 -2423
rect 107331 -2479 107387 -2423
rect 107441 -2479 107497 -2423
rect 107551 -2479 107607 -2423
rect 107661 -2479 107717 -2423
rect 107771 -2479 107827 -2423
rect 107881 -2479 107937 -2423
rect 107221 -2589 107277 -2533
rect 107331 -2589 107387 -2533
rect 107441 -2589 107497 -2533
rect 107551 -2589 107607 -2533
rect 107661 -2589 107717 -2533
rect 107771 -2589 107827 -2533
rect 107881 -2589 107937 -2533
rect 107221 -2699 107277 -2643
rect 107331 -2699 107387 -2643
rect 107441 -2699 107497 -2643
rect 107551 -2699 107607 -2643
rect 107661 -2699 107717 -2643
rect 107771 -2699 107827 -2643
rect 107881 -2699 107937 -2643
rect 107221 -2809 107277 -2753
rect 107331 -2809 107387 -2753
rect 107441 -2809 107497 -2753
rect 107551 -2809 107607 -2753
rect 107661 -2809 107717 -2753
rect 107771 -2809 107827 -2753
rect 107881 -2809 107937 -2753
rect 107221 -2919 107277 -2863
rect 107331 -2919 107387 -2863
rect 107441 -2919 107497 -2863
rect 107551 -2919 107607 -2863
rect 107661 -2919 107717 -2863
rect 107771 -2919 107827 -2863
rect 107881 -2919 107937 -2863
rect 107221 -3029 107277 -2973
rect 107331 -3029 107387 -2973
rect 107441 -3029 107497 -2973
rect 107551 -3029 107607 -2973
rect 107661 -3029 107717 -2973
rect 107771 -3029 107827 -2973
rect 107881 -3029 107937 -2973
rect 107221 -3139 107277 -3083
rect 107331 -3139 107387 -3083
rect 107441 -3139 107497 -3083
rect 107551 -3139 107607 -3083
rect 107661 -3139 107717 -3083
rect 107771 -3139 107827 -3083
rect 107881 -3139 107937 -3083
rect 31255 -11684 31311 -11628
rect 31365 -11684 31421 -11628
rect 31475 -11684 31531 -11628
rect 31585 -11684 31641 -11628
rect 31695 -11684 31751 -11628
rect 31255 -11794 31311 -11738
rect 31365 -11794 31421 -11738
rect 31475 -11794 31531 -11738
rect 31585 -11794 31641 -11738
rect 31695 -11794 31751 -11738
rect 31255 -11904 31311 -11848
rect 31365 -11904 31421 -11848
rect 31475 -11904 31531 -11848
rect 31585 -11904 31641 -11848
rect 31695 -11904 31751 -11848
rect 31255 -12014 31311 -11958
rect 31365 -12014 31421 -11958
rect 31475 -12014 31531 -11958
rect 31585 -12014 31641 -11958
rect 31695 -12014 31751 -11958
rect 31255 -12124 31311 -12068
rect 31365 -12124 31421 -12068
rect 31475 -12124 31531 -12068
rect 31585 -12124 31641 -12068
rect 31695 -12124 31751 -12068
rect 29533 -13720 29589 -13664
rect 29643 -13720 29699 -13664
rect 29753 -13720 29809 -13664
rect 29863 -13720 29919 -13664
rect 29973 -13720 30029 -13664
rect 30083 -13720 30139 -13664
rect 30193 -13712 30249 -13656
rect 30303 -13712 30359 -13656
rect 30413 -13712 30469 -13656
rect 29533 -13830 29589 -13774
rect 29643 -13830 29699 -13774
rect 29753 -13830 29809 -13774
rect 29863 -13830 29919 -13774
rect 29973 -13830 30029 -13774
rect 30083 -13830 30139 -13774
rect 30193 -13822 30249 -13766
rect 30303 -13822 30359 -13766
rect 30413 -13822 30469 -13766
rect 29852 -14525 29908 -14469
rect 29962 -14525 30018 -14469
rect 30072 -14525 30128 -14469
rect 30249 -14525 30305 -14469
rect 30359 -14525 30415 -14469
rect 30469 -14525 30525 -14469
rect 29852 -14635 29908 -14579
rect 29962 -14635 30018 -14579
rect 30072 -14635 30128 -14579
rect 30249 -14635 30305 -14579
rect 30359 -14635 30415 -14579
rect 30469 -14635 30525 -14579
rect 34121 -12438 34177 -12382
rect 34231 -12438 34287 -12382
rect 34341 -12438 34397 -12382
rect 34451 -12438 34507 -12382
rect 34121 -12548 34177 -12492
rect 34231 -12548 34287 -12492
rect 34341 -12548 34397 -12492
rect 34451 -12548 34507 -12492
rect 34121 -12658 34177 -12602
rect 34231 -12658 34287 -12602
rect 34341 -12658 34397 -12602
rect 34451 -12658 34507 -12602
rect 34121 -12768 34177 -12712
rect 34231 -12768 34287 -12712
rect 34341 -12768 34397 -12712
rect 34451 -12768 34507 -12712
rect 36056 -12443 36112 -12387
rect 36166 -12443 36222 -12387
rect 36276 -12443 36332 -12387
rect 36386 -12443 36442 -12387
rect 36496 -12443 36552 -12387
rect 36606 -12443 36662 -12387
rect 36716 -12443 36772 -12387
rect 36056 -12553 36112 -12497
rect 36166 -12553 36222 -12497
rect 36276 -12553 36332 -12497
rect 36386 -12553 36442 -12497
rect 36496 -12553 36552 -12497
rect 36606 -12553 36662 -12497
rect 36716 -12553 36772 -12497
rect 36056 -12663 36112 -12607
rect 36166 -12663 36222 -12607
rect 36276 -12663 36332 -12607
rect 36386 -12663 36442 -12607
rect 36496 -12663 36552 -12607
rect 36606 -12663 36662 -12607
rect 36716 -12663 36772 -12607
rect 36056 -12773 36112 -12717
rect 36166 -12773 36222 -12717
rect 36276 -12773 36332 -12717
rect 36386 -12773 36442 -12717
rect 36496 -12773 36552 -12717
rect 36606 -12773 36662 -12717
rect 36716 -12773 36772 -12717
rect 28388 -16618 28444 -16562
rect 28498 -16618 28554 -16562
rect 28608 -16618 28664 -16562
rect 28718 -16618 28774 -16562
rect 28873 -16614 28929 -16558
rect 28983 -16614 29039 -16558
rect 29093 -16614 29149 -16558
rect 29203 -16614 29259 -16558
rect 28388 -16728 28444 -16672
rect 28498 -16728 28554 -16672
rect 28608 -16728 28664 -16672
rect 28718 -16728 28774 -16672
rect 28873 -16724 28929 -16668
rect 28983 -16724 29039 -16668
rect 29093 -16724 29149 -16668
rect 29203 -16724 29259 -16668
rect 28388 -16838 28444 -16782
rect 28498 -16838 28554 -16782
rect 28608 -16838 28664 -16782
rect 28718 -16838 28774 -16782
rect 28873 -16834 28929 -16778
rect 28983 -16834 29039 -16778
rect 29093 -16834 29149 -16778
rect 29203 -16834 29259 -16778
rect 28388 -16948 28444 -16892
rect 28498 -16948 28554 -16892
rect 28608 -16948 28664 -16892
rect 28718 -16948 28774 -16892
rect 28873 -16944 28929 -16888
rect 28983 -16944 29039 -16888
rect 29093 -16944 29149 -16888
rect 29203 -16944 29259 -16888
rect 30894 -16612 30950 -16556
rect 31004 -16612 31060 -16556
rect 31114 -16612 31170 -16556
rect 31224 -16612 31280 -16556
rect 30894 -16722 30950 -16666
rect 31004 -16722 31060 -16666
rect 31114 -16722 31170 -16666
rect 31224 -16722 31280 -16666
rect 30894 -16832 30950 -16776
rect 31004 -16832 31060 -16776
rect 31114 -16832 31170 -16776
rect 31224 -16832 31280 -16776
rect 30894 -16942 30950 -16886
rect 31004 -16942 31060 -16886
rect 31114 -16942 31170 -16886
rect 31224 -16942 31280 -16886
rect 30249 -17512 30305 -17456
rect 30359 -17512 30415 -17456
rect 30469 -17512 30525 -17456
rect 30579 -17512 30635 -17456
rect 30249 -17622 30305 -17566
rect 30359 -17622 30415 -17566
rect 30469 -17622 30525 -17566
rect 30579 -17622 30635 -17566
rect 30249 -17732 30305 -17676
rect 30359 -17732 30415 -17676
rect 30469 -17732 30525 -17676
rect 30579 -17732 30635 -17676
rect 30249 -17842 30305 -17786
rect 30359 -17842 30415 -17786
rect 30469 -17842 30525 -17786
rect 30579 -17842 30635 -17786
rect 29788 -18391 29844 -18335
rect 29898 -18391 29954 -18335
rect 30008 -18391 30064 -18335
rect 30118 -18391 30174 -18335
rect 29788 -18501 29844 -18445
rect 29898 -18501 29954 -18445
rect 30008 -18501 30064 -18445
rect 30118 -18501 30174 -18445
rect 29782 -18629 29838 -18573
rect 29892 -18629 29948 -18573
rect 30002 -18629 30058 -18573
rect 30112 -18629 30168 -18573
rect 29782 -18739 29838 -18683
rect 29892 -18739 29948 -18683
rect 30002 -18739 30058 -18683
rect 30112 -18739 30168 -18683
rect 29782 -18849 29838 -18793
rect 29892 -18849 29948 -18793
rect 30002 -18849 30058 -18793
rect 30112 -18849 30168 -18793
rect 29782 -18959 29838 -18903
rect 29892 -18959 29948 -18903
rect 30002 -18959 30058 -18903
rect 30112 -18959 30168 -18903
rect 31488 -18729 31544 -18673
rect 31598 -18729 31654 -18673
rect 31708 -18729 31764 -18673
rect 31818 -18729 31874 -18673
rect 31488 -18839 31544 -18783
rect 31598 -18839 31654 -18783
rect 31708 -18839 31764 -18783
rect 31818 -18839 31874 -18783
rect 31488 -18949 31544 -18893
rect 31598 -18949 31654 -18893
rect 31708 -18949 31764 -18893
rect 31818 -18949 31874 -18893
rect 31488 -19059 31544 -19003
rect 31598 -19059 31654 -19003
rect 31708 -19059 31764 -19003
rect 31818 -19059 31874 -19003
rect 109095 -1058 109151 -1002
rect 109205 -1058 109261 -1002
rect 109315 -1058 109371 -1002
rect 109425 -1058 109481 -1002
rect 109535 -1058 109591 -1002
rect 109645 -1058 109701 -1002
rect 109755 -1058 109811 -1002
rect 109095 -1168 109151 -1112
rect 109205 -1168 109261 -1112
rect 109315 -1168 109371 -1112
rect 109425 -1168 109481 -1112
rect 109535 -1168 109591 -1112
rect 109645 -1168 109701 -1112
rect 109755 -1168 109811 -1112
rect 109095 -1278 109151 -1222
rect 109205 -1278 109261 -1222
rect 109315 -1278 109371 -1222
rect 109425 -1278 109481 -1222
rect 109535 -1278 109591 -1222
rect 109645 -1278 109701 -1222
rect 109755 -1278 109811 -1222
rect 109095 -1388 109151 -1332
rect 109205 -1388 109261 -1332
rect 109315 -1388 109371 -1332
rect 109425 -1388 109481 -1332
rect 109535 -1388 109591 -1332
rect 109645 -1388 109701 -1332
rect 109755 -1388 109811 -1332
rect 109095 -1498 109151 -1442
rect 109205 -1498 109261 -1442
rect 109315 -1498 109371 -1442
rect 109425 -1498 109481 -1442
rect 109535 -1498 109591 -1442
rect 109645 -1498 109701 -1442
rect 109755 -1498 109811 -1442
rect 109095 -1608 109151 -1552
rect 109205 -1608 109261 -1552
rect 109315 -1608 109371 -1552
rect 109425 -1608 109481 -1552
rect 109535 -1608 109591 -1552
rect 109645 -1608 109701 -1552
rect 109755 -1608 109811 -1552
rect 109095 -1718 109151 -1662
rect 109205 -1718 109261 -1662
rect 109315 -1718 109371 -1662
rect 109425 -1718 109481 -1662
rect 109535 -1718 109591 -1662
rect 109645 -1718 109701 -1662
rect 109755 -1718 109811 -1662
rect 109096 -14958 109152 -14902
rect 109206 -14958 109262 -14902
rect 109316 -14958 109372 -14902
rect 109426 -14958 109482 -14902
rect 109536 -14958 109592 -14902
rect 109646 -14958 109702 -14902
rect 109756 -14958 109812 -14902
rect 109096 -15068 109152 -15012
rect 109206 -15068 109262 -15012
rect 109316 -15068 109372 -15012
rect 109426 -15068 109482 -15012
rect 109536 -15068 109592 -15012
rect 109646 -15068 109702 -15012
rect 109756 -15068 109812 -15012
rect 109096 -15178 109152 -15122
rect 109206 -15178 109262 -15122
rect 109316 -15178 109372 -15122
rect 109426 -15178 109482 -15122
rect 109536 -15178 109592 -15122
rect 109646 -15178 109702 -15122
rect 109756 -15178 109812 -15122
rect 109096 -15288 109152 -15232
rect 109206 -15288 109262 -15232
rect 109316 -15288 109372 -15232
rect 109426 -15288 109482 -15232
rect 109536 -15288 109592 -15232
rect 109646 -15288 109702 -15232
rect 109756 -15288 109812 -15232
rect 109096 -15398 109152 -15342
rect 109206 -15398 109262 -15342
rect 109316 -15398 109372 -15342
rect 109426 -15398 109482 -15342
rect 109536 -15398 109592 -15342
rect 109646 -15398 109702 -15342
rect 109756 -15398 109812 -15342
rect 109096 -15508 109152 -15452
rect 109206 -15508 109262 -15452
rect 109316 -15508 109372 -15452
rect 109426 -15508 109482 -15452
rect 109536 -15508 109592 -15452
rect 109646 -15508 109702 -15452
rect 109756 -15508 109812 -15452
rect 109096 -15618 109152 -15562
rect 109206 -15618 109262 -15562
rect 109316 -15618 109372 -15562
rect 109426 -15618 109482 -15562
rect 109536 -15618 109592 -15562
rect 109646 -15618 109702 -15562
rect 109756 -15618 109812 -15562
rect 107210 -16327 107266 -16271
rect 107320 -16327 107376 -16271
rect 107430 -16327 107486 -16271
rect 107540 -16327 107596 -16271
rect 107650 -16327 107706 -16271
rect 107760 -16327 107816 -16271
rect 107870 -16327 107926 -16271
rect 107210 -16437 107266 -16381
rect 107320 -16437 107376 -16381
rect 107430 -16437 107486 -16381
rect 107540 -16437 107596 -16381
rect 107650 -16437 107706 -16381
rect 107760 -16437 107816 -16381
rect 107870 -16437 107926 -16381
rect 107210 -16547 107266 -16491
rect 107320 -16547 107376 -16491
rect 107430 -16547 107486 -16491
rect 107540 -16547 107596 -16491
rect 107650 -16547 107706 -16491
rect 107760 -16547 107816 -16491
rect 107870 -16547 107926 -16491
rect 107210 -16657 107266 -16601
rect 107320 -16657 107376 -16601
rect 107430 -16657 107486 -16601
rect 107540 -16657 107596 -16601
rect 107650 -16657 107706 -16601
rect 107760 -16657 107816 -16601
rect 107870 -16657 107926 -16601
rect 107210 -16767 107266 -16711
rect 107320 -16767 107376 -16711
rect 107430 -16767 107486 -16711
rect 107540 -16767 107596 -16711
rect 107650 -16767 107706 -16711
rect 107760 -16767 107816 -16711
rect 107870 -16767 107926 -16711
rect 107210 -16877 107266 -16821
rect 107320 -16877 107376 -16821
rect 107430 -16877 107486 -16821
rect 107540 -16877 107596 -16821
rect 107650 -16877 107706 -16821
rect 107760 -16877 107816 -16821
rect 107870 -16877 107926 -16821
rect 107210 -16987 107266 -16931
rect 107320 -16987 107376 -16931
rect 107430 -16987 107486 -16931
rect 107540 -16987 107596 -16931
rect 107650 -16987 107706 -16931
rect 107760 -16987 107816 -16931
rect 107870 -16987 107926 -16931
rect 34132 -18781 34188 -18725
rect 34242 -18781 34298 -18725
rect 34352 -18781 34408 -18725
rect 34462 -18781 34518 -18725
rect 34132 -18891 34188 -18835
rect 34242 -18891 34298 -18835
rect 34352 -18891 34408 -18835
rect 34462 -18891 34518 -18835
rect 34132 -19001 34188 -18945
rect 34242 -19001 34298 -18945
rect 34352 -19001 34408 -18945
rect 34462 -19001 34518 -18945
rect 34132 -19111 34188 -19055
rect 34242 -19111 34298 -19055
rect 34352 -19111 34408 -19055
rect 34462 -19111 34518 -19055
rect 94359 -18731 94415 -18675
rect 94469 -18731 94525 -18675
rect 94579 -18731 94635 -18675
rect 94689 -18731 94745 -18675
rect 94359 -18841 94415 -18785
rect 94469 -18841 94525 -18785
rect 94579 -18841 94635 -18785
rect 94689 -18841 94745 -18785
rect 94359 -18951 94415 -18895
rect 94469 -18951 94525 -18895
rect 94579 -18951 94635 -18895
rect 94689 -18951 94745 -18895
rect 94359 -19061 94415 -19005
rect 94469 -19061 94525 -19005
rect 94579 -19061 94635 -19005
rect 94689 -19061 94745 -19005
rect 94359 -19171 94415 -19115
rect 94469 -19171 94525 -19115
rect 94579 -19171 94635 -19115
rect 94689 -19171 94745 -19115
rect 94359 -19281 94415 -19225
rect 94469 -19281 94525 -19225
rect 94579 -19281 94635 -19225
rect 94689 -19281 94745 -19225
rect 94359 -19391 94415 -19335
rect 94469 -19391 94525 -19335
rect 94579 -19391 94635 -19335
rect 94689 -19391 94745 -19335
rect 28803 -20007 28859 -19951
rect 28913 -20007 28969 -19951
rect 29023 -20007 29079 -19951
rect 29133 -20007 29189 -19951
rect 28803 -20117 28859 -20061
rect 28913 -20117 28969 -20061
rect 29023 -20117 29079 -20061
rect 29133 -20117 29189 -20061
rect 28797 -20245 28853 -20189
rect 28907 -20245 28963 -20189
rect 29017 -20245 29073 -20189
rect 29127 -20245 29183 -20189
rect 28797 -20355 28853 -20299
rect 28907 -20355 28963 -20299
rect 29017 -20355 29073 -20299
rect 29127 -20355 29183 -20299
rect 28797 -20465 28853 -20409
rect 28907 -20465 28963 -20409
rect 29017 -20465 29073 -20409
rect 29127 -20465 29183 -20409
rect 28797 -20575 28853 -20519
rect 28907 -20575 28963 -20519
rect 29017 -20575 29073 -20519
rect 29127 -20575 29183 -20519
rect 28796 -20861 28852 -20805
rect 28906 -20861 28962 -20805
rect 29016 -20861 29072 -20805
rect 29126 -20861 29182 -20805
rect 94101 -19961 94157 -19905
rect 94211 -19961 94267 -19905
rect 94321 -19961 94377 -19905
rect 94431 -19961 94487 -19905
rect 94101 -20071 94157 -20015
rect 94211 -20071 94267 -20015
rect 94321 -20071 94377 -20015
rect 94431 -20071 94487 -20015
rect 94101 -20181 94157 -20125
rect 94211 -20181 94267 -20125
rect 94321 -20181 94377 -20125
rect 94431 -20181 94487 -20125
rect 94101 -20291 94157 -20235
rect 94211 -20291 94267 -20235
rect 94321 -20291 94377 -20235
rect 94431 -20291 94487 -20235
rect 94101 -20401 94157 -20345
rect 94211 -20401 94267 -20345
rect 94321 -20401 94377 -20345
rect 94431 -20401 94487 -20345
rect 94101 -20511 94157 -20455
rect 94211 -20511 94267 -20455
rect 94321 -20511 94377 -20455
rect 94431 -20511 94487 -20455
rect 94101 -20621 94157 -20565
rect 94211 -20621 94267 -20565
rect 94321 -20621 94377 -20565
rect 94431 -20621 94487 -20565
rect 28796 -20971 28852 -20915
rect 28906 -20971 28962 -20915
rect 29016 -20971 29072 -20915
rect 29126 -20971 29182 -20915
rect 28790 -21099 28846 -21043
rect 28900 -21099 28956 -21043
rect 29010 -21099 29066 -21043
rect 29120 -21099 29176 -21043
rect 28790 -21209 28846 -21153
rect 28900 -21209 28956 -21153
rect 29010 -21209 29066 -21153
rect 29120 -21209 29176 -21153
rect 28790 -21319 28846 -21263
rect 28900 -21319 28956 -21263
rect 29010 -21319 29066 -21263
rect 29120 -21319 29176 -21263
rect 28790 -21429 28846 -21373
rect 28900 -21429 28956 -21373
rect 29010 -21429 29066 -21373
rect 29120 -21429 29176 -21373
rect 93836 -20938 93892 -20882
rect 93946 -20938 94002 -20882
rect 94056 -20938 94112 -20882
rect 94166 -20938 94222 -20882
rect 93836 -21048 93892 -20992
rect 93946 -21048 94002 -20992
rect 94056 -21048 94112 -20992
rect 94166 -21048 94222 -20992
rect 93836 -21158 93892 -21102
rect 93946 -21158 94002 -21102
rect 94056 -21158 94112 -21102
rect 94166 -21158 94222 -21102
rect 93836 -21268 93892 -21212
rect 93946 -21268 94002 -21212
rect 94056 -21268 94112 -21212
rect 94166 -21268 94222 -21212
rect 93836 -21378 93892 -21322
rect 93946 -21378 94002 -21322
rect 94056 -21378 94112 -21322
rect 94166 -21378 94222 -21322
rect 93836 -21488 93892 -21432
rect 93946 -21488 94002 -21432
rect 94056 -21488 94112 -21432
rect 94166 -21488 94222 -21432
rect 93836 -21598 93892 -21542
rect 93946 -21598 94002 -21542
rect 94056 -21598 94112 -21542
rect 94166 -21598 94222 -21542
rect 27330 -22741 27386 -22685
rect 27440 -22741 27496 -22685
rect 27550 -22741 27606 -22685
rect 27660 -22741 27716 -22685
rect 27330 -22851 27386 -22795
rect 27440 -22851 27496 -22795
rect 27550 -22851 27606 -22795
rect 27660 -22851 27716 -22795
rect 27324 -22979 27380 -22923
rect 27434 -22979 27490 -22923
rect 27544 -22979 27600 -22923
rect 27654 -22979 27710 -22923
rect 27324 -23089 27380 -23033
rect 27434 -23089 27490 -23033
rect 27544 -23089 27600 -23033
rect 27654 -23089 27710 -23033
rect 27324 -23199 27380 -23143
rect 27434 -23199 27490 -23143
rect 27544 -23199 27600 -23143
rect 27654 -23199 27710 -23143
rect 27324 -23309 27380 -23253
rect 27434 -23309 27490 -23253
rect 27544 -23309 27600 -23253
rect 27654 -23309 27710 -23253
rect 56591 -27874 56647 -27818
rect 56701 -27874 56757 -27818
rect 56811 -27874 56867 -27818
rect 56921 -27874 56977 -27818
rect 57031 -27874 57087 -27818
rect 57141 -27874 57197 -27818
rect 57251 -27874 57307 -27818
rect 56591 -27984 56647 -27928
rect 56701 -27984 56757 -27928
rect 56811 -27984 56867 -27928
rect 56921 -27984 56977 -27928
rect 57031 -27984 57087 -27928
rect 57141 -27984 57197 -27928
rect 57251 -27984 57307 -27928
rect 56591 -28094 56647 -28038
rect 56701 -28094 56757 -28038
rect 56811 -28094 56867 -28038
rect 56921 -28094 56977 -28038
rect 57031 -28094 57087 -28038
rect 57141 -28094 57197 -28038
rect 57251 -28094 57307 -28038
rect 56591 -28204 56647 -28148
rect 56701 -28204 56757 -28148
rect 56811 -28204 56867 -28148
rect 56921 -28204 56977 -28148
rect 57031 -28204 57087 -28148
rect 57141 -28204 57197 -28148
rect 57251 -28204 57307 -28148
rect 56591 -28314 56647 -28258
rect 56701 -28314 56757 -28258
rect 56811 -28314 56867 -28258
rect 56921 -28314 56977 -28258
rect 57031 -28314 57087 -28258
rect 57141 -28314 57197 -28258
rect 57251 -28314 57307 -28258
rect 56591 -28424 56647 -28368
rect 56701 -28424 56757 -28368
rect 56811 -28424 56867 -28368
rect 56921 -28424 56977 -28368
rect 57031 -28424 57087 -28368
rect 57141 -28424 57197 -28368
rect 57251 -28424 57307 -28368
rect 56591 -28534 56647 -28478
rect 56701 -28534 56757 -28478
rect 56811 -28534 56867 -28478
rect 56921 -28534 56977 -28478
rect 57031 -28534 57087 -28478
rect 57141 -28534 57197 -28478
rect 57251 -28534 57307 -28478
rect 56591 -28644 56647 -28588
rect 56701 -28644 56757 -28588
rect 56811 -28644 56867 -28588
rect 56921 -28644 56977 -28588
rect 57031 -28644 57087 -28588
rect 57141 -28644 57197 -28588
rect 57251 -28644 57307 -28588
rect 39307 -29003 39363 -28947
rect 39417 -29003 39473 -28947
rect 39527 -29003 39583 -28947
rect 39637 -29003 39693 -28947
rect 39747 -29003 39803 -28947
rect 39857 -29003 39913 -28947
rect 39967 -29003 40023 -28947
rect 39307 -29113 39363 -29057
rect 39417 -29113 39473 -29057
rect 39527 -29113 39583 -29057
rect 39637 -29113 39693 -29057
rect 39747 -29113 39803 -29057
rect 39857 -29113 39913 -29057
rect 39967 -29113 40023 -29057
rect 39307 -29223 39363 -29167
rect 39417 -29223 39473 -29167
rect 39527 -29223 39583 -29167
rect 39637 -29223 39693 -29167
rect 39747 -29223 39803 -29167
rect 39857 -29223 39913 -29167
rect 39967 -29223 40023 -29167
rect 39307 -29333 39363 -29277
rect 39417 -29333 39473 -29277
rect 39527 -29333 39583 -29277
rect 39637 -29333 39693 -29277
rect 39747 -29333 39803 -29277
rect 39857 -29333 39913 -29277
rect 39967 -29333 40023 -29277
rect 39307 -29443 39363 -29387
rect 39417 -29443 39473 -29387
rect 39527 -29443 39583 -29387
rect 39637 -29443 39693 -29387
rect 39747 -29443 39803 -29387
rect 39857 -29443 39913 -29387
rect 39967 -29443 40023 -29387
rect 39307 -29553 39363 -29497
rect 39417 -29553 39473 -29497
rect 39527 -29553 39583 -29497
rect 39637 -29553 39693 -29497
rect 39747 -29553 39803 -29497
rect 39857 -29553 39913 -29497
rect 39967 -29553 40023 -29497
rect 39307 -29663 39363 -29607
rect 39417 -29663 39473 -29607
rect 39527 -29663 39583 -29607
rect 39637 -29663 39693 -29607
rect 39747 -29663 39803 -29607
rect 39857 -29663 39913 -29607
rect 39967 -29663 40023 -29607
rect 39307 -29773 39363 -29717
rect 39417 -29773 39473 -29717
rect 39527 -29773 39583 -29717
rect 39637 -29773 39693 -29717
rect 39747 -29773 39803 -29717
rect 39857 -29773 39913 -29717
rect 39967 -29773 40023 -29717
rect 112129 -27914 112185 -27858
rect 112239 -27914 112295 -27858
rect 112349 -27914 112405 -27858
rect 112459 -27914 112515 -27858
rect 112569 -27914 112625 -27858
rect 112679 -27914 112735 -27858
rect 112789 -27914 112845 -27858
rect 112129 -28024 112185 -27968
rect 112239 -28024 112295 -27968
rect 112349 -28024 112405 -27968
rect 112459 -28024 112515 -27968
rect 112569 -28024 112625 -27968
rect 112679 -28024 112735 -27968
rect 112789 -28024 112845 -27968
rect 112129 -28134 112185 -28078
rect 112239 -28134 112295 -28078
rect 112349 -28134 112405 -28078
rect 112459 -28134 112515 -28078
rect 112569 -28134 112625 -28078
rect 112679 -28134 112735 -28078
rect 112789 -28134 112845 -28078
rect 112129 -28244 112185 -28188
rect 112239 -28244 112295 -28188
rect 112349 -28244 112405 -28188
rect 112459 -28244 112515 -28188
rect 112569 -28244 112625 -28188
rect 112679 -28244 112735 -28188
rect 112789 -28244 112845 -28188
rect 112129 -28354 112185 -28298
rect 112239 -28354 112295 -28298
rect 112349 -28354 112405 -28298
rect 112459 -28354 112515 -28298
rect 112569 -28354 112625 -28298
rect 112679 -28354 112735 -28298
rect 112789 -28354 112845 -28298
rect 112129 -28464 112185 -28408
rect 112239 -28464 112295 -28408
rect 112349 -28464 112405 -28408
rect 112459 -28464 112515 -28408
rect 112569 -28464 112625 -28408
rect 112679 -28464 112735 -28408
rect 112789 -28464 112845 -28408
rect 112129 -28574 112185 -28518
rect 112239 -28574 112295 -28518
rect 112349 -28574 112405 -28518
rect 112459 -28574 112515 -28518
rect 112569 -28574 112625 -28518
rect 112679 -28574 112735 -28518
rect 112789 -28574 112845 -28518
rect 110768 -29080 110824 -29024
rect 110878 -29080 110934 -29024
rect 110988 -29080 111044 -29024
rect 111098 -29080 111154 -29024
rect 111208 -29080 111264 -29024
rect 111318 -29080 111374 -29024
rect 111428 -29080 111484 -29024
rect 110768 -29190 110824 -29134
rect 110878 -29190 110934 -29134
rect 110988 -29190 111044 -29134
rect 111098 -29190 111154 -29134
rect 111208 -29190 111264 -29134
rect 111318 -29190 111374 -29134
rect 111428 -29190 111484 -29134
rect 110768 -29300 110824 -29244
rect 110878 -29300 110934 -29244
rect 110988 -29300 111044 -29244
rect 111098 -29300 111154 -29244
rect 111208 -29300 111264 -29244
rect 111318 -29300 111374 -29244
rect 111428 -29300 111484 -29244
rect 110768 -29410 110824 -29354
rect 110878 -29410 110934 -29354
rect 110988 -29410 111044 -29354
rect 111098 -29410 111154 -29354
rect 111208 -29410 111264 -29354
rect 111318 -29410 111374 -29354
rect 111428 -29410 111484 -29354
rect 110768 -29520 110824 -29464
rect 110878 -29520 110934 -29464
rect 110988 -29520 111044 -29464
rect 111098 -29520 111154 -29464
rect 111208 -29520 111264 -29464
rect 111318 -29520 111374 -29464
rect 111428 -29520 111484 -29464
rect 110768 -29630 110824 -29574
rect 110878 -29630 110934 -29574
rect 110988 -29630 111044 -29574
rect 111098 -29630 111154 -29574
rect 111208 -29630 111264 -29574
rect 111318 -29630 111374 -29574
rect 111428 -29630 111484 -29574
rect 110768 -29740 110824 -29684
rect 110878 -29740 110934 -29684
rect 110988 -29740 111044 -29684
rect 111098 -29740 111154 -29684
rect 111208 -29740 111264 -29684
rect 111318 -29740 111374 -29684
rect 111428 -29740 111484 -29684
rect 129566 962 129622 1018
rect 129676 962 129732 1018
rect 129566 852 129622 908
rect 129676 852 129732 908
rect 129566 742 129622 798
rect 129676 742 129732 798
rect 129566 632 129622 688
rect 129676 632 129732 688
rect 129566 522 129622 578
rect 129676 522 129732 578
rect 129566 412 129622 468
rect 129676 412 129732 468
rect 129891 1647 129947 1703
rect 130001 1647 130057 1703
rect 129891 1537 129947 1593
rect 130001 1537 130057 1593
rect 129891 1427 129947 1483
rect 130001 1427 130057 1483
rect 129891 1317 129947 1373
rect 130001 1317 130057 1373
rect 129891 1207 129947 1263
rect 130001 1207 130057 1263
rect 129891 1097 129947 1153
rect 130001 1097 130057 1153
rect 130234 2320 130290 2376
rect 130344 2320 130400 2376
rect 130234 2210 130290 2266
rect 130344 2210 130400 2266
rect 130234 2100 130290 2156
rect 130344 2100 130400 2156
rect 130234 1990 130290 2046
rect 130344 1990 130400 2046
rect 130234 1880 130290 1936
rect 130344 1880 130400 1936
rect 130234 1770 130290 1826
rect 130344 1770 130400 1826
rect 130581 3063 130637 3119
rect 130691 3063 130747 3119
rect 130581 2953 130637 3009
rect 130691 2953 130747 3009
rect 130581 2843 130637 2899
rect 130691 2843 130747 2899
rect 130581 2733 130637 2789
rect 130691 2733 130747 2789
rect 130581 2623 130637 2679
rect 130691 2623 130747 2679
rect 130581 2513 130637 2569
rect 130691 2513 130747 2569
<< metal3 >>
rect 20909 17651 21799 17663
rect 1612 16822 21799 17651
rect 5559 11279 6443 11604
rect 6118 10608 6443 11279
rect 20909 10608 21799 16822
rect 44608 17222 112987 17411
rect 44608 17166 112156 17222
rect 112212 17166 112266 17222
rect 112322 17166 112376 17222
rect 112432 17166 112486 17222
rect 112542 17166 112596 17222
rect 112652 17166 112706 17222
rect 112762 17166 112816 17222
rect 112872 17166 112987 17222
rect 44608 17112 112987 17166
rect 44608 17056 112156 17112
rect 112212 17056 112266 17112
rect 112322 17056 112376 17112
rect 112432 17056 112486 17112
rect 112542 17056 112596 17112
rect 112652 17056 112706 17112
rect 112762 17056 112816 17112
rect 112872 17056 112987 17112
rect 44608 17002 112987 17056
rect 44608 16946 112156 17002
rect 112212 16946 112266 17002
rect 112322 16946 112376 17002
rect 112432 16946 112486 17002
rect 112542 16946 112596 17002
rect 112652 16946 112706 17002
rect 112762 16946 112816 17002
rect 112872 16946 112987 17002
rect 44608 16892 112987 16946
rect 44608 16836 112156 16892
rect 112212 16836 112266 16892
rect 112322 16836 112376 16892
rect 112432 16836 112486 16892
rect 112542 16836 112596 16892
rect 112652 16836 112706 16892
rect 112762 16836 112816 16892
rect 112872 16836 112987 16892
rect 44608 16782 112987 16836
rect 44608 16726 112156 16782
rect 112212 16726 112266 16782
rect 112322 16726 112376 16782
rect 112432 16726 112486 16782
rect 112542 16726 112596 16782
rect 112652 16726 112706 16782
rect 112762 16726 112816 16782
rect 112872 16726 112987 16782
rect 44608 16672 112987 16726
rect 44608 16616 112156 16672
rect 112212 16616 112266 16672
rect 112322 16616 112376 16672
rect 112432 16616 112486 16672
rect 112542 16616 112596 16672
rect 112652 16616 112706 16672
rect 112762 16616 112816 16672
rect 112872 16616 112987 16672
rect 44608 16562 112987 16616
rect 44608 16506 112156 16562
rect 112212 16506 112266 16562
rect 112322 16506 112376 16562
rect 112432 16506 112486 16562
rect 112542 16506 112596 16562
rect 112652 16506 112706 16562
rect 112762 16506 112816 16562
rect 112872 16506 112987 16562
rect 44608 16215 112987 16506
rect 44608 16094 47382 16215
rect 74833 16094 75735 16215
rect 27299 10665 27726 10700
rect 27299 10609 27330 10665
rect 27386 10609 27440 10665
rect 27496 10609 27550 10665
rect 27606 10609 27660 10665
rect 27716 10609 27726 10665
rect 27299 10608 27726 10609
rect 6118 10283 11003 10608
rect 17718 10555 27726 10608
rect 17718 10499 27330 10555
rect 27386 10499 27440 10555
rect 27496 10499 27550 10555
rect 27606 10499 27660 10555
rect 27716 10499 27726 10555
rect 17718 10445 27726 10499
rect 17718 10389 27330 10445
rect 27386 10389 27440 10445
rect 27496 10389 27550 10445
rect 27606 10389 27660 10445
rect 27716 10389 27726 10445
rect 17718 10335 27726 10389
rect 17718 10283 27330 10335
rect 27299 10279 27330 10283
rect 27386 10279 27440 10335
rect 27496 10279 27550 10335
rect 27606 10279 27660 10335
rect 27716 10279 27726 10335
rect 27299 10225 27726 10279
rect 27299 10169 27330 10225
rect 27386 10169 27440 10225
rect 27496 10169 27550 10225
rect 27606 10169 27660 10225
rect 27716 10169 27726 10225
rect 27299 10115 27726 10169
rect 27299 10059 27330 10115
rect 27386 10059 27440 10115
rect 27496 10059 27550 10115
rect 27606 10059 27660 10115
rect 27716 10059 27726 10115
rect 27299 10005 27726 10059
rect 27299 9949 27330 10005
rect 27386 9949 27440 10005
rect 27496 9949 27550 10005
rect 27606 9949 27660 10005
rect 27716 9949 27726 10005
rect 27299 9895 27726 9949
rect 27299 9839 27330 9895
rect 27386 9839 27440 9895
rect 27496 9839 27550 9895
rect 27606 9839 27660 9895
rect 27716 9839 27726 9895
rect 27299 9773 27726 9839
rect 40945 6904 54699 7056
rect 40945 6771 51065 6904
rect 24251 6004 27844 6164
rect 30984 6135 31774 6185
rect 30984 6095 31032 6135
rect 30704 6079 31032 6095
rect 31088 6079 31142 6135
rect 31198 6079 31252 6135
rect 31308 6079 31362 6135
rect 31418 6079 31472 6135
rect 31528 6079 31582 6135
rect 31638 6079 31692 6135
rect 31748 6095 31774 6135
rect 40945 6095 41230 6771
rect 46392 6309 46957 6314
rect 31748 6079 41230 6095
rect 30704 6025 41230 6079
rect 24251 1827 24411 6004
rect 30704 5969 31032 6025
rect 31088 5969 31142 6025
rect 31198 5969 31252 6025
rect 31308 5969 31362 6025
rect 31418 5969 31472 6025
rect 31528 5969 31582 6025
rect 31638 5969 31692 6025
rect 31748 5969 41230 6025
rect 30704 5915 41230 5969
rect 43879 6293 44495 6294
rect 43879 6290 44498 6293
rect 46392 6290 46418 6309
rect 43879 6253 46418 6290
rect 46474 6253 46528 6309
rect 46584 6253 46638 6309
rect 46694 6253 46748 6309
rect 46804 6253 46858 6309
rect 46914 6290 46957 6309
rect 46914 6253 46958 6290
rect 43879 6250 46958 6253
rect 43879 6194 43928 6250
rect 43984 6194 44038 6250
rect 44094 6194 44148 6250
rect 44204 6194 44258 6250
rect 44314 6194 44368 6250
rect 44424 6199 46958 6250
rect 44424 6198 46638 6199
rect 44424 6197 46530 6198
rect 44424 6194 46421 6197
rect 43879 6141 46421 6194
rect 46477 6142 46530 6197
rect 46586 6143 46638 6198
rect 46694 6143 46748 6199
rect 46804 6143 46858 6199
rect 46914 6143 46958 6199
rect 46586 6142 46958 6143
rect 46477 6141 46958 6142
rect 43879 6140 46958 6141
rect 43879 6084 43928 6140
rect 43984 6084 44038 6140
rect 44094 6084 44148 6140
rect 44204 6084 44258 6140
rect 44314 6084 44368 6140
rect 44424 6092 46958 6140
rect 44424 6091 46527 6092
rect 44424 6084 46421 6091
rect 43879 6035 46421 6084
rect 46477 6036 46527 6091
rect 46583 6089 46958 6092
rect 46583 6036 46638 6089
rect 46477 6035 46638 6036
rect 43879 6033 46638 6035
rect 46694 6033 46748 6089
rect 46804 6033 46858 6089
rect 46914 6033 46958 6089
rect 43879 6030 46958 6033
rect 43879 5974 43928 6030
rect 43984 5974 44038 6030
rect 44094 5974 44148 6030
rect 44204 5974 44258 6030
rect 44314 5974 44368 6030
rect 44424 5996 46958 6030
rect 44424 5974 44495 5996
rect 43879 5958 44495 5974
rect 30704 5859 31032 5915
rect 31088 5859 31142 5915
rect 31198 5859 31252 5915
rect 31308 5859 31362 5915
rect 31418 5859 31472 5915
rect 31528 5859 31582 5915
rect 31638 5859 31692 5915
rect 31748 5859 41230 5915
rect 30704 5810 41230 5859
rect 30984 5805 31774 5810
rect 30984 5749 31032 5805
rect 31088 5749 31142 5805
rect 31198 5749 31252 5805
rect 31308 5749 31362 5805
rect 31418 5749 31472 5805
rect 31528 5749 31582 5805
rect 31638 5749 31692 5805
rect 31748 5749 31774 5805
rect 30984 5695 31774 5749
rect 30984 5639 31032 5695
rect 31088 5639 31142 5695
rect 31198 5639 31252 5695
rect 31308 5639 31362 5695
rect 31418 5639 31472 5695
rect 31528 5639 31582 5695
rect 31638 5639 31692 5695
rect 31748 5639 31774 5695
rect 30984 5585 31774 5639
rect 30984 5529 31032 5585
rect 31088 5529 31142 5585
rect 31198 5529 31252 5585
rect 31308 5529 31362 5585
rect 31418 5529 31472 5585
rect 31528 5529 31582 5585
rect 31638 5529 31692 5585
rect 31748 5529 31774 5585
rect 30984 5475 31774 5529
rect 30984 5419 31032 5475
rect 31088 5419 31142 5475
rect 31198 5419 31252 5475
rect 31308 5419 31362 5475
rect 31418 5419 31472 5475
rect 31528 5419 31582 5475
rect 31638 5419 31692 5475
rect 31748 5419 31774 5475
rect 30984 5383 31774 5419
rect 30986 5382 31774 5383
rect 130565 3119 130761 3136
rect 130565 3063 130581 3119
rect 130637 3063 130691 3119
rect 130747 3063 130761 3119
rect 130565 3043 130761 3063
rect 130560 3009 132511 3043
rect 130560 2953 130581 3009
rect 130637 2953 130691 3009
rect 130747 2953 132511 3009
rect 130560 2899 132511 2953
rect 130560 2843 130581 2899
rect 130637 2843 130691 2899
rect 130747 2843 132511 2899
rect 130560 2789 132511 2843
rect 130560 2733 130581 2789
rect 130637 2733 130691 2789
rect 130747 2733 132511 2789
rect 130560 2679 132511 2733
rect 130560 2623 130581 2679
rect 130637 2623 130691 2679
rect 130747 2623 132511 2679
rect 130560 2569 132511 2623
rect 130560 2513 130581 2569
rect 130637 2513 130691 2569
rect 130747 2513 132511 2569
rect 130560 2494 132511 2513
rect 130218 2376 130414 2393
rect 130218 2320 130234 2376
rect 130290 2320 130344 2376
rect 130400 2320 130414 2376
rect 130218 2301 130414 2320
rect 8402 1667 24411 1827
rect 130207 2266 132158 2301
rect 130207 2210 130234 2266
rect 130290 2210 130344 2266
rect 130400 2210 132158 2266
rect 130207 2156 132158 2210
rect 130207 2100 130234 2156
rect 130290 2100 130344 2156
rect 130400 2100 132158 2156
rect 130207 2046 132158 2100
rect 130207 1990 130234 2046
rect 130290 1990 130344 2046
rect 130400 1990 132158 2046
rect 130207 1936 132158 1990
rect 130207 1880 130234 1936
rect 130290 1880 130344 1936
rect 130400 1880 132158 1936
rect 130207 1826 132158 1880
rect 93840 1746 111579 1814
rect 130207 1770 130234 1826
rect 130290 1770 130344 1826
rect 130400 1770 132158 1826
rect 130207 1752 132158 1770
rect 93840 1690 110643 1746
rect 110699 1690 110753 1746
rect 110809 1690 110863 1746
rect 110919 1690 110973 1746
rect 111029 1690 111083 1746
rect 111139 1690 111193 1746
rect 111249 1690 111303 1746
rect 111359 1690 111579 1746
rect 93840 1636 111579 1690
rect 93840 1580 110643 1636
rect 110699 1580 110753 1636
rect 110809 1580 110863 1636
rect 110919 1580 110973 1636
rect 111029 1580 111083 1636
rect 111139 1580 111193 1636
rect 111249 1580 111303 1636
rect 111359 1580 111579 1636
rect 129875 1703 130071 1720
rect 129875 1647 129891 1703
rect 129947 1647 130001 1703
rect 130057 1647 130071 1703
rect 129875 1625 130071 1647
rect 93840 1526 111579 1580
rect 93840 1470 110643 1526
rect 110699 1470 110753 1526
rect 110809 1470 110863 1526
rect 110919 1470 110973 1526
rect 111029 1470 111083 1526
rect 111139 1470 111193 1526
rect 111249 1470 111303 1526
rect 111359 1470 111579 1526
rect 93840 1416 111579 1470
rect 93840 1360 110643 1416
rect 110699 1360 110753 1416
rect 110809 1360 110863 1416
rect 110919 1360 110973 1416
rect 111029 1360 111083 1416
rect 111139 1360 111193 1416
rect 111249 1360 111303 1416
rect 111359 1360 111579 1416
rect 93840 1306 111579 1360
rect 93840 1250 110643 1306
rect 110699 1250 110753 1306
rect 110809 1250 110863 1306
rect 110919 1250 110973 1306
rect 111029 1250 111083 1306
rect 111139 1250 111193 1306
rect 111249 1250 111303 1306
rect 111359 1250 111579 1306
rect 93840 1196 111579 1250
rect 93840 1140 110643 1196
rect 110699 1140 110753 1196
rect 110809 1140 110863 1196
rect 110919 1140 110973 1196
rect 111029 1140 111083 1196
rect 111139 1140 111193 1196
rect 111249 1140 111303 1196
rect 111359 1140 111579 1196
rect 93840 1086 111579 1140
rect 93840 1030 110643 1086
rect 110699 1030 110753 1086
rect 110809 1030 110863 1086
rect 110919 1030 110973 1086
rect 111029 1030 111083 1086
rect 111139 1030 111193 1086
rect 111249 1030 111303 1086
rect 111359 1030 111579 1086
rect 129864 1593 131815 1625
rect 129864 1537 129891 1593
rect 129947 1537 130001 1593
rect 130057 1537 131815 1593
rect 129864 1483 131815 1537
rect 129864 1427 129891 1483
rect 129947 1427 130001 1483
rect 130057 1427 131815 1483
rect 129864 1373 131815 1427
rect 129864 1317 129891 1373
rect 129947 1317 130001 1373
rect 130057 1317 131815 1373
rect 129864 1263 131815 1317
rect 129864 1207 129891 1263
rect 129947 1207 130001 1263
rect 130057 1207 131815 1263
rect 129864 1153 131815 1207
rect 129864 1097 129891 1153
rect 129947 1097 130001 1153
rect 130057 1097 131815 1153
rect 129864 1076 131815 1097
rect 93840 992 111579 1030
rect 129550 1018 129746 1035
rect 129550 962 129566 1018
rect 129622 962 129676 1018
rect 129732 962 129746 1018
rect 129550 943 129746 962
rect 129546 908 131497 943
rect 129546 852 129566 908
rect 129622 852 129676 908
rect 129732 852 131497 908
rect 129546 798 131497 852
rect 129546 742 129566 798
rect 129622 742 129676 798
rect 129732 742 131497 798
rect 129546 688 131497 742
rect 129546 632 129566 688
rect 129622 632 129676 688
rect 129732 632 131497 688
rect 129546 578 131497 632
rect 129546 522 129566 578
rect 129622 522 129676 578
rect 129732 522 131497 578
rect 129546 468 131497 522
rect 129546 412 129566 468
rect 129622 412 129676 468
rect 129732 412 131497 468
rect 129546 394 131497 412
rect 4289 -643 4702 -639
rect 4263 -658 4702 -643
rect 4263 -714 4298 -658
rect 4354 -714 4408 -658
rect 4464 -714 4518 -658
rect 4574 -714 4628 -658
rect 4684 -714 4702 -658
rect 4263 -768 4702 -714
rect 4263 -824 4298 -768
rect 4354 -824 4408 -768
rect 4464 -824 4518 -768
rect 4574 -824 4628 -768
rect 4684 -824 4702 -768
rect 4263 -1423 4702 -824
rect 64971 -959 109855 -951
rect 64799 -1002 109855 -959
rect 64799 -1058 109095 -1002
rect 109151 -1058 109205 -1002
rect 109261 -1058 109315 -1002
rect 109371 -1058 109425 -1002
rect 109481 -1058 109535 -1002
rect 109591 -1058 109645 -1002
rect 109701 -1058 109755 -1002
rect 109811 -1058 109855 -1002
rect 64799 -1112 109855 -1058
rect 64799 -1168 109095 -1112
rect 109151 -1168 109205 -1112
rect 109261 -1168 109315 -1112
rect 109371 -1168 109425 -1112
rect 109481 -1168 109535 -1112
rect 109591 -1168 109645 -1112
rect 109701 -1168 109755 -1112
rect 109811 -1168 109855 -1112
rect 64799 -1222 109855 -1168
rect 64799 -1278 109095 -1222
rect 109151 -1278 109205 -1222
rect 109261 -1278 109315 -1222
rect 109371 -1278 109425 -1222
rect 109481 -1278 109535 -1222
rect 109591 -1278 109645 -1222
rect 109701 -1278 109755 -1222
rect 109811 -1278 109855 -1222
rect 64799 -1332 109855 -1278
rect 64799 -1388 109095 -1332
rect 109151 -1388 109205 -1332
rect 109261 -1388 109315 -1332
rect 109371 -1388 109425 -1332
rect 109481 -1388 109535 -1332
rect 109591 -1388 109645 -1332
rect 109701 -1388 109755 -1332
rect 109811 -1388 109855 -1332
rect 4263 -1458 12429 -1423
rect 4263 -1514 10881 -1458
rect 10937 -1514 10991 -1458
rect 11047 -1514 11101 -1458
rect 11157 -1514 11211 -1458
rect 11267 -1514 11321 -1458
rect 11377 -1514 11431 -1458
rect 11487 -1514 11541 -1458
rect 11597 -1514 11670 -1458
rect 11726 -1514 11780 -1458
rect 11836 -1514 11890 -1458
rect 11946 -1514 12000 -1458
rect 12056 -1514 12110 -1458
rect 12166 -1514 12220 -1458
rect 12276 -1514 12330 -1458
rect 12386 -1514 12429 -1458
rect 4263 -1568 12429 -1514
rect 4263 -1624 10881 -1568
rect 10937 -1624 10991 -1568
rect 11047 -1624 11101 -1568
rect 11157 -1624 11211 -1568
rect 11267 -1624 11321 -1568
rect 11377 -1624 11431 -1568
rect 11487 -1624 11541 -1568
rect 11597 -1624 11670 -1568
rect 11726 -1624 11780 -1568
rect 11836 -1624 11890 -1568
rect 11946 -1624 12000 -1568
rect 12056 -1624 12110 -1568
rect 12166 -1624 12220 -1568
rect 12276 -1624 12330 -1568
rect 12386 -1624 12429 -1568
rect 4263 -1678 12429 -1624
rect 4263 -1734 10881 -1678
rect 10937 -1734 10991 -1678
rect 11047 -1734 11101 -1678
rect 11157 -1734 11211 -1678
rect 11267 -1734 11321 -1678
rect 11377 -1734 11431 -1678
rect 11487 -1734 11541 -1678
rect 11597 -1734 11670 -1678
rect 11726 -1734 11780 -1678
rect 11836 -1734 11890 -1678
rect 11946 -1734 12000 -1678
rect 12056 -1734 12110 -1678
rect 12166 -1734 12220 -1678
rect 12276 -1734 12330 -1678
rect 12386 -1734 12429 -1678
rect 4263 -1860 12429 -1734
rect 4805 -1862 12429 -1860
rect 64799 -1442 109855 -1388
rect 64799 -1498 109095 -1442
rect 109151 -1498 109205 -1442
rect 109261 -1498 109315 -1442
rect 109371 -1498 109425 -1442
rect 109481 -1498 109535 -1442
rect 109591 -1498 109645 -1442
rect 109701 -1498 109755 -1442
rect 109811 -1498 109855 -1442
rect 64799 -1552 109855 -1498
rect 64799 -1608 109095 -1552
rect 109151 -1608 109205 -1552
rect 109261 -1608 109315 -1552
rect 109371 -1608 109425 -1552
rect 109481 -1608 109535 -1552
rect 109591 -1608 109645 -1552
rect 109701 -1608 109755 -1552
rect 109811 -1608 109855 -1552
rect 64799 -1662 109855 -1608
rect 64799 -1718 109095 -1662
rect 109151 -1718 109205 -1662
rect 109261 -1718 109315 -1662
rect 109371 -1718 109425 -1662
rect 109481 -1718 109535 -1662
rect 109591 -1718 109645 -1662
rect 109701 -1718 109755 -1662
rect 109811 -1718 109855 -1662
rect 64799 -1755 109855 -1718
rect 25865 -4126 30790 -4105
rect 25865 -4146 30811 -4126
rect 25865 -4147 26470 -4146
rect 25865 -4203 25883 -4147
rect 25939 -4203 25993 -4147
rect 26049 -4203 26103 -4147
rect 26159 -4203 26213 -4147
rect 26269 -4203 26323 -4147
rect 26379 -4202 26470 -4147
rect 26526 -4202 26580 -4146
rect 26636 -4202 26690 -4146
rect 26746 -4151 30811 -4146
rect 26746 -4202 30166 -4151
rect 26379 -4203 30166 -4202
rect 25865 -4207 30166 -4203
rect 30222 -4207 30276 -4151
rect 30332 -4207 30386 -4151
rect 30442 -4207 30496 -4151
rect 30552 -4207 30606 -4151
rect 30662 -4207 30716 -4151
rect 30772 -4207 30811 -4151
rect 25865 -4256 30811 -4207
rect 25865 -4257 26470 -4256
rect 25865 -4313 25883 -4257
rect 25939 -4313 25993 -4257
rect 26049 -4313 26103 -4257
rect 26159 -4313 26213 -4257
rect 26269 -4313 26323 -4257
rect 26379 -4312 26470 -4257
rect 26526 -4312 26580 -4256
rect 26636 -4312 26690 -4256
rect 26746 -4261 30811 -4256
rect 26746 -4312 30166 -4261
rect 26379 -4313 30166 -4312
rect 25865 -4317 30166 -4313
rect 30222 -4317 30276 -4261
rect 30332 -4317 30386 -4261
rect 30442 -4317 30496 -4261
rect 30552 -4317 30606 -4261
rect 30662 -4317 30716 -4261
rect 30772 -4317 30811 -4261
rect 25865 -4352 30811 -4317
rect 30146 -4376 30811 -4352
rect 64799 -4729 65536 -1755
rect 107175 -2423 107963 -2372
rect 107175 -2434 107221 -2423
rect 65941 -2479 107221 -2434
rect 107277 -2479 107331 -2423
rect 107387 -2479 107441 -2423
rect 107497 -2479 107551 -2423
rect 107607 -2479 107661 -2423
rect 107717 -2479 107771 -2423
rect 107827 -2479 107881 -2423
rect 107937 -2479 107963 -2423
rect 65941 -2533 107963 -2479
rect 65941 -2589 107221 -2533
rect 107277 -2589 107331 -2533
rect 107387 -2589 107441 -2533
rect 107497 -2589 107551 -2533
rect 107607 -2589 107661 -2533
rect 107717 -2589 107771 -2533
rect 107827 -2589 107881 -2533
rect 107937 -2589 107963 -2533
rect 65941 -2643 107963 -2589
rect 65941 -2699 107221 -2643
rect 107277 -2699 107331 -2643
rect 107387 -2699 107441 -2643
rect 107497 -2699 107551 -2643
rect 107607 -2699 107661 -2643
rect 107717 -2699 107771 -2643
rect 107827 -2699 107881 -2643
rect 107937 -2699 107963 -2643
rect 65941 -2753 107963 -2699
rect 65941 -2809 107221 -2753
rect 107277 -2809 107331 -2753
rect 107387 -2809 107441 -2753
rect 107497 -2809 107551 -2753
rect 107607 -2809 107661 -2753
rect 107717 -2809 107771 -2753
rect 107827 -2809 107881 -2753
rect 107937 -2809 107963 -2753
rect 65941 -2863 107963 -2809
rect 65941 -2919 107221 -2863
rect 107277 -2919 107331 -2863
rect 107387 -2919 107441 -2863
rect 107497 -2919 107551 -2863
rect 107607 -2919 107661 -2863
rect 107717 -2919 107771 -2863
rect 107827 -2919 107881 -2863
rect 107937 -2919 107963 -2863
rect 65941 -2973 107963 -2919
rect 65941 -3029 107221 -2973
rect 107277 -3029 107331 -2973
rect 107387 -3029 107441 -2973
rect 107497 -3029 107551 -2973
rect 107607 -3029 107661 -2973
rect 107717 -3029 107771 -2973
rect 107827 -3029 107881 -2973
rect 107937 -3029 107963 -2973
rect 65941 -3083 107963 -3029
rect 65941 -3139 107221 -3083
rect 107277 -3139 107331 -3083
rect 107387 -3139 107441 -3083
rect 107497 -3139 107551 -3083
rect 107607 -3139 107661 -3083
rect 107717 -3139 107771 -3083
rect 107827 -3139 107881 -3083
rect 107937 -3139 107963 -3083
rect 65941 -3176 107963 -3139
rect 64799 -4803 65255 -4729
rect 65941 -5208 66683 -3176
rect 5458 -7125 6386 -6800
rect 6061 -7795 6386 -7125
rect 27247 -7685 27774 -7670
rect 27247 -7741 27262 -7685
rect 27318 -7741 27372 -7685
rect 27428 -7741 27482 -7685
rect 27538 -7741 27592 -7685
rect 27648 -7741 27702 -7685
rect 27758 -7741 27774 -7685
rect 27247 -7795 27774 -7741
rect 6061 -8120 12430 -7795
rect 17702 -7851 27262 -7795
rect 27318 -7851 27372 -7795
rect 27428 -7851 27482 -7795
rect 27538 -7851 27592 -7795
rect 27648 -7851 27702 -7795
rect 27758 -7851 27775 -7795
rect 17702 -7905 27775 -7851
rect 17702 -7961 27262 -7905
rect 27318 -7961 27372 -7905
rect 27428 -7961 27482 -7905
rect 27538 -7961 27592 -7905
rect 27648 -7961 27702 -7905
rect 27758 -7961 27775 -7905
rect 17702 -8015 27775 -7961
rect 17702 -8071 27262 -8015
rect 27318 -8071 27372 -8015
rect 27428 -8071 27482 -8015
rect 27538 -8071 27592 -8015
rect 27648 -8071 27702 -8015
rect 27758 -8071 27775 -8015
rect 17702 -8120 27775 -8071
rect 27247 -8121 27774 -8120
rect 31244 -11628 31777 -11619
rect 31244 -11684 31255 -11628
rect 31311 -11684 31365 -11628
rect 31421 -11684 31475 -11628
rect 31531 -11684 31585 -11628
rect 31641 -11684 31695 -11628
rect 31751 -11667 31777 -11628
rect 31751 -11684 44491 -11667
rect 31244 -11738 44491 -11684
rect 31244 -11794 31255 -11738
rect 31311 -11794 31365 -11738
rect 31421 -11794 31475 -11738
rect 31531 -11794 31585 -11738
rect 31641 -11794 31695 -11738
rect 31751 -11794 44491 -11738
rect 31244 -11848 44491 -11794
rect 31244 -11904 31255 -11848
rect 31311 -11904 31365 -11848
rect 31421 -11904 31475 -11848
rect 31531 -11904 31585 -11848
rect 31641 -11904 31695 -11848
rect 31751 -11904 44491 -11848
rect 31244 -11915 44491 -11904
rect 31244 -11958 40884 -11915
rect 31244 -12014 31255 -11958
rect 31311 -12014 31365 -11958
rect 31421 -12014 31475 -11958
rect 31531 -12014 31585 -11958
rect 31641 -12014 31695 -11958
rect 31751 -12014 40884 -11958
rect 31244 -12068 40884 -12014
rect 31244 -12124 31255 -12068
rect 31311 -12124 31365 -12068
rect 31421 -12124 31475 -12068
rect 31531 -12124 31585 -12068
rect 31641 -12124 31695 -12068
rect 31751 -12124 40884 -12068
rect 31244 -12148 40884 -12124
rect 31244 -12161 31777 -12148
rect 34037 -12353 34633 -12318
rect 36010 -12353 36795 -12344
rect 34035 -12382 36795 -12353
rect 34035 -12438 34121 -12382
rect 34177 -12438 34231 -12382
rect 34287 -12438 34341 -12382
rect 34397 -12438 34451 -12382
rect 34507 -12387 36795 -12382
rect 34507 -12438 36056 -12387
rect 34035 -12443 36056 -12438
rect 36112 -12443 36166 -12387
rect 36222 -12443 36276 -12387
rect 36332 -12443 36386 -12387
rect 36442 -12443 36496 -12387
rect 36552 -12443 36606 -12387
rect 36662 -12443 36716 -12387
rect 36772 -12443 36795 -12387
rect 34035 -12492 36795 -12443
rect 34035 -12548 34121 -12492
rect 34177 -12548 34231 -12492
rect 34287 -12548 34341 -12492
rect 34397 -12548 34451 -12492
rect 34507 -12497 36795 -12492
rect 34507 -12548 36056 -12497
rect 34035 -12553 36056 -12548
rect 36112 -12553 36166 -12497
rect 36222 -12553 36276 -12497
rect 36332 -12553 36386 -12497
rect 36442 -12553 36496 -12497
rect 36552 -12553 36606 -12497
rect 36662 -12553 36716 -12497
rect 36772 -12553 36795 -12497
rect 34035 -12602 36795 -12553
rect 34035 -12658 34121 -12602
rect 34177 -12658 34231 -12602
rect 34287 -12658 34341 -12602
rect 34397 -12658 34451 -12602
rect 34507 -12607 36795 -12602
rect 34507 -12658 36056 -12607
rect 34035 -12663 36056 -12658
rect 36112 -12663 36166 -12607
rect 36222 -12663 36276 -12607
rect 36332 -12663 36386 -12607
rect 36442 -12663 36496 -12607
rect 36552 -12663 36606 -12607
rect 36662 -12663 36716 -12607
rect 36772 -12663 36795 -12607
rect 34035 -12712 36795 -12663
rect 34035 -12768 34121 -12712
rect 34177 -12768 34231 -12712
rect 34287 -12768 34341 -12712
rect 34397 -12768 34451 -12712
rect 34507 -12717 36795 -12712
rect 34507 -12768 36056 -12717
rect 34035 -12773 36056 -12768
rect 36112 -12773 36166 -12717
rect 36222 -12773 36276 -12717
rect 36332 -12773 36386 -12717
rect 36442 -12773 36496 -12717
rect 36552 -12773 36606 -12717
rect 36662 -12773 36716 -12717
rect 36772 -12773 36795 -12717
rect 34035 -12788 36795 -12773
rect 34037 -12827 34633 -12788
rect 36010 -12810 36795 -12788
rect 29479 -13569 30536 -13568
rect 24625 -13596 30536 -13569
rect 24625 -13652 24679 -13596
rect 24735 -13652 24789 -13596
rect 24845 -13652 24899 -13596
rect 24955 -13652 25009 -13596
rect 25065 -13652 25119 -13596
rect 25175 -13652 25229 -13596
rect 25285 -13652 25339 -13596
rect 25395 -13652 30536 -13596
rect 24625 -13656 30536 -13652
rect 24625 -13664 30193 -13656
rect 24625 -13706 29533 -13664
rect 24625 -13762 24679 -13706
rect 24735 -13762 24789 -13706
rect 24845 -13762 24899 -13706
rect 24955 -13762 25009 -13706
rect 25065 -13762 25119 -13706
rect 25175 -13762 25229 -13706
rect 25285 -13762 25339 -13706
rect 25395 -13720 29533 -13706
rect 29589 -13720 29643 -13664
rect 29699 -13720 29753 -13664
rect 29809 -13720 29863 -13664
rect 29919 -13720 29973 -13664
rect 30029 -13720 30083 -13664
rect 30139 -13712 30193 -13664
rect 30249 -13712 30303 -13656
rect 30359 -13712 30413 -13656
rect 30469 -13712 30536 -13656
rect 30139 -13720 30536 -13712
rect 25395 -13762 30536 -13720
rect 24625 -13766 30536 -13762
rect 24625 -13774 30193 -13766
rect 24625 -13816 29533 -13774
rect 24625 -13872 24679 -13816
rect 24735 -13872 24789 -13816
rect 24845 -13872 24899 -13816
rect 24955 -13872 25009 -13816
rect 25065 -13872 25119 -13816
rect 25175 -13872 25229 -13816
rect 25285 -13872 25339 -13816
rect 25395 -13830 29533 -13816
rect 29589 -13830 29643 -13774
rect 29699 -13830 29753 -13774
rect 29809 -13830 29863 -13774
rect 29919 -13830 29973 -13774
rect 30029 -13830 30083 -13774
rect 30139 -13822 30193 -13774
rect 30249 -13822 30303 -13766
rect 30359 -13822 30413 -13766
rect 30469 -13822 30536 -13766
rect 30139 -13830 30536 -13822
rect 25395 -13872 30536 -13830
rect 24625 -13895 30536 -13872
rect 24636 -13896 25419 -13895
rect 29479 -13897 30536 -13895
rect 25861 -14409 26644 -14408
rect 29799 -14409 30669 -14407
rect 25861 -14420 30669 -14409
rect 25861 -14476 25904 -14420
rect 25960 -14476 26014 -14420
rect 26070 -14476 26124 -14420
rect 26180 -14476 26234 -14420
rect 26290 -14476 26344 -14420
rect 26400 -14476 26454 -14420
rect 26510 -14476 26564 -14420
rect 26620 -14469 30669 -14420
rect 26620 -14476 29852 -14469
rect 25861 -14525 29852 -14476
rect 29908 -14525 29962 -14469
rect 30018 -14525 30072 -14469
rect 30128 -14525 30249 -14469
rect 30305 -14525 30359 -14469
rect 30415 -14525 30469 -14469
rect 30525 -14525 30669 -14469
rect 25861 -14530 30669 -14525
rect 25861 -14586 25904 -14530
rect 25960 -14586 26014 -14530
rect 26070 -14586 26124 -14530
rect 26180 -14586 26234 -14530
rect 26290 -14586 26344 -14530
rect 26400 -14586 26454 -14530
rect 26510 -14586 26564 -14530
rect 26620 -14579 30669 -14530
rect 26620 -14586 29852 -14579
rect 25861 -14635 29852 -14586
rect 29908 -14635 29962 -14579
rect 30018 -14635 30072 -14579
rect 30128 -14635 30249 -14579
rect 30305 -14635 30359 -14579
rect 30415 -14635 30469 -14579
rect 30525 -14635 30669 -14579
rect 25861 -14640 30669 -14635
rect 25861 -14696 25904 -14640
rect 25960 -14696 26014 -14640
rect 26070 -14696 26124 -14640
rect 26180 -14696 26234 -14640
rect 26290 -14696 26344 -14640
rect 26400 -14696 26454 -14640
rect 26510 -14696 26564 -14640
rect 26620 -14696 30669 -14640
rect 25861 -14720 30669 -14696
rect 29799 -14722 30669 -14720
rect 109049 -14902 127801 -14868
rect 109049 -14958 109096 -14902
rect 109152 -14958 109206 -14902
rect 109262 -14958 109316 -14902
rect 109372 -14958 109426 -14902
rect 109482 -14958 109536 -14902
rect 109592 -14958 109646 -14902
rect 109702 -14958 109756 -14902
rect 109812 -14958 127801 -14902
rect 109049 -15012 127801 -14958
rect 109049 -15068 109096 -15012
rect 109152 -15068 109206 -15012
rect 109262 -15068 109316 -15012
rect 109372 -15068 109426 -15012
rect 109482 -15068 109536 -15012
rect 109592 -15068 109646 -15012
rect 109702 -15068 109756 -15012
rect 109812 -15068 127801 -15012
rect 109049 -15122 127801 -15068
rect 109049 -15178 109096 -15122
rect 109152 -15178 109206 -15122
rect 109262 -15178 109316 -15122
rect 109372 -15178 109426 -15122
rect 109482 -15178 109536 -15122
rect 109592 -15178 109646 -15122
rect 109702 -15178 109756 -15122
rect 109812 -15178 127801 -15122
rect 109049 -15232 127801 -15178
rect 109049 -15288 109096 -15232
rect 109152 -15288 109206 -15232
rect 109262 -15288 109316 -15232
rect 109372 -15288 109426 -15232
rect 109482 -15288 109536 -15232
rect 109592 -15288 109646 -15232
rect 109702 -15288 109756 -15232
rect 109812 -15288 127801 -15232
rect 109049 -15342 127801 -15288
rect 109049 -15398 109096 -15342
rect 109152 -15398 109206 -15342
rect 109262 -15398 109316 -15342
rect 109372 -15398 109426 -15342
rect 109482 -15398 109536 -15342
rect 109592 -15398 109646 -15342
rect 109702 -15398 109756 -15342
rect 109812 -15398 127801 -15342
rect 109049 -15452 127801 -15398
rect 109049 -15508 109096 -15452
rect 109152 -15508 109206 -15452
rect 109262 -15508 109316 -15452
rect 109372 -15508 109426 -15452
rect 109482 -15508 109536 -15452
rect 109592 -15508 109646 -15452
rect 109702 -15508 109756 -15452
rect 109812 -15508 127801 -15452
rect 109049 -15562 127801 -15508
rect 109049 -15618 109096 -15562
rect 109152 -15618 109206 -15562
rect 109262 -15618 109316 -15562
rect 109372 -15618 109426 -15562
rect 109482 -15618 109536 -15562
rect 109592 -15618 109646 -15562
rect 109702 -15618 109756 -15562
rect 109812 -15618 127801 -15562
rect 109049 -15656 127801 -15618
rect 107175 -16271 127459 -16235
rect 107175 -16327 107210 -16271
rect 107266 -16327 107320 -16271
rect 107376 -16327 107430 -16271
rect 107486 -16327 107540 -16271
rect 107596 -16327 107650 -16271
rect 107706 -16327 107760 -16271
rect 107816 -16327 107870 -16271
rect 107926 -16327 127459 -16271
rect 107175 -16381 127459 -16327
rect -832 -16409 -70 -16389
rect -832 -16413 22477 -16409
rect -832 -16469 -814 -16413
rect -758 -16469 -704 -16413
rect -648 -16469 -594 -16413
rect -538 -16469 -484 -16413
rect -428 -16469 -374 -16413
rect -318 -16469 -264 -16413
rect -208 -16469 -154 -16413
rect -98 -16439 22477 -16413
rect -98 -16469 21746 -16439
rect -832 -16495 21746 -16469
rect 21802 -16495 21856 -16439
rect 21912 -16495 21966 -16439
rect 22022 -16495 22076 -16439
rect 22132 -16495 22186 -16439
rect 22242 -16495 22296 -16439
rect 22352 -16495 22406 -16439
rect 22462 -16495 22477 -16439
rect 107175 -16437 107210 -16381
rect 107266 -16437 107320 -16381
rect 107376 -16437 107430 -16381
rect 107486 -16437 107540 -16381
rect 107596 -16437 107650 -16381
rect 107706 -16437 107760 -16381
rect 107816 -16437 107870 -16381
rect 107926 -16437 127459 -16381
rect -832 -16523 22477 -16495
rect -832 -16579 -814 -16523
rect -758 -16579 -704 -16523
rect -648 -16579 -594 -16523
rect -538 -16579 -484 -16523
rect -428 -16579 -374 -16523
rect -318 -16579 -264 -16523
rect -208 -16579 -154 -16523
rect -98 -16549 22477 -16523
rect 28339 -16519 31322 -16459
rect 107175 -16491 127459 -16437
rect 28339 -16525 31325 -16519
rect -98 -16579 21746 -16549
rect -832 -16605 21746 -16579
rect 21802 -16605 21856 -16549
rect 21912 -16605 21966 -16549
rect 22022 -16605 22076 -16549
rect 22132 -16605 22186 -16549
rect 22242 -16605 22296 -16549
rect 22352 -16605 22406 -16549
rect 22462 -16605 22477 -16549
rect -832 -16633 22477 -16605
rect -832 -16689 -814 -16633
rect -758 -16689 -704 -16633
rect -648 -16689 -594 -16633
rect -538 -16689 -484 -16633
rect -428 -16689 -374 -16633
rect -318 -16689 -264 -16633
rect -208 -16689 -154 -16633
rect -98 -16659 22477 -16633
rect -98 -16689 21746 -16659
rect -832 -16715 21746 -16689
rect 21802 -16715 21856 -16659
rect 21912 -16715 21966 -16659
rect 22022 -16715 22076 -16659
rect 22132 -16715 22186 -16659
rect 22242 -16715 22296 -16659
rect 22352 -16715 22406 -16659
rect 22462 -16715 22477 -16659
rect -832 -16743 22477 -16715
rect -832 -16799 -814 -16743
rect -758 -16799 -704 -16743
rect -648 -16799 -594 -16743
rect -538 -16799 -484 -16743
rect -428 -16799 -374 -16743
rect -318 -16799 -264 -16743
rect -208 -16799 -154 -16743
rect -98 -16769 22477 -16743
rect -98 -16799 21746 -16769
rect -832 -16825 21746 -16799
rect 21802 -16825 21856 -16769
rect 21912 -16825 21966 -16769
rect 22022 -16825 22076 -16769
rect 22132 -16825 22186 -16769
rect 22242 -16825 22296 -16769
rect 22352 -16825 22406 -16769
rect 22462 -16825 22477 -16769
rect -832 -16853 22477 -16825
rect -832 -16909 -814 -16853
rect -758 -16909 -704 -16853
rect -648 -16909 -594 -16853
rect -538 -16909 -484 -16853
rect -428 -16909 -374 -16853
rect -318 -16909 -264 -16853
rect -208 -16909 -154 -16853
rect -98 -16879 22477 -16853
rect -98 -16909 21746 -16879
rect -832 -16935 21746 -16909
rect 21802 -16935 21856 -16879
rect 21912 -16935 21966 -16879
rect 22022 -16935 22076 -16879
rect 22132 -16935 22186 -16879
rect 22242 -16935 22296 -16879
rect 22352 -16935 22406 -16879
rect 22462 -16935 22477 -16879
rect -832 -16963 22477 -16935
rect -832 -17019 -814 -16963
rect -758 -17019 -704 -16963
rect -648 -17019 -594 -16963
rect -538 -17019 -484 -16963
rect -428 -17019 -374 -16963
rect -318 -17019 -264 -16963
rect -208 -17019 -154 -16963
rect -98 -16989 22477 -16963
rect -98 -17019 21746 -16989
rect -832 -17045 21746 -17019
rect 21802 -17045 21856 -16989
rect 21912 -17045 21966 -16989
rect 22022 -17045 22076 -16989
rect 22132 -17045 22186 -16989
rect 22242 -17045 22296 -16989
rect 22352 -17045 22406 -16989
rect 22462 -17045 22477 -16989
rect 28338 -16556 31325 -16525
rect 28338 -16558 30894 -16556
rect 28338 -16562 28873 -16558
rect 28338 -16618 28388 -16562
rect 28444 -16618 28498 -16562
rect 28554 -16618 28608 -16562
rect 28664 -16618 28718 -16562
rect 28774 -16614 28873 -16562
rect 28929 -16614 28983 -16558
rect 29039 -16614 29093 -16558
rect 29149 -16614 29203 -16558
rect 29259 -16612 30894 -16558
rect 30950 -16612 31004 -16556
rect 31060 -16612 31114 -16556
rect 31170 -16612 31224 -16556
rect 31280 -16612 31325 -16556
rect 29259 -16614 31325 -16612
rect 28774 -16618 31325 -16614
rect 28338 -16666 31325 -16618
rect 28338 -16668 30894 -16666
rect 28338 -16672 28873 -16668
rect 28338 -16728 28388 -16672
rect 28444 -16728 28498 -16672
rect 28554 -16728 28608 -16672
rect 28664 -16728 28718 -16672
rect 28774 -16724 28873 -16672
rect 28929 -16724 28983 -16668
rect 29039 -16724 29093 -16668
rect 29149 -16724 29203 -16668
rect 29259 -16722 30894 -16668
rect 30950 -16722 31004 -16666
rect 31060 -16722 31114 -16666
rect 31170 -16722 31224 -16666
rect 31280 -16722 31325 -16666
rect 29259 -16724 31325 -16722
rect 28774 -16728 31325 -16724
rect 28338 -16776 31325 -16728
rect 28338 -16778 30894 -16776
rect 28338 -16782 28873 -16778
rect 28338 -16838 28388 -16782
rect 28444 -16838 28498 -16782
rect 28554 -16838 28608 -16782
rect 28664 -16838 28718 -16782
rect 28774 -16834 28873 -16782
rect 28929 -16834 28983 -16778
rect 29039 -16834 29093 -16778
rect 29149 -16834 29203 -16778
rect 29259 -16832 30894 -16778
rect 30950 -16832 31004 -16776
rect 31060 -16832 31114 -16776
rect 31170 -16832 31224 -16776
rect 31280 -16832 31325 -16776
rect 29259 -16834 31325 -16832
rect 28774 -16838 31325 -16834
rect 28338 -16886 31325 -16838
rect 28338 -16888 30894 -16886
rect 28338 -16892 28873 -16888
rect 28338 -16948 28388 -16892
rect 28444 -16948 28498 -16892
rect 28554 -16948 28608 -16892
rect 28664 -16948 28718 -16892
rect 28774 -16944 28873 -16892
rect 28929 -16944 28983 -16888
rect 29039 -16944 29093 -16888
rect 29149 -16944 29203 -16888
rect 29259 -16942 30894 -16888
rect 30950 -16942 31004 -16886
rect 31060 -16942 31114 -16886
rect 31170 -16942 31224 -16886
rect 31280 -16942 31325 -16886
rect 29259 -16944 31325 -16942
rect 28774 -16948 31325 -16944
rect 28338 -17012 31325 -16948
rect 107175 -16547 107210 -16491
rect 107266 -16547 107320 -16491
rect 107376 -16547 107430 -16491
rect 107486 -16547 107540 -16491
rect 107596 -16547 107650 -16491
rect 107706 -16547 107760 -16491
rect 107816 -16547 107870 -16491
rect 107926 -16547 127459 -16491
rect 107175 -16601 127459 -16547
rect 107175 -16657 107210 -16601
rect 107266 -16657 107320 -16601
rect 107376 -16657 107430 -16601
rect 107486 -16657 107540 -16601
rect 107596 -16657 107650 -16601
rect 107706 -16657 107760 -16601
rect 107816 -16657 107870 -16601
rect 107926 -16657 127459 -16601
rect 107175 -16711 127459 -16657
rect 107175 -16767 107210 -16711
rect 107266 -16767 107320 -16711
rect 107376 -16767 107430 -16711
rect 107486 -16767 107540 -16711
rect 107596 -16767 107650 -16711
rect 107706 -16767 107760 -16711
rect 107816 -16767 107870 -16711
rect 107926 -16767 127459 -16711
rect 107175 -16821 127459 -16767
rect 107175 -16877 107210 -16821
rect 107266 -16877 107320 -16821
rect 107376 -16877 107430 -16821
rect 107486 -16877 107540 -16821
rect 107596 -16877 107650 -16821
rect 107706 -16877 107760 -16821
rect 107816 -16877 107870 -16821
rect 107926 -16877 127459 -16821
rect 107175 -16931 127459 -16877
rect 107175 -16987 107210 -16931
rect 107266 -16987 107320 -16931
rect 107376 -16987 107430 -16931
rect 107486 -16987 107540 -16931
rect 107596 -16987 107650 -16931
rect 107706 -16987 107760 -16931
rect 107816 -16987 107870 -16931
rect 107926 -16987 127459 -16931
rect 28338 -17018 31322 -17012
rect 28339 -17020 31322 -17018
rect 107175 -17023 127459 -16987
rect -832 -17073 22477 -17045
rect -832 -17129 -814 -17073
rect -758 -17129 -704 -17073
rect -648 -17129 -594 -17073
rect -538 -17129 -484 -17073
rect -428 -17129 -374 -17073
rect -318 -17129 -264 -17073
rect -208 -17129 -154 -17073
rect -98 -17099 22477 -17073
rect -98 -17129 21746 -17099
rect -832 -17143 21746 -17129
rect -545 -17155 21746 -17143
rect 21802 -17155 21856 -17099
rect 21912 -17155 21966 -17099
rect 22022 -17155 22076 -17099
rect 22132 -17155 22186 -17099
rect 22242 -17155 22296 -17099
rect 22352 -17155 22406 -17099
rect 22462 -17155 22477 -17099
rect -545 -17163 22477 -17155
rect 107 -17330 876 -17322
rect 106 -17348 16453 -17330
rect 106 -17404 121 -17348
rect 177 -17404 231 -17348
rect 287 -17404 341 -17348
rect 397 -17404 451 -17348
rect 507 -17404 561 -17348
rect 617 -17404 671 -17348
rect 727 -17404 781 -17348
rect 837 -17358 16453 -17348
rect 837 -17404 15724 -17358
rect 106 -17414 15724 -17404
rect 15780 -17414 15834 -17358
rect 15890 -17414 15944 -17358
rect 16000 -17414 16054 -17358
rect 16110 -17414 16164 -17358
rect 16220 -17414 16274 -17358
rect 16330 -17414 16384 -17358
rect 16440 -17414 16453 -17358
rect 30162 -17411 30769 -17390
rect 106 -17458 16453 -17414
rect 106 -17514 121 -17458
rect 177 -17514 231 -17458
rect 287 -17514 341 -17458
rect 397 -17514 451 -17458
rect 507 -17514 561 -17458
rect 617 -17514 671 -17458
rect 727 -17514 781 -17458
rect 837 -17468 16453 -17458
rect 837 -17514 15724 -17468
rect 106 -17524 15724 -17514
rect 15780 -17524 15834 -17468
rect 15890 -17524 15944 -17468
rect 16000 -17524 16054 -17468
rect 16110 -17524 16164 -17468
rect 16220 -17524 16274 -17468
rect 16330 -17524 16384 -17468
rect 16440 -17524 16453 -17468
rect 106 -17568 16453 -17524
rect 106 -17624 121 -17568
rect 177 -17624 231 -17568
rect 287 -17624 341 -17568
rect 397 -17624 451 -17568
rect 507 -17624 561 -17568
rect 617 -17624 671 -17568
rect 727 -17624 781 -17568
rect 837 -17578 16453 -17568
rect 837 -17624 15724 -17578
rect 106 -17634 15724 -17624
rect 15780 -17634 15834 -17578
rect 15890 -17634 15944 -17578
rect 16000 -17634 16054 -17578
rect 16110 -17634 16164 -17578
rect 16220 -17634 16274 -17578
rect 16330 -17634 16384 -17578
rect 16440 -17634 16453 -17578
rect 106 -17678 16453 -17634
rect 106 -17734 121 -17678
rect 177 -17734 231 -17678
rect 287 -17734 341 -17678
rect 397 -17734 451 -17678
rect 507 -17734 561 -17678
rect 617 -17734 671 -17678
rect 727 -17734 781 -17678
rect 837 -17688 16453 -17678
rect 837 -17734 15724 -17688
rect 106 -17744 15724 -17734
rect 15780 -17744 15834 -17688
rect 15890 -17744 15944 -17688
rect 16000 -17744 16054 -17688
rect 16110 -17744 16164 -17688
rect 16220 -17744 16274 -17688
rect 16330 -17744 16384 -17688
rect 16440 -17744 16453 -17688
rect 106 -17788 16453 -17744
rect 106 -17844 121 -17788
rect 177 -17844 231 -17788
rect 287 -17844 341 -17788
rect 397 -17844 451 -17788
rect 507 -17844 561 -17788
rect 617 -17844 671 -17788
rect 727 -17844 781 -17788
rect 837 -17798 16453 -17788
rect 837 -17844 15724 -17798
rect 106 -17854 15724 -17844
rect 15780 -17854 15834 -17798
rect 15890 -17854 15944 -17798
rect 16000 -17854 16054 -17798
rect 16110 -17854 16164 -17798
rect 16220 -17854 16274 -17798
rect 16330 -17854 16384 -17798
rect 16440 -17854 16453 -17798
rect 106 -17898 16453 -17854
rect 22870 -17450 30771 -17411
rect 22870 -17454 23387 -17450
rect 22870 -17510 22902 -17454
rect 22958 -17510 23012 -17454
rect 23068 -17510 23122 -17454
rect 23178 -17510 23232 -17454
rect 23288 -17506 23387 -17454
rect 23443 -17506 23497 -17450
rect 23553 -17506 23607 -17450
rect 23663 -17506 23717 -17450
rect 23773 -17456 30771 -17450
rect 23773 -17506 30249 -17456
rect 23288 -17510 30249 -17506
rect 22870 -17512 30249 -17510
rect 30305 -17512 30359 -17456
rect 30415 -17512 30469 -17456
rect 30525 -17512 30579 -17456
rect 30635 -17512 30771 -17456
rect 22870 -17560 30771 -17512
rect 22870 -17564 23387 -17560
rect 22870 -17620 22902 -17564
rect 22958 -17620 23012 -17564
rect 23068 -17620 23122 -17564
rect 23178 -17620 23232 -17564
rect 23288 -17616 23387 -17564
rect 23443 -17616 23497 -17560
rect 23553 -17616 23607 -17560
rect 23663 -17616 23717 -17560
rect 23773 -17566 30771 -17560
rect 23773 -17616 30249 -17566
rect 23288 -17620 30249 -17616
rect 22870 -17622 30249 -17620
rect 30305 -17622 30359 -17566
rect 30415 -17622 30469 -17566
rect 30525 -17622 30579 -17566
rect 30635 -17622 30771 -17566
rect 22870 -17670 30771 -17622
rect 22870 -17674 23387 -17670
rect 22870 -17730 22902 -17674
rect 22958 -17730 23012 -17674
rect 23068 -17730 23122 -17674
rect 23178 -17730 23232 -17674
rect 23288 -17726 23387 -17674
rect 23443 -17726 23497 -17670
rect 23553 -17726 23607 -17670
rect 23663 -17726 23717 -17670
rect 23773 -17676 30771 -17670
rect 23773 -17726 30249 -17676
rect 23288 -17730 30249 -17726
rect 22870 -17732 30249 -17730
rect 30305 -17732 30359 -17676
rect 30415 -17732 30469 -17676
rect 30525 -17732 30579 -17676
rect 30635 -17732 30771 -17676
rect 22870 -17780 30771 -17732
rect 22870 -17784 23387 -17780
rect 22870 -17840 22902 -17784
rect 22958 -17840 23012 -17784
rect 23068 -17840 23122 -17784
rect 23178 -17840 23232 -17784
rect 23288 -17836 23387 -17784
rect 23443 -17836 23497 -17780
rect 23553 -17836 23607 -17780
rect 23663 -17836 23717 -17780
rect 23773 -17786 30771 -17780
rect 23773 -17836 30249 -17786
rect 23288 -17840 30249 -17836
rect 22870 -17842 30249 -17840
rect 30305 -17842 30359 -17786
rect 30415 -17842 30469 -17786
rect 30525 -17842 30579 -17786
rect 30635 -17842 30771 -17786
rect 22870 -17878 30771 -17842
rect 106 -17954 121 -17898
rect 177 -17954 231 -17898
rect 287 -17954 341 -17898
rect 397 -17954 451 -17898
rect 507 -17954 561 -17898
rect 617 -17954 671 -17898
rect 727 -17954 781 -17898
rect 837 -17908 16453 -17898
rect 837 -17954 15724 -17908
rect 106 -17964 15724 -17954
rect 15780 -17964 15834 -17908
rect 15890 -17964 15944 -17908
rect 16000 -17964 16054 -17908
rect 16110 -17964 16164 -17908
rect 16220 -17964 16274 -17908
rect 16330 -17964 16384 -17908
rect 16440 -17964 16453 -17908
rect 30162 -17957 30769 -17878
rect 106 -18008 16453 -17964
rect 106 -18064 121 -18008
rect 177 -18064 231 -18008
rect 287 -18064 341 -18008
rect 397 -18064 451 -18008
rect 507 -18064 561 -18008
rect 617 -18064 671 -18008
rect 727 -18064 781 -18008
rect 837 -18018 16453 -18008
rect 837 -18064 15724 -18018
rect 106 -18074 15724 -18064
rect 15780 -18074 15834 -18018
rect 15890 -18074 15944 -18018
rect 16000 -18074 16054 -18018
rect 16110 -18074 16164 -18018
rect 16220 -18074 16274 -18018
rect 16330 -18074 16384 -18018
rect 16440 -18074 16453 -18018
rect 106 -18084 16453 -18074
rect 1189 -18275 1952 -18266
rect 1182 -18281 30211 -18275
rect 1182 -18337 1236 -18281
rect 1292 -18337 1346 -18281
rect 1402 -18337 1456 -18281
rect 1512 -18337 1566 -18281
rect 1622 -18337 1676 -18281
rect 1732 -18337 1786 -18281
rect 1842 -18337 1896 -18281
rect 1952 -18335 30211 -18281
rect 1952 -18337 29788 -18335
rect 1182 -18391 29788 -18337
rect 29844 -18391 29898 -18335
rect 29954 -18391 30008 -18335
rect 30064 -18391 30118 -18335
rect 30174 -18391 30211 -18335
rect 1182 -18447 1236 -18391
rect 1292 -18447 1346 -18391
rect 1402 -18447 1456 -18391
rect 1512 -18447 1566 -18391
rect 1622 -18447 1676 -18391
rect 1732 -18447 1786 -18391
rect 1842 -18447 1896 -18391
rect 1952 -18445 30211 -18391
rect 1952 -18447 29788 -18445
rect 1182 -18501 29788 -18447
rect 29844 -18501 29898 -18445
rect 29954 -18501 30008 -18445
rect 30064 -18501 30118 -18445
rect 30174 -18501 30211 -18445
rect 1182 -18557 1236 -18501
rect 1292 -18557 1346 -18501
rect 1402 -18557 1456 -18501
rect 1512 -18557 1566 -18501
rect 1622 -18557 1676 -18501
rect 1732 -18557 1786 -18501
rect 1842 -18557 1896 -18501
rect 1952 -18557 30211 -18501
rect 1182 -18573 30211 -18557
rect 1182 -18611 29782 -18573
rect 1182 -18667 1236 -18611
rect 1292 -18667 1346 -18611
rect 1402 -18667 1456 -18611
rect 1512 -18667 1566 -18611
rect 1622 -18667 1676 -18611
rect 1732 -18667 1786 -18611
rect 1842 -18667 1896 -18611
rect 1952 -18629 29782 -18611
rect 29838 -18629 29892 -18573
rect 29948 -18629 30002 -18573
rect 30058 -18629 30112 -18573
rect 30168 -18629 30211 -18573
rect 31430 -18619 31941 -18617
rect 1952 -18667 30211 -18629
rect 1182 -18683 30211 -18667
rect 1182 -18721 29782 -18683
rect 1182 -18777 1236 -18721
rect 1292 -18777 1346 -18721
rect 1402 -18777 1456 -18721
rect 1512 -18777 1566 -18721
rect 1622 -18777 1676 -18721
rect 1732 -18777 1786 -18721
rect 1842 -18777 1896 -18721
rect 1952 -18739 29782 -18721
rect 29838 -18739 29892 -18683
rect 29948 -18739 30002 -18683
rect 30058 -18739 30112 -18683
rect 30168 -18739 30211 -18683
rect 1952 -18777 30211 -18739
rect 1182 -18793 30211 -18777
rect 1182 -18831 29782 -18793
rect 1182 -18887 1236 -18831
rect 1292 -18887 1346 -18831
rect 1402 -18887 1456 -18831
rect 1512 -18887 1566 -18831
rect 1622 -18887 1676 -18831
rect 1732 -18887 1786 -18831
rect 1842 -18887 1896 -18831
rect 1952 -18849 29782 -18831
rect 29838 -18849 29892 -18793
rect 29948 -18849 30002 -18793
rect 30058 -18849 30112 -18793
rect 30168 -18849 30211 -18793
rect 1952 -18887 30211 -18849
rect 1182 -18903 30211 -18887
rect 1182 -18941 29782 -18903
rect 1182 -18997 1236 -18941
rect 1292 -18997 1346 -18941
rect 1402 -18997 1456 -18941
rect 1512 -18997 1566 -18941
rect 1622 -18997 1676 -18941
rect 1732 -18997 1786 -18941
rect 1842 -18997 1896 -18941
rect 1952 -18959 29782 -18941
rect 29838 -18959 29892 -18903
rect 29948 -18959 30002 -18903
rect 30058 -18959 30112 -18903
rect 30168 -18959 30211 -18903
rect 1952 -18997 30211 -18959
rect 1182 -19029 30211 -18997
rect 31386 -18623 31942 -18619
rect 31386 -18673 34621 -18623
rect 31386 -18729 31488 -18673
rect 31544 -18729 31598 -18673
rect 31654 -18729 31708 -18673
rect 31764 -18729 31818 -18673
rect 31874 -18725 34621 -18673
rect 31874 -18729 34132 -18725
rect 31386 -18781 34132 -18729
rect 34188 -18781 34242 -18725
rect 34298 -18781 34352 -18725
rect 34408 -18781 34462 -18725
rect 34518 -18781 34621 -18725
rect 31386 -18783 34621 -18781
rect 31386 -18839 31488 -18783
rect 31544 -18839 31598 -18783
rect 31654 -18839 31708 -18783
rect 31764 -18839 31818 -18783
rect 31874 -18835 34621 -18783
rect 31874 -18839 34132 -18835
rect 31386 -18891 34132 -18839
rect 34188 -18891 34242 -18835
rect 34298 -18891 34352 -18835
rect 34408 -18891 34462 -18835
rect 34518 -18891 34621 -18835
rect 31386 -18893 34621 -18891
rect 31386 -18949 31488 -18893
rect 31544 -18949 31598 -18893
rect 31654 -18949 31708 -18893
rect 31764 -18949 31818 -18893
rect 31874 -18945 34621 -18893
rect 31874 -18949 34132 -18945
rect 31386 -19001 34132 -18949
rect 34188 -19001 34242 -18945
rect 34298 -19001 34352 -18945
rect 34408 -19001 34462 -18945
rect 34518 -19001 34621 -18945
rect 31386 -19003 34621 -19001
rect 31386 -19059 31488 -19003
rect 31544 -19059 31598 -19003
rect 31654 -19059 31708 -19003
rect 31764 -19059 31818 -19003
rect 31874 -19055 34621 -19003
rect 31874 -19059 34132 -19055
rect 31386 -19111 34132 -19059
rect 34188 -19111 34242 -19055
rect 34298 -19111 34352 -19055
rect 34408 -19111 34462 -19055
rect 34518 -19111 34621 -19055
rect 31386 -19176 34621 -19111
rect 31388 -19184 34621 -19176
rect 94333 -18639 94715 -18638
rect 94333 -18642 94768 -18639
rect 94333 -18675 127319 -18642
rect 94333 -18731 94359 -18675
rect 94415 -18731 94469 -18675
rect 94525 -18731 94579 -18675
rect 94635 -18731 94689 -18675
rect 94745 -18731 127319 -18675
rect 94333 -18785 127319 -18731
rect 94333 -18841 94359 -18785
rect 94415 -18841 94469 -18785
rect 94525 -18841 94579 -18785
rect 94635 -18841 94689 -18785
rect 94745 -18841 127319 -18785
rect 94333 -18895 127319 -18841
rect 94333 -18951 94359 -18895
rect 94415 -18951 94469 -18895
rect 94525 -18951 94579 -18895
rect 94635 -18951 94689 -18895
rect 94745 -18951 127319 -18895
rect 94333 -19005 127319 -18951
rect 94333 -19061 94359 -19005
rect 94415 -19061 94469 -19005
rect 94525 -19061 94579 -19005
rect 94635 -19061 94689 -19005
rect 94745 -19061 127319 -19005
rect 94333 -19115 127319 -19061
rect 94333 -19171 94359 -19115
rect 94415 -19171 94469 -19115
rect 94525 -19171 94579 -19115
rect 94635 -19171 94689 -19115
rect 94745 -19171 127319 -19115
rect 94333 -19225 127319 -19171
rect 94333 -19281 94359 -19225
rect 94415 -19281 94469 -19225
rect 94525 -19281 94579 -19225
rect 94635 -19281 94689 -19225
rect 94745 -19281 127319 -19225
rect 94333 -19335 127319 -19281
rect 94333 -19391 94359 -19335
rect 94415 -19391 94469 -19335
rect 94525 -19391 94579 -19335
rect 94635 -19391 94689 -19335
rect 94745 -19391 127319 -19335
rect 94333 -19430 127319 -19391
rect 94333 -19432 94768 -19430
rect 28768 -19838 29207 -19837
rect 1177 -19871 29207 -19838
rect 1177 -19927 13167 -19871
rect 13223 -19927 13277 -19871
rect 13333 -19927 13387 -19871
rect 13443 -19927 13497 -19871
rect 13553 -19927 13607 -19871
rect 13663 -19927 13717 -19871
rect 13773 -19927 13827 -19871
rect 13883 -19872 29207 -19871
rect 13883 -19927 19494 -19872
rect 1177 -19928 19494 -19927
rect 19550 -19928 19604 -19872
rect 19660 -19928 19714 -19872
rect 19770 -19928 19824 -19872
rect 19880 -19928 19934 -19872
rect 19990 -19928 20044 -19872
rect 20100 -19928 20154 -19872
rect 20210 -19928 29207 -19872
rect 94075 -19873 94510 -19869
rect 1177 -19951 29207 -19928
rect 1177 -19981 28803 -19951
rect 1177 -20037 13167 -19981
rect 13223 -20037 13277 -19981
rect 13333 -20037 13387 -19981
rect 13443 -20037 13497 -19981
rect 13553 -20037 13607 -19981
rect 13663 -20037 13717 -19981
rect 13773 -20037 13827 -19981
rect 13883 -19982 28803 -19981
rect 13883 -20037 19494 -19982
rect 1177 -20038 19494 -20037
rect 19550 -20038 19604 -19982
rect 19660 -20038 19714 -19982
rect 19770 -20038 19824 -19982
rect 19880 -20038 19934 -19982
rect 19990 -20038 20044 -19982
rect 20100 -20038 20154 -19982
rect 20210 -20007 28803 -19982
rect 28859 -20007 28913 -19951
rect 28969 -20007 29023 -19951
rect 29079 -20007 29133 -19951
rect 29189 -20007 29207 -19951
rect 20210 -20038 29207 -20007
rect 1177 -20061 29207 -20038
rect 1177 -20091 28803 -20061
rect 1177 -20147 13167 -20091
rect 13223 -20147 13277 -20091
rect 13333 -20147 13387 -20091
rect 13443 -20147 13497 -20091
rect 13553 -20147 13607 -20091
rect 13663 -20147 13717 -20091
rect 13773 -20147 13827 -20091
rect 13883 -20092 28803 -20091
rect 13883 -20147 19494 -20092
rect 1177 -20148 19494 -20147
rect 19550 -20148 19604 -20092
rect 19660 -20148 19714 -20092
rect 19770 -20148 19824 -20092
rect 19880 -20148 19934 -20092
rect 19990 -20148 20044 -20092
rect 20100 -20148 20154 -20092
rect 20210 -20117 28803 -20092
rect 28859 -20117 28913 -20061
rect 28969 -20117 29023 -20061
rect 29079 -20117 29133 -20061
rect 29189 -20117 29207 -20061
rect 20210 -20148 29207 -20117
rect 1177 -20189 29207 -20148
rect 1177 -20201 28797 -20189
rect 1177 -20257 13167 -20201
rect 13223 -20257 13277 -20201
rect 13333 -20257 13387 -20201
rect 13443 -20257 13497 -20201
rect 13553 -20257 13607 -20201
rect 13663 -20257 13717 -20201
rect 13773 -20257 13827 -20201
rect 13883 -20202 28797 -20201
rect 13883 -20257 19494 -20202
rect 1177 -20258 19494 -20257
rect 19550 -20258 19604 -20202
rect 19660 -20258 19714 -20202
rect 19770 -20258 19824 -20202
rect 19880 -20258 19934 -20202
rect 19990 -20258 20044 -20202
rect 20100 -20258 20154 -20202
rect 20210 -20245 28797 -20202
rect 28853 -20245 28907 -20189
rect 28963 -20245 29017 -20189
rect 29073 -20245 29127 -20189
rect 29183 -20245 29207 -20189
rect 20210 -20258 29207 -20245
rect 1177 -20299 29207 -20258
rect 1177 -20311 28797 -20299
rect 1177 -20367 13167 -20311
rect 13223 -20367 13277 -20311
rect 13333 -20367 13387 -20311
rect 13443 -20367 13497 -20311
rect 13553 -20367 13607 -20311
rect 13663 -20367 13717 -20311
rect 13773 -20367 13827 -20311
rect 13883 -20312 28797 -20311
rect 13883 -20367 19494 -20312
rect 1177 -20368 19494 -20367
rect 19550 -20368 19604 -20312
rect 19660 -20368 19714 -20312
rect 19770 -20368 19824 -20312
rect 19880 -20368 19934 -20312
rect 19990 -20368 20044 -20312
rect 20100 -20368 20154 -20312
rect 20210 -20355 28797 -20312
rect 28853 -20355 28907 -20299
rect 28963 -20355 29017 -20299
rect 29073 -20355 29127 -20299
rect 29183 -20355 29207 -20299
rect 20210 -20368 29207 -20355
rect 1177 -20409 29207 -20368
rect 1177 -20421 28797 -20409
rect 1177 -20477 13167 -20421
rect 13223 -20477 13277 -20421
rect 13333 -20477 13387 -20421
rect 13443 -20477 13497 -20421
rect 13553 -20477 13607 -20421
rect 13663 -20477 13717 -20421
rect 13773 -20477 13827 -20421
rect 13883 -20422 28797 -20421
rect 13883 -20477 19494 -20422
rect 1177 -20478 19494 -20477
rect 19550 -20478 19604 -20422
rect 19660 -20478 19714 -20422
rect 19770 -20478 19824 -20422
rect 19880 -20478 19934 -20422
rect 19990 -20478 20044 -20422
rect 20100 -20478 20154 -20422
rect 20210 -20465 28797 -20422
rect 28853 -20465 28907 -20409
rect 28963 -20465 29017 -20409
rect 29073 -20465 29127 -20409
rect 29183 -20465 29207 -20409
rect 20210 -20478 29207 -20465
rect 1177 -20519 29207 -20478
rect 1177 -20531 28797 -20519
rect 1177 -20587 13167 -20531
rect 13223 -20587 13277 -20531
rect 13333 -20587 13387 -20531
rect 13443 -20587 13497 -20531
rect 13553 -20587 13607 -20531
rect 13663 -20587 13717 -20531
rect 13773 -20587 13827 -20531
rect 13883 -20532 28797 -20531
rect 13883 -20587 19494 -20532
rect 1177 -20588 19494 -20587
rect 19550 -20588 19604 -20532
rect 19660 -20588 19714 -20532
rect 19770 -20588 19824 -20532
rect 19880 -20588 19934 -20532
rect 19990 -20588 20044 -20532
rect 20100 -20588 20154 -20532
rect 20210 -20575 28797 -20532
rect 28853 -20575 28907 -20519
rect 28963 -20575 29017 -20519
rect 29073 -20575 29127 -20519
rect 29183 -20575 29207 -20519
rect 20210 -20588 29207 -20575
rect 1177 -20592 29207 -20588
rect 94074 -19905 127202 -19873
rect 94074 -19961 94101 -19905
rect 94157 -19961 94211 -19905
rect 94267 -19961 94321 -19905
rect 94377 -19961 94431 -19905
rect 94487 -19961 127202 -19905
rect 94074 -20015 127202 -19961
rect 94074 -20071 94101 -20015
rect 94157 -20071 94211 -20015
rect 94267 -20071 94321 -20015
rect 94377 -20071 94431 -20015
rect 94487 -20071 127202 -20015
rect 94074 -20125 127202 -20071
rect 94074 -20181 94101 -20125
rect 94157 -20181 94211 -20125
rect 94267 -20181 94321 -20125
rect 94377 -20181 94431 -20125
rect 94487 -20181 127202 -20125
rect 94074 -20235 127202 -20181
rect 94074 -20291 94101 -20235
rect 94157 -20291 94211 -20235
rect 94267 -20291 94321 -20235
rect 94377 -20291 94431 -20235
rect 94487 -20291 127202 -20235
rect 94074 -20345 127202 -20291
rect 94074 -20401 94101 -20345
rect 94157 -20401 94211 -20345
rect 94267 -20401 94321 -20345
rect 94377 -20401 94431 -20345
rect 94487 -20401 127202 -20345
rect 94074 -20455 127202 -20401
rect 94074 -20511 94101 -20455
rect 94157 -20511 94211 -20455
rect 94267 -20511 94321 -20455
rect 94377 -20511 94431 -20455
rect 94487 -20511 127202 -20455
rect 94074 -20565 127202 -20511
rect 13160 -20593 13888 -20592
rect 19486 -20593 20228 -20592
rect 94074 -20621 94101 -20565
rect 94157 -20621 94211 -20565
rect 94267 -20621 94321 -20565
rect 94377 -20621 94431 -20565
rect 94487 -20621 127202 -20565
rect 94074 -20661 127202 -20621
rect 94075 -20662 94510 -20661
rect 28837 -20718 29216 -20717
rect 28770 -20719 29216 -20718
rect 1117 -20752 29216 -20719
rect 1117 -20757 18599 -20752
rect 1117 -20813 12283 -20757
rect 12339 -20813 12393 -20757
rect 12449 -20813 12503 -20757
rect 12559 -20813 12613 -20757
rect 12669 -20813 12723 -20757
rect 12779 -20813 12833 -20757
rect 12889 -20813 12943 -20757
rect 12999 -20808 18599 -20757
rect 18655 -20808 18709 -20752
rect 18765 -20808 18819 -20752
rect 18875 -20808 18929 -20752
rect 18985 -20808 19039 -20752
rect 19095 -20808 19149 -20752
rect 19205 -20808 19259 -20752
rect 19315 -20805 29216 -20752
rect 19315 -20808 28796 -20805
rect 12999 -20813 28796 -20808
rect 1117 -20861 28796 -20813
rect 28852 -20861 28906 -20805
rect 28962 -20861 29016 -20805
rect 29072 -20861 29126 -20805
rect 29182 -20861 29216 -20805
rect 1117 -20862 29216 -20861
rect 1117 -20867 18599 -20862
rect 1117 -20923 12283 -20867
rect 12339 -20923 12393 -20867
rect 12449 -20923 12503 -20867
rect 12559 -20923 12613 -20867
rect 12669 -20923 12723 -20867
rect 12779 -20923 12833 -20867
rect 12889 -20923 12943 -20867
rect 12999 -20918 18599 -20867
rect 18655 -20918 18709 -20862
rect 18765 -20918 18819 -20862
rect 18875 -20918 18929 -20862
rect 18985 -20918 19039 -20862
rect 19095 -20918 19149 -20862
rect 19205 -20918 19259 -20862
rect 19315 -20915 29216 -20862
rect 19315 -20918 28796 -20915
rect 12999 -20923 28796 -20918
rect 1117 -20971 28796 -20923
rect 28852 -20971 28906 -20915
rect 28962 -20971 29016 -20915
rect 29072 -20971 29126 -20915
rect 29182 -20971 29216 -20915
rect 1117 -20972 29216 -20971
rect 1117 -20977 18599 -20972
rect 1117 -21033 12283 -20977
rect 12339 -21033 12393 -20977
rect 12449 -21033 12503 -20977
rect 12559 -21033 12613 -20977
rect 12669 -21033 12723 -20977
rect 12779 -21033 12833 -20977
rect 12889 -21033 12943 -20977
rect 12999 -21028 18599 -20977
rect 18655 -21028 18709 -20972
rect 18765 -21028 18819 -20972
rect 18875 -21028 18929 -20972
rect 18985 -21028 19039 -20972
rect 19095 -21028 19149 -20972
rect 19205 -21028 19259 -20972
rect 19315 -21028 29216 -20972
rect 12999 -21033 29216 -21028
rect 1117 -21043 29216 -21033
rect 1117 -21082 28790 -21043
rect 1117 -21087 18599 -21082
rect 1117 -21143 12283 -21087
rect 12339 -21143 12393 -21087
rect 12449 -21143 12503 -21087
rect 12559 -21143 12613 -21087
rect 12669 -21143 12723 -21087
rect 12779 -21143 12833 -21087
rect 12889 -21143 12943 -21087
rect 12999 -21138 18599 -21087
rect 18655 -21138 18709 -21082
rect 18765 -21138 18819 -21082
rect 18875 -21138 18929 -21082
rect 18985 -21138 19039 -21082
rect 19095 -21138 19149 -21082
rect 19205 -21138 19259 -21082
rect 19315 -21099 28790 -21082
rect 28846 -21099 28900 -21043
rect 28956 -21099 29010 -21043
rect 29066 -21099 29120 -21043
rect 29176 -21099 29216 -21043
rect 19315 -21138 29216 -21099
rect 12999 -21143 29216 -21138
rect 1117 -21153 29216 -21143
rect 1117 -21192 28790 -21153
rect 1117 -21197 18599 -21192
rect 1117 -21253 12283 -21197
rect 12339 -21253 12393 -21197
rect 12449 -21253 12503 -21197
rect 12559 -21253 12613 -21197
rect 12669 -21253 12723 -21197
rect 12779 -21253 12833 -21197
rect 12889 -21253 12943 -21197
rect 12999 -21248 18599 -21197
rect 18655 -21248 18709 -21192
rect 18765 -21248 18819 -21192
rect 18875 -21248 18929 -21192
rect 18985 -21248 19039 -21192
rect 19095 -21248 19149 -21192
rect 19205 -21248 19259 -21192
rect 19315 -21209 28790 -21192
rect 28846 -21209 28900 -21153
rect 28956 -21209 29010 -21153
rect 29066 -21209 29120 -21153
rect 29176 -21209 29216 -21153
rect 19315 -21248 29216 -21209
rect 12999 -21253 29216 -21248
rect 1117 -21263 29216 -21253
rect 1117 -21302 28790 -21263
rect 1117 -21307 18599 -21302
rect 1117 -21363 12283 -21307
rect 12339 -21363 12393 -21307
rect 12449 -21363 12503 -21307
rect 12559 -21363 12613 -21307
rect 12669 -21363 12723 -21307
rect 12779 -21363 12833 -21307
rect 12889 -21363 12943 -21307
rect 12999 -21358 18599 -21307
rect 18655 -21358 18709 -21302
rect 18765 -21358 18819 -21302
rect 18875 -21358 18929 -21302
rect 18985 -21358 19039 -21302
rect 19095 -21358 19149 -21302
rect 19205 -21358 19259 -21302
rect 19315 -21319 28790 -21302
rect 28846 -21319 28900 -21263
rect 28956 -21319 29010 -21263
rect 29066 -21319 29120 -21263
rect 29176 -21319 29216 -21263
rect 19315 -21358 29216 -21319
rect 12999 -21363 29216 -21358
rect 1117 -21373 29216 -21363
rect 1117 -21412 28790 -21373
rect 1117 -21417 18599 -21412
rect 1117 -21473 12283 -21417
rect 12339 -21473 12393 -21417
rect 12449 -21473 12503 -21417
rect 12559 -21473 12613 -21417
rect 12669 -21473 12723 -21417
rect 12779 -21473 12833 -21417
rect 12889 -21473 12943 -21417
rect 12999 -21468 18599 -21417
rect 18655 -21468 18709 -21412
rect 18765 -21468 18819 -21412
rect 18875 -21468 18929 -21412
rect 18985 -21468 19039 -21412
rect 19095 -21468 19149 -21412
rect 19205 -21468 19259 -21412
rect 19315 -21429 28790 -21412
rect 28846 -21429 28900 -21373
rect 28956 -21429 29010 -21373
rect 29066 -21429 29120 -21373
rect 29176 -21429 29216 -21373
rect 19315 -21468 29216 -21429
rect 12999 -21473 29216 -21468
rect 93809 -20882 127202 -20845
rect 93809 -20938 93836 -20882
rect 93892 -20938 93946 -20882
rect 94002 -20938 94056 -20882
rect 94112 -20938 94166 -20882
rect 94222 -20938 127202 -20882
rect 93809 -20992 127202 -20938
rect 93809 -21048 93836 -20992
rect 93892 -21048 93946 -20992
rect 94002 -21048 94056 -20992
rect 94112 -21048 94166 -20992
rect 94222 -21048 127202 -20992
rect 93809 -21102 127202 -21048
rect 93809 -21158 93836 -21102
rect 93892 -21158 93946 -21102
rect 94002 -21158 94056 -21102
rect 94112 -21158 94166 -21102
rect 94222 -21158 127202 -21102
rect 93809 -21212 127202 -21158
rect 93809 -21268 93836 -21212
rect 93892 -21268 93946 -21212
rect 94002 -21268 94056 -21212
rect 94112 -21268 94166 -21212
rect 94222 -21268 127202 -21212
rect 93809 -21322 127202 -21268
rect 93809 -21378 93836 -21322
rect 93892 -21378 93946 -21322
rect 94002 -21378 94056 -21322
rect 94112 -21378 94166 -21322
rect 94222 -21378 127202 -21322
rect 93809 -21432 127202 -21378
rect 12276 -21479 13004 -21473
rect 93809 -21488 93836 -21432
rect 93892 -21488 93946 -21432
rect 94002 -21488 94056 -21432
rect 94112 -21488 94166 -21432
rect 94222 -21488 127202 -21432
rect 93809 -21542 127202 -21488
rect 93809 -21598 93836 -21542
rect 93892 -21598 93946 -21542
rect 94002 -21598 94056 -21542
rect 94112 -21598 94166 -21542
rect 94222 -21598 127202 -21542
rect 93809 -21633 127202 -21598
rect 93810 -21639 94245 -21633
rect 597 -22685 27773 -22496
rect 597 -22741 27330 -22685
rect 27386 -22741 27440 -22685
rect 27496 -22741 27550 -22685
rect 27606 -22741 27660 -22685
rect 27716 -22741 27773 -22685
rect 597 -22795 27773 -22741
rect 597 -22851 27330 -22795
rect 27386 -22851 27440 -22795
rect 27496 -22851 27550 -22795
rect 27606 -22851 27660 -22795
rect 27716 -22851 27773 -22795
rect 597 -22883 27773 -22851
rect 597 -22923 27775 -22883
rect 597 -22979 27324 -22923
rect 27380 -22979 27434 -22923
rect 27490 -22979 27544 -22923
rect 27600 -22979 27654 -22923
rect 27710 -22979 27775 -22923
rect 597 -23025 27775 -22979
rect 599 -23033 27775 -23025
rect 599 -23089 27324 -23033
rect 27380 -23089 27434 -23033
rect 27490 -23089 27544 -23033
rect 27600 -23089 27654 -23033
rect 27710 -23089 27775 -23033
rect 599 -23143 27775 -23089
rect 599 -23199 27324 -23143
rect 27380 -23199 27434 -23143
rect 27490 -23199 27544 -23143
rect 27600 -23199 27654 -23143
rect 27710 -23199 27775 -23143
rect 599 -23253 27775 -23199
rect 599 -23309 27324 -23253
rect 27380 -23309 27434 -23253
rect 27490 -23309 27544 -23253
rect 27600 -23309 27654 -23253
rect 27710 -23309 27775 -23253
rect 599 -23412 27775 -23309
rect 56571 -27798 57329 -27796
rect 56571 -27818 125315 -27798
rect 56571 -27874 56591 -27818
rect 56647 -27874 56701 -27818
rect 56757 -27874 56811 -27818
rect 56867 -27874 56921 -27818
rect 56977 -27874 57031 -27818
rect 57087 -27874 57141 -27818
rect 57197 -27874 57251 -27818
rect 57307 -27858 125315 -27818
rect 57307 -27874 112129 -27858
rect 56571 -27914 112129 -27874
rect 112185 -27914 112239 -27858
rect 112295 -27914 112349 -27858
rect 112405 -27914 112459 -27858
rect 112515 -27914 112569 -27858
rect 112625 -27914 112679 -27858
rect 112735 -27914 112789 -27858
rect 112845 -27914 125315 -27858
rect 56571 -27928 125315 -27914
rect 56571 -27984 56591 -27928
rect 56647 -27984 56701 -27928
rect 56757 -27984 56811 -27928
rect 56867 -27984 56921 -27928
rect 56977 -27984 57031 -27928
rect 57087 -27984 57141 -27928
rect 57197 -27984 57251 -27928
rect 57307 -27968 125315 -27928
rect 57307 -27984 112129 -27968
rect 56571 -28024 112129 -27984
rect 112185 -28024 112239 -27968
rect 112295 -28024 112349 -27968
rect 112405 -28024 112459 -27968
rect 112515 -28024 112569 -27968
rect 112625 -28024 112679 -27968
rect 112735 -28024 112789 -27968
rect 112845 -28024 125315 -27968
rect 56571 -28038 125315 -28024
rect 56571 -28094 56591 -28038
rect 56647 -28094 56701 -28038
rect 56757 -28094 56811 -28038
rect 56867 -28094 56921 -28038
rect 56977 -28094 57031 -28038
rect 57087 -28094 57141 -28038
rect 57197 -28094 57251 -28038
rect 57307 -28078 125315 -28038
rect 57307 -28094 112129 -28078
rect 56571 -28134 112129 -28094
rect 112185 -28134 112239 -28078
rect 112295 -28134 112349 -28078
rect 112405 -28134 112459 -28078
rect 112515 -28134 112569 -28078
rect 112625 -28134 112679 -28078
rect 112735 -28134 112789 -28078
rect 112845 -28134 125315 -28078
rect 56571 -28148 125315 -28134
rect 56571 -28204 56591 -28148
rect 56647 -28204 56701 -28148
rect 56757 -28204 56811 -28148
rect 56867 -28204 56921 -28148
rect 56977 -28204 57031 -28148
rect 57087 -28204 57141 -28148
rect 57197 -28204 57251 -28148
rect 57307 -28188 125315 -28148
rect 57307 -28204 112129 -28188
rect 56571 -28244 112129 -28204
rect 112185 -28244 112239 -28188
rect 112295 -28244 112349 -28188
rect 112405 -28244 112459 -28188
rect 112515 -28244 112569 -28188
rect 112625 -28244 112679 -28188
rect 112735 -28244 112789 -28188
rect 112845 -28244 125315 -28188
rect 56571 -28258 125315 -28244
rect 56571 -28314 56591 -28258
rect 56647 -28314 56701 -28258
rect 56757 -28314 56811 -28258
rect 56867 -28314 56921 -28258
rect 56977 -28314 57031 -28258
rect 57087 -28314 57141 -28258
rect 57197 -28314 57251 -28258
rect 57307 -28298 125315 -28258
rect 57307 -28314 112129 -28298
rect 56571 -28354 112129 -28314
rect 112185 -28354 112239 -28298
rect 112295 -28354 112349 -28298
rect 112405 -28354 112459 -28298
rect 112515 -28354 112569 -28298
rect 112625 -28354 112679 -28298
rect 112735 -28354 112789 -28298
rect 112845 -28354 125315 -28298
rect 56571 -28368 125315 -28354
rect 56571 -28424 56591 -28368
rect 56647 -28424 56701 -28368
rect 56757 -28424 56811 -28368
rect 56867 -28424 56921 -28368
rect 56977 -28424 57031 -28368
rect 57087 -28424 57141 -28368
rect 57197 -28424 57251 -28368
rect 57307 -28408 125315 -28368
rect 57307 -28424 112129 -28408
rect 56571 -28464 112129 -28424
rect 112185 -28464 112239 -28408
rect 112295 -28464 112349 -28408
rect 112405 -28464 112459 -28408
rect 112515 -28464 112569 -28408
rect 112625 -28464 112679 -28408
rect 112735 -28464 112789 -28408
rect 112845 -28464 125315 -28408
rect 56571 -28478 125315 -28464
rect 56571 -28534 56591 -28478
rect 56647 -28534 56701 -28478
rect 56757 -28534 56811 -28478
rect 56867 -28534 56921 -28478
rect 56977 -28534 57031 -28478
rect 57087 -28534 57141 -28478
rect 57197 -28534 57251 -28478
rect 57307 -28518 125315 -28478
rect 57307 -28534 112129 -28518
rect 56571 -28574 112129 -28534
rect 112185 -28574 112239 -28518
rect 112295 -28574 112349 -28518
rect 112405 -28574 112459 -28518
rect 112515 -28574 112569 -28518
rect 112625 -28574 112679 -28518
rect 112735 -28574 112789 -28518
rect 112845 -28574 125315 -28518
rect 56571 -28588 125315 -28574
rect 56571 -28644 56591 -28588
rect 56647 -28644 56701 -28588
rect 56757 -28644 56811 -28588
rect 56867 -28644 56921 -28588
rect 56977 -28644 57031 -28588
rect 57087 -28644 57141 -28588
rect 57197 -28644 57251 -28588
rect 57307 -28644 125315 -28588
rect 56571 -28698 125315 -28644
rect 56571 -28703 57329 -28698
rect 39287 -28928 40045 -28925
rect 39287 -28947 125315 -28928
rect 39287 -29003 39307 -28947
rect 39363 -29003 39417 -28947
rect 39473 -29003 39527 -28947
rect 39583 -29003 39637 -28947
rect 39693 -29003 39747 -28947
rect 39803 -29003 39857 -28947
rect 39913 -29003 39967 -28947
rect 40023 -29003 125315 -28947
rect 39287 -29024 125315 -29003
rect 39287 -29057 110768 -29024
rect 39287 -29113 39307 -29057
rect 39363 -29113 39417 -29057
rect 39473 -29113 39527 -29057
rect 39583 -29113 39637 -29057
rect 39693 -29113 39747 -29057
rect 39803 -29113 39857 -29057
rect 39913 -29113 39967 -29057
rect 40023 -29080 110768 -29057
rect 110824 -29080 110878 -29024
rect 110934 -29080 110988 -29024
rect 111044 -29080 111098 -29024
rect 111154 -29080 111208 -29024
rect 111264 -29080 111318 -29024
rect 111374 -29080 111428 -29024
rect 111484 -29080 125315 -29024
rect 40023 -29113 125315 -29080
rect 39287 -29134 125315 -29113
rect 39287 -29167 110768 -29134
rect 39287 -29223 39307 -29167
rect 39363 -29223 39417 -29167
rect 39473 -29223 39527 -29167
rect 39583 -29223 39637 -29167
rect 39693 -29223 39747 -29167
rect 39803 -29223 39857 -29167
rect 39913 -29223 39967 -29167
rect 40023 -29190 110768 -29167
rect 110824 -29190 110878 -29134
rect 110934 -29190 110988 -29134
rect 111044 -29190 111098 -29134
rect 111154 -29190 111208 -29134
rect 111264 -29190 111318 -29134
rect 111374 -29190 111428 -29134
rect 111484 -29190 125315 -29134
rect 40023 -29223 125315 -29190
rect 39287 -29244 125315 -29223
rect 39287 -29277 110768 -29244
rect 39287 -29333 39307 -29277
rect 39363 -29333 39417 -29277
rect 39473 -29333 39527 -29277
rect 39583 -29333 39637 -29277
rect 39693 -29333 39747 -29277
rect 39803 -29333 39857 -29277
rect 39913 -29333 39967 -29277
rect 40023 -29300 110768 -29277
rect 110824 -29300 110878 -29244
rect 110934 -29300 110988 -29244
rect 111044 -29300 111098 -29244
rect 111154 -29300 111208 -29244
rect 111264 -29300 111318 -29244
rect 111374 -29300 111428 -29244
rect 111484 -29300 125315 -29244
rect 40023 -29333 125315 -29300
rect 39287 -29354 125315 -29333
rect 39287 -29387 110768 -29354
rect 39287 -29443 39307 -29387
rect 39363 -29443 39417 -29387
rect 39473 -29443 39527 -29387
rect 39583 -29443 39637 -29387
rect 39693 -29443 39747 -29387
rect 39803 -29443 39857 -29387
rect 39913 -29443 39967 -29387
rect 40023 -29410 110768 -29387
rect 110824 -29410 110878 -29354
rect 110934 -29410 110988 -29354
rect 111044 -29410 111098 -29354
rect 111154 -29410 111208 -29354
rect 111264 -29410 111318 -29354
rect 111374 -29410 111428 -29354
rect 111484 -29410 125315 -29354
rect 40023 -29443 125315 -29410
rect 39287 -29464 125315 -29443
rect 39287 -29497 110768 -29464
rect 39287 -29553 39307 -29497
rect 39363 -29553 39417 -29497
rect 39473 -29553 39527 -29497
rect 39583 -29553 39637 -29497
rect 39693 -29553 39747 -29497
rect 39803 -29553 39857 -29497
rect 39913 -29553 39967 -29497
rect 40023 -29520 110768 -29497
rect 110824 -29520 110878 -29464
rect 110934 -29520 110988 -29464
rect 111044 -29520 111098 -29464
rect 111154 -29520 111208 -29464
rect 111264 -29520 111318 -29464
rect 111374 -29520 111428 -29464
rect 111484 -29520 125315 -29464
rect 40023 -29553 125315 -29520
rect 39287 -29574 125315 -29553
rect 39287 -29607 110768 -29574
rect 39287 -29663 39307 -29607
rect 39363 -29663 39417 -29607
rect 39473 -29663 39527 -29607
rect 39583 -29663 39637 -29607
rect 39693 -29663 39747 -29607
rect 39803 -29663 39857 -29607
rect 39913 -29663 39967 -29607
rect 40023 -29630 110768 -29607
rect 110824 -29630 110878 -29574
rect 110934 -29630 110988 -29574
rect 111044 -29630 111098 -29574
rect 111154 -29630 111208 -29574
rect 111264 -29630 111318 -29574
rect 111374 -29630 111428 -29574
rect 111484 -29630 125315 -29574
rect 40023 -29663 125315 -29630
rect 39287 -29684 125315 -29663
rect 39287 -29717 110768 -29684
rect 39287 -29773 39307 -29717
rect 39363 -29773 39417 -29717
rect 39473 -29773 39527 -29717
rect 39583 -29773 39637 -29717
rect 39693 -29773 39747 -29717
rect 39803 -29773 39857 -29717
rect 39913 -29773 39967 -29717
rect 40023 -29740 110768 -29717
rect 110824 -29740 110878 -29684
rect 110934 -29740 110988 -29684
rect 111044 -29740 111098 -29684
rect 111154 -29740 111208 -29684
rect 111264 -29740 111318 -29684
rect 111374 -29740 111428 -29684
rect 111484 -29740 125315 -29684
rect 40023 -29773 125315 -29740
rect 39287 -29828 125315 -29773
rect 39287 -29832 40045 -29828
use 200_ohm_magic  200_ohm_magic_0
timestamp 1695102876
transform 0 -1 4473 1 0 -1241
box -260 -1592 3252 1626
use BIASING_1m_MAGIC  BIASING_1m_MAGIC_0
timestamp 1699967350
transform 1 0 14991 0 1 -28424
box -707 -1300 3491 4009
use BIASING_1m_MAGIC  BIASING_1m_MAGIC_1
timestamp 1699967350
transform 1 0 21019 0 1 -28424
box -707 -1300 3491 4009
use BIASING_CURRENT_MAGIC  BIASING_CURRENT_MAGIC_0
timestamp 1699939503
transform 1 0 29725 0 1 -20510
box -680 -1110 2693 998
use Filter_magic  Filter_magic_0
timestamp 1699872198
transform 1 0 44237 0 1 887
box -16674 0 67702 15718
use fold_cascode_opamp_mag  fold_cascode_opamp_mag_0
timestamp 1699707096
transform 1 0 7207 0 1 -4352
box -4063 -11248 17072 1731
use fold_cascode_opamp_mag  fold_cascode_opamp_mag_1
timestamp 1699707096
transform 1 0 7287 0 1 14051
box -4063 -11248 17072 1731
use MUX_1x8  MUX_1x8_0
timestamp 1698660008
transform -1 0 124030 0 1 -5401
box -5382 -7753 7936 2749
use MUX_1x8  MUX_1x8_1
timestamp 1698660008
transform -1 0 124135 0 1 9848
box -5382 -7753 7936 2749
use PGA_MAGIC  PGA_MAGIC_0
timestamp 1699683674
transform 1 0 34513 0 1 -8642
box -1790 -18792 67202 6560
use VCM_1.3V_magic  VCM_1.3V_magic_0
timestamp 1699891908
transform 1 0 29970 0 1 -4601
box -320 -320 2313 2408
use VCM_1.6_MAGIC  VCM_1.6_MAGIC_0
timestamp 1699896181
transform 1 0 29766 0 1 -15886
box -260 -260 2668 2179
<< labels >>
flabel metal1 131064 8868 131064 8869 0 FreeSans 3200 0 0 0 A0
port 0 nsew
flabel metal1 130927 4258 130927 4258 0 FreeSans 3200 0 0 0 A1
port 1 nsew
flabel metal1 130943 3706 130943 3706 0 FreeSans 3200 0 0 0 A5
port 2 nsew
flabel metal1 130963 5778 130963 5778 0 FreeSans 3200 0 0 0 A3
port 3 nsew
flabel metal1 130989 6444 130989 6444 0 FreeSans 3200 0 0 0 A7
port 4 nsew
flabel metal1 131037 8360 131037 8360 0 FreeSans 3200 0 0 0 A4
port 5 nsew
flabel metal1 131119 10464 131119 10464 0 FreeSans 3200 0 0 0 A2
port 6 nsew
flabel metal1 131041 10951 131041 10951 0 FreeSans 3200 0 0 0 A6
port 7 nsew
flabel metal1 130941 -4271 130941 -4271 0 FreeSans 3200 0 0 0 A6_B
port 8 nsew
flabel metal1 130930 -4798 130930 -4798 0 FreeSans 3200 0 0 0 A2_B
port 9 nsew
flabel metal1 130918 -6354 130918 -6354 0 FreeSans 3200 0 0 0 A0_B
port 10 nsew
flabel metal1 130988 -6908 130988 -6908 0 FreeSans 3200 0 0 0 A4_B
port 11 nsew
flabel metal1 130965 -8750 130965 -8750 0 FreeSans 3200 0 0 0 A7_B
port 12 nsew
flabel metal1 130946 -9427 130946 -9427 0 FreeSans 3200 0 0 0 A3_B
port 14 nsew
flabel metal1 130992 -11018 130992 -11018 0 FreeSans 3200 0 0 0 A1_B
port 15 nsew
flabel via2 130698 2568 130698 2568 0 FreeSans 3200 0 0 0 S2
port 17 nsew
flabel via2 130344 1901 130347 1901 0 FreeSans 3200 0 0 0 S1
port 18 nsew
flabel metal2 129985 1234 129985 1234 0 FreeSans 3200 0 0 0 S0
port 19 nsew
flabel metal2 129661 713 129661 713 0 FreeSans 3200 0 0 0 ENA
port 20 nsew
flabel metal1 472 2571 472 2571 0 FreeSans 3200 0 0 0 IN_P
port 27 nsew
flabel metal1 398 -2410 398 -2396 0 FreeSans 3200 0 0 0 IN_N
port 29 nsew
flabel metal2 1555 -15000 1555 -15000 0 FreeSans 3200 0 0 0 IBIAS
port 30 nsew
flabel metal1 48452 19431 48452 19431 0 FreeSans 4800 0 0 0 VDD
port 32 nsew
flabel metal1 48033 18338 48033 18338 0 FreeSans 4800 0 0 0 VSS
port 33 nsew
flabel metal3 1531 -20370 1531 -20370 0 FreeSans 4800 0 0 0 G_SINK_UP
port 35 nsew
flabel metal3 1548 -21230 1548 -21230 0 FreeSans 4800 0 0 0 G_SINK_DOWN
port 37 nsew
flabel metal3 96810 -18982 96810 -18982 0 FreeSans 4800 0 0 0 S_PGA_1
port 38 nsew
flabel metal3 96527 -20223 96527 -20223 0 FreeSans 4800 0 0 0 S_PGA_2
port 39 nsew
flabel metal3 96400 -21365 96400 -21365 0 FreeSans 4800 0 0 0 S_PGA_3
port 40 nsew
flabel metal3 126769 -15274 126790 -15274 0 FreeSans 4800 0 0 0 PGA_P_T
port 41 nsew
flabel metal3 126238 -16739 126259 -16739 0 FreeSans 4800 0 0 0 PGA_N_T
port 42 nsew
flabel metal3 124726 -28329 124726 -28329 0 FreeSans 4800 0 0 0 FIL_P_T
port 43 nsew
flabel metal3 124554 -29567 124554 -29567 0 FreeSans 4800 0 0 0 FIL_N_T
port 44 nsew
flabel metal1 131002 -11540 131002 -11540 0 FreeSans 3200 0 0 0 A5_B
port 16 nsew
flabel metal3 2004 17239 2004 17239 0 FreeSans 4800 0 0 0 IV_P_T
port 47 nsew
flabel metal3 1098 -23041 1098 -23041 0 FreeSans 4800 0 0 0 IV_N_T
port 48 nsew
<< end >>
