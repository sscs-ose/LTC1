* NGSPICE file created from pll_4_mag.ext - technology: gf180mcuC

.subckt pmos_3p3_MDMPD7 a_2804_n628# a_n968_24# a_n1784_24# a_152_68# a_1784_n628#
+ a_1072_24# a_n868_n628# a_356_n628# a_n1888_n628# a_2396_68# a_n2600_24# a_664_n672#
+ a_n256_68# a_868_24# a_n1072_68# a_764_68# a_560_n628# a_1684_24# a_n1376_24# a_n764_n672#
+ a_n52_68# a_1580_68# a_n2804_n672# a_2396_n628# a_52_24# a_n1784_n672# a_1376_n628#
+ a_2500_24# a_n868_68# a_n1684_68# a_2704_n672# a_n1988_24# a_356_68# a_1684_n672#
+ a_n2192_24# a_1276_24# a_256_n672# a_2600_n628# a_n2500_68# a_1172_68# a_1580_n628#
+ a_n664_n628# a_n2396_n672# a_152_n628# a_n2704_n628# a_n1684_n628# a_n560_24# a_n2804_24#
+ a_n356_n672# a_n1276_68# a_n1376_n672# a_460_n672# a_968_68# a_968_n628# a_1888_24#
+ a_2092_24# a_1784_68# a_2296_n672# a_n560_n672# a_2192_n628# a_460_24# a_n2600_n672#
+ a_1276_n672# a_2704_24# a_n1888_68# a_n1580_n672# a_n2092_68# a_n152_24# a_n2296_n628#
+ w_n2978_n758# a_2600_68# a_1172_n628# a_n256_n628# a_n2396_24# a_n1276_n628# a_2500_n672#
+ a_n2704_68# a_n460_68# a_1376_68# a_1480_n672# a_1988_n628# a_n764_24# a_n460_n628#
+ a_n1580_24# a_n2192_n672# a_52_n672# a_n2500_n628# a_n1480_n628# a_n152_n672# a_868_n672#
+ a_2296_24# a_1988_68# a_n1172_n672# a_2192_68# a_764_n628# a_2092_n672# a_664_24#
+ a_n968_n672# a_n2892_68# a_560_68# a_n2296_68# a_n1988_n672# a_n356_24# a_1480_24#
+ a_2804_68# a_n1172_24# a_1072_n672# a_n2092_n628# a_n664_68# a_n1480_68# a_n2892_n628#
+ a_1888_n672# a_n1072_n628# a_n52_n628# a_256_24#
X0 a_1172_68# a_1072_24# a_968_68# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1 a_2192_68# a_2092_24# a_1988_68# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X2 a_n256_n628# a_n356_n672# a_n460_n628# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X3 a_n1276_n628# a_n1376_n672# a_n1480_n628# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X4 a_1376_n628# a_1276_n672# a_1172_n628# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X5 a_356_n628# a_256_n672# a_152_n628# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X6 a_n1276_68# a_n1376_24# a_n1480_68# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X7 a_n664_68# a_n764_24# a_n868_68# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X8 a_968_68# a_868_24# a_764_68# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X9 a_1580_68# a_1480_24# a_1376_68# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X10 a_n2296_68# a_n2396_24# a_n2500_68# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X11 a_2600_68# a_2500_24# a_2396_68# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X12 a_n664_n628# a_n764_n672# a_n868_n628# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X13 a_n460_68# a_n560_24# a_n664_68# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X14 a_n1684_n628# a_n1784_n672# a_n1888_n628# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X15 a_152_n628# a_52_n672# a_n52_n628# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X16 a_1784_n628# a_1684_n672# a_1580_n628# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X17 a_1376_68# a_1276_24# a_1172_68# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X18 a_n2704_n628# a_n2804_n672# a_n2892_n628# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=1.232p ps=6.48u w=2.8u l=0.5u
X19 a_764_n628# a_664_n672# a_560_n628# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X20 a_2804_n628# a_2704_n672# a_2600_n628# w_n2978_n758# pfet_03v3 ad=1.232p pd=6.48u as=0.728p ps=3.32u w=2.8u l=0.5u
X21 a_n1684_68# a_n1784_24# a_n1888_68# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X22 a_2396_68# a_2296_24# a_2192_68# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X23 a_n2296_n628# a_n2396_n672# a_n2500_n628# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X24 a_2396_n628# a_2296_n672# a_2192_n628# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X25 a_n2704_68# a_n2804_24# a_n2892_68# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=1.232p ps=6.48u w=2.8u l=0.5u
X26 a_n1480_68# a_n1580_24# a_n1684_68# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X27 a_n868_68# a_n968_24# a_n1072_68# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X28 a_560_68# a_460_24# a_356_68# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X29 a_n460_n628# a_n560_n672# a_n664_n628# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X30 a_152_68# a_52_24# a_n52_68# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X31 a_1784_68# a_1684_24# a_1580_68# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X32 a_n1480_n628# a_n1580_n672# a_n1684_n628# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X33 a_n52_n628# a_n152_n672# a_n256_n628# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X34 a_n2500_68# a_n2600_24# a_n2704_68# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X35 a_2804_68# a_2704_24# a_2600_68# w_n2978_n758# pfet_03v3 ad=1.232p pd=6.48u as=0.728p ps=3.32u w=2.8u l=0.5u
X36 a_n1072_n628# a_n1172_n672# a_n1276_n628# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X37 a_1172_n628# a_1072_n672# a_968_n628# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X38 a_n52_68# a_n152_24# a_n256_68# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X39 a_356_68# a_256_24# a_152_68# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X40 a_n1888_68# a_n1988_24# a_n2092_68# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X41 a_n868_n628# a_n968_n672# a_n1072_n628# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X42 a_n1888_n628# a_n1988_n672# a_n2092_n628# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X43 a_1988_n628# a_1888_n672# a_1784_n628# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X44 a_n1072_68# a_n1172_24# a_n1276_68# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X45 a_1580_n628# a_1480_n672# a_1376_n628# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X46 a_764_68# a_664_24# a_560_68# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X47 a_n2500_n628# a_n2600_n672# a_n2704_n628# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X48 a_560_n628# a_460_n672# a_356_n628# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X49 a_968_n628# a_868_n672# a_764_n628# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X50 a_2600_n628# a_2500_n672# a_2396_n628# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X51 a_n2092_68# a_n2192_24# a_n2296_68# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X52 a_1988_68# a_1888_24# a_1784_68# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X53 a_n2092_n628# a_n2192_n672# a_n2296_n628# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X54 a_2192_n628# a_2092_n672# a_1988_n628# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X55 a_n256_68# a_n356_24# a_n460_68# w_n2978_n758# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
.ends

.subckt pmos_3p3_PPZSL5 a_n256_n280# a_52_n324# a_n460_n280# a_n152_n324# a_764_n280#
+ a_n52_n280# a_n852_n280# a_356_n280# a_664_n324# a_560_n280# a_n764_n324# a_256_n324#
+ w_n938_n410# a_152_n280# a_n664_n280# a_n356_n324# a_460_n324# a_n560_n324#
X0 a_560_n280# a_460_n324# a_356_n280# w_n938_n410# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1 a_n256_n280# a_n356_n324# a_n460_n280# w_n938_n410# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X2 a_356_n280# a_256_n324# a_152_n280# w_n938_n410# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X3 a_n664_n280# a_n764_n324# a_n852_n280# w_n938_n410# pfet_03v3 ad=0.728p pd=3.32u as=1.232p ps=6.48u w=2.8u l=0.5u
X4 a_152_n280# a_52_n324# a_n52_n280# w_n938_n410# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X5 a_764_n280# a_664_n324# a_560_n280# w_n938_n410# pfet_03v3 ad=1.232p pd=6.48u as=0.728p ps=3.32u w=2.8u l=0.5u
X6 a_n460_n280# a_n560_n324# a_n664_n280# w_n938_n410# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X7 a_n52_n280# a_n152_n324# a_n256_n280# w_n938_n410# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
.ends

.subckt nmos_3p3_JEEAMQ a_n256_n280# a_52_n324# a_n460_n280# a_n152_n324# a_764_n280#
+ a_n52_n280# a_n852_n280# a_356_n280# a_664_n324# a_560_n280# a_n764_n324# a_256_n324#
+ a_152_n280# a_n664_n280# a_n356_n324# a_460_n324# a_n560_n324# VSUBS
X0 a_560_n280# a_460_n324# a_356_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1 a_n256_n280# a_n356_n324# a_n460_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X2 a_356_n280# a_256_n324# a_152_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X3 a_n664_n280# a_n764_n324# a_n852_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=1.232p ps=6.48u w=2.8u l=0.5u
X4 a_152_n280# a_52_n324# a_n52_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X5 a_764_n280# a_664_n324# a_560_n280# VSUBS nfet_03v3 ad=1.232p pd=6.48u as=0.728p ps=3.32u w=2.8u l=0.5u
X6 a_n460_n280# a_n560_n324# a_n664_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X7 a_n52_n280# a_n152_n324# a_n256_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
.ends

.subckt pmos_3p3_MV44E7 a_n256_n280# a_n1276_n280# a_1480_n324# a_52_n324# a_n460_n280#
+ a_868_n324# a_n152_n324# a_n1480_n280# a_n1172_n324# a_764_n280# a_n968_n324# a_1072_n324#
+ a_n1668_n280# a_n52_n280# a_n1072_n280# a_356_n280# a_n868_n280# a_664_n324# a_560_n280#
+ a_n764_n324# w_n1754_n410# a_1376_n280# a_256_n324# a_1580_n280# a_152_n280# a_n664_n280#
+ a_n356_n324# a_460_n324# a_n1376_n324# a_968_n280# a_1276_n324# a_n560_n324# a_n1580_n324#
+ a_1172_n280#
X0 a_n868_n280# a_n968_n324# a_n1072_n280# w_n1754_n410# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1 a_1580_n280# a_1480_n324# a_1376_n280# w_n1754_n410# pfet_03v3 ad=1.232p pd=6.48u as=0.728p ps=3.32u w=2.8u l=0.5u
X2 a_560_n280# a_460_n324# a_356_n280# w_n1754_n410# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X3 a_968_n280# a_868_n324# a_764_n280# w_n1754_n410# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X4 a_n256_n280# a_n356_n324# a_n460_n280# w_n1754_n410# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X5 a_n1276_n280# a_n1376_n324# a_n1480_n280# w_n1754_n410# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X6 a_1376_n280# a_1276_n324# a_1172_n280# w_n1754_n410# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X7 a_356_n280# a_256_n324# a_152_n280# w_n1754_n410# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X8 a_n664_n280# a_n764_n324# a_n868_n280# w_n1754_n410# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X9 a_152_n280# a_52_n324# a_n52_n280# w_n1754_n410# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X10 a_764_n280# a_664_n324# a_560_n280# w_n1754_n410# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X11 a_n460_n280# a_n560_n324# a_n664_n280# w_n1754_n410# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X12 a_n52_n280# a_n152_n324# a_n256_n280# w_n1754_n410# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X13 a_n1480_n280# a_n1580_n324# a_n1668_n280# w_n1754_n410# pfet_03v3 ad=0.728p pd=3.32u as=1.232p ps=6.48u w=2.8u l=0.5u
X14 a_n1072_n280# a_n1172_n324# a_n1276_n280# w_n1754_n410# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X15 a_1172_n280# a_1072_n324# a_968_n280# w_n1754_n410# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
.ends

.subckt nmos_3p3_7NPLVN a_n256_n280# a_n1276_n280# a_2500_n324# a_1480_n324# a_1988_n280#
+ a_52_n324# a_n2192_n324# a_n460_n280# a_868_n324# a_n152_n324# a_n1480_n280# a_n2500_n280#
+ a_n1172_n324# a_2092_n324# a_764_n280# a_n968_n324# a_1072_n324# a_n1988_n324# a_n2092_n280#
+ a_1888_n324# a_n2892_n280# a_2804_n280# a_n52_n280# a_n1072_n280# a_1784_n280# a_356_n280#
+ a_n868_n280# a_n1888_n280# a_664_n324# a_560_n280# a_n764_n324# a_n2804_n324# a_2396_n280#
+ a_n1784_n324# a_1376_n280# a_2704_n324# a_1684_n324# a_256_n324# a_n2396_n324# a_2600_n280#
+ a_1580_n280# a_152_n280# a_n664_n280# a_n356_n324# a_n1684_n280# a_n2704_n280# a_460_n324#
+ a_n1376_n324# a_2296_n324# a_968_n280# a_1276_n324# a_n560_n324# a_n2600_n324# a_2192_n280#
+ a_n1580_n324# a_1172_n280# a_n2296_n280# VSUBS
X0 a_n868_n280# a_n968_n324# a_n1072_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1 a_n1888_n280# a_n1988_n324# a_n2092_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X2 a_1988_n280# a_1888_n324# a_1784_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X3 a_1580_n280# a_1480_n324# a_1376_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X4 a_968_n280# a_868_n324# a_764_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X5 a_n2500_n280# a_n2600_n324# a_n2704_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X6 a_n2092_n280# a_n2192_n324# a_n2296_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X7 a_560_n280# a_460_n324# a_356_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X8 a_2192_n280# a_2092_n324# a_1988_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X9 a_2600_n280# a_2500_n324# a_2396_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X10 a_n256_n280# a_n356_n324# a_n460_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X11 a_n1276_n280# a_n1376_n324# a_n1480_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X12 a_1376_n280# a_1276_n324# a_1172_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X13 a_356_n280# a_256_n324# a_152_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X14 a_n664_n280# a_n764_n324# a_n868_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X15 a_152_n280# a_52_n324# a_n52_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X16 a_n1684_n280# a_n1784_n324# a_n1888_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X17 a_1784_n280# a_1684_n324# a_1580_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X18 a_764_n280# a_664_n324# a_560_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X19 a_2804_n280# a_2704_n324# a_2600_n280# VSUBS nfet_03v3 ad=1.232p pd=6.48u as=0.728p ps=3.32u w=2.8u l=0.5u
X20 a_n2704_n280# a_n2804_n324# a_n2892_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=1.232p ps=6.48u w=2.8u l=0.5u
X21 a_n2296_n280# a_n2396_n324# a_n2500_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X22 a_2396_n280# a_2296_n324# a_2192_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X23 a_n460_n280# a_n560_n324# a_n664_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X24 a_n52_n280# a_n152_n324# a_n256_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X25 a_n1480_n280# a_n1580_n324# a_n1684_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X26 a_n1072_n280# a_n1172_n324# a_n1276_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X27 a_1172_n280# a_1072_n324# a_968_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
.ends

.subckt pmos_3p3_PPYSL5 a_n256_n280# a_52_n324# a_n152_n324# a_n52_n280# a_356_n280#
+ w_n530_n410# a_n444_n280# a_256_n324# a_152_n280# a_n356_n324#
X0 a_n256_n280# a_n356_n324# a_n444_n280# w_n530_n410# pfet_03v3 ad=0.728p pd=3.32u as=1.232p ps=6.48u w=2.8u l=0.5u
X1 a_356_n280# a_256_n324# a_152_n280# w_n530_n410# pfet_03v3 ad=1.232p pd=6.48u as=0.728p ps=3.32u w=2.8u l=0.5u
X2 a_152_n280# a_52_n324# a_n52_n280# w_n530_n410# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X3 a_n52_n280# a_n152_n324# a_n256_n280# w_n530_n410# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
.ends

.subckt nmos_3p3_PLQLVN a_n256_n280# a_n1276_n280# a_1480_n324# a_52_n324# a_n460_n280#
+ a_868_n324# a_n152_n324# a_n1480_n280# a_n1172_n324# a_764_n280# a_n968_n324# a_1072_n324#
+ a_n52_n280# a_n1072_n280# a_1784_n280# a_356_n280# a_n868_n280# a_n1872_n280# a_664_n324#
+ a_560_n280# a_n764_n324# a_n1784_n324# a_1376_n280# a_1684_n324# a_256_n324# a_1580_n280#
+ a_152_n280# a_n664_n280# a_n356_n324# a_n1684_n280# a_460_n324# a_n1376_n324# a_968_n280#
+ a_1276_n324# a_n560_n324# a_n1580_n324# a_1172_n280# VSUBS
X0 a_n868_n280# a_n968_n324# a_n1072_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1 a_1580_n280# a_1480_n324# a_1376_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X2 a_968_n280# a_868_n324# a_764_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X3 a_560_n280# a_460_n324# a_356_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X4 a_n256_n280# a_n356_n324# a_n460_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X5 a_n1276_n280# a_n1376_n324# a_n1480_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X6 a_1376_n280# a_1276_n324# a_1172_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X7 a_356_n280# a_256_n324# a_152_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X8 a_n664_n280# a_n764_n324# a_n868_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X9 a_152_n280# a_52_n324# a_n52_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X10 a_n1684_n280# a_n1784_n324# a_n1872_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=1.232p ps=6.48u w=2.8u l=0.5u
X11 a_1784_n280# a_1684_n324# a_1580_n280# VSUBS nfet_03v3 ad=1.232p pd=6.48u as=0.728p ps=3.32u w=2.8u l=0.5u
X12 a_764_n280# a_664_n324# a_560_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X13 a_n460_n280# a_n560_n324# a_n664_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X14 a_n52_n280# a_n152_n324# a_n256_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X15 a_n1480_n280# a_n1580_n324# a_n1684_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X16 a_n1072_n280# a_n1172_n324# a_n1276_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X17 a_1172_n280# a_1072_n324# a_968_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
.ends

.subckt nmos_3p3_8FEAMQ a_52_n324# a_n152_n324# a_n52_n280# a_152_n280# a_n240_n280#
+ VSUBS
X0 a_152_n280# a_52_n324# a_n52_n280# VSUBS nfet_03v3 ad=1.232p pd=6.48u as=0.728p ps=3.32u w=2.8u l=0.5u
X1 a_n52_n280# a_n152_n324# a_n240_n280# VSUBS nfet_03v3 ad=0.728p pd=3.32u as=1.232p ps=6.48u w=2.8u l=0.5u
.ends

.subckt Tappered_Buffer VDD IN OUT VSS
Xpmos_3p3_MDMPD7_0 VDD a_4254_n29# a_4254_n29# OUT OUT a_4254_n29# VDD VDD OUT VDD
+ a_4254_n29# a_4254_n29# OUT a_4254_n29# OUT VDD OUT a_4254_n29# a_4254_n29# a_4254_n29#
+ VDD VDD a_4254_n29# VDD a_4254_n29# a_4254_n29# OUT a_4254_n29# VDD VDD a_4254_n29#
+ a_4254_n29# VDD a_4254_n29# a_4254_n29# a_4254_n29# a_4254_n29# OUT VDD VDD VDD
+ OUT a_4254_n29# OUT OUT VDD a_4254_n29# a_4254_n29# a_4254_n29# VDD a_4254_n29#
+ a_4254_n29# OUT OUT a_4254_n29# a_4254_n29# OUT a_4254_n29# a_4254_n29# OUT a_4254_n29#
+ a_4254_n29# a_4254_n29# a_4254_n29# OUT a_4254_n29# VDD a_4254_n29# OUT VDD OUT
+ VDD OUT a_4254_n29# VDD a_4254_n29# OUT VDD OUT a_4254_n29# VDD a_4254_n29# VDD
+ a_4254_n29# a_4254_n29# a_4254_n29# VDD OUT a_4254_n29# a_4254_n29# a_4254_n29#
+ VDD a_4254_n29# OUT VDD a_4254_n29# a_4254_n29# a_4254_n29# VDD OUT OUT a_4254_n29#
+ a_4254_n29# a_4254_n29# VDD a_4254_n29# a_4254_n29# VDD OUT OUT VDD a_4254_n29#
+ OUT VDD a_4254_n29# pmos_3p3_MDMPD7
Xpmos_3p3_PPZSL5_0 OUT a_4254_n29# VDD a_4254_n29# VDD VDD VDD VDD a_4254_n29# OUT
+ a_4254_n29# a_4254_n29# VDD OUT OUT a_4254_n29# a_4254_n29# a_4254_n29# pmos_3p3_PPZSL5
Xnmos_3p3_JEEAMQ_0 a_4254_n29# a_548_n1560# VSS a_548_n1560# VSS VSS VSS VSS a_548_n1560#
+ a_4254_n29# a_548_n1560# a_548_n1560# a_4254_n29# a_4254_n29# a_548_n1560# a_548_n1560#
+ a_548_n1560# VSS nmos_3p3_JEEAMQ
Xpmos_3p3_MV44E7_0 a_4254_n29# VDD a_548_n1560# a_548_n1560# VDD a_548_n1560# a_548_n1560#
+ a_4254_n29# a_548_n1560# VDD a_548_n1560# a_548_n1560# VDD VDD a_4254_n29# VDD VDD
+ a_548_n1560# a_4254_n29# a_548_n1560# VDD a_4254_n29# a_548_n1560# VDD a_4254_n29#
+ a_4254_n29# a_548_n1560# a_548_n1560# a_548_n1560# a_4254_n29# a_548_n1560# a_548_n1560#
+ a_548_n1560# VDD pmos_3p3_MV44E7
Xnmos_3p3_7NPLVN_0 OUT VSS VSS VSS VSS VSS a_4254_n29# VSS VSS a_4254_n29# OUT VSS
+ a_4254_n29# VSS VSS a_4254_n29# VSS a_4254_n29# VSS VSS VSS VSS VSS OUT VSS VSS
+ VSS OUT VSS VSS a_4254_n29# a_4254_n29# VSS a_4254_n29# VSS VSS VSS VSS a_4254_n29#
+ VSS VSS VSS OUT a_4254_n29# VSS OUT VSS a_4254_n29# VSS VSS VSS a_4254_n29# a_4254_n29#
+ VSS a_4254_n29# VSS OUT VSS nmos_3p3_7NPLVN
Xpmos_3p3_PPYSL5_0 a_548_n1560# IN IN VDD VDD VDD VDD IN a_548_n1560# IN pmos_3p3_PPYSL5
Xnmos_3p3_PLQLVN_0 VSS OUT a_4254_n29# a_4254_n29# OUT a_4254_n29# a_4254_n29# VSS
+ a_4254_n29# OUT a_4254_n29# a_4254_n29# OUT VSS VSS OUT OUT VSS a_4254_n29# VSS
+ a_4254_n29# a_4254_n29# VSS a_4254_n29# a_4254_n29# OUT VSS VSS a_4254_n29# OUT
+ a_4254_n29# a_4254_n29# VSS a_4254_n29# a_4254_n29# a_4254_n29# OUT VSS nmos_3p3_PLQLVN
Xnmos_3p3_8FEAMQ_0 IN IN a_548_n1560# VSS VSS VSS nmos_3p3_8FEAMQ
.ends

.subckt pmos_3p3_DVJ9E7 a_764_n60# a_n664_n60# a_664_n104# a_560_n60# a_n460_n60#
+ a_n764_n104# a_256_n104# a_n256_n60# a_356_n60# a_n356_n104# a_460_n104# a_n1376_n104#
+ a_1580_n60# a_n1480_n60# a_152_n60# a_n1668_n60# a_1276_n104# a_n560_n104# a_n1580_n104#
+ a_n52_n60# a_1376_n60# a_n1276_n60# a_1480_n104# a_52_n104# a_868_n104# a_n152_n104#
+ a_1172_n60# a_n1072_n60# a_n1172_n104# a_n968_n104# a_1072_n104# a_968_n60# a_n868_n60#
+ w_n1754_n190#
X0 a_n52_n60# a_n152_n104# a_n256_n60# w_n1754_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X1 a_1172_n60# a_1072_n104# a_968_n60# w_n1754_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X2 a_n256_n60# a_n356_n104# a_n460_n60# w_n1754_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X3 a_1376_n60# a_1276_n104# a_1172_n60# w_n1754_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X4 a_1580_n60# a_1480_n104# a_1376_n60# w_n1754_n190# pfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X5 a_n460_n60# a_n560_n104# a_n664_n60# w_n1754_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X6 a_n664_n60# a_n764_n104# a_n868_n60# w_n1754_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X7 a_n1072_n60# a_n1172_n104# a_n1276_n60# w_n1754_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X8 a_n868_n60# a_n968_n104# a_n1072_n60# w_n1754_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X9 a_n1276_n60# a_n1376_n104# a_n1480_n60# w_n1754_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X10 a_356_n60# a_256_n104# a_152_n60# w_n1754_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X11 a_560_n60# a_460_n104# a_356_n60# w_n1754_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X12 a_n1480_n60# a_n1580_n104# a_n1668_n60# w_n1754_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X13 a_764_n60# a_664_n104# a_560_n60# w_n1754_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X14 a_152_n60# a_52_n104# a_n52_n60# w_n1754_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X15 a_968_n60# a_868_n104# a_764_n60# w_n1754_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
.ends

.subckt pmos_3p3_ZBCND7 a_n1276_n100# a_1072_n144# a_1988_n100# a_n460_n100# a_1888_n144#
+ a_n1480_n100# a_764_n100# a_664_n144# a_n764_n144# a_n1784_n144# a_n52_n100# a_n1072_n100#
+ a_1784_n100# a_356_n100# a_n868_n100# a_n1888_n100# a_1684_n144# a_256_n144# a_n356_n144#
+ a_560_n100# a_n1376_n144# a_460_n144# a_1376_n100# a_n560_n144# a_1276_n144# a_n1580_n144#
+ a_1580_n100# a_152_n100# a_n664_n100# a_n1684_n100# a_n2076_n100# a_1480_n144# a_968_n100#
+ a_52_n144# a_868_n144# a_n152_n144# a_n1172_n144# w_n2162_n230# a_n968_n144# a_1172_n100#
+ a_n256_n100# a_n1988_n144#
X0 a_n460_n100# a_n560_n144# a_n664_n100# w_n2162_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_1784_n100# a_1684_n144# a_1580_n100# w_n2162_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X2 a_n664_n100# a_n764_n144# a_n868_n100# w_n2162_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X3 a_n1072_n100# a_n1172_n144# a_n1276_n100# w_n2162_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X4 a_n868_n100# a_n968_n144# a_n1072_n100# w_n2162_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X5 a_1988_n100# a_1888_n144# a_1784_n100# w_n2162_n230# pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X6 a_n1276_n100# a_n1376_n144# a_n1480_n100# w_n2162_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X7 a_356_n100# a_256_n144# a_152_n100# w_n2162_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X8 a_560_n100# a_460_n144# a_356_n100# w_n2162_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X9 a_n1480_n100# a_n1580_n144# a_n1684_n100# w_n2162_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X10 a_n1684_n100# a_n1784_n144# a_n1888_n100# w_n2162_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X11 a_764_n100# a_664_n144# a_560_n100# w_n2162_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X12 a_152_n100# a_52_n144# a_n52_n100# w_n2162_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X13 a_968_n100# a_868_n144# a_764_n100# w_n2162_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X14 a_n1888_n100# a_n1988_n144# a_n2076_n100# w_n2162_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X15 a_n52_n100# a_n152_n144# a_n256_n100# w_n2162_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X16 a_1172_n100# a_1072_n144# a_968_n100# w_n2162_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X17 a_1376_n100# a_1276_n144# a_1172_n100# w_n2162_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X18 a_n256_n100# a_n356_n144# a_n460_n100# w_n2162_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X19 a_1580_n100# a_1480_n144# a_1376_n100# w_n2162_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
.ends

.subckt pmos_3p3_5QR9E7 a_560_n40# a_n460_n40# a_n764_n84# a_1988_n40# a_n1888_n40#
+ a_1072_n84# a_n2076_n40# a_n560_n84# a_1784_n40# a_n1684_n40# a_n1988_n84# a_356_n40#
+ a_n256_n40# a_868_n84# a_1580_n40# a_n1480_n40# a_n356_n84# a_n1784_n84# a_152_n40#
+ a_664_n84# w_n2162_n170# a_n152_n84# a_n1580_n84# a_n52_n40# a_1376_n40# a_n1276_n40#
+ a_460_n84# a_1888_n84# a_n1376_n84# a_1172_n40# a_n1072_n40# a_1684_n84# a_256_n84#
+ a_n1172_n84# a_n868_n40# a_1480_n84# a_968_n40# a_n664_n40# a_52_n84# a_n968_n84#
+ a_764_n40# a_1276_n84#
X0 a_n1072_n40# a_n1172_n84# a_n1276_n40# w_n2162_n170# pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X1 a_n868_n40# a_n968_n84# a_n1072_n40# w_n2162_n170# pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X2 a_1988_n40# a_1888_n84# a_1784_n40# w_n2162_n170# pfet_03v3 ad=0.176p pd=1.68u as=0.104p ps=0.92u w=0.4u l=0.5u
X3 a_n1276_n40# a_n1376_n84# a_n1480_n40# w_n2162_n170# pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X4 a_356_n40# a_256_n84# a_152_n40# w_n2162_n170# pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X5 a_560_n40# a_460_n84# a_356_n40# w_n2162_n170# pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X6 a_n1480_n40# a_n1580_n84# a_n1684_n40# w_n2162_n170# pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X7 a_n1684_n40# a_n1784_n84# a_n1888_n40# w_n2162_n170# pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X8 a_764_n40# a_664_n84# a_560_n40# w_n2162_n170# pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X9 a_152_n40# a_52_n84# a_n52_n40# w_n2162_n170# pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X10 a_968_n40# a_868_n84# a_764_n40# w_n2162_n170# pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X11 a_n1888_n40# a_n1988_n84# a_n2076_n40# w_n2162_n170# pfet_03v3 ad=0.104p pd=0.92u as=0.176p ps=1.68u w=0.4u l=0.5u
X12 a_n52_n40# a_n152_n84# a_n256_n40# w_n2162_n170# pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X13 a_1172_n40# a_1072_n84# a_968_n40# w_n2162_n170# pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X14 a_n256_n40# a_n356_n84# a_n460_n40# w_n2162_n170# pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X15 a_1376_n40# a_1276_n84# a_1172_n40# w_n2162_n170# pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X16 a_1580_n40# a_1480_n84# a_1376_n40# w_n2162_n170# pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X17 a_n460_n40# a_n560_n84# a_n664_n40# w_n2162_n170# pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X18 a_1784_n40# a_1684_n84# a_1580_n40# w_n2162_n170# pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X19 a_n664_n40# a_n764_n84# a_n868_n40# w_n2162_n170# pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
.ends

.subckt nmos_3p3_Z2JHD6 a_n1276_n100# a_1072_n144# a_1988_n100# a_n460_n100# a_1888_n144#
+ a_n1480_n100# a_764_n100# a_664_n144# a_n764_n144# a_n1784_n144# a_n52_n100# a_n1072_n100#
+ a_1784_n100# a_356_n100# a_n868_n100# a_n1888_n100# a_1684_n144# a_256_n144# a_n356_n144#
+ a_560_n100# a_n1376_n144# a_460_n144# a_1376_n100# a_n560_n144# a_1276_n144# a_n1580_n144#
+ a_1580_n100# a_152_n100# a_n664_n100# a_n1684_n100# a_n2076_n100# a_1480_n144# a_968_n100#
+ a_52_n144# a_868_n144# a_n152_n144# a_n1172_n144# a_n968_n144# a_1172_n100# a_n256_n100#
+ a_n1988_n144# VSUBS
X0 a_n664_n100# a_n764_n144# a_n868_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_1784_n100# a_1684_n144# a_1580_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X2 a_n1072_n100# a_n1172_n144# a_n1276_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X3 a_n868_n100# a_n968_n144# a_n1072_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X4 a_1988_n100# a_1888_n144# a_1784_n100# VSUBS nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X5 a_n1276_n100# a_n1376_n144# a_n1480_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X6 a_356_n100# a_256_n144# a_152_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X7 a_560_n100# a_460_n144# a_356_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X8 a_n1480_n100# a_n1580_n144# a_n1684_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X9 a_n1684_n100# a_n1784_n144# a_n1888_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X10 a_764_n100# a_664_n144# a_560_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X11 a_152_n100# a_52_n144# a_n52_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X12 a_n1888_n100# a_n1988_n144# a_n2076_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X13 a_968_n100# a_868_n144# a_764_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X14 a_n52_n100# a_n152_n144# a_n256_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X15 a_1172_n100# a_1072_n144# a_968_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X16 a_1376_n100# a_1276_n144# a_1172_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X17 a_n256_n100# a_n356_n144# a_n460_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X18 a_1580_n100# a_1480_n144# a_1376_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X19 a_n460_n100# a_n560_n144# a_n664_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
.ends

.subckt pfet_03v3_TTE2U8 a_764_n60# a_n664_n60# a_n852_n60# a_664_n104# w_n938_n190#
+ a_560_n60# a_n460_n60# a_n764_n104# a_256_n104# a_n256_n60# a_356_n60# a_n356_n104#
+ a_460_n104# a_152_n60# a_n560_n104# a_n52_n60# a_52_n104# a_n152_n104#
X0 a_n52_n60# a_n152_n104# a_n256_n60# w_n938_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X1 a_n256_n60# a_n356_n104# a_n460_n60# w_n938_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X2 a_n460_n60# a_n560_n104# a_n664_n60# w_n938_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X3 a_n664_n60# a_n764_n104# a_n852_n60# w_n938_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X4 a_356_n60# a_256_n104# a_152_n60# w_n938_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X5 a_560_n60# a_460_n104# a_356_n60# w_n938_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X6 a_764_n60# a_664_n104# a_560_n60# w_n938_n190# pfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X7 a_152_n60# a_52_n104# a_n52_n60# w_n938_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
.ends

.subckt nmos_3p3_AJEA3B a_764_n60# a_n664_n60# a_n852_n60# a_664_n104# a_560_n60#
+ a_n460_n60# a_n764_n104# a_256_n104# a_n256_n60# a_356_n60# a_n356_n104# a_460_n104#
+ a_152_n60# a_n560_n104# a_n52_n60# a_52_n104# a_n152_n104# VSUBS
X0 a_n256_n60# a_n356_n104# a_n460_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X1 a_n460_n60# a_n560_n104# a_n664_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X2 a_n664_n60# a_n764_n104# a_n852_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X3 a_356_n60# a_256_n104# a_152_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X4 a_560_n60# a_460_n104# a_356_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X5 a_764_n60# a_664_n104# a_560_n60# VSUBS nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X6 a_152_n60# a_52_n104# a_n52_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X7 a_n52_n60# a_n152_n104# a_n256_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
.ends

.subckt Current_Mirror_Top VDD G_source_up G_source_dn VSS G_sink_up G_sink_dn SD0_1
+ G1_2 G1_1 SD1_1 G2_1 SD2_1 ITAIL ITAIL_SINK ITAIL_SRC A1 A2
Xpmos_3p3_DVJ9E7_0 VDD G_source_up G_source_up G_source_up G_source_dn G_source_up
+ G_source_dn G_source_up G_source_dn G_source_dn G_source_dn G_source_dn VDD G_source_up
+ G_source_up VDD G_source_dn G_source_dn G_source_up VDD G_source_up G_source_dn
+ G_source_up G_source_up G_source_up G_source_up G_source_dn G_source_up G_source_dn
+ G_source_up G_source_dn G_source_up VDD VDD pmos_3p3_DVJ9E7
Xpmos_3p3_ZBCND7_0 VDD G1_2 VDD VDD G1_2 G1_2 G1_1 G1_1 G1_1 G1_1 G1_1 G1_2 G1_2 VDD
+ G1_1 G1_2 G1_1 G1_2 G1_2 G1_2 G1_2 G1_2 G1_2 G1_2 G1_2 G1_1 G1_1 G1_2 G1_2 G1_1
+ VDD G1_1 G1_2 G1_1 G1_1 G1_1 G1_2 VDD G1_1 VDD G1_2 G1_2 pmos_3p3_ZBCND7
Xpmos_3p3_5QR9E7_0 SD1_1 VDD G1_1 VDD SD1_1 G1_2 VDD G1_2 SD1_1 G_sink_up G1_2 VDD
+ SD1_1 G1_1 G_sink_up SD1_1 G1_2 G1_1 SD1_1 G1_1 VDD G1_1 G1_1 G_sink_up SD1_1 VDD
+ G1_2 G1_2 G1_2 VDD SD1_1 G1_1 G1_2 G1_2 G_sink_up G1_1 SD1_1 SD1_1 G1_1 G1_1 G_sink_up
+ G1_2 pmos_3p3_5QR9E7
Xpmos_3p3_ZBCND7_1 G1_1 G1_1 G1_1 G1_1 G1_1 G1_2 VDD G1_2 G1_2 G1_2 VDD G1_2 G1_2
+ G1_1 VDD G1_2 G1_2 G1_1 G1_1 G1_2 G1_1 G1_1 G1_2 G1_1 G1_1 G1_2 VDD G1_2 G1_2 VDD
+ G1_1 G1_2 G1_2 G1_2 G1_2 G1_2 G1_1 VDD G1_2 G1_1 G1_2 G1_1 pmos_3p3_ZBCND7
Xnmos_3p3_Z2JHD6_0 G1_1 ITAIL G1_1 G1_1 ITAIL SD2_1 VSS G2_1 G2_1 G2_1 VSS SD2_1 SD2_1
+ G1_1 VSS SD2_1 G2_1 ITAIL ITAIL SD2_1 ITAIL ITAIL SD2_1 ITAIL ITAIL G2_1 VSS SD2_1
+ SD2_1 VSS G1_1 G2_1 SD2_1 G2_1 G2_1 G2_1 ITAIL G2_1 G1_1 SD2_1 ITAIL VSS nmos_3p3_Z2JHD6
Xnmos_3p3_Z2JHD6_1 VSS G2_1 VSS VSS G2_1 G2_1 ITAIL ITAIL ITAIL ITAIL ITAIL G2_1 G2_1
+ VSS ITAIL G2_1 ITAIL G2_1 G2_1 G2_1 G2_1 G2_1 G2_1 G2_1 G2_1 ITAIL ITAIL G2_1 G2_1
+ ITAIL VSS ITAIL G2_1 ITAIL ITAIL ITAIL G2_1 ITAIL VSS G2_1 G2_1 VSS nmos_3p3_Z2JHD6
Xnmos_3p3_Z2JHD6_2 ITAIL ITAIL ITAIL ITAIL ITAIL G2_1 VSS G2_1 G2_1 G2_1 VSS G2_1
+ G2_1 ITAIL VSS G2_1 G2_1 ITAIL ITAIL G2_1 ITAIL ITAIL G2_1 ITAIL ITAIL G2_1 VSS
+ G2_1 G2_1 VSS ITAIL G2_1 G2_1 G2_1 G2_1 G2_1 ITAIL G2_1 ITAIL G2_1 ITAIL VSS nmos_3p3_Z2JHD6
Xpfet_03v3_TTE2U8_0 ITAIL_SRC A1 ITAIL_SRC G_source_dn VDD A1 VDD G_source_dn G_source_up
+ A1 VDD G_source_up G_source_up A1 G_source_up ITAIL_SRC G_source_dn G_source_dn
+ pfet_03v3_TTE2U8
Xnmos_3p3_AJEA3B_0 G_sink_up G_sink_dn G_sink_up G_sink_up G_sink_dn VSS G_sink_up
+ G_sink_dn G_sink_dn VSS G_sink_dn G_sink_dn G_sink_dn G_sink_dn G_sink_up G_sink_up
+ G_sink_up VSS nmos_3p3_AJEA3B
Xnmos_3p3_Z2JHD6_3 VSS G2_1 VSS VSS G2_1 SD2_1 G1_1 ITAIL ITAIL ITAIL G1_1 SD2_1 SD2_1
+ VSS G1_1 SD2_1 ITAIL G2_1 G2_1 SD2_1 G2_1 G2_1 SD2_1 G2_1 G2_1 ITAIL G1_1 SD2_1
+ SD2_1 G1_1 VSS ITAIL SD2_1 ITAIL ITAIL ITAIL G2_1 ITAIL VSS SD2_1 G2_1 VSS nmos_3p3_Z2JHD6
Xpfet_03v3_TTE2U8_1 VDD A1 VDD G_source_up VDD A1 ITAIL_SRC G_source_up G_source_dn
+ A1 ITAIL_SRC G_source_dn G_source_dn A1 G_source_dn VDD G_source_up G_source_up
+ pfet_03v3_TTE2U8
Xnmos_3p3_AJEA3B_1 VSS SD0_1 VSS G_sink_dn SD0_1 G_source_dn G_sink_dn G_sink_up SD0_1
+ G_source_dn G_sink_up G_sink_up SD0_1 G_sink_up VSS G_sink_dn G_sink_dn VSS nmos_3p3_AJEA3B
Xnmos_3p3_AJEA3B_2 ITAIL_SINK A2 ITAIL_SINK G_sink_up A2 VSS G_sink_up G_sink_dn A2
+ VSS G_sink_dn G_sink_dn A2 G_sink_dn ITAIL_SINK G_sink_up G_sink_up VSS nmos_3p3_AJEA3B
Xnmos_3p3_AJEA3B_4 VSS G_sink_dn VSS G_sink_dn G_sink_dn G_sink_up G_sink_dn G_sink_up
+ G_sink_dn G_sink_up G_sink_up G_sink_up G_sink_dn G_sink_up VSS G_sink_dn G_sink_dn
+ VSS nmos_3p3_AJEA3B
Xnmos_3p3_AJEA3B_3 G_source_dn SD0_1 G_source_dn G_sink_up SD0_1 VSS G_sink_up G_sink_dn
+ SD0_1 VSS G_sink_dn G_sink_dn SD0_1 G_sink_dn G_source_dn G_sink_up G_sink_up VSS
+ nmos_3p3_AJEA3B
Xnmos_3p3_AJEA3B_5 VSS A2 VSS G_sink_dn A2 ITAIL_SINK G_sink_dn G_sink_up A2 ITAIL_SINK
+ G_sink_up G_sink_up A2 G_sink_up VSS G_sink_dn G_sink_dn VSS nmos_3p3_AJEA3B
.ends

.subckt pmos_3p3_M8SWPS a_n28_n124# a_n116_n80# a_28_n80# w_n202_n210#
X0 a_28_n80# a_n28_n124# a_n116_n80# w_n202_n210# pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
.ends

.subckt nmos_3p3_5QNVWA a_n116_n44# a_28_n44# a_n28_n88# VSUBS
X0 a_28_n44# a_n28_n88# a_n116_n44# VSUBS nfet_03v3 ad=0.1936p pd=1.76u as=0.1936p ps=1.76u w=0.44u l=0.28u
.ends

.subckt nand2_ibr VDD IN2 IN1 OUT VSS
Xpmos_3p3_M8SWPS_0 IN1 OUT VDD VDD pmos_3p3_M8SWPS
Xpmos_3p3_M8SWPS_1 IN2 VDD OUT VDD pmos_3p3_M8SWPS
Xnmos_3p3_5QNVWA_0 VSS m1_186_70# IN2 VSS nmos_3p3_5QNVWA
Xnmos_3p3_5QNVWA_1 m1_186_70# OUT IN1 VSS nmos_3p3_5QNVWA
.ends

.subckt pmos_3p3_MQGBLR a_n28_n124# a_n116_n80# a_28_n80# w_n202_n210#
X0 a_28_n80# a_n28_n124# a_n116_n80# w_n202_n210# pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
.ends

.subckt nmos_3p3_DDNVWA a_n120_n36# a_28_n22# a_n28_n66# VSUBS
X0 a_28_n22# a_n28_n66# a_n120_n36# VSUBS nfet_03v3 ad=0.1516p pd=1.64u as=0.1516p ps=1.64u w=0.22u l=0.28u
.ends

.subckt nverterlayout_ibr VDD VSS OUT IN
Xpmos_3p3_MQGBLR_0 IN VDD OUT VDD pmos_3p3_MQGBLR
Xnmos_3p3_DDNVWA_0 VSS OUT IN VSS nmos_3p3_DDNVWA
.ends

.subckt mux_2x1_ibr Sel I1 OUT I0 VDD VSS
Xnand2_ibr_0 VDD I1 Sel nand2_ibr_1/IN2 VSS nand2_ibr
Xnand2_ibr_1 VDD nand2_ibr_1/IN2 nand2_ibr_2/OUT OUT VSS nand2_ibr
Xnand2_ibr_2 VDD nand2_ibr_2/IN2 I0 nand2_ibr_2/OUT VSS nand2_ibr
Xnverterlayout_ibr_0 VDD VSS nand2_ibr_2/IN2 Sel nverterlayout_ibr
.ends

.subckt mux_4x1_ibr I0 I1 I2 I3 S1 S0 OUT VSS VDD
Xmux_2x1_ibr_0 S0 I1 mux_2x1_ibr_2/I0 I0 VDD VSS mux_2x1_ibr
Xmux_2x1_ibr_1 S0 I3 mux_2x1_ibr_2/I1 I2 VDD VSS mux_2x1_ibr
Xmux_2x1_ibr_2 S1 mux_2x1_ibr_2/I1 OUT mux_2x1_ibr_2/I0 VDD VSS mux_2x1_ibr
.ends

.subckt nand2 IN2 IN1 OUT VSS VDD
Xpmos_3p3_M8SWPS_0 IN1 OUT VDD VDD pmos_3p3_M8SWPS
Xpmos_3p3_M8SWPS_1 IN2 VDD OUT VDD pmos_3p3_M8SWPS
Xnmos_3p3_5QNVWA_0 VSS m1_186_70# IN2 VSS nmos_3p3_5QNVWA
Xnmos_3p3_5QNVWA_1 m1_186_70# OUT IN1 VSS nmos_3p3_5QNVWA
.ends

.subckt nverterlayout VDD VSS OUT IN
Xpmos_3p3_MQGBLR_0 IN VDD OUT VDD pmos_3p3_MQGBLR
Xnmos_3p3_DDNVWA_0 VSS OUT IN VSS nmos_3p3_DDNVWA
.ends

.subckt mux_2x1 Sel I0 I1 VDD OUT VSS
Xnand2_0 I1 Sel nand2_1/IN2 VSS VDD nand2
Xnand2_1 nand2_1/IN2 nand2_2/OUT OUT VSS VDD nand2
Xnand2_2 nand2_2/IN2 I0 nand2_2/OUT VSS VDD nand2
Xnverterlayout_0 VDD VSS nand2_2/IN2 Sel nverterlayout
.ends

.subckt mux_4x1 I0 I1 I2 I3 S1 S0 OUT VSS mux_2x1_1/I0 VDD
Xmux_2x1_0 S0 I2 I3 VDD mux_2x1_1/I1 VSS mux_2x1
Xmux_2x1_1 S1 mux_2x1_1/I0 mux_2x1_1/I1 VDD OUT VSS mux_2x1
Xmux_2x1_2 S0 I0 I1 VDD mux_2x1_1/I0 VSS mux_2x1
.ends

.subckt and_2_ibr VDD IN2 OUT IN1 nand2_ibr_0/OUT VSS
Xnand2_ibr_0 VDD IN2 IN1 nand2_ibr_0/OUT VSS nand2_ibr
Xnverterlayout_ibr_0 VDD VSS OUT nand2_ibr_0/OUT nverterlayout_ibr
.ends

.subckt dec_2x4_ibr_mag IN1 IN2 D0 D1 D2 D3 VSS VDD
Xand_2_ibr_0 VDD and_2_ibr_2/IN2 D0 and_2_ibr_1/IN1 and_2_ibr_0/nand2_ibr_0/OUT VSS
+ and_2_ibr
Xand_2_ibr_1 VDD IN1 D1 and_2_ibr_1/IN1 and_2_ibr_1/nand2_ibr_0/OUT VSS and_2_ibr
Xand_2_ibr_2 VDD and_2_ibr_2/IN2 D2 IN2 and_2_ibr_2/nand2_ibr_0/OUT VSS and_2_ibr
Xand_2_ibr_3 VDD IN1 D3 IN2 and_2_ibr_3/nand2_ibr_0/OUT VSS and_2_ibr
Xnverterlayout_ibr_0 VDD VSS and_2_ibr_2/IN2 IN1 nverterlayout_ibr
Xnverterlayout_ibr_1 VDD VSS and_2_ibr_1/IN1 IN2 nverterlayout_ibr
.ends

.subckt nand2_mag IN2 IN1 VSS OUT m1_186_70# VDD
Xpmos_3p3_M8SWPS_0 IN1 OUT VDD VDD pmos_3p3_M8SWPS
Xpmos_3p3_M8SWPS_1 IN2 VDD OUT VDD pmos_3p3_M8SWPS
Xnmos_3p3_5QNVWA_0 VSS m1_186_70# IN2 VSS nmos_3p3_5QNVWA
Xnmos_3p3_5QNVWA_1 m1_186_70# OUT IN1 VSS nmos_3p3_5QNVWA
.ends

.subckt nmos_3p3_VGTVWA a_n116_n66# a_28_n66# a_n28_n110# VSUBS
X0 a_28_n66# a_n28_n110# a_n116_n66# VSUBS nfet_03v3 ad=0.2904p pd=2.2u as=0.2904p ps=2.2u w=0.66u l=0.28u
.ends

.subckt nand3_mag IN3 IN2 IN1 nmos_3p3_VGTVWA_1/a_28_n66# VSS nmos_3p3_VGTVWA_0/a_28_n66#
+ OUT VDD
Xnmos_3p3_VGTVWA_0 nmos_3p3_VGTVWA_1/a_28_n66# nmos_3p3_VGTVWA_0/a_28_n66# IN2 VSS
+ nmos_3p3_VGTVWA
Xnmos_3p3_VGTVWA_1 VSS nmos_3p3_VGTVWA_1/a_28_n66# IN3 VSS nmos_3p3_VGTVWA
Xnmos_3p3_VGTVWA_2 nmos_3p3_VGTVWA_0/a_28_n66# OUT IN1 VSS nmos_3p3_VGTVWA
Xpmos_3p3_M8SWPS_0 IN1 VDD OUT VDD pmos_3p3_M8SWPS
Xpmos_3p3_M8SWPS_1 IN3 VDD OUT VDD pmos_3p3_M8SWPS
Xpmos_3p3_M8SWPS_2 IN2 OUT VDD VDD pmos_3p3_M8SWPS
.ends

.subckt GF_INV_MAG IN OUT VSS w_n118_526#
Xpmos_3p3_MQGBLR_0 IN w_n118_526# OUT w_n118_526# pmos_3p3_MQGBLR
Xnmos_3p3_DDNVWA_0 VSS OUT IN VSS nmos_3p3_DDNVWA
.ends

.subckt JK_FF_mag RST J K nand2_mag_1/m1_186_70# nand3_mag_2/nmos_3p3_VGTVWA_1/a_28_n66#
+ nand2_mag_3/m1_186_70# nand3_mag_0/nmos_3p3_VGTVWA_0/a_28_n66# nand2_mag_2/m1_186_70#
+ nand2_mag_4/m1_186_70# nand3_mag_1/nmos_3p3_VGTVWA_0/a_28_n66# nand2_mag_4/IN2 nand3_mag_0/nmos_3p3_VGTVWA_1/a_28_n66#
+ nand3_mag_2/nmos_3p3_VGTVWA_0/a_28_n66# nand2_mag_1/IN2 nand3_mag_2/OUT nand3_mag_0/OUT
+ CLK QB nand3_mag_1/IN1 nand2_mag_3/IN1 nand3_mag_1/nmos_3p3_VGTVWA_1/a_28_n66# nand2_mag_0/m1_186_70#
+ Q nand3_mag_1/OUT VSS VDD
Xnand2_mag_1 nand2_mag_1/IN2 QB VSS Q nand2_mag_1/m1_186_70# VDD nand2_mag
Xnand3_mag_2 J CLK Q nand3_mag_2/nmos_3p3_VGTVWA_1/a_28_n66# VSS nand3_mag_2/nmos_3p3_VGTVWA_0/a_28_n66#
+ nand3_mag_2/OUT VDD nand3_mag
Xnand2_mag_2 nand3_mag_0/OUT nand3_mag_1/OUT VSS nand3_mag_1/IN1 nand2_mag_2/m1_186_70#
+ VDD nand2_mag
Xnand2_mag_3 nand3_mag_1/OUT nand2_mag_3/IN1 VSS nand2_mag_4/IN2 nand2_mag_3/m1_186_70#
+ VDD nand2_mag
Xnand2_mag_4 nand2_mag_4/IN2 Q VSS QB nand2_mag_4/m1_186_70# VDD nand2_mag
XGF_INV_MAG_0 CLK nand2_mag_3/IN1 VSS VDD GF_INV_MAG
Xnand3_mag_0 K CLK QB nand3_mag_0/nmos_3p3_VGTVWA_1/a_28_n66# VSS nand3_mag_0/nmos_3p3_VGTVWA_0/a_28_n66#
+ nand3_mag_0/OUT VDD nand3_mag
Xnand2_mag_0 nand3_mag_1/IN1 nand2_mag_3/IN1 VSS nand2_mag_1/IN2 nand2_mag_0/m1_186_70#
+ VDD nand2_mag
Xnand3_mag_1 nand3_mag_2/OUT RST nand3_mag_1/IN1 nand3_mag_1/nmos_3p3_VGTVWA_1/a_28_n66#
+ VSS nand3_mag_1/nmos_3p3_VGTVWA_0/a_28_n66# nand3_mag_1/OUT VDD nand3_mag
.ends

.subckt CLK_div_2_mag Vdiv2 CLK JK_FF_mag_0/nand3_mag_0/OUT JK_FF_mag_0/nand3_mag_1/OUT
+ VSS RST JK_FF_mag_0/nand3_mag_2/OUT VDD
XJK_FF_mag_0 RST VDD VDD JK_FF_mag_0/nand2_mag_1/m1_186_70# JK_FF_mag_0/nand3_mag_2/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_0/nand2_mag_3/m1_186_70# JK_FF_mag_0/nand3_mag_0/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_0/nand2_mag_2/m1_186_70# JK_FF_mag_0/nand2_mag_4/m1_186_70# JK_FF_mag_0/nand3_mag_1/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_0/nand2_mag_4/IN2 JK_FF_mag_0/nand3_mag_0/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_0/nand3_mag_2/nmos_3p3_VGTVWA_0/a_28_n66# JK_FF_mag_0/nand2_mag_1/IN2
+ JK_FF_mag_0/nand3_mag_2/OUT JK_FF_mag_0/nand3_mag_0/OUT CLK JK_FF_mag_0/QB JK_FF_mag_0/nand3_mag_1/IN1
+ JK_FF_mag_0/nand2_mag_3/IN1 JK_FF_mag_0/nand3_mag_1/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_0/nand2_mag_0/m1_186_70# Vdiv2 JK_FF_mag_0/nand3_mag_1/OUT VSS VDD JK_FF_mag
.ends

.subckt CLK_div_4_mag Vdiv4 VSS RST CLK CLK_div_2_mag_0/JK_FF_mag_0/nand3_mag_2/OUT
+ CLK_div_2_mag_1/JK_FF_mag_0/nand3_mag_1/OUT CLK_div_2_mag_1/JK_FF_mag_0/nand3_mag_2/OUT
+ CLK_div_2_mag_0/JK_FF_mag_0/nand3_mag_0/OUT VDD CLK_div_2_mag_0/JK_FF_mag_0/nand3_mag_1/OUT
+ CLK_div_2_mag_1/JK_FF_mag_0/nand3_mag_0/OUT
XCLK_div_2_mag_0 CLK_div_2_mag_1/CLK CLK CLK_div_2_mag_0/JK_FF_mag_0/nand3_mag_0/OUT
+ CLK_div_2_mag_0/JK_FF_mag_0/nand3_mag_1/OUT VSS RST CLK_div_2_mag_0/JK_FF_mag_0/nand3_mag_2/OUT
+ VDD CLK_div_2_mag
XCLK_div_2_mag_1 Vdiv4 CLK_div_2_mag_1/CLK CLK_div_2_mag_1/JK_FF_mag_0/nand3_mag_0/OUT
+ CLK_div_2_mag_1/JK_FF_mag_0/nand3_mag_1/OUT VSS RST CLK_div_2_mag_1/JK_FF_mag_0/nand3_mag_2/OUT
+ VDD CLK_div_2_mag
.ends

.subckt pmos_3p3_M8QNDR w_n202_n290# a_28_n160# a_n116_n160# a_n28_n204#
X0 a_28_n160# a_n28_n204# a_n116_n160# w_n202_n290# pfet_03v3 ad=0.704p pd=4.08u as=0.704p ps=4.08u w=1.6u l=0.28u
.ends

.subckt pmos_3p3_M4YALR w_n202_n290# a_28_n160# a_n116_n160# a_n28_n204#
X0 a_28_n160# a_n28_n204# a_n116_n160# w_n202_n290# pfet_03v3 ad=0.704p pd=4.08u as=0.704p ps=4.08u w=1.6u l=0.28u
.ends

.subckt or_2_mag VSS IN2 IN1 OUT w_721_942#
Xpmos_3p3_M8QNDR_0 w_721_942# pmos_3p3_M8QNDR_0/a_28_n160# w_721_942# IN2 pmos_3p3_M8QNDR
XGF_INV_MAG_1 GF_INV_MAG_1/IN OUT VSS w_721_942# GF_INV_MAG
Xpmos_3p3_M4YALR_0 w_721_942# GF_INV_MAG_1/IN pmos_3p3_M8QNDR_0/a_28_n160# IN1 pmos_3p3_M4YALR
Xnmos_3p3_DDNVWA_0 GF_INV_MAG_1/IN VSS IN1 VSS nmos_3p3_DDNVWA
Xnmos_3p3_DDNVWA_1 VSS GF_INV_MAG_1/IN IN2 VSS nmos_3p3_DDNVWA
.ends

.subckt and2_mag IN2 IN1 OUT VDD VSS
Xpmos_3p3_M8SWPS_0 IN1 GF_INV_MAG_0/IN VDD VDD pmos_3p3_M8SWPS
Xpmos_3p3_M8SWPS_1 IN2 VDD GF_INV_MAG_0/IN VDD pmos_3p3_M8SWPS
XGF_INV_MAG_0 GF_INV_MAG_0/IN OUT VSS VDD GF_INV_MAG
Xnmos_3p3_5QNVWA_0 VSS m1_186_70# IN2 VSS nmos_3p3_5QNVWA
Xnmos_3p3_5QNVWA_1 m1_186_70# GF_INV_MAG_0/IN IN1 VSS nmos_3p3_5QNVWA
.ends

.subckt CLK_div_3_mag Q1 Q0 Vdiv3 JK_FF_mag_1/nand3_mag_0/OUT JK_FF_mag_0/nand3_mag_0/OUT
+ JK_FF_mag_1/nand3_mag_1/OUT JK_FF_mag_0/nand3_mag_1/OUT JK_FF_mag_1/nand3_mag_2/OUT
+ VSS CLK RST JK_FF_mag_0/nand3_mag_2/OUT VDD
XJK_FF_mag_1 RST VDD JK_FF_mag_1/K JK_FF_mag_1/nand2_mag_1/m1_186_70# JK_FF_mag_1/nand3_mag_2/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_1/nand2_mag_3/m1_186_70# JK_FF_mag_1/nand3_mag_0/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_1/nand2_mag_2/m1_186_70# JK_FF_mag_1/nand2_mag_4/m1_186_70# JK_FF_mag_1/nand3_mag_1/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_1/nand2_mag_4/IN2 JK_FF_mag_1/nand3_mag_0/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_1/nand3_mag_2/nmos_3p3_VGTVWA_0/a_28_n66# JK_FF_mag_1/nand2_mag_1/IN2
+ JK_FF_mag_1/nand3_mag_2/OUT JK_FF_mag_1/nand3_mag_0/OUT CLK JK_FF_mag_1/QB JK_FF_mag_1/nand3_mag_1/IN1
+ JK_FF_mag_1/nand2_mag_3/IN1 JK_FF_mag_1/nand3_mag_1/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_1/nand2_mag_0/m1_186_70# Q1 JK_FF_mag_1/nand3_mag_1/OUT VSS VDD JK_FF_mag
XJK_FF_mag_0 RST VDD Q1 JK_FF_mag_0/nand2_mag_1/m1_186_70# JK_FF_mag_0/nand3_mag_2/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_0/nand2_mag_3/m1_186_70# JK_FF_mag_0/nand3_mag_0/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_0/nand2_mag_2/m1_186_70# JK_FF_mag_0/nand2_mag_4/m1_186_70# JK_FF_mag_0/nand3_mag_1/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_0/nand2_mag_4/IN2 JK_FF_mag_0/nand3_mag_0/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_0/nand3_mag_2/nmos_3p3_VGTVWA_0/a_28_n66# JK_FF_mag_0/nand2_mag_1/IN2
+ JK_FF_mag_0/nand3_mag_2/OUT JK_FF_mag_0/nand3_mag_0/OUT CLK JK_FF_mag_1/K JK_FF_mag_0/nand3_mag_1/IN1
+ JK_FF_mag_0/nand2_mag_3/IN1 JK_FF_mag_0/nand3_mag_1/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_0/nand2_mag_0/m1_186_70# Q0 JK_FF_mag_0/nand3_mag_1/OUT VSS VDD JK_FF_mag
Xor_2_mag_0 VSS or_2_mag_0/IN2 Q0 Vdiv3 VDD or_2_mag
Xand2_mag_0 CLK Q1 or_2_mag_0/IN2 VDD VSS and2_mag
.ends

.subckt pmos_3p3_MW53B7 a_n188_n80# a_n100_n124# a_100_n80# w_n274_n210#
X0 a_100_n80# a_n100_n124# a_n188_n80# w_n274_n210# pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
.ends

.subckt nmos_3p3_MGBSF7 a_100_n22# a_n100_n66# a_n192_n36# VSUBS
X0 a_100_n22# a_n100_n66# a_n192_n36# VSUBS nfet_03v3 ad=0.1516p pd=1.64u as=0.1516p ps=1.64u w=0.22u l=1u
.ends

.subckt Inverter_delayed_mag VSS IN OUT VDD
Xpmos_3p3_MW53B7_0 VDD IN OUT VDD pmos_3p3_MW53B7
Xnmos_3p3_MGBSF7_0 OUT IN VSS VSS nmos_3p3_MGBSF7
.ends

.subckt Buffer_delayed_mag IN OUT VDD VSS
Xpmos_3p3_MW53B7_0 VDD IN Inverter_delayed_mag_0/IN VDD pmos_3p3_MW53B7
XInverter_delayed_mag_0 VSS Inverter_delayed_mag_0/IN OUT VDD Inverter_delayed_mag
Xnmos_3p3_MGBSF7_0 Inverter_delayed_mag_0/IN IN VSS VSS nmos_3p3_MGBSF7
.ends

.subckt Output_Div_Mag OPA0 OPA1 Vdiv VDD RST CLK VSS
Xmux_4x1_0 mux_4x1_0/I0 mux_4x1_0/I1 mux_4x1_0/I2 mux_4x1_0/I3 OPA1 OPA0 Vdiv VSS
+ mux_4x1_0/mux_2x1_1/I0 VDD mux_4x1
Xdec_2x4_ibr_mag_0 OPA0 OPA1 dec_2x4_ibr_mag_0/D0 CLK_div_2_mag_0/VDD CLK_div_3_mag_0/VDD
+ CLK_div_4_mag_0/VDD VSS VDD dec_2x4_ibr_mag
XCLK_div_4_mag_0 mux_4x1_0/I3 VSS RST CLK CLK_div_4_mag_0/CLK_div_2_mag_0/JK_FF_mag_0/nand3_mag_2/OUT
+ CLK_div_4_mag_0/CLK_div_2_mag_1/JK_FF_mag_0/nand3_mag_1/OUT CLK_div_4_mag_0/CLK_div_2_mag_1/JK_FF_mag_0/nand3_mag_2/OUT
+ CLK_div_4_mag_0/CLK_div_2_mag_0/JK_FF_mag_0/nand3_mag_0/OUT CLK_div_4_mag_0/VDD
+ CLK_div_4_mag_0/CLK_div_2_mag_0/JK_FF_mag_0/nand3_mag_1/OUT CLK_div_4_mag_0/CLK_div_2_mag_1/JK_FF_mag_0/nand3_mag_0/OUT
+ CLK_div_4_mag
XCLK_div_3_mag_0 CLK_div_3_mag_0/Q1 CLK_div_3_mag_0/Q0 mux_4x1_0/I2 CLK_div_3_mag_0/JK_FF_mag_1/nand3_mag_0/OUT
+ CLK_div_3_mag_0/JK_FF_mag_0/nand3_mag_0/OUT CLK_div_3_mag_0/JK_FF_mag_1/nand3_mag_1/OUT
+ CLK_div_3_mag_0/JK_FF_mag_0/nand3_mag_1/OUT CLK_div_3_mag_0/JK_FF_mag_1/nand3_mag_2/OUT
+ VSS CLK RST CLK_div_3_mag_0/JK_FF_mag_0/nand3_mag_2/OUT CLK_div_3_mag_0/VDD CLK_div_3_mag
XCLK_div_2_mag_0 mux_4x1_0/I1 CLK CLK_div_2_mag_0/JK_FF_mag_0/nand3_mag_0/OUT CLK_div_2_mag_0/JK_FF_mag_0/nand3_mag_1/OUT
+ VSS RST CLK_div_2_mag_0/JK_FF_mag_0/nand3_mag_2/OUT CLK_div_2_mag_0/VDD CLK_div_2_mag
XBuffer_delayed_mag_0 CLK mux_4x1_0/I0 dec_2x4_ibr_mag_0/D0 VSS Buffer_delayed_mag
.ends

.subckt pmos_3p3_MYFUKR a_28_n240# a_n28_n284# a_n116_n240# w_n202_n370#
X0 a_28_n240# a_n28_n284# a_n116_n240# w_n202_n370# pfet_03v3 ad=1.056p pd=5.68u as=1.056p ps=5.68u w=2.4u l=0.28u
.ends

.subckt nor_3_mag IN3 IN2 IN1 OUT VSS w_801_880#
Xnmos_3p3_DDNVWA_2 OUT VSS IN2 VSS nmos_3p3_DDNVWA
Xpmos_3p3_MYFUKR_0 OUT IN1 pmos_3p3_MYFUKR_2/a_28_n240# w_801_880# pmos_3p3_MYFUKR
Xpmos_3p3_MYFUKR_1 pmos_3p3_MYFUKR_1/a_28_n240# IN3 w_801_880# w_801_880# pmos_3p3_MYFUKR
Xpmos_3p3_MYFUKR_2 pmos_3p3_MYFUKR_2/a_28_n240# IN2 pmos_3p3_MYFUKR_1/a_28_n240# w_801_880#
+ pmos_3p3_MYFUKR
Xnmos_3p3_DDNVWA_0 VSS OUT IN1 VSS nmos_3p3_DDNVWA
Xnmos_3p3_DDNVWA_1 VSS OUT IN3 VSS nmos_3p3_DDNVWA
.ends

.subckt CLK_DIV_11_mag_new CLK Vdiv11 Q3 Q2 Q1 Q0 VDD RST VSS
XJK_FF_mag_1 RST JK_FF_mag_1/K JK_FF_mag_1/K m1_7762_3820# m1_5915_5036# m1_7352_4917#
+ m1_6081_3939# m1_6634_3820# m1_7916_4917# m1_6799_5036# JK_FF_mag_1/nand2_mag_4/IN2
+ m1_5921_3939# m1_6075_5036# JK_FF_mag_1/nand2_mag_1/IN2 JK_FF_mag_1/nand3_mag_2/OUT
+ JK_FF_mag_1/nand3_mag_0/OUT CLK JK_FF_mag_1/QB JK_FF_mag_1/nand3_mag_1/IN1 JK_FF_mag_1/nand2_mag_3/IN1
+ m1_6639_5036# m1_7198_3820# Q2 JK_FF_mag_1/nand3_mag_1/OUT VSS VDD JK_FF_mag
XJK_FF_mag_0 RST JK_FF_mag_0/K JK_FF_mag_0/K m1_4627_3818# m1_2780_5034# m1_4217_4915#
+ m1_2946_3937# m1_3499_3818# m1_4781_4915# m1_3664_5034# JK_FF_mag_0/nand2_mag_4/IN2
+ m1_2786_3937# m1_2940_5034# JK_FF_mag_0/nand2_mag_1/IN2 JK_FF_mag_0/nand3_mag_2/OUT
+ JK_FF_mag_0/nand3_mag_0/OUT CLK or_2_mag_3/IN2 JK_FF_mag_0/nand3_mag_1/IN1 JK_FF_mag_0/nand2_mag_3/IN1
+ m1_3504_5034# m1_4063_3818# Q3 JK_FF_mag_0/nand3_mag_1/OUT VSS VDD JK_FF_mag
XJK_FF_mag_2 RST JK_FF_mag_2/K JK_FF_mag_2/K m1_10876_3818# m1_9029_5034# m1_10466_4915#
+ m1_9195_3937# m1_9748_3818# m1_11030_4915# m1_9913_5034# JK_FF_mag_2/nand2_mag_4/IN2
+ m1_9035_3937# m1_9189_5034# JK_FF_mag_2/nand2_mag_1/IN2 JK_FF_mag_2/nand3_mag_2/OUT
+ JK_FF_mag_2/nand3_mag_0/OUT CLK or_2_mag_3/IN1 JK_FF_mag_2/nand3_mag_1/IN1 JK_FF_mag_2/nand2_mag_3/IN1
+ m1_9753_5034# m1_10312_3818# Q1 JK_FF_mag_2/nand3_mag_1/OUT VSS VDD JK_FF_mag
XJK_FF_mag_3 RST JK_FF_mag_3/K JK_FF_mag_3/K m1_14035_3822# m1_12188_5038# m1_13625_4919#
+ m1_12354_3941# m1_12907_3822# m1_14189_4919# m1_13072_5038# JK_FF_mag_3/nand2_mag_4/IN2
+ m1_12194_3941# m1_12348_5038# JK_FF_mag_3/nand2_mag_1/IN2 JK_FF_mag_3/nand3_mag_2/OUT
+ JK_FF_mag_3/nand3_mag_0/OUT CLK JK_FF_mag_3/QB JK_FF_mag_3/nand3_mag_1/IN1 JK_FF_mag_3/nand2_mag_3/IN1
+ m1_12912_5038# m1_13471_3822# Q0 JK_FF_mag_3/nand3_mag_1/OUT VSS VDD JK_FF_mag
XGF_INV_MAG_0 nand3_mag_0/OUT or_2_mag_0/IN2 VSS VDD GF_INV_MAG
XGF_INV_MAG_1 nand3_mag_1/OUT GF_INV_MAG_1/OUT VSS VDD GF_INV_MAG
XGF_INV_MAG_2 nor_3_mag_0/OUT Vdiv11 VSS VDD GF_INV_MAG
Xor_2_mag_0 VSS or_2_mag_0/IN2 or_2_mag_0/IN1 JK_FF_mag_0/K VDD or_2_mag
Xor_2_mag_1 VSS Q0 or_2_mag_1/IN1 JK_FF_mag_2/K VDD or_2_mag
Xor_2_mag_3 VSS or_2_mag_3/IN2 or_2_mag_3/IN1 JK_FF_mag_3/K VDD or_2_mag
Xand2_mag_0 Q1 Q3 or_2_mag_0/IN1 VDD VSS and2_mag
Xand2_mag_1 Q0 Q1 JK_FF_mag_1/K VDD VSS and2_mag
Xand2_mag_2 Q1 Q3 or_2_mag_1/IN1 VDD VSS and2_mag
Xand2_mag_3 Q1 and2_mag_3/IN1 and2_mag_3/OUT VDD VSS and2_mag
XBuffer_delayed_mag_1 GF_INV_MAG_1/OUT nor_3_mag_0/IN3 VDD VSS Buffer_delayed_mag
XBuffer_delayed_mag_0 Q2 and2_mag_3/IN1 VDD VSS Buffer_delayed_mag
Xnor_3_mag_0 nor_3_mag_0/IN3 and2_mag_3/OUT Q3 nor_3_mag_0/OUT VSS VDD nor_3_mag
Xnand3_mag_0 Q1 Q0 Q2 nand3_mag_0/nmos_3p3_VGTVWA_1/a_28_n66# VSS nand3_mag_0/nmos_3p3_VGTVWA_0/a_28_n66#
+ nand3_mag_0/OUT VDD nand3_mag
Xnand3_mag_1 and2_mag_3/IN1 Q0 CLK nand3_mag_1/nmos_3p3_VGTVWA_1/a_28_n66# VSS nand3_mag_1/nmos_3p3_VGTVWA_0/a_28_n66#
+ nand3_mag_1/OUT VDD nand3_mag
.ends

.subckt CLK_div_99_mag VDD CLK Vdiv99 RST VSS
XCLK_DIV_11_mag_new_0 CLK_div_3_mag_0/Vdiv3 Vdiv99 CLK_DIV_11_mag_new_0/Q3 CLK_DIV_11_mag_new_0/Q2
+ CLK_DIV_11_mag_new_0/Q1 CLK_DIV_11_mag_new_0/Q0 VDD RST VSS CLK_DIV_11_mag_new
XCLK_div_3_mag_1 CLK_div_3_mag_1/Q1 CLK_div_3_mag_1/Q0 CLK_div_3_mag_0/CLK CLK_div_3_mag_1/JK_FF_mag_1/nand3_mag_0/OUT
+ CLK_div_3_mag_1/JK_FF_mag_0/nand3_mag_0/OUT CLK_div_3_mag_1/JK_FF_mag_1/nand3_mag_1/OUT
+ CLK_div_3_mag_1/JK_FF_mag_0/nand3_mag_1/OUT CLK_div_3_mag_1/JK_FF_mag_1/nand3_mag_2/OUT
+ VSS CLK RST CLK_div_3_mag_1/JK_FF_mag_0/nand3_mag_2/OUT VDD CLK_div_3_mag
XCLK_div_3_mag_0 CLK_div_3_mag_0/Q1 CLK_div_3_mag_0/Q0 CLK_div_3_mag_0/Vdiv3 CLK_div_3_mag_0/JK_FF_mag_1/nand3_mag_0/OUT
+ CLK_div_3_mag_0/JK_FF_mag_0/nand3_mag_0/OUT CLK_div_3_mag_0/JK_FF_mag_1/nand3_mag_1/OUT
+ CLK_div_3_mag_0/JK_FF_mag_0/nand3_mag_1/OUT CLK_div_3_mag_0/JK_FF_mag_1/nand3_mag_2/OUT
+ VSS CLK_div_3_mag_0/CLK RST CLK_div_3_mag_0/JK_FF_mag_0/nand3_mag_2/OUT VDD CLK_div_3_mag
.ends

.subckt mux_8x1_ibr I0 I1 I2 I3 I5 I6 I7 OUT S0 S1 S2 I4 VSS VDD
Xmux_4x1_ibr_0 I4 I5 I6 I7 S1 S0 mux_2x1_ibr_0/I1 VSS VDD mux_4x1_ibr
Xmux_4x1_ibr_1 I0 I1 I2 I3 S1 S0 mux_2x1_ibr_0/I0 VSS VDD mux_4x1_ibr
Xmux_2x1_ibr_0 S2 mux_2x1_ibr_0/I1 OUT mux_2x1_ibr_0/I0 VDD VSS mux_2x1_ibr
.ends

.subckt CLK_div_96_mag CLK Vdiv96 RST VSS VDD
XJK_FF_mag_0 RST VDD VDD JK_FF_mag_0/nand2_mag_1/m1_186_70# JK_FF_mag_0/nand3_mag_2/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_0/nand2_mag_3/m1_186_70# JK_FF_mag_0/nand3_mag_0/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_0/nand2_mag_2/m1_186_70# JK_FF_mag_0/nand2_mag_4/m1_186_70# JK_FF_mag_0/nand3_mag_1/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_0/nand2_mag_4/IN2 JK_FF_mag_0/nand3_mag_0/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_0/nand3_mag_2/nmos_3p3_VGTVWA_0/a_28_n66# JK_FF_mag_0/nand2_mag_1/IN2
+ JK_FF_mag_0/nand3_mag_2/OUT JK_FF_mag_0/nand3_mag_0/OUT JK_FF_mag_5/Q JK_FF_mag_0/QB
+ JK_FF_mag_0/nand3_mag_1/IN1 JK_FF_mag_0/nand2_mag_3/IN1 JK_FF_mag_0/nand3_mag_1/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_0/nand2_mag_0/m1_186_70# JK_FF_mag_0/Q JK_FF_mag_0/nand3_mag_1/OUT VSS
+ VDD JK_FF_mag
XJK_FF_mag_2 RST VDD VDD JK_FF_mag_2/nand2_mag_1/m1_186_70# JK_FF_mag_2/nand3_mag_2/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_2/nand2_mag_3/m1_186_70# JK_FF_mag_2/nand3_mag_0/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_2/nand2_mag_2/m1_186_70# JK_FF_mag_2/nand2_mag_4/m1_186_70# JK_FF_mag_2/nand3_mag_1/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_2/nand2_mag_4/IN2 JK_FF_mag_2/nand3_mag_0/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_2/nand3_mag_2/nmos_3p3_VGTVWA_0/a_28_n66# JK_FF_mag_2/nand2_mag_1/IN2
+ JK_FF_mag_2/nand3_mag_2/OUT JK_FF_mag_2/nand3_mag_0/OUT JK_FF_mag_0/Q JK_FF_mag_2/QB
+ JK_FF_mag_2/nand3_mag_1/IN1 JK_FF_mag_2/nand2_mag_3/IN1 JK_FF_mag_2/nand3_mag_1/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_2/nand2_mag_0/m1_186_70# JK_FF_mag_2/Q JK_FF_mag_2/nand3_mag_1/OUT VSS
+ VDD JK_FF_mag
XJK_FF_mag_3 RST VDD VDD JK_FF_mag_3/nand2_mag_1/m1_186_70# JK_FF_mag_3/nand3_mag_2/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_3/nand2_mag_3/m1_186_70# JK_FF_mag_3/nand3_mag_0/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_3/nand2_mag_2/m1_186_70# JK_FF_mag_3/nand2_mag_4/m1_186_70# JK_FF_mag_3/nand3_mag_1/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_3/nand2_mag_4/IN2 JK_FF_mag_3/nand3_mag_0/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_3/nand3_mag_2/nmos_3p3_VGTVWA_0/a_28_n66# JK_FF_mag_3/nand2_mag_1/IN2
+ JK_FF_mag_3/nand3_mag_2/OUT JK_FF_mag_3/nand3_mag_0/OUT JK_FF_mag_2/Q JK_FF_mag_3/QB
+ JK_FF_mag_3/nand3_mag_1/IN1 JK_FF_mag_3/nand2_mag_3/IN1 JK_FF_mag_3/nand3_mag_1/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_3/nand2_mag_0/m1_186_70# JK_FF_mag_3/Q JK_FF_mag_3/nand3_mag_1/OUT VSS
+ VDD JK_FF_mag
XJK_FF_mag_4 RST VDD VDD JK_FF_mag_4/nand2_mag_1/m1_186_70# JK_FF_mag_4/nand3_mag_2/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_4/nand2_mag_3/m1_186_70# JK_FF_mag_4/nand3_mag_0/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_4/nand2_mag_2/m1_186_70# JK_FF_mag_4/nand2_mag_4/m1_186_70# JK_FF_mag_4/nand3_mag_1/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_4/nand2_mag_4/IN2 JK_FF_mag_4/nand3_mag_0/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_4/nand3_mag_2/nmos_3p3_VGTVWA_0/a_28_n66# JK_FF_mag_4/nand2_mag_1/IN2
+ JK_FF_mag_4/nand3_mag_2/OUT JK_FF_mag_4/nand3_mag_0/OUT CLK JK_FF_mag_4/QB JK_FF_mag_4/nand3_mag_1/IN1
+ JK_FF_mag_4/nand2_mag_3/IN1 JK_FF_mag_4/nand3_mag_1/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_4/nand2_mag_0/m1_186_70# JK_FF_mag_4/Q JK_FF_mag_4/nand3_mag_1/OUT VSS
+ VDD JK_FF_mag
XJK_FF_mag_5 RST VDD VDD JK_FF_mag_5/nand2_mag_1/m1_186_70# JK_FF_mag_5/nand3_mag_2/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_5/nand2_mag_3/m1_186_70# JK_FF_mag_5/nand3_mag_0/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_5/nand2_mag_2/m1_186_70# JK_FF_mag_5/nand2_mag_4/m1_186_70# JK_FF_mag_5/nand3_mag_1/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_5/nand2_mag_4/IN2 JK_FF_mag_5/nand3_mag_0/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_5/nand3_mag_2/nmos_3p3_VGTVWA_0/a_28_n66# JK_FF_mag_5/nand2_mag_1/IN2
+ JK_FF_mag_5/nand3_mag_2/OUT JK_FF_mag_5/nand3_mag_0/OUT JK_FF_mag_4/Q JK_FF_mag_5/QB
+ JK_FF_mag_5/nand3_mag_1/IN1 JK_FF_mag_5/nand2_mag_3/IN1 JK_FF_mag_5/nand3_mag_1/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_5/nand2_mag_0/m1_186_70# JK_FF_mag_5/Q JK_FF_mag_5/nand3_mag_1/OUT VSS
+ VDD JK_FF_mag
XCLK_div_3_mag_0 CLK_div_3_mag_0/Q1 CLK_div_3_mag_0/Q0 Vdiv96 CLK_div_3_mag_0/JK_FF_mag_1/nand3_mag_0/OUT
+ CLK_div_3_mag_0/JK_FF_mag_0/nand3_mag_0/OUT CLK_div_3_mag_0/JK_FF_mag_1/nand3_mag_1/OUT
+ CLK_div_3_mag_0/JK_FF_mag_0/nand3_mag_1/OUT CLK_div_3_mag_0/JK_FF_mag_1/nand3_mag_2/OUT
+ VSS JK_FF_mag_3/Q RST CLK_div_3_mag_0/JK_FF_mag_0/nand3_mag_2/OUT VDD CLK_div_3_mag
.ends

.subckt Buffer_Delayed1_mag IN OUT VDD VSS
XInverter_delayed_mag_11 VSS Inverter_delayed_mag_11/IN Inverter_delayed_mag_10/IN
+ VDD Inverter_delayed_mag
XInverter_delayed_mag_13 VSS Inverter_delayed_mag_13/IN Inverter_delayed_mag_12/IN
+ VDD Inverter_delayed_mag
XInverter_delayed_mag_12 VSS Inverter_delayed_mag_12/IN Inverter_delayed_mag_11/IN
+ VDD Inverter_delayed_mag
XInverter_delayed_mag_14 VSS Inverter_delayed_mag_14/IN Inverter_delayed_mag_13/IN
+ VDD Inverter_delayed_mag
XInverter_delayed_mag_15 VSS IN Inverter_delayed_mag_14/IN VDD Inverter_delayed_mag
XInverter_delayed_mag_0 VSS Inverter_delayed_mag_0/IN Inverter_delayed_mag_3/IN VDD
+ Inverter_delayed_mag
XInverter_delayed_mag_1 VSS Inverter_delayed_mag_1/IN Inverter_delayed_mag_2/IN VDD
+ Inverter_delayed_mag
XInverter_delayed_mag_2 VSS Inverter_delayed_mag_2/IN Inverter_delayed_mag_0/IN VDD
+ Inverter_delayed_mag
XInverter_delayed_mag_3 VSS Inverter_delayed_mag_3/IN Inverter_delayed_mag_4/IN VDD
+ Inverter_delayed_mag
XInverter_delayed_mag_4 VSS Inverter_delayed_mag_4/IN Inverter_delayed_mag_5/IN VDD
+ Inverter_delayed_mag
XInverter_delayed_mag_5 VSS Inverter_delayed_mag_5/IN Inverter_delayed_mag_6/IN VDD
+ Inverter_delayed_mag
XInverter_delayed_mag_6 VSS Inverter_delayed_mag_6/IN Inverter_delayed_mag_7/IN VDD
+ Inverter_delayed_mag
XInverter_delayed_mag_7 VSS Inverter_delayed_mag_7/IN OUT VDD Inverter_delayed_mag
XInverter_delayed_mag_8 VSS Inverter_delayed_mag_8/IN Inverter_delayed_mag_1/IN VDD
+ Inverter_delayed_mag
XInverter_delayed_mag_9 VSS Inverter_delayed_mag_9/IN Inverter_delayed_mag_8/IN VDD
+ Inverter_delayed_mag
XInverter_delayed_mag_10 VSS Inverter_delayed_mag_10/IN Inverter_delayed_mag_9/IN
+ VDD Inverter_delayed_mag
.ends

.subckt and_5_mag A B C D E VOUT VDD VSS
Xand2_mag_1 and2_mag_1/IN2 C and2_mag_2/IN2 VDD VSS and2_mag
Xand2_mag_0 B A and2_mag_1/IN2 VDD VSS and2_mag
Xand2_mag_2 and2_mag_2/IN2 D and2_mag_3/IN2 VDD VSS and2_mag
Xand2_mag_3 and2_mag_3/IN2 E VOUT VDD VSS and2_mag
.ends

.subckt nand_5_mag A B D OUT E C VDD VSS
XGF_INV_MAG_0 GF_INV_MAG_0/IN OUT VSS VDD GF_INV_MAG
Xand_5_mag_0 A B C D E GF_INV_MAG_0/IN VDD VSS and_5_mag
.ends

.subckt CLK_div_31_mag Vdiv31 CLK Q0 Q1 Q2 Q3 Q4 RST VSS VDD
XJK_FF_mag_1 RST VDD VDD JK_FF_mag_1/nand2_mag_1/m1_186_70# JK_FF_mag_1/nand3_mag_2/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_1/nand2_mag_3/m1_186_70# JK_FF_mag_1/nand3_mag_0/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_1/nand2_mag_2/m1_186_70# JK_FF_mag_1/nand2_mag_4/m1_186_70# JK_FF_mag_1/nand3_mag_1/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_1/nand2_mag_4/IN2 JK_FF_mag_1/nand3_mag_0/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_1/nand3_mag_2/nmos_3p3_VGTVWA_0/a_28_n66# JK_FF_mag_1/nand2_mag_1/IN2
+ JK_FF_mag_1/nand3_mag_2/OUT JK_FF_mag_1/nand3_mag_0/OUT Q2 JK_FF_mag_1/QB JK_FF_mag_1/nand3_mag_1/IN1
+ JK_FF_mag_1/nand2_mag_3/IN1 JK_FF_mag_1/nand3_mag_1/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_1/nand2_mag_0/m1_186_70# Q3 JK_FF_mag_1/nand3_mag_1/OUT VSS VDD JK_FF_mag
XJK_FF_mag_0 RST VDD VDD JK_FF_mag_0/nand2_mag_1/m1_186_70# JK_FF_mag_0/nand3_mag_2/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_0/nand2_mag_3/m1_186_70# JK_FF_mag_0/nand3_mag_0/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_0/nand2_mag_2/m1_186_70# JK_FF_mag_0/nand2_mag_4/m1_186_70# JK_FF_mag_0/nand3_mag_1/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_0/nand2_mag_4/IN2 JK_FF_mag_0/nand3_mag_0/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_0/nand3_mag_2/nmos_3p3_VGTVWA_0/a_28_n66# JK_FF_mag_0/nand2_mag_1/IN2
+ JK_FF_mag_0/nand3_mag_2/OUT JK_FF_mag_0/nand3_mag_0/OUT Q1 JK_FF_mag_0/QB JK_FF_mag_0/nand3_mag_1/IN1
+ JK_FF_mag_0/nand2_mag_3/IN1 JK_FF_mag_0/nand3_mag_1/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_0/nand2_mag_0/m1_186_70# Q2 JK_FF_mag_0/nand3_mag_1/OUT VSS VDD JK_FF_mag
XJK_FF_mag_2 RST VDD VDD JK_FF_mag_2/nand2_mag_1/m1_186_70# JK_FF_mag_2/nand3_mag_2/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_2/nand2_mag_3/m1_186_70# JK_FF_mag_2/nand3_mag_0/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_2/nand2_mag_2/m1_186_70# JK_FF_mag_2/nand2_mag_4/m1_186_70# JK_FF_mag_2/nand3_mag_1/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_2/nand2_mag_4/IN2 JK_FF_mag_2/nand3_mag_0/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_2/nand3_mag_2/nmos_3p3_VGTVWA_0/a_28_n66# JK_FF_mag_2/nand2_mag_1/IN2
+ JK_FF_mag_2/nand3_mag_2/OUT JK_FF_mag_2/nand3_mag_0/OUT Q0 JK_FF_mag_2/QB JK_FF_mag_2/nand3_mag_1/IN1
+ JK_FF_mag_2/nand2_mag_3/IN1 JK_FF_mag_2/nand3_mag_1/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_2/nand2_mag_0/m1_186_70# Q1 JK_FF_mag_2/nand3_mag_1/OUT VSS VDD JK_FF_mag
XBuffer_Delayed1_mag_0 and_5_mag_0/VOUT or_2_mag_0/IN1 VDD VSS Buffer_Delayed1_mag
XJK_FF_mag_3 RST VDD VDD JK_FF_mag_3/nand2_mag_1/m1_186_70# JK_FF_mag_3/nand3_mag_2/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_3/nand2_mag_3/m1_186_70# JK_FF_mag_3/nand3_mag_0/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_3/nand2_mag_2/m1_186_70# JK_FF_mag_3/nand2_mag_4/m1_186_70# JK_FF_mag_3/nand3_mag_1/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_3/nand2_mag_4/IN2 JK_FF_mag_3/nand3_mag_0/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_3/nand3_mag_2/nmos_3p3_VGTVWA_0/a_28_n66# JK_FF_mag_3/nand2_mag_1/IN2
+ JK_FF_mag_3/nand3_mag_2/OUT JK_FF_mag_3/nand3_mag_0/OUT CLK JK_FF_mag_3/QB JK_FF_mag_3/nand3_mag_1/IN1
+ JK_FF_mag_3/nand2_mag_3/IN1 JK_FF_mag_3/nand3_mag_1/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_3/nand2_mag_0/m1_186_70# Q0 JK_FF_mag_3/nand3_mag_1/OUT VSS VDD JK_FF_mag
XJK_FF_mag_4 RST VDD VDD JK_FF_mag_4/nand2_mag_1/m1_186_70# JK_FF_mag_4/nand3_mag_2/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_4/nand2_mag_3/m1_186_70# JK_FF_mag_4/nand3_mag_0/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_4/nand2_mag_2/m1_186_70# JK_FF_mag_4/nand2_mag_4/m1_186_70# JK_FF_mag_4/nand3_mag_1/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_4/nand2_mag_4/IN2 JK_FF_mag_4/nand3_mag_0/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_4/nand3_mag_2/nmos_3p3_VGTVWA_0/a_28_n66# JK_FF_mag_4/nand2_mag_1/IN2
+ JK_FF_mag_4/nand3_mag_2/OUT JK_FF_mag_4/nand3_mag_0/OUT Q3 JK_FF_mag_4/QB JK_FF_mag_4/nand3_mag_1/IN1
+ JK_FF_mag_4/nand2_mag_3/IN1 JK_FF_mag_4/nand3_mag_1/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_4/nand2_mag_0/m1_186_70# Q4 JK_FF_mag_4/nand3_mag_1/OUT VSS VDD JK_FF_mag
Xor_2_mag_0 VSS Q4 or_2_mag_0/IN1 Vdiv31 VDD or_2_mag
Xand_5_mag_0 Q1 Q0 Q3 Q2 CLK and_5_mag_0/VOUT VDD VSS and_5_mag
Xnand_5_mag_0 Q4 Q0 Q3 RST Q1 Q2 VDD VSS nand_5_mag
.ends

.subckt CLK_div_93_mag VDD Vdiv93 RST CLK VSS
XCLK_div_31_mag_0 CLK_div_3_mag_0/CLK CLK CLK_div_31_mag_0/Q0 CLK_div_31_mag_0/Q1
+ CLK_div_31_mag_0/Q2 CLK_div_31_mag_0/Q3 CLK_div_31_mag_0/Q4 RST VSS VDD CLK_div_31_mag
XCLK_div_3_mag_0 CLK_div_3_mag_0/Q1 CLK_div_3_mag_0/Q0 Vdiv93 CLK_div_3_mag_0/JK_FF_mag_1/nand3_mag_0/OUT
+ CLK_div_3_mag_0/JK_FF_mag_0/nand3_mag_0/OUT CLK_div_3_mag_0/JK_FF_mag_1/nand3_mag_1/OUT
+ CLK_div_3_mag_0/JK_FF_mag_0/nand3_mag_1/OUT CLK_div_3_mag_0/JK_FF_mag_1/nand3_mag_2/OUT
+ VSS CLK_div_3_mag_0/CLK RST CLK_div_3_mag_0/JK_FF_mag_0/nand3_mag_2/OUT VDD CLK_div_3_mag
.ends

.subckt CLK_div_10_mag CLK Q0 Q1 Q2 Q3 Vdiv10 VDD VSS RST
XJK_FF_mag_1 RST VDD VDD JK_FF_mag_1/nand2_mag_1/m1_186_70# JK_FF_mag_1/nand3_mag_2/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_1/nand2_mag_3/m1_186_70# JK_FF_mag_1/nand3_mag_0/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_1/nand2_mag_2/m1_186_70# JK_FF_mag_1/nand2_mag_4/m1_186_70# JK_FF_mag_1/nand3_mag_1/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_1/nand2_mag_4/IN2 JK_FF_mag_1/nand3_mag_0/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_1/nand3_mag_2/nmos_3p3_VGTVWA_0/a_28_n66# JK_FF_mag_1/nand2_mag_1/IN2
+ JK_FF_mag_1/nand3_mag_2/OUT JK_FF_mag_1/nand3_mag_0/OUT CLK JK_FF_mag_1/QB JK_FF_mag_1/nand3_mag_1/IN1
+ JK_FF_mag_1/nand2_mag_3/IN1 JK_FF_mag_1/nand3_mag_1/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_1/nand2_mag_0/m1_186_70# Q0 JK_FF_mag_1/nand3_mag_1/OUT VSS VDD JK_FF_mag
XJK_FF_mag_0 RST VDD JK_FF_mag_0/K JK_FF_mag_0/nand2_mag_1/m1_186_70# JK_FF_mag_0/nand3_mag_2/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_0/nand2_mag_3/m1_186_70# JK_FF_mag_0/nand3_mag_0/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_0/nand2_mag_2/m1_186_70# JK_FF_mag_0/nand2_mag_4/m1_186_70# JK_FF_mag_0/nand3_mag_1/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_0/nand2_mag_4/IN2 JK_FF_mag_0/nand3_mag_0/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_0/nand3_mag_2/nmos_3p3_VGTVWA_0/a_28_n66# JK_FF_mag_0/nand2_mag_1/IN2
+ JK_FF_mag_0/nand3_mag_2/OUT JK_FF_mag_0/nand3_mag_0/OUT Q0 JK_FF_mag_2/K JK_FF_mag_0/nand3_mag_1/IN1
+ JK_FF_mag_0/nand2_mag_3/IN1 JK_FF_mag_0/nand3_mag_1/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_0/nand2_mag_0/m1_186_70# Q3 JK_FF_mag_0/nand3_mag_1/OUT VSS VDD JK_FF_mag
XJK_FF_mag_2 RST VDD JK_FF_mag_2/K JK_FF_mag_2/nand2_mag_1/m1_186_70# JK_FF_mag_2/nand3_mag_2/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_2/nand2_mag_3/m1_186_70# JK_FF_mag_2/nand3_mag_0/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_2/nand2_mag_2/m1_186_70# JK_FF_mag_2/nand2_mag_4/m1_186_70# JK_FF_mag_2/nand3_mag_1/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_2/nand2_mag_4/IN2 JK_FF_mag_2/nand3_mag_0/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_2/nand3_mag_2/nmos_3p3_VGTVWA_0/a_28_n66# JK_FF_mag_2/nand2_mag_1/IN2
+ JK_FF_mag_2/nand3_mag_2/OUT JK_FF_mag_2/nand3_mag_0/OUT Q0 JK_FF_mag_2/QB JK_FF_mag_2/nand3_mag_1/IN1
+ JK_FF_mag_2/nand2_mag_3/IN1 JK_FF_mag_2/nand3_mag_1/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_2/nand2_mag_0/m1_186_70# Q1 JK_FF_mag_2/nand3_mag_1/OUT VSS VDD JK_FF_mag
XJK_FF_mag_3 RST VDD VDD JK_FF_mag_3/nand2_mag_1/m1_186_70# JK_FF_mag_3/nand3_mag_2/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_3/nand2_mag_3/m1_186_70# JK_FF_mag_3/nand3_mag_0/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_3/nand2_mag_2/m1_186_70# JK_FF_mag_3/nand2_mag_4/m1_186_70# JK_FF_mag_3/nand3_mag_1/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_3/nand2_mag_4/IN2 JK_FF_mag_3/nand3_mag_0/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_3/nand3_mag_2/nmos_3p3_VGTVWA_0/a_28_n66# JK_FF_mag_3/nand2_mag_1/IN2
+ JK_FF_mag_3/nand3_mag_2/OUT JK_FF_mag_3/nand3_mag_0/OUT Q1 JK_FF_mag_3/QB JK_FF_mag_3/nand3_mag_1/IN1
+ JK_FF_mag_3/nand2_mag_3/IN1 JK_FF_mag_3/nand3_mag_1/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_3/nand2_mag_0/m1_186_70# Q2 JK_FF_mag_3/nand3_mag_1/OUT VSS VDD JK_FF_mag
Xand2_mag_1 Q0 Q2 and2_mag_1/OUT VDD VSS and2_mag
Xand2_mag_0 Q1 Q2 and2_mag_0/OUT VDD VSS and2_mag
Xand2_mag_2 Q2 Q1 JK_FF_mag_0/K VDD VSS and2_mag
XBuffer_delayed_mag_0 and2_mag_1/OUT nor_3_mag_0/IN3 VDD VSS Buffer_delayed_mag
Xnor_3_mag_0 nor_3_mag_0/IN3 and2_mag_0/OUT Q3 Vdiv10 VSS VDD nor_3_mag
.ends

.subckt CLK_div_105_mag CLK Vdiv100 RST VDD VSS
XCLK_div_10_mag_0 CLK CLK_div_10_mag_0/Q0 CLK_div_10_mag_0/Q1 CLK_div_10_mag_0/Q2
+ CLK_div_10_mag_0/Q3 CLK_div_10_mag_1/CLK VDD VSS RST CLK_div_10_mag
XCLK_div_10_mag_1 CLK_div_10_mag_1/CLK CLK_div_10_mag_1/Q0 CLK_div_10_mag_1/Q1 CLK_div_10_mag_1/Q2
+ CLK_div_10_mag_1/Q3 Vdiv100 VDD VSS RST CLK_div_10_mag
.ends

.subckt CLK_div_90_mag Vdiv90 VDD CLK RST VSS
XCLK_div_3_mag_1 CLK_div_3_mag_1/Q1 CLK_div_3_mag_1/Q0 CLK_div_3_mag_0/CLK CLK_div_3_mag_1/JK_FF_mag_1/nand3_mag_0/OUT
+ CLK_div_3_mag_1/JK_FF_mag_0/nand3_mag_0/OUT CLK_div_3_mag_1/JK_FF_mag_1/nand3_mag_1/OUT
+ CLK_div_3_mag_1/JK_FF_mag_0/nand3_mag_1/OUT CLK_div_3_mag_1/JK_FF_mag_1/nand3_mag_2/OUT
+ VSS CLK RST CLK_div_3_mag_1/JK_FF_mag_0/nand3_mag_2/OUT VDD CLK_div_3_mag
XCLK_div_3_mag_0 CLK_div_3_mag_0/Q1 CLK_div_3_mag_0/Q0 CLK_div_10_mag_0/CLK CLK_div_3_mag_0/JK_FF_mag_1/nand3_mag_0/OUT
+ CLK_div_3_mag_0/JK_FF_mag_0/nand3_mag_0/OUT CLK_div_3_mag_0/JK_FF_mag_1/nand3_mag_1/OUT
+ CLK_div_3_mag_0/JK_FF_mag_0/nand3_mag_1/OUT CLK_div_3_mag_0/JK_FF_mag_1/nand3_mag_2/OUT
+ VSS CLK_div_3_mag_0/CLK RST CLK_div_3_mag_0/JK_FF_mag_0/nand3_mag_2/OUT VDD CLK_div_3_mag
XCLK_div_10_mag_0 CLK_div_10_mag_0/CLK CLK_div_10_mag_0/Q0 CLK_div_10_mag_0/Q1 CLK_div_10_mag_0/Q2
+ CLK_div_10_mag_0/Q3 Vdiv90 VDD VSS RST CLK_div_10_mag
.ends

.subckt CLK_div_100_mag CLK Vdiv100 RST VDD VSS
XCLK_div_10_mag_0 CLK CLK_div_10_mag_0/Q0 CLK_div_10_mag_0/Q1 CLK_div_10_mag_0/Q2
+ CLK_div_10_mag_0/Q3 CLK_div_10_mag_1/CLK VDD VSS RST CLK_div_10_mag
XCLK_div_10_mag_1 CLK_div_10_mag_1/CLK CLK_div_10_mag_1/Q0 CLK_div_10_mag_1/Q1 CLK_div_10_mag_1/Q2
+ CLK_div_10_mag_1/Q3 Vdiv100 VDD VSS RST CLK_div_10_mag
.ends

.subckt nand3_mag_ibr IN3 IN2 IN1 VDD VSS OUT
Xnmos_3p3_VGTVWA_0 nmos_3p3_VGTVWA_1/a_28_n66# nmos_3p3_VGTVWA_0/a_28_n66# IN2 VSS
+ nmos_3p3_VGTVWA
Xnmos_3p3_VGTVWA_1 VSS nmos_3p3_VGTVWA_1/a_28_n66# IN3 VSS nmos_3p3_VGTVWA
Xnmos_3p3_VGTVWA_2 nmos_3p3_VGTVWA_0/a_28_n66# OUT IN1 VSS nmos_3p3_VGTVWA
Xpmos_3p3_M8SWPS_0 IN1 VDD OUT VDD pmos_3p3_M8SWPS
Xpmos_3p3_M8SWPS_1 IN3 VDD OUT VDD pmos_3p3_M8SWPS
Xpmos_3p3_M8SWPS_2 IN2 OUT VDD VDD pmos_3p3_M8SWPS
.ends

.subckt and_3_ibr IN2 IN3 VDD OUT IN1 nand3_mag_ibr_0/OUT VSS
Xnverterlayout_ibr_0 VDD VSS OUT nand3_mag_ibr_0/OUT nverterlayout_ibr
Xnand3_mag_ibr_0 IN3 IN2 IN1 VDD VSS nand3_mag_ibr_0/OUT nand3_mag_ibr
.ends

.subckt dec3x8_ibr_mag IN1 IN2 IN3 D0 D1 D2 D3 D4 D5 D6 VSS and_3_ibr_0/nand3_mag_ibr_0/OUT
+ and_3_ibr_2/nand3_mag_ibr_0/OUT and_3_ibr_4/nand3_mag_ibr_0/OUT and_3_ibr_6/nand3_mag_ibr_0/OUT
+ VDD D7 and_3_ibr_1/nand3_mag_ibr_0/OUT and_3_ibr_3/nand3_mag_ibr_0/OUT and_3_ibr_5/nand3_mag_ibr_0/OUT
+ and_3_ibr_7/nand3_mag_ibr_0/OUT
Xand_3_ibr_1 IN2 and_3_ibr_5/IN3 VDD D2 and_3_ibr_3/IN1 and_3_ibr_1/nand3_mag_ibr_0/OUT
+ VSS and_3_ibr
Xand_3_ibr_0 and_3_ibr_6/IN3 and_3_ibr_5/IN3 VDD D0 and_3_ibr_3/IN1 and_3_ibr_0/nand3_mag_ibr_0/OUT
+ VSS and_3_ibr
Xand_3_ibr_2 IN1 and_3_ibr_6/IN3 VDD D4 and_3_ibr_3/IN1 and_3_ibr_2/nand3_mag_ibr_0/OUT
+ VSS and_3_ibr
Xand_3_ibr_3 IN2 IN1 VDD D6 and_3_ibr_3/IN1 and_3_ibr_3/nand3_mag_ibr_0/OUT VSS and_3_ibr
Xand_3_ibr_4 and_3_ibr_5/IN3 and_3_ibr_6/IN3 VDD D1 IN3 and_3_ibr_4/nand3_mag_ibr_0/OUT
+ VSS and_3_ibr
Xand_3_ibr_5 IN2 and_3_ibr_5/IN3 VDD D3 IN3 and_3_ibr_5/nand3_mag_ibr_0/OUT VSS and_3_ibr
Xand_3_ibr_6 IN1 and_3_ibr_6/IN3 VDD D5 IN3 and_3_ibr_6/nand3_mag_ibr_0/OUT VSS and_3_ibr
Xand_3_ibr_7 IN2 IN1 VDD D7 IN3 and_3_ibr_7/nand3_mag_ibr_0/OUT VSS and_3_ibr
Xnverterlayout_ibr_0 VDD VSS and_3_ibr_3/IN1 IN3 nverterlayout_ibr
Xnverterlayout_ibr_2 VDD VSS and_3_ibr_5/IN3 IN1 nverterlayout_ibr
Xnverterlayout_ibr_1 VDD VSS and_3_ibr_6/IN3 IN2 nverterlayout_ibr
.ends

.subckt CLK_div_110_mag CLK Vdiv110 RST VDD VSS
XCLK_DIV_11_mag_new_0 CLK CLK_div_10_mag_0/CLK CLK_DIV_11_mag_new_0/Q3 CLK_DIV_11_mag_new_0/Q2
+ CLK_DIV_11_mag_new_0/Q1 CLK_DIV_11_mag_new_0/Q0 VDD RST VSS CLK_DIV_11_mag_new
XCLK_div_10_mag_0 CLK_div_10_mag_0/CLK CLK_div_10_mag_0/Q0 CLK_div_10_mag_0/Q1 CLK_div_10_mag_0/Q2
+ CLK_div_10_mag_0/Q3 Vdiv110 VDD VSS RST CLK_div_10_mag
.ends

.subckt CLK_div_108_new_mag VDD Vdiv108 CLK VSS RST
XJK_FF_mag_1 RST VDD VDD JK_FF_mag_1/nand2_mag_1/m1_186_70# JK_FF_mag_1/nand3_mag_2/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_1/nand2_mag_3/m1_186_70# JK_FF_mag_1/nand3_mag_0/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_1/nand2_mag_2/m1_186_70# JK_FF_mag_1/nand2_mag_4/m1_186_70# JK_FF_mag_1/nand3_mag_1/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_1/nand2_mag_4/IN2 JK_FF_mag_1/nand3_mag_0/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_1/nand3_mag_2/nmos_3p3_VGTVWA_0/a_28_n66# JK_FF_mag_1/nand2_mag_1/IN2
+ JK_FF_mag_1/nand3_mag_2/OUT JK_FF_mag_1/nand3_mag_0/OUT JK_FF_mag_1/CLK JK_FF_mag_1/QB
+ JK_FF_mag_1/nand3_mag_1/IN1 JK_FF_mag_1/nand2_mag_3/IN1 JK_FF_mag_1/nand3_mag_1/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_1/nand2_mag_0/m1_186_70# JK_FF_mag_1/Q JK_FF_mag_1/nand3_mag_1/OUT VSS
+ VDD JK_FF_mag
XJK_FF_mag_0 RST VDD VDD JK_FF_mag_0/nand2_mag_1/m1_186_70# JK_FF_mag_0/nand3_mag_2/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_0/nand2_mag_3/m1_186_70# JK_FF_mag_0/nand3_mag_0/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_0/nand2_mag_2/m1_186_70# JK_FF_mag_0/nand2_mag_4/m1_186_70# JK_FF_mag_0/nand3_mag_1/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_0/nand2_mag_4/IN2 JK_FF_mag_0/nand3_mag_0/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_0/nand3_mag_2/nmos_3p3_VGTVWA_0/a_28_n66# JK_FF_mag_0/nand2_mag_1/IN2
+ JK_FF_mag_0/nand3_mag_2/OUT JK_FF_mag_0/nand3_mag_0/OUT JK_FF_mag_1/Q JK_FF_mag_0/QB
+ JK_FF_mag_0/nand3_mag_1/IN1 JK_FF_mag_0/nand2_mag_3/IN1 JK_FF_mag_0/nand3_mag_1/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_0/nand2_mag_0/m1_186_70# Vdiv108 JK_FF_mag_0/nand3_mag_1/OUT VSS VDD JK_FF_mag
XCLK_div_3_mag_1 CLK_div_3_mag_1/Q1 CLK_div_3_mag_1/Q0 CLK_div_3_mag_0/CLK CLK_div_3_mag_1/JK_FF_mag_1/nand3_mag_0/OUT
+ CLK_div_3_mag_1/JK_FF_mag_0/nand3_mag_0/OUT CLK_div_3_mag_1/JK_FF_mag_1/nand3_mag_1/OUT
+ CLK_div_3_mag_1/JK_FF_mag_0/nand3_mag_1/OUT CLK_div_3_mag_1/JK_FF_mag_1/nand3_mag_2/OUT
+ VSS CLK_div_3_mag_1/CLK RST CLK_div_3_mag_1/JK_FF_mag_0/nand3_mag_2/OUT VDD CLK_div_3_mag
XCLK_div_3_mag_0 CLK_div_3_mag_0/Q1 CLK_div_3_mag_0/Q0 JK_FF_mag_1/CLK CLK_div_3_mag_0/JK_FF_mag_1/nand3_mag_0/OUT
+ CLK_div_3_mag_0/JK_FF_mag_0/nand3_mag_0/OUT CLK_div_3_mag_0/JK_FF_mag_1/nand3_mag_1/OUT
+ CLK_div_3_mag_0/JK_FF_mag_0/nand3_mag_1/OUT CLK_div_3_mag_0/JK_FF_mag_1/nand3_mag_2/OUT
+ VSS CLK_div_3_mag_0/CLK RST CLK_div_3_mag_0/JK_FF_mag_0/nand3_mag_2/OUT VDD CLK_div_3_mag
XCLK_div_3_mag_2 CLK_div_3_mag_2/Q1 CLK_div_3_mag_2/Q0 CLK_div_3_mag_1/CLK CLK_div_3_mag_2/JK_FF_mag_1/nand3_mag_0/OUT
+ CLK_div_3_mag_2/JK_FF_mag_0/nand3_mag_0/OUT CLK_div_3_mag_2/JK_FF_mag_1/nand3_mag_1/OUT
+ CLK_div_3_mag_2/JK_FF_mag_0/nand3_mag_1/OUT CLK_div_3_mag_2/JK_FF_mag_1/nand3_mag_2/OUT
+ VSS CLK RST CLK_div_3_mag_2/JK_FF_mag_0/nand3_mag_2/OUT VDD CLK_div_3_mag
.ends

.subckt Feedback_Divider_mag CLK RST F2 F1 F0 Vdiv VDD Vdiv90 Vdiv96 Vdiv93 Vdiv99
+ Vdiv110 Vdiv108 Vdiv100 Vdiv105 VDD90 VDD99 VDD108 VDD100 VDD105 VDD93 VDD96 VDD110
+ VSS
XCLK_div_99_mag_0 VDD99 CLK Vdiv99 RST VSS CLK_div_99_mag
Xmux_8x1_ibr_0 Vdiv90 Vdiv93 Vdiv96 Vdiv99 Vdiv105 Vdiv108 Vdiv110 Vdiv F0 F1 F2 Vdiv100
+ VSS VDD mux_8x1_ibr
XCLK_div_96_mag_0 CLK Vdiv96 RST VSS VDD96 CLK_div_96_mag
XCLK_div_93_mag_0 VDD93 Vdiv93 RST CLK VSS CLK_div_93_mag
XCLK_div_105_mag_0 CLK Vdiv105 RST VDD105 VSS CLK_div_105_mag
XCLK_div_90_mag_0 Vdiv90 VDD90 CLK RST VSS CLK_div_90_mag
XCLK_div_100_mag_0 CLK Vdiv100 RST VDD100 VSS CLK_div_100_mag
Xdec3x8_ibr_mag_0 F2 F1 F0 VDD90 VDD93 VDD96 VDD99 VDD100 VDD105 VDD108 VSS dec3x8_ibr_mag_0/and_3_ibr_0/nand3_mag_ibr_0/OUT
+ dec3x8_ibr_mag_0/and_3_ibr_2/nand3_mag_ibr_0/OUT dec3x8_ibr_mag_0/and_3_ibr_4/nand3_mag_ibr_0/OUT
+ dec3x8_ibr_mag_0/and_3_ibr_6/nand3_mag_ibr_0/OUT VDD VDD110 dec3x8_ibr_mag_0/and_3_ibr_1/nand3_mag_ibr_0/OUT
+ dec3x8_ibr_mag_0/and_3_ibr_3/nand3_mag_ibr_0/OUT dec3x8_ibr_mag_0/and_3_ibr_5/nand3_mag_ibr_0/OUT
+ dec3x8_ibr_mag_0/and_3_ibr_7/nand3_mag_ibr_0/OUT dec3x8_ibr_mag
XCLK_div_110_mag_0 CLK Vdiv110 RST VDD110 VSS CLK_div_110_mag
XCLK_div_108_new_mag_0 VDD108 Vdiv108 CLK VSS RST CLK_div_108_new_mag
.ends

.subckt nmos_3p3_6FEA4B a_n52_n50# a_256_n94# a_52_n94# a_356_n50# a_n256_n50# a_n444_n50#
+ a_152_n50# a_n356_n94# a_n152_n94# VSUBS
X0 a_152_n50# a_52_n94# a_n52_n50# VSUBS nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1 a_n52_n50# a_n152_n94# a_n256_n50# VSUBS nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X2 a_n256_n50# a_n356_n94# a_n444_n50# VSUBS nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X3 a_356_n50# a_256_n94# a_152_n50# VSUBS nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
.ends

.subckt pmos_3p3_KYEELV a_152_68# a_n444_n168# a_n256_68# a_n52_68# a_52_24# a_152_n168#
+ a_n444_68# a_356_68# a_256_n212# a_n256_n168# a_n356_n212# a_n152_24# w_n530_n298#
+ a_52_n212# a_n52_n168# a_n152_n212# a_n356_24# a_356_n168# a_256_24#
X0 a_n256_n168# a_n356_n212# a_n444_n168# w_n530_n298# pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X1 a_356_n168# a_256_n212# a_152_n168# w_n530_n298# pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X2 a_152_68# a_52_24# a_n52_68# w_n530_n298# pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X3 a_n52_68# a_n152_24# a_n256_68# w_n530_n298# pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X4 a_152_n168# a_52_n212# a_n52_n168# w_n530_n298# pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X5 a_356_68# a_256_24# a_152_68# w_n530_n298# pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X6 a_n52_n168# a_n152_n212# a_n256_n168# w_n530_n298# pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X7 a_n256_68# a_n356_24# a_n444_68# w_n530_n298# pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
.ends

.subckt INV_2 VDD VSS IN OUT
Xnmos_3p3_6FEA4B_0 VSS IN IN VSS OUT VSS OUT IN IN VSS nmos_3p3_6FEA4B
Xpmos_3p3_KYEELV_0 OUT VDD OUT VDD IN OUT VDD VDD IN OUT IN IN VDD IN VDD IN IN VDD
+ IN pmos_3p3_KYEELV
.ends

.subckt inv_my_mag VSS IN OUT w_n60_831#
Xpmos_3p3_MQGBLR_0 IN w_n60_831# OUT w_n60_831# pmos_3p3_MQGBLR
Xnmos_3p3_DDNVWA_0 VSS OUT IN VSS nmos_3p3_DDNVWA
.ends

.subckt inv VDD VSS IN OUT
Xpmos_3p3_MQGBLR_0 IN VDD OUT VDD pmos_3p3_MQGBLR
Xnmos_3p3_DDNVWA_0 VSS OUT IN VSS nmos_3p3_DDNVWA
.ends

.subckt DFF_ D VSS RST CLK Q QB nand2_4/IN2 VDD
Xnand2_6 Q nand2_7/IN1 QB VSS VDD nand2
Xnand2_7 D nand2_7/IN1 nand2_7/OUT VSS VDD nand2
Xinv_0 VDD VSS inv_0/IN inv_0/OUT inv
Xnand2_0 CLK RST nand2_5/IN2 VSS VDD nand2
Xnand2_1 inv_0/OUT nand2_5/IN2 nand2_4/IN2 VSS VDD nand2
Xnand2_2 nand2_4/IN2 nand2_7/OUT nand2_3/IN2 VSS VDD nand2
Xnand2_3 nand2_3/IN2 RST inv_0/IN VSS VDD nand2
Xnand2_4 nand2_4/IN2 QB Q VSS VDD nand2
Xnand2_5 nand2_5/IN2 inv_0/IN nand2_7/IN1 VSS VDD nand2
.ends

.subckt nmos_3p3_5GGST2 a_n52_n50# a_n212_n50# a_52_n94# a_108_n50# a_n356_n50# a_268_n50#
+ a_n108_n94# a_n268_n94# a_212_n94# VSUBS
X0 a_108_n50# a_52_n94# a_n52_n50# VSUBS nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X1 a_268_n50# a_212_n94# a_108_n50# VSUBS nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X2 a_n52_n50# a_n108_n94# a_n212_n50# VSUBS nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X3 a_n212_n50# a_n268_n94# a_n356_n50# VSUBS nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
.ends

.subckt pmos_3p3_MWXUAR a_212_n144# a_268_n100# a_n268_n144# a_n356_n100# a_n52_n100#
+ a_n212_n100# w_n442_n230# a_108_n100# a_52_n144# a_n108_n144#
X0 a_n52_n100# a_n108_n144# a_n212_n100# w_n442_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_n212_n100# a_n268_n144# a_n356_n100# w_n442_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X2 a_108_n100# a_52_n144# a_n52_n100# w_n442_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X3 a_268_n100# a_212_n144# a_108_n100# w_n442_n230# pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
.ends

.subckt buffer_loading_mag VDD VSS OUT IN
Xnmos_3p3_5GGST2_0 VSS a_876_227# IN a_876_227# VSS VSS IN IN IN VSS nmos_3p3_5GGST2
Xpmos_3p3_MWXUAR_0 IN VDD IN VDD VDD a_876_227# VDD a_876_227# IN IN pmos_3p3_MWXUAR
X0 OUT a_876_227# VDD VDD pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 OUT a_876_227# VSS VSS nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X2 OUT a_876_227# VDD VDD pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X3 VSS a_876_227# OUT VSS nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X4 VDD a_876_227# OUT VDD pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X5 OUT a_876_227# VSS VSS nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X6 VSS a_876_227# OUT VSS nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X7 VDD a_876_227# OUT VDD pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
.ends

.subckt nmos_3p3_EA23U2 a_122_n100# a_n52_n100# a_n122_n144# a_296_n100# a_n226_n100#
+ a_n296_n144# a_n384_n100# a_52_n144# a_226_n144# VSUBS
X0 a_296_n100# a_226_n144# a_122_n100# VSUBS nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.35u
X1 a_n226_n100# a_n296_n144# a_n384_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.35u
X2 a_n52_n100# a_n122_n144# a_n226_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.35u
X3 a_122_n100# a_52_n144# a_n52_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.35u
.ends

.subckt pmos_3p3_M6H3WS a_n52_n50# a_n384_n50# a_296_n50# a_226_n94# a_n296_n94# w_n470_n180#
+ a_52_n94# a_n226_n50# a_122_n50# a_n122_n94#
X0 a_n52_n50# a_n122_n94# a_n226_n50# w_n470_n180# pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.35u
X1 a_122_n50# a_52_n94# a_n52_n50# w_n470_n180# pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.35u
X2 a_296_n50# a_226_n94# a_122_n50# w_n470_n180# pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.35u
X3 a_n226_n50# a_n296_n94# a_n384_n50# w_n470_n180# pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.35u
.ends

.subckt gf_inv_mag VDD VSS OUT IN
Xnmos_3p3_EA23U2_0 OUT VSS IN VSS OUT IN VSS IN IN VSS nmos_3p3_EA23U2
Xpmos_3p3_M6H3WS_0 VDD VDD VDD IN IN VDD IN OUT OUT IN pmos_3p3_M6H3WS
.ends

.subckt buffer_mag VDD OUT IN VSS
Xgf_inv_mag_0 VDD VSS gf_inv_mag_1/IN IN gf_inv_mag
Xgf_inv_mag_1 VDD VSS OUT gf_inv_mag_1/IN gf_inv_mag
.ends

.subckt PFD_layout PD PU VDIV VREF VDD VSS
Xinv_my_mag_0 VSS VREF DFF__1/CLK VDD inv_my_mag
Xinv_my_mag_1 VSS VDIV DFF__0/CLK VDD inv_my_mag
XDFF__0 VDD VSS DFF__1/RST DFF__0/CLK DFF__0/Q DFF__0/QB DFF__0/nand2_4/IN2 VDD DFF_
XDFF__1 VDD VSS DFF__1/RST DFF__1/CLK DFF__1/Q DFF__1/QB DFF__1/nand2_4/IN2 VDD DFF_
Xbuffer_loading_mag_0 VDD VSS PU DFF__1/Q buffer_loading_mag
Xbuffer_loading_mag_1 VDD VSS PD DFF__0/Q buffer_loading_mag
Xbuffer_mag_0 VDD DFF__1/RST nand2_0/OUT VSS buffer_mag
Xnand2_0 DFF__0/Q DFF__1/Q nand2_0/OUT VSS VDD nand2
.ends

.subckt mim_2p0fF_WS3THJ m4_n4490_n4370# m4_n4370_n4250#
X0 m4_n4370_n4250# m4_n4490_n4370# cap_mim_2f0_m4m5_noshield c_width=42.5u c_length=42.5u
.ends

.subckt cap3p_layout Pp Nn
Xmim_2p0fF_WS3THJ_0 Nn Pp mim_2p0fF_WS3THJ
.ends

.subckt ppolyf_u_3D7VPB a_1000_n1102# a_280_1000# a_n440_1000# a_n920_n1102# a_n440_n1102#
+ a_520_n1102# a_40_1000# a_n200_1000# a_n1160_1000# a_n200_n1102# a_n1160_n1102#
+ a_1000_1000# a_760_1000# a_n680_n1102# a_n920_1000# w_n1376_n1318# a_760_n1102#
+ a_520_1000# a_280_n1102# a_n680_1000# a_40_n1102#
X0 a_n680_1000# a_n680_n1102# w_n1376_n1318# ppolyf_u r_width=0.8u r_length=10u
X1 a_n920_1000# a_n920_n1102# w_n1376_n1318# ppolyf_u r_width=0.8u r_length=10u
X2 a_280_1000# a_280_n1102# w_n1376_n1318# ppolyf_u r_width=0.8u r_length=10u
X3 a_520_1000# a_520_n1102# w_n1376_n1318# ppolyf_u r_width=0.8u r_length=10u
X4 a_40_1000# a_40_n1102# w_n1376_n1318# ppolyf_u r_width=0.8u r_length=10u
X5 a_n1160_1000# a_n1160_n1102# w_n1376_n1318# ppolyf_u r_width=0.8u r_length=10u
X6 a_760_1000# a_760_n1102# w_n1376_n1318# ppolyf_u r_width=0.8u r_length=10u
X7 a_1000_1000# a_1000_n1102# w_n1376_n1318# ppolyf_u r_width=0.8u r_length=10u
X8 a_n200_1000# a_n200_n1102# w_n1376_n1318# ppolyf_u r_width=0.8u r_length=10u
X9 a_n440_1000# a_n440_n1102# w_n1376_n1318# ppolyf_u r_width=0.8u r_length=10u
.ends

.subckt res_48k_mag VDD B A
Xppolyf_u_3D7VPB_0 m1_n2577_205# m1_n3297_2306# m1_n3777_2306# m1_n4497_204# m1_n4017_204#
+ m1_n3057_204# m1_n3297_2306# m1_n3777_2306# A m1_n3537_204# m1_n4497_204# B m1_n2817_2306#
+ m1_n4017_204# m1_n4257_2306# VDD m1_n2577_205# m1_n2817_2306# m1_n3057_204# m1_n4257_2306#
+ m1_n3537_204# ppolyf_u_3D7VPB
.ends

.subckt mim_2p0fF_Q67PCK m4_5681_n21380# m4_11295_n21380# m4_n16775_n21380# m4_n22389_n21380#
+ m4_n11041_n21260# m4_17029_n21260# m4_5801_n21260# m4_11415_n21260# m4_67_n21380#
+ m4_n16655_n21260# m4_187_n21260# m4_n5547_n21380# m4_n22269_n21260# m4_16909_n21380#
+ m4_n11161_n21380# m4_n5427_n21260#
X0 m4_11415_n21260# m4_11295_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X1 m4_n22269_n21260# m4_n22389_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X2 m4_n11041_n21260# m4_n11161_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X3 m4_n5427_n21260# m4_n5547_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X4 m4_17029_n21260# m4_16909_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X5 m4_187_n21260# m4_67_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X6 m4_187_n21260# m4_67_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X7 m4_11415_n21260# m4_11295_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X8 m4_17029_n21260# m4_16909_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X9 m4_n11041_n21260# m4_n11161_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X10 m4_5801_n21260# m4_5681_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X11 m4_5801_n21260# m4_5681_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X12 m4_n22269_n21260# m4_n22389_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X13 m4_n16655_n21260# m4_n16775_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X14 m4_187_n21260# m4_67_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X15 m4_5801_n21260# m4_5681_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X16 m4_17029_n21260# m4_16909_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X17 m4_n22269_n21260# m4_n22389_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X18 m4_n5427_n21260# m4_n5547_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X19 m4_n11041_n21260# m4_n11161_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X20 m4_11415_n21260# m4_11295_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X21 m4_5801_n21260# m4_5681_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X22 m4_n16655_n21260# m4_n16775_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X23 m4_11415_n21260# m4_11295_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X24 m4_17029_n21260# m4_16909_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X25 m4_n5427_n21260# m4_n5547_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X26 m4_n16655_n21260# m4_n16775_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X27 m4_n16655_n21260# m4_n16775_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X28 m4_11415_n21260# m4_11295_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X29 m4_187_n21260# m4_67_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X30 m4_n22269_n21260# m4_n22389_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X31 m4_n11041_n21260# m4_n11161_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X32 m4_187_n21260# m4_67_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X33 m4_n22269_n21260# m4_n22389_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X34 m4_n16655_n21260# m4_n16775_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X35 m4_187_n21260# m4_67_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X36 m4_n11041_n21260# m4_n11161_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X37 m4_n22269_n21260# m4_n22389_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X38 m4_n11041_n21260# m4_n11161_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X39 m4_187_n21260# m4_67_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X40 m4_5801_n21260# m4_5681_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X41 m4_n11041_n21260# m4_n11161_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X42 m4_n5427_n21260# m4_n5547_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X43 m4_n22269_n21260# m4_n22389_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X44 m4_5801_n21260# m4_5681_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X45 m4_n16655_n21260# m4_n16775_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X46 m4_n22269_n21260# m4_n22389_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X47 m4_n5427_n21260# m4_n5547_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X48 m4_17029_n21260# m4_16909_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X49 m4_11415_n21260# m4_11295_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X50 m4_11415_n21260# m4_11295_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X51 m4_n5427_n21260# m4_n5547_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X52 m4_11415_n21260# m4_11295_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X53 m4_5801_n21260# m4_5681_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X54 m4_17029_n21260# m4_16909_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X55 m4_n11041_n21260# m4_n11161_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X56 m4_187_n21260# m4_67_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X57 m4_n16655_n21260# m4_n16775_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X58 m4_n5427_n21260# m4_n5547_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X59 m4_n5427_n21260# m4_n5547_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X60 m4_5801_n21260# m4_5681_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X61 m4_17029_n21260# m4_16909_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X62 m4_17029_n21260# m4_16909_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X63 m4_n16655_n21260# m4_n16775_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
.ends

.subckt cap80p_mag P N
Xmim_2p0fF_Q67PCK_0 N N N N P P P P N P P N P N N P mim_2p0fF_Q67PCK
.ends

.subckt LF_mag VDD VSS VCNTL
Xcap3p_layout_0 VCNTL VSS cap3p_layout
Xres_48k_mag_0 VDD cap80p_mag_0/P VCNTL res_48k_mag
Xcap80p_mag_0 cap80p_mag_0/P VSS cap80p_mag
.ends

.subckt nmos_3p3_GYTGVN a_n260_n36# a_168_n28# a_56_n72# a_n168_n72# a_n56_n28# VSUBS
X0 a_n56_n28# a_n168_n72# a_n260_n36# VSUBS nfet_03v3 ad=92.799995f pd=0.92u as=0.1576p ps=1.64u w=0.28u l=0.56u
X1 a_168_n28# a_56_n72# a_n56_n28# VSUBS nfet_03v3 ad=0.1576p pd=1.64u as=92.799995f ps=0.92u w=0.28u l=0.56u
.ends

.subckt pmos_3p3_HVHFD7 a_n52_n50# w_n338_n180# a_52_n94# a_164_n50# a_n252_n50# a_n164_n94#
X0 a_164_n50# a_52_n94# a_n52_n50# w_n338_n180# pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.56u
X1 a_n52_n50# a_n164_n94# a_n252_n50# w_n338_n180# pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.56u
.ends

.subckt CP_mag VSS VCNTL PU PD IPD_ IPD+ inv_0/VDD
Xnmos_3p3_GYTGVN_0 m1_1391_990# m1_1391_990# PD PD VCNTL VSS nmos_3p3_GYTGVN
Xnmos_3p3_GYTGVN_1 VSS VSS IPD+ IPD+ IPD+ VSS nmos_3p3_GYTGVN
Xnmos_3p3_GYTGVN_2 VSS VSS IPD+ IPD+ m1_1391_990# VSS nmos_3p3_GYTGVN
Xpmos_3p3_HVHFD7_0 m1_1376_1265# inv_0/VDD IPD_ inv_0/VDD inv_0/VDD IPD_ pmos_3p3_HVHFD7
Xpmos_3p3_HVHFD7_1 VCNTL inv_0/VDD inv_0/OUT m1_1376_1265# m1_1376_1265# inv_0/OUT
+ pmos_3p3_HVHFD7
Xpmos_3p3_HVHFD7_2 IPD_ inv_0/VDD IPD_ inv_0/VDD inv_0/VDD IPD_ pmos_3p3_HVHFD7
Xinv_0 inv_0/VDD VSS PU inv_0/OUT inv
.ends

.subckt pre_div_mag OPA1 Vdiv VDD RST CLK OPA0 VSS
Xmux_4x1_0 mux_4x1_0/I0 mux_4x1_0/I1 mux_4x1_0/I2 mux_4x1_0/I3 OPA1 OPA0 Vdiv VSS
+ mux_4x1_0/mux_2x1_1/I0 VDD mux_4x1
Xdec_2x4_ibr_mag_0 OPA0 OPA1 dec_2x4_ibr_mag_0/D0 CLK_div_2_mag_0/VDD CLK_div_3_mag_0/VDD
+ CLK_div_4_mag_0/VDD VSS VDD dec_2x4_ibr_mag
XCLK_div_4_mag_0 mux_4x1_0/I3 VSS RST CLK CLK_div_4_mag_0/CLK_div_2_mag_0/JK_FF_mag_0/nand3_mag_2/OUT
+ CLK_div_4_mag_0/CLK_div_2_mag_1/JK_FF_mag_0/nand3_mag_1/OUT CLK_div_4_mag_0/CLK_div_2_mag_1/JK_FF_mag_0/nand3_mag_2/OUT
+ CLK_div_4_mag_0/CLK_div_2_mag_0/JK_FF_mag_0/nand3_mag_0/OUT CLK_div_4_mag_0/VDD
+ CLK_div_4_mag_0/CLK_div_2_mag_0/JK_FF_mag_0/nand3_mag_1/OUT CLK_div_4_mag_0/CLK_div_2_mag_1/JK_FF_mag_0/nand3_mag_0/OUT
+ CLK_div_4_mag
XCLK_div_3_mag_0 CLK_div_3_mag_0/Q1 CLK_div_3_mag_0/Q0 mux_4x1_0/I2 CLK_div_3_mag_0/JK_FF_mag_1/nand3_mag_0/OUT
+ CLK_div_3_mag_0/JK_FF_mag_0/nand3_mag_0/OUT CLK_div_3_mag_0/JK_FF_mag_1/nand3_mag_1/OUT
+ CLK_div_3_mag_0/JK_FF_mag_0/nand3_mag_1/OUT CLK_div_3_mag_0/JK_FF_mag_1/nand3_mag_2/OUT
+ VSS CLK RST CLK_div_3_mag_0/JK_FF_mag_0/nand3_mag_2/OUT CLK_div_3_mag_0/VDD CLK_div_3_mag
XCLK_div_2_mag_0 mux_4x1_0/I1 CLK CLK_div_2_mag_0/JK_FF_mag_0/nand3_mag_0/OUT CLK_div_2_mag_0/JK_FF_mag_0/nand3_mag_1/OUT
+ VSS RST CLK_div_2_mag_0/JK_FF_mag_0/nand3_mag_2/OUT CLK_div_2_mag_0/VDD CLK_div_2_mag
XBuffer_delayed_mag_0 CLK mux_4x1_0/I0 dec_2x4_ibr_mag_0/D0 VSS Buffer_delayed_mag
.ends

.subckt pmos_3p3_YMKZL5 a_n138_n84# a_50_n84# a_n50_n128# w_n224_n214#
X0 a_50_n84# a_n50_n128# a_n138_n84# w_n224_n214# pfet_03v3 ad=0.3696p pd=2.56u as=0.3696p ps=2.56u w=0.84u l=0.5u
.ends

.subckt nmos_3p3_UKFAHE a_n138_n84# a_50_n84# a_n50_n128# VSUBS
X0 a_50_n84# a_n50_n128# a_n138_n84# VSUBS nfet_03v3 ad=0.3696p pd=2.56u as=0.3696p ps=2.56u w=0.84u l=0.5u
.ends

.subckt Tr_Gate VSS OUT IN CLK VDD
Xpmos_3p3_YMKZL5_0 OUT IN a_174_n81# VDD pmos_3p3_YMKZL5
Xpmos_3p3_YMKZL5_1 IN OUT a_174_n81# VDD pmos_3p3_YMKZL5
Xpmos_3p3_YMKZL5_2 OUT IN a_174_n81# VDD pmos_3p3_YMKZL5
Xpmos_3p3_YMKZL5_3 IN OUT a_174_n81# VDD pmos_3p3_YMKZL5
Xpmos_3p3_YMKZL5_4 a_174_n81# VDD CLK VDD pmos_3p3_YMKZL5
Xpmos_3p3_YMKZL5_5 VDD a_174_n81# CLK VDD pmos_3p3_YMKZL5
Xnmos_3p3_UKFAHE_0 OUT IN CLK VSS nmos_3p3_UKFAHE
Xpmos_3p3_YMKZL5_6 a_174_n81# VDD CLK VDD pmos_3p3_YMKZL5
Xnmos_3p3_UKFAHE_1 IN OUT CLK VSS nmos_3p3_UKFAHE
Xpmos_3p3_YMKZL5_7 VDD a_174_n81# CLK VDD pmos_3p3_YMKZL5
Xnmos_3p3_UKFAHE_2 OUT IN CLK VSS nmos_3p3_UKFAHE
Xnmos_3p3_UKFAHE_3 OUT IN CLK VSS nmos_3p3_UKFAHE
Xnmos_3p3_UKFAHE_5 a_174_n81# VSS CLK VSS nmos_3p3_UKFAHE
Xnmos_3p3_UKFAHE_4 VSS a_174_n81# CLK VSS nmos_3p3_UKFAHE
.ends

.subckt A_MUX_mag SEL IN1 IN2 VSS OUT VDD
XINV_2_0 VDD VSS SEL INV_2_0/OUT INV_2
XTr_Gate_0 VSS OUT IN2 SEL VDD Tr_Gate
XTr_Gate_1 VSS OUT IN1 INV_2_0/OUT VDD Tr_Gate
.ends

.subckt nmos_3p3_9MTZEK a_n52_n70# a_52_n114# a_n122_n114# a_n210_n70# a_122_n70#
+ VSUBS
X0 a_n52_n70# a_n122_n114# a_n210_n70# VSUBS nfet_03v3 ad=0.182p pd=1.22u as=0.308p ps=2.28u w=0.7u l=0.35u
X1 a_122_n70# a_52_n114# a_n52_n70# VSUBS nfet_03v3 ad=0.308p pd=2.28u as=0.182p ps=1.22u w=0.7u l=0.35u
.ends

.subckt pmos_3p3_585UPK a_52_n184# a_122_n140# a_n52_n140# a_n122_n184# a_n210_n140#
+ w_n296_n270#
X0 a_122_n140# a_52_n184# a_n52_n140# w_n296_n270# pfet_03v3 ad=0.616p pd=3.68u as=0.364p ps=1.92u w=1.4u l=0.35u
X1 a_n52_n140# a_n122_n184# a_n210_n140# w_n296_n270# pfet_03v3 ad=0.364p pd=1.92u as=0.616p ps=3.68u w=1.4u l=0.35u
.ends

.subckt GF_INV4 VDD IN OUT VSS
Xnmos_3p3_9MTZEK_0 OUT IN IN VSS VSS VSS nmos_3p3_9MTZEK
Xpmos_3p3_585UPK_0 IN VDD OUT IN VDD VDD pmos_3p3_585UPK
.ends

.subckt pmos_3p3_ZB3RD7 a_268_n144# a_n52_n100# a_n468_n100# a_164_n100# a_380_n100#
+ a_n164_n144# a_n380_n144# a_52_n144# a_n268_n100# w_n554_n230#
X0 a_n268_n100# a_n380_n144# a_n468_n100# w_n554_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X1 a_380_n100# a_268_n144# a_164_n100# w_n554_n230# pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X2 a_164_n100# a_52_n144# a_n52_n100# w_n554_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X3 a_n52_n100# a_n164_n144# a_n268_n100# w_n554_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
.ends

.subckt nmos_3p3_FSHHD6 a_n52_n100# a_164_n100# a_n164_n144# a_n252_n100# a_52_n144#
+ VSUBS
X0 a_164_n100# a_52_n144# a_n52_n100# VSUBS nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X1 a_n52_n100# a_n164_n144# a_n252_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
.ends

.subckt nmos_3p3_VMHHD6 a_268_n144# a_n52_n100# a_n468_n100# a_164_n100# a_380_n100#
+ a_n164_n144# a_n380_n144# a_52_n144# a_n268_n100# VSUBS
X0 a_n268_n100# a_n380_n144# a_n468_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X1 a_380_n100# a_268_n144# a_164_n100# VSUBS nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X2 a_164_n100# a_52_n144# a_n52_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X3 a_n52_n100# a_n164_n144# a_n268_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
.ends

.subckt nmos_3p3_QNHHD6 a_56_n100# a_n56_n144# a_n144_n100# VSUBS
X0 a_56_n100# a_n56_n144# a_n144_n100# VSUBS nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.56u
.ends

.subckt Delay_Cell_mag OUT OUTB EN VCONT INB IN VSS VDD
Xpmos_3p3_ZB3RD7_5 OUT VDD VDD OUTB VDD OUT OUT OUT OUTB VDD pmos_3p3_ZB3RD7
Xpmos_3p3_ZB3RD7_4 OUTB VDD VDD OUT VDD OUTB OUTB OUTB OUT VDD pmos_3p3_ZB3RD7
Xnmos_3p3_FSHHD6_0 a_562_n2079# VSS EN VSS EN VSS nmos_3p3_FSHHD6
Xnmos_3p3_VMHHD6_0 VCONT VSS VSS a_2095_n808# VSS VCONT VCONT VCONT a_2095_n808# VSS
+ nmos_3p3_VMHHD6
Xnmos_3p3_VMHHD6_2 INB a_562_n2079# a_562_n2079# OUTB a_562_n2079# INB INB INB OUTB
+ VSS nmos_3p3_VMHHD6
Xnmos_3p3_VMHHD6_1 IN a_562_n2079# a_562_n2079# OUT a_562_n2079# IN IN IN OUT VSS
+ nmos_3p3_VMHHD6
Xnmos_3p3_QNHHD6_0 a_562_n2079# a_562_n2079# a_562_n2079# VSS nmos_3p3_QNHHD6
Xnmos_3p3_QNHHD6_1 a_562_n2079# a_562_n2079# a_562_n2079# VSS nmos_3p3_QNHHD6
Xpmos_3p3_ZB3RD7_0 a_2095_n808# VDD VDD a_2095_n808# VDD a_2095_n808# a_2095_n808#
+ a_2095_n808# a_2095_n808# VDD pmos_3p3_ZB3RD7
Xpmos_3p3_ZB3RD7_1 OUT m1_277_n67# m1_277_n67# OUT m1_277_n67# OUT OUT OUT OUT VDD
+ pmos_3p3_ZB3RD7
Xpmos_3p3_ZB3RD7_2 OUTB m1_277_n67# m1_277_n67# OUTB m1_277_n67# OUTB OUTB OUTB OUTB
+ VDD pmos_3p3_ZB3RD7
Xpmos_3p3_ZB3RD7_3 a_2095_n808# m1_277_n67# m1_277_n67# VDD m1_277_n67# a_2095_n808#
+ a_2095_n808# a_2095_n808# VDD VDD pmos_3p3_ZB3RD7
.ends

.subckt nmos_3p3_AQSZEK a_n123_n70# a_35_n70# a_n35_n114# VSUBS
X0 a_35_n70# a_n35_n114# a_n123_n70# VSUBS nfet_03v3 ad=0.308p pd=2.28u as=0.308p ps=2.28u w=0.7u l=0.35u
.ends

.subckt pmos_3p3_HBGRPK w_n213_n166# a_35_n35# a_n35_n79# a_n127_n36#
X0 a_35_n35# a_n35_n79# a_n127_n36# w_n213_n166# pfet_03v3 ad=0.1646p pd=1.64u as=0.1646p ps=1.64u w=0.35u l=0.35u
.ends

.subckt GF_INV1 VDD IN OUT VSS
Xnmos_3p3_AQSZEK_0 VSS OUT IN VSS nmos_3p3_AQSZEK
Xpmos_3p3_HBGRPK_0 VDD OUT IN VDD pmos_3p3_HBGRPK
.ends

.subckt pmos_3p3_MD4UPK a_52_n324# a_226_n324# a_122_n280# a_n52_n280# a_296_n280#
+ w_n470_n410# a_n226_n280# a_n384_n280# a_n122_n324# a_n296_n324#
X0 a_296_n280# a_226_n324# a_122_n280# w_n470_n410# pfet_03v3 ad=1.232p pd=6.48u as=0.728p ps=3.32u w=2.8u l=0.35u
X1 a_n226_n280# a_n296_n324# a_n384_n280# w_n470_n410# pfet_03v3 ad=0.728p pd=3.32u as=1.232p ps=6.48u w=2.8u l=0.35u
X2 a_122_n280# a_52_n324# a_n52_n280# w_n470_n410# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.35u
X3 a_n52_n280# a_n122_n324# a_n226_n280# w_n470_n410# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.35u
.ends

.subckt nmos_3p3_S7UZWU a_52_n184# a_226_n184# a_122_n140# a_n52_n140# a_n122_n184#
+ a_296_n140# a_n226_n140# a_n296_n184# a_n384_n140# VSUBS
X0 a_n226_n140# a_n296_n184# a_n384_n140# VSUBS nfet_03v3 ad=0.364p pd=1.92u as=0.616p ps=3.68u w=1.4u l=0.35u
X1 a_122_n140# a_52_n184# a_n52_n140# VSUBS nfet_03v3 ad=0.364p pd=1.92u as=0.364p ps=1.92u w=1.4u l=0.35u
X2 a_n52_n140# a_n122_n184# a_n226_n140# VSUBS nfet_03v3 ad=0.364p pd=1.92u as=0.364p ps=1.92u w=1.4u l=0.35u
X3 a_296_n140# a_226_n184# a_122_n140# VSUBS nfet_03v3 ad=0.616p pd=3.68u as=0.364p ps=1.92u w=1.4u l=0.35u
.ends

.subckt GF_INV16 VDD IN OUT VSS
Xpmos_3p3_MD4UPK_0 IN IN OUT VDD VDD VDD OUT VDD IN IN pmos_3p3_MD4UPK
Xnmos_3p3_S7UZWU_0 IN IN OUT VSS IN VSS OUT IN VSS VSS nmos_3p3_S7UZWU
.ends

.subckt pmos_3p3_HDJZPK a_n52_n50# a_n384_n50# a_296_n50# a_226_n94# a_n296_n94# w_n470_n180#
+ a_52_n94# a_n226_n50# a_122_n50# a_n122_n94#
X0 a_n52_n50# a_n122_n94# a_n226_n50# w_n470_n180# pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.35u
X1 a_122_n50# a_52_n94# a_n52_n50# w_n470_n180# pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.35u
X2 a_296_n50# a_226_n94# a_122_n50# w_n470_n180# pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.35u
X3 a_n226_n50# a_n296_n94# a_n384_n50# w_n470_n180# pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.35u
.ends

.subckt nmos_3p3_VDSZE6 a_122_n100# a_n52_n100# a_n122_n144# a_296_n100# a_n226_n100#
+ a_n296_n144# a_n384_n100# a_52_n144# a_226_n144# VSUBS
X0 a_296_n100# a_226_n144# a_122_n100# VSUBS nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.35u
X1 a_n226_n100# a_n296_n144# a_n384_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.35u
X2 a_n52_n100# a_n122_n144# a_n226_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.35u
X3 a_122_n100# a_52_n144# a_n52_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.35u
.ends

.subckt Stage_INV IN OUT VDD VSS
Xpmos_3p3_HDJZPK_0 VDD VDD VDD IN IN VDD IN OUT OUT IN pmos_3p3_HDJZPK
Xnmos_3p3_VDSZE6_0 OUT VSS IN VSS OUT IN VSS IN IN VSS nmos_3p3_VDSZE6
.ends

.subckt VCO_mag VCONT OUT OUTB VDD EN VSS
XGF_INV4_0 VDD GF_INV4_0/IN GF_INV4_0/OUT VSS GF_INV4
XGF_INV4_1 VDD GF_INV4_1/IN GF_INV4_1/OUT VSS GF_INV4
XDelay_Cell_mag_0 Delay_Cell_mag_3/INB Delay_Cell_mag_3/IN EN VCONT Stage_INV_0/OUT
+ Stage_INV_1/OUT VSS VDD Delay_Cell_mag
XGF_INV1_1 VDD GF_INV1_1/IN GF_INV4_1/IN VSS GF_INV1
XGF_INV1_0 VDD GF_INV1_0/IN GF_INV4_0/IN VSS GF_INV1
XDelay_Cell_mag_1 Delay_Cell_mag_2/INB Delay_Cell_mag_2/IN EN VCONT GF_INV1_0/IN GF_INV1_1/IN
+ VSS VDD Delay_Cell_mag
XGF_INV16_2 VDD GF_INV4_0/OUT OUT VSS GF_INV16
XGF_INV16_1 VDD GF_INV4_1/OUT OUTB VSS GF_INV16
XStage_INV_0 Stage_INV_0/IN Stage_INV_0/OUT VDD VSS Stage_INV
XDelay_Cell_mag_2 Stage_INV_0/IN Stage_INV_1/IN EN VCONT Delay_Cell_mag_2/INB Delay_Cell_mag_2/IN
+ VSS VDD Delay_Cell_mag
XDelay_Cell_mag_3 GF_INV1_0/IN GF_INV1_1/IN EN VCONT Delay_Cell_mag_3/INB Delay_Cell_mag_3/IN
+ VSS VDD Delay_Cell_mag
XStage_INV_1 Stage_INV_1/IN Stage_INV_1/OUT VDD VSS Stage_INV
.ends

.subckt pmos_3p3_Q354KU a_212_n144# a_268_n100# a_n692_n100# a_n268_n144# a_372_n144#
+ a_428_n100# a_n52_n100# a_n428_n144# a_532_n144# a_588_n100# w_n922_n230# a_n212_n100#
+ a_n588_n144# a_692_n144# a_748_n100# a_n372_n100# a_n748_n144# a_108_n100# a_52_n144#
+ a_n836_n100# a_n532_n100# a_n108_n144#
X0 a_n52_n100# a_n108_n144# a_n212_n100# w_n922_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_588_n100# a_532_n144# a_428_n100# w_n922_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X2 a_n212_n100# a_n268_n144# a_n372_n100# w_n922_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X3 a_n692_n100# a_n748_n144# a_n836_n100# w_n922_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X4 a_748_n100# a_692_n144# a_588_n100# w_n922_n230# pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X5 a_108_n100# a_52_n144# a_n52_n100# w_n922_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X6 a_268_n100# a_212_n144# a_108_n100# w_n922_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X7 a_n372_n100# a_n428_n144# a_n532_n100# w_n922_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X8 a_428_n100# a_372_n144# a_268_n100# w_n922_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X9 a_n532_n100# a_n588_n144# a_n692_n100# w_n922_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
.ends

.subckt nmos_3p3_W9BEG7 a_212_n144# a_268_n100# a_n692_n100# a_n268_n144# a_372_n144#
+ a_428_n100# a_n52_n100# a_n428_n144# a_532_n144# a_588_n100# a_n212_n100# a_n588_n144#
+ a_692_n144# a_748_n100# a_n372_n100# a_n748_n144# a_108_n100# a_52_n144# a_n836_n100#
+ a_n532_n100# a_n108_n144# VSUBS
X0 a_n52_n100# a_n108_n144# a_n212_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_588_n100# a_532_n144# a_428_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X2 a_n212_n100# a_n268_n144# a_n372_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X3 a_n692_n100# a_n748_n144# a_n836_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X4 a_748_n100# a_692_n144# a_588_n100# VSUBS nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X5 a_108_n100# a_52_n144# a_n52_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X6 a_268_n100# a_212_n144# a_108_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X7 a_n372_n100# a_n428_n144# a_n532_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X8 a_428_n100# a_372_n144# a_268_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X9 a_n532_n100# a_n588_n144# a_n692_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
.ends

.subckt Transmission_gate_mag CLK VDD VIN VOUT VSS
Xinv_my_mag_0 VSS CLK inv_my_mag_0/OUT VDD inv_my_mag
Xpmos_3p3_Q354KU_0 inv_my_mag_0/OUT VOUT VOUT inv_my_mag_0/OUT inv_my_mag_0/OUT VIN
+ VOUT inv_my_mag_0/OUT inv_my_mag_0/OUT VOUT VDD VIN inv_my_mag_0/OUT inv_my_mag_0/OUT
+ VIN VOUT inv_my_mag_0/OUT VIN inv_my_mag_0/OUT VIN VIN inv_my_mag_0/OUT pmos_3p3_Q354KU
Xnmos_3p3_W9BEG7_0 CLK VOUT VOUT CLK CLK VIN VOUT CLK CLK VOUT VIN CLK CLK VIN VOUT
+ CLK VIN CLK VIN VIN CLK VSS nmos_3p3_W9BEG7
.ends

.subckt a2x1mux_mag IN1 IN2 SEL VOUT VDD VSS
Xinv_my_mag_0 VSS SEL inv_my_mag_0/OUT VDD inv_my_mag
XTransmission_gate_mag_0 inv_my_mag_0/OUT VDD IN1 VOUT VSS Transmission_gate_mag
XTransmission_gate_mag_1 SEL VDD IN2 VOUT VSS Transmission_gate_mag
.ends

.subckt pll_4_mag IPD+ IPD_ VCO_op VCO_op_bar VSS Iref Output1 Output2 F2 F1 F0 T0
+ T1 LP_RES_CAP_INT Vdiv_FB_MUX_INT VCNT_MUX_INT VDD_BUFF_INT_2 INV_BUFF_INT_3 INV_BUFF_INT_2
+ INV_BUFF_INT_1 Output_2_INT Output_1_INT Test_Output_INT PRE_DIV_OP_INT PFD_Vdiv_IN_INT
+ PFD_Vref_IN_INT PU_INT PD_INT PU_MUX_OP_INT PD_MUX_OP_INT VDD_INT_8 P1 P0 Vref Vdiv_test
+ S0 S1 S2 PD_test PU_test LP_op_test LP_ext vcntl_test VDD_VCO Vo_test RST_DIV OPA0
+ OPA1 OPB0 OPB1 Test_output
XTappered_Buffer_0 VDD_BUFF_INT_2 INV_BUFF_INT_1 Output2 VSS Tappered_Buffer
XCurrent_Mirror_Top_0 VDD_INT_8 Current_Mirror_Top_0/G_source_up Current_Mirror_Top_0/G_source_dn
+ VSS Current_Mirror_Top_0/G_sink_up Current_Mirror_Top_0/G_sink_dn Current_Mirror_Top_0/SD0_1
+ Current_Mirror_Top_0/G1_2 Current_Mirror_Top_0/G1_1 Current_Mirror_Top_0/SD1_1 Current_Mirror_Top_0/G2_1
+ Current_Mirror_Top_0/SD2_1 Iref IPD_ IPD+ Current_Mirror_Top_0/A1 Current_Mirror_Top_0/A2
+ Current_Mirror_Top
XTappered_Buffer_1 VDD_BUFF_INT_2 INV_BUFF_INT_3 Test_output VSS Tappered_Buffer
XTappered_Buffer_2 VDD_BUFF_INT_2 INV_BUFF_INT_2 Output1 VSS Tappered_Buffer
Xmux_4x1_ibr_0 PU_INT PD_INT VCO_op Vdiv_FB_MUX_INT T1 T0 Test_Output_INT VSS VDD_INT_8
+ mux_4x1_ibr
XOutput_Div_Mag_0 OPA0 OPA1 Output_1_INT VDD_INT_8 RST_DIV VCO_op VSS Output_Div_Mag
XOutput_Div_Mag_1 OPB0 OPB1 Output_2_INT VDD_INT_8 RST_DIV VCO_op VSS Output_Div_Mag
XFeedback_Divider_mag_0 CLK_FB_IN_INT RST_DIV F2 F1 F0 Vdiv_FB_MUX_INT VDD_INT_8 Feedback_Divider_mag_0/Vdiv90
+ Feedback_Divider_mag_0/Vdiv96 Feedback_Divider_mag_0/Vdiv93 Feedback_Divider_mag_0/Vdiv99
+ Feedback_Divider_mag_0/Vdiv110 Feedback_Divider_mag_0/Vdiv108 Feedback_Divider_mag_0/Vdiv100
+ Feedback_Divider_mag_0/Vdiv105 Feedback_Divider_mag_0/VDD90 Feedback_Divider_mag_0/VDD99
+ Feedback_Divider_mag_0/VDD108 Feedback_Divider_mag_0/VDD100 Feedback_Divider_mag_0/VDD105
+ Feedback_Divider_mag_0/VDD93 Feedback_Divider_mag_0/VDD96 Feedback_Divider_mag_0/VDD110
+ VSS Feedback_Divider_mag
Xmux_2x1_ibr_0 S1 PD_INT PD_MUX_OP_INT PD_test VDD_INT_8 VSS mux_2x1_ibr
Xmux_2x1_ibr_1 S1 PU_INT PU_MUX_OP_INT PU_test VDD_INT_8 VSS mux_2x1_ibr
Xmux_2x1_ibr_3 S1 Vdiv_FB_MUX_INT PFD_Vdiv_IN_INT Vdiv_test VDD_INT_8 VSS mux_2x1_ibr
XINV_2_0 VDD_BUFF_INT_2 VSS Test_Output_INT INV_BUFF_INT_3 INV_2
XINV_2_2 VDD_BUFF_INT_2 VSS Output_2_INT INV_BUFF_INT_1 INV_2
XINV_2_1 VDD_BUFF_INT_2 VSS Output_1_INT INV_BUFF_INT_2 INV_2
Xmux_2x1_ibr_4 S0 PRE_DIV_OP_INT PFD_Vref_IN_INT Vref VDD_INT_8 VSS mux_2x1_ibr
XPFD_layout_0 PD_INT PU_INT PFD_Vdiv_IN_INT PFD_Vref_IN_INT VDD_INT_8 VSS PFD_layout
XLF_mag_0 VDD_INT_8 VSS LP_RES_CAP_INT LF_mag
XCP_mag_0 VSS LP_op_test PU_MUX_OP_INT PD_MUX_OP_INT IPD_ IPD+ VDD_INT_8 CP_mag
Xpre_div_mag_0 P1 PRE_DIV_OP_INT VDD_INT_8 RST_DIV Vref P0 VSS pre_div_mag
XA_MUX_mag_1 S1 Vo_test VCO_op VSS CLK_FB_IN_INT VDD_INT_8 A_MUX_mag
XVCO_mag_0 VCNT_MUX_INT VCO_op VCO_op_bar VDD_VCO VDD_INT_8 VSS VCO_mag
XA_MUX_mag_0 S1 vcntl_test LP_op_test VSS VCNT_MUX_INT VDD_INT_8 A_MUX_mag
Xa2x1mux_mag_0 LP_ext LP_RES_CAP_INT S2 LP_op_test VDD_INT_8 VSS a2x1mux_mag
.ends

