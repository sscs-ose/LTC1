magic
tech gf180mcuC
magscale 1 10
timestamp 1695206022
<< nwell >>
rect 15928 2099 16126 2153
<< psubdiff >>
rect 824 -34 1235 9
rect 824 -197 876 -34
rect 1187 -197 1235 -34
rect 824 -226 1235 -197
rect 1843 -29 2254 14
rect 1843 -192 1895 -29
rect 2206 -192 2254 -29
rect 1843 -221 2254 -192
rect 2910 -29 3321 14
rect 2910 -192 2962 -29
rect 3273 -192 3321 -29
rect 2910 -221 3321 -192
rect 4307 -22 4718 21
rect 4307 -185 4359 -22
rect 4670 -185 4718 -22
rect 4307 -214 4718 -185
rect 5960 -22 6371 21
rect 5960 -185 6012 -22
rect 6323 -185 6371 -22
rect 5960 -214 6371 -185
rect 7687 -27 8098 16
rect 7687 -190 7739 -27
rect 8050 -190 8098 -27
rect 7687 -219 8098 -190
rect 9340 -27 9751 16
rect 9340 -190 9392 -27
rect 9703 -190 9751 -27
rect 9340 -219 9751 -190
rect 11269 -27 11680 16
rect 11269 -190 11321 -27
rect 11632 -190 11680 -27
rect 11269 -219 11680 -190
rect 13198 -27 13609 16
rect 13198 -190 13250 -27
rect 13561 -190 13609 -27
rect 13198 -219 13609 -190
<< psubdiffcont >>
rect 876 -197 1187 -34
rect 1895 -192 2206 -29
rect 2962 -192 3273 -29
rect 4359 -185 4670 -22
rect 6012 -185 6323 -22
rect 7739 -190 8050 -27
rect 9392 -190 9703 -27
rect 11321 -190 11632 -27
rect 13250 -190 13561 -27
<< metal1 >>
rect 587 5156 20618 5340
rect 587 5147 18987 5156
rect 587 5132 18369 5147
rect 587 5121 17448 5132
rect 587 5101 16729 5121
rect 587 5088 15965 5101
rect 587 5014 15130 5088
rect 15236 5027 15965 5088
rect 16071 5047 16729 5101
rect 16835 5058 17448 5121
rect 17554 5073 18369 5132
rect 18475 5082 18987 5147
rect 19093 5145 20618 5156
rect 19093 5082 19678 5145
rect 18475 5073 19678 5082
rect 17554 5071 19678 5073
rect 19784 5135 20618 5145
rect 19784 5071 20077 5135
rect 17554 5058 20077 5071
rect 16835 5051 20077 5058
rect 20217 5051 20618 5135
rect 16835 5047 20618 5051
rect 16071 5027 20618 5047
rect 15236 5014 20618 5027
rect 587 5005 20618 5014
rect 6196 4538 6333 4704
rect 8927 4616 9134 5005
rect 9847 4616 10054 5005
rect 11106 4591 11337 5005
rect -502 4386 -188 4423
rect -502 4287 -451 4386
rect -321 4287 -188 4386
rect -502 4256 -188 4287
rect 12256 3186 12521 3431
rect 18187 3254 20352 3262
rect 18187 3243 18980 3254
rect 18187 3169 18371 3243
rect 18477 3180 18980 3243
rect 19086 3180 19681 3254
rect 19787 3180 20352 3254
rect 18477 3169 20352 3180
rect 18187 3082 20352 3169
rect 19948 2917 20352 3082
rect 20550 2581 20806 2632
rect 20294 2523 20806 2581
rect 20550 2502 20806 2523
rect -451 2404 -105 2441
rect -451 2288 -406 2404
rect -284 2288 -105 2404
rect 12876 2369 14508 2475
rect -451 2257 -105 2288
rect 14429 1654 14508 2369
rect 15939 2202 16098 2203
rect 14554 2199 18248 2202
rect 14554 2197 17435 2199
rect 14554 2195 15955 2197
rect 14554 2142 15132 2195
rect 15251 2142 15955 2195
rect 14554 2141 15955 2142
rect 16088 2141 16716 2197
rect 16849 2143 17435 2197
rect 17568 2143 18248 2199
rect 16849 2141 18248 2143
rect 14554 1979 18248 2141
rect 14429 1582 14695 1654
rect 14050 93 14899 357
rect 587 -22 20711 93
rect 587 -29 4359 -22
rect 587 -34 1895 -29
rect 587 -197 876 -34
rect 1187 -192 1895 -34
rect 2206 -192 2962 -29
rect 3273 -185 4359 -29
rect 4670 -185 6012 -22
rect 6323 -27 20711 -22
rect 6323 -185 7739 -27
rect 3273 -190 7739 -185
rect 8050 -190 9392 -27
rect 9703 -190 11321 -27
rect 11632 -190 13250 -27
rect 13561 -190 20711 -27
rect 3273 -192 20711 -190
rect 1187 -197 20711 -192
rect 587 -242 20711 -197
<< via1 >>
rect 15130 5014 15236 5088
rect 15965 5027 16071 5101
rect 16729 5047 16835 5121
rect 17448 5058 17554 5132
rect 18369 5073 18475 5147
rect 18987 5082 19093 5156
rect 19678 5071 19784 5145
rect 20077 5051 20217 5135
rect -451 4287 -321 4386
rect 18371 3169 18477 3243
rect 18980 3180 19086 3254
rect 19681 3180 19787 3254
rect -406 2288 -284 2404
rect 15132 2142 15251 2195
rect 15955 2141 16088 2197
rect 16716 2141 16849 2197
rect 17435 2143 17568 2199
<< metal2 >>
rect 16704 5121 16863 5148
rect 15939 5101 16098 5116
rect 15110 5088 15269 5100
rect 15110 5014 15130 5088
rect 15236 5014 15269 5088
rect -502 4411 -188 4423
rect -502 4275 -460 4411
rect -261 4275 -188 4411
rect -502 4256 -188 4275
rect -451 2410 -105 2441
rect -451 2279 -420 2410
rect -188 2279 -105 2410
rect -451 2257 -105 2279
rect 15110 2195 15269 5014
rect 15110 2142 15132 2195
rect 15251 2142 15269 2195
rect 15110 2139 15269 2142
rect 15939 5027 15965 5101
rect 16071 5027 16098 5101
rect 15939 2197 16098 5027
rect 15939 2141 15955 2197
rect 16088 2141 16098 2197
rect 15939 2129 16098 2141
rect 16704 5047 16729 5121
rect 16835 5047 16863 5121
rect 16704 2197 16863 5047
rect 16704 2141 16716 2197
rect 16849 2141 16863 2197
rect 16704 2136 16863 2141
rect 17421 5132 17580 5164
rect 17421 5058 17448 5132
rect 17554 5058 17580 5132
rect 17421 2199 17580 5058
rect 18329 5147 18536 5179
rect 18329 5073 18369 5147
rect 18475 5073 18536 5147
rect 18329 3243 18536 5073
rect 18329 3169 18371 3243
rect 18477 3169 18536 3243
rect 18934 5156 19141 5179
rect 18934 5082 18987 5156
rect 19093 5082 19141 5156
rect 18934 3254 19141 5082
rect 18934 3180 18980 3254
rect 19086 3180 19141 3254
rect 18934 3171 19141 3180
rect 19635 5145 19842 5163
rect 19635 5071 19678 5145
rect 19784 5071 19842 5145
rect 19635 3254 19842 5071
rect 19635 3180 19681 3254
rect 19787 3180 19842 3254
rect 19635 3171 19842 3180
rect 20051 5135 20258 5168
rect 20051 5051 20077 5135
rect 20217 5051 20258 5135
rect 18329 3158 18536 3169
rect 20051 3164 20258 5051
rect 17421 2143 17435 2199
rect 17568 2143 17580 2199
rect 17421 2138 17580 2143
<< via2 >>
rect -460 4386 -261 4411
rect -460 4287 -451 4386
rect -451 4287 -321 4386
rect -321 4287 -261 4386
rect -460 4275 -261 4287
rect -420 2404 -188 2410
rect -420 2288 -406 2404
rect -406 2288 -284 2404
rect -284 2288 -188 2404
rect -420 2279 -188 2288
<< metal3 >>
rect -502 4411 -188 4423
rect -502 4275 -460 4411
rect -261 4381 -188 4411
rect -261 4292 6307 4381
rect -261 4275 -188 4292
rect -502 4256 -188 4275
rect -451 2410 -105 2441
rect -451 2279 -420 2410
rect -188 2392 -105 2410
rect -188 2279 3825 2392
rect -451 2275 3825 2279
rect -451 2257 -105 2275
rect 11505 490 11562 2409
rect 11505 433 17697 490
use CLK_div_3_mag  CLK_div_3_mag_0
timestamp 1695206022
transform 1 0 14554 0 1 -4
box -34 -1 6461 3249
use CLK_div_31_mag  CLK_div_31_mag_0
timestamp 1695206022
transform 1 0 459 0 1 156
box -459 -156 13910 4667
<< labels >>
flabel metal1 8239 5167 8239 5167 0 FreeSans 960 0 0 0 VDD
port 0 nsew
flabel metal1 14374 62 14374 62 0 FreeSans 960 0 0 0 VSS
port 1 nsew
flabel metal1 20642 2582 20642 2582 0 FreeSans 960 0 0 0 Vdiv93
port 2 nsew
flabel via2 -274 2346 -274 2346 0 FreeSans 960 0 0 0 RST
port 3 nsew
flabel via2 -353 4344 -353 4344 0 FreeSans 960 0 0 0 CLK
port 4 nsew
<< end >>
