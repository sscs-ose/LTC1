magic
tech gf180mcuC
magscale 1 10
timestamp 1714492828
<< nwell >>
rect -15 429 577 545
rect -15 428 17 429
rect 540 428 577 429
rect 27 420 534 426
<< psubdiff >>
rect -32 -410 576 -391
rect -32 -463 0 -410
rect 52 -463 125 -410
rect 177 -463 250 -410
rect 302 -463 375 -410
rect 427 -463 500 -410
rect 552 -463 576 -410
rect -32 -481 576 -463
<< nsubdiff >>
rect 23 500 136 517
rect 23 454 38 500
rect 84 454 136 500
rect 23 445 136 454
rect 23 437 98 445
<< psubdiffcont >>
rect 0 -463 52 -410
rect 125 -463 177 -410
rect 250 -463 302 -410
rect 375 -463 427 -410
rect 500 -463 552 -410
<< nsubdiffcont >>
rect 38 454 84 500
<< polysilicon >>
rect 159 0 229 16
rect 79 -13 229 0
rect 333 -13 403 17
rect 79 -82 94 -13
rect 162 -82 403 -13
rect 79 -86 403 -82
rect 79 -95 229 -86
rect 159 -117 229 -95
rect 333 -116 403 -86
<< polycontact >>
rect 94 -82 162 -13
<< metal1 >>
rect -146 560 701 650
rect -146 -391 -54 560
rect 25 501 94 503
rect 25 500 135 501
rect 25 454 38 500
rect 84 454 534 500
rect 25 437 534 454
rect 27 412 534 437
rect 84 333 130 412
rect 432 334 478 412
rect 79 -13 173 0
rect 79 -22 94 -13
rect 10 -74 94 -22
rect 79 -82 94 -74
rect 162 -82 173 -13
rect 79 -95 173 -82
rect 258 -35 304 77
rect 258 -81 502 -35
rect 258 -175 304 -81
rect 84 -391 131 -263
rect 431 -391 478 -262
rect 611 -391 701 560
rect -146 -410 701 -391
rect -146 -463 0 -410
rect 52 -463 125 -410
rect 177 -463 250 -410
rect 302 -463 375 -410
rect 427 -463 500 -410
rect 552 -463 701 -410
rect -146 -481 701 -463
use nmos_3p3_9MTZEK  nmos_3p3_9MTZEK_0
timestamp 1714126980
transform 1 0 281 0 1 -229
box -234 -138 234 138
use pmos_3p3_585UPK  pmos_3p3_585UPK_0
timestamp 1714126980
transform 1 0 281 0 1 197
box -296 -270 296 270
<< labels >>
flabel metal1 25 -53 25 -53 0 FreeSans 320 0 0 0 IN
port 1 nsew
flabel metal1 452 -60 452 -60 0 FreeSans 320 0 0 0 OUT
port 2 nsew
flabel metal1 216 -425 216 -425 0 FreeSans 320 0 0 0 VSS
port 3 nsew
flabel metal1 121 455 121 455 0 FreeSans 320 0 0 0 VDD
port 0 nsew
<< end >>
