magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1073 -1289 1073 1289
<< metal1 >>
rect -73 283 73 289
rect -73 257 -67 283
rect -41 257 -13 283
rect 13 257 41 283
rect 67 257 73 283
rect -73 229 73 257
rect -73 203 -67 229
rect -41 203 -13 229
rect 13 203 41 229
rect 67 203 73 229
rect -73 175 73 203
rect -73 149 -67 175
rect -41 149 -13 175
rect 13 149 41 175
rect 67 149 73 175
rect -73 121 73 149
rect -73 95 -67 121
rect -41 95 -13 121
rect 13 95 41 121
rect 67 95 73 121
rect -73 67 73 95
rect -73 41 -67 67
rect -41 41 -13 67
rect 13 41 41 67
rect 67 41 73 67
rect -73 13 73 41
rect -73 -13 -67 13
rect -41 -13 -13 13
rect 13 -13 41 13
rect 67 -13 73 13
rect -73 -41 73 -13
rect -73 -67 -67 -41
rect -41 -67 -13 -41
rect 13 -67 41 -41
rect 67 -67 73 -41
rect -73 -95 73 -67
rect -73 -121 -67 -95
rect -41 -121 -13 -95
rect 13 -121 41 -95
rect 67 -121 73 -95
rect -73 -149 73 -121
rect -73 -175 -67 -149
rect -41 -175 -13 -149
rect 13 -175 41 -149
rect 67 -175 73 -149
rect -73 -203 73 -175
rect -73 -229 -67 -203
rect -41 -229 -13 -203
rect 13 -229 41 -203
rect 67 -229 73 -203
rect -73 -257 73 -229
rect -73 -283 -67 -257
rect -41 -283 -13 -257
rect 13 -283 41 -257
rect 67 -283 73 -257
rect -73 -289 73 -283
<< via1 >>
rect -67 257 -41 283
rect -13 257 13 283
rect 41 257 67 283
rect -67 203 -41 229
rect -13 203 13 229
rect 41 203 67 229
rect -67 149 -41 175
rect -13 149 13 175
rect 41 149 67 175
rect -67 95 -41 121
rect -13 95 13 121
rect 41 95 67 121
rect -67 41 -41 67
rect -13 41 13 67
rect 41 41 67 67
rect -67 -13 -41 13
rect -13 -13 13 13
rect 41 -13 67 13
rect -67 -67 -41 -41
rect -13 -67 13 -41
rect 41 -67 67 -41
rect -67 -121 -41 -95
rect -13 -121 13 -95
rect 41 -121 67 -95
rect -67 -175 -41 -149
rect -13 -175 13 -149
rect 41 -175 67 -149
rect -67 -229 -41 -203
rect -13 -229 13 -203
rect 41 -229 67 -203
rect -67 -283 -41 -257
rect -13 -283 13 -257
rect 41 -283 67 -257
<< metal2 >>
rect -73 283 73 289
rect -73 257 -67 283
rect -41 257 -13 283
rect 13 257 41 283
rect 67 257 73 283
rect -73 229 73 257
rect -73 203 -67 229
rect -41 203 -13 229
rect 13 203 41 229
rect 67 203 73 229
rect -73 175 73 203
rect -73 149 -67 175
rect -41 149 -13 175
rect 13 149 41 175
rect 67 149 73 175
rect -73 121 73 149
rect -73 95 -67 121
rect -41 95 -13 121
rect 13 95 41 121
rect 67 95 73 121
rect -73 67 73 95
rect -73 41 -67 67
rect -41 41 -13 67
rect 13 41 41 67
rect 67 41 73 67
rect -73 13 73 41
rect -73 -13 -67 13
rect -41 -13 -13 13
rect 13 -13 41 13
rect 67 -13 73 13
rect -73 -41 73 -13
rect -73 -67 -67 -41
rect -41 -67 -13 -41
rect 13 -67 41 -41
rect 67 -67 73 -41
rect -73 -95 73 -67
rect -73 -121 -67 -95
rect -41 -121 -13 -95
rect 13 -121 41 -95
rect 67 -121 73 -95
rect -73 -149 73 -121
rect -73 -175 -67 -149
rect -41 -175 -13 -149
rect 13 -175 41 -149
rect 67 -175 73 -149
rect -73 -203 73 -175
rect -73 -229 -67 -203
rect -41 -229 -13 -203
rect 13 -229 41 -203
rect 67 -229 73 -203
rect -73 -257 73 -229
rect -73 -283 -67 -257
rect -41 -283 -13 -257
rect 13 -283 41 -257
rect 67 -283 73 -257
rect -73 -289 73 -283
<< end >>
