magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -3037 -2045 3037 2045
<< psubdiff >>
rect -1037 23 1037 45
rect -1037 -23 -1015 23
rect -969 -23 -891 23
rect -845 -23 -767 23
rect -721 -23 -643 23
rect -597 -23 -519 23
rect -473 -23 -395 23
rect -349 -23 -271 23
rect -225 -23 -147 23
rect -101 -23 -23 23
rect 23 -23 101 23
rect 147 -23 225 23
rect 271 -23 349 23
rect 395 -23 473 23
rect 519 -23 597 23
rect 643 -23 721 23
rect 767 -23 845 23
rect 891 -23 969 23
rect 1015 -23 1037 23
rect -1037 -45 1037 -23
<< psubdiffcont >>
rect -1015 -23 -969 23
rect -891 -23 -845 23
rect -767 -23 -721 23
rect -643 -23 -597 23
rect -519 -23 -473 23
rect -395 -23 -349 23
rect -271 -23 -225 23
rect -147 -23 -101 23
rect -23 -23 23 23
rect 101 -23 147 23
rect 225 -23 271 23
rect 349 -23 395 23
rect 473 -23 519 23
rect 597 -23 643 23
rect 721 -23 767 23
rect 845 -23 891 23
rect 969 -23 1015 23
<< metal1 >>
rect -1026 23 1026 34
rect -1026 -23 -1015 23
rect -969 -23 -891 23
rect -845 -23 -767 23
rect -721 -23 -643 23
rect -597 -23 -519 23
rect -473 -23 -395 23
rect -349 -23 -271 23
rect -225 -23 -147 23
rect -101 -23 -23 23
rect 23 -23 101 23
rect 147 -23 225 23
rect 271 -23 349 23
rect 395 -23 473 23
rect 519 -23 597 23
rect 643 -23 721 23
rect 767 -23 845 23
rect 891 -23 969 23
rect 1015 -23 1026 23
rect -1026 -34 1026 -23
<< end >>
