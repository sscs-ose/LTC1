magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1236 -1205 1236 1205
<< metal1 >>
rect -236 199 236 205
rect -236 173 -230 199
rect -204 173 -168 199
rect -142 173 -106 199
rect -80 173 -44 199
rect -18 173 18 199
rect 44 173 80 199
rect 106 173 142 199
rect 168 173 204 199
rect 230 173 236 199
rect -236 137 236 173
rect -236 111 -230 137
rect -204 111 -168 137
rect -142 111 -106 137
rect -80 111 -44 137
rect -18 111 18 137
rect 44 111 80 137
rect 106 111 142 137
rect 168 111 204 137
rect 230 111 236 137
rect -236 75 236 111
rect -236 49 -230 75
rect -204 49 -168 75
rect -142 49 -106 75
rect -80 49 -44 75
rect -18 49 18 75
rect 44 49 80 75
rect 106 49 142 75
rect 168 49 204 75
rect 230 49 236 75
rect -236 13 236 49
rect -236 -13 -230 13
rect -204 -13 -168 13
rect -142 -13 -106 13
rect -80 -13 -44 13
rect -18 -13 18 13
rect 44 -13 80 13
rect 106 -13 142 13
rect 168 -13 204 13
rect 230 -13 236 13
rect -236 -49 236 -13
rect -236 -75 -230 -49
rect -204 -75 -168 -49
rect -142 -75 -106 -49
rect -80 -75 -44 -49
rect -18 -75 18 -49
rect 44 -75 80 -49
rect 106 -75 142 -49
rect 168 -75 204 -49
rect 230 -75 236 -49
rect -236 -111 236 -75
rect -236 -137 -230 -111
rect -204 -137 -168 -111
rect -142 -137 -106 -111
rect -80 -137 -44 -111
rect -18 -137 18 -111
rect 44 -137 80 -111
rect 106 -137 142 -111
rect 168 -137 204 -111
rect 230 -137 236 -111
rect -236 -173 236 -137
rect -236 -199 -230 -173
rect -204 -199 -168 -173
rect -142 -199 -106 -173
rect -80 -199 -44 -173
rect -18 -199 18 -173
rect 44 -199 80 -173
rect 106 -199 142 -173
rect 168 -199 204 -173
rect 230 -199 236 -173
rect -236 -205 236 -199
<< via1 >>
rect -230 173 -204 199
rect -168 173 -142 199
rect -106 173 -80 199
rect -44 173 -18 199
rect 18 173 44 199
rect 80 173 106 199
rect 142 173 168 199
rect 204 173 230 199
rect -230 111 -204 137
rect -168 111 -142 137
rect -106 111 -80 137
rect -44 111 -18 137
rect 18 111 44 137
rect 80 111 106 137
rect 142 111 168 137
rect 204 111 230 137
rect -230 49 -204 75
rect -168 49 -142 75
rect -106 49 -80 75
rect -44 49 -18 75
rect 18 49 44 75
rect 80 49 106 75
rect 142 49 168 75
rect 204 49 230 75
rect -230 -13 -204 13
rect -168 -13 -142 13
rect -106 -13 -80 13
rect -44 -13 -18 13
rect 18 -13 44 13
rect 80 -13 106 13
rect 142 -13 168 13
rect 204 -13 230 13
rect -230 -75 -204 -49
rect -168 -75 -142 -49
rect -106 -75 -80 -49
rect -44 -75 -18 -49
rect 18 -75 44 -49
rect 80 -75 106 -49
rect 142 -75 168 -49
rect 204 -75 230 -49
rect -230 -137 -204 -111
rect -168 -137 -142 -111
rect -106 -137 -80 -111
rect -44 -137 -18 -111
rect 18 -137 44 -111
rect 80 -137 106 -111
rect 142 -137 168 -111
rect 204 -137 230 -111
rect -230 -199 -204 -173
rect -168 -199 -142 -173
rect -106 -199 -80 -173
rect -44 -199 -18 -173
rect 18 -199 44 -173
rect 80 -199 106 -173
rect 142 -199 168 -173
rect 204 -199 230 -173
<< metal2 >>
rect -236 199 236 205
rect -236 173 -230 199
rect -204 173 -168 199
rect -142 173 -106 199
rect -80 173 -44 199
rect -18 173 18 199
rect 44 173 80 199
rect 106 173 142 199
rect 168 173 204 199
rect 230 173 236 199
rect -236 137 236 173
rect -236 111 -230 137
rect -204 111 -168 137
rect -142 111 -106 137
rect -80 111 -44 137
rect -18 111 18 137
rect 44 111 80 137
rect 106 111 142 137
rect 168 111 204 137
rect 230 111 236 137
rect -236 75 236 111
rect -236 49 -230 75
rect -204 49 -168 75
rect -142 49 -106 75
rect -80 49 -44 75
rect -18 49 18 75
rect 44 49 80 75
rect 106 49 142 75
rect 168 49 204 75
rect 230 49 236 75
rect -236 13 236 49
rect -236 -13 -230 13
rect -204 -13 -168 13
rect -142 -13 -106 13
rect -80 -13 -44 13
rect -18 -13 18 13
rect 44 -13 80 13
rect 106 -13 142 13
rect 168 -13 204 13
rect 230 -13 236 13
rect -236 -49 236 -13
rect -236 -75 -230 -49
rect -204 -75 -168 -49
rect -142 -75 -106 -49
rect -80 -75 -44 -49
rect -18 -75 18 -49
rect 44 -75 80 -49
rect 106 -75 142 -49
rect 168 -75 204 -49
rect 230 -75 236 -49
rect -236 -111 236 -75
rect -236 -137 -230 -111
rect -204 -137 -168 -111
rect -142 -137 -106 -111
rect -80 -137 -44 -111
rect -18 -137 18 -111
rect 44 -137 80 -111
rect 106 -137 142 -111
rect 168 -137 204 -111
rect 230 -137 236 -111
rect -236 -173 236 -137
rect -236 -199 -230 -173
rect -204 -199 -168 -173
rect -142 -199 -106 -173
rect -80 -199 -44 -173
rect -18 -199 18 -173
rect 44 -199 80 -173
rect 106 -199 142 -173
rect 168 -199 204 -173
rect 230 -199 236 -173
rect -236 -205 236 -199
<< end >>
