magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2045 -19811 2045 19811
<< psubdiff >>
rect -45 17789 45 17811
rect -45 -17789 -23 17789
rect 23 -17789 45 17789
rect -45 -17811 45 -17789
<< psubdiffcont >>
rect -23 -17789 23 17789
<< metal1 >>
rect -34 17789 34 17800
rect -34 -17789 -23 17789
rect 23 -17789 34 17789
rect -34 -17800 34 -17789
<< end >>
