* NGSPICE file created from and_5_mag_flat.ext - technology: gf180mcuC

.subckt and_5_mag_flat B C D E VDD VSS VOUT A
X0 VDD C.t0 and2_mag_1.GF_INV_MAG_0.IN VDD.t3 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1 and2_mag_0.GF_INV_MAG_0.IN A.t0 a_916_743# VSS.t19 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2 and2_mag_1.GF_INV_MAG_0.IN and2_mag_1.IN2 VDD.t27 VDD.t26 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X3 VOUT and2_mag_3.GF_INV_MAG_0.IN VDD.t23 VDD.t22 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X4 a_2813_727# and2_mag_2.IN2 VSS.t7 VSS.t6 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X5 VOUT and2_mag_3.GF_INV_MAG_0.IN VSS.t13 VSS.t12 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X6 VDD D.t0 and2_mag_2.GF_INV_MAG_0.IN VDD.t10 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X7 a_1862_738# and2_mag_1.IN2 VSS.t18 VSS.t17 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X8 and2_mag_0.GF_INV_MAG_0.IN B.t0 VDD.t16 VDD.t15 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X9 and2_mag_1.GF_INV_MAG_0.IN C.t1 a_1862_738# VSS.t0 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X10 and2_mag_2.GF_INV_MAG_0.IN and2_mag_2.IN2 VDD.t14 VDD.t13 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X11 a_916_743# B.t1 VSS.t9 VSS.t8 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X12 and2_mag_2.GF_INV_MAG_0.IN D.t1 a_2813_727# VSS.t5 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X13 and2_mag_2.IN2 and2_mag_1.GF_INV_MAG_0.IN VDD.t25 VDD.t24 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X14 and2_mag_1.IN2 and2_mag_0.GF_INV_MAG_0.IN VSS.t4 VSS.t3 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X15 a_3777_738# and2_mag_3.IN2 VSS.t11 VSS.t10 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X16 and2_mag_2.IN2 and2_mag_1.GF_INV_MAG_0.IN VSS.t16 VSS.t15 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X17 and2_mag_3.IN2 and2_mag_2.GF_INV_MAG_0.IN VDD.t7 VDD.t6 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X18 VDD E.t0 and2_mag_3.GF_INV_MAG_0.IN VDD.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X19 and2_mag_3.GF_INV_MAG_0.IN E.t1 a_3777_738# VSS.t14 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X20 and2_mag_3.GF_INV_MAG_0.IN and2_mag_3.IN2 VDD.t18 VDD.t17 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X21 and2_mag_3.IN2 and2_mag_2.GF_INV_MAG_0.IN VSS.t2 VSS.t1 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X22 VDD A.t1 and2_mag_0.GF_INV_MAG_0.IN VDD.t19 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X23 and2_mag_1.IN2 and2_mag_0.GF_INV_MAG_0.IN VDD.t9 VDD.t8 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
R0 C.n2 C.t1 31.528
R1 C.n2 C.t0 15.3826
R2 C.n3 C.n2 5.75592
R3 C.n7 C.n5 2.52047
R4 C.n7 C.n6 2.26996
R5 C.n1 C.n0 2.24713
R6 C.n5 C.n4 2.24658
R7 C.n0 C 0.0565142
R8 C C.n7 0.0199595
R9 C.n4 C.n3 0.0191207
R10 C.n5 C.n1 0.0105495
R11 VDD.n21 VDD.t26 13882.6
R12 VDD.n15 VDD.t13 12382.6
R13 VDD.n10 VDD.t17 7208.33
R14 VDD VDD.n21 451.327
R15 VDD VDD.n15 445.577
R16 VDD VDD.n10 431.3
R17 VDD VDD.n5 425.019
R18 VDD.n15 VDD.t3 378.788
R19 VDD.n10 VDD.t10 378.788
R20 VDD.n5 VDD.t0 378.788
R21 VDD.n23 VDD.t19 193.183
R22 VDD.n20 VDD.t3 193.183
R23 VDD.n14 VDD.t10 193.183
R24 VDD.n9 VDD.t0 193.183
R25 VDD.n23 VDD.t15 109.849
R26 VDD.t26 VDD.n20 109.849
R27 VDD.t13 VDD.n14 109.849
R28 VDD.t17 VDD.n9 109.849
R29 VDD.n21 VDD.t8 62.8277
R30 VDD.n15 VDD.t24 62.016
R31 VDD.n10 VDD.t6 60.0005
R32 VDD.n5 VDD.t22 59.1138
R33 VDD.n24 VDD.n23 6.3005
R34 VDD.n9 VDD.n8 6.3005
R35 VDD.n14 VDD.n13 6.3005
R36 VDD.n20 VDD.n19 6.3005
R37 VDD VDD.t16 5.1878
R38 VDD.n25 VDD.n22 5.13287
R39 VDD.n3 VDD.t18 5.13287
R40 VDD.n7 VDD.n4 5.13287
R41 VDD.n1 VDD.t14 5.13287
R42 VDD.n12 VDD.n2 5.13287
R43 VDD.n18 VDD.t27 5.13287
R44 VDD.n17 VDD.n0 5.13287
R45 VDD.n6 VDD.t23 5.09407
R46 VDD.n11 VDD.t7 5.09407
R47 VDD.n16 VDD.t25 5.09407
R48 VDD.n26 VDD.t9 5.09407
R49 VDD VDD.n3 0.126036
R50 VDD VDD.n1 0.12226
R51 VDD.n18 VDD 0.11887
R52 VDD.n26 VDD.n25 0.0984239
R53 VDD.n7 VDD.n6 0.0962255
R54 VDD.n17 VDD.n16 0.0962255
R55 VDD.n12 VDD.n11 0.0917202
R56 VDD.n25 VDD.n24 0.0782465
R57 VDD.n8 VDD.n7 0.0764633
R58 VDD.n19 VDD.n17 0.0764633
R59 VDD.n13 VDD.n12 0.0728144
R60 VDD VDD.n3 0.0541697
R61 VDD VDD.n18 0.0541697
R62 VDD VDD.n1 0.0515917
R63 VDD VDD.n26 0.0339978
R64 VDD.n6 VDD 0.0332632
R65 VDD.n16 VDD 0.0332632
R66 VDD.n11 VDD 0.0317552
R67 VDD.n24 VDD 0.00388028
R68 VDD.n8 VDD 0.00380275
R69 VDD.n19 VDD 0.00380275
R70 VDD.n13 VDD 0.0036441
R71 A.n0 A.t0 31.528
R72 A.n0 A.t1 15.3826
R73 A.n1 A.n0 7.63442
R74 A.n3 A.n2 2.25353
R75 A.n3 A.n1 1.48351
R76 A.n1 A 0.0831009
R77 A A.n3 0.00322727
R78 VSS.t1 VSS.t10 2179.77
R79 VSS.t15 VSS.t6 2109.58
R80 VSS.t3 VSS.t17 2054.29
R81 VSS.n11 VSS.t5 527.919
R82 VSS.n17 VSS.t0 518.273
R83 VSS.n5 VSS.t14 518.273
R84 VSS.n19 VSS.t19 514.004
R85 VSS.t6 VSS.n11 351.947
R86 VSS.t17 VSS.n17 345.515
R87 VSS.t10 VSS.n5 345.515
R88 VSS.n19 VSS.t8 342.67
R89 VSS.n6 VSS.t1 32.9954
R90 VSS.n12 VSS.t15 32.3925
R91 VSS.n0 VSS.t12 32.3925
R92 VSS.n18 VSS.t3 32.1257
R93 VSS.n2 VSS.t13 9.30652
R94 VSS.n8 VSS.t2 9.30652
R95 VSS.n14 VSS.t16 9.30652
R96 VSS.n21 VSS.t4 9.30652
R97 VSS VSS.t9 7.20535
R98 VSS.n3 VSS.t11 7.13989
R99 VSS.n15 VSS.t18 7.13989
R100 VSS.n9 VSS.t7 7.12156
R101 VSS.n20 VSS.n19 5.2005
R102 VSS.n1 VSS.n0 5.2005
R103 VSS.n5 VSS.n4 5.2005
R104 VSS.n7 VSS.n6 5.2005
R105 VSS.n11 VSS.n10 5.2005
R106 VSS.n13 VSS.n12 5.2005
R107 VSS.n17 VSS.n16 5.2005
R108 VSS.n22 VSS.n18 5.2005
R109 VSS.n10 VSS.n8 0.152216
R110 VSS.n4 VSS.n2 0.151517
R111 VSS.n16 VSS.n14 0.151517
R112 VSS.n21 VSS.n20 0.151143
R113 VSS.n3 VSS 0.100904
R114 VSS.n9 VSS 0.0940347
R115 VSS.n15 VSS 0.0799976
R116 VSS VSS.n3 0.0576233
R117 VSS VSS.n9 0.0576233
R118 VSS VSS.n15 0.0576233
R119 VSS.n8 VSS.n7 0.02025
R120 VSS.n2 VSS.n1 0.0196644
R121 VSS.n14 VSS.n13 0.0196644
R122 VSS.n22 VSS.n21 0.0194096
R123 VSS.n20 VSS 0.00214384
R124 VSS.n4 VSS 0.00214384
R125 VSS.n10 VSS 0.00214384
R126 VSS.n16 VSS 0.00214384
R127 VSS.n7 VSS 0.001
R128 VSS.n1 VSS 0.000985175
R129 VSS.n13 VSS 0.000985175
R130 VSS VSS.n22 0.000978723
R131 VOUT.n2 VOUT.n1 9.33985
R132 VOUT.n2 VOUT.n0 5.17836
R133 VOUT VOUT.n2 0.0594655
R134 D.n0 D.t1 31.528
R135 D.n0 D.t0 15.3826
R136 D.n1 D.n0 7.63656
R137 D.n3 D.n1 4.925
R138 D.n3 D.n2 2.26531
R139 D.n1 D 0.0809204
R140 D D.n3 0.0153101
R141 B.n0 B.t0 30.9379
R142 B.n0 B.t1 21.6422
R143 B B.n0 4.11094
R144 E.n0 E.t1 31.528
R145 E.n0 E.t0 15.3826
R146 E.n1 E.n0 7.622
R147 E.n3 E.n1 5.05815
R148 E.n3 E.n2 2.26269
R149 E.n1 E 0.0323803
R150 E E.n3 0.0095
C0 C and2_mag_0.GF_INV_MAG_0.IN 0.0724f
C1 C and2_mag_3.IN2 1.05e-20
C2 a_916_743# and2_mag_1.GF_INV_MAG_0.IN 4.6e-21
C3 D a_2813_727# 0.0193f
C4 VOUT and2_mag_2.GF_INV_MAG_0.IN 5.82e-21
C5 VOUT VDD 0.155f
C6 C a_1862_738# 0.00943f
C7 and2_mag_1.IN2 A 0.00841f
C8 D and2_mag_0.GF_INV_MAG_0.IN 0.0126f
C9 and2_mag_1.GF_INV_MAG_0.IN C 0.318f
C10 and2_mag_2.IN2 and2_mag_1.IN2 5.06e-21
C11 a_916_743# VDD 3.14e-19
C12 a_3777_738# and2_mag_3.IN2 0.00347f
C13 D and2_mag_3.IN2 0.0127f
C14 and2_mag_2.GF_INV_MAG_0.IN C 5.23e-19
C15 C VDD 0.254f
C16 E and2_mag_1.IN2 0.0502f
C17 D a_1862_738# 0.0114f
C18 and2_mag_2.IN2 A 9.39e-21
C19 D and2_mag_1.GF_INV_MAG_0.IN 0.0263f
C20 E and2_mag_3.GF_INV_MAG_0.IN 0.3f
C21 and2_mag_2.GF_INV_MAG_0.IN D 0.314f
C22 and2_mag_2.GF_INV_MAG_0.IN a_3777_738# 8.67e-20
C23 B A 0.169f
C24 a_2813_727# and2_mag_3.IN2 8.97e-21
C25 VDD a_3777_738# 3.14e-19
C26 D VDD 0.252f
C27 E A 0.287f
C28 E and2_mag_2.IN2 0.0512f
C29 and2_mag_1.GF_INV_MAG_0.IN a_2813_727# 1.05e-20
C30 VOUT and2_mag_3.GF_INV_MAG_0.IN 0.117f
C31 E B 0.0106f
C32 and2_mag_0.GF_INV_MAG_0.IN a_1862_738# 3.85e-20
C33 C and2_mag_1.IN2 0.101f
C34 and2_mag_1.GF_INV_MAG_0.IN and2_mag_0.GF_INV_MAG_0.IN 2.23e-19
C35 and2_mag_2.GF_INV_MAG_0.IN a_2813_727# 0.069f
C36 VDD a_2813_727# 3.14e-19
C37 and2_mag_1.GF_INV_MAG_0.IN and2_mag_3.IN2 1.97e-19
C38 a_916_743# A 0.00353f
C39 and2_mag_2.GF_INV_MAG_0.IN and2_mag_0.GF_INV_MAG_0.IN 1.9e-21
C40 and2_mag_0.GF_INV_MAG_0.IN VDD 0.428f
C41 and2_mag_1.GF_INV_MAG_0.IN a_1862_738# 0.069f
C42 VOUT E 0.00921f
C43 C A 0.164f
C44 and2_mag_2.GF_INV_MAG_0.IN and2_mag_3.IN2 0.127f
C45 D and2_mag_1.IN2 0.0053f
C46 and2_mag_2.IN2 C 0.0122f
C47 VDD and2_mag_3.IN2 0.384f
C48 a_916_743# B 0.00347f
C49 and2_mag_2.GF_INV_MAG_0.IN a_1862_738# 4.56e-21
C50 VDD a_1862_738# 3.14e-19
C51 and2_mag_2.GF_INV_MAG_0.IN and2_mag_1.GF_INV_MAG_0.IN 2.17e-19
C52 C B 0.15f
C53 and2_mag_1.GF_INV_MAG_0.IN VDD 0.43f
C54 a_3777_738# and2_mag_3.GF_INV_MAG_0.IN 0.069f
C55 D and2_mag_3.GF_INV_MAG_0.IN 0.00164f
C56 E C 0.176f
C57 D A 0.00372f
C58 D and2_mag_2.IN2 0.0782f
C59 and2_mag_2.GF_INV_MAG_0.IN VDD 0.429f
C60 D B 0.00833f
C61 and2_mag_1.IN2 and2_mag_0.GF_INV_MAG_0.IN 0.129f
C62 E D 0.143f
C63 E a_3777_738# 0.00479f
C64 a_916_743# C 0.00632f
C65 and2_mag_2.IN2 a_2813_727# 0.00347f
C66 and2_mag_1.IN2 a_1862_738# 0.00347f
C67 and2_mag_0.GF_INV_MAG_0.IN A 0.298f
C68 and2_mag_2.IN2 and2_mag_0.GF_INV_MAG_0.IN 3.34e-21
C69 and2_mag_1.GF_INV_MAG_0.IN and2_mag_1.IN2 0.12f
C70 VOUT D 3.02e-19
C71 and2_mag_3.IN2 and2_mag_3.GF_INV_MAG_0.IN 0.118f
C72 and2_mag_2.IN2 and2_mag_3.IN2 4.92e-21
C73 E a_2813_727# 7.37e-19
C74 a_916_743# D 0.0108f
C75 and2_mag_0.GF_INV_MAG_0.IN B 0.0929f
C76 and2_mag_1.IN2 VDD 0.387f
C77 A a_1862_738# 3.11e-21
C78 E and2_mag_0.GF_INV_MAG_0.IN 0.0441f
C79 and2_mag_1.GF_INV_MAG_0.IN A 1.88e-19
C80 D C 0.713f
C81 and2_mag_2.IN2 and2_mag_1.GF_INV_MAG_0.IN 0.128f
C82 E and2_mag_3.IN2 0.101f
C83 and2_mag_2.GF_INV_MAG_0.IN and2_mag_3.GF_INV_MAG_0.IN 2.8e-19
C84 VDD and2_mag_3.GF_INV_MAG_0.IN 0.422f
C85 and2_mag_2.GF_INV_MAG_0.IN and2_mag_2.IN2 0.119f
C86 VDD A 0.257f
C87 and2_mag_2.IN2 VDD 0.388f
C88 E and2_mag_1.GF_INV_MAG_0.IN 0.0477f
C89 D a_3777_738# 4.35e-19
C90 a_916_743# and2_mag_0.GF_INV_MAG_0.IN 0.069f
C91 C a_2813_727# 9.22e-21
C92 B VDD 0.174f
C93 E and2_mag_2.GF_INV_MAG_0.IN 0.046f
C94 E VDD 0.97f
C95 a_3777_738# VSS 0.073f
C96 a_2813_727# VSS 0.0757f
C97 a_1862_738# VSS 0.073f
C98 VOUT VSS 0.219f
C99 a_916_743# VSS 0.072f
C100 and2_mag_3.GF_INV_MAG_0.IN VSS 0.465f
C101 E VSS 0.873f
C102 and2_mag_3.IN2 VSS 0.401f
C103 and2_mag_2.GF_INV_MAG_0.IN VSS 0.451f
C104 D VSS 1.22f
C105 and2_mag_2.IN2 VSS 0.399f
C106 and2_mag_1.GF_INV_MAG_0.IN VSS 0.446f
C107 C VSS 0.372f
C108 and2_mag_1.IN2 VSS 0.396f
C109 and2_mag_0.GF_INV_MAG_0.IN VSS 0.45f
C110 A VSS 0.276f
C111 B VSS 0.337f
C112 VDD VSS 6.76f
.ends

