* NGSPICE file created from Delay_Cell_mag_flat.ext - technology: gf180mcuC

.subckt Delay_Cell_mag_flat OUT OUTB EN VCONT INB IN VSS VDD
X0 VDD OUTB.t16 OUT.t5 VDD.t21 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X1 a_474_n2321# EN.t0 VSS.t7 VSS.t6 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X2 OUT IN.t0 a_474_n2321# VSS.t16 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X3 a_474_n2321# IN.t1 OUT.t6 VSS.t6 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X4 a_279_n79# OUT.t13 OUT.t14 VDD.t15 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X5 OUT OUTB.t17 VDD.t20 VDD.t19 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X6 OUT OUT.t11 a_279_n79# VDD.t19 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X7 VDD a_1970_n1781.t9 a_1970_n1781.t10 VDD.t6 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X8 a_279_n79# a_1970_n1781.t12 VDD.t33 VDD.t32 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X9 OUTB OUTB.t10 a_279_n79# VDD.t18 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X10 a_474_n2321# a_474_n2321# a_474_n2321# VSS.t17 nfet_03v3 ad=0.44p pd=2.88u as=4p ps=24u w=1u l=0.56u
X11 OUT IN.t2 a_474_n2321# VSS.t0 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X12 OUTB OUT.t17 VDD.t30 VDD.t18 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X13 a_474_n2321# INB.t0 OUTB.t12 VSS.t8 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X14 a_279_n79# OUT.t9 OUT.t10 VDD.t21 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X15 VDD OUTB.t19 OUT.t4 VDD.t15 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X16 a_474_n2321# INB.t1 OUTB.t13 VSS.t15 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X17 VSS VCONT.t2 a_1970_n1781.t2 VSS.t12 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X18 VDD a_1970_n1781.t14 a_279_n79# VDD.t3 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X19 a_474_n2321# a_474_n2321# a_474_n2321# VSS.t12 nfet_03v3 ad=0.26p pd=1.52u as=0 ps=0 w=1u l=0.56u
X20 a_279_n79# OUTB.t8 OUTB.t9 VDD.t14 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X21 OUT OUT.t7 a_279_n79# VDD.t11 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X22 VDD a_1970_n1781.t5 a_1970_n1781.t6 VDD.t32 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X23 VSS EN.t1 a_474_n2321# VSS.t3 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X24 VDD OUT.t19 OUTB.t3 VDD.t10 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X25 a_474_n2321# IN.t3 OUT.t1 VSS.t2 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X26 OUTB INB.t2 a_474_n2321# VSS.t3 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X27 a_279_n79# a_1970_n1781.t15 VDD.t9 VDD.t6 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X28 OUTB OUTB.t6 a_279_n79# VDD.t13 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X29 OUT OUTB.t21 VDD.t12 VDD.t11 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X30 VSS VCONT.t3 a_1970_n1781.t1 VSS.t1 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X31 OUTB INB.t3 a_474_n2321# VSS.t1 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X32 VDD a_1970_n1781.t16 a_279_n79# VDD.t0 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X33 a_279_n79# OUTB.t4 OUTB.t5 VDD.t10 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X34 OUTB OUT.t20 VDD.t27 VDD.t13 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X35 VDD OUT.t21 OUTB.t15 VDD.t14 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
R0 OUTB.n20 OUTB.t19 22.2916
R1 OUTB.n6 OUTB.t10 22.1612
R2 OUTB.t19 OUTB.n19 17.311
R3 OUTB.n8 OUTB.t4 15.1219
R4 OUTB.n7 OUTB.n6 14.0791
R5 OUTB.n21 OUTB.n20 14.0791
R6 OUTB.n22 OUTB.n21 14.0791
R7 OUTB.n20 OUTB.t21 8.213
R8 OUTB.n21 OUTB.t16 8.213
R9 OUTB.n22 OUTB.t17 8.213
R10 OUTB.n7 OUTB.t6 8.08264
R11 OUTB.n6 OUTB.t8 8.08264
R12 OUTB.n8 OUTB.n7 7.03979
R13 OUTB OUTB.n22 5.02734
R14 OUTB.n16 OUTB.n15 4.70398
R15 OUTB.n17 OUTB.n16 4.4843
R16 OUTB.n9 OUTB.n8 4.0005
R17 OUTB.n19 OUTB.n1 3.3342
R18 OUTB.n16 OUTB.n13 3.1505
R19 OUTB.n9 OUTB.n5 2.94411
R20 OUTB.n19 OUTB.n3 2.9292
R21 OUTB.n17 OUTB.n11 2.6005
R22 OUTB.n11 OUTB.t3 1.8205
R23 OUTB.n11 OUTB.n10 1.8205
R24 OUTB.n5 OUTB.t5 1.8205
R25 OUTB.n5 OUTB.n4 1.8205
R26 OUTB.n3 OUTB.t15 1.8205
R27 OUTB.n3 OUTB.n2 1.8205
R28 OUTB.n1 OUTB.t9 1.8205
R29 OUTB.n1 OUTB.n0 1.8205
R30 OUTB.n13 OUTB.t13 1.6385
R31 OUTB.n13 OUTB.n12 1.6385
R32 OUTB.n15 OUTB.t12 1.6385
R33 OUTB.n15 OUTB.n14 1.6385
R34 OUTB.n19 OUTB.n18 0.845717
R35 OUTB.n18 OUTB.n9 0.335065
R36 OUTB.n18 OUTB.n17 0.329196
R37 OUT.n10 OUT.t19 22.3568
R38 OUT.n22 OUT.t13 22.096
R39 OUT.n9 OUT.t17 19.4889
R40 OUT.n23 OUT.n22 14.0791
R41 OUT.n24 OUT.n23 14.0791
R42 OUT.n11 OUT.n10 9.33211
R43 OUT.n10 OUT.t20 8.27818
R44 OUT.n8 OUT.t21 8.27818
R45 OUT.n22 OUT.t7 8.01746
R46 OUT.n23 OUT.t9 8.01746
R47 OUT.n24 OUT.t11 8.01746
R48 OUT.n25 OUT.n24 4.89822
R49 OUT.n16 OUT.n15 4.67659
R50 OUT.n17 OUT.n16 3.51328
R51 OUT.n21 OUT.n3 3.20507
R52 OUT.n16 OUT.n13 3.1505
R53 OUT.n20 OUT.n5 3.02311
R54 OUT.n21 OUT.n1 2.98985
R55 OUT.n9 OUT.n8 2.86836
R56 OUT.n19 OUT.n7 2.6005
R57 OUT.n18 OUT.n9 2.11815
R58 OUT.n7 OUT.t4 1.8205
R59 OUT.n7 OUT.n6 1.8205
R60 OUT.n5 OUT.t14 1.8205
R61 OUT.n5 OUT.n4 1.8205
R62 OUT.n3 OUT.t5 1.8205
R63 OUT.n3 OUT.n2 1.8205
R64 OUT.n1 OUT.t10 1.8205
R65 OUT.n1 OUT.n0 1.8205
R66 OUT.n13 OUT.t6 1.6385
R67 OUT.n13 OUT.n12 1.6385
R68 OUT.n15 OUT.t1 1.6385
R69 OUT.n15 OUT.n14 1.6385
R70 OUT.n17 OUT.n11 1.50108
R71 OUT.n19 OUT.n18 1.26616
R72 OUT.n21 OUT.n20 0.826273
R73 OUT.n20 OUT.n19 0.640283
R74 OUT OUT.n25 0.1605
R75 OUT.n25 OUT.n21 0.124944
R76 OUT.n18 OUT.n17 0.0603098
R77 VDD.n48 VDD.t6 42.1692
R78 VDD.n45 VDD.t3 35.5427
R79 VDD.n15 VDD.t19 30.7234
R80 VDD.n42 VDD.t32 28.9162
R81 VDD.n18 VDD.t21 24.0969
R82 VDD.n39 VDD.t0 22.2897
R83 VDD.n21 VDD.t11 17.4704
R84 VDD.n36 VDD.t10 15.6632
R85 VDD.n24 VDD.t15 10.8439
R86 VDD.n33 VDD.t13 9.03664
R87 VDD.n27 VDD.t18 4.21737
R88 VDD.n136 VDD.n135 3.9192
R89 VDD.n117 VDD.t20 3.80738
R90 VDD.n76 VDD.n66 3.1505
R91 VDD.n102 VDD.n101 3.1505
R92 VDD.n100 VDD.n99 3.1505
R93 VDD.n98 VDD.n97 3.1505
R94 VDD.n96 VDD.n95 3.1505
R95 VDD.n94 VDD.n93 3.1505
R96 VDD.n92 VDD.n91 3.1505
R97 VDD.n90 VDD.n89 3.1505
R98 VDD.n88 VDD.n87 3.1505
R99 VDD.n86 VDD.n85 3.1505
R100 VDD.n84 VDD.n83 3.1505
R101 VDD.n82 VDD.n81 3.1505
R102 VDD.n80 VDD.n79 3.1505
R103 VDD.n78 VDD.n77 3.1505
R104 VDD.n5 VDD.n4 3.1505
R105 VDD.n2 VDD.n1 3.1505
R106 VDD.n68 VDD.n67 3.1505
R107 VDD.n70 VDD.n69 3.1505
R108 VDD.n73 VDD.n72 3.1505
R109 VDD.n7 VDD.n6 3.1505
R110 VDD.n75 VDD.n74 3.1505
R111 VDD.n11 VDD.n10 3.1505
R112 VDD.n13 VDD.n12 3.1505
R113 VDD.n14 VDD.n13 3.1505
R114 VDD.n17 VDD.n16 3.1505
R115 VDD.n16 VDD.n15 3.1505
R116 VDD.n20 VDD.n19 3.1505
R117 VDD.n19 VDD.n18 3.1505
R118 VDD.n23 VDD.n22 3.1505
R119 VDD.n22 VDD.n21 3.1505
R120 VDD.n26 VDD.n25 3.1505
R121 VDD.n25 VDD.n24 3.1505
R122 VDD.n29 VDD.n28 3.1505
R123 VDD.n28 VDD.n27 3.1505
R124 VDD.n32 VDD.n31 3.1505
R125 VDD.n31 VDD.n30 3.1505
R126 VDD.n35 VDD.n34 3.1505
R127 VDD.n34 VDD.n33 3.1505
R128 VDD.n38 VDD.n37 3.1505
R129 VDD.n37 VDD.n36 3.1505
R130 VDD.n41 VDD.n40 3.1505
R131 VDD.n40 VDD.n39 3.1505
R132 VDD.n44 VDD.n43 3.1505
R133 VDD.n43 VDD.n42 3.1505
R134 VDD.n47 VDD.n46 3.1505
R135 VDD.n46 VDD.n45 3.1505
R136 VDD.n50 VDD.n49 3.1505
R137 VDD.n49 VDD.n48 3.1505
R138 VDD.n53 VDD.n52 3.1505
R139 VDD.n52 VDD.n51 3.1505
R140 VDD.n108 VDD.n107 3.1505
R141 VDD.n110 VDD.n109 3.1505
R142 VDD.n113 VDD.n112 3.1505
R143 VDD.n65 VDD.n64 3.1505
R144 VDD.n61 VDD.n60 3.1505
R145 VDD.n58 VDD.n57 3.1505
R146 VDD.n104 VDD.n103 3.1505
R147 VDD.n56 VDD.n55 3.1505
R148 VDD.n136 VDD.n133 3.07111
R149 VDD.n60 VDD.n59 3.001
R150 VDD.n64 VDD.n62 3.001
R151 VDD.n64 VDD.n63 3.001
R152 VDD.n112 VDD.n111 3.001
R153 VDD.n131 VDD.n130 2.64616
R154 VDD.n30 VDD.t14 2.41014
R155 VDD.n1 VDD.n0 2.03394
R156 VDD.n72 VDD.n71 2.03336
R157 VDD.n133 VDD.t9 1.8205
R158 VDD.n133 VDD.n132 1.8205
R159 VDD.n135 VDD.t33 1.8205
R160 VDD.n135 VDD.n134 1.8205
R161 VDD.n116 VDD.t12 1.8205
R162 VDD.n116 VDD.n115 1.8205
R163 VDD.n119 VDD.t30 1.8205
R164 VDD.n119 VDD.n118 1.8205
R165 VDD.n122 VDD.t27 1.8205
R166 VDD.n122 VDD.n121 1.8205
R167 VDD.n125 VDD.t24 1.8205
R168 VDD.n125 VDD.n124 1.8205
R169 VDD.n128 VDD.t31 1.8205
R170 VDD.n128 VDD.n127 1.8205
R171 VDD.n10 VDD.n9 1.72716
R172 VDD.n55 VDD.n54 1.72716
R173 VDD.n4 VDD.n3 1.72703
R174 VDD.n107 VDD.n106 1.72703
R175 VDD.n117 VDD.n116 1.42427
R176 VDD.n120 VDD.n119 1.42427
R177 VDD.n123 VDD.n122 1.42427
R178 VDD.n126 VDD.n125 1.42427
R179 VDD.n129 VDD.n128 1.42427
R180 VDD.n131 VDD.n129 1.16194
R181 VDD.n9 VDD.n8 0.950516
R182 VDD.n106 VDD.n105 0.950315
R183 VDD.n120 VDD.n117 0.562605
R184 VDD.n123 VDD.n120 0.562605
R185 VDD.n126 VDD.n123 0.562605
R186 VDD.n129 VDD.n126 0.562605
R187 VDD.n137 VDD.n136 0.418343
R188 VDD.n137 VDD.n131 0.41547
R189 VDD.n102 VDD.n100 0.185
R190 VDD.n100 VDD.n98 0.185
R191 VDD.n98 VDD.n96 0.185
R192 VDD.n96 VDD.n94 0.185
R193 VDD.n94 VDD.n92 0.185
R194 VDD.n92 VDD.n90 0.185
R195 VDD.n90 VDD.n88 0.185
R196 VDD.n88 VDD.n86 0.185
R197 VDD.n86 VDD.n84 0.185
R198 VDD.n84 VDD.n82 0.185
R199 VDD.n82 VDD.n80 0.185
R200 VDD.n80 VDD.n78 0.185
R201 VDD.n78 VDD.n76 0.185
R202 VDD.n53 VDD.n50 0.185
R203 VDD.n50 VDD.n47 0.185
R204 VDD.n47 VDD.n44 0.185
R205 VDD.n44 VDD.n41 0.185
R206 VDD.n41 VDD.n38 0.185
R207 VDD.n38 VDD.n35 0.185
R208 VDD.n35 VDD.n32 0.185
R209 VDD.n32 VDD.n29 0.185
R210 VDD.n29 VDD.n26 0.185
R211 VDD.n26 VDD.n23 0.185
R212 VDD.n23 VDD.n20 0.185
R213 VDD.n20 VDD.n17 0.185
R214 VDD.n17 VDD.n14 0.185
R215 VDD.n14 VDD.n11 0.172236
R216 VDD.n11 VDD.n7 0.164136
R217 VDD.n7 VDD.n5 0.164136
R218 VDD.n5 VDD.n2 0.164136
R219 VDD.n70 VDD.n68 0.164136
R220 VDD.n73 VDD.n70 0.164136
R221 VDD.n75 VDD.n73 0.164136
R222 VDD.n58 VDD.n56 0.164136
R223 VDD.n61 VDD.n58 0.164136
R224 VDD.n65 VDD.n61 0.164136
R225 VDD.n113 VDD.n110 0.164136
R226 VDD.n110 VDD.n108 0.164136
R227 VDD.n108 VDD.n104 0.164136
R228 VDD.n114 VDD.n113 0.161682
R229 VDD.n56 VDD.n53 0.151536
R230 VDD.n76 VDD.n75 0.137873
R231 VDD VDD.n114 0.130885
R232 VDD.n104 VDD.n102 0.117173
R233 VDD VDD.n137 0.0374231
R234 VDD.n114 VDD.n65 0.00295455
R235 EN EN.n0 60.8984
R236 EN.n0 EN.t1 22.6826
R237 EN.n0 EN.t0 8.60407
R238 VSS.n10 VSS.n9 513.072
R239 VSS.n61 VSS.n60 393.962
R240 VSS.n133 VSS.t12 144.998
R241 VSS.n136 VSS.t8 122.213
R242 VSS.n139 VSS.t1 99.4269
R243 VSS.n142 VSS.t15 76.6417
R244 VSS.n160 VSS.t17 60.0706
R245 VSS.n145 VSS.t3 53.8565
R246 VSS.n117 VSS.n116 45.5709
R247 VSS.n228 VSS.n227 43.4995
R248 VSS.n157 VSS.t16 37.2854
R249 VSS.n148 VSS.t6 31.0712
R250 VSS.n154 VSS.t2 14.5002
R251 VSS.n151 VSS.t0 8.28603
R252 VSS.n5 VSS.n4 5.99763
R253 VSS.n7 VSS.t7 5.0898
R254 VSS.n5 VSS.n3 3.51441
R255 VSS.n6 VSS.n1 3.51441
R256 VSS.n11 VSS.n10 2.60693
R257 VSS.n194 VSS.n186 2.60371
R258 VSS.n230 VSS.n229 2.60243
R259 VSS.n123 VSS.n122 2.60179
R260 VSS.n226 VSS.n225 2.6005
R261 VSS.n196 VSS.n195 2.6005
R262 VSS.n198 VSS.n197 2.6005
R263 VSS.n200 VSS.n199 2.6005
R264 VSS.n202 VSS.n201 2.6005
R265 VSS.n204 VSS.n203 2.6005
R266 VSS.n206 VSS.n205 2.6005
R267 VSS.n208 VSS.n207 2.6005
R268 VSS.n210 VSS.n209 2.6005
R269 VSS.n212 VSS.n211 2.6005
R270 VSS.n214 VSS.n213 2.6005
R271 VSS.n216 VSS.n215 2.6005
R272 VSS.n218 VSS.n217 2.6005
R273 VSS.n220 VSS.n219 2.6005
R274 VSS.n222 VSS.n221 2.6005
R275 VSS.n224 VSS.n223 2.6005
R276 VSS.n86 VSS.n85 2.6005
R277 VSS.n85 VSS.n84 2.6005
R278 VSS.n68 VSS.n67 2.6005
R279 VSS.n67 VSS.n66 2.6005
R280 VSS.n71 VSS.n70 2.6005
R281 VSS.n70 VSS.n69 2.6005
R282 VSS.n74 VSS.n73 2.6005
R283 VSS.n73 VSS.n72 2.6005
R284 VSS.n77 VSS.n76 2.6005
R285 VSS.n76 VSS.n75 2.6005
R286 VSS.n80 VSS.n79 2.6005
R287 VSS.n79 VSS.n78 2.6005
R288 VSS.n83 VSS.n82 2.6005
R289 VSS.n82 VSS.n81 2.6005
R290 VSS.n65 VSS.n64 2.6005
R291 VSS.n64 VSS.n63 2.6005
R292 VSS.n14 VSS.n13 2.6005
R293 VSS.n13 VSS.n12 2.6005
R294 VSS.n17 VSS.n16 2.6005
R295 VSS.n16 VSS.n15 2.6005
R296 VSS.n20 VSS.n19 2.6005
R297 VSS.n19 VSS.n18 2.6005
R298 VSS.n23 VSS.n22 2.6005
R299 VSS.n22 VSS.n21 2.6005
R300 VSS.n26 VSS.n25 2.6005
R301 VSS.n25 VSS.n24 2.6005
R302 VSS.n29 VSS.n28 2.6005
R303 VSS.n28 VSS.n27 2.6005
R304 VSS.n32 VSS.n31 2.6005
R305 VSS.n31 VSS.n30 2.6005
R306 VSS.n35 VSS.n34 2.6005
R307 VSS.n34 VSS.n33 2.6005
R308 VSS.n38 VSS.n37 2.6005
R309 VSS.n37 VSS.n36 2.6005
R310 VSS.n41 VSS.n40 2.6005
R311 VSS.n40 VSS.n39 2.6005
R312 VSS.n44 VSS.n43 2.6005
R313 VSS.n43 VSS.n42 2.6005
R314 VSS.n47 VSS.n46 2.6005
R315 VSS.n46 VSS.n45 2.6005
R316 VSS.n50 VSS.n49 2.6005
R317 VSS.n49 VSS.n48 2.6005
R318 VSS.n53 VSS.n52 2.6005
R319 VSS.n52 VSS.n51 2.6005
R320 VSS.n56 VSS.n55 2.6005
R321 VSS.n55 VSS.n54 2.6005
R322 VSS.n59 VSS.n58 2.6005
R323 VSS.n58 VSS.n57 2.6005
R324 VSS.n62 VSS.n61 2.6005
R325 VSS.n110 VSS.n109 2.6005
R326 VSS.n109 VSS.n108 2.6005
R327 VSS.n107 VSS.n106 2.6005
R328 VSS.n106 VSS.n105 2.6005
R329 VSS.n104 VSS.n103 2.6005
R330 VSS.n103 VSS.n102 2.6005
R331 VSS.n101 VSS.n100 2.6005
R332 VSS.n100 VSS.n99 2.6005
R333 VSS.n98 VSS.n97 2.6005
R334 VSS.n97 VSS.n96 2.6005
R335 VSS.n95 VSS.n94 2.6005
R336 VSS.n94 VSS.n93 2.6005
R337 VSS.n92 VSS.n91 2.6005
R338 VSS.n91 VSS.n90 2.6005
R339 VSS.n89 VSS.n88 2.6005
R340 VSS.n88 VSS.n87 2.6005
R341 VSS.n120 VSS.n119 2.6005
R342 VSS.n115 VSS.n114 2.6005
R343 VSS.n113 VSS.n112 2.6005
R344 VSS.n188 VSS.n187 2.6005
R345 VSS.n190 VSS.n189 2.6005
R346 VSS.n193 VSS.n192 2.6005
R347 VSS.n170 VSS.n169 2.6005
R348 VSS.n126 VSS.n125 2.6005
R349 VSS.n125 VSS.n124 2.6005
R350 VSS.n129 VSS.n128 2.6005
R351 VSS.n128 VSS.n127 2.6005
R352 VSS.n132 VSS.n131 2.6005
R353 VSS.n131 VSS.n130 2.6005
R354 VSS.n135 VSS.n134 2.6005
R355 VSS.n134 VSS.n133 2.6005
R356 VSS.n138 VSS.n137 2.6005
R357 VSS.n137 VSS.n136 2.6005
R358 VSS.n141 VSS.n140 2.6005
R359 VSS.n140 VSS.n139 2.6005
R360 VSS.n144 VSS.n143 2.6005
R361 VSS.n143 VSS.n142 2.6005
R362 VSS.n147 VSS.n146 2.6005
R363 VSS.n146 VSS.n145 2.6005
R364 VSS.n150 VSS.n149 2.6005
R365 VSS.n149 VSS.n148 2.6005
R366 VSS.n153 VSS.n152 2.6005
R367 VSS.n152 VSS.n151 2.6005
R368 VSS.n156 VSS.n155 2.6005
R369 VSS.n155 VSS.n154 2.6005
R370 VSS.n159 VSS.n158 2.6005
R371 VSS.n158 VSS.n157 2.6005
R372 VSS.n162 VSS.n161 2.6005
R373 VSS.n161 VSS.n160 2.6005
R374 VSS.n165 VSS.n164 2.6005
R375 VSS.n164 VSS.n163 2.6005
R376 VSS.n168 VSS.n167 2.6005
R377 VSS.n167 VSS.n166 2.6005
R378 VSS.n171 VSS.n170 2.6005
R379 VSS.n174 VSS.n173 2.6005
R380 VSS.n180 VSS.n179 2.6005
R381 VSS.n184 VSS.n183 2.6005
R382 VSS.n237 VSS.n236 2.6005
R383 VSS.n235 VSS.n234 2.6005
R384 VSS.n232 VSS.n231 2.6005
R385 VSS.n177 VSS.n176 2.6005
R386 VSS.n229 VSS.n228 2.6005
R387 VSS.n119 VSS.n118 1.7266
R388 VSS.n112 VSS.n111 1.7266
R389 VSS.n192 VSS.n191 1.72602
R390 VSS.n179 VSS.n178 1.72592
R391 VSS.n183 VSS.n182 1.72592
R392 VSS.n234 VSS.n233 1.72592
R393 VSS.n3 VSS.t9 1.6385
R394 VSS.n3 VSS.n2 1.6385
R395 VSS.n1 VSS.t18 1.6385
R396 VSS.n1 VSS.n0 1.6385
R397 VSS VSS.n7 1.46704
R398 VSS.n6 VSS.n5 0.845717
R399 VSS.n7 VSS.n6 0.827256
R400 VSS.n10 VSS.n8 0.5005
R401 VSS.n118 VSS.n117 0.438783
R402 VSS.n182 VSS.n181 0.43854
R403 VSS.n186 VSS.n185 0.2505
R404 VSS VSS.n238 0.224346
R405 VSS.n196 VSS.n194 0.149643
R406 VSS.n126 VSS.n123 0.149643
R407 VSS.n62 VSS.n59 0.147071
R408 VSS.n198 VSS.n196 0.132286
R409 VSS.n200 VSS.n198 0.132286
R410 VSS.n202 VSS.n200 0.132286
R411 VSS.n204 VSS.n202 0.132286
R412 VSS.n206 VSS.n204 0.132286
R413 VSS.n208 VSS.n206 0.132286
R414 VSS.n210 VSS.n208 0.132286
R415 VSS.n212 VSS.n210 0.132286
R416 VSS.n214 VSS.n212 0.132286
R417 VSS.n216 VSS.n214 0.132286
R418 VSS.n218 VSS.n216 0.132286
R419 VSS.n220 VSS.n218 0.132286
R420 VSS.n222 VSS.n220 0.132286
R421 VSS.n224 VSS.n222 0.132286
R422 VSS.n226 VSS.n224 0.132286
R423 VSS.n68 VSS.n65 0.132286
R424 VSS.n71 VSS.n68 0.132286
R425 VSS.n74 VSS.n71 0.132286
R426 VSS.n77 VSS.n74 0.132286
R427 VSS.n80 VSS.n77 0.132286
R428 VSS.n83 VSS.n80 0.132286
R429 VSS.n86 VSS.n83 0.132286
R430 VSS.n17 VSS.n14 0.132286
R431 VSS.n20 VSS.n17 0.132286
R432 VSS.n23 VSS.n20 0.132286
R433 VSS.n26 VSS.n23 0.132286
R434 VSS.n29 VSS.n26 0.132286
R435 VSS.n32 VSS.n29 0.132286
R436 VSS.n35 VSS.n32 0.132286
R437 VSS.n38 VSS.n35 0.132286
R438 VSS.n41 VSS.n38 0.132286
R439 VSS.n44 VSS.n41 0.132286
R440 VSS.n47 VSS.n44 0.132286
R441 VSS.n50 VSS.n47 0.132286
R442 VSS.n53 VSS.n50 0.132286
R443 VSS.n56 VSS.n53 0.132286
R444 VSS.n59 VSS.n56 0.132286
R445 VSS.n92 VSS.n89 0.132286
R446 VSS.n95 VSS.n92 0.132286
R447 VSS.n98 VSS.n95 0.132286
R448 VSS.n101 VSS.n98 0.132286
R449 VSS.n104 VSS.n101 0.132286
R450 VSS.n107 VSS.n104 0.132286
R451 VSS.n110 VSS.n107 0.132286
R452 VSS.n120 VSS.n115 0.132286
R453 VSS.n115 VSS.n113 0.132286
R454 VSS.n190 VSS.n188 0.132286
R455 VSS.n193 VSS.n190 0.132286
R456 VSS.n129 VSS.n126 0.132286
R457 VSS.n132 VSS.n129 0.132286
R458 VSS.n135 VSS.n132 0.132286
R459 VSS.n138 VSS.n135 0.132286
R460 VSS.n141 VSS.n138 0.132286
R461 VSS.n144 VSS.n141 0.132286
R462 VSS.n147 VSS.n144 0.132286
R463 VSS.n150 VSS.n147 0.132286
R464 VSS.n153 VSS.n150 0.132286
R465 VSS.n156 VSS.n153 0.132286
R466 VSS.n159 VSS.n156 0.132286
R467 VSS.n162 VSS.n159 0.132286
R468 VSS.n165 VSS.n162 0.132286
R469 VSS.n168 VSS.n165 0.132286
R470 VSS.n171 VSS.n168 0.132286
R471 VSS.n180 VSS.n177 0.132286
R472 VSS.n184 VSS.n180 0.132286
R473 VSS.n237 VSS.n235 0.132286
R474 VSS.n235 VSS.n232 0.132286
R475 VSS.n14 VSS.n11 0.125857
R476 VSS.n232 VSS.n230 0.124571
R477 VSS.n238 VSS.n237 0.123929
R478 VSS.n174 VSS.n171 0.123286
R479 VSS.n175 VSS.n86 0.102071
R480 VSS.n123 VSS.n110 0.102071
R481 VSS.n122 VSS.n121 0.1005
R482 VSS.n173 VSS.n172 0.1005
R483 VSS.n65 VSS.n62 0.0962857
R484 VSS.n230 VSS.n226 0.0795714
R485 VSS.n194 VSS.n193 0.0795714
R486 VSS.n123 VSS.n120 0.0725
R487 VSS.n177 VSS.n175 0.0725
R488 VSS.n238 VSS.n184 0.00885714
R489 VSS.n175 VSS.n174 0.00178571
R490 IN.n0 IN.t0 21.774
R491 IN.n1 IN.n0 12.7222
R492 IN.n2 IN.t1 11.9934
R493 IN.n2 IN.n1 9.78115
R494 IN.n0 IN.t3 6.51836
R495 IN.n1 IN.t2 6.51836
R496 IN IN.n2 4.47602
R497 a_1970_n1781.t9 a_1970_n1781.n5 22.8782
R498 a_1970_n1781.n6 a_1970_n1781.t9 22.4219
R499 a_1970_n1781.n3 a_1970_n1781.t16 22.2916
R500 a_1970_n1781.n5 a_1970_n1781.n4 14.0791
R501 a_1970_n1781.n4 a_1970_n1781.n3 14.0791
R502 a_1970_n1781.n7 a_1970_n1781.n6 14.0791
R503 a_1970_n1781.n1 a_1970_n1781.t3 11.3416
R504 a_1970_n1781.n6 a_1970_n1781.t7 8.34336
R505 a_1970_n1781.n7 a_1970_n1781.t5 8.34336
R506 a_1970_n1781.n5 a_1970_n1781.t15 8.213
R507 a_1970_n1781.n4 a_1970_n1781.t14 8.213
R508 a_1970_n1781.n3 a_1970_n1781.t12 8.213
R509 a_1970_n1781.n2 a_1970_n1781.n7 8.17193
R510 a_1970_n1781.n0 a_1970_n1781.n1 4.0005
R511 a_1970_n1781.n18 a_1970_n1781.n2 3.63045
R512 a_1970_n1781.n0 a_1970_n1781.n9 2.89398
R513 a_1970_n1781.n14 a_1970_n1781.n11 2.26392
R514 a_1970_n1781.n9 a_1970_n1781.t6 1.8205
R515 a_1970_n1781.n9 a_1970_n1781.n8 1.8205
R516 a_1970_n1781.t10 a_1970_n1781.n18 1.8205
R517 a_1970_n1781.n18 a_1970_n1781.n17 1.8205
R518 a_1970_n1781.n11 a_1970_n1781.t1 1.6385
R519 a_1970_n1781.n11 a_1970_n1781.n10 1.6385
R520 a_1970_n1781.n13 a_1970_n1781.t2 1.6385
R521 a_1970_n1781.n13 a_1970_n1781.n12 1.6385
R522 a_1970_n1781.n1 a_1970_n1781.n16 1.62996
R523 a_1970_n1781.n14 a_1970_n1781.n13 1.4936
R524 a_1970_n1781.n0 a_1970_n1781.n15 1.22554
R525 a_1970_n1781.n15 a_1970_n1781.n14 1.18673
R526 a_1970_n1781.n2 a_1970_n1781.n0 0.1505
R527 VCONT.n0 VCONT.t1 21.8873
R528 VCONT.n1 VCONT.n0 12.5576
R529 VCONT.n2 VCONT.t2 12.1889
R530 VCONT.n2 VCONT.n1 9.69888
R531 VCONT.n0 VCONT.t3 6.51836
R532 VCONT.n1 VCONT.t0 6.51836
R533 VCONT VCONT.n2 4.63297
R534 INB.n0 INB.t2 21.8182
R535 INB.n1 INB.n0 12.6801
R536 INB.n2 INB.t0 12.0585
R537 INB.n2 INB.n1 9.76014
R538 INB.n0 INB.t1 6.51836
R539 INB.n1 INB.t3 6.51836
R540 INB INB.n2 4.49657
C0 a_279_n79# OUTB 0.456f
C1 VCONT INB 0.0184f
C2 OUTB VCONT 0.0287f
C3 a_474_n2321# VCONT 0.0291f
C4 OUT IN 0.238f
C5 a_279_n79# VCONT 8.3e-20
C6 OUT EN 0.0484f
C7 IN EN 0.0168f
C8 OUT VDD 2.93f
C9 OUT INB 0.00336f
C10 VDD IN 2.07e-19
C11 OUT OUTB 0.828f
C12 OUT a_474_n2321# 0.499f
C13 IN INB 0.0297f
C14 VDD EN 0.051f
C15 IN OUTB 0.0201f
C16 IN a_474_n2321# 0.195f
C17 EN INB 0.00514f
C18 OUT a_279_n79# 0.5f
C19 EN OUTB 0.0276f
C20 a_474_n2321# EN 0.151f
C21 VDD INB 7.21e-19
C22 OUT VCONT 0.00241f
C23 VDD OUTB 3.04f
C24 VDD a_474_n2321# 0.0575f
C25 a_279_n79# EN 8.31e-20
C26 OUTB INB 0.243f
C27 a_474_n2321# INB 0.188f
C28 EN VCONT 0.023f
C29 a_474_n2321# OUTB 0.4f
C30 VDD a_279_n79# 1.15f
C31 VDD VCONT 0.0334f
.ends

