magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1484 -1019 1484 1019
<< metal1 >>
rect -484 13 484 19
rect -484 -13 -478 13
rect -452 -13 -416 13
rect -390 -13 -354 13
rect -328 -13 -292 13
rect -266 -13 -230 13
rect -204 -13 -168 13
rect -142 -13 -106 13
rect -80 -13 -44 13
rect -18 -13 18 13
rect 44 -13 80 13
rect 106 -13 142 13
rect 168 -13 204 13
rect 230 -13 266 13
rect 292 -13 328 13
rect 354 -13 390 13
rect 416 -13 452 13
rect 478 -13 484 13
rect -484 -19 484 -13
<< via1 >>
rect -478 -13 -452 13
rect -416 -13 -390 13
rect -354 -13 -328 13
rect -292 -13 -266 13
rect -230 -13 -204 13
rect -168 -13 -142 13
rect -106 -13 -80 13
rect -44 -13 -18 13
rect 18 -13 44 13
rect 80 -13 106 13
rect 142 -13 168 13
rect 204 -13 230 13
rect 266 -13 292 13
rect 328 -13 354 13
rect 390 -13 416 13
rect 452 -13 478 13
<< metal2 >>
rect -484 13 484 19
rect -484 -13 -478 13
rect -452 -13 -416 13
rect -390 -13 -354 13
rect -328 -13 -292 13
rect -266 -13 -230 13
rect -204 -13 -168 13
rect -142 -13 -106 13
rect -80 -13 -44 13
rect -18 -13 18 13
rect 44 -13 80 13
rect 106 -13 142 13
rect 168 -13 204 13
rect 230 -13 266 13
rect 292 -13 328 13
rect 354 -13 390 13
rect 416 -13 452 13
rect 478 -13 484 13
rect -484 -19 484 -13
<< end >>
