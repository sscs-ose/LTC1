magic
tech gf180mcuC
magscale 1 10
timestamp 1699891908
<< nwell >>
rect -320 2207 2313 2408
rect -320 2152 2310 2207
rect -320 -120 -120 2152
rect 2128 -120 2310 2152
rect -320 -320 2310 -120
<< nsubdiff >>
rect -270 2341 2260 2358
rect -270 2295 -253 2341
rect -207 2295 -155 2341
rect -109 2295 -57 2341
rect -11 2295 41 2341
rect 87 2295 139 2341
rect 185 2295 237 2341
rect 283 2295 335 2341
rect 381 2295 433 2341
rect 479 2295 531 2341
rect 577 2295 629 2341
rect 675 2295 727 2341
rect 773 2295 825 2341
rect 871 2295 923 2341
rect 969 2295 1021 2341
rect 1067 2295 1119 2341
rect 1165 2295 1217 2341
rect 1263 2295 1315 2341
rect 1361 2295 1413 2341
rect 1459 2295 1511 2341
rect 1557 2295 1609 2341
rect 1655 2295 1707 2341
rect 1753 2295 1805 2341
rect 1851 2295 1903 2341
rect 1949 2295 2001 2341
rect 2047 2295 2099 2341
rect 2145 2295 2197 2341
rect 2243 2295 2260 2341
rect -270 2278 2260 2295
rect -270 2243 -190 2278
rect -270 2197 -253 2243
rect -207 2197 -190 2243
rect -270 2145 -190 2197
rect -270 2099 -253 2145
rect -207 2099 -190 2145
rect -270 2047 -190 2099
rect -270 2001 -253 2047
rect -207 2001 -190 2047
rect -270 1949 -190 2001
rect -270 1903 -253 1949
rect -207 1903 -190 1949
rect -270 1851 -190 1903
rect -270 1805 -253 1851
rect -207 1805 -190 1851
rect -270 1753 -190 1805
rect -270 1707 -253 1753
rect -207 1707 -190 1753
rect -270 1655 -190 1707
rect -270 1609 -253 1655
rect -207 1609 -190 1655
rect -270 1557 -190 1609
rect -270 1511 -253 1557
rect -207 1511 -190 1557
rect -270 1459 -190 1511
rect -270 1413 -253 1459
rect -207 1413 -190 1459
rect -270 1361 -190 1413
rect -270 1315 -253 1361
rect -207 1315 -190 1361
rect -270 1263 -190 1315
rect -270 1217 -253 1263
rect -207 1217 -190 1263
rect -270 1165 -190 1217
rect -270 1119 -253 1165
rect -207 1119 -190 1165
rect -270 1067 -190 1119
rect -270 1021 -253 1067
rect -207 1021 -190 1067
rect -270 969 -190 1021
rect -270 923 -253 969
rect -207 923 -190 969
rect -270 871 -190 923
rect -270 825 -253 871
rect -207 825 -190 871
rect -270 773 -190 825
rect -270 727 -253 773
rect -207 727 -190 773
rect -270 675 -190 727
rect -270 629 -253 675
rect -207 629 -190 675
rect -270 577 -190 629
rect -270 531 -253 577
rect -207 531 -190 577
rect -270 479 -190 531
rect -270 433 -253 479
rect -207 433 -190 479
rect -270 381 -190 433
rect -270 335 -253 381
rect -207 335 -190 381
rect -270 283 -190 335
rect -270 237 -253 283
rect -207 237 -190 283
rect -270 185 -190 237
rect -270 139 -253 185
rect -207 139 -190 185
rect -270 87 -190 139
rect -270 41 -253 87
rect -207 41 -190 87
rect -270 -11 -190 41
rect -270 -57 -253 -11
rect -207 -57 -190 -11
rect -270 -109 -190 -57
rect -270 -155 -253 -109
rect -207 -155 -190 -109
rect -270 -190 -190 -155
rect 2180 2243 2260 2278
rect 2180 2197 2197 2243
rect 2243 2197 2260 2243
rect 2180 2145 2260 2197
rect 2180 2099 2197 2145
rect 2243 2099 2260 2145
rect 2180 2047 2260 2099
rect 2180 2001 2197 2047
rect 2243 2001 2260 2047
rect 2180 1949 2260 2001
rect 2180 1903 2197 1949
rect 2243 1903 2260 1949
rect 2180 1851 2260 1903
rect 2180 1805 2197 1851
rect 2243 1805 2260 1851
rect 2180 1753 2260 1805
rect 2180 1707 2197 1753
rect 2243 1707 2260 1753
rect 2180 1655 2260 1707
rect 2180 1609 2197 1655
rect 2243 1609 2260 1655
rect 2180 1557 2260 1609
rect 2180 1511 2197 1557
rect 2243 1511 2260 1557
rect 2180 1459 2260 1511
rect 2180 1413 2197 1459
rect 2243 1413 2260 1459
rect 2180 1361 2260 1413
rect 2180 1315 2197 1361
rect 2243 1315 2260 1361
rect 2180 1263 2260 1315
rect 2180 1217 2197 1263
rect 2243 1217 2260 1263
rect 2180 1165 2260 1217
rect 2180 1119 2197 1165
rect 2243 1119 2260 1165
rect 2180 1067 2260 1119
rect 2180 1021 2197 1067
rect 2243 1021 2260 1067
rect 2180 969 2260 1021
rect 2180 923 2197 969
rect 2243 923 2260 969
rect 2180 871 2260 923
rect 2180 825 2197 871
rect 2243 825 2260 871
rect 2180 773 2260 825
rect 2180 727 2197 773
rect 2243 727 2260 773
rect 2180 675 2260 727
rect 2180 629 2197 675
rect 2243 629 2260 675
rect 2180 577 2260 629
rect 2180 531 2197 577
rect 2243 531 2260 577
rect 2180 479 2260 531
rect 2180 433 2197 479
rect 2243 433 2260 479
rect 2180 381 2260 433
rect 2180 335 2197 381
rect 2243 335 2260 381
rect 2180 283 2260 335
rect 2180 237 2197 283
rect 2243 237 2260 283
rect 2180 185 2260 237
rect 2180 139 2197 185
rect 2243 139 2260 185
rect 2180 87 2260 139
rect 2180 41 2197 87
rect 2243 41 2260 87
rect 2180 -11 2260 41
rect 2180 -57 2197 -11
rect 2243 -57 2260 -11
rect 2180 -109 2260 -57
rect 2180 -155 2197 -109
rect 2243 -155 2260 -109
rect 2180 -190 2260 -155
rect -270 -207 2260 -190
rect -270 -253 -253 -207
rect -207 -253 -155 -207
rect -109 -253 -57 -207
rect -11 -253 41 -207
rect 87 -253 139 -207
rect 185 -253 237 -207
rect 283 -253 335 -207
rect 381 -253 433 -207
rect 479 -253 531 -207
rect 577 -253 629 -207
rect 675 -253 727 -207
rect 773 -253 825 -207
rect 871 -253 923 -207
rect 969 -253 1021 -207
rect 1067 -253 1119 -207
rect 1165 -253 1217 -207
rect 1263 -253 1315 -207
rect 1361 -253 1413 -207
rect 1459 -253 1511 -207
rect 1557 -253 1609 -207
rect 1655 -253 1707 -207
rect 1753 -253 1805 -207
rect 1851 -253 1903 -207
rect 1949 -253 2001 -207
rect 2047 -253 2099 -207
rect 2145 -253 2197 -207
rect 2243 -253 2260 -207
rect -270 -270 2260 -253
<< nsubdiffcont >>
rect -253 2295 -207 2341
rect -155 2295 -109 2341
rect -57 2295 -11 2341
rect 41 2295 87 2341
rect 139 2295 185 2341
rect 237 2295 283 2341
rect 335 2295 381 2341
rect 433 2295 479 2341
rect 531 2295 577 2341
rect 629 2295 675 2341
rect 727 2295 773 2341
rect 825 2295 871 2341
rect 923 2295 969 2341
rect 1021 2295 1067 2341
rect 1119 2295 1165 2341
rect 1217 2295 1263 2341
rect 1315 2295 1361 2341
rect 1413 2295 1459 2341
rect 1511 2295 1557 2341
rect 1609 2295 1655 2341
rect 1707 2295 1753 2341
rect 1805 2295 1851 2341
rect 1903 2295 1949 2341
rect 2001 2295 2047 2341
rect 2099 2295 2145 2341
rect 2197 2295 2243 2341
rect -253 2197 -207 2243
rect -253 2099 -207 2145
rect -253 2001 -207 2047
rect -253 1903 -207 1949
rect -253 1805 -207 1851
rect -253 1707 -207 1753
rect -253 1609 -207 1655
rect -253 1511 -207 1557
rect -253 1413 -207 1459
rect -253 1315 -207 1361
rect -253 1217 -207 1263
rect -253 1119 -207 1165
rect -253 1021 -207 1067
rect -253 923 -207 969
rect -253 825 -207 871
rect -253 727 -207 773
rect -253 629 -207 675
rect -253 531 -207 577
rect -253 433 -207 479
rect -253 335 -207 381
rect -253 237 -207 283
rect -253 139 -207 185
rect -253 41 -207 87
rect -253 -57 -207 -11
rect -253 -155 -207 -109
rect 2197 2197 2243 2243
rect 2197 2099 2243 2145
rect 2197 2001 2243 2047
rect 2197 1903 2243 1949
rect 2197 1805 2243 1851
rect 2197 1707 2243 1753
rect 2197 1609 2243 1655
rect 2197 1511 2243 1557
rect 2197 1413 2243 1459
rect 2197 1315 2243 1361
rect 2197 1217 2243 1263
rect 2197 1119 2243 1165
rect 2197 1021 2243 1067
rect 2197 923 2243 969
rect 2197 825 2243 871
rect 2197 727 2243 773
rect 2197 629 2243 675
rect 2197 531 2243 577
rect 2197 433 2243 479
rect 2197 335 2243 381
rect 2197 237 2243 283
rect 2197 139 2243 185
rect 2197 41 2243 87
rect 2197 -57 2243 -11
rect 2197 -155 2243 -109
rect -253 -253 -207 -207
rect -155 -253 -109 -207
rect -57 -253 -11 -207
rect 41 -253 87 -207
rect 139 -253 185 -207
rect 237 -253 283 -207
rect 335 -253 381 -207
rect 433 -253 479 -207
rect 531 -253 577 -207
rect 629 -253 675 -207
rect 727 -253 773 -207
rect 825 -253 871 -207
rect 923 -253 969 -207
rect 1021 -253 1067 -207
rect 1119 -253 1165 -207
rect 1217 -253 1263 -207
rect 1315 -253 1361 -207
rect 1413 -253 1459 -207
rect 1511 -253 1557 -207
rect 1609 -253 1655 -207
rect 1707 -253 1753 -207
rect 1805 -253 1851 -207
rect 1903 -253 1949 -207
rect 2001 -253 2047 -207
rect 2099 -253 2145 -207
rect 2197 -253 2243 -207
<< metal1 >>
rect -270 2341 2260 2358
rect -270 2295 -253 2341
rect -207 2295 -155 2341
rect -109 2295 -57 2341
rect -11 2295 41 2341
rect 87 2295 139 2341
rect 185 2295 237 2341
rect 283 2295 335 2341
rect 381 2295 433 2341
rect 479 2295 531 2341
rect 577 2295 629 2341
rect 675 2295 727 2341
rect 773 2295 825 2341
rect 871 2295 923 2341
rect 969 2295 1021 2341
rect 1067 2295 1119 2341
rect 1165 2295 1217 2341
rect 1263 2295 1315 2341
rect 1361 2295 1413 2341
rect 1459 2295 1511 2341
rect 1557 2295 1609 2341
rect 1655 2295 1707 2341
rect 1753 2295 1805 2341
rect 1851 2295 1903 2341
rect 1949 2295 2001 2341
rect 2047 2295 2099 2341
rect 2145 2295 2197 2341
rect 2243 2295 2260 2341
rect -270 2278 2260 2295
rect -270 2243 -190 2278
rect -270 2197 -253 2243
rect -207 2197 -190 2243
rect -270 2145 -190 2197
rect -270 2099 -253 2145
rect -207 2099 -190 2145
rect -270 2047 -190 2099
rect -270 2001 -253 2047
rect -207 2001 -190 2047
rect -270 1949 -190 2001
rect -270 1903 -253 1949
rect -207 1903 -190 1949
rect 67 1911 260 2278
rect 345 2052 542 2278
rect 345 1908 544 2052
rect 905 2023 1662 2152
rect -270 1851 -190 1903
rect -270 1805 -253 1851
rect -207 1805 -190 1851
rect 627 1840 823 1954
rect 906 1909 1102 2023
rect 1187 1840 1383 1954
rect 1466 1909 1662 2023
rect 1745 1906 1938 2278
rect 2180 2243 2260 2278
rect 2180 2197 2197 2243
rect 2243 2197 2260 2243
rect 2180 2145 2260 2197
rect 2180 2099 2197 2145
rect 2243 2099 2260 2145
rect 2180 2047 2260 2099
rect 2180 2001 2197 2047
rect 2243 2001 2260 2047
rect 2180 1949 2260 2001
rect -270 1753 -190 1805
rect -270 1707 -253 1753
rect -207 1707 -190 1753
rect -270 1655 -190 1707
rect -270 1609 -253 1655
rect -207 1609 -190 1655
rect -270 1557 -190 1609
rect 626 1599 1383 1840
rect 2180 1903 2197 1949
rect 2243 1903 2260 1949
rect 2180 1851 2260 1903
rect 2180 1805 2197 1851
rect 2243 1805 2260 1851
rect 2180 1753 2260 1805
rect 2180 1707 2197 1753
rect 2243 1707 2260 1753
rect 2180 1655 2260 1707
rect 2180 1609 2197 1655
rect 2243 1609 2260 1655
rect -270 1511 -253 1557
rect -207 1511 -190 1557
rect -270 1459 -190 1511
rect -270 1413 -253 1459
rect -207 1413 -190 1459
rect -270 1361 -190 1413
rect -270 1315 -253 1361
rect -207 1315 -190 1361
rect -270 1263 -190 1315
rect -270 1217 -253 1263
rect -207 1217 -190 1263
rect -270 1165 -190 1217
rect -270 1119 -253 1165
rect -207 1119 -190 1165
rect -270 1067 -190 1119
rect -270 1021 -253 1067
rect -207 1021 -190 1067
rect -270 969 -190 1021
rect -270 923 -253 969
rect -207 923 -190 969
rect -270 871 -190 923
rect -270 825 -253 871
rect -207 825 -190 871
rect -270 773 -190 825
rect -270 727 -253 773
rect -207 727 -190 773
rect -270 675 -190 727
rect -270 629 -253 675
rect -207 629 -190 675
rect -270 577 -190 629
rect -270 531 -253 577
rect -207 531 -190 577
rect -270 479 -190 531
rect -270 433 -253 479
rect -207 433 -190 479
rect -270 381 -190 433
rect 2180 1557 2260 1609
rect 2180 1511 2197 1557
rect 2243 1511 2260 1557
rect 2180 1459 2260 1511
rect 2180 1413 2197 1459
rect 2243 1413 2260 1459
rect 2180 1361 2260 1413
rect 2180 1315 2197 1361
rect 2243 1315 2260 1361
rect 2180 1263 2260 1315
rect 2180 1217 2197 1263
rect 2243 1217 2260 1263
rect 2180 1165 2260 1217
rect 2180 1119 2197 1165
rect 2243 1119 2260 1165
rect 2180 1067 2260 1119
rect 2180 1021 2197 1067
rect 2243 1021 2260 1067
rect 2180 969 2260 1021
rect 2180 923 2197 969
rect 2243 923 2260 969
rect 2180 871 2260 923
rect 2180 825 2197 871
rect 2243 825 2260 871
rect 2180 773 2260 825
rect 2180 727 2197 773
rect 2243 727 2260 773
rect 2180 675 2260 727
rect 2180 629 2197 675
rect 2243 629 2260 675
rect 2180 577 2260 629
rect 2180 531 2197 577
rect 2243 531 2260 577
rect 2180 479 2260 531
rect 2180 433 2197 479
rect 2243 433 2260 479
rect -270 335 -253 381
rect -207 335 -190 381
rect -270 283 -190 335
rect -270 237 -253 283
rect -207 237 -190 283
rect -270 185 -190 237
rect 175 191 822 423
rect -270 139 -253 185
rect -207 139 -190 185
rect -270 87 -190 139
rect -270 41 -253 87
rect -207 41 -190 87
rect -270 -11 -190 41
rect -270 -57 -253 -11
rect -207 -57 -190 -11
rect -270 -109 -190 -57
rect -270 -155 -253 -109
rect -207 -155 -190 -109
rect -270 -190 -190 -155
rect 68 -190 261 134
rect 346 9 542 123
rect 626 77 822 191
rect 2180 381 2260 433
rect 2180 335 2197 381
rect 2243 335 2260 381
rect 2180 283 2260 335
rect 2180 237 2197 283
rect 2243 237 2260 283
rect 2180 185 2260 237
rect 2180 139 2197 185
rect 2243 139 2260 185
rect 908 9 1104 123
rect 345 -120 1104 9
rect 1186 9 1382 123
rect 1465 9 1661 123
rect 1186 -120 1661 9
rect 1745 -190 1938 139
rect 2180 87 2260 139
rect 2180 41 2197 87
rect 2243 41 2260 87
rect 2180 -11 2260 41
rect 2180 -57 2197 -11
rect 2243 -57 2260 -11
rect 2180 -109 2260 -57
rect 2180 -155 2197 -109
rect 2243 -155 2260 -109
rect 2180 -190 2260 -155
rect -270 -207 2260 -190
rect -270 -253 -253 -207
rect -207 -253 -155 -207
rect -109 -253 -57 -207
rect -11 -253 41 -207
rect 87 -253 139 -207
rect 185 -253 237 -207
rect 283 -253 335 -207
rect 381 -253 433 -207
rect 479 -253 531 -207
rect 577 -253 629 -207
rect 675 -253 727 -207
rect 773 -253 825 -207
rect 871 -253 923 -207
rect 969 -253 1021 -207
rect 1067 -253 1119 -207
rect 1165 -253 1217 -207
rect 1263 -253 1315 -207
rect 1361 -253 1413 -207
rect 1459 -253 1511 -207
rect 1557 -253 1609 -207
rect 1655 -253 1707 -207
rect 1753 -253 1805 -207
rect 1851 -253 1903 -207
rect 1949 -253 2001 -207
rect 2047 -253 2099 -207
rect 2145 -253 2197 -207
rect 2243 -253 2260 -207
rect -270 -270 2260 -253
use ppolyf_u_3VY3SR  ppolyf_u_3VY3SR_0
timestamp 1699882188
transform 1 0 1004 0 1 1016
box -1124 -1136 1124 1136
<< labels >>
flabel metal1 418 2323 418 2323 0 FreeSans 1600 0 0 0 VDD
port 0 nsew
flabel metal1 301 267 301 267 0 FreeSans 1600 0 0 0 VSS
port 1 nsew
flabel metal1 1414 -11 1414 -11 0 FreeSans 800 0 0 0 VCM_1.3
port 4 nsew
<< end >>
