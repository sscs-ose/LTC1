magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1484 -1081 1484 1081
<< metal1 >>
rect -484 75 484 81
rect -484 49 -478 75
rect -452 49 -416 75
rect -390 49 -354 75
rect -328 49 -292 75
rect -266 49 -230 75
rect -204 49 -168 75
rect -142 49 -106 75
rect -80 49 -44 75
rect -18 49 18 75
rect 44 49 80 75
rect 106 49 142 75
rect 168 49 204 75
rect 230 49 266 75
rect 292 49 328 75
rect 354 49 390 75
rect 416 49 452 75
rect 478 49 484 75
rect -484 13 484 49
rect -484 -13 -478 13
rect -452 -13 -416 13
rect -390 -13 -354 13
rect -328 -13 -292 13
rect -266 -13 -230 13
rect -204 -13 -168 13
rect -142 -13 -106 13
rect -80 -13 -44 13
rect -18 -13 18 13
rect 44 -13 80 13
rect 106 -13 142 13
rect 168 -13 204 13
rect 230 -13 266 13
rect 292 -13 328 13
rect 354 -13 390 13
rect 416 -13 452 13
rect 478 -13 484 13
rect -484 -49 484 -13
rect -484 -75 -478 -49
rect -452 -75 -416 -49
rect -390 -75 -354 -49
rect -328 -75 -292 -49
rect -266 -75 -230 -49
rect -204 -75 -168 -49
rect -142 -75 -106 -49
rect -80 -75 -44 -49
rect -18 -75 18 -49
rect 44 -75 80 -49
rect 106 -75 142 -49
rect 168 -75 204 -49
rect 230 -75 266 -49
rect 292 -75 328 -49
rect 354 -75 390 -49
rect 416 -75 452 -49
rect 478 -75 484 -49
rect -484 -81 484 -75
<< via1 >>
rect -478 49 -452 75
rect -416 49 -390 75
rect -354 49 -328 75
rect -292 49 -266 75
rect -230 49 -204 75
rect -168 49 -142 75
rect -106 49 -80 75
rect -44 49 -18 75
rect 18 49 44 75
rect 80 49 106 75
rect 142 49 168 75
rect 204 49 230 75
rect 266 49 292 75
rect 328 49 354 75
rect 390 49 416 75
rect 452 49 478 75
rect -478 -13 -452 13
rect -416 -13 -390 13
rect -354 -13 -328 13
rect -292 -13 -266 13
rect -230 -13 -204 13
rect -168 -13 -142 13
rect -106 -13 -80 13
rect -44 -13 -18 13
rect 18 -13 44 13
rect 80 -13 106 13
rect 142 -13 168 13
rect 204 -13 230 13
rect 266 -13 292 13
rect 328 -13 354 13
rect 390 -13 416 13
rect 452 -13 478 13
rect -478 -75 -452 -49
rect -416 -75 -390 -49
rect -354 -75 -328 -49
rect -292 -75 -266 -49
rect -230 -75 -204 -49
rect -168 -75 -142 -49
rect -106 -75 -80 -49
rect -44 -75 -18 -49
rect 18 -75 44 -49
rect 80 -75 106 -49
rect 142 -75 168 -49
rect 204 -75 230 -49
rect 266 -75 292 -49
rect 328 -75 354 -49
rect 390 -75 416 -49
rect 452 -75 478 -49
<< metal2 >>
rect -484 75 484 81
rect -484 49 -478 75
rect -452 49 -416 75
rect -390 49 -354 75
rect -328 49 -292 75
rect -266 49 -230 75
rect -204 49 -168 75
rect -142 49 -106 75
rect -80 49 -44 75
rect -18 49 18 75
rect 44 49 80 75
rect 106 49 142 75
rect 168 49 204 75
rect 230 49 266 75
rect 292 49 328 75
rect 354 49 390 75
rect 416 49 452 75
rect 478 49 484 75
rect -484 13 484 49
rect -484 -13 -478 13
rect -452 -13 -416 13
rect -390 -13 -354 13
rect -328 -13 -292 13
rect -266 -13 -230 13
rect -204 -13 -168 13
rect -142 -13 -106 13
rect -80 -13 -44 13
rect -18 -13 18 13
rect 44 -13 80 13
rect 106 -13 142 13
rect 168 -13 204 13
rect 230 -13 266 13
rect 292 -13 328 13
rect 354 -13 390 13
rect 416 -13 452 13
rect 478 -13 484 13
rect -484 -49 484 -13
rect -484 -75 -478 -49
rect -452 -75 -416 -49
rect -390 -75 -354 -49
rect -328 -75 -292 -49
rect -266 -75 -230 -49
rect -204 -75 -168 -49
rect -142 -75 -106 -49
rect -80 -75 -44 -49
rect -18 -75 18 -49
rect 44 -75 80 -49
rect 106 -75 142 -49
rect 168 -75 204 -49
rect 230 -75 266 -49
rect 292 -75 328 -49
rect 354 -75 390 -49
rect 416 -75 452 -49
rect 478 -75 484 -49
rect -484 -81 484 -75
<< end >>
