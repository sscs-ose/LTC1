magic
tech gf180mcuC
magscale 1 10
timestamp 1692016228
<< nwell >>
rect 0 277 884 868
<< pwell >>
rect 222 0 662 236
<< nmos >>
rect 334 68 390 168
rect 494 68 550 168
<< pmos >>
rect 174 407 230 607
rect 334 407 390 607
rect 494 407 550 607
rect 654 407 710 607
<< ndiff >>
rect 246 155 334 168
rect 246 81 259 155
rect 305 81 334 155
rect 246 68 334 81
rect 390 155 494 168
rect 390 81 419 155
rect 465 81 494 155
rect 390 68 494 81
rect 550 155 638 168
rect 550 81 579 155
rect 625 81 638 155
rect 550 68 638 81
<< pdiff >>
rect 86 594 174 607
rect 86 420 99 594
rect 145 420 174 594
rect 86 407 174 420
rect 230 594 334 607
rect 230 420 259 594
rect 305 420 334 594
rect 230 407 334 420
rect 390 594 494 607
rect 390 420 419 594
rect 465 420 494 594
rect 390 407 494 420
rect 550 594 654 607
rect 550 420 579 594
rect 625 420 654 594
rect 550 407 654 420
rect 710 594 798 607
rect 710 420 739 594
rect 785 420 798 594
rect 710 407 798 420
<< ndiffc >>
rect 259 81 305 155
rect 419 81 465 155
rect 579 81 625 155
<< pdiffc >>
rect 99 420 145 594
rect 259 420 305 594
rect 419 420 465 594
rect 579 420 625 594
rect 739 420 785 594
<< psubdiff >>
rect 265 -33 619 -20
rect 265 -79 278 -33
rect 324 -79 372 -33
rect 418 -79 466 -33
rect 512 -79 560 -33
rect 606 -79 619 -33
rect 265 -92 619 -79
<< nsubdiff >>
rect 30 822 854 835
rect 30 776 43 822
rect 89 776 137 822
rect 183 776 231 822
rect 277 776 325 822
rect 371 776 419 822
rect 465 776 513 822
rect 559 776 607 822
rect 653 776 701 822
rect 747 776 795 822
rect 841 776 854 822
rect 30 763 854 776
<< psubdiffcont >>
rect 278 -79 324 -33
rect 372 -79 418 -33
rect 466 -79 512 -33
rect 560 -79 606 -33
<< nsubdiffcont >>
rect 43 776 89 822
rect 137 776 183 822
rect 231 776 277 822
rect 325 776 371 822
rect 419 776 465 822
rect 513 776 559 822
rect 607 776 653 822
rect 701 776 747 822
rect 795 776 841 822
<< polysilicon >>
rect 174 607 230 651
rect 334 607 390 651
rect 494 607 550 651
rect 654 607 710 651
rect 174 268 230 407
rect 155 260 230 268
rect 334 260 390 407
rect 155 255 390 260
rect 155 209 168 255
rect 214 209 390 255
rect 155 204 390 209
rect 155 196 227 204
rect 334 168 390 204
rect 494 343 550 407
rect 654 343 710 407
rect 494 287 714 343
rect 494 168 550 287
rect 658 230 714 287
rect 762 230 834 238
rect 658 225 834 230
rect 658 178 775 225
rect 821 178 834 225
rect 658 174 834 178
rect 762 165 834 174
rect 334 24 390 68
rect 494 24 550 68
<< polycontact >>
rect 168 209 214 255
rect 775 178 821 225
<< metal1 >>
rect 0 822 884 855
rect 0 776 43 822
rect 89 776 137 822
rect 183 776 231 822
rect 277 776 325 822
rect 371 776 419 822
rect 465 776 513 822
rect 559 776 607 822
rect 653 776 701 822
rect 747 776 795 822
rect 841 776 884 822
rect 0 743 884 776
rect 99 594 145 605
rect 99 363 145 420
rect 259 594 305 743
rect 259 409 305 420
rect 419 651 785 697
rect 419 594 465 651
rect 419 363 465 420
rect 99 317 465 363
rect 579 594 625 605
rect 579 363 625 420
rect 739 594 785 651
rect 739 409 785 420
rect 579 317 713 363
rect 157 255 225 266
rect 579 258 625 317
rect 113 209 168 255
rect 214 209 225 255
rect 157 198 225 209
rect 419 212 625 258
rect 764 225 832 236
rect 259 155 305 166
rect 259 0 305 81
rect 419 155 465 212
rect 764 178 775 225
rect 821 178 902 225
rect 764 167 832 178
rect 419 70 465 81
rect 579 155 625 166
rect 579 0 625 81
rect 222 -33 662 0
rect 222 -79 278 -33
rect 324 -79 372 -33
rect 418 -79 466 -33
rect 512 -79 560 -33
rect 606 -79 662 -33
rect 222 -112 662 -79
<< labels >>
flabel metal1 437 -56 437 -56 0 FreeSans 320 0 0 0 VSS
port 7 nsew
flabel nsubdiffcont 442 799 442 799 0 FreeSans 320 0 0 0 VDD
port 6 nsew
flabel metal1 123 232 123 232 0 FreeSans 320 0 0 0 A
port 0 nsew
flabel metal1 888 202 888 202 0 FreeSans 320 0 0 0 B
port 1 nsew
flabel metal1 681 340 681 340 0 FreeSans 320 0 0 0 OUT
port 4 nsew
<< end >>
