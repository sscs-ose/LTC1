magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1949 1019 1949
<< metal2 >>
rect -19 944 19 949
rect -19 916 -14 944
rect 14 916 19 944
rect -19 882 19 916
rect -19 854 -14 882
rect 14 854 19 882
rect -19 820 19 854
rect -19 792 -14 820
rect 14 792 19 820
rect -19 758 19 792
rect -19 730 -14 758
rect 14 730 19 758
rect -19 696 19 730
rect -19 668 -14 696
rect 14 668 19 696
rect -19 634 19 668
rect -19 606 -14 634
rect 14 606 19 634
rect -19 572 19 606
rect -19 544 -14 572
rect 14 544 19 572
rect -19 510 19 544
rect -19 482 -14 510
rect 14 482 19 510
rect -19 448 19 482
rect -19 420 -14 448
rect 14 420 19 448
rect -19 386 19 420
rect -19 358 -14 386
rect 14 358 19 386
rect -19 324 19 358
rect -19 296 -14 324
rect 14 296 19 324
rect -19 262 19 296
rect -19 234 -14 262
rect 14 234 19 262
rect -19 200 19 234
rect -19 172 -14 200
rect 14 172 19 200
rect -19 138 19 172
rect -19 110 -14 138
rect 14 110 19 138
rect -19 76 19 110
rect -19 48 -14 76
rect 14 48 19 76
rect -19 14 19 48
rect -19 -14 -14 14
rect 14 -14 19 14
rect -19 -48 19 -14
rect -19 -76 -14 -48
rect 14 -76 19 -48
rect -19 -110 19 -76
rect -19 -138 -14 -110
rect 14 -138 19 -110
rect -19 -172 19 -138
rect -19 -200 -14 -172
rect 14 -200 19 -172
rect -19 -234 19 -200
rect -19 -262 -14 -234
rect 14 -262 19 -234
rect -19 -296 19 -262
rect -19 -324 -14 -296
rect 14 -324 19 -296
rect -19 -358 19 -324
rect -19 -386 -14 -358
rect 14 -386 19 -358
rect -19 -420 19 -386
rect -19 -448 -14 -420
rect 14 -448 19 -420
rect -19 -482 19 -448
rect -19 -510 -14 -482
rect 14 -510 19 -482
rect -19 -544 19 -510
rect -19 -572 -14 -544
rect 14 -572 19 -544
rect -19 -606 19 -572
rect -19 -634 -14 -606
rect 14 -634 19 -606
rect -19 -668 19 -634
rect -19 -696 -14 -668
rect 14 -696 19 -668
rect -19 -730 19 -696
rect -19 -758 -14 -730
rect 14 -758 19 -730
rect -19 -792 19 -758
rect -19 -820 -14 -792
rect 14 -820 19 -792
rect -19 -854 19 -820
rect -19 -882 -14 -854
rect 14 -882 19 -854
rect -19 -916 19 -882
rect -19 -944 -14 -916
rect 14 -944 19 -916
rect -19 -949 19 -944
<< via2 >>
rect -14 916 14 944
rect -14 854 14 882
rect -14 792 14 820
rect -14 730 14 758
rect -14 668 14 696
rect -14 606 14 634
rect -14 544 14 572
rect -14 482 14 510
rect -14 420 14 448
rect -14 358 14 386
rect -14 296 14 324
rect -14 234 14 262
rect -14 172 14 200
rect -14 110 14 138
rect -14 48 14 76
rect -14 -14 14 14
rect -14 -76 14 -48
rect -14 -138 14 -110
rect -14 -200 14 -172
rect -14 -262 14 -234
rect -14 -324 14 -296
rect -14 -386 14 -358
rect -14 -448 14 -420
rect -14 -510 14 -482
rect -14 -572 14 -544
rect -14 -634 14 -606
rect -14 -696 14 -668
rect -14 -758 14 -730
rect -14 -820 14 -792
rect -14 -882 14 -854
rect -14 -944 14 -916
<< metal3 >>
rect -19 944 19 949
rect -19 916 -14 944
rect 14 916 19 944
rect -19 882 19 916
rect -19 854 -14 882
rect 14 854 19 882
rect -19 820 19 854
rect -19 792 -14 820
rect 14 792 19 820
rect -19 758 19 792
rect -19 730 -14 758
rect 14 730 19 758
rect -19 696 19 730
rect -19 668 -14 696
rect 14 668 19 696
rect -19 634 19 668
rect -19 606 -14 634
rect 14 606 19 634
rect -19 572 19 606
rect -19 544 -14 572
rect 14 544 19 572
rect -19 510 19 544
rect -19 482 -14 510
rect 14 482 19 510
rect -19 448 19 482
rect -19 420 -14 448
rect 14 420 19 448
rect -19 386 19 420
rect -19 358 -14 386
rect 14 358 19 386
rect -19 324 19 358
rect -19 296 -14 324
rect 14 296 19 324
rect -19 262 19 296
rect -19 234 -14 262
rect 14 234 19 262
rect -19 200 19 234
rect -19 172 -14 200
rect 14 172 19 200
rect -19 138 19 172
rect -19 110 -14 138
rect 14 110 19 138
rect -19 76 19 110
rect -19 48 -14 76
rect 14 48 19 76
rect -19 14 19 48
rect -19 -14 -14 14
rect 14 -14 19 14
rect -19 -48 19 -14
rect -19 -76 -14 -48
rect 14 -76 19 -48
rect -19 -110 19 -76
rect -19 -138 -14 -110
rect 14 -138 19 -110
rect -19 -172 19 -138
rect -19 -200 -14 -172
rect 14 -200 19 -172
rect -19 -234 19 -200
rect -19 -262 -14 -234
rect 14 -262 19 -234
rect -19 -296 19 -262
rect -19 -324 -14 -296
rect 14 -324 19 -296
rect -19 -358 19 -324
rect -19 -386 -14 -358
rect 14 -386 19 -358
rect -19 -420 19 -386
rect -19 -448 -14 -420
rect 14 -448 19 -420
rect -19 -482 19 -448
rect -19 -510 -14 -482
rect 14 -510 19 -482
rect -19 -544 19 -510
rect -19 -572 -14 -544
rect 14 -572 19 -544
rect -19 -606 19 -572
rect -19 -634 -14 -606
rect 14 -634 19 -606
rect -19 -668 19 -634
rect -19 -696 -14 -668
rect 14 -696 19 -668
rect -19 -730 19 -696
rect -19 -758 -14 -730
rect 14 -758 19 -730
rect -19 -792 19 -758
rect -19 -820 -14 -792
rect 14 -820 19 -792
rect -19 -854 19 -820
rect -19 -882 -14 -854
rect 14 -882 19 -854
rect -19 -916 19 -882
rect -19 -944 -14 -916
rect 14 -944 19 -916
rect -19 -949 19 -944
<< end >>
