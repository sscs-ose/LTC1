magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -70140 -70970 8839 10429
<< metal1 >>
rect -52012 8302 -51027 8429
rect -52012 8286 -51676 8302
rect -52012 8234 -51864 8286
rect -51812 8250 -51676 8286
rect -51624 8250 -51027 8302
rect -51812 8234 -51027 8250
rect -52012 8151 -51027 8234
rect -65244 7981 -64259 8149
rect -65244 7965 -64933 7981
rect -65244 7913 -65121 7965
rect -65069 7929 -64933 7965
rect -64881 7929 -64259 7981
rect -65069 7913 -64259 7929
rect -65244 7830 -64259 7913
rect -65244 7796 -64670 7830
rect -65244 7788 -64904 7796
rect -65244 7736 -65105 7788
rect -65053 7744 -64904 7788
rect -64852 7778 -64670 7796
rect -64618 7778 -64259 7830
rect -64852 7768 -64259 7778
rect -64852 7744 -64483 7768
rect -65053 7736 -64483 7744
rect -65244 7716 -64483 7736
rect -64431 7716 -64259 7768
rect -65244 7620 -64259 7716
rect -65244 7607 -64887 7620
rect -65244 7555 -65101 7607
rect -65049 7568 -64887 7607
rect -64835 7611 -64259 7620
rect -64835 7568 -64670 7611
rect -65049 7559 -64670 7568
rect -64618 7583 -64259 7611
rect -64618 7559 -64440 7583
rect -65049 7555 -64440 7559
rect -65244 7531 -64440 7555
rect -64388 7531 -64259 7583
rect -65244 7163 -64259 7531
rect -65244 7147 -64956 7163
rect -65244 7095 -65144 7147
rect -65092 7111 -64956 7147
rect -64904 7111 -64259 7163
rect -65092 7095 -64259 7111
rect -65244 7012 -64259 7095
rect -65244 6978 -64693 7012
rect -65244 6970 -64927 6978
rect -65244 6918 -65128 6970
rect -65076 6926 -64927 6970
rect -64875 6960 -64693 6978
rect -64641 6960 -64259 7012
rect -64875 6950 -64259 6960
rect -64875 6926 -64506 6950
rect -65076 6918 -64506 6926
rect -65244 6898 -64506 6918
rect -64454 6898 -64259 6950
rect -65244 6802 -64259 6898
rect -65244 6789 -64910 6802
rect -65244 6737 -65124 6789
rect -65072 6750 -64910 6789
rect -64858 6793 -64259 6802
rect -64858 6750 -64693 6793
rect -65072 6741 -64693 6750
rect -64641 6765 -64259 6793
rect -64641 6741 -64463 6765
rect -65072 6737 -64463 6741
rect -65244 6713 -64463 6737
rect -64411 6713 -64259 6765
rect -65244 6454 -64259 6713
rect -59062 8063 -58077 8149
rect -59062 8047 -58738 8063
rect -59062 7995 -58926 8047
rect -58874 8011 -58738 8047
rect -58686 8011 -58077 8063
rect -58874 7995 -58077 8011
rect -59062 7912 -58077 7995
rect -59062 7878 -58475 7912
rect -59062 7870 -58709 7878
rect -59062 7818 -58910 7870
rect -58858 7826 -58709 7870
rect -58657 7860 -58475 7878
rect -58423 7860 -58077 7912
rect -58657 7850 -58077 7860
rect -58657 7826 -58288 7850
rect -58858 7818 -58288 7826
rect -59062 7798 -58288 7818
rect -58236 7798 -58077 7850
rect -59062 7702 -58077 7798
rect -59062 7689 -58692 7702
rect -59062 7637 -58906 7689
rect -58854 7650 -58692 7689
rect -58640 7693 -58077 7702
rect -58640 7650 -58475 7693
rect -58854 7641 -58475 7650
rect -58423 7665 -58077 7693
rect -58423 7641 -58245 7665
rect -58854 7637 -58245 7641
rect -59062 7613 -58245 7637
rect -58193 7613 -58077 7665
rect -59062 7183 -58077 7613
rect -59062 7167 -58738 7183
rect -59062 7115 -58926 7167
rect -58874 7131 -58738 7167
rect -58686 7131 -58077 7183
rect -58874 7115 -58077 7131
rect -59062 7032 -58077 7115
rect -59062 6998 -58475 7032
rect -59062 6990 -58709 6998
rect -59062 6938 -58910 6990
rect -58858 6946 -58709 6990
rect -58657 6980 -58475 6998
rect -58423 6980 -58077 7032
rect -58657 6970 -58077 6980
rect -58657 6946 -58288 6970
rect -58858 6938 -58288 6946
rect -59062 6918 -58288 6938
rect -58236 6918 -58077 6970
rect -59062 6822 -58077 6918
rect -59062 6809 -58692 6822
rect -59062 6757 -58906 6809
rect -58854 6770 -58692 6809
rect -58640 6813 -58077 6822
rect -58640 6770 -58475 6813
rect -58854 6761 -58475 6770
rect -58423 6785 -58077 6813
rect -58423 6761 -58245 6785
rect -58854 6757 -58245 6761
rect -59062 6733 -58245 6757
rect -58193 6733 -58077 6785
rect -52012 8117 -51413 8151
rect -52012 8109 -51647 8117
rect -52012 8057 -51848 8109
rect -51796 8065 -51647 8109
rect -51595 8099 -51413 8117
rect -51361 8099 -51027 8151
rect -51595 8089 -51027 8099
rect -51595 8065 -51226 8089
rect -51796 8057 -51226 8065
rect -52012 8037 -51226 8057
rect -51174 8037 -51027 8089
rect -52012 7941 -51027 8037
rect -52012 7928 -51630 7941
rect -52012 7876 -51844 7928
rect -51792 7889 -51630 7928
rect -51578 7932 -51027 7941
rect -51578 7889 -51413 7932
rect -51792 7880 -51413 7889
rect -51361 7904 -51027 7932
rect -51361 7880 -51183 7904
rect -51792 7876 -51183 7880
rect -52012 7852 -51183 7876
rect -51131 7852 -51027 7904
rect -52012 7436 -51027 7852
rect -52012 7420 -51696 7436
rect -52012 7368 -51884 7420
rect -51832 7384 -51696 7420
rect -51644 7384 -51027 7436
rect -51832 7368 -51027 7384
rect -52012 7285 -51027 7368
rect -52012 7251 -51433 7285
rect -52012 7243 -51667 7251
rect -52012 7191 -51868 7243
rect -51816 7199 -51667 7243
rect -51615 7233 -51433 7251
rect -51381 7233 -51027 7285
rect -51615 7223 -51027 7233
rect -51615 7199 -51246 7223
rect -51816 7191 -51246 7199
rect -52012 7171 -51246 7191
rect -51194 7171 -51027 7223
rect -52012 7075 -51027 7171
rect -52012 7062 -51650 7075
rect -52012 7010 -51864 7062
rect -51812 7023 -51650 7062
rect -51598 7066 -51027 7075
rect -51598 7023 -51433 7066
rect -51812 7014 -51433 7023
rect -51381 7038 -51027 7066
rect -51381 7014 -51203 7038
rect -51812 7010 -51203 7014
rect -52012 6986 -51203 7010
rect -51151 6986 -51027 7038
rect -52012 6734 -51027 6986
rect -45475 8156 -44490 8254
rect -45475 8140 -45139 8156
rect -45475 8088 -45327 8140
rect -45275 8104 -45139 8140
rect -45087 8104 -44490 8156
rect -45275 8088 -44490 8104
rect -45475 8005 -44490 8088
rect -45475 7971 -44876 8005
rect -45475 7963 -45110 7971
rect -45475 7911 -45311 7963
rect -45259 7919 -45110 7963
rect -45058 7953 -44876 7971
rect -44824 7953 -44490 8005
rect -45058 7943 -44490 7953
rect -45058 7919 -44689 7943
rect -45259 7911 -44689 7919
rect -45475 7891 -44689 7911
rect -44637 7891 -44490 7943
rect -45475 7795 -44490 7891
rect -45475 7782 -45093 7795
rect -45475 7730 -45307 7782
rect -45255 7743 -45093 7782
rect -45041 7786 -44490 7795
rect -45041 7743 -44876 7786
rect -45255 7734 -44876 7743
rect -44824 7758 -44490 7786
rect -44824 7734 -44646 7758
rect -45255 7730 -44646 7734
rect -45475 7706 -44646 7730
rect -44594 7706 -44490 7758
rect -45475 7224 -44490 7706
rect -45475 7208 -45168 7224
rect -45475 7156 -45356 7208
rect -45304 7172 -45168 7208
rect -45116 7172 -44490 7224
rect -45304 7156 -44490 7172
rect -45475 7073 -44490 7156
rect -45475 7039 -44905 7073
rect -45475 7031 -45139 7039
rect -45475 6979 -45340 7031
rect -45288 6987 -45139 7031
rect -45087 7021 -44905 7039
rect -44853 7021 -44490 7073
rect -45087 7011 -44490 7021
rect -45087 6987 -44718 7011
rect -45288 6979 -44718 6987
rect -45475 6959 -44718 6979
rect -44666 6959 -44490 7011
rect -45475 6863 -44490 6959
rect -45475 6850 -45122 6863
rect -45475 6798 -45336 6850
rect -45284 6811 -45122 6850
rect -45070 6854 -44490 6863
rect -45070 6811 -44905 6854
rect -45284 6802 -44905 6811
rect -44853 6826 -44490 6854
rect -44853 6802 -44675 6826
rect -45284 6798 -44675 6802
rect -45475 6774 -44675 6798
rect -44623 6774 -44490 6826
rect -59062 6454 -58077 6733
rect -45475 6559 -44490 6774
rect -38757 8086 -37772 8237
rect -38757 8070 -38438 8086
rect -38757 8018 -38626 8070
rect -38574 8034 -38438 8070
rect -38386 8034 -37772 8086
rect -38574 8018 -37772 8034
rect -38757 7935 -37772 8018
rect -38757 7901 -38175 7935
rect -38757 7893 -38409 7901
rect -38757 7841 -38610 7893
rect -38558 7849 -38409 7893
rect -38357 7883 -38175 7901
rect -38123 7883 -37772 7935
rect -38357 7873 -37772 7883
rect -38357 7849 -37988 7873
rect -38558 7841 -37988 7849
rect -38757 7821 -37988 7841
rect -37936 7821 -37772 7873
rect -38757 7725 -37772 7821
rect -38757 7712 -38392 7725
rect -38757 7660 -38606 7712
rect -38554 7673 -38392 7712
rect -38340 7716 -37772 7725
rect -38340 7673 -38175 7716
rect -38554 7664 -38175 7673
rect -38123 7688 -37772 7716
rect -38123 7664 -37945 7688
rect -38554 7660 -37945 7664
rect -38757 7636 -37945 7660
rect -37893 7636 -37772 7688
rect -38757 7247 -37772 7636
rect -38757 7231 -38427 7247
rect -38757 7179 -38615 7231
rect -38563 7195 -38427 7231
rect -38375 7195 -37772 7247
rect -38563 7179 -37772 7195
rect -36350 7190 -33770 8380
rect -31724 8145 -30705 8360
rect -31724 8129 -31411 8145
rect -31724 8077 -31599 8129
rect -31547 8093 -31411 8129
rect -31359 8093 -30705 8145
rect -31547 8077 -30705 8093
rect -31724 7994 -30705 8077
rect -31724 7960 -31148 7994
rect -31724 7952 -31382 7960
rect -31724 7900 -31583 7952
rect -31531 7908 -31382 7952
rect -31330 7942 -31148 7960
rect -31096 7942 -30705 7994
rect -31330 7932 -30705 7942
rect -31330 7908 -30961 7932
rect -31531 7900 -30961 7908
rect -31724 7880 -30961 7900
rect -30909 7880 -30705 7932
rect -31724 7784 -30705 7880
rect -31724 7771 -31365 7784
rect -31724 7719 -31579 7771
rect -31527 7732 -31365 7771
rect -31313 7775 -30705 7784
rect -31313 7732 -31148 7775
rect -31527 7723 -31148 7732
rect -31096 7747 -30705 7775
rect -31096 7723 -30918 7747
rect -31527 7719 -30918 7723
rect -31724 7695 -30918 7719
rect -30866 7695 -30705 7747
rect -31724 7253 -30705 7695
rect -31724 7237 -31394 7253
rect -38757 7096 -37772 7179
rect -38757 7062 -38164 7096
rect -38757 7054 -38398 7062
rect -38757 7002 -38599 7054
rect -38547 7010 -38398 7054
rect -38346 7044 -38164 7062
rect -38112 7044 -37772 7096
rect -38346 7034 -37772 7044
rect -38346 7010 -37977 7034
rect -38547 7002 -37977 7010
rect -38757 6982 -37977 7002
rect -37925 6982 -37772 7034
rect -38757 6886 -37772 6982
rect -38757 6873 -38381 6886
rect -38757 6821 -38595 6873
rect -38543 6834 -38381 6873
rect -38329 6877 -37772 6886
rect -38329 6834 -38164 6877
rect -38543 6825 -38164 6834
rect -38112 6849 -37772 6877
rect -38112 6825 -37934 6849
rect -38543 6821 -37934 6825
rect -38757 6797 -37934 6821
rect -37882 6797 -37772 6849
rect -38757 6542 -37772 6797
rect -31724 7185 -31582 7237
rect -31530 7201 -31394 7237
rect -31342 7201 -30705 7253
rect -31530 7185 -30705 7201
rect -31724 7102 -30705 7185
rect -31724 7068 -31131 7102
rect -31724 7060 -31365 7068
rect -31724 7008 -31566 7060
rect -31514 7016 -31365 7060
rect -31313 7050 -31131 7068
rect -31079 7050 -30705 7102
rect -31313 7040 -30705 7050
rect -31313 7016 -30944 7040
rect -31514 7008 -30944 7016
rect -31724 6988 -30944 7008
rect -30892 6988 -30705 7040
rect -31724 6892 -30705 6988
rect -31724 6879 -31348 6892
rect -31724 6827 -31562 6879
rect -31510 6840 -31348 6879
rect -31296 6883 -30705 6892
rect -31296 6840 -31131 6883
rect -31510 6831 -31131 6840
rect -31079 6855 -30705 6883
rect -31079 6831 -30901 6855
rect -31510 6827 -30901 6831
rect -31724 6803 -30901 6827
rect -30849 6803 -30705 6855
rect -31724 6507 -30705 6803
rect -24931 8022 -23912 8238
rect -24931 8006 -24560 8022
rect -24931 7954 -24748 8006
rect -24696 7970 -24560 8006
rect -24508 7970 -23912 8022
rect -24696 7954 -23912 7970
rect -24931 7871 -23912 7954
rect -24931 7837 -24297 7871
rect -24931 7829 -24531 7837
rect -24931 7777 -24732 7829
rect -24680 7785 -24531 7829
rect -24479 7819 -24297 7837
rect -24245 7819 -23912 7871
rect -24479 7809 -23912 7819
rect -24479 7785 -24110 7809
rect -24680 7777 -24110 7785
rect -24931 7757 -24110 7777
rect -24058 7757 -23912 7809
rect -24931 7661 -23912 7757
rect -24931 7648 -24514 7661
rect -24931 7596 -24728 7648
rect -24676 7609 -24514 7648
rect -24462 7652 -23912 7661
rect -24462 7609 -24297 7652
rect -24676 7600 -24297 7609
rect -24245 7624 -23912 7652
rect -24245 7600 -24067 7624
rect -24676 7596 -24067 7600
rect -24931 7572 -24067 7596
rect -24015 7572 -23912 7624
rect -24931 7189 -23912 7572
rect -24931 7173 -24571 7189
rect -24931 7121 -24759 7173
rect -24707 7137 -24571 7173
rect -24519 7137 -23912 7189
rect -24707 7121 -23912 7137
rect -24931 7038 -23912 7121
rect -24931 7004 -24308 7038
rect -24931 6996 -24542 7004
rect -24931 6944 -24743 6996
rect -24691 6952 -24542 6996
rect -24490 6986 -24308 7004
rect -24256 6986 -23912 7038
rect -24490 6976 -23912 6986
rect -24490 6952 -24121 6976
rect -24691 6944 -24121 6952
rect -24931 6924 -24121 6944
rect -24069 6924 -23912 6976
rect -24931 6828 -23912 6924
rect -24931 6815 -24525 6828
rect -24931 6763 -24739 6815
rect -24687 6776 -24525 6815
rect -24473 6819 -23912 6828
rect -24473 6776 -24308 6819
rect -24687 6767 -24308 6776
rect -24256 6791 -23912 6819
rect -24256 6767 -24078 6791
rect -24687 6763 -24078 6767
rect -24931 6739 -24078 6763
rect -24026 6739 -23912 6791
rect -24931 6385 -23912 6739
rect -18061 8104 -17042 8354
rect -18061 8088 -17725 8104
rect -18061 8036 -17913 8088
rect -17861 8052 -17725 8088
rect -17673 8052 -17042 8104
rect -17861 8036 -17042 8052
rect -18061 7953 -17042 8036
rect -18061 7919 -17462 7953
rect -18061 7911 -17696 7919
rect -18061 7859 -17897 7911
rect -17845 7867 -17696 7911
rect -17644 7901 -17462 7919
rect -17410 7901 -17042 7953
rect -17644 7891 -17042 7901
rect -17644 7867 -17275 7891
rect -17845 7859 -17275 7867
rect -18061 7839 -17275 7859
rect -17223 7839 -17042 7891
rect -18061 7743 -17042 7839
rect -18061 7730 -17679 7743
rect -18061 7678 -17893 7730
rect -17841 7691 -17679 7730
rect -17627 7734 -17042 7743
rect -17627 7691 -17462 7734
rect -17841 7682 -17462 7691
rect -17410 7706 -17042 7734
rect -17410 7682 -17232 7706
rect -17841 7678 -17232 7682
rect -18061 7654 -17232 7678
rect -17180 7654 -17042 7706
rect -18061 7247 -17042 7654
rect -18061 7231 -17725 7247
rect -18061 7179 -17913 7231
rect -17861 7195 -17725 7231
rect -17673 7195 -17042 7247
rect -17861 7179 -17042 7195
rect -18061 7096 -17042 7179
rect -18061 7062 -17462 7096
rect -18061 7054 -17696 7062
rect -18061 7002 -17897 7054
rect -17845 7010 -17696 7054
rect -17644 7044 -17462 7062
rect -17410 7044 -17042 7096
rect -17644 7034 -17042 7044
rect -17644 7010 -17275 7034
rect -17845 7002 -17275 7010
rect -18061 6982 -17275 7002
rect -17223 6982 -17042 7034
rect -18061 6886 -17042 6982
rect -18061 6873 -17679 6886
rect -18061 6821 -17893 6873
rect -17841 6834 -17679 6873
rect -17627 6877 -17042 6886
rect -17627 6834 -17462 6877
rect -17841 6825 -17462 6834
rect -17410 6849 -17042 6877
rect -17410 6825 -17232 6849
rect -17841 6821 -17232 6825
rect -18061 6797 -17232 6821
rect -17180 6797 -17042 6849
rect -18061 6501 -17042 6797
rect -11069 8191 -10050 8319
rect -11069 8175 -10733 8191
rect -11069 8123 -10921 8175
rect -10869 8139 -10733 8175
rect -10681 8139 -10050 8191
rect -10869 8123 -10050 8139
rect -11069 8040 -10050 8123
rect -11069 8006 -10470 8040
rect -11069 7998 -10704 8006
rect -11069 7946 -10905 7998
rect -10853 7954 -10704 7998
rect -10652 7988 -10470 8006
rect -10418 7988 -10050 8040
rect -10652 7978 -10050 7988
rect -10652 7954 -10283 7978
rect -10853 7946 -10283 7954
rect -11069 7926 -10283 7946
rect -10231 7926 -10050 7978
rect -11069 7830 -10050 7926
rect -11069 7817 -10687 7830
rect -11069 7765 -10901 7817
rect -10849 7778 -10687 7817
rect -10635 7821 -10050 7830
rect -10635 7778 -10470 7821
rect -10849 7769 -10470 7778
rect -10418 7793 -10050 7821
rect -10418 7769 -10240 7793
rect -10849 7765 -10240 7769
rect -11069 7741 -10240 7765
rect -10188 7741 -10050 7793
rect -11069 7206 -10050 7741
rect -11069 7190 -10710 7206
rect -11069 7138 -10898 7190
rect -10846 7154 -10710 7190
rect -10658 7154 -10050 7206
rect -10846 7138 -10050 7154
rect -11069 7055 -10050 7138
rect -11069 7021 -10447 7055
rect -11069 7013 -10681 7021
rect -11069 6961 -10882 7013
rect -10830 6969 -10681 7013
rect -10629 7003 -10447 7021
rect -10395 7003 -10050 7055
rect -10629 6993 -10050 7003
rect -10629 6969 -10260 6993
rect -10830 6961 -10260 6969
rect -11069 6941 -10260 6961
rect -10208 6941 -10050 6993
rect -11069 6845 -10050 6941
rect -11069 6832 -10664 6845
rect -11069 6780 -10878 6832
rect -10826 6793 -10664 6832
rect -10612 6836 -10050 6845
rect -10612 6793 -10447 6836
rect -10826 6784 -10447 6793
rect -10395 6808 -10050 6836
rect -10395 6784 -10217 6808
rect -10826 6780 -10217 6784
rect -11069 6756 -10217 6780
rect -10165 6756 -10050 6808
rect -11069 6466 -10050 6756
rect -3635 8209 -2616 8337
rect -3635 8193 -3293 8209
rect -3635 8141 -3481 8193
rect -3429 8157 -3293 8193
rect -3241 8157 -2616 8209
rect -3429 8141 -2616 8157
rect -3635 8058 -2616 8141
rect -3635 8024 -3030 8058
rect -3635 8016 -3264 8024
rect -3635 7964 -3465 8016
rect -3413 7972 -3264 8016
rect -3212 8006 -3030 8024
rect -2978 8006 -2616 8058
rect -3212 7996 -2616 8006
rect -3212 7972 -2843 7996
rect -3413 7964 -2843 7972
rect -3635 7944 -2843 7964
rect -2791 7944 -2616 7996
rect -3635 7848 -2616 7944
rect -3635 7835 -3247 7848
rect -3635 7783 -3461 7835
rect -3409 7796 -3247 7835
rect -3195 7839 -2616 7848
rect -3195 7796 -3030 7839
rect -3409 7787 -3030 7796
rect -2978 7811 -2616 7839
rect -2978 7787 -2800 7811
rect -3409 7783 -2800 7787
rect -3635 7759 -2800 7783
rect -2748 7759 -2616 7811
rect -3635 7236 -2616 7759
rect -3635 7220 -3223 7236
rect -3635 7168 -3411 7220
rect -3359 7184 -3223 7220
rect -3171 7184 -2616 7236
rect -3359 7168 -2616 7184
rect -3635 7085 -2616 7168
rect -3635 7051 -2960 7085
rect -3635 7043 -3194 7051
rect -3635 6991 -3395 7043
rect -3343 6999 -3194 7043
rect -3142 7033 -2960 7051
rect -2908 7033 -2616 7085
rect -3142 7023 -2616 7033
rect -3142 6999 -2773 7023
rect -3343 6991 -2773 6999
rect -3635 6971 -2773 6991
rect -2721 6971 -2616 7023
rect -3635 6875 -2616 6971
rect -3635 6862 -3177 6875
rect -3635 6810 -3391 6862
rect -3339 6823 -3177 6862
rect -3125 6866 -2616 6875
rect -3125 6823 -2960 6866
rect -3339 6814 -2960 6823
rect -2908 6838 -2616 6866
rect -2908 6814 -2730 6838
rect -3339 6810 -2730 6814
rect -3635 6786 -2730 6810
rect -2678 6786 -2616 6838
rect -3635 6484 -2616 6786
rect 2058 8162 3077 8290
rect 2058 8146 2417 8162
rect 2058 8094 2229 8146
rect 2281 8110 2417 8146
rect 2469 8110 3077 8162
rect 2281 8094 3077 8110
rect 2058 8011 3077 8094
rect 2058 7977 2680 8011
rect 2058 7969 2446 7977
rect 2058 7917 2245 7969
rect 2297 7925 2446 7969
rect 2498 7959 2680 7977
rect 2732 7959 3077 8011
rect 2498 7949 3077 7959
rect 2498 7925 2867 7949
rect 2297 7917 2867 7925
rect 2058 7897 2867 7917
rect 2919 7897 3077 7949
rect 2058 7801 3077 7897
rect 2058 7788 2463 7801
rect 2058 7736 2249 7788
rect 2301 7749 2463 7788
rect 2515 7792 3077 7801
rect 2515 7749 2680 7792
rect 2301 7740 2680 7749
rect 2732 7764 3077 7792
rect 2732 7740 2910 7764
rect 2301 7736 2910 7740
rect 2058 7712 2910 7736
rect 2962 7712 3077 7764
rect 2058 7137 3077 7712
rect 2058 7121 2446 7137
rect 2058 7069 2258 7121
rect 2310 7085 2446 7121
rect 2498 7085 3077 7137
rect 2310 7069 3077 7085
rect 2058 6986 3077 7069
rect 2058 6952 2709 6986
rect 2058 6944 2475 6952
rect 2058 6892 2274 6944
rect 2326 6900 2475 6944
rect 2527 6934 2709 6952
rect 2761 6934 3077 6986
rect 2527 6924 3077 6934
rect 2527 6900 2896 6924
rect 2326 6892 2896 6900
rect 2058 6872 2896 6892
rect 2948 6872 3077 6924
rect 2058 6776 3077 6872
rect 2058 6763 2492 6776
rect 2058 6711 2278 6763
rect 2330 6724 2492 6763
rect 2544 6767 3077 6776
rect 2544 6724 2709 6767
rect 2330 6715 2709 6724
rect 2761 6739 3077 6767
rect 2761 6715 2939 6739
rect 2330 6711 2939 6715
rect 2058 6687 2939 6711
rect 2991 6687 3077 6739
rect 2058 6437 3077 6687
rect -61751 -68322 -60887 -68247
rect -61751 -68338 -61488 -68322
rect -61751 -68390 -61676 -68338
rect -61624 -68374 -61488 -68338
rect -61436 -68374 -60887 -68322
rect -61624 -68390 -60887 -68374
rect -61751 -68473 -60887 -68390
rect -61751 -68507 -61225 -68473
rect -61751 -68515 -61459 -68507
rect -61751 -68567 -61660 -68515
rect -61608 -68559 -61459 -68515
rect -61407 -68525 -61225 -68507
rect -61173 -68525 -60887 -68473
rect -61407 -68535 -60887 -68525
rect -61407 -68559 -61038 -68535
rect -61608 -68567 -61038 -68559
rect -61751 -68587 -61038 -68567
rect -60986 -68587 -60887 -68535
rect -61751 -68683 -60887 -68587
rect -61751 -68696 -61442 -68683
rect -61751 -68748 -61656 -68696
rect -61604 -68735 -61442 -68696
rect -61390 -68692 -60887 -68683
rect -61390 -68735 -61225 -68692
rect -61604 -68744 -61225 -68735
rect -61173 -68720 -60887 -68692
rect -61173 -68744 -60995 -68720
rect -61604 -68748 -60995 -68744
rect -61751 -68772 -60995 -68748
rect -60943 -68772 -60887 -68720
rect -61751 -68934 -60887 -68772
rect -55242 -68381 -54186 -68282
rect -55242 -68433 -54942 -68381
rect -54890 -68433 -54767 -68381
rect -54715 -68433 -54565 -68381
rect -54513 -68433 -54186 -68381
rect -55242 -68621 -54186 -68433
rect -55242 -68646 -54723 -68621
rect -55242 -68648 -54923 -68646
rect -55242 -68700 -55155 -68648
rect -55103 -68698 -54923 -68648
rect -54871 -68673 -54723 -68646
rect -54671 -68636 -54186 -68621
rect -54671 -68652 -54292 -68636
rect -54671 -68673 -54505 -68652
rect -54871 -68698 -54505 -68673
rect -55103 -68700 -54505 -68698
rect -55242 -68704 -54505 -68700
rect -54453 -68688 -54292 -68652
rect -54240 -68688 -54186 -68636
rect -54453 -68704 -54186 -68688
rect -55242 -68865 -54186 -68704
rect -55242 -68869 -54694 -68865
rect -55242 -68921 -54919 -68869
rect -54867 -68917 -54694 -68869
rect -54642 -68871 -54186 -68865
rect -54642 -68917 -54436 -68871
rect -54867 -68921 -54436 -68917
rect -55242 -68923 -54436 -68921
rect -54384 -68923 -54186 -68871
rect -48439 -68371 -47230 -68311
rect -48439 -68423 -48166 -68371
rect -48114 -68423 -47985 -68371
rect -47933 -68377 -47230 -68371
rect -47933 -68423 -47781 -68377
rect -48439 -68429 -47781 -68423
rect -47729 -68429 -47230 -68377
rect -48439 -68571 -47230 -68429
rect -48439 -68577 -47914 -68571
rect -48439 -68629 -48150 -68577
rect -48098 -68623 -47914 -68577
rect -47862 -68586 -47230 -68571
rect -47862 -68623 -47654 -68586
rect -48098 -68629 -47654 -68623
rect -48439 -68638 -47654 -68629
rect -47602 -68638 -47230 -68586
rect -48439 -68788 -47230 -68638
rect -48439 -68840 -48210 -68788
rect -48158 -68792 -47230 -68788
rect -48158 -68840 -47968 -68792
rect -48439 -68844 -47968 -68840
rect -47916 -68844 -47768 -68792
rect -47716 -68802 -47230 -68792
rect -47716 -68844 -47464 -68802
rect -48439 -68854 -47464 -68844
rect -47412 -68854 -47230 -68802
rect -48439 -68909 -47230 -68854
rect -41649 -68371 -40440 -68326
rect -21096 -68350 -20092 -68263
rect -41649 -68375 -41149 -68371
rect -41649 -68427 -41330 -68375
rect -41278 -68423 -41149 -68375
rect -41097 -68381 -40440 -68371
rect -41097 -68423 -40949 -68381
rect -41278 -68427 -40949 -68423
rect -41649 -68433 -40949 -68427
rect -40897 -68433 -40440 -68381
rect -41649 -68544 -40440 -68433
rect -41649 -68583 -41328 -68544
rect -41649 -68635 -41515 -68583
rect -41463 -68596 -41328 -68583
rect -41276 -68548 -40440 -68544
rect -41276 -68558 -40888 -68548
rect -41276 -68596 -41115 -68558
rect -41463 -68610 -41115 -68596
rect -41063 -68600 -40888 -68558
rect -40836 -68571 -40440 -68548
rect -40836 -68600 -40692 -68571
rect -41063 -68610 -40692 -68600
rect -41463 -68623 -40692 -68610
rect -40640 -68623 -40440 -68571
rect -41463 -68635 -40440 -68623
rect -41649 -68744 -40440 -68635
rect -41649 -68761 -41082 -68744
rect -41649 -68813 -41315 -68761
rect -41263 -68796 -41082 -68761
rect -41030 -68756 -40440 -68744
rect -41030 -68796 -40834 -68756
rect -41263 -68808 -40834 -68796
rect -40782 -68808 -40440 -68756
rect -41263 -68813 -40440 -68808
rect -55242 -68970 -54186 -68923
rect -41649 -68924 -40440 -68813
rect -34904 -68410 -33695 -68353
rect -34904 -68462 -34575 -68410
rect -34523 -68417 -33695 -68410
rect -34523 -68462 -34394 -68417
rect -34904 -68469 -34394 -68462
rect -34342 -68469 -34219 -68417
rect -34167 -68469 -33695 -68417
rect -34904 -68627 -33695 -68469
rect -34904 -68633 -33998 -68627
rect -34904 -68652 -34558 -68633
rect -34904 -68704 -34817 -68652
rect -34765 -68685 -34558 -68652
rect -34506 -68685 -34327 -68633
rect -34275 -68679 -33998 -68633
rect -33946 -68679 -33695 -68627
rect -34275 -68685 -33695 -68679
rect -34765 -68704 -33695 -68685
rect -34904 -68836 -33695 -68704
rect -34904 -68850 -33841 -68836
rect -34904 -68902 -34579 -68850
rect -34527 -68902 -34344 -68850
rect -34292 -68854 -33841 -68850
rect -34292 -68902 -34104 -68854
rect -34904 -68906 -34104 -68902
rect -34052 -68888 -33841 -68854
rect -33789 -68888 -33695 -68836
rect -34052 -68906 -33695 -68888
rect -34904 -68951 -33695 -68906
rect -28030 -68390 -26900 -68350
rect -28030 -68442 -27725 -68390
rect -27673 -68397 -26900 -68390
rect -27673 -68442 -27544 -68397
rect -28030 -68449 -27544 -68442
rect -27492 -68449 -27369 -68397
rect -27317 -68449 -26900 -68397
rect -28030 -68607 -26900 -68449
rect -28030 -68613 -27148 -68607
rect -28030 -68632 -27708 -68613
rect -28030 -68684 -27967 -68632
rect -27915 -68665 -27708 -68632
rect -27656 -68665 -27477 -68613
rect -27425 -68659 -27148 -68613
rect -27096 -68659 -26900 -68607
rect -27425 -68665 -26900 -68659
rect -27915 -68684 -26900 -68665
rect -28030 -68816 -26900 -68684
rect -28030 -68830 -26991 -68816
rect -28030 -68882 -27729 -68830
rect -27677 -68882 -27494 -68830
rect -27442 -68834 -26991 -68830
rect -27442 -68882 -27254 -68834
rect -28030 -68886 -27254 -68882
rect -27202 -68868 -26991 -68834
rect -26939 -68868 -26900 -68816
rect -27202 -68886 -26900 -68868
rect -28030 -68930 -26900 -68886
rect -21096 -68390 -19960 -68350
rect -21096 -68442 -20785 -68390
rect -20733 -68397 -19960 -68390
rect -20733 -68442 -20604 -68397
rect -21096 -68449 -20604 -68442
rect -20552 -68449 -20429 -68397
rect -20377 -68449 -19960 -68397
rect -21096 -68607 -19960 -68449
rect -21096 -68613 -20208 -68607
rect -21096 -68632 -20768 -68613
rect -21096 -68684 -21027 -68632
rect -20975 -68665 -20768 -68632
rect -20716 -68665 -20537 -68613
rect -20485 -68659 -20208 -68613
rect -20156 -68659 -19960 -68607
rect -20485 -68665 -19960 -68659
rect -20975 -68684 -19960 -68665
rect -21096 -68816 -19960 -68684
rect -21096 -68830 -20051 -68816
rect -21096 -68882 -20789 -68830
rect -20737 -68882 -20554 -68830
rect -20502 -68834 -20051 -68830
rect -20502 -68882 -20314 -68834
rect -21096 -68886 -20314 -68882
rect -20262 -68868 -20051 -68834
rect -19999 -68868 -19960 -68816
rect -20262 -68886 -19960 -68868
rect -21096 -68930 -19960 -68886
rect -14409 -68383 -13405 -68255
rect -14409 -68435 -14122 -68383
rect -14070 -68388 -13405 -68383
rect -14070 -68435 -13943 -68388
rect -14409 -68440 -13943 -68435
rect -13891 -68440 -13760 -68388
rect -13708 -68440 -13405 -68388
rect -14409 -68636 -13405 -68440
rect -14409 -68640 -13635 -68636
rect -14409 -68646 -13843 -68640
rect -14409 -68652 -14035 -68646
rect -14409 -68704 -14260 -68652
rect -14208 -68698 -14035 -68652
rect -13983 -68692 -13843 -68646
rect -13791 -68688 -13635 -68640
rect -13583 -68688 -13405 -68636
rect -13791 -68692 -13405 -68688
rect -13983 -68698 -13405 -68692
rect -14208 -68704 -13405 -68698
rect -14409 -68850 -13405 -68704
rect -14409 -68902 -14197 -68850
rect -14145 -68902 -13978 -68850
rect -13926 -68902 -13789 -68850
rect -13737 -68902 -13541 -68850
rect -13489 -68902 -13405 -68850
rect -21096 -68951 -20092 -68930
rect -14409 -68943 -13405 -68902
rect -7481 -68363 -6477 -68255
rect -7481 -68415 -7284 -68363
rect -7232 -68415 -7109 -68363
rect -7057 -68415 -6919 -68363
rect -6867 -68415 -6477 -68363
rect -7481 -68613 -6477 -68415
rect -7481 -68619 -6646 -68613
rect -7481 -68625 -6907 -68619
rect -7481 -68631 -7127 -68625
rect -7481 -68683 -7400 -68631
rect -7348 -68677 -7127 -68631
rect -7075 -68671 -6907 -68625
rect -6855 -68665 -6646 -68619
rect -6594 -68665 -6477 -68613
rect -6855 -68671 -6477 -68665
rect -7075 -68677 -6477 -68671
rect -7348 -68683 -6477 -68677
rect -7481 -68848 -6477 -68683
rect -7481 -68854 -6721 -68848
rect -7481 -68856 -7150 -68854
rect -7481 -68908 -7365 -68856
rect -7313 -68906 -7150 -68856
rect -7098 -68906 -6932 -68854
rect -6880 -68900 -6721 -68854
rect -6669 -68900 -6477 -68848
rect -6880 -68906 -6477 -68900
rect -7313 -68908 -6477 -68906
rect -7481 -68943 -6477 -68908
rect -676 -68360 328 -68259
rect -676 -68363 -68 -68360
rect -676 -68415 -474 -68363
rect -422 -68367 -68 -68363
rect -422 -68415 -281 -68367
rect -676 -68419 -281 -68415
rect -229 -68412 -68 -68367
rect -16 -68412 328 -68360
rect -229 -68419 328 -68412
rect -676 -68596 328 -68419
rect -676 -68600 147 -68596
rect -676 -68604 -343 -68600
rect -676 -68656 -593 -68604
rect -541 -68652 -343 -68604
rect -291 -68652 -110 -68600
rect -58 -68648 147 -68600
rect 199 -68648 328 -68596
rect -58 -68652 328 -68648
rect -541 -68656 328 -68652
rect -676 -68850 328 -68656
rect -676 -68854 -306 -68850
rect -676 -68906 -564 -68854
rect -512 -68902 -306 -68854
rect -254 -68854 328 -68850
rect -254 -68902 -68 -68854
rect -512 -68906 -68 -68902
rect -16 -68861 328 -68854
rect -16 -68906 186 -68861
rect -676 -68913 186 -68906
rect 238 -68913 328 -68861
rect -676 -68947 328 -68913
rect 5835 -68354 6839 -68257
rect 5835 -68406 6320 -68354
rect 6372 -68406 6508 -68354
rect 6560 -68360 6839 -68354
rect 6560 -68406 6710 -68360
rect 5835 -68412 6710 -68406
rect 6762 -68412 6839 -68360
rect 5835 -68575 6839 -68412
rect 5835 -68627 6145 -68575
rect 6197 -68579 6608 -68575
rect 6197 -68627 6397 -68579
rect 5835 -68631 6397 -68627
rect 6449 -68627 6608 -68579
rect 6660 -68627 6839 -68575
rect 6449 -68631 6839 -68627
rect 5835 -68690 6839 -68631
rect 5835 -68742 5933 -68690
rect 5985 -68742 6839 -68690
rect 5835 -68854 6839 -68742
rect 5835 -68856 6329 -68854
rect 5835 -68908 6141 -68856
rect 6193 -68906 6329 -68856
rect 6381 -68906 6535 -68854
rect 6587 -68856 6839 -68854
rect 6587 -68906 6739 -68856
rect 6193 -68908 6739 -68906
rect 6791 -68908 6839 -68856
rect 5835 -68945 6839 -68908
<< via1 >>
rect -51864 8234 -51812 8286
rect -51676 8250 -51624 8302
rect -65121 7913 -65069 7965
rect -64933 7929 -64881 7981
rect -65105 7736 -65053 7788
rect -64904 7744 -64852 7796
rect -64670 7778 -64618 7830
rect -64483 7716 -64431 7768
rect -65101 7555 -65049 7607
rect -64887 7568 -64835 7620
rect -64670 7559 -64618 7611
rect -64440 7531 -64388 7583
rect -65144 7095 -65092 7147
rect -64956 7111 -64904 7163
rect -65128 6918 -65076 6970
rect -64927 6926 -64875 6978
rect -64693 6960 -64641 7012
rect -64506 6898 -64454 6950
rect -65124 6737 -65072 6789
rect -64910 6750 -64858 6802
rect -64693 6741 -64641 6793
rect -64463 6713 -64411 6765
rect -58926 7995 -58874 8047
rect -58738 8011 -58686 8063
rect -58910 7818 -58858 7870
rect -58709 7826 -58657 7878
rect -58475 7860 -58423 7912
rect -58288 7798 -58236 7850
rect -58906 7637 -58854 7689
rect -58692 7650 -58640 7702
rect -58475 7641 -58423 7693
rect -58245 7613 -58193 7665
rect -58926 7115 -58874 7167
rect -58738 7131 -58686 7183
rect -58910 6938 -58858 6990
rect -58709 6946 -58657 6998
rect -58475 6980 -58423 7032
rect -58288 6918 -58236 6970
rect -58906 6757 -58854 6809
rect -58692 6770 -58640 6822
rect -58475 6761 -58423 6813
rect -58245 6733 -58193 6785
rect -51848 8057 -51796 8109
rect -51647 8065 -51595 8117
rect -51413 8099 -51361 8151
rect -51226 8037 -51174 8089
rect -51844 7876 -51792 7928
rect -51630 7889 -51578 7941
rect -51413 7880 -51361 7932
rect -51183 7852 -51131 7904
rect -51884 7368 -51832 7420
rect -51696 7384 -51644 7436
rect -51868 7191 -51816 7243
rect -51667 7199 -51615 7251
rect -51433 7233 -51381 7285
rect -51246 7171 -51194 7223
rect -51864 7010 -51812 7062
rect -51650 7023 -51598 7075
rect -51433 7014 -51381 7066
rect -51203 6986 -51151 7038
rect -45327 8088 -45275 8140
rect -45139 8104 -45087 8156
rect -45311 7911 -45259 7963
rect -45110 7919 -45058 7971
rect -44876 7953 -44824 8005
rect -44689 7891 -44637 7943
rect -45307 7730 -45255 7782
rect -45093 7743 -45041 7795
rect -44876 7734 -44824 7786
rect -44646 7706 -44594 7758
rect -45356 7156 -45304 7208
rect -45168 7172 -45116 7224
rect -45340 6979 -45288 7031
rect -45139 6987 -45087 7039
rect -44905 7021 -44853 7073
rect -44718 6959 -44666 7011
rect -45336 6798 -45284 6850
rect -45122 6811 -45070 6863
rect -44905 6802 -44853 6854
rect -44675 6774 -44623 6826
rect -38626 8018 -38574 8070
rect -38438 8034 -38386 8086
rect -38610 7841 -38558 7893
rect -38409 7849 -38357 7901
rect -38175 7883 -38123 7935
rect -37988 7821 -37936 7873
rect -38606 7660 -38554 7712
rect -38392 7673 -38340 7725
rect -38175 7664 -38123 7716
rect -37945 7636 -37893 7688
rect -38615 7179 -38563 7231
rect -38427 7195 -38375 7247
rect -31599 8077 -31547 8129
rect -31411 8093 -31359 8145
rect -31583 7900 -31531 7952
rect -31382 7908 -31330 7960
rect -31148 7942 -31096 7994
rect -30961 7880 -30909 7932
rect -31579 7719 -31527 7771
rect -31365 7732 -31313 7784
rect -31148 7723 -31096 7775
rect -30918 7695 -30866 7747
rect -38599 7002 -38547 7054
rect -38398 7010 -38346 7062
rect -38164 7044 -38112 7096
rect -37977 6982 -37925 7034
rect -38595 6821 -38543 6873
rect -38381 6834 -38329 6886
rect -38164 6825 -38112 6877
rect -37934 6797 -37882 6849
rect -31582 7185 -31530 7237
rect -31394 7201 -31342 7253
rect -31566 7008 -31514 7060
rect -31365 7016 -31313 7068
rect -31131 7050 -31079 7102
rect -30944 6988 -30892 7040
rect -31562 6827 -31510 6879
rect -31348 6840 -31296 6892
rect -31131 6831 -31079 6883
rect -30901 6803 -30849 6855
rect -24748 7954 -24696 8006
rect -24560 7970 -24508 8022
rect -24732 7777 -24680 7829
rect -24531 7785 -24479 7837
rect -24297 7819 -24245 7871
rect -24110 7757 -24058 7809
rect -24728 7596 -24676 7648
rect -24514 7609 -24462 7661
rect -24297 7600 -24245 7652
rect -24067 7572 -24015 7624
rect -24759 7121 -24707 7173
rect -24571 7137 -24519 7189
rect -24743 6944 -24691 6996
rect -24542 6952 -24490 7004
rect -24308 6986 -24256 7038
rect -24121 6924 -24069 6976
rect -24739 6763 -24687 6815
rect -24525 6776 -24473 6828
rect -24308 6767 -24256 6819
rect -24078 6739 -24026 6791
rect -17913 8036 -17861 8088
rect -17725 8052 -17673 8104
rect -17897 7859 -17845 7911
rect -17696 7867 -17644 7919
rect -17462 7901 -17410 7953
rect -17275 7839 -17223 7891
rect -17893 7678 -17841 7730
rect -17679 7691 -17627 7743
rect -17462 7682 -17410 7734
rect -17232 7654 -17180 7706
rect -17913 7179 -17861 7231
rect -17725 7195 -17673 7247
rect -17897 7002 -17845 7054
rect -17696 7010 -17644 7062
rect -17462 7044 -17410 7096
rect -17275 6982 -17223 7034
rect -17893 6821 -17841 6873
rect -17679 6834 -17627 6886
rect -17462 6825 -17410 6877
rect -17232 6797 -17180 6849
rect -10921 8123 -10869 8175
rect -10733 8139 -10681 8191
rect -10905 7946 -10853 7998
rect -10704 7954 -10652 8006
rect -10470 7988 -10418 8040
rect -10283 7926 -10231 7978
rect -10901 7765 -10849 7817
rect -10687 7778 -10635 7830
rect -10470 7769 -10418 7821
rect -10240 7741 -10188 7793
rect -10898 7138 -10846 7190
rect -10710 7154 -10658 7206
rect -10882 6961 -10830 7013
rect -10681 6969 -10629 7021
rect -10447 7003 -10395 7055
rect -10260 6941 -10208 6993
rect -10878 6780 -10826 6832
rect -10664 6793 -10612 6845
rect -10447 6784 -10395 6836
rect -10217 6756 -10165 6808
rect -3481 8141 -3429 8193
rect -3293 8157 -3241 8209
rect -3465 7964 -3413 8016
rect -3264 7972 -3212 8024
rect -3030 8006 -2978 8058
rect -2843 7944 -2791 7996
rect -3461 7783 -3409 7835
rect -3247 7796 -3195 7848
rect -3030 7787 -2978 7839
rect -2800 7759 -2748 7811
rect -3411 7168 -3359 7220
rect -3223 7184 -3171 7236
rect -3395 6991 -3343 7043
rect -3194 6999 -3142 7051
rect -2960 7033 -2908 7085
rect -2773 6971 -2721 7023
rect -3391 6810 -3339 6862
rect -3177 6823 -3125 6875
rect -2960 6814 -2908 6866
rect -2730 6786 -2678 6838
rect 2229 8094 2281 8146
rect 2417 8110 2469 8162
rect 2245 7917 2297 7969
rect 2446 7925 2498 7977
rect 2680 7959 2732 8011
rect 2867 7897 2919 7949
rect 2249 7736 2301 7788
rect 2463 7749 2515 7801
rect 2680 7740 2732 7792
rect 2910 7712 2962 7764
rect 2258 7069 2310 7121
rect 2446 7085 2498 7137
rect 2274 6892 2326 6944
rect 2475 6900 2527 6952
rect 2709 6934 2761 6986
rect 2896 6872 2948 6924
rect 2278 6711 2330 6763
rect 2492 6724 2544 6776
rect 2709 6715 2761 6767
rect 2939 6687 2991 6739
rect -61676 -68390 -61624 -68338
rect -61488 -68374 -61436 -68322
rect -61660 -68567 -61608 -68515
rect -61459 -68559 -61407 -68507
rect -61225 -68525 -61173 -68473
rect -61038 -68587 -60986 -68535
rect -61656 -68748 -61604 -68696
rect -61442 -68735 -61390 -68683
rect -61225 -68744 -61173 -68692
rect -60995 -68772 -60943 -68720
rect -54942 -68433 -54890 -68381
rect -54767 -68433 -54715 -68381
rect -54565 -68433 -54513 -68381
rect -55155 -68700 -55103 -68648
rect -54923 -68698 -54871 -68646
rect -54723 -68673 -54671 -68621
rect -54505 -68704 -54453 -68652
rect -54292 -68688 -54240 -68636
rect -54919 -68921 -54867 -68869
rect -54694 -68917 -54642 -68865
rect -54436 -68923 -54384 -68871
rect -48166 -68423 -48114 -68371
rect -47985 -68423 -47933 -68371
rect -47781 -68429 -47729 -68377
rect -48150 -68629 -48098 -68577
rect -47914 -68623 -47862 -68571
rect -47654 -68638 -47602 -68586
rect -48210 -68840 -48158 -68788
rect -47968 -68844 -47916 -68792
rect -47768 -68844 -47716 -68792
rect -47464 -68854 -47412 -68802
rect -41330 -68427 -41278 -68375
rect -41149 -68423 -41097 -68371
rect -40949 -68433 -40897 -68381
rect -41515 -68635 -41463 -68583
rect -41328 -68596 -41276 -68544
rect -41115 -68610 -41063 -68558
rect -40888 -68600 -40836 -68548
rect -40692 -68623 -40640 -68571
rect -41315 -68813 -41263 -68761
rect -41082 -68796 -41030 -68744
rect -40834 -68808 -40782 -68756
rect -34575 -68462 -34523 -68410
rect -34394 -68469 -34342 -68417
rect -34219 -68469 -34167 -68417
rect -34817 -68704 -34765 -68652
rect -34558 -68685 -34506 -68633
rect -34327 -68685 -34275 -68633
rect -33998 -68679 -33946 -68627
rect -34579 -68902 -34527 -68850
rect -34344 -68902 -34292 -68850
rect -34104 -68906 -34052 -68854
rect -33841 -68888 -33789 -68836
rect -27725 -68442 -27673 -68390
rect -27544 -68449 -27492 -68397
rect -27369 -68449 -27317 -68397
rect -27967 -68684 -27915 -68632
rect -27708 -68665 -27656 -68613
rect -27477 -68665 -27425 -68613
rect -27148 -68659 -27096 -68607
rect -27729 -68882 -27677 -68830
rect -27494 -68882 -27442 -68830
rect -27254 -68886 -27202 -68834
rect -26991 -68868 -26939 -68816
rect -20785 -68442 -20733 -68390
rect -20604 -68449 -20552 -68397
rect -20429 -68449 -20377 -68397
rect -21027 -68684 -20975 -68632
rect -20768 -68665 -20716 -68613
rect -20537 -68665 -20485 -68613
rect -20208 -68659 -20156 -68607
rect -20789 -68882 -20737 -68830
rect -20554 -68882 -20502 -68830
rect -20314 -68886 -20262 -68834
rect -20051 -68868 -19999 -68816
rect -14122 -68435 -14070 -68383
rect -13943 -68440 -13891 -68388
rect -13760 -68440 -13708 -68388
rect -14260 -68704 -14208 -68652
rect -14035 -68698 -13983 -68646
rect -13843 -68692 -13791 -68640
rect -13635 -68688 -13583 -68636
rect -14197 -68902 -14145 -68850
rect -13978 -68902 -13926 -68850
rect -13789 -68902 -13737 -68850
rect -13541 -68902 -13489 -68850
rect -7284 -68415 -7232 -68363
rect -7109 -68415 -7057 -68363
rect -6919 -68415 -6867 -68363
rect -7400 -68683 -7348 -68631
rect -7127 -68677 -7075 -68625
rect -6907 -68671 -6855 -68619
rect -6646 -68665 -6594 -68613
rect -7365 -68908 -7313 -68856
rect -7150 -68906 -7098 -68854
rect -6932 -68906 -6880 -68854
rect -6721 -68900 -6669 -68848
rect -474 -68415 -422 -68363
rect -281 -68419 -229 -68367
rect -68 -68412 -16 -68360
rect -593 -68656 -541 -68604
rect -343 -68652 -291 -68600
rect -110 -68652 -58 -68600
rect 147 -68648 199 -68596
rect -564 -68906 -512 -68854
rect -306 -68902 -254 -68850
rect -68 -68906 -16 -68854
rect 186 -68913 238 -68861
rect 6320 -68406 6372 -68354
rect 6508 -68406 6560 -68354
rect 6710 -68412 6762 -68360
rect 6145 -68627 6197 -68575
rect 6397 -68631 6449 -68579
rect 6608 -68627 6660 -68575
rect 5933 -68742 5985 -68690
rect 6141 -68908 6193 -68856
rect 6329 -68906 6381 -68854
rect 6535 -68906 6587 -68854
rect 6739 -68908 6791 -68856
<< metal2 >>
rect -52012 8304 -51027 8429
rect -52012 8288 -51678 8304
rect -52012 8232 -51866 8288
rect -51810 8248 -51678 8288
rect -51622 8248 -51027 8304
rect -51810 8232 -51027 8248
rect -52012 8153 -51027 8232
rect -65244 7983 -64259 8149
rect -65244 7967 -64935 7983
rect -65244 7911 -65123 7967
rect -65067 7927 -64935 7967
rect -64879 7927 -64259 7983
rect -65067 7911 -64259 7927
rect -65244 7832 -64259 7911
rect -65244 7798 -64672 7832
rect -65244 7790 -64906 7798
rect -65244 7734 -65107 7790
rect -65051 7742 -64906 7790
rect -64850 7776 -64672 7798
rect -64616 7776 -64259 7832
rect -64850 7770 -64259 7776
rect -64850 7742 -64485 7770
rect -65051 7734 -64485 7742
rect -65244 7714 -64485 7734
rect -64429 7714 -64259 7770
rect -65244 7622 -64259 7714
rect -65244 7609 -64889 7622
rect -65244 7553 -65103 7609
rect -65047 7566 -64889 7609
rect -64833 7613 -64259 7622
rect -64833 7566 -64672 7613
rect -65047 7557 -64672 7566
rect -64616 7585 -64259 7613
rect -64616 7557 -64442 7585
rect -65047 7553 -64442 7557
rect -65244 7529 -64442 7553
rect -64386 7529 -64259 7585
rect -65244 7165 -64259 7529
rect -65244 7149 -64958 7165
rect -65244 7093 -65146 7149
rect -65090 7109 -64958 7149
rect -64902 7109 -64259 7165
rect -65090 7093 -64259 7109
rect -65244 7014 -64259 7093
rect -65244 6980 -64695 7014
rect -65244 6972 -64929 6980
rect -65244 6916 -65130 6972
rect -65074 6924 -64929 6972
rect -64873 6958 -64695 6980
rect -64639 6958 -64259 7014
rect -64873 6952 -64259 6958
rect -64873 6924 -64508 6952
rect -65074 6916 -64508 6924
rect -65244 6896 -64508 6916
rect -64452 6896 -64259 6952
rect -65244 6804 -64259 6896
rect -65244 6791 -64912 6804
rect -65244 6735 -65126 6791
rect -65070 6748 -64912 6791
rect -64856 6795 -64259 6804
rect -64856 6748 -64695 6795
rect -65070 6739 -64695 6748
rect -64639 6767 -64259 6795
rect -64639 6739 -64465 6767
rect -65070 6735 -64465 6739
rect -65244 6711 -64465 6735
rect -64409 6711 -64259 6767
rect -65244 6454 -64259 6711
rect -59062 8065 -58077 8149
rect -59062 8049 -58740 8065
rect -59062 7993 -58928 8049
rect -58872 8009 -58740 8049
rect -58684 8009 -58077 8065
rect -58872 7993 -58077 8009
rect -59062 7914 -58077 7993
rect -59062 7880 -58477 7914
rect -59062 7872 -58711 7880
rect -59062 7816 -58912 7872
rect -58856 7824 -58711 7872
rect -58655 7858 -58477 7880
rect -58421 7858 -58077 7914
rect -58655 7852 -58077 7858
rect -58655 7824 -58290 7852
rect -58856 7816 -58290 7824
rect -59062 7796 -58290 7816
rect -58234 7796 -58077 7852
rect -59062 7704 -58077 7796
rect -59062 7691 -58694 7704
rect -59062 7635 -58908 7691
rect -58852 7648 -58694 7691
rect -58638 7695 -58077 7704
rect -58638 7648 -58477 7695
rect -58852 7639 -58477 7648
rect -58421 7667 -58077 7695
rect -58421 7639 -58247 7667
rect -58852 7635 -58247 7639
rect -59062 7611 -58247 7635
rect -58191 7611 -58077 7667
rect -59062 7185 -58077 7611
rect -59062 7169 -58740 7185
rect -59062 7113 -58928 7169
rect -58872 7129 -58740 7169
rect -58684 7129 -58077 7185
rect -58872 7113 -58077 7129
rect -59062 7034 -58077 7113
rect -59062 7000 -58477 7034
rect -59062 6992 -58711 7000
rect -59062 6936 -58912 6992
rect -58856 6944 -58711 6992
rect -58655 6978 -58477 7000
rect -58421 6978 -58077 7034
rect -58655 6972 -58077 6978
rect -58655 6944 -58290 6972
rect -58856 6936 -58290 6944
rect -59062 6916 -58290 6936
rect -58234 6916 -58077 6972
rect -59062 6824 -58077 6916
rect -59062 6811 -58694 6824
rect -59062 6755 -58908 6811
rect -58852 6768 -58694 6811
rect -58638 6815 -58077 6824
rect -58638 6768 -58477 6815
rect -58852 6759 -58477 6768
rect -58421 6787 -58077 6815
rect -58421 6759 -58247 6787
rect -58852 6755 -58247 6759
rect -59062 6731 -58247 6755
rect -58191 6731 -58077 6787
rect -52012 8119 -51415 8153
rect -52012 8111 -51649 8119
rect -52012 8055 -51850 8111
rect -51794 8063 -51649 8111
rect -51593 8097 -51415 8119
rect -51359 8097 -51027 8153
rect -51593 8091 -51027 8097
rect -51593 8063 -51228 8091
rect -51794 8055 -51228 8063
rect -52012 8035 -51228 8055
rect -51172 8035 -51027 8091
rect -52012 7943 -51027 8035
rect -52012 7930 -51632 7943
rect -52012 7874 -51846 7930
rect -51790 7887 -51632 7930
rect -51576 7934 -51027 7943
rect -51576 7887 -51415 7934
rect -51790 7878 -51415 7887
rect -51359 7906 -51027 7934
rect -51359 7878 -51185 7906
rect -51790 7874 -51185 7878
rect -52012 7850 -51185 7874
rect -51129 7850 -51027 7906
rect -52012 7438 -51027 7850
rect -52012 7422 -51698 7438
rect -52012 7366 -51886 7422
rect -51830 7382 -51698 7422
rect -51642 7382 -51027 7438
rect -51830 7366 -51027 7382
rect -52012 7287 -51027 7366
rect -52012 7253 -51435 7287
rect -52012 7245 -51669 7253
rect -52012 7189 -51870 7245
rect -51814 7197 -51669 7245
rect -51613 7231 -51435 7253
rect -51379 7231 -51027 7287
rect -51613 7225 -51027 7231
rect -51613 7197 -51248 7225
rect -51814 7189 -51248 7197
rect -52012 7169 -51248 7189
rect -51192 7169 -51027 7225
rect -52012 7077 -51027 7169
rect -52012 7064 -51652 7077
rect -52012 7008 -51866 7064
rect -51810 7021 -51652 7064
rect -51596 7068 -51027 7077
rect -51596 7021 -51435 7068
rect -51810 7012 -51435 7021
rect -51379 7040 -51027 7068
rect -51379 7012 -51205 7040
rect -51810 7008 -51205 7012
rect -52012 6984 -51205 7008
rect -51149 6984 -51027 7040
rect -52012 6734 -51027 6984
rect -45475 8158 -44490 8254
rect -45475 8142 -45141 8158
rect -45475 8086 -45329 8142
rect -45273 8102 -45141 8142
rect -45085 8102 -44490 8158
rect -45273 8086 -44490 8102
rect -45475 8007 -44490 8086
rect -45475 7973 -44878 8007
rect -45475 7965 -45112 7973
rect -45475 7909 -45313 7965
rect -45257 7917 -45112 7965
rect -45056 7951 -44878 7973
rect -44822 7951 -44490 8007
rect -45056 7945 -44490 7951
rect -45056 7917 -44691 7945
rect -45257 7909 -44691 7917
rect -45475 7889 -44691 7909
rect -44635 7889 -44490 7945
rect -45475 7797 -44490 7889
rect -45475 7784 -45095 7797
rect -45475 7728 -45309 7784
rect -45253 7741 -45095 7784
rect -45039 7788 -44490 7797
rect -45039 7741 -44878 7788
rect -45253 7732 -44878 7741
rect -44822 7760 -44490 7788
rect -44822 7732 -44648 7760
rect -45253 7728 -44648 7732
rect -45475 7704 -44648 7728
rect -44592 7704 -44490 7760
rect -45475 7226 -44490 7704
rect -45475 7210 -45170 7226
rect -45475 7154 -45358 7210
rect -45302 7170 -45170 7210
rect -45114 7170 -44490 7226
rect -45302 7154 -44490 7170
rect -45475 7075 -44490 7154
rect -45475 7041 -44907 7075
rect -45475 7033 -45141 7041
rect -45475 6977 -45342 7033
rect -45286 6985 -45141 7033
rect -45085 7019 -44907 7041
rect -44851 7019 -44490 7075
rect -45085 7013 -44490 7019
rect -45085 6985 -44720 7013
rect -45286 6977 -44720 6985
rect -45475 6957 -44720 6977
rect -44664 6957 -44490 7013
rect -45475 6865 -44490 6957
rect -45475 6852 -45124 6865
rect -45475 6796 -45338 6852
rect -45282 6809 -45124 6852
rect -45068 6856 -44490 6865
rect -45068 6809 -44907 6856
rect -45282 6800 -44907 6809
rect -44851 6828 -44490 6856
rect -44851 6800 -44677 6828
rect -45282 6796 -44677 6800
rect -45475 6772 -44677 6796
rect -44621 6772 -44490 6828
rect -59062 6454 -58077 6731
rect -45475 6559 -44490 6772
rect -38757 8088 -37772 8237
rect -38757 8072 -38440 8088
rect -38757 8016 -38628 8072
rect -38572 8032 -38440 8072
rect -38384 8032 -37772 8088
rect -38572 8016 -37772 8032
rect -38757 7937 -37772 8016
rect -38757 7903 -38177 7937
rect -38757 7895 -38411 7903
rect -38757 7839 -38612 7895
rect -38556 7847 -38411 7895
rect -38355 7881 -38177 7903
rect -38121 7881 -37772 7937
rect -38355 7875 -37772 7881
rect -38355 7847 -37990 7875
rect -38556 7839 -37990 7847
rect -38757 7819 -37990 7839
rect -37934 7819 -37772 7875
rect -38757 7727 -37772 7819
rect -38757 7714 -38394 7727
rect -38757 7658 -38608 7714
rect -38552 7671 -38394 7714
rect -38338 7718 -37772 7727
rect -38338 7671 -38177 7718
rect -38552 7662 -38177 7671
rect -38121 7690 -37772 7718
rect -38121 7662 -37947 7690
rect -38552 7658 -37947 7662
rect -38757 7634 -37947 7658
rect -37891 7634 -37772 7690
rect -38757 7249 -37772 7634
rect -38757 7233 -38429 7249
rect -38757 7177 -38617 7233
rect -38561 7193 -38429 7233
rect -38373 7193 -37772 7249
rect -38561 7177 -37772 7193
rect -38757 7098 -37772 7177
rect -38757 7064 -38166 7098
rect -38757 7056 -38400 7064
rect -38757 7000 -38601 7056
rect -38545 7008 -38400 7056
rect -38344 7042 -38166 7064
rect -38110 7042 -37772 7098
rect -38344 7036 -37772 7042
rect -38344 7008 -37979 7036
rect -38545 7000 -37979 7008
rect -38757 6980 -37979 7000
rect -37923 6980 -37772 7036
rect -38757 6888 -37772 6980
rect -38757 6875 -38383 6888
rect -38757 6819 -38597 6875
rect -38541 6832 -38383 6875
rect -38327 6879 -37772 6888
rect -38327 6832 -38166 6879
rect -38541 6823 -38166 6832
rect -38110 6851 -37772 6879
rect -38110 6823 -37936 6851
rect -38541 6819 -37936 6823
rect -38757 6795 -37936 6819
rect -37880 6795 -37772 6851
rect -38757 6542 -37772 6795
rect -31724 8147 -30705 8360
rect -31724 8131 -31413 8147
rect -31724 8075 -31601 8131
rect -31545 8091 -31413 8131
rect -31357 8091 -30705 8147
rect -31545 8075 -30705 8091
rect -31724 7996 -30705 8075
rect -31724 7962 -31150 7996
rect -31724 7954 -31384 7962
rect -31724 7898 -31585 7954
rect -31529 7906 -31384 7954
rect -31328 7940 -31150 7962
rect -31094 7940 -30705 7996
rect -31328 7934 -30705 7940
rect -31328 7906 -30963 7934
rect -31529 7898 -30963 7906
rect -31724 7878 -30963 7898
rect -30907 7878 -30705 7934
rect -31724 7786 -30705 7878
rect -31724 7773 -31367 7786
rect -31724 7717 -31581 7773
rect -31525 7730 -31367 7773
rect -31311 7777 -30705 7786
rect -31311 7730 -31150 7777
rect -31525 7721 -31150 7730
rect -31094 7749 -30705 7777
rect -31094 7721 -30920 7749
rect -31525 7717 -30920 7721
rect -31724 7693 -30920 7717
rect -30864 7693 -30705 7749
rect -31724 7255 -30705 7693
rect -31724 7239 -31396 7255
rect -31724 7183 -31584 7239
rect -31528 7199 -31396 7239
rect -31340 7199 -30705 7255
rect -31528 7183 -30705 7199
rect -31724 7104 -30705 7183
rect -31724 7070 -31133 7104
rect -31724 7062 -31367 7070
rect -31724 7006 -31568 7062
rect -31512 7014 -31367 7062
rect -31311 7048 -31133 7070
rect -31077 7048 -30705 7104
rect -31311 7042 -30705 7048
rect -31311 7014 -30946 7042
rect -31512 7006 -30946 7014
rect -31724 6986 -30946 7006
rect -30890 6986 -30705 7042
rect -31724 6894 -30705 6986
rect -31724 6881 -31350 6894
rect -31724 6825 -31564 6881
rect -31508 6838 -31350 6881
rect -31294 6885 -30705 6894
rect -31294 6838 -31133 6885
rect -31508 6829 -31133 6838
rect -31077 6857 -30705 6885
rect -31077 6829 -30903 6857
rect -31508 6825 -30903 6829
rect -31724 6801 -30903 6825
rect -30847 6801 -30705 6857
rect -31724 6507 -30705 6801
rect -24931 8024 -23912 8238
rect -24931 8008 -24562 8024
rect -24931 7952 -24750 8008
rect -24694 7968 -24562 8008
rect -24506 7968 -23912 8024
rect -24694 7952 -23912 7968
rect -24931 7873 -23912 7952
rect -24931 7839 -24299 7873
rect -24931 7831 -24533 7839
rect -24931 7775 -24734 7831
rect -24678 7783 -24533 7831
rect -24477 7817 -24299 7839
rect -24243 7817 -23912 7873
rect -24477 7811 -23912 7817
rect -24477 7783 -24112 7811
rect -24678 7775 -24112 7783
rect -24931 7755 -24112 7775
rect -24056 7755 -23912 7811
rect -24931 7663 -23912 7755
rect -24931 7650 -24516 7663
rect -24931 7594 -24730 7650
rect -24674 7607 -24516 7650
rect -24460 7654 -23912 7663
rect -24460 7607 -24299 7654
rect -24674 7598 -24299 7607
rect -24243 7626 -23912 7654
rect -24243 7598 -24069 7626
rect -24674 7594 -24069 7598
rect -24931 7570 -24069 7594
rect -24013 7570 -23912 7626
rect -24931 7191 -23912 7570
rect -24931 7175 -24573 7191
rect -24931 7119 -24761 7175
rect -24705 7135 -24573 7175
rect -24517 7135 -23912 7191
rect -24705 7119 -23912 7135
rect -24931 7040 -23912 7119
rect -24931 7006 -24310 7040
rect -24931 6998 -24544 7006
rect -24931 6942 -24745 6998
rect -24689 6950 -24544 6998
rect -24488 6984 -24310 7006
rect -24254 6984 -23912 7040
rect -24488 6978 -23912 6984
rect -24488 6950 -24123 6978
rect -24689 6942 -24123 6950
rect -24931 6922 -24123 6942
rect -24067 6922 -23912 6978
rect -24931 6830 -23912 6922
rect -24931 6817 -24527 6830
rect -24931 6761 -24741 6817
rect -24685 6774 -24527 6817
rect -24471 6821 -23912 6830
rect -24471 6774 -24310 6821
rect -24685 6765 -24310 6774
rect -24254 6793 -23912 6821
rect -24254 6765 -24080 6793
rect -24685 6761 -24080 6765
rect -24931 6737 -24080 6761
rect -24024 6737 -23912 6793
rect -24931 6385 -23912 6737
rect -18061 8106 -17042 8354
rect -18061 8090 -17727 8106
rect -18061 8034 -17915 8090
rect -17859 8050 -17727 8090
rect -17671 8050 -17042 8106
rect -17859 8034 -17042 8050
rect -18061 7955 -17042 8034
rect -18061 7921 -17464 7955
rect -18061 7913 -17698 7921
rect -18061 7857 -17899 7913
rect -17843 7865 -17698 7913
rect -17642 7899 -17464 7921
rect -17408 7899 -17042 7955
rect -17642 7893 -17042 7899
rect -17642 7865 -17277 7893
rect -17843 7857 -17277 7865
rect -18061 7837 -17277 7857
rect -17221 7837 -17042 7893
rect -18061 7745 -17042 7837
rect -18061 7732 -17681 7745
rect -18061 7676 -17895 7732
rect -17839 7689 -17681 7732
rect -17625 7736 -17042 7745
rect -17625 7689 -17464 7736
rect -17839 7680 -17464 7689
rect -17408 7708 -17042 7736
rect -17408 7680 -17234 7708
rect -17839 7676 -17234 7680
rect -18061 7652 -17234 7676
rect -17178 7652 -17042 7708
rect -18061 7249 -17042 7652
rect -18061 7233 -17727 7249
rect -18061 7177 -17915 7233
rect -17859 7193 -17727 7233
rect -17671 7193 -17042 7249
rect -17859 7177 -17042 7193
rect -18061 7098 -17042 7177
rect -18061 7064 -17464 7098
rect -18061 7056 -17698 7064
rect -18061 7000 -17899 7056
rect -17843 7008 -17698 7056
rect -17642 7042 -17464 7064
rect -17408 7042 -17042 7098
rect -17642 7036 -17042 7042
rect -17642 7008 -17277 7036
rect -17843 7000 -17277 7008
rect -18061 6980 -17277 7000
rect -17221 6980 -17042 7036
rect -18061 6888 -17042 6980
rect -18061 6875 -17681 6888
rect -18061 6819 -17895 6875
rect -17839 6832 -17681 6875
rect -17625 6879 -17042 6888
rect -17625 6832 -17464 6879
rect -17839 6823 -17464 6832
rect -17408 6851 -17042 6879
rect -17408 6823 -17234 6851
rect -17839 6819 -17234 6823
rect -18061 6795 -17234 6819
rect -17178 6795 -17042 6851
rect -18061 6501 -17042 6795
rect -11069 8193 -10050 8319
rect -11069 8177 -10735 8193
rect -11069 8121 -10923 8177
rect -10867 8137 -10735 8177
rect -10679 8137 -10050 8193
rect -10867 8121 -10050 8137
rect -11069 8042 -10050 8121
rect -11069 8008 -10472 8042
rect -11069 8000 -10706 8008
rect -11069 7944 -10907 8000
rect -10851 7952 -10706 8000
rect -10650 7986 -10472 8008
rect -10416 7986 -10050 8042
rect -10650 7980 -10050 7986
rect -10650 7952 -10285 7980
rect -10851 7944 -10285 7952
rect -11069 7924 -10285 7944
rect -10229 7924 -10050 7980
rect -11069 7832 -10050 7924
rect -11069 7819 -10689 7832
rect -11069 7763 -10903 7819
rect -10847 7776 -10689 7819
rect -10633 7823 -10050 7832
rect -10633 7776 -10472 7823
rect -10847 7767 -10472 7776
rect -10416 7795 -10050 7823
rect -10416 7767 -10242 7795
rect -10847 7763 -10242 7767
rect -11069 7739 -10242 7763
rect -10186 7739 -10050 7795
rect -11069 7208 -10050 7739
rect -11069 7192 -10712 7208
rect -11069 7136 -10900 7192
rect -10844 7152 -10712 7192
rect -10656 7152 -10050 7208
rect -10844 7136 -10050 7152
rect -11069 7057 -10050 7136
rect -11069 7023 -10449 7057
rect -11069 7015 -10683 7023
rect -11069 6959 -10884 7015
rect -10828 6967 -10683 7015
rect -10627 7001 -10449 7023
rect -10393 7001 -10050 7057
rect -10627 6995 -10050 7001
rect -10627 6967 -10262 6995
rect -10828 6959 -10262 6967
rect -11069 6939 -10262 6959
rect -10206 6939 -10050 6995
rect -11069 6847 -10050 6939
rect -11069 6834 -10666 6847
rect -11069 6778 -10880 6834
rect -10824 6791 -10666 6834
rect -10610 6838 -10050 6847
rect -10610 6791 -10449 6838
rect -10824 6782 -10449 6791
rect -10393 6810 -10050 6838
rect -10393 6782 -10219 6810
rect -10824 6778 -10219 6782
rect -11069 6754 -10219 6778
rect -10163 6754 -10050 6810
rect -11069 6466 -10050 6754
rect -3635 8211 -2616 8337
rect -3635 8195 -3295 8211
rect -3635 8139 -3483 8195
rect -3427 8155 -3295 8195
rect -3239 8155 -2616 8211
rect -3427 8139 -2616 8155
rect -3635 8060 -2616 8139
rect -3635 8026 -3032 8060
rect -3635 8018 -3266 8026
rect -3635 7962 -3467 8018
rect -3411 7970 -3266 8018
rect -3210 8004 -3032 8026
rect -2976 8004 -2616 8060
rect -3210 7998 -2616 8004
rect -3210 7970 -2845 7998
rect -3411 7962 -2845 7970
rect -3635 7942 -2845 7962
rect -2789 7942 -2616 7998
rect -3635 7850 -2616 7942
rect -3635 7837 -3249 7850
rect -3635 7781 -3463 7837
rect -3407 7794 -3249 7837
rect -3193 7841 -2616 7850
rect -3193 7794 -3032 7841
rect -3407 7785 -3032 7794
rect -2976 7813 -2616 7841
rect -2976 7785 -2802 7813
rect -3407 7781 -2802 7785
rect -3635 7757 -2802 7781
rect -2746 7757 -2616 7813
rect -3635 7238 -2616 7757
rect -3635 7222 -3225 7238
rect -3635 7166 -3413 7222
rect -3357 7182 -3225 7222
rect -3169 7182 -2616 7238
rect -3357 7166 -2616 7182
rect -3635 7087 -2616 7166
rect -3635 7053 -2962 7087
rect -3635 7045 -3196 7053
rect -3635 6989 -3397 7045
rect -3341 6997 -3196 7045
rect -3140 7031 -2962 7053
rect -2906 7031 -2616 7087
rect -3140 7025 -2616 7031
rect -3140 6997 -2775 7025
rect -3341 6989 -2775 6997
rect -3635 6969 -2775 6989
rect -2719 6969 -2616 7025
rect -3635 6877 -2616 6969
rect -3635 6864 -3179 6877
rect -3635 6808 -3393 6864
rect -3337 6821 -3179 6864
rect -3123 6868 -2616 6877
rect -3123 6821 -2962 6868
rect -3337 6812 -2962 6821
rect -2906 6840 -2616 6868
rect -2906 6812 -2732 6840
rect -3337 6808 -2732 6812
rect -3635 6784 -2732 6808
rect -2676 6784 -2616 6840
rect -3635 6484 -2616 6784
rect 2058 8164 3077 8290
rect 2058 8148 2415 8164
rect 2058 8092 2227 8148
rect 2283 8108 2415 8148
rect 2471 8108 3077 8164
rect 2283 8092 3077 8108
rect 2058 8013 3077 8092
rect 2058 7979 2678 8013
rect 2058 7971 2444 7979
rect 2058 7915 2243 7971
rect 2299 7923 2444 7971
rect 2500 7957 2678 7979
rect 2734 7957 3077 8013
rect 2500 7951 3077 7957
rect 2500 7923 2865 7951
rect 2299 7915 2865 7923
rect 2058 7895 2865 7915
rect 2921 7895 3077 7951
rect 2058 7803 3077 7895
rect 2058 7790 2461 7803
rect 2058 7734 2247 7790
rect 2303 7747 2461 7790
rect 2517 7794 3077 7803
rect 2517 7747 2678 7794
rect 2303 7738 2678 7747
rect 2734 7766 3077 7794
rect 2734 7738 2908 7766
rect 2303 7734 2908 7738
rect 2058 7710 2908 7734
rect 2964 7710 3077 7766
rect 2058 7139 3077 7710
rect 2058 7123 2444 7139
rect 2058 7067 2256 7123
rect 2312 7083 2444 7123
rect 2500 7083 3077 7139
rect 2312 7067 3077 7083
rect 2058 6988 3077 7067
rect 2058 6954 2707 6988
rect 2058 6946 2473 6954
rect 2058 6890 2272 6946
rect 2328 6898 2473 6946
rect 2529 6932 2707 6954
rect 2763 6932 3077 6988
rect 2529 6926 3077 6932
rect 2529 6898 2894 6926
rect 2328 6890 2894 6898
rect 2058 6870 2894 6890
rect 2950 6870 3077 6926
rect 2058 6778 3077 6870
rect 2058 6765 2490 6778
rect 2058 6709 2276 6765
rect 2332 6722 2490 6765
rect 2546 6769 3077 6778
rect 2546 6722 2707 6769
rect 2332 6713 2707 6722
rect 2763 6741 3077 6769
rect 2763 6713 2937 6741
rect 2332 6709 2937 6713
rect 2058 6685 2937 6709
rect 2993 6685 3077 6741
rect 2058 6437 3077 6685
rect -61751 -68320 -60887 -68247
rect -61751 -68336 -61490 -68320
rect -61751 -68392 -61678 -68336
rect -61622 -68376 -61490 -68336
rect -61434 -68376 -60887 -68320
rect -61622 -68392 -60887 -68376
rect -61751 -68471 -60887 -68392
rect -61751 -68505 -61227 -68471
rect -61751 -68513 -61461 -68505
rect -61751 -68569 -61662 -68513
rect -61606 -68561 -61461 -68513
rect -61405 -68527 -61227 -68505
rect -61171 -68527 -60887 -68471
rect -61405 -68533 -60887 -68527
rect -61405 -68561 -61040 -68533
rect -61606 -68569 -61040 -68561
rect -61751 -68589 -61040 -68569
rect -60984 -68589 -60887 -68533
rect -61751 -68681 -60887 -68589
rect -61751 -68694 -61444 -68681
rect -61751 -68750 -61658 -68694
rect -61602 -68737 -61444 -68694
rect -61388 -68690 -60887 -68681
rect -61388 -68737 -61227 -68690
rect -61602 -68746 -61227 -68737
rect -61171 -68718 -60887 -68690
rect -61171 -68746 -60997 -68718
rect -61602 -68750 -60997 -68746
rect -61751 -68774 -60997 -68750
rect -60941 -68774 -60887 -68718
rect -61751 -68934 -60887 -68774
rect -55242 -68379 -54186 -68282
rect -55242 -68435 -54944 -68379
rect -54888 -68435 -54769 -68379
rect -54713 -68435 -54567 -68379
rect -54511 -68435 -54186 -68379
rect -55242 -68619 -54186 -68435
rect -55242 -68644 -54725 -68619
rect -55242 -68646 -54925 -68644
rect -55242 -68702 -55157 -68646
rect -55101 -68700 -54925 -68646
rect -54869 -68675 -54725 -68644
rect -54669 -68634 -54186 -68619
rect -54669 -68650 -54294 -68634
rect -54669 -68675 -54507 -68650
rect -54869 -68700 -54507 -68675
rect -55101 -68702 -54507 -68700
rect -55242 -68706 -54507 -68702
rect -54451 -68690 -54294 -68650
rect -54238 -68690 -54186 -68634
rect -54451 -68706 -54186 -68690
rect -55242 -68863 -54186 -68706
rect -55242 -68867 -54696 -68863
rect -55242 -68923 -54921 -68867
rect -54865 -68919 -54696 -68867
rect -54640 -68869 -54186 -68863
rect -54640 -68919 -54438 -68869
rect -54865 -68923 -54438 -68919
rect -55242 -68925 -54438 -68923
rect -54382 -68925 -54186 -68869
rect -48439 -68369 -47230 -68311
rect -48439 -68425 -48168 -68369
rect -48112 -68425 -47987 -68369
rect -47931 -68375 -47230 -68369
rect -47931 -68425 -47783 -68375
rect -48439 -68431 -47783 -68425
rect -47727 -68431 -47230 -68375
rect -48439 -68569 -47230 -68431
rect -48439 -68575 -47916 -68569
rect -48439 -68631 -48152 -68575
rect -48096 -68625 -47916 -68575
rect -47860 -68584 -47230 -68569
rect -47860 -68625 -47656 -68584
rect -48096 -68631 -47656 -68625
rect -48439 -68640 -47656 -68631
rect -47600 -68640 -47230 -68584
rect -48439 -68786 -47230 -68640
rect -48439 -68842 -48212 -68786
rect -48156 -68790 -47230 -68786
rect -48156 -68842 -47970 -68790
rect -48439 -68846 -47970 -68842
rect -47914 -68846 -47770 -68790
rect -47714 -68800 -47230 -68790
rect -47714 -68846 -47466 -68800
rect -48439 -68856 -47466 -68846
rect -47410 -68856 -47230 -68800
rect -48439 -68909 -47230 -68856
rect -41649 -68369 -40440 -68326
rect -21096 -68350 -20092 -68263
rect -41649 -68373 -41151 -68369
rect -41649 -68429 -41332 -68373
rect -41276 -68425 -41151 -68373
rect -41095 -68379 -40440 -68369
rect -41095 -68425 -40951 -68379
rect -41276 -68429 -40951 -68425
rect -41649 -68435 -40951 -68429
rect -40895 -68435 -40440 -68379
rect -41649 -68542 -40440 -68435
rect -41649 -68581 -41330 -68542
rect -41649 -68637 -41517 -68581
rect -41461 -68598 -41330 -68581
rect -41274 -68546 -40440 -68542
rect -41274 -68556 -40890 -68546
rect -41274 -68598 -41117 -68556
rect -41461 -68612 -41117 -68598
rect -41061 -68602 -40890 -68556
rect -40834 -68569 -40440 -68546
rect -40834 -68602 -40694 -68569
rect -41061 -68612 -40694 -68602
rect -41461 -68625 -40694 -68612
rect -40638 -68625 -40440 -68569
rect -41461 -68637 -40440 -68625
rect -41649 -68742 -40440 -68637
rect -41649 -68759 -41084 -68742
rect -41649 -68815 -41317 -68759
rect -41261 -68798 -41084 -68759
rect -41028 -68754 -40440 -68742
rect -41028 -68798 -40836 -68754
rect -41261 -68810 -40836 -68798
rect -40780 -68810 -40440 -68754
rect -41261 -68815 -40440 -68810
rect -41649 -68924 -40440 -68815
rect -34904 -68408 -33695 -68353
rect -34904 -68464 -34577 -68408
rect -34521 -68415 -33695 -68408
rect -34521 -68464 -34396 -68415
rect -34904 -68471 -34396 -68464
rect -34340 -68471 -34221 -68415
rect -34165 -68471 -33695 -68415
rect -34904 -68625 -33695 -68471
rect -34904 -68631 -34000 -68625
rect -34904 -68650 -34560 -68631
rect -34904 -68706 -34819 -68650
rect -34763 -68687 -34560 -68650
rect -34504 -68687 -34329 -68631
rect -34273 -68681 -34000 -68631
rect -33944 -68681 -33695 -68625
rect -34273 -68687 -33695 -68681
rect -34763 -68706 -33695 -68687
rect -34904 -68834 -33695 -68706
rect -34904 -68848 -33843 -68834
rect -34904 -68904 -34581 -68848
rect -34525 -68904 -34346 -68848
rect -34290 -68852 -33843 -68848
rect -34290 -68904 -34106 -68852
rect -34904 -68908 -34106 -68904
rect -34050 -68890 -33843 -68852
rect -33787 -68890 -33695 -68834
rect -34050 -68908 -33695 -68890
rect -55242 -68970 -54186 -68925
rect -34904 -68951 -33695 -68908
rect -28030 -68388 -26900 -68350
rect -28030 -68444 -27727 -68388
rect -27671 -68395 -26900 -68388
rect -27671 -68444 -27546 -68395
rect -28030 -68451 -27546 -68444
rect -27490 -68451 -27371 -68395
rect -27315 -68451 -26900 -68395
rect -28030 -68605 -26900 -68451
rect -28030 -68611 -27150 -68605
rect -28030 -68630 -27710 -68611
rect -28030 -68686 -27969 -68630
rect -27913 -68667 -27710 -68630
rect -27654 -68667 -27479 -68611
rect -27423 -68661 -27150 -68611
rect -27094 -68661 -26900 -68605
rect -27423 -68667 -26900 -68661
rect -27913 -68686 -26900 -68667
rect -28030 -68814 -26900 -68686
rect -28030 -68828 -26993 -68814
rect -28030 -68884 -27731 -68828
rect -27675 -68884 -27496 -68828
rect -27440 -68832 -26993 -68828
rect -27440 -68884 -27256 -68832
rect -28030 -68888 -27256 -68884
rect -27200 -68870 -26993 -68832
rect -26937 -68870 -26900 -68814
rect -27200 -68888 -26900 -68870
rect -28030 -68930 -26900 -68888
rect -21096 -68388 -19960 -68350
rect -21096 -68444 -20787 -68388
rect -20731 -68395 -19960 -68388
rect -20731 -68444 -20606 -68395
rect -21096 -68451 -20606 -68444
rect -20550 -68451 -20431 -68395
rect -20375 -68451 -19960 -68395
rect -21096 -68605 -19960 -68451
rect -21096 -68611 -20210 -68605
rect -21096 -68630 -20770 -68611
rect -21096 -68686 -21029 -68630
rect -20973 -68667 -20770 -68630
rect -20714 -68667 -20539 -68611
rect -20483 -68661 -20210 -68611
rect -20154 -68661 -19960 -68605
rect -20483 -68667 -19960 -68661
rect -20973 -68686 -19960 -68667
rect -21096 -68814 -19960 -68686
rect -21096 -68828 -20053 -68814
rect -21096 -68884 -20791 -68828
rect -20735 -68884 -20556 -68828
rect -20500 -68832 -20053 -68828
rect -20500 -68884 -20316 -68832
rect -21096 -68888 -20316 -68884
rect -20260 -68870 -20053 -68832
rect -19997 -68870 -19960 -68814
rect -20260 -68888 -19960 -68870
rect -21096 -68930 -19960 -68888
rect -14409 -68381 -13405 -68255
rect -14409 -68437 -14124 -68381
rect -14068 -68386 -13405 -68381
rect -14068 -68437 -13945 -68386
rect -14409 -68442 -13945 -68437
rect -13889 -68442 -13762 -68386
rect -13706 -68442 -13405 -68386
rect -14409 -68634 -13405 -68442
rect -14409 -68638 -13637 -68634
rect -14409 -68644 -13845 -68638
rect -14409 -68650 -14037 -68644
rect -14409 -68706 -14262 -68650
rect -14206 -68700 -14037 -68650
rect -13981 -68694 -13845 -68644
rect -13789 -68690 -13637 -68638
rect -13581 -68690 -13405 -68634
rect -13789 -68694 -13405 -68690
rect -13981 -68700 -13405 -68694
rect -14206 -68706 -13405 -68700
rect -14409 -68848 -13405 -68706
rect -14409 -68904 -14199 -68848
rect -14143 -68904 -13980 -68848
rect -13924 -68904 -13791 -68848
rect -13735 -68904 -13543 -68848
rect -13487 -68904 -13405 -68848
rect -21096 -68951 -20092 -68930
rect -14409 -68943 -13405 -68904
rect -7481 -68361 -6477 -68255
rect -7481 -68417 -7286 -68361
rect -7230 -68417 -7111 -68361
rect -7055 -68417 -6921 -68361
rect -6865 -68417 -6477 -68361
rect -7481 -68611 -6477 -68417
rect -7481 -68617 -6648 -68611
rect -7481 -68623 -6909 -68617
rect -7481 -68629 -7129 -68623
rect -7481 -68685 -7402 -68629
rect -7346 -68679 -7129 -68629
rect -7073 -68673 -6909 -68623
rect -6853 -68667 -6648 -68617
rect -6592 -68667 -6477 -68611
rect -6853 -68673 -6477 -68667
rect -7073 -68679 -6477 -68673
rect -7346 -68685 -6477 -68679
rect -7481 -68846 -6477 -68685
rect -7481 -68852 -6723 -68846
rect -7481 -68854 -7152 -68852
rect -7481 -68910 -7367 -68854
rect -7311 -68908 -7152 -68854
rect -7096 -68908 -6934 -68852
rect -6878 -68902 -6723 -68852
rect -6667 -68902 -6477 -68846
rect -6878 -68908 -6477 -68902
rect -7311 -68910 -6477 -68908
rect -7481 -68943 -6477 -68910
rect -676 -68358 328 -68259
rect -676 -68361 -70 -68358
rect -676 -68417 -476 -68361
rect -420 -68365 -70 -68361
rect -420 -68417 -283 -68365
rect -676 -68421 -283 -68417
rect -227 -68414 -70 -68365
rect -14 -68414 328 -68358
rect -227 -68421 328 -68414
rect -676 -68594 328 -68421
rect -676 -68598 145 -68594
rect -676 -68602 -345 -68598
rect -676 -68658 -595 -68602
rect -539 -68654 -345 -68602
rect -289 -68654 -112 -68598
rect -56 -68650 145 -68598
rect 201 -68650 328 -68594
rect -56 -68654 328 -68650
rect -539 -68658 328 -68654
rect -676 -68848 328 -68658
rect -676 -68852 -308 -68848
rect -676 -68908 -566 -68852
rect -510 -68904 -308 -68852
rect -252 -68852 328 -68848
rect -252 -68904 -70 -68852
rect -510 -68908 -70 -68904
rect -14 -68859 328 -68852
rect -14 -68908 184 -68859
rect -676 -68915 184 -68908
rect 240 -68915 328 -68859
rect -676 -68947 328 -68915
rect 5835 -68352 6839 -68257
rect 5835 -68408 6318 -68352
rect 6374 -68408 6506 -68352
rect 6562 -68358 6839 -68352
rect 6562 -68408 6708 -68358
rect 5835 -68414 6708 -68408
rect 6764 -68414 6839 -68358
rect 5835 -68573 6839 -68414
rect 5835 -68629 6143 -68573
rect 6199 -68577 6606 -68573
rect 6199 -68629 6395 -68577
rect 5835 -68633 6395 -68629
rect 6451 -68629 6606 -68577
rect 6662 -68629 6839 -68573
rect 6451 -68633 6839 -68629
rect 5835 -68688 6839 -68633
rect 5835 -68744 5931 -68688
rect 5987 -68744 6839 -68688
rect 5835 -68852 6839 -68744
rect 5835 -68854 6327 -68852
rect 5835 -68910 6139 -68854
rect 6195 -68908 6327 -68854
rect 6383 -68908 6533 -68852
rect 6589 -68854 6839 -68852
rect 6589 -68908 6737 -68854
rect 6195 -68910 6737 -68908
rect 6793 -68910 6839 -68854
rect 5835 -68945 6839 -68910
<< via2 >>
rect -51678 8302 -51622 8304
rect -51866 8286 -51810 8288
rect -51866 8234 -51864 8286
rect -51864 8234 -51812 8286
rect -51812 8234 -51810 8286
rect -51678 8250 -51676 8302
rect -51676 8250 -51624 8302
rect -51624 8250 -51622 8302
rect -51678 8248 -51622 8250
rect -51866 8232 -51810 8234
rect -64935 7981 -64879 7983
rect -65123 7965 -65067 7967
rect -65123 7913 -65121 7965
rect -65121 7913 -65069 7965
rect -65069 7913 -65067 7965
rect -64935 7929 -64933 7981
rect -64933 7929 -64881 7981
rect -64881 7929 -64879 7981
rect -64935 7927 -64879 7929
rect -65123 7911 -65067 7913
rect -64672 7830 -64616 7832
rect -64906 7796 -64850 7798
rect -65107 7788 -65051 7790
rect -65107 7736 -65105 7788
rect -65105 7736 -65053 7788
rect -65053 7736 -65051 7788
rect -64906 7744 -64904 7796
rect -64904 7744 -64852 7796
rect -64852 7744 -64850 7796
rect -64672 7778 -64670 7830
rect -64670 7778 -64618 7830
rect -64618 7778 -64616 7830
rect -64672 7776 -64616 7778
rect -64906 7742 -64850 7744
rect -64485 7768 -64429 7770
rect -65107 7734 -65051 7736
rect -64485 7716 -64483 7768
rect -64483 7716 -64431 7768
rect -64431 7716 -64429 7768
rect -64485 7714 -64429 7716
rect -64889 7620 -64833 7622
rect -65103 7607 -65047 7609
rect -65103 7555 -65101 7607
rect -65101 7555 -65049 7607
rect -65049 7555 -65047 7607
rect -64889 7568 -64887 7620
rect -64887 7568 -64835 7620
rect -64835 7568 -64833 7620
rect -64889 7566 -64833 7568
rect -64672 7611 -64616 7613
rect -64672 7559 -64670 7611
rect -64670 7559 -64618 7611
rect -64618 7559 -64616 7611
rect -64672 7557 -64616 7559
rect -64442 7583 -64386 7585
rect -65103 7553 -65047 7555
rect -64442 7531 -64440 7583
rect -64440 7531 -64388 7583
rect -64388 7531 -64386 7583
rect -64442 7529 -64386 7531
rect -64958 7163 -64902 7165
rect -65146 7147 -65090 7149
rect -65146 7095 -65144 7147
rect -65144 7095 -65092 7147
rect -65092 7095 -65090 7147
rect -64958 7111 -64956 7163
rect -64956 7111 -64904 7163
rect -64904 7111 -64902 7163
rect -64958 7109 -64902 7111
rect -65146 7093 -65090 7095
rect -64695 7012 -64639 7014
rect -64929 6978 -64873 6980
rect -65130 6970 -65074 6972
rect -65130 6918 -65128 6970
rect -65128 6918 -65076 6970
rect -65076 6918 -65074 6970
rect -64929 6926 -64927 6978
rect -64927 6926 -64875 6978
rect -64875 6926 -64873 6978
rect -64695 6960 -64693 7012
rect -64693 6960 -64641 7012
rect -64641 6960 -64639 7012
rect -64695 6958 -64639 6960
rect -64929 6924 -64873 6926
rect -64508 6950 -64452 6952
rect -65130 6916 -65074 6918
rect -64508 6898 -64506 6950
rect -64506 6898 -64454 6950
rect -64454 6898 -64452 6950
rect -64508 6896 -64452 6898
rect -64912 6802 -64856 6804
rect -65126 6789 -65070 6791
rect -65126 6737 -65124 6789
rect -65124 6737 -65072 6789
rect -65072 6737 -65070 6789
rect -64912 6750 -64910 6802
rect -64910 6750 -64858 6802
rect -64858 6750 -64856 6802
rect -64912 6748 -64856 6750
rect -64695 6793 -64639 6795
rect -64695 6741 -64693 6793
rect -64693 6741 -64641 6793
rect -64641 6741 -64639 6793
rect -64695 6739 -64639 6741
rect -64465 6765 -64409 6767
rect -65126 6735 -65070 6737
rect -64465 6713 -64463 6765
rect -64463 6713 -64411 6765
rect -64411 6713 -64409 6765
rect -64465 6711 -64409 6713
rect -58740 8063 -58684 8065
rect -58928 8047 -58872 8049
rect -58928 7995 -58926 8047
rect -58926 7995 -58874 8047
rect -58874 7995 -58872 8047
rect -58740 8011 -58738 8063
rect -58738 8011 -58686 8063
rect -58686 8011 -58684 8063
rect -58740 8009 -58684 8011
rect -58928 7993 -58872 7995
rect -58477 7912 -58421 7914
rect -58711 7878 -58655 7880
rect -58912 7870 -58856 7872
rect -58912 7818 -58910 7870
rect -58910 7818 -58858 7870
rect -58858 7818 -58856 7870
rect -58711 7826 -58709 7878
rect -58709 7826 -58657 7878
rect -58657 7826 -58655 7878
rect -58477 7860 -58475 7912
rect -58475 7860 -58423 7912
rect -58423 7860 -58421 7912
rect -58477 7858 -58421 7860
rect -58711 7824 -58655 7826
rect -58290 7850 -58234 7852
rect -58912 7816 -58856 7818
rect -58290 7798 -58288 7850
rect -58288 7798 -58236 7850
rect -58236 7798 -58234 7850
rect -58290 7796 -58234 7798
rect -58694 7702 -58638 7704
rect -58908 7689 -58852 7691
rect -58908 7637 -58906 7689
rect -58906 7637 -58854 7689
rect -58854 7637 -58852 7689
rect -58694 7650 -58692 7702
rect -58692 7650 -58640 7702
rect -58640 7650 -58638 7702
rect -58694 7648 -58638 7650
rect -58477 7693 -58421 7695
rect -58477 7641 -58475 7693
rect -58475 7641 -58423 7693
rect -58423 7641 -58421 7693
rect -58477 7639 -58421 7641
rect -58247 7665 -58191 7667
rect -58908 7635 -58852 7637
rect -58247 7613 -58245 7665
rect -58245 7613 -58193 7665
rect -58193 7613 -58191 7665
rect -58247 7611 -58191 7613
rect -58740 7183 -58684 7185
rect -58928 7167 -58872 7169
rect -58928 7115 -58926 7167
rect -58926 7115 -58874 7167
rect -58874 7115 -58872 7167
rect -58740 7131 -58738 7183
rect -58738 7131 -58686 7183
rect -58686 7131 -58684 7183
rect -58740 7129 -58684 7131
rect -58928 7113 -58872 7115
rect -58477 7032 -58421 7034
rect -58711 6998 -58655 7000
rect -58912 6990 -58856 6992
rect -58912 6938 -58910 6990
rect -58910 6938 -58858 6990
rect -58858 6938 -58856 6990
rect -58711 6946 -58709 6998
rect -58709 6946 -58657 6998
rect -58657 6946 -58655 6998
rect -58477 6980 -58475 7032
rect -58475 6980 -58423 7032
rect -58423 6980 -58421 7032
rect -58477 6978 -58421 6980
rect -58711 6944 -58655 6946
rect -58290 6970 -58234 6972
rect -58912 6936 -58856 6938
rect -58290 6918 -58288 6970
rect -58288 6918 -58236 6970
rect -58236 6918 -58234 6970
rect -58290 6916 -58234 6918
rect -58694 6822 -58638 6824
rect -58908 6809 -58852 6811
rect -58908 6757 -58906 6809
rect -58906 6757 -58854 6809
rect -58854 6757 -58852 6809
rect -58694 6770 -58692 6822
rect -58692 6770 -58640 6822
rect -58640 6770 -58638 6822
rect -58694 6768 -58638 6770
rect -58477 6813 -58421 6815
rect -58477 6761 -58475 6813
rect -58475 6761 -58423 6813
rect -58423 6761 -58421 6813
rect -58477 6759 -58421 6761
rect -58247 6785 -58191 6787
rect -58908 6755 -58852 6757
rect -58247 6733 -58245 6785
rect -58245 6733 -58193 6785
rect -58193 6733 -58191 6785
rect -58247 6731 -58191 6733
rect -51415 8151 -51359 8153
rect -51649 8117 -51593 8119
rect -51850 8109 -51794 8111
rect -51850 8057 -51848 8109
rect -51848 8057 -51796 8109
rect -51796 8057 -51794 8109
rect -51649 8065 -51647 8117
rect -51647 8065 -51595 8117
rect -51595 8065 -51593 8117
rect -51415 8099 -51413 8151
rect -51413 8099 -51361 8151
rect -51361 8099 -51359 8151
rect -51415 8097 -51359 8099
rect -51649 8063 -51593 8065
rect -51228 8089 -51172 8091
rect -51850 8055 -51794 8057
rect -51228 8037 -51226 8089
rect -51226 8037 -51174 8089
rect -51174 8037 -51172 8089
rect -51228 8035 -51172 8037
rect -51632 7941 -51576 7943
rect -51846 7928 -51790 7930
rect -51846 7876 -51844 7928
rect -51844 7876 -51792 7928
rect -51792 7876 -51790 7928
rect -51632 7889 -51630 7941
rect -51630 7889 -51578 7941
rect -51578 7889 -51576 7941
rect -51632 7887 -51576 7889
rect -51415 7932 -51359 7934
rect -51415 7880 -51413 7932
rect -51413 7880 -51361 7932
rect -51361 7880 -51359 7932
rect -51415 7878 -51359 7880
rect -51185 7904 -51129 7906
rect -51846 7874 -51790 7876
rect -51185 7852 -51183 7904
rect -51183 7852 -51131 7904
rect -51131 7852 -51129 7904
rect -51185 7850 -51129 7852
rect -51698 7436 -51642 7438
rect -51886 7420 -51830 7422
rect -51886 7368 -51884 7420
rect -51884 7368 -51832 7420
rect -51832 7368 -51830 7420
rect -51698 7384 -51696 7436
rect -51696 7384 -51644 7436
rect -51644 7384 -51642 7436
rect -51698 7382 -51642 7384
rect -51886 7366 -51830 7368
rect -51435 7285 -51379 7287
rect -51669 7251 -51613 7253
rect -51870 7243 -51814 7245
rect -51870 7191 -51868 7243
rect -51868 7191 -51816 7243
rect -51816 7191 -51814 7243
rect -51669 7199 -51667 7251
rect -51667 7199 -51615 7251
rect -51615 7199 -51613 7251
rect -51435 7233 -51433 7285
rect -51433 7233 -51381 7285
rect -51381 7233 -51379 7285
rect -51435 7231 -51379 7233
rect -51669 7197 -51613 7199
rect -51248 7223 -51192 7225
rect -51870 7189 -51814 7191
rect -51248 7171 -51246 7223
rect -51246 7171 -51194 7223
rect -51194 7171 -51192 7223
rect -51248 7169 -51192 7171
rect -51652 7075 -51596 7077
rect -51866 7062 -51810 7064
rect -51866 7010 -51864 7062
rect -51864 7010 -51812 7062
rect -51812 7010 -51810 7062
rect -51652 7023 -51650 7075
rect -51650 7023 -51598 7075
rect -51598 7023 -51596 7075
rect -51652 7021 -51596 7023
rect -51435 7066 -51379 7068
rect -51435 7014 -51433 7066
rect -51433 7014 -51381 7066
rect -51381 7014 -51379 7066
rect -51435 7012 -51379 7014
rect -51205 7038 -51149 7040
rect -51866 7008 -51810 7010
rect -51205 6986 -51203 7038
rect -51203 6986 -51151 7038
rect -51151 6986 -51149 7038
rect -51205 6984 -51149 6986
rect -45141 8156 -45085 8158
rect -45329 8140 -45273 8142
rect -45329 8088 -45327 8140
rect -45327 8088 -45275 8140
rect -45275 8088 -45273 8140
rect -45141 8104 -45139 8156
rect -45139 8104 -45087 8156
rect -45087 8104 -45085 8156
rect -45141 8102 -45085 8104
rect -45329 8086 -45273 8088
rect -44878 8005 -44822 8007
rect -45112 7971 -45056 7973
rect -45313 7963 -45257 7965
rect -45313 7911 -45311 7963
rect -45311 7911 -45259 7963
rect -45259 7911 -45257 7963
rect -45112 7919 -45110 7971
rect -45110 7919 -45058 7971
rect -45058 7919 -45056 7971
rect -44878 7953 -44876 8005
rect -44876 7953 -44824 8005
rect -44824 7953 -44822 8005
rect -44878 7951 -44822 7953
rect -45112 7917 -45056 7919
rect -44691 7943 -44635 7945
rect -45313 7909 -45257 7911
rect -44691 7891 -44689 7943
rect -44689 7891 -44637 7943
rect -44637 7891 -44635 7943
rect -44691 7889 -44635 7891
rect -45095 7795 -45039 7797
rect -45309 7782 -45253 7784
rect -45309 7730 -45307 7782
rect -45307 7730 -45255 7782
rect -45255 7730 -45253 7782
rect -45095 7743 -45093 7795
rect -45093 7743 -45041 7795
rect -45041 7743 -45039 7795
rect -45095 7741 -45039 7743
rect -44878 7786 -44822 7788
rect -44878 7734 -44876 7786
rect -44876 7734 -44824 7786
rect -44824 7734 -44822 7786
rect -44878 7732 -44822 7734
rect -44648 7758 -44592 7760
rect -45309 7728 -45253 7730
rect -44648 7706 -44646 7758
rect -44646 7706 -44594 7758
rect -44594 7706 -44592 7758
rect -44648 7704 -44592 7706
rect -45170 7224 -45114 7226
rect -45358 7208 -45302 7210
rect -45358 7156 -45356 7208
rect -45356 7156 -45304 7208
rect -45304 7156 -45302 7208
rect -45170 7172 -45168 7224
rect -45168 7172 -45116 7224
rect -45116 7172 -45114 7224
rect -45170 7170 -45114 7172
rect -45358 7154 -45302 7156
rect -44907 7073 -44851 7075
rect -45141 7039 -45085 7041
rect -45342 7031 -45286 7033
rect -45342 6979 -45340 7031
rect -45340 6979 -45288 7031
rect -45288 6979 -45286 7031
rect -45141 6987 -45139 7039
rect -45139 6987 -45087 7039
rect -45087 6987 -45085 7039
rect -44907 7021 -44905 7073
rect -44905 7021 -44853 7073
rect -44853 7021 -44851 7073
rect -44907 7019 -44851 7021
rect -45141 6985 -45085 6987
rect -44720 7011 -44664 7013
rect -45342 6977 -45286 6979
rect -44720 6959 -44718 7011
rect -44718 6959 -44666 7011
rect -44666 6959 -44664 7011
rect -44720 6957 -44664 6959
rect -45124 6863 -45068 6865
rect -45338 6850 -45282 6852
rect -45338 6798 -45336 6850
rect -45336 6798 -45284 6850
rect -45284 6798 -45282 6850
rect -45124 6811 -45122 6863
rect -45122 6811 -45070 6863
rect -45070 6811 -45068 6863
rect -45124 6809 -45068 6811
rect -44907 6854 -44851 6856
rect -44907 6802 -44905 6854
rect -44905 6802 -44853 6854
rect -44853 6802 -44851 6854
rect -44907 6800 -44851 6802
rect -44677 6826 -44621 6828
rect -45338 6796 -45282 6798
rect -44677 6774 -44675 6826
rect -44675 6774 -44623 6826
rect -44623 6774 -44621 6826
rect -44677 6772 -44621 6774
rect -38440 8086 -38384 8088
rect -38628 8070 -38572 8072
rect -38628 8018 -38626 8070
rect -38626 8018 -38574 8070
rect -38574 8018 -38572 8070
rect -38440 8034 -38438 8086
rect -38438 8034 -38386 8086
rect -38386 8034 -38384 8086
rect -38440 8032 -38384 8034
rect -38628 8016 -38572 8018
rect -38177 7935 -38121 7937
rect -38411 7901 -38355 7903
rect -38612 7893 -38556 7895
rect -38612 7841 -38610 7893
rect -38610 7841 -38558 7893
rect -38558 7841 -38556 7893
rect -38411 7849 -38409 7901
rect -38409 7849 -38357 7901
rect -38357 7849 -38355 7901
rect -38177 7883 -38175 7935
rect -38175 7883 -38123 7935
rect -38123 7883 -38121 7935
rect -38177 7881 -38121 7883
rect -38411 7847 -38355 7849
rect -37990 7873 -37934 7875
rect -38612 7839 -38556 7841
rect -37990 7821 -37988 7873
rect -37988 7821 -37936 7873
rect -37936 7821 -37934 7873
rect -37990 7819 -37934 7821
rect -38394 7725 -38338 7727
rect -38608 7712 -38552 7714
rect -38608 7660 -38606 7712
rect -38606 7660 -38554 7712
rect -38554 7660 -38552 7712
rect -38394 7673 -38392 7725
rect -38392 7673 -38340 7725
rect -38340 7673 -38338 7725
rect -38394 7671 -38338 7673
rect -38177 7716 -38121 7718
rect -38177 7664 -38175 7716
rect -38175 7664 -38123 7716
rect -38123 7664 -38121 7716
rect -38177 7662 -38121 7664
rect -37947 7688 -37891 7690
rect -38608 7658 -38552 7660
rect -37947 7636 -37945 7688
rect -37945 7636 -37893 7688
rect -37893 7636 -37891 7688
rect -37947 7634 -37891 7636
rect -38429 7247 -38373 7249
rect -38617 7231 -38561 7233
rect -38617 7179 -38615 7231
rect -38615 7179 -38563 7231
rect -38563 7179 -38561 7231
rect -38429 7195 -38427 7247
rect -38427 7195 -38375 7247
rect -38375 7195 -38373 7247
rect -38429 7193 -38373 7195
rect -38617 7177 -38561 7179
rect -38166 7096 -38110 7098
rect -38400 7062 -38344 7064
rect -38601 7054 -38545 7056
rect -38601 7002 -38599 7054
rect -38599 7002 -38547 7054
rect -38547 7002 -38545 7054
rect -38400 7010 -38398 7062
rect -38398 7010 -38346 7062
rect -38346 7010 -38344 7062
rect -38166 7044 -38164 7096
rect -38164 7044 -38112 7096
rect -38112 7044 -38110 7096
rect -38166 7042 -38110 7044
rect -38400 7008 -38344 7010
rect -37979 7034 -37923 7036
rect -38601 7000 -38545 7002
rect -37979 6982 -37977 7034
rect -37977 6982 -37925 7034
rect -37925 6982 -37923 7034
rect -37979 6980 -37923 6982
rect -38383 6886 -38327 6888
rect -38597 6873 -38541 6875
rect -38597 6821 -38595 6873
rect -38595 6821 -38543 6873
rect -38543 6821 -38541 6873
rect -38383 6834 -38381 6886
rect -38381 6834 -38329 6886
rect -38329 6834 -38327 6886
rect -38383 6832 -38327 6834
rect -38166 6877 -38110 6879
rect -38166 6825 -38164 6877
rect -38164 6825 -38112 6877
rect -38112 6825 -38110 6877
rect -38166 6823 -38110 6825
rect -37936 6849 -37880 6851
rect -38597 6819 -38541 6821
rect -37936 6797 -37934 6849
rect -37934 6797 -37882 6849
rect -37882 6797 -37880 6849
rect -37936 6795 -37880 6797
rect -31413 8145 -31357 8147
rect -31601 8129 -31545 8131
rect -31601 8077 -31599 8129
rect -31599 8077 -31547 8129
rect -31547 8077 -31545 8129
rect -31413 8093 -31411 8145
rect -31411 8093 -31359 8145
rect -31359 8093 -31357 8145
rect -31413 8091 -31357 8093
rect -31601 8075 -31545 8077
rect -31150 7994 -31094 7996
rect -31384 7960 -31328 7962
rect -31585 7952 -31529 7954
rect -31585 7900 -31583 7952
rect -31583 7900 -31531 7952
rect -31531 7900 -31529 7952
rect -31384 7908 -31382 7960
rect -31382 7908 -31330 7960
rect -31330 7908 -31328 7960
rect -31150 7942 -31148 7994
rect -31148 7942 -31096 7994
rect -31096 7942 -31094 7994
rect -31150 7940 -31094 7942
rect -31384 7906 -31328 7908
rect -30963 7932 -30907 7934
rect -31585 7898 -31529 7900
rect -30963 7880 -30961 7932
rect -30961 7880 -30909 7932
rect -30909 7880 -30907 7932
rect -30963 7878 -30907 7880
rect -31367 7784 -31311 7786
rect -31581 7771 -31525 7773
rect -31581 7719 -31579 7771
rect -31579 7719 -31527 7771
rect -31527 7719 -31525 7771
rect -31367 7732 -31365 7784
rect -31365 7732 -31313 7784
rect -31313 7732 -31311 7784
rect -31367 7730 -31311 7732
rect -31150 7775 -31094 7777
rect -31150 7723 -31148 7775
rect -31148 7723 -31096 7775
rect -31096 7723 -31094 7775
rect -31150 7721 -31094 7723
rect -30920 7747 -30864 7749
rect -31581 7717 -31525 7719
rect -30920 7695 -30918 7747
rect -30918 7695 -30866 7747
rect -30866 7695 -30864 7747
rect -30920 7693 -30864 7695
rect -31396 7253 -31340 7255
rect -31584 7237 -31528 7239
rect -31584 7185 -31582 7237
rect -31582 7185 -31530 7237
rect -31530 7185 -31528 7237
rect -31396 7201 -31394 7253
rect -31394 7201 -31342 7253
rect -31342 7201 -31340 7253
rect -31396 7199 -31340 7201
rect -31584 7183 -31528 7185
rect -31133 7102 -31077 7104
rect -31367 7068 -31311 7070
rect -31568 7060 -31512 7062
rect -31568 7008 -31566 7060
rect -31566 7008 -31514 7060
rect -31514 7008 -31512 7060
rect -31367 7016 -31365 7068
rect -31365 7016 -31313 7068
rect -31313 7016 -31311 7068
rect -31133 7050 -31131 7102
rect -31131 7050 -31079 7102
rect -31079 7050 -31077 7102
rect -31133 7048 -31077 7050
rect -31367 7014 -31311 7016
rect -30946 7040 -30890 7042
rect -31568 7006 -31512 7008
rect -30946 6988 -30944 7040
rect -30944 6988 -30892 7040
rect -30892 6988 -30890 7040
rect -30946 6986 -30890 6988
rect -31350 6892 -31294 6894
rect -31564 6879 -31508 6881
rect -31564 6827 -31562 6879
rect -31562 6827 -31510 6879
rect -31510 6827 -31508 6879
rect -31350 6840 -31348 6892
rect -31348 6840 -31296 6892
rect -31296 6840 -31294 6892
rect -31350 6838 -31294 6840
rect -31133 6883 -31077 6885
rect -31133 6831 -31131 6883
rect -31131 6831 -31079 6883
rect -31079 6831 -31077 6883
rect -31133 6829 -31077 6831
rect -30903 6855 -30847 6857
rect -31564 6825 -31508 6827
rect -30903 6803 -30901 6855
rect -30901 6803 -30849 6855
rect -30849 6803 -30847 6855
rect -30903 6801 -30847 6803
rect -24562 8022 -24506 8024
rect -24750 8006 -24694 8008
rect -24750 7954 -24748 8006
rect -24748 7954 -24696 8006
rect -24696 7954 -24694 8006
rect -24562 7970 -24560 8022
rect -24560 7970 -24508 8022
rect -24508 7970 -24506 8022
rect -24562 7968 -24506 7970
rect -24750 7952 -24694 7954
rect -24299 7871 -24243 7873
rect -24533 7837 -24477 7839
rect -24734 7829 -24678 7831
rect -24734 7777 -24732 7829
rect -24732 7777 -24680 7829
rect -24680 7777 -24678 7829
rect -24533 7785 -24531 7837
rect -24531 7785 -24479 7837
rect -24479 7785 -24477 7837
rect -24299 7819 -24297 7871
rect -24297 7819 -24245 7871
rect -24245 7819 -24243 7871
rect -24299 7817 -24243 7819
rect -24533 7783 -24477 7785
rect -24112 7809 -24056 7811
rect -24734 7775 -24678 7777
rect -24112 7757 -24110 7809
rect -24110 7757 -24058 7809
rect -24058 7757 -24056 7809
rect -24112 7755 -24056 7757
rect -24516 7661 -24460 7663
rect -24730 7648 -24674 7650
rect -24730 7596 -24728 7648
rect -24728 7596 -24676 7648
rect -24676 7596 -24674 7648
rect -24516 7609 -24514 7661
rect -24514 7609 -24462 7661
rect -24462 7609 -24460 7661
rect -24516 7607 -24460 7609
rect -24299 7652 -24243 7654
rect -24299 7600 -24297 7652
rect -24297 7600 -24245 7652
rect -24245 7600 -24243 7652
rect -24299 7598 -24243 7600
rect -24069 7624 -24013 7626
rect -24730 7594 -24674 7596
rect -24069 7572 -24067 7624
rect -24067 7572 -24015 7624
rect -24015 7572 -24013 7624
rect -24069 7570 -24013 7572
rect -24573 7189 -24517 7191
rect -24761 7173 -24705 7175
rect -24761 7121 -24759 7173
rect -24759 7121 -24707 7173
rect -24707 7121 -24705 7173
rect -24573 7137 -24571 7189
rect -24571 7137 -24519 7189
rect -24519 7137 -24517 7189
rect -24573 7135 -24517 7137
rect -24761 7119 -24705 7121
rect -24310 7038 -24254 7040
rect -24544 7004 -24488 7006
rect -24745 6996 -24689 6998
rect -24745 6944 -24743 6996
rect -24743 6944 -24691 6996
rect -24691 6944 -24689 6996
rect -24544 6952 -24542 7004
rect -24542 6952 -24490 7004
rect -24490 6952 -24488 7004
rect -24310 6986 -24308 7038
rect -24308 6986 -24256 7038
rect -24256 6986 -24254 7038
rect -24310 6984 -24254 6986
rect -24544 6950 -24488 6952
rect -24123 6976 -24067 6978
rect -24745 6942 -24689 6944
rect -24123 6924 -24121 6976
rect -24121 6924 -24069 6976
rect -24069 6924 -24067 6976
rect -24123 6922 -24067 6924
rect -24527 6828 -24471 6830
rect -24741 6815 -24685 6817
rect -24741 6763 -24739 6815
rect -24739 6763 -24687 6815
rect -24687 6763 -24685 6815
rect -24527 6776 -24525 6828
rect -24525 6776 -24473 6828
rect -24473 6776 -24471 6828
rect -24527 6774 -24471 6776
rect -24310 6819 -24254 6821
rect -24310 6767 -24308 6819
rect -24308 6767 -24256 6819
rect -24256 6767 -24254 6819
rect -24310 6765 -24254 6767
rect -24080 6791 -24024 6793
rect -24741 6761 -24685 6763
rect -24080 6739 -24078 6791
rect -24078 6739 -24026 6791
rect -24026 6739 -24024 6791
rect -24080 6737 -24024 6739
rect -17727 8104 -17671 8106
rect -17915 8088 -17859 8090
rect -17915 8036 -17913 8088
rect -17913 8036 -17861 8088
rect -17861 8036 -17859 8088
rect -17727 8052 -17725 8104
rect -17725 8052 -17673 8104
rect -17673 8052 -17671 8104
rect -17727 8050 -17671 8052
rect -17915 8034 -17859 8036
rect -17464 7953 -17408 7955
rect -17698 7919 -17642 7921
rect -17899 7911 -17843 7913
rect -17899 7859 -17897 7911
rect -17897 7859 -17845 7911
rect -17845 7859 -17843 7911
rect -17698 7867 -17696 7919
rect -17696 7867 -17644 7919
rect -17644 7867 -17642 7919
rect -17464 7901 -17462 7953
rect -17462 7901 -17410 7953
rect -17410 7901 -17408 7953
rect -17464 7899 -17408 7901
rect -17698 7865 -17642 7867
rect -17277 7891 -17221 7893
rect -17899 7857 -17843 7859
rect -17277 7839 -17275 7891
rect -17275 7839 -17223 7891
rect -17223 7839 -17221 7891
rect -17277 7837 -17221 7839
rect -17681 7743 -17625 7745
rect -17895 7730 -17839 7732
rect -17895 7678 -17893 7730
rect -17893 7678 -17841 7730
rect -17841 7678 -17839 7730
rect -17681 7691 -17679 7743
rect -17679 7691 -17627 7743
rect -17627 7691 -17625 7743
rect -17681 7689 -17625 7691
rect -17464 7734 -17408 7736
rect -17464 7682 -17462 7734
rect -17462 7682 -17410 7734
rect -17410 7682 -17408 7734
rect -17464 7680 -17408 7682
rect -17234 7706 -17178 7708
rect -17895 7676 -17839 7678
rect -17234 7654 -17232 7706
rect -17232 7654 -17180 7706
rect -17180 7654 -17178 7706
rect -17234 7652 -17178 7654
rect -17727 7247 -17671 7249
rect -17915 7231 -17859 7233
rect -17915 7179 -17913 7231
rect -17913 7179 -17861 7231
rect -17861 7179 -17859 7231
rect -17727 7195 -17725 7247
rect -17725 7195 -17673 7247
rect -17673 7195 -17671 7247
rect -17727 7193 -17671 7195
rect -17915 7177 -17859 7179
rect -17464 7096 -17408 7098
rect -17698 7062 -17642 7064
rect -17899 7054 -17843 7056
rect -17899 7002 -17897 7054
rect -17897 7002 -17845 7054
rect -17845 7002 -17843 7054
rect -17698 7010 -17696 7062
rect -17696 7010 -17644 7062
rect -17644 7010 -17642 7062
rect -17464 7044 -17462 7096
rect -17462 7044 -17410 7096
rect -17410 7044 -17408 7096
rect -17464 7042 -17408 7044
rect -17698 7008 -17642 7010
rect -17277 7034 -17221 7036
rect -17899 7000 -17843 7002
rect -17277 6982 -17275 7034
rect -17275 6982 -17223 7034
rect -17223 6982 -17221 7034
rect -17277 6980 -17221 6982
rect -17681 6886 -17625 6888
rect -17895 6873 -17839 6875
rect -17895 6821 -17893 6873
rect -17893 6821 -17841 6873
rect -17841 6821 -17839 6873
rect -17681 6834 -17679 6886
rect -17679 6834 -17627 6886
rect -17627 6834 -17625 6886
rect -17681 6832 -17625 6834
rect -17464 6877 -17408 6879
rect -17464 6825 -17462 6877
rect -17462 6825 -17410 6877
rect -17410 6825 -17408 6877
rect -17464 6823 -17408 6825
rect -17234 6849 -17178 6851
rect -17895 6819 -17839 6821
rect -17234 6797 -17232 6849
rect -17232 6797 -17180 6849
rect -17180 6797 -17178 6849
rect -17234 6795 -17178 6797
rect -10735 8191 -10679 8193
rect -10923 8175 -10867 8177
rect -10923 8123 -10921 8175
rect -10921 8123 -10869 8175
rect -10869 8123 -10867 8175
rect -10735 8139 -10733 8191
rect -10733 8139 -10681 8191
rect -10681 8139 -10679 8191
rect -10735 8137 -10679 8139
rect -10923 8121 -10867 8123
rect -10472 8040 -10416 8042
rect -10706 8006 -10650 8008
rect -10907 7998 -10851 8000
rect -10907 7946 -10905 7998
rect -10905 7946 -10853 7998
rect -10853 7946 -10851 7998
rect -10706 7954 -10704 8006
rect -10704 7954 -10652 8006
rect -10652 7954 -10650 8006
rect -10472 7988 -10470 8040
rect -10470 7988 -10418 8040
rect -10418 7988 -10416 8040
rect -10472 7986 -10416 7988
rect -10706 7952 -10650 7954
rect -10285 7978 -10229 7980
rect -10907 7944 -10851 7946
rect -10285 7926 -10283 7978
rect -10283 7926 -10231 7978
rect -10231 7926 -10229 7978
rect -10285 7924 -10229 7926
rect -10689 7830 -10633 7832
rect -10903 7817 -10847 7819
rect -10903 7765 -10901 7817
rect -10901 7765 -10849 7817
rect -10849 7765 -10847 7817
rect -10689 7778 -10687 7830
rect -10687 7778 -10635 7830
rect -10635 7778 -10633 7830
rect -10689 7776 -10633 7778
rect -10472 7821 -10416 7823
rect -10472 7769 -10470 7821
rect -10470 7769 -10418 7821
rect -10418 7769 -10416 7821
rect -10472 7767 -10416 7769
rect -10242 7793 -10186 7795
rect -10903 7763 -10847 7765
rect -10242 7741 -10240 7793
rect -10240 7741 -10188 7793
rect -10188 7741 -10186 7793
rect -10242 7739 -10186 7741
rect -10712 7206 -10656 7208
rect -10900 7190 -10844 7192
rect -10900 7138 -10898 7190
rect -10898 7138 -10846 7190
rect -10846 7138 -10844 7190
rect -10712 7154 -10710 7206
rect -10710 7154 -10658 7206
rect -10658 7154 -10656 7206
rect -10712 7152 -10656 7154
rect -10900 7136 -10844 7138
rect -10449 7055 -10393 7057
rect -10683 7021 -10627 7023
rect -10884 7013 -10828 7015
rect -10884 6961 -10882 7013
rect -10882 6961 -10830 7013
rect -10830 6961 -10828 7013
rect -10683 6969 -10681 7021
rect -10681 6969 -10629 7021
rect -10629 6969 -10627 7021
rect -10449 7003 -10447 7055
rect -10447 7003 -10395 7055
rect -10395 7003 -10393 7055
rect -10449 7001 -10393 7003
rect -10683 6967 -10627 6969
rect -10262 6993 -10206 6995
rect -10884 6959 -10828 6961
rect -10262 6941 -10260 6993
rect -10260 6941 -10208 6993
rect -10208 6941 -10206 6993
rect -10262 6939 -10206 6941
rect -10666 6845 -10610 6847
rect -10880 6832 -10824 6834
rect -10880 6780 -10878 6832
rect -10878 6780 -10826 6832
rect -10826 6780 -10824 6832
rect -10666 6793 -10664 6845
rect -10664 6793 -10612 6845
rect -10612 6793 -10610 6845
rect -10666 6791 -10610 6793
rect -10449 6836 -10393 6838
rect -10449 6784 -10447 6836
rect -10447 6784 -10395 6836
rect -10395 6784 -10393 6836
rect -10449 6782 -10393 6784
rect -10219 6808 -10163 6810
rect -10880 6778 -10824 6780
rect -10219 6756 -10217 6808
rect -10217 6756 -10165 6808
rect -10165 6756 -10163 6808
rect -10219 6754 -10163 6756
rect -3295 8209 -3239 8211
rect -3483 8193 -3427 8195
rect -3483 8141 -3481 8193
rect -3481 8141 -3429 8193
rect -3429 8141 -3427 8193
rect -3295 8157 -3293 8209
rect -3293 8157 -3241 8209
rect -3241 8157 -3239 8209
rect -3295 8155 -3239 8157
rect -3483 8139 -3427 8141
rect -3032 8058 -2976 8060
rect -3266 8024 -3210 8026
rect -3467 8016 -3411 8018
rect -3467 7964 -3465 8016
rect -3465 7964 -3413 8016
rect -3413 7964 -3411 8016
rect -3266 7972 -3264 8024
rect -3264 7972 -3212 8024
rect -3212 7972 -3210 8024
rect -3032 8006 -3030 8058
rect -3030 8006 -2978 8058
rect -2978 8006 -2976 8058
rect -3032 8004 -2976 8006
rect -3266 7970 -3210 7972
rect -2845 7996 -2789 7998
rect -3467 7962 -3411 7964
rect -2845 7944 -2843 7996
rect -2843 7944 -2791 7996
rect -2791 7944 -2789 7996
rect -2845 7942 -2789 7944
rect -3249 7848 -3193 7850
rect -3463 7835 -3407 7837
rect -3463 7783 -3461 7835
rect -3461 7783 -3409 7835
rect -3409 7783 -3407 7835
rect -3249 7796 -3247 7848
rect -3247 7796 -3195 7848
rect -3195 7796 -3193 7848
rect -3249 7794 -3193 7796
rect -3032 7839 -2976 7841
rect -3032 7787 -3030 7839
rect -3030 7787 -2978 7839
rect -2978 7787 -2976 7839
rect -3032 7785 -2976 7787
rect -2802 7811 -2746 7813
rect -3463 7781 -3407 7783
rect -2802 7759 -2800 7811
rect -2800 7759 -2748 7811
rect -2748 7759 -2746 7811
rect -2802 7757 -2746 7759
rect -3225 7236 -3169 7238
rect -3413 7220 -3357 7222
rect -3413 7168 -3411 7220
rect -3411 7168 -3359 7220
rect -3359 7168 -3357 7220
rect -3225 7184 -3223 7236
rect -3223 7184 -3171 7236
rect -3171 7184 -3169 7236
rect -3225 7182 -3169 7184
rect -3413 7166 -3357 7168
rect -2962 7085 -2906 7087
rect -3196 7051 -3140 7053
rect -3397 7043 -3341 7045
rect -3397 6991 -3395 7043
rect -3395 6991 -3343 7043
rect -3343 6991 -3341 7043
rect -3196 6999 -3194 7051
rect -3194 6999 -3142 7051
rect -3142 6999 -3140 7051
rect -2962 7033 -2960 7085
rect -2960 7033 -2908 7085
rect -2908 7033 -2906 7085
rect -2962 7031 -2906 7033
rect -3196 6997 -3140 6999
rect -2775 7023 -2719 7025
rect -3397 6989 -3341 6991
rect -2775 6971 -2773 7023
rect -2773 6971 -2721 7023
rect -2721 6971 -2719 7023
rect -2775 6969 -2719 6971
rect -3179 6875 -3123 6877
rect -3393 6862 -3337 6864
rect -3393 6810 -3391 6862
rect -3391 6810 -3339 6862
rect -3339 6810 -3337 6862
rect -3179 6823 -3177 6875
rect -3177 6823 -3125 6875
rect -3125 6823 -3123 6875
rect -3179 6821 -3123 6823
rect -2962 6866 -2906 6868
rect -2962 6814 -2960 6866
rect -2960 6814 -2908 6866
rect -2908 6814 -2906 6866
rect -2962 6812 -2906 6814
rect -2732 6838 -2676 6840
rect -3393 6808 -3337 6810
rect -2732 6786 -2730 6838
rect -2730 6786 -2678 6838
rect -2678 6786 -2676 6838
rect -2732 6784 -2676 6786
rect 2415 8162 2471 8164
rect 2227 8146 2283 8148
rect 2227 8094 2229 8146
rect 2229 8094 2281 8146
rect 2281 8094 2283 8146
rect 2415 8110 2417 8162
rect 2417 8110 2469 8162
rect 2469 8110 2471 8162
rect 2415 8108 2471 8110
rect 2227 8092 2283 8094
rect 2678 8011 2734 8013
rect 2444 7977 2500 7979
rect 2243 7969 2299 7971
rect 2243 7917 2245 7969
rect 2245 7917 2297 7969
rect 2297 7917 2299 7969
rect 2444 7925 2446 7977
rect 2446 7925 2498 7977
rect 2498 7925 2500 7977
rect 2678 7959 2680 8011
rect 2680 7959 2732 8011
rect 2732 7959 2734 8011
rect 2678 7957 2734 7959
rect 2444 7923 2500 7925
rect 2865 7949 2921 7951
rect 2243 7915 2299 7917
rect 2865 7897 2867 7949
rect 2867 7897 2919 7949
rect 2919 7897 2921 7949
rect 2865 7895 2921 7897
rect 2461 7801 2517 7803
rect 2247 7788 2303 7790
rect 2247 7736 2249 7788
rect 2249 7736 2301 7788
rect 2301 7736 2303 7788
rect 2461 7749 2463 7801
rect 2463 7749 2515 7801
rect 2515 7749 2517 7801
rect 2461 7747 2517 7749
rect 2678 7792 2734 7794
rect 2678 7740 2680 7792
rect 2680 7740 2732 7792
rect 2732 7740 2734 7792
rect 2678 7738 2734 7740
rect 2908 7764 2964 7766
rect 2247 7734 2303 7736
rect 2908 7712 2910 7764
rect 2910 7712 2962 7764
rect 2962 7712 2964 7764
rect 2908 7710 2964 7712
rect 2444 7137 2500 7139
rect 2256 7121 2312 7123
rect 2256 7069 2258 7121
rect 2258 7069 2310 7121
rect 2310 7069 2312 7121
rect 2444 7085 2446 7137
rect 2446 7085 2498 7137
rect 2498 7085 2500 7137
rect 2444 7083 2500 7085
rect 2256 7067 2312 7069
rect 2707 6986 2763 6988
rect 2473 6952 2529 6954
rect 2272 6944 2328 6946
rect 2272 6892 2274 6944
rect 2274 6892 2326 6944
rect 2326 6892 2328 6944
rect 2473 6900 2475 6952
rect 2475 6900 2527 6952
rect 2527 6900 2529 6952
rect 2707 6934 2709 6986
rect 2709 6934 2761 6986
rect 2761 6934 2763 6986
rect 2707 6932 2763 6934
rect 2473 6898 2529 6900
rect 2894 6924 2950 6926
rect 2272 6890 2328 6892
rect 2894 6872 2896 6924
rect 2896 6872 2948 6924
rect 2948 6872 2950 6924
rect 2894 6870 2950 6872
rect 2490 6776 2546 6778
rect 2276 6763 2332 6765
rect 2276 6711 2278 6763
rect 2278 6711 2330 6763
rect 2330 6711 2332 6763
rect 2490 6724 2492 6776
rect 2492 6724 2544 6776
rect 2544 6724 2546 6776
rect 2490 6722 2546 6724
rect 2707 6767 2763 6769
rect 2707 6715 2709 6767
rect 2709 6715 2761 6767
rect 2761 6715 2763 6767
rect 2707 6713 2763 6715
rect 2937 6739 2993 6741
rect 2276 6709 2332 6711
rect 2937 6687 2939 6739
rect 2939 6687 2991 6739
rect 2991 6687 2993 6739
rect 2937 6685 2993 6687
rect -61490 -68322 -61434 -68320
rect -61678 -68338 -61622 -68336
rect -61678 -68390 -61676 -68338
rect -61676 -68390 -61624 -68338
rect -61624 -68390 -61622 -68338
rect -61490 -68374 -61488 -68322
rect -61488 -68374 -61436 -68322
rect -61436 -68374 -61434 -68322
rect -61490 -68376 -61434 -68374
rect -61678 -68392 -61622 -68390
rect -61227 -68473 -61171 -68471
rect -61461 -68507 -61405 -68505
rect -61662 -68515 -61606 -68513
rect -61662 -68567 -61660 -68515
rect -61660 -68567 -61608 -68515
rect -61608 -68567 -61606 -68515
rect -61461 -68559 -61459 -68507
rect -61459 -68559 -61407 -68507
rect -61407 -68559 -61405 -68507
rect -61227 -68525 -61225 -68473
rect -61225 -68525 -61173 -68473
rect -61173 -68525 -61171 -68473
rect -61227 -68527 -61171 -68525
rect -61461 -68561 -61405 -68559
rect -61040 -68535 -60984 -68533
rect -61662 -68569 -61606 -68567
rect -61040 -68587 -61038 -68535
rect -61038 -68587 -60986 -68535
rect -60986 -68587 -60984 -68535
rect -61040 -68589 -60984 -68587
rect -61444 -68683 -61388 -68681
rect -61658 -68696 -61602 -68694
rect -61658 -68748 -61656 -68696
rect -61656 -68748 -61604 -68696
rect -61604 -68748 -61602 -68696
rect -61444 -68735 -61442 -68683
rect -61442 -68735 -61390 -68683
rect -61390 -68735 -61388 -68683
rect -61444 -68737 -61388 -68735
rect -61227 -68692 -61171 -68690
rect -61227 -68744 -61225 -68692
rect -61225 -68744 -61173 -68692
rect -61173 -68744 -61171 -68692
rect -61227 -68746 -61171 -68744
rect -60997 -68720 -60941 -68718
rect -61658 -68750 -61602 -68748
rect -60997 -68772 -60995 -68720
rect -60995 -68772 -60943 -68720
rect -60943 -68772 -60941 -68720
rect -60997 -68774 -60941 -68772
rect -54944 -68381 -54888 -68379
rect -54944 -68433 -54942 -68381
rect -54942 -68433 -54890 -68381
rect -54890 -68433 -54888 -68381
rect -54944 -68435 -54888 -68433
rect -54769 -68381 -54713 -68379
rect -54769 -68433 -54767 -68381
rect -54767 -68433 -54715 -68381
rect -54715 -68433 -54713 -68381
rect -54769 -68435 -54713 -68433
rect -54567 -68381 -54511 -68379
rect -54567 -68433 -54565 -68381
rect -54565 -68433 -54513 -68381
rect -54513 -68433 -54511 -68381
rect -54567 -68435 -54511 -68433
rect -54725 -68621 -54669 -68619
rect -54925 -68646 -54869 -68644
rect -55157 -68648 -55101 -68646
rect -55157 -68700 -55155 -68648
rect -55155 -68700 -55103 -68648
rect -55103 -68700 -55101 -68648
rect -54925 -68698 -54923 -68646
rect -54923 -68698 -54871 -68646
rect -54871 -68698 -54869 -68646
rect -54725 -68673 -54723 -68621
rect -54723 -68673 -54671 -68621
rect -54671 -68673 -54669 -68621
rect -54294 -68636 -54238 -68634
rect -54725 -68675 -54669 -68673
rect -54507 -68652 -54451 -68650
rect -54925 -68700 -54869 -68698
rect -55157 -68702 -55101 -68700
rect -54507 -68704 -54505 -68652
rect -54505 -68704 -54453 -68652
rect -54453 -68704 -54451 -68652
rect -54294 -68688 -54292 -68636
rect -54292 -68688 -54240 -68636
rect -54240 -68688 -54238 -68636
rect -54294 -68690 -54238 -68688
rect -54507 -68706 -54451 -68704
rect -54696 -68865 -54640 -68863
rect -54921 -68869 -54865 -68867
rect -54921 -68921 -54919 -68869
rect -54919 -68921 -54867 -68869
rect -54867 -68921 -54865 -68869
rect -54696 -68917 -54694 -68865
rect -54694 -68917 -54642 -68865
rect -54642 -68917 -54640 -68865
rect -54696 -68919 -54640 -68917
rect -54438 -68871 -54382 -68869
rect -54921 -68923 -54865 -68921
rect -54438 -68923 -54436 -68871
rect -54436 -68923 -54384 -68871
rect -54384 -68923 -54382 -68871
rect -54438 -68925 -54382 -68923
rect -48168 -68371 -48112 -68369
rect -48168 -68423 -48166 -68371
rect -48166 -68423 -48114 -68371
rect -48114 -68423 -48112 -68371
rect -48168 -68425 -48112 -68423
rect -47987 -68371 -47931 -68369
rect -47987 -68423 -47985 -68371
rect -47985 -68423 -47933 -68371
rect -47933 -68423 -47931 -68371
rect -47987 -68425 -47931 -68423
rect -47783 -68377 -47727 -68375
rect -47783 -68429 -47781 -68377
rect -47781 -68429 -47729 -68377
rect -47729 -68429 -47727 -68377
rect -47783 -68431 -47727 -68429
rect -47916 -68571 -47860 -68569
rect -48152 -68577 -48096 -68575
rect -48152 -68629 -48150 -68577
rect -48150 -68629 -48098 -68577
rect -48098 -68629 -48096 -68577
rect -47916 -68623 -47914 -68571
rect -47914 -68623 -47862 -68571
rect -47862 -68623 -47860 -68571
rect -47916 -68625 -47860 -68623
rect -47656 -68586 -47600 -68584
rect -48152 -68631 -48096 -68629
rect -47656 -68638 -47654 -68586
rect -47654 -68638 -47602 -68586
rect -47602 -68638 -47600 -68586
rect -47656 -68640 -47600 -68638
rect -48212 -68788 -48156 -68786
rect -48212 -68840 -48210 -68788
rect -48210 -68840 -48158 -68788
rect -48158 -68840 -48156 -68788
rect -48212 -68842 -48156 -68840
rect -47970 -68792 -47914 -68790
rect -47970 -68844 -47968 -68792
rect -47968 -68844 -47916 -68792
rect -47916 -68844 -47914 -68792
rect -47970 -68846 -47914 -68844
rect -47770 -68792 -47714 -68790
rect -47770 -68844 -47768 -68792
rect -47768 -68844 -47716 -68792
rect -47716 -68844 -47714 -68792
rect -47770 -68846 -47714 -68844
rect -47466 -68802 -47410 -68800
rect -47466 -68854 -47464 -68802
rect -47464 -68854 -47412 -68802
rect -47412 -68854 -47410 -68802
rect -47466 -68856 -47410 -68854
rect -41151 -68371 -41095 -68369
rect -41332 -68375 -41276 -68373
rect -41332 -68427 -41330 -68375
rect -41330 -68427 -41278 -68375
rect -41278 -68427 -41276 -68375
rect -41151 -68423 -41149 -68371
rect -41149 -68423 -41097 -68371
rect -41097 -68423 -41095 -68371
rect -41151 -68425 -41095 -68423
rect -40951 -68381 -40895 -68379
rect -41332 -68429 -41276 -68427
rect -40951 -68433 -40949 -68381
rect -40949 -68433 -40897 -68381
rect -40897 -68433 -40895 -68381
rect -40951 -68435 -40895 -68433
rect -41330 -68544 -41274 -68542
rect -41517 -68583 -41461 -68581
rect -41517 -68635 -41515 -68583
rect -41515 -68635 -41463 -68583
rect -41463 -68635 -41461 -68583
rect -41330 -68596 -41328 -68544
rect -41328 -68596 -41276 -68544
rect -41276 -68596 -41274 -68544
rect -40890 -68548 -40834 -68546
rect -41330 -68598 -41274 -68596
rect -41117 -68558 -41061 -68556
rect -41117 -68610 -41115 -68558
rect -41115 -68610 -41063 -68558
rect -41063 -68610 -41061 -68558
rect -40890 -68600 -40888 -68548
rect -40888 -68600 -40836 -68548
rect -40836 -68600 -40834 -68548
rect -40890 -68602 -40834 -68600
rect -40694 -68571 -40638 -68569
rect -41117 -68612 -41061 -68610
rect -40694 -68623 -40692 -68571
rect -40692 -68623 -40640 -68571
rect -40640 -68623 -40638 -68571
rect -40694 -68625 -40638 -68623
rect -41517 -68637 -41461 -68635
rect -41084 -68744 -41028 -68742
rect -41317 -68761 -41261 -68759
rect -41317 -68813 -41315 -68761
rect -41315 -68813 -41263 -68761
rect -41263 -68813 -41261 -68761
rect -41084 -68796 -41082 -68744
rect -41082 -68796 -41030 -68744
rect -41030 -68796 -41028 -68744
rect -41084 -68798 -41028 -68796
rect -40836 -68756 -40780 -68754
rect -40836 -68808 -40834 -68756
rect -40834 -68808 -40782 -68756
rect -40782 -68808 -40780 -68756
rect -40836 -68810 -40780 -68808
rect -41317 -68815 -41261 -68813
rect -34577 -68410 -34521 -68408
rect -34577 -68462 -34575 -68410
rect -34575 -68462 -34523 -68410
rect -34523 -68462 -34521 -68410
rect -34577 -68464 -34521 -68462
rect -34396 -68417 -34340 -68415
rect -34396 -68469 -34394 -68417
rect -34394 -68469 -34342 -68417
rect -34342 -68469 -34340 -68417
rect -34396 -68471 -34340 -68469
rect -34221 -68417 -34165 -68415
rect -34221 -68469 -34219 -68417
rect -34219 -68469 -34167 -68417
rect -34167 -68469 -34165 -68417
rect -34221 -68471 -34165 -68469
rect -34000 -68627 -33944 -68625
rect -34560 -68633 -34504 -68631
rect -34819 -68652 -34763 -68650
rect -34819 -68704 -34817 -68652
rect -34817 -68704 -34765 -68652
rect -34765 -68704 -34763 -68652
rect -34560 -68685 -34558 -68633
rect -34558 -68685 -34506 -68633
rect -34506 -68685 -34504 -68633
rect -34560 -68687 -34504 -68685
rect -34329 -68633 -34273 -68631
rect -34329 -68685 -34327 -68633
rect -34327 -68685 -34275 -68633
rect -34275 -68685 -34273 -68633
rect -34000 -68679 -33998 -68627
rect -33998 -68679 -33946 -68627
rect -33946 -68679 -33944 -68627
rect -34000 -68681 -33944 -68679
rect -34329 -68687 -34273 -68685
rect -34819 -68706 -34763 -68704
rect -33843 -68836 -33787 -68834
rect -34581 -68850 -34525 -68848
rect -34581 -68902 -34579 -68850
rect -34579 -68902 -34527 -68850
rect -34527 -68902 -34525 -68850
rect -34581 -68904 -34525 -68902
rect -34346 -68850 -34290 -68848
rect -34346 -68902 -34344 -68850
rect -34344 -68902 -34292 -68850
rect -34292 -68902 -34290 -68850
rect -34346 -68904 -34290 -68902
rect -34106 -68854 -34050 -68852
rect -34106 -68906 -34104 -68854
rect -34104 -68906 -34052 -68854
rect -34052 -68906 -34050 -68854
rect -33843 -68888 -33841 -68836
rect -33841 -68888 -33789 -68836
rect -33789 -68888 -33787 -68836
rect -33843 -68890 -33787 -68888
rect -34106 -68908 -34050 -68906
rect -27727 -68390 -27671 -68388
rect -27727 -68442 -27725 -68390
rect -27725 -68442 -27673 -68390
rect -27673 -68442 -27671 -68390
rect -27727 -68444 -27671 -68442
rect -27546 -68397 -27490 -68395
rect -27546 -68449 -27544 -68397
rect -27544 -68449 -27492 -68397
rect -27492 -68449 -27490 -68397
rect -27546 -68451 -27490 -68449
rect -27371 -68397 -27315 -68395
rect -27371 -68449 -27369 -68397
rect -27369 -68449 -27317 -68397
rect -27317 -68449 -27315 -68397
rect -27371 -68451 -27315 -68449
rect -27150 -68607 -27094 -68605
rect -27710 -68613 -27654 -68611
rect -27969 -68632 -27913 -68630
rect -27969 -68684 -27967 -68632
rect -27967 -68684 -27915 -68632
rect -27915 -68684 -27913 -68632
rect -27710 -68665 -27708 -68613
rect -27708 -68665 -27656 -68613
rect -27656 -68665 -27654 -68613
rect -27710 -68667 -27654 -68665
rect -27479 -68613 -27423 -68611
rect -27479 -68665 -27477 -68613
rect -27477 -68665 -27425 -68613
rect -27425 -68665 -27423 -68613
rect -27150 -68659 -27148 -68607
rect -27148 -68659 -27096 -68607
rect -27096 -68659 -27094 -68607
rect -27150 -68661 -27094 -68659
rect -27479 -68667 -27423 -68665
rect -27969 -68686 -27913 -68684
rect -26993 -68816 -26937 -68814
rect -27731 -68830 -27675 -68828
rect -27731 -68882 -27729 -68830
rect -27729 -68882 -27677 -68830
rect -27677 -68882 -27675 -68830
rect -27731 -68884 -27675 -68882
rect -27496 -68830 -27440 -68828
rect -27496 -68882 -27494 -68830
rect -27494 -68882 -27442 -68830
rect -27442 -68882 -27440 -68830
rect -27496 -68884 -27440 -68882
rect -27256 -68834 -27200 -68832
rect -27256 -68886 -27254 -68834
rect -27254 -68886 -27202 -68834
rect -27202 -68886 -27200 -68834
rect -26993 -68868 -26991 -68816
rect -26991 -68868 -26939 -68816
rect -26939 -68868 -26937 -68816
rect -26993 -68870 -26937 -68868
rect -27256 -68888 -27200 -68886
rect -20787 -68390 -20731 -68388
rect -20787 -68442 -20785 -68390
rect -20785 -68442 -20733 -68390
rect -20733 -68442 -20731 -68390
rect -20787 -68444 -20731 -68442
rect -20606 -68397 -20550 -68395
rect -20606 -68449 -20604 -68397
rect -20604 -68449 -20552 -68397
rect -20552 -68449 -20550 -68397
rect -20606 -68451 -20550 -68449
rect -20431 -68397 -20375 -68395
rect -20431 -68449 -20429 -68397
rect -20429 -68449 -20377 -68397
rect -20377 -68449 -20375 -68397
rect -20431 -68451 -20375 -68449
rect -20210 -68607 -20154 -68605
rect -20770 -68613 -20714 -68611
rect -21029 -68632 -20973 -68630
rect -21029 -68684 -21027 -68632
rect -21027 -68684 -20975 -68632
rect -20975 -68684 -20973 -68632
rect -20770 -68665 -20768 -68613
rect -20768 -68665 -20716 -68613
rect -20716 -68665 -20714 -68613
rect -20770 -68667 -20714 -68665
rect -20539 -68613 -20483 -68611
rect -20539 -68665 -20537 -68613
rect -20537 -68665 -20485 -68613
rect -20485 -68665 -20483 -68613
rect -20210 -68659 -20208 -68607
rect -20208 -68659 -20156 -68607
rect -20156 -68659 -20154 -68607
rect -20210 -68661 -20154 -68659
rect -20539 -68667 -20483 -68665
rect -21029 -68686 -20973 -68684
rect -20053 -68816 -19997 -68814
rect -20791 -68830 -20735 -68828
rect -20791 -68882 -20789 -68830
rect -20789 -68882 -20737 -68830
rect -20737 -68882 -20735 -68830
rect -20791 -68884 -20735 -68882
rect -20556 -68830 -20500 -68828
rect -20556 -68882 -20554 -68830
rect -20554 -68882 -20502 -68830
rect -20502 -68882 -20500 -68830
rect -20556 -68884 -20500 -68882
rect -20316 -68834 -20260 -68832
rect -20316 -68886 -20314 -68834
rect -20314 -68886 -20262 -68834
rect -20262 -68886 -20260 -68834
rect -20053 -68868 -20051 -68816
rect -20051 -68868 -19999 -68816
rect -19999 -68868 -19997 -68816
rect -20053 -68870 -19997 -68868
rect -20316 -68888 -20260 -68886
rect -14124 -68383 -14068 -68381
rect -14124 -68435 -14122 -68383
rect -14122 -68435 -14070 -68383
rect -14070 -68435 -14068 -68383
rect -14124 -68437 -14068 -68435
rect -13945 -68388 -13889 -68386
rect -13945 -68440 -13943 -68388
rect -13943 -68440 -13891 -68388
rect -13891 -68440 -13889 -68388
rect -13945 -68442 -13889 -68440
rect -13762 -68388 -13706 -68386
rect -13762 -68440 -13760 -68388
rect -13760 -68440 -13708 -68388
rect -13708 -68440 -13706 -68388
rect -13762 -68442 -13706 -68440
rect -13637 -68636 -13581 -68634
rect -13845 -68640 -13789 -68638
rect -14037 -68646 -13981 -68644
rect -14262 -68652 -14206 -68650
rect -14262 -68704 -14260 -68652
rect -14260 -68704 -14208 -68652
rect -14208 -68704 -14206 -68652
rect -14037 -68698 -14035 -68646
rect -14035 -68698 -13983 -68646
rect -13983 -68698 -13981 -68646
rect -13845 -68692 -13843 -68640
rect -13843 -68692 -13791 -68640
rect -13791 -68692 -13789 -68640
rect -13637 -68688 -13635 -68636
rect -13635 -68688 -13583 -68636
rect -13583 -68688 -13581 -68636
rect -13637 -68690 -13581 -68688
rect -13845 -68694 -13789 -68692
rect -14037 -68700 -13981 -68698
rect -14262 -68706 -14206 -68704
rect -14199 -68850 -14143 -68848
rect -14199 -68902 -14197 -68850
rect -14197 -68902 -14145 -68850
rect -14145 -68902 -14143 -68850
rect -14199 -68904 -14143 -68902
rect -13980 -68850 -13924 -68848
rect -13980 -68902 -13978 -68850
rect -13978 -68902 -13926 -68850
rect -13926 -68902 -13924 -68850
rect -13980 -68904 -13924 -68902
rect -13791 -68850 -13735 -68848
rect -13791 -68902 -13789 -68850
rect -13789 -68902 -13737 -68850
rect -13737 -68902 -13735 -68850
rect -13791 -68904 -13735 -68902
rect -13543 -68850 -13487 -68848
rect -13543 -68902 -13541 -68850
rect -13541 -68902 -13489 -68850
rect -13489 -68902 -13487 -68850
rect -13543 -68904 -13487 -68902
rect -7286 -68363 -7230 -68361
rect -7286 -68415 -7284 -68363
rect -7284 -68415 -7232 -68363
rect -7232 -68415 -7230 -68363
rect -7286 -68417 -7230 -68415
rect -7111 -68363 -7055 -68361
rect -7111 -68415 -7109 -68363
rect -7109 -68415 -7057 -68363
rect -7057 -68415 -7055 -68363
rect -7111 -68417 -7055 -68415
rect -6921 -68363 -6865 -68361
rect -6921 -68415 -6919 -68363
rect -6919 -68415 -6867 -68363
rect -6867 -68415 -6865 -68363
rect -6921 -68417 -6865 -68415
rect -6648 -68613 -6592 -68611
rect -6909 -68619 -6853 -68617
rect -7129 -68625 -7073 -68623
rect -7402 -68631 -7346 -68629
rect -7402 -68683 -7400 -68631
rect -7400 -68683 -7348 -68631
rect -7348 -68683 -7346 -68631
rect -7129 -68677 -7127 -68625
rect -7127 -68677 -7075 -68625
rect -7075 -68677 -7073 -68625
rect -6909 -68671 -6907 -68619
rect -6907 -68671 -6855 -68619
rect -6855 -68671 -6853 -68619
rect -6648 -68665 -6646 -68613
rect -6646 -68665 -6594 -68613
rect -6594 -68665 -6592 -68613
rect -6648 -68667 -6592 -68665
rect -6909 -68673 -6853 -68671
rect -7129 -68679 -7073 -68677
rect -7402 -68685 -7346 -68683
rect -6723 -68848 -6667 -68846
rect -7152 -68854 -7096 -68852
rect -7367 -68856 -7311 -68854
rect -7367 -68908 -7365 -68856
rect -7365 -68908 -7313 -68856
rect -7313 -68908 -7311 -68856
rect -7152 -68906 -7150 -68854
rect -7150 -68906 -7098 -68854
rect -7098 -68906 -7096 -68854
rect -7152 -68908 -7096 -68906
rect -6934 -68854 -6878 -68852
rect -6934 -68906 -6932 -68854
rect -6932 -68906 -6880 -68854
rect -6880 -68906 -6878 -68854
rect -6723 -68900 -6721 -68848
rect -6721 -68900 -6669 -68848
rect -6669 -68900 -6667 -68848
rect -6723 -68902 -6667 -68900
rect -6934 -68908 -6878 -68906
rect -7367 -68910 -7311 -68908
rect -70 -68360 -14 -68358
rect -476 -68363 -420 -68361
rect -476 -68415 -474 -68363
rect -474 -68415 -422 -68363
rect -422 -68415 -420 -68363
rect -476 -68417 -420 -68415
rect -283 -68367 -227 -68365
rect -283 -68419 -281 -68367
rect -281 -68419 -229 -68367
rect -229 -68419 -227 -68367
rect -70 -68412 -68 -68360
rect -68 -68412 -16 -68360
rect -16 -68412 -14 -68360
rect -70 -68414 -14 -68412
rect -283 -68421 -227 -68419
rect 145 -68596 201 -68594
rect -345 -68600 -289 -68598
rect -595 -68604 -539 -68602
rect -595 -68656 -593 -68604
rect -593 -68656 -541 -68604
rect -541 -68656 -539 -68604
rect -345 -68652 -343 -68600
rect -343 -68652 -291 -68600
rect -291 -68652 -289 -68600
rect -345 -68654 -289 -68652
rect -112 -68600 -56 -68598
rect -112 -68652 -110 -68600
rect -110 -68652 -58 -68600
rect -58 -68652 -56 -68600
rect 145 -68648 147 -68596
rect 147 -68648 199 -68596
rect 199 -68648 201 -68596
rect 145 -68650 201 -68648
rect -112 -68654 -56 -68652
rect -595 -68658 -539 -68656
rect -308 -68850 -252 -68848
rect -566 -68854 -510 -68852
rect -566 -68906 -564 -68854
rect -564 -68906 -512 -68854
rect -512 -68906 -510 -68854
rect -308 -68902 -306 -68850
rect -306 -68902 -254 -68850
rect -254 -68902 -252 -68850
rect -308 -68904 -252 -68902
rect -70 -68854 -14 -68852
rect -566 -68908 -510 -68906
rect -70 -68906 -68 -68854
rect -68 -68906 -16 -68854
rect -16 -68906 -14 -68854
rect -70 -68908 -14 -68906
rect 184 -68861 240 -68859
rect 184 -68913 186 -68861
rect 186 -68913 238 -68861
rect 238 -68913 240 -68861
rect 184 -68915 240 -68913
rect 6318 -68354 6374 -68352
rect 6318 -68406 6320 -68354
rect 6320 -68406 6372 -68354
rect 6372 -68406 6374 -68354
rect 6318 -68408 6374 -68406
rect 6506 -68354 6562 -68352
rect 6506 -68406 6508 -68354
rect 6508 -68406 6560 -68354
rect 6560 -68406 6562 -68354
rect 6506 -68408 6562 -68406
rect 6708 -68360 6764 -68358
rect 6708 -68412 6710 -68360
rect 6710 -68412 6762 -68360
rect 6762 -68412 6764 -68360
rect 6708 -68414 6764 -68412
rect 6143 -68575 6199 -68573
rect 6143 -68627 6145 -68575
rect 6145 -68627 6197 -68575
rect 6197 -68627 6199 -68575
rect 6606 -68575 6662 -68573
rect 6143 -68629 6199 -68627
rect 6395 -68579 6451 -68577
rect 6395 -68631 6397 -68579
rect 6397 -68631 6449 -68579
rect 6449 -68631 6451 -68579
rect 6606 -68627 6608 -68575
rect 6608 -68627 6660 -68575
rect 6660 -68627 6662 -68575
rect 6606 -68629 6662 -68627
rect 6395 -68633 6451 -68631
rect 5931 -68690 5987 -68688
rect 5931 -68742 5933 -68690
rect 5933 -68742 5985 -68690
rect 5985 -68742 5987 -68690
rect 5931 -68744 5987 -68742
rect 6327 -68854 6383 -68852
rect 6139 -68856 6195 -68854
rect 6139 -68908 6141 -68856
rect 6141 -68908 6193 -68856
rect 6193 -68908 6195 -68856
rect 6327 -68906 6329 -68854
rect 6329 -68906 6381 -68854
rect 6381 -68906 6383 -68854
rect 6327 -68908 6383 -68906
rect 6533 -68854 6589 -68852
rect 6533 -68906 6535 -68854
rect 6535 -68906 6587 -68854
rect 6587 -68906 6589 -68854
rect 6533 -68908 6589 -68906
rect 6737 -68856 6793 -68854
rect 6737 -68908 6739 -68856
rect 6739 -68908 6791 -68856
rect 6791 -68908 6793 -68856
rect 6139 -68910 6195 -68908
rect 6737 -68910 6793 -68908
<< metal3 >>
rect -52012 8304 -51027 8429
rect -52012 8288 -51678 8304
rect -52012 8232 -51866 8288
rect -51810 8248 -51678 8288
rect -51622 8248 -51027 8304
rect -51810 8232 -51027 8248
rect -52012 8153 -51027 8232
rect -65244 7983 -64259 8149
rect -65244 7967 -64935 7983
rect -65244 7911 -65123 7967
rect -65067 7927 -64935 7967
rect -64879 7927 -64259 7983
rect -65067 7911 -64259 7927
rect -65244 7832 -64259 7911
rect -65244 7798 -64672 7832
rect -65244 7790 -64906 7798
rect -65244 7734 -65107 7790
rect -65051 7742 -64906 7790
rect -64850 7776 -64672 7798
rect -64616 7776 -64259 7832
rect -64850 7770 -64259 7776
rect -64850 7742 -64485 7770
rect -65051 7734 -64485 7742
rect -65244 7714 -64485 7734
rect -64429 7714 -64259 7770
rect -65244 7622 -64259 7714
rect -65244 7609 -64889 7622
rect -65244 7553 -65103 7609
rect -65047 7566 -64889 7609
rect -64833 7613 -64259 7622
rect -64833 7566 -64672 7613
rect -65047 7557 -64672 7566
rect -64616 7585 -64259 7613
rect -64616 7557 -64442 7585
rect -65047 7553 -64442 7557
rect -65244 7529 -64442 7553
rect -64386 7529 -64259 7585
rect -65244 7165 -64259 7529
rect -65244 7149 -64958 7165
rect -65244 7093 -65146 7149
rect -65090 7109 -64958 7149
rect -64902 7109 -64259 7165
rect -65090 7093 -64259 7109
rect -65244 7014 -64259 7093
rect -65244 6980 -64695 7014
rect -65244 6972 -64929 6980
rect -65244 6916 -65130 6972
rect -65074 6924 -64929 6972
rect -64873 6958 -64695 6980
rect -64639 6958 -64259 7014
rect -64873 6952 -64259 6958
rect -64873 6924 -64508 6952
rect -65074 6916 -64508 6924
rect -65244 6896 -64508 6916
rect -64452 6896 -64259 6952
rect -65244 6804 -64259 6896
rect -65244 6791 -64912 6804
rect -65244 6735 -65126 6791
rect -65070 6748 -64912 6791
rect -64856 6795 -64259 6804
rect -64856 6748 -64695 6795
rect -65070 6739 -64695 6748
rect -64639 6767 -64259 6795
rect -64639 6739 -64465 6767
rect -65070 6735 -64465 6739
rect -65244 6711 -64465 6735
rect -64409 6711 -64259 6767
rect -65244 6454 -64259 6711
rect -59062 8065 -58077 8149
rect -59062 8049 -58740 8065
rect -59062 7993 -58928 8049
rect -58872 8009 -58740 8049
rect -58684 8009 -58077 8065
rect -58872 7993 -58077 8009
rect -59062 7914 -58077 7993
rect -59062 7880 -58477 7914
rect -59062 7872 -58711 7880
rect -59062 7816 -58912 7872
rect -58856 7824 -58711 7872
rect -58655 7858 -58477 7880
rect -58421 7858 -58077 7914
rect -58655 7852 -58077 7858
rect -58655 7824 -58290 7852
rect -58856 7816 -58290 7824
rect -59062 7796 -58290 7816
rect -58234 7796 -58077 7852
rect -59062 7704 -58077 7796
rect -59062 7691 -58694 7704
rect -59062 7635 -58908 7691
rect -58852 7648 -58694 7691
rect -58638 7695 -58077 7704
rect -58638 7648 -58477 7695
rect -58852 7639 -58477 7648
rect -58421 7667 -58077 7695
rect -58421 7639 -58247 7667
rect -58852 7635 -58247 7639
rect -59062 7611 -58247 7635
rect -58191 7611 -58077 7667
rect -59062 7185 -58077 7611
rect -59062 7169 -58740 7185
rect -59062 7113 -58928 7169
rect -58872 7129 -58740 7169
rect -58684 7129 -58077 7185
rect -58872 7113 -58077 7129
rect -59062 7034 -58077 7113
rect -59062 7000 -58477 7034
rect -59062 6992 -58711 7000
rect -59062 6936 -58912 6992
rect -58856 6944 -58711 6992
rect -58655 6978 -58477 7000
rect -58421 6978 -58077 7034
rect -58655 6972 -58077 6978
rect -58655 6944 -58290 6972
rect -58856 6936 -58290 6944
rect -59062 6916 -58290 6936
rect -58234 6916 -58077 6972
rect -59062 6824 -58077 6916
rect -59062 6811 -58694 6824
rect -59062 6755 -58908 6811
rect -58852 6768 -58694 6811
rect -58638 6815 -58077 6824
rect -58638 6768 -58477 6815
rect -58852 6759 -58477 6768
rect -58421 6787 -58077 6815
rect -58421 6759 -58247 6787
rect -58852 6755 -58247 6759
rect -59062 6731 -58247 6755
rect -58191 6731 -58077 6787
rect -52012 8119 -51415 8153
rect -52012 8111 -51649 8119
rect -52012 8055 -51850 8111
rect -51794 8063 -51649 8111
rect -51593 8097 -51415 8119
rect -51359 8097 -51027 8153
rect -51593 8091 -51027 8097
rect -51593 8063 -51228 8091
rect -51794 8055 -51228 8063
rect -52012 8035 -51228 8055
rect -51172 8035 -51027 8091
rect -52012 7943 -51027 8035
rect -52012 7930 -51632 7943
rect -52012 7874 -51846 7930
rect -51790 7887 -51632 7930
rect -51576 7934 -51027 7943
rect -51576 7887 -51415 7934
rect -51790 7878 -51415 7887
rect -51359 7906 -51027 7934
rect -51359 7878 -51185 7906
rect -51790 7874 -51185 7878
rect -52012 7850 -51185 7874
rect -51129 7850 -51027 7906
rect -52012 7438 -51027 7850
rect -52012 7422 -51698 7438
rect -52012 7366 -51886 7422
rect -51830 7382 -51698 7422
rect -51642 7382 -51027 7438
rect -51830 7366 -51027 7382
rect -52012 7287 -51027 7366
rect -52012 7253 -51435 7287
rect -52012 7245 -51669 7253
rect -52012 7189 -51870 7245
rect -51814 7197 -51669 7245
rect -51613 7231 -51435 7253
rect -51379 7231 -51027 7287
rect -51613 7225 -51027 7231
rect -51613 7197 -51248 7225
rect -51814 7189 -51248 7197
rect -52012 7169 -51248 7189
rect -51192 7169 -51027 7225
rect -52012 7077 -51027 7169
rect -52012 7064 -51652 7077
rect -52012 7008 -51866 7064
rect -51810 7021 -51652 7064
rect -51596 7068 -51027 7077
rect -51596 7021 -51435 7068
rect -51810 7012 -51435 7021
rect -51379 7040 -51027 7068
rect -51379 7012 -51205 7040
rect -51810 7008 -51205 7012
rect -52012 6984 -51205 7008
rect -51149 6984 -51027 7040
rect -52012 6734 -51027 6984
rect -45475 8158 -44490 8254
rect -45475 8142 -45141 8158
rect -45475 8086 -45329 8142
rect -45273 8102 -45141 8142
rect -45085 8102 -44490 8158
rect -45273 8086 -44490 8102
rect -45475 8007 -44490 8086
rect -45475 7973 -44878 8007
rect -45475 7965 -45112 7973
rect -45475 7909 -45313 7965
rect -45257 7917 -45112 7965
rect -45056 7951 -44878 7973
rect -44822 7951 -44490 8007
rect -45056 7945 -44490 7951
rect -45056 7917 -44691 7945
rect -45257 7909 -44691 7917
rect -45475 7889 -44691 7909
rect -44635 7889 -44490 7945
rect -45475 7797 -44490 7889
rect -45475 7784 -45095 7797
rect -45475 7728 -45309 7784
rect -45253 7741 -45095 7784
rect -45039 7788 -44490 7797
rect -45039 7741 -44878 7788
rect -45253 7732 -44878 7741
rect -44822 7760 -44490 7788
rect -44822 7732 -44648 7760
rect -45253 7728 -44648 7732
rect -45475 7704 -44648 7728
rect -44592 7704 -44490 7760
rect -45475 7226 -44490 7704
rect -45475 7210 -45170 7226
rect -45475 7154 -45358 7210
rect -45302 7170 -45170 7210
rect -45114 7170 -44490 7226
rect -45302 7154 -44490 7170
rect -45475 7075 -44490 7154
rect -45475 7041 -44907 7075
rect -45475 7033 -45141 7041
rect -45475 6977 -45342 7033
rect -45286 6985 -45141 7033
rect -45085 7019 -44907 7041
rect -44851 7019 -44490 7075
rect -45085 7013 -44490 7019
rect -45085 6985 -44720 7013
rect -45286 6977 -44720 6985
rect -45475 6957 -44720 6977
rect -44664 6957 -44490 7013
rect -45475 6865 -44490 6957
rect -45475 6852 -45124 6865
rect -45475 6796 -45338 6852
rect -45282 6809 -45124 6852
rect -45068 6856 -44490 6865
rect -45068 6809 -44907 6856
rect -45282 6800 -44907 6809
rect -44851 6828 -44490 6856
rect -44851 6800 -44677 6828
rect -45282 6796 -44677 6800
rect -45475 6772 -44677 6796
rect -44621 6772 -44490 6828
rect -59062 6454 -58077 6731
rect -45475 6559 -44490 6772
rect -38757 8088 -37772 8237
rect -38757 8072 -38440 8088
rect -38757 8016 -38628 8072
rect -38572 8032 -38440 8072
rect -38384 8032 -37772 8088
rect -38572 8016 -37772 8032
rect -38757 7937 -37772 8016
rect -38757 7903 -38177 7937
rect -38757 7895 -38411 7903
rect -38757 7839 -38612 7895
rect -38556 7847 -38411 7895
rect -38355 7881 -38177 7903
rect -38121 7881 -37772 7937
rect -38355 7875 -37772 7881
rect -38355 7847 -37990 7875
rect -38556 7839 -37990 7847
rect -38757 7819 -37990 7839
rect -37934 7819 -37772 7875
rect -38757 7727 -37772 7819
rect -38757 7714 -38394 7727
rect -38757 7658 -38608 7714
rect -38552 7671 -38394 7714
rect -38338 7718 -37772 7727
rect -38338 7671 -38177 7718
rect -38552 7662 -38177 7671
rect -38121 7690 -37772 7718
rect -38121 7662 -37947 7690
rect -38552 7658 -37947 7662
rect -38757 7634 -37947 7658
rect -37891 7634 -37772 7690
rect -38757 7249 -37772 7634
rect -38757 7233 -38429 7249
rect -38757 7177 -38617 7233
rect -38561 7193 -38429 7233
rect -38373 7193 -37772 7249
rect -38561 7177 -37772 7193
rect -38757 7098 -37772 7177
rect -38757 7064 -38166 7098
rect -38757 7056 -38400 7064
rect -38757 7000 -38601 7056
rect -38545 7008 -38400 7056
rect -38344 7042 -38166 7064
rect -38110 7042 -37772 7098
rect -38344 7036 -37772 7042
rect -38344 7008 -37979 7036
rect -38545 7000 -37979 7008
rect -38757 6980 -37979 7000
rect -37923 6980 -37772 7036
rect -38757 6888 -37772 6980
rect -38757 6875 -38383 6888
rect -38757 6819 -38597 6875
rect -38541 6832 -38383 6875
rect -38327 6879 -37772 6888
rect -38327 6832 -38166 6879
rect -38541 6823 -38166 6832
rect -38110 6851 -37772 6879
rect -38110 6823 -37936 6851
rect -38541 6819 -37936 6823
rect -38757 6795 -37936 6819
rect -37880 6795 -37772 6851
rect -38757 6542 -37772 6795
rect -31724 8147 -30705 8360
rect -31724 8131 -31413 8147
rect -31724 8075 -31601 8131
rect -31545 8091 -31413 8131
rect -31357 8091 -30705 8147
rect -31545 8075 -30705 8091
rect -31724 7996 -30705 8075
rect -31724 7962 -31150 7996
rect -31724 7954 -31384 7962
rect -31724 7898 -31585 7954
rect -31529 7906 -31384 7954
rect -31328 7940 -31150 7962
rect -31094 7940 -30705 7996
rect -31328 7934 -30705 7940
rect -31328 7906 -30963 7934
rect -31529 7898 -30963 7906
rect -31724 7878 -30963 7898
rect -30907 7878 -30705 7934
rect -31724 7786 -30705 7878
rect -31724 7773 -31367 7786
rect -31724 7717 -31581 7773
rect -31525 7730 -31367 7773
rect -31311 7777 -30705 7786
rect -31311 7730 -31150 7777
rect -31525 7721 -31150 7730
rect -31094 7749 -30705 7777
rect -31094 7721 -30920 7749
rect -31525 7717 -30920 7721
rect -31724 7693 -30920 7717
rect -30864 7693 -30705 7749
rect -31724 7255 -30705 7693
rect -31724 7239 -31396 7255
rect -31724 7183 -31584 7239
rect -31528 7199 -31396 7239
rect -31340 7199 -30705 7255
rect -31528 7183 -30705 7199
rect -31724 7104 -30705 7183
rect -31724 7070 -31133 7104
rect -31724 7062 -31367 7070
rect -31724 7006 -31568 7062
rect -31512 7014 -31367 7062
rect -31311 7048 -31133 7070
rect -31077 7048 -30705 7104
rect -31311 7042 -30705 7048
rect -31311 7014 -30946 7042
rect -31512 7006 -30946 7014
rect -31724 6986 -30946 7006
rect -30890 6986 -30705 7042
rect -31724 6894 -30705 6986
rect -31724 6881 -31350 6894
rect -31724 6825 -31564 6881
rect -31508 6838 -31350 6881
rect -31294 6885 -30705 6894
rect -31294 6838 -31133 6885
rect -31508 6829 -31133 6838
rect -31077 6857 -30705 6885
rect -31077 6829 -30903 6857
rect -31508 6825 -30903 6829
rect -31724 6801 -30903 6825
rect -30847 6801 -30705 6857
rect -31724 6507 -30705 6801
rect -24931 8024 -23912 8238
rect -24931 8008 -24562 8024
rect -24931 7952 -24750 8008
rect -24694 7968 -24562 8008
rect -24506 7968 -23912 8024
rect -24694 7952 -23912 7968
rect -24931 7873 -23912 7952
rect -24931 7839 -24299 7873
rect -24931 7831 -24533 7839
rect -24931 7775 -24734 7831
rect -24678 7783 -24533 7831
rect -24477 7817 -24299 7839
rect -24243 7817 -23912 7873
rect -24477 7811 -23912 7817
rect -24477 7783 -24112 7811
rect -24678 7775 -24112 7783
rect -24931 7755 -24112 7775
rect -24056 7755 -23912 7811
rect -24931 7663 -23912 7755
rect -24931 7650 -24516 7663
rect -24931 7594 -24730 7650
rect -24674 7607 -24516 7650
rect -24460 7654 -23912 7663
rect -24460 7607 -24299 7654
rect -24674 7598 -24299 7607
rect -24243 7626 -23912 7654
rect -24243 7598 -24069 7626
rect -24674 7594 -24069 7598
rect -24931 7570 -24069 7594
rect -24013 7570 -23912 7626
rect -24931 7191 -23912 7570
rect -24931 7175 -24573 7191
rect -24931 7119 -24761 7175
rect -24705 7135 -24573 7175
rect -24517 7135 -23912 7191
rect -24705 7119 -23912 7135
rect -24931 7040 -23912 7119
rect -24931 7006 -24310 7040
rect -24931 6998 -24544 7006
rect -24931 6942 -24745 6998
rect -24689 6950 -24544 6998
rect -24488 6984 -24310 7006
rect -24254 6984 -23912 7040
rect -24488 6978 -23912 6984
rect -24488 6950 -24123 6978
rect -24689 6942 -24123 6950
rect -24931 6922 -24123 6942
rect -24067 6922 -23912 6978
rect -24931 6830 -23912 6922
rect -24931 6817 -24527 6830
rect -24931 6761 -24741 6817
rect -24685 6774 -24527 6817
rect -24471 6821 -23912 6830
rect -24471 6774 -24310 6821
rect -24685 6765 -24310 6774
rect -24254 6793 -23912 6821
rect -24254 6765 -24080 6793
rect -24685 6761 -24080 6765
rect -24931 6737 -24080 6761
rect -24024 6737 -23912 6793
rect -24931 6385 -23912 6737
rect -18061 8106 -17042 8354
rect -18061 8090 -17727 8106
rect -18061 8034 -17915 8090
rect -17859 8050 -17727 8090
rect -17671 8050 -17042 8106
rect -17859 8034 -17042 8050
rect -18061 7955 -17042 8034
rect -18061 7921 -17464 7955
rect -18061 7913 -17698 7921
rect -18061 7857 -17899 7913
rect -17843 7865 -17698 7913
rect -17642 7899 -17464 7921
rect -17408 7899 -17042 7955
rect -17642 7893 -17042 7899
rect -17642 7865 -17277 7893
rect -17843 7857 -17277 7865
rect -18061 7837 -17277 7857
rect -17221 7837 -17042 7893
rect -18061 7745 -17042 7837
rect -18061 7732 -17681 7745
rect -18061 7676 -17895 7732
rect -17839 7689 -17681 7732
rect -17625 7736 -17042 7745
rect -17625 7689 -17464 7736
rect -17839 7680 -17464 7689
rect -17408 7708 -17042 7736
rect -17408 7680 -17234 7708
rect -17839 7676 -17234 7680
rect -18061 7652 -17234 7676
rect -17178 7652 -17042 7708
rect -18061 7249 -17042 7652
rect -18061 7233 -17727 7249
rect -18061 7177 -17915 7233
rect -17859 7193 -17727 7233
rect -17671 7193 -17042 7249
rect -17859 7177 -17042 7193
rect -18061 7098 -17042 7177
rect -18061 7064 -17464 7098
rect -18061 7056 -17698 7064
rect -18061 7000 -17899 7056
rect -17843 7008 -17698 7056
rect -17642 7042 -17464 7064
rect -17408 7042 -17042 7098
rect -17642 7036 -17042 7042
rect -17642 7008 -17277 7036
rect -17843 7000 -17277 7008
rect -18061 6980 -17277 7000
rect -17221 6980 -17042 7036
rect -18061 6888 -17042 6980
rect -18061 6875 -17681 6888
rect -18061 6819 -17895 6875
rect -17839 6832 -17681 6875
rect -17625 6879 -17042 6888
rect -17625 6832 -17464 6879
rect -17839 6823 -17464 6832
rect -17408 6851 -17042 6879
rect -17408 6823 -17234 6851
rect -17839 6819 -17234 6823
rect -18061 6795 -17234 6819
rect -17178 6795 -17042 6851
rect -18061 6501 -17042 6795
rect -11069 8193 -10050 8319
rect -11069 8177 -10735 8193
rect -11069 8121 -10923 8177
rect -10867 8137 -10735 8177
rect -10679 8137 -10050 8193
rect -10867 8121 -10050 8137
rect -11069 8042 -10050 8121
rect -11069 8008 -10472 8042
rect -11069 8000 -10706 8008
rect -11069 7944 -10907 8000
rect -10851 7952 -10706 8000
rect -10650 7986 -10472 8008
rect -10416 7986 -10050 8042
rect -10650 7980 -10050 7986
rect -10650 7952 -10285 7980
rect -10851 7944 -10285 7952
rect -11069 7924 -10285 7944
rect -10229 7924 -10050 7980
rect -11069 7832 -10050 7924
rect -11069 7819 -10689 7832
rect -11069 7763 -10903 7819
rect -10847 7776 -10689 7819
rect -10633 7823 -10050 7832
rect -10633 7776 -10472 7823
rect -10847 7767 -10472 7776
rect -10416 7795 -10050 7823
rect -10416 7767 -10242 7795
rect -10847 7763 -10242 7767
rect -11069 7739 -10242 7763
rect -10186 7739 -10050 7795
rect -11069 7208 -10050 7739
rect -11069 7192 -10712 7208
rect -11069 7136 -10900 7192
rect -10844 7152 -10712 7192
rect -10656 7152 -10050 7208
rect -10844 7136 -10050 7152
rect -11069 7057 -10050 7136
rect -11069 7023 -10449 7057
rect -11069 7015 -10683 7023
rect -11069 6959 -10884 7015
rect -10828 6967 -10683 7015
rect -10627 7001 -10449 7023
rect -10393 7001 -10050 7057
rect -10627 6995 -10050 7001
rect -10627 6967 -10262 6995
rect -10828 6959 -10262 6967
rect -11069 6939 -10262 6959
rect -10206 6939 -10050 6995
rect -11069 6847 -10050 6939
rect -11069 6834 -10666 6847
rect -11069 6778 -10880 6834
rect -10824 6791 -10666 6834
rect -10610 6838 -10050 6847
rect -10610 6791 -10449 6838
rect -10824 6782 -10449 6791
rect -10393 6810 -10050 6838
rect -10393 6782 -10219 6810
rect -10824 6778 -10219 6782
rect -11069 6754 -10219 6778
rect -10163 6754 -10050 6810
rect -11069 6466 -10050 6754
rect -3635 8211 -2616 8337
rect -3635 8195 -3295 8211
rect -3635 8139 -3483 8195
rect -3427 8155 -3295 8195
rect -3239 8155 -2616 8211
rect -3427 8139 -2616 8155
rect -3635 8060 -2616 8139
rect -3635 8026 -3032 8060
rect -3635 8018 -3266 8026
rect -3635 7962 -3467 8018
rect -3411 7970 -3266 8018
rect -3210 8004 -3032 8026
rect -2976 8004 -2616 8060
rect -3210 7998 -2616 8004
rect -3210 7970 -2845 7998
rect -3411 7962 -2845 7970
rect -3635 7942 -2845 7962
rect -2789 7942 -2616 7998
rect -3635 7850 -2616 7942
rect -3635 7837 -3249 7850
rect -3635 7781 -3463 7837
rect -3407 7794 -3249 7837
rect -3193 7841 -2616 7850
rect -3193 7794 -3032 7841
rect -3407 7785 -3032 7794
rect -2976 7813 -2616 7841
rect -2976 7785 -2802 7813
rect -3407 7781 -2802 7785
rect -3635 7757 -2802 7781
rect -2746 7757 -2616 7813
rect -3635 7238 -2616 7757
rect -3635 7222 -3225 7238
rect -3635 7166 -3413 7222
rect -3357 7182 -3225 7222
rect -3169 7182 -2616 7238
rect -3357 7166 -2616 7182
rect -3635 7087 -2616 7166
rect -3635 7053 -2962 7087
rect -3635 7045 -3196 7053
rect -3635 6989 -3397 7045
rect -3341 6997 -3196 7045
rect -3140 7031 -2962 7053
rect -2906 7031 -2616 7087
rect -3140 7025 -2616 7031
rect -3140 6997 -2775 7025
rect -3341 6989 -2775 6997
rect -3635 6969 -2775 6989
rect -2719 6969 -2616 7025
rect -3635 6877 -2616 6969
rect -3635 6864 -3179 6877
rect -3635 6808 -3393 6864
rect -3337 6821 -3179 6864
rect -3123 6868 -2616 6877
rect -3123 6821 -2962 6868
rect -3337 6812 -2962 6821
rect -2906 6840 -2616 6868
rect -2906 6812 -2732 6840
rect -3337 6808 -2732 6812
rect -3635 6784 -2732 6808
rect -2676 6784 -2616 6840
rect -3635 6484 -2616 6784
rect 2058 8164 3077 8290
rect 2058 8148 2415 8164
rect 2058 8092 2227 8148
rect 2283 8108 2415 8148
rect 2471 8108 3077 8164
rect 2283 8092 3077 8108
rect 2058 8013 3077 8092
rect 2058 7979 2678 8013
rect 2058 7971 2444 7979
rect 2058 7915 2243 7971
rect 2299 7923 2444 7971
rect 2500 7957 2678 7979
rect 2734 7957 3077 8013
rect 2500 7951 3077 7957
rect 2500 7923 2865 7951
rect 2299 7915 2865 7923
rect 2058 7895 2865 7915
rect 2921 7895 3077 7951
rect 2058 7803 3077 7895
rect 2058 7790 2461 7803
rect 2058 7734 2247 7790
rect 2303 7747 2461 7790
rect 2517 7794 3077 7803
rect 2517 7747 2678 7794
rect 2303 7738 2678 7747
rect 2734 7766 3077 7794
rect 2734 7738 2908 7766
rect 2303 7734 2908 7738
rect 2058 7710 2908 7734
rect 2964 7710 3077 7766
rect 2058 7139 3077 7710
rect 2058 7123 2444 7139
rect 2058 7067 2256 7123
rect 2312 7083 2444 7123
rect 2500 7083 3077 7139
rect 2312 7067 3077 7083
rect 2058 6988 3077 7067
rect 2058 6954 2707 6988
rect 2058 6946 2473 6954
rect 2058 6890 2272 6946
rect 2328 6898 2473 6946
rect 2529 6932 2707 6954
rect 2763 6932 3077 6988
rect 2529 6926 3077 6932
rect 2529 6898 2894 6926
rect 2328 6890 2894 6898
rect 2058 6870 2894 6890
rect 2950 6870 3077 6926
rect 2058 6778 3077 6870
rect 2058 6765 2490 6778
rect 2058 6709 2276 6765
rect 2332 6722 2490 6765
rect 2546 6769 3077 6778
rect 2546 6722 2707 6769
rect 2332 6713 2707 6722
rect 2763 6741 3077 6769
rect 2763 6713 2937 6741
rect 2332 6709 2937 6713
rect 2058 6685 2937 6709
rect 2993 6685 3077 6741
rect 2058 6437 3077 6685
rect -61751 -68320 -60887 -68247
rect -61751 -68336 -61490 -68320
rect -61751 -68392 -61678 -68336
rect -61622 -68376 -61490 -68336
rect -61434 -68376 -60887 -68320
rect -61622 -68392 -60887 -68376
rect -61751 -68471 -60887 -68392
rect -61751 -68505 -61227 -68471
rect -61751 -68513 -61461 -68505
rect -61751 -68569 -61662 -68513
rect -61606 -68561 -61461 -68513
rect -61405 -68527 -61227 -68505
rect -61171 -68527 -60887 -68471
rect -61405 -68533 -60887 -68527
rect -61405 -68561 -61040 -68533
rect -61606 -68569 -61040 -68561
rect -61751 -68589 -61040 -68569
rect -60984 -68589 -60887 -68533
rect -61751 -68681 -60887 -68589
rect -61751 -68694 -61444 -68681
rect -61751 -68750 -61658 -68694
rect -61602 -68737 -61444 -68694
rect -61388 -68690 -60887 -68681
rect -61388 -68737 -61227 -68690
rect -61602 -68746 -61227 -68737
rect -61171 -68718 -60887 -68690
rect -61171 -68746 -60997 -68718
rect -61602 -68750 -60997 -68746
rect -61751 -68774 -60997 -68750
rect -60941 -68774 -60887 -68718
rect -61751 -68934 -60887 -68774
rect -55242 -68379 -54186 -68282
rect -55242 -68435 -54944 -68379
rect -54888 -68435 -54769 -68379
rect -54713 -68435 -54567 -68379
rect -54511 -68435 -54186 -68379
rect -55242 -68619 -54186 -68435
rect -55242 -68644 -54725 -68619
rect -55242 -68646 -54925 -68644
rect -55242 -68702 -55157 -68646
rect -55101 -68700 -54925 -68646
rect -54869 -68675 -54725 -68644
rect -54669 -68634 -54186 -68619
rect -54669 -68650 -54294 -68634
rect -54669 -68675 -54507 -68650
rect -54869 -68700 -54507 -68675
rect -55101 -68702 -54507 -68700
rect -55242 -68706 -54507 -68702
rect -54451 -68690 -54294 -68650
rect -54238 -68690 -54186 -68634
rect -54451 -68706 -54186 -68690
rect -55242 -68863 -54186 -68706
rect -55242 -68867 -54696 -68863
rect -55242 -68923 -54921 -68867
rect -54865 -68919 -54696 -68867
rect -54640 -68869 -54186 -68863
rect -54640 -68919 -54438 -68869
rect -54865 -68923 -54438 -68919
rect -55242 -68925 -54438 -68923
rect -54382 -68925 -54186 -68869
rect -48439 -68369 -47230 -68311
rect -48439 -68425 -48168 -68369
rect -48112 -68425 -47987 -68369
rect -47931 -68375 -47230 -68369
rect -47931 -68425 -47783 -68375
rect -48439 -68431 -47783 -68425
rect -47727 -68431 -47230 -68375
rect -48439 -68569 -47230 -68431
rect -48439 -68575 -47916 -68569
rect -48439 -68631 -48152 -68575
rect -48096 -68625 -47916 -68575
rect -47860 -68584 -47230 -68569
rect -47860 -68625 -47656 -68584
rect -48096 -68631 -47656 -68625
rect -48439 -68640 -47656 -68631
rect -47600 -68640 -47230 -68584
rect -48439 -68786 -47230 -68640
rect -48439 -68842 -48212 -68786
rect -48156 -68790 -47230 -68786
rect -48156 -68842 -47970 -68790
rect -48439 -68846 -47970 -68842
rect -47914 -68846 -47770 -68790
rect -47714 -68800 -47230 -68790
rect -47714 -68846 -47466 -68800
rect -48439 -68856 -47466 -68846
rect -47410 -68856 -47230 -68800
rect -48439 -68909 -47230 -68856
rect -41649 -68369 -40440 -68326
rect -21096 -68350 -20092 -68263
rect -41649 -68373 -41151 -68369
rect -41649 -68429 -41332 -68373
rect -41276 -68425 -41151 -68373
rect -41095 -68379 -40440 -68369
rect -41095 -68425 -40951 -68379
rect -41276 -68429 -40951 -68425
rect -41649 -68435 -40951 -68429
rect -40895 -68435 -40440 -68379
rect -41649 -68542 -40440 -68435
rect -41649 -68581 -41330 -68542
rect -41649 -68637 -41517 -68581
rect -41461 -68598 -41330 -68581
rect -41274 -68546 -40440 -68542
rect -41274 -68556 -40890 -68546
rect -41274 -68598 -41117 -68556
rect -41461 -68612 -41117 -68598
rect -41061 -68602 -40890 -68556
rect -40834 -68569 -40440 -68546
rect -40834 -68602 -40694 -68569
rect -41061 -68612 -40694 -68602
rect -41461 -68625 -40694 -68612
rect -40638 -68625 -40440 -68569
rect -41461 -68637 -40440 -68625
rect -41649 -68742 -40440 -68637
rect -41649 -68759 -41084 -68742
rect -41649 -68815 -41317 -68759
rect -41261 -68798 -41084 -68759
rect -41028 -68754 -40440 -68742
rect -41028 -68798 -40836 -68754
rect -41261 -68810 -40836 -68798
rect -40780 -68810 -40440 -68754
rect -41261 -68815 -40440 -68810
rect -41649 -68924 -40440 -68815
rect -34904 -68408 -33695 -68353
rect -34904 -68464 -34577 -68408
rect -34521 -68415 -33695 -68408
rect -34521 -68464 -34396 -68415
rect -34904 -68471 -34396 -68464
rect -34340 -68471 -34221 -68415
rect -34165 -68471 -33695 -68415
rect -34904 -68625 -33695 -68471
rect -34904 -68631 -34000 -68625
rect -34904 -68650 -34560 -68631
rect -34904 -68706 -34819 -68650
rect -34763 -68687 -34560 -68650
rect -34504 -68687 -34329 -68631
rect -34273 -68681 -34000 -68631
rect -33944 -68681 -33695 -68625
rect -34273 -68687 -33695 -68681
rect -34763 -68706 -33695 -68687
rect -34904 -68834 -33695 -68706
rect -34904 -68848 -33843 -68834
rect -34904 -68904 -34581 -68848
rect -34525 -68904 -34346 -68848
rect -34290 -68852 -33843 -68848
rect -34290 -68904 -34106 -68852
rect -34904 -68908 -34106 -68904
rect -34050 -68890 -33843 -68852
rect -33787 -68890 -33695 -68834
rect -34050 -68908 -33695 -68890
rect -55242 -68970 -54186 -68925
rect -34904 -68951 -33695 -68908
rect -28030 -68388 -26900 -68350
rect -28030 -68444 -27727 -68388
rect -27671 -68395 -26900 -68388
rect -27671 -68444 -27546 -68395
rect -28030 -68451 -27546 -68444
rect -27490 -68451 -27371 -68395
rect -27315 -68451 -26900 -68395
rect -28030 -68605 -26900 -68451
rect -28030 -68611 -27150 -68605
rect -28030 -68630 -27710 -68611
rect -28030 -68686 -27969 -68630
rect -27913 -68667 -27710 -68630
rect -27654 -68667 -27479 -68611
rect -27423 -68661 -27150 -68611
rect -27094 -68661 -26900 -68605
rect -27423 -68667 -26900 -68661
rect -27913 -68686 -26900 -68667
rect -28030 -68814 -26900 -68686
rect -28030 -68828 -26993 -68814
rect -28030 -68884 -27731 -68828
rect -27675 -68884 -27496 -68828
rect -27440 -68832 -26993 -68828
rect -27440 -68884 -27256 -68832
rect -28030 -68888 -27256 -68884
rect -27200 -68870 -26993 -68832
rect -26937 -68870 -26900 -68814
rect -27200 -68888 -26900 -68870
rect -28030 -68930 -26900 -68888
rect -21096 -68388 -19960 -68350
rect -21096 -68444 -20787 -68388
rect -20731 -68395 -19960 -68388
rect -20731 -68444 -20606 -68395
rect -21096 -68451 -20606 -68444
rect -20550 -68451 -20431 -68395
rect -20375 -68451 -19960 -68395
rect -21096 -68605 -19960 -68451
rect -21096 -68611 -20210 -68605
rect -21096 -68630 -20770 -68611
rect -21096 -68686 -21029 -68630
rect -20973 -68667 -20770 -68630
rect -20714 -68667 -20539 -68611
rect -20483 -68661 -20210 -68611
rect -20154 -68661 -19960 -68605
rect -20483 -68667 -19960 -68661
rect -20973 -68686 -19960 -68667
rect -21096 -68814 -19960 -68686
rect -21096 -68828 -20053 -68814
rect -21096 -68884 -20791 -68828
rect -20735 -68884 -20556 -68828
rect -20500 -68832 -20053 -68828
rect -20500 -68884 -20316 -68832
rect -21096 -68888 -20316 -68884
rect -20260 -68870 -20053 -68832
rect -19997 -68870 -19960 -68814
rect -20260 -68888 -19960 -68870
rect -21096 -68930 -19960 -68888
rect -14409 -68381 -13405 -68255
rect -14409 -68437 -14124 -68381
rect -14068 -68386 -13405 -68381
rect -14068 -68437 -13945 -68386
rect -14409 -68442 -13945 -68437
rect -13889 -68442 -13762 -68386
rect -13706 -68442 -13405 -68386
rect -14409 -68634 -13405 -68442
rect -14409 -68638 -13637 -68634
rect -14409 -68644 -13845 -68638
rect -14409 -68650 -14037 -68644
rect -14409 -68706 -14262 -68650
rect -14206 -68700 -14037 -68650
rect -13981 -68694 -13845 -68644
rect -13789 -68690 -13637 -68638
rect -13581 -68690 -13405 -68634
rect -13789 -68694 -13405 -68690
rect -13981 -68700 -13405 -68694
rect -14206 -68706 -13405 -68700
rect -14409 -68848 -13405 -68706
rect -14409 -68904 -14199 -68848
rect -14143 -68904 -13980 -68848
rect -13924 -68904 -13791 -68848
rect -13735 -68904 -13543 -68848
rect -13487 -68904 -13405 -68848
rect -21096 -68951 -20092 -68930
rect -14409 -68943 -13405 -68904
rect -7481 -68361 -6477 -68255
rect -7481 -68417 -7286 -68361
rect -7230 -68417 -7111 -68361
rect -7055 -68417 -6921 -68361
rect -6865 -68417 -6477 -68361
rect -7481 -68611 -6477 -68417
rect -7481 -68617 -6648 -68611
rect -7481 -68623 -6909 -68617
rect -7481 -68629 -7129 -68623
rect -7481 -68685 -7402 -68629
rect -7346 -68679 -7129 -68629
rect -7073 -68673 -6909 -68623
rect -6853 -68667 -6648 -68617
rect -6592 -68667 -6477 -68611
rect -6853 -68673 -6477 -68667
rect -7073 -68679 -6477 -68673
rect -7346 -68685 -6477 -68679
rect -7481 -68846 -6477 -68685
rect -7481 -68852 -6723 -68846
rect -7481 -68854 -7152 -68852
rect -7481 -68910 -7367 -68854
rect -7311 -68908 -7152 -68854
rect -7096 -68908 -6934 -68852
rect -6878 -68902 -6723 -68852
rect -6667 -68902 -6477 -68846
rect -6878 -68908 -6477 -68902
rect -7311 -68910 -6477 -68908
rect -7481 -68943 -6477 -68910
rect -676 -68358 328 -68259
rect -676 -68361 -70 -68358
rect -676 -68417 -476 -68361
rect -420 -68365 -70 -68361
rect -420 -68417 -283 -68365
rect -676 -68421 -283 -68417
rect -227 -68414 -70 -68365
rect -14 -68414 328 -68358
rect -227 -68421 328 -68414
rect -676 -68594 328 -68421
rect -676 -68598 145 -68594
rect -676 -68602 -345 -68598
rect -676 -68658 -595 -68602
rect -539 -68654 -345 -68602
rect -289 -68654 -112 -68598
rect -56 -68650 145 -68598
rect 201 -68650 328 -68594
rect -56 -68654 328 -68650
rect -539 -68658 328 -68654
rect -676 -68848 328 -68658
rect -676 -68852 -308 -68848
rect -676 -68908 -566 -68852
rect -510 -68904 -308 -68852
rect -252 -68852 328 -68848
rect -252 -68904 -70 -68852
rect -510 -68908 -70 -68904
rect -14 -68859 328 -68852
rect -14 -68908 184 -68859
rect -676 -68915 184 -68908
rect 240 -68915 328 -68859
rect -676 -68947 328 -68915
rect 5835 -68352 6839 -68257
rect 5835 -68408 6318 -68352
rect 6374 -68408 6506 -68352
rect 6562 -68358 6839 -68352
rect 6562 -68408 6708 -68358
rect 5835 -68414 6708 -68408
rect 6764 -68414 6839 -68358
rect 5835 -68573 6839 -68414
rect 5835 -68629 6143 -68573
rect 6199 -68577 6606 -68573
rect 6199 -68629 6395 -68577
rect 5835 -68633 6395 -68629
rect 6451 -68629 6606 -68577
rect 6662 -68629 6839 -68573
rect 6451 -68633 6839 -68629
rect 5835 -68688 6839 -68633
rect 5835 -68744 5931 -68688
rect 5987 -68744 6839 -68688
rect 5835 -68852 6839 -68744
rect 5835 -68854 6327 -68852
rect 5835 -68910 6139 -68854
rect 6195 -68908 6327 -68854
rect 6383 -68908 6533 -68852
rect 6589 -68854 6839 -68852
rect 6589 -68908 6737 -68854
rect 6195 -68910 6737 -68908
rect 6793 -68910 6839 -68854
rect 5835 -68945 6839 -68910
<< via3 >>
rect -51866 8232 -51810 8288
rect -51678 8248 -51622 8304
rect -65123 7911 -65067 7967
rect -64935 7927 -64879 7983
rect -65107 7734 -65051 7790
rect -64906 7742 -64850 7798
rect -64672 7776 -64616 7832
rect -64485 7714 -64429 7770
rect -65103 7553 -65047 7609
rect -64889 7566 -64833 7622
rect -64672 7557 -64616 7613
rect -64442 7529 -64386 7585
rect -65146 7093 -65090 7149
rect -64958 7109 -64902 7165
rect -65130 6916 -65074 6972
rect -64929 6924 -64873 6980
rect -64695 6958 -64639 7014
rect -64508 6896 -64452 6952
rect -65126 6735 -65070 6791
rect -64912 6748 -64856 6804
rect -64695 6739 -64639 6795
rect -64465 6711 -64409 6767
rect -58928 7993 -58872 8049
rect -58740 8009 -58684 8065
rect -58912 7816 -58856 7872
rect -58711 7824 -58655 7880
rect -58477 7858 -58421 7914
rect -58290 7796 -58234 7852
rect -58908 7635 -58852 7691
rect -58694 7648 -58638 7704
rect -58477 7639 -58421 7695
rect -58247 7611 -58191 7667
rect -58928 7113 -58872 7169
rect -58740 7129 -58684 7185
rect -58912 6936 -58856 6992
rect -58711 6944 -58655 7000
rect -58477 6978 -58421 7034
rect -58290 6916 -58234 6972
rect -58908 6755 -58852 6811
rect -58694 6768 -58638 6824
rect -58477 6759 -58421 6815
rect -58247 6731 -58191 6787
rect -51850 8055 -51794 8111
rect -51649 8063 -51593 8119
rect -51415 8097 -51359 8153
rect -51228 8035 -51172 8091
rect -51846 7874 -51790 7930
rect -51632 7887 -51576 7943
rect -51415 7878 -51359 7934
rect -51185 7850 -51129 7906
rect -51886 7366 -51830 7422
rect -51698 7382 -51642 7438
rect -51870 7189 -51814 7245
rect -51669 7197 -51613 7253
rect -51435 7231 -51379 7287
rect -51248 7169 -51192 7225
rect -51866 7008 -51810 7064
rect -51652 7021 -51596 7077
rect -51435 7012 -51379 7068
rect -51205 6984 -51149 7040
rect -45329 8086 -45273 8142
rect -45141 8102 -45085 8158
rect -45313 7909 -45257 7965
rect -45112 7917 -45056 7973
rect -44878 7951 -44822 8007
rect -44691 7889 -44635 7945
rect -45309 7728 -45253 7784
rect -45095 7741 -45039 7797
rect -44878 7732 -44822 7788
rect -44648 7704 -44592 7760
rect -45358 7154 -45302 7210
rect -45170 7170 -45114 7226
rect -45342 6977 -45286 7033
rect -45141 6985 -45085 7041
rect -44907 7019 -44851 7075
rect -44720 6957 -44664 7013
rect -45338 6796 -45282 6852
rect -45124 6809 -45068 6865
rect -44907 6800 -44851 6856
rect -44677 6772 -44621 6828
rect -38628 8016 -38572 8072
rect -38440 8032 -38384 8088
rect -38612 7839 -38556 7895
rect -38411 7847 -38355 7903
rect -38177 7881 -38121 7937
rect -37990 7819 -37934 7875
rect -38608 7658 -38552 7714
rect -38394 7671 -38338 7727
rect -38177 7662 -38121 7718
rect -37947 7634 -37891 7690
rect -38617 7177 -38561 7233
rect -38429 7193 -38373 7249
rect -38601 7000 -38545 7056
rect -38400 7008 -38344 7064
rect -38166 7042 -38110 7098
rect -37979 6980 -37923 7036
rect -38597 6819 -38541 6875
rect -38383 6832 -38327 6888
rect -38166 6823 -38110 6879
rect -37936 6795 -37880 6851
rect -31601 8075 -31545 8131
rect -31413 8091 -31357 8147
rect -31585 7898 -31529 7954
rect -31384 7906 -31328 7962
rect -31150 7940 -31094 7996
rect -30963 7878 -30907 7934
rect -31581 7717 -31525 7773
rect -31367 7730 -31311 7786
rect -31150 7721 -31094 7777
rect -30920 7693 -30864 7749
rect -31584 7183 -31528 7239
rect -31396 7199 -31340 7255
rect -31568 7006 -31512 7062
rect -31367 7014 -31311 7070
rect -31133 7048 -31077 7104
rect -30946 6986 -30890 7042
rect -31564 6825 -31508 6881
rect -31350 6838 -31294 6894
rect -31133 6829 -31077 6885
rect -30903 6801 -30847 6857
rect -24750 7952 -24694 8008
rect -24562 7968 -24506 8024
rect -24734 7775 -24678 7831
rect -24533 7783 -24477 7839
rect -24299 7817 -24243 7873
rect -24112 7755 -24056 7811
rect -24730 7594 -24674 7650
rect -24516 7607 -24460 7663
rect -24299 7598 -24243 7654
rect -24069 7570 -24013 7626
rect -24761 7119 -24705 7175
rect -24573 7135 -24517 7191
rect -24745 6942 -24689 6998
rect -24544 6950 -24488 7006
rect -24310 6984 -24254 7040
rect -24123 6922 -24067 6978
rect -24741 6761 -24685 6817
rect -24527 6774 -24471 6830
rect -24310 6765 -24254 6821
rect -24080 6737 -24024 6793
rect -17915 8034 -17859 8090
rect -17727 8050 -17671 8106
rect -17899 7857 -17843 7913
rect -17698 7865 -17642 7921
rect -17464 7899 -17408 7955
rect -17277 7837 -17221 7893
rect -17895 7676 -17839 7732
rect -17681 7689 -17625 7745
rect -17464 7680 -17408 7736
rect -17234 7652 -17178 7708
rect -17915 7177 -17859 7233
rect -17727 7193 -17671 7249
rect -17899 7000 -17843 7056
rect -17698 7008 -17642 7064
rect -17464 7042 -17408 7098
rect -17277 6980 -17221 7036
rect -17895 6819 -17839 6875
rect -17681 6832 -17625 6888
rect -17464 6823 -17408 6879
rect -17234 6795 -17178 6851
rect -10923 8121 -10867 8177
rect -10735 8137 -10679 8193
rect -10907 7944 -10851 8000
rect -10706 7952 -10650 8008
rect -10472 7986 -10416 8042
rect -10285 7924 -10229 7980
rect -10903 7763 -10847 7819
rect -10689 7776 -10633 7832
rect -10472 7767 -10416 7823
rect -10242 7739 -10186 7795
rect -10900 7136 -10844 7192
rect -10712 7152 -10656 7208
rect -10884 6959 -10828 7015
rect -10683 6967 -10627 7023
rect -10449 7001 -10393 7057
rect -10262 6939 -10206 6995
rect -10880 6778 -10824 6834
rect -10666 6791 -10610 6847
rect -10449 6782 -10393 6838
rect -10219 6754 -10163 6810
rect -3483 8139 -3427 8195
rect -3295 8155 -3239 8211
rect -3467 7962 -3411 8018
rect -3266 7970 -3210 8026
rect -3032 8004 -2976 8060
rect -2845 7942 -2789 7998
rect -3463 7781 -3407 7837
rect -3249 7794 -3193 7850
rect -3032 7785 -2976 7841
rect -2802 7757 -2746 7813
rect -3413 7166 -3357 7222
rect -3225 7182 -3169 7238
rect -3397 6989 -3341 7045
rect -3196 6997 -3140 7053
rect -2962 7031 -2906 7087
rect -2775 6969 -2719 7025
rect -3393 6808 -3337 6864
rect -3179 6821 -3123 6877
rect -2962 6812 -2906 6868
rect -2732 6784 -2676 6840
rect 2227 8092 2283 8148
rect 2415 8108 2471 8164
rect 2243 7915 2299 7971
rect 2444 7923 2500 7979
rect 2678 7957 2734 8013
rect 2865 7895 2921 7951
rect 2247 7734 2303 7790
rect 2461 7747 2517 7803
rect 2678 7738 2734 7794
rect 2908 7710 2964 7766
rect 2256 7067 2312 7123
rect 2444 7083 2500 7139
rect 2272 6890 2328 6946
rect 2473 6898 2529 6954
rect 2707 6932 2763 6988
rect 2894 6870 2950 6926
rect 2276 6709 2332 6765
rect 2490 6722 2546 6778
rect 2707 6713 2763 6769
rect 2937 6685 2993 6741
rect -61678 -68392 -61622 -68336
rect -61490 -68376 -61434 -68320
rect -61662 -68569 -61606 -68513
rect -61461 -68561 -61405 -68505
rect -61227 -68527 -61171 -68471
rect -61040 -68589 -60984 -68533
rect -61658 -68750 -61602 -68694
rect -61444 -68737 -61388 -68681
rect -61227 -68746 -61171 -68690
rect -60997 -68774 -60941 -68718
rect -54944 -68435 -54888 -68379
rect -54769 -68435 -54713 -68379
rect -54567 -68435 -54511 -68379
rect -55157 -68702 -55101 -68646
rect -54925 -68700 -54869 -68644
rect -54725 -68675 -54669 -68619
rect -54507 -68706 -54451 -68650
rect -54294 -68690 -54238 -68634
rect -54921 -68923 -54865 -68867
rect -54696 -68919 -54640 -68863
rect -54438 -68925 -54382 -68869
rect -48168 -68425 -48112 -68369
rect -47987 -68425 -47931 -68369
rect -47783 -68431 -47727 -68375
rect -48152 -68631 -48096 -68575
rect -47916 -68625 -47860 -68569
rect -47656 -68640 -47600 -68584
rect -48212 -68842 -48156 -68786
rect -47970 -68846 -47914 -68790
rect -47770 -68846 -47714 -68790
rect -47466 -68856 -47410 -68800
rect -41332 -68429 -41276 -68373
rect -41151 -68425 -41095 -68369
rect -40951 -68435 -40895 -68379
rect -41517 -68637 -41461 -68581
rect -41330 -68598 -41274 -68542
rect -41117 -68612 -41061 -68556
rect -40890 -68602 -40834 -68546
rect -40694 -68625 -40638 -68569
rect -41317 -68815 -41261 -68759
rect -41084 -68798 -41028 -68742
rect -40836 -68810 -40780 -68754
rect -34577 -68464 -34521 -68408
rect -34396 -68471 -34340 -68415
rect -34221 -68471 -34165 -68415
rect -34819 -68706 -34763 -68650
rect -34560 -68687 -34504 -68631
rect -34329 -68687 -34273 -68631
rect -34000 -68681 -33944 -68625
rect -34581 -68904 -34525 -68848
rect -34346 -68904 -34290 -68848
rect -34106 -68908 -34050 -68852
rect -33843 -68890 -33787 -68834
rect -27727 -68444 -27671 -68388
rect -27546 -68451 -27490 -68395
rect -27371 -68451 -27315 -68395
rect -27969 -68686 -27913 -68630
rect -27710 -68667 -27654 -68611
rect -27479 -68667 -27423 -68611
rect -27150 -68661 -27094 -68605
rect -27731 -68884 -27675 -68828
rect -27496 -68884 -27440 -68828
rect -27256 -68888 -27200 -68832
rect -26993 -68870 -26937 -68814
rect -20787 -68444 -20731 -68388
rect -20606 -68451 -20550 -68395
rect -20431 -68451 -20375 -68395
rect -21029 -68686 -20973 -68630
rect -20770 -68667 -20714 -68611
rect -20539 -68667 -20483 -68611
rect -20210 -68661 -20154 -68605
rect -20791 -68884 -20735 -68828
rect -20556 -68884 -20500 -68828
rect -20316 -68888 -20260 -68832
rect -20053 -68870 -19997 -68814
rect -14124 -68437 -14068 -68381
rect -13945 -68442 -13889 -68386
rect -13762 -68442 -13706 -68386
rect -14262 -68706 -14206 -68650
rect -14037 -68700 -13981 -68644
rect -13845 -68694 -13789 -68638
rect -13637 -68690 -13581 -68634
rect -14199 -68904 -14143 -68848
rect -13980 -68904 -13924 -68848
rect -13791 -68904 -13735 -68848
rect -13543 -68904 -13487 -68848
rect -7286 -68417 -7230 -68361
rect -7111 -68417 -7055 -68361
rect -6921 -68417 -6865 -68361
rect -7402 -68685 -7346 -68629
rect -7129 -68679 -7073 -68623
rect -6909 -68673 -6853 -68617
rect -6648 -68667 -6592 -68611
rect -7367 -68910 -7311 -68854
rect -7152 -68908 -7096 -68852
rect -6934 -68908 -6878 -68852
rect -6723 -68902 -6667 -68846
rect -476 -68417 -420 -68361
rect -283 -68421 -227 -68365
rect -70 -68414 -14 -68358
rect -595 -68658 -539 -68602
rect -345 -68654 -289 -68598
rect -112 -68654 -56 -68598
rect 145 -68650 201 -68594
rect -566 -68908 -510 -68852
rect -308 -68904 -252 -68848
rect -70 -68908 -14 -68852
rect 184 -68915 240 -68859
rect 6318 -68408 6374 -68352
rect 6506 -68408 6562 -68352
rect 6708 -68414 6764 -68358
rect 6143 -68629 6199 -68573
rect 6395 -68633 6451 -68577
rect 6606 -68629 6662 -68573
rect 5931 -68744 5987 -68688
rect 6139 -68910 6195 -68854
rect 6327 -68908 6383 -68852
rect 6533 -68908 6589 -68852
rect 6737 -68910 6793 -68854
<< metal4 >>
rect -52012 8306 -51027 8429
rect -52012 8290 -51678 8306
rect -52012 8232 -51866 8290
rect -51810 8248 -51678 8290
rect -51622 8248 -51027 8306
rect -51810 8232 -51027 8248
rect -52012 8155 -51027 8232
rect -65244 7985 -64259 8149
rect -65244 7969 -64935 7985
rect -65244 7911 -65123 7969
rect -65067 7927 -64935 7969
rect -64879 7927 -64259 7985
rect -65067 7911 -64259 7927
rect -65244 7834 -64259 7911
rect -65244 7800 -64672 7834
rect -65244 7792 -64906 7800
rect -65244 7734 -65107 7792
rect -65051 7742 -64906 7792
rect -64850 7776 -64672 7800
rect -64616 7776 -64259 7834
rect -64850 7772 -64259 7776
rect -64850 7742 -64485 7772
rect -65051 7734 -64485 7742
rect -65244 7714 -64485 7734
rect -64429 7714 -64259 7772
rect -65244 7624 -64259 7714
rect -65244 7611 -64889 7624
rect -65244 7553 -65103 7611
rect -65047 7566 -64889 7611
rect -64833 7615 -64259 7624
rect -64833 7566 -64672 7615
rect -65047 7557 -64672 7566
rect -64616 7587 -64259 7615
rect -64616 7557 -64442 7587
rect -65047 7553 -64442 7557
rect -65244 7529 -64442 7553
rect -64386 7529 -64259 7587
rect -65244 7167 -64259 7529
rect -65244 7151 -64958 7167
rect -65244 7093 -65146 7151
rect -65090 7109 -64958 7151
rect -64902 7109 -64259 7167
rect -65090 7093 -64259 7109
rect -65244 7016 -64259 7093
rect -65244 6982 -64695 7016
rect -65244 6974 -64929 6982
rect -65244 6916 -65130 6974
rect -65074 6924 -64929 6974
rect -64873 6958 -64695 6982
rect -64639 6958 -64259 7016
rect -64873 6954 -64259 6958
rect -64873 6924 -64508 6954
rect -65074 6916 -64508 6924
rect -65244 6896 -64508 6916
rect -64452 6896 -64259 6954
rect -65244 6806 -64259 6896
rect -65244 6793 -64912 6806
rect -65244 6735 -65126 6793
rect -65070 6748 -64912 6793
rect -64856 6797 -64259 6806
rect -64856 6748 -64695 6797
rect -65070 6739 -64695 6748
rect -64639 6769 -64259 6797
rect -64639 6739 -64465 6769
rect -65070 6735 -64465 6739
rect -65244 6711 -64465 6735
rect -64409 6711 -64259 6769
rect -65244 6454 -64259 6711
rect -59062 8067 -58077 8149
rect -59062 8051 -58740 8067
rect -59062 7993 -58928 8051
rect -58872 8009 -58740 8051
rect -58684 8009 -58077 8067
rect -58872 7993 -58077 8009
rect -59062 7916 -58077 7993
rect -59062 7882 -58477 7916
rect -59062 7874 -58711 7882
rect -59062 7816 -58912 7874
rect -58856 7824 -58711 7874
rect -58655 7858 -58477 7882
rect -58421 7858 -58077 7916
rect -58655 7854 -58077 7858
rect -58655 7824 -58290 7854
rect -58856 7816 -58290 7824
rect -59062 7796 -58290 7816
rect -58234 7796 -58077 7854
rect -59062 7706 -58077 7796
rect -59062 7693 -58694 7706
rect -59062 7635 -58908 7693
rect -58852 7648 -58694 7693
rect -58638 7697 -58077 7706
rect -58638 7648 -58477 7697
rect -58852 7639 -58477 7648
rect -58421 7669 -58077 7697
rect -58421 7639 -58247 7669
rect -58852 7635 -58247 7639
rect -59062 7611 -58247 7635
rect -58191 7611 -58077 7669
rect -59062 7187 -58077 7611
rect -59062 7171 -58740 7187
rect -59062 7113 -58928 7171
rect -58872 7129 -58740 7171
rect -58684 7129 -58077 7187
rect -58872 7113 -58077 7129
rect -59062 7036 -58077 7113
rect -59062 7002 -58477 7036
rect -59062 6994 -58711 7002
rect -59062 6936 -58912 6994
rect -58856 6944 -58711 6994
rect -58655 6978 -58477 7002
rect -58421 6978 -58077 7036
rect -58655 6974 -58077 6978
rect -58655 6944 -58290 6974
rect -58856 6936 -58290 6944
rect -59062 6916 -58290 6936
rect -58234 6916 -58077 6974
rect -59062 6826 -58077 6916
rect -59062 6813 -58694 6826
rect -59062 6755 -58908 6813
rect -58852 6768 -58694 6813
rect -58638 6817 -58077 6826
rect -58638 6768 -58477 6817
rect -58852 6759 -58477 6768
rect -58421 6789 -58077 6817
rect -58421 6759 -58247 6789
rect -58852 6755 -58247 6759
rect -59062 6731 -58247 6755
rect -58191 6731 -58077 6789
rect -52012 8121 -51415 8155
rect -52012 8113 -51649 8121
rect -52012 8055 -51850 8113
rect -51794 8063 -51649 8113
rect -51593 8097 -51415 8121
rect -51359 8097 -51027 8155
rect -51593 8093 -51027 8097
rect -51593 8063 -51228 8093
rect -51794 8055 -51228 8063
rect -52012 8035 -51228 8055
rect -51172 8035 -51027 8093
rect -52012 7945 -51027 8035
rect -52012 7932 -51632 7945
rect -52012 7874 -51846 7932
rect -51790 7887 -51632 7932
rect -51576 7936 -51027 7945
rect -51576 7887 -51415 7936
rect -51790 7878 -51415 7887
rect -51359 7908 -51027 7936
rect -51359 7878 -51185 7908
rect -51790 7874 -51185 7878
rect -52012 7850 -51185 7874
rect -51129 7850 -51027 7908
rect -52012 7440 -51027 7850
rect -52012 7424 -51698 7440
rect -52012 7366 -51886 7424
rect -51830 7382 -51698 7424
rect -51642 7382 -51027 7440
rect -51830 7366 -51027 7382
rect -52012 7289 -51027 7366
rect -52012 7255 -51435 7289
rect -52012 7247 -51669 7255
rect -52012 7189 -51870 7247
rect -51814 7197 -51669 7247
rect -51613 7231 -51435 7255
rect -51379 7231 -51027 7289
rect -51613 7227 -51027 7231
rect -51613 7197 -51248 7227
rect -51814 7189 -51248 7197
rect -52012 7169 -51248 7189
rect -51192 7169 -51027 7227
rect -52012 7079 -51027 7169
rect -52012 7066 -51652 7079
rect -52012 7008 -51866 7066
rect -51810 7021 -51652 7066
rect -51596 7070 -51027 7079
rect -51596 7021 -51435 7070
rect -51810 7012 -51435 7021
rect -51379 7042 -51027 7070
rect -51379 7012 -51205 7042
rect -51810 7008 -51205 7012
rect -52012 6984 -51205 7008
rect -51149 6984 -51027 7042
rect -52012 6734 -51027 6984
rect -45475 8160 -44490 8254
rect -45475 8144 -45141 8160
rect -45475 8086 -45329 8144
rect -45273 8102 -45141 8144
rect -45085 8102 -44490 8160
rect -45273 8086 -44490 8102
rect -45475 8009 -44490 8086
rect -45475 7975 -44878 8009
rect -45475 7967 -45112 7975
rect -45475 7909 -45313 7967
rect -45257 7917 -45112 7967
rect -45056 7951 -44878 7975
rect -44822 7951 -44490 8009
rect -45056 7947 -44490 7951
rect -45056 7917 -44691 7947
rect -45257 7909 -44691 7917
rect -45475 7889 -44691 7909
rect -44635 7889 -44490 7947
rect -45475 7799 -44490 7889
rect -45475 7786 -45095 7799
rect -45475 7728 -45309 7786
rect -45253 7741 -45095 7786
rect -45039 7790 -44490 7799
rect -45039 7741 -44878 7790
rect -45253 7732 -44878 7741
rect -44822 7762 -44490 7790
rect -44822 7732 -44648 7762
rect -45253 7728 -44648 7732
rect -45475 7704 -44648 7728
rect -44592 7704 -44490 7762
rect -45475 7228 -44490 7704
rect -45475 7212 -45170 7228
rect -45475 7154 -45358 7212
rect -45302 7170 -45170 7212
rect -45114 7170 -44490 7228
rect -45302 7154 -44490 7170
rect -45475 7077 -44490 7154
rect -45475 7043 -44907 7077
rect -45475 7035 -45141 7043
rect -45475 6977 -45342 7035
rect -45286 6985 -45141 7035
rect -45085 7019 -44907 7043
rect -44851 7019 -44490 7077
rect -45085 7015 -44490 7019
rect -45085 6985 -44720 7015
rect -45286 6977 -44720 6985
rect -45475 6957 -44720 6977
rect -44664 6957 -44490 7015
rect -45475 6867 -44490 6957
rect -45475 6854 -45124 6867
rect -45475 6796 -45338 6854
rect -45282 6809 -45124 6854
rect -45068 6858 -44490 6867
rect -45068 6809 -44907 6858
rect -45282 6800 -44907 6809
rect -44851 6830 -44490 6858
rect -44851 6800 -44677 6830
rect -45282 6796 -44677 6800
rect -45475 6772 -44677 6796
rect -44621 6772 -44490 6830
rect -59062 6454 -58077 6731
rect -45475 6559 -44490 6772
rect -38757 8090 -37772 8237
rect -38757 8074 -38440 8090
rect -38757 8016 -38628 8074
rect -38572 8032 -38440 8074
rect -38384 8032 -37772 8090
rect -38572 8016 -37772 8032
rect -38757 7939 -37772 8016
rect -38757 7905 -38177 7939
rect -38757 7897 -38411 7905
rect -38757 7839 -38612 7897
rect -38556 7847 -38411 7897
rect -38355 7881 -38177 7905
rect -38121 7881 -37772 7939
rect -38355 7877 -37772 7881
rect -38355 7847 -37990 7877
rect -38556 7839 -37990 7847
rect -38757 7819 -37990 7839
rect -37934 7819 -37772 7877
rect -38757 7729 -37772 7819
rect -38757 7716 -38394 7729
rect -38757 7658 -38608 7716
rect -38552 7671 -38394 7716
rect -38338 7720 -37772 7729
rect -38338 7671 -38177 7720
rect -38552 7662 -38177 7671
rect -38121 7692 -37772 7720
rect -38121 7662 -37947 7692
rect -38552 7658 -37947 7662
rect -38757 7634 -37947 7658
rect -37891 7634 -37772 7692
rect -38757 7251 -37772 7634
rect -38757 7235 -38429 7251
rect -38757 7177 -38617 7235
rect -38561 7193 -38429 7235
rect -38373 7193 -37772 7251
rect -38561 7177 -37772 7193
rect -38757 7100 -37772 7177
rect -38757 7066 -38166 7100
rect -38757 7058 -38400 7066
rect -38757 7000 -38601 7058
rect -38545 7008 -38400 7058
rect -38344 7042 -38166 7066
rect -38110 7042 -37772 7100
rect -38344 7038 -37772 7042
rect -38344 7008 -37979 7038
rect -38545 7000 -37979 7008
rect -38757 6980 -37979 7000
rect -37923 6980 -37772 7038
rect -38757 6890 -37772 6980
rect -38757 6877 -38383 6890
rect -38757 6819 -38597 6877
rect -38541 6832 -38383 6877
rect -38327 6881 -37772 6890
rect -38327 6832 -38166 6881
rect -38541 6823 -38166 6832
rect -38110 6853 -37772 6881
rect -38110 6823 -37936 6853
rect -38541 6819 -37936 6823
rect -38757 6795 -37936 6819
rect -37880 6795 -37772 6853
rect -38757 6542 -37772 6795
rect -31724 8149 -30705 8360
rect -31724 8133 -31413 8149
rect -31724 8075 -31601 8133
rect -31545 8091 -31413 8133
rect -31357 8091 -30705 8149
rect -31545 8075 -30705 8091
rect -31724 7998 -30705 8075
rect -31724 7964 -31150 7998
rect -31724 7956 -31384 7964
rect -31724 7898 -31585 7956
rect -31529 7906 -31384 7956
rect -31328 7940 -31150 7964
rect -31094 7940 -30705 7998
rect -31328 7936 -30705 7940
rect -31328 7906 -30963 7936
rect -31529 7898 -30963 7906
rect -31724 7878 -30963 7898
rect -30907 7878 -30705 7936
rect -31724 7788 -30705 7878
rect -31724 7775 -31367 7788
rect -31724 7717 -31581 7775
rect -31525 7730 -31367 7775
rect -31311 7779 -30705 7788
rect -31311 7730 -31150 7779
rect -31525 7721 -31150 7730
rect -31094 7751 -30705 7779
rect -31094 7721 -30920 7751
rect -31525 7717 -30920 7721
rect -31724 7693 -30920 7717
rect -30864 7693 -30705 7751
rect -31724 7257 -30705 7693
rect -31724 7241 -31396 7257
rect -31724 7183 -31584 7241
rect -31528 7199 -31396 7241
rect -31340 7199 -30705 7257
rect -31528 7183 -30705 7199
rect -31724 7106 -30705 7183
rect -31724 7072 -31133 7106
rect -31724 7064 -31367 7072
rect -31724 7006 -31568 7064
rect -31512 7014 -31367 7064
rect -31311 7048 -31133 7072
rect -31077 7048 -30705 7106
rect -31311 7044 -30705 7048
rect -31311 7014 -30946 7044
rect -31512 7006 -30946 7014
rect -31724 6986 -30946 7006
rect -30890 6986 -30705 7044
rect -31724 6896 -30705 6986
rect -31724 6883 -31350 6896
rect -31724 6825 -31564 6883
rect -31508 6838 -31350 6883
rect -31294 6887 -30705 6896
rect -31294 6838 -31133 6887
rect -31508 6829 -31133 6838
rect -31077 6859 -30705 6887
rect -31077 6829 -30903 6859
rect -31508 6825 -30903 6829
rect -31724 6801 -30903 6825
rect -30847 6801 -30705 6859
rect -31724 6507 -30705 6801
rect -24931 8026 -23912 8238
rect -24931 8010 -24562 8026
rect -24931 7952 -24750 8010
rect -24694 7968 -24562 8010
rect -24506 7968 -23912 8026
rect -24694 7952 -23912 7968
rect -24931 7875 -23912 7952
rect -24931 7841 -24299 7875
rect -24931 7833 -24533 7841
rect -24931 7775 -24734 7833
rect -24678 7783 -24533 7833
rect -24477 7817 -24299 7841
rect -24243 7817 -23912 7875
rect -24477 7813 -23912 7817
rect -24477 7783 -24112 7813
rect -24678 7775 -24112 7783
rect -24931 7755 -24112 7775
rect -24056 7755 -23912 7813
rect -24931 7665 -23912 7755
rect -24931 7652 -24516 7665
rect -24931 7594 -24730 7652
rect -24674 7607 -24516 7652
rect -24460 7656 -23912 7665
rect -24460 7607 -24299 7656
rect -24674 7598 -24299 7607
rect -24243 7628 -23912 7656
rect -24243 7598 -24069 7628
rect -24674 7594 -24069 7598
rect -24931 7570 -24069 7594
rect -24013 7570 -23912 7628
rect -24931 7193 -23912 7570
rect -24931 7177 -24573 7193
rect -24931 7119 -24761 7177
rect -24705 7135 -24573 7177
rect -24517 7135 -23912 7193
rect -24705 7119 -23912 7135
rect -24931 7042 -23912 7119
rect -24931 7008 -24310 7042
rect -24931 7000 -24544 7008
rect -24931 6942 -24745 7000
rect -24689 6950 -24544 7000
rect -24488 6984 -24310 7008
rect -24254 6984 -23912 7042
rect -24488 6980 -23912 6984
rect -24488 6950 -24123 6980
rect -24689 6942 -24123 6950
rect -24931 6922 -24123 6942
rect -24067 6922 -23912 6980
rect -24931 6832 -23912 6922
rect -24931 6819 -24527 6832
rect -24931 6761 -24741 6819
rect -24685 6774 -24527 6819
rect -24471 6823 -23912 6832
rect -24471 6774 -24310 6823
rect -24685 6765 -24310 6774
rect -24254 6795 -23912 6823
rect -24254 6765 -24080 6795
rect -24685 6761 -24080 6765
rect -24931 6737 -24080 6761
rect -24024 6737 -23912 6795
rect -24931 6385 -23912 6737
rect -18061 8108 -17042 8354
rect -18061 8092 -17727 8108
rect -18061 8034 -17915 8092
rect -17859 8050 -17727 8092
rect -17671 8050 -17042 8108
rect -17859 8034 -17042 8050
rect -18061 7957 -17042 8034
rect -18061 7923 -17464 7957
rect -18061 7915 -17698 7923
rect -18061 7857 -17899 7915
rect -17843 7865 -17698 7915
rect -17642 7899 -17464 7923
rect -17408 7899 -17042 7957
rect -17642 7895 -17042 7899
rect -17642 7865 -17277 7895
rect -17843 7857 -17277 7865
rect -18061 7837 -17277 7857
rect -17221 7837 -17042 7895
rect -18061 7747 -17042 7837
rect -18061 7734 -17681 7747
rect -18061 7676 -17895 7734
rect -17839 7689 -17681 7734
rect -17625 7738 -17042 7747
rect -17625 7689 -17464 7738
rect -17839 7680 -17464 7689
rect -17408 7710 -17042 7738
rect -17408 7680 -17234 7710
rect -17839 7676 -17234 7680
rect -18061 7652 -17234 7676
rect -17178 7652 -17042 7710
rect -18061 7251 -17042 7652
rect -18061 7235 -17727 7251
rect -18061 7177 -17915 7235
rect -17859 7193 -17727 7235
rect -17671 7193 -17042 7251
rect -17859 7177 -17042 7193
rect -18061 7100 -17042 7177
rect -18061 7066 -17464 7100
rect -18061 7058 -17698 7066
rect -18061 7000 -17899 7058
rect -17843 7008 -17698 7058
rect -17642 7042 -17464 7066
rect -17408 7042 -17042 7100
rect -17642 7038 -17042 7042
rect -17642 7008 -17277 7038
rect -17843 7000 -17277 7008
rect -18061 6980 -17277 7000
rect -17221 6980 -17042 7038
rect -18061 6890 -17042 6980
rect -18061 6877 -17681 6890
rect -18061 6819 -17895 6877
rect -17839 6832 -17681 6877
rect -17625 6881 -17042 6890
rect -17625 6832 -17464 6881
rect -17839 6823 -17464 6832
rect -17408 6853 -17042 6881
rect -17408 6823 -17234 6853
rect -17839 6819 -17234 6823
rect -18061 6795 -17234 6819
rect -17178 6795 -17042 6853
rect -18061 6501 -17042 6795
rect -11069 8195 -10050 8319
rect -11069 8179 -10735 8195
rect -11069 8121 -10923 8179
rect -10867 8137 -10735 8179
rect -10679 8137 -10050 8195
rect -10867 8121 -10050 8137
rect -11069 8044 -10050 8121
rect -11069 8010 -10472 8044
rect -11069 8002 -10706 8010
rect -11069 7944 -10907 8002
rect -10851 7952 -10706 8002
rect -10650 7986 -10472 8010
rect -10416 7986 -10050 8044
rect -10650 7982 -10050 7986
rect -10650 7952 -10285 7982
rect -10851 7944 -10285 7952
rect -11069 7924 -10285 7944
rect -10229 7924 -10050 7982
rect -11069 7834 -10050 7924
rect -11069 7821 -10689 7834
rect -11069 7763 -10903 7821
rect -10847 7776 -10689 7821
rect -10633 7825 -10050 7834
rect -10633 7776 -10472 7825
rect -10847 7767 -10472 7776
rect -10416 7797 -10050 7825
rect -10416 7767 -10242 7797
rect -10847 7763 -10242 7767
rect -11069 7739 -10242 7763
rect -10186 7739 -10050 7797
rect -11069 7210 -10050 7739
rect -11069 7194 -10712 7210
rect -11069 7136 -10900 7194
rect -10844 7152 -10712 7194
rect -10656 7152 -10050 7210
rect -10844 7136 -10050 7152
rect -11069 7059 -10050 7136
rect -11069 7025 -10449 7059
rect -11069 7017 -10683 7025
rect -11069 6959 -10884 7017
rect -10828 6967 -10683 7017
rect -10627 7001 -10449 7025
rect -10393 7001 -10050 7059
rect -10627 6997 -10050 7001
rect -10627 6967 -10262 6997
rect -10828 6959 -10262 6967
rect -11069 6939 -10262 6959
rect -10206 6939 -10050 6997
rect -11069 6849 -10050 6939
rect -11069 6836 -10666 6849
rect -11069 6778 -10880 6836
rect -10824 6791 -10666 6836
rect -10610 6840 -10050 6849
rect -10610 6791 -10449 6840
rect -10824 6782 -10449 6791
rect -10393 6812 -10050 6840
rect -10393 6782 -10219 6812
rect -10824 6778 -10219 6782
rect -11069 6754 -10219 6778
rect -10163 6754 -10050 6812
rect -11069 6466 -10050 6754
rect -3635 8213 -2616 8337
rect -3635 8197 -3295 8213
rect -3635 8139 -3483 8197
rect -3427 8155 -3295 8197
rect -3239 8155 -2616 8213
rect -3427 8139 -2616 8155
rect -3635 8062 -2616 8139
rect -3635 8028 -3032 8062
rect -3635 8020 -3266 8028
rect -3635 7962 -3467 8020
rect -3411 7970 -3266 8020
rect -3210 8004 -3032 8028
rect -2976 8004 -2616 8062
rect -3210 8000 -2616 8004
rect -3210 7970 -2845 8000
rect -3411 7962 -2845 7970
rect -3635 7942 -2845 7962
rect -2789 7942 -2616 8000
rect -3635 7852 -2616 7942
rect -3635 7839 -3249 7852
rect -3635 7781 -3463 7839
rect -3407 7794 -3249 7839
rect -3193 7843 -2616 7852
rect -3193 7794 -3032 7843
rect -3407 7785 -3032 7794
rect -2976 7815 -2616 7843
rect -2976 7785 -2802 7815
rect -3407 7781 -2802 7785
rect -3635 7757 -2802 7781
rect -2746 7757 -2616 7815
rect -3635 7240 -2616 7757
rect -3635 7224 -3225 7240
rect -3635 7166 -3413 7224
rect -3357 7182 -3225 7224
rect -3169 7182 -2616 7240
rect -3357 7166 -2616 7182
rect -3635 7089 -2616 7166
rect -3635 7055 -2962 7089
rect -3635 7047 -3196 7055
rect -3635 6989 -3397 7047
rect -3341 6997 -3196 7047
rect -3140 7031 -2962 7055
rect -2906 7031 -2616 7089
rect -3140 7027 -2616 7031
rect -3140 6997 -2775 7027
rect -3341 6989 -2775 6997
rect -3635 6969 -2775 6989
rect -2719 6969 -2616 7027
rect -3635 6879 -2616 6969
rect -3635 6866 -3179 6879
rect -3635 6808 -3393 6866
rect -3337 6821 -3179 6866
rect -3123 6870 -2616 6879
rect -3123 6821 -2962 6870
rect -3337 6812 -2962 6821
rect -2906 6842 -2616 6870
rect -2906 6812 -2732 6842
rect -3337 6808 -2732 6812
rect -3635 6784 -2732 6808
rect -2676 6784 -2616 6842
rect -3635 6484 -2616 6784
rect 2058 8166 3077 8290
rect 2058 8150 2415 8166
rect 2058 8092 2227 8150
rect 2283 8108 2415 8150
rect 2471 8108 3077 8166
rect 2283 8092 3077 8108
rect 2058 8015 3077 8092
rect 2058 7981 2678 8015
rect 2058 7973 2444 7981
rect 2058 7915 2243 7973
rect 2299 7923 2444 7973
rect 2500 7957 2678 7981
rect 2734 7957 3077 8015
rect 2500 7953 3077 7957
rect 2500 7923 2865 7953
rect 2299 7915 2865 7923
rect 2058 7895 2865 7915
rect 2921 7895 3077 7953
rect 2058 7805 3077 7895
rect 2058 7792 2461 7805
rect 2058 7734 2247 7792
rect 2303 7747 2461 7792
rect 2517 7796 3077 7805
rect 2517 7747 2678 7796
rect 2303 7738 2678 7747
rect 2734 7768 3077 7796
rect 2734 7738 2908 7768
rect 2303 7734 2908 7738
rect 2058 7710 2908 7734
rect 2964 7710 3077 7768
rect 2058 7141 3077 7710
rect 2058 7125 2444 7141
rect 2058 7067 2256 7125
rect 2312 7083 2444 7125
rect 2500 7083 3077 7141
rect 2312 7067 3077 7083
rect 2058 6990 3077 7067
rect 2058 6956 2707 6990
rect 2058 6948 2473 6956
rect 2058 6890 2272 6948
rect 2328 6898 2473 6948
rect 2529 6932 2707 6956
rect 2763 6932 3077 6990
rect 2529 6928 3077 6932
rect 2529 6898 2894 6928
rect 2328 6890 2894 6898
rect 2058 6870 2894 6890
rect 2950 6870 3077 6928
rect 2058 6780 3077 6870
rect 2058 6767 2490 6780
rect 2058 6709 2276 6767
rect 2332 6722 2490 6767
rect 2546 6771 3077 6780
rect 2546 6722 2707 6771
rect 2332 6713 2707 6722
rect 2763 6743 3077 6771
rect 2763 6713 2937 6743
rect 2332 6709 2937 6713
rect 2058 6685 2937 6709
rect 2993 6685 3077 6743
rect 2058 6437 3077 6685
rect -61751 -68318 -60887 -68247
rect -61751 -68334 -61490 -68318
rect -61751 -68392 -61678 -68334
rect -61622 -68376 -61490 -68334
rect -61434 -68376 -60887 -68318
rect -61622 -68392 -60887 -68376
rect -61751 -68469 -60887 -68392
rect -61751 -68503 -61227 -68469
rect -61751 -68511 -61461 -68503
rect -61751 -68569 -61662 -68511
rect -61606 -68561 -61461 -68511
rect -61405 -68527 -61227 -68503
rect -61171 -68527 -60887 -68469
rect -61405 -68531 -60887 -68527
rect -61405 -68561 -61040 -68531
rect -61606 -68569 -61040 -68561
rect -61751 -68589 -61040 -68569
rect -60984 -68589 -60887 -68531
rect -61751 -68679 -60887 -68589
rect -61751 -68692 -61444 -68679
rect -61751 -68750 -61658 -68692
rect -61602 -68737 -61444 -68692
rect -61388 -68688 -60887 -68679
rect -61388 -68737 -61227 -68688
rect -61602 -68746 -61227 -68737
rect -61171 -68716 -60887 -68688
rect -61171 -68746 -60997 -68716
rect -61602 -68750 -60997 -68746
rect -61751 -68774 -60997 -68750
rect -60941 -68774 -60887 -68716
rect -61751 -68934 -60887 -68774
rect -55242 -68377 -54186 -68282
rect -55242 -68435 -54944 -68377
rect -54888 -68435 -54769 -68377
rect -54713 -68435 -54567 -68377
rect -54511 -68435 -54186 -68377
rect -55242 -68617 -54186 -68435
rect -55242 -68642 -54725 -68617
rect -55242 -68644 -54925 -68642
rect -55242 -68702 -55157 -68644
rect -55101 -68700 -54925 -68644
rect -54869 -68675 -54725 -68642
rect -54669 -68632 -54186 -68617
rect -54669 -68648 -54294 -68632
rect -54669 -68675 -54507 -68648
rect -54869 -68700 -54507 -68675
rect -55101 -68702 -54507 -68700
rect -55242 -68706 -54507 -68702
rect -54451 -68690 -54294 -68648
rect -54238 -68690 -54186 -68632
rect -54451 -68706 -54186 -68690
rect -55242 -68861 -54186 -68706
rect -55242 -68865 -54696 -68861
rect -55242 -68923 -54921 -68865
rect -54865 -68919 -54696 -68865
rect -54640 -68867 -54186 -68861
rect -54640 -68919 -54438 -68867
rect -54865 -68923 -54438 -68919
rect -55242 -68925 -54438 -68923
rect -54382 -68925 -54186 -68867
rect -48439 -68367 -47230 -68311
rect -48439 -68425 -48168 -68367
rect -48112 -68425 -47987 -68367
rect -47931 -68373 -47230 -68367
rect -47931 -68425 -47783 -68373
rect -48439 -68431 -47783 -68425
rect -47727 -68431 -47230 -68373
rect -48439 -68567 -47230 -68431
rect -48439 -68573 -47916 -68567
rect -48439 -68631 -48152 -68573
rect -48096 -68625 -47916 -68573
rect -47860 -68582 -47230 -68567
rect -47860 -68625 -47656 -68582
rect -48096 -68631 -47656 -68625
rect -48439 -68640 -47656 -68631
rect -47600 -68640 -47230 -68582
rect -48439 -68784 -47230 -68640
rect -48439 -68842 -48212 -68784
rect -48156 -68788 -47230 -68784
rect -48156 -68842 -47970 -68788
rect -48439 -68846 -47970 -68842
rect -47914 -68846 -47770 -68788
rect -47714 -68798 -47230 -68788
rect -47714 -68846 -47466 -68798
rect -48439 -68856 -47466 -68846
rect -47410 -68856 -47230 -68798
rect -48439 -68909 -47230 -68856
rect -41649 -68367 -40440 -68326
rect -21096 -68350 -20092 -68263
rect -41649 -68371 -41151 -68367
rect -41649 -68429 -41332 -68371
rect -41276 -68425 -41151 -68371
rect -41095 -68377 -40440 -68367
rect -41095 -68425 -40951 -68377
rect -41276 -68429 -40951 -68425
rect -41649 -68435 -40951 -68429
rect -40895 -68435 -40440 -68377
rect -41649 -68540 -40440 -68435
rect -41649 -68579 -41330 -68540
rect -41649 -68637 -41517 -68579
rect -41461 -68598 -41330 -68579
rect -41274 -68544 -40440 -68540
rect -41274 -68554 -40890 -68544
rect -41274 -68598 -41117 -68554
rect -41461 -68612 -41117 -68598
rect -41061 -68602 -40890 -68554
rect -40834 -68567 -40440 -68544
rect -40834 -68602 -40694 -68567
rect -41061 -68612 -40694 -68602
rect -41461 -68625 -40694 -68612
rect -40638 -68625 -40440 -68567
rect -41461 -68637 -40440 -68625
rect -41649 -68740 -40440 -68637
rect -41649 -68757 -41084 -68740
rect -41649 -68815 -41317 -68757
rect -41261 -68798 -41084 -68757
rect -41028 -68752 -40440 -68740
rect -41028 -68798 -40836 -68752
rect -41261 -68810 -40836 -68798
rect -40780 -68810 -40440 -68752
rect -41261 -68815 -40440 -68810
rect -41649 -68924 -40440 -68815
rect -34904 -68406 -33695 -68353
rect -34904 -68464 -34577 -68406
rect -34521 -68413 -33695 -68406
rect -34521 -68464 -34396 -68413
rect -34904 -68471 -34396 -68464
rect -34340 -68471 -34221 -68413
rect -34165 -68471 -33695 -68413
rect -34904 -68623 -33695 -68471
rect -34904 -68629 -34000 -68623
rect -34904 -68648 -34560 -68629
rect -34904 -68706 -34819 -68648
rect -34763 -68687 -34560 -68648
rect -34504 -68687 -34329 -68629
rect -34273 -68681 -34000 -68629
rect -33944 -68681 -33695 -68623
rect -34273 -68687 -33695 -68681
rect -34763 -68706 -33695 -68687
rect -34904 -68832 -33695 -68706
rect -34904 -68846 -33843 -68832
rect -34904 -68904 -34581 -68846
rect -34525 -68904 -34346 -68846
rect -34290 -68850 -33843 -68846
rect -34290 -68904 -34106 -68850
rect -34904 -68908 -34106 -68904
rect -34050 -68890 -33843 -68850
rect -33787 -68890 -33695 -68832
rect -34050 -68908 -33695 -68890
rect -55242 -68970 -54186 -68925
rect -34904 -68951 -33695 -68908
rect -28030 -68386 -26900 -68350
rect -28030 -68444 -27727 -68386
rect -27671 -68393 -26900 -68386
rect -27671 -68444 -27546 -68393
rect -28030 -68451 -27546 -68444
rect -27490 -68451 -27371 -68393
rect -27315 -68451 -26900 -68393
rect -28030 -68603 -26900 -68451
rect -28030 -68609 -27150 -68603
rect -28030 -68628 -27710 -68609
rect -28030 -68686 -27969 -68628
rect -27913 -68667 -27710 -68628
rect -27654 -68667 -27479 -68609
rect -27423 -68661 -27150 -68609
rect -27094 -68661 -26900 -68603
rect -27423 -68667 -26900 -68661
rect -27913 -68686 -26900 -68667
rect -28030 -68812 -26900 -68686
rect -28030 -68826 -26993 -68812
rect -28030 -68884 -27731 -68826
rect -27675 -68884 -27496 -68826
rect -27440 -68830 -26993 -68826
rect -27440 -68884 -27256 -68830
rect -28030 -68888 -27256 -68884
rect -27200 -68870 -26993 -68830
rect -26937 -68870 -26900 -68812
rect -27200 -68888 -26900 -68870
rect -28030 -68930 -26900 -68888
rect -21096 -68386 -19960 -68350
rect -21096 -68444 -20787 -68386
rect -20731 -68393 -19960 -68386
rect -20731 -68444 -20606 -68393
rect -21096 -68451 -20606 -68444
rect -20550 -68451 -20431 -68393
rect -20375 -68451 -19960 -68393
rect -21096 -68603 -19960 -68451
rect -21096 -68609 -20210 -68603
rect -21096 -68628 -20770 -68609
rect -21096 -68686 -21029 -68628
rect -20973 -68667 -20770 -68628
rect -20714 -68667 -20539 -68609
rect -20483 -68661 -20210 -68609
rect -20154 -68661 -19960 -68603
rect -20483 -68667 -19960 -68661
rect -20973 -68686 -19960 -68667
rect -21096 -68812 -19960 -68686
rect -21096 -68826 -20053 -68812
rect -21096 -68884 -20791 -68826
rect -20735 -68884 -20556 -68826
rect -20500 -68830 -20053 -68826
rect -20500 -68884 -20316 -68830
rect -21096 -68888 -20316 -68884
rect -20260 -68870 -20053 -68830
rect -19997 -68870 -19960 -68812
rect -20260 -68888 -19960 -68870
rect -21096 -68930 -19960 -68888
rect -14409 -68379 -13405 -68255
rect -14409 -68437 -14124 -68379
rect -14068 -68384 -13405 -68379
rect -14068 -68437 -13945 -68384
rect -14409 -68442 -13945 -68437
rect -13889 -68442 -13762 -68384
rect -13706 -68442 -13405 -68384
rect -14409 -68632 -13405 -68442
rect -14409 -68636 -13637 -68632
rect -14409 -68642 -13845 -68636
rect -14409 -68648 -14037 -68642
rect -14409 -68706 -14262 -68648
rect -14206 -68700 -14037 -68648
rect -13981 -68694 -13845 -68642
rect -13789 -68690 -13637 -68636
rect -13581 -68690 -13405 -68632
rect -13789 -68694 -13405 -68690
rect -13981 -68700 -13405 -68694
rect -14206 -68706 -13405 -68700
rect -14409 -68846 -13405 -68706
rect -14409 -68904 -14199 -68846
rect -14143 -68904 -13980 -68846
rect -13924 -68904 -13791 -68846
rect -13735 -68904 -13543 -68846
rect -13487 -68904 -13405 -68846
rect -21096 -68951 -20092 -68930
rect -14409 -68943 -13405 -68904
rect -7481 -68359 -6477 -68255
rect -7481 -68417 -7286 -68359
rect -7230 -68417 -7111 -68359
rect -7055 -68417 -6921 -68359
rect -6865 -68417 -6477 -68359
rect -7481 -68609 -6477 -68417
rect -7481 -68615 -6648 -68609
rect -7481 -68621 -6909 -68615
rect -7481 -68627 -7129 -68621
rect -7481 -68685 -7402 -68627
rect -7346 -68679 -7129 -68627
rect -7073 -68673 -6909 -68621
rect -6853 -68667 -6648 -68615
rect -6592 -68667 -6477 -68609
rect -6853 -68673 -6477 -68667
rect -7073 -68679 -6477 -68673
rect -7346 -68685 -6477 -68679
rect -7481 -68844 -6477 -68685
rect -7481 -68850 -6723 -68844
rect -7481 -68852 -7152 -68850
rect -7481 -68910 -7367 -68852
rect -7311 -68908 -7152 -68852
rect -7096 -68908 -6934 -68850
rect -6878 -68902 -6723 -68850
rect -6667 -68902 -6477 -68844
rect -6878 -68908 -6477 -68902
rect -7311 -68910 -6477 -68908
rect -7481 -68943 -6477 -68910
rect -676 -68356 328 -68259
rect -676 -68359 -70 -68356
rect -676 -68417 -476 -68359
rect -420 -68363 -70 -68359
rect -420 -68417 -283 -68363
rect -676 -68421 -283 -68417
rect -227 -68414 -70 -68363
rect -14 -68414 328 -68356
rect -227 -68421 328 -68414
rect -676 -68592 328 -68421
rect -676 -68596 145 -68592
rect -676 -68600 -345 -68596
rect -676 -68658 -595 -68600
rect -539 -68654 -345 -68600
rect -289 -68654 -112 -68596
rect -56 -68650 145 -68596
rect 201 -68650 328 -68592
rect -56 -68654 328 -68650
rect -539 -68658 328 -68654
rect -676 -68846 328 -68658
rect -676 -68850 -308 -68846
rect -676 -68908 -566 -68850
rect -510 -68904 -308 -68850
rect -252 -68850 328 -68846
rect -252 -68904 -70 -68850
rect -510 -68908 -70 -68904
rect -14 -68857 328 -68850
rect -14 -68908 184 -68857
rect -676 -68915 184 -68908
rect 240 -68915 328 -68857
rect -676 -68947 328 -68915
rect 5835 -68350 6839 -68257
rect 5835 -68408 6318 -68350
rect 6374 -68408 6506 -68350
rect 6562 -68356 6839 -68350
rect 6562 -68408 6708 -68356
rect 5835 -68414 6708 -68408
rect 6764 -68414 6839 -68356
rect 5835 -68571 6839 -68414
rect 5835 -68629 6143 -68571
rect 6199 -68575 6606 -68571
rect 6199 -68629 6395 -68575
rect 5835 -68633 6395 -68629
rect 6451 -68629 6606 -68575
rect 6662 -68629 6839 -68571
rect 6451 -68633 6839 -68629
rect 5835 -68686 6839 -68633
rect 5835 -68744 5931 -68686
rect 5987 -68744 6839 -68686
rect 5835 -68850 6839 -68744
rect 5835 -68852 6327 -68850
rect 5835 -68910 6139 -68852
rect 6195 -68908 6327 -68852
rect 6383 -68908 6533 -68850
rect 6589 -68852 6839 -68850
rect 6589 -68908 6737 -68852
rect 6195 -68910 6737 -68908
rect 6793 -68910 6839 -68852
rect 5835 -68945 6839 -68910
<< via4 >>
rect -51678 8304 -51622 8306
rect -51866 8288 -51810 8290
rect -51866 8234 -51810 8288
rect -51678 8250 -51622 8304
rect -64935 7983 -64879 7985
rect -65123 7967 -65067 7969
rect -65123 7913 -65067 7967
rect -64935 7929 -64879 7983
rect -64672 7832 -64616 7834
rect -64906 7798 -64850 7800
rect -65107 7790 -65051 7792
rect -65107 7736 -65051 7790
rect -64906 7744 -64850 7798
rect -64672 7778 -64616 7832
rect -64485 7770 -64429 7772
rect -64485 7716 -64429 7770
rect -64889 7622 -64833 7624
rect -65103 7609 -65047 7611
rect -65103 7555 -65047 7609
rect -64889 7568 -64833 7622
rect -64672 7613 -64616 7615
rect -64672 7559 -64616 7613
rect -64442 7585 -64386 7587
rect -64442 7531 -64386 7585
rect -64958 7165 -64902 7167
rect -65146 7149 -65090 7151
rect -65146 7095 -65090 7149
rect -64958 7111 -64902 7165
rect -64695 7014 -64639 7016
rect -64929 6980 -64873 6982
rect -65130 6972 -65074 6974
rect -65130 6918 -65074 6972
rect -64929 6926 -64873 6980
rect -64695 6960 -64639 7014
rect -64508 6952 -64452 6954
rect -64508 6898 -64452 6952
rect -64912 6804 -64856 6806
rect -65126 6791 -65070 6793
rect -65126 6737 -65070 6791
rect -64912 6750 -64856 6804
rect -64695 6795 -64639 6797
rect -64695 6741 -64639 6795
rect -64465 6767 -64409 6769
rect -64465 6713 -64409 6767
rect -58740 8065 -58684 8067
rect -58928 8049 -58872 8051
rect -58928 7995 -58872 8049
rect -58740 8011 -58684 8065
rect -58477 7914 -58421 7916
rect -58711 7880 -58655 7882
rect -58912 7872 -58856 7874
rect -58912 7818 -58856 7872
rect -58711 7826 -58655 7880
rect -58477 7860 -58421 7914
rect -58290 7852 -58234 7854
rect -58290 7798 -58234 7852
rect -58694 7704 -58638 7706
rect -58908 7691 -58852 7693
rect -58908 7637 -58852 7691
rect -58694 7650 -58638 7704
rect -58477 7695 -58421 7697
rect -58477 7641 -58421 7695
rect -58247 7667 -58191 7669
rect -58247 7613 -58191 7667
rect -58740 7185 -58684 7187
rect -58928 7169 -58872 7171
rect -58928 7115 -58872 7169
rect -58740 7131 -58684 7185
rect -58477 7034 -58421 7036
rect -58711 7000 -58655 7002
rect -58912 6992 -58856 6994
rect -58912 6938 -58856 6992
rect -58711 6946 -58655 7000
rect -58477 6980 -58421 7034
rect -58290 6972 -58234 6974
rect -58290 6918 -58234 6972
rect -58694 6824 -58638 6826
rect -58908 6811 -58852 6813
rect -58908 6757 -58852 6811
rect -58694 6770 -58638 6824
rect -58477 6815 -58421 6817
rect -58477 6761 -58421 6815
rect -58247 6787 -58191 6789
rect -58247 6733 -58191 6787
rect -51415 8153 -51359 8155
rect -51649 8119 -51593 8121
rect -51850 8111 -51794 8113
rect -51850 8057 -51794 8111
rect -51649 8065 -51593 8119
rect -51415 8099 -51359 8153
rect -51228 8091 -51172 8093
rect -51228 8037 -51172 8091
rect -51632 7943 -51576 7945
rect -51846 7930 -51790 7932
rect -51846 7876 -51790 7930
rect -51632 7889 -51576 7943
rect -51415 7934 -51359 7936
rect -51415 7880 -51359 7934
rect -51185 7906 -51129 7908
rect -51185 7852 -51129 7906
rect -51698 7438 -51642 7440
rect -51886 7422 -51830 7424
rect -51886 7368 -51830 7422
rect -51698 7384 -51642 7438
rect -51435 7287 -51379 7289
rect -51669 7253 -51613 7255
rect -51870 7245 -51814 7247
rect -51870 7191 -51814 7245
rect -51669 7199 -51613 7253
rect -51435 7233 -51379 7287
rect -51248 7225 -51192 7227
rect -51248 7171 -51192 7225
rect -51652 7077 -51596 7079
rect -51866 7064 -51810 7066
rect -51866 7010 -51810 7064
rect -51652 7023 -51596 7077
rect -51435 7068 -51379 7070
rect -51435 7014 -51379 7068
rect -51205 7040 -51149 7042
rect -51205 6986 -51149 7040
rect -45141 8158 -45085 8160
rect -45329 8142 -45273 8144
rect -45329 8088 -45273 8142
rect -45141 8104 -45085 8158
rect -44878 8007 -44822 8009
rect -45112 7973 -45056 7975
rect -45313 7965 -45257 7967
rect -45313 7911 -45257 7965
rect -45112 7919 -45056 7973
rect -44878 7953 -44822 8007
rect -44691 7945 -44635 7947
rect -44691 7891 -44635 7945
rect -45095 7797 -45039 7799
rect -45309 7784 -45253 7786
rect -45309 7730 -45253 7784
rect -45095 7743 -45039 7797
rect -44878 7788 -44822 7790
rect -44878 7734 -44822 7788
rect -44648 7760 -44592 7762
rect -44648 7706 -44592 7760
rect -45170 7226 -45114 7228
rect -45358 7210 -45302 7212
rect -45358 7156 -45302 7210
rect -45170 7172 -45114 7226
rect -44907 7075 -44851 7077
rect -45141 7041 -45085 7043
rect -45342 7033 -45286 7035
rect -45342 6979 -45286 7033
rect -45141 6987 -45085 7041
rect -44907 7021 -44851 7075
rect -44720 7013 -44664 7015
rect -44720 6959 -44664 7013
rect -45124 6865 -45068 6867
rect -45338 6852 -45282 6854
rect -45338 6798 -45282 6852
rect -45124 6811 -45068 6865
rect -44907 6856 -44851 6858
rect -44907 6802 -44851 6856
rect -44677 6828 -44621 6830
rect -44677 6774 -44621 6828
rect -38440 8088 -38384 8090
rect -38628 8072 -38572 8074
rect -38628 8018 -38572 8072
rect -38440 8034 -38384 8088
rect -38177 7937 -38121 7939
rect -38411 7903 -38355 7905
rect -38612 7895 -38556 7897
rect -38612 7841 -38556 7895
rect -38411 7849 -38355 7903
rect -38177 7883 -38121 7937
rect -37990 7875 -37934 7877
rect -37990 7821 -37934 7875
rect -38394 7727 -38338 7729
rect -38608 7714 -38552 7716
rect -38608 7660 -38552 7714
rect -38394 7673 -38338 7727
rect -38177 7718 -38121 7720
rect -38177 7664 -38121 7718
rect -37947 7690 -37891 7692
rect -37947 7636 -37891 7690
rect -38429 7249 -38373 7251
rect -38617 7233 -38561 7235
rect -38617 7179 -38561 7233
rect -38429 7195 -38373 7249
rect -38166 7098 -38110 7100
rect -38400 7064 -38344 7066
rect -38601 7056 -38545 7058
rect -38601 7002 -38545 7056
rect -38400 7010 -38344 7064
rect -38166 7044 -38110 7098
rect -37979 7036 -37923 7038
rect -37979 6982 -37923 7036
rect -38383 6888 -38327 6890
rect -38597 6875 -38541 6877
rect -38597 6821 -38541 6875
rect -38383 6834 -38327 6888
rect -38166 6879 -38110 6881
rect -38166 6825 -38110 6879
rect -37936 6851 -37880 6853
rect -37936 6797 -37880 6851
rect -31413 8147 -31357 8149
rect -31601 8131 -31545 8133
rect -31601 8077 -31545 8131
rect -31413 8093 -31357 8147
rect -31150 7996 -31094 7998
rect -31384 7962 -31328 7964
rect -31585 7954 -31529 7956
rect -31585 7900 -31529 7954
rect -31384 7908 -31328 7962
rect -31150 7942 -31094 7996
rect -30963 7934 -30907 7936
rect -30963 7880 -30907 7934
rect -31367 7786 -31311 7788
rect -31581 7773 -31525 7775
rect -31581 7719 -31525 7773
rect -31367 7732 -31311 7786
rect -31150 7777 -31094 7779
rect -31150 7723 -31094 7777
rect -30920 7749 -30864 7751
rect -30920 7695 -30864 7749
rect -31396 7255 -31340 7257
rect -31584 7239 -31528 7241
rect -31584 7185 -31528 7239
rect -31396 7201 -31340 7255
rect -31133 7104 -31077 7106
rect -31367 7070 -31311 7072
rect -31568 7062 -31512 7064
rect -31568 7008 -31512 7062
rect -31367 7016 -31311 7070
rect -31133 7050 -31077 7104
rect -30946 7042 -30890 7044
rect -30946 6988 -30890 7042
rect -31350 6894 -31294 6896
rect -31564 6881 -31508 6883
rect -31564 6827 -31508 6881
rect -31350 6840 -31294 6894
rect -31133 6885 -31077 6887
rect -31133 6831 -31077 6885
rect -30903 6857 -30847 6859
rect -30903 6803 -30847 6857
rect -24562 8024 -24506 8026
rect -24750 8008 -24694 8010
rect -24750 7954 -24694 8008
rect -24562 7970 -24506 8024
rect -24299 7873 -24243 7875
rect -24533 7839 -24477 7841
rect -24734 7831 -24678 7833
rect -24734 7777 -24678 7831
rect -24533 7785 -24477 7839
rect -24299 7819 -24243 7873
rect -24112 7811 -24056 7813
rect -24112 7757 -24056 7811
rect -24516 7663 -24460 7665
rect -24730 7650 -24674 7652
rect -24730 7596 -24674 7650
rect -24516 7609 -24460 7663
rect -24299 7654 -24243 7656
rect -24299 7600 -24243 7654
rect -24069 7626 -24013 7628
rect -24069 7572 -24013 7626
rect -24573 7191 -24517 7193
rect -24761 7175 -24705 7177
rect -24761 7121 -24705 7175
rect -24573 7137 -24517 7191
rect -24310 7040 -24254 7042
rect -24544 7006 -24488 7008
rect -24745 6998 -24689 7000
rect -24745 6944 -24689 6998
rect -24544 6952 -24488 7006
rect -24310 6986 -24254 7040
rect -24123 6978 -24067 6980
rect -24123 6924 -24067 6978
rect -24527 6830 -24471 6832
rect -24741 6817 -24685 6819
rect -24741 6763 -24685 6817
rect -24527 6776 -24471 6830
rect -24310 6821 -24254 6823
rect -24310 6767 -24254 6821
rect -24080 6793 -24024 6795
rect -24080 6739 -24024 6793
rect -17727 8106 -17671 8108
rect -17915 8090 -17859 8092
rect -17915 8036 -17859 8090
rect -17727 8052 -17671 8106
rect -17464 7955 -17408 7957
rect -17698 7921 -17642 7923
rect -17899 7913 -17843 7915
rect -17899 7859 -17843 7913
rect -17698 7867 -17642 7921
rect -17464 7901 -17408 7955
rect -17277 7893 -17221 7895
rect -17277 7839 -17221 7893
rect -17681 7745 -17625 7747
rect -17895 7732 -17839 7734
rect -17895 7678 -17839 7732
rect -17681 7691 -17625 7745
rect -17464 7736 -17408 7738
rect -17464 7682 -17408 7736
rect -17234 7708 -17178 7710
rect -17234 7654 -17178 7708
rect -17727 7249 -17671 7251
rect -17915 7233 -17859 7235
rect -17915 7179 -17859 7233
rect -17727 7195 -17671 7249
rect -17464 7098 -17408 7100
rect -17698 7064 -17642 7066
rect -17899 7056 -17843 7058
rect -17899 7002 -17843 7056
rect -17698 7010 -17642 7064
rect -17464 7044 -17408 7098
rect -17277 7036 -17221 7038
rect -17277 6982 -17221 7036
rect -17681 6888 -17625 6890
rect -17895 6875 -17839 6877
rect -17895 6821 -17839 6875
rect -17681 6834 -17625 6888
rect -17464 6879 -17408 6881
rect -17464 6825 -17408 6879
rect -17234 6851 -17178 6853
rect -17234 6797 -17178 6851
rect -10735 8193 -10679 8195
rect -10923 8177 -10867 8179
rect -10923 8123 -10867 8177
rect -10735 8139 -10679 8193
rect -10472 8042 -10416 8044
rect -10706 8008 -10650 8010
rect -10907 8000 -10851 8002
rect -10907 7946 -10851 8000
rect -10706 7954 -10650 8008
rect -10472 7988 -10416 8042
rect -10285 7980 -10229 7982
rect -10285 7926 -10229 7980
rect -10689 7832 -10633 7834
rect -10903 7819 -10847 7821
rect -10903 7765 -10847 7819
rect -10689 7778 -10633 7832
rect -10472 7823 -10416 7825
rect -10472 7769 -10416 7823
rect -10242 7795 -10186 7797
rect -10242 7741 -10186 7795
rect -10712 7208 -10656 7210
rect -10900 7192 -10844 7194
rect -10900 7138 -10844 7192
rect -10712 7154 -10656 7208
rect -10449 7057 -10393 7059
rect -10683 7023 -10627 7025
rect -10884 7015 -10828 7017
rect -10884 6961 -10828 7015
rect -10683 6969 -10627 7023
rect -10449 7003 -10393 7057
rect -10262 6995 -10206 6997
rect -10262 6941 -10206 6995
rect -10666 6847 -10610 6849
rect -10880 6834 -10824 6836
rect -10880 6780 -10824 6834
rect -10666 6793 -10610 6847
rect -10449 6838 -10393 6840
rect -10449 6784 -10393 6838
rect -10219 6810 -10163 6812
rect -10219 6756 -10163 6810
rect -3295 8211 -3239 8213
rect -3483 8195 -3427 8197
rect -3483 8141 -3427 8195
rect -3295 8157 -3239 8211
rect -3032 8060 -2976 8062
rect -3266 8026 -3210 8028
rect -3467 8018 -3411 8020
rect -3467 7964 -3411 8018
rect -3266 7972 -3210 8026
rect -3032 8006 -2976 8060
rect -2845 7998 -2789 8000
rect -2845 7944 -2789 7998
rect -3249 7850 -3193 7852
rect -3463 7837 -3407 7839
rect -3463 7783 -3407 7837
rect -3249 7796 -3193 7850
rect -3032 7841 -2976 7843
rect -3032 7787 -2976 7841
rect -2802 7813 -2746 7815
rect -2802 7759 -2746 7813
rect -3225 7238 -3169 7240
rect -3413 7222 -3357 7224
rect -3413 7168 -3357 7222
rect -3225 7184 -3169 7238
rect -2962 7087 -2906 7089
rect -3196 7053 -3140 7055
rect -3397 7045 -3341 7047
rect -3397 6991 -3341 7045
rect -3196 6999 -3140 7053
rect -2962 7033 -2906 7087
rect -2775 7025 -2719 7027
rect -2775 6971 -2719 7025
rect -3179 6877 -3123 6879
rect -3393 6864 -3337 6866
rect -3393 6810 -3337 6864
rect -3179 6823 -3123 6877
rect -2962 6868 -2906 6870
rect -2962 6814 -2906 6868
rect -2732 6840 -2676 6842
rect -2732 6786 -2676 6840
rect 2415 8164 2471 8166
rect 2227 8148 2283 8150
rect 2227 8094 2283 8148
rect 2415 8110 2471 8164
rect 2678 8013 2734 8015
rect 2444 7979 2500 7981
rect 2243 7971 2299 7973
rect 2243 7917 2299 7971
rect 2444 7925 2500 7979
rect 2678 7959 2734 8013
rect 2865 7951 2921 7953
rect 2865 7897 2921 7951
rect 2461 7803 2517 7805
rect 2247 7790 2303 7792
rect 2247 7736 2303 7790
rect 2461 7749 2517 7803
rect 2678 7794 2734 7796
rect 2678 7740 2734 7794
rect 2908 7766 2964 7768
rect 2908 7712 2964 7766
rect 2444 7139 2500 7141
rect 2256 7123 2312 7125
rect 2256 7069 2312 7123
rect 2444 7085 2500 7139
rect 2707 6988 2763 6990
rect 2473 6954 2529 6956
rect 2272 6946 2328 6948
rect 2272 6892 2328 6946
rect 2473 6900 2529 6954
rect 2707 6934 2763 6988
rect 2894 6926 2950 6928
rect 2894 6872 2950 6926
rect 2490 6778 2546 6780
rect 2276 6765 2332 6767
rect 2276 6711 2332 6765
rect 2490 6724 2546 6778
rect 2707 6769 2763 6771
rect 2707 6715 2763 6769
rect 2937 6741 2993 6743
rect 2937 6687 2993 6741
rect -61490 -68320 -61434 -68318
rect -61678 -68336 -61622 -68334
rect -61678 -68390 -61622 -68336
rect -61490 -68374 -61434 -68320
rect -61227 -68471 -61171 -68469
rect -61461 -68505 -61405 -68503
rect -61662 -68513 -61606 -68511
rect -61662 -68567 -61606 -68513
rect -61461 -68559 -61405 -68505
rect -61227 -68525 -61171 -68471
rect -61040 -68533 -60984 -68531
rect -61040 -68587 -60984 -68533
rect -61444 -68681 -61388 -68679
rect -61658 -68694 -61602 -68692
rect -61658 -68748 -61602 -68694
rect -61444 -68735 -61388 -68681
rect -61227 -68690 -61171 -68688
rect -61227 -68744 -61171 -68690
rect -60997 -68718 -60941 -68716
rect -60997 -68772 -60941 -68718
rect -54944 -68379 -54888 -68377
rect -54944 -68433 -54888 -68379
rect -54769 -68379 -54713 -68377
rect -54769 -68433 -54713 -68379
rect -54567 -68379 -54511 -68377
rect -54567 -68433 -54511 -68379
rect -54725 -68619 -54669 -68617
rect -54925 -68644 -54869 -68642
rect -55157 -68646 -55101 -68644
rect -55157 -68700 -55101 -68646
rect -54925 -68698 -54869 -68644
rect -54725 -68673 -54669 -68619
rect -54294 -68634 -54238 -68632
rect -54507 -68650 -54451 -68648
rect -54507 -68704 -54451 -68650
rect -54294 -68688 -54238 -68634
rect -54696 -68863 -54640 -68861
rect -54921 -68867 -54865 -68865
rect -54921 -68921 -54865 -68867
rect -54696 -68917 -54640 -68863
rect -54438 -68869 -54382 -68867
rect -54438 -68923 -54382 -68869
rect -48168 -68369 -48112 -68367
rect -48168 -68423 -48112 -68369
rect -47987 -68369 -47931 -68367
rect -47987 -68423 -47931 -68369
rect -47783 -68375 -47727 -68373
rect -47783 -68429 -47727 -68375
rect -47916 -68569 -47860 -68567
rect -48152 -68575 -48096 -68573
rect -48152 -68629 -48096 -68575
rect -47916 -68623 -47860 -68569
rect -47656 -68584 -47600 -68582
rect -47656 -68638 -47600 -68584
rect -48212 -68786 -48156 -68784
rect -48212 -68840 -48156 -68786
rect -47970 -68790 -47914 -68788
rect -47970 -68844 -47914 -68790
rect -47770 -68790 -47714 -68788
rect -47770 -68844 -47714 -68790
rect -47466 -68800 -47410 -68798
rect -47466 -68854 -47410 -68800
rect -41151 -68369 -41095 -68367
rect -41332 -68373 -41276 -68371
rect -41332 -68427 -41276 -68373
rect -41151 -68423 -41095 -68369
rect -40951 -68379 -40895 -68377
rect -40951 -68433 -40895 -68379
rect -41330 -68542 -41274 -68540
rect -41517 -68581 -41461 -68579
rect -41517 -68635 -41461 -68581
rect -41330 -68596 -41274 -68542
rect -40890 -68546 -40834 -68544
rect -41117 -68556 -41061 -68554
rect -41117 -68610 -41061 -68556
rect -40890 -68600 -40834 -68546
rect -40694 -68569 -40638 -68567
rect -40694 -68623 -40638 -68569
rect -41084 -68742 -41028 -68740
rect -41317 -68759 -41261 -68757
rect -41317 -68813 -41261 -68759
rect -41084 -68796 -41028 -68742
rect -40836 -68754 -40780 -68752
rect -40836 -68808 -40780 -68754
rect -34577 -68408 -34521 -68406
rect -34577 -68462 -34521 -68408
rect -34396 -68415 -34340 -68413
rect -34396 -68469 -34340 -68415
rect -34221 -68415 -34165 -68413
rect -34221 -68469 -34165 -68415
rect -34000 -68625 -33944 -68623
rect -34560 -68631 -34504 -68629
rect -34819 -68650 -34763 -68648
rect -34819 -68704 -34763 -68650
rect -34560 -68685 -34504 -68631
rect -34329 -68631 -34273 -68629
rect -34329 -68685 -34273 -68631
rect -34000 -68679 -33944 -68625
rect -33843 -68834 -33787 -68832
rect -34581 -68848 -34525 -68846
rect -34581 -68902 -34525 -68848
rect -34346 -68848 -34290 -68846
rect -34346 -68902 -34290 -68848
rect -34106 -68852 -34050 -68850
rect -34106 -68906 -34050 -68852
rect -33843 -68888 -33787 -68834
rect -27727 -68388 -27671 -68386
rect -27727 -68442 -27671 -68388
rect -27546 -68395 -27490 -68393
rect -27546 -68449 -27490 -68395
rect -27371 -68395 -27315 -68393
rect -27371 -68449 -27315 -68395
rect -27150 -68605 -27094 -68603
rect -27710 -68611 -27654 -68609
rect -27969 -68630 -27913 -68628
rect -27969 -68684 -27913 -68630
rect -27710 -68665 -27654 -68611
rect -27479 -68611 -27423 -68609
rect -27479 -68665 -27423 -68611
rect -27150 -68659 -27094 -68605
rect -26993 -68814 -26937 -68812
rect -27731 -68828 -27675 -68826
rect -27731 -68882 -27675 -68828
rect -27496 -68828 -27440 -68826
rect -27496 -68882 -27440 -68828
rect -27256 -68832 -27200 -68830
rect -27256 -68886 -27200 -68832
rect -26993 -68868 -26937 -68814
rect -20787 -68388 -20731 -68386
rect -20787 -68442 -20731 -68388
rect -20606 -68395 -20550 -68393
rect -20606 -68449 -20550 -68395
rect -20431 -68395 -20375 -68393
rect -20431 -68449 -20375 -68395
rect -20210 -68605 -20154 -68603
rect -20770 -68611 -20714 -68609
rect -21029 -68630 -20973 -68628
rect -21029 -68684 -20973 -68630
rect -20770 -68665 -20714 -68611
rect -20539 -68611 -20483 -68609
rect -20539 -68665 -20483 -68611
rect -20210 -68659 -20154 -68605
rect -20053 -68814 -19997 -68812
rect -20791 -68828 -20735 -68826
rect -20791 -68882 -20735 -68828
rect -20556 -68828 -20500 -68826
rect -20556 -68882 -20500 -68828
rect -20316 -68832 -20260 -68830
rect -20316 -68886 -20260 -68832
rect -20053 -68868 -19997 -68814
rect -14124 -68381 -14068 -68379
rect -14124 -68435 -14068 -68381
rect -13945 -68386 -13889 -68384
rect -13945 -68440 -13889 -68386
rect -13762 -68386 -13706 -68384
rect -13762 -68440 -13706 -68386
rect -13637 -68634 -13581 -68632
rect -13845 -68638 -13789 -68636
rect -14037 -68644 -13981 -68642
rect -14262 -68650 -14206 -68648
rect -14262 -68704 -14206 -68650
rect -14037 -68698 -13981 -68644
rect -13845 -68692 -13789 -68638
rect -13637 -68688 -13581 -68634
rect -14199 -68848 -14143 -68846
rect -14199 -68902 -14143 -68848
rect -13980 -68848 -13924 -68846
rect -13980 -68902 -13924 -68848
rect -13791 -68848 -13735 -68846
rect -13791 -68902 -13735 -68848
rect -13543 -68848 -13487 -68846
rect -13543 -68902 -13487 -68848
rect -7286 -68361 -7230 -68359
rect -7286 -68415 -7230 -68361
rect -7111 -68361 -7055 -68359
rect -7111 -68415 -7055 -68361
rect -6921 -68361 -6865 -68359
rect -6921 -68415 -6865 -68361
rect -6648 -68611 -6592 -68609
rect -6909 -68617 -6853 -68615
rect -7129 -68623 -7073 -68621
rect -7402 -68629 -7346 -68627
rect -7402 -68683 -7346 -68629
rect -7129 -68677 -7073 -68623
rect -6909 -68671 -6853 -68617
rect -6648 -68665 -6592 -68611
rect -6723 -68846 -6667 -68844
rect -7152 -68852 -7096 -68850
rect -7367 -68854 -7311 -68852
rect -7367 -68908 -7311 -68854
rect -7152 -68906 -7096 -68852
rect -6934 -68852 -6878 -68850
rect -6934 -68906 -6878 -68852
rect -6723 -68900 -6667 -68846
rect -70 -68358 -14 -68356
rect -476 -68361 -420 -68359
rect -476 -68415 -420 -68361
rect -283 -68365 -227 -68363
rect -283 -68419 -227 -68365
rect -70 -68412 -14 -68358
rect 145 -68594 201 -68592
rect -345 -68598 -289 -68596
rect -595 -68602 -539 -68600
rect -595 -68656 -539 -68602
rect -345 -68652 -289 -68598
rect -112 -68598 -56 -68596
rect -112 -68652 -56 -68598
rect 145 -68648 201 -68594
rect -308 -68848 -252 -68846
rect -566 -68852 -510 -68850
rect -566 -68906 -510 -68852
rect -308 -68902 -252 -68848
rect -70 -68852 -14 -68850
rect -70 -68906 -14 -68852
rect 184 -68859 240 -68857
rect 184 -68913 240 -68859
rect 6318 -68352 6374 -68350
rect 6318 -68406 6374 -68352
rect 6506 -68352 6562 -68350
rect 6506 -68406 6562 -68352
rect 6708 -68358 6764 -68356
rect 6708 -68412 6764 -68358
rect 6143 -68573 6199 -68571
rect 6143 -68627 6199 -68573
rect 6606 -68573 6662 -68571
rect 6395 -68577 6451 -68575
rect 6395 -68631 6451 -68577
rect 6606 -68627 6662 -68573
rect 5931 -68688 5987 -68686
rect 5931 -68742 5987 -68688
rect 6327 -68852 6383 -68850
rect 6139 -68854 6195 -68852
rect 6139 -68908 6195 -68854
rect 6327 -68906 6383 -68852
rect 6533 -68852 6589 -68850
rect 6533 -68906 6589 -68852
rect 6737 -68854 6793 -68852
rect 6737 -68908 6793 -68854
<< metal5 >>
rect -52012 8390 -51027 8429
rect -65240 8306 3710 8390
rect -65240 8290 -51678 8306
rect -65240 8234 -51866 8290
rect -51810 8250 -51678 8290
rect -51622 8250 3710 8306
rect -51810 8234 3710 8250
rect -65240 8213 3710 8234
rect -65240 8197 -3295 8213
rect -65240 8195 -3483 8197
rect -65240 8179 -10735 8195
rect -65240 8160 -10923 8179
rect -65240 8155 -45141 8160
rect -65240 8149 -51415 8155
rect -65244 8121 -51415 8149
rect -65244 8113 -51649 8121
rect -65244 8067 -51850 8113
rect -65244 8051 -58740 8067
rect -65244 7995 -58928 8051
rect -58872 8011 -58740 8051
rect -58684 8057 -51850 8067
rect -51794 8065 -51649 8113
rect -51593 8099 -51415 8121
rect -51359 8144 -45141 8155
rect -51359 8099 -45329 8144
rect -51593 8093 -45329 8099
rect -51593 8065 -51228 8093
rect -51794 8057 -51228 8065
rect -58684 8037 -51228 8057
rect -51172 8088 -45329 8093
rect -45273 8104 -45141 8144
rect -45085 8149 -10923 8160
rect -45085 8133 -31413 8149
rect -45085 8104 -31601 8133
rect -45273 8090 -31601 8104
rect -45273 8088 -38440 8090
rect -51172 8074 -38440 8088
rect -51172 8037 -38628 8074
rect -58684 8018 -38628 8037
rect -38572 8034 -38440 8074
rect -38384 8077 -31601 8090
rect -31545 8093 -31413 8133
rect -31357 8123 -10923 8149
rect -10867 8139 -10735 8179
rect -10679 8141 -3483 8195
rect -3427 8157 -3295 8197
rect -3239 8166 3710 8213
rect -3239 8157 2415 8166
rect -3427 8150 2415 8157
rect -3427 8141 2227 8150
rect -10679 8139 2227 8141
rect -10867 8123 2227 8139
rect -31357 8108 2227 8123
rect -31357 8093 -17727 8108
rect -31545 8092 -17727 8093
rect -31545 8077 -17915 8092
rect -38384 8036 -17915 8077
rect -17859 8052 -17727 8092
rect -17671 8094 2227 8108
rect 2283 8110 2415 8150
rect 2471 8110 3710 8166
rect 2283 8094 3710 8110
rect -17671 8062 3710 8094
rect -17671 8052 -3032 8062
rect -17859 8044 -3032 8052
rect -17859 8036 -10472 8044
rect -38384 8034 -10472 8036
rect -38572 8026 -10472 8034
rect -38572 8018 -24562 8026
rect -58684 8011 -24562 8018
rect -58872 8010 -24562 8011
rect -58872 8009 -24750 8010
rect -58872 7995 -44878 8009
rect -65244 7985 -44878 7995
rect -65244 7969 -64935 7985
rect -65244 7913 -65123 7969
rect -65067 7929 -64935 7969
rect -64879 7975 -44878 7985
rect -64879 7967 -45112 7975
rect -64879 7945 -45313 7967
rect -64879 7932 -51632 7945
rect -64879 7929 -51846 7932
rect -65067 7916 -51846 7929
rect -65067 7913 -58477 7916
rect -65244 7882 -58477 7913
rect -65244 7874 -58711 7882
rect -65244 7834 -58912 7874
rect -65244 7800 -64672 7834
rect -65244 7792 -64906 7800
rect -65244 7736 -65107 7792
rect -65051 7744 -64906 7792
rect -64850 7778 -64672 7800
rect -64616 7818 -58912 7834
rect -58856 7826 -58711 7874
rect -58655 7860 -58477 7882
rect -58421 7876 -51846 7916
rect -51790 7889 -51632 7932
rect -51576 7936 -45313 7945
rect -51576 7889 -51415 7936
rect -51790 7880 -51415 7889
rect -51359 7911 -45313 7936
rect -45257 7919 -45112 7967
rect -45056 7953 -44878 7975
rect -44822 7998 -24750 8009
rect -44822 7964 -31150 7998
rect -44822 7956 -31384 7964
rect -44822 7953 -31585 7956
rect -45056 7947 -31585 7953
rect -45056 7919 -44691 7947
rect -45257 7911 -44691 7919
rect -51359 7908 -44691 7911
rect -51359 7880 -51185 7908
rect -51790 7876 -51185 7880
rect -58421 7860 -51185 7876
rect -58655 7854 -51185 7860
rect -58655 7826 -58290 7854
rect -58856 7818 -58290 7826
rect -64616 7798 -58290 7818
rect -58234 7852 -51185 7854
rect -51129 7891 -44691 7908
rect -44635 7939 -31585 7947
rect -44635 7905 -38177 7939
rect -44635 7897 -38411 7905
rect -44635 7891 -38612 7897
rect -51129 7852 -38612 7891
rect -58234 7841 -38612 7852
rect -38556 7849 -38411 7897
rect -38355 7883 -38177 7905
rect -38121 7900 -31585 7939
rect -31529 7908 -31384 7956
rect -31328 7942 -31150 7964
rect -31094 7954 -24750 7998
rect -24694 7970 -24562 8010
rect -24506 8010 -10472 8026
rect -24506 8002 -10706 8010
rect -24506 7970 -10907 8002
rect -24694 7957 -10907 7970
rect -24694 7954 -17464 7957
rect -31094 7942 -17464 7954
rect -31328 7936 -17464 7942
rect -31328 7908 -30963 7936
rect -31529 7900 -30963 7908
rect -38121 7883 -30963 7900
rect -38355 7880 -30963 7883
rect -30907 7923 -17464 7936
rect -30907 7915 -17698 7923
rect -30907 7880 -17899 7915
rect -38355 7877 -17899 7880
rect -38355 7849 -37990 7877
rect -38556 7841 -37990 7849
rect -58234 7821 -37990 7841
rect -37934 7875 -17899 7877
rect -37934 7841 -24299 7875
rect -37934 7833 -24533 7841
rect -37934 7821 -24734 7833
rect -58234 7799 -24734 7821
rect -58234 7798 -45095 7799
rect -64616 7786 -45095 7798
rect -64616 7778 -45309 7786
rect -64850 7772 -45309 7778
rect -64850 7744 -64485 7772
rect -65051 7736 -64485 7744
rect -65244 7716 -64485 7736
rect -64429 7730 -45309 7772
rect -45253 7743 -45095 7786
rect -45039 7790 -24734 7799
rect -45039 7743 -44878 7790
rect -45253 7734 -44878 7743
rect -44822 7788 -24734 7790
rect -44822 7775 -31367 7788
rect -44822 7762 -31581 7775
rect -44822 7734 -44648 7762
rect -45253 7730 -44648 7734
rect -64429 7716 -44648 7730
rect -65244 7706 -44648 7716
rect -44592 7729 -31581 7762
rect -44592 7716 -38394 7729
rect -44592 7706 -38608 7716
rect -65244 7693 -58694 7706
rect -65244 7637 -58908 7693
rect -58852 7650 -58694 7693
rect -58638 7697 -38608 7706
rect -58638 7650 -58477 7697
rect -58852 7641 -58477 7650
rect -58421 7669 -38608 7697
rect -58421 7641 -58247 7669
rect -58852 7637 -58247 7641
rect -65244 7624 -58247 7637
rect -65244 7611 -64889 7624
rect -65244 7555 -65103 7611
rect -65047 7568 -64889 7611
rect -64833 7615 -58247 7624
rect -64833 7568 -64672 7615
rect -65047 7559 -64672 7568
rect -64616 7613 -58247 7615
rect -58191 7660 -38608 7669
rect -38552 7673 -38394 7716
rect -38338 7720 -31581 7729
rect -38338 7673 -38177 7720
rect -38552 7664 -38177 7673
rect -38121 7719 -31581 7720
rect -31525 7732 -31367 7775
rect -31311 7779 -24734 7788
rect -31311 7732 -31150 7779
rect -31525 7723 -31150 7732
rect -31094 7777 -24734 7779
rect -24678 7785 -24533 7833
rect -24477 7819 -24299 7841
rect -24243 7859 -17899 7875
rect -17843 7867 -17698 7915
rect -17642 7901 -17464 7923
rect -17408 7946 -10907 7957
rect -10851 7954 -10706 8002
rect -10650 7988 -10472 8010
rect -10416 8028 -3032 8044
rect -10416 8020 -3266 8028
rect -10416 7988 -3467 8020
rect -10650 7982 -3467 7988
rect -10650 7954 -10285 7982
rect -10851 7946 -10285 7954
rect -17408 7926 -10285 7946
rect -10229 7964 -3467 7982
rect -3411 7972 -3266 8020
rect -3210 8006 -3032 8028
rect -2976 8015 3710 8062
rect -2976 8006 2678 8015
rect -3210 8000 2678 8006
rect -3210 7972 -2845 8000
rect -3411 7964 -2845 7972
rect -10229 7944 -2845 7964
rect -2789 7981 2678 8000
rect -2789 7973 2444 7981
rect -2789 7944 2243 7973
rect -10229 7926 2243 7944
rect -17408 7917 2243 7926
rect 2299 7925 2444 7973
rect 2500 7959 2678 7981
rect 2734 7959 3710 8015
rect 2500 7953 3710 7959
rect 2500 7925 2865 7953
rect 2299 7917 2865 7925
rect -17408 7901 2865 7917
rect -17642 7897 2865 7901
rect 2921 7897 3710 7953
rect -17642 7895 3710 7897
rect -17642 7867 -17277 7895
rect -17843 7859 -17277 7867
rect -24243 7839 -17277 7859
rect -17221 7852 3710 7895
rect -17221 7839 -3249 7852
rect -24243 7834 -3463 7839
rect -24243 7821 -10689 7834
rect -24243 7819 -10903 7821
rect -24477 7813 -10903 7819
rect -24477 7785 -24112 7813
rect -24678 7777 -24112 7785
rect -31094 7757 -24112 7777
rect -24056 7765 -10903 7813
rect -10847 7778 -10689 7821
rect -10633 7825 -3463 7834
rect -10633 7778 -10472 7825
rect -10847 7769 -10472 7778
rect -10416 7797 -3463 7825
rect -10416 7769 -10242 7797
rect -10847 7765 -10242 7769
rect -24056 7757 -10242 7765
rect -31094 7751 -10242 7757
rect -31094 7723 -30920 7751
rect -31525 7719 -30920 7723
rect -38121 7695 -30920 7719
rect -30864 7747 -10242 7751
rect -30864 7734 -17681 7747
rect -30864 7695 -17895 7734
rect -38121 7692 -17895 7695
rect -38121 7664 -37947 7692
rect -38552 7660 -37947 7664
rect -58191 7636 -37947 7660
rect -37891 7678 -17895 7692
rect -17839 7691 -17681 7734
rect -17625 7741 -10242 7747
rect -10186 7783 -3463 7797
rect -3407 7796 -3249 7839
rect -3193 7843 3710 7852
rect -3193 7796 -3032 7843
rect -3407 7787 -3032 7796
rect -2976 7815 3710 7843
rect -2976 7787 -2802 7815
rect -3407 7783 -2802 7787
rect -10186 7759 -2802 7783
rect -2746 7805 3710 7815
rect -2746 7792 2461 7805
rect -2746 7759 2247 7792
rect -10186 7741 2247 7759
rect -17625 7738 2247 7741
rect -17625 7691 -17464 7738
rect -17839 7682 -17464 7691
rect -17408 7736 2247 7738
rect 2303 7749 2461 7792
rect 2517 7796 3710 7805
rect 2517 7749 2678 7796
rect 2303 7740 2678 7749
rect 2734 7768 3710 7796
rect 2734 7740 2908 7768
rect 2303 7736 2908 7740
rect -17408 7712 2908 7736
rect 2964 7712 3710 7768
rect -17408 7710 3710 7712
rect -17408 7682 -17234 7710
rect -17839 7678 -17234 7682
rect -37891 7665 -17234 7678
rect -37891 7652 -24516 7665
rect -37891 7636 -24730 7652
rect -58191 7613 -24730 7636
rect -64616 7596 -24730 7613
rect -24674 7609 -24516 7652
rect -24460 7656 -17234 7665
rect -24460 7609 -24299 7656
rect -24674 7600 -24299 7609
rect -24243 7654 -17234 7656
rect -17178 7654 3710 7710
rect -24243 7628 3710 7654
rect -24243 7600 -24069 7628
rect -24674 7596 -24069 7600
rect -64616 7587 -24069 7596
rect -64616 7559 -64442 7587
rect -65047 7555 -64442 7559
rect -65244 7531 -64442 7555
rect -64386 7572 -24069 7587
rect -24013 7572 3710 7628
rect -64386 7531 3710 7572
rect -65244 7440 3710 7531
rect -65244 7424 -51698 7440
rect -65244 7368 -51886 7424
rect -51830 7384 -51698 7424
rect -51642 7384 3710 7440
rect -51830 7368 3710 7384
rect -65244 7289 3710 7368
rect -65244 7255 -51435 7289
rect -65244 7247 -51669 7255
rect -65244 7191 -51870 7247
rect -51814 7199 -51669 7247
rect -51613 7233 -51435 7255
rect -51379 7257 3710 7289
rect -51379 7251 -31396 7257
rect -51379 7235 -38429 7251
rect -51379 7233 -38617 7235
rect -51613 7228 -38617 7233
rect -51613 7227 -45170 7228
rect -51613 7199 -51248 7227
rect -51814 7191 -51248 7199
rect -65244 7187 -51248 7191
rect -65244 7171 -58740 7187
rect -65244 7167 -58928 7171
rect -65244 7151 -64958 7167
rect -65244 7095 -65146 7151
rect -65090 7111 -64958 7151
rect -64902 7115 -58928 7167
rect -58872 7131 -58740 7171
rect -58684 7171 -51248 7187
rect -51192 7212 -45170 7227
rect -51192 7171 -45358 7212
rect -58684 7156 -45358 7171
rect -45302 7172 -45170 7212
rect -45114 7179 -38617 7228
rect -38561 7195 -38429 7235
rect -38373 7241 -31396 7251
rect -38373 7195 -31584 7241
rect -38561 7185 -31584 7195
rect -31528 7201 -31396 7241
rect -31340 7251 3710 7257
rect -31340 7235 -17727 7251
rect -31340 7201 -17915 7235
rect -31528 7193 -17915 7201
rect -31528 7185 -24573 7193
rect -38561 7179 -24573 7185
rect -45114 7177 -24573 7179
rect -45114 7172 -24761 7177
rect -45302 7156 -24761 7172
rect -58684 7131 -24761 7156
rect -58872 7121 -24761 7131
rect -24705 7137 -24573 7177
rect -24517 7179 -17915 7193
rect -17859 7195 -17727 7235
rect -17671 7240 3710 7251
rect -17671 7224 -3225 7240
rect -17671 7210 -3413 7224
rect -17671 7195 -10712 7210
rect -17859 7194 -10712 7195
rect -17859 7179 -10900 7194
rect -24517 7138 -10900 7179
rect -10844 7154 -10712 7194
rect -10656 7168 -3413 7210
rect -3357 7184 -3225 7224
rect -3169 7184 3710 7240
rect -3357 7168 3710 7184
rect -10656 7154 3710 7168
rect -10844 7141 3710 7154
rect -10844 7138 2444 7141
rect -24517 7137 2444 7138
rect -24705 7125 2444 7137
rect -24705 7121 2256 7125
rect -58872 7115 2256 7121
rect -64902 7111 2256 7115
rect -65090 7106 2256 7111
rect -65090 7100 -31133 7106
rect -65090 7095 -38166 7100
rect -65244 7079 -38166 7095
rect -65244 7066 -51652 7079
rect -65244 7036 -51866 7066
rect -65244 7016 -58477 7036
rect -65244 6982 -64695 7016
rect -65244 6974 -64929 6982
rect -65244 6918 -65130 6974
rect -65074 6926 -64929 6974
rect -64873 6960 -64695 6982
rect -64639 7002 -58477 7016
rect -64639 6994 -58711 7002
rect -64639 6960 -58912 6994
rect -64873 6954 -58912 6960
rect -64873 6926 -64508 6954
rect -65074 6918 -64508 6926
rect -65244 6898 -64508 6918
rect -64452 6938 -58912 6954
rect -58856 6946 -58711 6994
rect -58655 6980 -58477 7002
rect -58421 7010 -51866 7036
rect -51810 7023 -51652 7066
rect -51596 7077 -38166 7079
rect -51596 7070 -44907 7077
rect -51596 7023 -51435 7070
rect -51810 7014 -51435 7023
rect -51379 7043 -44907 7070
rect -51379 7042 -45141 7043
rect -51379 7014 -51205 7042
rect -51810 7010 -51205 7014
rect -58421 6986 -51205 7010
rect -51149 7035 -45141 7042
rect -51149 6986 -45342 7035
rect -58421 6980 -45342 6986
rect -58655 6979 -45342 6980
rect -45286 6987 -45141 7035
rect -45085 7021 -44907 7043
rect -44851 7066 -38166 7077
rect -44851 7058 -38400 7066
rect -44851 7021 -38601 7058
rect -45085 7015 -38601 7021
rect -45085 6987 -44720 7015
rect -45286 6979 -44720 6987
rect -58655 6974 -44720 6979
rect -58655 6946 -58290 6974
rect -58856 6938 -58290 6946
rect -64452 6918 -58290 6938
rect -58234 6959 -44720 6974
rect -44664 7002 -38601 7015
rect -38545 7010 -38400 7058
rect -38344 7044 -38166 7066
rect -38110 7072 -31133 7100
rect -38110 7064 -31367 7072
rect -38110 7044 -31568 7064
rect -38344 7038 -31568 7044
rect -38344 7010 -37979 7038
rect -38545 7002 -37979 7010
rect -44664 6982 -37979 7002
rect -37923 7008 -31568 7038
rect -31512 7016 -31367 7064
rect -31311 7050 -31133 7072
rect -31077 7100 2256 7106
rect -31077 7066 -17464 7100
rect -31077 7058 -17698 7066
rect -31077 7050 -17899 7058
rect -31311 7044 -17899 7050
rect -31311 7016 -30946 7044
rect -31512 7008 -30946 7016
rect -37923 6988 -30946 7008
rect -30890 7042 -17899 7044
rect -30890 7008 -24310 7042
rect -30890 7000 -24544 7008
rect -30890 6988 -24745 7000
rect -37923 6982 -24745 6988
rect -44664 6959 -24745 6982
rect -58234 6944 -24745 6959
rect -24689 6952 -24544 7000
rect -24488 6986 -24310 7008
rect -24254 7002 -17899 7042
rect -17843 7010 -17698 7058
rect -17642 7044 -17464 7066
rect -17408 7089 2256 7100
rect -17408 7059 -2962 7089
rect -17408 7044 -10449 7059
rect -17642 7038 -10449 7044
rect -17642 7010 -17277 7038
rect -17843 7002 -17277 7010
rect -24254 6986 -17277 7002
rect -24488 6982 -17277 6986
rect -17221 7025 -10449 7038
rect -17221 7017 -10683 7025
rect -17221 6982 -10884 7017
rect -24488 6980 -10884 6982
rect -24488 6952 -24123 6980
rect -24689 6944 -24123 6952
rect -58234 6924 -24123 6944
rect -24067 6961 -10884 6980
rect -10828 6969 -10683 7017
rect -10627 7003 -10449 7025
rect -10393 7055 -2962 7059
rect -10393 7047 -3196 7055
rect -10393 7003 -3397 7047
rect -10627 6997 -3397 7003
rect -10627 6969 -10262 6997
rect -10828 6961 -10262 6969
rect -24067 6941 -10262 6961
rect -10206 6991 -3397 6997
rect -3341 6999 -3196 7047
rect -3140 7033 -2962 7055
rect -2906 7069 2256 7089
rect 2312 7085 2444 7125
rect 2500 7085 3710 7141
rect 2312 7069 3710 7085
rect -2906 7033 3710 7069
rect -3140 7027 3710 7033
rect -3140 6999 -2775 7027
rect -3341 6991 -2775 6999
rect -10206 6971 -2775 6991
rect -2719 6990 3710 7027
rect -2719 6971 2707 6990
rect -10206 6956 2707 6971
rect -10206 6948 2473 6956
rect -10206 6941 2272 6948
rect -24067 6924 2272 6941
rect -58234 6918 2272 6924
rect -64452 6898 2272 6918
rect -65244 6896 2272 6898
rect -65244 6890 -31350 6896
rect -65244 6877 -38383 6890
rect -65244 6867 -38597 6877
rect -65244 6854 -45124 6867
rect -65244 6826 -45338 6854
rect -65244 6813 -58694 6826
rect -65244 6806 -58908 6813
rect -65244 6793 -64912 6806
rect -65244 6737 -65126 6793
rect -65070 6750 -64912 6793
rect -64856 6797 -58908 6806
rect -64856 6750 -64695 6797
rect -65070 6741 -64695 6750
rect -64639 6769 -58908 6797
rect -64639 6741 -64465 6769
rect -65070 6737 -64465 6741
rect -65244 6713 -64465 6737
rect -64409 6757 -58908 6769
rect -58852 6770 -58694 6813
rect -58638 6817 -45338 6826
rect -58638 6770 -58477 6817
rect -58852 6761 -58477 6770
rect -58421 6798 -45338 6817
rect -45282 6811 -45124 6854
rect -45068 6858 -38597 6867
rect -45068 6811 -44907 6858
rect -45282 6802 -44907 6811
rect -44851 6830 -38597 6858
rect -44851 6802 -44677 6830
rect -45282 6798 -44677 6802
rect -58421 6789 -44677 6798
rect -58421 6761 -58247 6789
rect -58852 6757 -58247 6761
rect -64409 6733 -58247 6757
rect -58191 6774 -44677 6789
rect -44621 6821 -38597 6830
rect -38541 6834 -38383 6877
rect -38327 6883 -31350 6890
rect -38327 6881 -31564 6883
rect -38327 6834 -38166 6881
rect -38541 6825 -38166 6834
rect -38110 6853 -31564 6881
rect -38110 6825 -37936 6853
rect -38541 6821 -37936 6825
rect -44621 6797 -37936 6821
rect -37880 6827 -31564 6853
rect -31508 6840 -31350 6883
rect -31294 6892 2272 6896
rect 2328 6900 2473 6948
rect 2529 6934 2707 6956
rect 2763 6934 3710 6990
rect 2529 6928 3710 6934
rect 2529 6900 2894 6928
rect 2328 6892 2894 6900
rect -31294 6890 2894 6892
rect -31294 6887 -17681 6890
rect -31294 6840 -31133 6887
rect -31508 6831 -31133 6840
rect -31077 6877 -17681 6887
rect -31077 6859 -17895 6877
rect -31077 6831 -30903 6859
rect -31508 6827 -30903 6831
rect -37880 6803 -30903 6827
rect -30847 6832 -17895 6859
rect -30847 6819 -24527 6832
rect -30847 6803 -24741 6819
rect -37880 6797 -24741 6803
rect -44621 6774 -24741 6797
rect -58191 6763 -24741 6774
rect -24685 6776 -24527 6819
rect -24471 6823 -17895 6832
rect -24471 6776 -24310 6823
rect -24685 6767 -24310 6776
rect -24254 6821 -17895 6823
rect -17839 6834 -17681 6877
rect -17625 6881 2894 6890
rect -17625 6834 -17464 6881
rect -17839 6825 -17464 6834
rect -17408 6879 2894 6881
rect -17408 6866 -3179 6879
rect -17408 6853 -3393 6866
rect -17408 6825 -17234 6853
rect -17839 6821 -17234 6825
rect -24254 6797 -17234 6821
rect -17178 6849 -3393 6853
rect -17178 6836 -10666 6849
rect -17178 6797 -10880 6836
rect -24254 6795 -10880 6797
rect -24254 6767 -24080 6795
rect -24685 6763 -24080 6767
rect -58191 6739 -24080 6763
rect -24024 6780 -10880 6795
rect -10824 6793 -10666 6836
rect -10610 6840 -3393 6849
rect -10610 6793 -10449 6840
rect -10824 6784 -10449 6793
rect -10393 6812 -3393 6840
rect -10393 6784 -10219 6812
rect -10824 6780 -10219 6784
rect -24024 6756 -10219 6780
rect -10163 6810 -3393 6812
rect -3337 6823 -3179 6866
rect -3123 6872 2894 6879
rect 2950 6872 3710 6928
rect -3123 6870 3710 6872
rect -3123 6823 -2962 6870
rect -3337 6814 -2962 6823
rect -2906 6842 3710 6870
rect -2906 6814 -2732 6842
rect -3337 6810 -2732 6814
rect -10163 6786 -2732 6810
rect -2676 6786 3710 6842
rect -10163 6780 3710 6786
rect -10163 6767 2490 6780
rect -10163 6756 2276 6767
rect -24024 6739 2276 6756
rect -58191 6733 2276 6739
rect -64409 6713 2276 6733
rect -65244 6711 2276 6713
rect 2332 6724 2490 6767
rect 2546 6771 3710 6780
rect 2546 6724 2707 6771
rect 2332 6715 2707 6724
rect 2763 6743 3710 6771
rect 2763 6715 2937 6743
rect 2332 6711 2937 6715
rect -65244 6687 2937 6711
rect 2993 6687 3710 6743
rect -65244 6530 3710 6687
rect -65244 6454 -63380 6530
rect -65240 4790 -63380 6454
rect -59200 5290 -57340 6530
rect -52179 4941 -50481 6530
rect -45510 4800 -43650 6530
rect -38810 4430 -36950 6530
rect -31760 4950 -29900 6530
rect -24990 4680 -23130 6530
rect -18260 4690 -16400 6530
rect -11400 4460 -9540 6530
rect -3930 4740 -2070 6530
rect 1670 4690 3530 6530
rect -61760 -68247 -61250 -67625
rect -61760 -68318 -60887 -68247
rect -55014 -68282 -54504 -67720
rect -48002 -67728 -47875 -67719
rect -61760 -68334 -61490 -68318
rect -61760 -68390 -61678 -68334
rect -61622 -68374 -61490 -68334
rect -61434 -68374 -60887 -68318
rect -61622 -68390 -60887 -68374
rect -61760 -68437 -60887 -68390
rect -55242 -68377 -54186 -68282
rect -48212 -68311 -47702 -67728
rect -41153 -67756 -41026 -67746
rect -55242 -68433 -54944 -68377
rect -54888 -68433 -54769 -68377
rect -54713 -68433 -54567 -68377
rect -54511 -68433 -54186 -68377
rect -55242 -68437 -54186 -68433
rect -48439 -68367 -47230 -68311
rect -41369 -68326 -40859 -67756
rect -48439 -68423 -48168 -68367
rect -48112 -68423 -47987 -68367
rect -47931 -68373 -47230 -68367
rect -47931 -68423 -47783 -68373
rect -48439 -68429 -47783 -68423
rect -47727 -68429 -47230 -68373
rect -48439 -68437 -47230 -68429
rect -41649 -68367 -40440 -68326
rect -34628 -68353 -34118 -67748
rect -27812 -68160 -27302 -67756
rect -28040 -68350 -26990 -68160
rect -20957 -68263 -20447 -67748
rect -14161 -68255 -13651 -67736
rect -7318 -68255 -6808 -67728
rect -21096 -68350 -20092 -68263
rect -41649 -68371 -41151 -68367
rect -41649 -68427 -41332 -68371
rect -41276 -68423 -41151 -68371
rect -41095 -68377 -40440 -68367
rect -41095 -68423 -40951 -68377
rect -41276 -68427 -40951 -68423
rect -41649 -68433 -40951 -68427
rect -40895 -68433 -40440 -68377
rect -41649 -68437 -40440 -68433
rect -34904 -68406 -33695 -68353
rect -34904 -68437 -34577 -68406
rect -61760 -68462 -34577 -68437
rect -34521 -68413 -33695 -68406
rect -34521 -68462 -34396 -68413
rect -61760 -68469 -34396 -68462
rect -34340 -68469 -34221 -68413
rect -34165 -68437 -33695 -68413
rect -28040 -68386 -26900 -68350
rect -28040 -68437 -27727 -68386
rect -34165 -68442 -27727 -68437
rect -27671 -68393 -26900 -68386
rect -27671 -68442 -27546 -68393
rect -34165 -68449 -27546 -68442
rect -27490 -68449 -27371 -68393
rect -27315 -68437 -26900 -68393
rect -21096 -68386 -19960 -68350
rect -21096 -68437 -20787 -68386
rect -27315 -68442 -20787 -68437
rect -20731 -68393 -19960 -68386
rect -20731 -68442 -20606 -68393
rect -27315 -68449 -20606 -68442
rect -20550 -68449 -20431 -68393
rect -20375 -68437 -19960 -68393
rect -14409 -68379 -13405 -68255
rect -14409 -68435 -14124 -68379
rect -14068 -68384 -13405 -68379
rect -14068 -68435 -13945 -68384
rect -14409 -68437 -13945 -68435
rect -20375 -68440 -13945 -68437
rect -13889 -68440 -13762 -68384
rect -13706 -68437 -13405 -68384
rect -7481 -68359 -6477 -68255
rect -510 -68259 0 -67756
rect 6404 -67829 6681 -67602
rect 6287 -68257 6797 -67829
rect -7481 -68415 -7286 -68359
rect -7230 -68415 -7111 -68359
rect -7055 -68415 -6921 -68359
rect -6865 -68415 -6477 -68359
rect -7481 -68437 -6477 -68415
rect -676 -68356 328 -68259
rect -676 -68359 -70 -68356
rect -676 -68415 -476 -68359
rect -420 -68363 -70 -68359
rect -420 -68415 -283 -68363
rect -676 -68419 -283 -68415
rect -227 -68412 -70 -68363
rect -14 -68412 328 -68356
rect -227 -68419 328 -68412
rect -676 -68437 328 -68419
rect 5835 -68350 6839 -68257
rect 5835 -68406 6318 -68350
rect 6374 -68406 6506 -68350
rect 6562 -68356 6839 -68350
rect 6562 -68406 6708 -68356
rect 5835 -68412 6708 -68406
rect 6764 -68412 6839 -68356
rect 5835 -68437 6839 -68412
rect -13706 -68440 6839 -68437
rect -20375 -68449 6839 -68440
rect -34165 -68469 6839 -68449
rect -61760 -68503 -61227 -68469
rect -61760 -68511 -61461 -68503
rect -61760 -68567 -61662 -68511
rect -61606 -68559 -61461 -68511
rect -61405 -68525 -61227 -68503
rect -61171 -68525 6839 -68469
rect -61405 -68531 6839 -68525
rect -61405 -68559 -61040 -68531
rect -61606 -68567 -61040 -68559
rect -61760 -68587 -61040 -68567
rect -60984 -68540 6839 -68531
rect -60984 -68567 -41330 -68540
rect -60984 -68573 -47916 -68567
rect -60984 -68587 -48152 -68573
rect -61760 -68617 -48152 -68587
rect -61760 -68642 -54725 -68617
rect -61760 -68644 -54925 -68642
rect -61760 -68679 -55157 -68644
rect -61760 -68692 -61444 -68679
rect -61760 -68748 -61658 -68692
rect -61602 -68735 -61444 -68692
rect -61388 -68688 -55157 -68679
rect -61388 -68735 -61227 -68688
rect -61602 -68744 -61227 -68735
rect -61171 -68700 -55157 -68688
rect -55101 -68698 -54925 -68644
rect -54869 -68673 -54725 -68642
rect -54669 -68629 -48152 -68617
rect -48096 -68623 -47916 -68573
rect -47860 -68579 -41330 -68567
rect -47860 -68582 -41517 -68579
rect -47860 -68623 -47656 -68582
rect -48096 -68629 -47656 -68623
rect -54669 -68632 -47656 -68629
rect -54669 -68648 -54294 -68632
rect -54669 -68673 -54507 -68648
rect -54869 -68698 -54507 -68673
rect -55101 -68700 -54507 -68698
rect -61171 -68704 -54507 -68700
rect -54451 -68688 -54294 -68648
rect -54238 -68638 -47656 -68632
rect -47600 -68635 -41517 -68582
rect -41461 -68596 -41330 -68579
rect -41274 -68544 6839 -68540
rect -41274 -68554 -40890 -68544
rect -41274 -68596 -41117 -68554
rect -41461 -68610 -41117 -68596
rect -41061 -68600 -40890 -68554
rect -40834 -68567 6839 -68544
rect -40834 -68600 -40694 -68567
rect -41061 -68610 -40694 -68600
rect -41461 -68623 -40694 -68610
rect -40638 -68571 6839 -68567
rect -40638 -68592 6143 -68571
rect -40638 -68596 145 -68592
rect -40638 -68600 -345 -68596
rect -40638 -68603 -595 -68600
rect -40638 -68609 -27150 -68603
rect -40638 -68623 -27710 -68609
rect -41461 -68629 -34000 -68623
rect -41461 -68635 -34560 -68629
rect -47600 -68638 -34560 -68635
rect -54238 -68648 -34560 -68638
rect -54238 -68688 -34819 -68648
rect -54451 -68704 -34819 -68688
rect -34763 -68685 -34560 -68648
rect -34504 -68685 -34329 -68629
rect -34273 -68679 -34000 -68629
rect -33944 -68628 -27710 -68623
rect -33944 -68679 -27969 -68628
rect -34273 -68684 -27969 -68679
rect -27913 -68665 -27710 -68628
rect -27654 -68665 -27479 -68609
rect -27423 -68659 -27150 -68609
rect -27094 -68609 -20210 -68603
rect -27094 -68628 -20770 -68609
rect -27094 -68659 -21029 -68628
rect -27423 -68665 -21029 -68659
rect -27913 -68684 -21029 -68665
rect -20973 -68665 -20770 -68628
rect -20714 -68665 -20539 -68609
rect -20483 -68659 -20210 -68609
rect -20154 -68609 -595 -68603
rect -20154 -68615 -6648 -68609
rect -20154 -68621 -6909 -68615
rect -20154 -68627 -7129 -68621
rect -20154 -68632 -7402 -68627
rect -20154 -68636 -13637 -68632
rect -20154 -68642 -13845 -68636
rect -20154 -68648 -14037 -68642
rect -20154 -68659 -14262 -68648
rect -20483 -68665 -14262 -68659
rect -20973 -68684 -14262 -68665
rect -34273 -68685 -14262 -68684
rect -34763 -68704 -14262 -68685
rect -14206 -68698 -14037 -68648
rect -13981 -68692 -13845 -68642
rect -13789 -68688 -13637 -68636
rect -13581 -68683 -7402 -68632
rect -7346 -68677 -7129 -68627
rect -7073 -68671 -6909 -68621
rect -6853 -68665 -6648 -68615
rect -6592 -68656 -595 -68609
rect -539 -68652 -345 -68600
rect -289 -68652 -112 -68596
rect -56 -68648 145 -68596
rect 201 -68627 6143 -68592
rect 6199 -68575 6606 -68571
rect 6199 -68627 6395 -68575
rect 201 -68631 6395 -68627
rect 6451 -68627 6606 -68575
rect 6662 -68627 6839 -68571
rect 6451 -68631 6839 -68627
rect 201 -68648 6839 -68631
rect -56 -68652 6839 -68648
rect -539 -68656 6839 -68652
rect -6592 -68665 6839 -68656
rect -6853 -68671 6839 -68665
rect -7073 -68677 6839 -68671
rect -7346 -68683 6839 -68677
rect -13581 -68686 6839 -68683
rect -13581 -68688 5931 -68686
rect -13789 -68692 5931 -68688
rect -13981 -68698 5931 -68692
rect -14206 -68704 5931 -68698
rect -61171 -68716 5931 -68704
rect -61171 -68744 -60997 -68716
rect -61602 -68748 -60997 -68744
rect -61760 -68772 -60997 -68748
rect -60941 -68740 5931 -68716
rect -60941 -68757 -41084 -68740
rect -60941 -68772 -41317 -68757
rect -61760 -68784 -41317 -68772
rect -61760 -68840 -48212 -68784
rect -48156 -68788 -41317 -68784
rect -48156 -68840 -47970 -68788
rect -61760 -68844 -47970 -68840
rect -47914 -68844 -47770 -68788
rect -47714 -68798 -41317 -68788
rect -47714 -68844 -47466 -68798
rect -61760 -68854 -47466 -68844
rect -47410 -68813 -41317 -68798
rect -41261 -68796 -41084 -68757
rect -41028 -68742 5931 -68740
rect 5987 -68742 6839 -68686
rect -41028 -68752 6839 -68742
rect -41028 -68796 -40836 -68752
rect -41261 -68808 -40836 -68796
rect -40780 -68808 6839 -68752
rect -41261 -68812 6839 -68808
rect -41261 -68813 -26993 -68812
rect -47410 -68826 -26993 -68813
rect -47410 -68832 -27731 -68826
rect -47410 -68846 -33843 -68832
rect -47410 -68854 -34581 -68846
rect -61760 -68861 -34581 -68854
rect -61760 -68865 -54696 -68861
rect -61760 -68921 -54921 -68865
rect -54865 -68917 -54696 -68865
rect -54640 -68867 -34581 -68861
rect -54640 -68917 -54438 -68867
rect -54865 -68921 -54438 -68917
rect -61760 -68923 -54438 -68921
rect -54382 -68902 -34581 -68867
rect -34525 -68902 -34346 -68846
rect -34290 -68850 -33843 -68846
rect -34290 -68902 -34106 -68850
rect -54382 -68906 -34106 -68902
rect -34050 -68888 -33843 -68850
rect -33787 -68882 -27731 -68832
rect -27675 -68882 -27496 -68826
rect -27440 -68830 -26993 -68826
rect -27440 -68882 -27256 -68830
rect -33787 -68886 -27256 -68882
rect -27200 -68868 -26993 -68830
rect -26937 -68826 -20053 -68812
rect -26937 -68868 -20791 -68826
rect -27200 -68882 -20791 -68868
rect -20735 -68882 -20556 -68826
rect -20500 -68830 -20053 -68826
rect -20500 -68882 -20316 -68830
rect -27200 -68886 -20316 -68882
rect -20260 -68868 -20053 -68830
rect -19997 -68844 6839 -68812
rect -19997 -68846 -6723 -68844
rect -19997 -68868 -14199 -68846
rect -20260 -68886 -14199 -68868
rect -33787 -68888 -14199 -68886
rect -34050 -68902 -14199 -68888
rect -14143 -68902 -13980 -68846
rect -13924 -68902 -13791 -68846
rect -13735 -68902 -13543 -68846
rect -13487 -68850 -6723 -68846
rect -13487 -68852 -7152 -68850
rect -13487 -68902 -7367 -68852
rect -34050 -68906 -7367 -68902
rect -54382 -68908 -7367 -68906
rect -7311 -68906 -7152 -68852
rect -7096 -68906 -6934 -68850
rect -6878 -68900 -6723 -68850
rect -6667 -68846 6839 -68844
rect -6667 -68850 -308 -68846
rect -6667 -68900 -566 -68850
rect -6878 -68906 -566 -68900
rect -510 -68902 -308 -68850
rect -252 -68850 6839 -68846
rect -252 -68902 -70 -68850
rect -510 -68906 -70 -68902
rect -14 -68852 6327 -68850
rect -14 -68857 6139 -68852
rect -14 -68906 184 -68857
rect -7311 -68908 184 -68906
rect -54382 -68913 184 -68908
rect 240 -68908 6139 -68857
rect 6195 -68906 6327 -68852
rect 6383 -68906 6533 -68850
rect 6589 -68852 6839 -68850
rect 6589 -68906 6737 -68852
rect 6195 -68908 6737 -68906
rect 6793 -68908 6839 -68852
rect 240 -68913 6839 -68908
rect -54382 -68923 6839 -68913
rect -61760 -68945 6839 -68923
rect -61760 -68947 6797 -68945
rect -55242 -68970 -54186 -68947
rect -34904 -68951 -33695 -68947
rect -28040 -68950 -26990 -68947
rect -21096 -68951 -20092 -68947
use cap_mim_2p0fF_CAMMVY  cap_mim_2p0fF_CAMMVY_0
timestamp 1713185578
transform 1 0 -30730 0 1 -30860
box -37410 -36960 37410 36960
<< labels >>
flabel metal5 s -29850 -68800 -29850 -68800 0 FreeSans 17500 0 0 0 M
port 1 nsew
flabel metal5 s -35200 7930 -35200 7930 0 FreeSans 25000 0 0 0 P
port 2 nsew
<< end >>
