magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1343 1019 1343
<< metal1 >>
rect -19 337 19 343
rect -19 311 -13 337
rect 13 311 19 337
rect -19 283 19 311
rect -19 257 -13 283
rect 13 257 19 283
rect -19 229 19 257
rect -19 203 -13 229
rect 13 203 19 229
rect -19 175 19 203
rect -19 149 -13 175
rect 13 149 19 175
rect -19 121 19 149
rect -19 95 -13 121
rect 13 95 19 121
rect -19 67 19 95
rect -19 41 -13 67
rect 13 41 19 67
rect -19 13 19 41
rect -19 -13 -13 13
rect 13 -13 19 13
rect -19 -41 19 -13
rect -19 -67 -13 -41
rect 13 -67 19 -41
rect -19 -95 19 -67
rect -19 -121 -13 -95
rect 13 -121 19 -95
rect -19 -149 19 -121
rect -19 -175 -13 -149
rect 13 -175 19 -149
rect -19 -203 19 -175
rect -19 -229 -13 -203
rect 13 -229 19 -203
rect -19 -257 19 -229
rect -19 -283 -13 -257
rect 13 -283 19 -257
rect -19 -311 19 -283
rect -19 -337 -13 -311
rect 13 -337 19 -311
rect -19 -343 19 -337
<< via1 >>
rect -13 311 13 337
rect -13 257 13 283
rect -13 203 13 229
rect -13 149 13 175
rect -13 95 13 121
rect -13 41 13 67
rect -13 -13 13 13
rect -13 -67 13 -41
rect -13 -121 13 -95
rect -13 -175 13 -149
rect -13 -229 13 -203
rect -13 -283 13 -257
rect -13 -337 13 -311
<< metal2 >>
rect -19 337 19 343
rect -19 311 -13 337
rect 13 311 19 337
rect -19 283 19 311
rect -19 257 -13 283
rect 13 257 19 283
rect -19 229 19 257
rect -19 203 -13 229
rect 13 203 19 229
rect -19 175 19 203
rect -19 149 -13 175
rect 13 149 19 175
rect -19 121 19 149
rect -19 95 -13 121
rect 13 95 19 121
rect -19 67 19 95
rect -19 41 -13 67
rect 13 41 19 67
rect -19 13 19 41
rect -19 -13 -13 13
rect 13 -13 19 13
rect -19 -41 19 -13
rect -19 -67 -13 -41
rect 13 -67 19 -41
rect -19 -95 19 -67
rect -19 -121 -13 -95
rect 13 -121 19 -95
rect -19 -149 19 -121
rect -19 -175 -13 -149
rect 13 -175 19 -149
rect -19 -203 19 -175
rect -19 -229 -13 -203
rect 13 -229 19 -203
rect -19 -257 19 -229
rect -19 -283 -13 -257
rect 13 -283 19 -257
rect -19 -311 19 -283
rect -19 -337 -13 -311
rect 13 -337 19 -311
rect -19 -343 19 -337
<< end >>
