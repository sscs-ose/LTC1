magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -2876 -2128 2876 2128
<< pwell >>
rect -876 -128 876 128
<< nmos >>
rect -764 -60 -664 60
rect -560 -60 -460 60
rect -356 -60 -256 60
rect -152 -60 -52 60
rect 52 -60 152 60
rect 256 -60 356 60
rect 460 -60 560 60
rect 664 -60 764 60
<< ndiff >>
rect -852 23 -764 60
rect -852 -23 -839 23
rect -793 -23 -764 23
rect -852 -60 -764 -23
rect -664 23 -560 60
rect -664 -23 -635 23
rect -589 -23 -560 23
rect -664 -60 -560 -23
rect -460 23 -356 60
rect -460 -23 -431 23
rect -385 -23 -356 23
rect -460 -60 -356 -23
rect -256 23 -152 60
rect -256 -23 -227 23
rect -181 -23 -152 23
rect -256 -60 -152 -23
rect -52 23 52 60
rect -52 -23 -23 23
rect 23 -23 52 23
rect -52 -60 52 -23
rect 152 23 256 60
rect 152 -23 181 23
rect 227 -23 256 23
rect 152 -60 256 -23
rect 356 23 460 60
rect 356 -23 385 23
rect 431 -23 460 23
rect 356 -60 460 -23
rect 560 23 664 60
rect 560 -23 589 23
rect 635 -23 664 23
rect 560 -60 664 -23
rect 764 23 852 60
rect 764 -23 793 23
rect 839 -23 852 23
rect 764 -60 852 -23
<< ndiffc >>
rect -839 -23 -793 23
rect -635 -23 -589 23
rect -431 -23 -385 23
rect -227 -23 -181 23
rect -23 -23 23 23
rect 181 -23 227 23
rect 385 -23 431 23
rect 589 -23 635 23
rect 793 -23 839 23
<< polysilicon >>
rect -764 60 -664 104
rect -560 60 -460 104
rect -356 60 -256 104
rect -152 60 -52 104
rect 52 60 152 104
rect 256 60 356 104
rect 460 60 560 104
rect 664 60 764 104
rect -764 -104 -664 -60
rect -560 -104 -460 -60
rect -356 -104 -256 -60
rect -152 -104 -52 -60
rect 52 -104 152 -60
rect 256 -104 356 -60
rect 460 -104 560 -60
rect 664 -104 764 -60
<< metal1 >>
rect -839 23 -793 58
rect -839 -58 -793 -23
rect -635 23 -589 58
rect -635 -58 -589 -23
rect -431 23 -385 58
rect -431 -58 -385 -23
rect -227 23 -181 58
rect -227 -58 -181 -23
rect -23 23 23 58
rect -23 -58 23 -23
rect 181 23 227 58
rect 181 -58 227 -23
rect 385 23 431 58
rect 385 -58 431 -23
rect 589 23 635 58
rect 589 -58 635 -23
rect 793 23 839 58
rect 793 -58 839 -23
<< end >>
