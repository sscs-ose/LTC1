magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -7937 -2115 7937 2115
<< metal4 >>
rect -5931 99 5931 109
rect -5931 43 -5921 99
rect -5865 43 -5779 99
rect -5723 43 -5637 99
rect -5581 43 -5495 99
rect -5439 43 -5353 99
rect -5297 43 -5211 99
rect -5155 43 -5069 99
rect -5013 43 -4927 99
rect -4871 43 -4785 99
rect -4729 43 -4643 99
rect -4587 43 -4501 99
rect -4445 43 -4359 99
rect -4303 43 -4217 99
rect -4161 43 -4075 99
rect -4019 43 -3933 99
rect -3877 43 -3791 99
rect -3735 43 -3649 99
rect -3593 43 -3507 99
rect -3451 43 -3365 99
rect -3309 43 -3223 99
rect -3167 43 -3081 99
rect -3025 43 -2939 99
rect -2883 43 -2797 99
rect -2741 43 -2655 99
rect -2599 43 -2513 99
rect -2457 43 -2371 99
rect -2315 43 -2229 99
rect -2173 43 -2087 99
rect -2031 43 -1945 99
rect -1889 43 -1803 99
rect -1747 43 -1661 99
rect -1605 43 -1519 99
rect -1463 43 -1377 99
rect -1321 43 -1235 99
rect -1179 43 -1093 99
rect -1037 43 -951 99
rect -895 43 -809 99
rect -753 43 -667 99
rect -611 43 -525 99
rect -469 43 -383 99
rect -327 43 -241 99
rect -185 43 -99 99
rect -43 43 43 99
rect 99 43 185 99
rect 241 43 327 99
rect 383 43 469 99
rect 525 43 611 99
rect 667 43 753 99
rect 809 43 895 99
rect 951 43 1037 99
rect 1093 43 1179 99
rect 1235 43 1321 99
rect 1377 43 1463 99
rect 1519 43 1605 99
rect 1661 43 1747 99
rect 1803 43 1889 99
rect 1945 43 2031 99
rect 2087 43 2173 99
rect 2229 43 2315 99
rect 2371 43 2457 99
rect 2513 43 2599 99
rect 2655 43 2741 99
rect 2797 43 2883 99
rect 2939 43 3025 99
rect 3081 43 3167 99
rect 3223 43 3309 99
rect 3365 43 3451 99
rect 3507 43 3593 99
rect 3649 43 3735 99
rect 3791 43 3877 99
rect 3933 43 4019 99
rect 4075 43 4161 99
rect 4217 43 4303 99
rect 4359 43 4445 99
rect 4501 43 4587 99
rect 4643 43 4729 99
rect 4785 43 4871 99
rect 4927 43 5013 99
rect 5069 43 5155 99
rect 5211 43 5297 99
rect 5353 43 5439 99
rect 5495 43 5581 99
rect 5637 43 5723 99
rect 5779 43 5865 99
rect 5921 43 5931 99
rect -5931 -43 5931 43
rect -5931 -99 -5921 -43
rect -5865 -99 -5779 -43
rect -5723 -99 -5637 -43
rect -5581 -99 -5495 -43
rect -5439 -99 -5353 -43
rect -5297 -99 -5211 -43
rect -5155 -99 -5069 -43
rect -5013 -99 -4927 -43
rect -4871 -99 -4785 -43
rect -4729 -99 -4643 -43
rect -4587 -99 -4501 -43
rect -4445 -99 -4359 -43
rect -4303 -99 -4217 -43
rect -4161 -99 -4075 -43
rect -4019 -99 -3933 -43
rect -3877 -99 -3791 -43
rect -3735 -99 -3649 -43
rect -3593 -99 -3507 -43
rect -3451 -99 -3365 -43
rect -3309 -99 -3223 -43
rect -3167 -99 -3081 -43
rect -3025 -99 -2939 -43
rect -2883 -99 -2797 -43
rect -2741 -99 -2655 -43
rect -2599 -99 -2513 -43
rect -2457 -99 -2371 -43
rect -2315 -99 -2229 -43
rect -2173 -99 -2087 -43
rect -2031 -99 -1945 -43
rect -1889 -99 -1803 -43
rect -1747 -99 -1661 -43
rect -1605 -99 -1519 -43
rect -1463 -99 -1377 -43
rect -1321 -99 -1235 -43
rect -1179 -99 -1093 -43
rect -1037 -99 -951 -43
rect -895 -99 -809 -43
rect -753 -99 -667 -43
rect -611 -99 -525 -43
rect -469 -99 -383 -43
rect -327 -99 -241 -43
rect -185 -99 -99 -43
rect -43 -99 43 -43
rect 99 -99 185 -43
rect 241 -99 327 -43
rect 383 -99 469 -43
rect 525 -99 611 -43
rect 667 -99 753 -43
rect 809 -99 895 -43
rect 951 -99 1037 -43
rect 1093 -99 1179 -43
rect 1235 -99 1321 -43
rect 1377 -99 1463 -43
rect 1519 -99 1605 -43
rect 1661 -99 1747 -43
rect 1803 -99 1889 -43
rect 1945 -99 2031 -43
rect 2087 -99 2173 -43
rect 2229 -99 2315 -43
rect 2371 -99 2457 -43
rect 2513 -99 2599 -43
rect 2655 -99 2741 -43
rect 2797 -99 2883 -43
rect 2939 -99 3025 -43
rect 3081 -99 3167 -43
rect 3223 -99 3309 -43
rect 3365 -99 3451 -43
rect 3507 -99 3593 -43
rect 3649 -99 3735 -43
rect 3791 -99 3877 -43
rect 3933 -99 4019 -43
rect 4075 -99 4161 -43
rect 4217 -99 4303 -43
rect 4359 -99 4445 -43
rect 4501 -99 4587 -43
rect 4643 -99 4729 -43
rect 4785 -99 4871 -43
rect 4927 -99 5013 -43
rect 5069 -99 5155 -43
rect 5211 -99 5297 -43
rect 5353 -99 5439 -43
rect 5495 -99 5581 -43
rect 5637 -99 5723 -43
rect 5779 -99 5865 -43
rect 5921 -99 5931 -43
rect -5931 -109 5931 -99
<< via4 >>
rect -5921 43 -5865 99
rect -5779 43 -5723 99
rect -5637 43 -5581 99
rect -5495 43 -5439 99
rect -5353 43 -5297 99
rect -5211 43 -5155 99
rect -5069 43 -5013 99
rect -4927 43 -4871 99
rect -4785 43 -4729 99
rect -4643 43 -4587 99
rect -4501 43 -4445 99
rect -4359 43 -4303 99
rect -4217 43 -4161 99
rect -4075 43 -4019 99
rect -3933 43 -3877 99
rect -3791 43 -3735 99
rect -3649 43 -3593 99
rect -3507 43 -3451 99
rect -3365 43 -3309 99
rect -3223 43 -3167 99
rect -3081 43 -3025 99
rect -2939 43 -2883 99
rect -2797 43 -2741 99
rect -2655 43 -2599 99
rect -2513 43 -2457 99
rect -2371 43 -2315 99
rect -2229 43 -2173 99
rect -2087 43 -2031 99
rect -1945 43 -1889 99
rect -1803 43 -1747 99
rect -1661 43 -1605 99
rect -1519 43 -1463 99
rect -1377 43 -1321 99
rect -1235 43 -1179 99
rect -1093 43 -1037 99
rect -951 43 -895 99
rect -809 43 -753 99
rect -667 43 -611 99
rect -525 43 -469 99
rect -383 43 -327 99
rect -241 43 -185 99
rect -99 43 -43 99
rect 43 43 99 99
rect 185 43 241 99
rect 327 43 383 99
rect 469 43 525 99
rect 611 43 667 99
rect 753 43 809 99
rect 895 43 951 99
rect 1037 43 1093 99
rect 1179 43 1235 99
rect 1321 43 1377 99
rect 1463 43 1519 99
rect 1605 43 1661 99
rect 1747 43 1803 99
rect 1889 43 1945 99
rect 2031 43 2087 99
rect 2173 43 2229 99
rect 2315 43 2371 99
rect 2457 43 2513 99
rect 2599 43 2655 99
rect 2741 43 2797 99
rect 2883 43 2939 99
rect 3025 43 3081 99
rect 3167 43 3223 99
rect 3309 43 3365 99
rect 3451 43 3507 99
rect 3593 43 3649 99
rect 3735 43 3791 99
rect 3877 43 3933 99
rect 4019 43 4075 99
rect 4161 43 4217 99
rect 4303 43 4359 99
rect 4445 43 4501 99
rect 4587 43 4643 99
rect 4729 43 4785 99
rect 4871 43 4927 99
rect 5013 43 5069 99
rect 5155 43 5211 99
rect 5297 43 5353 99
rect 5439 43 5495 99
rect 5581 43 5637 99
rect 5723 43 5779 99
rect 5865 43 5921 99
rect -5921 -99 -5865 -43
rect -5779 -99 -5723 -43
rect -5637 -99 -5581 -43
rect -5495 -99 -5439 -43
rect -5353 -99 -5297 -43
rect -5211 -99 -5155 -43
rect -5069 -99 -5013 -43
rect -4927 -99 -4871 -43
rect -4785 -99 -4729 -43
rect -4643 -99 -4587 -43
rect -4501 -99 -4445 -43
rect -4359 -99 -4303 -43
rect -4217 -99 -4161 -43
rect -4075 -99 -4019 -43
rect -3933 -99 -3877 -43
rect -3791 -99 -3735 -43
rect -3649 -99 -3593 -43
rect -3507 -99 -3451 -43
rect -3365 -99 -3309 -43
rect -3223 -99 -3167 -43
rect -3081 -99 -3025 -43
rect -2939 -99 -2883 -43
rect -2797 -99 -2741 -43
rect -2655 -99 -2599 -43
rect -2513 -99 -2457 -43
rect -2371 -99 -2315 -43
rect -2229 -99 -2173 -43
rect -2087 -99 -2031 -43
rect -1945 -99 -1889 -43
rect -1803 -99 -1747 -43
rect -1661 -99 -1605 -43
rect -1519 -99 -1463 -43
rect -1377 -99 -1321 -43
rect -1235 -99 -1179 -43
rect -1093 -99 -1037 -43
rect -951 -99 -895 -43
rect -809 -99 -753 -43
rect -667 -99 -611 -43
rect -525 -99 -469 -43
rect -383 -99 -327 -43
rect -241 -99 -185 -43
rect -99 -99 -43 -43
rect 43 -99 99 -43
rect 185 -99 241 -43
rect 327 -99 383 -43
rect 469 -99 525 -43
rect 611 -99 667 -43
rect 753 -99 809 -43
rect 895 -99 951 -43
rect 1037 -99 1093 -43
rect 1179 -99 1235 -43
rect 1321 -99 1377 -43
rect 1463 -99 1519 -43
rect 1605 -99 1661 -43
rect 1747 -99 1803 -43
rect 1889 -99 1945 -43
rect 2031 -99 2087 -43
rect 2173 -99 2229 -43
rect 2315 -99 2371 -43
rect 2457 -99 2513 -43
rect 2599 -99 2655 -43
rect 2741 -99 2797 -43
rect 2883 -99 2939 -43
rect 3025 -99 3081 -43
rect 3167 -99 3223 -43
rect 3309 -99 3365 -43
rect 3451 -99 3507 -43
rect 3593 -99 3649 -43
rect 3735 -99 3791 -43
rect 3877 -99 3933 -43
rect 4019 -99 4075 -43
rect 4161 -99 4217 -43
rect 4303 -99 4359 -43
rect 4445 -99 4501 -43
rect 4587 -99 4643 -43
rect 4729 -99 4785 -43
rect 4871 -99 4927 -43
rect 5013 -99 5069 -43
rect 5155 -99 5211 -43
rect 5297 -99 5353 -43
rect 5439 -99 5495 -43
rect 5581 -99 5637 -43
rect 5723 -99 5779 -43
rect 5865 -99 5921 -43
<< metal5 >>
rect -5937 99 5937 115
rect -5937 43 -5921 99
rect -5865 43 -5779 99
rect -5723 43 -5637 99
rect -5581 43 -5495 99
rect -5439 43 -5353 99
rect -5297 43 -5211 99
rect -5155 43 -5069 99
rect -5013 43 -4927 99
rect -4871 43 -4785 99
rect -4729 43 -4643 99
rect -4587 43 -4501 99
rect -4445 43 -4359 99
rect -4303 43 -4217 99
rect -4161 43 -4075 99
rect -4019 43 -3933 99
rect -3877 43 -3791 99
rect -3735 43 -3649 99
rect -3593 43 -3507 99
rect -3451 43 -3365 99
rect -3309 43 -3223 99
rect -3167 43 -3081 99
rect -3025 43 -2939 99
rect -2883 43 -2797 99
rect -2741 43 -2655 99
rect -2599 43 -2513 99
rect -2457 43 -2371 99
rect -2315 43 -2229 99
rect -2173 43 -2087 99
rect -2031 43 -1945 99
rect -1889 43 -1803 99
rect -1747 43 -1661 99
rect -1605 43 -1519 99
rect -1463 43 -1377 99
rect -1321 43 -1235 99
rect -1179 43 -1093 99
rect -1037 43 -951 99
rect -895 43 -809 99
rect -753 43 -667 99
rect -611 43 -525 99
rect -469 43 -383 99
rect -327 43 -241 99
rect -185 43 -99 99
rect -43 43 43 99
rect 99 43 185 99
rect 241 43 327 99
rect 383 43 469 99
rect 525 43 611 99
rect 667 43 753 99
rect 809 43 895 99
rect 951 43 1037 99
rect 1093 43 1179 99
rect 1235 43 1321 99
rect 1377 43 1463 99
rect 1519 43 1605 99
rect 1661 43 1747 99
rect 1803 43 1889 99
rect 1945 43 2031 99
rect 2087 43 2173 99
rect 2229 43 2315 99
rect 2371 43 2457 99
rect 2513 43 2599 99
rect 2655 43 2741 99
rect 2797 43 2883 99
rect 2939 43 3025 99
rect 3081 43 3167 99
rect 3223 43 3309 99
rect 3365 43 3451 99
rect 3507 43 3593 99
rect 3649 43 3735 99
rect 3791 43 3877 99
rect 3933 43 4019 99
rect 4075 43 4161 99
rect 4217 43 4303 99
rect 4359 43 4445 99
rect 4501 43 4587 99
rect 4643 43 4729 99
rect 4785 43 4871 99
rect 4927 43 5013 99
rect 5069 43 5155 99
rect 5211 43 5297 99
rect 5353 43 5439 99
rect 5495 43 5581 99
rect 5637 43 5723 99
rect 5779 43 5865 99
rect 5921 43 5937 99
rect -5937 -43 5937 43
rect -5937 -99 -5921 -43
rect -5865 -99 -5779 -43
rect -5723 -99 -5637 -43
rect -5581 -99 -5495 -43
rect -5439 -99 -5353 -43
rect -5297 -99 -5211 -43
rect -5155 -99 -5069 -43
rect -5013 -99 -4927 -43
rect -4871 -99 -4785 -43
rect -4729 -99 -4643 -43
rect -4587 -99 -4501 -43
rect -4445 -99 -4359 -43
rect -4303 -99 -4217 -43
rect -4161 -99 -4075 -43
rect -4019 -99 -3933 -43
rect -3877 -99 -3791 -43
rect -3735 -99 -3649 -43
rect -3593 -99 -3507 -43
rect -3451 -99 -3365 -43
rect -3309 -99 -3223 -43
rect -3167 -99 -3081 -43
rect -3025 -99 -2939 -43
rect -2883 -99 -2797 -43
rect -2741 -99 -2655 -43
rect -2599 -99 -2513 -43
rect -2457 -99 -2371 -43
rect -2315 -99 -2229 -43
rect -2173 -99 -2087 -43
rect -2031 -99 -1945 -43
rect -1889 -99 -1803 -43
rect -1747 -99 -1661 -43
rect -1605 -99 -1519 -43
rect -1463 -99 -1377 -43
rect -1321 -99 -1235 -43
rect -1179 -99 -1093 -43
rect -1037 -99 -951 -43
rect -895 -99 -809 -43
rect -753 -99 -667 -43
rect -611 -99 -525 -43
rect -469 -99 -383 -43
rect -327 -99 -241 -43
rect -185 -99 -99 -43
rect -43 -99 43 -43
rect 99 -99 185 -43
rect 241 -99 327 -43
rect 383 -99 469 -43
rect 525 -99 611 -43
rect 667 -99 753 -43
rect 809 -99 895 -43
rect 951 -99 1037 -43
rect 1093 -99 1179 -43
rect 1235 -99 1321 -43
rect 1377 -99 1463 -43
rect 1519 -99 1605 -43
rect 1661 -99 1747 -43
rect 1803 -99 1889 -43
rect 1945 -99 2031 -43
rect 2087 -99 2173 -43
rect 2229 -99 2315 -43
rect 2371 -99 2457 -43
rect 2513 -99 2599 -43
rect 2655 -99 2741 -43
rect 2797 -99 2883 -43
rect 2939 -99 3025 -43
rect 3081 -99 3167 -43
rect 3223 -99 3309 -43
rect 3365 -99 3451 -43
rect 3507 -99 3593 -43
rect 3649 -99 3735 -43
rect 3791 -99 3877 -43
rect 3933 -99 4019 -43
rect 4075 -99 4161 -43
rect 4217 -99 4303 -43
rect 4359 -99 4445 -43
rect 4501 -99 4587 -43
rect 4643 -99 4729 -43
rect 4785 -99 4871 -43
rect 4927 -99 5013 -43
rect 5069 -99 5155 -43
rect 5211 -99 5297 -43
rect 5353 -99 5439 -43
rect 5495 -99 5581 -43
rect 5637 -99 5723 -43
rect 5779 -99 5865 -43
rect 5921 -99 5937 -43
rect -5937 -115 5937 -99
<< end >>
