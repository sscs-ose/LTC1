magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2045 -3314 2045 3314
<< psubdiff >>
rect -45 1292 45 1314
rect -45 -1292 -23 1292
rect 23 -1292 45 1292
rect -45 -1314 45 -1292
<< psubdiffcont >>
rect -23 -1292 23 1292
<< metal1 >>
rect -34 1292 34 1303
rect -34 -1292 -23 1292
rect 23 -1292 34 1292
rect -34 -1303 34 -1292
<< end >>
