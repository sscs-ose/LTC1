** sch_path: /home/shahid/GF180Projects/PFD/xschem/4x1_mux_test.sch
**.subckt 4x1_mux_test
V1 VDD VSS 3.3
.save i(v1)
V2 VSS GND 0
.save i(v2)
V4 S0 VSS pulse(3.3 0 0 100p 100p 400n 800n)
.save i(v4)
V6 I0 VSS pulse(0 3.3 0 100p 100p 200n 400n)3.3
.save i(v6)
V7 I1 VSS pulse(0 3.3 0 100p 100p 100n 200n)
.save i(v7)
x1 VDD S1 VSS I0 I1 S0 I0 I1 OUT 4x1_mux
V5 S1 VSS pulse(3.3 0 0 100p 100p 200n 400n)
.save i(v5)
**** begin user architecture code

.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical



.control
save all
tran 50p 800n
plot v(S0) v(S1)+4  v(I0)+8 v(I1)+12  v(OUT)+16


*write test_nfet_03v3.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  4x1_mux.sym # of pins=9
** sym_path: /home/shahid/GF180Projects/PFD/xschem/4x1_mux.sym
** sch_path: /home/shahid/GF180Projects/PFD/xschem/4x1_mux.sch
.subckt 4x1_mux VDD S1 VSS I2 I3 S0 I0 I1 OUT
*.iopin VDD
*.iopin VSS
*.ipin S1
*.opin OUT
*.ipin I2
*.ipin I3
*.ipin S0
*.ipin I0
*.ipin I1
x1 VSS S0 net1 I0 I1 VDD 2x1_mux
x2 VSS S0 net2 I2 I3 VDD 2x1_mux
x3 VSS S1 OUT net1 net2 VDD 2x1_mux
.ends


* expanding   symbol:  2x1_mux.sym # of pins=6
** sym_path: /home/shahid/GF180Projects/PFD/xschem/2x1_mux.sym
** sch_path: /home/shahid/GF180Projects/PFD/xschem/2x1_mux.sch
.subckt 2x1_mux VSS Sel OUT I0 I1 VDD
*.iopin VDD
*.iopin VSS
*.ipin Sel
*.opin OUT
*.ipin I0
*.ipin I1
x1 net1 VSS VDD net2 I0 NAND
x2 Sel VSS VDD net3 I1 NAND
x3 net2 VSS VDD OUT net3 NAND
x4 VSS Sel net1 VDD inv_my
.ends


* expanding   symbol:  NAND.sym # of pins=5
** sym_path: /home/shahid/GF180Projects/PFD/xschem/NAND.sym
** sch_path: /home/shahid/GF180Projects/PFD/xschem/NAND.sch
.subckt NAND IN1 VSS VDD OUT IN2
*.ipin IN2
*.ipin IN1
*.iopin VSS
*.iopin VDD
*.opin OUT
XM1 OUT IN2 VDD VDD pfet_03v3_dss L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM2 OUT IN1 VDD VDD pfet_03v3_dss L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM3 net1 IN2 VSS VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM4 OUT IN1 net1 VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
.ends


* expanding   symbol:  inv_my.sym # of pins=4
** sym_path: /home/shahid/GF180Projects/PFD/xschem/inv_my.sym
** sch_path: /home/shahid/GF180Projects/PFD/xschem/inv_my.sch
.subckt inv_my VSS IN OUT VDD
*.iopin VDD
*.iopin VSS
*.ipin IN
*.opin OUT
XM1 OUT IN VSS VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 OUT IN VDD VDD pfet_03v3 L=0.28u W=0.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends

.GLOBAL GND
.end
