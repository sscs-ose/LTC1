magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -6369 -2045 6369 2045
<< psubdiff >>
rect -4369 23 4369 45
rect -4369 -23 -4347 23
rect 4347 -23 4369 23
rect -4369 -45 4369 -23
<< psubdiffcont >>
rect -4347 -23 4347 23
<< metal1 >>
rect -4358 23 4358 34
rect -4358 -23 -4347 23
rect 4347 -23 4358 23
rect -4358 -34 4358 -23
<< end >>
