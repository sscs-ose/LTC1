magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1100 -1046 1100 1046
<< metal1 >>
rect -100 40 100 46
rect -100 14 -94 40
rect -68 14 -40 40
rect -14 14 14 40
rect 40 14 68 40
rect 94 14 100 40
rect -100 -14 100 14
rect -100 -40 -94 -14
rect -68 -40 -40 -14
rect -14 -40 14 -14
rect 40 -40 68 -14
rect 94 -40 100 -14
rect -100 -46 100 -40
<< via1 >>
rect -94 14 -68 40
rect -40 14 -14 40
rect 14 14 40 40
rect 68 14 94 40
rect -94 -40 -68 -14
rect -40 -40 -14 -14
rect 14 -40 40 -14
rect 68 -40 94 -14
<< metal2 >>
rect -100 40 100 46
rect -100 14 -94 40
rect -68 14 -40 40
rect -14 14 14 40
rect 40 14 68 40
rect 94 14 100 40
rect -100 -14 100 14
rect -100 -40 -94 -14
rect -68 -40 -40 -14
rect -14 -40 14 -14
rect 40 -40 68 -14
rect 94 -40 100 -14
rect -100 -46 100 -40
<< end >>
