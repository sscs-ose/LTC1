magic
tech gf180mcuC
magscale 1 10
timestamp 1692806124
<< nwell >>
rect -64 804 500 863
rect -64 763 685 804
rect -64 708 681 763
rect -64 682 500 708
rect 295 365 304 418
rect 345 366 354 417
rect 386 361 388 418
rect 485 417 528 421
rect 436 414 484 417
rect 485 414 529 417
rect 436 365 447 414
rect 485 364 528 414
<< psubdiff >>
rect 13 -105 402 -91
rect 13 -151 75 -105
rect 333 -151 402 -105
rect 13 -167 402 -151
<< nsubdiff >>
rect 41 774 395 826
rect 41 728 85 774
rect 312 728 395 774
rect 41 710 395 728
<< psubdiffcont >>
rect 75 -151 333 -105
<< nsubdiffcont >>
rect 85 728 312 774
<< polysilicon >>
rect 289 421 369 427
rect 112 334 166 421
rect 63 318 166 334
rect 63 268 81 318
rect 130 268 166 318
rect 63 254 166 268
rect 112 200 166 254
rect 272 414 369 421
rect 272 366 300 414
rect 348 366 369 414
rect 272 360 369 366
rect 432 414 528 427
rect 432 366 447 414
rect 495 366 528 414
rect 272 350 368 360
rect 432 350 528 366
rect 272 200 328 350
rect 432 200 488 350
<< polycontact >>
rect 81 268 130 318
rect 300 366 348 414
rect 447 366 495 414
<< metal1 >>
rect -64 804 500 863
rect -64 774 685 804
rect -64 728 85 774
rect 312 763 685 774
rect 312 728 681 763
rect -64 708 681 728
rect 32 471 89 708
rect 186 470 253 545
rect 354 473 411 708
rect 63 325 144 334
rect 10 318 144 325
rect 10 278 81 318
rect 63 268 81 278
rect 130 268 144 318
rect 63 254 144 268
rect 191 314 243 470
rect 515 465 634 630
rect 289 414 388 418
rect 289 366 300 414
rect 348 366 388 414
rect 289 361 388 366
rect 436 414 537 417
rect 436 366 447 414
rect 495 366 537 414
rect 289 360 369 361
rect 436 360 537 366
rect 583 373 634 465
rect 583 314 680 373
rect 191 301 671 314
rect 191 265 634 301
rect 980 300 1066 362
rect 34 -79 88 149
rect 517 25 566 265
rect 662 -79 720 7
rect -70 -105 720 -79
rect -70 -151 75 -105
rect 333 -151 720 -105
rect -70 -188 720 -151
use GF_INV_MAG  GF_INV_MAG_0
timestamp 1692764011
transform 1 0 780 0 1 173
box -118 -175 286 631
use nmos_3p3_VGTVWA  nmos_3p3_VGTVWA_0
timestamp 1692764011
transform 1 0 300 0 1 90
box -140 -134 140 134
use nmos_3p3_VGTVWA  nmos_3p3_VGTVWA_1
timestamp 1692764011
transform 1 0 140 0 1 90
box -140 -134 140 134
use nmos_3p3_VGTVWA  nmos_3p3_VGTVWA_2
timestamp 1692764011
transform 1 0 460 0 1 90
box -140 -134 140 134
use pmos_3p3_M8SWPS  pmos_3p3_M8SWPS_0
timestamp 1692764011
transform 1 0 460 0 1 545
box -202 -210 202 210
use pmos_3p3_M8SWPS  pmos_3p3_M8SWPS_1
timestamp 1692764011
transform 1 0 140 0 1 545
box -202 -210 202 210
use pmos_3p3_M8SWPS  pmos_3p3_M8SWPS_2
timestamp 1692764011
transform 1 0 300 0 1 545
box -202 -210 202 210
<< labels >>
flabel nsubdiffcont 196 756 196 756 0 FreeSans 480 0 0 0 VDD
port 3 nsew
flabel psubdiffcont 200 -126 200 -126 0 FreeSans 480 0 0 0 VSS
port 4 nsew
flabel space 200 -126 571 44 0 FreeSans 480 0 0 0 VSS
port 5 nsew
flabel metal1 24 302 24 302 0 FreeSans 320 0 0 0 IN3
port 8 nsew
flabel metal1 375 388 375 388 0 FreeSans 320 0 0 0 IN2
port 9 nsew
flabel metal1 529 390 529 390 0 FreeSans 320 0 0 0 IN1
port 11 nsew
flabel metal1 1057 325 1057 325 0 FreeSans 320 0 0 0 OUT
port 12 nsew
<< end >>
