* NGSPICE file created from TG_Layout_flat.ext - technology: gf180mcuC

.subckt TG_Layout_flat CLK VIN VOUT VDD VSS
X0 VOUT Inverter_Layout_0.OUT.t0 VIN.t48 VDD.t15 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1 VOUT Inverter_Layout_0.OUT.t1 VIN.t47 VDD.t14 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X2 VIN CLK.t0 VOUT.t59 VSS.t7 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X3 VOUT CLK.t1 VIN.t4 VSS.t6 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X4 VOUT CLK.t2 VIN.t5 VSS.t5 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X5 VSS CLK.t3 Inverter_Layout_0.OUT VSS.t8 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X6 VIN Inverter_Layout_0.OUT.t2 VOUT.t54 VDD.t7 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X7 VOUT Inverter_Layout_0.OUT.t3 VIN.t46 VDD.t12 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X8 VOUT Inverter_Layout_0.OUT.t4 VIN.t45 VDD.t6 pfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X9 VOUT Inverter_Layout_0.OUT.t5 VIN.t44 VDD.t5 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X10 VIN Inverter_Layout_0.OUT.t6 VOUT.t50 VDD.t9 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X11 VOUT CLK.t4 VIN.t2 VSS.t3 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X12 VIN CLK.t5 VOUT.t6 VSS.t2 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X13 VIN Inverter_Layout_0.OUT.t7 VOUT.t49 VDD.t3 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X14 VIN Inverter_Layout_0.OUT.t8 VOUT.t48 VDD.t1 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X15 VIN CLK.t6 VOUT.t61 VSS.t4 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X16 VOUT CLK.t7 VIN.t57 VSS.t1 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X17 VOUT Inverter_Layout_0.OUT.t9 VIN.t43 VDD.t2 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X18 VOUT Inverter_Layout_0.OUT.t10 VIN.t42 VDD.t13 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X19 VOUT Inverter_Layout_0.OUT.t11 VIN.t41 VDD.t15 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X20 VOUT Inverter_Layout_0.OUT.t12 VIN.t40 VDD.t14 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X21 VIN Inverter_Layout_0.OUT.t13 VOUT.t43 VDD.t0 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X22 VIN Inverter_Layout_0.OUT.t14 VOUT.t42 VDD.t10 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X23 VIN CLK.t8 VOUT.t60 VSS.t7 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X24 VIN Inverter_Layout_0.OUT.t15 VOUT.t41 VDD.t11 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X25 VOUT CLK.t9 VIN.t66 VSS.t6 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X26 VOUT Inverter_Layout_0.OUT.t16 VIN.t39 VDD.t8 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X27 VIN Inverter_Layout_0.OUT.t17 VOUT.t39 VDD.t4 pfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X28 VIN Inverter_Layout_0.OUT.t18 VOUT.t38 VDD.t7 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X29 VIN CLK.t10 VOUT.t69 VSS.t0 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X30 VOUT Inverter_Layout_0.OUT.t19 VIN.t38 VDD.t6 pfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X31 VOUT Inverter_Layout_0.OUT.t20 VIN.t37 VDD.t5 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X32 VOUT CLK.t11 VIN.t68 VSS.t5 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X33 VDD CLK.t12 Inverter_Layout_0.OUT VDD.t16 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X34 VIN Inverter_Layout_0.OUT.t21 VOUT.t35 VDD.t3 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X35 VIN CLK.t13 VOUT.t64 VSS.t4 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X36 VOUT CLK.t14 VIN.t3 VSS.t1 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X37 VOUT Inverter_Layout_0.OUT.t22 VIN.t36 VDD.t13 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X38 VIN Inverter_Layout_0.OUT.t23 VOUT.t33 VDD.t1 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X39 VIN Inverter_Layout_0.OUT.t24 VOUT.t32 VDD.t11 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X40 VIN Inverter_Layout_0.OUT.t25 VOUT.t31 VDD.t10 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X41 VOUT Inverter_Layout_0.OUT.t26 VIN.t35 VDD.t15 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X42 VOUT Inverter_Layout_0.OUT.t27 VIN.t34 VDD.t14 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X43 VOUT Inverter_Layout_0.OUT.t28 VIN.t33 VDD.t8 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X44 VOUT CLK.t15 VIN.t0 VSS.t3 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X45 VIN CLK.t16 VOUT.t1 VSS.t7 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X46 VOUT Inverter_Layout_0.OUT.t29 VIN.t32 VDD.t12 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X47 VIN CLK.t17 VOUT.t63 VSS.t2 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X48 VOUT CLK.t18 VIN.t62 VSS.t6 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X49 VIN Inverter_Layout_0.OUT.t30 VOUT.t26 VDD.t9 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X50 VIN Inverter_Layout_0.OUT.t31 VOUT.t25 VDD.t4 pfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X51 VOUT Inverter_Layout_0.OUT.t32 VIN.t31 VDD.t2 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X52 VIN CLK.t19 VOUT.t71 VSS.t0 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X53 VIN Inverter_Layout_0.OUT.t33 VOUT.t23 VDD.t0 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X54 VOUT CLK.t20 VIN.t58 VSS.t5 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X55 VIN CLK.t21 VOUT.t65 VSS.t4 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X56 VOUT Inverter_Layout_0.OUT.t34 VIN.t30 VDD.t13 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X57 VOUT Inverter_Layout_0.OUT.t35 VIN.t29 VDD.t12 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X58 VIN Inverter_Layout_0.OUT.t36 VOUT.t20 VDD.t11 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X59 VIN Inverter_Layout_0.OUT.t37 VOUT.t19 VDD.t10 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X60 VIN Inverter_Layout_0.OUT.t38 VOUT.t18 VDD.t9 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X61 VOUT Inverter_Layout_0.OUT.t39 VIN.t28 VDD.t8 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X62 VOUT CLK.t22 VIN.t8 VSS.t3 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X63 VIN Inverter_Layout_0.OUT.t40 VOUT.t16 VDD.t7 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X64 VIN CLK.t23 VOUT.t7 VSS.t2 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X65 VOUT Inverter_Layout_0.OUT.t41 VIN.t27 VDD.t6 pfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X66 VOUT Inverter_Layout_0.OUT.t42 VIN.t26 VDD.t5 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X67 VIN Inverter_Layout_0.OUT.t43 VOUT.t13 VDD.t4 pfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X68 VOUT CLK.t24 VIN.t67 VSS.t1 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X69 VIN Inverter_Layout_0.OUT.t44 VOUT.t12 VDD.t3 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X70 VOUT Inverter_Layout_0.OUT.t45 VIN.t25 VDD.t2 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X71 VIN Inverter_Layout_0.OUT.t46 VOUT.t10 VDD.t1 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X72 VIN Inverter_Layout_0.OUT.t47 VOUT.t9 VDD.t0 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X73 VIN CLK.t25 VOUT.t70 VSS.t0 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
R0 Inverter_Layout_0.OUT.t2 Inverter_Layout_0.OUT.t18 50.3184
R1 Inverter_Layout_0.OUT.t40 Inverter_Layout_0.OUT.t2 50.3184
R2 Inverter_Layout_0.OUT.t35 Inverter_Layout_0.OUT.t3 50.3184
R3 Inverter_Layout_0.OUT.t29 Inverter_Layout_0.OUT.t35 50.3184
R4 Inverter_Layout_0.OUT.t24 Inverter_Layout_0.OUT.t36 50.3184
R5 Inverter_Layout_0.OUT.t15 Inverter_Layout_0.OUT.t24 50.3184
R6 Inverter_Layout_0.OUT.t22 Inverter_Layout_0.OUT.t34 50.3184
R7 Inverter_Layout_0.OUT.t10 Inverter_Layout_0.OUT.t22 50.3184
R8 Inverter_Layout_0.OUT.t7 Inverter_Layout_0.OUT.t21 50.3184
R9 Inverter_Layout_0.OUT.t44 Inverter_Layout_0.OUT.t7 50.3184
R10 Inverter_Layout_0.OUT.t5 Inverter_Layout_0.OUT.t20 50.3184
R11 Inverter_Layout_0.OUT.t42 Inverter_Layout_0.OUT.t5 50.3184
R12 Inverter_Layout_0.OUT.t38 Inverter_Layout_0.OUT.t6 50.3184
R13 Inverter_Layout_0.OUT.t30 Inverter_Layout_0.OUT.t38 50.3184
R14 Inverter_Layout_0.OUT.t28 Inverter_Layout_0.OUT.t39 50.3184
R15 Inverter_Layout_0.OUT.t16 Inverter_Layout_0.OUT.t28 50.3184
R16 Inverter_Layout_0.OUT.t25 Inverter_Layout_0.OUT.t37 50.3184
R17 Inverter_Layout_0.OUT.t14 Inverter_Layout_0.OUT.t25 50.3184
R18 Inverter_Layout_0.OUT.t11 Inverter_Layout_0.OUT.t26 50.3184
R19 Inverter_Layout_0.OUT.t0 Inverter_Layout_0.OUT.t11 50.3184
R20 Inverter_Layout_0.OUT.t8 Inverter_Layout_0.OUT.t23 50.3184
R21 Inverter_Layout_0.OUT.t46 Inverter_Layout_0.OUT.t8 50.3184
R22 Inverter_Layout_0.OUT.t12 Inverter_Layout_0.OUT.t27 50.3184
R23 Inverter_Layout_0.OUT.t1 Inverter_Layout_0.OUT.t12 50.3184
R24 Inverter_Layout_0.OUT.t47 Inverter_Layout_0.OUT.t13 50.3184
R25 Inverter_Layout_0.OUT.t33 Inverter_Layout_0.OUT.t47 50.3184
R26 Inverter_Layout_0.OUT.t45 Inverter_Layout_0.OUT.t9 50.3184
R27 Inverter_Layout_0.OUT.t32 Inverter_Layout_0.OUT.t45 50.3184
R28 Inverter_Layout_0.OUT.t31 Inverter_Layout_0.OUT.t43 50.3184
R29 Inverter_Layout_0.OUT.t17 Inverter_Layout_0.OUT.t31 50.3184
R30 Inverter_Layout_0.OUT.t4 Inverter_Layout_0.OUT.t41 50.3184
R31 Inverter_Layout_0.OUT.t19 Inverter_Layout_0.OUT.t4 50.3184
R32 Inverter_Layout_0.OUT Inverter_Layout_0.OUT.t19 49.2314
R33 Inverter_Layout_0.OUT.n0 Inverter_Layout_0.OUT.t17 39.7594
R34 Inverter_Layout_0.OUT.t41 Inverter_Layout_0.OUT.n13 39.7594
R35 Inverter_Layout_0.OUT.n1 Inverter_Layout_0.OUT.n0 20.8576
R36 Inverter_Layout_0.OUT.n2 Inverter_Layout_0.OUT.n1 20.8576
R37 Inverter_Layout_0.OUT.n3 Inverter_Layout_0.OUT.n2 20.8576
R38 Inverter_Layout_0.OUT.n4 Inverter_Layout_0.OUT.n3 20.8576
R39 Inverter_Layout_0.OUT.n5 Inverter_Layout_0.OUT.n4 20.8576
R40 Inverter_Layout_0.OUT.n6 Inverter_Layout_0.OUT.n5 20.8576
R41 Inverter_Layout_0.OUT.n7 Inverter_Layout_0.OUT.n6 20.8576
R42 Inverter_Layout_0.OUT.n8 Inverter_Layout_0.OUT.n7 20.8576
R43 Inverter_Layout_0.OUT.n9 Inverter_Layout_0.OUT.n8 20.8576
R44 Inverter_Layout_0.OUT.n10 Inverter_Layout_0.OUT.n9 20.8576
R45 Inverter_Layout_0.OUT.n11 Inverter_Layout_0.OUT.n10 20.8576
R46 Inverter_Layout_0.OUT.n12 Inverter_Layout_0.OUT.n11 20.8576
R47 Inverter_Layout_0.OUT.n13 Inverter_Layout_0.OUT.n12 20.8576
R48 Inverter_Layout_0.OUT.n13 Inverter_Layout_0.OUT.t40 18.9023
R49 Inverter_Layout_0.OUT.n12 Inverter_Layout_0.OUT.t29 18.9023
R50 Inverter_Layout_0.OUT.n11 Inverter_Layout_0.OUT.t15 18.9023
R51 Inverter_Layout_0.OUT.n10 Inverter_Layout_0.OUT.t10 18.9023
R52 Inverter_Layout_0.OUT.n9 Inverter_Layout_0.OUT.t44 18.9023
R53 Inverter_Layout_0.OUT.n8 Inverter_Layout_0.OUT.t42 18.9023
R54 Inverter_Layout_0.OUT.n7 Inverter_Layout_0.OUT.t30 18.9023
R55 Inverter_Layout_0.OUT.n6 Inverter_Layout_0.OUT.t16 18.9023
R56 Inverter_Layout_0.OUT.n5 Inverter_Layout_0.OUT.t14 18.9023
R57 Inverter_Layout_0.OUT.n4 Inverter_Layout_0.OUT.t0 18.9023
R58 Inverter_Layout_0.OUT.n3 Inverter_Layout_0.OUT.t46 18.9023
R59 Inverter_Layout_0.OUT.n2 Inverter_Layout_0.OUT.t1 18.9023
R60 Inverter_Layout_0.OUT.n1 Inverter_Layout_0.OUT.t33 18.9023
R61 Inverter_Layout_0.OUT.n0 Inverter_Layout_0.OUT.t32 18.9023
R62 VIN.n73 VIN.n72 4.81172
R63 VIN.n104 VIN.n2 4.4609
R64 VIN.n105 VIN.n1 4.4609
R65 VIN.n106 VIN.n0 4.4609
R66 VIN.n100 VIN.t67 4.4609
R67 VIN.n101 VIN.t57 4.4609
R68 VIN.n102 VIN.t3 4.4609
R69 VIN.n95 VIN.t27 4.0565
R70 VIN.n96 VIN.t45 4.0565
R71 VIN.n97 VIN.t38 4.0565
R72 VIN.n74 VIN.n70 4.0565
R73 VIN.n73 VIN.n71 4.0565
R74 VIN.n26 VIN.n25 3.90572
R75 VIN.n9 VIN.n8 3.90572
R76 VIN.n32 VIN.n29 3.35572
R77 VIN.n46 VIN.n43 3.35572
R78 VIN.n86 VIN.n83 3.35572
R79 VIN.n63 VIN.n60 3.35572
R80 VIN.n26 VIN.n23 3.1505
R81 VIN.n27 VIN.n21 3.1505
R82 VIN.n9 VIN.n6 3.1505
R83 VIN.n10 VIN.n4 3.1505
R84 VIN.n13 VIN.n12 3.1505
R85 VIN.n16 VIN.n15 3.1505
R86 VIN.n19 VIN.n18 3.1505
R87 VIN.n32 VIN.n31 2.6005
R88 VIN.n35 VIN.n34 2.6005
R89 VIN.n46 VIN.n45 2.6005
R90 VIN.n49 VIN.n48 2.6005
R91 VIN.n50 VIN.n41 2.6005
R92 VIN.n51 VIN.n39 2.6005
R93 VIN.n52 VIN.n37 2.6005
R94 VIN.n86 VIN.n85 2.6005
R95 VIN.n89 VIN.n88 2.6005
R96 VIN.n63 VIN.n62 2.6005
R97 VIN.n66 VIN.n65 2.6005
R98 VIN.n67 VIN.n58 2.6005
R99 VIN.n68 VIN.n56 2.6005
R100 VIN.n69 VIN.n54 2.6005
R101 VIN.n90 VIN.n81 2.6005
R102 VIN.n91 VIN.n79 2.6005
R103 VIN.n92 VIN.n77 2.6005
R104 VIN.n95 VIN.n94 2.47941
R105 VIN.n103 VIN.n102 2.47941
R106 VIN.n93 VIN.n75 2.05876
R107 VIN.n34 VIN.t46 1.4565
R108 VIN.n34 VIN.n33 1.4565
R109 VIN.n31 VIN.t29 1.4565
R110 VIN.n31 VIN.n30 1.4565
R111 VIN.n29 VIN.t32 1.4565
R112 VIN.n29 VIN.n28 1.4565
R113 VIN.n37 VIN.t26 1.4565
R114 VIN.n37 VIN.n36 1.4565
R115 VIN.n39 VIN.t44 1.4565
R116 VIN.n39 VIN.n38 1.4565
R117 VIN.n41 VIN.t37 1.4565
R118 VIN.n41 VIN.n40 1.4565
R119 VIN.n48 VIN.t30 1.4565
R120 VIN.n48 VIN.n47 1.4565
R121 VIN.n45 VIN.t36 1.4565
R122 VIN.n45 VIN.n44 1.4565
R123 VIN.n43 VIN.t42 1.4565
R124 VIN.n43 VIN.n42 1.4565
R125 VIN.n77 VIN.t39 1.4565
R126 VIN.n77 VIN.n76 1.4565
R127 VIN.n79 VIN.t33 1.4565
R128 VIN.n79 VIN.n78 1.4565
R129 VIN.n81 VIN.t28 1.4565
R130 VIN.n81 VIN.n80 1.4565
R131 VIN.n88 VIN.t35 1.4565
R132 VIN.n88 VIN.n87 1.4565
R133 VIN.n85 VIN.t41 1.4565
R134 VIN.n85 VIN.n84 1.4565
R135 VIN.n83 VIN.t48 1.4565
R136 VIN.n83 VIN.n82 1.4565
R137 VIN.n54 VIN.t31 1.4565
R138 VIN.n54 VIN.n53 1.4565
R139 VIN.n56 VIN.t25 1.4565
R140 VIN.n56 VIN.n55 1.4565
R141 VIN.n58 VIN.t43 1.4565
R142 VIN.n58 VIN.n57 1.4565
R143 VIN.n65 VIN.t34 1.4565
R144 VIN.n65 VIN.n64 1.4565
R145 VIN.n62 VIN.t40 1.4565
R146 VIN.n62 VIN.n61 1.4565
R147 VIN.n60 VIN.t47 1.4565
R148 VIN.n60 VIN.n59 1.4565
R149 VIN.n21 VIN.t0 1.3109
R150 VIN.n21 VIN.n20 1.3109
R151 VIN.n23 VIN.t8 1.3109
R152 VIN.n23 VIN.n22 1.3109
R153 VIN.n25 VIN.t2 1.3109
R154 VIN.n25 VIN.n24 1.3109
R155 VIN.n18 VIN.t62 1.3109
R156 VIN.n18 VIN.n17 1.3109
R157 VIN.n15 VIN.t66 1.3109
R158 VIN.n15 VIN.n14 1.3109
R159 VIN.n12 VIN.t4 1.3109
R160 VIN.n12 VIN.n11 1.3109
R161 VIN.n4 VIN.t68 1.3109
R162 VIN.n4 VIN.n3 1.3109
R163 VIN.n6 VIN.t58 1.3109
R164 VIN.n6 VIN.n5 1.3109
R165 VIN.n8 VIN.t5 1.3109
R166 VIN.n8 VIN.n7 1.3109
R167 VIN.n50 VIN.n49 1.28789
R168 VIN.n90 VIN.n89 1.28789
R169 VIN.n67 VIN.n66 1.28789
R170 VIN.n13 VIN.n10 1.28789
R171 VIN.n75 VIN.n74 0.957239
R172 VIN.n98 VIN.n97 0.957239
R173 VIN.n99 VIN.n27 0.957239
R174 VIN.n104 VIN.n103 0.957239
R175 VIN.n99 VIN.n98 0.896587
R176 VIN.n35 VIN.n32 0.755717
R177 VIN.n49 VIN.n46 0.755717
R178 VIN.n52 VIN.n51 0.755717
R179 VIN.n51 VIN.n50 0.755717
R180 VIN.n89 VIN.n86 0.755717
R181 VIN.n66 VIN.n63 0.755717
R182 VIN.n69 VIN.n68 0.755717
R183 VIN.n68 VIN.n67 0.755717
R184 VIN.n74 VIN.n73 0.755717
R185 VIN.n92 VIN.n91 0.755717
R186 VIN.n91 VIN.n90 0.755717
R187 VIN.n96 VIN.n95 0.755717
R188 VIN.n97 VIN.n96 0.755717
R189 VIN.n27 VIN.n26 0.755717
R190 VIN.n101 VIN.n100 0.755717
R191 VIN.n102 VIN.n101 0.755717
R192 VIN.n10 VIN.n9 0.755717
R193 VIN.n16 VIN.n13 0.755717
R194 VIN.n19 VIN.n16 0.755717
R195 VIN.n106 VIN.n105 0.755717
R196 VIN.n105 VIN.n104 0.755717
R197 VIN.n94 VIN.n93 0.626587
R198 VIN VIN.n106 0.513109
R199 VIN.n98 VIN.n35 0.331152
R200 VIN.n94 VIN.n52 0.331152
R201 VIN.n75 VIN.n69 0.331152
R202 VIN.n93 VIN.n92 0.331152
R203 VIN.n100 VIN.n99 0.331152
R204 VIN.n103 VIN.n19 0.331152
R205 VOUT.n40 VOUT.n39 3.90572
R206 VOUT.n60 VOUT.n57 3.90572
R207 VOUT.n68 VOUT.n65 3.90572
R208 VOUT.n4 VOUT.n1 3.35572
R209 VOUT.n22 VOUT.n21 3.35572
R210 VOUT.n14 VOUT.n13 3.35572
R211 VOUT.n46 VOUT.n43 3.35572
R212 VOUT.n90 VOUT.n89 3.35572
R213 VOUT.n82 VOUT.n81 3.35572
R214 VOUT.n40 VOUT.n37 3.1505
R215 VOUT.n41 VOUT.n35 3.1505
R216 VOUT.n60 VOUT.n59 3.1505
R217 VOUT.n63 VOUT.n62 3.1505
R218 VOUT.n68 VOUT.n67 3.1505
R219 VOUT.n71 VOUT.n70 3.1505
R220 VOUT.n73 VOUT.n55 3.1505
R221 VOUT.n74 VOUT.n53 3.1505
R222 VOUT.n75 VOUT.n51 3.1505
R223 VOUT.n4 VOUT.n3 2.6005
R224 VOUT.n7 VOUT.n6 2.6005
R225 VOUT.n22 VOUT.n19 2.6005
R226 VOUT.n23 VOUT.n17 2.6005
R227 VOUT.n14 VOUT.n11 2.6005
R228 VOUT.n15 VOUT.n9 2.6005
R229 VOUT.n27 VOUT.n26 2.6005
R230 VOUT.n30 VOUT.n29 2.6005
R231 VOUT.n33 VOUT.n32 2.6005
R232 VOUT.n46 VOUT.n45 2.6005
R233 VOUT.n49 VOUT.n48 2.6005
R234 VOUT.n90 VOUT.n87 2.6005
R235 VOUT.n91 VOUT.n85 2.6005
R236 VOUT.n82 VOUT.n79 2.6005
R237 VOUT.n83 VOUT.n77 2.6005
R238 VOUT.n101 VOUT.n100 2.6005
R239 VOUT.n98 VOUT.n97 2.6005
R240 VOUT.n95 VOUT.n94 2.6005
R241 VOUT.n102 VOUT.n101 1.76333
R242 VOUT.n6 VOUT.t13 1.4565
R243 VOUT.n6 VOUT.n5 1.4565
R244 VOUT.n3 VOUT.t25 1.4565
R245 VOUT.n3 VOUT.n2 1.4565
R246 VOUT.n1 VOUT.t39 1.4565
R247 VOUT.n1 VOUT.n0 1.4565
R248 VOUT.n32 VOUT.t33 1.4565
R249 VOUT.n32 VOUT.n31 1.4565
R250 VOUT.n29 VOUT.t48 1.4565
R251 VOUT.n29 VOUT.n28 1.4565
R252 VOUT.n26 VOUT.t10 1.4565
R253 VOUT.n26 VOUT.n25 1.4565
R254 VOUT.n17 VOUT.t42 1.4565
R255 VOUT.n17 VOUT.n16 1.4565
R256 VOUT.n19 VOUT.t31 1.4565
R257 VOUT.n19 VOUT.n18 1.4565
R258 VOUT.n21 VOUT.t19 1.4565
R259 VOUT.n21 VOUT.n20 1.4565
R260 VOUT.n9 VOUT.t23 1.4565
R261 VOUT.n9 VOUT.n8 1.4565
R262 VOUT.n11 VOUT.t9 1.4565
R263 VOUT.n11 VOUT.n10 1.4565
R264 VOUT.n13 VOUT.t43 1.4565
R265 VOUT.n13 VOUT.n12 1.4565
R266 VOUT.n48 VOUT.t50 1.4565
R267 VOUT.n48 VOUT.n47 1.4565
R268 VOUT.n45 VOUT.t18 1.4565
R269 VOUT.n45 VOUT.n44 1.4565
R270 VOUT.n43 VOUT.t26 1.4565
R271 VOUT.n43 VOUT.n42 1.4565
R272 VOUT.n94 VOUT.t41 1.4565
R273 VOUT.n94 VOUT.n93 1.4565
R274 VOUT.n97 VOUT.t32 1.4565
R275 VOUT.n97 VOUT.n96 1.4565
R276 VOUT.n100 VOUT.t20 1.4565
R277 VOUT.n100 VOUT.n99 1.4565
R278 VOUT.n85 VOUT.t16 1.4565
R279 VOUT.n85 VOUT.n84 1.4565
R280 VOUT.n87 VOUT.t54 1.4565
R281 VOUT.n87 VOUT.n86 1.4565
R282 VOUT.n89 VOUT.t38 1.4565
R283 VOUT.n89 VOUT.n88 1.4565
R284 VOUT.n77 VOUT.t12 1.4565
R285 VOUT.n77 VOUT.n76 1.4565
R286 VOUT.n79 VOUT.t49 1.4565
R287 VOUT.n79 VOUT.n78 1.4565
R288 VOUT.n81 VOUT.t35 1.4565
R289 VOUT.n81 VOUT.n80 1.4565
R290 VOUT.n35 VOUT.t61 1.3109
R291 VOUT.n35 VOUT.n34 1.3109
R292 VOUT.n37 VOUT.t64 1.3109
R293 VOUT.n37 VOUT.n36 1.3109
R294 VOUT.n39 VOUT.t65 1.3109
R295 VOUT.n39 VOUT.n38 1.3109
R296 VOUT.n51 VOUT.t59 1.3109
R297 VOUT.n51 VOUT.n50 1.3109
R298 VOUT.n53 VOUT.t60 1.3109
R299 VOUT.n53 VOUT.n52 1.3109
R300 VOUT.n55 VOUT.t1 1.3109
R301 VOUT.n55 VOUT.n54 1.3109
R302 VOUT.n62 VOUT.t6 1.3109
R303 VOUT.n62 VOUT.n61 1.3109
R304 VOUT.n59 VOUT.t7 1.3109
R305 VOUT.n59 VOUT.n58 1.3109
R306 VOUT.n57 VOUT.t63 1.3109
R307 VOUT.n57 VOUT.n56 1.3109
R308 VOUT.n70 VOUT.t70 1.3109
R309 VOUT.n70 VOUT.n69 1.3109
R310 VOUT.n67 VOUT.t71 1.3109
R311 VOUT.n67 VOUT.n66 1.3109
R312 VOUT.n65 VOUT.t69 1.3109
R313 VOUT.n65 VOUT.n64 1.3109
R314 VOUT.n104 VOUT.n103 1.25267
R315 VOUT.n103 VOUT.n102 1.25267
R316 VOUT.n24 VOUT.n23 0.957239
R317 VOUT.n24 VOUT.n15 0.957239
R318 VOUT.n72 VOUT.n63 0.957239
R319 VOUT.n72 VOUT.n71 0.957239
R320 VOUT.n92 VOUT.n91 0.957239
R321 VOUT.n92 VOUT.n83 0.957239
R322 VOUT.n7 VOUT.n4 0.755717
R323 VOUT.n23 VOUT.n22 0.755717
R324 VOUT.n15 VOUT.n14 0.755717
R325 VOUT.n30 VOUT.n27 0.755717
R326 VOUT.n33 VOUT.n30 0.755717
R327 VOUT.n41 VOUT.n40 0.755717
R328 VOUT.n63 VOUT.n60 0.755717
R329 VOUT.n71 VOUT.n68 0.755717
R330 VOUT.n49 VOUT.n46 0.755717
R331 VOUT.n75 VOUT.n74 0.755717
R332 VOUT.n74 VOUT.n73 0.755717
R333 VOUT.n91 VOUT.n90 0.755717
R334 VOUT.n83 VOUT.n82 0.755717
R335 VOUT.n98 VOUT.n95 0.755717
R336 VOUT.n101 VOUT.n98 0.755717
R337 VOUT.n104 VOUT.n7 0.511152
R338 VOUT.n103 VOUT.n33 0.511152
R339 VOUT.n103 VOUT.n41 0.511152
R340 VOUT.n102 VOUT.n49 0.511152
R341 VOUT.n102 VOUT.n75 0.511152
R342 VOUT.n27 VOUT.n24 0.331152
R343 VOUT.n73 VOUT.n72 0.331152
R344 VOUT.n95 VOUT.n92 0.331152
R345 VOUT VOUT.n104 0.0885435
R346 VDD.n5 VDD.n0 577.115
R347 VDD.n5 VDD.t16 409.62
R348 VDD.t2 VDD.t4 124.805
R349 VDD.t0 VDD.t2 124.805
R350 VDD.t14 VDD.t0 124.805
R351 VDD.t1 VDD.t14 124.805
R352 VDD.t15 VDD.t1 124.805
R353 VDD.t10 VDD.t15 124.805
R354 VDD.t8 VDD.t10 124.805
R355 VDD.t9 VDD.t8 124.805
R356 VDD.t5 VDD.t9 124.805
R357 VDD.t3 VDD.t5 124.805
R358 VDD.t13 VDD.t3 124.805
R359 VDD.t11 VDD.t13 124.805
R360 VDD.t12 VDD.t11 124.805
R361 VDD.t7 VDD.t12 124.805
R362 VDD.n0 VDD.t6 77.2236
R363 VDD.n0 VDD.t7 47.5824
R364 VDD.n4 VDD.n3 4.98375
R365 VDD.n3 VDD.n2 4.7942
R366 VDD.n1 VDD 3.1505
R367 VDD.n4 VDD.n1 1.78473
R368 VDD VDD.n6 1.62573
R369 VDD.n6 VDD.n5 1.58353
R370 VDD.n5 VDD.n4 0.684132
R371 VDD.n3 VDD 0.0270179
R372 CLK.t13 CLK.t6 50.3184
R373 CLK.t21 CLK.t13 50.3184
R374 CLK.t9 CLK.t1 50.3184
R375 CLK.t18 CLK.t9 50.3184
R376 CLK.t23 CLK.t17 50.3184
R377 CLK.t5 CLK.t23 50.3184
R378 CLK.t20 CLK.t11 50.3184
R379 CLK.t2 CLK.t20 50.3184
R380 CLK.t8 CLK.t0 50.3184
R381 CLK.t16 CLK.t8 50.3184
R382 CLK.t22 CLK.t15 50.3184
R383 CLK.t4 CLK.t22 50.3184
R384 CLK.t19 CLK.t10 50.3184
R385 CLK.t25 CLK.t19 50.3184
R386 CLK.t7 CLK.t24 50.3184
R387 CLK.t14 CLK.t7 50.3184
R388 CLK CLK.n6 48.0321
R389 CLK.n0 CLK.t21 39.7594
R390 CLK.n7 CLK.t12 34.6755
R391 CLK.n1 CLK.n0 20.8576
R392 CLK.n2 CLK.n1 20.8576
R393 CLK.n3 CLK.n2 20.8576
R394 CLK.n4 CLK.n3 20.8576
R395 CLK.n5 CLK.n4 20.8576
R396 CLK.n6 CLK.n5 20.8576
R397 CLK.n0 CLK.t18 18.9023
R398 CLK.n1 CLK.t5 18.9023
R399 CLK.n2 CLK.t2 18.9023
R400 CLK.n3 CLK.t16 18.9023
R401 CLK.n4 CLK.t4 18.9023
R402 CLK.n5 CLK.t25 18.9023
R403 CLK.n6 CLK.t14 18.9023
R404 CLK CLK.n7 17.6692
R405 CLK.n7 CLK.t3 13.0362
R406 VSS.n2 VSS.t1 558.01
R407 VSS.n3 VSS.n2 506.635
R408 VSS.n2 VSS.t8 495.854
R409 VSS.t6 VSS.t4 373.563
R410 VSS.t2 VSS.t6 373.563
R411 VSS.t5 VSS.t2 373.563
R412 VSS.t7 VSS.t5 373.563
R413 VSS.t3 VSS.t7 373.563
R414 VSS.t0 VSS.t3 373.563
R415 VSS.t1 VSS.t0 373.563
R416 VSS.n1 VSS.n0 6.68085
R417 VSS VSS.n6 2.67604
R418 VSS VSS.n5 2.6005
R419 VSS.n5 VSS.n4 1.65811
R420 VSS.n4 VSS.n3 0.472445
R421 VSS VSS.n1 0.0647857
C0 VDD CLK 0.198f
C1 VOUT VIN 15.9f
C2 Inverter_Layout_0.OUT VOUT 0.623f
C3 Inverter_Layout_0.OUT VIN 0.755f
C4 VOUT CLK 0.318f
C5 VDD VOUT 0.379f
C6 VIN CLK 0.543f
C7 Inverter_Layout_0.OUT CLK 0.0739f
C8 VDD VIN 0.722f
C9 Inverter_Layout_0.OUT VDD 4.02f
C10 VOUT VSS 1.1f
C11 VIN VSS 2.77f
C12 CLK VSS 3.37f
C13 Inverter_Layout_0.OUT VSS 2.63f
C14 VDD VSS 12.3f
C15 VDD.t4 VSS 0.345f
C16 VDD.t2 VSS 0.196f
C17 VDD.t0 VSS 0.196f
C18 VDD.t14 VSS 0.196f
C19 VDD.t1 VSS 0.196f
C20 VDD.t15 VSS 0.196f
C21 VDD.t10 VSS 0.196f
C22 VDD.t8 VSS 0.196f
C23 VDD.t9 VSS 0.196f
C24 VDD.t5 VSS 0.196f
C25 VDD.t3 VSS 0.196f
C26 VDD.t13 VSS 0.196f
C27 VDD.t11 VSS 0.196f
C28 VDD.t12 VSS 0.196f
C29 VDD.t7 VSS 0.135f
C30 VDD.t6 VSS 0.308f
C31 VDD.n0 VSS 0.198f
C32 VDD.t16 VSS 0.203f
C33 VDD.n1 VSS 0.00687f
C34 VDD.n2 VSS 0.013f
C35 VDD.n3 VSS 0.0332f
C36 VDD.n4 VSS 0.00376f
C37 VDD.n5 VSS 0.173f
C38 VDD.n6 VSS 0.00819f
C39 VOUT.t39 VSS 0.0592f
C40 VOUT.n0 VSS 0.0592f
C41 VOUT.n1 VSS 0.148f
C42 VOUT.t25 VSS 0.0592f
C43 VOUT.n2 VSS 0.0592f
C44 VOUT.n3 VSS 0.118f
C45 VOUT.n4 VSS 0.264f
C46 VOUT.t13 VSS 0.0592f
C47 VOUT.n5 VSS 0.0592f
C48 VOUT.n6 VSS 0.118f
C49 VOUT.n7 VSS 0.136f
C50 VOUT.t23 VSS 0.0592f
C51 VOUT.n8 VSS 0.0592f
C52 VOUT.n9 VSS 0.118f
C53 VOUT.t9 VSS 0.0592f
C54 VOUT.n10 VSS 0.0592f
C55 VOUT.n11 VSS 0.118f
C56 VOUT.t43 VSS 0.0592f
C57 VOUT.n12 VSS 0.0592f
C58 VOUT.n13 VSS 0.148f
C59 VOUT.n14 VSS 0.264f
C60 VOUT.n15 VSS 0.19f
C61 VOUT.t42 VSS 0.0592f
C62 VOUT.n16 VSS 0.0592f
C63 VOUT.n17 VSS 0.118f
C64 VOUT.t31 VSS 0.0592f
C65 VOUT.n18 VSS 0.0592f
C66 VOUT.n19 VSS 0.118f
C67 VOUT.t19 VSS 0.0592f
C68 VOUT.n20 VSS 0.0592f
C69 VOUT.n21 VSS 0.148f
C70 VOUT.n22 VSS 0.264f
C71 VOUT.n23 VSS 0.19f
C72 VOUT.n24 VSS 0.247f
C73 VOUT.t10 VSS 0.0592f
C74 VOUT.n25 VSS 0.0592f
C75 VOUT.n26 VSS 0.118f
C76 VOUT.n27 VSS 0.116f
C77 VOUT.t48 VSS 0.0592f
C78 VOUT.n28 VSS 0.0592f
C79 VOUT.n29 VSS 0.118f
C80 VOUT.n30 VSS 0.162f
C81 VOUT.t33 VSS 0.0592f
C82 VOUT.n31 VSS 0.0592f
C83 VOUT.n32 VSS 0.118f
C84 VOUT.n33 VSS 0.136f
C85 VOUT.t61 VSS 0.0592f
C86 VOUT.n34 VSS 0.0592f
C87 VOUT.n35 VSS 0.118f
C88 VOUT.t64 VSS 0.0592f
C89 VOUT.n36 VSS 0.0592f
C90 VOUT.n37 VSS 0.118f
C91 VOUT.t65 VSS 0.0592f
C92 VOUT.n38 VSS 0.0592f
C93 VOUT.n39 VSS 0.144f
C94 VOUT.n40 VSS 0.269f
C95 VOUT.n41 VSS 0.136f
C96 VOUT.t26 VSS 0.0592f
C97 VOUT.n42 VSS 0.0592f
C98 VOUT.n43 VSS 0.148f
C99 VOUT.t18 VSS 0.0592f
C100 VOUT.n44 VSS 0.0592f
C101 VOUT.n45 VSS 0.118f
C102 VOUT.n46 VSS 0.264f
C103 VOUT.t50 VSS 0.0592f
C104 VOUT.n47 VSS 0.0592f
C105 VOUT.n48 VSS 0.118f
C106 VOUT.n49 VSS 0.136f
C107 VOUT.t59 VSS 0.0592f
C108 VOUT.n50 VSS 0.0592f
C109 VOUT.n51 VSS 0.118f
C110 VOUT.t60 VSS 0.0592f
C111 VOUT.n52 VSS 0.0592f
C112 VOUT.n53 VSS 0.118f
C113 VOUT.t1 VSS 0.0592f
C114 VOUT.n54 VSS 0.0592f
C115 VOUT.n55 VSS 0.118f
C116 VOUT.t63 VSS 0.0592f
C117 VOUT.n56 VSS 0.0592f
C118 VOUT.n57 VSS 0.144f
C119 VOUT.t7 VSS 0.0592f
C120 VOUT.n58 VSS 0.0592f
C121 VOUT.n59 VSS 0.118f
C122 VOUT.n60 VSS 0.269f
C123 VOUT.t6 VSS 0.0592f
C124 VOUT.n61 VSS 0.0592f
C125 VOUT.n62 VSS 0.118f
C126 VOUT.n63 VSS 0.19f
C127 VOUT.t69 VSS 0.0592f
C128 VOUT.n64 VSS 0.0592f
C129 VOUT.n65 VSS 0.144f
C130 VOUT.t71 VSS 0.0592f
C131 VOUT.n66 VSS 0.0592f
C132 VOUT.n67 VSS 0.118f
C133 VOUT.n68 VSS 0.269f
C134 VOUT.t70 VSS 0.0592f
C135 VOUT.n69 VSS 0.0592f
C136 VOUT.n70 VSS 0.118f
C137 VOUT.n71 VSS 0.19f
C138 VOUT.n72 VSS 0.247f
C139 VOUT.n73 VSS 0.116f
C140 VOUT.n74 VSS 0.162f
C141 VOUT.n75 VSS 0.136f
C142 VOUT.t12 VSS 0.0592f
C143 VOUT.n76 VSS 0.0592f
C144 VOUT.n77 VSS 0.118f
C145 VOUT.t49 VSS 0.0592f
C146 VOUT.n78 VSS 0.0592f
C147 VOUT.n79 VSS 0.118f
C148 VOUT.t35 VSS 0.0592f
C149 VOUT.n80 VSS 0.0592f
C150 VOUT.n81 VSS 0.148f
C151 VOUT.n82 VSS 0.264f
C152 VOUT.n83 VSS 0.19f
C153 VOUT.t16 VSS 0.0592f
C154 VOUT.n84 VSS 0.0592f
C155 VOUT.n85 VSS 0.118f
C156 VOUT.t54 VSS 0.0592f
C157 VOUT.n86 VSS 0.0592f
C158 VOUT.n87 VSS 0.118f
C159 VOUT.t38 VSS 0.0592f
C160 VOUT.n88 VSS 0.0592f
C161 VOUT.n89 VSS 0.148f
C162 VOUT.n90 VSS 0.264f
C163 VOUT.n91 VSS 0.19f
C164 VOUT.n92 VSS 0.247f
C165 VOUT.t41 VSS 0.0592f
C166 VOUT.n93 VSS 0.0592f
C167 VOUT.n94 VSS 0.118f
C168 VOUT.n95 VSS 0.116f
C169 VOUT.t32 VSS 0.0592f
C170 VOUT.n96 VSS 0.0592f
C171 VOUT.n97 VSS 0.118f
C172 VOUT.n98 VSS 0.162f
C173 VOUT.t20 VSS 0.0592f
C174 VOUT.n99 VSS 0.0592f
C175 VOUT.n100 VSS 0.118f
C176 VOUT.n101 VSS 0.277f
C177 VOUT.n102 VSS 0.435f
C178 VOUT.n103 VSS 0.378f
C179 VOUT.n104 VSS 0.198f
C180 VIN.n0 VSS 0.133f
C181 VIN.n1 VSS 0.133f
C182 VIN.n2 VSS 0.133f
C183 VIN.t68 VSS 0.0496f
C184 VIN.n3 VSS 0.0496f
C185 VIN.n4 VSS 0.0993f
C186 VIN.t58 VSS 0.0496f
C187 VIN.n5 VSS 0.0496f
C188 VIN.n6 VSS 0.0993f
C189 VIN.t5 VSS 0.0496f
C190 VIN.n7 VSS 0.0496f
C191 VIN.n8 VSS 0.121f
C192 VIN.n9 VSS 0.225f
C193 VIN.n10 VSS 0.191f
C194 VIN.t4 VSS 0.0496f
C195 VIN.n11 VSS 0.0496f
C196 VIN.n12 VSS 0.0993f
C197 VIN.n13 VSS 0.191f
C198 VIN.t66 VSS 0.0496f
C199 VIN.n14 VSS 0.0496f
C200 VIN.n15 VSS 0.0993f
C201 VIN.n16 VSS 0.136f
C202 VIN.t62 VSS 0.0496f
C203 VIN.n17 VSS 0.0496f
C204 VIN.n18 VSS 0.0993f
C205 VIN.n19 VSS 0.0975f
C206 VIN.t0 VSS 0.0496f
C207 VIN.n20 VSS 0.0496f
C208 VIN.n21 VSS 0.0993f
C209 VIN.t8 VSS 0.0496f
C210 VIN.n22 VSS 0.0496f
C211 VIN.n23 VSS 0.0993f
C212 VIN.t2 VSS 0.0496f
C213 VIN.n24 VSS 0.0496f
C214 VIN.n25 VSS 0.121f
C215 VIN.n26 VSS 0.225f
C216 VIN.n27 VSS 0.159f
C217 VIN.t32 VSS 0.0496f
C218 VIN.n28 VSS 0.0496f
C219 VIN.n29 VSS 0.124f
C220 VIN.t29 VSS 0.0496f
C221 VIN.n30 VSS 0.0496f
C222 VIN.n31 VSS 0.0993f
C223 VIN.n32 VSS 0.222f
C224 VIN.t46 VSS 0.0496f
C225 VIN.n33 VSS 0.0496f
C226 VIN.n34 VSS 0.0993f
C227 VIN.n35 VSS 0.0975f
C228 VIN.t26 VSS 0.0496f
C229 VIN.n36 VSS 0.0496f
C230 VIN.n37 VSS 0.0993f
C231 VIN.t44 VSS 0.0496f
C232 VIN.n38 VSS 0.0496f
C233 VIN.n39 VSS 0.0993f
C234 VIN.t37 VSS 0.0496f
C235 VIN.n40 VSS 0.0496f
C236 VIN.n41 VSS 0.0993f
C237 VIN.t42 VSS 0.0496f
C238 VIN.n42 VSS 0.0496f
C239 VIN.n43 VSS 0.124f
C240 VIN.t36 VSS 0.0496f
C241 VIN.n44 VSS 0.0496f
C242 VIN.n45 VSS 0.0993f
C243 VIN.n46 VSS 0.222f
C244 VIN.t30 VSS 0.0496f
C245 VIN.n47 VSS 0.0496f
C246 VIN.n48 VSS 0.0993f
C247 VIN.n49 VSS 0.191f
C248 VIN.n50 VSS 0.191f
C249 VIN.n51 VSS 0.136f
C250 VIN.n52 VSS 0.0975f
C251 VIN.t31 VSS 0.0496f
C252 VIN.n53 VSS 0.0496f
C253 VIN.n54 VSS 0.0993f
C254 VIN.t25 VSS 0.0496f
C255 VIN.n55 VSS 0.0496f
C256 VIN.n56 VSS 0.0993f
C257 VIN.t43 VSS 0.0496f
C258 VIN.n57 VSS 0.0496f
C259 VIN.n58 VSS 0.0993f
C260 VIN.t47 VSS 0.0496f
C261 VIN.n59 VSS 0.0496f
C262 VIN.n60 VSS 0.124f
C263 VIN.t40 VSS 0.0496f
C264 VIN.n61 VSS 0.0496f
C265 VIN.n62 VSS 0.0993f
C266 VIN.n63 VSS 0.222f
C267 VIN.t34 VSS 0.0496f
C268 VIN.n64 VSS 0.0496f
C269 VIN.n65 VSS 0.0993f
C270 VIN.n66 VSS 0.192f
C271 VIN.n67 VSS 0.192f
C272 VIN.n68 VSS 0.136f
C273 VIN.n69 VSS 0.0975f
C274 VIN.n70 VSS 0.126f
C275 VIN.n71 VSS 0.126f
C276 VIN.n72 VSS 0.15f
C277 VIN.n73 VSS 0.307f
C278 VIN.n74 VSS 0.201f
C279 VIN.n75 VSS 0.319f
C280 VIN.t39 VSS 0.0496f
C281 VIN.n76 VSS 0.0496f
C282 VIN.n77 VSS 0.0993f
C283 VIN.t33 VSS 0.0496f
C284 VIN.n78 VSS 0.0496f
C285 VIN.n79 VSS 0.0993f
C286 VIN.t28 VSS 0.0496f
C287 VIN.n80 VSS 0.0496f
C288 VIN.n81 VSS 0.0993f
C289 VIN.t48 VSS 0.0496f
C290 VIN.n82 VSS 0.0496f
C291 VIN.n83 VSS 0.124f
C292 VIN.t41 VSS 0.0496f
C293 VIN.n84 VSS 0.0496f
C294 VIN.n85 VSS 0.0993f
C295 VIN.n86 VSS 0.222f
C296 VIN.t35 VSS 0.0496f
C297 VIN.n87 VSS 0.0496f
C298 VIN.n88 VSS 0.0993f
C299 VIN.n89 VSS 0.191f
C300 VIN.n90 VSS 0.191f
C301 VIN.n91 VSS 0.136f
C302 VIN.n92 VSS 0.0975f
C303 VIN.n93 VSS 0.287f
C304 VIN.n94 VSS 0.326f
C305 VIN.t27 VSS 0.126f
C306 VIN.n95 VSS 0.34f
C307 VIN.t45 VSS 0.126f
C308 VIN.n96 VSS 0.178f
C309 VIN.t38 VSS 0.126f
C310 VIN.n97 VSS 0.201f
C311 VIN.n98 VSS 0.213f
C312 VIN.n99 VSS 0.201f
C313 VIN.t67 VSS 0.133f
C314 VIN.n100 VSS 0.132f
C315 VIN.t57 VSS 0.133f
C316 VIN.n101 VSS 0.17f
C317 VIN.t3 VSS 0.133f
C318 VIN.n102 VSS 0.332f
C319 VIN.n103 VSS 0.358f
C320 VIN.n104 VSS 0.194f
C321 VIN.n105 VSS 0.17f
C322 VIN.n106 VSS 0.152f
C323 Inverter_Layout_0.OUT.t18 VSS 0.0535f
C324 Inverter_Layout_0.OUT.t2 VSS 0.0754f
C325 Inverter_Layout_0.OUT.t40 VSS 0.0518f
C326 Inverter_Layout_0.OUT.t3 VSS 0.0535f
C327 Inverter_Layout_0.OUT.t35 VSS 0.0754f
C328 Inverter_Layout_0.OUT.t29 VSS 0.0518f
C329 Inverter_Layout_0.OUT.t36 VSS 0.0535f
C330 Inverter_Layout_0.OUT.t24 VSS 0.0754f
C331 Inverter_Layout_0.OUT.t15 VSS 0.0518f
C332 Inverter_Layout_0.OUT.t34 VSS 0.0535f
C333 Inverter_Layout_0.OUT.t22 VSS 0.0754f
C334 Inverter_Layout_0.OUT.t10 VSS 0.0518f
C335 Inverter_Layout_0.OUT.t21 VSS 0.0535f
C336 Inverter_Layout_0.OUT.t7 VSS 0.0754f
C337 Inverter_Layout_0.OUT.t44 VSS 0.0518f
C338 Inverter_Layout_0.OUT.t20 VSS 0.0535f
C339 Inverter_Layout_0.OUT.t5 VSS 0.0754f
C340 Inverter_Layout_0.OUT.t42 VSS 0.0518f
C341 Inverter_Layout_0.OUT.t6 VSS 0.0535f
C342 Inverter_Layout_0.OUT.t38 VSS 0.0754f
C343 Inverter_Layout_0.OUT.t30 VSS 0.0518f
C344 Inverter_Layout_0.OUT.t39 VSS 0.0535f
C345 Inverter_Layout_0.OUT.t28 VSS 0.0754f
C346 Inverter_Layout_0.OUT.t16 VSS 0.0518f
C347 Inverter_Layout_0.OUT.t37 VSS 0.0535f
C348 Inverter_Layout_0.OUT.t25 VSS 0.0754f
C349 Inverter_Layout_0.OUT.t14 VSS 0.0518f
C350 Inverter_Layout_0.OUT.t26 VSS 0.0535f
C351 Inverter_Layout_0.OUT.t11 VSS 0.0754f
C352 Inverter_Layout_0.OUT.t0 VSS 0.0518f
C353 Inverter_Layout_0.OUT.t23 VSS 0.0535f
C354 Inverter_Layout_0.OUT.t8 VSS 0.0754f
C355 Inverter_Layout_0.OUT.t46 VSS 0.0518f
C356 Inverter_Layout_0.OUT.t27 VSS 0.0535f
C357 Inverter_Layout_0.OUT.t12 VSS 0.0754f
C358 Inverter_Layout_0.OUT.t1 VSS 0.0518f
C359 Inverter_Layout_0.OUT.t13 VSS 0.0535f
C360 Inverter_Layout_0.OUT.t47 VSS 0.0754f
C361 Inverter_Layout_0.OUT.t33 VSS 0.0518f
C362 Inverter_Layout_0.OUT.t9 VSS 0.0535f
C363 Inverter_Layout_0.OUT.t45 VSS 0.0754f
C364 Inverter_Layout_0.OUT.t32 VSS 0.0518f
C365 Inverter_Layout_0.OUT.t43 VSS 0.0535f
C366 Inverter_Layout_0.OUT.t31 VSS 0.0754f
C367 Inverter_Layout_0.OUT.t17 VSS 0.0703f
C368 Inverter_Layout_0.OUT.n0 VSS 0.0622f
C369 Inverter_Layout_0.OUT.n1 VSS 0.0454f
C370 Inverter_Layout_0.OUT.n2 VSS 0.0454f
C371 Inverter_Layout_0.OUT.n3 VSS 0.0454f
C372 Inverter_Layout_0.OUT.n4 VSS 0.0454f
C373 Inverter_Layout_0.OUT.n5 VSS 0.0454f
C374 Inverter_Layout_0.OUT.n6 VSS 0.0454f
C375 Inverter_Layout_0.OUT.n7 VSS 0.0454f
C376 Inverter_Layout_0.OUT.n8 VSS 0.0454f
C377 Inverter_Layout_0.OUT.n9 VSS 0.0454f
C378 Inverter_Layout_0.OUT.n10 VSS 0.0454f
C379 Inverter_Layout_0.OUT.n11 VSS 0.0454f
C380 Inverter_Layout_0.OUT.n12 VSS 0.0454f
C381 Inverter_Layout_0.OUT.n13 VSS 0.0622f
C382 Inverter_Layout_0.OUT.t41 VSS 0.0703f
C383 Inverter_Layout_0.OUT.t4 VSS 0.0754f
C384 Inverter_Layout_0.OUT.t19 VSS 0.0783f
.ends

