magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2045 -2797 2045 2797
<< psubdiff >>
rect -45 775 45 797
rect -45 -775 -23 775
rect 23 -775 45 775
rect -45 -797 45 -775
<< psubdiffcont >>
rect -23 -775 23 775
<< metal1 >>
rect -34 775 34 786
rect -34 -775 -23 775
rect 23 -775 34 775
rect -34 -786 34 -775
<< end >>
