* NGSPICE file created from mux_2x1_flat.ext - technology: gf180mcuC

.subckt mux_2x1_flat I0 I1 VDD VSS OUT Sel
X0 nand2_2.OUT I0.t0 a_801_n344# VSS.t0 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1 nand2_1.IN2 Sel.t0 a_238_256# VSS.t6 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2 VDD I0.t1 nand2_2.OUT VDD.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3 OUT nand2_1.IN2 VDD.t4 VDD.t3 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X4 a_801_n344# nand2_2.IN2 VSS.t5 VSS.t1 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X5 nand2_2.IN2 Sel.t1 VSS.t4 VSS.t3 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X6 nand2_2.OUT nand2_2.IN2 VDD.t6 VDD.t5 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X7 nand2_1.IN2 I1.t0 VDD.t16 VDD.t15 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X8 a_801_256# nand2_1.IN2 VSS.t2 VSS.t1 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X9 nand2_2.IN2 Sel.t2 VDD.t14 VDD.t13 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X10 VDD nand2_2.OUT OUT.t2 VDD.t7 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X11 a_238_256# I1.t1 VSS.t8 VSS.t7 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X12 VDD Sel.t3 nand2_1.IN2 VDD.t10 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X13 OUT nand2_2.OUT a_801_256# VSS.t0 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
R0 I0.n0 I0.t0 31.528
R1 I0.n0 I0.t1 15.3826
R2 I0.n1 I0.n0 8.74076
R3 I0 I0.n1 0.116779
R4 I0.n1 I0 0.00355085
R5 VSS.t6 VSS.t1 1483.3
R6 VSS.n3 VSS.t0 353.341
R7 VSS.t1 VSS.n3 235.561
R8 VSS.n5 VSS.t7 235.561
R9 VSS.n0 VSS.t4 9.34566
R10 VSS VSS.t8 7.24801
R11 VSS.n2 VSS.t2 7.19156
R12 VSS.n2 VSS.t5 7.19156
R13 VSS.t3 VSS.t6 3.68113
R14 VSS.n6 VSS.n4 3.37613
R15 VSS.n3 VSS 2.60269
R16 VSS VSS.n6 2.6005
R17 VSS.n6 VSS.n5 2.6005
R18 VSS.n4 VSS.n1 2.6005
R19 VSS.n4 VSS.t3 2.6005
R20 VSS.n2 VSS 0.117596
R21 VSS VSS.n2 0.0595367
R22 VSS VSS.n0 0.0340526
R23 VSS VSS.n1 0.0139211
R24 VSS VSS.n0 0.00405263
R25 VSS.n1 VSS 0.000894737
R26 Sel.n2 Sel.t0 31.528
R27 Sel.n1 Sel.t2 25.7638
R28 Sel.n2 Sel.t3 15.3826
R29 Sel.n1 Sel.t1 13.2969
R30 Sel.n3 Sel.n2 7.62851
R31 Sel.n4 Sel.n0 4.52555
R32 Sel.n4 Sel.n3 2.2324
R33 Sel.n5 Sel.n1 2.11815
R34 Sel.n5 Sel 1.13555
R35 Sel.n3 Sel 0.107918
R36 Sel Sel.n4 0.0252959
R37 Sel Sel.n0 0.00328351
R38 Sel Sel.n5 0.00142783
R39 VDD.t10 VDD.t3 763.259
R40 VDD.n12 VDD.t5 386.348
R41 VDD.n12 VDD.t13 362.409
R42 VDD.n13 VDD.n12 319.75
R43 VDD.n1 VDD.t0 193.183
R44 VDD.n5 VDD.t7 193.183
R45 VDD.n6 VDD.t10 193.183
R46 VDD.t5 VDD.n1 109.849
R47 VDD.t3 VDD.n5 109.849
R48 VDD.n6 VDD.t15 109.849
R49 VDD.n14 VDD 11.7877
R50 VDD.n5 VDD.n3 6.3005
R51 VDD.n7 VDD.n6 6.3005
R52 VDD.n15 VDD.n1 6.3005
R53 VDD VDD.n0 5.23855
R54 VDD VDD.n2 5.23855
R55 VDD.n7 VDD.t16 5.21701
R56 VDD.n13 VDD.t14 5.19258
R57 VDD.n8 VDD.n4 5.13287
R58 VDD.n10 VDD.t4 3.91303
R59 VDD.n11 VDD.n10 3.87579
R60 VDD.n11 VDD.t6 3.51066
R61 VDD.n14 VDD.n11 0.272933
R62 VDD.n10 VDD.n9 0.22389
R63 VDD.n9 VDD.n8 0.141016
R64 VDD.n8 VDD 0.106177
R65 VDD.n9 VDD.n3 0.0800484
R66 VDD VDD.n14 0.0783065
R67 VDD.n15 VDD 0.00224194
R68 VDD.n3 VDD 0.00166129
R69 VDD VDD.n7 0.00166129
R70 VDD VDD.n15 0.00166129
R71 VDD VDD.n13 0.00105556
R72 OUT OUT.n3 7.15141
R73 OUT.n2 OUT.n1 3.2163
R74 OUT.n1 OUT.t2 2.2755
R75 OUT.n1 OUT.n0 2.2755
R76 OUT.n2 OUT 0.0445816
R77 OUT OUT.n2 0.0119545
R78 I1.n0 I1.t0 30.9379
R79 I1.n0 I1.t1 21.6422
R80 I1 I1.n0 4.00388
C0 nand2_1.IN2 a_801_256# 0.00372f
C1 I0 nand2_2.OUT 0.202f
C2 Sel OUT 0.00946f
C3 OUT VDD 0.234f
C4 Sel nand2_1.IN2 0.341f
C5 nand2_1.IN2 nand2_2.IN2 0.00212f
C6 Sel a_238_256# 0.0144f
C7 nand2_1.IN2 VDD 0.458f
C8 a_238_256# VDD 3.14e-19
C9 I0 a_801_n344# 0.00293f
C10 nand2_2.IN2 I0 0.0473f
C11 I0 VDD 0.233f
C12 nand2_2.OUT a_801_256# 0.00949f
C13 I1 nand2_1.IN2 0.0959f
C14 I1 a_238_256# 0.00347f
C15 nand2_2.OUT a_801_n344# 0.0964f
C16 Sel nand2_2.OUT 4.46e-19
C17 nand2_2.IN2 nand2_2.OUT 0.12f
C18 nand2_2.OUT VDD 0.637f
C19 nand2_1.IN2 OUT 0.109f
C20 VDD a_801_256# 0.00444f
C21 Sel a_801_n344# 2.62e-19
C22 nand2_2.IN2 a_801_n344# 0.00372f
C23 nand2_1.IN2 a_238_256# 0.069f
C24 Sel nand2_2.IN2 0.136f
C25 VDD a_801_n344# 0.00444f
C26 I0 OUT 1.36e-19
C27 Sel VDD 0.587f
C28 nand2_2.IN2 VDD 0.401f
C29 nand2_2.OUT OUT 0.303f
C30 Sel I1 0.055f
C31 nand2_1.IN2 nand2_2.OUT 0.053f
C32 I1 VDD 0.147f
C33 OUT a_801_256# 0.069f
C34 a_801_n344# VSS 0.0676f
C35 I0 VSS 0.256f
C36 nand2_2.IN2 VSS 0.437f
C37 a_801_256# VSS 0.0676f
C38 a_238_256# VSS 0.0678f
C39 OUT VSS 0.14f
C40 nand2_2.OUT VSS 0.659f
C41 nand2_1.IN2 VSS 0.435f
C42 Sel VSS 0.842f
C43 I1 VSS 0.292f
C44 VDD VSS 4.29f
.ends

