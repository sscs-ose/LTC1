magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -3754 -2410 3754 2410
<< nwell >>
rect -1754 -410 1754 410
<< pmos >>
rect -1580 -280 -1480 280
rect -1376 -280 -1276 280
rect -1172 -280 -1072 280
rect -968 -280 -868 280
rect -764 -280 -664 280
rect -560 -280 -460 280
rect -356 -280 -256 280
rect -152 -280 -52 280
rect 52 -280 152 280
rect 256 -280 356 280
rect 460 -280 560 280
rect 664 -280 764 280
rect 868 -280 968 280
rect 1072 -280 1172 280
rect 1276 -280 1376 280
rect 1480 -280 1580 280
<< pdiff >>
rect -1668 258 -1580 280
rect -1668 -258 -1655 258
rect -1609 -258 -1580 258
rect -1668 -280 -1580 -258
rect -1480 258 -1376 280
rect -1480 -258 -1451 258
rect -1405 -258 -1376 258
rect -1480 -280 -1376 -258
rect -1276 258 -1172 280
rect -1276 -258 -1247 258
rect -1201 -258 -1172 258
rect -1276 -280 -1172 -258
rect -1072 258 -968 280
rect -1072 -258 -1043 258
rect -997 -258 -968 258
rect -1072 -280 -968 -258
rect -868 258 -764 280
rect -868 -258 -839 258
rect -793 -258 -764 258
rect -868 -280 -764 -258
rect -664 258 -560 280
rect -664 -258 -635 258
rect -589 -258 -560 258
rect -664 -280 -560 -258
rect -460 258 -356 280
rect -460 -258 -431 258
rect -385 -258 -356 258
rect -460 -280 -356 -258
rect -256 258 -152 280
rect -256 -258 -227 258
rect -181 -258 -152 258
rect -256 -280 -152 -258
rect -52 258 52 280
rect -52 -258 -23 258
rect 23 -258 52 258
rect -52 -280 52 -258
rect 152 258 256 280
rect 152 -258 181 258
rect 227 -258 256 258
rect 152 -280 256 -258
rect 356 258 460 280
rect 356 -258 385 258
rect 431 -258 460 258
rect 356 -280 460 -258
rect 560 258 664 280
rect 560 -258 589 258
rect 635 -258 664 258
rect 560 -280 664 -258
rect 764 258 868 280
rect 764 -258 793 258
rect 839 -258 868 258
rect 764 -280 868 -258
rect 968 258 1072 280
rect 968 -258 997 258
rect 1043 -258 1072 258
rect 968 -280 1072 -258
rect 1172 258 1276 280
rect 1172 -258 1201 258
rect 1247 -258 1276 258
rect 1172 -280 1276 -258
rect 1376 258 1480 280
rect 1376 -258 1405 258
rect 1451 -258 1480 258
rect 1376 -280 1480 -258
rect 1580 258 1668 280
rect 1580 -258 1609 258
rect 1655 -258 1668 258
rect 1580 -280 1668 -258
<< pdiffc >>
rect -1655 -258 -1609 258
rect -1451 -258 -1405 258
rect -1247 -258 -1201 258
rect -1043 -258 -997 258
rect -839 -258 -793 258
rect -635 -258 -589 258
rect -431 -258 -385 258
rect -227 -258 -181 258
rect -23 -258 23 258
rect 181 -258 227 258
rect 385 -258 431 258
rect 589 -258 635 258
rect 793 -258 839 258
rect 997 -258 1043 258
rect 1201 -258 1247 258
rect 1405 -258 1451 258
rect 1609 -258 1655 258
<< polysilicon >>
rect -1580 280 -1480 324
rect -1376 280 -1276 324
rect -1172 280 -1072 324
rect -968 280 -868 324
rect -764 280 -664 324
rect -560 280 -460 324
rect -356 280 -256 324
rect -152 280 -52 324
rect 52 280 152 324
rect 256 280 356 324
rect 460 280 560 324
rect 664 280 764 324
rect 868 280 968 324
rect 1072 280 1172 324
rect 1276 280 1376 324
rect 1480 280 1580 324
rect -1580 -324 -1480 -280
rect -1376 -324 -1276 -280
rect -1172 -324 -1072 -280
rect -968 -324 -868 -280
rect -764 -324 -664 -280
rect -560 -324 -460 -280
rect -356 -324 -256 -280
rect -152 -324 -52 -280
rect 52 -324 152 -280
rect 256 -324 356 -280
rect 460 -324 560 -280
rect 664 -324 764 -280
rect 868 -324 968 -280
rect 1072 -324 1172 -280
rect 1276 -324 1376 -280
rect 1480 -324 1580 -280
<< metal1 >>
rect -1655 258 -1609 278
rect -1655 -278 -1609 -258
rect -1451 258 -1405 278
rect -1451 -278 -1405 -258
rect -1247 258 -1201 278
rect -1247 -278 -1201 -258
rect -1043 258 -997 278
rect -1043 -278 -997 -258
rect -839 258 -793 278
rect -839 -278 -793 -258
rect -635 258 -589 278
rect -635 -278 -589 -258
rect -431 258 -385 278
rect -431 -278 -385 -258
rect -227 258 -181 278
rect -227 -278 -181 -258
rect -23 258 23 278
rect -23 -278 23 -258
rect 181 258 227 278
rect 181 -278 227 -258
rect 385 258 431 278
rect 385 -278 431 -258
rect 589 258 635 278
rect 589 -278 635 -258
rect 793 258 839 278
rect 793 -278 839 -258
rect 997 258 1043 278
rect 997 -278 1043 -258
rect 1201 258 1247 278
rect 1201 -278 1247 -258
rect 1405 258 1451 278
rect 1405 -278 1451 -258
rect 1609 258 1655 278
rect 1609 -278 1655 -258
<< end >>
