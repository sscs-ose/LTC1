magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -3626 -1382 3626 1382
<< metal2 >>
rect -2626 377 2626 382
rect -2626 349 -2621 377
rect -2593 349 -2555 377
rect -2527 349 -2489 377
rect -2461 349 -2423 377
rect -2395 349 -2357 377
rect -2329 349 -2291 377
rect -2263 349 -2225 377
rect -2197 349 -2159 377
rect -2131 349 -2093 377
rect -2065 349 -2027 377
rect -1999 349 -1961 377
rect -1933 349 -1895 377
rect -1867 349 -1829 377
rect -1801 349 -1763 377
rect -1735 349 -1697 377
rect -1669 349 -1631 377
rect -1603 349 -1565 377
rect -1537 349 -1499 377
rect -1471 349 -1433 377
rect -1405 349 -1367 377
rect -1339 349 -1301 377
rect -1273 349 -1235 377
rect -1207 349 -1169 377
rect -1141 349 -1103 377
rect -1075 349 -1037 377
rect -1009 349 -971 377
rect -943 349 -905 377
rect -877 349 -839 377
rect -811 349 -773 377
rect -745 349 -707 377
rect -679 349 -641 377
rect -613 349 -575 377
rect -547 349 -509 377
rect -481 349 -443 377
rect -415 349 -377 377
rect -349 349 -311 377
rect -283 349 -245 377
rect -217 349 -179 377
rect -151 349 -113 377
rect -85 349 -47 377
rect -19 349 19 377
rect 47 349 85 377
rect 113 349 151 377
rect 179 349 217 377
rect 245 349 283 377
rect 311 349 349 377
rect 377 349 415 377
rect 443 349 481 377
rect 509 349 547 377
rect 575 349 613 377
rect 641 349 679 377
rect 707 349 745 377
rect 773 349 811 377
rect 839 349 877 377
rect 905 349 943 377
rect 971 349 1009 377
rect 1037 349 1075 377
rect 1103 349 1141 377
rect 1169 349 1207 377
rect 1235 349 1273 377
rect 1301 349 1339 377
rect 1367 349 1405 377
rect 1433 349 1471 377
rect 1499 349 1537 377
rect 1565 349 1603 377
rect 1631 349 1669 377
rect 1697 349 1735 377
rect 1763 349 1801 377
rect 1829 349 1867 377
rect 1895 349 1933 377
rect 1961 349 1999 377
rect 2027 349 2065 377
rect 2093 349 2131 377
rect 2159 349 2197 377
rect 2225 349 2263 377
rect 2291 349 2329 377
rect 2357 349 2395 377
rect 2423 349 2461 377
rect 2489 349 2527 377
rect 2555 349 2593 377
rect 2621 349 2626 377
rect -2626 311 2626 349
rect -2626 283 -2621 311
rect -2593 283 -2555 311
rect -2527 283 -2489 311
rect -2461 283 -2423 311
rect -2395 283 -2357 311
rect -2329 283 -2291 311
rect -2263 283 -2225 311
rect -2197 283 -2159 311
rect -2131 283 -2093 311
rect -2065 283 -2027 311
rect -1999 283 -1961 311
rect -1933 283 -1895 311
rect -1867 283 -1829 311
rect -1801 283 -1763 311
rect -1735 283 -1697 311
rect -1669 283 -1631 311
rect -1603 283 -1565 311
rect -1537 283 -1499 311
rect -1471 283 -1433 311
rect -1405 283 -1367 311
rect -1339 283 -1301 311
rect -1273 283 -1235 311
rect -1207 283 -1169 311
rect -1141 283 -1103 311
rect -1075 283 -1037 311
rect -1009 283 -971 311
rect -943 283 -905 311
rect -877 283 -839 311
rect -811 283 -773 311
rect -745 283 -707 311
rect -679 283 -641 311
rect -613 283 -575 311
rect -547 283 -509 311
rect -481 283 -443 311
rect -415 283 -377 311
rect -349 283 -311 311
rect -283 283 -245 311
rect -217 283 -179 311
rect -151 283 -113 311
rect -85 283 -47 311
rect -19 283 19 311
rect 47 283 85 311
rect 113 283 151 311
rect 179 283 217 311
rect 245 283 283 311
rect 311 283 349 311
rect 377 283 415 311
rect 443 283 481 311
rect 509 283 547 311
rect 575 283 613 311
rect 641 283 679 311
rect 707 283 745 311
rect 773 283 811 311
rect 839 283 877 311
rect 905 283 943 311
rect 971 283 1009 311
rect 1037 283 1075 311
rect 1103 283 1141 311
rect 1169 283 1207 311
rect 1235 283 1273 311
rect 1301 283 1339 311
rect 1367 283 1405 311
rect 1433 283 1471 311
rect 1499 283 1537 311
rect 1565 283 1603 311
rect 1631 283 1669 311
rect 1697 283 1735 311
rect 1763 283 1801 311
rect 1829 283 1867 311
rect 1895 283 1933 311
rect 1961 283 1999 311
rect 2027 283 2065 311
rect 2093 283 2131 311
rect 2159 283 2197 311
rect 2225 283 2263 311
rect 2291 283 2329 311
rect 2357 283 2395 311
rect 2423 283 2461 311
rect 2489 283 2527 311
rect 2555 283 2593 311
rect 2621 283 2626 311
rect -2626 245 2626 283
rect -2626 217 -2621 245
rect -2593 217 -2555 245
rect -2527 217 -2489 245
rect -2461 217 -2423 245
rect -2395 217 -2357 245
rect -2329 217 -2291 245
rect -2263 217 -2225 245
rect -2197 217 -2159 245
rect -2131 217 -2093 245
rect -2065 217 -2027 245
rect -1999 217 -1961 245
rect -1933 217 -1895 245
rect -1867 217 -1829 245
rect -1801 217 -1763 245
rect -1735 217 -1697 245
rect -1669 217 -1631 245
rect -1603 217 -1565 245
rect -1537 217 -1499 245
rect -1471 217 -1433 245
rect -1405 217 -1367 245
rect -1339 217 -1301 245
rect -1273 217 -1235 245
rect -1207 217 -1169 245
rect -1141 217 -1103 245
rect -1075 217 -1037 245
rect -1009 217 -971 245
rect -943 217 -905 245
rect -877 217 -839 245
rect -811 217 -773 245
rect -745 217 -707 245
rect -679 217 -641 245
rect -613 217 -575 245
rect -547 217 -509 245
rect -481 217 -443 245
rect -415 217 -377 245
rect -349 217 -311 245
rect -283 217 -245 245
rect -217 217 -179 245
rect -151 217 -113 245
rect -85 217 -47 245
rect -19 217 19 245
rect 47 217 85 245
rect 113 217 151 245
rect 179 217 217 245
rect 245 217 283 245
rect 311 217 349 245
rect 377 217 415 245
rect 443 217 481 245
rect 509 217 547 245
rect 575 217 613 245
rect 641 217 679 245
rect 707 217 745 245
rect 773 217 811 245
rect 839 217 877 245
rect 905 217 943 245
rect 971 217 1009 245
rect 1037 217 1075 245
rect 1103 217 1141 245
rect 1169 217 1207 245
rect 1235 217 1273 245
rect 1301 217 1339 245
rect 1367 217 1405 245
rect 1433 217 1471 245
rect 1499 217 1537 245
rect 1565 217 1603 245
rect 1631 217 1669 245
rect 1697 217 1735 245
rect 1763 217 1801 245
rect 1829 217 1867 245
rect 1895 217 1933 245
rect 1961 217 1999 245
rect 2027 217 2065 245
rect 2093 217 2131 245
rect 2159 217 2197 245
rect 2225 217 2263 245
rect 2291 217 2329 245
rect 2357 217 2395 245
rect 2423 217 2461 245
rect 2489 217 2527 245
rect 2555 217 2593 245
rect 2621 217 2626 245
rect -2626 179 2626 217
rect -2626 151 -2621 179
rect -2593 151 -2555 179
rect -2527 151 -2489 179
rect -2461 151 -2423 179
rect -2395 151 -2357 179
rect -2329 151 -2291 179
rect -2263 151 -2225 179
rect -2197 151 -2159 179
rect -2131 151 -2093 179
rect -2065 151 -2027 179
rect -1999 151 -1961 179
rect -1933 151 -1895 179
rect -1867 151 -1829 179
rect -1801 151 -1763 179
rect -1735 151 -1697 179
rect -1669 151 -1631 179
rect -1603 151 -1565 179
rect -1537 151 -1499 179
rect -1471 151 -1433 179
rect -1405 151 -1367 179
rect -1339 151 -1301 179
rect -1273 151 -1235 179
rect -1207 151 -1169 179
rect -1141 151 -1103 179
rect -1075 151 -1037 179
rect -1009 151 -971 179
rect -943 151 -905 179
rect -877 151 -839 179
rect -811 151 -773 179
rect -745 151 -707 179
rect -679 151 -641 179
rect -613 151 -575 179
rect -547 151 -509 179
rect -481 151 -443 179
rect -415 151 -377 179
rect -349 151 -311 179
rect -283 151 -245 179
rect -217 151 -179 179
rect -151 151 -113 179
rect -85 151 -47 179
rect -19 151 19 179
rect 47 151 85 179
rect 113 151 151 179
rect 179 151 217 179
rect 245 151 283 179
rect 311 151 349 179
rect 377 151 415 179
rect 443 151 481 179
rect 509 151 547 179
rect 575 151 613 179
rect 641 151 679 179
rect 707 151 745 179
rect 773 151 811 179
rect 839 151 877 179
rect 905 151 943 179
rect 971 151 1009 179
rect 1037 151 1075 179
rect 1103 151 1141 179
rect 1169 151 1207 179
rect 1235 151 1273 179
rect 1301 151 1339 179
rect 1367 151 1405 179
rect 1433 151 1471 179
rect 1499 151 1537 179
rect 1565 151 1603 179
rect 1631 151 1669 179
rect 1697 151 1735 179
rect 1763 151 1801 179
rect 1829 151 1867 179
rect 1895 151 1933 179
rect 1961 151 1999 179
rect 2027 151 2065 179
rect 2093 151 2131 179
rect 2159 151 2197 179
rect 2225 151 2263 179
rect 2291 151 2329 179
rect 2357 151 2395 179
rect 2423 151 2461 179
rect 2489 151 2527 179
rect 2555 151 2593 179
rect 2621 151 2626 179
rect -2626 113 2626 151
rect -2626 85 -2621 113
rect -2593 85 -2555 113
rect -2527 85 -2489 113
rect -2461 85 -2423 113
rect -2395 85 -2357 113
rect -2329 85 -2291 113
rect -2263 85 -2225 113
rect -2197 85 -2159 113
rect -2131 85 -2093 113
rect -2065 85 -2027 113
rect -1999 85 -1961 113
rect -1933 85 -1895 113
rect -1867 85 -1829 113
rect -1801 85 -1763 113
rect -1735 85 -1697 113
rect -1669 85 -1631 113
rect -1603 85 -1565 113
rect -1537 85 -1499 113
rect -1471 85 -1433 113
rect -1405 85 -1367 113
rect -1339 85 -1301 113
rect -1273 85 -1235 113
rect -1207 85 -1169 113
rect -1141 85 -1103 113
rect -1075 85 -1037 113
rect -1009 85 -971 113
rect -943 85 -905 113
rect -877 85 -839 113
rect -811 85 -773 113
rect -745 85 -707 113
rect -679 85 -641 113
rect -613 85 -575 113
rect -547 85 -509 113
rect -481 85 -443 113
rect -415 85 -377 113
rect -349 85 -311 113
rect -283 85 -245 113
rect -217 85 -179 113
rect -151 85 -113 113
rect -85 85 -47 113
rect -19 85 19 113
rect 47 85 85 113
rect 113 85 151 113
rect 179 85 217 113
rect 245 85 283 113
rect 311 85 349 113
rect 377 85 415 113
rect 443 85 481 113
rect 509 85 547 113
rect 575 85 613 113
rect 641 85 679 113
rect 707 85 745 113
rect 773 85 811 113
rect 839 85 877 113
rect 905 85 943 113
rect 971 85 1009 113
rect 1037 85 1075 113
rect 1103 85 1141 113
rect 1169 85 1207 113
rect 1235 85 1273 113
rect 1301 85 1339 113
rect 1367 85 1405 113
rect 1433 85 1471 113
rect 1499 85 1537 113
rect 1565 85 1603 113
rect 1631 85 1669 113
rect 1697 85 1735 113
rect 1763 85 1801 113
rect 1829 85 1867 113
rect 1895 85 1933 113
rect 1961 85 1999 113
rect 2027 85 2065 113
rect 2093 85 2131 113
rect 2159 85 2197 113
rect 2225 85 2263 113
rect 2291 85 2329 113
rect 2357 85 2395 113
rect 2423 85 2461 113
rect 2489 85 2527 113
rect 2555 85 2593 113
rect 2621 85 2626 113
rect -2626 47 2626 85
rect -2626 19 -2621 47
rect -2593 19 -2555 47
rect -2527 19 -2489 47
rect -2461 19 -2423 47
rect -2395 19 -2357 47
rect -2329 19 -2291 47
rect -2263 19 -2225 47
rect -2197 19 -2159 47
rect -2131 19 -2093 47
rect -2065 19 -2027 47
rect -1999 19 -1961 47
rect -1933 19 -1895 47
rect -1867 19 -1829 47
rect -1801 19 -1763 47
rect -1735 19 -1697 47
rect -1669 19 -1631 47
rect -1603 19 -1565 47
rect -1537 19 -1499 47
rect -1471 19 -1433 47
rect -1405 19 -1367 47
rect -1339 19 -1301 47
rect -1273 19 -1235 47
rect -1207 19 -1169 47
rect -1141 19 -1103 47
rect -1075 19 -1037 47
rect -1009 19 -971 47
rect -943 19 -905 47
rect -877 19 -839 47
rect -811 19 -773 47
rect -745 19 -707 47
rect -679 19 -641 47
rect -613 19 -575 47
rect -547 19 -509 47
rect -481 19 -443 47
rect -415 19 -377 47
rect -349 19 -311 47
rect -283 19 -245 47
rect -217 19 -179 47
rect -151 19 -113 47
rect -85 19 -47 47
rect -19 19 19 47
rect 47 19 85 47
rect 113 19 151 47
rect 179 19 217 47
rect 245 19 283 47
rect 311 19 349 47
rect 377 19 415 47
rect 443 19 481 47
rect 509 19 547 47
rect 575 19 613 47
rect 641 19 679 47
rect 707 19 745 47
rect 773 19 811 47
rect 839 19 877 47
rect 905 19 943 47
rect 971 19 1009 47
rect 1037 19 1075 47
rect 1103 19 1141 47
rect 1169 19 1207 47
rect 1235 19 1273 47
rect 1301 19 1339 47
rect 1367 19 1405 47
rect 1433 19 1471 47
rect 1499 19 1537 47
rect 1565 19 1603 47
rect 1631 19 1669 47
rect 1697 19 1735 47
rect 1763 19 1801 47
rect 1829 19 1867 47
rect 1895 19 1933 47
rect 1961 19 1999 47
rect 2027 19 2065 47
rect 2093 19 2131 47
rect 2159 19 2197 47
rect 2225 19 2263 47
rect 2291 19 2329 47
rect 2357 19 2395 47
rect 2423 19 2461 47
rect 2489 19 2527 47
rect 2555 19 2593 47
rect 2621 19 2626 47
rect -2626 -19 2626 19
rect -2626 -47 -2621 -19
rect -2593 -47 -2555 -19
rect -2527 -47 -2489 -19
rect -2461 -47 -2423 -19
rect -2395 -47 -2357 -19
rect -2329 -47 -2291 -19
rect -2263 -47 -2225 -19
rect -2197 -47 -2159 -19
rect -2131 -47 -2093 -19
rect -2065 -47 -2027 -19
rect -1999 -47 -1961 -19
rect -1933 -47 -1895 -19
rect -1867 -47 -1829 -19
rect -1801 -47 -1763 -19
rect -1735 -47 -1697 -19
rect -1669 -47 -1631 -19
rect -1603 -47 -1565 -19
rect -1537 -47 -1499 -19
rect -1471 -47 -1433 -19
rect -1405 -47 -1367 -19
rect -1339 -47 -1301 -19
rect -1273 -47 -1235 -19
rect -1207 -47 -1169 -19
rect -1141 -47 -1103 -19
rect -1075 -47 -1037 -19
rect -1009 -47 -971 -19
rect -943 -47 -905 -19
rect -877 -47 -839 -19
rect -811 -47 -773 -19
rect -745 -47 -707 -19
rect -679 -47 -641 -19
rect -613 -47 -575 -19
rect -547 -47 -509 -19
rect -481 -47 -443 -19
rect -415 -47 -377 -19
rect -349 -47 -311 -19
rect -283 -47 -245 -19
rect -217 -47 -179 -19
rect -151 -47 -113 -19
rect -85 -47 -47 -19
rect -19 -47 19 -19
rect 47 -47 85 -19
rect 113 -47 151 -19
rect 179 -47 217 -19
rect 245 -47 283 -19
rect 311 -47 349 -19
rect 377 -47 415 -19
rect 443 -47 481 -19
rect 509 -47 547 -19
rect 575 -47 613 -19
rect 641 -47 679 -19
rect 707 -47 745 -19
rect 773 -47 811 -19
rect 839 -47 877 -19
rect 905 -47 943 -19
rect 971 -47 1009 -19
rect 1037 -47 1075 -19
rect 1103 -47 1141 -19
rect 1169 -47 1207 -19
rect 1235 -47 1273 -19
rect 1301 -47 1339 -19
rect 1367 -47 1405 -19
rect 1433 -47 1471 -19
rect 1499 -47 1537 -19
rect 1565 -47 1603 -19
rect 1631 -47 1669 -19
rect 1697 -47 1735 -19
rect 1763 -47 1801 -19
rect 1829 -47 1867 -19
rect 1895 -47 1933 -19
rect 1961 -47 1999 -19
rect 2027 -47 2065 -19
rect 2093 -47 2131 -19
rect 2159 -47 2197 -19
rect 2225 -47 2263 -19
rect 2291 -47 2329 -19
rect 2357 -47 2395 -19
rect 2423 -47 2461 -19
rect 2489 -47 2527 -19
rect 2555 -47 2593 -19
rect 2621 -47 2626 -19
rect -2626 -85 2626 -47
rect -2626 -113 -2621 -85
rect -2593 -113 -2555 -85
rect -2527 -113 -2489 -85
rect -2461 -113 -2423 -85
rect -2395 -113 -2357 -85
rect -2329 -113 -2291 -85
rect -2263 -113 -2225 -85
rect -2197 -113 -2159 -85
rect -2131 -113 -2093 -85
rect -2065 -113 -2027 -85
rect -1999 -113 -1961 -85
rect -1933 -113 -1895 -85
rect -1867 -113 -1829 -85
rect -1801 -113 -1763 -85
rect -1735 -113 -1697 -85
rect -1669 -113 -1631 -85
rect -1603 -113 -1565 -85
rect -1537 -113 -1499 -85
rect -1471 -113 -1433 -85
rect -1405 -113 -1367 -85
rect -1339 -113 -1301 -85
rect -1273 -113 -1235 -85
rect -1207 -113 -1169 -85
rect -1141 -113 -1103 -85
rect -1075 -113 -1037 -85
rect -1009 -113 -971 -85
rect -943 -113 -905 -85
rect -877 -113 -839 -85
rect -811 -113 -773 -85
rect -745 -113 -707 -85
rect -679 -113 -641 -85
rect -613 -113 -575 -85
rect -547 -113 -509 -85
rect -481 -113 -443 -85
rect -415 -113 -377 -85
rect -349 -113 -311 -85
rect -283 -113 -245 -85
rect -217 -113 -179 -85
rect -151 -113 -113 -85
rect -85 -113 -47 -85
rect -19 -113 19 -85
rect 47 -113 85 -85
rect 113 -113 151 -85
rect 179 -113 217 -85
rect 245 -113 283 -85
rect 311 -113 349 -85
rect 377 -113 415 -85
rect 443 -113 481 -85
rect 509 -113 547 -85
rect 575 -113 613 -85
rect 641 -113 679 -85
rect 707 -113 745 -85
rect 773 -113 811 -85
rect 839 -113 877 -85
rect 905 -113 943 -85
rect 971 -113 1009 -85
rect 1037 -113 1075 -85
rect 1103 -113 1141 -85
rect 1169 -113 1207 -85
rect 1235 -113 1273 -85
rect 1301 -113 1339 -85
rect 1367 -113 1405 -85
rect 1433 -113 1471 -85
rect 1499 -113 1537 -85
rect 1565 -113 1603 -85
rect 1631 -113 1669 -85
rect 1697 -113 1735 -85
rect 1763 -113 1801 -85
rect 1829 -113 1867 -85
rect 1895 -113 1933 -85
rect 1961 -113 1999 -85
rect 2027 -113 2065 -85
rect 2093 -113 2131 -85
rect 2159 -113 2197 -85
rect 2225 -113 2263 -85
rect 2291 -113 2329 -85
rect 2357 -113 2395 -85
rect 2423 -113 2461 -85
rect 2489 -113 2527 -85
rect 2555 -113 2593 -85
rect 2621 -113 2626 -85
rect -2626 -151 2626 -113
rect -2626 -179 -2621 -151
rect -2593 -179 -2555 -151
rect -2527 -179 -2489 -151
rect -2461 -179 -2423 -151
rect -2395 -179 -2357 -151
rect -2329 -179 -2291 -151
rect -2263 -179 -2225 -151
rect -2197 -179 -2159 -151
rect -2131 -179 -2093 -151
rect -2065 -179 -2027 -151
rect -1999 -179 -1961 -151
rect -1933 -179 -1895 -151
rect -1867 -179 -1829 -151
rect -1801 -179 -1763 -151
rect -1735 -179 -1697 -151
rect -1669 -179 -1631 -151
rect -1603 -179 -1565 -151
rect -1537 -179 -1499 -151
rect -1471 -179 -1433 -151
rect -1405 -179 -1367 -151
rect -1339 -179 -1301 -151
rect -1273 -179 -1235 -151
rect -1207 -179 -1169 -151
rect -1141 -179 -1103 -151
rect -1075 -179 -1037 -151
rect -1009 -179 -971 -151
rect -943 -179 -905 -151
rect -877 -179 -839 -151
rect -811 -179 -773 -151
rect -745 -179 -707 -151
rect -679 -179 -641 -151
rect -613 -179 -575 -151
rect -547 -179 -509 -151
rect -481 -179 -443 -151
rect -415 -179 -377 -151
rect -349 -179 -311 -151
rect -283 -179 -245 -151
rect -217 -179 -179 -151
rect -151 -179 -113 -151
rect -85 -179 -47 -151
rect -19 -179 19 -151
rect 47 -179 85 -151
rect 113 -179 151 -151
rect 179 -179 217 -151
rect 245 -179 283 -151
rect 311 -179 349 -151
rect 377 -179 415 -151
rect 443 -179 481 -151
rect 509 -179 547 -151
rect 575 -179 613 -151
rect 641 -179 679 -151
rect 707 -179 745 -151
rect 773 -179 811 -151
rect 839 -179 877 -151
rect 905 -179 943 -151
rect 971 -179 1009 -151
rect 1037 -179 1075 -151
rect 1103 -179 1141 -151
rect 1169 -179 1207 -151
rect 1235 -179 1273 -151
rect 1301 -179 1339 -151
rect 1367 -179 1405 -151
rect 1433 -179 1471 -151
rect 1499 -179 1537 -151
rect 1565 -179 1603 -151
rect 1631 -179 1669 -151
rect 1697 -179 1735 -151
rect 1763 -179 1801 -151
rect 1829 -179 1867 -151
rect 1895 -179 1933 -151
rect 1961 -179 1999 -151
rect 2027 -179 2065 -151
rect 2093 -179 2131 -151
rect 2159 -179 2197 -151
rect 2225 -179 2263 -151
rect 2291 -179 2329 -151
rect 2357 -179 2395 -151
rect 2423 -179 2461 -151
rect 2489 -179 2527 -151
rect 2555 -179 2593 -151
rect 2621 -179 2626 -151
rect -2626 -217 2626 -179
rect -2626 -245 -2621 -217
rect -2593 -245 -2555 -217
rect -2527 -245 -2489 -217
rect -2461 -245 -2423 -217
rect -2395 -245 -2357 -217
rect -2329 -245 -2291 -217
rect -2263 -245 -2225 -217
rect -2197 -245 -2159 -217
rect -2131 -245 -2093 -217
rect -2065 -245 -2027 -217
rect -1999 -245 -1961 -217
rect -1933 -245 -1895 -217
rect -1867 -245 -1829 -217
rect -1801 -245 -1763 -217
rect -1735 -245 -1697 -217
rect -1669 -245 -1631 -217
rect -1603 -245 -1565 -217
rect -1537 -245 -1499 -217
rect -1471 -245 -1433 -217
rect -1405 -245 -1367 -217
rect -1339 -245 -1301 -217
rect -1273 -245 -1235 -217
rect -1207 -245 -1169 -217
rect -1141 -245 -1103 -217
rect -1075 -245 -1037 -217
rect -1009 -245 -971 -217
rect -943 -245 -905 -217
rect -877 -245 -839 -217
rect -811 -245 -773 -217
rect -745 -245 -707 -217
rect -679 -245 -641 -217
rect -613 -245 -575 -217
rect -547 -245 -509 -217
rect -481 -245 -443 -217
rect -415 -245 -377 -217
rect -349 -245 -311 -217
rect -283 -245 -245 -217
rect -217 -245 -179 -217
rect -151 -245 -113 -217
rect -85 -245 -47 -217
rect -19 -245 19 -217
rect 47 -245 85 -217
rect 113 -245 151 -217
rect 179 -245 217 -217
rect 245 -245 283 -217
rect 311 -245 349 -217
rect 377 -245 415 -217
rect 443 -245 481 -217
rect 509 -245 547 -217
rect 575 -245 613 -217
rect 641 -245 679 -217
rect 707 -245 745 -217
rect 773 -245 811 -217
rect 839 -245 877 -217
rect 905 -245 943 -217
rect 971 -245 1009 -217
rect 1037 -245 1075 -217
rect 1103 -245 1141 -217
rect 1169 -245 1207 -217
rect 1235 -245 1273 -217
rect 1301 -245 1339 -217
rect 1367 -245 1405 -217
rect 1433 -245 1471 -217
rect 1499 -245 1537 -217
rect 1565 -245 1603 -217
rect 1631 -245 1669 -217
rect 1697 -245 1735 -217
rect 1763 -245 1801 -217
rect 1829 -245 1867 -217
rect 1895 -245 1933 -217
rect 1961 -245 1999 -217
rect 2027 -245 2065 -217
rect 2093 -245 2131 -217
rect 2159 -245 2197 -217
rect 2225 -245 2263 -217
rect 2291 -245 2329 -217
rect 2357 -245 2395 -217
rect 2423 -245 2461 -217
rect 2489 -245 2527 -217
rect 2555 -245 2593 -217
rect 2621 -245 2626 -217
rect -2626 -283 2626 -245
rect -2626 -311 -2621 -283
rect -2593 -311 -2555 -283
rect -2527 -311 -2489 -283
rect -2461 -311 -2423 -283
rect -2395 -311 -2357 -283
rect -2329 -311 -2291 -283
rect -2263 -311 -2225 -283
rect -2197 -311 -2159 -283
rect -2131 -311 -2093 -283
rect -2065 -311 -2027 -283
rect -1999 -311 -1961 -283
rect -1933 -311 -1895 -283
rect -1867 -311 -1829 -283
rect -1801 -311 -1763 -283
rect -1735 -311 -1697 -283
rect -1669 -311 -1631 -283
rect -1603 -311 -1565 -283
rect -1537 -311 -1499 -283
rect -1471 -311 -1433 -283
rect -1405 -311 -1367 -283
rect -1339 -311 -1301 -283
rect -1273 -311 -1235 -283
rect -1207 -311 -1169 -283
rect -1141 -311 -1103 -283
rect -1075 -311 -1037 -283
rect -1009 -311 -971 -283
rect -943 -311 -905 -283
rect -877 -311 -839 -283
rect -811 -311 -773 -283
rect -745 -311 -707 -283
rect -679 -311 -641 -283
rect -613 -311 -575 -283
rect -547 -311 -509 -283
rect -481 -311 -443 -283
rect -415 -311 -377 -283
rect -349 -311 -311 -283
rect -283 -311 -245 -283
rect -217 -311 -179 -283
rect -151 -311 -113 -283
rect -85 -311 -47 -283
rect -19 -311 19 -283
rect 47 -311 85 -283
rect 113 -311 151 -283
rect 179 -311 217 -283
rect 245 -311 283 -283
rect 311 -311 349 -283
rect 377 -311 415 -283
rect 443 -311 481 -283
rect 509 -311 547 -283
rect 575 -311 613 -283
rect 641 -311 679 -283
rect 707 -311 745 -283
rect 773 -311 811 -283
rect 839 -311 877 -283
rect 905 -311 943 -283
rect 971 -311 1009 -283
rect 1037 -311 1075 -283
rect 1103 -311 1141 -283
rect 1169 -311 1207 -283
rect 1235 -311 1273 -283
rect 1301 -311 1339 -283
rect 1367 -311 1405 -283
rect 1433 -311 1471 -283
rect 1499 -311 1537 -283
rect 1565 -311 1603 -283
rect 1631 -311 1669 -283
rect 1697 -311 1735 -283
rect 1763 -311 1801 -283
rect 1829 -311 1867 -283
rect 1895 -311 1933 -283
rect 1961 -311 1999 -283
rect 2027 -311 2065 -283
rect 2093 -311 2131 -283
rect 2159 -311 2197 -283
rect 2225 -311 2263 -283
rect 2291 -311 2329 -283
rect 2357 -311 2395 -283
rect 2423 -311 2461 -283
rect 2489 -311 2527 -283
rect 2555 -311 2593 -283
rect 2621 -311 2626 -283
rect -2626 -349 2626 -311
rect -2626 -377 -2621 -349
rect -2593 -377 -2555 -349
rect -2527 -377 -2489 -349
rect -2461 -377 -2423 -349
rect -2395 -377 -2357 -349
rect -2329 -377 -2291 -349
rect -2263 -377 -2225 -349
rect -2197 -377 -2159 -349
rect -2131 -377 -2093 -349
rect -2065 -377 -2027 -349
rect -1999 -377 -1961 -349
rect -1933 -377 -1895 -349
rect -1867 -377 -1829 -349
rect -1801 -377 -1763 -349
rect -1735 -377 -1697 -349
rect -1669 -377 -1631 -349
rect -1603 -377 -1565 -349
rect -1537 -377 -1499 -349
rect -1471 -377 -1433 -349
rect -1405 -377 -1367 -349
rect -1339 -377 -1301 -349
rect -1273 -377 -1235 -349
rect -1207 -377 -1169 -349
rect -1141 -377 -1103 -349
rect -1075 -377 -1037 -349
rect -1009 -377 -971 -349
rect -943 -377 -905 -349
rect -877 -377 -839 -349
rect -811 -377 -773 -349
rect -745 -377 -707 -349
rect -679 -377 -641 -349
rect -613 -377 -575 -349
rect -547 -377 -509 -349
rect -481 -377 -443 -349
rect -415 -377 -377 -349
rect -349 -377 -311 -349
rect -283 -377 -245 -349
rect -217 -377 -179 -349
rect -151 -377 -113 -349
rect -85 -377 -47 -349
rect -19 -377 19 -349
rect 47 -377 85 -349
rect 113 -377 151 -349
rect 179 -377 217 -349
rect 245 -377 283 -349
rect 311 -377 349 -349
rect 377 -377 415 -349
rect 443 -377 481 -349
rect 509 -377 547 -349
rect 575 -377 613 -349
rect 641 -377 679 -349
rect 707 -377 745 -349
rect 773 -377 811 -349
rect 839 -377 877 -349
rect 905 -377 943 -349
rect 971 -377 1009 -349
rect 1037 -377 1075 -349
rect 1103 -377 1141 -349
rect 1169 -377 1207 -349
rect 1235 -377 1273 -349
rect 1301 -377 1339 -349
rect 1367 -377 1405 -349
rect 1433 -377 1471 -349
rect 1499 -377 1537 -349
rect 1565 -377 1603 -349
rect 1631 -377 1669 -349
rect 1697 -377 1735 -349
rect 1763 -377 1801 -349
rect 1829 -377 1867 -349
rect 1895 -377 1933 -349
rect 1961 -377 1999 -349
rect 2027 -377 2065 -349
rect 2093 -377 2131 -349
rect 2159 -377 2197 -349
rect 2225 -377 2263 -349
rect 2291 -377 2329 -349
rect 2357 -377 2395 -349
rect 2423 -377 2461 -349
rect 2489 -377 2527 -349
rect 2555 -377 2593 -349
rect 2621 -377 2626 -349
rect -2626 -382 2626 -377
<< via2 >>
rect -2621 349 -2593 377
rect -2555 349 -2527 377
rect -2489 349 -2461 377
rect -2423 349 -2395 377
rect -2357 349 -2329 377
rect -2291 349 -2263 377
rect -2225 349 -2197 377
rect -2159 349 -2131 377
rect -2093 349 -2065 377
rect -2027 349 -1999 377
rect -1961 349 -1933 377
rect -1895 349 -1867 377
rect -1829 349 -1801 377
rect -1763 349 -1735 377
rect -1697 349 -1669 377
rect -1631 349 -1603 377
rect -1565 349 -1537 377
rect -1499 349 -1471 377
rect -1433 349 -1405 377
rect -1367 349 -1339 377
rect -1301 349 -1273 377
rect -1235 349 -1207 377
rect -1169 349 -1141 377
rect -1103 349 -1075 377
rect -1037 349 -1009 377
rect -971 349 -943 377
rect -905 349 -877 377
rect -839 349 -811 377
rect -773 349 -745 377
rect -707 349 -679 377
rect -641 349 -613 377
rect -575 349 -547 377
rect -509 349 -481 377
rect -443 349 -415 377
rect -377 349 -349 377
rect -311 349 -283 377
rect -245 349 -217 377
rect -179 349 -151 377
rect -113 349 -85 377
rect -47 349 -19 377
rect 19 349 47 377
rect 85 349 113 377
rect 151 349 179 377
rect 217 349 245 377
rect 283 349 311 377
rect 349 349 377 377
rect 415 349 443 377
rect 481 349 509 377
rect 547 349 575 377
rect 613 349 641 377
rect 679 349 707 377
rect 745 349 773 377
rect 811 349 839 377
rect 877 349 905 377
rect 943 349 971 377
rect 1009 349 1037 377
rect 1075 349 1103 377
rect 1141 349 1169 377
rect 1207 349 1235 377
rect 1273 349 1301 377
rect 1339 349 1367 377
rect 1405 349 1433 377
rect 1471 349 1499 377
rect 1537 349 1565 377
rect 1603 349 1631 377
rect 1669 349 1697 377
rect 1735 349 1763 377
rect 1801 349 1829 377
rect 1867 349 1895 377
rect 1933 349 1961 377
rect 1999 349 2027 377
rect 2065 349 2093 377
rect 2131 349 2159 377
rect 2197 349 2225 377
rect 2263 349 2291 377
rect 2329 349 2357 377
rect 2395 349 2423 377
rect 2461 349 2489 377
rect 2527 349 2555 377
rect 2593 349 2621 377
rect -2621 283 -2593 311
rect -2555 283 -2527 311
rect -2489 283 -2461 311
rect -2423 283 -2395 311
rect -2357 283 -2329 311
rect -2291 283 -2263 311
rect -2225 283 -2197 311
rect -2159 283 -2131 311
rect -2093 283 -2065 311
rect -2027 283 -1999 311
rect -1961 283 -1933 311
rect -1895 283 -1867 311
rect -1829 283 -1801 311
rect -1763 283 -1735 311
rect -1697 283 -1669 311
rect -1631 283 -1603 311
rect -1565 283 -1537 311
rect -1499 283 -1471 311
rect -1433 283 -1405 311
rect -1367 283 -1339 311
rect -1301 283 -1273 311
rect -1235 283 -1207 311
rect -1169 283 -1141 311
rect -1103 283 -1075 311
rect -1037 283 -1009 311
rect -971 283 -943 311
rect -905 283 -877 311
rect -839 283 -811 311
rect -773 283 -745 311
rect -707 283 -679 311
rect -641 283 -613 311
rect -575 283 -547 311
rect -509 283 -481 311
rect -443 283 -415 311
rect -377 283 -349 311
rect -311 283 -283 311
rect -245 283 -217 311
rect -179 283 -151 311
rect -113 283 -85 311
rect -47 283 -19 311
rect 19 283 47 311
rect 85 283 113 311
rect 151 283 179 311
rect 217 283 245 311
rect 283 283 311 311
rect 349 283 377 311
rect 415 283 443 311
rect 481 283 509 311
rect 547 283 575 311
rect 613 283 641 311
rect 679 283 707 311
rect 745 283 773 311
rect 811 283 839 311
rect 877 283 905 311
rect 943 283 971 311
rect 1009 283 1037 311
rect 1075 283 1103 311
rect 1141 283 1169 311
rect 1207 283 1235 311
rect 1273 283 1301 311
rect 1339 283 1367 311
rect 1405 283 1433 311
rect 1471 283 1499 311
rect 1537 283 1565 311
rect 1603 283 1631 311
rect 1669 283 1697 311
rect 1735 283 1763 311
rect 1801 283 1829 311
rect 1867 283 1895 311
rect 1933 283 1961 311
rect 1999 283 2027 311
rect 2065 283 2093 311
rect 2131 283 2159 311
rect 2197 283 2225 311
rect 2263 283 2291 311
rect 2329 283 2357 311
rect 2395 283 2423 311
rect 2461 283 2489 311
rect 2527 283 2555 311
rect 2593 283 2621 311
rect -2621 217 -2593 245
rect -2555 217 -2527 245
rect -2489 217 -2461 245
rect -2423 217 -2395 245
rect -2357 217 -2329 245
rect -2291 217 -2263 245
rect -2225 217 -2197 245
rect -2159 217 -2131 245
rect -2093 217 -2065 245
rect -2027 217 -1999 245
rect -1961 217 -1933 245
rect -1895 217 -1867 245
rect -1829 217 -1801 245
rect -1763 217 -1735 245
rect -1697 217 -1669 245
rect -1631 217 -1603 245
rect -1565 217 -1537 245
rect -1499 217 -1471 245
rect -1433 217 -1405 245
rect -1367 217 -1339 245
rect -1301 217 -1273 245
rect -1235 217 -1207 245
rect -1169 217 -1141 245
rect -1103 217 -1075 245
rect -1037 217 -1009 245
rect -971 217 -943 245
rect -905 217 -877 245
rect -839 217 -811 245
rect -773 217 -745 245
rect -707 217 -679 245
rect -641 217 -613 245
rect -575 217 -547 245
rect -509 217 -481 245
rect -443 217 -415 245
rect -377 217 -349 245
rect -311 217 -283 245
rect -245 217 -217 245
rect -179 217 -151 245
rect -113 217 -85 245
rect -47 217 -19 245
rect 19 217 47 245
rect 85 217 113 245
rect 151 217 179 245
rect 217 217 245 245
rect 283 217 311 245
rect 349 217 377 245
rect 415 217 443 245
rect 481 217 509 245
rect 547 217 575 245
rect 613 217 641 245
rect 679 217 707 245
rect 745 217 773 245
rect 811 217 839 245
rect 877 217 905 245
rect 943 217 971 245
rect 1009 217 1037 245
rect 1075 217 1103 245
rect 1141 217 1169 245
rect 1207 217 1235 245
rect 1273 217 1301 245
rect 1339 217 1367 245
rect 1405 217 1433 245
rect 1471 217 1499 245
rect 1537 217 1565 245
rect 1603 217 1631 245
rect 1669 217 1697 245
rect 1735 217 1763 245
rect 1801 217 1829 245
rect 1867 217 1895 245
rect 1933 217 1961 245
rect 1999 217 2027 245
rect 2065 217 2093 245
rect 2131 217 2159 245
rect 2197 217 2225 245
rect 2263 217 2291 245
rect 2329 217 2357 245
rect 2395 217 2423 245
rect 2461 217 2489 245
rect 2527 217 2555 245
rect 2593 217 2621 245
rect -2621 151 -2593 179
rect -2555 151 -2527 179
rect -2489 151 -2461 179
rect -2423 151 -2395 179
rect -2357 151 -2329 179
rect -2291 151 -2263 179
rect -2225 151 -2197 179
rect -2159 151 -2131 179
rect -2093 151 -2065 179
rect -2027 151 -1999 179
rect -1961 151 -1933 179
rect -1895 151 -1867 179
rect -1829 151 -1801 179
rect -1763 151 -1735 179
rect -1697 151 -1669 179
rect -1631 151 -1603 179
rect -1565 151 -1537 179
rect -1499 151 -1471 179
rect -1433 151 -1405 179
rect -1367 151 -1339 179
rect -1301 151 -1273 179
rect -1235 151 -1207 179
rect -1169 151 -1141 179
rect -1103 151 -1075 179
rect -1037 151 -1009 179
rect -971 151 -943 179
rect -905 151 -877 179
rect -839 151 -811 179
rect -773 151 -745 179
rect -707 151 -679 179
rect -641 151 -613 179
rect -575 151 -547 179
rect -509 151 -481 179
rect -443 151 -415 179
rect -377 151 -349 179
rect -311 151 -283 179
rect -245 151 -217 179
rect -179 151 -151 179
rect -113 151 -85 179
rect -47 151 -19 179
rect 19 151 47 179
rect 85 151 113 179
rect 151 151 179 179
rect 217 151 245 179
rect 283 151 311 179
rect 349 151 377 179
rect 415 151 443 179
rect 481 151 509 179
rect 547 151 575 179
rect 613 151 641 179
rect 679 151 707 179
rect 745 151 773 179
rect 811 151 839 179
rect 877 151 905 179
rect 943 151 971 179
rect 1009 151 1037 179
rect 1075 151 1103 179
rect 1141 151 1169 179
rect 1207 151 1235 179
rect 1273 151 1301 179
rect 1339 151 1367 179
rect 1405 151 1433 179
rect 1471 151 1499 179
rect 1537 151 1565 179
rect 1603 151 1631 179
rect 1669 151 1697 179
rect 1735 151 1763 179
rect 1801 151 1829 179
rect 1867 151 1895 179
rect 1933 151 1961 179
rect 1999 151 2027 179
rect 2065 151 2093 179
rect 2131 151 2159 179
rect 2197 151 2225 179
rect 2263 151 2291 179
rect 2329 151 2357 179
rect 2395 151 2423 179
rect 2461 151 2489 179
rect 2527 151 2555 179
rect 2593 151 2621 179
rect -2621 85 -2593 113
rect -2555 85 -2527 113
rect -2489 85 -2461 113
rect -2423 85 -2395 113
rect -2357 85 -2329 113
rect -2291 85 -2263 113
rect -2225 85 -2197 113
rect -2159 85 -2131 113
rect -2093 85 -2065 113
rect -2027 85 -1999 113
rect -1961 85 -1933 113
rect -1895 85 -1867 113
rect -1829 85 -1801 113
rect -1763 85 -1735 113
rect -1697 85 -1669 113
rect -1631 85 -1603 113
rect -1565 85 -1537 113
rect -1499 85 -1471 113
rect -1433 85 -1405 113
rect -1367 85 -1339 113
rect -1301 85 -1273 113
rect -1235 85 -1207 113
rect -1169 85 -1141 113
rect -1103 85 -1075 113
rect -1037 85 -1009 113
rect -971 85 -943 113
rect -905 85 -877 113
rect -839 85 -811 113
rect -773 85 -745 113
rect -707 85 -679 113
rect -641 85 -613 113
rect -575 85 -547 113
rect -509 85 -481 113
rect -443 85 -415 113
rect -377 85 -349 113
rect -311 85 -283 113
rect -245 85 -217 113
rect -179 85 -151 113
rect -113 85 -85 113
rect -47 85 -19 113
rect 19 85 47 113
rect 85 85 113 113
rect 151 85 179 113
rect 217 85 245 113
rect 283 85 311 113
rect 349 85 377 113
rect 415 85 443 113
rect 481 85 509 113
rect 547 85 575 113
rect 613 85 641 113
rect 679 85 707 113
rect 745 85 773 113
rect 811 85 839 113
rect 877 85 905 113
rect 943 85 971 113
rect 1009 85 1037 113
rect 1075 85 1103 113
rect 1141 85 1169 113
rect 1207 85 1235 113
rect 1273 85 1301 113
rect 1339 85 1367 113
rect 1405 85 1433 113
rect 1471 85 1499 113
rect 1537 85 1565 113
rect 1603 85 1631 113
rect 1669 85 1697 113
rect 1735 85 1763 113
rect 1801 85 1829 113
rect 1867 85 1895 113
rect 1933 85 1961 113
rect 1999 85 2027 113
rect 2065 85 2093 113
rect 2131 85 2159 113
rect 2197 85 2225 113
rect 2263 85 2291 113
rect 2329 85 2357 113
rect 2395 85 2423 113
rect 2461 85 2489 113
rect 2527 85 2555 113
rect 2593 85 2621 113
rect -2621 19 -2593 47
rect -2555 19 -2527 47
rect -2489 19 -2461 47
rect -2423 19 -2395 47
rect -2357 19 -2329 47
rect -2291 19 -2263 47
rect -2225 19 -2197 47
rect -2159 19 -2131 47
rect -2093 19 -2065 47
rect -2027 19 -1999 47
rect -1961 19 -1933 47
rect -1895 19 -1867 47
rect -1829 19 -1801 47
rect -1763 19 -1735 47
rect -1697 19 -1669 47
rect -1631 19 -1603 47
rect -1565 19 -1537 47
rect -1499 19 -1471 47
rect -1433 19 -1405 47
rect -1367 19 -1339 47
rect -1301 19 -1273 47
rect -1235 19 -1207 47
rect -1169 19 -1141 47
rect -1103 19 -1075 47
rect -1037 19 -1009 47
rect -971 19 -943 47
rect -905 19 -877 47
rect -839 19 -811 47
rect -773 19 -745 47
rect -707 19 -679 47
rect -641 19 -613 47
rect -575 19 -547 47
rect -509 19 -481 47
rect -443 19 -415 47
rect -377 19 -349 47
rect -311 19 -283 47
rect -245 19 -217 47
rect -179 19 -151 47
rect -113 19 -85 47
rect -47 19 -19 47
rect 19 19 47 47
rect 85 19 113 47
rect 151 19 179 47
rect 217 19 245 47
rect 283 19 311 47
rect 349 19 377 47
rect 415 19 443 47
rect 481 19 509 47
rect 547 19 575 47
rect 613 19 641 47
rect 679 19 707 47
rect 745 19 773 47
rect 811 19 839 47
rect 877 19 905 47
rect 943 19 971 47
rect 1009 19 1037 47
rect 1075 19 1103 47
rect 1141 19 1169 47
rect 1207 19 1235 47
rect 1273 19 1301 47
rect 1339 19 1367 47
rect 1405 19 1433 47
rect 1471 19 1499 47
rect 1537 19 1565 47
rect 1603 19 1631 47
rect 1669 19 1697 47
rect 1735 19 1763 47
rect 1801 19 1829 47
rect 1867 19 1895 47
rect 1933 19 1961 47
rect 1999 19 2027 47
rect 2065 19 2093 47
rect 2131 19 2159 47
rect 2197 19 2225 47
rect 2263 19 2291 47
rect 2329 19 2357 47
rect 2395 19 2423 47
rect 2461 19 2489 47
rect 2527 19 2555 47
rect 2593 19 2621 47
rect -2621 -47 -2593 -19
rect -2555 -47 -2527 -19
rect -2489 -47 -2461 -19
rect -2423 -47 -2395 -19
rect -2357 -47 -2329 -19
rect -2291 -47 -2263 -19
rect -2225 -47 -2197 -19
rect -2159 -47 -2131 -19
rect -2093 -47 -2065 -19
rect -2027 -47 -1999 -19
rect -1961 -47 -1933 -19
rect -1895 -47 -1867 -19
rect -1829 -47 -1801 -19
rect -1763 -47 -1735 -19
rect -1697 -47 -1669 -19
rect -1631 -47 -1603 -19
rect -1565 -47 -1537 -19
rect -1499 -47 -1471 -19
rect -1433 -47 -1405 -19
rect -1367 -47 -1339 -19
rect -1301 -47 -1273 -19
rect -1235 -47 -1207 -19
rect -1169 -47 -1141 -19
rect -1103 -47 -1075 -19
rect -1037 -47 -1009 -19
rect -971 -47 -943 -19
rect -905 -47 -877 -19
rect -839 -47 -811 -19
rect -773 -47 -745 -19
rect -707 -47 -679 -19
rect -641 -47 -613 -19
rect -575 -47 -547 -19
rect -509 -47 -481 -19
rect -443 -47 -415 -19
rect -377 -47 -349 -19
rect -311 -47 -283 -19
rect -245 -47 -217 -19
rect -179 -47 -151 -19
rect -113 -47 -85 -19
rect -47 -47 -19 -19
rect 19 -47 47 -19
rect 85 -47 113 -19
rect 151 -47 179 -19
rect 217 -47 245 -19
rect 283 -47 311 -19
rect 349 -47 377 -19
rect 415 -47 443 -19
rect 481 -47 509 -19
rect 547 -47 575 -19
rect 613 -47 641 -19
rect 679 -47 707 -19
rect 745 -47 773 -19
rect 811 -47 839 -19
rect 877 -47 905 -19
rect 943 -47 971 -19
rect 1009 -47 1037 -19
rect 1075 -47 1103 -19
rect 1141 -47 1169 -19
rect 1207 -47 1235 -19
rect 1273 -47 1301 -19
rect 1339 -47 1367 -19
rect 1405 -47 1433 -19
rect 1471 -47 1499 -19
rect 1537 -47 1565 -19
rect 1603 -47 1631 -19
rect 1669 -47 1697 -19
rect 1735 -47 1763 -19
rect 1801 -47 1829 -19
rect 1867 -47 1895 -19
rect 1933 -47 1961 -19
rect 1999 -47 2027 -19
rect 2065 -47 2093 -19
rect 2131 -47 2159 -19
rect 2197 -47 2225 -19
rect 2263 -47 2291 -19
rect 2329 -47 2357 -19
rect 2395 -47 2423 -19
rect 2461 -47 2489 -19
rect 2527 -47 2555 -19
rect 2593 -47 2621 -19
rect -2621 -113 -2593 -85
rect -2555 -113 -2527 -85
rect -2489 -113 -2461 -85
rect -2423 -113 -2395 -85
rect -2357 -113 -2329 -85
rect -2291 -113 -2263 -85
rect -2225 -113 -2197 -85
rect -2159 -113 -2131 -85
rect -2093 -113 -2065 -85
rect -2027 -113 -1999 -85
rect -1961 -113 -1933 -85
rect -1895 -113 -1867 -85
rect -1829 -113 -1801 -85
rect -1763 -113 -1735 -85
rect -1697 -113 -1669 -85
rect -1631 -113 -1603 -85
rect -1565 -113 -1537 -85
rect -1499 -113 -1471 -85
rect -1433 -113 -1405 -85
rect -1367 -113 -1339 -85
rect -1301 -113 -1273 -85
rect -1235 -113 -1207 -85
rect -1169 -113 -1141 -85
rect -1103 -113 -1075 -85
rect -1037 -113 -1009 -85
rect -971 -113 -943 -85
rect -905 -113 -877 -85
rect -839 -113 -811 -85
rect -773 -113 -745 -85
rect -707 -113 -679 -85
rect -641 -113 -613 -85
rect -575 -113 -547 -85
rect -509 -113 -481 -85
rect -443 -113 -415 -85
rect -377 -113 -349 -85
rect -311 -113 -283 -85
rect -245 -113 -217 -85
rect -179 -113 -151 -85
rect -113 -113 -85 -85
rect -47 -113 -19 -85
rect 19 -113 47 -85
rect 85 -113 113 -85
rect 151 -113 179 -85
rect 217 -113 245 -85
rect 283 -113 311 -85
rect 349 -113 377 -85
rect 415 -113 443 -85
rect 481 -113 509 -85
rect 547 -113 575 -85
rect 613 -113 641 -85
rect 679 -113 707 -85
rect 745 -113 773 -85
rect 811 -113 839 -85
rect 877 -113 905 -85
rect 943 -113 971 -85
rect 1009 -113 1037 -85
rect 1075 -113 1103 -85
rect 1141 -113 1169 -85
rect 1207 -113 1235 -85
rect 1273 -113 1301 -85
rect 1339 -113 1367 -85
rect 1405 -113 1433 -85
rect 1471 -113 1499 -85
rect 1537 -113 1565 -85
rect 1603 -113 1631 -85
rect 1669 -113 1697 -85
rect 1735 -113 1763 -85
rect 1801 -113 1829 -85
rect 1867 -113 1895 -85
rect 1933 -113 1961 -85
rect 1999 -113 2027 -85
rect 2065 -113 2093 -85
rect 2131 -113 2159 -85
rect 2197 -113 2225 -85
rect 2263 -113 2291 -85
rect 2329 -113 2357 -85
rect 2395 -113 2423 -85
rect 2461 -113 2489 -85
rect 2527 -113 2555 -85
rect 2593 -113 2621 -85
rect -2621 -179 -2593 -151
rect -2555 -179 -2527 -151
rect -2489 -179 -2461 -151
rect -2423 -179 -2395 -151
rect -2357 -179 -2329 -151
rect -2291 -179 -2263 -151
rect -2225 -179 -2197 -151
rect -2159 -179 -2131 -151
rect -2093 -179 -2065 -151
rect -2027 -179 -1999 -151
rect -1961 -179 -1933 -151
rect -1895 -179 -1867 -151
rect -1829 -179 -1801 -151
rect -1763 -179 -1735 -151
rect -1697 -179 -1669 -151
rect -1631 -179 -1603 -151
rect -1565 -179 -1537 -151
rect -1499 -179 -1471 -151
rect -1433 -179 -1405 -151
rect -1367 -179 -1339 -151
rect -1301 -179 -1273 -151
rect -1235 -179 -1207 -151
rect -1169 -179 -1141 -151
rect -1103 -179 -1075 -151
rect -1037 -179 -1009 -151
rect -971 -179 -943 -151
rect -905 -179 -877 -151
rect -839 -179 -811 -151
rect -773 -179 -745 -151
rect -707 -179 -679 -151
rect -641 -179 -613 -151
rect -575 -179 -547 -151
rect -509 -179 -481 -151
rect -443 -179 -415 -151
rect -377 -179 -349 -151
rect -311 -179 -283 -151
rect -245 -179 -217 -151
rect -179 -179 -151 -151
rect -113 -179 -85 -151
rect -47 -179 -19 -151
rect 19 -179 47 -151
rect 85 -179 113 -151
rect 151 -179 179 -151
rect 217 -179 245 -151
rect 283 -179 311 -151
rect 349 -179 377 -151
rect 415 -179 443 -151
rect 481 -179 509 -151
rect 547 -179 575 -151
rect 613 -179 641 -151
rect 679 -179 707 -151
rect 745 -179 773 -151
rect 811 -179 839 -151
rect 877 -179 905 -151
rect 943 -179 971 -151
rect 1009 -179 1037 -151
rect 1075 -179 1103 -151
rect 1141 -179 1169 -151
rect 1207 -179 1235 -151
rect 1273 -179 1301 -151
rect 1339 -179 1367 -151
rect 1405 -179 1433 -151
rect 1471 -179 1499 -151
rect 1537 -179 1565 -151
rect 1603 -179 1631 -151
rect 1669 -179 1697 -151
rect 1735 -179 1763 -151
rect 1801 -179 1829 -151
rect 1867 -179 1895 -151
rect 1933 -179 1961 -151
rect 1999 -179 2027 -151
rect 2065 -179 2093 -151
rect 2131 -179 2159 -151
rect 2197 -179 2225 -151
rect 2263 -179 2291 -151
rect 2329 -179 2357 -151
rect 2395 -179 2423 -151
rect 2461 -179 2489 -151
rect 2527 -179 2555 -151
rect 2593 -179 2621 -151
rect -2621 -245 -2593 -217
rect -2555 -245 -2527 -217
rect -2489 -245 -2461 -217
rect -2423 -245 -2395 -217
rect -2357 -245 -2329 -217
rect -2291 -245 -2263 -217
rect -2225 -245 -2197 -217
rect -2159 -245 -2131 -217
rect -2093 -245 -2065 -217
rect -2027 -245 -1999 -217
rect -1961 -245 -1933 -217
rect -1895 -245 -1867 -217
rect -1829 -245 -1801 -217
rect -1763 -245 -1735 -217
rect -1697 -245 -1669 -217
rect -1631 -245 -1603 -217
rect -1565 -245 -1537 -217
rect -1499 -245 -1471 -217
rect -1433 -245 -1405 -217
rect -1367 -245 -1339 -217
rect -1301 -245 -1273 -217
rect -1235 -245 -1207 -217
rect -1169 -245 -1141 -217
rect -1103 -245 -1075 -217
rect -1037 -245 -1009 -217
rect -971 -245 -943 -217
rect -905 -245 -877 -217
rect -839 -245 -811 -217
rect -773 -245 -745 -217
rect -707 -245 -679 -217
rect -641 -245 -613 -217
rect -575 -245 -547 -217
rect -509 -245 -481 -217
rect -443 -245 -415 -217
rect -377 -245 -349 -217
rect -311 -245 -283 -217
rect -245 -245 -217 -217
rect -179 -245 -151 -217
rect -113 -245 -85 -217
rect -47 -245 -19 -217
rect 19 -245 47 -217
rect 85 -245 113 -217
rect 151 -245 179 -217
rect 217 -245 245 -217
rect 283 -245 311 -217
rect 349 -245 377 -217
rect 415 -245 443 -217
rect 481 -245 509 -217
rect 547 -245 575 -217
rect 613 -245 641 -217
rect 679 -245 707 -217
rect 745 -245 773 -217
rect 811 -245 839 -217
rect 877 -245 905 -217
rect 943 -245 971 -217
rect 1009 -245 1037 -217
rect 1075 -245 1103 -217
rect 1141 -245 1169 -217
rect 1207 -245 1235 -217
rect 1273 -245 1301 -217
rect 1339 -245 1367 -217
rect 1405 -245 1433 -217
rect 1471 -245 1499 -217
rect 1537 -245 1565 -217
rect 1603 -245 1631 -217
rect 1669 -245 1697 -217
rect 1735 -245 1763 -217
rect 1801 -245 1829 -217
rect 1867 -245 1895 -217
rect 1933 -245 1961 -217
rect 1999 -245 2027 -217
rect 2065 -245 2093 -217
rect 2131 -245 2159 -217
rect 2197 -245 2225 -217
rect 2263 -245 2291 -217
rect 2329 -245 2357 -217
rect 2395 -245 2423 -217
rect 2461 -245 2489 -217
rect 2527 -245 2555 -217
rect 2593 -245 2621 -217
rect -2621 -311 -2593 -283
rect -2555 -311 -2527 -283
rect -2489 -311 -2461 -283
rect -2423 -311 -2395 -283
rect -2357 -311 -2329 -283
rect -2291 -311 -2263 -283
rect -2225 -311 -2197 -283
rect -2159 -311 -2131 -283
rect -2093 -311 -2065 -283
rect -2027 -311 -1999 -283
rect -1961 -311 -1933 -283
rect -1895 -311 -1867 -283
rect -1829 -311 -1801 -283
rect -1763 -311 -1735 -283
rect -1697 -311 -1669 -283
rect -1631 -311 -1603 -283
rect -1565 -311 -1537 -283
rect -1499 -311 -1471 -283
rect -1433 -311 -1405 -283
rect -1367 -311 -1339 -283
rect -1301 -311 -1273 -283
rect -1235 -311 -1207 -283
rect -1169 -311 -1141 -283
rect -1103 -311 -1075 -283
rect -1037 -311 -1009 -283
rect -971 -311 -943 -283
rect -905 -311 -877 -283
rect -839 -311 -811 -283
rect -773 -311 -745 -283
rect -707 -311 -679 -283
rect -641 -311 -613 -283
rect -575 -311 -547 -283
rect -509 -311 -481 -283
rect -443 -311 -415 -283
rect -377 -311 -349 -283
rect -311 -311 -283 -283
rect -245 -311 -217 -283
rect -179 -311 -151 -283
rect -113 -311 -85 -283
rect -47 -311 -19 -283
rect 19 -311 47 -283
rect 85 -311 113 -283
rect 151 -311 179 -283
rect 217 -311 245 -283
rect 283 -311 311 -283
rect 349 -311 377 -283
rect 415 -311 443 -283
rect 481 -311 509 -283
rect 547 -311 575 -283
rect 613 -311 641 -283
rect 679 -311 707 -283
rect 745 -311 773 -283
rect 811 -311 839 -283
rect 877 -311 905 -283
rect 943 -311 971 -283
rect 1009 -311 1037 -283
rect 1075 -311 1103 -283
rect 1141 -311 1169 -283
rect 1207 -311 1235 -283
rect 1273 -311 1301 -283
rect 1339 -311 1367 -283
rect 1405 -311 1433 -283
rect 1471 -311 1499 -283
rect 1537 -311 1565 -283
rect 1603 -311 1631 -283
rect 1669 -311 1697 -283
rect 1735 -311 1763 -283
rect 1801 -311 1829 -283
rect 1867 -311 1895 -283
rect 1933 -311 1961 -283
rect 1999 -311 2027 -283
rect 2065 -311 2093 -283
rect 2131 -311 2159 -283
rect 2197 -311 2225 -283
rect 2263 -311 2291 -283
rect 2329 -311 2357 -283
rect 2395 -311 2423 -283
rect 2461 -311 2489 -283
rect 2527 -311 2555 -283
rect 2593 -311 2621 -283
rect -2621 -377 -2593 -349
rect -2555 -377 -2527 -349
rect -2489 -377 -2461 -349
rect -2423 -377 -2395 -349
rect -2357 -377 -2329 -349
rect -2291 -377 -2263 -349
rect -2225 -377 -2197 -349
rect -2159 -377 -2131 -349
rect -2093 -377 -2065 -349
rect -2027 -377 -1999 -349
rect -1961 -377 -1933 -349
rect -1895 -377 -1867 -349
rect -1829 -377 -1801 -349
rect -1763 -377 -1735 -349
rect -1697 -377 -1669 -349
rect -1631 -377 -1603 -349
rect -1565 -377 -1537 -349
rect -1499 -377 -1471 -349
rect -1433 -377 -1405 -349
rect -1367 -377 -1339 -349
rect -1301 -377 -1273 -349
rect -1235 -377 -1207 -349
rect -1169 -377 -1141 -349
rect -1103 -377 -1075 -349
rect -1037 -377 -1009 -349
rect -971 -377 -943 -349
rect -905 -377 -877 -349
rect -839 -377 -811 -349
rect -773 -377 -745 -349
rect -707 -377 -679 -349
rect -641 -377 -613 -349
rect -575 -377 -547 -349
rect -509 -377 -481 -349
rect -443 -377 -415 -349
rect -377 -377 -349 -349
rect -311 -377 -283 -349
rect -245 -377 -217 -349
rect -179 -377 -151 -349
rect -113 -377 -85 -349
rect -47 -377 -19 -349
rect 19 -377 47 -349
rect 85 -377 113 -349
rect 151 -377 179 -349
rect 217 -377 245 -349
rect 283 -377 311 -349
rect 349 -377 377 -349
rect 415 -377 443 -349
rect 481 -377 509 -349
rect 547 -377 575 -349
rect 613 -377 641 -349
rect 679 -377 707 -349
rect 745 -377 773 -349
rect 811 -377 839 -349
rect 877 -377 905 -349
rect 943 -377 971 -349
rect 1009 -377 1037 -349
rect 1075 -377 1103 -349
rect 1141 -377 1169 -349
rect 1207 -377 1235 -349
rect 1273 -377 1301 -349
rect 1339 -377 1367 -349
rect 1405 -377 1433 -349
rect 1471 -377 1499 -349
rect 1537 -377 1565 -349
rect 1603 -377 1631 -349
rect 1669 -377 1697 -349
rect 1735 -377 1763 -349
rect 1801 -377 1829 -349
rect 1867 -377 1895 -349
rect 1933 -377 1961 -349
rect 1999 -377 2027 -349
rect 2065 -377 2093 -349
rect 2131 -377 2159 -349
rect 2197 -377 2225 -349
rect 2263 -377 2291 -349
rect 2329 -377 2357 -349
rect 2395 -377 2423 -349
rect 2461 -377 2489 -349
rect 2527 -377 2555 -349
rect 2593 -377 2621 -349
<< metal3 >>
rect -2626 377 2626 382
rect -2626 349 -2621 377
rect -2593 349 -2555 377
rect -2527 349 -2489 377
rect -2461 349 -2423 377
rect -2395 349 -2357 377
rect -2329 349 -2291 377
rect -2263 349 -2225 377
rect -2197 349 -2159 377
rect -2131 349 -2093 377
rect -2065 349 -2027 377
rect -1999 349 -1961 377
rect -1933 349 -1895 377
rect -1867 349 -1829 377
rect -1801 349 -1763 377
rect -1735 349 -1697 377
rect -1669 349 -1631 377
rect -1603 349 -1565 377
rect -1537 349 -1499 377
rect -1471 349 -1433 377
rect -1405 349 -1367 377
rect -1339 349 -1301 377
rect -1273 349 -1235 377
rect -1207 349 -1169 377
rect -1141 349 -1103 377
rect -1075 349 -1037 377
rect -1009 349 -971 377
rect -943 349 -905 377
rect -877 349 -839 377
rect -811 349 -773 377
rect -745 349 -707 377
rect -679 349 -641 377
rect -613 349 -575 377
rect -547 349 -509 377
rect -481 349 -443 377
rect -415 349 -377 377
rect -349 349 -311 377
rect -283 349 -245 377
rect -217 349 -179 377
rect -151 349 -113 377
rect -85 349 -47 377
rect -19 349 19 377
rect 47 349 85 377
rect 113 349 151 377
rect 179 349 217 377
rect 245 349 283 377
rect 311 349 349 377
rect 377 349 415 377
rect 443 349 481 377
rect 509 349 547 377
rect 575 349 613 377
rect 641 349 679 377
rect 707 349 745 377
rect 773 349 811 377
rect 839 349 877 377
rect 905 349 943 377
rect 971 349 1009 377
rect 1037 349 1075 377
rect 1103 349 1141 377
rect 1169 349 1207 377
rect 1235 349 1273 377
rect 1301 349 1339 377
rect 1367 349 1405 377
rect 1433 349 1471 377
rect 1499 349 1537 377
rect 1565 349 1603 377
rect 1631 349 1669 377
rect 1697 349 1735 377
rect 1763 349 1801 377
rect 1829 349 1867 377
rect 1895 349 1933 377
rect 1961 349 1999 377
rect 2027 349 2065 377
rect 2093 349 2131 377
rect 2159 349 2197 377
rect 2225 349 2263 377
rect 2291 349 2329 377
rect 2357 349 2395 377
rect 2423 349 2461 377
rect 2489 349 2527 377
rect 2555 349 2593 377
rect 2621 349 2626 377
rect -2626 311 2626 349
rect -2626 283 -2621 311
rect -2593 283 -2555 311
rect -2527 283 -2489 311
rect -2461 283 -2423 311
rect -2395 283 -2357 311
rect -2329 283 -2291 311
rect -2263 283 -2225 311
rect -2197 283 -2159 311
rect -2131 283 -2093 311
rect -2065 283 -2027 311
rect -1999 283 -1961 311
rect -1933 283 -1895 311
rect -1867 283 -1829 311
rect -1801 283 -1763 311
rect -1735 283 -1697 311
rect -1669 283 -1631 311
rect -1603 283 -1565 311
rect -1537 283 -1499 311
rect -1471 283 -1433 311
rect -1405 283 -1367 311
rect -1339 283 -1301 311
rect -1273 283 -1235 311
rect -1207 283 -1169 311
rect -1141 283 -1103 311
rect -1075 283 -1037 311
rect -1009 283 -971 311
rect -943 283 -905 311
rect -877 283 -839 311
rect -811 283 -773 311
rect -745 283 -707 311
rect -679 283 -641 311
rect -613 283 -575 311
rect -547 283 -509 311
rect -481 283 -443 311
rect -415 283 -377 311
rect -349 283 -311 311
rect -283 283 -245 311
rect -217 283 -179 311
rect -151 283 -113 311
rect -85 283 -47 311
rect -19 283 19 311
rect 47 283 85 311
rect 113 283 151 311
rect 179 283 217 311
rect 245 283 283 311
rect 311 283 349 311
rect 377 283 415 311
rect 443 283 481 311
rect 509 283 547 311
rect 575 283 613 311
rect 641 283 679 311
rect 707 283 745 311
rect 773 283 811 311
rect 839 283 877 311
rect 905 283 943 311
rect 971 283 1009 311
rect 1037 283 1075 311
rect 1103 283 1141 311
rect 1169 283 1207 311
rect 1235 283 1273 311
rect 1301 283 1339 311
rect 1367 283 1405 311
rect 1433 283 1471 311
rect 1499 283 1537 311
rect 1565 283 1603 311
rect 1631 283 1669 311
rect 1697 283 1735 311
rect 1763 283 1801 311
rect 1829 283 1867 311
rect 1895 283 1933 311
rect 1961 283 1999 311
rect 2027 283 2065 311
rect 2093 283 2131 311
rect 2159 283 2197 311
rect 2225 283 2263 311
rect 2291 283 2329 311
rect 2357 283 2395 311
rect 2423 283 2461 311
rect 2489 283 2527 311
rect 2555 283 2593 311
rect 2621 283 2626 311
rect -2626 245 2626 283
rect -2626 217 -2621 245
rect -2593 217 -2555 245
rect -2527 217 -2489 245
rect -2461 217 -2423 245
rect -2395 217 -2357 245
rect -2329 217 -2291 245
rect -2263 217 -2225 245
rect -2197 217 -2159 245
rect -2131 217 -2093 245
rect -2065 217 -2027 245
rect -1999 217 -1961 245
rect -1933 217 -1895 245
rect -1867 217 -1829 245
rect -1801 217 -1763 245
rect -1735 217 -1697 245
rect -1669 217 -1631 245
rect -1603 217 -1565 245
rect -1537 217 -1499 245
rect -1471 217 -1433 245
rect -1405 217 -1367 245
rect -1339 217 -1301 245
rect -1273 217 -1235 245
rect -1207 217 -1169 245
rect -1141 217 -1103 245
rect -1075 217 -1037 245
rect -1009 217 -971 245
rect -943 217 -905 245
rect -877 217 -839 245
rect -811 217 -773 245
rect -745 217 -707 245
rect -679 217 -641 245
rect -613 217 -575 245
rect -547 217 -509 245
rect -481 217 -443 245
rect -415 217 -377 245
rect -349 217 -311 245
rect -283 217 -245 245
rect -217 217 -179 245
rect -151 217 -113 245
rect -85 217 -47 245
rect -19 217 19 245
rect 47 217 85 245
rect 113 217 151 245
rect 179 217 217 245
rect 245 217 283 245
rect 311 217 349 245
rect 377 217 415 245
rect 443 217 481 245
rect 509 217 547 245
rect 575 217 613 245
rect 641 217 679 245
rect 707 217 745 245
rect 773 217 811 245
rect 839 217 877 245
rect 905 217 943 245
rect 971 217 1009 245
rect 1037 217 1075 245
rect 1103 217 1141 245
rect 1169 217 1207 245
rect 1235 217 1273 245
rect 1301 217 1339 245
rect 1367 217 1405 245
rect 1433 217 1471 245
rect 1499 217 1537 245
rect 1565 217 1603 245
rect 1631 217 1669 245
rect 1697 217 1735 245
rect 1763 217 1801 245
rect 1829 217 1867 245
rect 1895 217 1933 245
rect 1961 217 1999 245
rect 2027 217 2065 245
rect 2093 217 2131 245
rect 2159 217 2197 245
rect 2225 217 2263 245
rect 2291 217 2329 245
rect 2357 217 2395 245
rect 2423 217 2461 245
rect 2489 217 2527 245
rect 2555 217 2593 245
rect 2621 217 2626 245
rect -2626 179 2626 217
rect -2626 151 -2621 179
rect -2593 151 -2555 179
rect -2527 151 -2489 179
rect -2461 151 -2423 179
rect -2395 151 -2357 179
rect -2329 151 -2291 179
rect -2263 151 -2225 179
rect -2197 151 -2159 179
rect -2131 151 -2093 179
rect -2065 151 -2027 179
rect -1999 151 -1961 179
rect -1933 151 -1895 179
rect -1867 151 -1829 179
rect -1801 151 -1763 179
rect -1735 151 -1697 179
rect -1669 151 -1631 179
rect -1603 151 -1565 179
rect -1537 151 -1499 179
rect -1471 151 -1433 179
rect -1405 151 -1367 179
rect -1339 151 -1301 179
rect -1273 151 -1235 179
rect -1207 151 -1169 179
rect -1141 151 -1103 179
rect -1075 151 -1037 179
rect -1009 151 -971 179
rect -943 151 -905 179
rect -877 151 -839 179
rect -811 151 -773 179
rect -745 151 -707 179
rect -679 151 -641 179
rect -613 151 -575 179
rect -547 151 -509 179
rect -481 151 -443 179
rect -415 151 -377 179
rect -349 151 -311 179
rect -283 151 -245 179
rect -217 151 -179 179
rect -151 151 -113 179
rect -85 151 -47 179
rect -19 151 19 179
rect 47 151 85 179
rect 113 151 151 179
rect 179 151 217 179
rect 245 151 283 179
rect 311 151 349 179
rect 377 151 415 179
rect 443 151 481 179
rect 509 151 547 179
rect 575 151 613 179
rect 641 151 679 179
rect 707 151 745 179
rect 773 151 811 179
rect 839 151 877 179
rect 905 151 943 179
rect 971 151 1009 179
rect 1037 151 1075 179
rect 1103 151 1141 179
rect 1169 151 1207 179
rect 1235 151 1273 179
rect 1301 151 1339 179
rect 1367 151 1405 179
rect 1433 151 1471 179
rect 1499 151 1537 179
rect 1565 151 1603 179
rect 1631 151 1669 179
rect 1697 151 1735 179
rect 1763 151 1801 179
rect 1829 151 1867 179
rect 1895 151 1933 179
rect 1961 151 1999 179
rect 2027 151 2065 179
rect 2093 151 2131 179
rect 2159 151 2197 179
rect 2225 151 2263 179
rect 2291 151 2329 179
rect 2357 151 2395 179
rect 2423 151 2461 179
rect 2489 151 2527 179
rect 2555 151 2593 179
rect 2621 151 2626 179
rect -2626 113 2626 151
rect -2626 85 -2621 113
rect -2593 85 -2555 113
rect -2527 85 -2489 113
rect -2461 85 -2423 113
rect -2395 85 -2357 113
rect -2329 85 -2291 113
rect -2263 85 -2225 113
rect -2197 85 -2159 113
rect -2131 85 -2093 113
rect -2065 85 -2027 113
rect -1999 85 -1961 113
rect -1933 85 -1895 113
rect -1867 85 -1829 113
rect -1801 85 -1763 113
rect -1735 85 -1697 113
rect -1669 85 -1631 113
rect -1603 85 -1565 113
rect -1537 85 -1499 113
rect -1471 85 -1433 113
rect -1405 85 -1367 113
rect -1339 85 -1301 113
rect -1273 85 -1235 113
rect -1207 85 -1169 113
rect -1141 85 -1103 113
rect -1075 85 -1037 113
rect -1009 85 -971 113
rect -943 85 -905 113
rect -877 85 -839 113
rect -811 85 -773 113
rect -745 85 -707 113
rect -679 85 -641 113
rect -613 85 -575 113
rect -547 85 -509 113
rect -481 85 -443 113
rect -415 85 -377 113
rect -349 85 -311 113
rect -283 85 -245 113
rect -217 85 -179 113
rect -151 85 -113 113
rect -85 85 -47 113
rect -19 85 19 113
rect 47 85 85 113
rect 113 85 151 113
rect 179 85 217 113
rect 245 85 283 113
rect 311 85 349 113
rect 377 85 415 113
rect 443 85 481 113
rect 509 85 547 113
rect 575 85 613 113
rect 641 85 679 113
rect 707 85 745 113
rect 773 85 811 113
rect 839 85 877 113
rect 905 85 943 113
rect 971 85 1009 113
rect 1037 85 1075 113
rect 1103 85 1141 113
rect 1169 85 1207 113
rect 1235 85 1273 113
rect 1301 85 1339 113
rect 1367 85 1405 113
rect 1433 85 1471 113
rect 1499 85 1537 113
rect 1565 85 1603 113
rect 1631 85 1669 113
rect 1697 85 1735 113
rect 1763 85 1801 113
rect 1829 85 1867 113
rect 1895 85 1933 113
rect 1961 85 1999 113
rect 2027 85 2065 113
rect 2093 85 2131 113
rect 2159 85 2197 113
rect 2225 85 2263 113
rect 2291 85 2329 113
rect 2357 85 2395 113
rect 2423 85 2461 113
rect 2489 85 2527 113
rect 2555 85 2593 113
rect 2621 85 2626 113
rect -2626 47 2626 85
rect -2626 19 -2621 47
rect -2593 19 -2555 47
rect -2527 19 -2489 47
rect -2461 19 -2423 47
rect -2395 19 -2357 47
rect -2329 19 -2291 47
rect -2263 19 -2225 47
rect -2197 19 -2159 47
rect -2131 19 -2093 47
rect -2065 19 -2027 47
rect -1999 19 -1961 47
rect -1933 19 -1895 47
rect -1867 19 -1829 47
rect -1801 19 -1763 47
rect -1735 19 -1697 47
rect -1669 19 -1631 47
rect -1603 19 -1565 47
rect -1537 19 -1499 47
rect -1471 19 -1433 47
rect -1405 19 -1367 47
rect -1339 19 -1301 47
rect -1273 19 -1235 47
rect -1207 19 -1169 47
rect -1141 19 -1103 47
rect -1075 19 -1037 47
rect -1009 19 -971 47
rect -943 19 -905 47
rect -877 19 -839 47
rect -811 19 -773 47
rect -745 19 -707 47
rect -679 19 -641 47
rect -613 19 -575 47
rect -547 19 -509 47
rect -481 19 -443 47
rect -415 19 -377 47
rect -349 19 -311 47
rect -283 19 -245 47
rect -217 19 -179 47
rect -151 19 -113 47
rect -85 19 -47 47
rect -19 19 19 47
rect 47 19 85 47
rect 113 19 151 47
rect 179 19 217 47
rect 245 19 283 47
rect 311 19 349 47
rect 377 19 415 47
rect 443 19 481 47
rect 509 19 547 47
rect 575 19 613 47
rect 641 19 679 47
rect 707 19 745 47
rect 773 19 811 47
rect 839 19 877 47
rect 905 19 943 47
rect 971 19 1009 47
rect 1037 19 1075 47
rect 1103 19 1141 47
rect 1169 19 1207 47
rect 1235 19 1273 47
rect 1301 19 1339 47
rect 1367 19 1405 47
rect 1433 19 1471 47
rect 1499 19 1537 47
rect 1565 19 1603 47
rect 1631 19 1669 47
rect 1697 19 1735 47
rect 1763 19 1801 47
rect 1829 19 1867 47
rect 1895 19 1933 47
rect 1961 19 1999 47
rect 2027 19 2065 47
rect 2093 19 2131 47
rect 2159 19 2197 47
rect 2225 19 2263 47
rect 2291 19 2329 47
rect 2357 19 2395 47
rect 2423 19 2461 47
rect 2489 19 2527 47
rect 2555 19 2593 47
rect 2621 19 2626 47
rect -2626 -19 2626 19
rect -2626 -47 -2621 -19
rect -2593 -47 -2555 -19
rect -2527 -47 -2489 -19
rect -2461 -47 -2423 -19
rect -2395 -47 -2357 -19
rect -2329 -47 -2291 -19
rect -2263 -47 -2225 -19
rect -2197 -47 -2159 -19
rect -2131 -47 -2093 -19
rect -2065 -47 -2027 -19
rect -1999 -47 -1961 -19
rect -1933 -47 -1895 -19
rect -1867 -47 -1829 -19
rect -1801 -47 -1763 -19
rect -1735 -47 -1697 -19
rect -1669 -47 -1631 -19
rect -1603 -47 -1565 -19
rect -1537 -47 -1499 -19
rect -1471 -47 -1433 -19
rect -1405 -47 -1367 -19
rect -1339 -47 -1301 -19
rect -1273 -47 -1235 -19
rect -1207 -47 -1169 -19
rect -1141 -47 -1103 -19
rect -1075 -47 -1037 -19
rect -1009 -47 -971 -19
rect -943 -47 -905 -19
rect -877 -47 -839 -19
rect -811 -47 -773 -19
rect -745 -47 -707 -19
rect -679 -47 -641 -19
rect -613 -47 -575 -19
rect -547 -47 -509 -19
rect -481 -47 -443 -19
rect -415 -47 -377 -19
rect -349 -47 -311 -19
rect -283 -47 -245 -19
rect -217 -47 -179 -19
rect -151 -47 -113 -19
rect -85 -47 -47 -19
rect -19 -47 19 -19
rect 47 -47 85 -19
rect 113 -47 151 -19
rect 179 -47 217 -19
rect 245 -47 283 -19
rect 311 -47 349 -19
rect 377 -47 415 -19
rect 443 -47 481 -19
rect 509 -47 547 -19
rect 575 -47 613 -19
rect 641 -47 679 -19
rect 707 -47 745 -19
rect 773 -47 811 -19
rect 839 -47 877 -19
rect 905 -47 943 -19
rect 971 -47 1009 -19
rect 1037 -47 1075 -19
rect 1103 -47 1141 -19
rect 1169 -47 1207 -19
rect 1235 -47 1273 -19
rect 1301 -47 1339 -19
rect 1367 -47 1405 -19
rect 1433 -47 1471 -19
rect 1499 -47 1537 -19
rect 1565 -47 1603 -19
rect 1631 -47 1669 -19
rect 1697 -47 1735 -19
rect 1763 -47 1801 -19
rect 1829 -47 1867 -19
rect 1895 -47 1933 -19
rect 1961 -47 1999 -19
rect 2027 -47 2065 -19
rect 2093 -47 2131 -19
rect 2159 -47 2197 -19
rect 2225 -47 2263 -19
rect 2291 -47 2329 -19
rect 2357 -47 2395 -19
rect 2423 -47 2461 -19
rect 2489 -47 2527 -19
rect 2555 -47 2593 -19
rect 2621 -47 2626 -19
rect -2626 -85 2626 -47
rect -2626 -113 -2621 -85
rect -2593 -113 -2555 -85
rect -2527 -113 -2489 -85
rect -2461 -113 -2423 -85
rect -2395 -113 -2357 -85
rect -2329 -113 -2291 -85
rect -2263 -113 -2225 -85
rect -2197 -113 -2159 -85
rect -2131 -113 -2093 -85
rect -2065 -113 -2027 -85
rect -1999 -113 -1961 -85
rect -1933 -113 -1895 -85
rect -1867 -113 -1829 -85
rect -1801 -113 -1763 -85
rect -1735 -113 -1697 -85
rect -1669 -113 -1631 -85
rect -1603 -113 -1565 -85
rect -1537 -113 -1499 -85
rect -1471 -113 -1433 -85
rect -1405 -113 -1367 -85
rect -1339 -113 -1301 -85
rect -1273 -113 -1235 -85
rect -1207 -113 -1169 -85
rect -1141 -113 -1103 -85
rect -1075 -113 -1037 -85
rect -1009 -113 -971 -85
rect -943 -113 -905 -85
rect -877 -113 -839 -85
rect -811 -113 -773 -85
rect -745 -113 -707 -85
rect -679 -113 -641 -85
rect -613 -113 -575 -85
rect -547 -113 -509 -85
rect -481 -113 -443 -85
rect -415 -113 -377 -85
rect -349 -113 -311 -85
rect -283 -113 -245 -85
rect -217 -113 -179 -85
rect -151 -113 -113 -85
rect -85 -113 -47 -85
rect -19 -113 19 -85
rect 47 -113 85 -85
rect 113 -113 151 -85
rect 179 -113 217 -85
rect 245 -113 283 -85
rect 311 -113 349 -85
rect 377 -113 415 -85
rect 443 -113 481 -85
rect 509 -113 547 -85
rect 575 -113 613 -85
rect 641 -113 679 -85
rect 707 -113 745 -85
rect 773 -113 811 -85
rect 839 -113 877 -85
rect 905 -113 943 -85
rect 971 -113 1009 -85
rect 1037 -113 1075 -85
rect 1103 -113 1141 -85
rect 1169 -113 1207 -85
rect 1235 -113 1273 -85
rect 1301 -113 1339 -85
rect 1367 -113 1405 -85
rect 1433 -113 1471 -85
rect 1499 -113 1537 -85
rect 1565 -113 1603 -85
rect 1631 -113 1669 -85
rect 1697 -113 1735 -85
rect 1763 -113 1801 -85
rect 1829 -113 1867 -85
rect 1895 -113 1933 -85
rect 1961 -113 1999 -85
rect 2027 -113 2065 -85
rect 2093 -113 2131 -85
rect 2159 -113 2197 -85
rect 2225 -113 2263 -85
rect 2291 -113 2329 -85
rect 2357 -113 2395 -85
rect 2423 -113 2461 -85
rect 2489 -113 2527 -85
rect 2555 -113 2593 -85
rect 2621 -113 2626 -85
rect -2626 -151 2626 -113
rect -2626 -179 -2621 -151
rect -2593 -179 -2555 -151
rect -2527 -179 -2489 -151
rect -2461 -179 -2423 -151
rect -2395 -179 -2357 -151
rect -2329 -179 -2291 -151
rect -2263 -179 -2225 -151
rect -2197 -179 -2159 -151
rect -2131 -179 -2093 -151
rect -2065 -179 -2027 -151
rect -1999 -179 -1961 -151
rect -1933 -179 -1895 -151
rect -1867 -179 -1829 -151
rect -1801 -179 -1763 -151
rect -1735 -179 -1697 -151
rect -1669 -179 -1631 -151
rect -1603 -179 -1565 -151
rect -1537 -179 -1499 -151
rect -1471 -179 -1433 -151
rect -1405 -179 -1367 -151
rect -1339 -179 -1301 -151
rect -1273 -179 -1235 -151
rect -1207 -179 -1169 -151
rect -1141 -179 -1103 -151
rect -1075 -179 -1037 -151
rect -1009 -179 -971 -151
rect -943 -179 -905 -151
rect -877 -179 -839 -151
rect -811 -179 -773 -151
rect -745 -179 -707 -151
rect -679 -179 -641 -151
rect -613 -179 -575 -151
rect -547 -179 -509 -151
rect -481 -179 -443 -151
rect -415 -179 -377 -151
rect -349 -179 -311 -151
rect -283 -179 -245 -151
rect -217 -179 -179 -151
rect -151 -179 -113 -151
rect -85 -179 -47 -151
rect -19 -179 19 -151
rect 47 -179 85 -151
rect 113 -179 151 -151
rect 179 -179 217 -151
rect 245 -179 283 -151
rect 311 -179 349 -151
rect 377 -179 415 -151
rect 443 -179 481 -151
rect 509 -179 547 -151
rect 575 -179 613 -151
rect 641 -179 679 -151
rect 707 -179 745 -151
rect 773 -179 811 -151
rect 839 -179 877 -151
rect 905 -179 943 -151
rect 971 -179 1009 -151
rect 1037 -179 1075 -151
rect 1103 -179 1141 -151
rect 1169 -179 1207 -151
rect 1235 -179 1273 -151
rect 1301 -179 1339 -151
rect 1367 -179 1405 -151
rect 1433 -179 1471 -151
rect 1499 -179 1537 -151
rect 1565 -179 1603 -151
rect 1631 -179 1669 -151
rect 1697 -179 1735 -151
rect 1763 -179 1801 -151
rect 1829 -179 1867 -151
rect 1895 -179 1933 -151
rect 1961 -179 1999 -151
rect 2027 -179 2065 -151
rect 2093 -179 2131 -151
rect 2159 -179 2197 -151
rect 2225 -179 2263 -151
rect 2291 -179 2329 -151
rect 2357 -179 2395 -151
rect 2423 -179 2461 -151
rect 2489 -179 2527 -151
rect 2555 -179 2593 -151
rect 2621 -179 2626 -151
rect -2626 -217 2626 -179
rect -2626 -245 -2621 -217
rect -2593 -245 -2555 -217
rect -2527 -245 -2489 -217
rect -2461 -245 -2423 -217
rect -2395 -245 -2357 -217
rect -2329 -245 -2291 -217
rect -2263 -245 -2225 -217
rect -2197 -245 -2159 -217
rect -2131 -245 -2093 -217
rect -2065 -245 -2027 -217
rect -1999 -245 -1961 -217
rect -1933 -245 -1895 -217
rect -1867 -245 -1829 -217
rect -1801 -245 -1763 -217
rect -1735 -245 -1697 -217
rect -1669 -245 -1631 -217
rect -1603 -245 -1565 -217
rect -1537 -245 -1499 -217
rect -1471 -245 -1433 -217
rect -1405 -245 -1367 -217
rect -1339 -245 -1301 -217
rect -1273 -245 -1235 -217
rect -1207 -245 -1169 -217
rect -1141 -245 -1103 -217
rect -1075 -245 -1037 -217
rect -1009 -245 -971 -217
rect -943 -245 -905 -217
rect -877 -245 -839 -217
rect -811 -245 -773 -217
rect -745 -245 -707 -217
rect -679 -245 -641 -217
rect -613 -245 -575 -217
rect -547 -245 -509 -217
rect -481 -245 -443 -217
rect -415 -245 -377 -217
rect -349 -245 -311 -217
rect -283 -245 -245 -217
rect -217 -245 -179 -217
rect -151 -245 -113 -217
rect -85 -245 -47 -217
rect -19 -245 19 -217
rect 47 -245 85 -217
rect 113 -245 151 -217
rect 179 -245 217 -217
rect 245 -245 283 -217
rect 311 -245 349 -217
rect 377 -245 415 -217
rect 443 -245 481 -217
rect 509 -245 547 -217
rect 575 -245 613 -217
rect 641 -245 679 -217
rect 707 -245 745 -217
rect 773 -245 811 -217
rect 839 -245 877 -217
rect 905 -245 943 -217
rect 971 -245 1009 -217
rect 1037 -245 1075 -217
rect 1103 -245 1141 -217
rect 1169 -245 1207 -217
rect 1235 -245 1273 -217
rect 1301 -245 1339 -217
rect 1367 -245 1405 -217
rect 1433 -245 1471 -217
rect 1499 -245 1537 -217
rect 1565 -245 1603 -217
rect 1631 -245 1669 -217
rect 1697 -245 1735 -217
rect 1763 -245 1801 -217
rect 1829 -245 1867 -217
rect 1895 -245 1933 -217
rect 1961 -245 1999 -217
rect 2027 -245 2065 -217
rect 2093 -245 2131 -217
rect 2159 -245 2197 -217
rect 2225 -245 2263 -217
rect 2291 -245 2329 -217
rect 2357 -245 2395 -217
rect 2423 -245 2461 -217
rect 2489 -245 2527 -217
rect 2555 -245 2593 -217
rect 2621 -245 2626 -217
rect -2626 -283 2626 -245
rect -2626 -311 -2621 -283
rect -2593 -311 -2555 -283
rect -2527 -311 -2489 -283
rect -2461 -311 -2423 -283
rect -2395 -311 -2357 -283
rect -2329 -311 -2291 -283
rect -2263 -311 -2225 -283
rect -2197 -311 -2159 -283
rect -2131 -311 -2093 -283
rect -2065 -311 -2027 -283
rect -1999 -311 -1961 -283
rect -1933 -311 -1895 -283
rect -1867 -311 -1829 -283
rect -1801 -311 -1763 -283
rect -1735 -311 -1697 -283
rect -1669 -311 -1631 -283
rect -1603 -311 -1565 -283
rect -1537 -311 -1499 -283
rect -1471 -311 -1433 -283
rect -1405 -311 -1367 -283
rect -1339 -311 -1301 -283
rect -1273 -311 -1235 -283
rect -1207 -311 -1169 -283
rect -1141 -311 -1103 -283
rect -1075 -311 -1037 -283
rect -1009 -311 -971 -283
rect -943 -311 -905 -283
rect -877 -311 -839 -283
rect -811 -311 -773 -283
rect -745 -311 -707 -283
rect -679 -311 -641 -283
rect -613 -311 -575 -283
rect -547 -311 -509 -283
rect -481 -311 -443 -283
rect -415 -311 -377 -283
rect -349 -311 -311 -283
rect -283 -311 -245 -283
rect -217 -311 -179 -283
rect -151 -311 -113 -283
rect -85 -311 -47 -283
rect -19 -311 19 -283
rect 47 -311 85 -283
rect 113 -311 151 -283
rect 179 -311 217 -283
rect 245 -311 283 -283
rect 311 -311 349 -283
rect 377 -311 415 -283
rect 443 -311 481 -283
rect 509 -311 547 -283
rect 575 -311 613 -283
rect 641 -311 679 -283
rect 707 -311 745 -283
rect 773 -311 811 -283
rect 839 -311 877 -283
rect 905 -311 943 -283
rect 971 -311 1009 -283
rect 1037 -311 1075 -283
rect 1103 -311 1141 -283
rect 1169 -311 1207 -283
rect 1235 -311 1273 -283
rect 1301 -311 1339 -283
rect 1367 -311 1405 -283
rect 1433 -311 1471 -283
rect 1499 -311 1537 -283
rect 1565 -311 1603 -283
rect 1631 -311 1669 -283
rect 1697 -311 1735 -283
rect 1763 -311 1801 -283
rect 1829 -311 1867 -283
rect 1895 -311 1933 -283
rect 1961 -311 1999 -283
rect 2027 -311 2065 -283
rect 2093 -311 2131 -283
rect 2159 -311 2197 -283
rect 2225 -311 2263 -283
rect 2291 -311 2329 -283
rect 2357 -311 2395 -283
rect 2423 -311 2461 -283
rect 2489 -311 2527 -283
rect 2555 -311 2593 -283
rect 2621 -311 2626 -283
rect -2626 -349 2626 -311
rect -2626 -377 -2621 -349
rect -2593 -377 -2555 -349
rect -2527 -377 -2489 -349
rect -2461 -377 -2423 -349
rect -2395 -377 -2357 -349
rect -2329 -377 -2291 -349
rect -2263 -377 -2225 -349
rect -2197 -377 -2159 -349
rect -2131 -377 -2093 -349
rect -2065 -377 -2027 -349
rect -1999 -377 -1961 -349
rect -1933 -377 -1895 -349
rect -1867 -377 -1829 -349
rect -1801 -377 -1763 -349
rect -1735 -377 -1697 -349
rect -1669 -377 -1631 -349
rect -1603 -377 -1565 -349
rect -1537 -377 -1499 -349
rect -1471 -377 -1433 -349
rect -1405 -377 -1367 -349
rect -1339 -377 -1301 -349
rect -1273 -377 -1235 -349
rect -1207 -377 -1169 -349
rect -1141 -377 -1103 -349
rect -1075 -377 -1037 -349
rect -1009 -377 -971 -349
rect -943 -377 -905 -349
rect -877 -377 -839 -349
rect -811 -377 -773 -349
rect -745 -377 -707 -349
rect -679 -377 -641 -349
rect -613 -377 -575 -349
rect -547 -377 -509 -349
rect -481 -377 -443 -349
rect -415 -377 -377 -349
rect -349 -377 -311 -349
rect -283 -377 -245 -349
rect -217 -377 -179 -349
rect -151 -377 -113 -349
rect -85 -377 -47 -349
rect -19 -377 19 -349
rect 47 -377 85 -349
rect 113 -377 151 -349
rect 179 -377 217 -349
rect 245 -377 283 -349
rect 311 -377 349 -349
rect 377 -377 415 -349
rect 443 -377 481 -349
rect 509 -377 547 -349
rect 575 -377 613 -349
rect 641 -377 679 -349
rect 707 -377 745 -349
rect 773 -377 811 -349
rect 839 -377 877 -349
rect 905 -377 943 -349
rect 971 -377 1009 -349
rect 1037 -377 1075 -349
rect 1103 -377 1141 -349
rect 1169 -377 1207 -349
rect 1235 -377 1273 -349
rect 1301 -377 1339 -349
rect 1367 -377 1405 -349
rect 1433 -377 1471 -349
rect 1499 -377 1537 -349
rect 1565 -377 1603 -349
rect 1631 -377 1669 -349
rect 1697 -377 1735 -349
rect 1763 -377 1801 -349
rect 1829 -377 1867 -349
rect 1895 -377 1933 -349
rect 1961 -377 1999 -349
rect 2027 -377 2065 -349
rect 2093 -377 2131 -349
rect 2159 -377 2197 -349
rect 2225 -377 2263 -349
rect 2291 -377 2329 -349
rect 2357 -377 2395 -349
rect 2423 -377 2461 -349
rect 2489 -377 2527 -349
rect 2555 -377 2593 -349
rect 2621 -377 2626 -349
rect -2626 -382 2626 -377
<< end >>
