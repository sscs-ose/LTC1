magic
tech gf180mcuC
magscale 1 10
timestamp 1695206022
<< metal1 >>
rect 6936 5743 19892 6076
rect 13218 5585 19892 5743
rect 13218 5521 19896 5585
rect 13222 5313 19896 5521
rect 19046 5294 19896 5313
rect 13088 4982 13247 4985
rect 13088 4968 13248 4982
rect 13088 4882 13107 4968
rect 13194 4954 13248 4968
rect 13194 4882 13347 4954
rect 16286 4934 16469 4959
rect 13673 4900 13754 4901
rect 13673 4896 13769 4900
rect 13088 4862 13247 4882
rect 13673 4842 13686 4896
rect 13742 4849 13769 4896
rect 13742 4842 13754 4849
rect 13673 4834 13754 4842
rect 16286 4806 16307 4934
rect 16369 4887 16469 4934
rect 16817 4899 16918 4906
rect 16369 4806 16394 4887
rect 16817 4846 16829 4899
rect 16905 4846 16918 4899
rect 16817 4841 16918 4846
rect 16286 4787 16394 4806
rect 6575 4199 6920 4250
rect 6575 2308 6680 4199
rect 6742 3885 6975 3957
rect 6742 2588 6800 3885
rect 13653 3821 13761 3835
rect 13653 3762 13663 3821
rect 13747 3762 13761 3821
rect 13653 3745 13761 3762
rect 16803 3812 16899 3814
rect 16803 3759 16817 3812
rect 16872 3759 16899 3812
rect 16803 3752 16899 3759
rect 6868 3208 10622 3467
rect 12952 3298 19360 3442
rect 8066 3172 8514 3208
rect 13073 3041 13234 3064
rect 13073 3016 13086 3041
rect 12597 2958 13086 3016
rect 13073 2946 13086 2958
rect 13216 2946 13234 3041
rect 13073 2934 13234 2946
rect 6742 2530 7173 2588
rect 12955 2569 13562 2587
rect 12954 2529 13562 2569
rect 6575 2203 6907 2308
rect 10507 2145 12345 2363
rect 12954 1661 13026 2529
rect 19478 2165 19658 5294
rect 19786 4817 19881 4834
rect 19786 4754 19803 4817
rect 19867 4754 19881 4817
rect 19786 4735 19881 4754
rect 15808 2021 19658 2165
rect 15780 1991 19658 2021
rect 19069 1985 19658 1991
rect 12749 1589 13026 1661
rect 19378 1660 19564 1704
rect 19168 1588 19564 1660
rect 19378 1526 19564 1588
rect 6480 504 6601 523
rect 6480 446 6506 504
rect 6577 446 6601 504
rect 6480 415 6601 446
rect 19204 13 19296 1328
rect 6735 -290 19854 13
<< via1 >>
rect 13107 4882 13194 4968
rect 13686 4842 13742 4896
rect 16307 4806 16369 4934
rect 16829 4846 16905 4899
rect 13660 4233 13716 4287
rect 16814 4239 16877 4328
rect 14710 3848 14771 3902
rect 17858 3853 17927 3905
rect 13663 3762 13747 3821
rect 16817 3759 16872 3812
rect 13086 2946 13216 3041
rect 19803 4754 19867 4817
rect 12421 919 12485 1035
rect 13344 918 13408 1034
rect 6506 446 6577 504
<< metal2 >>
rect 13088 4982 13247 4985
rect 13088 4968 13248 4982
rect 13088 4882 13107 4968
rect 13194 4909 13248 4968
rect 16286 4934 16394 4959
rect 13194 4882 13247 4909
rect 13088 4862 13247 4882
rect 13656 4901 13722 4904
rect 13656 4896 13754 4901
rect 13089 3064 13220 4862
rect 13656 4842 13686 4896
rect 13742 4842 13754 4896
rect 16286 4857 16307 4934
rect 13656 4834 13754 4842
rect 13656 4287 13722 4834
rect 15972 4806 16307 4857
rect 16369 4806 16394 4934
rect 15972 4801 16394 4806
rect 16286 4787 16394 4801
rect 16807 4899 16918 4906
rect 16807 4846 16829 4899
rect 16905 4846 16918 4899
rect 16807 4841 16918 4846
rect 13656 4233 13660 4287
rect 13716 4233 13722 4287
rect 13656 3835 13722 4233
rect 16807 4328 16885 4841
rect 19786 4820 19881 4834
rect 19111 4817 19881 4820
rect 19111 4764 19803 4817
rect 19786 4754 19803 4764
rect 19867 4754 19881 4817
rect 19786 4735 19881 4754
rect 16807 4239 16814 4328
rect 16877 4239 16885 4328
rect 14694 3905 14787 3917
rect 14694 3843 14704 3905
rect 14782 3843 14787 3905
rect 13653 3821 13761 3835
rect 14694 3833 14787 3843
rect 13653 3762 13663 3821
rect 13747 3762 13761 3821
rect 16807 3814 16885 4239
rect 17835 3923 17929 3926
rect 17835 3916 17930 3923
rect 17835 3843 17846 3916
rect 17922 3905 17930 3916
rect 17927 3853 17930 3905
rect 17922 3843 17930 3853
rect 17835 3839 17930 3843
rect 17835 3832 17929 3839
rect 13653 3745 13761 3762
rect 16803 3812 16885 3814
rect 16803 3759 16817 3812
rect 16872 3759 16885 3812
rect 16803 3752 16885 3759
rect 13073 3041 13234 3064
rect 13073 2946 13086 3041
rect 13216 2946 13234 3041
rect 13073 2934 13234 2946
rect 12404 1035 13427 1053
rect 12404 919 12421 1035
rect 12485 1034 13427 1035
rect 12485 919 13344 1034
rect 12404 918 13344 919
rect 13408 918 13427 1034
rect 12404 899 13427 918
rect 6480 508 6601 523
rect 6480 440 6503 508
rect 6579 440 6601 508
rect 6480 415 6601 440
<< via2 >>
rect 14704 3902 14782 3905
rect 14704 3848 14710 3902
rect 14710 3848 14771 3902
rect 14771 3848 14782 3902
rect 14704 3843 14782 3848
rect 17846 3905 17922 3916
rect 17846 3853 17858 3905
rect 17858 3853 17922 3905
rect 17846 3843 17922 3853
rect 6503 504 6579 508
rect 6503 446 6506 504
rect 6506 446 6577 504
rect 6577 446 6579 504
rect 6503 440 6579 446
<< metal3 >>
rect 6480 508 6601 523
rect 6480 440 6503 508
rect 6579 497 6601 508
rect 6579 440 9698 497
rect 9701 440 9758 5102
rect 17835 3923 17933 3927
rect 14694 3907 14791 3917
rect 17835 3916 17934 3923
rect 17835 3907 17846 3916
rect 14694 3905 17846 3907
rect 14694 3843 14704 3905
rect 14782 3843 17846 3905
rect 17922 3907 17934 3916
rect 17922 3843 17939 3907
rect 14694 3839 17939 3843
rect 14694 3833 14791 3839
rect 16095 497 16163 3839
rect 17835 3832 17933 3839
rect 9855 440 16177 497
rect 6480 415 6601 440
use CLK_div_3_mag  CLK_div_3_mag_0
timestamp 1695206022
transform 1 0 6869 0 -1 5543
box -34 -1 6461 3249
use CLK_div_3_mag  CLK_div_3_mag_1
timestamp 1695206022
transform -1 0 12896 0 1 3
box -34 -1 6461 3249
use CLK_div_3_mag  CLK_div_3_mag_2
timestamp 1695206022
transform -1 0 19302 0 1 2
box -34 -1 6461 3249
use JK_FF_mag  JK_FF_mag_0
timestamp 1695127730
transform 1 0 16757 0 1 3301
box -390 0 2603 2148
use JK_FF_mag  JK_FF_mag_1
timestamp 1695127730
transform 1 0 13613 0 1 3298
box -390 0 2603 2148
<< labels >>
flabel via1 19821 4789 19821 4789 0 FreeSans 640 0 0 0 Vdiv108
port 0 nsew
flabel metal1 16191 5515 16191 5515 0 FreeSans 640 0 0 0 VDD
port 1 nsew
flabel metal1 12790 -69 12790 -69 0 FreeSans 640 0 0 0 VSS
port 2 nsew
flabel metal1 19462 1610 19462 1610 0 FreeSans 640 0 0 0 CLK
port 3 nsew
flabel via2 6532 469 6532 469 0 FreeSans 640 0 0 0 RST
port 4 nsew
<< end >>
