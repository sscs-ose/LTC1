magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1227 -1019 1227 1019
<< metal1 >>
rect -227 13 227 19
rect -227 -13 -221 13
rect 221 -13 227 13
rect -227 -19 227 -13
<< via1 >>
rect -221 -13 221 13
<< metal2 >>
rect -227 13 227 19
rect -227 -13 -221 13
rect 221 -13 227 13
rect -227 -19 227 -13
<< end >>
