magic
tech gf180mcuC
magscale 1 10
timestamp 1694584912
<< nwell >>
rect 1738 2353 1814 2427
<< metal1 >>
rect 75 2845 190 2846
rect -304 2802 -208 2817
rect 75 2802 2212 2845
rect -304 2735 -289 2802
rect -222 2735 2212 2802
rect -304 2729 -208 2735
rect 75 2730 2212 2735
rect 2280 2437 2361 2451
rect 74 2255 120 2395
rect 593 2391 883 2437
rect 2167 2435 2426 2437
rect 1738 2421 1814 2427
rect 837 2255 883 2391
rect 1299 2401 1380 2410
rect 1299 2345 1314 2401
rect 1370 2345 1380 2401
rect 1738 2365 1749 2421
rect 1805 2365 1814 2421
rect 2167 2391 2293 2435
rect 2280 2379 2293 2391
rect 2349 2391 2426 2435
rect 2349 2379 2361 2391
rect 2280 2369 2361 2379
rect 1738 2353 1814 2365
rect 1299 2333 1380 2345
rect 1599 2264 1681 2302
rect 1599 2208 1615 2264
rect 1671 2208 1681 2264
rect 1599 2197 1681 2208
rect -111 2028 -25 2042
rect 51 2028 2227 2037
rect -111 2027 2227 2028
rect -111 1962 -99 2027
rect -34 1970 2227 2027
rect -34 1962 118 1970
rect -111 1961 118 1962
rect -111 1955 -25 1961
rect -304 1871 -194 1872
rect -304 1851 2187 1871
rect -304 1784 -289 1851
rect -222 1784 2187 1851
rect -304 1756 2187 1784
rect 1893 1669 1971 1681
rect 687 1625 765 1635
rect 687 1571 699 1625
rect 753 1621 765 1625
rect 753 1575 883 1621
rect 1893 1615 1905 1669
rect 1959 1615 1971 1669
rect 1893 1603 1971 1615
rect 1909 1592 1955 1603
rect 753 1571 765 1575
rect 687 1559 765 1571
rect 74 1284 120 1424
rect 593 1213 639 1466
rect 837 1378 883 1575
rect 1560 1573 1643 1588
rect 1560 1519 1574 1573
rect 1628 1519 1643 1573
rect 1560 1504 1643 1519
rect 1325 1449 1371 1466
rect 1303 1437 1387 1449
rect 1303 1383 1321 1437
rect 1375 1383 1387 1437
rect 1303 1377 1387 1383
rect 1578 1424 1624 1504
rect 1578 1378 1694 1424
rect 2167 1420 2244 1466
rect 2198 1410 2244 1420
rect 2198 1364 2343 1410
rect 816 1319 886 1332
rect 816 1263 826 1319
rect 882 1263 886 1319
rect 1263 1284 1696 1330
rect 816 1251 886 1263
rect 593 1204 696 1213
rect 593 1154 630 1204
rect 618 1150 630 1154
rect 684 1150 696 1204
rect 618 1141 696 1150
rect -110 1057 -29 1064
rect 51 1057 2219 1064
rect -110 1056 2219 1057
rect -110 991 -98 1056
rect -33 997 2219 1056
rect -33 991 118 997
rect -110 990 118 991
rect -110 986 -29 990
rect -299 843 2196 883
rect -299 775 -289 843
rect -222 775 2196 843
rect -299 768 2196 775
rect -299 767 -208 768
rect -299 763 -210 767
rect 749 514 824 526
rect 74 309 120 449
rect 593 354 639 491
rect 749 460 758 514
rect 812 460 824 514
rect 1324 472 1370 490
rect 1319 466 1375 472
rect 749 448 824 460
rect 1303 463 1386 466
rect 2129 464 2175 490
rect 762 402 883 448
rect 1303 409 1320 463
rect 1374 409 1386 463
rect 2124 460 2180 464
rect 2112 455 2189 460
rect 1303 396 1386 409
rect 1648 380 1694 448
rect 2112 401 2125 455
rect 2179 401 2189 455
rect 2112 389 2189 401
rect 1586 373 1694 380
rect 593 308 885 354
rect 1586 319 1599 373
rect 1653 319 1694 373
rect 1586 309 1694 319
rect 1586 305 1655 309
rect -111 86 -18 96
rect -111 19 -99 86
rect -32 19 2229 86
rect -111 7 -18 19
<< via1 >>
rect -289 2735 -222 2802
rect 1314 2345 1370 2401
rect 1749 2365 1805 2421
rect 2293 2379 2349 2435
rect 1615 2208 1671 2264
rect -99 1962 -34 2027
rect -289 1784 -222 1851
rect 699 1571 753 1625
rect 1905 1615 1959 1669
rect 1574 1519 1628 1573
rect 1321 1383 1375 1437
rect 826 1263 882 1319
rect 630 1150 684 1204
rect -98 991 -33 1056
rect -289 775 -222 843
rect 758 460 812 514
rect 1320 409 1374 463
rect 2125 401 2179 455
rect 1599 319 1653 373
rect -99 19 -32 86
<< metal2 >>
rect -304 2802 -208 2817
rect -304 2735 -289 2802
rect -222 2735 -208 2802
rect -304 2729 -208 2735
rect -289 1872 -222 2729
rect 1749 2430 2180 2456
rect 1738 2421 2180 2430
rect 1304 2401 1380 2410
rect 697 2345 1314 2401
rect 1370 2345 1380 2401
rect 1738 2365 1749 2421
rect 1805 2400 2180 2421
rect 1805 2365 1819 2400
rect 1738 2349 1819 2365
rect -111 2027 -25 2042
rect -111 1962 -99 2027
rect -34 1962 -25 2027
rect -111 1955 -25 1962
rect -304 1851 -194 1872
rect -304 1784 -289 1851
rect -222 1784 -194 1851
rect -304 1756 -194 1784
rect -289 883 -222 1756
rect -99 1064 -32 1955
rect 697 1659 753 2345
rect 1304 2333 1380 2345
rect 1599 2293 1681 2302
rect 1599 2264 1960 2293
rect 1599 2208 1615 2264
rect 1671 2237 1960 2264
rect 1671 2208 1681 2237
rect 1599 2197 1681 2208
rect 1904 1681 1960 2237
rect 1893 1669 1971 1681
rect 697 1635 754 1659
rect 687 1625 765 1635
rect 687 1571 699 1625
rect 753 1571 765 1625
rect 1893 1615 1905 1669
rect 1959 1615 1971 1669
rect 1893 1603 1971 1615
rect 687 1559 765 1571
rect 1560 1574 1643 1588
rect 1560 1518 1573 1574
rect 1629 1518 1643 1574
rect 1560 1504 1643 1518
rect 1303 1437 1387 1449
rect 1303 1383 1321 1437
rect 1375 1383 1387 1437
rect 1303 1377 1387 1383
rect 1320 1346 1377 1377
rect 816 1319 886 1332
rect 816 1263 826 1319
rect 882 1263 1002 1319
rect 816 1251 886 1263
rect 616 1204 699 1214
rect 616 1191 630 1204
rect 548 1150 630 1191
rect 684 1150 699 1204
rect 548 1140 699 1150
rect 548 1135 660 1140
rect -110 1056 -29 1064
rect -110 991 -98 1056
rect -33 991 -29 1056
rect -110 986 -29 991
rect -299 843 -210 883
rect -299 775 -289 843
rect -222 775 -210 843
rect -299 763 -210 775
rect -99 96 -32 986
rect 548 640 604 1135
rect 548 584 813 640
rect 757 526 813 584
rect 749 514 824 526
rect 749 460 758 514
rect 812 460 824 514
rect 749 448 824 460
rect 946 464 1002 1263
rect 1321 1127 1377 1346
rect 1321 1071 1654 1127
rect 1303 464 1386 466
rect 946 463 1386 464
rect 946 409 1320 463
rect 1374 409 1386 463
rect 946 408 1386 409
rect 1303 396 1386 408
rect 1598 380 1654 1071
rect 2124 460 2180 2400
rect 2280 2435 2361 2451
rect 2280 2379 2293 2435
rect 2349 2379 2361 2435
rect 2280 2369 2361 2379
rect 2293 1583 2349 2369
rect 2284 1574 2360 1583
rect 2284 1518 2293 1574
rect 2349 1518 2360 1574
rect 2284 1506 2360 1518
rect 2112 455 2189 460
rect 2112 401 2125 455
rect 2179 401 2189 455
rect 2112 389 2189 401
rect 1586 373 1655 380
rect 1586 319 1599 373
rect 1653 319 1655 373
rect 1586 305 1655 319
rect -111 86 -18 96
rect -111 19 -99 86
rect -32 19 -18 86
rect -111 7 -18 19
<< via2 >>
rect 1573 1573 1629 1574
rect 1573 1519 1574 1573
rect 1574 1519 1628 1573
rect 1628 1519 1629 1573
rect 1573 1518 1629 1519
rect 2293 1518 2349 1574
<< metal3 >>
rect 1560 1574 1643 1588
rect 2284 1574 2360 1583
rect 1560 1518 1573 1574
rect 1629 1518 2293 1574
rect 2349 1518 2360 1574
rect 1560 1504 1643 1518
rect 2284 1506 2360 1518
use NAND  NAND_0
timestamp 1694584912
transform 1 0 137 0 1 2043
box -86 -97 530 818
use NAND  NAND_1
timestamp 1694584912
transform 1 0 900 0 1 2043
box -86 -97 530 818
use NAND  NAND_2
timestamp 1694584912
transform 1 0 137 0 1 1072
box -86 -97 530 818
use NAND  NAND_3
timestamp 1694584912
transform 1 0 137 0 1 97
box -86 -97 530 818
use NAND  NAND_4
timestamp 1694584912
transform 1 0 1711 0 1 2043
box -86 -97 530 818
use NAND  NAND_5
timestamp 1694584912
transform 1 0 900 0 1 1072
box -86 -97 530 818
use NAND  NAND_6
timestamp 1694584912
transform 1 0 900 0 1 96
box -86 -97 530 818
use NAND  NAND_7
timestamp 1694584912
transform 1 0 1711 0 1 96
box -86 -97 530 818
use NAND  NAND_8
timestamp 1694584912
transform 1 0 1711 0 1 1072
box -86 -97 530 818
<< labels >>
flabel metal1 93 2328 93 2328 0 FreeSans 480 0 0 0 Ri-1
port 0 nsew
flabel metal1 1098 2792 1098 2792 0 FreeSans 480 0 0 0 VDD
port 1 nsew
flabel metal1 1102 2005 1102 2005 0 FreeSans 480 0 0 0 VSS
port 2 nsew
flabel metal1 2322 1385 2322 1385 0 FreeSans 480 0 0 0 Q
port 3 nsew
flabel metal1 2396 2412 2396 2412 0 FreeSans 480 0 0 0 QB
port 4 nsew
flabel metal1 93 1350 93 1350 0 FreeSans 480 0 0 0 Ci
port 5 nsew
flabel metal1 92 377 92 377 0 FreeSans 480 0 0 0 Ri
port 6 nsew
<< end >>
