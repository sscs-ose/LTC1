magic
tech gf180mcuC
magscale 1 10
timestamp 1692057126
<< nwell >>
rect -2264 -1106 2264 1106
<< pmos >>
rect -2090 416 -1990 976
rect -1886 416 -1786 976
rect -1682 416 -1582 976
rect -1478 416 -1378 976
rect -1274 416 -1174 976
rect -1070 416 -970 976
rect -866 416 -766 976
rect -662 416 -562 976
rect -458 416 -358 976
rect -254 416 -154 976
rect -50 416 50 976
rect 154 416 254 976
rect 358 416 458 976
rect 562 416 662 976
rect 766 416 866 976
rect 970 416 1070 976
rect 1174 416 1274 976
rect 1378 416 1478 976
rect 1582 416 1682 976
rect 1786 416 1886 976
rect 1990 416 2090 976
rect -2090 -280 -1990 280
rect -1886 -280 -1786 280
rect -1682 -280 -1582 280
rect -1478 -280 -1378 280
rect -1274 -280 -1174 280
rect -1070 -280 -970 280
rect -866 -280 -766 280
rect -662 -280 -562 280
rect -458 -280 -358 280
rect -254 -280 -154 280
rect -50 -280 50 280
rect 154 -280 254 280
rect 358 -280 458 280
rect 562 -280 662 280
rect 766 -280 866 280
rect 970 -280 1070 280
rect 1174 -280 1274 280
rect 1378 -280 1478 280
rect 1582 -280 1682 280
rect 1786 -280 1886 280
rect 1990 -280 2090 280
rect -2090 -976 -1990 -416
rect -1886 -976 -1786 -416
rect -1682 -976 -1582 -416
rect -1478 -976 -1378 -416
rect -1274 -976 -1174 -416
rect -1070 -976 -970 -416
rect -866 -976 -766 -416
rect -662 -976 -562 -416
rect -458 -976 -358 -416
rect -254 -976 -154 -416
rect -50 -976 50 -416
rect 154 -976 254 -416
rect 358 -976 458 -416
rect 562 -976 662 -416
rect 766 -976 866 -416
rect 970 -976 1070 -416
rect 1174 -976 1274 -416
rect 1378 -976 1478 -416
rect 1582 -976 1682 -416
rect 1786 -976 1886 -416
rect 1990 -976 2090 -416
<< pdiff >>
rect -2178 963 -2090 976
rect -2178 429 -2165 963
rect -2119 429 -2090 963
rect -2178 416 -2090 429
rect -1990 963 -1886 976
rect -1990 429 -1961 963
rect -1915 429 -1886 963
rect -1990 416 -1886 429
rect -1786 963 -1682 976
rect -1786 429 -1757 963
rect -1711 429 -1682 963
rect -1786 416 -1682 429
rect -1582 963 -1478 976
rect -1582 429 -1553 963
rect -1507 429 -1478 963
rect -1582 416 -1478 429
rect -1378 963 -1274 976
rect -1378 429 -1349 963
rect -1303 429 -1274 963
rect -1378 416 -1274 429
rect -1174 963 -1070 976
rect -1174 429 -1145 963
rect -1099 429 -1070 963
rect -1174 416 -1070 429
rect -970 963 -866 976
rect -970 429 -941 963
rect -895 429 -866 963
rect -970 416 -866 429
rect -766 963 -662 976
rect -766 429 -737 963
rect -691 429 -662 963
rect -766 416 -662 429
rect -562 963 -458 976
rect -562 429 -533 963
rect -487 429 -458 963
rect -562 416 -458 429
rect -358 963 -254 976
rect -358 429 -329 963
rect -283 429 -254 963
rect -358 416 -254 429
rect -154 963 -50 976
rect -154 429 -125 963
rect -79 429 -50 963
rect -154 416 -50 429
rect 50 963 154 976
rect 50 429 79 963
rect 125 429 154 963
rect 50 416 154 429
rect 254 963 358 976
rect 254 429 283 963
rect 329 429 358 963
rect 254 416 358 429
rect 458 963 562 976
rect 458 429 487 963
rect 533 429 562 963
rect 458 416 562 429
rect 662 963 766 976
rect 662 429 691 963
rect 737 429 766 963
rect 662 416 766 429
rect 866 963 970 976
rect 866 429 895 963
rect 941 429 970 963
rect 866 416 970 429
rect 1070 963 1174 976
rect 1070 429 1099 963
rect 1145 429 1174 963
rect 1070 416 1174 429
rect 1274 963 1378 976
rect 1274 429 1303 963
rect 1349 429 1378 963
rect 1274 416 1378 429
rect 1478 963 1582 976
rect 1478 429 1507 963
rect 1553 429 1582 963
rect 1478 416 1582 429
rect 1682 963 1786 976
rect 1682 429 1711 963
rect 1757 429 1786 963
rect 1682 416 1786 429
rect 1886 963 1990 976
rect 1886 429 1915 963
rect 1961 429 1990 963
rect 1886 416 1990 429
rect 2090 963 2178 976
rect 2090 429 2119 963
rect 2165 429 2178 963
rect 2090 416 2178 429
rect -2178 267 -2090 280
rect -2178 -267 -2165 267
rect -2119 -267 -2090 267
rect -2178 -280 -2090 -267
rect -1990 267 -1886 280
rect -1990 -267 -1961 267
rect -1915 -267 -1886 267
rect -1990 -280 -1886 -267
rect -1786 267 -1682 280
rect -1786 -267 -1757 267
rect -1711 -267 -1682 267
rect -1786 -280 -1682 -267
rect -1582 267 -1478 280
rect -1582 -267 -1553 267
rect -1507 -267 -1478 267
rect -1582 -280 -1478 -267
rect -1378 267 -1274 280
rect -1378 -267 -1349 267
rect -1303 -267 -1274 267
rect -1378 -280 -1274 -267
rect -1174 267 -1070 280
rect -1174 -267 -1145 267
rect -1099 -267 -1070 267
rect -1174 -280 -1070 -267
rect -970 267 -866 280
rect -970 -267 -941 267
rect -895 -267 -866 267
rect -970 -280 -866 -267
rect -766 267 -662 280
rect -766 -267 -737 267
rect -691 -267 -662 267
rect -766 -280 -662 -267
rect -562 267 -458 280
rect -562 -267 -533 267
rect -487 -267 -458 267
rect -562 -280 -458 -267
rect -358 267 -254 280
rect -358 -267 -329 267
rect -283 -267 -254 267
rect -358 -280 -254 -267
rect -154 267 -50 280
rect -154 -267 -125 267
rect -79 -267 -50 267
rect -154 -280 -50 -267
rect 50 267 154 280
rect 50 -267 79 267
rect 125 -267 154 267
rect 50 -280 154 -267
rect 254 267 358 280
rect 254 -267 283 267
rect 329 -267 358 267
rect 254 -280 358 -267
rect 458 267 562 280
rect 458 -267 487 267
rect 533 -267 562 267
rect 458 -280 562 -267
rect 662 267 766 280
rect 662 -267 691 267
rect 737 -267 766 267
rect 662 -280 766 -267
rect 866 267 970 280
rect 866 -267 895 267
rect 941 -267 970 267
rect 866 -280 970 -267
rect 1070 267 1174 280
rect 1070 -267 1099 267
rect 1145 -267 1174 267
rect 1070 -280 1174 -267
rect 1274 267 1378 280
rect 1274 -267 1303 267
rect 1349 -267 1378 267
rect 1274 -280 1378 -267
rect 1478 267 1582 280
rect 1478 -267 1507 267
rect 1553 -267 1582 267
rect 1478 -280 1582 -267
rect 1682 267 1786 280
rect 1682 -267 1711 267
rect 1757 -267 1786 267
rect 1682 -280 1786 -267
rect 1886 267 1990 280
rect 1886 -267 1915 267
rect 1961 -267 1990 267
rect 1886 -280 1990 -267
rect 2090 267 2178 280
rect 2090 -267 2119 267
rect 2165 -267 2178 267
rect 2090 -280 2178 -267
rect -2178 -429 -2090 -416
rect -2178 -963 -2165 -429
rect -2119 -963 -2090 -429
rect -2178 -976 -2090 -963
rect -1990 -429 -1886 -416
rect -1990 -963 -1961 -429
rect -1915 -963 -1886 -429
rect -1990 -976 -1886 -963
rect -1786 -429 -1682 -416
rect -1786 -963 -1757 -429
rect -1711 -963 -1682 -429
rect -1786 -976 -1682 -963
rect -1582 -429 -1478 -416
rect -1582 -963 -1553 -429
rect -1507 -963 -1478 -429
rect -1582 -976 -1478 -963
rect -1378 -429 -1274 -416
rect -1378 -963 -1349 -429
rect -1303 -963 -1274 -429
rect -1378 -976 -1274 -963
rect -1174 -429 -1070 -416
rect -1174 -963 -1145 -429
rect -1099 -963 -1070 -429
rect -1174 -976 -1070 -963
rect -970 -429 -866 -416
rect -970 -963 -941 -429
rect -895 -963 -866 -429
rect -970 -976 -866 -963
rect -766 -429 -662 -416
rect -766 -963 -737 -429
rect -691 -963 -662 -429
rect -766 -976 -662 -963
rect -562 -429 -458 -416
rect -562 -963 -533 -429
rect -487 -963 -458 -429
rect -562 -976 -458 -963
rect -358 -429 -254 -416
rect -358 -963 -329 -429
rect -283 -963 -254 -429
rect -358 -976 -254 -963
rect -154 -429 -50 -416
rect -154 -963 -125 -429
rect -79 -963 -50 -429
rect -154 -976 -50 -963
rect 50 -429 154 -416
rect 50 -963 79 -429
rect 125 -963 154 -429
rect 50 -976 154 -963
rect 254 -429 358 -416
rect 254 -963 283 -429
rect 329 -963 358 -429
rect 254 -976 358 -963
rect 458 -429 562 -416
rect 458 -963 487 -429
rect 533 -963 562 -429
rect 458 -976 562 -963
rect 662 -429 766 -416
rect 662 -963 691 -429
rect 737 -963 766 -429
rect 662 -976 766 -963
rect 866 -429 970 -416
rect 866 -963 895 -429
rect 941 -963 970 -429
rect 866 -976 970 -963
rect 1070 -429 1174 -416
rect 1070 -963 1099 -429
rect 1145 -963 1174 -429
rect 1070 -976 1174 -963
rect 1274 -429 1378 -416
rect 1274 -963 1303 -429
rect 1349 -963 1378 -429
rect 1274 -976 1378 -963
rect 1478 -429 1582 -416
rect 1478 -963 1507 -429
rect 1553 -963 1582 -429
rect 1478 -976 1582 -963
rect 1682 -429 1786 -416
rect 1682 -963 1711 -429
rect 1757 -963 1786 -429
rect 1682 -976 1786 -963
rect 1886 -429 1990 -416
rect 1886 -963 1915 -429
rect 1961 -963 1990 -429
rect 1886 -976 1990 -963
rect 2090 -429 2178 -416
rect 2090 -963 2119 -429
rect 2165 -963 2178 -429
rect 2090 -976 2178 -963
<< pdiffc >>
rect -2165 429 -2119 963
rect -1961 429 -1915 963
rect -1757 429 -1711 963
rect -1553 429 -1507 963
rect -1349 429 -1303 963
rect -1145 429 -1099 963
rect -941 429 -895 963
rect -737 429 -691 963
rect -533 429 -487 963
rect -329 429 -283 963
rect -125 429 -79 963
rect 79 429 125 963
rect 283 429 329 963
rect 487 429 533 963
rect 691 429 737 963
rect 895 429 941 963
rect 1099 429 1145 963
rect 1303 429 1349 963
rect 1507 429 1553 963
rect 1711 429 1757 963
rect 1915 429 1961 963
rect 2119 429 2165 963
rect -2165 -267 -2119 267
rect -1961 -267 -1915 267
rect -1757 -267 -1711 267
rect -1553 -267 -1507 267
rect -1349 -267 -1303 267
rect -1145 -267 -1099 267
rect -941 -267 -895 267
rect -737 -267 -691 267
rect -533 -267 -487 267
rect -329 -267 -283 267
rect -125 -267 -79 267
rect 79 -267 125 267
rect 283 -267 329 267
rect 487 -267 533 267
rect 691 -267 737 267
rect 895 -267 941 267
rect 1099 -267 1145 267
rect 1303 -267 1349 267
rect 1507 -267 1553 267
rect 1711 -267 1757 267
rect 1915 -267 1961 267
rect 2119 -267 2165 267
rect -2165 -963 -2119 -429
rect -1961 -963 -1915 -429
rect -1757 -963 -1711 -429
rect -1553 -963 -1507 -429
rect -1349 -963 -1303 -429
rect -1145 -963 -1099 -429
rect -941 -963 -895 -429
rect -737 -963 -691 -429
rect -533 -963 -487 -429
rect -329 -963 -283 -429
rect -125 -963 -79 -429
rect 79 -963 125 -429
rect 283 -963 329 -429
rect 487 -963 533 -429
rect 691 -963 737 -429
rect 895 -963 941 -429
rect 1099 -963 1145 -429
rect 1303 -963 1349 -429
rect 1507 -963 1553 -429
rect 1711 -963 1757 -429
rect 1915 -963 1961 -429
rect 2119 -963 2165 -429
<< polysilicon >>
rect -2090 976 -1990 1020
rect -1886 976 -1786 1020
rect -1682 976 -1582 1020
rect -1478 976 -1378 1020
rect -1274 976 -1174 1020
rect -1070 976 -970 1020
rect -866 976 -766 1020
rect -662 976 -562 1020
rect -458 976 -358 1020
rect -254 976 -154 1020
rect -50 976 50 1020
rect 154 976 254 1020
rect 358 976 458 1020
rect 562 976 662 1020
rect 766 976 866 1020
rect 970 976 1070 1020
rect 1174 976 1274 1020
rect 1378 976 1478 1020
rect 1582 976 1682 1020
rect 1786 976 1886 1020
rect 1990 976 2090 1020
rect -2090 372 -1990 416
rect -1886 372 -1786 416
rect -1682 372 -1582 416
rect -1478 372 -1378 416
rect -1274 372 -1174 416
rect -1070 372 -970 416
rect -866 372 -766 416
rect -662 372 -562 416
rect -458 372 -358 416
rect -254 372 -154 416
rect -50 372 50 416
rect 154 372 254 416
rect 358 372 458 416
rect 562 372 662 416
rect 766 372 866 416
rect 970 372 1070 416
rect 1174 372 1274 416
rect 1378 372 1478 416
rect 1582 372 1682 416
rect 1786 372 1886 416
rect 1990 372 2090 416
rect -2090 280 -1990 324
rect -1886 280 -1786 324
rect -1682 280 -1582 324
rect -1478 280 -1378 324
rect -1274 280 -1174 324
rect -1070 280 -970 324
rect -866 280 -766 324
rect -662 280 -562 324
rect -458 280 -358 324
rect -254 280 -154 324
rect -50 280 50 324
rect 154 280 254 324
rect 358 280 458 324
rect 562 280 662 324
rect 766 280 866 324
rect 970 280 1070 324
rect 1174 280 1274 324
rect 1378 280 1478 324
rect 1582 280 1682 324
rect 1786 280 1886 324
rect 1990 280 2090 324
rect -2090 -324 -1990 -280
rect -1886 -324 -1786 -280
rect -1682 -324 -1582 -280
rect -1478 -324 -1378 -280
rect -1274 -324 -1174 -280
rect -1070 -324 -970 -280
rect -866 -324 -766 -280
rect -662 -324 -562 -280
rect -458 -324 -358 -280
rect -254 -324 -154 -280
rect -50 -324 50 -280
rect 154 -324 254 -280
rect 358 -324 458 -280
rect 562 -324 662 -280
rect 766 -324 866 -280
rect 970 -324 1070 -280
rect 1174 -324 1274 -280
rect 1378 -324 1478 -280
rect 1582 -324 1682 -280
rect 1786 -324 1886 -280
rect 1990 -324 2090 -280
rect -2090 -416 -1990 -372
rect -1886 -416 -1786 -372
rect -1682 -416 -1582 -372
rect -1478 -416 -1378 -372
rect -1274 -416 -1174 -372
rect -1070 -416 -970 -372
rect -866 -416 -766 -372
rect -662 -416 -562 -372
rect -458 -416 -358 -372
rect -254 -416 -154 -372
rect -50 -416 50 -372
rect 154 -416 254 -372
rect 358 -416 458 -372
rect 562 -416 662 -372
rect 766 -416 866 -372
rect 970 -416 1070 -372
rect 1174 -416 1274 -372
rect 1378 -416 1478 -372
rect 1582 -416 1682 -372
rect 1786 -416 1886 -372
rect 1990 -416 2090 -372
rect -2090 -1020 -1990 -976
rect -1886 -1020 -1786 -976
rect -1682 -1020 -1582 -976
rect -1478 -1020 -1378 -976
rect -1274 -1020 -1174 -976
rect -1070 -1020 -970 -976
rect -866 -1020 -766 -976
rect -662 -1020 -562 -976
rect -458 -1020 -358 -976
rect -254 -1020 -154 -976
rect -50 -1020 50 -976
rect 154 -1020 254 -976
rect 358 -1020 458 -976
rect 562 -1020 662 -976
rect 766 -1020 866 -976
rect 970 -1020 1070 -976
rect 1174 -1020 1274 -976
rect 1378 -1020 1478 -976
rect 1582 -1020 1682 -976
rect 1786 -1020 1886 -976
rect 1990 -1020 2090 -976
<< metal1 >>
rect -2165 963 -2119 974
rect -2165 418 -2119 429
rect -1961 963 -1915 974
rect -1961 418 -1915 429
rect -1757 963 -1711 974
rect -1757 418 -1711 429
rect -1553 963 -1507 974
rect -1553 418 -1507 429
rect -1349 963 -1303 974
rect -1349 418 -1303 429
rect -1145 963 -1099 974
rect -1145 418 -1099 429
rect -941 963 -895 974
rect -941 418 -895 429
rect -737 963 -691 974
rect -737 418 -691 429
rect -533 963 -487 974
rect -533 418 -487 429
rect -329 963 -283 974
rect -329 418 -283 429
rect -125 963 -79 974
rect -125 418 -79 429
rect 79 963 125 974
rect 79 418 125 429
rect 283 963 329 974
rect 283 418 329 429
rect 487 963 533 974
rect 487 418 533 429
rect 691 963 737 974
rect 691 418 737 429
rect 895 963 941 974
rect 895 418 941 429
rect 1099 963 1145 974
rect 1099 418 1145 429
rect 1303 963 1349 974
rect 1303 418 1349 429
rect 1507 963 1553 974
rect 1507 418 1553 429
rect 1711 963 1757 974
rect 1711 418 1757 429
rect 1915 963 1961 974
rect 1915 418 1961 429
rect 2119 963 2165 974
rect 2119 418 2165 429
rect -2165 267 -2119 278
rect -2165 -278 -2119 -267
rect -1961 267 -1915 278
rect -1961 -278 -1915 -267
rect -1757 267 -1711 278
rect -1757 -278 -1711 -267
rect -1553 267 -1507 278
rect -1553 -278 -1507 -267
rect -1349 267 -1303 278
rect -1349 -278 -1303 -267
rect -1145 267 -1099 278
rect -1145 -278 -1099 -267
rect -941 267 -895 278
rect -941 -278 -895 -267
rect -737 267 -691 278
rect -737 -278 -691 -267
rect -533 267 -487 278
rect -533 -278 -487 -267
rect -329 267 -283 278
rect -329 -278 -283 -267
rect -125 267 -79 278
rect -125 -278 -79 -267
rect 79 267 125 278
rect 79 -278 125 -267
rect 283 267 329 278
rect 283 -278 329 -267
rect 487 267 533 278
rect 487 -278 533 -267
rect 691 267 737 278
rect 691 -278 737 -267
rect 895 267 941 278
rect 895 -278 941 -267
rect 1099 267 1145 278
rect 1099 -278 1145 -267
rect 1303 267 1349 278
rect 1303 -278 1349 -267
rect 1507 267 1553 278
rect 1507 -278 1553 -267
rect 1711 267 1757 278
rect 1711 -278 1757 -267
rect 1915 267 1961 278
rect 1915 -278 1961 -267
rect 2119 267 2165 278
rect 2119 -278 2165 -267
rect -2165 -429 -2119 -418
rect -2165 -974 -2119 -963
rect -1961 -429 -1915 -418
rect -1961 -974 -1915 -963
rect -1757 -429 -1711 -418
rect -1757 -974 -1711 -963
rect -1553 -429 -1507 -418
rect -1553 -974 -1507 -963
rect -1349 -429 -1303 -418
rect -1349 -974 -1303 -963
rect -1145 -429 -1099 -418
rect -1145 -974 -1099 -963
rect -941 -429 -895 -418
rect -941 -974 -895 -963
rect -737 -429 -691 -418
rect -737 -974 -691 -963
rect -533 -429 -487 -418
rect -533 -974 -487 -963
rect -329 -429 -283 -418
rect -329 -974 -283 -963
rect -125 -429 -79 -418
rect -125 -974 -79 -963
rect 79 -429 125 -418
rect 79 -974 125 -963
rect 283 -429 329 -418
rect 283 -974 329 -963
rect 487 -429 533 -418
rect 487 -974 533 -963
rect 691 -429 737 -418
rect 691 -974 737 -963
rect 895 -429 941 -418
rect 895 -974 941 -963
rect 1099 -429 1145 -418
rect 1099 -974 1145 -963
rect 1303 -429 1349 -418
rect 1303 -974 1349 -963
rect 1507 -429 1553 -418
rect 1507 -974 1553 -963
rect 1711 -429 1757 -418
rect 1711 -974 1757 -963
rect 1915 -429 1961 -418
rect 1915 -974 1961 -963
rect 2119 -429 2165 -418
rect 2119 -974 2165 -963
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 2.8 l 0.5 m 3 nf 21 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
