magic
tech gf180mcuC
magscale 1 10
timestamp 1714559211
<< nsubdiff >>
rect 12139 16031 12422 16032
rect 12139 16000 12429 16031
rect 12139 15970 12449 16000
rect 12139 15960 12298 15970
rect 3928 13170 4184 13250
<< metal1 >>
rect 1317 16101 17677 16746
rect 1317 16075 9653 16101
rect 1317 15657 3173 16075
rect 1317 15649 2510 15657
rect 1368 8107 1617 15649
rect 14970 15586 15130 15670
rect 14751 15528 15130 15586
rect 14970 15480 15130 15528
rect 3050 11490 3260 11530
rect 3050 11340 3090 11490
rect 3220 11340 3260 11490
rect 6398 11389 17640 11685
rect 3050 11300 3260 11340
rect 3441 11256 17640 11389
rect 3441 11239 15730 11256
rect 3441 11130 15727 11239
rect 9500 10715 9624 10727
rect 9500 10641 9514 10715
rect 9608 10641 9624 10715
rect 9500 10631 9624 10641
rect 16051 9653 16259 9723
rect 9465 9581 9726 9653
rect 15843 9581 16259 9653
rect 3440 8712 3720 8740
rect 3440 8710 3861 8712
rect 3440 8580 3490 8710
rect 3670 8654 3861 8710
rect 3670 8580 3720 8654
rect 3440 8560 3720 8580
rect 6724 8107 6888 9128
rect 7281 8107 7445 9154
rect 7876 8107 8040 9147
rect 8393 8107 8557 9121
rect 8863 8107 9027 9134
rect 9267 8107 9431 9167
rect 9668 8712 9726 9581
rect 16051 9510 16259 9581
rect 9668 8654 10254 8712
rect 13002 8107 13166 9143
rect 13482 8107 13646 9143
rect 14015 8107 14179 9170
rect 14416 8107 14580 9163
rect 14817 8107 14981 9150
rect 15316 8107 15480 9170
rect 1317 7658 17710 8107
<< via1 >>
rect 3090 11340 3220 11490
rect 9514 10641 9608 10715
rect 3490 8580 3670 8710
<< metal2 >>
rect 3490 11590 4570 11750
rect 3050 11490 3260 11530
rect 3050 11340 3090 11490
rect 3220 11340 3260 11490
rect 3050 11300 3260 11340
rect 3490 8740 3650 11590
rect 9500 10720 9624 10727
rect 9500 10638 9506 10720
rect 9616 10638 9624 10720
rect 9500 10631 9624 10638
rect 3440 8710 3720 8740
rect 3440 8580 3490 8710
rect 3670 8580 3720 8710
rect 3440 8560 3720 8580
<< via2 >>
rect 3090 11340 3220 11490
rect 9506 10715 9616 10720
rect 9506 10641 9514 10715
rect 9514 10641 9608 10715
rect 9608 10641 9616 10715
rect 9506 10638 9616 10641
<< metal3 >>
rect 3050 11490 3260 11530
rect 3050 11340 3090 11490
rect 3220 11455 3260 11490
rect 6212 11455 6293 11705
rect 3220 11374 6293 11455
rect 3220 11340 3260 11374
rect 3050 11300 3260 11340
rect 6212 10750 6293 11374
rect 6461 10966 12885 11009
rect 6460 10909 12885 10966
rect 6461 10739 6518 10909
rect 9512 10746 9612 10909
rect 9486 10720 9641 10746
rect 12828 10745 12885 10909
rect 9486 10638 9506 10720
rect 9616 10638 9641 10720
rect 9486 10616 9641 10638
use CLK_div_3_mag  CLK_div_3_mag_0
timestamp 1714558796
transform -1 0 9601 0 -1 11239
box -40 -1 6461 3249
use CLK_div_3_mag  CLK_div_3_mag_1
timestamp 1714558796
transform -1 0 15970 0 -1 11239
box -40 -1 6461 3249
use CLK_DIV_11_mag_new  CLK_DIV_11_mag_new_0
timestamp 1714559059
transform 1 0 2617 0 -1 16936
box -827 763 15023 5476
<< labels >>
flabel metal1 9843 7982 9843 7982 0 FreeSans 640 0 0 0 VDD
port 0 nsew
flabel metal1 16004 11498 16004 11498 0 FreeSans 640 0 0 0 VSS
port 1 nsew
flabel metal1 16088 9631 16088 9631 0 FreeSans 640 0 0 0 CLK
port 2 nsew
flabel metal1 15033 15585 15033 15585 0 FreeSans 640 0 0 0 Vdiv99
port 3 nsew
flabel via2 3141 11415 3141 11415 0 FreeSans 640 0 0 0 RST
port 4 nsew
<< end >>
