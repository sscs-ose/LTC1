magic
tech gf180mcuC
magscale 1 10
timestamp 1693911244
<< nwell >>
rect -202 -1902 202 1902
<< pmos >>
rect -28 1172 28 1772
rect -28 436 28 1036
rect -28 -300 28 300
rect -28 -1036 28 -436
rect -28 -1772 28 -1172
<< pdiff >>
rect -116 1759 -28 1772
rect -116 1185 -103 1759
rect -57 1185 -28 1759
rect -116 1172 -28 1185
rect 28 1759 116 1772
rect 28 1185 57 1759
rect 103 1185 116 1759
rect 28 1172 116 1185
rect -116 1023 -28 1036
rect -116 449 -103 1023
rect -57 449 -28 1023
rect -116 436 -28 449
rect 28 1023 116 1036
rect 28 449 57 1023
rect 103 449 116 1023
rect 28 436 116 449
rect -116 287 -28 300
rect -116 -287 -103 287
rect -57 -287 -28 287
rect -116 -300 -28 -287
rect 28 287 116 300
rect 28 -287 57 287
rect 103 -287 116 287
rect 28 -300 116 -287
rect -116 -449 -28 -436
rect -116 -1023 -103 -449
rect -57 -1023 -28 -449
rect -116 -1036 -28 -1023
rect 28 -449 116 -436
rect 28 -1023 57 -449
rect 103 -1023 116 -449
rect 28 -1036 116 -1023
rect -116 -1185 -28 -1172
rect -116 -1759 -103 -1185
rect -57 -1759 -28 -1185
rect -116 -1772 -28 -1759
rect 28 -1185 116 -1172
rect 28 -1759 57 -1185
rect 103 -1759 116 -1185
rect 28 -1772 116 -1759
<< pdiffc >>
rect -103 1185 -57 1759
rect 57 1185 103 1759
rect -103 449 -57 1023
rect 57 449 103 1023
rect -103 -287 -57 287
rect 57 -287 103 287
rect -103 -1023 -57 -449
rect 57 -1023 103 -449
rect -103 -1759 -57 -1185
rect 57 -1759 103 -1185
<< polysilicon >>
rect -28 1772 28 1816
rect -28 1128 28 1172
rect -28 1036 28 1080
rect -28 392 28 436
rect -28 300 28 344
rect -28 -344 28 -300
rect -28 -436 28 -392
rect -28 -1080 28 -1036
rect -28 -1172 28 -1128
rect -28 -1816 28 -1772
<< metal1 >>
rect -103 1759 -57 1770
rect -103 1174 -57 1185
rect 57 1759 103 1770
rect 57 1174 103 1185
rect -103 1023 -57 1034
rect -103 438 -57 449
rect 57 1023 103 1034
rect 57 438 103 449
rect -103 287 -57 298
rect -103 -298 -57 -287
rect 57 287 103 298
rect 57 -298 103 -287
rect -103 -449 -57 -438
rect -103 -1034 -57 -1023
rect 57 -449 103 -438
rect 57 -1034 103 -1023
rect -103 -1185 -57 -1174
rect -103 -1770 -57 -1759
rect 57 -1185 103 -1174
rect 57 -1770 103 -1759
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 3 l 0.280 m 5 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
