magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1391 1019 1391
<< metal2 >>
rect -19 386 19 391
rect -19 358 -14 386
rect 14 358 19 386
rect -19 324 19 358
rect -19 296 -14 324
rect 14 296 19 324
rect -19 262 19 296
rect -19 234 -14 262
rect 14 234 19 262
rect -19 200 19 234
rect -19 172 -14 200
rect 14 172 19 200
rect -19 138 19 172
rect -19 110 -14 138
rect 14 110 19 138
rect -19 76 19 110
rect -19 48 -14 76
rect 14 48 19 76
rect -19 14 19 48
rect -19 -14 -14 14
rect 14 -14 19 14
rect -19 -48 19 -14
rect -19 -76 -14 -48
rect 14 -76 19 -48
rect -19 -110 19 -76
rect -19 -138 -14 -110
rect 14 -138 19 -110
rect -19 -172 19 -138
rect -19 -200 -14 -172
rect 14 -200 19 -172
rect -19 -234 19 -200
rect -19 -262 -14 -234
rect 14 -262 19 -234
rect -19 -296 19 -262
rect -19 -324 -14 -296
rect 14 -324 19 -296
rect -19 -358 19 -324
rect -19 -386 -14 -358
rect 14 -386 19 -358
rect -19 -391 19 -386
<< via2 >>
rect -14 358 14 386
rect -14 296 14 324
rect -14 234 14 262
rect -14 172 14 200
rect -14 110 14 138
rect -14 48 14 76
rect -14 -14 14 14
rect -14 -76 14 -48
rect -14 -138 14 -110
rect -14 -200 14 -172
rect -14 -262 14 -234
rect -14 -324 14 -296
rect -14 -386 14 -358
<< metal3 >>
rect -19 386 19 391
rect -19 358 -14 386
rect 14 358 19 386
rect -19 324 19 358
rect -19 296 -14 324
rect 14 296 19 324
rect -19 262 19 296
rect -19 234 -14 262
rect 14 234 19 262
rect -19 200 19 234
rect -19 172 -14 200
rect 14 172 19 200
rect -19 138 19 172
rect -19 110 -14 138
rect 14 110 19 138
rect -19 76 19 110
rect -19 48 -14 76
rect 14 48 19 76
rect -19 14 19 48
rect -19 -14 -14 14
rect 14 -14 19 14
rect -19 -48 19 -14
rect -19 -76 -14 -48
rect 14 -76 19 -48
rect -19 -110 19 -76
rect -19 -138 -14 -110
rect 14 -138 19 -110
rect -19 -172 19 -138
rect -19 -200 -14 -172
rect 14 -200 19 -172
rect -19 -234 19 -200
rect -19 -262 -14 -234
rect 14 -262 19 -234
rect -19 -296 19 -262
rect -19 -324 -14 -296
rect 14 -324 19 -296
rect -19 -358 19 -324
rect -19 -386 -14 -358
rect 14 -386 19 -358
rect -19 -391 19 -386
<< end >>
