magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2495 -2795 2495 2795
<< psubdiff >>
rect -495 773 495 795
rect -495 -773 -473 773
rect 473 -773 495 773
rect -495 -795 495 -773
<< psubdiffcont >>
rect -473 -773 473 773
<< metal1 >>
rect -484 773 484 784
rect -484 -773 -473 773
rect 473 -773 484 773
rect -484 -784 484 -773
<< end >>
