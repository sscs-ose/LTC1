magic
tech gf180mcuC
magscale 1 10
timestamp 1695096662
<< nwell >>
rect -424 -786 424 786
<< nsubdiff >>
rect -400 690 400 762
rect -400 -690 -328 690
rect 328 -690 400 690
rect -400 -762 400 -690
<< polysilicon >>
rect -240 589 -40 602
rect -240 543 -227 589
rect -53 543 -40 589
rect -240 500 -40 543
rect -240 -543 -40 -500
rect -240 -589 -227 -543
rect -53 -589 -40 -543
rect -240 -602 -40 -589
rect 40 589 240 602
rect 40 543 53 589
rect 227 543 240 589
rect 40 500 240 543
rect 40 -543 240 -500
rect 40 -589 53 -543
rect 227 -589 240 -543
rect 40 -602 240 -589
<< polycontact >>
rect -227 543 -53 589
rect -227 -589 -53 -543
rect 53 543 227 589
rect 53 -589 227 -543
<< ppolyres >>
rect -240 -500 -40 500
rect 40 -500 240 500
<< metal1 >>
rect -238 543 -227 589
rect -53 543 -42 589
rect 42 543 53 589
rect 227 543 238 589
rect -238 -589 -227 -543
rect -53 -589 -42 -543
rect 42 -589 53 -543
rect 227 -589 238 -543
<< properties >>
string FIXED_BBOX -364 -726 364 726
string gencell ppolyf_u
string library gf180mcu
string parameters w 1.0 l 5.0 m 1 nx 2 wmin 0.80 lmin 1.00 rho 315 val 1.693k dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 0 grc 0 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 0
<< end >>
