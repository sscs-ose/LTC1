** sch_path: /home/shahid/GF180Projects/inv/Xschem/untitled.sch
**.subckt untitled
x1 VSS IN OUT VDD inv_my
C1 OUT VSS 50f m=1
V1 IN VSS pulse (0 3.3 0 100p 100p 100n 200n)
.save i(v1)
V2 VSS GND 0
.save i(v2)
V3 VDD VSS 3.3
.save i(v3)
**** begin user architecture code

.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical



.control
save all
dc v1 0 3.3 0.1
plot v(IN) v(OUT)

tran 10p 1u
plot v(IN) v(OUT)
plot ()
*write test_nfet_03v3.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  inv_my.sym # of pins=4
** sym_path: /home/shahid/GF180Projects/inv/Xschem/inv_my.sym
** sch_path: /home/shahid/GF180Projects/inv/Xschem/inv_my.sch
.subckt inv_my VSS IN OUT VDD
*.iopin VDD
*.iopin VSS
*.ipin IN
*.opin OUT
XM1 OUT IN VSS VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 OUT IN VDD VDD pfet_03v3 L=0.28u W=0.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends

.GLOBAL GND
.end
