magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -989 -1022 2639 1022
<< metal4 >>
rect 14 14 1636 19
rect 14 -14 19 14
rect 47 -14 85 14
rect 113 -14 151 14
rect 179 -14 217 14
rect 245 -14 283 14
rect 311 -14 349 14
rect 377 -14 415 14
rect 443 -14 481 14
rect 509 -14 547 14
rect 575 -14 613 14
rect 641 -14 679 14
rect 707 -14 745 14
rect 773 -14 811 14
rect 839 -14 877 14
rect 905 -14 943 14
rect 971 -14 1009 14
rect 1037 -14 1075 14
rect 1103 -14 1141 14
rect 1169 -14 1207 14
rect 1235 -14 1273 14
rect 1301 -14 1339 14
rect 1367 -14 1405 14
rect 1433 -14 1471 14
rect 1499 -14 1537 14
rect 1565 -14 1603 14
rect 1631 -14 1636 14
rect 14 -19 1636 -14
<< via4 >>
rect 19 -14 47 14
rect 85 -14 113 14
rect 151 -14 179 14
rect 217 -14 245 14
rect 283 -14 311 14
rect 349 -14 377 14
rect 415 -14 443 14
rect 481 -14 509 14
rect 547 -14 575 14
rect 613 -14 641 14
rect 679 -14 707 14
rect 745 -14 773 14
rect 811 -14 839 14
rect 877 -14 905 14
rect 943 -14 971 14
rect 1009 -14 1037 14
rect 1075 -14 1103 14
rect 1141 -14 1169 14
rect 1207 -14 1235 14
rect 1273 -14 1301 14
rect 1339 -14 1367 14
rect 1405 -14 1433 14
rect 1471 -14 1499 14
rect 1537 -14 1565 14
rect 1603 -14 1631 14
<< metal5 >>
rect 11 14 1639 22
rect 11 -14 19 14
rect 47 -14 85 14
rect 113 -14 151 14
rect 179 -14 217 14
rect 245 -14 283 14
rect 311 -14 349 14
rect 377 -14 415 14
rect 443 -14 481 14
rect 509 -14 547 14
rect 575 -14 613 14
rect 641 -14 679 14
rect 707 -14 745 14
rect 773 -14 811 14
rect 839 -14 877 14
rect 905 -14 943 14
rect 971 -14 1009 14
rect 1037 -14 1075 14
rect 1103 -14 1141 14
rect 1169 -14 1207 14
rect 1235 -14 1273 14
rect 1301 -14 1339 14
rect 1367 -14 1405 14
rect 1433 -14 1471 14
rect 1499 -14 1537 14
rect 1565 -14 1603 14
rect 1631 -14 1639 14
rect 11 -22 1639 -14
<< end >>
