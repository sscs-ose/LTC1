** sch_path: /home/shahid/GF180Projects/PGA_Decoder/Resis_cap/xschem/resis_PGA.sch
**.subckt resis_PGA VDD A B C D E F G H
*.iopin VDD
*.iopin A
*.iopin B
*.iopin C
*.iopin D
*.iopin E
*.iopin F
*.iopin G
*.iopin H
XR1 A net1 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR2 net1 net2 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR3 net2 net3 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR4 net3 net4 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR5 net4 net5 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR6 net5 net6 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR7 net6 net7 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR8 net7 net8 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR9 net8 net9 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR10 net9 B VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR11 C net10 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR12 net10 net11 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR13 net11 net12 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR14 net12 net13 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR15 net13 net14 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR16 net14 net15 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR17 net15 net16 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR18 net16 B VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR19 C net17 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR20 net17 net18 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR21 net18 net19 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR22 net19 net20 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR23 net20 net21 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR24 net21 net22 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR25 net22 net23 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR26 net23 net24 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR27 net24 net25 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR28 net25 net26 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR29 net26 net27 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR30 net27 D VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR31 E net28 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR32 net28 net29 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR33 net29 net30 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR34 net30 net31 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR35 net31 net32 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR36 net32 net33 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR37 net33 net34 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR38 net34 net35 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR39 net35 net36 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR40 net36 net37 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR41 net37 net38 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR42 net38 net39 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR43 net39 net40 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR44 net40 net41 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR45 net41 D VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR46 E net42 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR47 net42 net43 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR48 net43 net44 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR49 net44 net45 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR50 net45 net46 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR51 net46 net47 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR52 net47 net48 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR53 net48 net49 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR54 net49 net50 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR55 net50 net51 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR56 net51 net52 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR57 net52 net53 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR58 net53 net54 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR59 net54 net55 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR60 net55 F VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR61 G net56 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR62 net56 net57 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR63 net57 net58 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR64 net58 net59 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR65 net59 net60 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR66 net60 net61 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR67 net61 net62 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR68 net62 net63 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR69 net63 net64 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR70 net64 net65 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR71 net65 net66 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR72 net66 F VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR73 G net67 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR74 net67 net68 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR75 net68 net69 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR76 net69 net70 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR77 net70 net71 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR78 net71 net72 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR79 net72 net73 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR80 net73 net74 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR81 net74 net75 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR82 net75 net76 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR83 net76 net77 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR84 net77 net78 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR85 net78 net79 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR86 net79 net80 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR87 net80 net81 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR88 net81 net82 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR89 net82 net83 VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR90 net83 H VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR91 VDD VDD VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR92 VDD VDD VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR93 VDD VDD VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR94 VDD VDD VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR95 VDD VDD VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR96 VDD VDD VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR97 VDD VDD VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR98 VDD VDD VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR99 B B VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR103 H H VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR105 A A VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR100 G G VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR101 E E VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
XR102 E E VDD ppolyf_u r_width=1.2e-6 r_length=1e-6 m=1
**.ends
.end
