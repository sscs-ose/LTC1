magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1097 -1071 1097 1071
<< metal1 >>
rect -97 65 97 71
rect -97 -65 -91 65
rect 91 -65 97 65
rect -97 -71 97 -65
<< via1 >>
rect -91 -65 91 65
<< metal2 >>
rect -97 65 97 71
rect -97 -65 -91 65
rect 91 -65 97 65
rect -97 -71 97 -65
<< end >>
