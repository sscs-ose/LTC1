** sch_path: /home/shahid/Downloads/PLL_pakistan2/top/xschem/pex_Feedback_Divider_mag_TB.sch
**.subckt pex_Feedback_Divider_mag_TB
V1 VDD VSS 3.3
.save i(v1)
V2 VSS GND 0
.save i(v2)
V3 CLK VSS pulse(3.3 0 0 100p 100p 2.50n 5n)
.save i(v3)
C5 Vdiv VSS 1p m=1
V5 RST VSS PWL( 0 0 10n 0 10.001n 3)
.save i(v5)
V4 F0 VSS pulse(3.3 0 0 100p 100p 1u 2u)
.save i(v4)
V6 F1 VSS pulse(3.3 0 0 100p 100p 2u 4u)
.save i(v6)
V7 F2 VSS pulse(3.3 0 0 100p 100p 4u 8u)
.save i(v7)
x1 VSS VDD RST Vdiv F2 F1 F0 CLK pex_Feedback_Divider_mag
**** begin user architecture code

.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical



.include pex_Feedback_Divider_mag.spice
.control
ave F2  F1  F0  CLK  Vdiv  Output2  RST_DIV  x1.net1  x1.net2  x1.PU

tran 1n 10u
plot v(CLK) v(Vdiv)+3.5 v(RST)+7 v(F0)+10.5 v(F1)+14 v(F2)+17.5
write pex_Feedback_Divider_mag_TB.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
