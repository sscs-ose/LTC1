magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2045 -3267 2045 3267
<< psubdiff >>
rect -45 1245 45 1267
rect -45 -1245 -23 1245
rect 23 -1245 45 1245
rect -45 -1267 45 -1245
<< psubdiffcont >>
rect -23 -1245 23 1245
<< metal1 >>
rect -34 1245 34 1256
rect -34 -1245 -23 1245
rect 23 -1245 34 1245
rect -34 -1256 34 -1245
<< end >>
