magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1073 -1073 1073 1073
<< metal1 >>
rect -73 67 73 73
rect -73 41 -67 67
rect -41 41 -13 67
rect 13 41 41 67
rect 67 41 73 67
rect -73 13 73 41
rect -73 -13 -67 13
rect -41 -13 -13 13
rect 13 -13 41 13
rect 67 -13 73 13
rect -73 -41 73 -13
rect -73 -67 -67 -41
rect -41 -67 -13 -41
rect 13 -67 41 -41
rect 67 -67 73 -41
rect -73 -73 73 -67
<< via1 >>
rect -67 41 -41 67
rect -13 41 13 67
rect 41 41 67 67
rect -67 -13 -41 13
rect -13 -13 13 13
rect 41 -13 67 13
rect -67 -67 -41 -41
rect -13 -67 13 -41
rect 41 -67 67 -41
<< metal2 >>
rect -73 67 73 73
rect -73 41 -67 67
rect -41 41 -13 67
rect 13 41 41 67
rect 67 41 73 67
rect -73 13 73 41
rect -73 -13 -67 13
rect -41 -13 -13 13
rect 13 -13 41 13
rect 67 -13 73 13
rect -73 -41 73 -13
rect -73 -67 -67 -41
rect -41 -67 -13 -41
rect 13 -67 41 -41
rect 67 -67 73 -41
rect -73 -73 73 -67
<< end >>
