magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1279 1019 1279
<< metal1 >>
rect -19 273 19 279
rect -19 -273 -13 273
rect 13 -273 19 273
rect -19 -279 19 -273
<< via1 >>
rect -13 -273 13 273
<< metal2 >>
rect -19 273 19 279
rect -19 -273 -13 273
rect 13 -273 19 273
rect -19 -279 19 -273
<< end >>
