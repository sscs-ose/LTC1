magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -2224 -2214 2224 2214
<< nwell >>
rect -224 -214 224 214
<< pmos >>
rect -50 -84 50 84
<< pdiff >>
rect -138 70 -50 84
rect -138 -70 -125 70
rect -79 -70 -50 70
rect -138 -84 -50 -70
rect 50 70 138 84
rect 50 -70 79 70
rect 125 -70 138 70
rect 50 -84 138 -70
<< pdiffc >>
rect -125 -70 -79 70
rect 79 -70 125 70
<< polysilicon >>
rect -50 84 50 128
rect -50 -128 50 -84
<< metal1 >>
rect -125 70 -79 82
rect -125 -82 -79 -70
rect 79 70 125 82
rect 79 -82 125 -70
<< end >>
