magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1071 -1253 1071 1253
<< metal1 >>
rect -71 247 71 253
rect -71 -247 -65 247
rect 65 -247 71 247
rect -71 -253 71 -247
<< via1 >>
rect -65 -247 65 247
<< metal2 >>
rect -71 247 71 253
rect -71 -247 -65 247
rect 65 -247 71 247
rect -71 -253 71 -247
<< end >>
