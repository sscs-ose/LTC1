* NGSPICE file created from and_3_flat.ext - technology: gf180mcuC

.subckt and_3_PEX IN1 VSS VDD OUT IN3 IN2
X0 a_398_212# IN2.t0 a_238_212# VSS.t0 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1 OUT nand3_mag_0.OUT VSS.t4 VSS.t3 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2 nand3_mag_0.OUT IN1.t0 VDD.t1 VDD.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3 nand3_mag_0.OUT IN1.t1 a_398_212# VSS.t5 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X4 nand3_mag_0.OUT IN3.t0 VDD.t2 VDD.t0 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X5 a_238_212# IN3.t1 VSS.t2 VSS.t1 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X6 OUT nand3_mag_0.OUT VDD.t6 VDD.t5 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X7 VDD IN2.t1 nand3_mag_0.OUT VDD.t0 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
R0 IN2.n0 IN2.t0 36.935
R1 IN2.n0 IN2.t1 18.1962
R2 IN2.n1 IN2.n0 4.0005
R3 IN2 IN2.n1 0.087696
R4 IN2.n1 IN2 0.00205172
R5 VSS.t5 VSS.n1 1255.26
R6 VSS.n1 VSS.t3 1037.75
R7 VSS.t0 VSS.t5 994.264
R8 VSS.n2 VSS.t0 596.558
R9 VSS.n2 VSS.t1 397.707
R10 VSS.n1 VSS 391.339
R11 VSS.n0 VSS.t4 9.34566
R12 VSS VSS.t2 6.02545
R13 VSS.n3 VSS.n2 5.2005
R14 VSS.n3 VSS.n0 0.533184
R15 VSS VSS.n0 0.0647857
R16 VSS VSS.n3 0.00380275
R17 OUT OUT.n1 9.36021
R18 OUT OUT.n0 5.13104
R19 IN1.n0 IN1.t1 36.935
R20 IN1.n0 IN1.t0 18.1962
R21 IN1.n1 IN1.n0 4.0005
R22 IN1 IN1.n1 0.0936579
R23 IN1.n1 IN1 0.00365789
R24 VDD.n6 VDD.n5 182.94
R25 VDD.n5 VDD.t5 19.5347
R26 VDD.n7 VDD.n6 6.3005
R27 VDD VDD.t2 5.21184
R28 VDD.n3 VDD.t6 5.14703
R29 VDD.n4 VDD.n1 2.85787
R30 VDD.n1 VDD.t1 2.2755
R31 VDD.n1 VDD.n0 2.2755
R32 VDD.n4 VDD.n3 0.230303
R33 VDD VDD.n4 0.106177
R34 VDD.n3 VDD.n2 0.0460556
R35 VDD.n5 VDD.t0 0.00414464
R36 VDD VDD.n7 0.00166129
R37 VDD.n7 VDD 0.00166129
R38 VDD.n2 VDD 0.00105556
R39 IN3.n0 IN3.t0 30.9379
R40 IN3.n0 IN3.t1 24.5101
R41 IN3 IN3.n0 4.0005
C0 IN1 IN2 0.115f
C1 IN1 nand3_mag_0.OUT 0.257f
C2 a_398_212# IN1 8.64e-19
C3 IN3 VDD 0.158f
C4 OUT IN1 1.89e-19
C5 IN3 IN2 0.0466f
C6 IN3 nand3_mag_0.OUT 0.0908f
C7 IN3 a_238_212# 8.64e-19
C8 VDD IN2 0.171f
C9 VDD nand3_mag_0.OUT 0.663f
C10 VDD a_238_212# 2.21e-19
C11 IN2 nand3_mag_0.OUT 0.21f
C12 a_238_212# IN2 8.64e-19
C13 a_238_212# nand3_mag_0.OUT 0.0202f
C14 a_398_212# IN2 0.00103f
C15 a_398_212# nand3_mag_0.OUT 0.0732f
C16 a_398_212# a_238_212# 0.0504f
C17 VDD OUT 0.121f
C18 OUT nand3_mag_0.OUT 0.135f
C19 IN3 IN1 1.3e-19
C20 VDD IN1 0.149f
C21 a_398_212# VSS 0.0343f
C22 a_238_212# VSS 0.0881f
C23 OUT VSS 0.148f
C24 nand3_mag_0.OUT VSS 0.543f
C25 IN1 VSS 0.213f
C26 IN2 VSS 0.192f
C27 IN3 VSS 0.31f
C28 VDD VSS 2.12f
.ends

