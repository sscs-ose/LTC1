magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -3788 -1090 3788 1090
<< metal2 >>
rect -2788 85 2788 90
rect -2788 57 -2783 85
rect -2755 57 -2712 85
rect -2684 57 -2641 85
rect -2613 57 -2570 85
rect -2542 57 -2499 85
rect -2471 57 -2428 85
rect -2400 57 -2357 85
rect -2329 57 -2286 85
rect -2258 57 -2215 85
rect -2187 57 -2144 85
rect -2116 57 -2073 85
rect -2045 57 -2002 85
rect -1974 57 -1931 85
rect -1903 57 -1860 85
rect -1832 57 -1789 85
rect -1761 57 -1718 85
rect -1690 57 -1647 85
rect -1619 57 -1576 85
rect -1548 57 -1505 85
rect -1477 57 -1434 85
rect -1406 57 -1363 85
rect -1335 57 -1292 85
rect -1264 57 -1221 85
rect -1193 57 -1150 85
rect -1122 57 -1079 85
rect -1051 57 -1008 85
rect -980 57 -937 85
rect -909 57 -866 85
rect -838 57 -795 85
rect -767 57 -724 85
rect -696 57 -653 85
rect -625 57 -582 85
rect -554 57 -511 85
rect -483 57 -440 85
rect -412 57 -369 85
rect -341 57 -298 85
rect -270 57 -227 85
rect -199 57 -156 85
rect -128 57 -85 85
rect -57 57 -14 85
rect 14 57 57 85
rect 85 57 128 85
rect 156 57 199 85
rect 227 57 270 85
rect 298 57 341 85
rect 369 57 412 85
rect 440 57 483 85
rect 511 57 554 85
rect 582 57 625 85
rect 653 57 696 85
rect 724 57 767 85
rect 795 57 838 85
rect 866 57 909 85
rect 937 57 980 85
rect 1008 57 1051 85
rect 1079 57 1122 85
rect 1150 57 1193 85
rect 1221 57 1264 85
rect 1292 57 1335 85
rect 1363 57 1406 85
rect 1434 57 1477 85
rect 1505 57 1548 85
rect 1576 57 1619 85
rect 1647 57 1690 85
rect 1718 57 1761 85
rect 1789 57 1832 85
rect 1860 57 1903 85
rect 1931 57 1974 85
rect 2002 57 2045 85
rect 2073 57 2116 85
rect 2144 57 2187 85
rect 2215 57 2258 85
rect 2286 57 2329 85
rect 2357 57 2400 85
rect 2428 57 2471 85
rect 2499 57 2542 85
rect 2570 57 2613 85
rect 2641 57 2684 85
rect 2712 57 2755 85
rect 2783 57 2788 85
rect -2788 14 2788 57
rect -2788 -14 -2783 14
rect -2755 -14 -2712 14
rect -2684 -14 -2641 14
rect -2613 -14 -2570 14
rect -2542 -14 -2499 14
rect -2471 -14 -2428 14
rect -2400 -14 -2357 14
rect -2329 -14 -2286 14
rect -2258 -14 -2215 14
rect -2187 -14 -2144 14
rect -2116 -14 -2073 14
rect -2045 -14 -2002 14
rect -1974 -14 -1931 14
rect -1903 -14 -1860 14
rect -1832 -14 -1789 14
rect -1761 -14 -1718 14
rect -1690 -14 -1647 14
rect -1619 -14 -1576 14
rect -1548 -14 -1505 14
rect -1477 -14 -1434 14
rect -1406 -14 -1363 14
rect -1335 -14 -1292 14
rect -1264 -14 -1221 14
rect -1193 -14 -1150 14
rect -1122 -14 -1079 14
rect -1051 -14 -1008 14
rect -980 -14 -937 14
rect -909 -14 -866 14
rect -838 -14 -795 14
rect -767 -14 -724 14
rect -696 -14 -653 14
rect -625 -14 -582 14
rect -554 -14 -511 14
rect -483 -14 -440 14
rect -412 -14 -369 14
rect -341 -14 -298 14
rect -270 -14 -227 14
rect -199 -14 -156 14
rect -128 -14 -85 14
rect -57 -14 -14 14
rect 14 -14 57 14
rect 85 -14 128 14
rect 156 -14 199 14
rect 227 -14 270 14
rect 298 -14 341 14
rect 369 -14 412 14
rect 440 -14 483 14
rect 511 -14 554 14
rect 582 -14 625 14
rect 653 -14 696 14
rect 724 -14 767 14
rect 795 -14 838 14
rect 866 -14 909 14
rect 937 -14 980 14
rect 1008 -14 1051 14
rect 1079 -14 1122 14
rect 1150 -14 1193 14
rect 1221 -14 1264 14
rect 1292 -14 1335 14
rect 1363 -14 1406 14
rect 1434 -14 1477 14
rect 1505 -14 1548 14
rect 1576 -14 1619 14
rect 1647 -14 1690 14
rect 1718 -14 1761 14
rect 1789 -14 1832 14
rect 1860 -14 1903 14
rect 1931 -14 1974 14
rect 2002 -14 2045 14
rect 2073 -14 2116 14
rect 2144 -14 2187 14
rect 2215 -14 2258 14
rect 2286 -14 2329 14
rect 2357 -14 2400 14
rect 2428 -14 2471 14
rect 2499 -14 2542 14
rect 2570 -14 2613 14
rect 2641 -14 2684 14
rect 2712 -14 2755 14
rect 2783 -14 2788 14
rect -2788 -57 2788 -14
rect -2788 -85 -2783 -57
rect -2755 -85 -2712 -57
rect -2684 -85 -2641 -57
rect -2613 -85 -2570 -57
rect -2542 -85 -2499 -57
rect -2471 -85 -2428 -57
rect -2400 -85 -2357 -57
rect -2329 -85 -2286 -57
rect -2258 -85 -2215 -57
rect -2187 -85 -2144 -57
rect -2116 -85 -2073 -57
rect -2045 -85 -2002 -57
rect -1974 -85 -1931 -57
rect -1903 -85 -1860 -57
rect -1832 -85 -1789 -57
rect -1761 -85 -1718 -57
rect -1690 -85 -1647 -57
rect -1619 -85 -1576 -57
rect -1548 -85 -1505 -57
rect -1477 -85 -1434 -57
rect -1406 -85 -1363 -57
rect -1335 -85 -1292 -57
rect -1264 -85 -1221 -57
rect -1193 -85 -1150 -57
rect -1122 -85 -1079 -57
rect -1051 -85 -1008 -57
rect -980 -85 -937 -57
rect -909 -85 -866 -57
rect -838 -85 -795 -57
rect -767 -85 -724 -57
rect -696 -85 -653 -57
rect -625 -85 -582 -57
rect -554 -85 -511 -57
rect -483 -85 -440 -57
rect -412 -85 -369 -57
rect -341 -85 -298 -57
rect -270 -85 -227 -57
rect -199 -85 -156 -57
rect -128 -85 -85 -57
rect -57 -85 -14 -57
rect 14 -85 57 -57
rect 85 -85 128 -57
rect 156 -85 199 -57
rect 227 -85 270 -57
rect 298 -85 341 -57
rect 369 -85 412 -57
rect 440 -85 483 -57
rect 511 -85 554 -57
rect 582 -85 625 -57
rect 653 -85 696 -57
rect 724 -85 767 -57
rect 795 -85 838 -57
rect 866 -85 909 -57
rect 937 -85 980 -57
rect 1008 -85 1051 -57
rect 1079 -85 1122 -57
rect 1150 -85 1193 -57
rect 1221 -85 1264 -57
rect 1292 -85 1335 -57
rect 1363 -85 1406 -57
rect 1434 -85 1477 -57
rect 1505 -85 1548 -57
rect 1576 -85 1619 -57
rect 1647 -85 1690 -57
rect 1718 -85 1761 -57
rect 1789 -85 1832 -57
rect 1860 -85 1903 -57
rect 1931 -85 1974 -57
rect 2002 -85 2045 -57
rect 2073 -85 2116 -57
rect 2144 -85 2187 -57
rect 2215 -85 2258 -57
rect 2286 -85 2329 -57
rect 2357 -85 2400 -57
rect 2428 -85 2471 -57
rect 2499 -85 2542 -57
rect 2570 -85 2613 -57
rect 2641 -85 2684 -57
rect 2712 -85 2755 -57
rect 2783 -85 2788 -57
rect -2788 -90 2788 -85
<< via2 >>
rect -2783 57 -2755 85
rect -2712 57 -2684 85
rect -2641 57 -2613 85
rect -2570 57 -2542 85
rect -2499 57 -2471 85
rect -2428 57 -2400 85
rect -2357 57 -2329 85
rect -2286 57 -2258 85
rect -2215 57 -2187 85
rect -2144 57 -2116 85
rect -2073 57 -2045 85
rect -2002 57 -1974 85
rect -1931 57 -1903 85
rect -1860 57 -1832 85
rect -1789 57 -1761 85
rect -1718 57 -1690 85
rect -1647 57 -1619 85
rect -1576 57 -1548 85
rect -1505 57 -1477 85
rect -1434 57 -1406 85
rect -1363 57 -1335 85
rect -1292 57 -1264 85
rect -1221 57 -1193 85
rect -1150 57 -1122 85
rect -1079 57 -1051 85
rect -1008 57 -980 85
rect -937 57 -909 85
rect -866 57 -838 85
rect -795 57 -767 85
rect -724 57 -696 85
rect -653 57 -625 85
rect -582 57 -554 85
rect -511 57 -483 85
rect -440 57 -412 85
rect -369 57 -341 85
rect -298 57 -270 85
rect -227 57 -199 85
rect -156 57 -128 85
rect -85 57 -57 85
rect -14 57 14 85
rect 57 57 85 85
rect 128 57 156 85
rect 199 57 227 85
rect 270 57 298 85
rect 341 57 369 85
rect 412 57 440 85
rect 483 57 511 85
rect 554 57 582 85
rect 625 57 653 85
rect 696 57 724 85
rect 767 57 795 85
rect 838 57 866 85
rect 909 57 937 85
rect 980 57 1008 85
rect 1051 57 1079 85
rect 1122 57 1150 85
rect 1193 57 1221 85
rect 1264 57 1292 85
rect 1335 57 1363 85
rect 1406 57 1434 85
rect 1477 57 1505 85
rect 1548 57 1576 85
rect 1619 57 1647 85
rect 1690 57 1718 85
rect 1761 57 1789 85
rect 1832 57 1860 85
rect 1903 57 1931 85
rect 1974 57 2002 85
rect 2045 57 2073 85
rect 2116 57 2144 85
rect 2187 57 2215 85
rect 2258 57 2286 85
rect 2329 57 2357 85
rect 2400 57 2428 85
rect 2471 57 2499 85
rect 2542 57 2570 85
rect 2613 57 2641 85
rect 2684 57 2712 85
rect 2755 57 2783 85
rect -2783 -14 -2755 14
rect -2712 -14 -2684 14
rect -2641 -14 -2613 14
rect -2570 -14 -2542 14
rect -2499 -14 -2471 14
rect -2428 -14 -2400 14
rect -2357 -14 -2329 14
rect -2286 -14 -2258 14
rect -2215 -14 -2187 14
rect -2144 -14 -2116 14
rect -2073 -14 -2045 14
rect -2002 -14 -1974 14
rect -1931 -14 -1903 14
rect -1860 -14 -1832 14
rect -1789 -14 -1761 14
rect -1718 -14 -1690 14
rect -1647 -14 -1619 14
rect -1576 -14 -1548 14
rect -1505 -14 -1477 14
rect -1434 -14 -1406 14
rect -1363 -14 -1335 14
rect -1292 -14 -1264 14
rect -1221 -14 -1193 14
rect -1150 -14 -1122 14
rect -1079 -14 -1051 14
rect -1008 -14 -980 14
rect -937 -14 -909 14
rect -866 -14 -838 14
rect -795 -14 -767 14
rect -724 -14 -696 14
rect -653 -14 -625 14
rect -582 -14 -554 14
rect -511 -14 -483 14
rect -440 -14 -412 14
rect -369 -14 -341 14
rect -298 -14 -270 14
rect -227 -14 -199 14
rect -156 -14 -128 14
rect -85 -14 -57 14
rect -14 -14 14 14
rect 57 -14 85 14
rect 128 -14 156 14
rect 199 -14 227 14
rect 270 -14 298 14
rect 341 -14 369 14
rect 412 -14 440 14
rect 483 -14 511 14
rect 554 -14 582 14
rect 625 -14 653 14
rect 696 -14 724 14
rect 767 -14 795 14
rect 838 -14 866 14
rect 909 -14 937 14
rect 980 -14 1008 14
rect 1051 -14 1079 14
rect 1122 -14 1150 14
rect 1193 -14 1221 14
rect 1264 -14 1292 14
rect 1335 -14 1363 14
rect 1406 -14 1434 14
rect 1477 -14 1505 14
rect 1548 -14 1576 14
rect 1619 -14 1647 14
rect 1690 -14 1718 14
rect 1761 -14 1789 14
rect 1832 -14 1860 14
rect 1903 -14 1931 14
rect 1974 -14 2002 14
rect 2045 -14 2073 14
rect 2116 -14 2144 14
rect 2187 -14 2215 14
rect 2258 -14 2286 14
rect 2329 -14 2357 14
rect 2400 -14 2428 14
rect 2471 -14 2499 14
rect 2542 -14 2570 14
rect 2613 -14 2641 14
rect 2684 -14 2712 14
rect 2755 -14 2783 14
rect -2783 -85 -2755 -57
rect -2712 -85 -2684 -57
rect -2641 -85 -2613 -57
rect -2570 -85 -2542 -57
rect -2499 -85 -2471 -57
rect -2428 -85 -2400 -57
rect -2357 -85 -2329 -57
rect -2286 -85 -2258 -57
rect -2215 -85 -2187 -57
rect -2144 -85 -2116 -57
rect -2073 -85 -2045 -57
rect -2002 -85 -1974 -57
rect -1931 -85 -1903 -57
rect -1860 -85 -1832 -57
rect -1789 -85 -1761 -57
rect -1718 -85 -1690 -57
rect -1647 -85 -1619 -57
rect -1576 -85 -1548 -57
rect -1505 -85 -1477 -57
rect -1434 -85 -1406 -57
rect -1363 -85 -1335 -57
rect -1292 -85 -1264 -57
rect -1221 -85 -1193 -57
rect -1150 -85 -1122 -57
rect -1079 -85 -1051 -57
rect -1008 -85 -980 -57
rect -937 -85 -909 -57
rect -866 -85 -838 -57
rect -795 -85 -767 -57
rect -724 -85 -696 -57
rect -653 -85 -625 -57
rect -582 -85 -554 -57
rect -511 -85 -483 -57
rect -440 -85 -412 -57
rect -369 -85 -341 -57
rect -298 -85 -270 -57
rect -227 -85 -199 -57
rect -156 -85 -128 -57
rect -85 -85 -57 -57
rect -14 -85 14 -57
rect 57 -85 85 -57
rect 128 -85 156 -57
rect 199 -85 227 -57
rect 270 -85 298 -57
rect 341 -85 369 -57
rect 412 -85 440 -57
rect 483 -85 511 -57
rect 554 -85 582 -57
rect 625 -85 653 -57
rect 696 -85 724 -57
rect 767 -85 795 -57
rect 838 -85 866 -57
rect 909 -85 937 -57
rect 980 -85 1008 -57
rect 1051 -85 1079 -57
rect 1122 -85 1150 -57
rect 1193 -85 1221 -57
rect 1264 -85 1292 -57
rect 1335 -85 1363 -57
rect 1406 -85 1434 -57
rect 1477 -85 1505 -57
rect 1548 -85 1576 -57
rect 1619 -85 1647 -57
rect 1690 -85 1718 -57
rect 1761 -85 1789 -57
rect 1832 -85 1860 -57
rect 1903 -85 1931 -57
rect 1974 -85 2002 -57
rect 2045 -85 2073 -57
rect 2116 -85 2144 -57
rect 2187 -85 2215 -57
rect 2258 -85 2286 -57
rect 2329 -85 2357 -57
rect 2400 -85 2428 -57
rect 2471 -85 2499 -57
rect 2542 -85 2570 -57
rect 2613 -85 2641 -57
rect 2684 -85 2712 -57
rect 2755 -85 2783 -57
<< metal3 >>
rect -2788 85 2788 90
rect -2788 57 -2783 85
rect -2755 57 -2712 85
rect -2684 57 -2641 85
rect -2613 57 -2570 85
rect -2542 57 -2499 85
rect -2471 57 -2428 85
rect -2400 57 -2357 85
rect -2329 57 -2286 85
rect -2258 57 -2215 85
rect -2187 57 -2144 85
rect -2116 57 -2073 85
rect -2045 57 -2002 85
rect -1974 57 -1931 85
rect -1903 57 -1860 85
rect -1832 57 -1789 85
rect -1761 57 -1718 85
rect -1690 57 -1647 85
rect -1619 57 -1576 85
rect -1548 57 -1505 85
rect -1477 57 -1434 85
rect -1406 57 -1363 85
rect -1335 57 -1292 85
rect -1264 57 -1221 85
rect -1193 57 -1150 85
rect -1122 57 -1079 85
rect -1051 57 -1008 85
rect -980 57 -937 85
rect -909 57 -866 85
rect -838 57 -795 85
rect -767 57 -724 85
rect -696 57 -653 85
rect -625 57 -582 85
rect -554 57 -511 85
rect -483 57 -440 85
rect -412 57 -369 85
rect -341 57 -298 85
rect -270 57 -227 85
rect -199 57 -156 85
rect -128 57 -85 85
rect -57 57 -14 85
rect 14 57 57 85
rect 85 57 128 85
rect 156 57 199 85
rect 227 57 270 85
rect 298 57 341 85
rect 369 57 412 85
rect 440 57 483 85
rect 511 57 554 85
rect 582 57 625 85
rect 653 57 696 85
rect 724 57 767 85
rect 795 57 838 85
rect 866 57 909 85
rect 937 57 980 85
rect 1008 57 1051 85
rect 1079 57 1122 85
rect 1150 57 1193 85
rect 1221 57 1264 85
rect 1292 57 1335 85
rect 1363 57 1406 85
rect 1434 57 1477 85
rect 1505 57 1548 85
rect 1576 57 1619 85
rect 1647 57 1690 85
rect 1718 57 1761 85
rect 1789 57 1832 85
rect 1860 57 1903 85
rect 1931 57 1974 85
rect 2002 57 2045 85
rect 2073 57 2116 85
rect 2144 57 2187 85
rect 2215 57 2258 85
rect 2286 57 2329 85
rect 2357 57 2400 85
rect 2428 57 2471 85
rect 2499 57 2542 85
rect 2570 57 2613 85
rect 2641 57 2684 85
rect 2712 57 2755 85
rect 2783 57 2788 85
rect -2788 14 2788 57
rect -2788 -14 -2783 14
rect -2755 -14 -2712 14
rect -2684 -14 -2641 14
rect -2613 -14 -2570 14
rect -2542 -14 -2499 14
rect -2471 -14 -2428 14
rect -2400 -14 -2357 14
rect -2329 -14 -2286 14
rect -2258 -14 -2215 14
rect -2187 -14 -2144 14
rect -2116 -14 -2073 14
rect -2045 -14 -2002 14
rect -1974 -14 -1931 14
rect -1903 -14 -1860 14
rect -1832 -14 -1789 14
rect -1761 -14 -1718 14
rect -1690 -14 -1647 14
rect -1619 -14 -1576 14
rect -1548 -14 -1505 14
rect -1477 -14 -1434 14
rect -1406 -14 -1363 14
rect -1335 -14 -1292 14
rect -1264 -14 -1221 14
rect -1193 -14 -1150 14
rect -1122 -14 -1079 14
rect -1051 -14 -1008 14
rect -980 -14 -937 14
rect -909 -14 -866 14
rect -838 -14 -795 14
rect -767 -14 -724 14
rect -696 -14 -653 14
rect -625 -14 -582 14
rect -554 -14 -511 14
rect -483 -14 -440 14
rect -412 -14 -369 14
rect -341 -14 -298 14
rect -270 -14 -227 14
rect -199 -14 -156 14
rect -128 -14 -85 14
rect -57 -14 -14 14
rect 14 -14 57 14
rect 85 -14 128 14
rect 156 -14 199 14
rect 227 -14 270 14
rect 298 -14 341 14
rect 369 -14 412 14
rect 440 -14 483 14
rect 511 -14 554 14
rect 582 -14 625 14
rect 653 -14 696 14
rect 724 -14 767 14
rect 795 -14 838 14
rect 866 -14 909 14
rect 937 -14 980 14
rect 1008 -14 1051 14
rect 1079 -14 1122 14
rect 1150 -14 1193 14
rect 1221 -14 1264 14
rect 1292 -14 1335 14
rect 1363 -14 1406 14
rect 1434 -14 1477 14
rect 1505 -14 1548 14
rect 1576 -14 1619 14
rect 1647 -14 1690 14
rect 1718 -14 1761 14
rect 1789 -14 1832 14
rect 1860 -14 1903 14
rect 1931 -14 1974 14
rect 2002 -14 2045 14
rect 2073 -14 2116 14
rect 2144 -14 2187 14
rect 2215 -14 2258 14
rect 2286 -14 2329 14
rect 2357 -14 2400 14
rect 2428 -14 2471 14
rect 2499 -14 2542 14
rect 2570 -14 2613 14
rect 2641 -14 2684 14
rect 2712 -14 2755 14
rect 2783 -14 2788 14
rect -2788 -57 2788 -14
rect -2788 -85 -2783 -57
rect -2755 -85 -2712 -57
rect -2684 -85 -2641 -57
rect -2613 -85 -2570 -57
rect -2542 -85 -2499 -57
rect -2471 -85 -2428 -57
rect -2400 -85 -2357 -57
rect -2329 -85 -2286 -57
rect -2258 -85 -2215 -57
rect -2187 -85 -2144 -57
rect -2116 -85 -2073 -57
rect -2045 -85 -2002 -57
rect -1974 -85 -1931 -57
rect -1903 -85 -1860 -57
rect -1832 -85 -1789 -57
rect -1761 -85 -1718 -57
rect -1690 -85 -1647 -57
rect -1619 -85 -1576 -57
rect -1548 -85 -1505 -57
rect -1477 -85 -1434 -57
rect -1406 -85 -1363 -57
rect -1335 -85 -1292 -57
rect -1264 -85 -1221 -57
rect -1193 -85 -1150 -57
rect -1122 -85 -1079 -57
rect -1051 -85 -1008 -57
rect -980 -85 -937 -57
rect -909 -85 -866 -57
rect -838 -85 -795 -57
rect -767 -85 -724 -57
rect -696 -85 -653 -57
rect -625 -85 -582 -57
rect -554 -85 -511 -57
rect -483 -85 -440 -57
rect -412 -85 -369 -57
rect -341 -85 -298 -57
rect -270 -85 -227 -57
rect -199 -85 -156 -57
rect -128 -85 -85 -57
rect -57 -85 -14 -57
rect 14 -85 57 -57
rect 85 -85 128 -57
rect 156 -85 199 -57
rect 227 -85 270 -57
rect 298 -85 341 -57
rect 369 -85 412 -57
rect 440 -85 483 -57
rect 511 -85 554 -57
rect 582 -85 625 -57
rect 653 -85 696 -57
rect 724 -85 767 -57
rect 795 -85 838 -57
rect 866 -85 909 -57
rect 937 -85 980 -57
rect 1008 -85 1051 -57
rect 1079 -85 1122 -57
rect 1150 -85 1193 -57
rect 1221 -85 1264 -57
rect 1292 -85 1335 -57
rect 1363 -85 1406 -57
rect 1434 -85 1477 -57
rect 1505 -85 1548 -57
rect 1576 -85 1619 -57
rect 1647 -85 1690 -57
rect 1718 -85 1761 -57
rect 1789 -85 1832 -57
rect 1860 -85 1903 -57
rect 1931 -85 1974 -57
rect 2002 -85 2045 -57
rect 2073 -85 2116 -57
rect 2144 -85 2187 -57
rect 2215 -85 2258 -57
rect 2286 -85 2329 -57
rect 2357 -85 2400 -57
rect 2428 -85 2471 -57
rect 2499 -85 2542 -57
rect 2570 -85 2613 -57
rect 2641 -85 2684 -57
rect 2712 -85 2755 -57
rect 2783 -85 2788 -57
rect -2788 -90 2788 -85
<< end >>
