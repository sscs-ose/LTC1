magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1123 -1019 1123 1019
<< metal1 >>
rect -123 13 123 19
rect -123 -13 -117 13
rect 117 -13 123 13
rect -123 -19 123 -13
<< via1 >>
rect -117 -13 117 13
<< metal2 >>
rect -123 13 123 19
rect -123 -13 -117 13
rect 117 -13 123 13
rect -123 -19 123 -13
<< end >>
