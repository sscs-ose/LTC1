magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2083 -1989 3139 4586
<< nwell >>
rect -83 1292 1139 2586
<< polysilicon >>
rect 336 925 476 1883
rect 580 925 720 1883
<< metal1 >>
rect 79 2424 165 2492
rect 246 1633 322 2476
rect 490 1088 566 2233
rect 734 1633 810 2476
rect 891 2424 977 2492
rect 490 1012 810 1088
rect 79 22 165 90
rect 246 35 322 881
rect 734 281 810 1012
rect 891 22 977 90
use M1_NWELL_CDNS_40661953145218  M1_NWELL_CDNS_40661953145218_0
timestamp 1713338890
transform 1 0 528 0 1 2458
box -457 -128 457 128
use M1_NWELL_CDNS_40661953145315  M1_NWELL_CDNS_40661953145315_0
timestamp 1713338890
transform 1 0 45 0 1 1988
box -128 -598 128 598
use M1_NWELL_CDNS_40661953145315  M1_NWELL_CDNS_40661953145315_1
timestamp 1713338890
transform 1 0 1011 0 1 1988
box -128 -598 128 598
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_0
timestamp 1713338890
transform 1 0 406 0 1 1263
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_1
timestamp 1713338890
transform 1 0 650 0 1 1263
box -42 -89 42 89
use M1_PSUB_CDNS_69033583165609  M1_PSUB_CDNS_69033583165609_0
timestamp 1713338890
transform 1 0 45 0 -1 526
box -45 -515 45 515
use M1_PSUB_CDNS_69033583165609  M1_PSUB_CDNS_69033583165609_1
timestamp 1713338890
transform 1 0 1011 0 -1 526
box -45 -515 45 515
use M1_PSUB_CDNS_69033583165613  M1_PSUB_CDNS_69033583165613_0
timestamp 1713338890
transform 1 0 528 0 -1 56
box -374 -45 374 45
use nmos_6p0_CDNS_4066195314511  nmos_6p0_CDNS_4066195314511_0
timestamp 1713338890
transform 1 0 580 0 1 281
box -88 -44 228 644
use nmos_6p0_CDNS_4066195314511  nmos_6p0_CDNS_4066195314511_1
timestamp 1713338890
transform 1 0 336 0 1 281
box -88 -44 228 644
use pmos_6p0_CDNS_4066195314512  pmos_6p0_CDNS_4066195314512_0
timestamp 1713338890
transform 1 0 336 0 1 1633
box -208 -120 348 720
use pmos_6p0_CDNS_4066195314512  pmos_6p0_CDNS_4066195314512_1
timestamp 1713338890
transform -1 0 720 0 1 1633
box -208 -120 348 720
<< labels >>
rlabel metal1 s 528 1268 528 1268 4 Z
port 1 nsew
rlabel metal1 s 652 1268 652 1268 4 B
port 2 nsew
rlabel metal1 s 407 1268 407 1268 4 A
port 3 nsew
rlabel metal1 s 244 56 244 56 4 VSS
port 4 nsew
rlabel metal1 s 75 2463 75 2463 4 VDD
port 5 nsew
<< end >>
