magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -2276 -2180 2276 2180
<< pwell >>
rect -276 -180 276 180
<< nmos >>
rect -164 -112 -52 112
rect 52 -112 164 112
<< ndiff >>
rect -252 70 -164 112
rect -252 -70 -239 70
rect -193 -70 -164 70
rect -252 -112 -164 -70
rect -52 70 52 112
rect -52 -70 -23 70
rect 23 -70 52 70
rect -52 -112 52 -70
rect 164 70 252 112
rect 164 -70 193 70
rect 239 -70 252 70
rect 164 -112 252 -70
<< ndiffc >>
rect -239 -70 -193 70
rect -23 -70 23 70
rect 193 -70 239 70
<< polysilicon >>
rect -164 112 -52 156
rect 52 112 164 156
rect -164 -156 -52 -112
rect 52 -156 164 -112
<< metal1 >>
rect -239 70 -193 110
rect -239 -110 -193 -70
rect -23 70 23 110
rect -23 -110 23 -70
rect 193 70 239 110
rect 193 -110 239 -70
<< end >>
