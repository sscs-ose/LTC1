magic
tech gf180mcuC
magscale 1 10
timestamp 1695206022
<< metal1 >>
rect -2010 5830 12900 6270
rect 10384 5333 12913 5371
rect 10384 5275 12765 5333
rect 12842 5275 12913 5333
rect 10384 5239 12913 5275
rect -424 2955 -351 2968
rect -424 2889 -411 2955
rect -356 2889 -351 2955
rect -424 2880 -351 2889
rect 40 1375 303 1521
rect 500 1097 620 1110
rect 500 1045 518 1097
rect 606 1045 620 1097
rect 500 1039 620 1045
rect 488 1038 620 1039
rect 107 575 312 596
rect 107 441 128 575
rect 279 441 312 575
rect 107 432 312 441
rect 488 -483 623 1038
rect 2430 994 2539 1512
rect 3374 1365 3699 1537
rect 3754 994 3863 1512
rect 4672 994 4781 1521
rect 5369 994 5478 1518
rect 6104 994 6213 1509
rect 6916 994 7025 1526
rect 7709 994 7818 1490
rect 8487 994 8596 1524
rect 9602 994 9711 1490
rect 10822 994 10931 1466
rect 11519 994 11628 1490
rect 12146 994 12255 1490
rect 488 -555 862 -483
rect 493 -556 623 -555
rect -419 -881 740 -880
rect -419 -890 1140 -881
rect -430 -893 7738 -890
rect -430 -975 -412 -893
rect -360 -975 7884 -893
rect -430 -1046 7884 -975
rect -430 -1060 7897 -1046
rect -430 -1070 5030 -1060
rect -430 -1090 3020 -1070
rect -430 -1100 880 -1090
rect -430 -1220 -180 -1100
rect -30 -1220 320 -1100
rect 470 -1210 880 -1100
rect 1030 -1210 1350 -1090
rect 1500 -1210 1900 -1090
rect 2050 -1210 2460 -1090
rect 2610 -1190 3020 -1090
rect 3170 -1190 3640 -1070
rect 3790 -1080 5030 -1070
rect 3790 -1190 4260 -1080
rect 2610 -1200 4260 -1190
rect 4410 -1180 5030 -1080
rect 5180 -1080 7897 -1060
rect 5180 -1180 5710 -1080
rect 4410 -1200 5710 -1180
rect 5860 -1200 6380 -1080
rect 6530 -1100 7897 -1080
rect 6530 -1200 7050 -1100
rect 2610 -1210 7050 -1200
rect 470 -1220 7050 -1210
rect 7200 -1220 7897 -1100
rect -430 -1229 7897 -1220
rect 7757 -1990 7897 -1229
rect 12667 -1530 12911 -1461
rect 11184 -1990 11991 -1960
rect -1850 -2050 12040 -1990
rect -1850 -2070 3650 -2050
rect -1850 -2090 2450 -2070
rect -1850 -2100 880 -2090
rect -1850 -2110 320 -2100
rect -1850 -2230 -180 -2110
rect -30 -2220 320 -2110
rect 470 -2210 880 -2100
rect 1030 -2210 1340 -2090
rect 1490 -2210 1900 -2090
rect 2050 -2190 2450 -2090
rect 2600 -2080 3650 -2070
rect 2600 -2190 3020 -2080
rect 2050 -2200 3020 -2190
rect 3170 -2170 3650 -2080
rect 3800 -2170 4260 -2050
rect 4410 -2060 12040 -2050
rect 4410 -2070 6380 -2060
rect 4410 -2170 5020 -2070
rect 3170 -2190 5020 -2170
rect 5170 -2190 5710 -2070
rect 5860 -2180 6380 -2070
rect 6530 -2180 7060 -2060
rect 7210 -2180 12040 -2060
rect 5860 -2190 12040 -2180
rect 3170 -2200 12040 -2190
rect 2050 -2210 12040 -2200
rect 470 -2220 12040 -2210
rect -30 -2230 12040 -2220
rect -1850 -2330 12040 -2230
<< via1 >>
rect 12765 5275 12842 5333
rect -411 2889 -356 2955
rect 518 1045 606 1097
rect 128 441 279 575
rect -412 -975 -360 -893
rect -180 -1220 -30 -1100
rect 320 -1220 470 -1100
rect 880 -1210 1030 -1090
rect 1350 -1210 1500 -1090
rect 1900 -1210 2050 -1090
rect 2460 -1210 2610 -1090
rect 3020 -1190 3170 -1070
rect 3640 -1190 3790 -1070
rect 4260 -1200 4410 -1080
rect 5030 -1180 5180 -1060
rect 5710 -1200 5860 -1080
rect 6380 -1200 6530 -1080
rect 7050 -1220 7200 -1100
rect -180 -2230 -30 -2110
rect 320 -2220 470 -2100
rect 880 -2210 1030 -2090
rect 1340 -2210 1490 -2090
rect 1900 -2210 2050 -2090
rect 2450 -2190 2600 -2070
rect 3020 -2200 3170 -2080
rect 3650 -2170 3800 -2050
rect 4260 -2170 4410 -2050
rect 5020 -2190 5170 -2070
rect 5710 -2190 5860 -2070
rect 6380 -2180 6530 -2060
rect 7060 -2180 7210 -2060
<< metal2 >>
rect 12790 5345 12903 5347
rect 12748 5333 12903 5345
rect 12748 5275 12765 5333
rect 12842 5275 12903 5333
rect 12748 5255 12903 5275
rect -434 2955 -291 2977
rect -434 2889 -411 2955
rect -356 2889 -291 2955
rect -434 -893 -291 2889
rect 12766 1314 12903 5255
rect 500 1223 1787 1314
rect 2023 1258 12903 1314
rect 2021 1223 12903 1258
rect 500 1137 12903 1223
rect 500 1097 620 1137
rect 500 1045 518 1097
rect 606 1045 620 1097
rect 1786 1091 2036 1137
rect 500 1020 620 1045
rect 107 575 312 596
rect 107 441 128 575
rect 279 441 312 575
rect 107 432 312 441
rect -434 -975 -412 -893
rect -360 -975 -291 -893
rect -434 -1033 -291 -975
rect -190 -1100 -10 -1080
rect -190 -1220 -180 -1100
rect -30 -1220 -10 -1100
rect -190 -2110 -10 -1220
rect -190 -2230 -180 -2110
rect -30 -2230 -10 -2110
rect -190 -2260 -10 -2230
rect 310 -1100 490 -1080
rect 310 -1220 320 -1100
rect 470 -1220 490 -1100
rect 310 -2100 490 -1220
rect 310 -2220 320 -2100
rect 470 -2220 490 -2100
rect 310 -2260 490 -2220
rect 870 -1090 1050 -1060
rect 870 -1210 880 -1090
rect 1030 -1210 1050 -1090
rect 870 -2090 1050 -1210
rect 870 -2210 880 -2090
rect 1030 -2210 1050 -2090
rect 870 -2240 1050 -2210
rect 1330 -1090 1510 -1080
rect 1330 -1210 1350 -1090
rect 1500 -1210 1510 -1090
rect 1330 -2090 1510 -1210
rect 1330 -2210 1340 -2090
rect 1490 -2210 1510 -2090
rect 1330 -2260 1510 -2210
rect 1880 -1090 2060 -1060
rect 1880 -1210 1900 -1090
rect 2050 -1210 2060 -1090
rect 1880 -2090 2060 -1210
rect 1880 -2210 1900 -2090
rect 2050 -2210 2060 -2090
rect 1880 -2240 2060 -2210
rect 2440 -1090 2620 -1060
rect 2440 -1210 2460 -1090
rect 2610 -1210 2620 -1090
rect 2440 -2070 2620 -1210
rect 2440 -2190 2450 -2070
rect 2600 -2190 2620 -2070
rect 2440 -2240 2620 -2190
rect 3010 -1070 3190 -1060
rect 3010 -1190 3020 -1070
rect 3170 -1190 3190 -1070
rect 3010 -2080 3190 -1190
rect 3010 -2200 3020 -2080
rect 3170 -2200 3190 -2080
rect 3010 -2240 3190 -2200
rect 3630 -1070 3810 -1050
rect 3630 -1190 3640 -1070
rect 3790 -1190 3810 -1070
rect 3630 -2050 3810 -1190
rect 3630 -2170 3650 -2050
rect 3800 -2170 3810 -2050
rect 3630 -2230 3810 -2170
rect 4250 -1080 4430 -1050
rect 4250 -1200 4260 -1080
rect 4410 -1200 4430 -1080
rect 4250 -2050 4430 -1200
rect 4250 -2170 4260 -2050
rect 4410 -2170 4430 -2050
rect 4250 -2230 4430 -2170
rect 5010 -1060 5190 -1040
rect 5010 -1180 5030 -1060
rect 5180 -1180 5190 -1060
rect 5010 -2070 5190 -1180
rect 5010 -2190 5020 -2070
rect 5170 -2190 5190 -2070
rect 5010 -2220 5190 -2190
rect 5700 -1080 5880 -1060
rect 5700 -1200 5710 -1080
rect 5860 -1200 5880 -1080
rect 5700 -2070 5880 -1200
rect 5700 -2190 5710 -2070
rect 5860 -2190 5880 -2070
rect 5700 -2240 5880 -2190
rect 6370 -1080 6550 -1070
rect 6370 -1200 6380 -1080
rect 6530 -1200 6550 -1080
rect 6370 -2060 6550 -1200
rect 6370 -2180 6380 -2060
rect 6530 -2180 6550 -2060
rect 6370 -2250 6550 -2180
rect 7040 -1100 7220 -1090
rect 7040 -1220 7050 -1100
rect 7200 -1220 7220 -1100
rect 7040 -2060 7220 -1220
rect 7040 -2180 7060 -2060
rect 7210 -2180 7220 -2060
rect 7040 -2270 7220 -2180
<< via2 >>
rect 128 441 279 575
<< metal3 >>
rect 1865 1493 1946 1581
rect 1860 1165 1946 1493
rect 107 575 312 596
rect 107 441 128 575
rect 279 558 312 575
rect 1865 558 1946 1165
rect 279 554 1946 558
rect 279 477 2623 554
rect 279 441 312 477
rect 107 432 312 441
use CLK_div_10_mag  CLK_div_10_mag_0
timestamp 1695206022
transform 1 0 740 0 -1 1103
box -34 0 12197 3533
use CLK_DIV_11_mag_new  CLK_DIV_11_mag_new_0
timestamp 1695206022
transform 1 0 -1735 0 -1 6681
box -827 763 15023 5476
<< labels >>
flabel metal1 4142 -1057 4142 -1057 0 FreeSans 640 0 0 0 VDD
port 0 nsew
flabel via2 194 515 194 515 0 FreeSans 640 0 0 0 RST
port 1 nsew
flabel metal1 143 1406 143 1406 0 FreeSans 640 0 0 0 CLK
port 2 nsew
flabel metal1 12846 -1493 12846 -1491 0 FreeSans 640 0 0 0 Vdiv110
port 3 nsew
flabel metal1 3512 1475 3512 1477 0 FreeSans 640 0 0 0 VSS
port 4 nsew
<< end >>
