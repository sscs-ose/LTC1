magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -3730 -2583 13766 12481
<< nwell >>
rect -1730 -583 -500 10481
rect 10573 -583 11766 10481
<< ndiff >>
rect -458 -500 10532 -98
<< psubdiff >>
rect -458 8756 10536 9430
rect -458 322 -118 8756
rect 10146 322 10536 8756
rect -458 254 254 322
rect 9819 254 10536 322
rect -458 32 10536 254
<< nsubdiff >>
rect -1647 9580 -500 10398
rect 10573 9580 11683 10398
rect -1647 8339 -583 9580
rect -1647 -449 -1587 8339
rect -1541 -449 -1483 8339
rect -1437 -449 -1379 8339
rect -1333 -449 -1275 8339
rect -1229 -449 -1171 8339
rect -1125 -449 -1067 8339
rect -1021 -449 -963 8339
rect -917 -449 -859 8339
rect -813 -449 -755 8339
rect -709 -449 -651 8339
rect -605 -98 -583 8339
rect 10656 8339 11683 9580
rect 10656 -98 10678 8339
rect -605 -449 -500 -98
rect -1647 -500 -500 -449
rect 10573 -449 10678 -98
rect 10724 -449 10782 8339
rect 10828 -449 10886 8339
rect 10932 -449 10990 8339
rect 11036 -449 11094 8339
rect 11140 -449 11198 8339
rect 11244 -449 11302 8339
rect 11348 -449 11406 8339
rect 11452 -449 11510 8339
rect 11556 -449 11614 8339
rect 11660 -449 11683 8339
rect 10573 -500 11683 -449
<< nsubdiffcont >>
rect -1587 -449 -1541 8339
rect -1483 -449 -1437 8339
rect -1379 -449 -1333 8339
rect -1275 -449 -1229 8339
rect -1171 -449 -1125 8339
rect -1067 -449 -1021 8339
rect -963 -449 -917 8339
rect -859 -449 -813 8339
rect -755 -449 -709 8339
rect -651 -449 -605 8339
rect 10678 -449 10724 8339
rect 10782 -449 10828 8339
rect 10886 -449 10932 8339
rect 10990 -449 11036 8339
rect 11094 -449 11140 8339
rect 11198 -449 11244 8339
rect 11302 -449 11348 8339
rect 11406 -449 11452 8339
rect 11510 -449 11556 8339
rect 11614 -449 11660 8339
<< metal1 >>
rect -1598 8339 -594 8388
rect -1598 -449 -1587 8339
rect -1541 -449 -1483 8339
rect -1437 -449 -1379 8339
rect -1333 -449 -1275 8339
rect -1229 -449 -1171 8339
rect -1125 -449 -1067 8339
rect -1021 -449 -963 8339
rect -917 -449 -859 8339
rect -813 -449 -755 8339
rect -709 -449 -651 8339
rect -605 -109 -594 8339
rect -457 311 111 8396
rect 9962 311 10530 8397
rect -457 43 10530 311
rect 10666 8339 11670 8410
rect 10666 -109 10678 8339
rect -605 -449 10678 -109
rect 10724 -449 10782 8339
rect 10828 -449 10886 8339
rect 10932 -449 10990 8339
rect 11036 -449 11094 8339
rect 11140 -449 11198 8339
rect 11244 -449 11302 8339
rect 11348 -449 11406 8339
rect 11452 -449 11510 8339
rect 11556 -449 11614 8339
rect 11660 -449 11670 8339
rect -1598 -489 11670 -449
use M1_NWELL_CDNS_40661953145373  M1_NWELL_CDNS_40661953145373_0
timestamp 1713338890
transform 1 0 5037 0 1 -299
box -5578 -284 5578 284
use M1_NWELL_CDNS_40661953145374  M1_NWELL_CDNS_40661953145374_0
timestamp 1713338890
transform 1 0 5037 0 1 9989
box -5578 -492 5578 492
use M1_PSUB_CDNS_69033583165667  M1_PSUB_CDNS_69033583165667_0
timestamp 1713338890
transform 0 -1 5034 1 0 177
box -145 -5045 145 5045
use M1_PSUB_CDNS_69033583165668  M1_PSUB_CDNS_69033583165668_0
timestamp 1713338890
transform 1 0 10346 0 1 4177
box -195 -4145 195 4145
use M1_PSUB_CDNS_69033583165669  M1_PSUB_CDNS_69033583165669_0
timestamp 1713338890
transform 1 0 -273 0 1 4177
box -145 -4145 145 4145
<< end >>
