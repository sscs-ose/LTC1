magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1349 -4385 1349 4385
<< metal3 >>
rect -349 3380 349 3385
rect -349 3352 -344 3380
rect -316 3352 -278 3380
rect -250 3352 -212 3380
rect -184 3352 -146 3380
rect -118 3352 -80 3380
rect -52 3352 -14 3380
rect 14 3352 52 3380
rect 80 3352 118 3380
rect 146 3352 184 3380
rect 212 3352 250 3380
rect 278 3352 316 3380
rect 344 3352 349 3380
rect -349 3314 349 3352
rect -349 3286 -344 3314
rect -316 3286 -278 3314
rect -250 3286 -212 3314
rect -184 3286 -146 3314
rect -118 3286 -80 3314
rect -52 3286 -14 3314
rect 14 3286 52 3314
rect 80 3286 118 3314
rect 146 3286 184 3314
rect 212 3286 250 3314
rect 278 3286 316 3314
rect 344 3286 349 3314
rect -349 3248 349 3286
rect -349 3220 -344 3248
rect -316 3220 -278 3248
rect -250 3220 -212 3248
rect -184 3220 -146 3248
rect -118 3220 -80 3248
rect -52 3220 -14 3248
rect 14 3220 52 3248
rect 80 3220 118 3248
rect 146 3220 184 3248
rect 212 3220 250 3248
rect 278 3220 316 3248
rect 344 3220 349 3248
rect -349 3182 349 3220
rect -349 3154 -344 3182
rect -316 3154 -278 3182
rect -250 3154 -212 3182
rect -184 3154 -146 3182
rect -118 3154 -80 3182
rect -52 3154 -14 3182
rect 14 3154 52 3182
rect 80 3154 118 3182
rect 146 3154 184 3182
rect 212 3154 250 3182
rect 278 3154 316 3182
rect 344 3154 349 3182
rect -349 3116 349 3154
rect -349 3088 -344 3116
rect -316 3088 -278 3116
rect -250 3088 -212 3116
rect -184 3088 -146 3116
rect -118 3088 -80 3116
rect -52 3088 -14 3116
rect 14 3088 52 3116
rect 80 3088 118 3116
rect 146 3088 184 3116
rect 212 3088 250 3116
rect 278 3088 316 3116
rect 344 3088 349 3116
rect -349 3050 349 3088
rect -349 3022 -344 3050
rect -316 3022 -278 3050
rect -250 3022 -212 3050
rect -184 3022 -146 3050
rect -118 3022 -80 3050
rect -52 3022 -14 3050
rect 14 3022 52 3050
rect 80 3022 118 3050
rect 146 3022 184 3050
rect 212 3022 250 3050
rect 278 3022 316 3050
rect 344 3022 349 3050
rect -349 2984 349 3022
rect -349 2956 -344 2984
rect -316 2956 -278 2984
rect -250 2956 -212 2984
rect -184 2956 -146 2984
rect -118 2956 -80 2984
rect -52 2956 -14 2984
rect 14 2956 52 2984
rect 80 2956 118 2984
rect 146 2956 184 2984
rect 212 2956 250 2984
rect 278 2956 316 2984
rect 344 2956 349 2984
rect -349 2918 349 2956
rect -349 2890 -344 2918
rect -316 2890 -278 2918
rect -250 2890 -212 2918
rect -184 2890 -146 2918
rect -118 2890 -80 2918
rect -52 2890 -14 2918
rect 14 2890 52 2918
rect 80 2890 118 2918
rect 146 2890 184 2918
rect 212 2890 250 2918
rect 278 2890 316 2918
rect 344 2890 349 2918
rect -349 2852 349 2890
rect -349 2824 -344 2852
rect -316 2824 -278 2852
rect -250 2824 -212 2852
rect -184 2824 -146 2852
rect -118 2824 -80 2852
rect -52 2824 -14 2852
rect 14 2824 52 2852
rect 80 2824 118 2852
rect 146 2824 184 2852
rect 212 2824 250 2852
rect 278 2824 316 2852
rect 344 2824 349 2852
rect -349 2786 349 2824
rect -349 2758 -344 2786
rect -316 2758 -278 2786
rect -250 2758 -212 2786
rect -184 2758 -146 2786
rect -118 2758 -80 2786
rect -52 2758 -14 2786
rect 14 2758 52 2786
rect 80 2758 118 2786
rect 146 2758 184 2786
rect 212 2758 250 2786
rect 278 2758 316 2786
rect 344 2758 349 2786
rect -349 2720 349 2758
rect -349 2692 -344 2720
rect -316 2692 -278 2720
rect -250 2692 -212 2720
rect -184 2692 -146 2720
rect -118 2692 -80 2720
rect -52 2692 -14 2720
rect 14 2692 52 2720
rect 80 2692 118 2720
rect 146 2692 184 2720
rect 212 2692 250 2720
rect 278 2692 316 2720
rect 344 2692 349 2720
rect -349 2654 349 2692
rect -349 2626 -344 2654
rect -316 2626 -278 2654
rect -250 2626 -212 2654
rect -184 2626 -146 2654
rect -118 2626 -80 2654
rect -52 2626 -14 2654
rect 14 2626 52 2654
rect 80 2626 118 2654
rect 146 2626 184 2654
rect 212 2626 250 2654
rect 278 2626 316 2654
rect 344 2626 349 2654
rect -349 2588 349 2626
rect -349 2560 -344 2588
rect -316 2560 -278 2588
rect -250 2560 -212 2588
rect -184 2560 -146 2588
rect -118 2560 -80 2588
rect -52 2560 -14 2588
rect 14 2560 52 2588
rect 80 2560 118 2588
rect 146 2560 184 2588
rect 212 2560 250 2588
rect 278 2560 316 2588
rect 344 2560 349 2588
rect -349 2522 349 2560
rect -349 2494 -344 2522
rect -316 2494 -278 2522
rect -250 2494 -212 2522
rect -184 2494 -146 2522
rect -118 2494 -80 2522
rect -52 2494 -14 2522
rect 14 2494 52 2522
rect 80 2494 118 2522
rect 146 2494 184 2522
rect 212 2494 250 2522
rect 278 2494 316 2522
rect 344 2494 349 2522
rect -349 2456 349 2494
rect -349 2428 -344 2456
rect -316 2428 -278 2456
rect -250 2428 -212 2456
rect -184 2428 -146 2456
rect -118 2428 -80 2456
rect -52 2428 -14 2456
rect 14 2428 52 2456
rect 80 2428 118 2456
rect 146 2428 184 2456
rect 212 2428 250 2456
rect 278 2428 316 2456
rect 344 2428 349 2456
rect -349 2390 349 2428
rect -349 2362 -344 2390
rect -316 2362 -278 2390
rect -250 2362 -212 2390
rect -184 2362 -146 2390
rect -118 2362 -80 2390
rect -52 2362 -14 2390
rect 14 2362 52 2390
rect 80 2362 118 2390
rect 146 2362 184 2390
rect 212 2362 250 2390
rect 278 2362 316 2390
rect 344 2362 349 2390
rect -349 2324 349 2362
rect -349 2296 -344 2324
rect -316 2296 -278 2324
rect -250 2296 -212 2324
rect -184 2296 -146 2324
rect -118 2296 -80 2324
rect -52 2296 -14 2324
rect 14 2296 52 2324
rect 80 2296 118 2324
rect 146 2296 184 2324
rect 212 2296 250 2324
rect 278 2296 316 2324
rect 344 2296 349 2324
rect -349 2258 349 2296
rect -349 2230 -344 2258
rect -316 2230 -278 2258
rect -250 2230 -212 2258
rect -184 2230 -146 2258
rect -118 2230 -80 2258
rect -52 2230 -14 2258
rect 14 2230 52 2258
rect 80 2230 118 2258
rect 146 2230 184 2258
rect 212 2230 250 2258
rect 278 2230 316 2258
rect 344 2230 349 2258
rect -349 2192 349 2230
rect -349 2164 -344 2192
rect -316 2164 -278 2192
rect -250 2164 -212 2192
rect -184 2164 -146 2192
rect -118 2164 -80 2192
rect -52 2164 -14 2192
rect 14 2164 52 2192
rect 80 2164 118 2192
rect 146 2164 184 2192
rect 212 2164 250 2192
rect 278 2164 316 2192
rect 344 2164 349 2192
rect -349 2126 349 2164
rect -349 2098 -344 2126
rect -316 2098 -278 2126
rect -250 2098 -212 2126
rect -184 2098 -146 2126
rect -118 2098 -80 2126
rect -52 2098 -14 2126
rect 14 2098 52 2126
rect 80 2098 118 2126
rect 146 2098 184 2126
rect 212 2098 250 2126
rect 278 2098 316 2126
rect 344 2098 349 2126
rect -349 2060 349 2098
rect -349 2032 -344 2060
rect -316 2032 -278 2060
rect -250 2032 -212 2060
rect -184 2032 -146 2060
rect -118 2032 -80 2060
rect -52 2032 -14 2060
rect 14 2032 52 2060
rect 80 2032 118 2060
rect 146 2032 184 2060
rect 212 2032 250 2060
rect 278 2032 316 2060
rect 344 2032 349 2060
rect -349 1994 349 2032
rect -349 1966 -344 1994
rect -316 1966 -278 1994
rect -250 1966 -212 1994
rect -184 1966 -146 1994
rect -118 1966 -80 1994
rect -52 1966 -14 1994
rect 14 1966 52 1994
rect 80 1966 118 1994
rect 146 1966 184 1994
rect 212 1966 250 1994
rect 278 1966 316 1994
rect 344 1966 349 1994
rect -349 1928 349 1966
rect -349 1900 -344 1928
rect -316 1900 -278 1928
rect -250 1900 -212 1928
rect -184 1900 -146 1928
rect -118 1900 -80 1928
rect -52 1900 -14 1928
rect 14 1900 52 1928
rect 80 1900 118 1928
rect 146 1900 184 1928
rect 212 1900 250 1928
rect 278 1900 316 1928
rect 344 1900 349 1928
rect -349 1862 349 1900
rect -349 1834 -344 1862
rect -316 1834 -278 1862
rect -250 1834 -212 1862
rect -184 1834 -146 1862
rect -118 1834 -80 1862
rect -52 1834 -14 1862
rect 14 1834 52 1862
rect 80 1834 118 1862
rect 146 1834 184 1862
rect 212 1834 250 1862
rect 278 1834 316 1862
rect 344 1834 349 1862
rect -349 1796 349 1834
rect -349 1768 -344 1796
rect -316 1768 -278 1796
rect -250 1768 -212 1796
rect -184 1768 -146 1796
rect -118 1768 -80 1796
rect -52 1768 -14 1796
rect 14 1768 52 1796
rect 80 1768 118 1796
rect 146 1768 184 1796
rect 212 1768 250 1796
rect 278 1768 316 1796
rect 344 1768 349 1796
rect -349 1730 349 1768
rect -349 1702 -344 1730
rect -316 1702 -278 1730
rect -250 1702 -212 1730
rect -184 1702 -146 1730
rect -118 1702 -80 1730
rect -52 1702 -14 1730
rect 14 1702 52 1730
rect 80 1702 118 1730
rect 146 1702 184 1730
rect 212 1702 250 1730
rect 278 1702 316 1730
rect 344 1702 349 1730
rect -349 1664 349 1702
rect -349 1636 -344 1664
rect -316 1636 -278 1664
rect -250 1636 -212 1664
rect -184 1636 -146 1664
rect -118 1636 -80 1664
rect -52 1636 -14 1664
rect 14 1636 52 1664
rect 80 1636 118 1664
rect 146 1636 184 1664
rect 212 1636 250 1664
rect 278 1636 316 1664
rect 344 1636 349 1664
rect -349 1598 349 1636
rect -349 1570 -344 1598
rect -316 1570 -278 1598
rect -250 1570 -212 1598
rect -184 1570 -146 1598
rect -118 1570 -80 1598
rect -52 1570 -14 1598
rect 14 1570 52 1598
rect 80 1570 118 1598
rect 146 1570 184 1598
rect 212 1570 250 1598
rect 278 1570 316 1598
rect 344 1570 349 1598
rect -349 1532 349 1570
rect -349 1504 -344 1532
rect -316 1504 -278 1532
rect -250 1504 -212 1532
rect -184 1504 -146 1532
rect -118 1504 -80 1532
rect -52 1504 -14 1532
rect 14 1504 52 1532
rect 80 1504 118 1532
rect 146 1504 184 1532
rect 212 1504 250 1532
rect 278 1504 316 1532
rect 344 1504 349 1532
rect -349 1466 349 1504
rect -349 1438 -344 1466
rect -316 1438 -278 1466
rect -250 1438 -212 1466
rect -184 1438 -146 1466
rect -118 1438 -80 1466
rect -52 1438 -14 1466
rect 14 1438 52 1466
rect 80 1438 118 1466
rect 146 1438 184 1466
rect 212 1438 250 1466
rect 278 1438 316 1466
rect 344 1438 349 1466
rect -349 1400 349 1438
rect -349 1372 -344 1400
rect -316 1372 -278 1400
rect -250 1372 -212 1400
rect -184 1372 -146 1400
rect -118 1372 -80 1400
rect -52 1372 -14 1400
rect 14 1372 52 1400
rect 80 1372 118 1400
rect 146 1372 184 1400
rect 212 1372 250 1400
rect 278 1372 316 1400
rect 344 1372 349 1400
rect -349 1334 349 1372
rect -349 1306 -344 1334
rect -316 1306 -278 1334
rect -250 1306 -212 1334
rect -184 1306 -146 1334
rect -118 1306 -80 1334
rect -52 1306 -14 1334
rect 14 1306 52 1334
rect 80 1306 118 1334
rect 146 1306 184 1334
rect 212 1306 250 1334
rect 278 1306 316 1334
rect 344 1306 349 1334
rect -349 1268 349 1306
rect -349 1240 -344 1268
rect -316 1240 -278 1268
rect -250 1240 -212 1268
rect -184 1240 -146 1268
rect -118 1240 -80 1268
rect -52 1240 -14 1268
rect 14 1240 52 1268
rect 80 1240 118 1268
rect 146 1240 184 1268
rect 212 1240 250 1268
rect 278 1240 316 1268
rect 344 1240 349 1268
rect -349 1202 349 1240
rect -349 1174 -344 1202
rect -316 1174 -278 1202
rect -250 1174 -212 1202
rect -184 1174 -146 1202
rect -118 1174 -80 1202
rect -52 1174 -14 1202
rect 14 1174 52 1202
rect 80 1174 118 1202
rect 146 1174 184 1202
rect 212 1174 250 1202
rect 278 1174 316 1202
rect 344 1174 349 1202
rect -349 1136 349 1174
rect -349 1108 -344 1136
rect -316 1108 -278 1136
rect -250 1108 -212 1136
rect -184 1108 -146 1136
rect -118 1108 -80 1136
rect -52 1108 -14 1136
rect 14 1108 52 1136
rect 80 1108 118 1136
rect 146 1108 184 1136
rect 212 1108 250 1136
rect 278 1108 316 1136
rect 344 1108 349 1136
rect -349 1070 349 1108
rect -349 1042 -344 1070
rect -316 1042 -278 1070
rect -250 1042 -212 1070
rect -184 1042 -146 1070
rect -118 1042 -80 1070
rect -52 1042 -14 1070
rect 14 1042 52 1070
rect 80 1042 118 1070
rect 146 1042 184 1070
rect 212 1042 250 1070
rect 278 1042 316 1070
rect 344 1042 349 1070
rect -349 1004 349 1042
rect -349 976 -344 1004
rect -316 976 -278 1004
rect -250 976 -212 1004
rect -184 976 -146 1004
rect -118 976 -80 1004
rect -52 976 -14 1004
rect 14 976 52 1004
rect 80 976 118 1004
rect 146 976 184 1004
rect 212 976 250 1004
rect 278 976 316 1004
rect 344 976 349 1004
rect -349 938 349 976
rect -349 910 -344 938
rect -316 910 -278 938
rect -250 910 -212 938
rect -184 910 -146 938
rect -118 910 -80 938
rect -52 910 -14 938
rect 14 910 52 938
rect 80 910 118 938
rect 146 910 184 938
rect 212 910 250 938
rect 278 910 316 938
rect 344 910 349 938
rect -349 872 349 910
rect -349 844 -344 872
rect -316 844 -278 872
rect -250 844 -212 872
rect -184 844 -146 872
rect -118 844 -80 872
rect -52 844 -14 872
rect 14 844 52 872
rect 80 844 118 872
rect 146 844 184 872
rect 212 844 250 872
rect 278 844 316 872
rect 344 844 349 872
rect -349 806 349 844
rect -349 778 -344 806
rect -316 778 -278 806
rect -250 778 -212 806
rect -184 778 -146 806
rect -118 778 -80 806
rect -52 778 -14 806
rect 14 778 52 806
rect 80 778 118 806
rect 146 778 184 806
rect 212 778 250 806
rect 278 778 316 806
rect 344 778 349 806
rect -349 740 349 778
rect -349 712 -344 740
rect -316 712 -278 740
rect -250 712 -212 740
rect -184 712 -146 740
rect -118 712 -80 740
rect -52 712 -14 740
rect 14 712 52 740
rect 80 712 118 740
rect 146 712 184 740
rect 212 712 250 740
rect 278 712 316 740
rect 344 712 349 740
rect -349 674 349 712
rect -349 646 -344 674
rect -316 646 -278 674
rect -250 646 -212 674
rect -184 646 -146 674
rect -118 646 -80 674
rect -52 646 -14 674
rect 14 646 52 674
rect 80 646 118 674
rect 146 646 184 674
rect 212 646 250 674
rect 278 646 316 674
rect 344 646 349 674
rect -349 608 349 646
rect -349 580 -344 608
rect -316 580 -278 608
rect -250 580 -212 608
rect -184 580 -146 608
rect -118 580 -80 608
rect -52 580 -14 608
rect 14 580 52 608
rect 80 580 118 608
rect 146 580 184 608
rect 212 580 250 608
rect 278 580 316 608
rect 344 580 349 608
rect -349 542 349 580
rect -349 514 -344 542
rect -316 514 -278 542
rect -250 514 -212 542
rect -184 514 -146 542
rect -118 514 -80 542
rect -52 514 -14 542
rect 14 514 52 542
rect 80 514 118 542
rect 146 514 184 542
rect 212 514 250 542
rect 278 514 316 542
rect 344 514 349 542
rect -349 476 349 514
rect -349 448 -344 476
rect -316 448 -278 476
rect -250 448 -212 476
rect -184 448 -146 476
rect -118 448 -80 476
rect -52 448 -14 476
rect 14 448 52 476
rect 80 448 118 476
rect 146 448 184 476
rect 212 448 250 476
rect 278 448 316 476
rect 344 448 349 476
rect -349 410 349 448
rect -349 382 -344 410
rect -316 382 -278 410
rect -250 382 -212 410
rect -184 382 -146 410
rect -118 382 -80 410
rect -52 382 -14 410
rect 14 382 52 410
rect 80 382 118 410
rect 146 382 184 410
rect 212 382 250 410
rect 278 382 316 410
rect 344 382 349 410
rect -349 344 349 382
rect -349 316 -344 344
rect -316 316 -278 344
rect -250 316 -212 344
rect -184 316 -146 344
rect -118 316 -80 344
rect -52 316 -14 344
rect 14 316 52 344
rect 80 316 118 344
rect 146 316 184 344
rect 212 316 250 344
rect 278 316 316 344
rect 344 316 349 344
rect -349 278 349 316
rect -349 250 -344 278
rect -316 250 -278 278
rect -250 250 -212 278
rect -184 250 -146 278
rect -118 250 -80 278
rect -52 250 -14 278
rect 14 250 52 278
rect 80 250 118 278
rect 146 250 184 278
rect 212 250 250 278
rect 278 250 316 278
rect 344 250 349 278
rect -349 212 349 250
rect -349 184 -344 212
rect -316 184 -278 212
rect -250 184 -212 212
rect -184 184 -146 212
rect -118 184 -80 212
rect -52 184 -14 212
rect 14 184 52 212
rect 80 184 118 212
rect 146 184 184 212
rect 212 184 250 212
rect 278 184 316 212
rect 344 184 349 212
rect -349 146 349 184
rect -349 118 -344 146
rect -316 118 -278 146
rect -250 118 -212 146
rect -184 118 -146 146
rect -118 118 -80 146
rect -52 118 -14 146
rect 14 118 52 146
rect 80 118 118 146
rect 146 118 184 146
rect 212 118 250 146
rect 278 118 316 146
rect 344 118 349 146
rect -349 80 349 118
rect -349 52 -344 80
rect -316 52 -278 80
rect -250 52 -212 80
rect -184 52 -146 80
rect -118 52 -80 80
rect -52 52 -14 80
rect 14 52 52 80
rect 80 52 118 80
rect 146 52 184 80
rect 212 52 250 80
rect 278 52 316 80
rect 344 52 349 80
rect -349 14 349 52
rect -349 -14 -344 14
rect -316 -14 -278 14
rect -250 -14 -212 14
rect -184 -14 -146 14
rect -118 -14 -80 14
rect -52 -14 -14 14
rect 14 -14 52 14
rect 80 -14 118 14
rect 146 -14 184 14
rect 212 -14 250 14
rect 278 -14 316 14
rect 344 -14 349 14
rect -349 -52 349 -14
rect -349 -80 -344 -52
rect -316 -80 -278 -52
rect -250 -80 -212 -52
rect -184 -80 -146 -52
rect -118 -80 -80 -52
rect -52 -80 -14 -52
rect 14 -80 52 -52
rect 80 -80 118 -52
rect 146 -80 184 -52
rect 212 -80 250 -52
rect 278 -80 316 -52
rect 344 -80 349 -52
rect -349 -118 349 -80
rect -349 -146 -344 -118
rect -316 -146 -278 -118
rect -250 -146 -212 -118
rect -184 -146 -146 -118
rect -118 -146 -80 -118
rect -52 -146 -14 -118
rect 14 -146 52 -118
rect 80 -146 118 -118
rect 146 -146 184 -118
rect 212 -146 250 -118
rect 278 -146 316 -118
rect 344 -146 349 -118
rect -349 -184 349 -146
rect -349 -212 -344 -184
rect -316 -212 -278 -184
rect -250 -212 -212 -184
rect -184 -212 -146 -184
rect -118 -212 -80 -184
rect -52 -212 -14 -184
rect 14 -212 52 -184
rect 80 -212 118 -184
rect 146 -212 184 -184
rect 212 -212 250 -184
rect 278 -212 316 -184
rect 344 -212 349 -184
rect -349 -250 349 -212
rect -349 -278 -344 -250
rect -316 -278 -278 -250
rect -250 -278 -212 -250
rect -184 -278 -146 -250
rect -118 -278 -80 -250
rect -52 -278 -14 -250
rect 14 -278 52 -250
rect 80 -278 118 -250
rect 146 -278 184 -250
rect 212 -278 250 -250
rect 278 -278 316 -250
rect 344 -278 349 -250
rect -349 -316 349 -278
rect -349 -344 -344 -316
rect -316 -344 -278 -316
rect -250 -344 -212 -316
rect -184 -344 -146 -316
rect -118 -344 -80 -316
rect -52 -344 -14 -316
rect 14 -344 52 -316
rect 80 -344 118 -316
rect 146 -344 184 -316
rect 212 -344 250 -316
rect 278 -344 316 -316
rect 344 -344 349 -316
rect -349 -382 349 -344
rect -349 -410 -344 -382
rect -316 -410 -278 -382
rect -250 -410 -212 -382
rect -184 -410 -146 -382
rect -118 -410 -80 -382
rect -52 -410 -14 -382
rect 14 -410 52 -382
rect 80 -410 118 -382
rect 146 -410 184 -382
rect 212 -410 250 -382
rect 278 -410 316 -382
rect 344 -410 349 -382
rect -349 -448 349 -410
rect -349 -476 -344 -448
rect -316 -476 -278 -448
rect -250 -476 -212 -448
rect -184 -476 -146 -448
rect -118 -476 -80 -448
rect -52 -476 -14 -448
rect 14 -476 52 -448
rect 80 -476 118 -448
rect 146 -476 184 -448
rect 212 -476 250 -448
rect 278 -476 316 -448
rect 344 -476 349 -448
rect -349 -514 349 -476
rect -349 -542 -344 -514
rect -316 -542 -278 -514
rect -250 -542 -212 -514
rect -184 -542 -146 -514
rect -118 -542 -80 -514
rect -52 -542 -14 -514
rect 14 -542 52 -514
rect 80 -542 118 -514
rect 146 -542 184 -514
rect 212 -542 250 -514
rect 278 -542 316 -514
rect 344 -542 349 -514
rect -349 -580 349 -542
rect -349 -608 -344 -580
rect -316 -608 -278 -580
rect -250 -608 -212 -580
rect -184 -608 -146 -580
rect -118 -608 -80 -580
rect -52 -608 -14 -580
rect 14 -608 52 -580
rect 80 -608 118 -580
rect 146 -608 184 -580
rect 212 -608 250 -580
rect 278 -608 316 -580
rect 344 -608 349 -580
rect -349 -646 349 -608
rect -349 -674 -344 -646
rect -316 -674 -278 -646
rect -250 -674 -212 -646
rect -184 -674 -146 -646
rect -118 -674 -80 -646
rect -52 -674 -14 -646
rect 14 -674 52 -646
rect 80 -674 118 -646
rect 146 -674 184 -646
rect 212 -674 250 -646
rect 278 -674 316 -646
rect 344 -674 349 -646
rect -349 -712 349 -674
rect -349 -740 -344 -712
rect -316 -740 -278 -712
rect -250 -740 -212 -712
rect -184 -740 -146 -712
rect -118 -740 -80 -712
rect -52 -740 -14 -712
rect 14 -740 52 -712
rect 80 -740 118 -712
rect 146 -740 184 -712
rect 212 -740 250 -712
rect 278 -740 316 -712
rect 344 -740 349 -712
rect -349 -778 349 -740
rect -349 -806 -344 -778
rect -316 -806 -278 -778
rect -250 -806 -212 -778
rect -184 -806 -146 -778
rect -118 -806 -80 -778
rect -52 -806 -14 -778
rect 14 -806 52 -778
rect 80 -806 118 -778
rect 146 -806 184 -778
rect 212 -806 250 -778
rect 278 -806 316 -778
rect 344 -806 349 -778
rect -349 -844 349 -806
rect -349 -872 -344 -844
rect -316 -872 -278 -844
rect -250 -872 -212 -844
rect -184 -872 -146 -844
rect -118 -872 -80 -844
rect -52 -872 -14 -844
rect 14 -872 52 -844
rect 80 -872 118 -844
rect 146 -872 184 -844
rect 212 -872 250 -844
rect 278 -872 316 -844
rect 344 -872 349 -844
rect -349 -910 349 -872
rect -349 -938 -344 -910
rect -316 -938 -278 -910
rect -250 -938 -212 -910
rect -184 -938 -146 -910
rect -118 -938 -80 -910
rect -52 -938 -14 -910
rect 14 -938 52 -910
rect 80 -938 118 -910
rect 146 -938 184 -910
rect 212 -938 250 -910
rect 278 -938 316 -910
rect 344 -938 349 -910
rect -349 -976 349 -938
rect -349 -1004 -344 -976
rect -316 -1004 -278 -976
rect -250 -1004 -212 -976
rect -184 -1004 -146 -976
rect -118 -1004 -80 -976
rect -52 -1004 -14 -976
rect 14 -1004 52 -976
rect 80 -1004 118 -976
rect 146 -1004 184 -976
rect 212 -1004 250 -976
rect 278 -1004 316 -976
rect 344 -1004 349 -976
rect -349 -1042 349 -1004
rect -349 -1070 -344 -1042
rect -316 -1070 -278 -1042
rect -250 -1070 -212 -1042
rect -184 -1070 -146 -1042
rect -118 -1070 -80 -1042
rect -52 -1070 -14 -1042
rect 14 -1070 52 -1042
rect 80 -1070 118 -1042
rect 146 -1070 184 -1042
rect 212 -1070 250 -1042
rect 278 -1070 316 -1042
rect 344 -1070 349 -1042
rect -349 -1108 349 -1070
rect -349 -1136 -344 -1108
rect -316 -1136 -278 -1108
rect -250 -1136 -212 -1108
rect -184 -1136 -146 -1108
rect -118 -1136 -80 -1108
rect -52 -1136 -14 -1108
rect 14 -1136 52 -1108
rect 80 -1136 118 -1108
rect 146 -1136 184 -1108
rect 212 -1136 250 -1108
rect 278 -1136 316 -1108
rect 344 -1136 349 -1108
rect -349 -1174 349 -1136
rect -349 -1202 -344 -1174
rect -316 -1202 -278 -1174
rect -250 -1202 -212 -1174
rect -184 -1202 -146 -1174
rect -118 -1202 -80 -1174
rect -52 -1202 -14 -1174
rect 14 -1202 52 -1174
rect 80 -1202 118 -1174
rect 146 -1202 184 -1174
rect 212 -1202 250 -1174
rect 278 -1202 316 -1174
rect 344 -1202 349 -1174
rect -349 -1240 349 -1202
rect -349 -1268 -344 -1240
rect -316 -1268 -278 -1240
rect -250 -1268 -212 -1240
rect -184 -1268 -146 -1240
rect -118 -1268 -80 -1240
rect -52 -1268 -14 -1240
rect 14 -1268 52 -1240
rect 80 -1268 118 -1240
rect 146 -1268 184 -1240
rect 212 -1268 250 -1240
rect 278 -1268 316 -1240
rect 344 -1268 349 -1240
rect -349 -1306 349 -1268
rect -349 -1334 -344 -1306
rect -316 -1334 -278 -1306
rect -250 -1334 -212 -1306
rect -184 -1334 -146 -1306
rect -118 -1334 -80 -1306
rect -52 -1334 -14 -1306
rect 14 -1334 52 -1306
rect 80 -1334 118 -1306
rect 146 -1334 184 -1306
rect 212 -1334 250 -1306
rect 278 -1334 316 -1306
rect 344 -1334 349 -1306
rect -349 -1372 349 -1334
rect -349 -1400 -344 -1372
rect -316 -1400 -278 -1372
rect -250 -1400 -212 -1372
rect -184 -1400 -146 -1372
rect -118 -1400 -80 -1372
rect -52 -1400 -14 -1372
rect 14 -1400 52 -1372
rect 80 -1400 118 -1372
rect 146 -1400 184 -1372
rect 212 -1400 250 -1372
rect 278 -1400 316 -1372
rect 344 -1400 349 -1372
rect -349 -1438 349 -1400
rect -349 -1466 -344 -1438
rect -316 -1466 -278 -1438
rect -250 -1466 -212 -1438
rect -184 -1466 -146 -1438
rect -118 -1466 -80 -1438
rect -52 -1466 -14 -1438
rect 14 -1466 52 -1438
rect 80 -1466 118 -1438
rect 146 -1466 184 -1438
rect 212 -1466 250 -1438
rect 278 -1466 316 -1438
rect 344 -1466 349 -1438
rect -349 -1504 349 -1466
rect -349 -1532 -344 -1504
rect -316 -1532 -278 -1504
rect -250 -1532 -212 -1504
rect -184 -1532 -146 -1504
rect -118 -1532 -80 -1504
rect -52 -1532 -14 -1504
rect 14 -1532 52 -1504
rect 80 -1532 118 -1504
rect 146 -1532 184 -1504
rect 212 -1532 250 -1504
rect 278 -1532 316 -1504
rect 344 -1532 349 -1504
rect -349 -1570 349 -1532
rect -349 -1598 -344 -1570
rect -316 -1598 -278 -1570
rect -250 -1598 -212 -1570
rect -184 -1598 -146 -1570
rect -118 -1598 -80 -1570
rect -52 -1598 -14 -1570
rect 14 -1598 52 -1570
rect 80 -1598 118 -1570
rect 146 -1598 184 -1570
rect 212 -1598 250 -1570
rect 278 -1598 316 -1570
rect 344 -1598 349 -1570
rect -349 -1636 349 -1598
rect -349 -1664 -344 -1636
rect -316 -1664 -278 -1636
rect -250 -1664 -212 -1636
rect -184 -1664 -146 -1636
rect -118 -1664 -80 -1636
rect -52 -1664 -14 -1636
rect 14 -1664 52 -1636
rect 80 -1664 118 -1636
rect 146 -1664 184 -1636
rect 212 -1664 250 -1636
rect 278 -1664 316 -1636
rect 344 -1664 349 -1636
rect -349 -1702 349 -1664
rect -349 -1730 -344 -1702
rect -316 -1730 -278 -1702
rect -250 -1730 -212 -1702
rect -184 -1730 -146 -1702
rect -118 -1730 -80 -1702
rect -52 -1730 -14 -1702
rect 14 -1730 52 -1702
rect 80 -1730 118 -1702
rect 146 -1730 184 -1702
rect 212 -1730 250 -1702
rect 278 -1730 316 -1702
rect 344 -1730 349 -1702
rect -349 -1768 349 -1730
rect -349 -1796 -344 -1768
rect -316 -1796 -278 -1768
rect -250 -1796 -212 -1768
rect -184 -1796 -146 -1768
rect -118 -1796 -80 -1768
rect -52 -1796 -14 -1768
rect 14 -1796 52 -1768
rect 80 -1796 118 -1768
rect 146 -1796 184 -1768
rect 212 -1796 250 -1768
rect 278 -1796 316 -1768
rect 344 -1796 349 -1768
rect -349 -1834 349 -1796
rect -349 -1862 -344 -1834
rect -316 -1862 -278 -1834
rect -250 -1862 -212 -1834
rect -184 -1862 -146 -1834
rect -118 -1862 -80 -1834
rect -52 -1862 -14 -1834
rect 14 -1862 52 -1834
rect 80 -1862 118 -1834
rect 146 -1862 184 -1834
rect 212 -1862 250 -1834
rect 278 -1862 316 -1834
rect 344 -1862 349 -1834
rect -349 -1900 349 -1862
rect -349 -1928 -344 -1900
rect -316 -1928 -278 -1900
rect -250 -1928 -212 -1900
rect -184 -1928 -146 -1900
rect -118 -1928 -80 -1900
rect -52 -1928 -14 -1900
rect 14 -1928 52 -1900
rect 80 -1928 118 -1900
rect 146 -1928 184 -1900
rect 212 -1928 250 -1900
rect 278 -1928 316 -1900
rect 344 -1928 349 -1900
rect -349 -1966 349 -1928
rect -349 -1994 -344 -1966
rect -316 -1994 -278 -1966
rect -250 -1994 -212 -1966
rect -184 -1994 -146 -1966
rect -118 -1994 -80 -1966
rect -52 -1994 -14 -1966
rect 14 -1994 52 -1966
rect 80 -1994 118 -1966
rect 146 -1994 184 -1966
rect 212 -1994 250 -1966
rect 278 -1994 316 -1966
rect 344 -1994 349 -1966
rect -349 -2032 349 -1994
rect -349 -2060 -344 -2032
rect -316 -2060 -278 -2032
rect -250 -2060 -212 -2032
rect -184 -2060 -146 -2032
rect -118 -2060 -80 -2032
rect -52 -2060 -14 -2032
rect 14 -2060 52 -2032
rect 80 -2060 118 -2032
rect 146 -2060 184 -2032
rect 212 -2060 250 -2032
rect 278 -2060 316 -2032
rect 344 -2060 349 -2032
rect -349 -2098 349 -2060
rect -349 -2126 -344 -2098
rect -316 -2126 -278 -2098
rect -250 -2126 -212 -2098
rect -184 -2126 -146 -2098
rect -118 -2126 -80 -2098
rect -52 -2126 -14 -2098
rect 14 -2126 52 -2098
rect 80 -2126 118 -2098
rect 146 -2126 184 -2098
rect 212 -2126 250 -2098
rect 278 -2126 316 -2098
rect 344 -2126 349 -2098
rect -349 -2164 349 -2126
rect -349 -2192 -344 -2164
rect -316 -2192 -278 -2164
rect -250 -2192 -212 -2164
rect -184 -2192 -146 -2164
rect -118 -2192 -80 -2164
rect -52 -2192 -14 -2164
rect 14 -2192 52 -2164
rect 80 -2192 118 -2164
rect 146 -2192 184 -2164
rect 212 -2192 250 -2164
rect 278 -2192 316 -2164
rect 344 -2192 349 -2164
rect -349 -2230 349 -2192
rect -349 -2258 -344 -2230
rect -316 -2258 -278 -2230
rect -250 -2258 -212 -2230
rect -184 -2258 -146 -2230
rect -118 -2258 -80 -2230
rect -52 -2258 -14 -2230
rect 14 -2258 52 -2230
rect 80 -2258 118 -2230
rect 146 -2258 184 -2230
rect 212 -2258 250 -2230
rect 278 -2258 316 -2230
rect 344 -2258 349 -2230
rect -349 -2296 349 -2258
rect -349 -2324 -344 -2296
rect -316 -2324 -278 -2296
rect -250 -2324 -212 -2296
rect -184 -2324 -146 -2296
rect -118 -2324 -80 -2296
rect -52 -2324 -14 -2296
rect 14 -2324 52 -2296
rect 80 -2324 118 -2296
rect 146 -2324 184 -2296
rect 212 -2324 250 -2296
rect 278 -2324 316 -2296
rect 344 -2324 349 -2296
rect -349 -2362 349 -2324
rect -349 -2390 -344 -2362
rect -316 -2390 -278 -2362
rect -250 -2390 -212 -2362
rect -184 -2390 -146 -2362
rect -118 -2390 -80 -2362
rect -52 -2390 -14 -2362
rect 14 -2390 52 -2362
rect 80 -2390 118 -2362
rect 146 -2390 184 -2362
rect 212 -2390 250 -2362
rect 278 -2390 316 -2362
rect 344 -2390 349 -2362
rect -349 -2428 349 -2390
rect -349 -2456 -344 -2428
rect -316 -2456 -278 -2428
rect -250 -2456 -212 -2428
rect -184 -2456 -146 -2428
rect -118 -2456 -80 -2428
rect -52 -2456 -14 -2428
rect 14 -2456 52 -2428
rect 80 -2456 118 -2428
rect 146 -2456 184 -2428
rect 212 -2456 250 -2428
rect 278 -2456 316 -2428
rect 344 -2456 349 -2428
rect -349 -2494 349 -2456
rect -349 -2522 -344 -2494
rect -316 -2522 -278 -2494
rect -250 -2522 -212 -2494
rect -184 -2522 -146 -2494
rect -118 -2522 -80 -2494
rect -52 -2522 -14 -2494
rect 14 -2522 52 -2494
rect 80 -2522 118 -2494
rect 146 -2522 184 -2494
rect 212 -2522 250 -2494
rect 278 -2522 316 -2494
rect 344 -2522 349 -2494
rect -349 -2560 349 -2522
rect -349 -2588 -344 -2560
rect -316 -2588 -278 -2560
rect -250 -2588 -212 -2560
rect -184 -2588 -146 -2560
rect -118 -2588 -80 -2560
rect -52 -2588 -14 -2560
rect 14 -2588 52 -2560
rect 80 -2588 118 -2560
rect 146 -2588 184 -2560
rect 212 -2588 250 -2560
rect 278 -2588 316 -2560
rect 344 -2588 349 -2560
rect -349 -2626 349 -2588
rect -349 -2654 -344 -2626
rect -316 -2654 -278 -2626
rect -250 -2654 -212 -2626
rect -184 -2654 -146 -2626
rect -118 -2654 -80 -2626
rect -52 -2654 -14 -2626
rect 14 -2654 52 -2626
rect 80 -2654 118 -2626
rect 146 -2654 184 -2626
rect 212 -2654 250 -2626
rect 278 -2654 316 -2626
rect 344 -2654 349 -2626
rect -349 -2692 349 -2654
rect -349 -2720 -344 -2692
rect -316 -2720 -278 -2692
rect -250 -2720 -212 -2692
rect -184 -2720 -146 -2692
rect -118 -2720 -80 -2692
rect -52 -2720 -14 -2692
rect 14 -2720 52 -2692
rect 80 -2720 118 -2692
rect 146 -2720 184 -2692
rect 212 -2720 250 -2692
rect 278 -2720 316 -2692
rect 344 -2720 349 -2692
rect -349 -2758 349 -2720
rect -349 -2786 -344 -2758
rect -316 -2786 -278 -2758
rect -250 -2786 -212 -2758
rect -184 -2786 -146 -2758
rect -118 -2786 -80 -2758
rect -52 -2786 -14 -2758
rect 14 -2786 52 -2758
rect 80 -2786 118 -2758
rect 146 -2786 184 -2758
rect 212 -2786 250 -2758
rect 278 -2786 316 -2758
rect 344 -2786 349 -2758
rect -349 -2824 349 -2786
rect -349 -2852 -344 -2824
rect -316 -2852 -278 -2824
rect -250 -2852 -212 -2824
rect -184 -2852 -146 -2824
rect -118 -2852 -80 -2824
rect -52 -2852 -14 -2824
rect 14 -2852 52 -2824
rect 80 -2852 118 -2824
rect 146 -2852 184 -2824
rect 212 -2852 250 -2824
rect 278 -2852 316 -2824
rect 344 -2852 349 -2824
rect -349 -2890 349 -2852
rect -349 -2918 -344 -2890
rect -316 -2918 -278 -2890
rect -250 -2918 -212 -2890
rect -184 -2918 -146 -2890
rect -118 -2918 -80 -2890
rect -52 -2918 -14 -2890
rect 14 -2918 52 -2890
rect 80 -2918 118 -2890
rect 146 -2918 184 -2890
rect 212 -2918 250 -2890
rect 278 -2918 316 -2890
rect 344 -2918 349 -2890
rect -349 -2956 349 -2918
rect -349 -2984 -344 -2956
rect -316 -2984 -278 -2956
rect -250 -2984 -212 -2956
rect -184 -2984 -146 -2956
rect -118 -2984 -80 -2956
rect -52 -2984 -14 -2956
rect 14 -2984 52 -2956
rect 80 -2984 118 -2956
rect 146 -2984 184 -2956
rect 212 -2984 250 -2956
rect 278 -2984 316 -2956
rect 344 -2984 349 -2956
rect -349 -3022 349 -2984
rect -349 -3050 -344 -3022
rect -316 -3050 -278 -3022
rect -250 -3050 -212 -3022
rect -184 -3050 -146 -3022
rect -118 -3050 -80 -3022
rect -52 -3050 -14 -3022
rect 14 -3050 52 -3022
rect 80 -3050 118 -3022
rect 146 -3050 184 -3022
rect 212 -3050 250 -3022
rect 278 -3050 316 -3022
rect 344 -3050 349 -3022
rect -349 -3088 349 -3050
rect -349 -3116 -344 -3088
rect -316 -3116 -278 -3088
rect -250 -3116 -212 -3088
rect -184 -3116 -146 -3088
rect -118 -3116 -80 -3088
rect -52 -3116 -14 -3088
rect 14 -3116 52 -3088
rect 80 -3116 118 -3088
rect 146 -3116 184 -3088
rect 212 -3116 250 -3088
rect 278 -3116 316 -3088
rect 344 -3116 349 -3088
rect -349 -3154 349 -3116
rect -349 -3182 -344 -3154
rect -316 -3182 -278 -3154
rect -250 -3182 -212 -3154
rect -184 -3182 -146 -3154
rect -118 -3182 -80 -3154
rect -52 -3182 -14 -3154
rect 14 -3182 52 -3154
rect 80 -3182 118 -3154
rect 146 -3182 184 -3154
rect 212 -3182 250 -3154
rect 278 -3182 316 -3154
rect 344 -3182 349 -3154
rect -349 -3220 349 -3182
rect -349 -3248 -344 -3220
rect -316 -3248 -278 -3220
rect -250 -3248 -212 -3220
rect -184 -3248 -146 -3220
rect -118 -3248 -80 -3220
rect -52 -3248 -14 -3220
rect 14 -3248 52 -3220
rect 80 -3248 118 -3220
rect 146 -3248 184 -3220
rect 212 -3248 250 -3220
rect 278 -3248 316 -3220
rect 344 -3248 349 -3220
rect -349 -3286 349 -3248
rect -349 -3314 -344 -3286
rect -316 -3314 -278 -3286
rect -250 -3314 -212 -3286
rect -184 -3314 -146 -3286
rect -118 -3314 -80 -3286
rect -52 -3314 -14 -3286
rect 14 -3314 52 -3286
rect 80 -3314 118 -3286
rect 146 -3314 184 -3286
rect 212 -3314 250 -3286
rect 278 -3314 316 -3286
rect 344 -3314 349 -3286
rect -349 -3352 349 -3314
rect -349 -3380 -344 -3352
rect -316 -3380 -278 -3352
rect -250 -3380 -212 -3352
rect -184 -3380 -146 -3352
rect -118 -3380 -80 -3352
rect -52 -3380 -14 -3352
rect 14 -3380 52 -3352
rect 80 -3380 118 -3352
rect 146 -3380 184 -3352
rect 212 -3380 250 -3352
rect 278 -3380 316 -3352
rect 344 -3380 349 -3352
rect -349 -3385 349 -3380
<< via3 >>
rect -344 3352 -316 3380
rect -278 3352 -250 3380
rect -212 3352 -184 3380
rect -146 3352 -118 3380
rect -80 3352 -52 3380
rect -14 3352 14 3380
rect 52 3352 80 3380
rect 118 3352 146 3380
rect 184 3352 212 3380
rect 250 3352 278 3380
rect 316 3352 344 3380
rect -344 3286 -316 3314
rect -278 3286 -250 3314
rect -212 3286 -184 3314
rect -146 3286 -118 3314
rect -80 3286 -52 3314
rect -14 3286 14 3314
rect 52 3286 80 3314
rect 118 3286 146 3314
rect 184 3286 212 3314
rect 250 3286 278 3314
rect 316 3286 344 3314
rect -344 3220 -316 3248
rect -278 3220 -250 3248
rect -212 3220 -184 3248
rect -146 3220 -118 3248
rect -80 3220 -52 3248
rect -14 3220 14 3248
rect 52 3220 80 3248
rect 118 3220 146 3248
rect 184 3220 212 3248
rect 250 3220 278 3248
rect 316 3220 344 3248
rect -344 3154 -316 3182
rect -278 3154 -250 3182
rect -212 3154 -184 3182
rect -146 3154 -118 3182
rect -80 3154 -52 3182
rect -14 3154 14 3182
rect 52 3154 80 3182
rect 118 3154 146 3182
rect 184 3154 212 3182
rect 250 3154 278 3182
rect 316 3154 344 3182
rect -344 3088 -316 3116
rect -278 3088 -250 3116
rect -212 3088 -184 3116
rect -146 3088 -118 3116
rect -80 3088 -52 3116
rect -14 3088 14 3116
rect 52 3088 80 3116
rect 118 3088 146 3116
rect 184 3088 212 3116
rect 250 3088 278 3116
rect 316 3088 344 3116
rect -344 3022 -316 3050
rect -278 3022 -250 3050
rect -212 3022 -184 3050
rect -146 3022 -118 3050
rect -80 3022 -52 3050
rect -14 3022 14 3050
rect 52 3022 80 3050
rect 118 3022 146 3050
rect 184 3022 212 3050
rect 250 3022 278 3050
rect 316 3022 344 3050
rect -344 2956 -316 2984
rect -278 2956 -250 2984
rect -212 2956 -184 2984
rect -146 2956 -118 2984
rect -80 2956 -52 2984
rect -14 2956 14 2984
rect 52 2956 80 2984
rect 118 2956 146 2984
rect 184 2956 212 2984
rect 250 2956 278 2984
rect 316 2956 344 2984
rect -344 2890 -316 2918
rect -278 2890 -250 2918
rect -212 2890 -184 2918
rect -146 2890 -118 2918
rect -80 2890 -52 2918
rect -14 2890 14 2918
rect 52 2890 80 2918
rect 118 2890 146 2918
rect 184 2890 212 2918
rect 250 2890 278 2918
rect 316 2890 344 2918
rect -344 2824 -316 2852
rect -278 2824 -250 2852
rect -212 2824 -184 2852
rect -146 2824 -118 2852
rect -80 2824 -52 2852
rect -14 2824 14 2852
rect 52 2824 80 2852
rect 118 2824 146 2852
rect 184 2824 212 2852
rect 250 2824 278 2852
rect 316 2824 344 2852
rect -344 2758 -316 2786
rect -278 2758 -250 2786
rect -212 2758 -184 2786
rect -146 2758 -118 2786
rect -80 2758 -52 2786
rect -14 2758 14 2786
rect 52 2758 80 2786
rect 118 2758 146 2786
rect 184 2758 212 2786
rect 250 2758 278 2786
rect 316 2758 344 2786
rect -344 2692 -316 2720
rect -278 2692 -250 2720
rect -212 2692 -184 2720
rect -146 2692 -118 2720
rect -80 2692 -52 2720
rect -14 2692 14 2720
rect 52 2692 80 2720
rect 118 2692 146 2720
rect 184 2692 212 2720
rect 250 2692 278 2720
rect 316 2692 344 2720
rect -344 2626 -316 2654
rect -278 2626 -250 2654
rect -212 2626 -184 2654
rect -146 2626 -118 2654
rect -80 2626 -52 2654
rect -14 2626 14 2654
rect 52 2626 80 2654
rect 118 2626 146 2654
rect 184 2626 212 2654
rect 250 2626 278 2654
rect 316 2626 344 2654
rect -344 2560 -316 2588
rect -278 2560 -250 2588
rect -212 2560 -184 2588
rect -146 2560 -118 2588
rect -80 2560 -52 2588
rect -14 2560 14 2588
rect 52 2560 80 2588
rect 118 2560 146 2588
rect 184 2560 212 2588
rect 250 2560 278 2588
rect 316 2560 344 2588
rect -344 2494 -316 2522
rect -278 2494 -250 2522
rect -212 2494 -184 2522
rect -146 2494 -118 2522
rect -80 2494 -52 2522
rect -14 2494 14 2522
rect 52 2494 80 2522
rect 118 2494 146 2522
rect 184 2494 212 2522
rect 250 2494 278 2522
rect 316 2494 344 2522
rect -344 2428 -316 2456
rect -278 2428 -250 2456
rect -212 2428 -184 2456
rect -146 2428 -118 2456
rect -80 2428 -52 2456
rect -14 2428 14 2456
rect 52 2428 80 2456
rect 118 2428 146 2456
rect 184 2428 212 2456
rect 250 2428 278 2456
rect 316 2428 344 2456
rect -344 2362 -316 2390
rect -278 2362 -250 2390
rect -212 2362 -184 2390
rect -146 2362 -118 2390
rect -80 2362 -52 2390
rect -14 2362 14 2390
rect 52 2362 80 2390
rect 118 2362 146 2390
rect 184 2362 212 2390
rect 250 2362 278 2390
rect 316 2362 344 2390
rect -344 2296 -316 2324
rect -278 2296 -250 2324
rect -212 2296 -184 2324
rect -146 2296 -118 2324
rect -80 2296 -52 2324
rect -14 2296 14 2324
rect 52 2296 80 2324
rect 118 2296 146 2324
rect 184 2296 212 2324
rect 250 2296 278 2324
rect 316 2296 344 2324
rect -344 2230 -316 2258
rect -278 2230 -250 2258
rect -212 2230 -184 2258
rect -146 2230 -118 2258
rect -80 2230 -52 2258
rect -14 2230 14 2258
rect 52 2230 80 2258
rect 118 2230 146 2258
rect 184 2230 212 2258
rect 250 2230 278 2258
rect 316 2230 344 2258
rect -344 2164 -316 2192
rect -278 2164 -250 2192
rect -212 2164 -184 2192
rect -146 2164 -118 2192
rect -80 2164 -52 2192
rect -14 2164 14 2192
rect 52 2164 80 2192
rect 118 2164 146 2192
rect 184 2164 212 2192
rect 250 2164 278 2192
rect 316 2164 344 2192
rect -344 2098 -316 2126
rect -278 2098 -250 2126
rect -212 2098 -184 2126
rect -146 2098 -118 2126
rect -80 2098 -52 2126
rect -14 2098 14 2126
rect 52 2098 80 2126
rect 118 2098 146 2126
rect 184 2098 212 2126
rect 250 2098 278 2126
rect 316 2098 344 2126
rect -344 2032 -316 2060
rect -278 2032 -250 2060
rect -212 2032 -184 2060
rect -146 2032 -118 2060
rect -80 2032 -52 2060
rect -14 2032 14 2060
rect 52 2032 80 2060
rect 118 2032 146 2060
rect 184 2032 212 2060
rect 250 2032 278 2060
rect 316 2032 344 2060
rect -344 1966 -316 1994
rect -278 1966 -250 1994
rect -212 1966 -184 1994
rect -146 1966 -118 1994
rect -80 1966 -52 1994
rect -14 1966 14 1994
rect 52 1966 80 1994
rect 118 1966 146 1994
rect 184 1966 212 1994
rect 250 1966 278 1994
rect 316 1966 344 1994
rect -344 1900 -316 1928
rect -278 1900 -250 1928
rect -212 1900 -184 1928
rect -146 1900 -118 1928
rect -80 1900 -52 1928
rect -14 1900 14 1928
rect 52 1900 80 1928
rect 118 1900 146 1928
rect 184 1900 212 1928
rect 250 1900 278 1928
rect 316 1900 344 1928
rect -344 1834 -316 1862
rect -278 1834 -250 1862
rect -212 1834 -184 1862
rect -146 1834 -118 1862
rect -80 1834 -52 1862
rect -14 1834 14 1862
rect 52 1834 80 1862
rect 118 1834 146 1862
rect 184 1834 212 1862
rect 250 1834 278 1862
rect 316 1834 344 1862
rect -344 1768 -316 1796
rect -278 1768 -250 1796
rect -212 1768 -184 1796
rect -146 1768 -118 1796
rect -80 1768 -52 1796
rect -14 1768 14 1796
rect 52 1768 80 1796
rect 118 1768 146 1796
rect 184 1768 212 1796
rect 250 1768 278 1796
rect 316 1768 344 1796
rect -344 1702 -316 1730
rect -278 1702 -250 1730
rect -212 1702 -184 1730
rect -146 1702 -118 1730
rect -80 1702 -52 1730
rect -14 1702 14 1730
rect 52 1702 80 1730
rect 118 1702 146 1730
rect 184 1702 212 1730
rect 250 1702 278 1730
rect 316 1702 344 1730
rect -344 1636 -316 1664
rect -278 1636 -250 1664
rect -212 1636 -184 1664
rect -146 1636 -118 1664
rect -80 1636 -52 1664
rect -14 1636 14 1664
rect 52 1636 80 1664
rect 118 1636 146 1664
rect 184 1636 212 1664
rect 250 1636 278 1664
rect 316 1636 344 1664
rect -344 1570 -316 1598
rect -278 1570 -250 1598
rect -212 1570 -184 1598
rect -146 1570 -118 1598
rect -80 1570 -52 1598
rect -14 1570 14 1598
rect 52 1570 80 1598
rect 118 1570 146 1598
rect 184 1570 212 1598
rect 250 1570 278 1598
rect 316 1570 344 1598
rect -344 1504 -316 1532
rect -278 1504 -250 1532
rect -212 1504 -184 1532
rect -146 1504 -118 1532
rect -80 1504 -52 1532
rect -14 1504 14 1532
rect 52 1504 80 1532
rect 118 1504 146 1532
rect 184 1504 212 1532
rect 250 1504 278 1532
rect 316 1504 344 1532
rect -344 1438 -316 1466
rect -278 1438 -250 1466
rect -212 1438 -184 1466
rect -146 1438 -118 1466
rect -80 1438 -52 1466
rect -14 1438 14 1466
rect 52 1438 80 1466
rect 118 1438 146 1466
rect 184 1438 212 1466
rect 250 1438 278 1466
rect 316 1438 344 1466
rect -344 1372 -316 1400
rect -278 1372 -250 1400
rect -212 1372 -184 1400
rect -146 1372 -118 1400
rect -80 1372 -52 1400
rect -14 1372 14 1400
rect 52 1372 80 1400
rect 118 1372 146 1400
rect 184 1372 212 1400
rect 250 1372 278 1400
rect 316 1372 344 1400
rect -344 1306 -316 1334
rect -278 1306 -250 1334
rect -212 1306 -184 1334
rect -146 1306 -118 1334
rect -80 1306 -52 1334
rect -14 1306 14 1334
rect 52 1306 80 1334
rect 118 1306 146 1334
rect 184 1306 212 1334
rect 250 1306 278 1334
rect 316 1306 344 1334
rect -344 1240 -316 1268
rect -278 1240 -250 1268
rect -212 1240 -184 1268
rect -146 1240 -118 1268
rect -80 1240 -52 1268
rect -14 1240 14 1268
rect 52 1240 80 1268
rect 118 1240 146 1268
rect 184 1240 212 1268
rect 250 1240 278 1268
rect 316 1240 344 1268
rect -344 1174 -316 1202
rect -278 1174 -250 1202
rect -212 1174 -184 1202
rect -146 1174 -118 1202
rect -80 1174 -52 1202
rect -14 1174 14 1202
rect 52 1174 80 1202
rect 118 1174 146 1202
rect 184 1174 212 1202
rect 250 1174 278 1202
rect 316 1174 344 1202
rect -344 1108 -316 1136
rect -278 1108 -250 1136
rect -212 1108 -184 1136
rect -146 1108 -118 1136
rect -80 1108 -52 1136
rect -14 1108 14 1136
rect 52 1108 80 1136
rect 118 1108 146 1136
rect 184 1108 212 1136
rect 250 1108 278 1136
rect 316 1108 344 1136
rect -344 1042 -316 1070
rect -278 1042 -250 1070
rect -212 1042 -184 1070
rect -146 1042 -118 1070
rect -80 1042 -52 1070
rect -14 1042 14 1070
rect 52 1042 80 1070
rect 118 1042 146 1070
rect 184 1042 212 1070
rect 250 1042 278 1070
rect 316 1042 344 1070
rect -344 976 -316 1004
rect -278 976 -250 1004
rect -212 976 -184 1004
rect -146 976 -118 1004
rect -80 976 -52 1004
rect -14 976 14 1004
rect 52 976 80 1004
rect 118 976 146 1004
rect 184 976 212 1004
rect 250 976 278 1004
rect 316 976 344 1004
rect -344 910 -316 938
rect -278 910 -250 938
rect -212 910 -184 938
rect -146 910 -118 938
rect -80 910 -52 938
rect -14 910 14 938
rect 52 910 80 938
rect 118 910 146 938
rect 184 910 212 938
rect 250 910 278 938
rect 316 910 344 938
rect -344 844 -316 872
rect -278 844 -250 872
rect -212 844 -184 872
rect -146 844 -118 872
rect -80 844 -52 872
rect -14 844 14 872
rect 52 844 80 872
rect 118 844 146 872
rect 184 844 212 872
rect 250 844 278 872
rect 316 844 344 872
rect -344 778 -316 806
rect -278 778 -250 806
rect -212 778 -184 806
rect -146 778 -118 806
rect -80 778 -52 806
rect -14 778 14 806
rect 52 778 80 806
rect 118 778 146 806
rect 184 778 212 806
rect 250 778 278 806
rect 316 778 344 806
rect -344 712 -316 740
rect -278 712 -250 740
rect -212 712 -184 740
rect -146 712 -118 740
rect -80 712 -52 740
rect -14 712 14 740
rect 52 712 80 740
rect 118 712 146 740
rect 184 712 212 740
rect 250 712 278 740
rect 316 712 344 740
rect -344 646 -316 674
rect -278 646 -250 674
rect -212 646 -184 674
rect -146 646 -118 674
rect -80 646 -52 674
rect -14 646 14 674
rect 52 646 80 674
rect 118 646 146 674
rect 184 646 212 674
rect 250 646 278 674
rect 316 646 344 674
rect -344 580 -316 608
rect -278 580 -250 608
rect -212 580 -184 608
rect -146 580 -118 608
rect -80 580 -52 608
rect -14 580 14 608
rect 52 580 80 608
rect 118 580 146 608
rect 184 580 212 608
rect 250 580 278 608
rect 316 580 344 608
rect -344 514 -316 542
rect -278 514 -250 542
rect -212 514 -184 542
rect -146 514 -118 542
rect -80 514 -52 542
rect -14 514 14 542
rect 52 514 80 542
rect 118 514 146 542
rect 184 514 212 542
rect 250 514 278 542
rect 316 514 344 542
rect -344 448 -316 476
rect -278 448 -250 476
rect -212 448 -184 476
rect -146 448 -118 476
rect -80 448 -52 476
rect -14 448 14 476
rect 52 448 80 476
rect 118 448 146 476
rect 184 448 212 476
rect 250 448 278 476
rect 316 448 344 476
rect -344 382 -316 410
rect -278 382 -250 410
rect -212 382 -184 410
rect -146 382 -118 410
rect -80 382 -52 410
rect -14 382 14 410
rect 52 382 80 410
rect 118 382 146 410
rect 184 382 212 410
rect 250 382 278 410
rect 316 382 344 410
rect -344 316 -316 344
rect -278 316 -250 344
rect -212 316 -184 344
rect -146 316 -118 344
rect -80 316 -52 344
rect -14 316 14 344
rect 52 316 80 344
rect 118 316 146 344
rect 184 316 212 344
rect 250 316 278 344
rect 316 316 344 344
rect -344 250 -316 278
rect -278 250 -250 278
rect -212 250 -184 278
rect -146 250 -118 278
rect -80 250 -52 278
rect -14 250 14 278
rect 52 250 80 278
rect 118 250 146 278
rect 184 250 212 278
rect 250 250 278 278
rect 316 250 344 278
rect -344 184 -316 212
rect -278 184 -250 212
rect -212 184 -184 212
rect -146 184 -118 212
rect -80 184 -52 212
rect -14 184 14 212
rect 52 184 80 212
rect 118 184 146 212
rect 184 184 212 212
rect 250 184 278 212
rect 316 184 344 212
rect -344 118 -316 146
rect -278 118 -250 146
rect -212 118 -184 146
rect -146 118 -118 146
rect -80 118 -52 146
rect -14 118 14 146
rect 52 118 80 146
rect 118 118 146 146
rect 184 118 212 146
rect 250 118 278 146
rect 316 118 344 146
rect -344 52 -316 80
rect -278 52 -250 80
rect -212 52 -184 80
rect -146 52 -118 80
rect -80 52 -52 80
rect -14 52 14 80
rect 52 52 80 80
rect 118 52 146 80
rect 184 52 212 80
rect 250 52 278 80
rect 316 52 344 80
rect -344 -14 -316 14
rect -278 -14 -250 14
rect -212 -14 -184 14
rect -146 -14 -118 14
rect -80 -14 -52 14
rect -14 -14 14 14
rect 52 -14 80 14
rect 118 -14 146 14
rect 184 -14 212 14
rect 250 -14 278 14
rect 316 -14 344 14
rect -344 -80 -316 -52
rect -278 -80 -250 -52
rect -212 -80 -184 -52
rect -146 -80 -118 -52
rect -80 -80 -52 -52
rect -14 -80 14 -52
rect 52 -80 80 -52
rect 118 -80 146 -52
rect 184 -80 212 -52
rect 250 -80 278 -52
rect 316 -80 344 -52
rect -344 -146 -316 -118
rect -278 -146 -250 -118
rect -212 -146 -184 -118
rect -146 -146 -118 -118
rect -80 -146 -52 -118
rect -14 -146 14 -118
rect 52 -146 80 -118
rect 118 -146 146 -118
rect 184 -146 212 -118
rect 250 -146 278 -118
rect 316 -146 344 -118
rect -344 -212 -316 -184
rect -278 -212 -250 -184
rect -212 -212 -184 -184
rect -146 -212 -118 -184
rect -80 -212 -52 -184
rect -14 -212 14 -184
rect 52 -212 80 -184
rect 118 -212 146 -184
rect 184 -212 212 -184
rect 250 -212 278 -184
rect 316 -212 344 -184
rect -344 -278 -316 -250
rect -278 -278 -250 -250
rect -212 -278 -184 -250
rect -146 -278 -118 -250
rect -80 -278 -52 -250
rect -14 -278 14 -250
rect 52 -278 80 -250
rect 118 -278 146 -250
rect 184 -278 212 -250
rect 250 -278 278 -250
rect 316 -278 344 -250
rect -344 -344 -316 -316
rect -278 -344 -250 -316
rect -212 -344 -184 -316
rect -146 -344 -118 -316
rect -80 -344 -52 -316
rect -14 -344 14 -316
rect 52 -344 80 -316
rect 118 -344 146 -316
rect 184 -344 212 -316
rect 250 -344 278 -316
rect 316 -344 344 -316
rect -344 -410 -316 -382
rect -278 -410 -250 -382
rect -212 -410 -184 -382
rect -146 -410 -118 -382
rect -80 -410 -52 -382
rect -14 -410 14 -382
rect 52 -410 80 -382
rect 118 -410 146 -382
rect 184 -410 212 -382
rect 250 -410 278 -382
rect 316 -410 344 -382
rect -344 -476 -316 -448
rect -278 -476 -250 -448
rect -212 -476 -184 -448
rect -146 -476 -118 -448
rect -80 -476 -52 -448
rect -14 -476 14 -448
rect 52 -476 80 -448
rect 118 -476 146 -448
rect 184 -476 212 -448
rect 250 -476 278 -448
rect 316 -476 344 -448
rect -344 -542 -316 -514
rect -278 -542 -250 -514
rect -212 -542 -184 -514
rect -146 -542 -118 -514
rect -80 -542 -52 -514
rect -14 -542 14 -514
rect 52 -542 80 -514
rect 118 -542 146 -514
rect 184 -542 212 -514
rect 250 -542 278 -514
rect 316 -542 344 -514
rect -344 -608 -316 -580
rect -278 -608 -250 -580
rect -212 -608 -184 -580
rect -146 -608 -118 -580
rect -80 -608 -52 -580
rect -14 -608 14 -580
rect 52 -608 80 -580
rect 118 -608 146 -580
rect 184 -608 212 -580
rect 250 -608 278 -580
rect 316 -608 344 -580
rect -344 -674 -316 -646
rect -278 -674 -250 -646
rect -212 -674 -184 -646
rect -146 -674 -118 -646
rect -80 -674 -52 -646
rect -14 -674 14 -646
rect 52 -674 80 -646
rect 118 -674 146 -646
rect 184 -674 212 -646
rect 250 -674 278 -646
rect 316 -674 344 -646
rect -344 -740 -316 -712
rect -278 -740 -250 -712
rect -212 -740 -184 -712
rect -146 -740 -118 -712
rect -80 -740 -52 -712
rect -14 -740 14 -712
rect 52 -740 80 -712
rect 118 -740 146 -712
rect 184 -740 212 -712
rect 250 -740 278 -712
rect 316 -740 344 -712
rect -344 -806 -316 -778
rect -278 -806 -250 -778
rect -212 -806 -184 -778
rect -146 -806 -118 -778
rect -80 -806 -52 -778
rect -14 -806 14 -778
rect 52 -806 80 -778
rect 118 -806 146 -778
rect 184 -806 212 -778
rect 250 -806 278 -778
rect 316 -806 344 -778
rect -344 -872 -316 -844
rect -278 -872 -250 -844
rect -212 -872 -184 -844
rect -146 -872 -118 -844
rect -80 -872 -52 -844
rect -14 -872 14 -844
rect 52 -872 80 -844
rect 118 -872 146 -844
rect 184 -872 212 -844
rect 250 -872 278 -844
rect 316 -872 344 -844
rect -344 -938 -316 -910
rect -278 -938 -250 -910
rect -212 -938 -184 -910
rect -146 -938 -118 -910
rect -80 -938 -52 -910
rect -14 -938 14 -910
rect 52 -938 80 -910
rect 118 -938 146 -910
rect 184 -938 212 -910
rect 250 -938 278 -910
rect 316 -938 344 -910
rect -344 -1004 -316 -976
rect -278 -1004 -250 -976
rect -212 -1004 -184 -976
rect -146 -1004 -118 -976
rect -80 -1004 -52 -976
rect -14 -1004 14 -976
rect 52 -1004 80 -976
rect 118 -1004 146 -976
rect 184 -1004 212 -976
rect 250 -1004 278 -976
rect 316 -1004 344 -976
rect -344 -1070 -316 -1042
rect -278 -1070 -250 -1042
rect -212 -1070 -184 -1042
rect -146 -1070 -118 -1042
rect -80 -1070 -52 -1042
rect -14 -1070 14 -1042
rect 52 -1070 80 -1042
rect 118 -1070 146 -1042
rect 184 -1070 212 -1042
rect 250 -1070 278 -1042
rect 316 -1070 344 -1042
rect -344 -1136 -316 -1108
rect -278 -1136 -250 -1108
rect -212 -1136 -184 -1108
rect -146 -1136 -118 -1108
rect -80 -1136 -52 -1108
rect -14 -1136 14 -1108
rect 52 -1136 80 -1108
rect 118 -1136 146 -1108
rect 184 -1136 212 -1108
rect 250 -1136 278 -1108
rect 316 -1136 344 -1108
rect -344 -1202 -316 -1174
rect -278 -1202 -250 -1174
rect -212 -1202 -184 -1174
rect -146 -1202 -118 -1174
rect -80 -1202 -52 -1174
rect -14 -1202 14 -1174
rect 52 -1202 80 -1174
rect 118 -1202 146 -1174
rect 184 -1202 212 -1174
rect 250 -1202 278 -1174
rect 316 -1202 344 -1174
rect -344 -1268 -316 -1240
rect -278 -1268 -250 -1240
rect -212 -1268 -184 -1240
rect -146 -1268 -118 -1240
rect -80 -1268 -52 -1240
rect -14 -1268 14 -1240
rect 52 -1268 80 -1240
rect 118 -1268 146 -1240
rect 184 -1268 212 -1240
rect 250 -1268 278 -1240
rect 316 -1268 344 -1240
rect -344 -1334 -316 -1306
rect -278 -1334 -250 -1306
rect -212 -1334 -184 -1306
rect -146 -1334 -118 -1306
rect -80 -1334 -52 -1306
rect -14 -1334 14 -1306
rect 52 -1334 80 -1306
rect 118 -1334 146 -1306
rect 184 -1334 212 -1306
rect 250 -1334 278 -1306
rect 316 -1334 344 -1306
rect -344 -1400 -316 -1372
rect -278 -1400 -250 -1372
rect -212 -1400 -184 -1372
rect -146 -1400 -118 -1372
rect -80 -1400 -52 -1372
rect -14 -1400 14 -1372
rect 52 -1400 80 -1372
rect 118 -1400 146 -1372
rect 184 -1400 212 -1372
rect 250 -1400 278 -1372
rect 316 -1400 344 -1372
rect -344 -1466 -316 -1438
rect -278 -1466 -250 -1438
rect -212 -1466 -184 -1438
rect -146 -1466 -118 -1438
rect -80 -1466 -52 -1438
rect -14 -1466 14 -1438
rect 52 -1466 80 -1438
rect 118 -1466 146 -1438
rect 184 -1466 212 -1438
rect 250 -1466 278 -1438
rect 316 -1466 344 -1438
rect -344 -1532 -316 -1504
rect -278 -1532 -250 -1504
rect -212 -1532 -184 -1504
rect -146 -1532 -118 -1504
rect -80 -1532 -52 -1504
rect -14 -1532 14 -1504
rect 52 -1532 80 -1504
rect 118 -1532 146 -1504
rect 184 -1532 212 -1504
rect 250 -1532 278 -1504
rect 316 -1532 344 -1504
rect -344 -1598 -316 -1570
rect -278 -1598 -250 -1570
rect -212 -1598 -184 -1570
rect -146 -1598 -118 -1570
rect -80 -1598 -52 -1570
rect -14 -1598 14 -1570
rect 52 -1598 80 -1570
rect 118 -1598 146 -1570
rect 184 -1598 212 -1570
rect 250 -1598 278 -1570
rect 316 -1598 344 -1570
rect -344 -1664 -316 -1636
rect -278 -1664 -250 -1636
rect -212 -1664 -184 -1636
rect -146 -1664 -118 -1636
rect -80 -1664 -52 -1636
rect -14 -1664 14 -1636
rect 52 -1664 80 -1636
rect 118 -1664 146 -1636
rect 184 -1664 212 -1636
rect 250 -1664 278 -1636
rect 316 -1664 344 -1636
rect -344 -1730 -316 -1702
rect -278 -1730 -250 -1702
rect -212 -1730 -184 -1702
rect -146 -1730 -118 -1702
rect -80 -1730 -52 -1702
rect -14 -1730 14 -1702
rect 52 -1730 80 -1702
rect 118 -1730 146 -1702
rect 184 -1730 212 -1702
rect 250 -1730 278 -1702
rect 316 -1730 344 -1702
rect -344 -1796 -316 -1768
rect -278 -1796 -250 -1768
rect -212 -1796 -184 -1768
rect -146 -1796 -118 -1768
rect -80 -1796 -52 -1768
rect -14 -1796 14 -1768
rect 52 -1796 80 -1768
rect 118 -1796 146 -1768
rect 184 -1796 212 -1768
rect 250 -1796 278 -1768
rect 316 -1796 344 -1768
rect -344 -1862 -316 -1834
rect -278 -1862 -250 -1834
rect -212 -1862 -184 -1834
rect -146 -1862 -118 -1834
rect -80 -1862 -52 -1834
rect -14 -1862 14 -1834
rect 52 -1862 80 -1834
rect 118 -1862 146 -1834
rect 184 -1862 212 -1834
rect 250 -1862 278 -1834
rect 316 -1862 344 -1834
rect -344 -1928 -316 -1900
rect -278 -1928 -250 -1900
rect -212 -1928 -184 -1900
rect -146 -1928 -118 -1900
rect -80 -1928 -52 -1900
rect -14 -1928 14 -1900
rect 52 -1928 80 -1900
rect 118 -1928 146 -1900
rect 184 -1928 212 -1900
rect 250 -1928 278 -1900
rect 316 -1928 344 -1900
rect -344 -1994 -316 -1966
rect -278 -1994 -250 -1966
rect -212 -1994 -184 -1966
rect -146 -1994 -118 -1966
rect -80 -1994 -52 -1966
rect -14 -1994 14 -1966
rect 52 -1994 80 -1966
rect 118 -1994 146 -1966
rect 184 -1994 212 -1966
rect 250 -1994 278 -1966
rect 316 -1994 344 -1966
rect -344 -2060 -316 -2032
rect -278 -2060 -250 -2032
rect -212 -2060 -184 -2032
rect -146 -2060 -118 -2032
rect -80 -2060 -52 -2032
rect -14 -2060 14 -2032
rect 52 -2060 80 -2032
rect 118 -2060 146 -2032
rect 184 -2060 212 -2032
rect 250 -2060 278 -2032
rect 316 -2060 344 -2032
rect -344 -2126 -316 -2098
rect -278 -2126 -250 -2098
rect -212 -2126 -184 -2098
rect -146 -2126 -118 -2098
rect -80 -2126 -52 -2098
rect -14 -2126 14 -2098
rect 52 -2126 80 -2098
rect 118 -2126 146 -2098
rect 184 -2126 212 -2098
rect 250 -2126 278 -2098
rect 316 -2126 344 -2098
rect -344 -2192 -316 -2164
rect -278 -2192 -250 -2164
rect -212 -2192 -184 -2164
rect -146 -2192 -118 -2164
rect -80 -2192 -52 -2164
rect -14 -2192 14 -2164
rect 52 -2192 80 -2164
rect 118 -2192 146 -2164
rect 184 -2192 212 -2164
rect 250 -2192 278 -2164
rect 316 -2192 344 -2164
rect -344 -2258 -316 -2230
rect -278 -2258 -250 -2230
rect -212 -2258 -184 -2230
rect -146 -2258 -118 -2230
rect -80 -2258 -52 -2230
rect -14 -2258 14 -2230
rect 52 -2258 80 -2230
rect 118 -2258 146 -2230
rect 184 -2258 212 -2230
rect 250 -2258 278 -2230
rect 316 -2258 344 -2230
rect -344 -2324 -316 -2296
rect -278 -2324 -250 -2296
rect -212 -2324 -184 -2296
rect -146 -2324 -118 -2296
rect -80 -2324 -52 -2296
rect -14 -2324 14 -2296
rect 52 -2324 80 -2296
rect 118 -2324 146 -2296
rect 184 -2324 212 -2296
rect 250 -2324 278 -2296
rect 316 -2324 344 -2296
rect -344 -2390 -316 -2362
rect -278 -2390 -250 -2362
rect -212 -2390 -184 -2362
rect -146 -2390 -118 -2362
rect -80 -2390 -52 -2362
rect -14 -2390 14 -2362
rect 52 -2390 80 -2362
rect 118 -2390 146 -2362
rect 184 -2390 212 -2362
rect 250 -2390 278 -2362
rect 316 -2390 344 -2362
rect -344 -2456 -316 -2428
rect -278 -2456 -250 -2428
rect -212 -2456 -184 -2428
rect -146 -2456 -118 -2428
rect -80 -2456 -52 -2428
rect -14 -2456 14 -2428
rect 52 -2456 80 -2428
rect 118 -2456 146 -2428
rect 184 -2456 212 -2428
rect 250 -2456 278 -2428
rect 316 -2456 344 -2428
rect -344 -2522 -316 -2494
rect -278 -2522 -250 -2494
rect -212 -2522 -184 -2494
rect -146 -2522 -118 -2494
rect -80 -2522 -52 -2494
rect -14 -2522 14 -2494
rect 52 -2522 80 -2494
rect 118 -2522 146 -2494
rect 184 -2522 212 -2494
rect 250 -2522 278 -2494
rect 316 -2522 344 -2494
rect -344 -2588 -316 -2560
rect -278 -2588 -250 -2560
rect -212 -2588 -184 -2560
rect -146 -2588 -118 -2560
rect -80 -2588 -52 -2560
rect -14 -2588 14 -2560
rect 52 -2588 80 -2560
rect 118 -2588 146 -2560
rect 184 -2588 212 -2560
rect 250 -2588 278 -2560
rect 316 -2588 344 -2560
rect -344 -2654 -316 -2626
rect -278 -2654 -250 -2626
rect -212 -2654 -184 -2626
rect -146 -2654 -118 -2626
rect -80 -2654 -52 -2626
rect -14 -2654 14 -2626
rect 52 -2654 80 -2626
rect 118 -2654 146 -2626
rect 184 -2654 212 -2626
rect 250 -2654 278 -2626
rect 316 -2654 344 -2626
rect -344 -2720 -316 -2692
rect -278 -2720 -250 -2692
rect -212 -2720 -184 -2692
rect -146 -2720 -118 -2692
rect -80 -2720 -52 -2692
rect -14 -2720 14 -2692
rect 52 -2720 80 -2692
rect 118 -2720 146 -2692
rect 184 -2720 212 -2692
rect 250 -2720 278 -2692
rect 316 -2720 344 -2692
rect -344 -2786 -316 -2758
rect -278 -2786 -250 -2758
rect -212 -2786 -184 -2758
rect -146 -2786 -118 -2758
rect -80 -2786 -52 -2758
rect -14 -2786 14 -2758
rect 52 -2786 80 -2758
rect 118 -2786 146 -2758
rect 184 -2786 212 -2758
rect 250 -2786 278 -2758
rect 316 -2786 344 -2758
rect -344 -2852 -316 -2824
rect -278 -2852 -250 -2824
rect -212 -2852 -184 -2824
rect -146 -2852 -118 -2824
rect -80 -2852 -52 -2824
rect -14 -2852 14 -2824
rect 52 -2852 80 -2824
rect 118 -2852 146 -2824
rect 184 -2852 212 -2824
rect 250 -2852 278 -2824
rect 316 -2852 344 -2824
rect -344 -2918 -316 -2890
rect -278 -2918 -250 -2890
rect -212 -2918 -184 -2890
rect -146 -2918 -118 -2890
rect -80 -2918 -52 -2890
rect -14 -2918 14 -2890
rect 52 -2918 80 -2890
rect 118 -2918 146 -2890
rect 184 -2918 212 -2890
rect 250 -2918 278 -2890
rect 316 -2918 344 -2890
rect -344 -2984 -316 -2956
rect -278 -2984 -250 -2956
rect -212 -2984 -184 -2956
rect -146 -2984 -118 -2956
rect -80 -2984 -52 -2956
rect -14 -2984 14 -2956
rect 52 -2984 80 -2956
rect 118 -2984 146 -2956
rect 184 -2984 212 -2956
rect 250 -2984 278 -2956
rect 316 -2984 344 -2956
rect -344 -3050 -316 -3022
rect -278 -3050 -250 -3022
rect -212 -3050 -184 -3022
rect -146 -3050 -118 -3022
rect -80 -3050 -52 -3022
rect -14 -3050 14 -3022
rect 52 -3050 80 -3022
rect 118 -3050 146 -3022
rect 184 -3050 212 -3022
rect 250 -3050 278 -3022
rect 316 -3050 344 -3022
rect -344 -3116 -316 -3088
rect -278 -3116 -250 -3088
rect -212 -3116 -184 -3088
rect -146 -3116 -118 -3088
rect -80 -3116 -52 -3088
rect -14 -3116 14 -3088
rect 52 -3116 80 -3088
rect 118 -3116 146 -3088
rect 184 -3116 212 -3088
rect 250 -3116 278 -3088
rect 316 -3116 344 -3088
rect -344 -3182 -316 -3154
rect -278 -3182 -250 -3154
rect -212 -3182 -184 -3154
rect -146 -3182 -118 -3154
rect -80 -3182 -52 -3154
rect -14 -3182 14 -3154
rect 52 -3182 80 -3154
rect 118 -3182 146 -3154
rect 184 -3182 212 -3154
rect 250 -3182 278 -3154
rect 316 -3182 344 -3154
rect -344 -3248 -316 -3220
rect -278 -3248 -250 -3220
rect -212 -3248 -184 -3220
rect -146 -3248 -118 -3220
rect -80 -3248 -52 -3220
rect -14 -3248 14 -3220
rect 52 -3248 80 -3220
rect 118 -3248 146 -3220
rect 184 -3248 212 -3220
rect 250 -3248 278 -3220
rect 316 -3248 344 -3220
rect -344 -3314 -316 -3286
rect -278 -3314 -250 -3286
rect -212 -3314 -184 -3286
rect -146 -3314 -118 -3286
rect -80 -3314 -52 -3286
rect -14 -3314 14 -3286
rect 52 -3314 80 -3286
rect 118 -3314 146 -3286
rect 184 -3314 212 -3286
rect 250 -3314 278 -3286
rect 316 -3314 344 -3286
rect -344 -3380 -316 -3352
rect -278 -3380 -250 -3352
rect -212 -3380 -184 -3352
rect -146 -3380 -118 -3352
rect -80 -3380 -52 -3352
rect -14 -3380 14 -3352
rect 52 -3380 80 -3352
rect 118 -3380 146 -3352
rect 184 -3380 212 -3352
rect 250 -3380 278 -3352
rect 316 -3380 344 -3352
<< metal4 >>
rect -349 3380 349 3385
rect -349 3352 -344 3380
rect -316 3352 -278 3380
rect -250 3352 -212 3380
rect -184 3352 -146 3380
rect -118 3352 -80 3380
rect -52 3352 -14 3380
rect 14 3352 52 3380
rect 80 3352 118 3380
rect 146 3352 184 3380
rect 212 3352 250 3380
rect 278 3352 316 3380
rect 344 3352 349 3380
rect -349 3314 349 3352
rect -349 3286 -344 3314
rect -316 3286 -278 3314
rect -250 3286 -212 3314
rect -184 3286 -146 3314
rect -118 3286 -80 3314
rect -52 3286 -14 3314
rect 14 3286 52 3314
rect 80 3286 118 3314
rect 146 3286 184 3314
rect 212 3286 250 3314
rect 278 3286 316 3314
rect 344 3286 349 3314
rect -349 3248 349 3286
rect -349 3220 -344 3248
rect -316 3220 -278 3248
rect -250 3220 -212 3248
rect -184 3220 -146 3248
rect -118 3220 -80 3248
rect -52 3220 -14 3248
rect 14 3220 52 3248
rect 80 3220 118 3248
rect 146 3220 184 3248
rect 212 3220 250 3248
rect 278 3220 316 3248
rect 344 3220 349 3248
rect -349 3182 349 3220
rect -349 3154 -344 3182
rect -316 3154 -278 3182
rect -250 3154 -212 3182
rect -184 3154 -146 3182
rect -118 3154 -80 3182
rect -52 3154 -14 3182
rect 14 3154 52 3182
rect 80 3154 118 3182
rect 146 3154 184 3182
rect 212 3154 250 3182
rect 278 3154 316 3182
rect 344 3154 349 3182
rect -349 3116 349 3154
rect -349 3088 -344 3116
rect -316 3088 -278 3116
rect -250 3088 -212 3116
rect -184 3088 -146 3116
rect -118 3088 -80 3116
rect -52 3088 -14 3116
rect 14 3088 52 3116
rect 80 3088 118 3116
rect 146 3088 184 3116
rect 212 3088 250 3116
rect 278 3088 316 3116
rect 344 3088 349 3116
rect -349 3050 349 3088
rect -349 3022 -344 3050
rect -316 3022 -278 3050
rect -250 3022 -212 3050
rect -184 3022 -146 3050
rect -118 3022 -80 3050
rect -52 3022 -14 3050
rect 14 3022 52 3050
rect 80 3022 118 3050
rect 146 3022 184 3050
rect 212 3022 250 3050
rect 278 3022 316 3050
rect 344 3022 349 3050
rect -349 2984 349 3022
rect -349 2956 -344 2984
rect -316 2956 -278 2984
rect -250 2956 -212 2984
rect -184 2956 -146 2984
rect -118 2956 -80 2984
rect -52 2956 -14 2984
rect 14 2956 52 2984
rect 80 2956 118 2984
rect 146 2956 184 2984
rect 212 2956 250 2984
rect 278 2956 316 2984
rect 344 2956 349 2984
rect -349 2918 349 2956
rect -349 2890 -344 2918
rect -316 2890 -278 2918
rect -250 2890 -212 2918
rect -184 2890 -146 2918
rect -118 2890 -80 2918
rect -52 2890 -14 2918
rect 14 2890 52 2918
rect 80 2890 118 2918
rect 146 2890 184 2918
rect 212 2890 250 2918
rect 278 2890 316 2918
rect 344 2890 349 2918
rect -349 2852 349 2890
rect -349 2824 -344 2852
rect -316 2824 -278 2852
rect -250 2824 -212 2852
rect -184 2824 -146 2852
rect -118 2824 -80 2852
rect -52 2824 -14 2852
rect 14 2824 52 2852
rect 80 2824 118 2852
rect 146 2824 184 2852
rect 212 2824 250 2852
rect 278 2824 316 2852
rect 344 2824 349 2852
rect -349 2786 349 2824
rect -349 2758 -344 2786
rect -316 2758 -278 2786
rect -250 2758 -212 2786
rect -184 2758 -146 2786
rect -118 2758 -80 2786
rect -52 2758 -14 2786
rect 14 2758 52 2786
rect 80 2758 118 2786
rect 146 2758 184 2786
rect 212 2758 250 2786
rect 278 2758 316 2786
rect 344 2758 349 2786
rect -349 2720 349 2758
rect -349 2692 -344 2720
rect -316 2692 -278 2720
rect -250 2692 -212 2720
rect -184 2692 -146 2720
rect -118 2692 -80 2720
rect -52 2692 -14 2720
rect 14 2692 52 2720
rect 80 2692 118 2720
rect 146 2692 184 2720
rect 212 2692 250 2720
rect 278 2692 316 2720
rect 344 2692 349 2720
rect -349 2654 349 2692
rect -349 2626 -344 2654
rect -316 2626 -278 2654
rect -250 2626 -212 2654
rect -184 2626 -146 2654
rect -118 2626 -80 2654
rect -52 2626 -14 2654
rect 14 2626 52 2654
rect 80 2626 118 2654
rect 146 2626 184 2654
rect 212 2626 250 2654
rect 278 2626 316 2654
rect 344 2626 349 2654
rect -349 2588 349 2626
rect -349 2560 -344 2588
rect -316 2560 -278 2588
rect -250 2560 -212 2588
rect -184 2560 -146 2588
rect -118 2560 -80 2588
rect -52 2560 -14 2588
rect 14 2560 52 2588
rect 80 2560 118 2588
rect 146 2560 184 2588
rect 212 2560 250 2588
rect 278 2560 316 2588
rect 344 2560 349 2588
rect -349 2522 349 2560
rect -349 2494 -344 2522
rect -316 2494 -278 2522
rect -250 2494 -212 2522
rect -184 2494 -146 2522
rect -118 2494 -80 2522
rect -52 2494 -14 2522
rect 14 2494 52 2522
rect 80 2494 118 2522
rect 146 2494 184 2522
rect 212 2494 250 2522
rect 278 2494 316 2522
rect 344 2494 349 2522
rect -349 2456 349 2494
rect -349 2428 -344 2456
rect -316 2428 -278 2456
rect -250 2428 -212 2456
rect -184 2428 -146 2456
rect -118 2428 -80 2456
rect -52 2428 -14 2456
rect 14 2428 52 2456
rect 80 2428 118 2456
rect 146 2428 184 2456
rect 212 2428 250 2456
rect 278 2428 316 2456
rect 344 2428 349 2456
rect -349 2390 349 2428
rect -349 2362 -344 2390
rect -316 2362 -278 2390
rect -250 2362 -212 2390
rect -184 2362 -146 2390
rect -118 2362 -80 2390
rect -52 2362 -14 2390
rect 14 2362 52 2390
rect 80 2362 118 2390
rect 146 2362 184 2390
rect 212 2362 250 2390
rect 278 2362 316 2390
rect 344 2362 349 2390
rect -349 2324 349 2362
rect -349 2296 -344 2324
rect -316 2296 -278 2324
rect -250 2296 -212 2324
rect -184 2296 -146 2324
rect -118 2296 -80 2324
rect -52 2296 -14 2324
rect 14 2296 52 2324
rect 80 2296 118 2324
rect 146 2296 184 2324
rect 212 2296 250 2324
rect 278 2296 316 2324
rect 344 2296 349 2324
rect -349 2258 349 2296
rect -349 2230 -344 2258
rect -316 2230 -278 2258
rect -250 2230 -212 2258
rect -184 2230 -146 2258
rect -118 2230 -80 2258
rect -52 2230 -14 2258
rect 14 2230 52 2258
rect 80 2230 118 2258
rect 146 2230 184 2258
rect 212 2230 250 2258
rect 278 2230 316 2258
rect 344 2230 349 2258
rect -349 2192 349 2230
rect -349 2164 -344 2192
rect -316 2164 -278 2192
rect -250 2164 -212 2192
rect -184 2164 -146 2192
rect -118 2164 -80 2192
rect -52 2164 -14 2192
rect 14 2164 52 2192
rect 80 2164 118 2192
rect 146 2164 184 2192
rect 212 2164 250 2192
rect 278 2164 316 2192
rect 344 2164 349 2192
rect -349 2126 349 2164
rect -349 2098 -344 2126
rect -316 2098 -278 2126
rect -250 2098 -212 2126
rect -184 2098 -146 2126
rect -118 2098 -80 2126
rect -52 2098 -14 2126
rect 14 2098 52 2126
rect 80 2098 118 2126
rect 146 2098 184 2126
rect 212 2098 250 2126
rect 278 2098 316 2126
rect 344 2098 349 2126
rect -349 2060 349 2098
rect -349 2032 -344 2060
rect -316 2032 -278 2060
rect -250 2032 -212 2060
rect -184 2032 -146 2060
rect -118 2032 -80 2060
rect -52 2032 -14 2060
rect 14 2032 52 2060
rect 80 2032 118 2060
rect 146 2032 184 2060
rect 212 2032 250 2060
rect 278 2032 316 2060
rect 344 2032 349 2060
rect -349 1994 349 2032
rect -349 1966 -344 1994
rect -316 1966 -278 1994
rect -250 1966 -212 1994
rect -184 1966 -146 1994
rect -118 1966 -80 1994
rect -52 1966 -14 1994
rect 14 1966 52 1994
rect 80 1966 118 1994
rect 146 1966 184 1994
rect 212 1966 250 1994
rect 278 1966 316 1994
rect 344 1966 349 1994
rect -349 1928 349 1966
rect -349 1900 -344 1928
rect -316 1900 -278 1928
rect -250 1900 -212 1928
rect -184 1900 -146 1928
rect -118 1900 -80 1928
rect -52 1900 -14 1928
rect 14 1900 52 1928
rect 80 1900 118 1928
rect 146 1900 184 1928
rect 212 1900 250 1928
rect 278 1900 316 1928
rect 344 1900 349 1928
rect -349 1862 349 1900
rect -349 1834 -344 1862
rect -316 1834 -278 1862
rect -250 1834 -212 1862
rect -184 1834 -146 1862
rect -118 1834 -80 1862
rect -52 1834 -14 1862
rect 14 1834 52 1862
rect 80 1834 118 1862
rect 146 1834 184 1862
rect 212 1834 250 1862
rect 278 1834 316 1862
rect 344 1834 349 1862
rect -349 1796 349 1834
rect -349 1768 -344 1796
rect -316 1768 -278 1796
rect -250 1768 -212 1796
rect -184 1768 -146 1796
rect -118 1768 -80 1796
rect -52 1768 -14 1796
rect 14 1768 52 1796
rect 80 1768 118 1796
rect 146 1768 184 1796
rect 212 1768 250 1796
rect 278 1768 316 1796
rect 344 1768 349 1796
rect -349 1730 349 1768
rect -349 1702 -344 1730
rect -316 1702 -278 1730
rect -250 1702 -212 1730
rect -184 1702 -146 1730
rect -118 1702 -80 1730
rect -52 1702 -14 1730
rect 14 1702 52 1730
rect 80 1702 118 1730
rect 146 1702 184 1730
rect 212 1702 250 1730
rect 278 1702 316 1730
rect 344 1702 349 1730
rect -349 1664 349 1702
rect -349 1636 -344 1664
rect -316 1636 -278 1664
rect -250 1636 -212 1664
rect -184 1636 -146 1664
rect -118 1636 -80 1664
rect -52 1636 -14 1664
rect 14 1636 52 1664
rect 80 1636 118 1664
rect 146 1636 184 1664
rect 212 1636 250 1664
rect 278 1636 316 1664
rect 344 1636 349 1664
rect -349 1598 349 1636
rect -349 1570 -344 1598
rect -316 1570 -278 1598
rect -250 1570 -212 1598
rect -184 1570 -146 1598
rect -118 1570 -80 1598
rect -52 1570 -14 1598
rect 14 1570 52 1598
rect 80 1570 118 1598
rect 146 1570 184 1598
rect 212 1570 250 1598
rect 278 1570 316 1598
rect 344 1570 349 1598
rect -349 1532 349 1570
rect -349 1504 -344 1532
rect -316 1504 -278 1532
rect -250 1504 -212 1532
rect -184 1504 -146 1532
rect -118 1504 -80 1532
rect -52 1504 -14 1532
rect 14 1504 52 1532
rect 80 1504 118 1532
rect 146 1504 184 1532
rect 212 1504 250 1532
rect 278 1504 316 1532
rect 344 1504 349 1532
rect -349 1466 349 1504
rect -349 1438 -344 1466
rect -316 1438 -278 1466
rect -250 1438 -212 1466
rect -184 1438 -146 1466
rect -118 1438 -80 1466
rect -52 1438 -14 1466
rect 14 1438 52 1466
rect 80 1438 118 1466
rect 146 1438 184 1466
rect 212 1438 250 1466
rect 278 1438 316 1466
rect 344 1438 349 1466
rect -349 1400 349 1438
rect -349 1372 -344 1400
rect -316 1372 -278 1400
rect -250 1372 -212 1400
rect -184 1372 -146 1400
rect -118 1372 -80 1400
rect -52 1372 -14 1400
rect 14 1372 52 1400
rect 80 1372 118 1400
rect 146 1372 184 1400
rect 212 1372 250 1400
rect 278 1372 316 1400
rect 344 1372 349 1400
rect -349 1334 349 1372
rect -349 1306 -344 1334
rect -316 1306 -278 1334
rect -250 1306 -212 1334
rect -184 1306 -146 1334
rect -118 1306 -80 1334
rect -52 1306 -14 1334
rect 14 1306 52 1334
rect 80 1306 118 1334
rect 146 1306 184 1334
rect 212 1306 250 1334
rect 278 1306 316 1334
rect 344 1306 349 1334
rect -349 1268 349 1306
rect -349 1240 -344 1268
rect -316 1240 -278 1268
rect -250 1240 -212 1268
rect -184 1240 -146 1268
rect -118 1240 -80 1268
rect -52 1240 -14 1268
rect 14 1240 52 1268
rect 80 1240 118 1268
rect 146 1240 184 1268
rect 212 1240 250 1268
rect 278 1240 316 1268
rect 344 1240 349 1268
rect -349 1202 349 1240
rect -349 1174 -344 1202
rect -316 1174 -278 1202
rect -250 1174 -212 1202
rect -184 1174 -146 1202
rect -118 1174 -80 1202
rect -52 1174 -14 1202
rect 14 1174 52 1202
rect 80 1174 118 1202
rect 146 1174 184 1202
rect 212 1174 250 1202
rect 278 1174 316 1202
rect 344 1174 349 1202
rect -349 1136 349 1174
rect -349 1108 -344 1136
rect -316 1108 -278 1136
rect -250 1108 -212 1136
rect -184 1108 -146 1136
rect -118 1108 -80 1136
rect -52 1108 -14 1136
rect 14 1108 52 1136
rect 80 1108 118 1136
rect 146 1108 184 1136
rect 212 1108 250 1136
rect 278 1108 316 1136
rect 344 1108 349 1136
rect -349 1070 349 1108
rect -349 1042 -344 1070
rect -316 1042 -278 1070
rect -250 1042 -212 1070
rect -184 1042 -146 1070
rect -118 1042 -80 1070
rect -52 1042 -14 1070
rect 14 1042 52 1070
rect 80 1042 118 1070
rect 146 1042 184 1070
rect 212 1042 250 1070
rect 278 1042 316 1070
rect 344 1042 349 1070
rect -349 1004 349 1042
rect -349 976 -344 1004
rect -316 976 -278 1004
rect -250 976 -212 1004
rect -184 976 -146 1004
rect -118 976 -80 1004
rect -52 976 -14 1004
rect 14 976 52 1004
rect 80 976 118 1004
rect 146 976 184 1004
rect 212 976 250 1004
rect 278 976 316 1004
rect 344 976 349 1004
rect -349 938 349 976
rect -349 910 -344 938
rect -316 910 -278 938
rect -250 910 -212 938
rect -184 910 -146 938
rect -118 910 -80 938
rect -52 910 -14 938
rect 14 910 52 938
rect 80 910 118 938
rect 146 910 184 938
rect 212 910 250 938
rect 278 910 316 938
rect 344 910 349 938
rect -349 872 349 910
rect -349 844 -344 872
rect -316 844 -278 872
rect -250 844 -212 872
rect -184 844 -146 872
rect -118 844 -80 872
rect -52 844 -14 872
rect 14 844 52 872
rect 80 844 118 872
rect 146 844 184 872
rect 212 844 250 872
rect 278 844 316 872
rect 344 844 349 872
rect -349 806 349 844
rect -349 778 -344 806
rect -316 778 -278 806
rect -250 778 -212 806
rect -184 778 -146 806
rect -118 778 -80 806
rect -52 778 -14 806
rect 14 778 52 806
rect 80 778 118 806
rect 146 778 184 806
rect 212 778 250 806
rect 278 778 316 806
rect 344 778 349 806
rect -349 740 349 778
rect -349 712 -344 740
rect -316 712 -278 740
rect -250 712 -212 740
rect -184 712 -146 740
rect -118 712 -80 740
rect -52 712 -14 740
rect 14 712 52 740
rect 80 712 118 740
rect 146 712 184 740
rect 212 712 250 740
rect 278 712 316 740
rect 344 712 349 740
rect -349 674 349 712
rect -349 646 -344 674
rect -316 646 -278 674
rect -250 646 -212 674
rect -184 646 -146 674
rect -118 646 -80 674
rect -52 646 -14 674
rect 14 646 52 674
rect 80 646 118 674
rect 146 646 184 674
rect 212 646 250 674
rect 278 646 316 674
rect 344 646 349 674
rect -349 608 349 646
rect -349 580 -344 608
rect -316 580 -278 608
rect -250 580 -212 608
rect -184 580 -146 608
rect -118 580 -80 608
rect -52 580 -14 608
rect 14 580 52 608
rect 80 580 118 608
rect 146 580 184 608
rect 212 580 250 608
rect 278 580 316 608
rect 344 580 349 608
rect -349 542 349 580
rect -349 514 -344 542
rect -316 514 -278 542
rect -250 514 -212 542
rect -184 514 -146 542
rect -118 514 -80 542
rect -52 514 -14 542
rect 14 514 52 542
rect 80 514 118 542
rect 146 514 184 542
rect 212 514 250 542
rect 278 514 316 542
rect 344 514 349 542
rect -349 476 349 514
rect -349 448 -344 476
rect -316 448 -278 476
rect -250 448 -212 476
rect -184 448 -146 476
rect -118 448 -80 476
rect -52 448 -14 476
rect 14 448 52 476
rect 80 448 118 476
rect 146 448 184 476
rect 212 448 250 476
rect 278 448 316 476
rect 344 448 349 476
rect -349 410 349 448
rect -349 382 -344 410
rect -316 382 -278 410
rect -250 382 -212 410
rect -184 382 -146 410
rect -118 382 -80 410
rect -52 382 -14 410
rect 14 382 52 410
rect 80 382 118 410
rect 146 382 184 410
rect 212 382 250 410
rect 278 382 316 410
rect 344 382 349 410
rect -349 344 349 382
rect -349 316 -344 344
rect -316 316 -278 344
rect -250 316 -212 344
rect -184 316 -146 344
rect -118 316 -80 344
rect -52 316 -14 344
rect 14 316 52 344
rect 80 316 118 344
rect 146 316 184 344
rect 212 316 250 344
rect 278 316 316 344
rect 344 316 349 344
rect -349 278 349 316
rect -349 250 -344 278
rect -316 250 -278 278
rect -250 250 -212 278
rect -184 250 -146 278
rect -118 250 -80 278
rect -52 250 -14 278
rect 14 250 52 278
rect 80 250 118 278
rect 146 250 184 278
rect 212 250 250 278
rect 278 250 316 278
rect 344 250 349 278
rect -349 212 349 250
rect -349 184 -344 212
rect -316 184 -278 212
rect -250 184 -212 212
rect -184 184 -146 212
rect -118 184 -80 212
rect -52 184 -14 212
rect 14 184 52 212
rect 80 184 118 212
rect 146 184 184 212
rect 212 184 250 212
rect 278 184 316 212
rect 344 184 349 212
rect -349 146 349 184
rect -349 118 -344 146
rect -316 118 -278 146
rect -250 118 -212 146
rect -184 118 -146 146
rect -118 118 -80 146
rect -52 118 -14 146
rect 14 118 52 146
rect 80 118 118 146
rect 146 118 184 146
rect 212 118 250 146
rect 278 118 316 146
rect 344 118 349 146
rect -349 80 349 118
rect -349 52 -344 80
rect -316 52 -278 80
rect -250 52 -212 80
rect -184 52 -146 80
rect -118 52 -80 80
rect -52 52 -14 80
rect 14 52 52 80
rect 80 52 118 80
rect 146 52 184 80
rect 212 52 250 80
rect 278 52 316 80
rect 344 52 349 80
rect -349 14 349 52
rect -349 -14 -344 14
rect -316 -14 -278 14
rect -250 -14 -212 14
rect -184 -14 -146 14
rect -118 -14 -80 14
rect -52 -14 -14 14
rect 14 -14 52 14
rect 80 -14 118 14
rect 146 -14 184 14
rect 212 -14 250 14
rect 278 -14 316 14
rect 344 -14 349 14
rect -349 -52 349 -14
rect -349 -80 -344 -52
rect -316 -80 -278 -52
rect -250 -80 -212 -52
rect -184 -80 -146 -52
rect -118 -80 -80 -52
rect -52 -80 -14 -52
rect 14 -80 52 -52
rect 80 -80 118 -52
rect 146 -80 184 -52
rect 212 -80 250 -52
rect 278 -80 316 -52
rect 344 -80 349 -52
rect -349 -118 349 -80
rect -349 -146 -344 -118
rect -316 -146 -278 -118
rect -250 -146 -212 -118
rect -184 -146 -146 -118
rect -118 -146 -80 -118
rect -52 -146 -14 -118
rect 14 -146 52 -118
rect 80 -146 118 -118
rect 146 -146 184 -118
rect 212 -146 250 -118
rect 278 -146 316 -118
rect 344 -146 349 -118
rect -349 -184 349 -146
rect -349 -212 -344 -184
rect -316 -212 -278 -184
rect -250 -212 -212 -184
rect -184 -212 -146 -184
rect -118 -212 -80 -184
rect -52 -212 -14 -184
rect 14 -212 52 -184
rect 80 -212 118 -184
rect 146 -212 184 -184
rect 212 -212 250 -184
rect 278 -212 316 -184
rect 344 -212 349 -184
rect -349 -250 349 -212
rect -349 -278 -344 -250
rect -316 -278 -278 -250
rect -250 -278 -212 -250
rect -184 -278 -146 -250
rect -118 -278 -80 -250
rect -52 -278 -14 -250
rect 14 -278 52 -250
rect 80 -278 118 -250
rect 146 -278 184 -250
rect 212 -278 250 -250
rect 278 -278 316 -250
rect 344 -278 349 -250
rect -349 -316 349 -278
rect -349 -344 -344 -316
rect -316 -344 -278 -316
rect -250 -344 -212 -316
rect -184 -344 -146 -316
rect -118 -344 -80 -316
rect -52 -344 -14 -316
rect 14 -344 52 -316
rect 80 -344 118 -316
rect 146 -344 184 -316
rect 212 -344 250 -316
rect 278 -344 316 -316
rect 344 -344 349 -316
rect -349 -382 349 -344
rect -349 -410 -344 -382
rect -316 -410 -278 -382
rect -250 -410 -212 -382
rect -184 -410 -146 -382
rect -118 -410 -80 -382
rect -52 -410 -14 -382
rect 14 -410 52 -382
rect 80 -410 118 -382
rect 146 -410 184 -382
rect 212 -410 250 -382
rect 278 -410 316 -382
rect 344 -410 349 -382
rect -349 -448 349 -410
rect -349 -476 -344 -448
rect -316 -476 -278 -448
rect -250 -476 -212 -448
rect -184 -476 -146 -448
rect -118 -476 -80 -448
rect -52 -476 -14 -448
rect 14 -476 52 -448
rect 80 -476 118 -448
rect 146 -476 184 -448
rect 212 -476 250 -448
rect 278 -476 316 -448
rect 344 -476 349 -448
rect -349 -514 349 -476
rect -349 -542 -344 -514
rect -316 -542 -278 -514
rect -250 -542 -212 -514
rect -184 -542 -146 -514
rect -118 -542 -80 -514
rect -52 -542 -14 -514
rect 14 -542 52 -514
rect 80 -542 118 -514
rect 146 -542 184 -514
rect 212 -542 250 -514
rect 278 -542 316 -514
rect 344 -542 349 -514
rect -349 -580 349 -542
rect -349 -608 -344 -580
rect -316 -608 -278 -580
rect -250 -608 -212 -580
rect -184 -608 -146 -580
rect -118 -608 -80 -580
rect -52 -608 -14 -580
rect 14 -608 52 -580
rect 80 -608 118 -580
rect 146 -608 184 -580
rect 212 -608 250 -580
rect 278 -608 316 -580
rect 344 -608 349 -580
rect -349 -646 349 -608
rect -349 -674 -344 -646
rect -316 -674 -278 -646
rect -250 -674 -212 -646
rect -184 -674 -146 -646
rect -118 -674 -80 -646
rect -52 -674 -14 -646
rect 14 -674 52 -646
rect 80 -674 118 -646
rect 146 -674 184 -646
rect 212 -674 250 -646
rect 278 -674 316 -646
rect 344 -674 349 -646
rect -349 -712 349 -674
rect -349 -740 -344 -712
rect -316 -740 -278 -712
rect -250 -740 -212 -712
rect -184 -740 -146 -712
rect -118 -740 -80 -712
rect -52 -740 -14 -712
rect 14 -740 52 -712
rect 80 -740 118 -712
rect 146 -740 184 -712
rect 212 -740 250 -712
rect 278 -740 316 -712
rect 344 -740 349 -712
rect -349 -778 349 -740
rect -349 -806 -344 -778
rect -316 -806 -278 -778
rect -250 -806 -212 -778
rect -184 -806 -146 -778
rect -118 -806 -80 -778
rect -52 -806 -14 -778
rect 14 -806 52 -778
rect 80 -806 118 -778
rect 146 -806 184 -778
rect 212 -806 250 -778
rect 278 -806 316 -778
rect 344 -806 349 -778
rect -349 -844 349 -806
rect -349 -872 -344 -844
rect -316 -872 -278 -844
rect -250 -872 -212 -844
rect -184 -872 -146 -844
rect -118 -872 -80 -844
rect -52 -872 -14 -844
rect 14 -872 52 -844
rect 80 -872 118 -844
rect 146 -872 184 -844
rect 212 -872 250 -844
rect 278 -872 316 -844
rect 344 -872 349 -844
rect -349 -910 349 -872
rect -349 -938 -344 -910
rect -316 -938 -278 -910
rect -250 -938 -212 -910
rect -184 -938 -146 -910
rect -118 -938 -80 -910
rect -52 -938 -14 -910
rect 14 -938 52 -910
rect 80 -938 118 -910
rect 146 -938 184 -910
rect 212 -938 250 -910
rect 278 -938 316 -910
rect 344 -938 349 -910
rect -349 -976 349 -938
rect -349 -1004 -344 -976
rect -316 -1004 -278 -976
rect -250 -1004 -212 -976
rect -184 -1004 -146 -976
rect -118 -1004 -80 -976
rect -52 -1004 -14 -976
rect 14 -1004 52 -976
rect 80 -1004 118 -976
rect 146 -1004 184 -976
rect 212 -1004 250 -976
rect 278 -1004 316 -976
rect 344 -1004 349 -976
rect -349 -1042 349 -1004
rect -349 -1070 -344 -1042
rect -316 -1070 -278 -1042
rect -250 -1070 -212 -1042
rect -184 -1070 -146 -1042
rect -118 -1070 -80 -1042
rect -52 -1070 -14 -1042
rect 14 -1070 52 -1042
rect 80 -1070 118 -1042
rect 146 -1070 184 -1042
rect 212 -1070 250 -1042
rect 278 -1070 316 -1042
rect 344 -1070 349 -1042
rect -349 -1108 349 -1070
rect -349 -1136 -344 -1108
rect -316 -1136 -278 -1108
rect -250 -1136 -212 -1108
rect -184 -1136 -146 -1108
rect -118 -1136 -80 -1108
rect -52 -1136 -14 -1108
rect 14 -1136 52 -1108
rect 80 -1136 118 -1108
rect 146 -1136 184 -1108
rect 212 -1136 250 -1108
rect 278 -1136 316 -1108
rect 344 -1136 349 -1108
rect -349 -1174 349 -1136
rect -349 -1202 -344 -1174
rect -316 -1202 -278 -1174
rect -250 -1202 -212 -1174
rect -184 -1202 -146 -1174
rect -118 -1202 -80 -1174
rect -52 -1202 -14 -1174
rect 14 -1202 52 -1174
rect 80 -1202 118 -1174
rect 146 -1202 184 -1174
rect 212 -1202 250 -1174
rect 278 -1202 316 -1174
rect 344 -1202 349 -1174
rect -349 -1240 349 -1202
rect -349 -1268 -344 -1240
rect -316 -1268 -278 -1240
rect -250 -1268 -212 -1240
rect -184 -1268 -146 -1240
rect -118 -1268 -80 -1240
rect -52 -1268 -14 -1240
rect 14 -1268 52 -1240
rect 80 -1268 118 -1240
rect 146 -1268 184 -1240
rect 212 -1268 250 -1240
rect 278 -1268 316 -1240
rect 344 -1268 349 -1240
rect -349 -1306 349 -1268
rect -349 -1334 -344 -1306
rect -316 -1334 -278 -1306
rect -250 -1334 -212 -1306
rect -184 -1334 -146 -1306
rect -118 -1334 -80 -1306
rect -52 -1334 -14 -1306
rect 14 -1334 52 -1306
rect 80 -1334 118 -1306
rect 146 -1334 184 -1306
rect 212 -1334 250 -1306
rect 278 -1334 316 -1306
rect 344 -1334 349 -1306
rect -349 -1372 349 -1334
rect -349 -1400 -344 -1372
rect -316 -1400 -278 -1372
rect -250 -1400 -212 -1372
rect -184 -1400 -146 -1372
rect -118 -1400 -80 -1372
rect -52 -1400 -14 -1372
rect 14 -1400 52 -1372
rect 80 -1400 118 -1372
rect 146 -1400 184 -1372
rect 212 -1400 250 -1372
rect 278 -1400 316 -1372
rect 344 -1400 349 -1372
rect -349 -1438 349 -1400
rect -349 -1466 -344 -1438
rect -316 -1466 -278 -1438
rect -250 -1466 -212 -1438
rect -184 -1466 -146 -1438
rect -118 -1466 -80 -1438
rect -52 -1466 -14 -1438
rect 14 -1466 52 -1438
rect 80 -1466 118 -1438
rect 146 -1466 184 -1438
rect 212 -1466 250 -1438
rect 278 -1466 316 -1438
rect 344 -1466 349 -1438
rect -349 -1504 349 -1466
rect -349 -1532 -344 -1504
rect -316 -1532 -278 -1504
rect -250 -1532 -212 -1504
rect -184 -1532 -146 -1504
rect -118 -1532 -80 -1504
rect -52 -1532 -14 -1504
rect 14 -1532 52 -1504
rect 80 -1532 118 -1504
rect 146 -1532 184 -1504
rect 212 -1532 250 -1504
rect 278 -1532 316 -1504
rect 344 -1532 349 -1504
rect -349 -1570 349 -1532
rect -349 -1598 -344 -1570
rect -316 -1598 -278 -1570
rect -250 -1598 -212 -1570
rect -184 -1598 -146 -1570
rect -118 -1598 -80 -1570
rect -52 -1598 -14 -1570
rect 14 -1598 52 -1570
rect 80 -1598 118 -1570
rect 146 -1598 184 -1570
rect 212 -1598 250 -1570
rect 278 -1598 316 -1570
rect 344 -1598 349 -1570
rect -349 -1636 349 -1598
rect -349 -1664 -344 -1636
rect -316 -1664 -278 -1636
rect -250 -1664 -212 -1636
rect -184 -1664 -146 -1636
rect -118 -1664 -80 -1636
rect -52 -1664 -14 -1636
rect 14 -1664 52 -1636
rect 80 -1664 118 -1636
rect 146 -1664 184 -1636
rect 212 -1664 250 -1636
rect 278 -1664 316 -1636
rect 344 -1664 349 -1636
rect -349 -1702 349 -1664
rect -349 -1730 -344 -1702
rect -316 -1730 -278 -1702
rect -250 -1730 -212 -1702
rect -184 -1730 -146 -1702
rect -118 -1730 -80 -1702
rect -52 -1730 -14 -1702
rect 14 -1730 52 -1702
rect 80 -1730 118 -1702
rect 146 -1730 184 -1702
rect 212 -1730 250 -1702
rect 278 -1730 316 -1702
rect 344 -1730 349 -1702
rect -349 -1768 349 -1730
rect -349 -1796 -344 -1768
rect -316 -1796 -278 -1768
rect -250 -1796 -212 -1768
rect -184 -1796 -146 -1768
rect -118 -1796 -80 -1768
rect -52 -1796 -14 -1768
rect 14 -1796 52 -1768
rect 80 -1796 118 -1768
rect 146 -1796 184 -1768
rect 212 -1796 250 -1768
rect 278 -1796 316 -1768
rect 344 -1796 349 -1768
rect -349 -1834 349 -1796
rect -349 -1862 -344 -1834
rect -316 -1862 -278 -1834
rect -250 -1862 -212 -1834
rect -184 -1862 -146 -1834
rect -118 -1862 -80 -1834
rect -52 -1862 -14 -1834
rect 14 -1862 52 -1834
rect 80 -1862 118 -1834
rect 146 -1862 184 -1834
rect 212 -1862 250 -1834
rect 278 -1862 316 -1834
rect 344 -1862 349 -1834
rect -349 -1900 349 -1862
rect -349 -1928 -344 -1900
rect -316 -1928 -278 -1900
rect -250 -1928 -212 -1900
rect -184 -1928 -146 -1900
rect -118 -1928 -80 -1900
rect -52 -1928 -14 -1900
rect 14 -1928 52 -1900
rect 80 -1928 118 -1900
rect 146 -1928 184 -1900
rect 212 -1928 250 -1900
rect 278 -1928 316 -1900
rect 344 -1928 349 -1900
rect -349 -1966 349 -1928
rect -349 -1994 -344 -1966
rect -316 -1994 -278 -1966
rect -250 -1994 -212 -1966
rect -184 -1994 -146 -1966
rect -118 -1994 -80 -1966
rect -52 -1994 -14 -1966
rect 14 -1994 52 -1966
rect 80 -1994 118 -1966
rect 146 -1994 184 -1966
rect 212 -1994 250 -1966
rect 278 -1994 316 -1966
rect 344 -1994 349 -1966
rect -349 -2032 349 -1994
rect -349 -2060 -344 -2032
rect -316 -2060 -278 -2032
rect -250 -2060 -212 -2032
rect -184 -2060 -146 -2032
rect -118 -2060 -80 -2032
rect -52 -2060 -14 -2032
rect 14 -2060 52 -2032
rect 80 -2060 118 -2032
rect 146 -2060 184 -2032
rect 212 -2060 250 -2032
rect 278 -2060 316 -2032
rect 344 -2060 349 -2032
rect -349 -2098 349 -2060
rect -349 -2126 -344 -2098
rect -316 -2126 -278 -2098
rect -250 -2126 -212 -2098
rect -184 -2126 -146 -2098
rect -118 -2126 -80 -2098
rect -52 -2126 -14 -2098
rect 14 -2126 52 -2098
rect 80 -2126 118 -2098
rect 146 -2126 184 -2098
rect 212 -2126 250 -2098
rect 278 -2126 316 -2098
rect 344 -2126 349 -2098
rect -349 -2164 349 -2126
rect -349 -2192 -344 -2164
rect -316 -2192 -278 -2164
rect -250 -2192 -212 -2164
rect -184 -2192 -146 -2164
rect -118 -2192 -80 -2164
rect -52 -2192 -14 -2164
rect 14 -2192 52 -2164
rect 80 -2192 118 -2164
rect 146 -2192 184 -2164
rect 212 -2192 250 -2164
rect 278 -2192 316 -2164
rect 344 -2192 349 -2164
rect -349 -2230 349 -2192
rect -349 -2258 -344 -2230
rect -316 -2258 -278 -2230
rect -250 -2258 -212 -2230
rect -184 -2258 -146 -2230
rect -118 -2258 -80 -2230
rect -52 -2258 -14 -2230
rect 14 -2258 52 -2230
rect 80 -2258 118 -2230
rect 146 -2258 184 -2230
rect 212 -2258 250 -2230
rect 278 -2258 316 -2230
rect 344 -2258 349 -2230
rect -349 -2296 349 -2258
rect -349 -2324 -344 -2296
rect -316 -2324 -278 -2296
rect -250 -2324 -212 -2296
rect -184 -2324 -146 -2296
rect -118 -2324 -80 -2296
rect -52 -2324 -14 -2296
rect 14 -2324 52 -2296
rect 80 -2324 118 -2296
rect 146 -2324 184 -2296
rect 212 -2324 250 -2296
rect 278 -2324 316 -2296
rect 344 -2324 349 -2296
rect -349 -2362 349 -2324
rect -349 -2390 -344 -2362
rect -316 -2390 -278 -2362
rect -250 -2390 -212 -2362
rect -184 -2390 -146 -2362
rect -118 -2390 -80 -2362
rect -52 -2390 -14 -2362
rect 14 -2390 52 -2362
rect 80 -2390 118 -2362
rect 146 -2390 184 -2362
rect 212 -2390 250 -2362
rect 278 -2390 316 -2362
rect 344 -2390 349 -2362
rect -349 -2428 349 -2390
rect -349 -2456 -344 -2428
rect -316 -2456 -278 -2428
rect -250 -2456 -212 -2428
rect -184 -2456 -146 -2428
rect -118 -2456 -80 -2428
rect -52 -2456 -14 -2428
rect 14 -2456 52 -2428
rect 80 -2456 118 -2428
rect 146 -2456 184 -2428
rect 212 -2456 250 -2428
rect 278 -2456 316 -2428
rect 344 -2456 349 -2428
rect -349 -2494 349 -2456
rect -349 -2522 -344 -2494
rect -316 -2522 -278 -2494
rect -250 -2522 -212 -2494
rect -184 -2522 -146 -2494
rect -118 -2522 -80 -2494
rect -52 -2522 -14 -2494
rect 14 -2522 52 -2494
rect 80 -2522 118 -2494
rect 146 -2522 184 -2494
rect 212 -2522 250 -2494
rect 278 -2522 316 -2494
rect 344 -2522 349 -2494
rect -349 -2560 349 -2522
rect -349 -2588 -344 -2560
rect -316 -2588 -278 -2560
rect -250 -2588 -212 -2560
rect -184 -2588 -146 -2560
rect -118 -2588 -80 -2560
rect -52 -2588 -14 -2560
rect 14 -2588 52 -2560
rect 80 -2588 118 -2560
rect 146 -2588 184 -2560
rect 212 -2588 250 -2560
rect 278 -2588 316 -2560
rect 344 -2588 349 -2560
rect -349 -2626 349 -2588
rect -349 -2654 -344 -2626
rect -316 -2654 -278 -2626
rect -250 -2654 -212 -2626
rect -184 -2654 -146 -2626
rect -118 -2654 -80 -2626
rect -52 -2654 -14 -2626
rect 14 -2654 52 -2626
rect 80 -2654 118 -2626
rect 146 -2654 184 -2626
rect 212 -2654 250 -2626
rect 278 -2654 316 -2626
rect 344 -2654 349 -2626
rect -349 -2692 349 -2654
rect -349 -2720 -344 -2692
rect -316 -2720 -278 -2692
rect -250 -2720 -212 -2692
rect -184 -2720 -146 -2692
rect -118 -2720 -80 -2692
rect -52 -2720 -14 -2692
rect 14 -2720 52 -2692
rect 80 -2720 118 -2692
rect 146 -2720 184 -2692
rect 212 -2720 250 -2692
rect 278 -2720 316 -2692
rect 344 -2720 349 -2692
rect -349 -2758 349 -2720
rect -349 -2786 -344 -2758
rect -316 -2786 -278 -2758
rect -250 -2786 -212 -2758
rect -184 -2786 -146 -2758
rect -118 -2786 -80 -2758
rect -52 -2786 -14 -2758
rect 14 -2786 52 -2758
rect 80 -2786 118 -2758
rect 146 -2786 184 -2758
rect 212 -2786 250 -2758
rect 278 -2786 316 -2758
rect 344 -2786 349 -2758
rect -349 -2824 349 -2786
rect -349 -2852 -344 -2824
rect -316 -2852 -278 -2824
rect -250 -2852 -212 -2824
rect -184 -2852 -146 -2824
rect -118 -2852 -80 -2824
rect -52 -2852 -14 -2824
rect 14 -2852 52 -2824
rect 80 -2852 118 -2824
rect 146 -2852 184 -2824
rect 212 -2852 250 -2824
rect 278 -2852 316 -2824
rect 344 -2852 349 -2824
rect -349 -2890 349 -2852
rect -349 -2918 -344 -2890
rect -316 -2918 -278 -2890
rect -250 -2918 -212 -2890
rect -184 -2918 -146 -2890
rect -118 -2918 -80 -2890
rect -52 -2918 -14 -2890
rect 14 -2918 52 -2890
rect 80 -2918 118 -2890
rect 146 -2918 184 -2890
rect 212 -2918 250 -2890
rect 278 -2918 316 -2890
rect 344 -2918 349 -2890
rect -349 -2956 349 -2918
rect -349 -2984 -344 -2956
rect -316 -2984 -278 -2956
rect -250 -2984 -212 -2956
rect -184 -2984 -146 -2956
rect -118 -2984 -80 -2956
rect -52 -2984 -14 -2956
rect 14 -2984 52 -2956
rect 80 -2984 118 -2956
rect 146 -2984 184 -2956
rect 212 -2984 250 -2956
rect 278 -2984 316 -2956
rect 344 -2984 349 -2956
rect -349 -3022 349 -2984
rect -349 -3050 -344 -3022
rect -316 -3050 -278 -3022
rect -250 -3050 -212 -3022
rect -184 -3050 -146 -3022
rect -118 -3050 -80 -3022
rect -52 -3050 -14 -3022
rect 14 -3050 52 -3022
rect 80 -3050 118 -3022
rect 146 -3050 184 -3022
rect 212 -3050 250 -3022
rect 278 -3050 316 -3022
rect 344 -3050 349 -3022
rect -349 -3088 349 -3050
rect -349 -3116 -344 -3088
rect -316 -3116 -278 -3088
rect -250 -3116 -212 -3088
rect -184 -3116 -146 -3088
rect -118 -3116 -80 -3088
rect -52 -3116 -14 -3088
rect 14 -3116 52 -3088
rect 80 -3116 118 -3088
rect 146 -3116 184 -3088
rect 212 -3116 250 -3088
rect 278 -3116 316 -3088
rect 344 -3116 349 -3088
rect -349 -3154 349 -3116
rect -349 -3182 -344 -3154
rect -316 -3182 -278 -3154
rect -250 -3182 -212 -3154
rect -184 -3182 -146 -3154
rect -118 -3182 -80 -3154
rect -52 -3182 -14 -3154
rect 14 -3182 52 -3154
rect 80 -3182 118 -3154
rect 146 -3182 184 -3154
rect 212 -3182 250 -3154
rect 278 -3182 316 -3154
rect 344 -3182 349 -3154
rect -349 -3220 349 -3182
rect -349 -3248 -344 -3220
rect -316 -3248 -278 -3220
rect -250 -3248 -212 -3220
rect -184 -3248 -146 -3220
rect -118 -3248 -80 -3220
rect -52 -3248 -14 -3220
rect 14 -3248 52 -3220
rect 80 -3248 118 -3220
rect 146 -3248 184 -3220
rect 212 -3248 250 -3220
rect 278 -3248 316 -3220
rect 344 -3248 349 -3220
rect -349 -3286 349 -3248
rect -349 -3314 -344 -3286
rect -316 -3314 -278 -3286
rect -250 -3314 -212 -3286
rect -184 -3314 -146 -3286
rect -118 -3314 -80 -3286
rect -52 -3314 -14 -3286
rect 14 -3314 52 -3286
rect 80 -3314 118 -3286
rect 146 -3314 184 -3286
rect 212 -3314 250 -3286
rect 278 -3314 316 -3286
rect 344 -3314 349 -3286
rect -349 -3352 349 -3314
rect -349 -3380 -344 -3352
rect -316 -3380 -278 -3352
rect -250 -3380 -212 -3352
rect -184 -3380 -146 -3352
rect -118 -3380 -80 -3352
rect -52 -3380 -14 -3352
rect 14 -3380 52 -3352
rect 80 -3380 118 -3352
rect 146 -3380 184 -3352
rect 212 -3380 250 -3352
rect 278 -3380 316 -3352
rect 344 -3380 349 -3352
rect -349 -3385 349 -3380
<< end >>
