* NGSPICE file created from TG_Layout_flat_flat.ext - technology: gf180mcuC

.subckt TG_Layout_flat_flat VSS CLK VIN VOUT VDD
X0 VOUT Inverter_Layout_0.OUT.t1 VIN.t38 VDD.t15 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1 VOUT Inverter_Layout_0.OUT.t2 VIN.t37 VDD.t14 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X2 VIN CLK.t0 VOUT.t56 VSS.t7 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X3 VOUT CLK.t1 VIN.t59 VSS.t6 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X4 VOUT CLK.t2 VIN.t0 VSS.t5 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X5 VIN Inverter_Layout_0.OUT.t3 VOUT.t50 VDD.t7 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X6 VOUT Inverter_Layout_0.OUT.t4 VIN.t36 VDD.t12 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X7 VOUT Inverter_Layout_0.OUT.t5 VIN.t35 VDD.t6 pfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X8 VOUT Inverter_Layout_0.OUT.t6 VIN.t34 VDD.t5 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X9 VIN Inverter_Layout_0.OUT.t7 VOUT.t46 VDD.t9 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X10 VOUT CLK.t4 VIN.t66 VSS.t3 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X11 VIN CLK.t5 VOUT.t70 VSS.t2 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X12 VIN Inverter_Layout_0.OUT.t8 VOUT.t45 VDD.t3 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X13 VIN Inverter_Layout_0.OUT.t9 VOUT.t44 VDD.t1 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X14 VIN CLK.t6 VOUT.t54 VSS.t4 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X15 VOUT CLK.t7 VIN.t60 VSS.t1 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X16 VOUT Inverter_Layout_0.OUT.t10 VIN.t33 VDD.t2 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X17 VOUT Inverter_Layout_0.OUT.t11 VIN.t32 VDD.t13 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X18 VOUT Inverter_Layout_0.OUT.t12 VIN.t31 VDD.t15 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X19 VOUT Inverter_Layout_0.OUT.t13 VIN.t30 VDD.t14 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X20 VIN Inverter_Layout_0.OUT.t14 VOUT.t39 VDD.t0 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X21 VIN Inverter_Layout_0.OUT.t15 VOUT.t38 VDD.t10 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X22 VIN CLK.t8 VOUT.t64 VSS.t7 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X23 VIN Inverter_Layout_0.OUT.t16 VOUT.t37 VDD.t11 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X24 VOUT CLK.t9 VIN.t61 VSS.t6 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X25 VOUT Inverter_Layout_0.OUT.t17 VIN.t29 VDD.t8 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X26 VIN Inverter_Layout_0.OUT.t18 VOUT.t35 VDD.t4 pfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X27 VIN Inverter_Layout_0.OUT.t19 VOUT.t34 VDD.t7 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X28 VIN CLK.t10 VOUT.t68 VSS.t0 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X29 VOUT Inverter_Layout_0.OUT.t20 VIN.t28 VDD.t6 pfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X30 VOUT Inverter_Layout_0.OUT.t21 VIN.t27 VDD.t5 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X31 VOUT CLK.t11 VIN.t4 VSS.t5 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X32 VIN Inverter_Layout_0.OUT.t22 VOUT.t31 VDD.t3 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X33 VIN CLK.t13 VOUT.t62 VSS.t4 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X34 VOUT CLK.t14 VIN.t53 VSS.t1 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X35 VOUT Inverter_Layout_0.OUT.t23 VIN.t26 VDD.t13 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X36 VIN Inverter_Layout_0.OUT.t24 VOUT.t29 VDD.t1 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X37 VIN Inverter_Layout_0.OUT.t25 VOUT.t28 VDD.t11 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X38 VIN Inverter_Layout_0.OUT.t26 VOUT.t27 VDD.t10 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X39 VOUT Inverter_Layout_0.OUT.t27 VIN.t25 VDD.t15 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X40 VOUT Inverter_Layout_0.OUT.t28 VIN.t24 VDD.t14 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X41 VOUT Inverter_Layout_0.OUT.t29 VIN.t23 VDD.t8 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X42 VOUT CLK.t15 VIN.t71 VSS.t3 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X43 VIN CLK.t16 VOUT.t69 VSS.t7 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X44 VOUT Inverter_Layout_0.OUT.t30 VIN.t22 VDD.t12 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X45 VIN CLK.t17 VOUT.t58 VSS.t2 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X46 VOUT CLK.t18 VIN.t63 VSS.t6 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X47 VIN Inverter_Layout_0.OUT.t31 VOUT.t22 VDD.t9 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X48 VIN Inverter_Layout_0.OUT.t32 VOUT.t21 VDD.t4 pfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X49 VOUT Inverter_Layout_0.OUT.t33 VIN.t21 VDD.t2 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X50 VIN CLK.t19 VOUT.t3 VSS.t0 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X51 VIN Inverter_Layout_0.OUT.t34 VOUT.t19 VDD.t0 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X52 VOUT CLK.t20 VIN.t55 VSS.t5 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X53 VIN CLK.t21 VOUT.t57 VSS.t4 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X54 VOUT Inverter_Layout_0.OUT.t35 VIN.t20 VDD.t13 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X55 VOUT Inverter_Layout_0.OUT.t36 VIN.t19 VDD.t12 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X56 VIN Inverter_Layout_0.OUT.t37 VOUT.t16 VDD.t11 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X57 VIN Inverter_Layout_0.OUT.t38 VOUT.t15 VDD.t10 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X58 VIN Inverter_Layout_0.OUT.t39 VOUT.t14 VDD.t9 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X59 VOUT Inverter_Layout_0.OUT.t40 VIN.t18 VDD.t8 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X60 VOUT CLK.t22 VIN.t65 VSS.t3 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X61 VIN Inverter_Layout_0.OUT.t41 VOUT.t12 VDD.t7 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X62 VIN CLK.t23 VOUT.t1 VSS.t2 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X63 VOUT Inverter_Layout_0.OUT.t42 VIN.t17 VDD.t6 pfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X64 VOUT Inverter_Layout_0.OUT.t43 VIN.t16 VDD.t5 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X65 VIN Inverter_Layout_0.OUT.t44 VOUT.t9 VDD.t4 pfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X66 VOUT CLK.t24 VIN.t67 VSS.t1 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X67 VIN Inverter_Layout_0.OUT.t45 VOUT.t8 VDD.t3 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X68 VOUT Inverter_Layout_0.OUT.t46 VIN.t15 VDD.t2 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X69 VIN Inverter_Layout_0.OUT.t47 VOUT.t6 VDD.t1 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X70 VIN Inverter_Layout_0.OUT.t48 VOUT.t5 VDD.t0 pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X71 VIN CLK.t25 VOUT.t2 VSS.t0 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
R0 Inverter_Layout_0.OUT.t3 Inverter_Layout_0.OUT.t19 50.3184
R1 Inverter_Layout_0.OUT.t41 Inverter_Layout_0.OUT.t3 50.3184
R2 Inverter_Layout_0.OUT.t36 Inverter_Layout_0.OUT.t4 50.3184
R3 Inverter_Layout_0.OUT.t30 Inverter_Layout_0.OUT.t36 50.3184
R4 Inverter_Layout_0.OUT.t25 Inverter_Layout_0.OUT.t37 50.3184
R5 Inverter_Layout_0.OUT.t16 Inverter_Layout_0.OUT.t25 50.3184
R6 Inverter_Layout_0.OUT.t23 Inverter_Layout_0.OUT.t35 50.3184
R7 Inverter_Layout_0.OUT.t11 Inverter_Layout_0.OUT.t23 50.3184
R8 Inverter_Layout_0.OUT.t8 Inverter_Layout_0.OUT.t22 50.3184
R9 Inverter_Layout_0.OUT.t45 Inverter_Layout_0.OUT.t8 50.3184
R10 Inverter_Layout_0.OUT.t6 Inverter_Layout_0.OUT.t21 50.3184
R11 Inverter_Layout_0.OUT.t43 Inverter_Layout_0.OUT.t6 50.3184
R12 Inverter_Layout_0.OUT.t39 Inverter_Layout_0.OUT.t7 50.3184
R13 Inverter_Layout_0.OUT.t31 Inverter_Layout_0.OUT.t39 50.3184
R14 Inverter_Layout_0.OUT.t29 Inverter_Layout_0.OUT.t40 50.3184
R15 Inverter_Layout_0.OUT.t17 Inverter_Layout_0.OUT.t29 50.3184
R16 Inverter_Layout_0.OUT.t26 Inverter_Layout_0.OUT.t38 50.3184
R17 Inverter_Layout_0.OUT.t15 Inverter_Layout_0.OUT.t26 50.3184
R18 Inverter_Layout_0.OUT.t12 Inverter_Layout_0.OUT.t27 50.3184
R19 Inverter_Layout_0.OUT.t1 Inverter_Layout_0.OUT.t12 50.3184
R20 Inverter_Layout_0.OUT.t9 Inverter_Layout_0.OUT.t24 50.3184
R21 Inverter_Layout_0.OUT.t47 Inverter_Layout_0.OUT.t9 50.3184
R22 Inverter_Layout_0.OUT.t13 Inverter_Layout_0.OUT.t28 50.3184
R23 Inverter_Layout_0.OUT.t2 Inverter_Layout_0.OUT.t13 50.3184
R24 Inverter_Layout_0.OUT.t48 Inverter_Layout_0.OUT.t14 50.3184
R25 Inverter_Layout_0.OUT.t34 Inverter_Layout_0.OUT.t48 50.3184
R26 Inverter_Layout_0.OUT.t46 Inverter_Layout_0.OUT.t10 50.3184
R27 Inverter_Layout_0.OUT.t33 Inverter_Layout_0.OUT.t46 50.3184
R28 Inverter_Layout_0.OUT.t32 Inverter_Layout_0.OUT.t44 50.3184
R29 Inverter_Layout_0.OUT.t18 Inverter_Layout_0.OUT.t32 50.3184
R30 Inverter_Layout_0.OUT.t5 Inverter_Layout_0.OUT.t42 50.3184
R31 Inverter_Layout_0.OUT.t20 Inverter_Layout_0.OUT.t5 50.3184
R32 Inverter_Layout_0.OUT.n14 Inverter_Layout_0.OUT.t20 48.7834
R33 Inverter_Layout_0.OUT.n0 Inverter_Layout_0.OUT.t18 39.7594
R34 Inverter_Layout_0.OUT.t42 Inverter_Layout_0.OUT.n13 39.7594
R35 Inverter_Layout_0.OUT.n1 Inverter_Layout_0.OUT.n0 20.8576
R36 Inverter_Layout_0.OUT.n2 Inverter_Layout_0.OUT.n1 20.8576
R37 Inverter_Layout_0.OUT.n3 Inverter_Layout_0.OUT.n2 20.8576
R38 Inverter_Layout_0.OUT.n4 Inverter_Layout_0.OUT.n3 20.8576
R39 Inverter_Layout_0.OUT.n5 Inverter_Layout_0.OUT.n4 20.8576
R40 Inverter_Layout_0.OUT.n6 Inverter_Layout_0.OUT.n5 20.8576
R41 Inverter_Layout_0.OUT.n7 Inverter_Layout_0.OUT.n6 20.8576
R42 Inverter_Layout_0.OUT.n8 Inverter_Layout_0.OUT.n7 20.8576
R43 Inverter_Layout_0.OUT.n9 Inverter_Layout_0.OUT.n8 20.8576
R44 Inverter_Layout_0.OUT.n10 Inverter_Layout_0.OUT.n9 20.8576
R45 Inverter_Layout_0.OUT.n11 Inverter_Layout_0.OUT.n10 20.8576
R46 Inverter_Layout_0.OUT.n12 Inverter_Layout_0.OUT.n11 20.8576
R47 Inverter_Layout_0.OUT.n13 Inverter_Layout_0.OUT.n12 20.8576
R48 Inverter_Layout_0.OUT.n13 Inverter_Layout_0.OUT.t41 18.9023
R49 Inverter_Layout_0.OUT.n12 Inverter_Layout_0.OUT.t30 18.9023
R50 Inverter_Layout_0.OUT.n11 Inverter_Layout_0.OUT.t16 18.9023
R51 Inverter_Layout_0.OUT.n10 Inverter_Layout_0.OUT.t11 18.9023
R52 Inverter_Layout_0.OUT.n9 Inverter_Layout_0.OUT.t45 18.9023
R53 Inverter_Layout_0.OUT.n8 Inverter_Layout_0.OUT.t43 18.9023
R54 Inverter_Layout_0.OUT.n7 Inverter_Layout_0.OUT.t31 18.9023
R55 Inverter_Layout_0.OUT.n6 Inverter_Layout_0.OUT.t17 18.9023
R56 Inverter_Layout_0.OUT.n5 Inverter_Layout_0.OUT.t15 18.9023
R57 Inverter_Layout_0.OUT.n4 Inverter_Layout_0.OUT.t1 18.9023
R58 Inverter_Layout_0.OUT.n3 Inverter_Layout_0.OUT.t47 18.9023
R59 Inverter_Layout_0.OUT.n2 Inverter_Layout_0.OUT.t2 18.9023
R60 Inverter_Layout_0.OUT.n1 Inverter_Layout_0.OUT.t34 18.9023
R61 Inverter_Layout_0.OUT.n0 Inverter_Layout_0.OUT.t33 18.9023
R62 Inverter_Layout_0.OUT.n14 Inverter_Layout_0.OUT.t0 4.4205
R63 Inverter_Layout_0.OUT Inverter_Layout_0.OUT.n14 0.4505
R64 VIN.n73 VIN.n72 4.81172
R65 VIN.n104 VIN.n2 4.4609
R66 VIN.n105 VIN.n1 4.4609
R67 VIN.n106 VIN.n0 4.4609
R68 VIN.n100 VIN.t67 4.4609
R69 VIN.n101 VIN.t60 4.4609
R70 VIN.n102 VIN.t53 4.4609
R71 VIN.n95 VIN.t17 4.0565
R72 VIN.n96 VIN.t35 4.0565
R73 VIN.n97 VIN.t28 4.0565
R74 VIN.n74 VIN.n70 4.0565
R75 VIN.n73 VIN.n71 4.0565
R76 VIN.n26 VIN.n25 3.90572
R77 VIN.n9 VIN.n8 3.90572
R78 VIN.n32 VIN.n29 3.35572
R79 VIN.n46 VIN.n43 3.35572
R80 VIN.n86 VIN.n83 3.35572
R81 VIN.n63 VIN.n60 3.35572
R82 VIN.n26 VIN.n23 3.1505
R83 VIN.n27 VIN.n21 3.1505
R84 VIN.n9 VIN.n6 3.1505
R85 VIN.n10 VIN.n4 3.1505
R86 VIN.n13 VIN.n12 3.1505
R87 VIN.n16 VIN.n15 3.1505
R88 VIN.n19 VIN.n18 3.1505
R89 VIN.n32 VIN.n31 2.6005
R90 VIN.n35 VIN.n34 2.6005
R91 VIN.n46 VIN.n45 2.6005
R92 VIN.n49 VIN.n48 2.6005
R93 VIN.n50 VIN.n41 2.6005
R94 VIN.n51 VIN.n39 2.6005
R95 VIN.n52 VIN.n37 2.6005
R96 VIN.n86 VIN.n85 2.6005
R97 VIN.n89 VIN.n88 2.6005
R98 VIN.n63 VIN.n62 2.6005
R99 VIN.n66 VIN.n65 2.6005
R100 VIN.n67 VIN.n58 2.6005
R101 VIN.n68 VIN.n56 2.6005
R102 VIN.n69 VIN.n54 2.6005
R103 VIN.n90 VIN.n81 2.6005
R104 VIN.n91 VIN.n79 2.6005
R105 VIN.n92 VIN.n77 2.6005
R106 VIN.n95 VIN.n94 2.47941
R107 VIN.n103 VIN.n102 2.47941
R108 VIN.n93 VIN.n75 2.05876
R109 VIN.n34 VIN.t36 1.4565
R110 VIN.n34 VIN.n33 1.4565
R111 VIN.n31 VIN.t19 1.4565
R112 VIN.n31 VIN.n30 1.4565
R113 VIN.n29 VIN.t22 1.4565
R114 VIN.n29 VIN.n28 1.4565
R115 VIN.n37 VIN.t16 1.4565
R116 VIN.n37 VIN.n36 1.4565
R117 VIN.n39 VIN.t34 1.4565
R118 VIN.n39 VIN.n38 1.4565
R119 VIN.n41 VIN.t27 1.4565
R120 VIN.n41 VIN.n40 1.4565
R121 VIN.n48 VIN.t20 1.4565
R122 VIN.n48 VIN.n47 1.4565
R123 VIN.n45 VIN.t26 1.4565
R124 VIN.n45 VIN.n44 1.4565
R125 VIN.n43 VIN.t32 1.4565
R126 VIN.n43 VIN.n42 1.4565
R127 VIN.n77 VIN.t29 1.4565
R128 VIN.n77 VIN.n76 1.4565
R129 VIN.n79 VIN.t23 1.4565
R130 VIN.n79 VIN.n78 1.4565
R131 VIN.n81 VIN.t18 1.4565
R132 VIN.n81 VIN.n80 1.4565
R133 VIN.n88 VIN.t25 1.4565
R134 VIN.n88 VIN.n87 1.4565
R135 VIN.n85 VIN.t31 1.4565
R136 VIN.n85 VIN.n84 1.4565
R137 VIN.n83 VIN.t38 1.4565
R138 VIN.n83 VIN.n82 1.4565
R139 VIN.n54 VIN.t21 1.4565
R140 VIN.n54 VIN.n53 1.4565
R141 VIN.n56 VIN.t15 1.4565
R142 VIN.n56 VIN.n55 1.4565
R143 VIN.n58 VIN.t33 1.4565
R144 VIN.n58 VIN.n57 1.4565
R145 VIN.n65 VIN.t24 1.4565
R146 VIN.n65 VIN.n64 1.4565
R147 VIN.n62 VIN.t30 1.4565
R148 VIN.n62 VIN.n61 1.4565
R149 VIN.n60 VIN.t37 1.4565
R150 VIN.n60 VIN.n59 1.4565
R151 VIN.n21 VIN.t71 1.3109
R152 VIN.n21 VIN.n20 1.3109
R153 VIN.n23 VIN.t65 1.3109
R154 VIN.n23 VIN.n22 1.3109
R155 VIN.n25 VIN.t66 1.3109
R156 VIN.n25 VIN.n24 1.3109
R157 VIN.n18 VIN.t63 1.3109
R158 VIN.n18 VIN.n17 1.3109
R159 VIN.n15 VIN.t61 1.3109
R160 VIN.n15 VIN.n14 1.3109
R161 VIN.n12 VIN.t59 1.3109
R162 VIN.n12 VIN.n11 1.3109
R163 VIN.n4 VIN.t4 1.3109
R164 VIN.n4 VIN.n3 1.3109
R165 VIN.n6 VIN.t55 1.3109
R166 VIN.n6 VIN.n5 1.3109
R167 VIN.n8 VIN.t0 1.3109
R168 VIN.n8 VIN.n7 1.3109
R169 VIN.n50 VIN.n49 1.28789
R170 VIN.n90 VIN.n89 1.28789
R171 VIN.n67 VIN.n66 1.28789
R172 VIN.n13 VIN.n10 1.28789
R173 VIN.n75 VIN.n74 0.957239
R174 VIN.n98 VIN.n97 0.957239
R175 VIN.n99 VIN.n27 0.957239
R176 VIN.n104 VIN.n103 0.957239
R177 VIN.n99 VIN.n98 0.896587
R178 VIN.n35 VIN.n32 0.755717
R179 VIN.n49 VIN.n46 0.755717
R180 VIN.n52 VIN.n51 0.755717
R181 VIN.n51 VIN.n50 0.755717
R182 VIN.n89 VIN.n86 0.755717
R183 VIN.n66 VIN.n63 0.755717
R184 VIN.n69 VIN.n68 0.755717
R185 VIN.n68 VIN.n67 0.755717
R186 VIN.n74 VIN.n73 0.755717
R187 VIN.n92 VIN.n91 0.755717
R188 VIN.n91 VIN.n90 0.755717
R189 VIN.n96 VIN.n95 0.755717
R190 VIN.n97 VIN.n96 0.755717
R191 VIN.n27 VIN.n26 0.755717
R192 VIN.n101 VIN.n100 0.755717
R193 VIN.n102 VIN.n101 0.755717
R194 VIN.n10 VIN.n9 0.755717
R195 VIN.n16 VIN.n13 0.755717
R196 VIN.n19 VIN.n16 0.755717
R197 VIN.n106 VIN.n105 0.755717
R198 VIN.n105 VIN.n104 0.755717
R199 VIN.n94 VIN.n93 0.626587
R200 VIN VIN.n106 0.513109
R201 VIN.n98 VIN.n35 0.331152
R202 VIN.n94 VIN.n52 0.331152
R203 VIN.n75 VIN.n69 0.331152
R204 VIN.n93 VIN.n92 0.331152
R205 VIN.n100 VIN.n99 0.331152
R206 VIN.n103 VIN.n19 0.331152
R207 VOUT.n40 VOUT.n39 3.90572
R208 VOUT.n60 VOUT.n57 3.90572
R209 VOUT.n68 VOUT.n65 3.90572
R210 VOUT.n4 VOUT.n1 3.35572
R211 VOUT.n22 VOUT.n21 3.35572
R212 VOUT.n14 VOUT.n13 3.35572
R213 VOUT.n46 VOUT.n43 3.35572
R214 VOUT.n90 VOUT.n89 3.35572
R215 VOUT.n82 VOUT.n81 3.35572
R216 VOUT.n40 VOUT.n37 3.1505
R217 VOUT.n41 VOUT.n35 3.1505
R218 VOUT.n60 VOUT.n59 3.1505
R219 VOUT.n63 VOUT.n62 3.1505
R220 VOUT.n68 VOUT.n67 3.1505
R221 VOUT.n71 VOUT.n70 3.1505
R222 VOUT.n73 VOUT.n55 3.1505
R223 VOUT.n74 VOUT.n53 3.1505
R224 VOUT.n75 VOUT.n51 3.1505
R225 VOUT.n4 VOUT.n3 2.6005
R226 VOUT.n7 VOUT.n6 2.6005
R227 VOUT.n22 VOUT.n19 2.6005
R228 VOUT.n23 VOUT.n17 2.6005
R229 VOUT.n14 VOUT.n11 2.6005
R230 VOUT.n15 VOUT.n9 2.6005
R231 VOUT.n27 VOUT.n26 2.6005
R232 VOUT.n30 VOUT.n29 2.6005
R233 VOUT.n33 VOUT.n32 2.6005
R234 VOUT.n46 VOUT.n45 2.6005
R235 VOUT.n49 VOUT.n48 2.6005
R236 VOUT.n90 VOUT.n87 2.6005
R237 VOUT.n91 VOUT.n85 2.6005
R238 VOUT.n82 VOUT.n79 2.6005
R239 VOUT.n83 VOUT.n77 2.6005
R240 VOUT.n101 VOUT.n100 2.6005
R241 VOUT.n98 VOUT.n97 2.6005
R242 VOUT.n95 VOUT.n94 2.6005
R243 VOUT.n102 VOUT.n101 1.76333
R244 VOUT.n6 VOUT.t9 1.4565
R245 VOUT.n6 VOUT.n5 1.4565
R246 VOUT.n3 VOUT.t21 1.4565
R247 VOUT.n3 VOUT.n2 1.4565
R248 VOUT.n1 VOUT.t35 1.4565
R249 VOUT.n1 VOUT.n0 1.4565
R250 VOUT.n32 VOUT.t29 1.4565
R251 VOUT.n32 VOUT.n31 1.4565
R252 VOUT.n29 VOUT.t44 1.4565
R253 VOUT.n29 VOUT.n28 1.4565
R254 VOUT.n26 VOUT.t6 1.4565
R255 VOUT.n26 VOUT.n25 1.4565
R256 VOUT.n17 VOUT.t38 1.4565
R257 VOUT.n17 VOUT.n16 1.4565
R258 VOUT.n19 VOUT.t27 1.4565
R259 VOUT.n19 VOUT.n18 1.4565
R260 VOUT.n21 VOUT.t15 1.4565
R261 VOUT.n21 VOUT.n20 1.4565
R262 VOUT.n9 VOUT.t19 1.4565
R263 VOUT.n9 VOUT.n8 1.4565
R264 VOUT.n11 VOUT.t5 1.4565
R265 VOUT.n11 VOUT.n10 1.4565
R266 VOUT.n13 VOUT.t39 1.4565
R267 VOUT.n13 VOUT.n12 1.4565
R268 VOUT.n48 VOUT.t46 1.4565
R269 VOUT.n48 VOUT.n47 1.4565
R270 VOUT.n45 VOUT.t14 1.4565
R271 VOUT.n45 VOUT.n44 1.4565
R272 VOUT.n43 VOUT.t22 1.4565
R273 VOUT.n43 VOUT.n42 1.4565
R274 VOUT.n94 VOUT.t37 1.4565
R275 VOUT.n94 VOUT.n93 1.4565
R276 VOUT.n97 VOUT.t28 1.4565
R277 VOUT.n97 VOUT.n96 1.4565
R278 VOUT.n100 VOUT.t16 1.4565
R279 VOUT.n100 VOUT.n99 1.4565
R280 VOUT.n85 VOUT.t12 1.4565
R281 VOUT.n85 VOUT.n84 1.4565
R282 VOUT.n87 VOUT.t50 1.4565
R283 VOUT.n87 VOUT.n86 1.4565
R284 VOUT.n89 VOUT.t34 1.4565
R285 VOUT.n89 VOUT.n88 1.4565
R286 VOUT.n77 VOUT.t8 1.4565
R287 VOUT.n77 VOUT.n76 1.4565
R288 VOUT.n79 VOUT.t45 1.4565
R289 VOUT.n79 VOUT.n78 1.4565
R290 VOUT.n81 VOUT.t31 1.4565
R291 VOUT.n81 VOUT.n80 1.4565
R292 VOUT.n35 VOUT.t54 1.3109
R293 VOUT.n35 VOUT.n34 1.3109
R294 VOUT.n37 VOUT.t62 1.3109
R295 VOUT.n37 VOUT.n36 1.3109
R296 VOUT.n39 VOUT.t57 1.3109
R297 VOUT.n39 VOUT.n38 1.3109
R298 VOUT.n51 VOUT.t56 1.3109
R299 VOUT.n51 VOUT.n50 1.3109
R300 VOUT.n53 VOUT.t64 1.3109
R301 VOUT.n53 VOUT.n52 1.3109
R302 VOUT.n55 VOUT.t69 1.3109
R303 VOUT.n55 VOUT.n54 1.3109
R304 VOUT.n62 VOUT.t70 1.3109
R305 VOUT.n62 VOUT.n61 1.3109
R306 VOUT.n59 VOUT.t1 1.3109
R307 VOUT.n59 VOUT.n58 1.3109
R308 VOUT.n57 VOUT.t58 1.3109
R309 VOUT.n57 VOUT.n56 1.3109
R310 VOUT.n70 VOUT.t2 1.3109
R311 VOUT.n70 VOUT.n69 1.3109
R312 VOUT.n67 VOUT.t3 1.3109
R313 VOUT.n67 VOUT.n66 1.3109
R314 VOUT.n65 VOUT.t68 1.3109
R315 VOUT.n65 VOUT.n64 1.3109
R316 VOUT.n104 VOUT.n103 1.25267
R317 VOUT.n103 VOUT.n102 1.25267
R318 VOUT.n24 VOUT.n23 0.957239
R319 VOUT.n24 VOUT.n15 0.957239
R320 VOUT.n72 VOUT.n63 0.957239
R321 VOUT.n72 VOUT.n71 0.957239
R322 VOUT.n92 VOUT.n91 0.957239
R323 VOUT.n92 VOUT.n83 0.957239
R324 VOUT.n7 VOUT.n4 0.755717
R325 VOUT.n23 VOUT.n22 0.755717
R326 VOUT.n15 VOUT.n14 0.755717
R327 VOUT.n30 VOUT.n27 0.755717
R328 VOUT.n33 VOUT.n30 0.755717
R329 VOUT.n41 VOUT.n40 0.755717
R330 VOUT.n63 VOUT.n60 0.755717
R331 VOUT.n71 VOUT.n68 0.755717
R332 VOUT.n49 VOUT.n46 0.755717
R333 VOUT.n75 VOUT.n74 0.755717
R334 VOUT.n74 VOUT.n73 0.755717
R335 VOUT.n91 VOUT.n90 0.755717
R336 VOUT.n83 VOUT.n82 0.755717
R337 VOUT.n98 VOUT.n95 0.755717
R338 VOUT.n101 VOUT.n98 0.755717
R339 VOUT.n104 VOUT.n7 0.511152
R340 VOUT.n103 VOUT.n33 0.511152
R341 VOUT.n103 VOUT.n41 0.511152
R342 VOUT.n102 VOUT.n49 0.511152
R343 VOUT.n102 VOUT.n75 0.511152
R344 VOUT.n27 VOUT.n24 0.331152
R345 VOUT.n73 VOUT.n72 0.331152
R346 VOUT.n95 VOUT.n92 0.331152
R347 VOUT VOUT.n104 0.0885435
R348 VDD.n2 VDD.n1 945.545
R349 VDD.n2 VDD.t16 527.229
R350 VDD.t2 VDD.t4 124.805
R351 VDD.t0 VDD.t2 124.805
R352 VDD.t14 VDD.t0 124.805
R353 VDD.t1 VDD.t14 124.805
R354 VDD.t15 VDD.t1 124.805
R355 VDD.t10 VDD.t15 124.805
R356 VDD.t8 VDD.t10 124.805
R357 VDD.t9 VDD.t8 124.805
R358 VDD.t5 VDD.t9 124.805
R359 VDD.t3 VDD.t5 124.805
R360 VDD.t13 VDD.t3 124.805
R361 VDD.t11 VDD.t13 124.805
R362 VDD.t12 VDD.t11 124.805
R363 VDD.t7 VDD.t6 124.805
R364 VDD.n1 VDD.t12 94.3843
R365 VDD.n1 VDD.t7 30.4217
R366 VDD VDD.n2 6.3005
R367 VDD VDD.n0 4.78572
R368 CLK.t13 CLK.t6 50.3184
R369 CLK.t21 CLK.t13 50.3184
R370 CLK.t9 CLK.t1 50.3184
R371 CLK.t18 CLK.t9 50.3184
R372 CLK.t23 CLK.t17 50.3184
R373 CLK.t5 CLK.t23 50.3184
R374 CLK.t20 CLK.t11 50.3184
R375 CLK.t2 CLK.t20 50.3184
R376 CLK.t8 CLK.t0 50.3184
R377 CLK.t16 CLK.t8 50.3184
R378 CLK.t22 CLK.t15 50.3184
R379 CLK.t4 CLK.t22 50.3184
R380 CLK.t19 CLK.t10 50.3184
R381 CLK.t25 CLK.t19 50.3184
R382 CLK.t7 CLK.t24 50.3184
R383 CLK.t14 CLK.t7 50.3184
R384 CLK CLK.n6 48.1123
R385 CLK.n0 CLK.t21 39.7594
R386 CLK.n7 CLK.t12 29.3309
R387 CLK.n1 CLK.n0 20.8576
R388 CLK.n2 CLK.n1 20.8576
R389 CLK.n3 CLK.n2 20.8576
R390 CLK.n4 CLK.n3 20.8576
R391 CLK.n5 CLK.n4 20.8576
R392 CLK.n6 CLK.n5 20.8576
R393 CLK.n0 CLK.t18 18.9023
R394 CLK.n1 CLK.t5 18.9023
R395 CLK.n2 CLK.t2 18.9023
R396 CLK.n3 CLK.t16 18.9023
R397 CLK.n4 CLK.t4 18.9023
R398 CLK.n5 CLK.t25 18.9023
R399 CLK.n6 CLK.t14 18.9023
R400 CLK.n7 CLK.t3 18.3809
R401 CLK CLK.n7 17.6692
R402 VSS.n1 VSS.t1 558.01
R403 VSS.n1 VSS.t8 495.854
R404 VSS VSS.n1 414.82
R405 VSS.t6 VSS.t4 373.563
R406 VSS.t2 VSS.t6 373.563
R407 VSS.t5 VSS.t2 373.563
R408 VSS.t7 VSS.t5 373.563
R409 VSS.t3 VSS.t7 373.563
R410 VSS.t0 VSS.t3 373.563
R411 VSS.t1 VSS.t0 373.563
R412 VSS VSS.n0 6.68867
C0 VOUT VIN 15.9f
C1 CLK VIN 0.575f
C2 Inverter_Layout_0.OUT VIN 0.753f
C3 CLK VOUT 0.318f
C4 Inverter_Layout_0.OUT VOUT 0.623f
C5 CLK Inverter_Layout_0.OUT 0.0797f
C6 VOUT 0 1.1f
C7 VIN 0 2.79f
C8 CLK 0 3.35f
C9 Inverter_Layout_0.OUT 0 2.39f
C10 VDD.n0 0 0.0129f
C11 VDD.t4 0 0.345f
C12 VDD.t2 0 0.196f
C13 VDD.t0 0 0.196f
C14 VDD.t14 0 0.196f
C15 VDD.t1 0 0.196f
C16 VDD.t15 0 0.196f
C17 VDD.t10 0 0.196f
C18 VDD.t8 0 0.196f
C19 VDD.t9 0 0.196f
C20 VDD.t5 0 0.196f
C21 VDD.t3 0 0.196f
C22 VDD.t13 0 0.196f
C23 VDD.t11 0 0.196f
C24 VDD.t12 0 0.172f
C25 VDD.t6 0 0.345f
C26 VDD.t7 0 0.122f
C27 VDD.n1 0 0.172f
C28 VDD.t16 0 0.13f
C29 VDD.n2 0 0.119f
C30 VOUT.t35 0 0.0592f
C31 VOUT.n0 0 0.0592f
C32 VOUT.n1 0 0.148f
C33 VOUT.t21 0 0.0592f
C34 VOUT.n2 0 0.0592f
C35 VOUT.n3 0 0.118f
C36 VOUT.n4 0 0.264f
C37 VOUT.t9 0 0.0592f
C38 VOUT.n5 0 0.0592f
C39 VOUT.n6 0 0.118f
C40 VOUT.n7 0 0.136f
C41 VOUT.t19 0 0.0592f
C42 VOUT.n8 0 0.0592f
C43 VOUT.n9 0 0.118f
C44 VOUT.t5 0 0.0592f
C45 VOUT.n10 0 0.0592f
C46 VOUT.n11 0 0.118f
C47 VOUT.t39 0 0.0592f
C48 VOUT.n12 0 0.0592f
C49 VOUT.n13 0 0.148f
C50 VOUT.n14 0 0.264f
C51 VOUT.n15 0 0.19f
C52 VOUT.t38 0 0.0592f
C53 VOUT.n16 0 0.0592f
C54 VOUT.n17 0 0.118f
C55 VOUT.t27 0 0.0592f
C56 VOUT.n18 0 0.0592f
C57 VOUT.n19 0 0.118f
C58 VOUT.t15 0 0.0592f
C59 VOUT.n20 0 0.0592f
C60 VOUT.n21 0 0.148f
C61 VOUT.n22 0 0.264f
C62 VOUT.n23 0 0.19f
C63 VOUT.n24 0 0.247f
C64 VOUT.t6 0 0.0592f
C65 VOUT.n25 0 0.0592f
C66 VOUT.n26 0 0.118f
C67 VOUT.n27 0 0.116f
C68 VOUT.t44 0 0.0592f
C69 VOUT.n28 0 0.0592f
C70 VOUT.n29 0 0.118f
C71 VOUT.n30 0 0.162f
C72 VOUT.t29 0 0.0592f
C73 VOUT.n31 0 0.0592f
C74 VOUT.n32 0 0.118f
C75 VOUT.n33 0 0.136f
C76 VOUT.t54 0 0.0592f
C77 VOUT.n34 0 0.0592f
C78 VOUT.n35 0 0.118f
C79 VOUT.t62 0 0.0592f
C80 VOUT.n36 0 0.0592f
C81 VOUT.n37 0 0.118f
C82 VOUT.t57 0 0.0592f
C83 VOUT.n38 0 0.0592f
C84 VOUT.n39 0 0.144f
C85 VOUT.n40 0 0.269f
C86 VOUT.n41 0 0.136f
C87 VOUT.t22 0 0.0592f
C88 VOUT.n42 0 0.0592f
C89 VOUT.n43 0 0.148f
C90 VOUT.t14 0 0.0592f
C91 VOUT.n44 0 0.0592f
C92 VOUT.n45 0 0.118f
C93 VOUT.n46 0 0.264f
C94 VOUT.t46 0 0.0592f
C95 VOUT.n47 0 0.0592f
C96 VOUT.n48 0 0.118f
C97 VOUT.n49 0 0.136f
C98 VOUT.t56 0 0.0592f
C99 VOUT.n50 0 0.0592f
C100 VOUT.n51 0 0.118f
C101 VOUT.t64 0 0.0592f
C102 VOUT.n52 0 0.0592f
C103 VOUT.n53 0 0.118f
C104 VOUT.t69 0 0.0592f
C105 VOUT.n54 0 0.0592f
C106 VOUT.n55 0 0.118f
C107 VOUT.t58 0 0.0592f
C108 VOUT.n56 0 0.0592f
C109 VOUT.n57 0 0.144f
C110 VOUT.t1 0 0.0592f
C111 VOUT.n58 0 0.0592f
C112 VOUT.n59 0 0.118f
C113 VOUT.n60 0 0.269f
C114 VOUT.t70 0 0.0592f
C115 VOUT.n61 0 0.0592f
C116 VOUT.n62 0 0.118f
C117 VOUT.n63 0 0.19f
C118 VOUT.t68 0 0.0592f
C119 VOUT.n64 0 0.0592f
C120 VOUT.n65 0 0.144f
C121 VOUT.t3 0 0.0592f
C122 VOUT.n66 0 0.0592f
C123 VOUT.n67 0 0.118f
C124 VOUT.n68 0 0.269f
C125 VOUT.t2 0 0.0592f
C126 VOUT.n69 0 0.0592f
C127 VOUT.n70 0 0.118f
C128 VOUT.n71 0 0.19f
C129 VOUT.n72 0 0.247f
C130 VOUT.n73 0 0.116f
C131 VOUT.n74 0 0.162f
C132 VOUT.n75 0 0.136f
C133 VOUT.t8 0 0.0592f
C134 VOUT.n76 0 0.0592f
C135 VOUT.n77 0 0.118f
C136 VOUT.t45 0 0.0592f
C137 VOUT.n78 0 0.0592f
C138 VOUT.n79 0 0.118f
C139 VOUT.t31 0 0.0592f
C140 VOUT.n80 0 0.0592f
C141 VOUT.n81 0 0.148f
C142 VOUT.n82 0 0.264f
C143 VOUT.n83 0 0.19f
C144 VOUT.t12 0 0.0592f
C145 VOUT.n84 0 0.0592f
C146 VOUT.n85 0 0.118f
C147 VOUT.t50 0 0.0592f
C148 VOUT.n86 0 0.0592f
C149 VOUT.n87 0 0.118f
C150 VOUT.t34 0 0.0592f
C151 VOUT.n88 0 0.0592f
C152 VOUT.n89 0 0.148f
C153 VOUT.n90 0 0.264f
C154 VOUT.n91 0 0.19f
C155 VOUT.n92 0 0.247f
C156 VOUT.t37 0 0.0592f
C157 VOUT.n93 0 0.0592f
C158 VOUT.n94 0 0.118f
C159 VOUT.n95 0 0.116f
C160 VOUT.t28 0 0.0592f
C161 VOUT.n96 0 0.0592f
C162 VOUT.n97 0 0.118f
C163 VOUT.n98 0 0.162f
C164 VOUT.t16 0 0.0592f
C165 VOUT.n99 0 0.0592f
C166 VOUT.n100 0 0.118f
C167 VOUT.n101 0 0.277f
C168 VOUT.n102 0 0.435f
C169 VOUT.n103 0 0.378f
C170 VOUT.n104 0 0.198f
C171 VIN.n0 0 0.133f
C172 VIN.n1 0 0.133f
C173 VIN.n2 0 0.133f
C174 VIN.t4 0 0.0496f
C175 VIN.n3 0 0.0496f
C176 VIN.n4 0 0.0993f
C177 VIN.t55 0 0.0496f
C178 VIN.n5 0 0.0496f
C179 VIN.n6 0 0.0993f
C180 VIN.t0 0 0.0496f
C181 VIN.n7 0 0.0496f
C182 VIN.n8 0 0.121f
C183 VIN.n9 0 0.225f
C184 VIN.n10 0 0.191f
C185 VIN.t59 0 0.0496f
C186 VIN.n11 0 0.0496f
C187 VIN.n12 0 0.0993f
C188 VIN.n13 0 0.191f
C189 VIN.t61 0 0.0496f
C190 VIN.n14 0 0.0496f
C191 VIN.n15 0 0.0993f
C192 VIN.n16 0 0.136f
C193 VIN.t63 0 0.0496f
C194 VIN.n17 0 0.0496f
C195 VIN.n18 0 0.0993f
C196 VIN.n19 0 0.0975f
C197 VIN.t71 0 0.0496f
C198 VIN.n20 0 0.0496f
C199 VIN.n21 0 0.0993f
C200 VIN.t65 0 0.0496f
C201 VIN.n22 0 0.0496f
C202 VIN.n23 0 0.0993f
C203 VIN.t66 0 0.0496f
C204 VIN.n24 0 0.0496f
C205 VIN.n25 0 0.121f
C206 VIN.n26 0 0.225f
C207 VIN.n27 0 0.159f
C208 VIN.t22 0 0.0496f
C209 VIN.n28 0 0.0496f
C210 VIN.n29 0 0.124f
C211 VIN.t19 0 0.0496f
C212 VIN.n30 0 0.0496f
C213 VIN.n31 0 0.0993f
C214 VIN.n32 0 0.222f
C215 VIN.t36 0 0.0496f
C216 VIN.n33 0 0.0496f
C217 VIN.n34 0 0.0993f
C218 VIN.n35 0 0.0975f
C219 VIN.t16 0 0.0496f
C220 VIN.n36 0 0.0496f
C221 VIN.n37 0 0.0993f
C222 VIN.t34 0 0.0496f
C223 VIN.n38 0 0.0496f
C224 VIN.n39 0 0.0993f
C225 VIN.t27 0 0.0496f
C226 VIN.n40 0 0.0496f
C227 VIN.n41 0 0.0993f
C228 VIN.t32 0 0.0496f
C229 VIN.n42 0 0.0496f
C230 VIN.n43 0 0.124f
C231 VIN.t26 0 0.0496f
C232 VIN.n44 0 0.0496f
C233 VIN.n45 0 0.0993f
C234 VIN.n46 0 0.222f
C235 VIN.t20 0 0.0496f
C236 VIN.n47 0 0.0496f
C237 VIN.n48 0 0.0993f
C238 VIN.n49 0 0.191f
C239 VIN.n50 0 0.191f
C240 VIN.n51 0 0.136f
C241 VIN.n52 0 0.0975f
C242 VIN.t21 0 0.0496f
C243 VIN.n53 0 0.0496f
C244 VIN.n54 0 0.0993f
C245 VIN.t15 0 0.0496f
C246 VIN.n55 0 0.0496f
C247 VIN.n56 0 0.0993f
C248 VIN.t33 0 0.0496f
C249 VIN.n57 0 0.0496f
C250 VIN.n58 0 0.0993f
C251 VIN.t37 0 0.0496f
C252 VIN.n59 0 0.0496f
C253 VIN.n60 0 0.124f
C254 VIN.t30 0 0.0496f
C255 VIN.n61 0 0.0496f
C256 VIN.n62 0 0.0993f
C257 VIN.n63 0 0.222f
C258 VIN.t24 0 0.0496f
C259 VIN.n64 0 0.0496f
C260 VIN.n65 0 0.0993f
C261 VIN.n66 0 0.192f
C262 VIN.n67 0 0.192f
C263 VIN.n68 0 0.136f
C264 VIN.n69 0 0.0975f
C265 VIN.n70 0 0.126f
C266 VIN.n71 0 0.126f
C267 VIN.n72 0 0.15f
C268 VIN.n73 0 0.307f
C269 VIN.n74 0 0.201f
C270 VIN.n75 0 0.319f
C271 VIN.t29 0 0.0496f
C272 VIN.n76 0 0.0496f
C273 VIN.n77 0 0.0993f
C274 VIN.t23 0 0.0496f
C275 VIN.n78 0 0.0496f
C276 VIN.n79 0 0.0993f
C277 VIN.t18 0 0.0496f
C278 VIN.n80 0 0.0496f
C279 VIN.n81 0 0.0993f
C280 VIN.t38 0 0.0496f
C281 VIN.n82 0 0.0496f
C282 VIN.n83 0 0.124f
C283 VIN.t31 0 0.0496f
C284 VIN.n84 0 0.0496f
C285 VIN.n85 0 0.0993f
C286 VIN.n86 0 0.222f
C287 VIN.t25 0 0.0496f
C288 VIN.n87 0 0.0496f
C289 VIN.n88 0 0.0993f
C290 VIN.n89 0 0.191f
C291 VIN.n90 0 0.191f
C292 VIN.n91 0 0.136f
C293 VIN.n92 0 0.0975f
C294 VIN.n93 0 0.287f
C295 VIN.n94 0 0.326f
C296 VIN.t17 0 0.126f
C297 VIN.n95 0 0.34f
C298 VIN.t35 0 0.126f
C299 VIN.n96 0 0.178f
C300 VIN.t28 0 0.126f
C301 VIN.n97 0 0.201f
C302 VIN.n98 0 0.213f
C303 VIN.n99 0 0.201f
C304 VIN.t67 0 0.133f
C305 VIN.n100 0 0.132f
C306 VIN.t60 0 0.133f
C307 VIN.n101 0 0.17f
C308 VIN.t53 0 0.133f
C309 VIN.n102 0 0.332f
C310 VIN.n103 0 0.358f
C311 VIN.n104 0 0.194f
C312 VIN.n105 0 0.17f
C313 VIN.n106 0 0.152f
C314 Inverter_Layout_0.OUT.t19 0 0.0514f
C315 Inverter_Layout_0.OUT.t3 0 0.0724f
C316 Inverter_Layout_0.OUT.t41 0 0.0498f
C317 Inverter_Layout_0.OUT.t4 0 0.0514f
C318 Inverter_Layout_0.OUT.t36 0 0.0724f
C319 Inverter_Layout_0.OUT.t30 0 0.0498f
C320 Inverter_Layout_0.OUT.t37 0 0.0514f
C321 Inverter_Layout_0.OUT.t25 0 0.0724f
C322 Inverter_Layout_0.OUT.t16 0 0.0498f
C323 Inverter_Layout_0.OUT.t35 0 0.0514f
C324 Inverter_Layout_0.OUT.t23 0 0.0724f
C325 Inverter_Layout_0.OUT.t11 0 0.0498f
C326 Inverter_Layout_0.OUT.t22 0 0.0514f
C327 Inverter_Layout_0.OUT.t8 0 0.0724f
C328 Inverter_Layout_0.OUT.t45 0 0.0498f
C329 Inverter_Layout_0.OUT.t21 0 0.0514f
C330 Inverter_Layout_0.OUT.t6 0 0.0724f
C331 Inverter_Layout_0.OUT.t43 0 0.0498f
C332 Inverter_Layout_0.OUT.t7 0 0.0514f
C333 Inverter_Layout_0.OUT.t39 0 0.0724f
C334 Inverter_Layout_0.OUT.t31 0 0.0498f
C335 Inverter_Layout_0.OUT.t40 0 0.0514f
C336 Inverter_Layout_0.OUT.t29 0 0.0724f
C337 Inverter_Layout_0.OUT.t17 0 0.0498f
C338 Inverter_Layout_0.OUT.t38 0 0.0514f
C339 Inverter_Layout_0.OUT.t26 0 0.0724f
C340 Inverter_Layout_0.OUT.t15 0 0.0498f
C341 Inverter_Layout_0.OUT.t27 0 0.0514f
C342 Inverter_Layout_0.OUT.t12 0 0.0724f
C343 Inverter_Layout_0.OUT.t1 0 0.0498f
C344 Inverter_Layout_0.OUT.t24 0 0.0514f
C345 Inverter_Layout_0.OUT.t9 0 0.0724f
C346 Inverter_Layout_0.OUT.t47 0 0.0498f
C347 Inverter_Layout_0.OUT.t28 0 0.0514f
C348 Inverter_Layout_0.OUT.t13 0 0.0724f
C349 Inverter_Layout_0.OUT.t2 0 0.0498f
C350 Inverter_Layout_0.OUT.t14 0 0.0514f
C351 Inverter_Layout_0.OUT.t48 0 0.0724f
C352 Inverter_Layout_0.OUT.t34 0 0.0498f
C353 Inverter_Layout_0.OUT.t10 0 0.0514f
C354 Inverter_Layout_0.OUT.t46 0 0.0724f
C355 Inverter_Layout_0.OUT.t33 0 0.0498f
C356 Inverter_Layout_0.OUT.t44 0 0.0514f
C357 Inverter_Layout_0.OUT.t32 0 0.0724f
C358 Inverter_Layout_0.OUT.t18 0 0.0676f
C359 Inverter_Layout_0.OUT.n0 0 0.0597f
C360 Inverter_Layout_0.OUT.n1 0 0.0436f
C361 Inverter_Layout_0.OUT.n2 0 0.0436f
C362 Inverter_Layout_0.OUT.n3 0 0.0436f
C363 Inverter_Layout_0.OUT.n4 0 0.0436f
C364 Inverter_Layout_0.OUT.n5 0 0.0436f
C365 Inverter_Layout_0.OUT.n6 0 0.0436f
C366 Inverter_Layout_0.OUT.n7 0 0.0436f
C367 Inverter_Layout_0.OUT.n8 0 0.0436f
C368 Inverter_Layout_0.OUT.n9 0 0.0436f
C369 Inverter_Layout_0.OUT.n10 0 0.0436f
C370 Inverter_Layout_0.OUT.n11 0 0.0436f
C371 Inverter_Layout_0.OUT.n12 0 0.0436f
C372 Inverter_Layout_0.OUT.n13 0 0.0597f
C373 Inverter_Layout_0.OUT.t42 0 0.0676f
C374 Inverter_Layout_0.OUT.t5 0 0.0724f
C375 Inverter_Layout_0.OUT.t20 0 0.0737f
C376 Inverter_Layout_0.OUT.t0 0 0.0419f
C377 Inverter_Layout_0.OUT.n14 0 0.179f
.ends

