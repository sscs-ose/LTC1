magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2045 -30395 2045 30395
<< psubdiff >>
rect -45 28364 45 28395
rect -45 -28364 -23 28364
rect 23 -28364 45 28364
rect -45 -28395 45 -28364
<< psubdiffcont >>
rect -23 -28364 23 28364
<< metal1 >>
rect -34 28364 34 28384
rect -34 -28364 -23 28364
rect 23 -28364 34 28364
rect -34 -28384 34 -28364
<< end >>
