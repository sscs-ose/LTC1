* NGSPICE file created from folded_cascode_check3_flat.ext - technology: gf180mcuC


* Top level circuit folded_cascode_check3_flat

C0 m1_n2767_n4043# m3_n1726_n4250# 0.0166f
C1 m1_n2607_n3890# m3_n1726_n4250# 0.00594f
C2 w_n3327_n4250# m1_n3088_n4204# 0.348f
C3 m1_n2767_n4043# w_n3327_n4250# 0.38f
C4 m1_n2607_n3890# w_n3327_n4250# 0.162f
C5 m1_n2767_n4043# a_n2438_n4035# 0.00347f
C6 w_n3327_n4250# m3_n2833_n4250# 0.0389f
C7 w_n3327_n4250# m3_n1726_n4250# 0.0434f
C8 m1_n2767_n4043# m1_n3088_n4204# 0.524f
C9 m1_n2607_n3890# m1_n3088_n4204# 0.166f
C10 m1_n2767_n4043# m1_n2607_n3890# 0.315f
C11 m1_n3088_n4204# m3_n2833_n4250# 0.0355f
C12 m1_n2767_n4043# m3_n2833_n4250# 0.048f
C13 m1_n2607_n3890# m3_n2833_n4250# 0.0958f
C14 m1_n3088_n4204# m3_n1726_n4250# 0.133f
C15 m3_n1726_n4250# VSUBS 0.0741f $ **FLOATING
C16 m3_n2833_n4250# VSUBS 0.0693f $ **FLOATING
C17 m1_n3088_n4204# VSUBS 0.479f $ **FLOATING
C18 m1_n2767_n4043# VSUBS 0.413f $ **FLOATING
C19 m1_n2607_n3890# VSUBS 0.216f $ **FLOATING
C20 w_n3327_n4250# VSUBS 3.59f $ **FLOATING
.end

