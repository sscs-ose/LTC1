magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2995 -4495 2995 4495
<< psubdiff >>
rect -995 2473 995 2495
rect -995 -2473 -973 2473
rect 973 -2473 995 2473
rect -995 -2495 995 -2473
<< psubdiffcont >>
rect -973 -2473 973 2473
<< metal1 >>
rect -984 2473 984 2484
rect -984 -2473 -973 2473
rect 973 -2473 984 2473
rect -984 -2484 984 -2473
<< end >>
