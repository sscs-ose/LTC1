magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1045 -2972 1045 2972
<< metal1 >>
rect -45 1966 45 1972
rect -45 1940 -39 1966
rect 39 1940 45 1966
rect -45 1904 45 1940
rect -45 1878 -39 1904
rect 39 1878 45 1904
rect -45 1842 45 1878
rect -45 1816 -39 1842
rect 39 1816 45 1842
rect -45 1780 45 1816
rect -45 1754 -39 1780
rect 39 1754 45 1780
rect -45 1718 45 1754
rect -45 1692 -39 1718
rect 39 1692 45 1718
rect -45 1656 45 1692
rect -45 1630 -39 1656
rect 39 1630 45 1656
rect -45 1594 45 1630
rect -45 1568 -39 1594
rect 39 1568 45 1594
rect -45 1532 45 1568
rect -45 1506 -39 1532
rect 39 1506 45 1532
rect -45 1470 45 1506
rect -45 1444 -39 1470
rect 39 1444 45 1470
rect -45 1408 45 1444
rect -45 1382 -39 1408
rect 39 1382 45 1408
rect -45 1346 45 1382
rect -45 1320 -39 1346
rect 39 1320 45 1346
rect -45 1284 45 1320
rect -45 1258 -39 1284
rect 39 1258 45 1284
rect -45 1222 45 1258
rect -45 1196 -39 1222
rect 39 1196 45 1222
rect -45 1160 45 1196
rect -45 1134 -39 1160
rect 39 1134 45 1160
rect -45 1098 45 1134
rect -45 1072 -39 1098
rect 39 1072 45 1098
rect -45 1036 45 1072
rect -45 1010 -39 1036
rect 39 1010 45 1036
rect -45 974 45 1010
rect -45 948 -39 974
rect 39 948 45 974
rect -45 912 45 948
rect -45 886 -39 912
rect 39 886 45 912
rect -45 850 45 886
rect -45 824 -39 850
rect 39 824 45 850
rect -45 788 45 824
rect -45 762 -39 788
rect 39 762 45 788
rect -45 726 45 762
rect -45 700 -39 726
rect 39 700 45 726
rect -45 664 45 700
rect -45 638 -39 664
rect 39 638 45 664
rect -45 602 45 638
rect -45 576 -39 602
rect 39 576 45 602
rect -45 540 45 576
rect -45 514 -39 540
rect 39 514 45 540
rect -45 478 45 514
rect -45 452 -39 478
rect 39 452 45 478
rect -45 416 45 452
rect -45 390 -39 416
rect 39 390 45 416
rect -45 354 45 390
rect -45 328 -39 354
rect 39 328 45 354
rect -45 292 45 328
rect -45 266 -39 292
rect 39 266 45 292
rect -45 230 45 266
rect -45 204 -39 230
rect 39 204 45 230
rect -45 168 45 204
rect -45 142 -39 168
rect 39 142 45 168
rect -45 106 45 142
rect -45 80 -39 106
rect 39 80 45 106
rect -45 44 45 80
rect -45 18 -39 44
rect 39 18 45 44
rect -45 -18 45 18
rect -45 -44 -39 -18
rect 39 -44 45 -18
rect -45 -80 45 -44
rect -45 -106 -39 -80
rect 39 -106 45 -80
rect -45 -142 45 -106
rect -45 -168 -39 -142
rect 39 -168 45 -142
rect -45 -204 45 -168
rect -45 -230 -39 -204
rect 39 -230 45 -204
rect -45 -266 45 -230
rect -45 -292 -39 -266
rect 39 -292 45 -266
rect -45 -328 45 -292
rect -45 -354 -39 -328
rect 39 -354 45 -328
rect -45 -390 45 -354
rect -45 -416 -39 -390
rect 39 -416 45 -390
rect -45 -452 45 -416
rect -45 -478 -39 -452
rect 39 -478 45 -452
rect -45 -514 45 -478
rect -45 -540 -39 -514
rect 39 -540 45 -514
rect -45 -576 45 -540
rect -45 -602 -39 -576
rect 39 -602 45 -576
rect -45 -638 45 -602
rect -45 -664 -39 -638
rect 39 -664 45 -638
rect -45 -700 45 -664
rect -45 -726 -39 -700
rect 39 -726 45 -700
rect -45 -762 45 -726
rect -45 -788 -39 -762
rect 39 -788 45 -762
rect -45 -824 45 -788
rect -45 -850 -39 -824
rect 39 -850 45 -824
rect -45 -886 45 -850
rect -45 -912 -39 -886
rect 39 -912 45 -886
rect -45 -948 45 -912
rect -45 -974 -39 -948
rect 39 -974 45 -948
rect -45 -1010 45 -974
rect -45 -1036 -39 -1010
rect 39 -1036 45 -1010
rect -45 -1072 45 -1036
rect -45 -1098 -39 -1072
rect 39 -1098 45 -1072
rect -45 -1134 45 -1098
rect -45 -1160 -39 -1134
rect 39 -1160 45 -1134
rect -45 -1196 45 -1160
rect -45 -1222 -39 -1196
rect 39 -1222 45 -1196
rect -45 -1258 45 -1222
rect -45 -1284 -39 -1258
rect 39 -1284 45 -1258
rect -45 -1320 45 -1284
rect -45 -1346 -39 -1320
rect 39 -1346 45 -1320
rect -45 -1382 45 -1346
rect -45 -1408 -39 -1382
rect 39 -1408 45 -1382
rect -45 -1444 45 -1408
rect -45 -1470 -39 -1444
rect 39 -1470 45 -1444
rect -45 -1506 45 -1470
rect -45 -1532 -39 -1506
rect 39 -1532 45 -1506
rect -45 -1568 45 -1532
rect -45 -1594 -39 -1568
rect 39 -1594 45 -1568
rect -45 -1630 45 -1594
rect -45 -1656 -39 -1630
rect 39 -1656 45 -1630
rect -45 -1692 45 -1656
rect -45 -1718 -39 -1692
rect 39 -1718 45 -1692
rect -45 -1754 45 -1718
rect -45 -1780 -39 -1754
rect 39 -1780 45 -1754
rect -45 -1816 45 -1780
rect -45 -1842 -39 -1816
rect 39 -1842 45 -1816
rect -45 -1878 45 -1842
rect -45 -1904 -39 -1878
rect 39 -1904 45 -1878
rect -45 -1940 45 -1904
rect -45 -1966 -39 -1940
rect 39 -1966 45 -1940
rect -45 -1972 45 -1966
<< via1 >>
rect -39 1940 39 1966
rect -39 1878 39 1904
rect -39 1816 39 1842
rect -39 1754 39 1780
rect -39 1692 39 1718
rect -39 1630 39 1656
rect -39 1568 39 1594
rect -39 1506 39 1532
rect -39 1444 39 1470
rect -39 1382 39 1408
rect -39 1320 39 1346
rect -39 1258 39 1284
rect -39 1196 39 1222
rect -39 1134 39 1160
rect -39 1072 39 1098
rect -39 1010 39 1036
rect -39 948 39 974
rect -39 886 39 912
rect -39 824 39 850
rect -39 762 39 788
rect -39 700 39 726
rect -39 638 39 664
rect -39 576 39 602
rect -39 514 39 540
rect -39 452 39 478
rect -39 390 39 416
rect -39 328 39 354
rect -39 266 39 292
rect -39 204 39 230
rect -39 142 39 168
rect -39 80 39 106
rect -39 18 39 44
rect -39 -44 39 -18
rect -39 -106 39 -80
rect -39 -168 39 -142
rect -39 -230 39 -204
rect -39 -292 39 -266
rect -39 -354 39 -328
rect -39 -416 39 -390
rect -39 -478 39 -452
rect -39 -540 39 -514
rect -39 -602 39 -576
rect -39 -664 39 -638
rect -39 -726 39 -700
rect -39 -788 39 -762
rect -39 -850 39 -824
rect -39 -912 39 -886
rect -39 -974 39 -948
rect -39 -1036 39 -1010
rect -39 -1098 39 -1072
rect -39 -1160 39 -1134
rect -39 -1222 39 -1196
rect -39 -1284 39 -1258
rect -39 -1346 39 -1320
rect -39 -1408 39 -1382
rect -39 -1470 39 -1444
rect -39 -1532 39 -1506
rect -39 -1594 39 -1568
rect -39 -1656 39 -1630
rect -39 -1718 39 -1692
rect -39 -1780 39 -1754
rect -39 -1842 39 -1816
rect -39 -1904 39 -1878
rect -39 -1966 39 -1940
<< metal2 >>
rect -45 1966 45 1972
rect -45 1940 -39 1966
rect 39 1940 45 1966
rect -45 1904 45 1940
rect -45 1878 -39 1904
rect 39 1878 45 1904
rect -45 1842 45 1878
rect -45 1816 -39 1842
rect 39 1816 45 1842
rect -45 1780 45 1816
rect -45 1754 -39 1780
rect 39 1754 45 1780
rect -45 1718 45 1754
rect -45 1692 -39 1718
rect 39 1692 45 1718
rect -45 1656 45 1692
rect -45 1630 -39 1656
rect 39 1630 45 1656
rect -45 1594 45 1630
rect -45 1568 -39 1594
rect 39 1568 45 1594
rect -45 1532 45 1568
rect -45 1506 -39 1532
rect 39 1506 45 1532
rect -45 1470 45 1506
rect -45 1444 -39 1470
rect 39 1444 45 1470
rect -45 1408 45 1444
rect -45 1382 -39 1408
rect 39 1382 45 1408
rect -45 1346 45 1382
rect -45 1320 -39 1346
rect 39 1320 45 1346
rect -45 1284 45 1320
rect -45 1258 -39 1284
rect 39 1258 45 1284
rect -45 1222 45 1258
rect -45 1196 -39 1222
rect 39 1196 45 1222
rect -45 1160 45 1196
rect -45 1134 -39 1160
rect 39 1134 45 1160
rect -45 1098 45 1134
rect -45 1072 -39 1098
rect 39 1072 45 1098
rect -45 1036 45 1072
rect -45 1010 -39 1036
rect 39 1010 45 1036
rect -45 974 45 1010
rect -45 948 -39 974
rect 39 948 45 974
rect -45 912 45 948
rect -45 886 -39 912
rect 39 886 45 912
rect -45 850 45 886
rect -45 824 -39 850
rect 39 824 45 850
rect -45 788 45 824
rect -45 762 -39 788
rect 39 762 45 788
rect -45 726 45 762
rect -45 700 -39 726
rect 39 700 45 726
rect -45 664 45 700
rect -45 638 -39 664
rect 39 638 45 664
rect -45 602 45 638
rect -45 576 -39 602
rect 39 576 45 602
rect -45 540 45 576
rect -45 514 -39 540
rect 39 514 45 540
rect -45 478 45 514
rect -45 452 -39 478
rect 39 452 45 478
rect -45 416 45 452
rect -45 390 -39 416
rect 39 390 45 416
rect -45 354 45 390
rect -45 328 -39 354
rect 39 328 45 354
rect -45 292 45 328
rect -45 266 -39 292
rect 39 266 45 292
rect -45 230 45 266
rect -45 204 -39 230
rect 39 204 45 230
rect -45 168 45 204
rect -45 142 -39 168
rect 39 142 45 168
rect -45 106 45 142
rect -45 80 -39 106
rect 39 80 45 106
rect -45 44 45 80
rect -45 18 -39 44
rect 39 18 45 44
rect -45 -18 45 18
rect -45 -44 -39 -18
rect 39 -44 45 -18
rect -45 -80 45 -44
rect -45 -106 -39 -80
rect 39 -106 45 -80
rect -45 -142 45 -106
rect -45 -168 -39 -142
rect 39 -168 45 -142
rect -45 -204 45 -168
rect -45 -230 -39 -204
rect 39 -230 45 -204
rect -45 -266 45 -230
rect -45 -292 -39 -266
rect 39 -292 45 -266
rect -45 -328 45 -292
rect -45 -354 -39 -328
rect 39 -354 45 -328
rect -45 -390 45 -354
rect -45 -416 -39 -390
rect 39 -416 45 -390
rect -45 -452 45 -416
rect -45 -478 -39 -452
rect 39 -478 45 -452
rect -45 -514 45 -478
rect -45 -540 -39 -514
rect 39 -540 45 -514
rect -45 -576 45 -540
rect -45 -602 -39 -576
rect 39 -602 45 -576
rect -45 -638 45 -602
rect -45 -664 -39 -638
rect 39 -664 45 -638
rect -45 -700 45 -664
rect -45 -726 -39 -700
rect 39 -726 45 -700
rect -45 -762 45 -726
rect -45 -788 -39 -762
rect 39 -788 45 -762
rect -45 -824 45 -788
rect -45 -850 -39 -824
rect 39 -850 45 -824
rect -45 -886 45 -850
rect -45 -912 -39 -886
rect 39 -912 45 -886
rect -45 -948 45 -912
rect -45 -974 -39 -948
rect 39 -974 45 -948
rect -45 -1010 45 -974
rect -45 -1036 -39 -1010
rect 39 -1036 45 -1010
rect -45 -1072 45 -1036
rect -45 -1098 -39 -1072
rect 39 -1098 45 -1072
rect -45 -1134 45 -1098
rect -45 -1160 -39 -1134
rect 39 -1160 45 -1134
rect -45 -1196 45 -1160
rect -45 -1222 -39 -1196
rect 39 -1222 45 -1196
rect -45 -1258 45 -1222
rect -45 -1284 -39 -1258
rect 39 -1284 45 -1258
rect -45 -1320 45 -1284
rect -45 -1346 -39 -1320
rect 39 -1346 45 -1320
rect -45 -1382 45 -1346
rect -45 -1408 -39 -1382
rect 39 -1408 45 -1382
rect -45 -1444 45 -1408
rect -45 -1470 -39 -1444
rect 39 -1470 45 -1444
rect -45 -1506 45 -1470
rect -45 -1532 -39 -1506
rect 39 -1532 45 -1506
rect -45 -1568 45 -1532
rect -45 -1594 -39 -1568
rect 39 -1594 45 -1568
rect -45 -1630 45 -1594
rect -45 -1656 -39 -1630
rect 39 -1656 45 -1630
rect -45 -1692 45 -1656
rect -45 -1718 -39 -1692
rect 39 -1718 45 -1692
rect -45 -1754 45 -1718
rect -45 -1780 -39 -1754
rect 39 -1780 45 -1754
rect -45 -1816 45 -1780
rect -45 -1842 -39 -1816
rect 39 -1842 45 -1816
rect -45 -1878 45 -1842
rect -45 -1904 -39 -1878
rect 39 -1904 45 -1878
rect -45 -1940 45 -1904
rect -45 -1966 -39 -1940
rect 39 -1966 45 -1940
rect -45 -1972 45 -1966
<< end >>
