* NGSPICE file created from Transmission_Gate_Layout.ext - technology: gf180mcuC

.subckt pmos_3p3_METUKR a_n28_n930# a_n28_342# a_28_n886# a_n116_n886# w_n202_n1016#
+ a_n116_386# a_28_n250# a_28_386# a_n28_n294# a_n116_n250#
X0 a_28_386# a_n28_342# a_n116_386# w_n202_n1016# pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X1 a_28_n250# a_n28_n294# a_n116_n250# w_n202_n1016# pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X2 a_28_n886# a_n28_n930# a_n116_n886# w_n202_n1016# pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
.ends

.subckt nmos_3p3_Y4JRT2 a_n28_217# a_28_n511# a_28_n125# a_n28_n555# a_n28_n169# a_n116_n511#
+ a_n116_n125# a_n116_261# a_28_261# VSUBS
X0 a_28_n511# a_n28_n555# a_n116_n511# VSUBS nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X1 a_28_261# a_n28_217# a_n116_261# VSUBS nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X2 a_28_n125# a_n28_n169# a_n116_n125# VSUBS nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
.ends

.subckt nmos_3p3_RZHRT2 a_372_217# a_52_n555# a_428_261# a_108_n511# a_52_n169# a_588_261#
+ a_n676_261# a_108_n125# a_n532_n511# a_n108_n555# a_n532_n125# a_n108_n169# a_212_n555#
+ a_212_n169# a_268_n511# a_268_n125# a_n428_217# a_n212_261# a_n372_261# a_n588_217#
+ a_n268_n555# a_n268_n169# a_372_n555# a_372_n169# a_428_n511# a_428_n125# a_108_261#
+ a_532_217# a_268_261# a_n52_n511# a_52_217# a_n428_n555# a_n52_n125# a_n428_n169#
+ a_532_n555# a_588_n511# a_532_n169# a_588_n125# a_n212_n511# a_n108_217# a_n588_n555#
+ a_n212_n125# a_n588_n169# a_n268_217# a_n676_n511# a_n532_261# a_n676_n125# a_n372_n511#
+ a_n52_261# a_n372_n125# a_212_217# VSUBS
X0 a_108_261# a_52_217# a_n52_261# VSUBS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1 a_268_261# a_212_217# a_108_261# VSUBS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X2 a_588_n511# a_532_n555# a_428_n511# VSUBS nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X3 a_n372_261# a_n428_217# a_n532_261# VSUBS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X4 a_n532_n511# a_n588_n555# a_n676_n511# VSUBS nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X5 a_428_261# a_372_217# a_268_261# VSUBS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X6 a_n372_n511# a_n428_n555# a_n532_n511# VSUBS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X7 a_n532_261# a_n588_217# a_n676_261# VSUBS nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X8 a_588_n125# a_532_n169# a_428_n125# VSUBS nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X9 a_108_n511# a_52_n555# a_n52_n511# VSUBS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X10 a_428_n511# a_372_n555# a_268_n511# VSUBS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X11 a_268_n511# a_212_n555# a_108_n511# VSUBS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X12 a_n532_n125# a_n588_n169# a_n676_n125# VSUBS nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X13 a_n372_n125# a_n428_n169# a_n532_n125# VSUBS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X14 a_n212_n511# a_n268_n555# a_n372_n511# VSUBS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X15 a_n52_n511# a_n108_n555# a_n212_n511# VSUBS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X16 a_n52_261# a_n108_217# a_n212_261# VSUBS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X17 a_108_n125# a_52_n169# a_n52_n125# VSUBS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X18 a_428_n125# a_372_n169# a_268_n125# VSUBS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X19 a_588_261# a_532_217# a_428_261# VSUBS nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X20 a_268_n125# a_212_n169# a_108_n125# VSUBS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X21 a_n212_261# a_n268_217# a_n372_261# VSUBS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X22 a_n212_n125# a_n268_n169# a_n372_n125# VSUBS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X23 a_n52_n125# a_n108_n169# a_n212_n125# VSUBS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
.ends

.subckt pmos_3p3_M6SUKR a_108_n886# a_n428_n930# a_532_n930# a_n676_n250# a_n532_n886#
+ a_n372_n250# a_212_342# a_372_342# a_268_n886# a_n588_n930# a_108_n250# a_52_n294#
+ a_n212_386# a_n372_386# a_n532_n250# a_n108_n294# a_212_n294# a_428_n886# a_268_n250#
+ a_108_386# a_268_386# a_n428_342# a_52_n930# a_n588_342# a_n52_n886# a_n268_n294#
+ a_372_n294# a_588_n886# a_n108_n930# a_212_n930# w_n762_n1016# a_428_n250# a_532_342#
+ a_n212_n886# a_52_342# a_n52_n250# a_n428_n294# a_n532_386# a_n676_n886# a_n268_n930#
+ a_532_n294# a_372_n930# a_588_n250# a_n52_386# a_n372_n886# a_n108_342# a_n212_n250#
+ a_n588_n294# a_428_386# a_n676_386# a_n268_342# a_588_386#
X0 a_268_386# a_212_342# a_108_386# w_n762_n1016# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_n372_n886# a_n428_n930# a_n532_n886# w_n762_n1016# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_n372_386# a_n428_342# a_n532_386# w_n762_n1016# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X3 a_108_n886# a_52_n930# a_n52_n886# w_n762_n1016# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X4 a_428_n886# a_372_n930# a_268_n886# w_n762_n1016# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X5 a_428_386# a_372_342# a_268_386# w_n762_n1016# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X6 a_268_n886# a_212_n930# a_108_n886# w_n762_n1016# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X7 a_n532_386# a_n588_342# a_n676_386# w_n762_n1016# pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X8 a_588_n250# a_532_n294# a_428_n250# w_n762_n1016# pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X9 a_n212_n886# a_n268_n930# a_n372_n886# w_n762_n1016# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X10 a_n52_n886# a_n108_n930# a_n212_n886# w_n762_n1016# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X11 a_n532_n250# a_n588_n294# a_n676_n250# w_n762_n1016# pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X12 a_n372_n250# a_n428_n294# a_n532_n250# w_n762_n1016# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X13 a_n52_386# a_n108_342# a_n212_386# w_n762_n1016# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X14 a_108_n250# a_52_n294# a_n52_n250# w_n762_n1016# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X15 a_428_n250# a_372_n294# a_268_n250# w_n762_n1016# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X16 a_588_386# a_532_342# a_428_386# w_n762_n1016# pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X17 a_268_n250# a_212_n294# a_108_n250# w_n762_n1016# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X18 a_n212_386# a_n268_342# a_n372_386# w_n762_n1016# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X19 a_n212_n250# a_n268_n294# a_n372_n250# w_n762_n1016# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X20 a_n52_n250# a_n108_n294# a_n212_n250# w_n762_n1016# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X21 a_588_n886# a_532_n930# a_428_n886# w_n762_n1016# pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X22 a_108_386# a_52_342# a_n52_386# w_n762_n1016# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X23 a_n532_n886# a_n588_n930# a_n676_n886# w_n762_n1016# pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
.ends

.subckt Transmission_Gate_Layout VSS VDD CLK VIN VOUT
Xpmos_3p3_METUKR_0 CLK CLK a_n72_1206# VDD VDD VDD a_n72_1206# a_n72_1206# CLK VDD
+ pmos_3p3_METUKR
Xnmos_3p3_Y4JRT2_0 CLK a_n72_1206# a_n72_1206# CLK CLK VSS VSS VSS a_n72_1206# VSS
+ nmos_3p3_Y4JRT2
Xnmos_3p3_RZHRT2_0 CLK CLK VOUT VOUT CLK VIN VIN VOUT VOUT CLK VOUT CLK CLK CLK VIN
+ VIN CLK VOUT VIN CLK CLK CLK CLK CLK VOUT VOUT VOUT CLK VIN VIN CLK CLK VIN CLK
+ CLK VIN CLK VIN VOUT CLK CLK VOUT CLK CLK VIN VOUT VIN VIN VIN VIN CLK VSS nmos_3p3_RZHRT2
Xpmos_3p3_M6SUKR_1 VOUT a_n72_1206# a_n72_1206# VIN VOUT VIN a_n72_1206# a_n72_1206#
+ VIN a_n72_1206# VOUT a_n72_1206# VOUT VIN VOUT a_n72_1206# a_n72_1206# VOUT VIN
+ VOUT VIN a_n72_1206# a_n72_1206# a_n72_1206# VIN a_n72_1206# a_n72_1206# VIN a_n72_1206#
+ a_n72_1206# VDD VOUT a_n72_1206# VOUT a_n72_1206# VIN a_n72_1206# VOUT VIN a_n72_1206#
+ a_n72_1206# a_n72_1206# VIN VIN VIN a_n72_1206# VOUT a_n72_1206# VOUT VIN a_n72_1206#
+ VIN pmos_3p3_M6SUKR
.ends

