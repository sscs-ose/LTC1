magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2277 -2042 2277 2042
<< polysilicon >>
rect -277 23 277 42
rect -277 -23 -258 23
rect 258 -23 277 23
rect -277 -42 277 -23
<< polycontact >>
rect -258 -23 258 23
<< metal1 >>
rect -269 23 269 34
rect -269 -23 -258 23
rect 258 -23 269 23
rect -269 -34 269 -23
<< end >>
