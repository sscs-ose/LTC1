* NGSPICE file created from mux_2x1_ibr_flat.ext - technology: gf180mcuC

.subckt pex_mux_2x1_ibr VSS Sel OUT I0 I1 VDD
X0 nand2_ibr_2.OUT I0.t0 a_801_n344# VSS.t2 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1 nand2_ibr_1.IN2 Sel.t0 a_238_256# VSS.t8 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2 VDD I0.t1 nand2_ibr_2.OUT VDD.t5 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3 OUT nand2_ibr_1.IN2 VDD.t1 VDD.t0 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X4 a_801_n344# nand2_ibr_2.IN2 VSS.t5 VSS.t0 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X5 nand2_ibr_2.IN2 Sel.t1 VSS.t4 VSS.t3 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X6 nand2_ibr_2.OUT nand2_ibr_2.IN2 VDD.t9 VDD.t8 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X7 nand2_ibr_1.IN2 I1.t0 VDD.t16 VDD.t15 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X8 a_801_256# nand2_ibr_1.IN2 VSS.t1 VSS.t0 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X9 nand2_ibr_2.IN2 Sel.t2 VDD.t14 VDD.t13 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X10 VDD nand2_ibr_2.OUT OUT.t1 VDD.t2 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X11 a_238_256# I1.t1 VSS.t7 VSS.t6 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X12 VDD Sel.t3 nand2_ibr_1.IN2 VDD.t10 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X13 OUT nand2_ibr_2.OUT a_801_256# VSS.t2 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
R0 I0.n0 I0.t0 31.528
R1 I0.n0 I0.t1 15.3826
R2 I0.n1 I0.n0 8.74076
R3 I0 I0.n1 0.116779
R4 I0.n1 I0 0.00202542
R5 VSS.t8 VSS.t0 1483.3
R6 VSS.n3 VSS.t2 353.341
R7 VSS.t0 VSS.n3 235.561
R8 VSS.n5 VSS.t6 235.561
R9 VSS.n0 VSS.t4 9.34566
R10 VSS.n2 VSS.t1 7.19156
R11 VSS.n2 VSS.t5 7.19156
R12 VSS.n7 VSS.t7 7.19156
R13 VSS.t3 VSS.t8 3.68113
R14 VSS.n6 VSS.n4 3.37613
R15 VSS.n3 VSS 2.60269
R16 VSS VSS.n6 2.6005
R17 VSS.n6 VSS.n5 2.6005
R18 VSS.n4 VSS.n1 2.6005
R19 VSS.n4 VSS.t3 2.6005
R20 VSS.n2 VSS.n1 0.131017
R21 VSS VSS.n2 0.0595367
R22 VSS VSS.n7 0.0569474
R23 VSS VSS.n0 0.0340526
R24 VSS.n7 VSS 0.0158947
R25 VSS VSS.n0 0.00405263
R26 VSS.n1 VSS 0.000894737
R27 Sel.n1 Sel.t0 31.528
R28 Sel.n0 Sel.t2 25.7638
R29 Sel.n1 Sel.t3 15.3826
R30 Sel.n0 Sel.t1 13.2969
R31 Sel.n2 Sel.n1 7.62851
R32 Sel.n5 Sel 2.26841
R33 Sel.n6 Sel.n4 2.2505
R34 Sel.n3 Sel.n2 2.2324
R35 Sel.n6 Sel.n0 2.11815
R36 Sel.n2 Sel 0.107918
R37 Sel.n4 Sel.n3 0.0289694
R38 Sel.n6 Sel.n5 0.00235567
R39 Sel Sel.n4 0.00233673
R40 Sel Sel.n6 0.00142783
R41 VDD.t10 VDD.t0 763.259
R42 VDD.n5 VDD.t8 386.348
R43 VDD.n5 VDD.t13 362.409
R44 VDD.n6 VDD.n5 319.75
R45 VDD.n1 VDD.t2 193.183
R46 VDD.n11 VDD.t10 193.183
R47 VDD.n4 VDD.t5 193.183
R48 VDD.t0 VDD.n1 109.849
R49 VDD.n11 VDD.t15 109.849
R50 VDD.t8 VDD.n4 109.849
R51 VDD.n7 VDD 11.7877
R52 VDD.n4 VDD.n3 6.3005
R53 VDD.n15 VDD.n1 6.3005
R54 VDD.n12 VDD.n11 6.3005
R55 VDD VDD.n2 5.23855
R56 VDD VDD.n0 5.23855
R57 VDD.n12 VDD.t16 5.21701
R58 VDD.n6 VDD.t14 5.19258
R59 VDD.n13 VDD.n10 5.13287
R60 VDD.n9 VDD.t1 3.91303
R61 VDD.n9 VDD.n8 3.87523
R62 VDD.n8 VDD.t9 3.51093
R63 VDD.n8 VDD.n7 0.272927
R64 VDD.n14 VDD.n9 0.22389
R65 VDD.n13 VDD 0.106177
R66 VDD.n7 VDD.n3 0.0800484
R67 VDD.n15 VDD.n14 0.0800484
R68 VDD.n14 VDD 0.0713387
R69 VDD VDD.n13 0.0701774
R70 VDD.n3 VDD 0.00166129
R71 VDD VDD.n15 0.00166129
R72 VDD VDD.n12 0.00166129
R73 VDD VDD.n6 0.00105556
R74 OUT OUT.n3 7.15141
R75 OUT.n2 OUT.n1 3.2163
R76 OUT.n1 OUT.t1 2.2755
R77 OUT.n1 OUT.n0 2.2755
R78 OUT.n2 OUT 0.0574388
R79 OUT OUT.n2 0.0119545
R80 I1.n0 I1.t0 30.9379
R81 I1.n0 I1.t1 21.6422
R82 I1 I1.n0 4.005
C0 a_801_256# nand2_ibr_1.IN2 0.00372f
C1 a_801_256# VDD 0.00444f
C2 nand2_ibr_2.OUT nand2_ibr_1.IN2 0.053f
C3 nand2_ibr_2.OUT VDD 0.637f
C4 OUT Sel 0.00946f
C5 nand2_ibr_2.OUT a_801_n344# 0.0964f
C6 Sel nand2_ibr_2.IN2 0.136f
C7 I1 nand2_ibr_1.IN2 0.0959f
C8 I1 VDD 0.147f
C9 OUT I0 1.36e-19
C10 I0 nand2_ibr_2.IN2 0.0473f
C11 I1 a_238_256# 0.00347f
C12 a_801_256# OUT 0.069f
C13 nand2_ibr_2.OUT Sel 4.46e-19
C14 nand2_ibr_2.OUT OUT 0.303f
C15 nand2_ibr_2.OUT nand2_ibr_2.IN2 0.12f
C16 nand2_ibr_2.OUT I0 0.202f
C17 I1 Sel 0.055f
C18 VDD nand2_ibr_1.IN2 0.458f
C19 a_801_n344# VDD 0.00444f
C20 a_238_256# nand2_ibr_1.IN2 0.069f
C21 VDD a_238_256# 3.14e-19
C22 a_801_256# nand2_ibr_2.OUT 0.00949f
C23 Sel nand2_ibr_1.IN2 0.341f
C24 Sel VDD 0.588f
C25 OUT nand2_ibr_1.IN2 0.109f
C26 OUT VDD 0.234f
C27 Sel a_801_n344# 2.62e-19
C28 nand2_ibr_2.IN2 nand2_ibr_1.IN2 0.00212f
C29 VDD nand2_ibr_2.IN2 0.401f
C30 Sel a_238_256# 0.0144f
C31 I0 VDD 0.233f
C32 a_801_n344# nand2_ibr_2.IN2 0.00372f
C33 I0 a_801_n344# 0.00293f
C34 a_801_n344# VSS 0.0676f
C35 I0 VSS 0.256f
C36 nand2_ibr_2.IN2 VSS 0.436f
C37 a_801_256# VSS 0.0676f
C38 a_238_256# VSS 0.0678f
C39 OUT VSS 0.14f
C40 nand2_ibr_2.OUT VSS 0.659f
C41 nand2_ibr_1.IN2 VSS 0.435f
C42 Sel VSS 0.842f
C43 I1 VSS 0.292f
C44 VDD VSS 4.29f
.ends

