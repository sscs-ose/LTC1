magic
tech gf180mcuC
magscale 1 10
timestamp 1694088685
<< nwell >>
rect 2736 3570 2863 3599
rect 2736 3551 2873 3570
rect 2736 3479 2863 3551
rect 3331 3455 3339 3923
rect 3706 3480 3839 3576
rect 3326 3454 3339 3455
rect 4307 3454 4315 3923
rect 6388 3738 6391 3930
rect 5252 3737 5354 3738
rect 6388 3737 6389 3738
rect 5252 3686 5386 3737
rect 5283 3685 5386 3686
rect 5283 3454 5288 3685
rect 6339 3684 6394 3737
rect 6979 3700 7146 3931
rect 6384 3267 6393 3684
rect 7104 3463 7126 3700
rect 7113 3462 7118 3463
rect 6384 3265 6392 3267
<< metal1 >>
rect 3331 3817 3339 3923
rect 4307 3817 4314 3923
rect 5258 3630 5411 3922
rect 6330 3636 6491 3818
rect 6979 3700 7146 3931
rect 7508 3769 7854 3940
rect 2736 3535 2862 3540
rect 2736 3482 2748 3535
rect 2801 3482 2862 3535
rect 2736 3479 2862 3482
rect 3706 3537 3839 3540
rect 3706 3483 3724 3537
rect 3778 3483 3839 3537
rect 3706 3480 3839 3483
rect 4690 3535 4812 3537
rect 4690 3481 4701 3535
rect 4754 3481 4812 3535
rect 3727 3479 3794 3480
rect 4690 3479 4812 3481
rect 2478 3439 2567 3461
rect 2478 3380 2494 3439
rect 2557 3380 2567 3439
rect 2478 3372 2567 3380
rect 3416 3441 3543 3450
rect 4433 3442 4497 3443
rect 3416 3379 3450 3441
rect 3513 3379 3543 3441
rect 3416 3370 3543 3379
rect 4421 3438 4500 3442
rect 4421 3384 4434 3438
rect 4487 3384 4500 3438
rect 6995 3433 7202 3499
rect 4141 3365 4280 3376
rect 4421 3373 4500 3384
rect 3186 3355 3271 3362
rect 3186 3300 3198 3355
rect 3250 3300 3271 3355
rect 3186 3296 3271 3300
rect 4141 3301 4163 3365
rect 4227 3301 4280 3365
rect 4141 3288 4280 3301
rect -14 2870 2407 3041
rect 3273 2930 3372 3222
rect 4252 2932 4351 3224
rect 5242 3180 5341 3223
rect 5242 3038 5374 3180
rect 6234 3174 6300 3179
rect 6234 3120 6240 3174
rect 6292 3120 6300 3174
rect 6234 3107 6300 3120
rect 6540 3093 6618 3105
rect 6540 3040 6553 3093
rect 6607 3040 6618 3093
rect 5242 2931 5421 3038
rect -14 2464 157 2870
rect 6308 2593 6410 3037
rect 6540 3032 6618 3040
rect 6683 3095 6771 3104
rect 6683 3040 6706 3095
rect 6759 3040 6771 3095
rect 6683 3033 6771 3040
rect 6831 3094 6921 3105
rect 6831 3041 6854 3094
rect 6907 3041 6921 3094
rect 6831 3032 6921 3041
rect 7172 2712 7301 3206
rect 6963 2592 7301 2712
rect 7172 2591 7301 2592
rect -336 2293 157 2464
rect -336 1459 -165 2293
rect 2897 1989 3686 2150
rect 6163 1994 7178 2155
rect 7683 2069 7854 3769
rect 6164 1991 7013 1994
rect 6164 1990 6953 1991
rect 494 1607 607 1616
rect 493 1595 607 1607
rect 493 1538 512 1595
rect 569 1538 607 1595
rect 493 1537 607 1538
rect 3735 1596 3846 1608
rect 3735 1538 3751 1596
rect 3815 1538 3846 1596
rect 6655 1588 6792 1667
rect 7086 1620 7143 1935
rect 7079 1605 7200 1620
rect 493 1528 606 1537
rect 3735 1528 3846 1538
rect 7079 1541 7107 1605
rect 7171 1541 7200 1605
rect 7079 1535 7200 1541
rect 7086 1531 7143 1535
rect -336 1288 147 1459
rect 4711 611 4810 613
rect 1474 607 1567 609
rect 1474 551 1487 607
rect 1544 551 1567 607
rect 4711 555 4722 611
rect 4778 555 4810 611
rect 4711 553 4810 555
rect 8064 611 8160 614
rect 8064 557 8075 611
rect 8131 557 8160 611
rect 8064 553 8160 557
rect 1474 549 1567 551
rect 494 512 601 522
rect 494 450 523 512
rect 588 450 601 512
rect 494 439 601 450
rect 3727 519 3842 528
rect 3727 456 3752 519
rect 3810 456 3842 519
rect 3727 446 3842 456
rect 7048 516 7189 532
rect 7048 459 7102 516
rect 7164 459 7189 516
rect 7048 453 7189 459
rect 9529 478 9641 506
rect 9529 410 9551 478
rect 9620 410 9641 478
rect 9529 386 9641 410
rect 2865 11 3598 118
rect 6135 11 6868 118
<< via1 >>
rect 5141 3656 5193 3709
rect 2748 3482 2801 3535
rect 3724 3483 3778 3537
rect 4701 3481 4754 3535
rect 2494 3380 2557 3439
rect 3450 3379 3513 3441
rect 4434 3384 4487 3438
rect 3198 3300 3250 3355
rect 4163 3301 4227 3365
rect 5466 3235 5530 3299
rect 6240 3120 6292 3174
rect 6553 3040 6607 3093
rect 6706 3040 6759 3095
rect 6854 3041 6907 3094
rect 512 1538 569 1595
rect 3751 1538 3815 1596
rect 7107 1541 7171 1605
rect 1487 551 1544 607
rect 4722 555 4778 611
rect 8075 557 8131 611
rect 523 450 588 512
rect 3752 456 3810 519
rect 7102 459 7164 516
rect 9551 410 9620 478
<< metal2 >>
rect 2476 3734 4764 3823
rect 2476 3460 2565 3734
rect 2740 3623 3794 3630
rect 2740 3599 4500 3623
rect 2736 3562 4500 3599
rect 2736 3552 2873 3562
rect 2735 3551 2873 3552
rect 3706 3555 4500 3562
rect 2735 3535 2863 3551
rect 2735 3484 2748 3535
rect 2736 3482 2748 3484
rect 2801 3482 2863 3535
rect 2736 3479 2863 3482
rect 3706 3537 3839 3555
rect 3706 3483 3724 3537
rect 3778 3483 3839 3537
rect 3706 3480 3839 3483
rect 4432 3466 4500 3555
rect 4675 3546 4764 3734
rect 5123 3709 6940 3724
rect 5123 3656 5141 3709
rect 5193 3656 6940 3709
rect 5123 3641 6940 3656
rect 4675 3535 4768 3546
rect 4675 3481 4701 3535
rect 4754 3481 4768 3535
rect 4675 3475 4768 3481
rect 2448 3439 2585 3460
rect 3416 3444 3543 3450
rect 2448 3380 2494 3439
rect 2557 3380 2585 3439
rect 2448 3059 2585 3380
rect 3414 3441 3543 3444
rect 3414 3379 3450 3441
rect 3513 3379 3543 3441
rect 3414 3370 3543 3379
rect 4417 3438 4516 3466
rect 4417 3384 4434 3438
rect 4487 3384 4516 3438
rect 3186 3361 3271 3362
rect 3179 3355 3304 3361
rect 3179 3300 3198 3355
rect 3250 3300 3304 3355
rect 68 2100 2313 2129
rect 68 2025 2179 2100
rect 2259 2025 2313 2100
rect 68 2008 2313 2025
rect 68 1581 189 2008
rect 2451 1936 2582 3059
rect 3179 2423 3304 3300
rect 3179 2365 3203 2423
rect 3260 2365 3304 2423
rect 3179 2340 3304 2365
rect 3414 2137 3538 3370
rect 4141 3365 4280 3376
rect 4141 3301 4163 3365
rect 4227 3301 4280 3365
rect 4141 3288 4280 3301
rect 4149 3285 4280 3288
rect 3648 2430 4303 2458
rect 3648 2424 4184 2430
rect 3648 2366 3685 2424
rect 3742 2372 4184 2424
rect 4241 2372 4303 2430
rect 3742 2366 4303 2372
rect 3648 2333 4303 2366
rect 2704 2107 4313 2137
rect 2704 2032 2731 2107
rect 2811 2032 4210 2107
rect 4286 2032 4313 2107
rect 2704 2016 4313 2032
rect 2451 1805 3022 1936
rect 493 1595 606 1607
rect 493 1538 512 1595
rect 569 1538 606 1595
rect 2891 1593 3022 1805
rect 3324 1664 3425 2016
rect 4417 2013 4516 3384
rect 4702 3369 5321 3385
rect 4702 3305 4762 3369
rect 4826 3310 5321 3369
rect 4826 3305 5597 3310
rect 4702 3299 5597 3305
rect 4702 3293 5466 3299
rect 5234 3235 5466 3293
rect 5530 3235 5597 3299
rect 5234 3226 5597 3235
rect 6228 3174 6307 3179
rect 6228 3120 6240 3174
rect 6292 3120 6307 3174
rect 6228 3107 6307 3120
rect 6234 3104 6307 3107
rect 6502 3104 6618 3105
rect 6234 3093 6618 3104
rect 6234 3040 6553 3093
rect 6607 3040 6618 3093
rect 6234 3039 6618 3040
rect 6346 3038 6618 3039
rect 6540 3032 6618 3038
rect 6683 3095 6773 3109
rect 6857 3105 6940 3641
rect 6683 3040 6706 3095
rect 6759 3040 6773 3095
rect 4612 2416 6401 2451
rect 4612 2358 4654 2416
rect 4711 2358 6315 2416
rect 6372 2358 6401 2416
rect 6683 2374 6773 3040
rect 6831 3094 6940 3105
rect 6831 3041 6854 3094
rect 6907 3041 6940 3094
rect 6831 3032 6940 3041
rect 6857 3016 6940 3032
rect 4612 2326 6401 2358
rect 6679 2274 6975 2374
rect 4612 2172 6779 2204
rect 4612 2097 4631 2172
rect 4707 2097 6779 2172
rect 4612 2083 6779 2097
rect 4417 1914 6182 2013
rect 3357 1663 3425 1664
rect 6083 1630 6182 1914
rect 6004 1613 6182 1630
rect 3727 1596 3846 1608
rect 5996 1597 6182 1613
rect 3727 1593 3751 1596
rect 493 1528 606 1538
rect 2748 1498 3293 1593
rect 3198 1467 3293 1498
rect 3517 1538 3751 1593
rect 3815 1538 3846 1596
rect 3517 1498 3846 1538
rect 3517 1467 3612 1498
rect 3198 1372 3612 1467
rect 1468 608 1564 609
rect 1468 551 1482 608
rect 1539 607 1564 608
rect 1544 551 1564 607
rect 1468 549 1564 551
rect 503 522 600 525
rect 494 512 601 522
rect 494 450 523 512
rect 588 450 601 512
rect 494 439 601 450
rect 3727 519 3846 1498
rect 5963 1494 6182 1597
rect 5996 1493 6182 1494
rect 6281 1933 6406 1976
rect 6281 1875 6312 1933
rect 6369 1875 6406 1933
rect 4698 611 4797 613
rect 4698 555 4719 611
rect 4778 555 4797 611
rect 4698 553 4797 555
rect 6281 562 6406 1875
rect 6650 1588 6777 2083
rect 6875 2011 6975 2274
rect 6875 1911 9530 2011
rect 7079 1605 7200 1612
rect 7079 1541 7107 1605
rect 7171 1541 7200 1605
rect 9430 1600 9530 1911
rect 7079 1535 7200 1541
rect 9326 1500 9530 1600
rect 9326 1499 9398 1500
rect 3727 456 3752 519
rect 3810 456 3846 519
rect 3727 445 3846 456
rect 6281 516 7201 562
rect 8056 557 8072 613
rect 8128 611 8151 613
rect 8131 557 8151 611
rect 8056 552 8151 557
rect 6281 459 7102 516
rect 7164 459 7201 516
rect 9542 506 9637 514
rect 503 430 600 439
rect 6281 438 7201 459
rect 9529 478 9641 506
rect 503 152 598 430
rect 9529 410 9551 478
rect 9620 410 9641 478
rect 9529 386 9641 410
rect 9542 152 9637 386
rect 503 57 9637 152
<< via2 >>
rect 2179 2025 2259 2100
rect 3203 2365 3260 2423
rect 4163 3301 4227 3365
rect 3685 2366 3742 2424
rect 4184 2372 4241 2430
rect 2731 2032 2811 2107
rect 4210 2032 4286 2107
rect 512 1538 569 1595
rect 4762 3305 4826 3369
rect 4654 2358 4711 2416
rect 6315 2358 6372 2416
rect 4631 2097 4707 2172
rect 1482 607 1539 608
rect 1482 551 1487 607
rect 1487 551 1539 607
rect 6312 1875 6369 1933
rect 4719 555 4722 611
rect 4722 555 4775 611
rect 7107 1541 7171 1605
rect 8072 611 8128 613
rect 8072 557 8075 611
rect 8075 557 8128 611
<< metal3 >>
rect 4144 3369 4861 3380
rect 4144 3365 4762 3369
rect 4144 3301 4163 3365
rect 4227 3305 4762 3365
rect 4826 3305 4861 3369
rect 4227 3301 4861 3305
rect 4144 3288 4861 3301
rect 3178 2424 3784 2461
rect 3178 2423 3685 2424
rect 3178 2365 3203 2423
rect 3260 2366 3685 2423
rect 3742 2366 3784 2424
rect 3260 2365 3784 2366
rect 3178 2332 3784 2365
rect 4145 2430 4751 2456
rect 4145 2372 4184 2430
rect 4241 2416 4751 2430
rect 4241 2372 4654 2416
rect 4145 2358 4654 2372
rect 4711 2358 4751 2416
rect 4145 2327 4751 2358
rect 6279 2416 6413 2461
rect 6279 2358 6315 2416
rect 6372 2358 6413 2416
rect 4188 2172 4737 2204
rect 2302 2129 2830 2137
rect 2154 2107 2830 2129
rect 2154 2100 2731 2107
rect 2154 2025 2179 2100
rect 2259 2032 2731 2100
rect 2811 2032 2830 2107
rect 2259 2025 2830 2032
rect 2154 2009 2830 2025
rect 4188 2107 4631 2172
rect 4188 2032 4210 2107
rect 4286 2097 4631 2107
rect 4707 2097 4737 2172
rect 4286 2084 4737 2097
rect 4286 2032 4313 2084
rect 4188 2017 4313 2032
rect 2302 2008 2830 2009
rect 6279 1933 6413 2358
rect 6279 1875 6312 1933
rect 6369 1875 6413 1933
rect 6279 1827 6413 1875
rect 477 1595 641 1645
rect 477 1538 512 1595
rect 569 1538 641 1595
rect 477 978 641 1538
rect 7049 1605 7213 1638
rect 7049 1541 7107 1605
rect 7171 1541 7213 1605
rect 7049 978 7213 1541
rect 477 814 7213 978
rect 1448 613 8182 650
rect 1448 611 8072 613
rect 1448 608 4719 611
rect 1448 551 1482 608
rect 1539 555 4719 608
rect 4775 557 8072 611
rect 8128 557 8182 613
rect 4775 555 8182 557
rect 1539 551 8182 555
rect 1448 520 8182 551
use and2_mag  and2_mag_0
timestamp 1694088685
transform 1 0 2425 0 1 3119
box -70 -188 1009 863
use and2_mag  and2_mag_1
timestamp 1694088685
transform 1 0 3401 0 1 3119
box -70 -188 1009 863
use and2_mag  and2_mag_2
timestamp 1694088685
transform 1 0 4377 0 1 3119
box -70 -188 1009 863
use Buffer_delayed_mag  Buffer_delayed_mag_0
timestamp 1692973937
transform 1 0 5506 0 1 3106
box -218 -175 878 631
use GF_INV_MAG  GF_INV_MAG_0
timestamp 1694086208
transform 1 0 7235 0 1 3300
box -118 -175 286 631
use JK_FF_mag  JK_FF_mag_0
timestamp 1694088685
transform 1 0 390 0 1 0
box -390 0 2603 2148
use JK_FF_mag  JK_FF_mag_1
timestamp 1694088685
transform 1 0 3627 0 1 5
box -390 0 2603 2148
use JK_FF_mag  JK_FF_mag_2
timestamp 1694088685
transform 1 0 6980 0 1 5
box -390 0 2603 2148
use nor_3_mag  nor_3_mag_0
timestamp 1694086208
transform 1 0 6059 0 1 2152
box 329 440 1054 1778
<< labels >>
flabel via2 1517 576 1517 576 0 FreeSans 800 0 0 0 RST
port 0 nsew
flabel metal2 174 1621 174 1621 0 FreeSans 800 0 0 0 CLK
port 1 nsew
flabel metal1 3281 25 3281 25 0 FreeSans 800 0 0 0 VSS
port 2 nsew
flabel metal1 7762 2582 7762 2582 0 FreeSans 800 0 0 0 VDD
port 3 nsew
flabel via1 2784 3509 2784 3509 0 FreeSans 800 0 0 0 Q1
port 6 nsew
flabel via1 2528 3416 2528 3416 0 FreeSans 800 0 0 0 Q0
port 7 nsew
flabel via1 6739 3067 6739 3067 0 FreeSans 800 0 0 0 Q2
port 8 nsew
<< end >>
