magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect 11097 11097 73000 73000
<< metal4 >>
rect 14000 47020 17000 71000
rect 17200 48366 20200 71000
rect 20400 49774 23400 71000
rect 23600 50362 25000 71000
rect 25200 51120 26600 71000
rect 26800 52360 29800 71000
rect 30000 53704 33000 71000
rect 33200 55027 36200 71000
rect 36400 56465 39400 71000
rect 39600 57132 41000 71000
rect 41200 57810 42600 71000
rect 42800 59044 45800 71000
rect 46000 60708 49000 71000
rect 49200 61091 50600 71000
rect 50800 61751 52200 71000
rect 52400 62421 53800 71000
rect 54000 63320 55400 71000
rect 55600 63753 57000 71000
rect 57200 64540 58600 71000
rect 58800 65081 60200 71000
rect 60400 65760 61800 71000
rect 62000 66402 63400 71000
rect 63600 67263 65000 71000
rect 65200 67745 66600 71000
rect 66800 68493 68200 71000
rect 68400 69678 69678 71000
rect 68400 68769 71000 69678
tri 68400 68693 68476 68769 ne
rect 68476 68693 71000 68769
tri 68200 68493 68400 68693 sw
tri 68476 68493 68676 68693 ne
rect 68676 68493 71000 68693
rect 66800 68400 68400 68493
tri 68400 68400 68493 68493 sw
tri 68676 68400 68769 68493 ne
rect 68769 68400 71000 68493
rect 66800 68200 68493 68400
tri 68493 68200 68693 68400 sw
rect 66800 68113 71000 68200
tri 66800 68029 66884 68113 ne
rect 66884 68029 71000 68113
tri 66600 67745 66884 68029 sw
tri 66884 67745 67168 68029 ne
rect 67168 67745 71000 68029
rect 65200 67461 66884 67745
tri 66884 67461 67168 67745 sw
tri 67168 67461 67452 67745 ne
rect 67452 67461 71000 67745
rect 65200 67452 67168 67461
tri 67168 67452 67177 67461 sw
tri 67452 67452 67461 67461 ne
rect 67461 67452 71000 67461
rect 65200 67449 67177 67452
tri 65200 67366 65283 67449 ne
rect 65283 67366 67177 67449
tri 65000 67263 65103 67366 sw
tri 65283 67263 65386 67366 ne
rect 65386 67263 67177 67366
rect 63600 66980 65103 67263
tri 65103 66980 65386 67263 sw
tri 65386 66980 65669 67263 ne
rect 65669 67168 67177 67263
tri 67177 67168 67461 67452 sw
tri 67461 67168 67745 67452 ne
rect 67745 67168 71000 67452
rect 65669 66980 67461 67168
rect 63600 66786 65386 66980
tri 63600 66694 63692 66786 ne
rect 63692 66697 65386 66786
tri 65386 66697 65669 66980 sw
tri 65669 66697 65952 66980 ne
rect 65952 66884 67461 66980
tri 67461 66884 67745 67168 sw
tri 67745 66884 68029 67168 ne
rect 68029 66884 71000 67168
rect 65952 66697 67745 66884
rect 63692 66694 65669 66697
tri 63400 66402 63692 66694 sw
tri 63692 66402 63984 66694 ne
rect 63984 66414 65669 66694
tri 65669 66414 65952 66697 sw
tri 65952 66414 66235 66697 ne
rect 66235 66600 67745 66697
tri 67745 66600 68029 66884 sw
tri 68029 66800 68113 66884 ne
rect 68113 66800 71000 66884
rect 66235 66414 71000 66600
rect 63984 66402 65952 66414
rect 62000 66114 63692 66402
tri 62000 66031 62083 66114 ne
rect 62083 66110 63692 66114
tri 63692 66110 63984 66402 sw
tri 63984 66110 64276 66402 ne
rect 64276 66332 65952 66402
tri 65952 66332 66034 66414 sw
tri 66235 66332 66317 66414 ne
rect 66317 66332 71000 66414
rect 64276 66110 66034 66332
rect 62083 66031 63984 66110
tri 61800 65760 62071 66031 sw
tri 62083 65760 62354 66031 ne
rect 62354 65964 63984 66031
tri 63984 65964 64130 66110 sw
tri 64276 65964 64422 66110 ne
rect 64422 66049 66034 66110
tri 66034 66049 66317 66332 sw
tri 66317 66049 66600 66332 ne
rect 66600 66049 71000 66332
rect 64422 65964 66317 66049
rect 62354 65760 64130 65964
rect 60400 65477 62071 65760
tri 62071 65477 62354 65760 sw
tri 62354 65477 62637 65760 ne
rect 62637 65672 64130 65760
tri 64130 65672 64422 65964 sw
tri 64422 65672 64714 65964 ne
rect 64714 65766 66317 65964
tri 66317 65766 66600 66049 sw
tri 66600 65766 66883 66049 ne
rect 66883 65766 71000 66049
rect 64714 65672 66600 65766
rect 62637 65477 64422 65672
rect 60400 65451 62354 65477
tri 60400 65366 60485 65451 ne
rect 60485 65366 62354 65451
tri 60200 65081 60485 65366 sw
tri 60485 65081 60770 65366 ne
rect 60770 65194 62354 65366
tri 62354 65194 62637 65477 sw
tri 62637 65194 62920 65477 ne
rect 62920 65380 64422 65477
tri 64422 65380 64714 65672 sw
tri 64714 65380 65006 65672 ne
rect 65006 65566 66600 65672
tri 66600 65566 66800 65766 sw
tri 66883 65566 67083 65766 ne
rect 67083 65566 71000 65766
rect 65006 65380 66800 65566
rect 62920 65194 64714 65380
rect 60770 65081 62637 65194
rect 58800 64796 60485 65081
tri 60485 64796 60770 65081 sw
tri 60770 64796 61055 65081 ne
rect 61055 64997 62637 65081
tri 62637 64997 62834 65194 sw
tri 62920 64997 63117 65194 ne
rect 63117 65088 64714 65194
tri 64714 65088 65006 65380 sw
tri 65006 65088 65298 65380 ne
rect 65298 65283 66800 65380
tri 66800 65283 67083 65566 sw
tri 67083 65283 67366 65566 ne
rect 67366 65283 71000 65566
rect 65298 65088 67083 65283
rect 63117 65000 65006 65088
tri 65006 65000 65094 65088 sw
tri 65298 65000 65386 65088 ne
rect 65386 65000 67083 65088
tri 67083 65000 67366 65283 sw
tri 67366 65200 67449 65283 ne
rect 67449 65200 71000 65283
rect 63117 64997 65094 65000
rect 61055 64796 62834 64997
rect 58800 64786 60770 64796
tri 58800 64699 58887 64786 ne
rect 58887 64730 60770 64786
tri 60770 64730 60836 64796 sw
tri 61055 64730 61121 64796 ne
rect 61121 64730 62834 64796
rect 58887 64699 60836 64730
tri 58600 64540 58759 64699 sw
tri 58887 64540 59046 64699 ne
rect 59046 64540 60836 64699
rect 57200 64253 58759 64540
tri 58759 64253 59046 64540 sw
tri 59046 64253 59333 64540 ne
rect 59333 64445 60836 64540
tri 60836 64445 61121 64730 sw
tri 61121 64445 61406 64730 ne
rect 61406 64714 62834 64730
tri 62834 64714 63117 64997 sw
tri 63117 64714 63400 64997 ne
rect 63400 64714 65094 64997
rect 61406 64445 63117 64714
rect 59333 64253 61121 64445
rect 57200 64119 59046 64253
tri 57200 64036 57283 64119 ne
rect 57283 64036 59046 64119
tri 57000 63753 57283 64036 sw
tri 57283 63753 57566 64036 ne
rect 57566 63966 59046 64036
tri 59046 63966 59333 64253 sw
tri 59333 63966 59620 64253 ne
rect 59620 64160 61121 64253
tri 61121 64160 61406 64445 sw
tri 61406 64160 61691 64445 ne
rect 61691 64431 63117 64445
tri 63117 64431 63400 64714 sw
tri 63400 64431 63683 64714 ne
rect 63683 64708 65094 64714
tri 65094 64708 65386 65000 sw
tri 65386 64708 65678 65000 ne
rect 65678 64708 71000 65000
rect 63683 64431 65386 64708
rect 61691 64346 63400 64431
tri 63400 64346 63485 64431 sw
tri 63683 64346 63768 64431 ne
rect 63768 64416 65386 64431
tri 65386 64416 65678 64708 sw
tri 65678 64416 65970 64708 ne
rect 65970 64416 71000 64708
rect 63768 64346 65678 64416
rect 61691 64160 63485 64346
rect 59620 63966 61406 64160
rect 57566 63960 59333 63966
tri 59333 63960 59339 63966 sw
tri 59620 63960 59626 63966 ne
rect 59626 63960 61406 63966
rect 57566 63753 59339 63960
rect 55600 63506 57283 63753
tri 57283 63506 57530 63753 sw
tri 57566 63506 57813 63753 ne
rect 57813 63673 59339 63753
tri 59339 63673 59626 63960 sw
tri 59626 63673 59913 63960 ne
rect 59913 63875 61406 63960
tri 61406 63875 61691 64160 sw
tri 61691 63875 61976 64160 ne
rect 61976 64063 63485 64160
tri 63485 64063 63768 64346 sw
tri 63768 64063 64051 64346 ne
rect 64051 64276 65678 64346
tri 65678 64276 65818 64416 sw
tri 65970 64276 66110 64416 ne
rect 66110 64276 71000 64416
rect 64051 64063 65818 64276
rect 61976 63875 63768 64063
rect 59913 63780 61691 63875
tri 61691 63780 61786 63875 sw
tri 61976 63780 62071 63875 ne
rect 62071 63780 63768 63875
tri 63768 63780 64051 64063 sw
tri 64051 63780 64334 64063 ne
rect 64334 63984 65818 64063
tri 65818 63984 66110 64276 sw
tri 66110 63984 66402 64276 ne
rect 66402 63984 71000 64276
rect 64334 63780 66110 63984
rect 59913 63673 61786 63780
rect 57813 63506 59626 63673
rect 55600 63456 57530 63506
tri 55600 63373 55683 63456 ne
rect 55683 63373 57530 63456
tri 55400 63320 55453 63373 sw
tri 55683 63320 55736 63373 ne
rect 55736 63320 57530 63373
rect 54000 63037 55453 63320
tri 55453 63037 55736 63320 sw
tri 55736 63037 56019 63320 ne
rect 56019 63223 57530 63320
tri 57530 63223 57813 63506 sw
tri 57813 63223 58096 63506 ne
rect 58096 63386 59626 63506
tri 59626 63386 59913 63673 sw
tri 59913 63386 60200 63673 ne
rect 60200 63495 61786 63673
tri 61786 63495 62071 63780 sw
tri 62071 63495 62356 63780 ne
rect 62356 63497 64051 63780
tri 64051 63497 64334 63780 sw
tri 64334 63497 64617 63780 ne
rect 64617 63692 66110 63780
tri 66110 63692 66402 63984 sw
tri 66402 63692 66694 63984 ne
rect 66694 63692 71000 63984
rect 64617 63497 66402 63692
rect 62356 63495 64334 63497
rect 60200 63386 62071 63495
rect 58096 63223 59913 63386
rect 56019 63037 57813 63223
rect 54000 62793 55736 63037
tri 54000 62707 54086 62793 ne
rect 54086 62754 55736 62793
tri 55736 62754 56019 63037 sw
tri 56019 62754 56302 63037 ne
rect 56302 62940 57813 63037
tri 57813 62940 58096 63223 sw
tri 58096 62940 58379 63223 ne
rect 58379 63099 59913 63223
tri 59913 63099 60200 63386 sw
tri 60200 63099 60487 63386 ne
rect 60487 63210 62071 63386
tri 62071 63210 62356 63495 sw
tri 62356 63210 62641 63495 ne
rect 62641 63400 64334 63495
tri 64334 63400 64431 63497 sw
tri 64617 63400 64714 63497 ne
rect 64714 63400 66402 63497
tri 66402 63400 66694 63692 sw
tri 66694 63600 66786 63692 ne
rect 66786 63600 71000 63692
rect 62641 63210 64431 63400
rect 60487 63099 62356 63210
rect 58379 62940 60200 63099
rect 56302 62754 58096 62940
rect 54086 62707 56019 62754
tri 53800 62421 54086 62707 sw
tri 54086 62421 54372 62707 ne
rect 54372 62622 56019 62707
tri 56019 62622 56151 62754 sw
tri 56302 62622 56434 62754 ne
rect 56434 62657 58096 62754
tri 58096 62657 58379 62940 sw
tri 58379 62657 58662 62940 ne
rect 58662 62847 60200 62940
tri 60200 62847 60452 63099 sw
tri 60487 62847 60739 63099 ne
rect 60739 63035 62356 63099
tri 62356 63035 62531 63210 sw
tri 62641 63035 62816 63210 ne
rect 62816 63117 64431 63210
tri 64431 63117 64714 63400 sw
tri 64714 63117 64997 63400 ne
rect 64997 63117 71000 63400
rect 62816 63035 64714 63117
rect 60739 62847 62531 63035
rect 58662 62657 60452 62847
rect 56434 62622 58379 62657
rect 54372 62421 56151 62622
rect 52400 62292 54086 62421
tri 54086 62292 54215 62421 sw
tri 54372 62292 54501 62421 ne
rect 54501 62339 56151 62421
tri 56151 62339 56434 62622 sw
tri 56434 62339 56717 62622 ne
rect 56717 62560 58379 62622
tri 58379 62560 58476 62657 sw
tri 58662 62560 58759 62657 ne
rect 58759 62560 60452 62657
tri 60452 62560 60739 62847 sw
tri 60739 62560 61026 62847 ne
rect 61026 62750 62531 62847
tri 62531 62750 62816 63035 sw
tri 62816 62750 63101 63035 ne
rect 63101 62834 64714 63035
tri 64714 62834 64997 63117 sw
tri 64997 62834 65280 63117 ne
rect 65280 62834 71000 63117
rect 63101 62750 64997 62834
rect 61026 62560 62816 62750
rect 56717 62339 58476 62560
rect 54501 62292 56434 62339
rect 52400 62127 54215 62292
tri 52400 62039 52488 62127 ne
rect 52488 62039 54215 62127
tri 52200 61751 52488 62039 sw
tri 52488 61751 52776 62039 ne
rect 52776 62006 54215 62039
tri 54215 62006 54501 62292 sw
tri 54501 62006 54787 62292 ne
rect 54787 62056 56434 62292
tri 56434 62056 56717 62339 sw
tri 56717 62056 57000 62339 ne
rect 57000 62277 58476 62339
tri 58476 62277 58759 62560 sw
tri 58759 62277 59042 62560 ne
rect 59042 62277 60739 62560
rect 57000 62056 58759 62277
rect 54787 62006 56717 62056
rect 52776 61751 54501 62006
rect 50800 61463 52488 61751
tri 52488 61463 52776 61751 sw
tri 52776 61463 53064 61751 ne
rect 53064 61720 54501 61751
tri 54501 61720 54787 62006 sw
tri 54787 61720 55073 62006 ne
rect 55073 61773 56717 62006
tri 56717 61773 57000 62056 sw
tri 57000 61773 57283 62056 ne
rect 57283 61994 58759 62056
tri 58759 61994 59042 62277 sw
tri 59042 61994 59325 62277 ne
rect 59325 62273 60739 62277
tri 60739 62273 61026 62560 sw
tri 61026 62273 61313 62560 ne
rect 61313 62465 62816 62560
tri 62816 62465 63101 62750 sw
tri 63101 62465 63386 62750 ne
rect 63386 62649 64997 62750
tri 64997 62649 65182 62834 sw
tri 65280 62649 65465 62834 ne
rect 65465 62649 71000 62834
rect 63386 62465 65182 62649
rect 61313 62273 63101 62465
rect 59325 62180 61026 62273
tri 61026 62180 61119 62273 sw
tri 61313 62180 61406 62273 ne
rect 61406 62180 63101 62273
tri 63101 62180 63386 62465 sw
tri 63386 62180 63671 62465 ne
rect 63671 62366 65182 62465
tri 65182 62366 65465 62649 sw
tri 65465 62366 65748 62649 ne
rect 65748 62366 71000 62649
rect 63671 62180 65465 62366
rect 59325 61994 61119 62180
rect 57283 61809 59042 61994
tri 59042 61809 59227 61994 sw
tri 59325 61809 59510 61994 ne
rect 59510 61893 61119 61994
tri 61119 61893 61406 62180 sw
tri 61406 61893 61693 62180 ne
rect 61693 61895 63386 62180
tri 63386 61895 63671 62180 sw
tri 63671 61895 63956 62180 ne
rect 63956 62083 65465 62180
tri 65465 62083 65748 62366 sw
tri 65748 62083 66031 62366 ne
rect 66031 62083 71000 62366
rect 63956 61895 65748 62083
rect 61693 61893 63671 61895
rect 59510 61809 61406 61893
rect 57283 61773 59227 61809
rect 55073 61720 57000 61773
rect 53064 61463 54787 61720
rect 50800 61459 52776 61463
tri 50800 61375 50884 61459 ne
rect 50884 61375 52776 61459
tri 50600 61091 50884 61375 sw
tri 50884 61091 51168 61375 ne
rect 51168 61303 52776 61375
tri 52776 61303 52936 61463 sw
tri 53064 61303 53224 61463 ne
rect 53224 61434 54787 61463
tri 54787 61434 55073 61720 sw
tri 55073 61434 55359 61720 ne
rect 55359 61623 57000 61720
tri 57000 61623 57150 61773 sw
tri 57283 61623 57433 61773 ne
rect 57433 61623 59227 61773
rect 55359 61434 57150 61623
rect 53224 61340 55073 61434
tri 55073 61340 55167 61434 sw
tri 55359 61340 55453 61434 ne
rect 55453 61340 57150 61434
tri 57150 61340 57433 61623 sw
tri 57433 61340 57716 61623 ne
rect 57716 61526 59227 61623
tri 59227 61526 59510 61809 sw
tri 59510 61526 59793 61809 ne
rect 59793 61606 61406 61809
tri 61406 61606 61693 61893 sw
tri 61693 61606 61980 61893 ne
rect 61980 61800 63671 61893
tri 63671 61800 63766 61895 sw
tri 63956 61800 64051 61895 ne
rect 64051 61800 65748 61895
tri 65748 61800 66031 62083 sw
tri 66031 62000 66114 62083 ne
rect 66114 62000 71000 62083
rect 61980 61606 63766 61800
rect 59793 61526 61693 61606
rect 57716 61340 59510 61526
rect 53224 61303 55167 61340
rect 51168 61091 52936 61303
rect 49200 61068 50884 61091
tri 50884 61068 50907 61091 sw
tri 51168 61068 51191 61091 ne
rect 51191 61068 52936 61091
rect 49200 60795 50907 61068
tri 49200 60710 49285 60795 ne
rect 49285 60784 50907 60795
tri 50907 60784 51191 61068 sw
tri 51191 60784 51475 61068 ne
rect 51475 61015 52936 61068
tri 52936 61015 53224 61303 sw
tri 53224 61015 53512 61303 ne
rect 53512 61054 55167 61303
tri 55167 61054 55453 61340 sw
tri 55453 61054 55739 61340 ne
rect 55739 61057 57433 61340
tri 57433 61057 57716 61340 sw
tri 57716 61057 57999 61340 ne
rect 57999 61243 59510 61340
tri 59510 61243 59793 61526 sw
tri 59793 61243 60076 61526 ne
rect 60076 61441 61693 61526
tri 61693 61441 61858 61606 sw
tri 61980 61441 62145 61606 ne
rect 62145 61515 63766 61606
tri 63766 61515 64051 61800 sw
tri 64051 61515 64336 61800 ne
rect 64336 61515 71000 61800
rect 62145 61441 64051 61515
rect 60076 61243 61858 61441
rect 57999 61057 59793 61243
rect 55739 61054 57716 61057
rect 53512 61015 55453 61054
rect 51475 60784 53224 61015
rect 49285 60710 51191 60784
tri 49000 60708 49002 60710 sw
tri 49285 60708 49287 60710 ne
rect 49287 60708 51191 60710
rect 46000 60423 49002 60708
tri 49002 60423 49287 60708 sw
tri 49287 60423 49572 60708 ne
rect 49572 60500 51191 60708
tri 51191 60500 51475 60784 sw
tri 51475 60500 51759 60784 ne
rect 51759 60727 53224 60784
tri 53224 60727 53512 61015 sw
tri 53512 60727 53800 61015 ne
rect 53800 60768 55453 61015
tri 55453 60768 55739 61054 sw
tri 55739 60768 56025 61054 ne
rect 56025 60960 57716 61054
tri 57716 60960 57813 61057 sw
tri 57999 60960 58096 61057 ne
rect 58096 60960 59793 61057
tri 59793 60960 60076 61243 sw
tri 60076 60960 60359 61243 ne
rect 60359 61154 61858 61243
tri 61858 61154 62145 61441 sw
tri 62145 61154 62432 61441 ne
rect 62432 61230 64051 61441
tri 64051 61230 64336 61515 sw
tri 64336 61230 64621 61515 ne
rect 64621 61230 71000 61515
rect 62432 61154 64336 61230
rect 60359 60960 62145 61154
rect 56025 60768 57813 60960
rect 53800 60727 55739 60768
rect 51759 60500 53512 60727
rect 49572 60423 51475 60500
rect 46000 60138 49287 60423
tri 49287 60138 49572 60423 sw
tri 49572 60138 49857 60423 ne
rect 49857 60216 51475 60423
tri 51475 60216 51759 60500 sw
tri 51759 60216 52043 60500 ne
rect 52043 60439 53512 60500
tri 53512 60439 53800 60727 sw
tri 53800 60439 54088 60727 ne
rect 54088 60598 55739 60727
tri 55739 60598 55909 60768 sw
tri 56025 60598 56195 60768 ne
rect 56195 60677 57813 60768
tri 57813 60677 58096 60960 sw
tri 58096 60677 58379 60960 ne
rect 58379 60677 60076 60960
tri 60076 60677 60359 60960 sw
tri 60359 60677 60642 60960 ne
rect 60642 60867 62145 60960
tri 62145 60867 62432 61154 sw
tri 62432 60867 62719 61154 ne
rect 62719 61055 64336 61154
tri 64336 61055 64511 61230 sw
tri 64621 61055 64796 61230 ne
rect 64796 61055 71000 61230
rect 62719 60867 64511 61055
rect 60642 60677 62432 60867
rect 56195 60598 58096 60677
rect 54088 60439 55909 60598
rect 52043 60408 53800 60439
tri 53800 60408 53831 60439 sw
tri 54088 60408 54119 60439 ne
rect 54119 60408 55909 60439
rect 52043 60216 53831 60408
rect 49857 60138 51759 60216
rect 46000 59853 49572 60138
tri 49572 59853 49857 60138 sw
tri 49857 59853 50142 60138 ne
rect 50142 60059 51759 60138
tri 51759 60059 51916 60216 sw
tri 52043 60059 52200 60216 ne
rect 52200 60120 53831 60216
tri 53831 60120 54119 60408 sw
tri 54119 60120 54407 60408 ne
rect 54407 60312 55909 60408
tri 55909 60312 56195 60598 sw
tri 56195 60312 56481 60598 ne
rect 56481 60394 58096 60598
tri 58096 60394 58379 60677 sw
tri 58379 60394 58662 60677 ne
rect 58662 60580 60359 60677
tri 60359 60580 60456 60677 sw
tri 60642 60580 60739 60677 ne
rect 60739 60580 62432 60677
tri 62432 60580 62719 60867 sw
tri 62719 60580 63006 60867 ne
rect 63006 60770 64511 60867
tri 64511 60770 64796 61055 sw
tri 64796 60770 65081 61055 ne
rect 65081 60770 71000 61055
rect 63006 60580 64796 60770
rect 58662 60394 60456 60580
rect 56481 60312 58379 60394
rect 54407 60120 56195 60312
rect 52200 60059 54119 60120
rect 50142 59853 51916 60059
rect 46000 59683 49857 59853
tri 49857 59683 50027 59853 sw
tri 50142 59683 50312 59853 ne
rect 50312 59775 51916 59853
tri 51916 59775 52200 60059 sw
tri 52200 59775 52484 60059 ne
rect 52484 59832 54119 60059
tri 54119 59832 54407 60120 sw
tri 54407 59832 54695 60120 ne
rect 54695 60026 56195 60120
tri 56195 60026 56481 60312 sw
tri 56481 60026 56767 60312 ne
rect 56767 60209 58379 60312
tri 58379 60209 58564 60394 sw
tri 58662 60209 58847 60394 ne
rect 58847 60297 60456 60394
tri 60456 60297 60739 60580 sw
tri 60739 60297 61022 60580 ne
rect 61022 60297 62719 60580
rect 58847 60209 60739 60297
rect 56767 60026 58564 60209
rect 54695 59832 56481 60026
rect 52484 59775 54407 59832
rect 50312 59683 52200 59775
rect 46000 59461 50027 59683
tri 46000 59350 46111 59461 ne
rect 46111 59398 50027 59461
tri 50027 59398 50312 59683 sw
tri 50312 59398 50597 59683 ne
rect 50597 59491 52200 59683
tri 52200 59491 52484 59775 sw
tri 52484 59491 52768 59775 ne
rect 52768 59740 54407 59775
tri 54407 59740 54499 59832 sw
tri 54695 59740 54787 59832 ne
rect 54787 59740 56481 59832
tri 56481 59740 56767 60026 sw
tri 56767 59740 57053 60026 ne
rect 57053 59926 58564 60026
tri 58564 59926 58847 60209 sw
tri 58847 59926 59130 60209 ne
rect 59130 60014 60739 60209
tri 60739 60014 61022 60297 sw
tri 61022 60014 61305 60297 ne
rect 61305 60293 62719 60297
tri 62719 60293 63006 60580 sw
tri 63006 60293 63293 60580 ne
rect 63293 60485 64796 60580
tri 64796 60485 65081 60770 sw
tri 65081 60485 65366 60770 ne
rect 65366 60485 71000 60770
rect 63293 60293 65081 60485
rect 61305 60200 63006 60293
tri 63006 60200 63099 60293 sw
tri 63293 60200 63386 60293 ne
rect 63386 60200 65081 60293
tri 65081 60200 65366 60485 sw
tri 65366 60400 65451 60485 ne
rect 65451 60400 71000 60485
rect 61305 60014 63099 60200
rect 59130 59926 61022 60014
rect 57053 59740 58847 59926
rect 52768 59491 54499 59740
rect 50597 59398 52484 59491
rect 46111 59397 50312 59398
tri 50312 59397 50313 59398 sw
tri 50597 59397 50598 59398 ne
rect 50598 59397 52484 59398
rect 46111 59350 50313 59397
tri 45800 59044 46106 59350 sw
tri 46111 59044 46417 59350 ne
rect 46417 59112 50313 59350
tri 50313 59112 50598 59397 sw
tri 50598 59112 50883 59397 ne
rect 50883 59372 52484 59397
tri 52484 59372 52603 59491 sw
tri 52768 59372 52887 59491 ne
rect 52887 59452 54499 59491
tri 54499 59452 54787 59740 sw
tri 54787 59452 55075 59740 ne
rect 55075 59454 56767 59740
tri 56767 59454 57053 59740 sw
tri 57053 59454 57339 59740 ne
rect 57339 59643 58847 59740
tri 58847 59643 59130 59926 sw
tri 59130 59643 59413 59926 ne
rect 59413 59829 61022 59926
tri 61022 59829 61207 60014 sw
tri 61305 59829 61490 60014 ne
rect 61490 59913 63099 60014
tri 63099 59913 63386 60200 sw
tri 63386 59913 63673 60200 ne
rect 63673 59913 71000 60200
rect 61490 59829 63386 59913
rect 59413 59643 61207 59829
rect 57339 59454 59130 59643
rect 55075 59452 57053 59454
rect 52887 59372 54787 59452
rect 50883 59112 52603 59372
rect 46417 59110 50598 59112
tri 50598 59110 50600 59112 sw
tri 50883 59110 50885 59112 ne
rect 50885 59110 52603 59112
rect 46417 59044 50600 59110
rect 42800 58834 46106 59044
tri 46106 58834 46316 59044 sw
tri 46417 58834 46627 59044 ne
rect 46627 58834 50600 59044
rect 42800 58551 46316 58834
tri 46316 58551 46599 58834 sw
tri 46627 58551 46910 58834 ne
rect 46910 58825 50600 58834
tri 50600 58825 50885 59110 sw
tri 50885 58825 51170 59110 ne
rect 51170 59088 52603 59110
tri 52603 59088 52887 59372 sw
tri 52887 59088 53171 59372 ne
rect 53171 59164 54787 59372
tri 54787 59164 55075 59452 sw
tri 55075 59164 55363 59452 ne
rect 55363 59360 57053 59452
tri 57053 59360 57147 59454 sw
tri 57339 59360 57433 59454 ne
rect 57433 59360 59130 59454
tri 59130 59360 59413 59643 sw
tri 59413 59360 59696 59643 ne
rect 59696 59546 61207 59643
tri 61207 59546 61490 59829 sw
tri 61490 59546 61773 59829 ne
rect 61773 59626 63386 59829
tri 63386 59626 63673 59913 sw
tri 63673 59626 63960 59913 ne
rect 63960 59626 71000 59913
rect 61773 59546 63673 59626
rect 59696 59360 61490 59546
rect 55363 59164 57147 59360
rect 53171 59088 55075 59164
rect 51170 58825 52887 59088
rect 46910 58551 50885 58825
rect 42800 58436 46599 58551
tri 46599 58436 46714 58551 sw
tri 46910 58436 47025 58551 ne
rect 47025 58541 50885 58551
tri 50885 58541 51169 58825 sw
tri 51170 58541 51454 58825 ne
rect 51454 58804 52887 58825
tri 52887 58804 53171 59088 sw
tri 53171 58804 53455 59088 ne
rect 53455 59004 55075 59088
tri 55075 59004 55235 59164 sw
tri 55363 59004 55523 59164 ne
rect 55523 59074 57147 59164
tri 57147 59074 57433 59360 sw
tri 57433 59074 57719 59360 ne
rect 57719 59077 59413 59360
tri 59413 59077 59696 59360 sw
tri 59696 59077 59979 59360 ne
rect 59979 59263 61490 59360
tri 61490 59263 61773 59546 sw
tri 61773 59263 62056 59546 ne
rect 62056 59461 63673 59546
tri 63673 59461 63838 59626 sw
tri 63960 59461 64125 59626 ne
rect 64125 59461 71000 59626
rect 62056 59263 63838 59461
rect 59979 59077 61773 59263
rect 57719 59074 59696 59077
rect 55523 59004 57433 59074
rect 53455 58804 55235 59004
rect 51454 58541 53171 58804
rect 47025 58520 51169 58541
tri 51169 58520 51190 58541 sw
tri 51454 58520 51475 58541 ne
rect 51475 58520 53171 58541
tri 53171 58520 53455 58804 sw
tri 53455 58520 53739 58804 ne
rect 53739 58716 55235 58804
tri 55235 58716 55523 59004 sw
tri 55523 58716 55811 59004 ne
rect 55811 58788 57433 59004
tri 57433 58788 57719 59074 sw
tri 57719 58788 58005 59074 ne
rect 58005 58980 59696 59074
tri 59696 58980 59793 59077 sw
tri 59979 58980 60076 59077 ne
rect 60076 58980 61773 59077
tri 61773 58980 62056 59263 sw
tri 62056 58980 62339 59263 ne
rect 62339 59174 63838 59263
tri 63838 59174 64125 59461 sw
tri 64125 59174 64412 59461 ne
rect 64412 59174 71000 59461
rect 62339 58980 64125 59174
rect 58005 58788 59793 58980
rect 55811 58716 57719 58788
rect 53739 58520 55523 58716
rect 47025 58436 51190 58520
rect 42800 58131 46714 58436
tri 46714 58131 47019 58436 sw
tri 47025 58131 47330 58436 ne
rect 47330 58235 51190 58436
tri 51190 58235 51475 58520 sw
tri 51475 58235 51760 58520 ne
rect 51760 58236 53455 58520
tri 53455 58236 53739 58520 sw
tri 53739 58236 54023 58520 ne
rect 54023 58428 55523 58520
tri 55523 58428 55811 58716 sw
tri 55811 58428 56099 58716 ne
rect 56099 58618 57719 58716
tri 57719 58618 57889 58788 sw
tri 58005 58618 58175 58788 ne
rect 58175 58697 59793 58788
tri 59793 58697 60076 58980 sw
tri 60076 58697 60359 58980 ne
rect 60359 58697 62056 58980
tri 62056 58697 62339 58980 sw
tri 62339 58697 62622 58980 ne
rect 62622 58887 64125 58980
tri 64125 58887 64412 59174 sw
tri 64412 58887 64699 59174 ne
rect 64699 58887 71000 59174
rect 62622 58697 64412 58887
rect 58175 58618 60076 58697
rect 56099 58428 57889 58618
rect 54023 58236 55811 58428
rect 51760 58235 53739 58236
rect 47330 58131 51475 58235
rect 42800 58097 47019 58131
tri 42800 58010 42887 58097 ne
rect 42887 58010 47019 58097
tri 42600 57810 42800 58010 sw
tri 42887 57810 43087 58010 ne
rect 43087 57888 47019 58010
tri 47019 57888 47262 58131 sw
tri 47330 57888 47573 58131 ne
rect 47573 57950 51475 58131
tri 51475 57950 51760 58235 sw
tri 51760 57950 52045 58235 ne
rect 52045 58140 53739 58235
tri 53739 58140 53835 58236 sw
tri 54023 58140 54119 58236 ne
rect 54119 58140 55811 58236
tri 55811 58140 56099 58428 sw
tri 56099 58140 56387 58428 ne
rect 56387 58332 57889 58428
tri 57889 58332 58175 58618 sw
tri 58175 58332 58461 58618 ne
rect 58461 58414 60076 58618
tri 60076 58414 60359 58697 sw
tri 60359 58414 60642 58697 ne
rect 60642 58600 62339 58697
tri 62339 58600 62436 58697 sw
tri 62622 58600 62719 58697 ne
rect 62719 58600 64412 58697
tri 64412 58600 64699 58887 sw
tri 64699 58800 64786 58887 ne
rect 64786 58800 71000 58887
rect 60642 58414 62436 58600
rect 58461 58332 60359 58414
rect 56387 58140 58175 58332
rect 52045 57950 53835 58140
rect 47573 57888 51760 57950
rect 43087 57810 47262 57888
rect 41200 57722 42800 57810
tri 42800 57722 42888 57810 sw
tri 43087 57722 43175 57810 ne
rect 43175 57722 47262 57810
rect 41200 57435 42888 57722
tri 42888 57435 43175 57722 sw
tri 43175 57435 43462 57722 ne
rect 43462 57582 47262 57722
tri 47262 57582 47568 57888 sw
tri 47573 57582 47879 57888 ne
rect 47879 57774 51760 57888
tri 51760 57774 51936 57950 sw
tri 52045 57774 52221 57950 ne
rect 52221 57856 53835 57950
tri 53835 57856 54119 58140 sw
tri 54119 57856 54403 58140 ne
rect 54403 57856 56099 58140
rect 52221 57774 54119 57856
rect 47879 57582 51936 57774
rect 43462 57562 47568 57582
tri 47568 57562 47588 57582 sw
tri 47879 57562 47899 57582 ne
rect 47899 57562 51936 57582
rect 43462 57435 47588 57562
rect 41200 57430 43175 57435
tri 41200 57338 41292 57430 ne
rect 41292 57338 43175 57430
tri 41000 57132 41206 57338 sw
tri 41292 57132 41498 57338 ne
rect 41498 57322 43175 57338
tri 43175 57322 43288 57435 sw
tri 43462 57322 43575 57435 ne
rect 43575 57322 47588 57435
rect 41498 57132 43288 57322
rect 39600 56840 41206 57132
tri 41206 56840 41498 57132 sw
tri 41498 56840 41790 57132 ne
rect 41790 57035 43288 57132
tri 43288 57035 43575 57322 sw
tri 43575 57035 43862 57322 ne
rect 43862 57260 47588 57322
tri 47588 57260 47890 57562 sw
tri 47899 57260 48201 57562 ne
rect 48201 57489 51936 57562
tri 51936 57489 52221 57774 sw
tri 52221 57489 52506 57774 ne
rect 52506 57572 54119 57774
tri 54119 57572 54403 57856 sw
tri 54403 57572 54687 57856 ne
rect 54687 57852 56099 57856
tri 56099 57852 56387 58140 sw
tri 56387 57852 56675 58140 ne
rect 56675 58046 58175 58140
tri 58175 58046 58461 58332 sw
tri 58461 58046 58747 58332 ne
rect 58747 58229 60359 58332
tri 60359 58229 60544 58414 sw
tri 60642 58229 60827 58414 ne
rect 60827 58317 62436 58414
tri 62436 58317 62719 58600 sw
tri 62719 58317 63002 58600 ne
rect 63002 58317 71000 58600
rect 60827 58229 62719 58317
rect 58747 58046 60544 58229
rect 56675 57852 58461 58046
rect 54687 57760 56387 57852
tri 56387 57760 56479 57852 sw
tri 56675 57760 56767 57852 ne
rect 56767 57760 58461 57852
tri 58461 57760 58747 58046 sw
tri 58747 57760 59033 58046 ne
rect 59033 57946 60544 58046
tri 60544 57946 60827 58229 sw
tri 60827 57946 61110 58229 ne
rect 61110 58034 62719 58229
tri 62719 58034 63002 58317 sw
tri 63002 58034 63285 58317 ne
rect 63285 58034 71000 58317
rect 61110 57946 63002 58034
rect 59033 57760 60827 57946
rect 54687 57572 56479 57760
rect 52506 57489 54403 57572
rect 48201 57487 52221 57489
tri 52221 57487 52223 57489 sw
tri 52506 57487 52508 57489 ne
rect 52508 57487 54403 57489
rect 48201 57260 52223 57487
rect 43862 57126 47890 57260
tri 47890 57126 48024 57260 sw
tri 48201 57126 48335 57260 ne
rect 48335 57202 52223 57260
tri 52223 57202 52508 57487 sw
tri 52508 57202 52793 57487 ne
rect 52793 57392 54403 57487
tri 54403 57392 54583 57572 sw
tri 54687 57392 54867 57572 ne
rect 54867 57472 56479 57572
tri 56479 57472 56767 57760 sw
tri 56767 57472 57055 57760 ne
rect 57055 57474 58747 57760
tri 58747 57474 59033 57760 sw
tri 59033 57474 59319 57760 ne
rect 59319 57663 60827 57760
tri 60827 57663 61110 57946 sw
tri 61110 57663 61393 57946 ne
rect 61393 57849 63002 57946
tri 63002 57849 63187 58034 sw
tri 63285 57849 63470 58034 ne
rect 63470 57849 71000 58034
rect 61393 57663 63187 57849
rect 59319 57474 61110 57663
rect 57055 57472 59033 57474
rect 54867 57392 56767 57472
rect 52793 57202 54583 57392
rect 48335 57201 52508 57202
tri 52508 57201 52509 57202 sw
tri 52793 57201 52794 57202 ne
rect 52794 57201 54583 57202
rect 48335 57126 52509 57201
rect 43862 57035 48024 57126
rect 41790 56840 43575 57035
rect 39600 56758 41498 56840
tri 39600 56665 39693 56758 ne
rect 39693 56665 41498 56758
tri 39400 56465 39600 56665 sw
tri 39693 56465 39893 56665 ne
rect 39893 56548 41498 56665
tri 41498 56548 41790 56840 sw
tri 41790 56548 42082 56840 ne
rect 42082 56748 43575 56840
tri 43575 56748 43862 57035 sw
tri 43862 56748 44149 57035 ne
rect 44149 56820 48024 57035
tri 48024 56820 48330 57126 sw
tri 48335 56820 48641 57126 ne
rect 48641 56916 52509 57126
tri 52509 56916 52794 57201 sw
tri 52794 56916 53079 57201 ne
rect 53079 57108 54583 57201
tri 54583 57108 54867 57392 sw
tri 54867 57108 55151 57392 ne
rect 55151 57184 56767 57392
tri 56767 57184 57055 57472 sw
tri 57055 57184 57343 57472 ne
rect 57343 57380 59033 57472
tri 59033 57380 59127 57474 sw
tri 59319 57380 59413 57474 ne
rect 59413 57380 61110 57474
tri 61110 57380 61393 57663 sw
tri 61393 57380 61676 57663 ne
rect 61676 57566 63187 57663
tri 63187 57566 63470 57849 sw
tri 63470 57566 63753 57849 ne
rect 63753 57566 71000 57849
rect 61676 57380 63470 57566
rect 57343 57184 59127 57380
rect 55151 57108 57055 57184
rect 53079 56916 54867 57108
rect 48641 56914 52794 56916
tri 52794 56914 52796 56916 sw
tri 53079 56914 53081 56916 ne
rect 53081 56914 54867 56916
rect 48641 56820 52796 56914
rect 44149 56800 48330 56820
tri 48330 56800 48350 56820 sw
tri 48641 56800 48661 56820 ne
rect 48661 56800 52796 56820
rect 44149 56748 48350 56800
rect 42082 56747 43862 56748
tri 43862 56747 43863 56748 sw
tri 44149 56747 44150 56748 ne
rect 44150 56747 48350 56748
rect 42082 56548 43863 56747
rect 39893 56465 41790 56548
rect 36400 56371 39600 56465
tri 39600 56371 39694 56465 sw
tri 39893 56371 39987 56465 ne
rect 39987 56371 41790 56465
rect 36400 56078 39694 56371
tri 39694 56078 39987 56371 sw
tri 39987 56078 40280 56371 ne
rect 40280 56322 41790 56371
tri 41790 56322 42016 56548 sw
tri 42082 56322 42308 56548 ne
rect 42308 56460 43863 56548
tri 43863 56460 44150 56747 sw
tri 44150 56460 44437 56747 ne
rect 44437 56494 48350 56747
tri 48350 56494 48656 56800 sw
tri 48661 56494 48967 56800 ne
rect 48967 56630 52796 56800
tri 52796 56630 53080 56914 sw
tri 53081 56630 53365 56914 ne
rect 53365 56824 54867 56914
tri 54867 56824 55151 57108 sw
tri 55151 56824 55435 57108 ne
rect 55435 57024 57055 57108
tri 57055 57024 57215 57184 sw
tri 57343 57024 57503 57184 ne
rect 57503 57094 59127 57184
tri 59127 57094 59413 57380 sw
tri 59413 57094 59699 57380 ne
rect 59699 57097 61393 57380
tri 61393 57097 61676 57380 sw
tri 61676 57097 61959 57380 ne
rect 61959 57283 63470 57380
tri 63470 57283 63753 57566 sw
tri 63753 57283 64036 57566 ne
rect 64036 57283 71000 57566
rect 61959 57097 63753 57283
rect 59699 57094 61676 57097
rect 57503 57024 59413 57094
rect 55435 56824 57215 57024
rect 53365 56630 55151 56824
rect 48967 56540 53080 56630
tri 53080 56540 53170 56630 sw
tri 53365 56540 53455 56630 ne
rect 53455 56540 55151 56630
tri 55151 56540 55435 56824 sw
tri 55435 56540 55719 56824 ne
rect 55719 56736 57215 56824
tri 57215 56736 57503 57024 sw
tri 57503 56736 57791 57024 ne
rect 57791 56808 59413 57024
tri 59413 56808 59699 57094 sw
tri 59699 56808 59985 57094 ne
rect 59985 57000 61676 57094
tri 61676 57000 61773 57097 sw
tri 61959 57000 62056 57097 ne
rect 62056 57000 63753 57097
tri 63753 57000 64036 57283 sw
tri 64036 57200 64119 57283 ne
rect 64119 57200 71000 57283
rect 59985 56808 61773 57000
rect 57791 56736 59699 56808
rect 55719 56540 57503 56736
rect 48967 56494 53170 56540
rect 44437 56475 48656 56494
tri 48656 56475 48675 56494 sw
tri 48967 56475 48986 56494 ne
rect 48986 56475 53170 56494
rect 44437 56460 48675 56475
rect 42308 56459 44150 56460
tri 44150 56459 44151 56460 sw
tri 44437 56459 44438 56460 ne
rect 44438 56459 48675 56460
rect 42308 56322 44151 56459
rect 40280 56078 42016 56322
rect 36400 55785 39987 56078
tri 39987 55785 40280 56078 sw
tri 40280 55785 40573 56078 ne
rect 40573 56030 42016 56078
tri 42016 56030 42308 56322 sw
tri 42308 56030 42600 56322 ne
rect 42600 56172 44151 56322
tri 44151 56172 44438 56459 sw
tri 44438 56172 44725 56459 ne
rect 44725 56172 48675 56459
rect 42600 56030 44438 56172
rect 40573 55785 42308 56030
rect 36400 55492 40280 55785
tri 40280 55492 40573 55785 sw
tri 40573 55492 40866 55785 ne
rect 40866 55738 42308 55785
tri 42308 55738 42600 56030 sw
tri 42600 55738 42892 56030 ne
rect 42892 55885 44438 56030
tri 44438 55885 44725 56172 sw
tri 44725 55885 45012 56172 ne
rect 45012 56169 48675 56172
tri 48675 56169 48981 56475 sw
tri 48986 56169 49292 56475 ne
rect 49292 56255 53170 56475
tri 53170 56255 53455 56540 sw
tri 53455 56255 53740 56540 ne
rect 53740 56256 55435 56540
tri 55435 56256 55719 56540 sw
tri 55719 56256 56003 56540 ne
rect 56003 56448 57503 56540
tri 57503 56448 57791 56736 sw
tri 57791 56448 58079 56736 ne
rect 58079 56638 59699 56736
tri 59699 56638 59869 56808 sw
tri 59985 56638 60155 56808 ne
rect 60155 56717 61773 56808
tri 61773 56717 62056 57000 sw
tri 62056 56717 62339 57000 ne
rect 62339 56717 71000 57000
rect 60155 56638 62056 56717
rect 58079 56448 59869 56638
rect 56003 56256 57791 56448
rect 53740 56255 55719 56256
rect 49292 56169 53455 56255
rect 45012 56150 48981 56169
tri 48981 56150 49000 56169 sw
tri 49292 56150 49311 56169 ne
rect 49311 56150 53455 56169
rect 45012 55885 49000 56150
rect 42892 55884 44725 55885
tri 44725 55884 44726 55885 sw
tri 45012 55884 45013 55885 ne
rect 45013 55884 49000 55885
rect 42892 55738 44726 55884
rect 40866 55492 42600 55738
rect 36400 55421 40573 55492
tri 36400 55324 36497 55421 ne
rect 36497 55324 40573 55421
tri 36200 55027 36497 55324 sw
tri 36497 55027 36794 55324 ne
rect 36794 55199 40573 55324
tri 40573 55199 40866 55492 sw
tri 40866 55199 41159 55492 ne
rect 41159 55446 42600 55492
tri 42600 55446 42892 55738 sw
tri 42892 55446 43184 55738 ne
rect 43184 55597 44726 55738
tri 44726 55597 45013 55884 sw
tri 45013 55597 45300 55884 ne
rect 45300 55844 49000 55884
tri 49000 55844 49306 56150 sw
tri 49311 55844 49617 56150 ne
rect 49617 55970 53455 56150
tri 53455 55970 53740 56255 sw
tri 53740 55970 54025 56255 ne
rect 54025 56160 55719 56255
tri 55719 56160 55815 56256 sw
tri 56003 56160 56099 56256 ne
rect 56099 56160 57791 56256
tri 57791 56160 58079 56448 sw
tri 58079 56160 58367 56448 ne
rect 58367 56352 59869 56448
tri 59869 56352 60155 56638 sw
tri 60155 56352 60441 56638 ne
rect 60441 56434 62056 56638
tri 62056 56434 62339 56717 sw
tri 62339 56434 62622 56717 ne
rect 62622 56434 71000 56717
rect 60441 56352 62339 56434
rect 58367 56160 60155 56352
rect 54025 55970 55815 56160
rect 49617 55968 53740 55970
tri 53740 55968 53742 55970 sw
tri 54025 55968 54027 55970 ne
rect 54027 55968 55815 55970
rect 49617 55844 53742 55968
rect 45300 55597 49306 55844
rect 43184 55446 45013 55597
rect 41159 55444 42892 55446
tri 42892 55444 42894 55446 sw
tri 43184 55444 43186 55446 ne
rect 43186 55444 45013 55446
rect 41159 55199 42894 55444
rect 36794 55154 40866 55199
tri 40866 55154 40911 55199 sw
tri 41159 55154 41204 55199 ne
rect 41204 55154 42894 55199
rect 36794 55027 40911 55154
rect 33200 54827 36497 55027
tri 36497 54827 36697 55027 sw
tri 36794 54827 36994 55027 ne
rect 36994 54861 40911 55027
tri 40911 54861 41204 55154 sw
tri 41204 54861 41497 55154 ne
rect 41497 55152 42894 55154
tri 42894 55152 43186 55444 sw
tri 43186 55152 43478 55444 ne
rect 43478 55343 45013 55444
tri 45013 55343 45267 55597 sw
tri 45300 55343 45554 55597 ne
rect 45554 55559 49306 55597
tri 49306 55559 49591 55844 sw
tri 49617 55559 49902 55844 ne
rect 49902 55683 53742 55844
tri 53742 55683 54027 55968 sw
tri 54027 55683 54312 55968 ne
rect 54312 55876 55815 55968
tri 55815 55876 56099 56160 sw
tri 56099 55876 56383 56160 ne
rect 56383 55876 58079 56160
rect 54312 55683 56099 55876
rect 49902 55682 54027 55683
tri 54027 55682 54028 55683 sw
tri 54312 55682 54313 55683 ne
rect 54313 55682 56099 55683
rect 49902 55559 54028 55682
rect 45554 55343 49591 55559
rect 43478 55272 45267 55343
tri 45267 55272 45338 55343 sw
tri 45554 55272 45625 55343 ne
rect 45625 55272 49591 55343
rect 43478 55152 45338 55272
rect 41497 54861 43186 55152
rect 36994 54827 41204 54861
rect 33200 54728 36697 54827
tri 36697 54728 36796 54827 sw
tri 36994 54728 37093 54827 ne
rect 37093 54728 41204 54827
rect 33200 54431 36796 54728
tri 36796 54431 37093 54728 sw
tri 37093 54431 37390 54728 ne
rect 37390 54568 41204 54728
tri 41204 54568 41497 54861 sw
tri 41497 54568 41790 54861 ne
rect 41790 54860 43186 54861
tri 43186 54860 43478 55152 sw
tri 43478 54860 43770 55152 ne
rect 43770 55055 45338 55152
tri 45338 55055 45555 55272 sw
tri 45625 55055 45842 55272 ne
rect 45842 55257 49591 55272
tri 49591 55257 49893 55559 sw
tri 49902 55257 50204 55559 ne
rect 50204 55397 54028 55559
tri 54028 55397 54313 55682 sw
tri 54313 55397 54598 55682 ne
rect 54598 55592 56099 55682
tri 56099 55592 56383 55876 sw
tri 56383 55592 56667 55876 ne
rect 56667 55872 58079 55876
tri 58079 55872 58367 56160 sw
tri 58367 55872 58655 56160 ne
rect 58655 56066 60155 56160
tri 60155 56066 60441 56352 sw
tri 60441 56066 60727 56352 ne
rect 60727 56249 62339 56352
tri 62339 56249 62524 56434 sw
tri 62622 56249 62807 56434 ne
rect 62807 56249 71000 56434
rect 60727 56066 62524 56249
rect 58655 55872 60441 56066
rect 56667 55780 58367 55872
tri 58367 55780 58459 55872 sw
tri 58655 55780 58747 55872 ne
rect 58747 55780 60441 55872
tri 60441 55780 60727 56066 sw
tri 60727 55780 61013 56066 ne
rect 61013 55966 62524 56066
tri 62524 55966 62807 56249 sw
tri 62807 55966 63090 56249 ne
rect 63090 55966 71000 56249
rect 61013 55780 62807 55966
rect 56667 55592 58459 55780
rect 54598 55412 56383 55592
tri 56383 55412 56563 55592 sw
tri 56667 55412 56847 55592 ne
rect 56847 55492 58459 55592
tri 58459 55492 58747 55780 sw
tri 58747 55492 59035 55780 ne
rect 59035 55494 60727 55780
tri 60727 55494 61013 55780 sw
tri 61013 55494 61299 55780 ne
rect 61299 55683 62807 55780
tri 62807 55683 63090 55966 sw
tri 63090 55683 63373 55966 ne
rect 63373 55683 71000 55966
rect 61299 55494 63090 55683
rect 59035 55492 61013 55494
rect 56847 55412 58747 55492
rect 54598 55397 56563 55412
rect 50204 55257 54313 55397
rect 45842 55055 49893 55257
rect 43770 54860 45555 55055
rect 41790 54568 43478 54860
tri 43478 54568 43770 54860 sw
tri 43770 54568 44062 54860 ne
rect 44062 54768 45555 54860
tri 45555 54768 45842 55055 sw
tri 45842 54768 46129 55055 ne
rect 46129 54946 49893 55055
tri 49893 54946 50204 55257 sw
tri 50204 54946 50515 55257 ne
rect 50515 55135 54313 55257
tri 54313 55135 54575 55397 sw
tri 54598 55135 54860 55397 ne
rect 54860 55135 56563 55397
rect 50515 54946 54575 55135
rect 46129 54768 50204 54946
rect 44062 54767 45842 54768
tri 45842 54767 45843 54768 sw
tri 46129 54767 46130 54768 ne
rect 46130 54767 50204 54768
rect 44062 54568 45843 54767
rect 37390 54567 41497 54568
tri 41497 54567 41498 54568 sw
tri 41790 54567 41791 54568 ne
rect 41791 54567 43770 54568
rect 37390 54431 41498 54567
rect 33200 54429 37093 54431
tri 37093 54429 37095 54431 sw
tri 37390 54429 37392 54431 ne
rect 37392 54429 41498 54431
rect 33200 54133 37095 54429
tri 37095 54133 37391 54429 sw
tri 37392 54133 37688 54429 ne
rect 37688 54274 41498 54429
tri 41498 54274 41791 54567 sw
tri 41791 54274 42084 54567 ne
rect 42084 54402 43770 54567
tri 43770 54402 43936 54568 sw
tri 44062 54402 44228 54568 ne
rect 44228 54480 45843 54568
tri 45843 54480 46130 54767 sw
tri 46130 54480 46417 54767 ne
rect 46417 54640 50204 54767
tri 50204 54640 50510 54946 sw
tri 50515 54640 50821 54946 ne
rect 50821 54850 54575 54946
tri 54575 54850 54860 55135 sw
tri 54860 54850 55145 55135 ne
rect 55145 55128 56563 55135
tri 56563 55128 56847 55412 sw
tri 56847 55128 57131 55412 ne
rect 57131 55204 58747 55412
tri 58747 55204 59035 55492 sw
tri 59035 55204 59323 55492 ne
rect 59323 55400 61013 55492
tri 61013 55400 61107 55494 sw
tri 61299 55400 61393 55494 ne
rect 61393 55400 63090 55494
tri 63090 55400 63373 55683 sw
tri 63373 55600 63456 55683 ne
rect 63456 55600 71000 55683
rect 59323 55204 61107 55400
rect 57131 55128 59035 55204
rect 55145 54850 56847 55128
rect 50821 54848 54860 54850
tri 54860 54848 54862 54850 sw
tri 55145 54848 55147 54850 ne
rect 55147 54848 56847 54850
rect 50821 54640 54862 54848
rect 46417 54620 50510 54640
tri 50510 54620 50530 54640 sw
tri 50821 54620 50841 54640 ne
rect 50841 54620 54862 54640
rect 46417 54480 50530 54620
rect 44228 54402 46130 54480
rect 42084 54274 43936 54402
rect 37688 54273 41791 54274
tri 41791 54273 41792 54274 sw
tri 42084 54273 42085 54274 ne
rect 42085 54273 43936 54274
rect 37688 54133 41792 54273
rect 33200 54080 37391 54133
tri 37391 54080 37444 54133 sw
tri 37688 54080 37741 54133 ne
rect 37741 54080 41792 54133
tri 33200 53992 33288 54080 ne
rect 33288 53992 37444 54080
tri 33000 53704 33288 53992 sw
tri 33288 53704 33576 53992 ne
rect 33576 53783 37444 53992
tri 37444 53783 37741 54080 sw
tri 37741 53783 38038 54080 ne
rect 38038 53980 41792 54080
tri 41792 53980 42085 54273 sw
tri 42085 53980 42378 54273 ne
rect 42378 54188 43936 54273
tri 43936 54188 44150 54402 sw
tri 44228 54188 44442 54402 ne
rect 44442 54285 46130 54402
tri 46130 54285 46325 54480 sw
tri 46417 54285 46612 54480 ne
rect 46612 54312 50530 54480
tri 50530 54312 50838 54620 sw
tri 50841 54312 51149 54620 ne
rect 51149 54563 54862 54620
tri 54862 54563 55147 54848 sw
tri 55147 54563 55432 54848 ne
rect 55432 54844 56847 54848
tri 56847 54844 57131 55128 sw
tri 57131 54844 57415 55128 ne
rect 57415 55044 59035 55128
tri 59035 55044 59195 55204 sw
tri 59323 55044 59483 55204 ne
rect 59483 55114 61107 55204
tri 61107 55114 61393 55400 sw
tri 61393 55114 61679 55400 ne
rect 61679 55114 71000 55400
rect 59483 55044 61393 55114
rect 57415 54844 59195 55044
rect 55432 54563 57131 54844
rect 51149 54312 55147 54563
rect 46612 54285 50838 54312
rect 44442 54188 46325 54285
rect 42378 53980 44150 54188
rect 38038 53783 42085 53980
rect 33576 53768 37741 53783
tri 37741 53768 37756 53783 sw
tri 38038 53768 38053 53783 ne
rect 38053 53768 42085 53783
rect 33576 53704 37756 53768
rect 30000 53504 33288 53704
tri 33288 53504 33488 53704 sw
tri 33576 53504 33776 53704 ne
rect 33776 53504 37756 53704
rect 30000 53414 33488 53504
tri 33488 53414 33578 53504 sw
tri 33776 53414 33866 53504 ne
rect 33866 53471 37756 53504
tri 37756 53471 38053 53768 sw
tri 38053 53471 38350 53768 ne
rect 38350 53687 42085 53768
tri 42085 53687 42378 53980 sw
tri 42378 53687 42671 53980 ne
rect 42671 53896 44150 53980
tri 44150 53896 44442 54188 sw
tri 44442 53896 44734 54188 ne
rect 44734 53998 46325 54188
tri 46325 53998 46612 54285 sw
tri 46612 53998 46899 54285 ne
rect 46899 54187 50838 54285
tri 50838 54187 50963 54312 sw
tri 51149 54187 51274 54312 ne
rect 51274 54278 55147 54312
tri 55147 54278 55432 54563 sw
tri 55432 54278 55717 54563 ne
rect 55717 54560 57131 54563
tri 57131 54560 57415 54844 sw
tri 57415 54560 57699 54844 ne
rect 57699 54756 59195 54844
tri 59195 54756 59483 55044 sw
tri 59483 54756 59771 55044 ne
rect 59771 54828 61393 55044
tri 61393 54828 61679 55114 sw
tri 61679 54828 61965 55114 ne
rect 61965 54828 71000 55114
rect 59771 54756 61679 54828
rect 57699 54560 59483 54756
rect 55717 54278 57415 54560
rect 51274 54273 55432 54278
tri 55432 54273 55437 54278 sw
tri 55717 54273 55722 54278 ne
rect 55722 54276 57415 54278
tri 57415 54276 57699 54560 sw
tri 57699 54276 57983 54560 ne
rect 57983 54468 59483 54560
tri 59483 54468 59771 54756 sw
tri 59771 54468 60059 54756 ne
rect 60059 54658 61679 54756
tri 61679 54658 61849 54828 sw
tri 61965 54658 62135 54828 ne
rect 62135 54658 71000 54828
rect 60059 54468 61849 54658
rect 57983 54276 59771 54468
rect 55722 54273 57699 54276
rect 51274 54187 55437 54273
rect 46899 53998 50963 54187
rect 44734 53997 46612 53998
tri 46612 53997 46613 53998 sw
tri 46899 53997 46900 53998 ne
rect 46900 53997 50963 53998
rect 44734 53896 46613 53997
rect 42671 53756 44442 53896
tri 44442 53756 44582 53896 sw
tri 44734 53756 44874 53896 ne
rect 44874 53756 46613 53896
rect 42671 53687 44582 53756
rect 38350 53471 42378 53687
rect 33866 53470 38053 53471
tri 38053 53470 38054 53471 sw
tri 38350 53470 38351 53471 ne
rect 38351 53470 42378 53471
rect 33866 53414 38054 53470
rect 30000 53126 33578 53414
tri 33578 53126 33866 53414 sw
tri 33866 53126 34154 53414 ne
rect 34154 53173 38054 53414
tri 38054 53173 38351 53470 sw
tri 38351 53173 38648 53470 ne
rect 38648 53468 42378 53470
tri 42378 53468 42597 53687 sw
tri 42671 53468 42890 53687 ne
rect 42890 53468 44582 53687
rect 38648 53175 42597 53468
tri 42597 53175 42890 53468 sw
tri 42890 53175 43183 53468 ne
rect 43183 53464 44582 53468
tri 44582 53464 44874 53756 sw
tri 44874 53464 45166 53756 ne
rect 45166 53710 46613 53756
tri 46613 53710 46900 53997 sw
tri 46900 53710 47187 53997 ne
rect 47187 53879 50963 53997
tri 50963 53879 51271 54187 sw
tri 51274 53879 51582 54187 ne
rect 51582 53988 55437 54187
tri 55437 53988 55722 54273 sw
tri 55722 53988 56007 54273 ne
rect 56007 54180 57699 54273
tri 57699 54180 57795 54276 sw
tri 57983 54180 58079 54276 ne
rect 58079 54180 59771 54276
tri 59771 54180 60059 54468 sw
tri 60059 54180 60347 54468 ne
rect 60347 54372 61849 54468
tri 61849 54372 62135 54658 sw
tri 62135 54372 62421 54658 ne
rect 62421 54372 71000 54658
rect 60347 54180 62135 54372
rect 56007 53988 57795 54180
rect 51582 53879 55722 53988
rect 47187 53710 51271 53879
rect 45166 53464 46900 53710
rect 43183 53175 44874 53464
rect 38648 53173 42890 53175
rect 34154 53126 38351 53173
rect 30000 53124 33866 53126
tri 33866 53124 33868 53126 sw
tri 34154 53124 34156 53126 ne
rect 34156 53124 38351 53126
rect 30000 52836 33868 53124
tri 33868 52836 34156 53124 sw
tri 34156 52836 34444 53124 ne
rect 34444 53079 38351 53124
tri 38351 53079 38445 53173 sw
tri 38648 53079 38742 53173 ne
rect 38742 53079 42890 53173
rect 34444 52836 38445 53079
rect 30000 52835 34156 52836
tri 34156 52835 34157 52836 sw
tri 34444 52835 34445 52836 ne
rect 34445 52835 38445 52836
rect 30000 52748 34157 52835
tri 30000 52654 30094 52748 ne
rect 30094 52654 34157 52748
tri 29800 52360 30094 52654 sw
tri 30094 52360 30388 52654 ne
rect 30388 52547 34157 52654
tri 34157 52547 34445 52835 sw
tri 34445 52547 34733 52835 ne
rect 34733 52782 38445 52835
tri 38445 52782 38742 53079 sw
tri 38742 52782 39039 53079 ne
rect 39039 52882 42890 53079
tri 42890 52882 43183 53175 sw
tri 43183 52882 43476 53175 ne
rect 43476 53172 44874 53175
tri 44874 53172 45166 53464 sw
tri 45166 53172 45458 53464 ne
rect 45458 53423 46900 53464
tri 46900 53423 47187 53710 sw
tri 47187 53423 47474 53710 ne
rect 47474 53645 51271 53710
tri 51271 53645 51505 53879 sw
tri 51582 53645 51816 53879 ne
rect 51816 53704 55722 53879
tri 55722 53704 56006 53988 sw
tri 56007 53704 56291 53988 ne
rect 56291 53896 57795 53988
tri 57795 53896 58079 54180 sw
tri 58079 53896 58363 54180 ne
rect 58363 53896 60059 54180
rect 56291 53704 58079 53896
rect 51816 53645 56006 53704
rect 47474 53423 51505 53645
rect 45458 53362 47187 53423
tri 47187 53362 47248 53423 sw
tri 47474 53362 47535 53423 ne
rect 47535 53362 51505 53423
rect 45458 53172 47248 53362
rect 43476 52882 45166 53172
rect 39039 52881 43183 52882
tri 43183 52881 43184 52882 sw
tri 43476 52881 43477 52882 ne
rect 43477 52881 45166 52882
rect 39039 52782 43184 52881
rect 34733 52575 38742 52782
tri 38742 52575 38949 52782 sw
tri 39039 52575 39246 52782 ne
rect 39246 52588 43184 52782
tri 43184 52588 43477 52881 sw
tri 43477 52588 43770 52881 ne
rect 43770 52880 45166 52881
tri 45166 52880 45458 53172 sw
tri 45458 52880 45750 53172 ne
rect 45750 53075 47248 53172
tri 47248 53075 47535 53362 sw
tri 47535 53075 47822 53362 ne
rect 47822 53339 51505 53362
tri 51505 53339 51811 53645 sw
tri 51816 53339 52122 53645 ne
rect 52122 53531 56006 53645
tri 56006 53531 56179 53704 sw
tri 56291 53531 56464 53704 ne
rect 56464 53612 58079 53704
tri 58079 53612 58363 53896 sw
tri 58363 53612 58647 53896 ne
rect 58647 53892 60059 53896
tri 60059 53892 60347 54180 sw
tri 60347 53892 60635 54180 ne
rect 60635 54086 62135 54180
tri 62135 54086 62421 54372 sw
tri 62421 54086 62707 54372 ne
rect 62707 54086 71000 54372
rect 60635 53892 62421 54086
rect 58647 53800 60347 53892
tri 60347 53800 60439 53892 sw
tri 60635 53800 60727 53892 ne
rect 60727 53800 62421 53892
tri 62421 53800 62707 54086 sw
tri 62707 54000 62793 54086 ne
rect 62793 54000 71000 54086
rect 58647 53612 60439 53800
rect 56464 53531 58363 53612
rect 52122 53339 56179 53531
rect 47822 53252 51811 53339
tri 51811 53252 51898 53339 sw
tri 52122 53252 52209 53339 ne
rect 52209 53252 56179 53339
rect 47822 53075 51898 53252
rect 45750 52880 47535 53075
rect 43770 52588 45458 52880
tri 45458 52588 45750 52880 sw
tri 45750 52588 46042 52880 ne
rect 46042 52788 47535 52880
tri 47535 52788 47822 53075 sw
tri 47822 52788 48109 53075 ne
rect 48109 52946 51898 53075
tri 51898 52946 52204 53252 sw
tri 52209 52946 52515 53252 ne
rect 52515 53246 56179 53252
tri 56179 53246 56464 53531 sw
tri 56464 53246 56749 53531 ne
rect 56749 53432 58363 53531
tri 58363 53432 58543 53612 sw
tri 58647 53432 58827 53612 ne
rect 58827 53512 60439 53612
tri 60439 53512 60727 53800 sw
tri 60727 53512 61015 53800 ne
rect 61015 53512 71000 53800
rect 58827 53432 60727 53512
rect 56749 53246 58543 53432
rect 52515 53244 56464 53246
tri 56464 53244 56466 53246 sw
tri 56749 53244 56751 53246 ne
rect 56751 53244 58543 53246
rect 52515 52959 56466 53244
tri 56466 52959 56751 53244 sw
tri 56751 52959 57036 53244 ne
rect 57036 53148 58543 53244
tri 58543 53148 58827 53432 sw
tri 58827 53148 59111 53432 ne
rect 59111 53224 60727 53432
tri 60727 53224 61015 53512 sw
tri 61015 53224 61303 53512 ne
rect 61303 53224 71000 53512
rect 59111 53148 61015 53224
rect 57036 52959 58827 53148
rect 52515 52958 56751 52959
tri 56751 52958 56752 52959 sw
tri 57036 52958 57037 52959 ne
rect 57037 52958 58827 52959
rect 52515 52946 56752 52958
rect 48109 52927 52204 52946
tri 52204 52927 52223 52946 sw
tri 52515 52927 52534 52946 ne
rect 52534 52927 56752 52946
rect 48109 52788 52223 52927
rect 46042 52787 47822 52788
tri 47822 52787 47823 52788 sw
tri 48109 52787 48110 52788 ne
rect 48110 52787 52223 52788
rect 46042 52588 47823 52787
rect 39246 52587 43477 52588
tri 43477 52587 43478 52588 sw
tri 43770 52587 43771 52588 ne
rect 43771 52587 45750 52588
rect 39246 52575 43478 52587
rect 34733 52547 38949 52575
rect 30388 52546 34445 52547
tri 34445 52546 34446 52547 sw
tri 34733 52546 34734 52547 ne
rect 34734 52546 38949 52547
rect 30388 52360 34446 52546
rect 26800 52160 30094 52360
tri 30094 52160 30294 52360 sw
tri 30388 52160 30588 52360 ne
rect 30588 52258 34446 52360
tri 34446 52258 34734 52546 sw
tri 34734 52258 35022 52546 ne
rect 35022 52278 38949 52546
tri 38949 52278 39246 52575 sw
tri 39246 52278 39543 52575 ne
rect 39543 52294 43478 52575
tri 43478 52294 43771 52587 sw
tri 43771 52294 44064 52587 ne
rect 44064 52500 45750 52587
tri 45750 52500 45838 52588 sw
tri 46042 52500 46130 52588 ne
rect 46130 52500 47823 52588
tri 47823 52500 48110 52787 sw
tri 48110 52500 48397 52787 ne
rect 48397 52621 52223 52787
tri 52223 52621 52529 52927 sw
tri 52534 52621 52840 52927 ne
rect 52840 52673 56752 52927
tri 56752 52673 57037 52958 sw
tri 57037 52673 57322 52958 ne
rect 57322 52864 58827 52958
tri 58827 52864 59111 53148 sw
tri 59111 52864 59395 53148 ne
rect 59395 53064 61015 53148
tri 61015 53064 61175 53224 sw
tri 61303 53064 61463 53224 ne
rect 61463 53064 71000 53224
rect 59395 52864 61175 53064
rect 57322 52673 59111 52864
rect 52840 52621 57037 52673
rect 48397 52602 52529 52621
tri 52529 52602 52548 52621 sw
tri 52840 52602 52859 52621 ne
rect 52859 52602 57037 52621
rect 48397 52500 52548 52602
rect 44064 52294 45838 52500
rect 39543 52278 43771 52294
rect 35022 52258 39246 52278
rect 30588 52238 34734 52258
tri 34734 52238 34754 52258 sw
tri 35022 52238 35042 52258 ne
rect 35042 52238 39246 52258
rect 30588 52160 34754 52238
rect 26800 52064 30294 52160
tri 30294 52064 30390 52160 sw
tri 30588 52064 30684 52160 ne
rect 30684 52064 34754 52160
rect 26800 51770 30390 52064
tri 30390 51770 30684 52064 sw
tri 30684 51770 30978 52064 ne
rect 30978 51950 34754 52064
tri 34754 51950 35042 52238 sw
tri 35042 51950 35330 52238 ne
rect 35330 52129 39246 52238
tri 39246 52129 39395 52278 sw
tri 39543 52129 39692 52278 ne
rect 39692 52129 43771 52278
tri 43771 52129 43936 52294 sw
tri 44064 52129 44229 52294 ne
rect 44229 52208 45838 52294
tri 45838 52208 46130 52500 sw
tri 46130 52208 46422 52500 ne
rect 46422 52499 48110 52500
tri 48110 52499 48111 52500 sw
tri 48397 52499 48398 52500 ne
rect 48398 52499 52548 52500
rect 46422 52212 48111 52499
tri 48111 52212 48398 52499 sw
tri 48398 52212 48685 52499 ne
rect 48685 52296 52548 52499
tri 52548 52296 52854 52602 sw
tri 52859 52296 53165 52602 ne
rect 53165 52582 57037 52602
tri 57037 52582 57128 52673 sw
tri 57322 52582 57413 52673 ne
rect 57413 52582 59111 52673
rect 53165 52297 57128 52582
tri 57128 52297 57413 52582 sw
tri 57413 52297 57698 52582 ne
rect 57698 52580 59111 52582
tri 59111 52580 59395 52864 sw
tri 59395 52580 59679 52864 ne
rect 59679 52776 61175 52864
tri 61175 52776 61463 53064 sw
tri 61463 52776 61751 53064 ne
rect 61751 52776 71000 53064
rect 59679 52580 61463 52776
rect 57698 52297 59395 52580
rect 53165 52296 57413 52297
rect 48685 52277 52854 52296
tri 52854 52277 52873 52296 sw
tri 53165 52277 53184 52296 ne
rect 53184 52295 57413 52296
tri 57413 52295 57415 52297 sw
tri 57698 52295 57700 52297 ne
rect 57700 52296 59395 52297
tri 59395 52296 59679 52580 sw
tri 59679 52296 59963 52580 ne
rect 59963 52488 61463 52580
tri 61463 52488 61751 52776 sw
tri 61751 52488 62039 52776 ne
rect 62039 52488 71000 52776
rect 59963 52296 61751 52488
rect 57700 52295 59679 52296
rect 53184 52277 57415 52295
rect 48685 52212 52873 52277
rect 46422 52208 48398 52212
rect 44229 52129 46130 52208
rect 35330 51950 39395 52129
rect 30978 51949 35042 51950
tri 35042 51949 35043 51950 sw
tri 35330 51949 35331 51950 ne
rect 35331 51949 39395 51950
rect 30978 51770 35043 51949
rect 26800 51605 30684 51770
tri 30684 51605 30849 51770 sw
tri 30978 51605 31143 51770 ne
rect 31143 51661 35043 51770
tri 35043 51661 35331 51949 sw
tri 35331 51661 35619 51949 ne
rect 35619 51832 39395 51949
tri 39395 51832 39692 52129 sw
tri 39692 51832 39989 52129 ne
rect 39989 51836 43936 52129
tri 43936 51836 44229 52129 sw
tri 44229 51836 44522 52129 ne
rect 44522 51916 46130 52129
tri 46130 51916 46422 52208 sw
tri 46422 51916 46714 52208 ne
rect 46714 51925 48398 52208
tri 48398 51925 48685 52212 sw
tri 48685 51925 48972 52212 ne
rect 48972 51971 52873 52212
tri 52873 51971 53179 52277 sw
tri 53184 51971 53490 52277 ne
rect 53490 52010 57415 52277
tri 57415 52010 57700 52295 sw
tri 57700 52010 57985 52295 ne
rect 57985 52200 59679 52295
tri 59679 52200 59775 52296 sw
tri 59963 52200 60059 52296 ne
rect 60059 52200 61751 52296
tri 61751 52200 62039 52488 sw
tri 62039 52400 62127 52488 ne
rect 62127 52400 71000 52488
rect 57985 52010 59775 52200
rect 53490 52008 57700 52010
tri 57700 52008 57702 52010 sw
tri 57985 52008 57987 52010 ne
rect 57987 52008 59775 52010
rect 53490 51971 57702 52008
rect 48972 51952 53179 51971
tri 53179 51952 53198 51971 sw
tri 53490 51952 53509 51971 ne
rect 53509 51952 57702 51971
rect 48972 51925 53198 51952
rect 46714 51924 48685 51925
tri 48685 51924 48686 51925 sw
tri 48972 51924 48973 51925 ne
rect 48973 51924 53198 51925
rect 46714 51916 48686 51924
rect 44522 51836 46422 51916
rect 39989 51835 44229 51836
tri 44229 51835 44230 51836 sw
tri 44522 51835 44523 51836 ne
rect 44523 51835 46422 51836
rect 39989 51832 44230 51835
rect 35619 51831 39692 51832
tri 39692 51831 39693 51832 sw
tri 39989 51831 39990 51832 ne
rect 39990 51831 44230 51832
rect 35619 51661 39693 51831
rect 31143 51660 35331 51661
tri 35331 51660 35332 51661 sw
tri 35619 51660 35620 51661 ne
rect 35620 51660 39693 51661
rect 31143 51605 35332 51660
rect 26800 51410 30849 51605
tri 30849 51410 31044 51605 sw
tri 31143 51410 31338 51605 ne
rect 31338 51410 35332 51605
tri 26800 51320 26890 51410 ne
rect 26890 51320 31044 51410
tri 26600 51120 26800 51320 sw
tri 26890 51120 27090 51320 ne
rect 27090 51120 31044 51320
rect 25200 50941 26800 51120
tri 26800 50941 26979 51120 sw
tri 27090 50941 27269 51120 ne
rect 27269 51116 31044 51120
tri 31044 51116 31338 51410 sw
tri 31338 51116 31632 51410 ne
rect 31632 51372 35332 51410
tri 35332 51372 35620 51660 sw
tri 35620 51372 35908 51660 ne
rect 35908 51534 39693 51660
tri 39693 51534 39990 51831 sw
tri 39990 51534 40287 51831 ne
rect 40287 51542 44230 51831
tri 44230 51542 44523 51835 sw
tri 44523 51542 44816 51835 ne
rect 44816 51776 46422 51835
tri 46422 51776 46562 51916 sw
tri 46714 51776 46854 51916 ne
rect 46854 51776 48686 51916
rect 44816 51542 46562 51776
rect 40287 51534 44523 51542
rect 35908 51533 39990 51534
tri 39990 51533 39991 51534 sw
tri 40287 51533 40288 51534 ne
rect 40288 51533 44523 51534
rect 35908 51372 39991 51533
rect 31632 51220 35620 51372
tri 35620 51220 35772 51372 sw
tri 35908 51220 36060 51372 ne
rect 36060 51236 39991 51372
tri 39991 51236 40288 51533 sw
tri 40288 51236 40585 51533 ne
rect 40585 51249 44523 51533
tri 44523 51249 44816 51542 sw
tri 44816 51249 45109 51542 ne
rect 45109 51484 46562 51542
tri 46562 51484 46854 51776 sw
tri 46854 51484 47146 51776 ne
rect 47146 51637 48686 51776
tri 48686 51637 48973 51924 sw
tri 48973 51637 49260 51924 ne
rect 49260 51645 53198 51924
tri 53198 51645 53505 51952 sw
tri 53509 51645 53816 51952 ne
rect 53816 51723 57702 51952
tri 57702 51723 57987 52008 sw
tri 57987 51723 58272 52008 ne
rect 58272 51916 59775 52008
tri 59775 51916 60059 52200 sw
tri 60059 51916 60343 52200 ne
rect 60343 51916 71000 52200
rect 58272 51723 60059 51916
rect 53816 51722 57987 51723
tri 57987 51722 57988 51723 sw
tri 58272 51722 58273 51723 ne
rect 58273 51722 60059 51723
rect 53816 51645 57988 51722
rect 49260 51637 53505 51645
rect 47146 51484 48973 51637
rect 45109 51249 46854 51484
rect 40585 51236 44816 51249
rect 36060 51234 40288 51236
tri 40288 51234 40290 51236 sw
tri 40585 51234 40587 51236 ne
rect 40587 51234 44816 51236
rect 36060 51220 40290 51234
rect 31632 51116 35772 51220
rect 27269 50941 31338 51116
rect 25200 50740 26979 50941
tri 25200 50651 25289 50740 ne
rect 25289 50651 26979 50740
tri 26979 50651 27269 50941 sw
tri 27269 50651 27559 50941 ne
rect 27559 50926 31338 50941
tri 31338 50926 31528 51116 sw
tri 31632 50926 31822 51116 ne
rect 31822 50932 35772 51116
tri 35772 50932 36060 51220 sw
tri 36060 50932 36348 51220 ne
rect 36348 50937 40290 51220
tri 40290 50937 40587 51234 sw
tri 40587 50937 40884 51234 ne
rect 40884 50956 44816 51234
tri 44816 50956 45109 51249 sw
tri 45109 50956 45402 51249 ne
rect 45402 51192 46854 51249
tri 46854 51192 47146 51484 sw
tri 47146 51192 47438 51484 ne
rect 47438 51383 48973 51484
tri 48973 51383 49227 51637 sw
tri 49260 51383 49514 51637 ne
rect 49514 51383 53505 51637
rect 47438 51306 49227 51383
tri 49227 51306 49304 51383 sw
tri 49514 51306 49591 51383 ne
rect 49591 51353 53505 51383
tri 53505 51353 53797 51645 sw
tri 53816 51353 54108 51645 ne
rect 54108 51437 57988 51645
tri 57988 51437 58273 51722 sw
tri 58273 51437 58558 51722 ne
rect 58558 51632 60059 51722
tri 60059 51632 60343 51916 sw
tri 60343 51632 60627 51916 ne
rect 60627 51632 71000 51916
rect 58558 51452 60343 51632
tri 60343 51452 60523 51632 sw
tri 60627 51452 60807 51632 ne
rect 60807 51452 71000 51632
rect 58558 51437 60523 51452
rect 54108 51353 58273 51437
rect 49591 51306 53797 51353
tri 53797 51306 53844 51353 sw
tri 54108 51306 54155 51353 ne
rect 54155 51306 58273 51353
rect 47438 51192 49304 51306
rect 45402 50956 47146 51192
rect 40884 50937 45109 50956
rect 36348 50936 40587 50937
tri 40587 50936 40588 50937 sw
tri 40884 50936 40885 50937 ne
rect 40885 50936 45109 50937
rect 36348 50932 40588 50936
rect 31822 50926 36060 50932
rect 27559 50651 31528 50926
tri 25000 50362 25289 50651 sw
tri 25289 50362 25578 50651 ne
rect 25578 50650 27269 50651
tri 27269 50650 27270 50651 sw
tri 27559 50650 27560 50651 ne
rect 27560 50650 31528 50651
rect 25578 50362 27270 50650
rect 23600 50073 25289 50362
tri 25289 50073 25578 50362 sw
tri 25578 50073 25867 50362 ne
rect 25867 50360 27270 50362
tri 27270 50360 27560 50650 sw
tri 27560 50360 27850 50650 ne
rect 27850 50632 31528 50650
tri 31528 50632 31822 50926 sw
tri 31822 50632 32116 50926 ne
rect 32116 50792 36060 50926
tri 36060 50792 36200 50932 sw
tri 36348 50792 36488 50932 ne
rect 36488 50792 40588 50932
rect 32116 50632 36200 50792
rect 27850 50424 31822 50632
tri 31822 50424 32030 50632 sw
tri 32116 50424 32324 50632 ne
rect 32324 50504 36200 50632
tri 36200 50504 36488 50792 sw
tri 36488 50504 36776 50792 ne
rect 36776 50639 40588 50792
tri 40588 50639 40885 50936 sw
tri 40885 50639 41182 50936 ne
rect 41182 50901 45109 50936
tri 45109 50901 45164 50956 sw
tri 45402 50901 45457 50956 ne
rect 45457 50901 47146 50956
rect 41182 50639 45164 50901
rect 36776 50638 40885 50639
tri 40885 50638 40886 50639 sw
tri 41182 50638 41183 50639 ne
rect 41183 50638 45164 50639
rect 36776 50504 40886 50638
rect 32324 50424 36488 50504
rect 27850 50360 32030 50424
rect 25867 50359 27560 50360
tri 27560 50359 27561 50360 sw
tri 27850 50359 27851 50360 ne
rect 27851 50359 32030 50360
rect 25867 50073 27561 50359
rect 23600 50071 25578 50073
tri 23600 49974 23697 50071 ne
rect 23697 49974 25578 50071
tri 23400 49774 23600 49974 sw
tri 23697 49774 23897 49974 ne
rect 23897 49918 25578 49974
tri 25578 49918 25733 50073 sw
tri 25867 49918 26022 50073 ne
rect 26022 50069 27561 50073
tri 27561 50069 27851 50359 sw
tri 27851 50069 28141 50359 ne
rect 28141 50130 32030 50359
tri 32030 50130 32324 50424 sw
tri 32324 50130 32618 50424 ne
rect 32618 50261 36488 50424
tri 36488 50261 36731 50504 sw
tri 36776 50261 37019 50504 ne
rect 37019 50341 40886 50504
tri 40886 50341 41183 50638 sw
tri 41183 50341 41480 50638 ne
rect 41480 50608 45164 50638
tri 45164 50608 45457 50901 sw
tri 45457 50608 45750 50901 ne
rect 45750 50900 47146 50901
tri 47146 50900 47438 51192 sw
tri 47438 50900 47730 51192 ne
rect 47730 51019 49304 51192
tri 49304 51019 49591 51306 sw
tri 49591 51019 49878 51306 ne
rect 49878 51019 53844 51306
rect 47730 50900 49591 51019
rect 45750 50608 47438 50900
tri 47438 50608 47730 50900 sw
tri 47730 50608 48022 50900 ne
rect 48022 50807 49591 50900
tri 49591 50807 49803 51019 sw
tri 49878 50807 50090 51019 ne
rect 50090 51004 53844 51019
tri 53844 51004 54146 51306 sw
tri 54155 51004 54457 51306 ne
rect 54457 51175 58273 51306
tri 58273 51175 58535 51437 sw
tri 58558 51175 58820 51437 ne
rect 58820 51175 60523 51437
rect 54457 51004 58535 51175
rect 50090 50807 54146 51004
rect 48022 50608 49803 50807
rect 41480 50607 45457 50608
tri 45457 50607 45458 50608 sw
tri 45750 50607 45751 50608 ne
rect 45751 50607 47730 50608
rect 41480 50341 45458 50607
rect 37019 50261 41183 50341
rect 32618 50130 36731 50261
rect 28141 50069 32324 50130
rect 26022 49918 27851 50069
rect 23897 49774 25733 49918
rect 20400 49676 23600 49774
tri 23600 49676 23698 49774 sw
tri 23897 49676 23995 49774 ne
rect 23995 49676 25733 49774
rect 20400 49379 23698 49676
tri 23698 49379 23995 49676 sw
tri 23995 49379 24292 49676 ne
rect 24292 49629 25733 49676
tri 25733 49629 26022 49918 sw
tri 26022 49629 26311 49918 ne
rect 26311 49779 27851 49918
tri 27851 49779 28141 50069 sw
tri 28141 49779 28431 50069 ne
rect 28431 50044 32324 50069
tri 32324 50044 32410 50130 sw
tri 32618 50044 32704 50130 ne
rect 32704 50044 36731 50130
rect 28431 49779 32410 50044
rect 26311 49778 28141 49779
tri 28141 49778 28142 49779 sw
tri 28431 49778 28432 49779 ne
rect 28432 49778 32410 49779
rect 26311 49629 28142 49778
rect 24292 49379 26022 49629
rect 20400 49155 23995 49379
tri 23995 49155 24219 49379 sw
tri 24292 49155 24516 49379 ne
rect 24516 49340 26022 49379
tri 26022 49340 26311 49629 sw
tri 26311 49340 26600 49629 ne
rect 26600 49488 28142 49629
tri 28142 49488 28432 49778 sw
tri 28432 49488 28722 49778 ne
rect 28722 49750 32410 49778
tri 32410 49750 32704 50044 sw
tri 32704 49750 32998 50044 ne
rect 32998 49973 36731 50044
tri 36731 49973 37019 50261 sw
tri 37019 49973 37307 50261 ne
rect 37307 50122 41183 50261
tri 41183 50122 41402 50341 sw
tri 41480 50122 41699 50341 ne
rect 41699 50314 45458 50341
tri 45458 50314 45751 50607 sw
tri 45751 50314 46044 50607 ne
rect 46044 50520 47730 50607
tri 47730 50520 47818 50608 sw
tri 48022 50520 48110 50608 ne
rect 48110 50520 49803 50608
tri 49803 50520 50090 50807 sw
tri 50090 50520 50377 50807 ne
rect 50377 50703 54146 50807
tri 54146 50703 54447 51004 sw
tri 54457 50703 54758 51004 ne
rect 54758 50890 58535 51004
tri 58535 50890 58820 51175 sw
tri 58820 50890 59105 51175 ne
rect 59105 51168 60523 51175
tri 60523 51168 60807 51452 sw
tri 60807 51168 61091 51452 ne
rect 61091 51168 71000 51452
rect 59105 50890 60807 51168
rect 54758 50888 58820 50890
tri 58820 50888 58822 50890 sw
tri 59105 50888 59107 50890 ne
rect 59107 50888 60807 50890
rect 54758 50703 58822 50888
rect 50377 50520 54447 50703
rect 46044 50314 47818 50520
rect 41699 50313 45751 50314
tri 45751 50313 45752 50314 sw
tri 46044 50313 46045 50314 ne
rect 46045 50313 47818 50314
rect 41699 50122 45752 50313
rect 37307 49973 41402 50122
rect 32998 49888 37019 49973
tri 37019 49888 37104 49973 sw
tri 37307 49888 37392 49973 ne
rect 37392 49888 41402 49973
rect 32998 49750 37104 49888
rect 28722 49749 32704 49750
tri 32704 49749 32705 49750 sw
tri 32998 49749 32999 49750 ne
rect 32999 49749 37104 49750
rect 28722 49488 32705 49749
rect 26600 49340 28432 49488
rect 24516 49155 26311 49340
rect 20400 48858 24219 49155
tri 24219 48858 24516 49155 sw
tri 24516 48858 24813 49155 ne
rect 24813 49051 26311 49155
tri 26311 49051 26600 49340 sw
tri 26600 49051 26889 49340 ne
rect 26889 49251 28432 49340
tri 28432 49251 28669 49488 sw
tri 28722 49251 28959 49488 ne
rect 28959 49455 32705 49488
tri 32705 49455 32999 49749 sw
tri 32999 49455 33293 49749 ne
rect 33293 49600 37104 49749
tri 37104 49600 37392 49888 sw
tri 37392 49600 37680 49888 ne
rect 37680 49879 41402 49888
tri 41402 49879 41645 50122 sw
tri 41699 49879 41942 50122 ne
rect 41942 50020 45752 50122
tri 45752 50020 46045 50313 sw
tri 46045 50020 46338 50313 ne
rect 46338 50228 47818 50313
tri 47818 50228 48110 50520 sw
tri 48110 50228 48402 50520 ne
rect 48402 50519 50090 50520
tri 50090 50519 50091 50520 sw
tri 50377 50519 50378 50520 ne
rect 50378 50519 54447 50520
rect 48402 50232 50091 50519
tri 50091 50232 50378 50519 sw
tri 50378 50232 50665 50519 ne
rect 50665 50397 54447 50519
tri 54447 50397 54753 50703 sw
tri 54758 50397 55064 50703 ne
rect 55064 50603 58822 50703
tri 58822 50603 59107 50888 sw
tri 59107 50603 59392 50888 ne
rect 59392 50884 60807 50888
tri 60807 50884 61091 51168 sw
tri 61091 50884 61375 51168 ne
rect 61375 50884 71000 51168
rect 59392 50603 61091 50884
rect 55064 50602 59107 50603
tri 59107 50602 59108 50603 sw
tri 59392 50602 59393 50603 ne
rect 59393 50602 61091 50603
rect 55064 50397 59108 50602
rect 50665 50378 54753 50397
tri 54753 50378 54772 50397 sw
tri 55064 50378 55083 50397 ne
rect 55083 50378 59108 50397
rect 50665 50232 54772 50378
rect 48402 50228 50378 50232
rect 46338 50020 48110 50228
rect 41942 49879 46045 50020
rect 37680 49824 41645 49879
tri 41645 49824 41700 49879 sw
tri 41942 49824 41997 49879 ne
rect 41997 49824 46045 49879
rect 37680 49600 41700 49824
rect 33293 49455 37392 49600
rect 28959 49454 32999 49455
tri 32999 49454 33000 49455 sw
tri 33293 49454 33294 49455 ne
rect 33294 49454 37392 49455
rect 28959 49251 33000 49454
rect 26889 49051 28669 49251
rect 24813 49049 26600 49051
tri 26600 49049 26602 49051 sw
tri 26889 49049 26891 49051 ne
rect 26891 49049 28669 49051
rect 24813 48858 26602 49049
rect 20400 48730 24516 48858
tri 20400 48648 20482 48730 ne
rect 20482 48648 24516 48730
tri 20200 48366 20482 48648 sw
tri 20482 48366 20764 48648 ne
rect 20764 48561 24516 48648
tri 24516 48561 24813 48858 sw
tri 24813 48561 25110 48858 ne
rect 25110 48760 26602 48858
tri 26602 48760 26891 49049 sw
tri 26891 48760 27180 49049 ne
rect 27180 48961 28669 49049
tri 28669 48961 28959 49251 sw
tri 28959 48961 29249 49251 ne
rect 29249 49160 33000 49251
tri 33000 49160 33294 49454 sw
tri 33294 49160 33588 49454 ne
rect 33588 49393 37392 49454
tri 37392 49393 37599 49600 sw
tri 37680 49393 37887 49600 ne
rect 37887 49527 41700 49600
tri 41700 49527 41997 49824 sw
tri 41997 49527 42294 49824 ne
rect 42294 49727 46045 49824
tri 46045 49727 46338 50020 sw
tri 46338 49727 46631 50020 ne
rect 46631 49936 48110 50020
tri 48110 49936 48402 50228 sw
tri 48402 49936 48694 50228 ne
rect 48694 50042 50378 50228
tri 50378 50042 50568 50232 sw
tri 50665 50042 50855 50232 ne
rect 50855 50072 54772 50232
tri 54772 50072 55078 50378 sw
tri 55083 50072 55389 50378 ne
rect 55389 50317 59108 50378
tri 59108 50317 59393 50602 sw
tri 59393 50317 59678 50602 ne
rect 59678 50600 61091 50602
tri 61091 50600 61375 50884 sw
tri 61375 50800 61459 50884 ne
rect 61459 50800 71000 50884
rect 59678 50317 71000 50600
rect 55389 50249 59393 50317
tri 59393 50249 59461 50317 sw
tri 59678 50249 59746 50317 ne
rect 59746 50249 71000 50317
rect 55389 50072 59461 50249
rect 50855 50042 55078 50072
rect 48694 49936 50568 50042
rect 46631 49796 48402 49936
tri 48402 49796 48542 49936 sw
tri 48694 49796 48834 49936 ne
rect 48834 49796 50568 49936
rect 46631 49727 48542 49796
rect 42294 49527 46338 49727
rect 37887 49525 41997 49527
tri 41997 49525 41999 49527 sw
tri 42294 49525 42296 49527 ne
rect 42296 49525 46338 49527
rect 37887 49393 41999 49525
rect 33588 49160 37599 49393
rect 29249 49159 33294 49160
tri 33294 49159 33295 49160 sw
tri 33588 49159 33589 49160 ne
rect 33589 49159 37599 49160
rect 29249 48961 33295 49159
rect 27180 48760 28959 48961
rect 25110 48561 26891 48760
rect 20764 48374 24813 48561
tri 24813 48374 25000 48561 sw
tri 25110 48374 25297 48561 ne
rect 25297 48471 26891 48561
tri 26891 48471 27180 48760 sw
tri 27180 48471 27469 48760 ne
rect 27469 48671 28959 48760
tri 28959 48671 29249 48961 sw
tri 29249 48671 29539 48961 ne
rect 29539 48865 33295 48961
tri 33295 48865 33589 49159 sw
tri 33589 48865 33883 49159 ne
rect 33883 49105 37599 49159
tri 37599 49105 37887 49393 sw
tri 37887 49105 38175 49393 ne
rect 38175 49228 41999 49393
tri 41999 49228 42296 49525 sw
tri 42296 49228 42593 49525 ne
rect 42593 49508 46338 49525
tri 46338 49508 46557 49727 sw
tri 46631 49508 46850 49727 ne
rect 46850 49508 48542 49727
rect 42593 49228 46557 49508
rect 38175 49227 42296 49228
tri 42296 49227 42297 49228 sw
tri 42593 49227 42594 49228 ne
rect 42594 49227 46557 49228
rect 38175 49105 42297 49227
rect 33883 48929 37887 49105
tri 37887 48929 38063 49105 sw
tri 38175 48929 38351 49105 ne
rect 38351 48930 42297 49105
tri 42297 48930 42594 49227 sw
tri 42594 48930 42891 49227 ne
rect 42891 49215 46557 49227
tri 46557 49215 46850 49508 sw
tri 46850 49215 47143 49508 ne
rect 47143 49504 48542 49508
tri 48542 49504 48834 49796 sw
tri 48834 49504 49126 49796 ne
rect 49126 49755 50568 49796
tri 50568 49755 50855 50042 sw
tri 50855 49755 51142 50042 ne
rect 51142 49938 55078 50042
tri 55078 49938 55212 50072 sw
tri 55389 49938 55523 50072 ne
rect 55523 49964 59461 50072
tri 59461 49964 59746 50249 sw
tri 59746 49964 60031 50249 ne
rect 60031 49964 71000 50249
rect 55523 49938 59746 49964
rect 51142 49755 55212 49938
rect 49126 49504 50855 49755
rect 47143 49215 48834 49504
rect 42891 48930 46850 49215
rect 38351 48929 42594 48930
rect 33883 48865 38063 48929
rect 29539 48864 33589 48865
tri 33589 48864 33590 48865 sw
tri 33883 48864 33884 48865 ne
rect 33884 48864 38063 48865
rect 29539 48671 33590 48864
rect 27469 48670 29249 48671
tri 29249 48670 29250 48671 sw
tri 29539 48670 29540 48671 ne
rect 29540 48670 33590 48671
rect 27469 48471 29250 48670
rect 25297 48380 27180 48471
tri 27180 48380 27271 48471 sw
tri 27469 48380 27560 48471 ne
rect 27560 48380 29250 48471
tri 29250 48380 29540 48670 sw
tri 29540 48380 29830 48670 ne
rect 29830 48570 33590 48670
tri 33590 48570 33884 48864 sw
tri 33884 48570 34178 48864 ne
rect 34178 48641 38063 48864
tri 38063 48641 38351 48929 sw
tri 38351 48641 38639 48929 ne
rect 38639 48835 42594 48929
tri 42594 48835 42689 48930 sw
tri 42891 48835 42986 48930 ne
rect 42986 48922 46850 48930
tri 46850 48922 47143 49215 sw
tri 47143 48922 47436 49215 ne
rect 47436 49212 48834 49215
tri 48834 49212 49126 49504 sw
tri 49126 49212 49418 49504 ne
rect 49418 49468 50855 49504
tri 50855 49468 51142 49755 sw
tri 51142 49468 51429 49755 ne
rect 51429 49636 55212 49755
tri 55212 49636 55514 49938 sw
tri 55523 49636 55825 49938 ne
rect 55825 49743 59746 49938
tri 59746 49743 59967 49964 sw
tri 60031 49743 60252 49964 ne
rect 60252 49743 71000 49964
rect 55825 49636 59967 49743
rect 51429 49468 55514 49636
rect 49418 49402 51142 49468
tri 51142 49402 51208 49468 sw
tri 51429 49402 51495 49468 ne
rect 51495 49402 55514 49468
tri 55514 49402 55748 49636 sw
tri 55825 49402 56059 49636 ne
rect 56059 49575 59967 49636
tri 59967 49575 60135 49743 sw
tri 60252 49575 60420 49743 ne
rect 60420 49575 71000 49743
rect 56059 49402 60135 49575
rect 49418 49212 51208 49402
rect 47436 48922 49126 49212
rect 42986 48920 47143 48922
tri 47143 48920 47145 48922 sw
tri 47436 48920 47438 48922 ne
rect 47438 48920 49126 48922
tri 49126 48920 49418 49212 sw
tri 49418 48920 49710 49212 ne
rect 49710 49115 51208 49212
tri 51208 49115 51495 49402 sw
tri 51495 49115 51782 49402 ne
rect 51782 49115 55748 49402
rect 49710 48920 51495 49115
rect 42986 48835 47145 48920
rect 38639 48641 42689 48835
rect 34178 48640 38351 48641
tri 38351 48640 38352 48641 sw
tri 38639 48640 38640 48641 ne
rect 38640 48640 42689 48641
rect 34178 48570 38352 48640
rect 29830 48568 33884 48570
tri 33884 48568 33886 48570 sw
tri 34178 48568 34180 48570 ne
rect 34180 48568 38352 48570
rect 29830 48380 33886 48568
rect 25297 48374 27271 48380
rect 20764 48366 25000 48374
rect 17200 48166 20482 48366
tri 20482 48166 20682 48366 sw
tri 20764 48166 20964 48366 ne
rect 20964 48166 25000 48366
rect 17200 48082 20682 48166
tri 20682 48082 20766 48166 sw
tri 20964 48082 21048 48166 ne
rect 21048 48082 25000 48166
rect 17200 47800 20766 48082
tri 20766 47800 21048 48082 sw
tri 21048 47800 21330 48082 ne
rect 21330 48077 25000 48082
tri 25000 48077 25297 48374 sw
tri 25297 48077 25594 48374 ne
rect 25594 48091 27271 48374
tri 27271 48091 27560 48380 sw
tri 27560 48091 27849 48380 ne
rect 27849 48379 29540 48380
tri 29540 48379 29541 48380 sw
tri 29830 48379 29831 48380 ne
rect 29831 48379 33886 48380
rect 27849 48091 29541 48379
rect 25594 48077 27560 48091
rect 21330 48076 25297 48077
tri 25297 48076 25298 48077 sw
tri 25594 48076 25595 48077 ne
rect 25595 48076 27560 48077
rect 21330 47800 25298 48076
rect 17200 47798 21048 47800
tri 21048 47798 21050 47800 sw
tri 21330 47798 21332 47800 ne
rect 21332 47798 25298 47800
rect 17200 47516 21050 47798
tri 21050 47516 21332 47798 sw
tri 21332 47516 21614 47798 ne
rect 21614 47779 25298 47798
tri 25298 47779 25595 48076 sw
tri 25595 47779 25892 48076 ne
rect 25892 47802 27560 48076
tri 27560 47802 27849 48091 sw
tri 27849 47802 28138 48091 ne
rect 28138 48089 29541 48091
tri 29541 48089 29831 48379 sw
tri 29831 48089 30121 48379 ne
rect 30121 48274 33886 48379
tri 33886 48274 34180 48568 sw
tri 34180 48274 34474 48568 ne
rect 34474 48352 38352 48568
tri 38352 48352 38640 48640 sw
tri 38640 48352 38928 48640 ne
rect 38928 48538 42689 48640
tri 42689 48538 42986 48835 sw
tri 42986 48538 43283 48835 ne
rect 43283 48627 47145 48835
tri 47145 48627 47438 48920 sw
tri 47438 48627 47731 48920 ne
rect 47731 48628 49418 48920
tri 49418 48628 49710 48920 sw
tri 49710 48628 50002 48920 ne
rect 50002 48828 51495 48920
tri 51495 48828 51782 49115 sw
tri 51782 48828 52069 49115 ne
rect 52069 49096 55748 49115
tri 55748 49096 56054 49402 sw
tri 56059 49096 56365 49402 ne
rect 56365 49290 60135 49402
tri 60135 49290 60420 49575 sw
tri 60420 49290 60705 49575 ne
rect 60705 49290 71000 49575
rect 56365 49288 60420 49290
tri 60420 49288 60422 49290 sw
tri 60705 49288 60707 49290 ne
rect 60707 49288 71000 49290
rect 56365 49096 60422 49288
rect 52069 49010 56054 49096
tri 56054 49010 56140 49096 sw
tri 56365 49010 56451 49096 ne
rect 56451 49010 60422 49096
rect 52069 48828 56140 49010
rect 50002 48827 51782 48828
tri 51782 48827 51783 48828 sw
tri 52069 48827 52070 48828 ne
rect 52070 48827 56140 48828
rect 50002 48628 51783 48827
rect 47731 48627 49710 48628
rect 43283 48538 47438 48627
rect 38928 48352 42986 48538
rect 34474 48351 38640 48352
tri 38640 48351 38641 48352 sw
tri 38928 48351 38929 48352 ne
rect 38929 48351 42986 48352
rect 34474 48274 38641 48351
rect 30121 48089 34180 48274
rect 28138 48020 29831 48089
tri 29831 48020 29900 48089 sw
tri 30121 48020 30190 48089 ne
rect 30190 48020 34180 48089
tri 34180 48020 34434 48274 sw
tri 34474 48020 34728 48274 ne
rect 34728 48063 38641 48274
tri 38641 48063 38929 48351 sw
tri 38929 48063 39217 48351 ne
rect 39217 48333 42986 48351
tri 42986 48333 43191 48538 sw
tri 43283 48333 43488 48538 ne
rect 43488 48334 47438 48538
tri 47438 48334 47731 48627 sw
tri 47731 48334 48024 48627 ne
rect 48024 48540 49710 48627
tri 49710 48540 49798 48628 sw
tri 50002 48540 50090 48628 ne
rect 50090 48540 51783 48628
tri 51783 48540 52070 48827 sw
tri 52070 48540 52357 48827 ne
rect 52357 48704 56140 48827
tri 56140 48704 56446 49010 sw
tri 56451 48704 56757 49010 ne
rect 56757 49003 60422 49010
tri 60422 49003 60707 49288 sw
tri 60707 49200 60795 49288 ne
rect 60795 49200 71000 49288
rect 56757 49000 60707 49003
tri 60707 49000 60710 49003 sw
rect 56757 48704 71000 49000
rect 52357 48684 56446 48704
tri 56446 48684 56466 48704 sw
tri 56757 48684 56777 48704 ne
rect 56777 48684 71000 48704
rect 52357 48540 56466 48684
rect 48024 48334 49798 48540
rect 43488 48333 47731 48334
rect 39217 48063 43191 48333
rect 34728 48061 38929 48063
tri 38929 48061 38931 48063 sw
tri 39217 48061 39219 48063 ne
rect 39219 48061 43191 48063
rect 34728 48020 38931 48061
rect 28138 47802 29900 48020
rect 25892 47779 27849 47802
rect 21614 47516 25595 47779
rect 17200 47515 21332 47516
tri 21332 47515 21333 47516 sw
tri 21614 47515 21615 47516 ne
rect 21615 47515 25595 47516
rect 17200 47404 21333 47515
tri 17200 47312 17292 47404 ne
rect 17292 47312 21333 47404
tri 17000 47020 17292 47312 sw
tri 17292 47020 17584 47312 ne
rect 17584 47233 21333 47312
tri 21333 47233 21615 47515 sw
tri 21615 47233 21897 47515 ne
rect 21897 47482 25595 47515
tri 25595 47482 25892 47779 sw
tri 25892 47482 26189 47779 ne
rect 26189 47647 27849 47779
tri 27849 47647 28004 47802 sw
tri 28138 47647 28293 47802 ne
rect 28293 47730 29900 47802
tri 29900 47730 30190 48020 sw
tri 30190 47730 30480 48020 ne
rect 30480 47730 34434 48020
rect 28293 47647 30190 47730
rect 26189 47482 28004 47647
rect 21897 47376 25892 47482
tri 25892 47376 25998 47482 sw
tri 26189 47376 26295 47482 ne
rect 26295 47376 28004 47482
rect 21897 47233 25998 47376
rect 17584 47232 21615 47233
tri 21615 47232 21616 47233 sw
tri 21897 47232 21898 47233 ne
rect 21898 47232 25998 47233
rect 17584 47020 21616 47232
rect 14000 46820 17292 47020
tri 17292 46820 17492 47020 sw
tri 17584 46820 17784 47020 ne
rect 17784 46950 21616 47020
tri 21616 46950 21898 47232 sw
tri 21898 46950 22180 47232 ne
rect 22180 47079 25998 47232
tri 25998 47079 26295 47376 sw
tri 26295 47079 26592 47376 ne
rect 26592 47358 28004 47376
tri 28004 47358 28293 47647 sw
tri 28293 47358 28582 47647 ne
rect 28582 47508 30190 47647
tri 30190 47508 30412 47730 sw
tri 30480 47508 30702 47730 ne
rect 30702 47726 34434 47730
tri 34434 47726 34728 48020 sw
tri 34728 47726 35022 48020 ne
rect 35022 47773 38931 48020
tri 38931 47773 39219 48061 sw
tri 39219 47773 39507 48061 ne
rect 39507 48036 43191 48061
tri 43191 48036 43488 48333 sw
tri 43488 48036 43785 48333 ne
rect 43785 48180 47731 48333
tri 47731 48180 47885 48334 sw
tri 48024 48180 48178 48334 ne
rect 48178 48248 49798 48334
tri 49798 48248 50090 48540 sw
tri 50090 48248 50382 48540 ne
rect 50382 48539 52070 48540
tri 52070 48539 52071 48540 sw
tri 52357 48539 52358 48540 ne
rect 52358 48539 56466 48540
rect 50382 48252 52071 48539
tri 52071 48252 52358 48539 sw
tri 52358 48252 52645 48539 ne
rect 52645 48378 56466 48539
tri 56466 48378 56772 48684 sw
tri 56777 48378 57083 48684 ne
rect 57083 48378 71000 48684
rect 52645 48359 56772 48378
tri 56772 48359 56791 48378 sw
tri 57083 48359 57102 48378 ne
rect 57102 48359 71000 48378
rect 52645 48252 56791 48359
rect 50382 48248 52358 48252
rect 48178 48180 50090 48248
rect 43785 48036 47885 48180
rect 39507 47886 43488 48036
tri 43488 47886 43638 48036 sw
tri 43785 47886 43935 48036 ne
rect 43935 47887 47885 48036
tri 47885 47887 48178 48180 sw
tri 48178 47887 48471 48180 ne
rect 48471 47956 50090 48180
tri 50090 47956 50382 48248 sw
tri 50382 47956 50674 48248 ne
rect 50674 47965 52358 48248
tri 52358 47965 52645 48252 sw
tri 52645 47965 52932 48252 ne
rect 52932 48053 56791 48252
tri 56791 48053 57097 48359 sw
tri 57102 48053 57408 48359 ne
rect 57408 48053 71000 48359
rect 52932 48034 57097 48053
tri 57097 48034 57116 48053 sw
tri 57408 48034 57427 48053 ne
rect 57427 48034 71000 48053
rect 52932 47965 57116 48034
rect 50674 47964 52645 47965
tri 52645 47964 52646 47965 sw
tri 52932 47964 52933 47965 ne
rect 52933 47964 57116 47965
rect 50674 47956 52646 47964
rect 48471 47887 50382 47956
rect 43935 47886 48178 47887
tri 48178 47886 48179 47887 sw
tri 48471 47886 48472 47887 ne
rect 48472 47886 50382 47887
rect 39507 47773 43638 47886
rect 35022 47772 39219 47773
tri 39219 47772 39220 47773 sw
tri 39507 47772 39508 47773 ne
rect 39508 47772 43638 47773
rect 35022 47726 39220 47772
rect 30702 47657 34728 47726
tri 34728 47657 34797 47726 sw
tri 35022 47657 35091 47726 ne
rect 35091 47657 39220 47726
rect 30702 47508 34797 47657
rect 28582 47358 30412 47508
rect 26592 47079 28293 47358
rect 22180 47078 26295 47079
tri 26295 47078 26296 47079 sw
tri 26592 47078 26593 47079 ne
rect 26593 47078 28293 47079
rect 22180 46950 26296 47078
rect 17784 46820 21898 46950
rect 14000 46616 17492 46820
tri 17492 46616 17696 46820 sw
tri 17784 46616 17988 46820 ne
rect 17988 46790 21898 46820
tri 21898 46790 22058 46950 sw
tri 22180 46790 22340 46950 ne
rect 22340 46790 26296 46950
rect 17988 46626 22058 46790
tri 22058 46626 22222 46790 sw
tri 22340 46626 22504 46790 ne
rect 22504 46781 26296 46790
tri 26296 46781 26593 47078 sw
tri 26593 46781 26890 47078 ne
rect 26890 47069 28293 47078
tri 28293 47069 28582 47358 sw
tri 28582 47069 28871 47358 ne
rect 28871 47352 30412 47358
tri 30412 47352 30568 47508 sw
tri 30702 47352 30858 47508 ne
rect 30858 47363 34797 47508
tri 34797 47363 35091 47657 sw
tri 35091 47363 35385 47657 ne
rect 35385 47484 39220 47657
tri 39220 47484 39508 47772 sw
tri 39508 47484 39796 47772 ne
rect 39796 47589 43638 47772
tri 43638 47589 43935 47886 sw
tri 43935 47589 44232 47886 ne
rect 44232 47593 48179 47886
tri 48179 47593 48472 47886 sw
tri 48472 47593 48765 47886 ne
rect 48765 47816 50382 47886
tri 50382 47816 50522 47956 sw
tri 50674 47816 50814 47956 ne
rect 50814 47816 52646 47956
rect 48765 47593 50522 47816
rect 44232 47589 48472 47593
rect 39796 47588 43935 47589
tri 43935 47588 43936 47589 sw
tri 44232 47588 44233 47589 ne
rect 44233 47588 48472 47589
rect 39796 47484 43936 47588
rect 35385 47483 39508 47484
tri 39508 47483 39509 47484 sw
tri 39796 47483 39797 47484 ne
rect 39797 47483 43936 47484
rect 35385 47363 39509 47483
rect 30858 47362 35091 47363
tri 35091 47362 35092 47363 sw
tri 35385 47362 35386 47363 ne
rect 35386 47362 39509 47363
rect 30858 47352 35092 47362
rect 28871 47069 30568 47352
rect 26890 46781 28582 47069
rect 22504 46626 26593 46781
rect 17988 46616 22222 46626
rect 14000 46324 17696 46616
tri 17696 46324 17988 46616 sw
tri 17988 46324 18280 46616 ne
rect 18280 46507 22222 46616
tri 22222 46507 22341 46626 sw
tri 22504 46507 22623 46626 ne
rect 22623 46507 26593 46626
rect 18280 46324 22341 46507
rect 14000 46114 17988 46324
tri 17988 46114 18198 46324 sw
tri 18280 46114 18490 46324 ne
rect 18490 46225 22341 46324
tri 22341 46225 22623 46507 sw
tri 22623 46225 22905 46507 ne
rect 22905 46484 26593 46507
tri 26593 46484 26890 46781 sw
tri 26890 46484 27187 46781 ne
rect 27187 46780 28582 46781
tri 28582 46780 28871 47069 sw
tri 28871 46780 29160 47069 ne
rect 29160 47062 30568 47069
tri 30568 47062 30858 47352 sw
tri 30858 47062 31148 47352 ne
rect 31148 47068 35092 47352
tri 35092 47068 35386 47362 sw
tri 35386 47068 35680 47362 ne
rect 35680 47195 39509 47362
tri 39509 47195 39797 47483 sw
tri 39797 47195 40085 47483 ne
rect 40085 47291 43936 47483
tri 43936 47291 44233 47588 sw
tri 44233 47291 44530 47588 ne
rect 44530 47300 48472 47588
tri 48472 47300 48765 47593 sw
tri 48765 47300 49058 47593 ne
rect 49058 47524 50522 47593
tri 50522 47524 50814 47816 sw
tri 50814 47524 51106 47816 ne
rect 51106 47677 52646 47816
tri 52646 47677 52933 47964 sw
tri 52933 47677 53220 47964 ne
rect 53220 47728 57116 47964
tri 57116 47728 57422 48034 sw
tri 57427 47728 57733 48034 ne
rect 57733 47728 71000 48034
rect 53220 47709 57422 47728
tri 57422 47709 57441 47728 sw
tri 57733 47709 57752 47728 ne
rect 57752 47709 71000 47728
rect 53220 47677 57441 47709
rect 51106 47524 52933 47677
rect 49058 47300 50814 47524
rect 44530 47299 48765 47300
tri 48765 47299 48766 47300 sw
tri 49058 47299 49059 47300 ne
rect 49059 47299 50814 47300
rect 44530 47291 48766 47299
rect 40085 47290 44233 47291
tri 44233 47290 44234 47291 sw
tri 44530 47290 44531 47291 ne
rect 44531 47290 48766 47291
rect 40085 47195 44234 47290
rect 35680 47068 39797 47195
rect 31148 47067 35386 47068
tri 35386 47067 35387 47068 sw
tri 35680 47067 35681 47068 ne
rect 35681 47067 39797 47068
rect 31148 47062 35387 47067
rect 29160 47061 30858 47062
tri 30858 47061 30859 47062 sw
tri 31148 47061 31149 47062 ne
rect 31149 47061 35387 47062
rect 29160 46780 30859 47061
rect 27187 46491 28871 46780
tri 28871 46491 29160 46780 sw
tri 29160 46491 29449 46780 ne
rect 29449 46771 30859 46780
tri 30859 46771 31149 47061 sw
tri 31149 46771 31439 47061 ne
rect 31439 46773 35387 47061
tri 35387 46773 35681 47067 sw
tri 35681 46773 35975 47067 ne
rect 35975 46976 39797 47067
tri 39797 46976 40016 47195 sw
tri 40085 46976 40304 47195 ne
rect 40304 46993 44234 47195
tri 44234 46993 44531 47290 sw
tri 44531 46993 44828 47290 ne
rect 44828 47006 48766 47290
tri 48766 47006 49059 47299 sw
tri 49059 47006 49352 47299 ne
rect 49352 47232 50814 47299
tri 50814 47232 51106 47524 sw
tri 51106 47232 51398 47524 ne
rect 51398 47422 52933 47524
tri 52933 47422 53188 47677 sw
tri 53220 47422 53475 47677 ne
rect 53475 47422 57441 47677
rect 51398 47232 53188 47422
rect 49352 47006 51106 47232
rect 44828 46993 49059 47006
rect 40304 46992 44531 46993
tri 44531 46992 44532 46993 sw
tri 44828 46992 44829 46993 ne
rect 44829 46992 49059 46993
rect 40304 46976 44532 46992
rect 35975 46773 40016 46976
rect 31439 46771 35681 46773
rect 29449 46690 31149 46771
tri 31149 46690 31230 46771 sw
tri 31439 46690 31520 46771 ne
rect 31520 46690 35681 46771
rect 29449 46491 31230 46690
rect 27187 46484 29160 46491
rect 22905 46483 26890 46484
tri 26890 46483 26891 46484 sw
tri 27187 46483 27188 46484 ne
rect 27188 46483 29160 46484
rect 22905 46225 26891 46483
rect 18490 46224 22623 46225
tri 22623 46224 22624 46225 sw
tri 22905 46224 22906 46225 ne
rect 22906 46224 26891 46225
rect 18490 46114 22624 46224
rect 14000 46068 18198 46114
tri 14000 43708 16360 46068 ne
rect 16360 45822 18198 46068
tri 18198 45822 18490 46114 sw
tri 18490 45822 18782 46114 ne
rect 18782 45942 22624 46114
tri 22624 45942 22906 46224 sw
tri 22906 45942 23188 46224 ne
rect 23188 46186 26891 46224
tri 26891 46186 27188 46483 sw
tri 27188 46186 27485 46483 ne
rect 27485 46400 29160 46483
tri 29160 46400 29251 46491 sw
tri 29449 46400 29540 46491 ne
rect 29540 46400 31230 46491
tri 31230 46400 31520 46690 sw
tri 31520 46400 31810 46690 ne
rect 31810 46682 35681 46690
tri 35681 46682 35772 46773 sw
tri 35975 46682 36066 46773 ne
rect 36066 46688 40016 46773
tri 40016 46688 40304 46976 sw
tri 40304 46688 40592 46976 ne
rect 40592 46695 44532 46976
tri 44532 46695 44829 46992 sw
tri 44829 46695 45126 46992 ne
rect 45126 46940 49059 46992
tri 49059 46940 49125 47006 sw
tri 49352 46940 49418 47006 ne
rect 49418 46940 51106 47006
tri 51106 46940 51398 47232 sw
tri 51398 46940 51690 47232 ne
rect 51690 47135 53188 47232
tri 53188 47135 53475 47422 sw
tri 53475 47135 53762 47422 ne
rect 53762 47402 57441 47422
tri 57441 47402 57748 47709 sw
tri 57752 47402 58059 47709 ne
rect 58059 47402 71000 47709
rect 53762 47135 57748 47402
rect 51690 47053 53475 47135
tri 53475 47053 53557 47135 sw
tri 53762 47053 53844 47135 ne
rect 53844 47110 57748 47135
tri 57748 47110 58040 47402 sw
tri 58059 47110 58351 47402 ne
rect 58351 47110 71000 47402
rect 53844 47053 58040 47110
tri 58040 47053 58097 47110 sw
tri 58351 47053 58408 47110 ne
rect 58408 47053 71000 47110
rect 51690 46940 53557 47053
rect 45126 46695 49125 46940
rect 40592 46693 44829 46695
tri 44829 46693 44831 46695 sw
tri 45126 46693 45128 46695 ne
rect 45128 46693 49125 46695
rect 40592 46688 44831 46693
rect 36066 46682 40304 46688
rect 31810 46400 35772 46682
rect 27485 46186 29251 46400
rect 23188 46185 27188 46186
tri 27188 46185 27189 46186 sw
tri 27485 46185 27486 46186 ne
rect 27486 46185 29251 46186
rect 23188 45942 27189 46185
rect 18782 45941 22906 45942
tri 22906 45941 22907 45942 sw
tri 23188 45941 23189 45942 ne
rect 23189 45941 27189 45942
rect 18782 45822 22907 45941
rect 16360 45821 18490 45822
tri 18490 45821 18491 45822 sw
tri 18782 45821 18783 45822 ne
rect 18783 45821 22907 45822
rect 16360 45529 18491 45821
tri 18491 45529 18783 45821 sw
tri 18783 45529 19075 45821 ne
rect 19075 45659 22907 45821
tri 22907 45659 23189 45941 sw
tri 23189 45659 23471 45941 ne
rect 23471 45888 27189 45941
tri 27189 45888 27486 46185 sw
tri 27486 45888 27783 46185 ne
rect 27783 46111 29251 46185
tri 29251 46111 29540 46400 sw
tri 29540 46111 29829 46400 ne
rect 29829 46399 31520 46400
tri 31520 46399 31521 46400 sw
tri 31810 46399 31811 46400 ne
rect 31811 46399 35772 46400
rect 29829 46111 31521 46399
rect 27783 45888 29540 46111
rect 23471 45804 27486 45888
tri 27486 45804 27570 45888 sw
tri 27783 45804 27867 45888 ne
rect 27867 45822 29540 45888
tri 29540 45822 29829 46111 sw
tri 29829 45822 30118 46111 ne
rect 30118 46109 31521 46111
tri 31521 46109 31811 46399 sw
tri 31811 46109 32101 46399 ne
rect 32101 46388 35772 46399
tri 35772 46388 36066 46682 sw
tri 36066 46388 36360 46682 ne
rect 36360 46597 40304 46682
tri 40304 46597 40395 46688 sw
tri 40592 46597 40683 46688 ne
rect 40683 46597 44831 46688
rect 36360 46388 40395 46597
rect 32101 46181 36066 46388
tri 36066 46181 36273 46388 sw
tri 36360 46181 36567 46388 ne
rect 36567 46309 40395 46388
tri 40395 46309 40683 46597 sw
tri 40683 46309 40971 46597 ne
rect 40971 46396 44831 46597
tri 44831 46396 45128 46693 sw
tri 45128 46396 45425 46693 ne
rect 45425 46647 49125 46693
tri 49125 46647 49418 46940 sw
tri 49418 46647 49711 46940 ne
rect 49711 46648 51398 46940
tri 51398 46648 51690 46940 sw
tri 51690 46648 51982 46940 ne
rect 51982 46766 53557 46940
tri 53557 46766 53844 47053 sw
tri 53844 46766 54131 47053 ne
rect 54131 46766 58097 47053
rect 51982 46648 53844 46766
rect 49711 46647 51690 46648
rect 45425 46396 49418 46647
rect 40971 46309 45128 46396
rect 36567 46307 40683 46309
tri 40683 46307 40685 46309 sw
tri 40971 46307 40973 46309 ne
rect 40973 46307 45128 46309
rect 36567 46181 40685 46307
rect 32101 46109 36273 46181
rect 30118 45822 31811 46109
rect 27867 45804 29829 45822
rect 23471 45659 27570 45804
rect 19075 45582 23189 45659
tri 23189 45582 23266 45659 sw
tri 23471 45582 23548 45659 ne
rect 23548 45582 27570 45659
rect 19075 45529 23266 45582
rect 16360 45527 18783 45529
tri 18783 45527 18785 45529 sw
tri 19075 45527 19077 45529 ne
rect 19077 45527 23266 45529
rect 16360 45236 18785 45527
tri 18785 45236 19076 45527 sw
tri 19077 45236 19368 45527 ne
rect 19368 45300 23266 45527
tri 23266 45300 23548 45582 sw
tri 23548 45300 23830 45582 ne
rect 23830 45507 27570 45582
tri 27570 45507 27867 45804 sw
tri 27867 45507 28164 45804 ne
rect 28164 45667 29829 45804
tri 29829 45667 29984 45822 sw
tri 30118 45667 30273 45822 ne
rect 30273 45819 31811 45822
tri 31811 45819 32101 46109 sw
tri 32101 45819 32391 46109 ne
rect 32391 45887 36273 46109
tri 36273 45887 36567 46181 sw
tri 36567 45887 36861 46181 ne
rect 36861 46019 40685 46181
tri 40685 46019 40973 46307 sw
tri 40973 46019 41261 46307 ne
rect 41261 46099 45128 46307
tri 45128 46099 45425 46396 sw
tri 45425 46099 45722 46396 ne
rect 45722 46354 49418 46396
tri 49418 46354 49711 46647 sw
tri 49711 46354 50004 46647 ne
rect 50004 46560 51690 46647
tri 51690 46560 51778 46648 sw
tri 51982 46560 52070 46648 ne
rect 52070 46560 53844 46648
rect 50004 46354 51778 46560
rect 45722 46353 49711 46354
tri 49711 46353 49712 46354 sw
tri 50004 46353 50005 46354 ne
rect 50005 46353 51778 46354
rect 45722 46099 49712 46353
rect 41261 46019 45425 46099
rect 36861 46018 40973 46019
tri 40973 46018 40974 46019 sw
tri 41261 46018 41262 46019 ne
rect 41262 46018 45425 46019
rect 36861 45887 40974 46018
rect 32391 45819 36567 45887
rect 30273 45818 32101 45819
tri 32101 45818 32102 45819 sw
tri 32391 45818 32392 45819 ne
rect 32392 45818 36567 45819
rect 30273 45667 32102 45818
rect 28164 45507 29984 45667
rect 23830 45300 27867 45507
rect 19368 45236 23548 45300
rect 16360 44992 19076 45236
tri 19076 44992 19320 45236 sw
tri 19368 44992 19612 45236 ne
rect 19612 45091 23548 45236
tri 23548 45091 23757 45300 sw
tri 23830 45091 24039 45300 ne
rect 24039 45210 27867 45300
tri 27867 45210 28164 45507 sw
tri 28164 45210 28461 45507 ne
rect 28461 45378 29984 45507
tri 29984 45378 30273 45667 sw
tri 30273 45378 30562 45667 ne
rect 30562 45528 32102 45667
tri 32102 45528 32392 45818 sw
tri 32392 45528 32682 45818 ne
rect 32682 45729 36567 45818
tri 36567 45729 36725 45887 sw
tri 36861 45729 37019 45887 ne
rect 37019 45730 40974 45887
tri 40974 45730 41262 46018 sw
tri 41262 45730 41550 46018 ne
rect 41550 45879 45425 46018
tri 45425 45879 45645 46099 sw
tri 45722 45879 45942 46099 ne
rect 45942 46060 49712 46099
tri 49712 46060 50005 46353 sw
tri 50005 46060 50298 46353 ne
rect 50298 46268 51778 46353
tri 51778 46268 52070 46560 sw
tri 52070 46268 52362 46560 ne
rect 52362 46559 53844 46560
tri 53844 46559 54051 46766 sw
tri 54131 46559 54338 46766 ne
rect 54338 46742 58097 46766
tri 58097 46742 58408 47053 sw
tri 58408 46742 58719 47053 ne
rect 58719 46742 71000 47053
rect 54338 46559 58408 46742
rect 52362 46272 54051 46559
tri 54051 46272 54338 46559 sw
tri 54338 46272 54625 46559 ne
rect 54625 46460 58408 46559
tri 58408 46460 58690 46742 sw
tri 58719 46460 59001 46742 ne
rect 59001 46460 71000 46742
rect 54625 46272 58690 46460
rect 52362 46268 54338 46272
rect 50298 46060 52070 46268
rect 45942 45879 50005 46060
rect 41550 45730 45645 45879
rect 37019 45729 41262 45730
rect 32682 45528 36725 45729
rect 30562 45378 32392 45528
rect 28461 45210 30273 45378
rect 24039 45091 28164 45210
rect 19612 44992 23757 45091
rect 16360 44700 19320 44992
tri 19320 44700 19612 44992 sw
tri 19612 44700 19904 44992 ne
rect 19904 44809 23757 44992
tri 23757 44809 24039 45091 sw
tri 24039 44809 24321 45091 ne
rect 24321 44913 28164 45091
tri 28164 44913 28461 45210 sw
tri 28461 44913 28758 45210 ne
rect 28758 45089 30273 45210
tri 30273 45089 30562 45378 sw
tri 30562 45089 30851 45378 ne
rect 30851 45291 32392 45378
tri 32392 45291 32629 45528 sw
tri 32682 45291 32919 45528 ne
rect 32919 45435 36725 45528
tri 36725 45435 37019 45729 sw
tri 37019 45435 37313 45729 ne
rect 37313 45644 41262 45729
tri 41262 45644 41348 45730 sw
tri 41550 45644 41636 45730 ne
rect 41636 45644 45645 45730
rect 37313 45435 41348 45644
rect 32919 45434 37019 45435
tri 37019 45434 37020 45435 sw
tri 37313 45434 37314 45435 ne
rect 37314 45434 41348 45435
rect 32919 45291 37020 45434
rect 30851 45089 32629 45291
rect 28758 44913 30562 45089
rect 24321 44912 28461 44913
tri 28461 44912 28462 44913 sw
tri 28758 44912 28759 44913 ne
rect 28759 44912 30562 44913
rect 24321 44809 28462 44912
rect 19904 44700 24039 44809
rect 16360 44698 19612 44700
tri 19612 44698 19614 44700 sw
tri 19904 44698 19906 44700 ne
rect 19906 44698 24039 44700
rect 16360 44406 19614 44698
tri 19614 44406 19906 44698 sw
tri 19906 44406 20198 44698 ne
rect 20198 44615 24039 44698
tri 24039 44615 24233 44809 sw
tri 24321 44615 24515 44809 ne
rect 24515 44615 28462 44809
tri 28462 44615 28759 44912 sw
tri 28759 44615 29056 44912 ne
rect 29056 44800 30562 44912
tri 30562 44800 30851 45089 sw
tri 30851 44800 31140 45089 ne
rect 31140 45001 32629 45089
tri 32629 45001 32919 45291 sw
tri 32919 45001 33209 45291 ne
rect 33209 45140 37020 45291
tri 37020 45140 37314 45434 sw
tri 37314 45140 37608 45434 ne
rect 37608 45356 41348 45434
tri 41348 45356 41636 45644 sw
tri 41636 45356 41924 45644 ne
rect 41924 45635 45645 45644
tri 45645 45635 45889 45879 sw
tri 45942 45635 46186 45879 ne
rect 46186 45767 50005 45879
tri 50005 45767 50298 46060 sw
tri 50298 45767 50591 46060 ne
rect 50591 45976 52070 46060
tri 52070 45976 52362 46268 sw
tri 52362 45976 52654 46268 ne
rect 52654 46087 54338 46268
tri 54338 46087 54523 46272 sw
tri 54625 46087 54810 46272 ne
rect 54810 46154 58690 46272
tri 58690 46154 58996 46460 sw
tri 59001 46154 59307 46460 ne
rect 59307 46154 71000 46460
rect 54810 46135 58996 46154
tri 58996 46135 59015 46154 sw
tri 59307 46135 59326 46154 ne
rect 59326 46135 71000 46154
rect 54810 46087 59015 46135
rect 52654 45976 54523 46087
rect 50591 45836 52362 45976
tri 52362 45836 52502 45976 sw
tri 52654 45836 52794 45976 ne
rect 52794 45836 54523 45976
rect 50591 45767 52502 45836
rect 46186 45635 50298 45767
rect 41924 45581 45889 45635
tri 45889 45581 45943 45635 sw
tri 46186 45581 46240 45635 ne
rect 46240 45581 50298 45635
rect 41924 45356 45943 45581
rect 37608 45151 41636 45356
tri 41636 45151 41841 45356 sw
tri 41924 45151 42129 45356 ne
rect 42129 45284 45943 45356
tri 45943 45284 46240 45581 sw
tri 46240 45284 46537 45581 ne
rect 46537 45548 50298 45581
tri 50298 45548 50517 45767 sw
tri 50591 45548 50810 45767 ne
rect 50810 45548 52502 45767
rect 46537 45284 50517 45548
rect 42129 45283 46240 45284
tri 46240 45283 46241 45284 sw
tri 46537 45283 46538 45284 ne
rect 46538 45283 50517 45284
rect 42129 45151 46241 45283
rect 37608 45140 41841 45151
rect 33209 45139 37314 45140
tri 37314 45139 37315 45140 sw
tri 37608 45139 37609 45140 ne
rect 37609 45139 41841 45140
rect 33209 45001 37315 45139
rect 31140 44800 32919 45001
rect 29056 44615 30851 44800
rect 20198 44406 24233 44615
rect 16360 44405 19906 44406
tri 19906 44405 19907 44406 sw
tri 20198 44405 20199 44406 ne
rect 20199 44405 24233 44406
rect 16360 44113 19907 44405
tri 19907 44113 20199 44405 sw
tri 20199 44113 20491 44405 ne
rect 20491 44333 24233 44405
tri 24233 44333 24515 44615 sw
tri 24515 44333 24797 44615 ne
rect 24797 44333 28759 44615
rect 20491 44331 24515 44333
tri 24515 44331 24517 44333 sw
tri 24797 44331 24799 44333 ne
rect 24799 44331 28759 44333
rect 20491 44113 24517 44331
rect 16360 44112 20199 44113
tri 20199 44112 20200 44113 sw
tri 20491 44112 20492 44113 ne
rect 20492 44112 24517 44113
rect 16360 43820 20200 44112
tri 20200 43820 20492 44112 sw
tri 20492 43820 20784 44112 ne
rect 20784 44049 24517 44112
tri 24517 44049 24799 44331 sw
tri 24799 44049 25081 44331 ne
rect 25081 44318 28759 44331
tri 28759 44318 29056 44615 sw
tri 29056 44318 29353 44615 ne
rect 29353 44511 30851 44615
tri 30851 44511 31140 44800 sw
tri 31140 44511 31429 44800 ne
rect 31429 44711 32919 44800
tri 32919 44711 33209 45001 sw
tri 33209 44711 33499 45001 ne
rect 33499 44845 37315 45001
tri 37315 44845 37609 45139 sw
tri 37609 44845 37903 45139 ne
rect 37903 44863 41841 45139
tri 41841 44863 42129 45151 sw
tri 42129 44863 42417 45151 ne
rect 42417 44986 46241 45151
tri 46241 44986 46538 45283 sw
tri 46538 44986 46835 45283 ne
rect 46835 45255 50517 45283
tri 50517 45255 50810 45548 sw
tri 50810 45255 51103 45548 ne
rect 51103 45544 52502 45548
tri 52502 45544 52794 45836 sw
tri 52794 45544 53086 45836 ne
rect 53086 45800 54523 45836
tri 54523 45800 54810 46087 sw
tri 54810 45800 55097 46087 ne
rect 55097 45829 59015 46087
tri 59015 45829 59321 46135 sw
tri 59326 46000 59461 46135 ne
rect 59461 46000 71000 46135
rect 55097 45800 59321 45829
tri 59321 45800 59350 45829 sw
rect 53086 45799 54810 45800
tri 54810 45799 54811 45800 sw
tri 55097 45799 55098 45800 ne
rect 55098 45799 71000 45800
rect 53086 45544 54811 45799
rect 51103 45255 52794 45544
rect 46835 45254 50810 45255
tri 50810 45254 50811 45255 sw
tri 51103 45254 51104 45255 ne
rect 51104 45254 52794 45255
rect 46835 44986 50811 45254
rect 42417 44984 46538 44986
tri 46538 44984 46540 44986 sw
tri 46835 44984 46837 44986 ne
rect 46837 44984 50811 44986
rect 42417 44863 46540 44984
rect 37903 44845 42129 44863
rect 33499 44843 37609 44845
tri 37609 44843 37611 44845 sw
tri 37903 44843 37905 44845 ne
rect 37905 44843 42129 44845
rect 33499 44711 37611 44843
rect 31429 44710 33209 44711
tri 33209 44710 33210 44711 sw
tri 33499 44710 33500 44711 ne
rect 33500 44710 37611 44711
rect 31429 44511 33210 44710
rect 29353 44420 31140 44511
tri 31140 44420 31231 44511 sw
tri 31429 44420 31520 44511 ne
rect 31520 44420 33210 44511
tri 33210 44420 33500 44710 sw
tri 33500 44420 33790 44710 ne
rect 33790 44549 37611 44710
tri 37611 44549 37905 44843 sw
tri 37905 44549 38199 44843 ne
rect 38199 44686 42129 44843
tri 42129 44686 42306 44863 sw
tri 42417 44686 42594 44863 ne
rect 42594 44688 46540 44863
tri 46540 44688 46836 44984 sw
tri 46837 44688 47133 44984 ne
rect 47133 44961 50811 44984
tri 50811 44961 51104 45254 sw
tri 51104 44961 51397 45254 ne
rect 51397 45252 52794 45254
tri 52794 45252 53086 45544 sw
tri 53086 45252 53378 45544 ne
rect 53378 45512 54811 45544
tri 54811 45512 55098 45799 sw
tri 55098 45512 55385 45799 ne
rect 55385 45512 71000 45799
rect 53378 45252 55098 45512
rect 51397 44961 53086 45252
rect 47133 44688 51104 44961
rect 42594 44686 46836 44688
rect 38199 44549 42306 44686
rect 33790 44548 37905 44549
tri 37905 44548 37906 44549 sw
tri 38199 44548 38200 44549 ne
rect 38200 44548 42306 44549
rect 33790 44420 37906 44548
rect 29353 44318 31231 44420
rect 25081 44317 29056 44318
tri 29056 44317 29057 44318 sw
tri 29353 44317 29354 44318 ne
rect 29354 44317 31231 44318
rect 25081 44049 29057 44317
rect 20784 44048 24799 44049
tri 24799 44048 24800 44049 sw
tri 25081 44048 25082 44049 ne
rect 25082 44048 29057 44049
rect 20784 43820 24800 44048
rect 16360 43708 20492 43820
tri 20492 43708 20604 43820 sw
tri 20784 43708 20896 43820 ne
rect 20896 43766 24800 43820
tri 24800 43766 25082 44048 sw
tri 25082 43766 25364 44048 ne
rect 25364 44020 29057 44048
tri 29057 44020 29354 44317 sw
tri 29354 44020 29651 44317 ne
rect 29651 44131 31231 44317
tri 31231 44131 31520 44420 sw
tri 31520 44131 31809 44420 ne
rect 31809 44419 33500 44420
tri 33500 44419 33501 44420 sw
tri 33790 44419 33791 44420 ne
rect 33791 44419 37906 44420
rect 31809 44131 33501 44419
rect 29651 44020 31520 44131
rect 25364 44019 29354 44020
tri 29354 44019 29355 44020 sw
tri 29651 44019 29652 44020 ne
rect 29652 44019 31520 44020
rect 25364 43766 29355 44019
rect 20896 43765 25082 43766
tri 25082 43765 25083 43766 sw
tri 25364 43765 25365 43766 ne
rect 25365 43765 29355 43766
rect 20896 43708 25083 43765
tri 16360 39464 20604 43708 ne
tri 20604 43416 20896 43708 sw
tri 20896 43416 21188 43708 ne
rect 21188 43483 25083 43708
tri 25083 43483 25365 43765 sw
tri 25365 43483 25647 43765 ne
rect 25647 43722 29355 43765
tri 29355 43722 29652 44019 sw
tri 29652 43722 29949 44019 ne
rect 29949 43842 31520 44019
tri 31520 43842 31809 44131 sw
tri 31809 43842 32098 44131 ne
rect 32098 44129 33501 44131
tri 33501 44129 33791 44419 sw
tri 33791 44129 34081 44419 ne
rect 34081 44254 37906 44419
tri 37906 44254 38200 44548 sw
tri 38200 44254 38494 44548 ne
rect 38494 44398 42306 44548
tri 42306 44398 42594 44686 sw
tri 42594 44398 42882 44686 ne
rect 42882 44591 46836 44686
tri 46836 44591 46933 44688 sw
tri 47133 44591 47230 44688 ne
rect 47230 44668 51104 44688
tri 51104 44668 51397 44961 sw
tri 51397 44668 51690 44961 ne
rect 51690 44960 53086 44961
tri 53086 44960 53378 45252 sw
tri 53378 44960 53670 45252 ne
rect 53670 45225 55098 45252
tri 55098 45225 55385 45512 sw
tri 55385 45225 55672 45512 ne
rect 55672 45225 71000 45512
rect 53670 45155 55385 45225
tri 55385 45155 55455 45225 sw
tri 55672 45155 55742 45225 ne
rect 55742 45155 71000 45225
rect 53670 44960 55455 45155
rect 51690 44668 53378 44960
tri 53378 44668 53670 44960 sw
tri 53670 44668 53962 44960 ne
rect 53962 44868 55455 44960
tri 55455 44868 55742 45155 sw
tri 55742 44868 56029 45155 ne
rect 56029 44868 71000 45155
rect 53962 44867 55742 44868
tri 55742 44867 55743 44868 sw
tri 56029 44867 56030 44868 ne
rect 56030 44867 71000 44868
rect 53962 44668 55743 44867
rect 47230 44666 51397 44668
tri 51397 44666 51399 44668 sw
tri 51690 44666 51692 44668 ne
rect 51692 44666 53670 44668
rect 47230 44591 51399 44666
rect 42882 44398 46933 44591
rect 38494 44397 42594 44398
tri 42594 44397 42595 44398 sw
tri 42882 44397 42883 44398 ne
rect 42883 44397 46933 44398
rect 38494 44254 42595 44397
rect 34081 44253 38200 44254
tri 38200 44253 38201 44254 sw
tri 38494 44253 38495 44254 ne
rect 38495 44253 42595 44254
rect 34081 44129 38201 44253
rect 32098 43842 33791 44129
rect 29949 43722 31809 43842
rect 25647 43483 29652 43722
rect 21188 43482 25365 43483
tri 25365 43482 25366 43483 sw
tri 25647 43482 25648 43483 ne
rect 25648 43482 29652 43483
rect 21188 43416 25366 43482
rect 20604 43233 20896 43416
tri 20896 43233 21079 43416 sw
tri 21188 43233 21371 43416 ne
rect 21371 43233 25366 43416
rect 20604 43044 21079 43233
tri 21079 43044 21268 43233 sw
tri 21371 43044 21560 43233 ne
rect 21560 43200 25366 43233
tri 25366 43200 25648 43482 sw
tri 25648 43200 25930 43482 ne
rect 25930 43425 29652 43482
tri 29652 43425 29949 43722 sw
tri 29949 43425 30246 43722 ne
rect 30246 43687 31809 43722
tri 31809 43687 31964 43842 sw
tri 32098 43687 32253 43842 ne
rect 32253 43839 33791 43842
tri 33791 43839 34081 44129 sw
tri 34081 43839 34371 44129 ne
rect 34371 43959 38201 44129
tri 38201 43959 38495 44253 sw
tri 38495 43959 38789 44253 ne
rect 38789 44109 42595 44253
tri 42595 44109 42883 44397 sw
tri 42883 44109 43171 44397 ne
rect 43171 44294 46933 44397
tri 46933 44294 47230 44591 sw
tri 47230 44294 47527 44591 ne
rect 47527 44373 51399 44591
tri 51399 44373 51692 44666 sw
tri 51692 44373 51985 44666 ne
rect 51985 44580 53670 44666
tri 53670 44580 53758 44668 sw
tri 53962 44580 54050 44668 ne
rect 54050 44580 55743 44668
tri 55743 44580 56030 44867 sw
tri 56030 44580 56317 44867 ne
rect 56317 44580 71000 44867
rect 51985 44373 53758 44580
rect 47527 44294 51692 44373
rect 43171 44109 47230 44294
rect 38789 44108 42883 44109
tri 42883 44108 42884 44109 sw
tri 43171 44108 43172 44109 ne
rect 43172 44108 47230 44109
rect 38789 43959 42884 44108
rect 34371 43839 38495 43959
rect 32253 43776 34081 43839
tri 34081 43776 34144 43839 sw
tri 34371 43776 34434 43839 ne
rect 34434 43776 38495 43839
rect 32253 43687 34144 43776
rect 30246 43425 31964 43687
rect 25930 43416 29949 43425
tri 29949 43416 29958 43425 sw
tri 30246 43416 30255 43425 ne
rect 30255 43416 31964 43425
rect 25930 43200 29958 43416
rect 21560 43199 25648 43200
tri 25648 43199 25649 43200 sw
tri 25930 43199 25931 43200 ne
rect 25931 43199 29958 43200
rect 21560 43044 25649 43199
rect 20604 42752 21268 43044
tri 21268 42752 21560 43044 sw
tri 21560 42752 21852 43044 ne
rect 21852 42917 25649 43044
tri 25649 42917 25931 43199 sw
tri 25931 42917 26213 43199 ne
rect 26213 43119 29958 43199
tri 29958 43119 30255 43416 sw
tri 30255 43119 30552 43416 ne
rect 30552 43398 31964 43416
tri 31964 43398 32253 43687 sw
tri 32253 43398 32542 43687 ne
rect 32542 43486 34144 43687
tri 34144 43486 34434 43776 sw
tri 34434 43486 34724 43776 ne
rect 34724 43710 38495 43776
tri 38495 43710 38744 43959 sw
tri 38789 43710 39038 43959 ne
rect 39038 43820 42884 43959
tri 42884 43820 43172 44108 sw
tri 43172 43820 43460 44108 ne
rect 43460 44090 47230 44108
tri 47230 44090 47434 44294 sw
tri 47527 44090 47731 44294 ne
rect 47731 44090 51692 44294
rect 43460 43820 47434 44090
rect 39038 43819 43172 43820
tri 43172 43819 43173 43820 sw
tri 43460 43819 43461 43820 ne
rect 43461 43819 47434 43820
rect 39038 43710 43173 43819
rect 34724 43486 38744 43710
rect 32542 43398 34434 43486
rect 30552 43119 32253 43398
rect 26213 43118 30255 43119
tri 30255 43118 30256 43119 sw
tri 30552 43118 30553 43119 ne
rect 30553 43118 32253 43119
rect 26213 42917 30256 43118
rect 21852 42752 25931 42917
rect 20604 42751 21560 42752
tri 21560 42751 21561 42752 sw
tri 21852 42751 21853 42752 ne
rect 21853 42751 25931 42752
rect 20604 42459 21561 42751
tri 21561 42459 21853 42751 sw
tri 21853 42459 22145 42751 ne
rect 22145 42664 25931 42751
tri 25931 42664 26184 42917 sw
tri 26213 42664 26466 42917 ne
rect 26466 42821 30256 42917
tri 30256 42821 30553 43118 sw
tri 30553 42821 30850 43118 ne
rect 30850 43109 32253 43118
tri 32253 43109 32542 43398 sw
tri 32542 43109 32831 43398 ne
rect 32831 43311 34434 43398
tri 34434 43311 34609 43486 sw
tri 34724 43311 34899 43486 ne
rect 34899 43482 38744 43486
tri 38744 43482 38972 43710 sw
tri 39038 43482 39266 43710 ne
rect 39266 43531 43173 43710
tri 43173 43531 43461 43819 sw
tri 43461 43531 43749 43819 ne
rect 43749 43793 47434 43819
tri 47434 43793 47731 44090 sw
tri 47731 43793 48028 44090 ne
rect 48028 44080 51692 44090
tri 51692 44080 51985 44373 sw
tri 51985 44080 52278 44373 ne
rect 52278 44288 53758 44373
tri 53758 44288 54050 44580 sw
tri 54050 44288 54342 44580 ne
rect 54342 44579 56030 44580
tri 56030 44579 56031 44580 sw
tri 56317 44579 56318 44580 ne
rect 56318 44579 71000 44580
rect 54342 44292 56031 44579
tri 56031 44292 56318 44579 sw
tri 56318 44292 56605 44579 ne
rect 56605 44292 71000 44579
rect 54342 44288 56318 44292
rect 52278 44080 54050 44288
rect 48028 43937 51985 44080
tri 51985 43937 52128 44080 sw
tri 52278 43937 52421 44080 ne
rect 52421 43996 54050 44080
tri 54050 43996 54342 44288 sw
tri 54342 43996 54634 44288 ne
rect 54634 44005 56318 44288
tri 56318 44005 56605 44292 sw
tri 56605 44005 56892 44292 ne
rect 56892 44005 71000 44292
rect 54634 44004 56605 44005
tri 56605 44004 56606 44005 sw
tri 56892 44004 56893 44005 ne
rect 56893 44004 71000 44005
rect 54634 43996 56606 44004
rect 52421 43937 54342 43996
rect 48028 43793 52128 43937
rect 43749 43643 47731 43793
tri 47731 43643 47881 43793 sw
tri 48028 43643 48178 43793 ne
rect 48178 43644 52128 43793
tri 52128 43644 52421 43937 sw
tri 52421 43644 52714 43937 ne
rect 52714 43856 54342 43937
tri 54342 43856 54482 43996 sw
tri 54634 43856 54774 43996 ne
rect 54774 43856 56606 43996
rect 52714 43644 54482 43856
rect 48178 43643 52421 43644
tri 52421 43643 52422 43644 sw
tri 52714 43643 52715 43644 ne
rect 52715 43643 54482 43644
rect 43749 43531 47881 43643
rect 39266 43529 43461 43531
tri 43461 43529 43463 43531 sw
tri 43749 43529 43751 43531 ne
rect 43751 43529 47881 43531
rect 39266 43482 43463 43529
rect 34899 43415 38972 43482
tri 38972 43415 39039 43482 sw
tri 39266 43415 39333 43482 ne
rect 39333 43415 43463 43482
rect 34899 43311 39039 43415
rect 32831 43109 34609 43311
rect 30850 42821 32542 43109
rect 26466 42664 30553 42821
rect 22145 42459 26184 42664
rect 20604 42372 21853 42459
tri 21853 42372 21940 42459 sw
tri 22145 42372 22232 42459 ne
rect 22232 42382 26184 42459
tri 26184 42382 26466 42664 sw
tri 26466 42382 26748 42664 ne
rect 26748 42524 30553 42664
tri 30553 42524 30850 42821 sw
tri 30850 42524 31147 42821 ne
rect 31147 42820 32542 42821
tri 32542 42820 32831 43109 sw
tri 32831 42820 33120 43109 ne
rect 33120 43021 34609 43109
tri 34609 43021 34899 43311 sw
tri 34899 43021 35189 43311 ne
rect 35189 43121 39039 43311
tri 39039 43121 39333 43415 sw
tri 39333 43121 39627 43415 ne
rect 39627 43241 43463 43415
tri 43463 43241 43751 43529 sw
tri 43751 43241 44039 43529 ne
rect 44039 43346 47881 43529
tri 47881 43346 48178 43643 sw
tri 48178 43346 48475 43643 ne
rect 48475 43350 52422 43643
tri 52422 43350 52715 43643 sw
tri 52715 43350 53008 43643 ne
rect 53008 43564 54482 43643
tri 54482 43564 54774 43856 sw
tri 54774 43564 55066 43856 ne
rect 55066 43717 56606 43856
tri 56606 43717 56893 44004 sw
tri 56893 43717 57180 44004 ne
rect 57180 43717 71000 44004
rect 55066 43564 56893 43717
rect 53008 43350 54774 43564
rect 48475 43346 52715 43350
rect 44039 43345 48178 43346
tri 48178 43345 48179 43346 sw
tri 48475 43345 48476 43346 ne
rect 48476 43345 52715 43346
rect 44039 43241 48179 43345
rect 39627 43121 43751 43241
rect 35189 43119 39333 43121
tri 39333 43119 39335 43121 sw
tri 39627 43119 39629 43121 ne
rect 39629 43119 43751 43121
rect 35189 43021 39335 43119
rect 33120 42820 34899 43021
rect 31147 42531 32831 42820
tri 32831 42531 33120 42820 sw
tri 33120 42531 33409 42820 ne
rect 33409 42731 34899 42820
tri 34899 42731 35189 43021 sw
tri 35189 42731 35479 43021 ne
rect 35479 42825 39335 43021
tri 39335 42825 39629 43119 sw
tri 39629 42825 39923 43119 ne
rect 39923 42953 43751 43119
tri 43751 42953 44039 43241 sw
tri 44039 42953 44327 43241 ne
rect 44327 43048 48179 43241
tri 48179 43048 48476 43345 sw
tri 48476 43048 48773 43345 ne
rect 48773 43057 52715 43345
tri 52715 43057 53008 43350 sw
tri 53008 43057 53301 43350 ne
rect 53301 43272 54774 43350
tri 54774 43272 55066 43564 sw
tri 55066 43272 55358 43564 ne
rect 55358 43462 56893 43564
tri 56893 43462 57148 43717 sw
tri 57180 43462 57435 43717 ne
rect 57435 43462 71000 43717
rect 55358 43272 57148 43462
rect 53301 43057 55066 43272
rect 48773 43048 53008 43057
rect 44327 43047 48476 43048
tri 48476 43047 48477 43048 sw
tri 48773 43047 48774 43048 ne
rect 48774 43047 53008 43048
rect 44327 42953 48477 43047
rect 39923 42825 44039 42953
rect 35479 42824 39629 42825
tri 39629 42824 39630 42825 sw
tri 39923 42824 39924 42825 ne
rect 39924 42824 44039 42825
rect 35479 42731 39630 42824
rect 33409 42730 35189 42731
tri 35189 42730 35190 42731 sw
tri 35479 42730 35480 42731 ne
rect 35480 42730 39630 42731
rect 33409 42531 35190 42730
rect 31147 42524 33120 42531
rect 26748 42523 30850 42524
tri 30850 42523 30851 42524 sw
tri 31147 42523 31148 42524 ne
rect 31148 42523 33120 42524
rect 26748 42382 30851 42523
rect 22232 42372 26466 42382
rect 20604 42080 21940 42372
tri 21940 42080 22232 42372 sw
tri 22232 42080 22524 42372 ne
rect 22524 42264 26466 42372
tri 26466 42264 26584 42382 sw
tri 26748 42264 26866 42382 ne
rect 26866 42264 30851 42382
rect 22524 42080 26584 42264
rect 20604 41871 22232 42080
tri 22232 41871 22441 42080 sw
tri 22524 41871 22733 42080 ne
rect 22733 41982 26584 42080
tri 26584 41982 26866 42264 sw
tri 26866 41982 27148 42264 ne
rect 27148 42226 30851 42264
tri 30851 42226 31148 42523 sw
tri 31148 42226 31445 42523 ne
rect 31445 42440 33120 42523
tri 33120 42440 33211 42531 sw
tri 33409 42440 33500 42531 ne
rect 33500 42440 35190 42531
tri 35190 42440 35480 42730 sw
tri 35480 42440 35770 42730 ne
rect 35770 42530 39630 42730
tri 39630 42530 39924 42824 sw
tri 39924 42530 40218 42824 ne
rect 40218 42732 44039 42824
tri 44039 42732 44260 42953 sw
tri 44327 42732 44548 42953 ne
rect 44548 42750 48477 42953
tri 48477 42750 48774 43047 sw
tri 48774 42750 49071 43047 ne
rect 49071 42981 53008 43047
tri 53008 42981 53084 43057 sw
tri 53301 42981 53377 43057 ne
rect 53377 42981 55066 43057
rect 49071 42750 53084 42981
rect 44548 42749 48774 42750
tri 48774 42749 48775 42750 sw
tri 49071 42749 49072 42750 ne
rect 49072 42749 53084 42750
rect 44548 42732 48775 42749
rect 40218 42530 44260 42732
rect 35770 42440 39924 42530
rect 31445 42226 33211 42440
rect 27148 42225 31148 42226
tri 31148 42225 31149 42226 sw
tri 31445 42225 31446 42226 ne
rect 31446 42225 33211 42226
rect 27148 41982 31149 42225
rect 22733 41981 26866 41982
tri 26866 41981 26867 41982 sw
tri 27148 41981 27149 41982 ne
rect 27149 41981 31149 41982
rect 22733 41871 26867 41981
rect 20604 41579 22441 41871
tri 22441 41579 22733 41871 sw
tri 22733 41579 23025 41871 ne
rect 23025 41699 26867 41871
tri 26867 41699 27149 41981 sw
tri 27149 41699 27431 41981 ne
rect 27431 41928 31149 41981
tri 31149 41928 31446 42225 sw
tri 31446 41928 31743 42225 ne
rect 31743 42151 33211 42225
tri 33211 42151 33500 42440 sw
tri 33500 42151 33789 42440 ne
rect 33789 42439 35480 42440
tri 35480 42439 35481 42440 sw
tri 35770 42439 35771 42440 ne
rect 35771 42439 39924 42440
rect 33789 42151 35481 42439
rect 31743 41928 33500 42151
rect 27431 41699 31446 41928
rect 23025 41698 27149 41699
tri 27149 41698 27150 41699 sw
tri 27431 41698 27432 41699 ne
rect 27432 41698 31446 41699
rect 23025 41579 27150 41698
rect 20604 41415 22733 41579
tri 22733 41415 22897 41579 sw
tri 23025 41415 23189 41579 ne
rect 23189 41416 27150 41579
tri 27150 41416 27432 41698 sw
tri 27432 41416 27714 41698 ne
rect 27714 41631 31446 41698
tri 31446 41631 31743 41928 sw
tri 31743 41631 32040 41928 ne
rect 32040 41862 33500 41928
tri 33500 41862 33789 42151 sw
tri 33789 41862 34078 42151 ne
rect 34078 42149 35481 42151
tri 35481 42149 35771 42439 sw
tri 35771 42149 36061 42439 ne
rect 36061 42438 39924 42439
tri 39924 42438 40016 42530 sw
tri 40218 42438 40310 42530 ne
rect 40310 42444 44260 42530
tri 44260 42444 44548 42732 sw
tri 44548 42444 44836 42732 ne
rect 44836 42452 48775 42732
tri 48775 42452 49072 42749 sw
tri 49072 42452 49369 42749 ne
rect 49369 42688 53084 42749
tri 53084 42688 53377 42981 sw
tri 53377 42688 53670 42981 ne
rect 53670 42980 55066 42981
tri 55066 42980 55358 43272 sw
tri 55358 42980 55650 43272 ne
rect 55650 43175 57148 43272
tri 57148 43175 57435 43462 sw
tri 57435 43175 57722 43462 ne
rect 57722 43175 71000 43462
rect 55650 42980 57435 43175
rect 53670 42688 55358 42980
tri 55358 42688 55650 42980 sw
tri 55650 42688 55942 42980 ne
rect 55942 42888 57435 42980
tri 57435 42888 57722 43175 sw
tri 57722 42888 58009 43175 ne
rect 58009 42888 71000 43175
rect 55942 42800 57722 42888
tri 57722 42800 57810 42888 sw
tri 58009 42800 58097 42888 ne
rect 58097 42800 71000 42888
rect 55942 42688 57810 42800
rect 49369 42687 53377 42688
tri 53377 42687 53378 42688 sw
tri 53670 42687 53671 42688 ne
rect 53671 42687 55650 42688
rect 49369 42452 53378 42687
rect 44836 42451 49072 42452
tri 49072 42451 49073 42452 sw
tri 49369 42451 49370 42452 ne
rect 49370 42451 53378 42452
rect 44836 42444 49073 42451
rect 40310 42438 44548 42444
rect 36061 42149 40016 42438
rect 34078 41862 35771 42149
rect 32040 41707 33789 41862
tri 33789 41707 33944 41862 sw
tri 34078 41707 34233 41862 ne
rect 34233 41859 35771 41862
tri 35771 41859 36061 42149 sw
tri 36061 41859 36351 42149 ne
rect 36351 42144 40016 42149
tri 40016 42144 40310 42438 sw
tri 40310 42144 40604 42438 ne
rect 40604 42354 44548 42438
tri 44548 42354 44638 42444 sw
tri 44836 42354 44926 42444 ne
rect 44926 42354 49073 42444
rect 40604 42144 44638 42354
rect 36351 41939 40310 42144
tri 40310 41939 40515 42144 sw
tri 40604 41939 40809 42144 ne
rect 40809 42066 44638 42144
tri 44638 42066 44926 42354 sw
tri 44926 42066 45214 42354 ne
rect 45214 42154 49073 42354
tri 49073 42154 49370 42451 sw
tri 49370 42154 49667 42451 ne
rect 49667 42394 53378 42451
tri 53378 42394 53671 42687 sw
tri 53671 42394 53964 42687 ne
rect 53964 42600 55650 42687
tri 55650 42600 55738 42688 sw
tri 55942 42600 56030 42688 ne
rect 56030 42600 57810 42688
tri 57810 42600 58010 42800 sw
rect 53964 42394 55738 42600
rect 49667 42393 53671 42394
tri 53671 42393 53672 42394 sw
tri 53964 42393 53965 42394 ne
rect 53965 42393 55738 42394
rect 49667 42154 53672 42393
rect 45214 42152 49370 42154
tri 49370 42152 49372 42154 sw
tri 49667 42152 49669 42154 ne
rect 49669 42152 53672 42154
rect 45214 42066 49372 42152
rect 40809 42065 44926 42066
tri 44926 42065 44927 42066 sw
tri 45214 42065 45215 42066 ne
rect 45215 42065 49372 42066
rect 40809 41939 44927 42065
rect 36351 41859 40515 41939
rect 34233 41858 36061 41859
tri 36061 41858 36062 41859 sw
tri 36351 41858 36352 41859 ne
rect 36352 41858 40515 41859
rect 34233 41707 36062 41858
rect 32040 41631 33944 41707
rect 27714 41416 31743 41631
rect 23189 41415 27432 41416
rect 20604 41123 22897 41415
tri 22897 41123 23189 41415 sw
tri 23189 41123 23481 41415 ne
rect 23481 41338 27432 41415
tri 27432 41338 27510 41416 sw
tri 27714 41338 27792 41416 ne
rect 27792 41338 31743 41416
rect 23481 41123 27510 41338
rect 20604 41121 23189 41123
tri 23189 41121 23191 41123 sw
tri 23481 41121 23483 41123 ne
rect 23483 41121 27510 41123
rect 20604 40829 23191 41121
tri 23191 40829 23483 41121 sw
tri 23483 40829 23775 41121 ne
rect 23775 41056 27510 41121
tri 27510 41056 27792 41338 sw
tri 27792 41056 28074 41338 ne
rect 28074 41334 31743 41338
tri 31743 41334 32040 41631 sw
tri 32040 41334 32337 41631 ne
rect 32337 41418 33944 41631
tri 33944 41418 34233 41707 sw
tri 34233 41418 34522 41707 ne
rect 34522 41568 36062 41707
tri 36062 41568 36352 41858 sw
tri 36352 41568 36642 41858 ne
rect 36642 41645 40515 41858
tri 40515 41645 40809 41939 sw
tri 40809 41645 41103 41939 ne
rect 41103 41777 44927 41939
tri 44927 41777 45215 42065 sw
tri 45215 41777 45503 42065 ne
rect 45503 41856 49372 42065
tri 49372 41856 49668 42152 sw
tri 49669 41856 49965 42152 ne
rect 49965 42100 53672 42152
tri 53672 42100 53965 42393 sw
tri 53965 42100 54258 42393 ne
rect 54258 42308 55738 42393
tri 55738 42308 56030 42600 sw
tri 56030 42308 56322 42600 ne
rect 56322 42308 71000 42600
rect 54258 42100 56030 42308
rect 49965 41856 53965 42100
rect 45503 41777 49668 41856
rect 41103 41775 45215 41777
tri 45215 41775 45217 41777 sw
tri 45503 41775 45505 41777 ne
rect 45505 41775 49668 41777
rect 41103 41645 45217 41775
rect 36642 41568 40809 41645
rect 34522 41418 36352 41568
rect 32337 41334 34233 41418
rect 28074 41138 32040 41334
tri 32040 41138 32236 41334 sw
tri 32337 41138 32533 41334 ne
rect 32533 41138 34233 41334
rect 28074 41056 32236 41138
rect 23775 40848 27792 41056
tri 27792 40848 28000 41056 sw
tri 28074 40848 28282 41056 ne
rect 28282 40848 32236 41056
rect 23775 40829 28000 40848
rect 20604 40828 23483 40829
tri 23483 40828 23484 40829 sw
tri 23775 40828 23776 40829 ne
rect 23776 40828 28000 40829
rect 20604 40536 23484 40828
tri 23484 40536 23776 40828 sw
tri 23776 40536 24068 40828 ne
rect 24068 40566 28000 40828
tri 28000 40566 28282 40848 sw
tri 28282 40566 28564 40848 ne
rect 28564 40841 32236 40848
tri 32236 40841 32533 41138 sw
tri 32533 40841 32830 41138 ne
rect 32830 41129 34233 41138
tri 34233 41129 34522 41418 sw
tri 34522 41129 34811 41418 ne
rect 34811 41331 36352 41418
tri 36352 41331 36589 41568 sw
tri 36642 41331 36879 41568 ne
rect 36879 41486 40809 41568
tri 40809 41486 40968 41645 sw
tri 41103 41486 41262 41645 ne
rect 41262 41488 45217 41645
tri 45217 41488 45504 41775 sw
tri 45505 41488 45792 41775 ne
rect 45792 41636 49668 41775
tri 49668 41636 49888 41856 sw
tri 49965 41636 50185 41856 ne
rect 50185 41807 53965 41856
tri 53965 41807 54258 42100 sw
tri 54258 41807 54551 42100 ne
rect 54551 42016 56030 42100
tri 56030 42016 56322 42308 sw
tri 56322 42016 56614 42308 ne
rect 56614 42016 71000 42308
rect 54551 41876 56322 42016
tri 56322 41876 56462 42016 sw
tri 56614 41876 56754 42016 ne
rect 56754 41876 71000 42016
rect 54551 41807 56462 41876
rect 50185 41636 54258 41807
rect 45792 41488 49888 41636
rect 41262 41486 45504 41488
rect 36879 41331 40968 41486
rect 34811 41129 36589 41331
rect 32830 40841 34522 41129
rect 28564 40566 32533 40841
rect 24068 40536 28282 40566
rect 20604 40535 23776 40536
tri 23776 40535 23777 40536 sw
tri 24068 40535 24069 40536 ne
rect 24069 40535 28282 40536
rect 20604 40243 23777 40535
tri 23777 40243 24069 40535 sw
tri 24069 40243 24361 40535 ne
rect 24361 40372 28282 40535
tri 28282 40372 28476 40566 sw
tri 28564 40372 28758 40566 ne
rect 28758 40544 32533 40566
tri 32533 40544 32830 40841 sw
tri 32830 40544 33127 40841 ne
rect 33127 40840 34522 40841
tri 34522 40840 34811 41129 sw
tri 34811 40840 35100 41129 ne
rect 35100 41041 36589 41129
tri 36589 41041 36879 41331 sw
tri 36879 41041 37169 41331 ne
rect 37169 41192 40968 41331
tri 40968 41192 41262 41486 sw
tri 41262 41192 41556 41486 ne
rect 41556 41400 45504 41486
tri 45504 41400 45592 41488 sw
tri 45792 41400 45880 41488 ne
rect 45880 41400 49888 41488
rect 41556 41192 45592 41400
rect 37169 41191 41262 41192
tri 41262 41191 41263 41192 sw
tri 41556 41191 41557 41192 ne
rect 41557 41191 45592 41192
rect 37169 41041 41263 41191
rect 35100 40840 36879 41041
rect 33127 40551 34811 40840
tri 34811 40551 35100 40840 sw
tri 35100 40551 35389 40840 ne
rect 35389 40751 36879 40840
tri 36879 40751 37169 41041 sw
tri 37169 40751 37459 41041 ne
rect 37459 40897 41263 41041
tri 41263 40897 41557 41191 sw
tri 41557 40897 41851 41191 ne
rect 41851 41112 45592 41191
tri 45592 41112 45880 41400 sw
tri 45880 41112 46168 41400 ne
rect 46168 41391 49888 41400
tri 49888 41391 50133 41636 sw
tri 50185 41391 50430 41636 ne
rect 50430 41588 54258 41636
tri 54258 41588 54477 41807 sw
tri 54551 41588 54770 41807 ne
rect 54770 41588 56462 41807
rect 50430 41391 54477 41588
rect 46168 41338 50133 41391
tri 50133 41338 50186 41391 sw
tri 50430 41338 50483 41391 ne
rect 50483 41338 54477 41391
rect 46168 41112 50186 41338
rect 41851 40908 45880 41112
tri 45880 40908 46084 41112 sw
tri 46168 40908 46372 41112 ne
rect 46372 41041 50186 41112
tri 50186 41041 50483 41338 sw
tri 50483 41041 50780 41338 ne
rect 50780 41295 54477 41338
tri 54477 41295 54770 41588 sw
tri 54770 41295 55063 41588 ne
rect 55063 41584 56462 41588
tri 56462 41584 56754 41876 sw
tri 56754 41584 57046 41876 ne
rect 57046 41584 71000 41876
rect 55063 41295 56754 41584
rect 50780 41294 54770 41295
tri 54770 41294 54771 41295 sw
tri 55063 41294 55064 41295 ne
rect 55064 41294 56754 41295
rect 50780 41041 54771 41294
rect 46372 41040 50483 41041
tri 50483 41040 50484 41041 sw
tri 50780 41040 50781 41041 ne
rect 50781 41040 54771 41041
rect 46372 40908 50484 41040
rect 41851 40897 46084 40908
rect 37459 40896 41557 40897
tri 41557 40896 41558 40897 sw
tri 41851 40896 41852 40897 ne
rect 41852 40896 46084 40897
rect 37459 40751 41558 40896
rect 35389 40750 37169 40751
tri 37169 40750 37170 40751 sw
tri 37459 40750 37460 40751 ne
rect 37460 40750 41558 40751
rect 35389 40551 37170 40750
rect 33127 40544 35100 40551
rect 28758 40372 32830 40544
tri 32830 40372 33002 40544 sw
tri 33127 40372 33299 40544 ne
rect 33299 40460 35100 40544
tri 35100 40460 35191 40551 sw
tri 35389 40460 35480 40551 ne
rect 35480 40460 37170 40551
tri 37170 40460 37460 40750 sw
tri 37460 40460 37750 40750 ne
rect 37750 40602 41558 40750
tri 41558 40602 41852 40896 sw
tri 41852 40602 42146 40896 ne
rect 42146 40620 46084 40896
tri 46084 40620 46372 40908 sw
tri 46372 40620 46660 40908 ne
rect 46660 40743 50484 40908
tri 50484 40743 50781 41040 sw
tri 50781 40743 51078 41040 ne
rect 51078 41001 54771 41040
tri 54771 41001 55064 41294 sw
tri 55064 41001 55357 41294 ne
rect 55357 41292 56754 41294
tri 56754 41292 57046 41584 sw
tri 57046 41292 57338 41584 ne
rect 57338 41292 71000 41584
rect 55357 41001 57046 41292
rect 51078 40743 55064 41001
rect 46660 40742 50781 40743
tri 50781 40742 50782 40743 sw
tri 51078 40742 51079 40743 ne
rect 51079 40742 55064 40743
rect 46660 40620 50782 40742
rect 42146 40602 46372 40620
rect 37750 40601 41852 40602
tri 41852 40601 41853 40602 sw
tri 42146 40601 42147 40602 ne
rect 42147 40601 46372 40602
rect 37750 40460 41853 40601
rect 33299 40372 35191 40460
rect 24361 40243 28476 40372
rect 20604 40242 24069 40243
tri 24069 40242 24070 40243 sw
tri 24361 40242 24362 40243 ne
rect 24362 40242 28476 40243
rect 20604 39950 24070 40242
tri 24070 39950 24362 40242 sw
tri 24362 39950 24654 40242 ne
rect 24654 40090 28476 40242
tri 28476 40090 28758 40372 sw
tri 28758 40090 29040 40372 ne
rect 29040 40090 33002 40372
rect 24654 40089 28758 40090
tri 28758 40089 28759 40090 sw
tri 29040 40089 29041 40090 ne
rect 29041 40089 33002 40090
rect 24654 39950 28759 40089
rect 20604 39949 24362 39950
tri 24362 39949 24363 39950 sw
tri 24654 39949 24655 39950 ne
rect 24655 39949 28759 39950
rect 20604 39657 24363 39949
tri 24363 39657 24655 39949 sw
tri 24655 39657 24947 39949 ne
rect 24947 39807 28759 39949
tri 28759 39807 29041 40089 sw
tri 29041 39807 29323 40089 ne
rect 29323 40075 33002 40089
tri 33002 40075 33299 40372 sw
tri 33299 40075 33596 40372 ne
rect 33596 40171 35191 40372
tri 35191 40171 35480 40460 sw
tri 35480 40171 35769 40460 ne
rect 35769 40459 37460 40460
tri 37460 40459 37461 40460 sw
tri 37750 40459 37751 40460 ne
rect 37751 40459 41853 40460
rect 35769 40171 37461 40459
rect 33596 40075 35480 40171
rect 29323 40074 33299 40075
tri 33299 40074 33300 40075 sw
tri 33596 40074 33597 40075 ne
rect 33597 40074 35480 40075
rect 29323 39807 33300 40074
rect 24947 39805 29041 39807
tri 29041 39805 29043 39807 sw
tri 29323 39805 29325 39807 ne
rect 29325 39805 33300 39807
rect 24947 39657 29043 39805
rect 20604 39464 24655 39657
tri 24655 39464 24848 39657 sw
tri 24947 39464 25140 39657 ne
rect 25140 39523 29043 39657
tri 29043 39523 29325 39805 sw
tri 29325 39523 29607 39805 ne
rect 29607 39777 33300 39805
tri 33300 39777 33597 40074 sw
tri 33597 39777 33894 40074 ne
rect 33894 39882 35480 40074
tri 35480 39882 35769 40171 sw
tri 35769 39882 36058 40171 ne
rect 36058 40169 37461 40171
tri 37461 40169 37751 40459 sw
tri 37751 40169 38041 40459 ne
rect 38041 40307 41853 40459
tri 41853 40307 42147 40601 sw
tri 42147 40307 42441 40601 ne
rect 42441 40443 46372 40601
tri 46372 40443 46549 40620 sw
tri 46660 40443 46837 40620 ne
rect 46837 40445 50782 40620
tri 50782 40445 51079 40742 sw
tri 51079 40445 51376 40742 ne
rect 51376 40708 55064 40742
tri 55064 40708 55357 41001 sw
tri 55357 40708 55650 41001 ne
rect 55650 41000 57046 41001
tri 57046 41000 57338 41292 sw
tri 57338 41200 57430 41292 ne
rect 57430 41200 71000 41292
rect 55650 40708 71000 41000
rect 51376 40644 55357 40708
tri 55357 40644 55421 40708 sw
tri 55650 40644 55714 40708 ne
rect 55714 40644 71000 40708
rect 51376 40445 55421 40644
rect 46837 40443 51079 40445
rect 42441 40307 46549 40443
rect 38041 40305 42147 40307
tri 42147 40305 42149 40307 sw
tri 42441 40305 42443 40307 ne
rect 42443 40305 46549 40307
rect 38041 40169 42149 40305
rect 36058 39882 37751 40169
rect 33894 39777 35769 39882
rect 29607 39523 33597 39777
rect 25140 39522 29325 39523
tri 29325 39522 29326 39523 sw
tri 29607 39522 29608 39523 ne
rect 29608 39522 33597 39523
rect 25140 39464 29326 39522
tri 20604 35220 24848 39464 ne
tri 24848 39172 25140 39464 sw
tri 25140 39172 25432 39464 ne
rect 25432 39240 29326 39464
tri 29326 39240 29608 39522 sw
tri 29608 39240 29890 39522 ne
rect 29890 39480 33597 39522
tri 33597 39480 33894 39777 sw
tri 33894 39480 34191 39777 ne
rect 34191 39653 35769 39777
tri 35769 39653 35998 39882 sw
tri 36058 39653 36287 39882 ne
rect 36287 39879 37751 39882
tri 37751 39879 38041 40169 sw
tri 38041 39879 38331 40169 ne
rect 38331 40011 42149 40169
tri 42149 40011 42443 40305 sw
tri 42443 40011 42737 40305 ne
rect 42737 40155 46549 40305
tri 46549 40155 46837 40443 sw
tri 46837 40155 47125 40443 ne
rect 47125 40347 51079 40443
tri 51079 40347 51177 40445 sw
tri 51376 40347 51474 40445 ne
rect 51474 40351 55421 40445
tri 55421 40351 55714 40644 sw
tri 55714 40351 56007 40644 ne
rect 56007 40351 71000 40644
rect 51474 40347 55714 40351
rect 47125 40155 51177 40347
rect 42737 40154 46837 40155
tri 46837 40154 46838 40155 sw
tri 47125 40154 47126 40155 ne
rect 47126 40154 51177 40155
rect 42737 40011 46838 40154
rect 38331 39879 42443 40011
rect 36287 39878 38041 39879
tri 38041 39878 38042 39879 sw
tri 38331 39878 38332 39879 ne
rect 38332 39878 42443 39879
rect 36287 39653 38042 39878
rect 34191 39480 35998 39653
rect 29890 39479 33894 39480
tri 33894 39479 33895 39480 sw
tri 34191 39479 34192 39480 ne
rect 34192 39479 35998 39480
rect 29890 39240 33895 39479
rect 25432 39239 29608 39240
tri 29608 39239 29609 39240 sw
tri 29890 39239 29891 39240 ne
rect 29891 39239 33895 39240
rect 25432 39172 29609 39239
rect 24848 39094 25140 39172
tri 25140 39094 25218 39172 sw
tri 25432 39094 25510 39172 ne
rect 25510 39094 29609 39172
rect 24848 38802 25218 39094
tri 25218 38802 25510 39094 sw
tri 25510 38802 25802 39094 ne
rect 25802 38957 29609 39094
tri 29609 38957 29891 39239 sw
tri 29891 38957 30173 39239 ne
rect 30173 39182 33895 39239
tri 33895 39182 34192 39479 sw
tri 34192 39182 34489 39479 ne
rect 34489 39438 35998 39479
tri 35998 39438 36213 39653 sw
tri 36287 39438 36502 39653 ne
rect 36502 39588 38042 39653
tri 38042 39588 38332 39878 sw
tri 38332 39588 38622 39878 ne
rect 38622 39717 42443 39878
tri 42443 39717 42737 40011 sw
tri 42737 39717 43031 40011 ne
rect 43031 39866 46838 40011
tri 46838 39866 47126 40154 sw
tri 47126 39866 47414 40154 ne
rect 47414 40050 51177 40154
tri 51177 40050 51474 40347 sw
tri 51474 40050 51771 40347 ne
rect 51771 40120 55714 40347
tri 55714 40120 55945 40351 sw
tri 56007 40120 56238 40351 ne
rect 56238 40120 71000 40351
rect 51771 40050 55945 40120
rect 47414 39866 51474 40050
rect 43031 39865 47126 39866
tri 47126 39865 47127 39866 sw
tri 47414 39865 47415 39866 ne
rect 47415 39865 51474 39866
rect 43031 39717 47127 39865
rect 38622 39588 42737 39717
rect 36502 39438 38332 39588
rect 34489 39182 36213 39438
rect 30173 39158 34192 39182
tri 34192 39158 34216 39182 sw
tri 34489 39158 34513 39182 ne
rect 34513 39158 36213 39182
rect 30173 38957 34216 39158
rect 25802 38956 29891 38957
tri 29891 38956 29892 38957 sw
tri 30173 38956 30174 38957 ne
rect 30174 38956 34216 38957
rect 25802 38802 29892 38956
rect 24848 38801 25510 38802
tri 25510 38801 25511 38802 sw
tri 25802 38801 25803 38802 ne
rect 25803 38801 29892 38802
rect 24848 38509 25511 38801
tri 25511 38509 25803 38801 sw
tri 25803 38509 26095 38801 ne
rect 26095 38674 29892 38801
tri 29892 38674 30174 38956 sw
tri 30174 38674 30456 38956 ne
rect 30456 38861 34216 38956
tri 34216 38861 34513 39158 sw
tri 34513 38861 34810 39158 ne
rect 34810 39149 36213 39158
tri 36213 39149 36502 39438 sw
tri 36502 39149 36791 39438 ne
rect 36791 39352 38332 39438
tri 38332 39352 38568 39588 sw
tri 38622 39352 38858 39588 ne
rect 38858 39467 42737 39588
tri 42737 39467 42987 39717 sw
tri 43031 39467 43281 39717 ne
rect 43281 39577 47127 39717
tri 47127 39577 47415 39865 sw
tri 47415 39577 47703 39865 ne
rect 47703 39847 51474 39865
tri 51474 39847 51677 40050 sw
tri 51771 39847 51974 40050 ne
rect 51974 39988 55945 40050
tri 55945 39988 56077 40120 sw
tri 56238 39988 56370 40120 ne
rect 56370 39988 71000 40120
rect 51974 39847 56077 39988
rect 47703 39577 51677 39847
rect 43281 39576 47415 39577
tri 47415 39576 47416 39577 sw
tri 47703 39576 47704 39577 ne
rect 47704 39576 51677 39577
rect 43281 39467 47416 39576
rect 38858 39352 42987 39467
rect 36791 39242 38568 39352
tri 38568 39242 38678 39352 sw
tri 38858 39242 38968 39352 ne
rect 38968 39242 42987 39352
rect 36791 39149 38678 39242
rect 34810 38861 36502 39149
rect 30456 38674 34513 38861
rect 26095 38509 30174 38674
rect 24848 38508 25803 38509
tri 25803 38508 25804 38509 sw
tri 26095 38508 26096 38509 ne
rect 26096 38508 30174 38509
rect 24848 38216 25804 38508
tri 25804 38216 26096 38508 sw
tri 26096 38216 26388 38508 ne
rect 26388 38420 30174 38508
tri 30174 38420 30428 38674 sw
tri 30456 38420 30710 38674 ne
rect 30710 38564 34513 38674
tri 34513 38564 34810 38861 sw
tri 34810 38564 35107 38861 ne
rect 35107 38860 36502 38861
tri 36502 38860 36791 39149 sw
tri 36791 38860 37080 39149 ne
rect 37080 39061 38678 39149
tri 38678 39061 38859 39242 sw
tri 38968 39061 39149 39242 ne
rect 39149 39238 42987 39242
tri 42987 39238 43216 39467 sw
tri 43281 39238 43510 39467 ne
rect 43510 39288 47416 39467
tri 47416 39288 47704 39576 sw
tri 47704 39288 47992 39576 ne
rect 47992 39550 51677 39576
tri 51677 39550 51974 39847 sw
tri 51974 39550 52271 39847 ne
rect 52271 39695 56077 39847
tri 56077 39695 56370 39988 sw
tri 56370 39695 56663 39988 ne
rect 56663 39695 71000 39988
rect 52271 39694 56370 39695
tri 56370 39694 56371 39695 sw
tri 56663 39694 56664 39695 ne
rect 56664 39694 71000 39695
rect 52271 39550 56371 39694
rect 47992 39401 51974 39550
tri 51974 39401 52123 39550 sw
tri 52271 39401 52420 39550 ne
rect 52420 39401 56371 39550
tri 56371 39401 56664 39694 sw
tri 56664 39600 56758 39694 ne
rect 56758 39600 71000 39694
rect 47992 39288 52123 39401
rect 43510 39287 47704 39288
tri 47704 39287 47705 39288 sw
tri 47992 39287 47993 39288 ne
rect 47993 39287 52123 39288
rect 43510 39238 47705 39287
rect 39149 39172 43216 39238
tri 43216 39172 43282 39238 sw
tri 43510 39172 43576 39238 ne
rect 43576 39172 47705 39238
rect 39149 39061 43282 39172
rect 37080 38860 38859 39061
rect 35107 38571 36791 38860
tri 36791 38571 37080 38860 sw
tri 37080 38571 37369 38860 ne
rect 37369 38771 38859 38860
tri 38859 38771 39149 39061 sw
tri 39149 38771 39439 39061 ne
rect 39439 38878 43282 39061
tri 43282 38878 43576 39172 sw
tri 43576 38878 43870 39172 ne
rect 43870 38999 47705 39172
tri 47705 38999 47993 39287 sw
tri 47993 38999 48281 39287 ne
rect 48281 39104 52123 39287
tri 52123 39104 52420 39401 sw
tri 52420 39104 52717 39401 ne
rect 52717 39400 56664 39401
tri 56664 39400 56665 39401 sw
rect 52717 39104 71000 39400
rect 48281 39102 52420 39104
tri 52420 39102 52422 39104 sw
tri 52717 39102 52719 39104 ne
rect 52719 39102 71000 39104
rect 48281 38999 52422 39102
rect 43870 38997 47993 38999
tri 47993 38997 47995 38999 sw
tri 48281 38997 48283 38999 ne
rect 48283 38997 52422 38999
rect 43870 38878 47995 38997
rect 39439 38877 43576 38878
tri 43576 38877 43577 38878 sw
tri 43870 38877 43871 38878 ne
rect 43871 38877 47995 38878
rect 39439 38771 43577 38877
rect 37369 38770 39149 38771
tri 39149 38770 39150 38771 sw
tri 39439 38770 39440 38771 ne
rect 39440 38770 43577 38771
rect 37369 38571 39150 38770
rect 35107 38564 37080 38571
rect 30710 38563 34810 38564
tri 34810 38563 34811 38564 sw
tri 35107 38563 35108 38564 ne
rect 35108 38563 37080 38564
rect 30710 38420 34811 38563
rect 26388 38216 30428 38420
rect 24848 38128 26096 38216
tri 26096 38128 26184 38216 sw
tri 26388 38128 26476 38216 ne
rect 26476 38138 30428 38216
tri 30428 38138 30710 38420 sw
tri 30710 38138 30992 38420 ne
rect 30992 38266 34811 38420
tri 34811 38266 35108 38563 sw
tri 35108 38266 35405 38563 ne
rect 35405 38406 37080 38563
tri 37080 38406 37245 38571 sw
tri 37369 38406 37534 38571 ne
rect 37534 38480 39150 38571
tri 39150 38480 39440 38770 sw
tri 39440 38480 39730 38770 ne
rect 39730 38583 43577 38770
tri 43577 38583 43871 38877 sw
tri 43871 38583 44165 38877 ne
rect 44165 38710 47995 38877
tri 47995 38710 48282 38997 sw
tri 48283 38710 48570 38997 ne
rect 48570 38805 52422 38997
tri 52422 38805 52719 39102 sw
tri 52719 38805 53016 39102 ne
rect 53016 38805 71000 39102
rect 48570 38804 52719 38805
tri 52719 38804 52720 38805 sw
tri 53016 38804 53017 38805 ne
rect 53017 38804 71000 38805
rect 48570 38710 52720 38804
rect 44165 38583 48282 38710
rect 39730 38581 43871 38583
tri 43871 38581 43873 38583 sw
tri 44165 38581 44167 38583 ne
rect 44167 38581 48282 38583
rect 39730 38480 43873 38581
rect 37534 38406 39440 38480
rect 35405 38266 37245 38406
rect 30992 38265 35108 38266
tri 35108 38265 35109 38266 sw
tri 35405 38265 35406 38266 ne
rect 35406 38265 37245 38266
rect 30992 38138 35109 38265
rect 26476 38128 30710 38138
rect 24848 37836 26184 38128
tri 26184 37836 26476 38128 sw
tri 26476 37836 26768 38128 ne
rect 26768 38021 30710 38128
tri 30710 38021 30827 38138 sw
tri 30992 38021 31109 38138 ne
rect 31109 38021 35109 38138
rect 26768 37836 30827 38021
rect 24848 37628 26476 37836
tri 26476 37628 26684 37836 sw
tri 26768 37628 26976 37836 ne
rect 26976 37739 30827 37836
tri 30827 37739 31109 38021 sw
tri 31109 37739 31391 38021 ne
rect 31391 37968 35109 38021
tri 35109 37968 35406 38265 sw
tri 35406 37968 35703 38265 ne
rect 35703 38191 37245 38265
tri 37245 38191 37460 38406 sw
tri 37534 38191 37749 38406 ne
rect 37749 38285 39440 38406
tri 39440 38285 39635 38480 sw
tri 39730 38285 39925 38480 ne
rect 39925 38288 43873 38480
tri 43873 38288 44166 38581 sw
tri 44167 38288 44460 38581 ne
rect 44460 38488 48282 38581
tri 48282 38488 48504 38710 sw
tri 48570 38488 48792 38710 ne
rect 48792 38507 52720 38710
tri 52720 38507 53017 38804 sw
tri 53017 38507 53314 38804 ne
rect 53314 38507 71000 38804
rect 48792 38506 53017 38507
tri 53017 38506 53018 38507 sw
tri 53314 38506 53315 38507 ne
rect 53315 38506 71000 38507
rect 48792 38488 53018 38506
rect 44460 38288 48504 38488
rect 39925 38285 44166 38288
rect 37749 38191 39635 38285
rect 35703 37968 37460 38191
rect 31391 37739 35406 37968
rect 26976 37738 31109 37739
tri 31109 37738 31110 37739 sw
tri 31391 37738 31392 37739 ne
rect 31392 37738 35406 37739
rect 26976 37628 31110 37738
rect 24848 37337 26684 37628
tri 26684 37337 26975 37628 sw
tri 26976 37337 27267 37628 ne
rect 27267 37456 31110 37628
tri 31110 37456 31392 37738 sw
tri 31392 37456 31674 37738 ne
rect 31674 37671 35406 37738
tri 35406 37671 35703 37968 sw
tri 35703 37671 36000 37968 ne
rect 36000 37902 37460 37968
tri 37460 37902 37749 38191 sw
tri 37749 37902 38038 38191 ne
rect 38038 37995 39635 38191
tri 39635 37995 39925 38285 sw
tri 39925 37995 40215 38285 ne
rect 40215 38194 44166 38285
tri 44166 38194 44260 38288 sw
tri 44460 38194 44554 38288 ne
rect 44554 38200 48504 38288
tri 48504 38200 48792 38488 sw
tri 48792 38200 49080 38488 ne
rect 49080 38209 53018 38488
tri 53018 38209 53315 38506 sw
tri 53315 38209 53612 38506 ne
rect 53612 38209 71000 38506
rect 49080 38208 53315 38209
tri 53315 38208 53316 38209 sw
tri 53612 38208 53613 38209 ne
rect 53613 38208 71000 38209
rect 49080 38200 53316 38208
rect 44554 38194 48792 38200
rect 40215 37995 44260 38194
rect 38038 37994 39925 37995
tri 39925 37994 39926 37995 sw
tri 40215 37994 40216 37995 ne
rect 40216 37994 44260 37995
rect 38038 37902 39926 37994
rect 36000 37747 37749 37902
tri 37749 37747 37904 37902 sw
tri 38038 37747 38193 37902 ne
rect 38193 37747 39926 37902
rect 36000 37671 37904 37747
rect 31674 37456 35703 37671
rect 27267 37455 31392 37456
tri 31392 37455 31393 37456 sw
tri 31674 37455 31675 37456 ne
rect 31675 37455 35703 37456
rect 27267 37337 31393 37455
rect 24848 37172 26975 37337
tri 26975 37172 27140 37337 sw
tri 27267 37172 27432 37337 ne
rect 27432 37173 31393 37337
tri 31393 37173 31675 37455 sw
tri 31675 37173 31957 37455 ne
rect 31957 37374 35703 37455
tri 35703 37374 36000 37671 sw
tri 36000 37374 36297 37671 ne
rect 36297 37458 37904 37671
tri 37904 37458 38193 37747 sw
tri 38193 37458 38482 37747 ne
rect 38482 37704 39926 37747
tri 39926 37704 40216 37994 sw
tri 40216 37704 40506 37994 ne
rect 40506 37900 44260 37994
tri 44260 37900 44554 38194 sw
tri 44554 37900 44848 38194 ne
rect 44848 38111 48792 38194
tri 48792 38111 48881 38200 sw
tri 49080 38111 49169 38200 ne
rect 49169 38111 53316 38200
rect 44848 37900 48881 38111
rect 40506 37704 44554 37900
rect 38482 37458 40216 37704
rect 36297 37374 38193 37458
rect 31957 37173 36000 37374
rect 27432 37172 31675 37173
rect 24848 36880 27140 37172
tri 27140 36880 27432 37172 sw
tri 27432 36880 27724 37172 ne
rect 27724 37094 31675 37172
tri 31675 37094 31754 37173 sw
tri 31957 37094 32036 37173 ne
rect 32036 37094 36000 37173
rect 27724 36880 31754 37094
rect 24848 36879 27432 36880
tri 27432 36879 27433 36880 sw
tri 27724 36879 27725 36880 ne
rect 27725 36879 31754 36880
rect 24848 36587 27433 36879
tri 27433 36587 27725 36879 sw
tri 27725 36587 28017 36879 ne
rect 28017 36812 31754 36879
tri 31754 36812 32036 37094 sw
tri 32036 36812 32318 37094 ne
rect 32318 37077 36000 37094
tri 36000 37077 36297 37374 sw
tri 36297 37077 36594 37374 ne
rect 36594 37169 38193 37374
tri 38193 37169 38482 37458 sw
tri 38482 37169 38771 37458 ne
rect 38771 37414 40216 37458
tri 40216 37414 40506 37704 sw
tri 40506 37414 40796 37704 ne
rect 40796 37696 44554 37704
tri 44554 37696 44758 37900 sw
tri 44848 37696 45052 37900 ne
rect 45052 37823 48881 37900
tri 48881 37823 49169 38111 sw
tri 49169 37823 49457 38111 ne
rect 49457 37911 53316 38111
tri 53316 37911 53613 38208 sw
tri 53613 37911 53910 38208 ne
rect 53910 37911 71000 38208
rect 49457 37910 53613 37911
tri 53613 37910 53614 37911 sw
tri 53910 37910 53911 37911 ne
rect 53911 37910 71000 37911
rect 49457 37823 53614 37910
rect 45052 37822 49169 37823
tri 49169 37822 49170 37823 sw
tri 49457 37822 49458 37823 ne
rect 49458 37822 53614 37823
rect 45052 37696 49170 37822
rect 40796 37414 44758 37696
rect 38771 37371 40506 37414
tri 40506 37371 40549 37414 sw
tri 40796 37371 40839 37414 ne
rect 40839 37402 44758 37414
tri 44758 37402 45052 37696 sw
tri 45052 37402 45346 37696 ne
rect 45346 37534 49170 37696
tri 49170 37534 49458 37822 sw
tri 49458 37534 49746 37822 ne
rect 49746 37613 53614 37822
tri 53614 37613 53911 37910 sw
tri 53911 37613 54208 37910 ne
rect 54208 37613 71000 37910
rect 49746 37534 53911 37613
rect 45346 37533 49458 37534
tri 49458 37533 49459 37534 sw
tri 49746 37533 49747 37534 ne
rect 49747 37533 53911 37534
rect 45346 37402 49459 37533
rect 40839 37371 45052 37402
rect 38771 37169 40549 37371
rect 36594 37077 38482 37169
rect 32318 36881 36297 37077
tri 36297 36881 36493 37077 sw
tri 36594 36881 36790 37077 ne
rect 36790 36881 38482 37077
rect 32318 36812 36493 36881
rect 28017 36605 32036 36812
tri 32036 36605 32243 36812 sw
tri 32318 36605 32525 36812 ne
rect 32525 36605 36493 36812
rect 28017 36587 32243 36605
rect 24848 36585 27725 36587
tri 27725 36585 27727 36587 sw
tri 28017 36585 28019 36587 ne
rect 28019 36585 32243 36587
rect 24848 36293 27727 36585
tri 27727 36293 28019 36585 sw
tri 28019 36293 28311 36585 ne
rect 28311 36323 32243 36585
tri 32243 36323 32525 36605 sw
tri 32525 36323 32807 36605 ne
rect 32807 36584 36493 36605
tri 36493 36584 36790 36881 sw
tri 36790 36584 37087 36881 ne
rect 37087 36880 38482 36881
tri 38482 36880 38771 37169 sw
tri 38771 36880 39060 37169 ne
rect 39060 37081 40549 37169
tri 40549 37081 40839 37371 sw
tri 40839 37081 41129 37371 ne
rect 41129 37243 45052 37371
tri 45052 37243 45211 37402 sw
tri 45346 37243 45505 37402 ne
rect 45505 37245 49459 37402
tri 49459 37245 49747 37533 sw
tri 49747 37245 50035 37533 ne
rect 50035 37393 53911 37533
tri 53911 37393 54131 37613 sw
tri 54208 37393 54428 37613 ne
rect 54428 37393 71000 37613
rect 50035 37245 54131 37393
rect 45505 37243 49747 37245
rect 41129 37081 45211 37243
rect 39060 36880 40839 37081
rect 37087 36591 38771 36880
tri 38771 36591 39060 36880 sw
tri 39060 36591 39349 36880 ne
rect 39349 36791 40839 36880
tri 40839 36791 41129 37081 sw
tri 41129 36791 41419 37081 ne
rect 41419 36949 45211 37081
tri 45211 36949 45505 37243 sw
tri 45505 36949 45799 37243 ne
rect 45799 37156 49747 37243
tri 49747 37156 49836 37245 sw
tri 50035 37156 50124 37245 ne
rect 50124 37156 54131 37245
rect 45799 36949 49836 37156
rect 41419 36948 45505 36949
tri 45505 36948 45506 36949 sw
tri 45799 36948 45800 36949 ne
rect 45800 36948 49836 36949
rect 41419 36791 45506 36948
rect 39349 36790 41129 36791
tri 41129 36790 41130 36791 sw
tri 41419 36790 41420 36791 ne
rect 41420 36790 45506 36791
rect 39349 36591 41130 36790
rect 37087 36584 39060 36591
rect 32807 36583 36790 36584
tri 36790 36583 36791 36584 sw
tri 37087 36583 37088 36584 ne
rect 37088 36583 39060 36584
rect 32807 36323 36791 36583
rect 28311 36293 32525 36323
rect 24848 36292 28019 36293
tri 28019 36292 28020 36293 sw
tri 28311 36292 28312 36293 ne
rect 28312 36292 32525 36293
rect 24848 36000 28020 36292
tri 28020 36000 28312 36292 sw
tri 28312 36000 28604 36292 ne
rect 28604 36129 32525 36292
tri 32525 36129 32719 36323 sw
tri 32807 36129 33001 36323 ne
rect 33001 36286 36791 36323
tri 36791 36286 37088 36583 sw
tri 37088 36286 37385 36583 ne
rect 37385 36500 39060 36583
tri 39060 36500 39151 36591 sw
tri 39349 36500 39440 36591 ne
rect 39440 36500 41130 36591
tri 41130 36500 41420 36790 sw
tri 41420 36500 41710 36790 ne
rect 41710 36654 45506 36790
tri 45506 36654 45800 36948 sw
tri 45800 36654 46094 36948 ne
rect 46094 36868 49836 36948
tri 49836 36868 50124 37156 sw
tri 50124 36868 50412 37156 ne
rect 50412 37147 54131 37156
tri 54131 37147 54377 37393 sw
tri 54428 37147 54674 37393 ne
rect 54674 37147 71000 37393
rect 50412 37095 54377 37147
tri 54377 37095 54429 37147 sw
tri 54674 37095 54726 37147 ne
rect 54726 37095 71000 37147
rect 50412 36868 54429 37095
rect 46094 36665 50124 36868
tri 50124 36665 50327 36868 sw
tri 50412 36665 50615 36868 ne
rect 50615 36798 54429 36868
tri 54429 36798 54726 37095 sw
tri 54726 36798 55023 37095 ne
rect 55023 36798 71000 37095
rect 50615 36797 54726 36798
tri 54726 36797 54727 36798 sw
tri 55023 36797 55024 36798 ne
rect 55024 36797 71000 36798
rect 50615 36665 54727 36797
rect 46094 36654 50327 36665
rect 41710 36653 45800 36654
tri 45800 36653 45801 36654 sw
tri 46094 36653 46095 36654 ne
rect 46095 36653 50327 36654
rect 41710 36500 45801 36653
rect 37385 36286 39151 36500
rect 33001 36129 37088 36286
tri 37088 36129 37245 36286 sw
tri 37385 36129 37542 36286 ne
rect 37542 36211 39151 36286
tri 39151 36211 39440 36500 sw
tri 39440 36211 39729 36500 ne
rect 39729 36499 41420 36500
tri 41420 36499 41421 36500 sw
tri 41710 36499 41711 36500 ne
rect 41711 36499 45801 36500
rect 39729 36211 41421 36499
rect 37542 36129 39440 36211
rect 28604 36000 32719 36129
rect 24848 35999 28312 36000
tri 28312 35999 28313 36000 sw
tri 28604 35999 28605 36000 ne
rect 28605 35999 32719 36000
rect 24848 35707 28313 35999
tri 28313 35707 28605 35999 sw
tri 28605 35707 28897 35999 ne
rect 28897 35847 32719 35999
tri 32719 35847 33001 36129 sw
tri 33001 35847 33283 36129 ne
rect 33283 35847 37245 36129
rect 28897 35846 33001 35847
tri 33001 35846 33002 35847 sw
tri 33283 35846 33284 35847 ne
rect 33284 35846 37245 35847
rect 28897 35707 33002 35846
rect 24848 35706 28605 35707
tri 28605 35706 28606 35707 sw
tri 28897 35706 28898 35707 ne
rect 28898 35706 33002 35707
rect 24848 35414 28606 35706
tri 28606 35414 28898 35706 sw
tri 28898 35414 29190 35706 ne
rect 29190 35564 33002 35706
tri 33002 35564 33284 35846 sw
tri 33284 35564 33566 35846 ne
rect 33566 35832 37245 35846
tri 37245 35832 37542 36129 sw
tri 37542 35832 37839 36129 ne
rect 37839 35922 39440 36129
tri 39440 35922 39729 36211 sw
tri 39729 35922 40018 36211 ne
rect 40018 36209 41421 36211
tri 41421 36209 41711 36499 sw
tri 41711 36209 42001 36499 ne
rect 42001 36359 45801 36499
tri 45801 36359 46095 36653 sw
tri 46095 36359 46389 36653 ne
rect 46389 36377 50327 36653
tri 50327 36377 50615 36665 sw
tri 50615 36377 50903 36665 ne
rect 50903 36500 54727 36665
tri 54727 36500 55024 36797 sw
tri 55024 36500 55321 36797 ne
rect 55321 36500 71000 36797
rect 50903 36499 55024 36500
tri 55024 36499 55025 36500 sw
tri 55321 36499 55322 36500 ne
rect 55322 36499 71000 36500
rect 50903 36377 55025 36499
rect 46389 36359 50615 36377
rect 42001 36358 46095 36359
tri 46095 36358 46096 36359 sw
tri 46389 36358 46390 36359 ne
rect 46390 36358 50615 36359
rect 42001 36209 46096 36358
rect 40018 35922 41711 36209
rect 37839 35832 39729 35922
rect 33566 35831 37542 35832
tri 37542 35831 37543 35832 sw
tri 37839 35831 37840 35832 ne
rect 37840 35831 39729 35832
rect 33566 35564 37543 35831
rect 29190 35563 33284 35564
tri 33284 35563 33285 35564 sw
tri 33566 35563 33567 35564 ne
rect 33567 35563 37543 35564
rect 29190 35414 33285 35563
rect 24848 35220 28898 35414
tri 28898 35220 29092 35414 sw
tri 29190 35220 29384 35414 ne
rect 29384 35281 33285 35414
tri 33285 35281 33567 35563 sw
tri 33567 35281 33849 35563 ne
rect 33849 35534 37543 35563
tri 37543 35534 37840 35831 sw
tri 37840 35534 38137 35831 ne
rect 38137 35767 39729 35831
tri 39729 35767 39884 35922 sw
tri 40018 35767 40173 35922 ne
rect 40173 35919 41711 35922
tri 41711 35919 42001 36209 sw
tri 42001 35919 42291 36209 ne
rect 42291 36064 46096 36209
tri 46096 36064 46390 36358 sw
tri 46390 36064 46684 36358 ne
rect 46684 36201 50615 36358
tri 50615 36201 50791 36377 sw
tri 50903 36201 51079 36377 ne
rect 51079 36202 55025 36377
tri 55025 36202 55322 36499 sw
tri 55322 36400 55421 36499 ne
rect 55421 36400 71000 36499
rect 51079 36201 55322 36202
rect 46684 36064 50791 36201
rect 42291 36063 46390 36064
tri 46390 36063 46391 36064 sw
tri 46684 36063 46685 36064 ne
rect 46685 36063 50791 36064
rect 42291 35919 46391 36063
rect 40173 35918 42001 35919
tri 42001 35918 42002 35919 sw
tri 42291 35918 42292 35919 ne
rect 42292 35918 46391 35919
rect 40173 35767 42002 35918
rect 38137 35534 39884 35767
rect 33849 35281 37840 35534
rect 29384 35279 33567 35281
tri 33567 35279 33569 35281 sw
tri 33849 35279 33851 35281 ne
rect 33851 35279 37840 35281
rect 29384 35220 33569 35279
tri 24848 30976 29092 35220 ne
tri 29092 34928 29384 35220 sw
tri 29384 34928 29676 35220 ne
rect 29676 34997 33569 35220
tri 33569 34997 33851 35279 sw
tri 33851 34997 34133 35279 ne
rect 34133 35237 37840 35279
tri 37840 35237 38137 35534 sw
tri 38137 35237 38434 35534 ne
rect 38434 35478 39884 35534
tri 39884 35478 40173 35767 sw
tri 40173 35478 40462 35767 ne
rect 40462 35628 42002 35767
tri 42002 35628 42292 35918 sw
tri 42292 35628 42582 35918 ne
rect 42582 35769 46391 35918
tri 46391 35769 46685 36063 sw
tri 46685 35769 46979 36063 ne
rect 46979 35913 50791 36063
tri 50791 35913 51079 36201 sw
tri 51079 35913 51367 36201 ne
rect 51367 36200 55322 36201
tri 55322 36200 55324 36202 sw
rect 51367 35913 71000 36200
rect 46979 35911 51079 35913
tri 51079 35911 51081 35913 sw
tri 51367 35911 51369 35913 ne
rect 51369 35911 71000 35913
rect 46979 35769 51081 35911
rect 42582 35767 46685 35769
tri 46685 35767 46687 35769 sw
tri 46979 35767 46981 35769 ne
rect 46981 35767 51081 35769
rect 42582 35628 46687 35767
rect 40462 35478 42292 35628
rect 38434 35237 40173 35478
rect 34133 34997 38137 35237
rect 29676 34996 33851 34997
tri 33851 34996 33852 34997 sw
tri 34133 34996 34134 34997 ne
rect 34134 34996 38137 34997
rect 29676 34928 33852 34996
rect 29092 34851 29384 34928
tri 29384 34851 29461 34928 sw
tri 29676 34851 29753 34928 ne
rect 29753 34851 33852 34928
rect 29092 34559 29461 34851
tri 29461 34559 29753 34851 sw
tri 29753 34559 30045 34851 ne
rect 30045 34714 33852 34851
tri 33852 34714 34134 34996 sw
tri 34134 34714 34416 34996 ne
rect 34416 34940 38137 34996
tri 38137 34940 38434 35237 sw
tri 38434 34940 38731 35237 ne
rect 38731 35189 40173 35237
tri 40173 35189 40462 35478 sw
tri 40462 35189 40751 35478 ne
rect 40751 35392 42292 35478
tri 42292 35392 42528 35628 sw
tri 42582 35392 42818 35628 ne
rect 42818 35474 46687 35628
tri 46687 35474 46980 35767 sw
tri 46981 35474 47274 35767 ne
rect 47274 35623 51081 35767
tri 51081 35623 51369 35911 sw
tri 51369 35623 51657 35911 ne
rect 51657 35623 71000 35911
rect 47274 35622 51369 35623
tri 51369 35622 51370 35623 sw
tri 51657 35622 51658 35623 ne
rect 51658 35622 71000 35623
rect 47274 35474 51370 35622
rect 42818 35392 46980 35474
rect 40751 35288 42528 35392
tri 42528 35288 42632 35392 sw
tri 42818 35288 42922 35392 ne
rect 42922 35288 46980 35392
rect 40751 35189 42632 35288
rect 38731 34940 40462 35189
rect 34416 34901 38434 34940
tri 38434 34901 38473 34940 sw
tri 38731 34901 38770 34940 ne
rect 38770 34901 40462 34940
rect 34416 34714 38473 34901
rect 30045 34713 34134 34714
tri 34134 34713 34135 34714 sw
tri 34416 34713 34417 34714 ne
rect 34417 34713 38473 34714
rect 30045 34559 34135 34713
rect 29092 34558 29753 34559
tri 29753 34558 29754 34559 sw
tri 30045 34558 30046 34559 ne
rect 30046 34558 34135 34559
rect 29092 34266 29754 34558
tri 29754 34266 30046 34558 sw
tri 30046 34266 30338 34558 ne
rect 30338 34431 34135 34558
tri 34135 34431 34417 34713 sw
tri 34417 34431 34699 34713 ne
rect 34699 34604 38473 34713
tri 38473 34604 38770 34901 sw
tri 38770 34604 39067 34901 ne
rect 39067 34900 40462 34901
tri 40462 34900 40751 35189 sw
tri 40751 34900 41040 35189 ne
rect 41040 34998 42632 35189
tri 42632 34998 42922 35288 sw
tri 42922 34998 43212 35288 ne
rect 43212 35224 46980 35288
tri 46980 35224 47230 35474 sw
tri 47274 35224 47524 35474 ne
rect 47524 35334 51370 35474
tri 51370 35334 51658 35622 sw
tri 51658 35334 51946 35622 ne
rect 51946 35334 71000 35622
rect 47524 35333 51658 35334
tri 51658 35333 51659 35334 sw
tri 51946 35333 51947 35334 ne
rect 51947 35333 71000 35334
rect 47524 35224 51659 35333
rect 43212 34998 47230 35224
rect 41040 34900 42922 34998
rect 39067 34611 40751 34900
tri 40751 34611 41040 34900 sw
tri 41040 34611 41329 34900 ne
rect 41329 34810 42922 34900
tri 42922 34810 43110 34998 sw
tri 43212 34810 43400 34998 ne
rect 43400 34994 47230 34998
tri 47230 34994 47460 35224 sw
tri 47524 34994 47754 35224 ne
rect 47754 35045 51659 35224
tri 51659 35045 51947 35333 sw
tri 51947 35045 52235 35333 ne
rect 52235 35045 71000 35333
rect 47754 35044 51947 35045
tri 51947 35044 51948 35045 sw
tri 52235 35044 52236 35045 ne
rect 52236 35044 71000 35045
rect 47754 34994 51948 35044
rect 43400 34929 47460 34994
tri 47460 34929 47525 34994 sw
tri 47754 34929 47819 34994 ne
rect 47819 34929 51948 34994
rect 43400 34810 47525 34929
rect 41329 34611 43110 34810
rect 39067 34604 41040 34611
rect 34699 34603 38770 34604
tri 38770 34603 38771 34604 sw
tri 39067 34603 39068 34604 ne
rect 39068 34603 41040 34604
rect 34699 34431 38771 34603
rect 30338 34266 34417 34431
rect 29092 34265 30046 34266
tri 30046 34265 30047 34266 sw
tri 30338 34265 30339 34266 ne
rect 30339 34265 34417 34266
rect 29092 33973 30047 34265
tri 30047 33973 30339 34265 sw
tri 30339 33973 30631 34265 ne
rect 30631 34176 34417 34265
tri 34417 34176 34672 34431 sw
tri 34699 34176 34954 34431 ne
rect 34954 34306 38771 34431
tri 38771 34306 39068 34603 sw
tri 39068 34306 39365 34603 ne
rect 39365 34520 41040 34603
tri 41040 34520 41131 34611 sw
tri 41329 34520 41420 34611 ne
rect 41420 34520 43110 34611
tri 43110 34520 43400 34810 sw
tri 43400 34520 43690 34810 ne
rect 43690 34635 47525 34810
tri 47525 34635 47819 34929 sw
tri 47819 34635 48113 34929 ne
rect 48113 34756 51948 34929
tri 51948 34756 52236 35044 sw
tri 52236 34756 52524 35044 ne
rect 52524 34756 71000 35044
rect 48113 34755 52236 34756
tri 52236 34755 52237 34756 sw
tri 52524 34755 52525 34756 ne
rect 52525 34755 71000 34756
rect 48113 34635 52237 34755
rect 43690 34634 47819 34635
tri 47819 34634 47820 34635 sw
tri 48113 34634 48114 34635 ne
rect 48114 34634 52237 34635
rect 43690 34520 47820 34634
rect 39365 34306 41131 34520
rect 34954 34305 39068 34306
tri 39068 34305 39069 34306 sw
tri 39365 34305 39366 34306 ne
rect 39366 34305 41131 34306
rect 34954 34176 39069 34305
rect 30631 33973 34672 34176
rect 29092 33884 30339 33973
tri 30339 33884 30428 33973 sw
tri 30631 33884 30720 33973 ne
rect 30720 33894 34672 33973
tri 34672 33894 34954 34176 sw
tri 34954 33894 35236 34176 ne
rect 35236 34008 39069 34176
tri 39069 34008 39366 34305 sw
tri 39366 34008 39663 34305 ne
rect 39663 34231 41131 34305
tri 41131 34231 41420 34520 sw
tri 41420 34231 41709 34520 ne
rect 41709 34519 43400 34520
tri 43400 34519 43401 34520 sw
tri 43690 34519 43691 34520 ne
rect 43691 34519 47820 34520
rect 41709 34231 43401 34519
rect 39663 34008 41420 34231
rect 35236 33894 39366 34008
rect 30720 33884 34954 33894
rect 29092 33592 30428 33884
tri 30428 33592 30720 33884 sw
tri 30720 33592 31012 33884 ne
rect 31012 33779 34954 33884
tri 34954 33779 35069 33894 sw
tri 35236 33779 35351 33894 ne
rect 35351 33779 39366 33894
rect 31012 33592 35069 33779
rect 29092 33385 30720 33592
tri 30720 33385 30927 33592 sw
tri 31012 33385 31219 33592 ne
rect 31219 33497 35069 33592
tri 35069 33497 35351 33779 sw
tri 35351 33497 35633 33779 ne
rect 35633 33711 39366 33779
tri 39366 33711 39663 34008 sw
tri 39663 33711 39960 34008 ne
rect 39960 33942 41420 34008
tri 41420 33942 41709 34231 sw
tri 41709 33942 41998 34231 ne
rect 41998 34229 43401 34231
tri 43401 34229 43691 34519 sw
tri 43691 34229 43981 34519 ne
rect 43981 34340 47820 34519
tri 47820 34340 48114 34634 sw
tri 48114 34340 48408 34634 ne
rect 48408 34467 52237 34634
tri 52237 34467 52525 34755 sw
tri 52525 34467 52813 34755 ne
rect 52813 34467 71000 34755
rect 48408 34340 52525 34467
rect 43981 34339 48114 34340
tri 48114 34339 48115 34340 sw
tri 48408 34339 48409 34340 ne
rect 48409 34339 52525 34340
rect 43981 34229 48115 34339
rect 41998 34042 43691 34229
tri 43691 34042 43878 34229 sw
tri 43981 34042 44168 34229 ne
rect 44168 34045 48115 34229
tri 48115 34045 48409 34339 sw
tri 48409 34045 48703 34339 ne
rect 48703 34244 52525 34339
tri 52525 34244 52748 34467 sw
tri 52813 34244 53036 34467 ne
rect 53036 34244 71000 34467
rect 48703 34045 52748 34244
rect 44168 34042 48409 34045
rect 41998 33942 43878 34042
rect 39960 33787 41709 33942
tri 41709 33787 41864 33942 sw
tri 41998 33787 42153 33942 ne
rect 42153 33787 43878 33942
rect 39960 33711 41864 33787
rect 35633 33516 39663 33711
tri 39663 33516 39858 33711 sw
tri 39960 33516 40155 33711 ne
rect 40155 33516 41864 33711
rect 35633 33497 39858 33516
rect 31219 33495 35351 33497
tri 35351 33495 35353 33497 sw
tri 35633 33495 35635 33497 ne
rect 35635 33495 39858 33497
rect 31219 33385 35353 33495
rect 29092 33094 30927 33385
tri 30927 33094 31218 33385 sw
tri 31219 33094 31510 33385 ne
rect 31510 33213 35353 33385
tri 35353 33213 35635 33495 sw
tri 35635 33213 35917 33495 ne
rect 35917 33219 39858 33495
tri 39858 33219 40155 33516 sw
tri 40155 33219 40452 33516 ne
rect 40452 33498 41864 33516
tri 41864 33498 42153 33787 sw
tri 42153 33498 42442 33787 ne
rect 42442 33752 43878 33787
tri 43878 33752 44168 34042 sw
tri 44168 33752 44458 34042 ne
rect 44458 33950 48409 34042
tri 48409 33950 48504 34045 sw
tri 48703 33950 48798 34045 ne
rect 48798 33956 52748 34045
tri 52748 33956 53036 34244 sw
tri 53036 33956 53324 34244 ne
rect 53324 33956 71000 34244
rect 48798 33950 53036 33956
rect 44458 33752 48504 33950
rect 42442 33498 44168 33752
rect 40452 33219 42153 33498
rect 35917 33213 40155 33219
rect 31510 33212 35635 33213
tri 35635 33212 35636 33213 sw
tri 35917 33212 35918 33213 ne
rect 35918 33212 40155 33213
rect 31510 33094 35636 33212
rect 29092 32929 31218 33094
tri 31218 32929 31383 33094 sw
tri 31510 32929 31675 33094 ne
rect 31675 32930 35636 33094
tri 35636 32930 35918 33212 sw
tri 35918 32930 36200 33212 ne
rect 36200 32930 40155 33212
rect 31675 32929 35918 32930
rect 29092 32637 31383 32929
tri 31383 32637 31675 32929 sw
tri 31675 32637 31967 32929 ne
rect 31967 32850 35918 32929
tri 35918 32850 35998 32930 sw
tri 36200 32850 36280 32930 ne
rect 36280 32922 40155 32930
tri 40155 32922 40452 33219 sw
tri 40452 32922 40749 33219 ne
rect 40749 33209 42153 33219
tri 42153 33209 42442 33498 sw
tri 42442 33209 42731 33498 ne
rect 42731 33462 44168 33498
tri 44168 33462 44458 33752 sw
tri 44458 33462 44748 33752 ne
rect 44748 33656 48504 33752
tri 48504 33656 48798 33950 sw
tri 48798 33656 49092 33950 ne
rect 49092 33868 53036 33950
tri 53036 33868 53124 33956 sw
tri 53324 33868 53412 33956 ne
rect 53412 33868 71000 33956
rect 49092 33656 53124 33868
rect 44748 33462 48798 33656
rect 42731 33411 44458 33462
tri 44458 33411 44509 33462 sw
tri 44748 33411 44799 33462 ne
rect 44799 33453 48798 33462
tri 48798 33453 49001 33656 sw
tri 49092 33453 49295 33656 ne
rect 49295 33580 53124 33656
tri 53124 33580 53412 33868 sw
tri 53412 33580 53700 33868 ne
rect 53700 33580 71000 33868
rect 49295 33579 53412 33580
tri 53412 33579 53413 33580 sw
tri 53700 33579 53701 33580 ne
rect 53701 33579 71000 33580
rect 49295 33453 53413 33579
rect 44799 33411 49001 33453
rect 42731 33209 44509 33411
rect 40749 32922 42442 33209
rect 36280 32920 40452 32922
tri 40452 32920 40454 32922 sw
tri 40749 32920 40751 32922 ne
rect 40751 32920 42442 32922
tri 42442 32920 42731 33209 sw
tri 42731 32920 43020 33209 ne
rect 43020 33121 44509 33209
tri 44509 33121 44799 33411 sw
tri 44799 33121 45089 33411 ne
rect 45089 33159 49001 33411
tri 49001 33159 49295 33453 sw
tri 49295 33159 49589 33453 ne
rect 49589 33291 53413 33453
tri 53413 33291 53701 33579 sw
tri 53701 33291 53989 33579 ne
rect 53989 33291 71000 33579
rect 49589 33290 53701 33291
tri 53701 33290 53702 33291 sw
tri 53989 33290 53990 33291 ne
rect 53990 33290 71000 33291
rect 49589 33159 53702 33290
rect 45089 33121 49295 33159
rect 43020 32920 44799 33121
rect 36280 32850 40454 32920
rect 31967 32637 35998 32850
rect 29092 32636 31675 32637
tri 31675 32636 31676 32637 sw
tri 31967 32636 31968 32637 ne
rect 31968 32636 35998 32637
rect 29092 32344 31676 32636
tri 31676 32344 31968 32636 sw
tri 31968 32344 32260 32636 ne
rect 32260 32568 35998 32636
tri 35998 32568 36280 32850 sw
tri 36280 32568 36562 32850 ne
rect 36562 32623 40454 32850
tri 40454 32623 40751 32920 sw
tri 40751 32623 41048 32920 ne
rect 41048 32631 42731 32920
tri 42731 32631 43020 32920 sw
tri 43020 32631 43309 32920 ne
rect 43309 32831 44799 32920
tri 44799 32831 45089 33121 sw
tri 45089 32831 45379 33121 ne
rect 45379 33001 49295 33121
tri 49295 33001 49453 33159 sw
tri 49589 33001 49747 33159 ne
rect 49747 33002 53702 33159
tri 53702 33002 53990 33290 sw
tri 53990 33200 54080 33290 ne
rect 54080 33200 71000 33290
rect 49747 33001 53990 33002
rect 45379 32831 49453 33001
rect 43309 32830 45089 32831
tri 45089 32830 45090 32831 sw
tri 45379 32830 45380 32831 ne
rect 45380 32830 49453 32831
rect 43309 32631 45090 32830
rect 41048 32623 43020 32631
rect 36562 32568 40751 32623
rect 32260 32363 36280 32568
tri 36280 32363 36485 32568 sw
tri 36562 32363 36767 32568 ne
rect 36767 32363 40751 32568
rect 32260 32344 36485 32363
rect 29092 32343 31968 32344
tri 31968 32343 31969 32344 sw
tri 32260 32343 32261 32344 ne
rect 32261 32343 36485 32344
rect 29092 32051 31969 32343
tri 31969 32051 32261 32343 sw
tri 32261 32051 32553 32343 ne
rect 32553 32081 36485 32343
tri 36485 32081 36767 32363 sw
tri 36767 32081 37049 32363 ne
rect 37049 32326 40751 32363
tri 40751 32326 41048 32623 sw
tri 41048 32326 41345 32623 ne
rect 41345 32540 43020 32623
tri 43020 32540 43111 32631 sw
tri 43309 32540 43400 32631 ne
rect 43400 32540 45090 32631
tri 45090 32540 45380 32830 sw
tri 45380 32540 45670 32830 ne
rect 45670 32707 49453 32830
tri 49453 32707 49747 33001 sw
tri 49747 32707 50041 33001 ne
rect 50041 33000 53990 33001
tri 53990 33000 53992 33002 sw
rect 50041 32707 71000 33000
rect 45670 32705 49747 32707
tri 49747 32705 49749 32707 sw
tri 50041 32705 50043 32707 ne
rect 50043 32705 71000 32707
rect 45670 32540 49749 32705
rect 41345 32326 43111 32540
rect 37049 32184 41048 32326
tri 41048 32184 41190 32326 sw
tri 41345 32184 41487 32326 ne
rect 41487 32251 43111 32326
tri 43111 32251 43400 32540 sw
tri 43400 32251 43689 32540 ne
rect 43689 32539 45380 32540
tri 45380 32539 45381 32540 sw
tri 45670 32539 45671 32540 ne
rect 45671 32539 49749 32540
rect 43689 32251 45381 32539
rect 41487 32184 43400 32251
rect 37049 32081 41190 32184
rect 32553 32051 36767 32081
rect 29092 32049 32261 32051
tri 32261 32049 32263 32051 sw
tri 32553 32049 32555 32051 ne
rect 32555 32049 36767 32051
rect 29092 31757 32263 32049
tri 32263 31757 32555 32049 sw
tri 32555 31757 32847 32049 ne
rect 32847 31886 36767 32049
tri 36767 31886 36962 32081 sw
tri 37049 31886 37244 32081 ne
rect 37244 31887 41190 32081
tri 41190 31887 41487 32184 sw
tri 41487 31887 41784 32184 ne
rect 41784 31962 43400 32184
tri 43400 31962 43689 32251 sw
tri 43689 31962 43978 32251 ne
rect 43978 32249 45381 32251
tri 45381 32249 45671 32539 sw
tri 45671 32249 45961 32539 ne
rect 45961 32411 49749 32539
tri 49749 32411 50043 32705 sw
tri 50043 32411 50337 32705 ne
rect 50337 32411 71000 32705
rect 45961 32410 50043 32411
tri 50043 32410 50044 32411 sw
tri 50337 32410 50338 32411 ne
rect 50338 32410 71000 32411
rect 45961 32249 50044 32410
rect 43978 31962 45671 32249
rect 41784 31887 43689 31962
rect 37244 31886 41487 31887
tri 41487 31886 41488 31887 sw
tri 41784 31886 41785 31887 ne
rect 41785 31886 43689 31887
rect 32847 31757 36962 31886
rect 29092 31756 32555 31757
tri 32555 31756 32556 31757 sw
tri 32847 31756 32848 31757 ne
rect 32848 31756 36962 31757
rect 29092 31464 32556 31756
tri 32556 31464 32848 31756 sw
tri 32848 31464 33140 31756 ne
rect 33140 31604 36962 31756
tri 36962 31604 37244 31886 sw
tri 37244 31604 37526 31886 ne
rect 37526 31604 41488 31886
rect 33140 31603 37244 31604
tri 37244 31603 37245 31604 sw
tri 37526 31603 37527 31604 ne
rect 37527 31603 41488 31604
rect 33140 31464 37245 31603
rect 29092 31463 32848 31464
tri 32848 31463 32849 31464 sw
tri 33140 31463 33141 31464 ne
rect 33141 31463 37245 31464
rect 29092 31171 32849 31463
tri 32849 31171 33141 31463 sw
tri 33141 31171 33433 31463 ne
rect 33433 31321 37245 31463
tri 37245 31321 37527 31603 sw
tri 37527 31321 37809 31603 ne
rect 37809 31589 41488 31603
tri 41488 31589 41785 31886 sw
tri 41785 31589 42082 31886 ne
rect 42082 31807 43689 31886
tri 43689 31807 43844 31962 sw
tri 43978 31807 44133 31962 ne
rect 44133 31959 45671 31962
tri 45671 31959 45961 32249 sw
tri 45961 31959 46251 32249 ne
rect 46251 32116 50044 32249
tri 50044 32116 50338 32410 sw
tri 50338 32116 50632 32410 ne
rect 50632 32116 71000 32410
rect 46251 32115 50338 32116
tri 50338 32115 50339 32116 sw
tri 50632 32115 50633 32116 ne
rect 50633 32115 71000 32116
rect 46251 31959 50339 32115
rect 44133 31958 45961 31959
tri 45961 31958 45962 31959 sw
tri 46251 31958 46252 31959 ne
rect 46252 31958 50339 31959
rect 44133 31807 45962 31958
rect 42082 31589 43844 31807
rect 37809 31321 41785 31589
rect 33433 31320 37527 31321
tri 37527 31320 37528 31321 sw
tri 37809 31320 37810 31321 ne
rect 37810 31320 41785 31321
rect 33433 31171 37528 31320
rect 29092 30976 33141 31171
tri 33141 30976 33336 31171 sw
tri 33433 30976 33628 31171 ne
rect 33628 31038 37528 31171
tri 37528 31038 37810 31320 sw
tri 37810 31038 38092 31320 ne
rect 38092 31292 41785 31320
tri 41785 31292 42082 31589 sw
tri 42082 31292 42379 31589 ne
rect 42379 31518 43844 31589
tri 43844 31518 44133 31807 sw
tri 44133 31518 44422 31807 ne
rect 44422 31668 45962 31807
tri 45962 31668 46252 31958 sw
tri 46252 31668 46542 31958 ne
rect 46542 31821 50339 31958
tri 50339 31821 50633 32115 sw
tri 50633 31821 50927 32115 ne
rect 50927 31821 71000 32115
rect 46542 31820 50633 31821
tri 50633 31820 50634 31821 sw
tri 50927 31820 50928 31821 ne
rect 50928 31820 71000 31821
rect 46542 31668 50634 31820
rect 44422 31518 46252 31668
rect 42379 31292 44133 31518
rect 38092 31291 42082 31292
tri 42082 31291 42083 31292 sw
tri 42379 31291 42380 31292 ne
rect 42380 31291 44133 31292
rect 38092 31038 42083 31291
rect 33628 31037 37810 31038
tri 37810 31037 37811 31038 sw
tri 38092 31037 38093 31038 ne
rect 38093 31037 42083 31038
rect 33628 30976 37811 31037
tri 29092 26732 33336 30976 ne
tri 33336 30684 33628 30976 sw
tri 33628 30684 33920 30976 ne
rect 33920 30755 37811 30976
tri 37811 30755 38093 31037 sw
tri 38093 30755 38375 31037 ne
rect 38375 30994 42083 31037
tri 42083 30994 42380 31291 sw
tri 42380 30994 42677 31291 ne
rect 42677 31229 44133 31291
tri 44133 31229 44422 31518 sw
tri 44422 31229 44711 31518 ne
rect 44711 31431 46252 31518
tri 46252 31431 46489 31668 sw
tri 46542 31431 46779 31668 ne
rect 46779 31526 50634 31668
tri 50634 31526 50928 31820 sw
tri 50928 31526 51222 31820 ne
rect 51222 31526 71000 31820
rect 46779 31525 50928 31526
tri 50928 31525 50929 31526 sw
tri 51222 31525 51223 31526 ne
rect 51223 31525 71000 31526
rect 46779 31431 50929 31525
rect 44711 31229 46489 31431
rect 42677 30994 44422 31229
rect 38375 30940 42380 30994
tri 42380 30940 42434 30994 sw
tri 42677 30940 42731 30994 ne
rect 42731 30940 44422 30994
tri 44422 30940 44711 31229 sw
tri 44711 30940 45000 31229 ne
rect 45000 31141 46489 31229
tri 46489 31141 46779 31431 sw
tri 46779 31141 47069 31431 ne
rect 47069 31231 50929 31431
tri 50929 31231 51223 31525 sw
tri 51223 31231 51517 31525 ne
rect 51517 31231 71000 31525
rect 47069 31141 51223 31231
rect 45000 31044 46779 31141
tri 46779 31044 46876 31141 sw
tri 47069 31044 47166 31141 ne
rect 47166 31044 51223 31141
rect 45000 30940 46876 31044
rect 38375 30755 42434 30940
rect 33920 30753 38093 30755
tri 38093 30753 38095 30755 sw
tri 38375 30753 38377 30755 ne
rect 38377 30753 42434 30755
rect 33920 30684 38095 30753
rect 33336 30609 33628 30684
tri 33628 30609 33703 30684 sw
tri 33920 30609 33995 30684 ne
rect 33995 30609 38095 30684
rect 33336 30317 33703 30609
tri 33703 30317 33995 30609 sw
tri 33995 30317 34287 30609 ne
rect 34287 30471 38095 30609
tri 38095 30471 38377 30753 sw
tri 38377 30471 38659 30753 ne
rect 38659 30643 42434 30753
tri 42434 30643 42731 30940 sw
tri 42731 30643 43028 30940 ne
rect 43028 30651 44711 30940
tri 44711 30651 45000 30940 sw
tri 45000 30651 45289 30940 ne
rect 45289 30754 46876 30940
tri 46876 30754 47166 31044 sw
tri 47166 30754 47456 31044 ne
rect 47456 30981 51223 31044
tri 51223 30981 51473 31231 sw
tri 51517 30981 51767 31231 ne
rect 51767 30981 71000 31231
rect 47456 30754 51473 30981
rect 45289 30651 47166 30754
rect 43028 30643 45000 30651
rect 38659 30471 42731 30643
rect 34287 30317 38377 30471
rect 33336 30315 33995 30317
tri 33995 30315 33997 30317 sw
tri 34287 30315 34289 30317 ne
rect 34289 30315 38377 30317
rect 33336 30023 33997 30315
tri 33997 30023 34289 30315 sw
tri 34289 30023 34581 30315 ne
rect 34581 30189 38377 30315
tri 38377 30189 38659 30471 sw
tri 38659 30189 38941 30471 ne
rect 38941 30346 42731 30471
tri 42731 30346 43028 30643 sw
tri 43028 30346 43325 30643 ne
rect 43325 30560 45000 30643
tri 45000 30560 45091 30651 sw
tri 45289 30560 45380 30651 ne
rect 45380 30560 47166 30651
rect 43325 30346 45091 30560
rect 38941 30345 43028 30346
tri 43028 30345 43029 30346 sw
tri 43325 30345 43326 30346 ne
rect 43326 30345 45091 30346
rect 38941 30189 43029 30345
rect 34581 30023 38659 30189
rect 33336 30022 34289 30023
tri 34289 30022 34290 30023 sw
tri 34581 30022 34582 30023 ne
rect 34582 30022 38659 30023
rect 33336 29730 34290 30022
tri 34290 29730 34582 30022 sw
tri 34582 29730 34874 30022 ne
rect 34874 29932 38659 30022
tri 38659 29932 38916 30189 sw
tri 38941 29932 39198 30189 ne
rect 39198 30048 43029 30189
tri 43029 30048 43326 30345 sw
tri 43326 30048 43623 30345 ne
rect 43623 30271 45091 30345
tri 45091 30271 45380 30560 sw
tri 45380 30271 45669 30560 ne
rect 45669 30559 47166 30560
tri 47166 30559 47361 30754 sw
tri 47456 30559 47651 30754 ne
rect 47651 30750 51473 30754
tri 51473 30750 51704 30981 sw
tri 51767 30750 51998 30981 ne
rect 51998 30750 71000 30981
rect 47651 30686 51704 30750
tri 51704 30686 51768 30750 sw
tri 51998 30686 52062 30750 ne
rect 52062 30686 71000 30750
rect 47651 30559 51768 30686
rect 45669 30271 47361 30559
rect 43623 30048 45380 30271
rect 39198 29932 43326 30048
rect 34874 29730 38916 29932
rect 33336 29640 34582 29730
tri 34582 29640 34672 29730 sw
tri 34874 29640 34964 29730 ne
rect 34964 29650 38916 29730
tri 38916 29650 39198 29932 sw
tri 39198 29650 39480 29932 ne
rect 39480 29751 43326 29932
tri 43326 29751 43623 30048 sw
tri 43623 29751 43920 30048 ne
rect 43920 29982 45380 30048
tri 45380 29982 45669 30271 sw
tri 45669 29982 45958 30271 ne
rect 45958 30269 47361 30271
tri 47361 30269 47651 30559 sw
tri 47651 30269 47941 30559 ne
rect 47941 30392 51768 30559
tri 51768 30392 52062 30686 sw
tri 52062 30392 52356 30686 ne
rect 52356 30392 71000 30686
rect 47941 30391 52062 30392
tri 52062 30391 52063 30392 sw
tri 52356 30391 52357 30392 ne
rect 52357 30391 71000 30392
rect 47941 30269 52063 30391
rect 45958 30090 47651 30269
tri 47651 30090 47830 30269 sw
tri 47941 30090 48120 30269 ne
rect 48120 30097 52063 30269
tri 52063 30097 52357 30391 sw
tri 52357 30097 52651 30391 ne
rect 52651 30097 71000 30391
rect 48120 30096 52357 30097
tri 52357 30096 52358 30097 sw
tri 52651 30096 52652 30097 ne
rect 52652 30096 71000 30097
rect 48120 30090 52358 30096
rect 45958 29982 47830 30090
rect 43920 29827 45669 29982
tri 45669 29827 45824 29982 sw
tri 45958 29827 46113 29982 ne
rect 46113 29827 47830 29982
rect 43920 29751 45824 29827
rect 39480 29650 43623 29751
rect 34964 29640 39198 29650
rect 33336 29348 34672 29640
tri 34672 29348 34964 29640 sw
tri 34964 29348 35256 29640 ne
rect 35256 29536 39198 29640
tri 39198 29536 39312 29650 sw
tri 39480 29536 39594 29650 ne
rect 39594 29556 43623 29650
tri 43623 29556 43818 29751 sw
tri 43920 29556 44115 29751 ne
rect 44115 29556 45824 29751
rect 39594 29536 43818 29556
rect 35256 29348 39312 29536
rect 33336 29143 34964 29348
tri 34964 29143 35169 29348 sw
tri 35256 29143 35461 29348 ne
rect 35461 29254 39312 29348
tri 39312 29254 39594 29536 sw
tri 39594 29254 39876 29536 ne
rect 39876 29259 43818 29536
tri 43818 29259 44115 29556 sw
tri 44115 29259 44412 29556 ne
rect 44412 29538 45824 29556
tri 45824 29538 46113 29827 sw
tri 46113 29538 46402 29827 ne
rect 46402 29800 47830 29827
tri 47830 29800 48120 30090 sw
tri 48120 29800 48410 30090 ne
rect 48410 29802 52358 30090
tri 52358 29802 52652 30096 sw
tri 52652 30000 52748 30096 ne
rect 52748 30000 71000 30096
rect 48410 29800 52652 29802
tri 52652 29800 52654 29802 sw
rect 46402 29799 48120 29800
tri 48120 29799 48121 29800 sw
tri 48410 29799 48411 29800 ne
rect 48411 29799 71000 29800
rect 46402 29538 48121 29799
rect 44412 29259 46113 29538
rect 39876 29258 44115 29259
tri 44115 29258 44116 29259 sw
tri 44412 29258 44413 29259 ne
rect 44413 29258 46113 29259
rect 39876 29254 44116 29258
rect 35461 29253 39594 29254
tri 39594 29253 39595 29254 sw
tri 39876 29253 39877 29254 ne
rect 39877 29253 44116 29254
rect 35461 29143 39595 29253
rect 33336 28851 35169 29143
tri 35169 28851 35461 29143 sw
tri 35461 28851 35753 29143 ne
rect 35753 28971 39595 29143
tri 39595 28971 39877 29253 sw
tri 39877 28971 40159 29253 ne
rect 40159 28971 44116 29253
rect 35753 28969 39877 28971
tri 39877 28969 39879 28971 sw
tri 40159 28969 40161 28971 ne
rect 40161 28969 44116 28971
rect 35753 28851 39879 28969
rect 33336 28686 35461 28851
tri 35461 28686 35626 28851 sw
tri 35753 28686 35918 28851 ne
rect 35918 28688 39879 28851
tri 39879 28688 40160 28969 sw
tri 40161 28688 40442 28969 ne
rect 40442 28961 44116 28969
tri 44116 28961 44413 29258 sw
tri 44413 28961 44710 29258 ne
rect 44710 29249 46113 29258
tri 46113 29249 46402 29538 sw
tri 46402 29249 46691 29538 ne
rect 46691 29509 48121 29538
tri 48121 29509 48411 29799 sw
tri 48411 29509 48701 29799 ne
rect 48701 29509 71000 29799
rect 46691 29249 48411 29509
rect 44710 28961 46402 29249
rect 40442 28688 44413 28961
rect 35918 28686 40160 28688
rect 33336 28394 35626 28686
tri 35626 28394 35918 28686 sw
tri 35918 28394 36210 28686 ne
rect 36210 28606 40160 28686
tri 40160 28606 40242 28688 sw
tri 40442 28606 40524 28688 ne
rect 40524 28664 44413 28688
tri 44413 28664 44710 28961 sw
tri 44710 28664 45007 28961 ne
rect 45007 28960 46402 28961
tri 46402 28960 46691 29249 sw
tri 46691 28960 46980 29249 ne
rect 46980 29219 48411 29249
tri 48411 29219 48701 29509 sw
tri 48701 29219 48991 29509 ne
rect 48991 29219 71000 29509
rect 46980 29161 48701 29219
tri 48701 29161 48759 29219 sw
tri 48991 29161 49049 29219 ne
rect 49049 29161 71000 29219
rect 46980 28960 48759 29161
rect 45007 28671 46691 28960
tri 46691 28671 46980 28960 sw
tri 46980 28671 47269 28960 ne
rect 47269 28871 48759 28960
tri 48759 28871 49049 29161 sw
tri 49049 28871 49339 29161 ne
rect 49339 28871 71000 29161
rect 47269 28870 49049 28871
tri 49049 28870 49050 28871 sw
tri 49339 28870 49340 28871 ne
rect 49340 28870 71000 28871
rect 47269 28671 49050 28870
rect 45007 28664 46980 28671
rect 40524 28662 44710 28664
tri 44710 28662 44712 28664 sw
tri 45007 28662 45009 28664 ne
rect 45009 28662 46980 28664
rect 40524 28606 44712 28662
rect 36210 28394 40242 28606
rect 33336 28393 35918 28394
tri 35918 28393 35919 28394 sw
tri 36210 28393 36211 28394 ne
rect 36211 28393 40242 28394
rect 33336 28101 35919 28393
tri 35919 28101 36211 28393 sw
tri 36211 28101 36503 28393 ne
rect 36503 28324 40242 28393
tri 40242 28324 40524 28606 sw
tri 40524 28324 40806 28606 ne
rect 40806 28365 44712 28606
tri 44712 28365 45009 28662 sw
tri 45009 28365 45306 28662 ne
rect 45306 28580 46980 28662
tri 46980 28580 47071 28671 sw
tri 47269 28580 47360 28671 ne
rect 47360 28580 49050 28671
tri 49050 28580 49340 28870 sw
tri 49340 28580 49630 28870 ne
rect 49630 28580 71000 28870
rect 45306 28365 47071 28580
rect 40806 28324 45009 28365
rect 36503 28120 40524 28324
tri 40524 28120 40728 28324 sw
tri 40806 28120 41010 28324 ne
rect 41010 28120 45009 28324
rect 36503 28101 40728 28120
rect 33336 28100 36211 28101
tri 36211 28100 36212 28101 sw
tri 36503 28100 36504 28101 ne
rect 36504 28100 40728 28101
rect 33336 27808 36212 28100
tri 36212 27808 36504 28100 sw
tri 36504 27808 36796 28100 ne
rect 36796 27838 40728 28100
tri 40728 27838 41010 28120 sw
tri 41010 27838 41292 28120 ne
rect 41292 28069 45009 28120
tri 45009 28069 45305 28365 sw
tri 45306 28069 45602 28365 ne
rect 45602 28291 47071 28365
tri 47071 28291 47360 28580 sw
tri 47360 28291 47649 28580 ne
rect 47649 28579 49340 28580
tri 49340 28579 49341 28580 sw
tri 49630 28579 49631 28580 ne
rect 49631 28579 71000 28580
rect 47649 28291 49341 28579
rect 45602 28069 47360 28291
rect 41292 27941 45305 28069
tri 45305 27941 45433 28069 sw
tri 45602 27941 45730 28069 ne
rect 45730 28002 47360 28069
tri 47360 28002 47649 28291 sw
tri 47649 28002 47938 28291 ne
rect 47938 28289 49341 28291
tri 49341 28289 49631 28579 sw
tri 49631 28289 49921 28579 ne
rect 49921 28289 71000 28579
rect 47938 28002 49631 28289
rect 45730 27941 47649 28002
rect 41292 27838 45433 27941
rect 36796 27808 41010 27838
rect 33336 27807 36504 27808
tri 36504 27807 36505 27808 sw
tri 36796 27807 36797 27808 ne
rect 36797 27807 41010 27808
rect 33336 27515 36505 27807
tri 36505 27515 36797 27807 sw
tri 36797 27515 37089 27807 ne
rect 37089 27643 41010 27807
tri 41010 27643 41205 27838 sw
tri 41292 27643 41487 27838 ne
rect 41487 27644 45433 27838
tri 45433 27644 45730 27941 sw
tri 45730 27644 46027 27941 ne
rect 46027 27847 47649 27941
tri 47649 27847 47804 28002 sw
tri 47938 27847 48093 28002 ne
rect 48093 27999 49631 28002
tri 49631 27999 49921 28289 sw
tri 49921 27999 50211 28289 ne
rect 50211 27999 71000 28289
rect 48093 27998 49921 27999
tri 49921 27998 49922 27999 sw
tri 50211 27998 50212 27999 ne
rect 50212 27998 71000 27999
rect 48093 27847 49922 27998
rect 46027 27644 47804 27847
rect 41487 27643 45730 27644
tri 45730 27643 45731 27644 sw
tri 46027 27643 46028 27644 ne
rect 46028 27643 47804 27644
rect 37089 27515 41205 27643
rect 33336 27513 36797 27515
tri 36797 27513 36799 27515 sw
tri 37089 27513 37091 27515 ne
rect 37091 27513 41205 27515
rect 33336 27221 36799 27513
tri 36799 27221 37091 27513 sw
tri 37091 27221 37383 27513 ne
rect 37383 27361 41205 27513
tri 41205 27361 41487 27643 sw
tri 41487 27361 41769 27643 ne
rect 41769 27361 45731 27643
rect 37383 27360 41487 27361
tri 41487 27360 41488 27361 sw
tri 41769 27360 41770 27361 ne
rect 41770 27360 45731 27361
rect 37383 27221 41488 27360
rect 33336 27220 37091 27221
tri 37091 27220 37092 27221 sw
tri 37383 27220 37384 27221 ne
rect 37384 27220 41488 27221
rect 33336 26928 37092 27220
tri 37092 26928 37384 27220 sw
tri 37384 26928 37676 27220 ne
rect 37676 27078 41488 27220
tri 41488 27078 41770 27360 sw
tri 41770 27078 42052 27360 ne
rect 42052 27346 45731 27360
tri 45731 27346 46028 27643 sw
tri 46028 27346 46325 27643 ne
rect 46325 27558 47804 27643
tri 47804 27558 48093 27847 sw
tri 48093 27558 48382 27847 ne
rect 48382 27708 49922 27847
tri 49922 27708 50212 27998 sw
tri 50212 27708 50502 27998 ne
rect 50502 27708 71000 27998
rect 48382 27558 50212 27708
rect 46325 27346 48093 27558
rect 42052 27078 46028 27346
rect 37676 27077 41770 27078
tri 41770 27077 41771 27078 sw
tri 42052 27077 42053 27078 ne
rect 42053 27077 46028 27078
rect 37676 26928 41771 27077
rect 33336 26732 37384 26928
tri 37384 26732 37580 26928 sw
tri 37676 26732 37872 26928 ne
rect 37872 26795 41771 26928
tri 41771 26795 42053 27077 sw
tri 42053 26795 42335 27077 ne
rect 42335 27049 46028 27077
tri 46028 27049 46325 27346 sw
tri 46325 27049 46622 27346 ne
rect 46622 27269 48093 27346
tri 48093 27269 48382 27558 sw
tri 48382 27269 48671 27558 ne
rect 48671 27471 50212 27558
tri 50212 27471 50449 27708 sw
tri 50502 27471 50739 27708 ne
rect 50739 27471 71000 27708
rect 48671 27269 50449 27471
rect 46622 27049 48382 27269
rect 42335 26981 46325 27049
tri 46325 26981 46393 27049 sw
tri 46622 26981 46690 27049 ne
rect 46690 26981 48382 27049
rect 42335 26795 46393 26981
rect 37872 26794 42053 26795
tri 42053 26794 42054 26795 sw
tri 42335 26794 42336 26795 ne
rect 42336 26794 46393 26795
rect 37872 26732 42054 26794
tri 33336 22488 37580 26732 ne
tri 37580 26440 37872 26732 sw
tri 37872 26440 38164 26732 ne
rect 38164 26512 42054 26732
tri 42054 26512 42336 26794 sw
tri 42336 26512 42618 26794 ne
rect 42618 26684 46393 26794
tri 46393 26684 46690 26981 sw
tri 46690 26684 46987 26981 ne
rect 46987 26980 48382 26981
tri 48382 26980 48671 27269 sw
tri 48671 26980 48960 27269 ne
rect 48960 27181 50449 27269
tri 50449 27181 50739 27471 sw
tri 50739 27181 51029 27471 ne
rect 51029 27181 71000 27471
rect 48960 26980 50739 27181
rect 46987 26691 48671 26980
tri 48671 26691 48960 26980 sw
tri 48960 26691 49249 26980 ne
rect 49249 26891 50739 26980
tri 50739 26891 51029 27181 sw
tri 51029 26891 51319 27181 ne
rect 51319 26891 71000 27181
rect 49249 26800 51029 26891
tri 51029 26800 51120 26891 sw
tri 51319 26800 51410 26891 ne
rect 51410 26800 71000 26891
rect 49249 26691 51120 26800
rect 46987 26684 48960 26691
rect 42618 26683 46690 26684
tri 46690 26683 46691 26684 sw
tri 46987 26683 46988 26684 ne
rect 46988 26683 48960 26684
rect 42618 26512 46691 26683
rect 38164 26511 42336 26512
tri 42336 26511 42337 26512 sw
tri 42618 26511 42619 26512 ne
rect 42619 26511 46691 26512
rect 38164 26440 42337 26511
rect 37580 26366 37872 26440
tri 37872 26366 37946 26440 sw
tri 38164 26366 38238 26440 ne
rect 38238 26366 42337 26440
rect 37580 26074 37946 26366
tri 37946 26074 38238 26366 sw
tri 38238 26074 38530 26366 ne
rect 38530 26229 42337 26366
tri 42337 26229 42619 26511 sw
tri 42619 26229 42901 26511 ne
rect 42901 26386 46691 26511
tri 46691 26386 46988 26683 sw
tri 46988 26386 47285 26683 ne
rect 47285 26600 48960 26683
tri 48960 26600 49051 26691 sw
tri 49249 26600 49340 26691 ne
rect 49340 26600 51120 26691
tri 51120 26600 51320 26800 sw
rect 47285 26386 49051 26600
rect 42901 26385 46988 26386
tri 46988 26385 46989 26386 sw
tri 47285 26385 47286 26386 ne
rect 47286 26385 49051 26386
rect 42901 26229 46989 26385
rect 38530 26227 42619 26229
tri 42619 26227 42621 26229 sw
tri 42901 26227 42903 26229 ne
rect 42903 26227 46989 26229
rect 38530 26074 42621 26227
rect 37580 26073 38238 26074
tri 38238 26073 38239 26074 sw
tri 38530 26073 38531 26074 ne
rect 38531 26073 42621 26074
rect 37580 25781 38239 26073
tri 38239 25781 38531 26073 sw
tri 38531 25781 38823 26073 ne
rect 38823 25946 42621 26073
tri 42621 25946 42902 26227 sw
tri 42903 25946 43184 26227 ne
rect 43184 26088 46989 26227
tri 46989 26088 47286 26385 sw
tri 47286 26088 47583 26385 ne
rect 47583 26311 49051 26385
tri 49051 26311 49340 26600 sw
tri 49340 26311 49629 26600 ne
rect 49629 26311 71000 26600
rect 47583 26088 49340 26311
rect 43184 25946 47286 26088
rect 38823 25781 42902 25946
rect 37580 25779 38531 25781
tri 38531 25779 38533 25781 sw
tri 38823 25779 38825 25781 ne
rect 38825 25779 42902 25781
rect 37580 25487 38533 25779
tri 38533 25487 38825 25779 sw
tri 38825 25487 39117 25779 ne
rect 39117 25688 42902 25779
tri 42902 25688 43160 25946 sw
tri 43184 25688 43442 25946 ne
rect 43442 25791 47286 25946
tri 47286 25791 47583 26088 sw
tri 47583 25791 47880 26088 ne
rect 47880 26022 49340 26088
tri 49340 26022 49629 26311 sw
tri 49629 26022 49918 26311 ne
rect 49918 26022 71000 26311
rect 47880 25867 49629 26022
tri 49629 25867 49784 26022 sw
tri 49918 25867 50073 26022 ne
rect 50073 25867 71000 26022
rect 47880 25791 49784 25867
rect 43442 25688 47583 25791
rect 39117 25487 43160 25688
rect 37580 25396 38825 25487
tri 38825 25396 38916 25487 sw
tri 39117 25396 39208 25487 ne
rect 39208 25406 43160 25487
tri 43160 25406 43442 25688 sw
tri 43442 25406 43724 25688 ne
rect 43724 25596 47583 25688
tri 47583 25596 47778 25791 sw
tri 47880 25596 48075 25791 ne
rect 48075 25596 49784 25791
rect 43724 25406 47778 25596
rect 39208 25396 43442 25406
rect 37580 25104 38916 25396
tri 38916 25104 39208 25396 sw
tri 39208 25104 39500 25396 ne
rect 39500 25293 43442 25396
tri 43442 25293 43555 25406 sw
tri 43724 25293 43837 25406 ne
rect 43837 25299 47778 25406
tri 47778 25299 48075 25596 sw
tri 48075 25299 48372 25596 ne
rect 48372 25578 49784 25596
tri 49784 25578 50073 25867 sw
tri 50073 25578 50362 25867 ne
rect 50362 25578 71000 25867
rect 48372 25299 50073 25578
rect 43837 25298 48075 25299
tri 48075 25298 48076 25299 sw
tri 48372 25298 48373 25299 ne
rect 48373 25298 50073 25299
rect 43837 25293 48076 25298
rect 39500 25104 43555 25293
rect 37580 24900 39208 25104
tri 39208 24900 39412 25104 sw
tri 39500 24900 39704 25104 ne
rect 39704 25011 43555 25104
tri 43555 25011 43837 25293 sw
tri 43837 25011 44119 25293 ne
rect 44119 25011 48076 25293
rect 39704 25010 43837 25011
tri 43837 25010 43838 25011 sw
tri 44119 25010 44120 25011 ne
rect 44120 25010 48076 25011
rect 39704 24900 43838 25010
rect 37580 24608 39412 24900
tri 39412 24608 39704 24900 sw
tri 39704 24608 39996 24900 ne
rect 39996 24728 43838 24900
tri 43838 24728 44120 25010 sw
tri 44120 24728 44402 25010 ne
rect 44402 25001 48076 25010
tri 48076 25001 48373 25298 sw
tri 48373 25001 48670 25298 ne
rect 48670 25289 50073 25298
tri 50073 25289 50362 25578 sw
tri 50362 25289 50651 25578 ne
rect 50651 25289 71000 25578
rect 48670 25001 50362 25289
rect 44402 24728 48373 25001
rect 39996 24727 44120 24728
tri 44120 24727 44121 24728 sw
tri 44402 24727 44403 24728 ne
rect 44403 24727 48373 24728
rect 39996 24608 44121 24727
rect 37580 24443 39704 24608
tri 39704 24443 39869 24608 sw
tri 39996 24443 40161 24608 ne
rect 40161 24445 44121 24608
tri 44121 24445 44403 24727 sw
tri 44403 24445 44685 24727 ne
rect 44685 24704 48373 24727
tri 48373 24704 48670 25001 sw
tri 48670 24704 48967 25001 ne
rect 48967 25000 50362 25001
tri 50362 25000 50651 25289 sw
tri 50651 25200 50740 25289 ne
rect 50740 25200 71000 25289
rect 48967 24704 71000 25000
rect 44685 24644 48670 24704
tri 48670 24644 48730 24704 sw
tri 48967 24644 49027 24704 ne
rect 49027 24644 71000 24704
rect 44685 24445 48730 24644
rect 40161 24443 44403 24445
rect 37580 24151 39869 24443
tri 39869 24151 40161 24443 sw
tri 40161 24151 40453 24443 ne
rect 40453 24362 44403 24443
tri 44403 24362 44486 24445 sw
tri 44685 24362 44768 24445 ne
rect 44768 24362 48730 24445
rect 40453 24151 44486 24362
rect 37580 24150 40161 24151
tri 40161 24150 40162 24151 sw
tri 40453 24150 40454 24151 ne
rect 40454 24150 44486 24151
rect 37580 23858 40162 24150
tri 40162 23858 40454 24150 sw
tri 40454 23858 40746 24150 ne
rect 40746 24080 44486 24150
tri 44486 24080 44768 24362 sw
tri 44768 24080 45050 24362 ne
rect 45050 24347 48730 24362
tri 48730 24347 49027 24644 sw
tri 49027 24347 49324 24644 ne
rect 49324 24347 71000 24644
rect 45050 24108 49027 24347
tri 49027 24108 49266 24347 sw
tri 49324 24108 49563 24347 ne
rect 49563 24108 71000 24347
rect 45050 24080 49266 24108
rect 40746 23877 44768 24080
tri 44768 23877 44971 24080 sw
tri 45050 23877 45253 24080 ne
rect 45253 23996 49266 24080
tri 49266 23996 49378 24108 sw
tri 49563 23996 49675 24108 ne
rect 49675 23996 71000 24108
rect 45253 23877 49378 23996
rect 40746 23858 44971 23877
rect 37580 23857 40454 23858
tri 40454 23857 40455 23858 sw
tri 40746 23857 40747 23858 ne
rect 40747 23857 44971 23858
rect 37580 23565 40455 23857
tri 40455 23565 40747 23857 sw
tri 40747 23565 41039 23857 ne
rect 41039 23595 44971 23857
tri 44971 23595 45253 23877 sw
tri 45253 23595 45535 23877 ne
rect 45535 23699 49378 23877
tri 49378 23699 49675 23996 sw
tri 49675 23699 49972 23996 ne
rect 49972 23699 71000 23996
rect 45535 23698 49675 23699
tri 49675 23698 49676 23699 sw
tri 49972 23698 49973 23699 ne
rect 49973 23698 71000 23699
rect 45535 23595 49676 23698
rect 41039 23565 45253 23595
rect 37580 23564 40747 23565
tri 40747 23564 40748 23565 sw
tri 41039 23564 41040 23565 ne
rect 41040 23564 45253 23565
rect 37580 23272 40748 23564
tri 40748 23272 41040 23564 sw
tri 41040 23272 41332 23564 ne
rect 41332 23401 45253 23564
tri 45253 23401 45447 23595 sw
tri 45535 23401 45729 23595 ne
rect 45729 23401 49676 23595
tri 49676 23401 49973 23698 sw
tri 49973 23600 50071 23698 ne
rect 50071 23600 71000 23698
rect 41332 23272 45447 23401
rect 37580 23271 41040 23272
tri 41040 23271 41041 23272 sw
tri 41332 23271 41333 23272 ne
rect 41333 23271 45447 23272
rect 37580 22979 41041 23271
tri 41041 22979 41333 23271 sw
tri 41333 22979 41625 23271 ne
rect 41625 23119 45447 23271
tri 45447 23119 45729 23401 sw
tri 45729 23119 46011 23401 ne
rect 46011 23400 49973 23401
tri 49973 23400 49974 23401 sw
rect 46011 23119 71000 23400
rect 41625 23117 45729 23119
tri 45729 23117 45731 23119 sw
tri 46011 23117 46013 23119 ne
rect 46013 23117 71000 23119
rect 41625 22979 45731 23117
rect 37580 22977 41333 22979
tri 41333 22977 41335 22979 sw
tri 41625 22977 41627 22979 ne
rect 41627 22977 45731 22979
rect 37580 22685 41335 22977
tri 41335 22685 41627 22977 sw
tri 41627 22685 41919 22977 ne
rect 41919 22835 45731 22977
tri 45731 22835 46013 23117 sw
tri 46013 22835 46295 23117 ne
rect 46295 22835 71000 23117
rect 41919 22834 46013 22835
tri 46013 22834 46014 22835 sw
tri 46295 22834 46296 22835 ne
rect 46296 22834 71000 22835
rect 41919 22685 46014 22834
rect 37580 22488 41627 22685
tri 41627 22488 41824 22685 sw
tri 41919 22488 42116 22685 ne
rect 42116 22552 46014 22685
tri 46014 22552 46296 22834 sw
tri 46296 22552 46578 22834 ne
rect 46578 22552 71000 22834
rect 42116 22551 46296 22552
tri 46296 22551 46297 22552 sw
tri 46578 22551 46579 22552 ne
rect 46579 22551 71000 22552
rect 42116 22488 46297 22551
tri 37580 18244 41824 22488 ne
tri 41824 22196 42116 22488 sw
tri 42116 22196 42408 22488 ne
rect 42408 22269 46297 22488
tri 46297 22269 46579 22551 sw
tri 46579 22269 46861 22551 ne
rect 46861 22269 71000 22551
rect 42408 22268 46579 22269
tri 46579 22268 46580 22269 sw
tri 46861 22268 46862 22269 ne
rect 46862 22268 71000 22269
rect 42408 22196 46580 22268
rect 41824 22123 42116 22196
tri 42116 22123 42189 22196 sw
tri 42408 22123 42481 22196 ne
rect 42481 22123 46580 22196
rect 41824 21831 42189 22123
tri 42189 21831 42481 22123 sw
tri 42481 21831 42773 22123 ne
rect 42773 21986 46580 22123
tri 46580 21986 46862 22268 sw
tri 46862 21986 47144 22268 ne
rect 47144 21986 71000 22268
rect 42773 21985 46862 21986
tri 46862 21985 46863 21986 sw
tri 47144 21985 47145 21986 ne
rect 47145 21985 71000 21986
rect 42773 21831 46863 21985
rect 41824 21830 42481 21831
tri 42481 21830 42482 21831 sw
tri 42773 21830 42774 21831 ne
rect 42774 21830 46863 21831
rect 41824 21538 42482 21830
tri 42482 21538 42774 21830 sw
tri 42774 21538 43066 21830 ne
rect 43066 21703 46863 21830
tri 46863 21703 47145 21985 sw
tri 47145 21703 47427 21985 ne
rect 47427 21703 71000 21985
rect 43066 21538 47145 21703
rect 41824 21537 42774 21538
tri 42774 21537 42775 21538 sw
tri 43066 21537 43067 21538 ne
rect 43067 21537 47145 21538
rect 41824 21245 42775 21537
tri 42775 21245 43067 21537 sw
tri 43067 21245 43359 21537 ne
rect 43359 21444 47145 21537
tri 47145 21444 47404 21703 sw
tri 47427 21444 47686 21703 ne
rect 47686 21444 71000 21703
rect 43359 21245 47404 21444
rect 41824 21152 43067 21245
tri 43067 21152 43160 21245 sw
tri 43359 21152 43452 21245 ne
rect 43452 21162 47404 21245
tri 47404 21162 47686 21444 sw
tri 47686 21162 47968 21444 ne
rect 47968 21162 71000 21444
rect 43452 21152 47686 21162
rect 41824 20860 43160 21152
tri 43160 20860 43452 21152 sw
tri 43452 20860 43744 21152 ne
rect 43744 21050 47686 21152
tri 47686 21050 47798 21162 sw
tri 47968 21050 48080 21162 ne
rect 48080 21050 71000 21162
rect 43744 20860 47798 21050
rect 41824 20657 43452 20860
tri 43452 20657 43655 20860 sw
tri 43744 20657 43947 20860 ne
rect 43947 20768 47798 20860
tri 47798 20768 48080 21050 sw
tri 48080 20768 48362 21050 ne
rect 48362 20768 71000 21050
rect 43947 20767 48080 20768
tri 48080 20767 48081 20768 sw
tri 48362 20767 48363 20768 ne
rect 48363 20767 71000 20768
rect 43947 20657 48081 20767
rect 41824 20365 43655 20657
tri 43655 20365 43947 20657 sw
tri 43947 20365 44239 20657 ne
rect 44239 20485 48081 20657
tri 48081 20485 48363 20767 sw
tri 48363 20485 48645 20767 ne
rect 48645 20485 71000 20767
rect 44239 20484 48363 20485
tri 48363 20484 48364 20485 sw
tri 48645 20484 48646 20485 ne
rect 48646 20484 71000 20485
rect 44239 20365 48364 20484
rect 41824 20201 43947 20365
tri 43947 20201 44111 20365 sw
tri 44239 20201 44403 20365 ne
rect 44403 20202 48364 20365
tri 48364 20202 48646 20484 sw
tri 48646 20400 48730 20484 ne
rect 48730 20400 71000 20484
rect 44403 20201 48646 20202
rect 41824 19909 44111 20201
tri 44111 19909 44403 20201 sw
tri 44403 19909 44695 20201 ne
rect 44695 20200 48646 20201
tri 48646 20200 48648 20202 sw
rect 44695 19909 71000 20200
rect 41824 19907 44403 19909
tri 44403 19907 44405 19909 sw
tri 44695 19907 44697 19909 ne
rect 44697 19907 71000 19909
rect 41824 19615 44405 19907
tri 44405 19615 44697 19907 sw
tri 44697 19615 44989 19907 ne
rect 44989 19615 71000 19907
rect 41824 19614 44697 19615
tri 44697 19614 44698 19615 sw
tri 44989 19614 44990 19615 ne
rect 44990 19614 71000 19615
rect 41824 19322 44698 19614
tri 44698 19322 44990 19614 sw
tri 44990 19322 45282 19614 ne
rect 45282 19322 71000 19614
rect 41824 19321 44990 19322
tri 44990 19321 44991 19322 sw
tri 45282 19321 45283 19322 ne
rect 45283 19321 71000 19322
rect 41824 19029 44991 19321
tri 44991 19029 45283 19321 sw
tri 45283 19029 45575 19321 ne
rect 45575 19029 71000 19321
rect 41824 19028 45283 19029
tri 45283 19028 45284 19029 sw
tri 45575 19028 45576 19029 ne
rect 45576 19028 71000 19029
rect 41824 18736 45284 19028
tri 45284 18736 45576 19028 sw
tri 45576 18736 45868 19028 ne
rect 45868 18736 71000 19028
rect 41824 18735 45576 18736
tri 45576 18735 45577 18736 sw
tri 45868 18735 45869 18736 ne
rect 45869 18735 71000 18736
rect 41824 18443 45577 18735
tri 45577 18443 45869 18735 sw
tri 45869 18443 46161 18735 ne
rect 46161 18443 71000 18735
rect 41824 18244 45869 18443
tri 45869 18244 46068 18443 sw
tri 46161 18244 46360 18443 ne
rect 46360 18244 71000 18443
tri 41824 14000 46068 18244 ne
tri 46068 17952 46360 18244 sw
tri 46360 17952 46652 18244 ne
rect 46652 17952 71000 18244
rect 46068 17880 46360 17952
tri 46360 17880 46432 17952 sw
tri 46652 17880 46724 17952 ne
rect 46724 17880 71000 17952
rect 46068 17588 46432 17880
tri 46432 17588 46724 17880 sw
tri 46724 17588 47016 17880 ne
rect 47016 17588 71000 17880
rect 46068 17587 46724 17588
tri 46724 17587 46725 17588 sw
tri 47016 17587 47017 17588 ne
rect 47017 17587 71000 17588
rect 46068 17295 46725 17587
tri 46725 17295 47017 17587 sw
tri 47017 17295 47309 17587 ne
rect 47309 17295 71000 17587
rect 46068 17294 47017 17295
tri 47017 17294 47018 17295 sw
tri 47309 17294 47310 17295 ne
rect 47310 17294 71000 17295
rect 46068 17002 47018 17294
tri 47018 17002 47310 17294 sw
tri 47310 17200 47404 17294 ne
rect 47404 17200 71000 17294
rect 46068 17000 47310 17002
tri 47310 17000 47312 17002 sw
rect 46068 14000 71000 17000
use M4_M3_CDNS_69033583165207  M4_M3_CDNS_69033583165207_0
timestamp 1713338890
transform 1 0 14032 0 1 47127
box 28 -38 3008 38
use M4_M3_CDNS_69033583165207  M4_M3_CDNS_69033583165207_1
timestamp 1713338890
transform 1 0 17232 0 1 48463
box 28 -38 3008 38
use M4_M3_CDNS_69033583165207  M4_M3_CDNS_69033583165207_2
timestamp 1713338890
transform 1 0 20432 0 1 49789
box 28 -38 3008 38
use M4_M3_CDNS_69033583165207  M4_M3_CDNS_69033583165207_3
timestamp 1713338890
transform 1 0 26832 0 1 52469
box 28 -38 3008 38
use M4_M3_CDNS_69033583165207  M4_M3_CDNS_69033583165207_4
timestamp 1713338890
transform 1 0 30032 0 1 53807
box 28 -38 3008 38
use M4_M3_CDNS_69033583165207  M4_M3_CDNS_69033583165207_5
timestamp 1713338890
transform 1 0 33232 0 1 55139
box 28 -38 3008 38
use M4_M3_CDNS_69033583165207  M4_M3_CDNS_69033583165207_6
timestamp 1713338890
transform 1 0 36432 0 1 56480
box 28 -38 3008 38
use M4_M3_CDNS_69033583165207  M4_M3_CDNS_69033583165207_7
timestamp 1713338890
transform 1 0 42832 0 1 59156
box 28 -38 3008 38
use M4_M3_CDNS_69033583165207  M4_M3_CDNS_69033583165207_8
timestamp 1713338890
transform 1 0 46032 0 1 60523
box 28 -38 3008 38
use M4_M3_CDNS_69033583165208  M4_M3_CDNS_69033583165208_0
timestamp 1713338890
transform 1 0 34700 0 1 63162
box -1490 -7760 1490 7760
use M4_M3_CDNS_69033583165209  M4_M3_CDNS_69033583165209_0
timestamp 1713338890
transform 1 0 63162 0 1 34700
box -7760 -1490 7760 1490
use M4_M3_CDNS_69033583165210  M4_M3_CDNS_69033583165210_0
timestamp 1713338890
transform 1 0 14032 0 1 46863
box 28 -38 3272 38
use M4_M3_CDNS_69033583165210  M4_M3_CDNS_69033583165210_1
timestamp 1713338890
transform 1 0 17232 0 1 48199
box 28 -38 3272 38
use M4_M3_CDNS_69033583165210  M4_M3_CDNS_69033583165210_2
timestamp 1713338890
transform 1 0 20432 0 1 49525
box 28 -38 3272 38
use M4_M3_CDNS_69033583165210  M4_M3_CDNS_69033583165210_3
timestamp 1713338890
transform 1 0 26832 0 1 52205
box 28 -38 3272 38
use M4_M3_CDNS_69033583165210  M4_M3_CDNS_69033583165210_4
timestamp 1713338890
transform 1 0 30032 0 1 53543
box 28 -38 3272 38
use M4_M3_CDNS_69033583165210  M4_M3_CDNS_69033583165210_5
timestamp 1713338890
transform 1 0 33232 0 1 54875
box 28 -38 3272 38
use M4_M3_CDNS_69033583165210  M4_M3_CDNS_69033583165210_6
timestamp 1713338890
transform 1 0 36432 0 1 56216
box 28 -38 3272 38
use M4_M3_CDNS_69033583165210  M4_M3_CDNS_69033583165210_7
timestamp 1713338890
transform 1 0 42832 0 1 58892
box 28 -38 3272 38
use M4_M3_CDNS_69033583165210  M4_M3_CDNS_69033583165210_8
timestamp 1713338890
transform 1 0 46032 0 1 60259
box 28 -38 3272 38
use M4_M3_CDNS_69033583165211  M4_M3_CDNS_69033583165211_0
timestamp 1713338890
transform 1 0 14032 0 1 46203
box 28 -38 3932 38
use M4_M3_CDNS_69033583165211  M4_M3_CDNS_69033583165211_1
timestamp 1713338890
transform 1 0 17232 0 1 47539
box 28 -38 3932 38
use M4_M3_CDNS_69033583165211  M4_M3_CDNS_69033583165211_2
timestamp 1713338890
transform 1 0 20432 0 1 48865
box 28 -38 3932 38
use M4_M3_CDNS_69033583165211  M4_M3_CDNS_69033583165211_3
timestamp 1713338890
transform 1 0 26832 0 1 51545
box 28 -38 3932 38
use M4_M3_CDNS_69033583165211  M4_M3_CDNS_69033583165211_4
timestamp 1713338890
transform 1 0 30032 0 1 52883
box 28 -38 3932 38
use M4_M3_CDNS_69033583165211  M4_M3_CDNS_69033583165211_5
timestamp 1713338890
transform 1 0 33232 0 1 54215
box 28 -38 3932 38
use M4_M3_CDNS_69033583165211  M4_M3_CDNS_69033583165211_6
timestamp 1713338890
transform 1 0 36432 0 1 55556
box 28 -38 3932 38
use M4_M3_CDNS_69033583165211  M4_M3_CDNS_69033583165211_7
timestamp 1713338890
transform 1 0 42832 0 1 58232
box 28 -38 3932 38
use M4_M3_CDNS_69033583165211  M4_M3_CDNS_69033583165211_8
timestamp 1713338890
transform 1 0 46032 0 1 59599
box 28 -38 3932 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_0
timestamp 1713338890
transform 1 0 49590 0 1 25071
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1
timestamp 1713338890
transform 1 0 49458 0 1 25203
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_2
timestamp 1713338890
transform 1 0 49194 0 1 25467
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_3
timestamp 1713338890
transform 1 0 49326 0 1 25335
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_4
timestamp 1713338890
transform 1 0 49062 0 1 25599
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_5
timestamp 1713338890
transform 1 0 48930 0 1 25731
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_6
timestamp 1713338890
transform 1 0 48798 0 1 25863
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_7
timestamp 1713338890
transform 1 0 48666 0 1 25995
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_8
timestamp 1713338890
transform 1 0 48534 0 1 26127
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_9
timestamp 1713338890
transform 1 0 48402 0 1 26259
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_10
timestamp 1713338890
transform 1 0 48138 0 1 26523
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_11
timestamp 1713338890
transform 1 0 48270 0 1 26391
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_12
timestamp 1713338890
transform 1 0 48006 0 1 26655
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_13
timestamp 1713338890
transform 1 0 50266 0 1 26664
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_14
timestamp 1713338890
transform 1 0 47874 0 1 26787
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_15
timestamp 1713338890
transform 1 0 47742 0 1 26919
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_16
timestamp 1713338890
transform 1 0 50134 0 1 26796
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_17
timestamp 1713338890
transform 1 0 47610 0 1 27051
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_18
timestamp 1713338890
transform 1 0 49870 0 1 27060
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_19
timestamp 1713338890
transform 1 0 50002 0 1 26928
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_20
timestamp 1713338890
transform 1 0 47478 0 1 27183
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_21
timestamp 1713338890
transform 1 0 49738 0 1 27192
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_22
timestamp 1713338890
transform 1 0 49606 0 1 27324
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_23
timestamp 1713338890
transform 1 0 49474 0 1 27456
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_24
timestamp 1713338890
transform 1 0 47346 0 1 27315
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_25
timestamp 1713338890
transform 1 0 47214 0 1 27447
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_26
timestamp 1713338890
transform 1 0 49342 0 1 27588
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_27
timestamp 1713338890
transform 1 0 47082 0 1 27579
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_28
timestamp 1713338890
transform 1 0 49210 0 1 27720
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_29
timestamp 1713338890
transform 1 0 46818 0 1 27843
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_30
timestamp 1713338890
transform 1 0 46950 0 1 27711
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_31
timestamp 1713338890
transform 1 0 49078 0 1 27852
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_32
timestamp 1713338890
transform 1 0 48946 0 1 27984
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_33
timestamp 1713338890
transform 1 0 46686 0 1 27975
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_34
timestamp 1713338890
transform 1 0 48814 0 1 28116
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_35
timestamp 1713338890
transform 1 0 48682 0 1 28248
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_36
timestamp 1713338890
transform 1 0 46554 0 1 28107
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_37
timestamp 1713338890
transform 1 0 46422 0 1 28239
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_38
timestamp 1713338890
transform 1 0 48550 0 1 28380
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_39
timestamp 1713338890
transform 1 0 46290 0 1 28371
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_40
timestamp 1713338890
transform 1 0 48418 0 1 28512
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_41
timestamp 1713338890
transform 1 0 48286 0 1 28644
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_42
timestamp 1713338890
transform 1 0 46026 0 1 28635
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_43
timestamp 1713338890
transform 1 0 46158 0 1 28503
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_44
timestamp 1713338890
transform 1 0 48154 0 1 28776
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_45
timestamp 1713338890
transform 1 0 45894 0 1 28767
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_46
timestamp 1713338890
transform 1 0 45630 0 1 29031
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_47
timestamp 1713338890
transform 1 0 48022 0 1 28908
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_48
timestamp 1713338890
transform 1 0 47890 0 1 29040
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_49
timestamp 1713338890
transform 1 0 45762 0 1 28899
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_50
timestamp 1713338890
transform 1 0 45366 0 1 29295
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_51
timestamp 1713338890
transform 1 0 45498 0 1 29163
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_52
timestamp 1713338890
transform 1 0 47758 0 1 29172
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_53
timestamp 1713338890
transform 1 0 47626 0 1 29304
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_54
timestamp 1713338890
transform 1 0 45234 0 1 29427
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_55
timestamp 1713338890
transform 1 0 47494 0 1 29436
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_56
timestamp 1713338890
transform 1 0 44970 0 1 29691
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_57
timestamp 1713338890
transform 1 0 45102 0 1 29559
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_58
timestamp 1713338890
transform 1 0 47362 0 1 29568
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_59
timestamp 1713338890
transform 1 0 47230 0 1 29700
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_60
timestamp 1713338890
transform 1 0 44838 0 1 29823
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_61
timestamp 1713338890
transform 1 0 47098 0 1 29832
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_62
timestamp 1713338890
transform 1 0 44574 0 1 30087
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_63
timestamp 1713338890
transform 1 0 44706 0 1 29955
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_64
timestamp 1713338890
transform 1 0 46966 0 1 29964
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_65
timestamp 1713338890
transform 1 0 44442 0 1 30219
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_66
timestamp 1713338890
transform 1 0 46702 0 1 30228
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_67
timestamp 1713338890
transform 1 0 46834 0 1 30096
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_68
timestamp 1713338890
transform 1 0 44310 0 1 30351
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_69
timestamp 1713338890
transform 1 0 46570 0 1 30360
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_70
timestamp 1713338890
transform 1 0 44178 0 1 30483
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_71
timestamp 1713338890
transform 1 0 44046 0 1 30615
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_72
timestamp 1713338890
transform 1 0 46306 0 1 30624
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_73
timestamp 1713338890
transform 1 0 46438 0 1 30492
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_74
timestamp 1713338890
transform 1 0 43914 0 1 30747
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_75
timestamp 1713338890
transform 1 0 46174 0 1 30756
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_76
timestamp 1713338890
transform 1 0 43782 0 1 30879
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_77
timestamp 1713338890
transform 1 0 43650 0 1 31011
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_78
timestamp 1713338890
transform 1 0 46042 0 1 30888
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_79
timestamp 1713338890
transform 1 0 45910 0 1 31020
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_80
timestamp 1713338890
transform 1 0 43518 0 1 31143
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_81
timestamp 1713338890
transform 1 0 45778 0 1 31152
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_82
timestamp 1713338890
transform 1 0 43386 0 1 31275
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_83
timestamp 1713338890
transform 1 0 45646 0 1 31284
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_84
timestamp 1713338890
transform 1 0 45514 0 1 31416
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_85
timestamp 1713338890
transform 1 0 43254 0 1 31407
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_86
timestamp 1713338890
transform 1 0 45250 0 1 31680
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_87
timestamp 1713338890
transform 1 0 45382 0 1 31548
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_88
timestamp 1713338890
transform 1 0 43122 0 1 31539
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_89
timestamp 1713338890
transform 1 0 42990 0 1 31671
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_90
timestamp 1713338890
transform 1 0 45118 0 1 31812
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_91
timestamp 1713338890
transform 1 0 42858 0 1 31803
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_92
timestamp 1713338890
transform 1 0 44986 0 1 31944
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_93
timestamp 1713338890
transform 1 0 42726 0 1 31935
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_94
timestamp 1713338890
transform 1 0 44854 0 1 32076
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_95
timestamp 1713338890
transform 1 0 42594 0 1 32067
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_96
timestamp 1713338890
transform 1 0 44722 0 1 32208
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_97
timestamp 1713338890
transform 1 0 44590 0 1 32340
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_98
timestamp 1713338890
transform 1 0 42462 0 1 32199
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_99
timestamp 1713338890
transform 1 0 42330 0 1 32331
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_100
timestamp 1713338890
transform 1 0 44458 0 1 32472
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_101
timestamp 1713338890
transform 1 0 42198 0 1 32463
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_102
timestamp 1713338890
transform 1 0 44326 0 1 32604
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_103
timestamp 1713338890
transform 1 0 42066 0 1 32595
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_104
timestamp 1713338890
transform 1 0 44194 0 1 32736
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_105
timestamp 1713338890
transform 1 0 44062 0 1 32868
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_106
timestamp 1713338890
transform 1 0 41802 0 1 32859
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_107
timestamp 1713338890
transform 1 0 41934 0 1 32727
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_108
timestamp 1713338890
transform 1 0 43930 0 1 33000
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_109
timestamp 1713338890
transform 1 0 41670 0 1 32991
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_110
timestamp 1713338890
transform 1 0 41406 0 1 33255
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_111
timestamp 1713338890
transform 1 0 41538 0 1 33123
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_112
timestamp 1713338890
transform 1 0 43798 0 1 33132
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_113
timestamp 1713338890
transform 1 0 41274 0 1 33387
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_114
timestamp 1713338890
transform 1 0 43534 0 1 33396
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_115
timestamp 1713338890
transform 1 0 43666 0 1 33264
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_116
timestamp 1713338890
transform 1 0 41142 0 1 33519
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_117
timestamp 1713338890
transform 1 0 43402 0 1 33528
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_118
timestamp 1713338890
transform 1 0 40878 0 1 33783
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_119
timestamp 1713338890
transform 1 0 41010 0 1 33651
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_120
timestamp 1713338890
transform 1 0 43270 0 1 33660
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_121
timestamp 1713338890
transform 1 0 43138 0 1 33792
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_122
timestamp 1713338890
transform 1 0 40746 0 1 33915
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_123
timestamp 1713338890
transform 1 0 43006 0 1 33924
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_124
timestamp 1713338890
transform 1 0 40614 0 1 34047
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_125
timestamp 1713338890
transform 1 0 42874 0 1 34056
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_126
timestamp 1713338890
transform 1 0 40350 0 1 34311
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_127
timestamp 1713338890
transform 1 0 40482 0 1 34179
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_128
timestamp 1713338890
transform 1 0 42742 0 1 34188
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_129
timestamp 1713338890
transform 1 0 42610 0 1 34320
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_130
timestamp 1713338890
transform 1 0 40218 0 1 34443
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_131
timestamp 1713338890
transform 1 0 42478 0 1 34452
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_132
timestamp 1713338890
transform 1 0 40086 0 1 34575
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_133
timestamp 1713338890
transform 1 0 42346 0 1 34584
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_134
timestamp 1713338890
transform 1 0 39954 0 1 34707
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_135
timestamp 1713338890
transform 1 0 42214 0 1 34716
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_136
timestamp 1713338890
transform 1 0 39822 0 1 34839
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_137
timestamp 1713338890
transform 1 0 39690 0 1 34971
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_138
timestamp 1713338890
transform 1 0 42082 0 1 34848
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_139
timestamp 1713338890
transform 1 0 41950 0 1 34980
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_140
timestamp 1713338890
transform 1 0 39558 0 1 35103
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_141
timestamp 1713338890
transform 1 0 41818 0 1 35112
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_142
timestamp 1713338890
transform 1 0 39426 0 1 35235
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_143
timestamp 1713338890
transform 1 0 41686 0 1 35244
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_144
timestamp 1713338890
transform 1 0 39294 0 1 35367
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_145
timestamp 1713338890
transform 1 0 41554 0 1 35376
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_146
timestamp 1713338890
transform 1 0 39162 0 1 35499
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_147
timestamp 1713338890
transform 1 0 41422 0 1 35508
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_148
timestamp 1713338890
transform 1 0 39030 0 1 35631
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_149
timestamp 1713338890
transform 1 0 41290 0 1 35640
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_150
timestamp 1713338890
transform 1 0 38898 0 1 35763
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_151
timestamp 1713338890
transform 1 0 41158 0 1 35772
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_152
timestamp 1713338890
transform 1 0 38766 0 1 35895
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_153
timestamp 1713338890
transform 1 0 41026 0 1 35904
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_154
timestamp 1713338890
transform 1 0 38634 0 1 36027
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_155
timestamp 1713338890
transform 1 0 40894 0 1 36036
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_156
timestamp 1713338890
transform 1 0 40762 0 1 36168
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_157
timestamp 1713338890
transform 1 0 38502 0 1 36159
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_158
timestamp 1713338890
transform 1 0 40630 0 1 36300
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_159
timestamp 1713338890
transform 1 0 38370 0 1 36291
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_160
timestamp 1713338890
transform 1 0 40498 0 1 36432
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_161
timestamp 1713338890
transform 1 0 38238 0 1 36423
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_162
timestamp 1713338890
transform 1 0 40366 0 1 36564
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_163
timestamp 1713338890
transform 1 0 38106 0 1 36555
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_164
timestamp 1713338890
transform 1 0 40102 0 1 36828
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_165
timestamp 1713338890
transform 1 0 40234 0 1 36696
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_166
timestamp 1713338890
transform 1 0 37842 0 1 36819
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_167
timestamp 1713338890
transform 1 0 37974 0 1 36687
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_168
timestamp 1713338890
transform 1 0 39970 0 1 36960
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_169
timestamp 1713338890
transform 1 0 37710 0 1 36951
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_170
timestamp 1713338890
transform 1 0 37314 0 1 37347
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_171
timestamp 1713338890
transform 1 0 37446 0 1 37215
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_172
timestamp 1713338890
transform 1 0 37182 0 1 37479
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_173
timestamp 1713338890
transform 1 0 36918 0 1 37743
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_174
timestamp 1713338890
transform 1 0 37050 0 1 37611
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_175
timestamp 1713338890
transform 1 0 36786 0 1 37875
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_176
timestamp 1713338890
transform 1 0 36522 0 1 38139
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_177
timestamp 1713338890
transform 1 0 36654 0 1 38007
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_178
timestamp 1713338890
transform 1 0 36390 0 1 38271
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_179
timestamp 1713338890
transform 1 0 36126 0 1 38535
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_180
timestamp 1713338890
transform 1 0 36258 0 1 38403
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_181
timestamp 1713338890
transform 1 0 35994 0 1 38667
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_182
timestamp 1713338890
transform 1 0 35730 0 1 38931
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_183
timestamp 1713338890
transform 1 0 35862 0 1 38799
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_184
timestamp 1713338890
transform 1 0 35598 0 1 39063
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_185
timestamp 1713338890
transform 1 0 35466 0 1 39195
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_186
timestamp 1713338890
transform 1 0 35334 0 1 39327
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_187
timestamp 1713338890
transform 1 0 35202 0 1 39459
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_188
timestamp 1713338890
transform 1 0 37462 0 1 39468
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_189
timestamp 1713338890
transform 1 0 35070 0 1 39591
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_190
timestamp 1713338890
transform 1 0 34938 0 1 39723
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_191
timestamp 1713338890
transform 1 0 37330 0 1 39600
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_192
timestamp 1713338890
transform 1 0 37198 0 1 39732
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_193
timestamp 1713338890
transform 1 0 34806 0 1 39855
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_194
timestamp 1713338890
transform 1 0 37066 0 1 39864
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_195
timestamp 1713338890
transform 1 0 39838 0 1 37092
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_196
timestamp 1713338890
transform 1 0 37578 0 1 37083
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_197
timestamp 1713338890
transform 1 0 39706 0 1 37224
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_198
timestamp 1713338890
transform 1 0 39442 0 1 37488
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_199
timestamp 1713338890
transform 1 0 39574 0 1 37356
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_200
timestamp 1713338890
transform 1 0 39310 0 1 37620
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_201
timestamp 1713338890
transform 1 0 39178 0 1 37752
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_202
timestamp 1713338890
transform 1 0 38914 0 1 38016
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_203
timestamp 1713338890
transform 1 0 39046 0 1 37884
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_204
timestamp 1713338890
transform 1 0 38782 0 1 38148
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_205
timestamp 1713338890
transform 1 0 38650 0 1 38280
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_206
timestamp 1713338890
transform 1 0 38386 0 1 38544
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_207
timestamp 1713338890
transform 1 0 38518 0 1 38412
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_208
timestamp 1713338890
transform 1 0 38254 0 1 38676
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_209
timestamp 1713338890
transform 1 0 38122 0 1 38808
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_210
timestamp 1713338890
transform 1 0 37990 0 1 38940
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_211
timestamp 1713338890
transform 1 0 37858 0 1 39072
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_212
timestamp 1713338890
transform 1 0 37726 0 1 39204
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_213
timestamp 1713338890
transform 1 0 37594 0 1 39336
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_214
timestamp 1713338890
transform 1 0 34674 0 1 39987
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_215
timestamp 1713338890
transform 1 0 36802 0 1 40128
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_216
timestamp 1713338890
transform 1 0 36934 0 1 39996
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_217
timestamp 1713338890
transform 1 0 34542 0 1 40119
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_218
timestamp 1713338890
transform 1 0 36670 0 1 40260
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_219
timestamp 1713338890
transform 1 0 34278 0 1 40383
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_220
timestamp 1713338890
transform 1 0 34410 0 1 40251
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_221
timestamp 1713338890
transform 1 0 34146 0 1 40515
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_222
timestamp 1713338890
transform 1 0 36406 0 1 40524
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_223
timestamp 1713338890
transform 1 0 36538 0 1 40392
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_224
timestamp 1713338890
transform 1 0 34014 0 1 40647
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_225
timestamp 1713338890
transform 1 0 33882 0 1 40779
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_226
timestamp 1713338890
transform 1 0 36142 0 1 40788
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_227
timestamp 1713338890
transform 1 0 36274 0 1 40656
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_228
timestamp 1713338890
transform 1 0 33750 0 1 40911
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_229
timestamp 1713338890
transform 1 0 36010 0 1 40920
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_230
timestamp 1713338890
transform 1 0 33618 0 1 41043
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_231
timestamp 1713338890
transform 1 0 33486 0 1 41175
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_232
timestamp 1713338890
transform 1 0 35746 0 1 41184
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_233
timestamp 1713338890
transform 1 0 35878 0 1 41052
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_234
timestamp 1713338890
transform 1 0 33222 0 1 41439
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_235
timestamp 1713338890
transform 1 0 33354 0 1 41307
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_236
timestamp 1713338890
transform 1 0 35482 0 1 41448
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_237
timestamp 1713338890
transform 1 0 35614 0 1 41316
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_238
timestamp 1713338890
transform 1 0 33090 0 1 41571
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_239
timestamp 1713338890
transform 1 0 35350 0 1 41580
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_240
timestamp 1713338890
transform 1 0 32958 0 1 41703
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_241
timestamp 1713338890
transform 1 0 32826 0 1 41835
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_242
timestamp 1713338890
transform 1 0 35086 0 1 41844
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_243
timestamp 1713338890
transform 1 0 35218 0 1 41712
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_244
timestamp 1713338890
transform 1 0 32694 0 1 41967
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_245
timestamp 1713338890
transform 1 0 34954 0 1 41976
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_246
timestamp 1713338890
transform 1 0 56218 0 1 41130
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_247
timestamp 1713338890
transform 1 0 56086 0 1 41262
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_248
timestamp 1713338890
transform 1 0 55690 0 1 41658
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_249
timestamp 1713338890
transform 1 0 55822 0 1 41526
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_250
timestamp 1713338890
transform 1 0 55954 0 1 41394
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_251
timestamp 1713338890
transform 1 0 55294 0 1 42054
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_252
timestamp 1713338890
transform 1 0 55426 0 1 41922
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_253
timestamp 1713338890
transform 1 0 55558 0 1 41790
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_254
timestamp 1713338890
transform 1 0 25434 0 1 49227
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_255
timestamp 1713338890
transform 1 0 25302 0 1 49359
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_256
timestamp 1713338890
transform 1 0 25038 0 1 49623
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_257
timestamp 1713338890
transform 1 0 24906 0 1 49755
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_258
timestamp 1713338890
transform 1 0 25170 0 1 49491
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_259
timestamp 1713338890
transform 1 0 24642 0 1 50019
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_260
timestamp 1713338890
transform 1 0 24774 0 1 49887
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_261
timestamp 1713338890
transform 1 0 29526 0 1 45135
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_262
timestamp 1713338890
transform 1 0 29394 0 1 45267
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_263
timestamp 1713338890
transform 1 0 29262 0 1 45399
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_264
timestamp 1713338890
transform 1 0 29130 0 1 45531
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_265
timestamp 1713338890
transform 1 0 28998 0 1 45663
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_266
timestamp 1713338890
transform 1 0 28866 0 1 45795
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_267
timestamp 1713338890
transform 1 0 28734 0 1 45927
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_268
timestamp 1713338890
transform 1 0 28602 0 1 46059
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_269
timestamp 1713338890
transform 1 0 28470 0 1 46191
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_270
timestamp 1713338890
transform 1 0 28206 0 1 46455
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_271
timestamp 1713338890
transform 1 0 28338 0 1 46323
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_272
timestamp 1713338890
transform 1 0 28074 0 1 46587
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_273
timestamp 1713338890
transform 1 0 27942 0 1 46719
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_274
timestamp 1713338890
transform 1 0 27810 0 1 46851
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_275
timestamp 1713338890
transform 1 0 27678 0 1 46983
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_276
timestamp 1713338890
transform 1 0 27546 0 1 47115
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_277
timestamp 1713338890
transform 1 0 27414 0 1 47247
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_278
timestamp 1713338890
transform 1 0 27282 0 1 47379
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_279
timestamp 1713338890
transform 1 0 29542 0 1 47388
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_280
timestamp 1713338890
transform 1 0 27150 0 1 47511
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_281
timestamp 1713338890
transform 1 0 29410 0 1 47520
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_282
timestamp 1713338890
transform 1 0 27018 0 1 47643
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_283
timestamp 1713338890
transform 1 0 29278 0 1 47652
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_284
timestamp 1713338890
transform 1 0 26886 0 1 47775
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_285
timestamp 1713338890
transform 1 0 29146 0 1 47784
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_286
timestamp 1713338890
transform 1 0 26754 0 1 47907
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_287
timestamp 1713338890
transform 1 0 29014 0 1 47916
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_288
timestamp 1713338890
transform 1 0 26622 0 1 48039
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_289
timestamp 1713338890
transform 1 0 28882 0 1 48048
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_290
timestamp 1713338890
transform 1 0 26490 0 1 48171
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_291
timestamp 1713338890
transform 1 0 28750 0 1 48180
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_292
timestamp 1713338890
transform 1 0 26358 0 1 48303
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_293
timestamp 1713338890
transform 1 0 28618 0 1 48312
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_294
timestamp 1713338890
transform 1 0 26226 0 1 48435
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_295
timestamp 1713338890
transform 1 0 26094 0 1 48567
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_296
timestamp 1713338890
transform 1 0 28486 0 1 48444
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_297
timestamp 1713338890
transform 1 0 25962 0 1 48699
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_298
timestamp 1713338890
transform 1 0 28222 0 1 48708
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_299
timestamp 1713338890
transform 1 0 28354 0 1 48576
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_300
timestamp 1713338890
transform 1 0 25830 0 1 48831
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_301
timestamp 1713338890
transform 1 0 28090 0 1 48840
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_302
timestamp 1713338890
transform 1 0 27958 0 1 48972
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_303
timestamp 1713338890
transform 1 0 25698 0 1 48963
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_304
timestamp 1713338890
transform 1 0 27826 0 1 49104
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_305
timestamp 1713338890
transform 1 0 25566 0 1 49095
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_306
timestamp 1713338890
transform 1 0 27694 0 1 49236
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_307
timestamp 1713338890
transform 1 0 27562 0 1 49368
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_308
timestamp 1713338890
transform 1 0 27430 0 1 49500
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_309
timestamp 1713338890
transform 1 0 27298 0 1 49632
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_310
timestamp 1713338890
transform 1 0 27166 0 1 49764
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_311
timestamp 1713338890
transform 1 0 27034 0 1 49896
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_312
timestamp 1713338890
transform 1 0 26902 0 1 50028
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_313
timestamp 1713338890
transform 1 0 26770 0 1 50160
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_314
timestamp 1713338890
transform 1 0 26638 0 1 50292
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_315
timestamp 1713338890
transform 1 0 26506 0 1 50424
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_316
timestamp 1713338890
transform 1 0 26374 0 1 50556
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_317
timestamp 1713338890
transform 1 0 26242 0 1 50688
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_318
timestamp 1713338890
transform 1 0 32562 0 1 42099
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_319
timestamp 1713338890
transform 1 0 32430 0 1 42231
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_320
timestamp 1713338890
transform 1 0 32298 0 1 42363
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_321
timestamp 1713338890
transform 1 0 32166 0 1 42495
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_322
timestamp 1713338890
transform 1 0 32034 0 1 42627
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_323
timestamp 1713338890
transform 1 0 31902 0 1 42759
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_324
timestamp 1713338890
transform 1 0 31770 0 1 42891
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_325
timestamp 1713338890
transform 1 0 31638 0 1 43023
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_326
timestamp 1713338890
transform 1 0 31506 0 1 43155
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_327
timestamp 1713338890
transform 1 0 31374 0 1 43287
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_328
timestamp 1713338890
transform 1 0 31242 0 1 43419
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_329
timestamp 1713338890
transform 1 0 33502 0 1 43428
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_330
timestamp 1713338890
transform 1 0 31110 0 1 43551
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_331
timestamp 1713338890
transform 1 0 33370 0 1 43560
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_332
timestamp 1713338890
transform 1 0 30978 0 1 43683
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_333
timestamp 1713338890
transform 1 0 33238 0 1 43692
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_334
timestamp 1713338890
transform 1 0 30846 0 1 43815
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_335
timestamp 1713338890
transform 1 0 33106 0 1 43824
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_336
timestamp 1713338890
transform 1 0 30714 0 1 43947
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_337
timestamp 1713338890
transform 1 0 32974 0 1 43956
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_338
timestamp 1713338890
transform 1 0 30582 0 1 44079
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_339
timestamp 1713338890
transform 1 0 32842 0 1 44088
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_340
timestamp 1713338890
transform 1 0 30450 0 1 44211
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_341
timestamp 1713338890
transform 1 0 32710 0 1 44220
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_342
timestamp 1713338890
transform 1 0 30318 0 1 44343
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_343
timestamp 1713338890
transform 1 0 32578 0 1 44352
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_344
timestamp 1713338890
transform 1 0 30186 0 1 44475
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_345
timestamp 1713338890
transform 1 0 32446 0 1 44484
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_346
timestamp 1713338890
transform 1 0 30054 0 1 44607
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_347
timestamp 1713338890
transform 1 0 32314 0 1 44616
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_348
timestamp 1713338890
transform 1 0 29922 0 1 44739
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_349
timestamp 1713338890
transform 1 0 32182 0 1 44748
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_350
timestamp 1713338890
transform 1 0 29790 0 1 44871
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_351
timestamp 1713338890
transform 1 0 32050 0 1 44880
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_352
timestamp 1713338890
transform 1 0 31918 0 1 45012
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_353
timestamp 1713338890
transform 1 0 29658 0 1 45003
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_354
timestamp 1713338890
transform 1 0 31786 0 1 45144
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_355
timestamp 1713338890
transform 1 0 31654 0 1 45276
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_356
timestamp 1713338890
transform 1 0 31522 0 1 45408
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_357
timestamp 1713338890
transform 1 0 31390 0 1 45540
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_358
timestamp 1713338890
transform 1 0 31258 0 1 45672
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_359
timestamp 1713338890
transform 1 0 31126 0 1 45804
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_360
timestamp 1713338890
transform 1 0 30994 0 1 45936
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_361
timestamp 1713338890
transform 1 0 30862 0 1 46068
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_362
timestamp 1713338890
transform 1 0 30730 0 1 46200
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_363
timestamp 1713338890
transform 1 0 30598 0 1 46332
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_364
timestamp 1713338890
transform 1 0 30466 0 1 46464
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_365
timestamp 1713338890
transform 1 0 30334 0 1 46596
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_366
timestamp 1713338890
transform 1 0 30202 0 1 46728
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_367
timestamp 1713338890
transform 1 0 30070 0 1 46860
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_368
timestamp 1713338890
transform 1 0 29938 0 1 46992
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_369
timestamp 1713338890
transform 1 0 29806 0 1 47124
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_370
timestamp 1713338890
transform 1 0 29674 0 1 47256
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_371
timestamp 1713338890
transform 1 0 34690 0 1 42240
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_372
timestamp 1713338890
transform 1 0 34822 0 1 42108
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_373
timestamp 1713338890
transform 1 0 34558 0 1 42372
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_374
timestamp 1713338890
transform 1 0 34426 0 1 42504
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_375
timestamp 1713338890
transform 1 0 34294 0 1 42636
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_376
timestamp 1713338890
transform 1 0 34162 0 1 42768
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_377
timestamp 1713338890
transform 1 0 34030 0 1 42900
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_378
timestamp 1713338890
transform 1 0 33898 0 1 43032
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_379
timestamp 1713338890
transform 1 0 33766 0 1 43164
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_380
timestamp 1713338890
transform 1 0 33634 0 1 43296
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_381
timestamp 1713338890
transform 1 0 45130 0 1 52218
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_382
timestamp 1713338890
transform 1 0 44998 0 1 52350
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_383
timestamp 1713338890
transform 1 0 44866 0 1 52482
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_384
timestamp 1713338890
transform 1 0 44734 0 1 52614
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_385
timestamp 1713338890
transform 1 0 44602 0 1 52746
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_386
timestamp 1713338890
transform 1 0 44470 0 1 52878
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_387
timestamp 1713338890
transform 1 0 44338 0 1 53010
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_388
timestamp 1713338890
transform 1 0 44206 0 1 53142
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_389
timestamp 1713338890
transform 1 0 44074 0 1 53274
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_390
timestamp 1713338890
transform 1 0 43942 0 1 53406
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_391
timestamp 1713338890
transform 1 0 43810 0 1 53538
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_392
timestamp 1713338890
transform 1 0 43678 0 1 53670
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_393
timestamp 1713338890
transform 1 0 43546 0 1 53802
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_394
timestamp 1713338890
transform 1 0 43414 0 1 53934
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_395
timestamp 1713338890
transform 1 0 43282 0 1 54066
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_396
timestamp 1713338890
transform 1 0 43150 0 1 54198
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_397
timestamp 1713338890
transform 1 0 43018 0 1 54330
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_398
timestamp 1713338890
transform 1 0 45146 0 1 54474
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_399
timestamp 1713338890
transform 1 0 42886 0 1 54462
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_400
timestamp 1713338890
transform 1 0 45014 0 1 54606
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_401
timestamp 1713338890
transform 1 0 42754 0 1 54594
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_402
timestamp 1713338890
transform 1 0 44882 0 1 54738
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_403
timestamp 1713338890
transform 1 0 42622 0 1 54726
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_404
timestamp 1713338890
transform 1 0 44750 0 1 54870
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_405
timestamp 1713338890
transform 1 0 42490 0 1 54858
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_406
timestamp 1713338890
transform 1 0 44618 0 1 55002
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_407
timestamp 1713338890
transform 1 0 42358 0 1 54990
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_408
timestamp 1713338890
transform 1 0 44486 0 1 55134
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_409
timestamp 1713338890
transform 1 0 42226 0 1 55122
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_410
timestamp 1713338890
transform 1 0 44354 0 1 55266
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_411
timestamp 1713338890
transform 1 0 42094 0 1 55254
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_412
timestamp 1713338890
transform 1 0 44222 0 1 55398
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_413
timestamp 1713338890
transform 1 0 41962 0 1 55386
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_414
timestamp 1713338890
transform 1 0 44090 0 1 55530
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_415
timestamp 1713338890
transform 1 0 41830 0 1 55518
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_416
timestamp 1713338890
transform 1 0 43958 0 1 55662
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_417
timestamp 1713338890
transform 1 0 41698 0 1 55650
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_418
timestamp 1713338890
transform 1 0 43826 0 1 55794
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_419
timestamp 1713338890
transform 1 0 41566 0 1 55782
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_420
timestamp 1713338890
transform 1 0 43694 0 1 55926
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_421
timestamp 1713338890
transform 1 0 41434 0 1 55914
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_422
timestamp 1713338890
transform 1 0 43562 0 1 56058
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_423
timestamp 1713338890
transform 1 0 41302 0 1 56046
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_424
timestamp 1713338890
transform 1 0 41170 0 1 56178
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_425
timestamp 1713338890
transform 1 0 43430 0 1 56190
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_426
timestamp 1713338890
transform 1 0 48562 0 1 48786
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_427
timestamp 1713338890
transform 1 0 48430 0 1 48918
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_428
timestamp 1713338890
transform 1 0 48298 0 1 49050
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_429
timestamp 1713338890
transform 1 0 48166 0 1 49182
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_430
timestamp 1713338890
transform 1 0 48034 0 1 49314
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_431
timestamp 1713338890
transform 1 0 47902 0 1 49446
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_432
timestamp 1713338890
transform 1 0 47770 0 1 49578
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_433
timestamp 1713338890
transform 1 0 47638 0 1 49710
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_434
timestamp 1713338890
transform 1 0 47506 0 1 49842
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_435
timestamp 1713338890
transform 1 0 47374 0 1 49974
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_436
timestamp 1713338890
transform 1 0 47242 0 1 50106
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_437
timestamp 1713338890
transform 1 0 47110 0 1 50238
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_438
timestamp 1713338890
transform 1 0 46978 0 1 50370
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_439
timestamp 1713338890
transform 1 0 46846 0 1 50502
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_440
timestamp 1713338890
transform 1 0 46714 0 1 50634
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_441
timestamp 1713338890
transform 1 0 46582 0 1 50766
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_442
timestamp 1713338890
transform 1 0 46450 0 1 50898
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_443
timestamp 1713338890
transform 1 0 48578 0 1 51042
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_444
timestamp 1713338890
transform 1 0 46318 0 1 51030
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_445
timestamp 1713338890
transform 1 0 48446 0 1 51174
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_446
timestamp 1713338890
transform 1 0 46186 0 1 51162
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_447
timestamp 1713338890
transform 1 0 48314 0 1 51306
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_448
timestamp 1713338890
transform 1 0 46054 0 1 51294
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_449
timestamp 1713338890
transform 1 0 48182 0 1 51438
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_450
timestamp 1713338890
transform 1 0 45922 0 1 51426
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_451
timestamp 1713338890
transform 1 0 48050 0 1 51570
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_452
timestamp 1713338890
transform 1 0 45790 0 1 51558
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_453
timestamp 1713338890
transform 1 0 45658 0 1 51690
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_454
timestamp 1713338890
transform 1 0 47918 0 1 51702
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_455
timestamp 1713338890
transform 1 0 45526 0 1 51822
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_456
timestamp 1713338890
transform 1 0 47786 0 1 51834
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_457
timestamp 1713338890
transform 1 0 45394 0 1 51954
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_458
timestamp 1713338890
transform 1 0 47654 0 1 51966
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_459
timestamp 1713338890
transform 1 0 45262 0 1 52086
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_460
timestamp 1713338890
transform 1 0 47522 0 1 52098
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_461
timestamp 1713338890
transform 1 0 47390 0 1 52230
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_462
timestamp 1713338890
transform 1 0 47258 0 1 52362
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_463
timestamp 1713338890
transform 1 0 47126 0 1 52494
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_464
timestamp 1713338890
transform 1 0 46994 0 1 52626
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_465
timestamp 1713338890
transform 1 0 46862 0 1 52758
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_466
timestamp 1713338890
transform 1 0 46730 0 1 52890
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_467
timestamp 1713338890
transform 1 0 46598 0 1 53022
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_468
timestamp 1713338890
transform 1 0 46466 0 1 53154
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_469
timestamp 1713338890
transform 1 0 46334 0 1 53286
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_470
timestamp 1713338890
transform 1 0 46202 0 1 53418
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_471
timestamp 1713338890
transform 1 0 46070 0 1 53550
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_472
timestamp 1713338890
transform 1 0 45938 0 1 53682
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_473
timestamp 1713338890
transform 1 0 45806 0 1 53814
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_474
timestamp 1713338890
transform 1 0 45674 0 1 53946
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_475
timestamp 1713338890
transform 1 0 45542 0 1 54078
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_476
timestamp 1713338890
transform 1 0 45410 0 1 54210
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_477
timestamp 1713338890
transform 1 0 45278 0 1 54342
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_478
timestamp 1713338890
transform 1 0 41038 0 1 56310
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_479
timestamp 1713338890
transform 1 0 40906 0 1 56442
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_480
timestamp 1713338890
transform 1 0 40774 0 1 56574
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_481
timestamp 1713338890
transform 1 0 40642 0 1 56706
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_482
timestamp 1713338890
transform 1 0 43298 0 1 56322
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_483
timestamp 1713338890
transform 1 0 43166 0 1 56454
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_484
timestamp 1713338890
transform 1 0 43034 0 1 56586
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_485
timestamp 1713338890
transform 1 0 42902 0 1 56718
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_486
timestamp 1713338890
transform 1 0 42770 0 1 56850
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_487
timestamp 1713338890
transform 1 0 42506 0 1 57114
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_488
timestamp 1713338890
transform 1 0 42638 0 1 56982
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_489
timestamp 1713338890
transform 1 0 42374 0 1 57246
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_490
timestamp 1713338890
transform 1 0 42242 0 1 57378
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_491
timestamp 1713338890
transform 1 0 52654 0 1 44694
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_492
timestamp 1713338890
transform 1 0 52522 0 1 44826
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_493
timestamp 1713338890
transform 1 0 52390 0 1 44958
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_494
timestamp 1713338890
transform 1 0 52258 0 1 45090
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_495
timestamp 1713338890
transform 1 0 52126 0 1 45222
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_496
timestamp 1713338890
transform 1 0 51994 0 1 45354
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_497
timestamp 1713338890
transform 1 0 51862 0 1 45486
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_498
timestamp 1713338890
transform 1 0 51730 0 1 45618
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_499
timestamp 1713338890
transform 1 0 51598 0 1 45750
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_500
timestamp 1713338890
transform 1 0 51466 0 1 45882
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_501
timestamp 1713338890
transform 1 0 51334 0 1 46014
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_502
timestamp 1713338890
transform 1 0 51202 0 1 46146
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_503
timestamp 1713338890
transform 1 0 51070 0 1 46278
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_504
timestamp 1713338890
transform 1 0 50938 0 1 46410
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_505
timestamp 1713338890
transform 1 0 50806 0 1 46542
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_506
timestamp 1713338890
transform 1 0 50674 0 1 46674
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_507
timestamp 1713338890
transform 1 0 50542 0 1 46806
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_508
timestamp 1713338890
transform 1 0 52670 0 1 46950
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_509
timestamp 1713338890
transform 1 0 50410 0 1 46938
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_510
timestamp 1713338890
transform 1 0 52538 0 1 47082
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_511
timestamp 1713338890
transform 1 0 50278 0 1 47070
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_512
timestamp 1713338890
transform 1 0 52406 0 1 47214
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_513
timestamp 1713338890
transform 1 0 50146 0 1 47202
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_514
timestamp 1713338890
transform 1 0 50014 0 1 47334
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_515
timestamp 1713338890
transform 1 0 52274 0 1 47346
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_516
timestamp 1713338890
transform 1 0 52142 0 1 47478
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_517
timestamp 1713338890
transform 1 0 49882 0 1 47466
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_518
timestamp 1713338890
transform 1 0 52010 0 1 47610
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_519
timestamp 1713338890
transform 1 0 49750 0 1 47598
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_520
timestamp 1713338890
transform 1 0 49618 0 1 47730
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_521
timestamp 1713338890
transform 1 0 51878 0 1 47742
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_522
timestamp 1713338890
transform 1 0 49486 0 1 47862
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_523
timestamp 1713338890
transform 1 0 51746 0 1 47874
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_524
timestamp 1713338890
transform 1 0 49354 0 1 47994
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_525
timestamp 1713338890
transform 1 0 51614 0 1 48006
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_526
timestamp 1713338890
transform 1 0 49222 0 1 48126
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_527
timestamp 1713338890
transform 1 0 51482 0 1 48138
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_528
timestamp 1713338890
transform 1 0 49090 0 1 48258
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_529
timestamp 1713338890
transform 1 0 51350 0 1 48270
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_530
timestamp 1713338890
transform 1 0 48958 0 1 48390
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_531
timestamp 1713338890
transform 1 0 51218 0 1 48402
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_532
timestamp 1713338890
transform 1 0 48826 0 1 48522
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_533
timestamp 1713338890
transform 1 0 51086 0 1 48534
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_534
timestamp 1713338890
transform 1 0 48694 0 1 48654
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_535
timestamp 1713338890
transform 1 0 50954 0 1 48666
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_536
timestamp 1713338890
transform 1 0 50822 0 1 48798
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_537
timestamp 1713338890
transform 1 0 50690 0 1 48930
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_538
timestamp 1713338890
transform 1 0 50558 0 1 49062
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_539
timestamp 1713338890
transform 1 0 50426 0 1 49194
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_540
timestamp 1713338890
transform 1 0 50294 0 1 49326
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_541
timestamp 1713338890
transform 1 0 50162 0 1 49458
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_542
timestamp 1713338890
transform 1 0 50030 0 1 49590
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_543
timestamp 1713338890
transform 1 0 49898 0 1 49722
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_544
timestamp 1713338890
transform 1 0 49766 0 1 49854
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_545
timestamp 1713338890
transform 1 0 49634 0 1 49986
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_546
timestamp 1713338890
transform 1 0 49502 0 1 50118
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_547
timestamp 1713338890
transform 1 0 49370 0 1 50250
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_548
timestamp 1713338890
transform 1 0 49238 0 1 50382
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_549
timestamp 1713338890
transform 1 0 49106 0 1 50514
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_550
timestamp 1713338890
transform 1 0 48974 0 1 50646
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_551
timestamp 1713338890
transform 1 0 48842 0 1 50778
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_552
timestamp 1713338890
transform 1 0 48710 0 1 50910
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_553
timestamp 1713338890
transform 1 0 55162 0 1 42186
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_554
timestamp 1713338890
transform 1 0 55030 0 1 42318
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_555
timestamp 1713338890
transform 1 0 54898 0 1 42450
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_556
timestamp 1713338890
transform 1 0 54766 0 1 42582
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_557
timestamp 1713338890
transform 1 0 54634 0 1 42714
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_558
timestamp 1713338890
transform 1 0 54502 0 1 42846
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_559
timestamp 1713338890
transform 1 0 56630 0 1 42990
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_560
timestamp 1713338890
transform 1 0 54370 0 1 42978
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_561
timestamp 1713338890
transform 1 0 56498 0 1 43122
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_562
timestamp 1713338890
transform 1 0 54238 0 1 43110
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_563
timestamp 1713338890
transform 1 0 54106 0 1 43242
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_564
timestamp 1713338890
transform 1 0 56366 0 1 43254
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_565
timestamp 1713338890
transform 1 0 53974 0 1 43374
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_566
timestamp 1713338890
transform 1 0 56234 0 1 43386
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_567
timestamp 1713338890
transform 1 0 53842 0 1 43506
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_568
timestamp 1713338890
transform 1 0 56102 0 1 43518
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_569
timestamp 1713338890
transform 1 0 53710 0 1 43638
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_570
timestamp 1713338890
transform 1 0 55970 0 1 43650
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_571
timestamp 1713338890
transform 1 0 53578 0 1 43770
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_572
timestamp 1713338890
transform 1 0 55838 0 1 43782
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_573
timestamp 1713338890
transform 1 0 53446 0 1 43902
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_574
timestamp 1713338890
transform 1 0 55706 0 1 43914
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_575
timestamp 1713338890
transform 1 0 53314 0 1 44034
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_576
timestamp 1713338890
transform 1 0 55574 0 1 44046
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_577
timestamp 1713338890
transform 1 0 53182 0 1 44166
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_578
timestamp 1713338890
transform 1 0 55442 0 1 44178
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_579
timestamp 1713338890
transform 1 0 53050 0 1 44298
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_580
timestamp 1713338890
transform 1 0 55310 0 1 44310
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_581
timestamp 1713338890
transform 1 0 52918 0 1 44430
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_582
timestamp 1713338890
transform 1 0 55178 0 1 44442
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_583
timestamp 1713338890
transform 1 0 52786 0 1 44562
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_584
timestamp 1713338890
transform 1 0 55046 0 1 44574
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_585
timestamp 1713338890
transform 1 0 54914 0 1 44706
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_586
timestamp 1713338890
transform 1 0 54782 0 1 44838
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_587
timestamp 1713338890
transform 1 0 54650 0 1 44970
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_588
timestamp 1713338890
transform 1 0 54518 0 1 45102
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_589
timestamp 1713338890
transform 1 0 54386 0 1 45234
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_590
timestamp 1713338890
transform 1 0 54254 0 1 45366
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_591
timestamp 1713338890
transform 1 0 54122 0 1 45498
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_592
timestamp 1713338890
transform 1 0 53990 0 1 45630
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_593
timestamp 1713338890
transform 1 0 53858 0 1 45762
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_594
timestamp 1713338890
transform 1 0 53726 0 1 45894
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_595
timestamp 1713338890
transform 1 0 53594 0 1 46026
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_596
timestamp 1713338890
transform 1 0 53462 0 1 46158
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_597
timestamp 1713338890
transform 1 0 53330 0 1 46290
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_598
timestamp 1713338890
transform 1 0 53198 0 1 46422
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_599
timestamp 1713338890
transform 1 0 53066 0 1 46554
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_600
timestamp 1713338890
transform 1 0 52934 0 1 46686
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_601
timestamp 1713338890
transform 1 0 52802 0 1 46818
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_602
timestamp 1713338890
transform 1 0 56894 0 1 42726
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_603
timestamp 1713338890
transform 1 0 56762 0 1 42858
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_604
timestamp 1713338890
transform 1 0 60142 0 1 50843
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_605
timestamp 1713338890
transform 1 0 60010 0 1 50975
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_606
timestamp 1713338890
transform 1 0 59878 0 1 51107
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_607
timestamp 1713338890
transform 1 0 59746 0 1 51239
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_608
timestamp 1713338890
transform 1 0 59614 0 1 51371
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_609
timestamp 1713338890
transform 1 0 59482 0 1 51503
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_610
timestamp 1713338890
transform 1 0 59350 0 1 51635
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_611
timestamp 1713338890
transform 1 0 52618 0 1 58367
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_612
timestamp 1713338890
transform 1 0 52486 0 1 58499
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_613
timestamp 1713338890
transform 1 0 52354 0 1 58631
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_614
timestamp 1713338890
transform 1 0 52222 0 1 58763
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_615
timestamp 1713338890
transform 1 0 52090 0 1 58895
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_616
timestamp 1713338890
transform 1 0 51958 0 1 59027
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_617
timestamp 1713338890
transform 1 0 51826 0 1 59159
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_618
timestamp 1713338890
transform 1 0 51694 0 1 59291
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_619
timestamp 1713338890
transform 1 0 51562 0 1 59423
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_620
timestamp 1713338890
transform 1 0 51430 0 1 59555
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_621
timestamp 1713338890
transform 1 0 51298 0 1 59687
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_622
timestamp 1713338890
transform 1 0 51166 0 1 59819
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_623
timestamp 1713338890
transform 1 0 50902 0 1 60083
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_624
timestamp 1713338890
transform 1 0 51034 0 1 59951
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_625
timestamp 1713338890
transform 1 0 50770 0 1 60215
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_626
timestamp 1713338890
transform 1 0 50638 0 1 60347
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_627
timestamp 1713338890
transform 1 0 50506 0 1 60479
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_628
timestamp 1713338890
transform 1 0 52634 0 1 60615
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_629
timestamp 1713338890
transform 1 0 50374 0 1 60611
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_630
timestamp 1713338890
transform 1 0 52502 0 1 60747
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_631
timestamp 1713338890
transform 1 0 50242 0 1 60743
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_632
timestamp 1713338890
transform 1 0 52370 0 1 60879
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_633
timestamp 1713338890
transform 1 0 52238 0 1 61011
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_634
timestamp 1713338890
transform 1 0 52106 0 1 61143
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_635
timestamp 1713338890
transform 1 0 56710 0 1 54275
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_636
timestamp 1713338890
transform 1 0 56578 0 1 54407
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_637
timestamp 1713338890
transform 1 0 56446 0 1 54539
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_638
timestamp 1713338890
transform 1 0 56314 0 1 54671
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_639
timestamp 1713338890
transform 1 0 56182 0 1 54803
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_640
timestamp 1713338890
transform 1 0 56050 0 1 54935
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_641
timestamp 1713338890
transform 1 0 55918 0 1 55067
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_642
timestamp 1713338890
transform 1 0 55786 0 1 55199
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_643
timestamp 1713338890
transform 1 0 55654 0 1 55331
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_644
timestamp 1713338890
transform 1 0 55522 0 1 55463
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_645
timestamp 1713338890
transform 1 0 55390 0 1 55595
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_646
timestamp 1713338890
transform 1 0 55258 0 1 55727
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_647
timestamp 1713338890
transform 1 0 55126 0 1 55859
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_648
timestamp 1713338890
transform 1 0 54994 0 1 55991
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_649
timestamp 1713338890
transform 1 0 54862 0 1 56123
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_650
timestamp 1713338890
transform 1 0 54730 0 1 56255
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_651
timestamp 1713338890
transform 1 0 54598 0 1 56387
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_652
timestamp 1713338890
transform 1 0 56726 0 1 56523
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_653
timestamp 1713338890
transform 1 0 54466 0 1 56519
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_654
timestamp 1713338890
transform 1 0 56594 0 1 56655
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_655
timestamp 1713338890
transform 1 0 54334 0 1 56651
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_656
timestamp 1713338890
transform 1 0 56462 0 1 56787
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_657
timestamp 1713338890
transform 1 0 54202 0 1 56783
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_658
timestamp 1713338890
transform 1 0 54070 0 1 56915
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_659
timestamp 1713338890
transform 1 0 56330 0 1 56919
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_660
timestamp 1713338890
transform 1 0 53938 0 1 57047
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_661
timestamp 1713338890
transform 1 0 56198 0 1 57051
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_662
timestamp 1713338890
transform 1 0 53806 0 1 57179
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_663
timestamp 1713338890
transform 1 0 56066 0 1 57183
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_664
timestamp 1713338890
transform 1 0 53674 0 1 57311
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_665
timestamp 1713338890
transform 1 0 55934 0 1 57315
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_666
timestamp 1713338890
transform 1 0 53542 0 1 57443
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_667
timestamp 1713338890
transform 1 0 55802 0 1 57447
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_668
timestamp 1713338890
transform 1 0 53410 0 1 57575
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_669
timestamp 1713338890
transform 1 0 55670 0 1 57579
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_670
timestamp 1713338890
transform 1 0 53278 0 1 57707
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_671
timestamp 1713338890
transform 1 0 55538 0 1 57711
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_672
timestamp 1713338890
transform 1 0 53146 0 1 57839
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_673
timestamp 1713338890
transform 1 0 55406 0 1 57843
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_674
timestamp 1713338890
transform 1 0 53014 0 1 57971
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_675
timestamp 1713338890
transform 1 0 55274 0 1 57975
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_676
timestamp 1713338890
transform 1 0 52882 0 1 58103
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_677
timestamp 1713338890
transform 1 0 55142 0 1 58107
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_678
timestamp 1713338890
transform 1 0 52750 0 1 58235
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_679
timestamp 1713338890
transform 1 0 55010 0 1 58239
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_680
timestamp 1713338890
transform 1 0 54878 0 1 58371
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_681
timestamp 1713338890
transform 1 0 54746 0 1 58503
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_682
timestamp 1713338890
transform 1 0 54614 0 1 58635
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_683
timestamp 1713338890
transform 1 0 54482 0 1 58767
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_684
timestamp 1713338890
transform 1 0 56742 0 1 58775
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_685
timestamp 1713338890
transform 1 0 54350 0 1 58899
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_686
timestamp 1713338890
transform 1 0 56610 0 1 58907
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_687
timestamp 1713338890
transform 1 0 56478 0 1 59039
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_688
timestamp 1713338890
transform 1 0 54218 0 1 59031
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_689
timestamp 1713338890
transform 1 0 54086 0 1 59163
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_690
timestamp 1713338890
transform 1 0 56346 0 1 59171
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_691
timestamp 1713338890
transform 1 0 53954 0 1 59295
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_692
timestamp 1713338890
transform 1 0 56214 0 1 59303
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_693
timestamp 1713338890
transform 1 0 53822 0 1 59427
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_694
timestamp 1713338890
transform 1 0 56082 0 1 59435
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_695
timestamp 1713338890
transform 1 0 53690 0 1 59559
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_696
timestamp 1713338890
transform 1 0 55950 0 1 59567
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_697
timestamp 1713338890
transform 1 0 53558 0 1 59691
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_698
timestamp 1713338890
transform 1 0 55818 0 1 59699
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_699
timestamp 1713338890
transform 1 0 53426 0 1 59823
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_700
timestamp 1713338890
transform 1 0 55686 0 1 59831
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_701
timestamp 1713338890
transform 1 0 53294 0 1 59955
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_702
timestamp 1713338890
transform 1 0 55554 0 1 59963
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_703
timestamp 1713338890
transform 1 0 53162 0 1 60087
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_704
timestamp 1713338890
transform 1 0 55422 0 1 60095
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_705
timestamp 1713338890
transform 1 0 53030 0 1 60219
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_706
timestamp 1713338890
transform 1 0 55290 0 1 60227
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_707
timestamp 1713338890
transform 1 0 52898 0 1 60351
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_708
timestamp 1713338890
transform 1 0 55158 0 1 60359
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_709
timestamp 1713338890
transform 1 0 52766 0 1 60483
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_710
timestamp 1713338890
transform 1 0 55026 0 1 60491
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_711
timestamp 1713338890
transform 1 0 54894 0 1 60623
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_712
timestamp 1713338890
transform 1 0 54762 0 1 60755
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_713
timestamp 1713338890
transform 1 0 54630 0 1 60887
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_714
timestamp 1713338890
transform 1 0 54498 0 1 61019
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_715
timestamp 1713338890
transform 1 0 56626 0 1 61157
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_716
timestamp 1713338890
transform 1 0 54366 0 1 61151
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_717
timestamp 1713338890
transform 1 0 59218 0 1 51767
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_718
timestamp 1713338890
transform 1 0 59086 0 1 51899
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_719
timestamp 1713338890
transform 1 0 58822 0 1 52163
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_720
timestamp 1713338890
transform 1 0 58954 0 1 52031
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_721
timestamp 1713338890
transform 1 0 58558 0 1 52427
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_722
timestamp 1713338890
transform 1 0 58690 0 1 52295
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_723
timestamp 1713338890
transform 1 0 58426 0 1 52559
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_724
timestamp 1713338890
transform 1 0 58294 0 1 52691
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_725
timestamp 1713338890
transform 1 0 58162 0 1 52823
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_726
timestamp 1713338890
transform 1 0 58030 0 1 52955
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_727
timestamp 1713338890
transform 1 0 57766 0 1 53219
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_728
timestamp 1713338890
transform 1 0 57898 0 1 53087
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_729
timestamp 1713338890
transform 1 0 60026 0 1 53223
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_730
timestamp 1713338890
transform 1 0 60158 0 1 53091
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_731
timestamp 1713338890
transform 1 0 57502 0 1 53483
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_732
timestamp 1713338890
transform 1 0 57634 0 1 53351
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_733
timestamp 1713338890
transform 1 0 59762 0 1 53487
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_734
timestamp 1713338890
transform 1 0 59894 0 1 53355
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_735
timestamp 1713338890
transform 1 0 57238 0 1 53747
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_736
timestamp 1713338890
transform 1 0 57370 0 1 53615
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_737
timestamp 1713338890
transform 1 0 59630 0 1 53619
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_738
timestamp 1713338890
transform 1 0 59498 0 1 53751
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_739
timestamp 1713338890
transform 1 0 56974 0 1 54011
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_740
timestamp 1713338890
transform 1 0 57106 0 1 53879
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_741
timestamp 1713338890
transform 1 0 59234 0 1 54015
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_742
timestamp 1713338890
transform 1 0 59366 0 1 53883
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_743
timestamp 1713338890
transform 1 0 56842 0 1 54143
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_744
timestamp 1713338890
transform 1 0 59102 0 1 54147
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_745
timestamp 1713338890
transform 1 0 58970 0 1 54279
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_746
timestamp 1713338890
transform 1 0 58838 0 1 54411
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_747
timestamp 1713338890
transform 1 0 58706 0 1 54543
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_748
timestamp 1713338890
transform 1 0 58442 0 1 54807
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_749
timestamp 1713338890
transform 1 0 58574 0 1 54675
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_750
timestamp 1713338890
transform 1 0 58310 0 1 54939
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_751
timestamp 1713338890
transform 1 0 58178 0 1 55071
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_752
timestamp 1713338890
transform 1 0 57914 0 1 55335
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_753
timestamp 1713338890
transform 1 0 58046 0 1 55203
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_754
timestamp 1713338890
transform 1 0 60174 0 1 55343
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_755
timestamp 1713338890
transform 1 0 57650 0 1 55599
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_756
timestamp 1713338890
transform 1 0 57782 0 1 55467
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_757
timestamp 1713338890
transform 1 0 60042 0 1 55475
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_758
timestamp 1713338890
transform 1 0 59910 0 1 55607
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_759
timestamp 1713338890
transform 1 0 57386 0 1 55863
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_760
timestamp 1713338890
transform 1 0 57518 0 1 55731
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_761
timestamp 1713338890
transform 1 0 59778 0 1 55739
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_762
timestamp 1713338890
transform 1 0 59646 0 1 55871
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_763
timestamp 1713338890
transform 1 0 57122 0 1 56127
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_764
timestamp 1713338890
transform 1 0 57254 0 1 55995
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_765
timestamp 1713338890
transform 1 0 59514 0 1 56003
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_766
timestamp 1713338890
transform 1 0 59382 0 1 56135
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_767
timestamp 1713338890
transform 1 0 56858 0 1 56391
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_768
timestamp 1713338890
transform 1 0 56990 0 1 56259
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_769
timestamp 1713338890
transform 1 0 59118 0 1 56399
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_770
timestamp 1713338890
transform 1 0 59250 0 1 56267
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_771
timestamp 1713338890
transform 1 0 58854 0 1 56663
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_772
timestamp 1713338890
transform 1 0 58986 0 1 56531
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_773
timestamp 1713338890
transform 1 0 58590 0 1 56927
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_774
timestamp 1713338890
transform 1 0 58722 0 1 56795
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_775
timestamp 1713338890
transform 1 0 58326 0 1 57191
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_776
timestamp 1713338890
transform 1 0 58458 0 1 57059
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_777
timestamp 1713338890
transform 1 0 58062 0 1 57455
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_778
timestamp 1713338890
transform 1 0 58194 0 1 57323
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_779
timestamp 1713338890
transform 1 0 57930 0 1 57587
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_780
timestamp 1713338890
transform 1 0 57798 0 1 57719
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_781
timestamp 1713338890
transform 1 0 60058 0 1 57725
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_782
timestamp 1713338890
transform 1 0 60190 0 1 57593
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_783
timestamp 1713338890
transform 1 0 57534 0 1 57983
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_784
timestamp 1713338890
transform 1 0 57666 0 1 57851
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_785
timestamp 1713338890
transform 1 0 59794 0 1 57989
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_786
timestamp 1713338890
transform 1 0 59926 0 1 57857
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_787
timestamp 1713338890
transform 1 0 57270 0 1 58247
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_788
timestamp 1713338890
transform 1 0 57402 0 1 58115
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_789
timestamp 1713338890
transform 1 0 59530 0 1 58253
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_790
timestamp 1713338890
transform 1 0 59662 0 1 58121
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_791
timestamp 1713338890
transform 1 0 57138 0 1 58379
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_792
timestamp 1713338890
transform 1 0 57006 0 1 58511
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_793
timestamp 1713338890
transform 1 0 59266 0 1 58517
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_794
timestamp 1713338890
transform 1 0 59398 0 1 58385
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_795
timestamp 1713338890
transform 1 0 56874 0 1 58643
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_796
timestamp 1713338890
transform 1 0 59002 0 1 58781
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_797
timestamp 1713338890
transform 1 0 59134 0 1 58649
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_798
timestamp 1713338890
transform 1 0 58870 0 1 58913
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_799
timestamp 1713338890
transform 1 0 58738 0 1 59045
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_800
timestamp 1713338890
transform 1 0 58474 0 1 59309
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_801
timestamp 1713338890
transform 1 0 58606 0 1 59177
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_802
timestamp 1713338890
transform 1 0 58342 0 1 59441
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_803
timestamp 1713338890
transform 1 0 58210 0 1 59573
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_804
timestamp 1713338890
transform 1 0 57946 0 1 59837
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_805
timestamp 1713338890
transform 1 0 58078 0 1 59705
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_806
timestamp 1713338890
transform 1 0 60206 0 1 59840
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_807
timestamp 1713338890
transform 1 0 57814 0 1 59969
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_808
timestamp 1713338890
transform 1 0 57682 0 1 60101
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_809
timestamp 1713338890
transform 1 0 60074 0 1 59972
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_810
timestamp 1713338890
transform 1 0 59942 0 1 60104
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_811
timestamp 1713338890
transform 1 0 57550 0 1 60233
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_812
timestamp 1713338890
transform 1 0 57418 0 1 60365
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_813
timestamp 1713338890
transform 1 0 59678 0 1 60368
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_814
timestamp 1713338890
transform 1 0 59810 0 1 60236
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_815
timestamp 1713338890
transform 1 0 57286 0 1 60497
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_816
timestamp 1713338890
transform 1 0 57154 0 1 60629
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_817
timestamp 1713338890
transform 1 0 59414 0 1 60632
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_818
timestamp 1713338890
transform 1 0 59546 0 1 60500
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_819
timestamp 1713338890
transform 1 0 57022 0 1 60761
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_820
timestamp 1713338890
transform 1 0 56890 0 1 60893
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_821
timestamp 1713338890
transform 1 0 59150 0 1 60896
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_822
timestamp 1713338890
transform 1 0 59282 0 1 60764
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_823
timestamp 1713338890
transform 1 0 56758 0 1 61025
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_824
timestamp 1713338890
transform 1 0 58886 0 1 61160
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_825
timestamp 1713338890
transform 1 0 59018 0 1 61028
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_826
timestamp 1713338890
transform 1 0 51974 0 1 61275
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_827
timestamp 1713338890
transform 1 0 51842 0 1 61407
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_828
timestamp 1713338890
transform 1 0 53838 0 1 61679
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_829
timestamp 1713338890
transform 1 0 53970 0 1 61547
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_830
timestamp 1713338890
transform 1 0 54102 0 1 61415
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_831
timestamp 1713338890
transform 1 0 54234 0 1 61283
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_832
timestamp 1713338890
transform 1 0 53442 0 1 62075
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_833
timestamp 1713338890
transform 1 0 53574 0 1 61943
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_834
timestamp 1713338890
transform 1 0 53706 0 1 61811
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_835
timestamp 1713338890
transform 1 0 56230 0 1 61553
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_836
timestamp 1713338890
transform 1 0 56098 0 1 61685
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_837
timestamp 1713338890
transform 1 0 55966 0 1 61817
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_838
timestamp 1713338890
transform 1 0 55570 0 1 62213
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_839
timestamp 1713338890
transform 1 0 55702 0 1 62081
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_840
timestamp 1713338890
transform 1 0 55834 0 1 61949
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_841
timestamp 1713338890
transform 1 0 55174 0 1 62609
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_842
timestamp 1713338890
transform 1 0 55306 0 1 62477
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_843
timestamp 1713338890
transform 1 0 55438 0 1 62345
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_844
timestamp 1713338890
transform 1 0 55042 0 1 62741
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_845
timestamp 1713338890
transform 1 0 56642 0 1 63404
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_846
timestamp 1713338890
transform 1 0 56362 0 1 61421
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_847
timestamp 1713338890
transform 1 0 56494 0 1 61289
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_848
timestamp 1713338890
transform 1 0 58358 0 1 61688
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_849
timestamp 1713338890
transform 1 0 58490 0 1 61556
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_850
timestamp 1713338890
transform 1 0 58226 0 1 61820
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_851
timestamp 1713338890
transform 1 0 57962 0 1 62084
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_852
timestamp 1713338890
transform 1 0 58094 0 1 61952
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_853
timestamp 1713338890
transform 1 0 57698 0 1 62348
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_854
timestamp 1713338890
transform 1 0 57830 0 1 62216
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_855
timestamp 1713338890
transform 1 0 57566 0 1 62480
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_856
timestamp 1713338890
transform 1 0 57434 0 1 62612
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_857
timestamp 1713338890
transform 1 0 57302 0 1 62744
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_858
timestamp 1713338890
transform 1 0 57170 0 1 62876
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_859
timestamp 1713338890
transform 1 0 57038 0 1 63008
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_860
timestamp 1713338890
transform 1 0 56774 0 1 63272
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_861
timestamp 1713338890
transform 1 0 56906 0 1 63140
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_862
timestamp 1713338890
transform 1 0 58374 0 1 63935
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_863
timestamp 1713338890
transform 1 0 58506 0 1 63803
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_864
timestamp 1713338890
transform 1 0 58242 0 1 64067
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_865
timestamp 1713338890
transform 1 0 58622 0 1 61424
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_866
timestamp 1713338890
transform 1 0 58754 0 1 61292
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_867
timestamp 1713338890
transform 1 0 60222 0 1 62087
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_868
timestamp 1713338890
transform 1 0 60090 0 1 62219
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_869
timestamp 1713338890
transform 1 0 59958 0 1 62351
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_870
timestamp 1713338890
transform 1 0 59826 0 1 62483
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_871
timestamp 1713338890
transform 1 0 59694 0 1 62615
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_872
timestamp 1713338890
transform 1 0 59562 0 1 62747
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_873
timestamp 1713338890
transform 1 0 59430 0 1 62879
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_874
timestamp 1713338890
transform 1 0 59166 0 1 63143
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_875
timestamp 1713338890
transform 1 0 59298 0 1 63011
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_876
timestamp 1713338890
transform 1 0 58902 0 1 63407
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_877
timestamp 1713338890
transform 1 0 59034 0 1 63275
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_878
timestamp 1713338890
transform 1 0 58770 0 1 63539
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_879
timestamp 1713338890
transform 1 0 58638 0 1 63671
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_880
timestamp 1713338890
transform 1 0 60106 0 1 64470
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_881
timestamp 1713338890
transform 1 0 59974 0 1 64602
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_882
timestamp 1713338890
transform 1 0 59842 0 1 64734
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_883
timestamp 1713338890
transform 1 0 60274 0 1 50711
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_884
timestamp 1713338890
transform 1 0 60818 0 1 52431
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_885
timestamp 1713338890
transform 1 0 60950 0 1 52299
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_886
timestamp 1713338890
transform 1 0 60554 0 1 52695
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_887
timestamp 1713338890
transform 1 0 60422 0 1 52827
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_888
timestamp 1713338890
transform 1 0 60290 0 1 52959
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_889
timestamp 1713338890
transform 1 0 60686 0 1 52563
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_890
timestamp 1713338890
transform 1 0 61362 0 1 54155
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_891
timestamp 1713338890
transform 1 0 61494 0 1 54023
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_892
timestamp 1713338890
transform 1 0 61626 0 1 53891
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_893
timestamp 1713338890
transform 1 0 61230 0 1 54287
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_894
timestamp 1713338890
transform 1 0 61098 0 1 54419
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_895
timestamp 1713338890
transform 1 0 60966 0 1 54551
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_896
timestamp 1713338890
transform 1 0 60834 0 1 54683
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_897
timestamp 1713338890
transform 1 0 60702 0 1 54815
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_898
timestamp 1713338890
transform 1 0 60306 0 1 55211
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_899
timestamp 1713338890
transform 1 0 60570 0 1 54947
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_900
timestamp 1713338890
transform 1 0 60438 0 1 55079
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_901
timestamp 1713338890
transform 1 0 62302 0 1 55481
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_902
timestamp 1713338890
transform 1 0 62170 0 1 55613
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_903
timestamp 1713338890
transform 1 0 62038 0 1 55745
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_904
timestamp 1713338890
transform 1 0 61906 0 1 55877
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_905
timestamp 1713338890
transform 1 0 61774 0 1 56009
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_906
timestamp 1713338890
transform 1 0 61642 0 1 56141
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_907
timestamp 1713338890
transform 1 0 61510 0 1 56273
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_908
timestamp 1713338890
transform 1 0 61378 0 1 56405
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_909
timestamp 1713338890
transform 1 0 61246 0 1 56537
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_910
timestamp 1713338890
transform 1 0 60982 0 1 56801
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_911
timestamp 1713338890
transform 1 0 61114 0 1 56669
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_912
timestamp 1713338890
transform 1 0 60718 0 1 57065
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_913
timestamp 1713338890
transform 1 0 60850 0 1 56933
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_914
timestamp 1713338890
transform 1 0 60586 0 1 57197
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_915
timestamp 1713338890
transform 1 0 62846 0 1 57200
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_916
timestamp 1713338890
transform 1 0 62978 0 1 57068
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_917
timestamp 1713338890
transform 1 0 60322 0 1 57461
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_918
timestamp 1713338890
transform 1 0 60454 0 1 57329
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_919
timestamp 1713338890
transform 1 0 62450 0 1 57596
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_920
timestamp 1713338890
transform 1 0 62582 0 1 57464
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_921
timestamp 1713338890
transform 1 0 62714 0 1 57332
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_922
timestamp 1713338890
transform 1 0 62186 0 1 57860
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_923
timestamp 1713338890
transform 1 0 62318 0 1 57728
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_924
timestamp 1713338890
transform 1 0 61922 0 1 58124
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_925
timestamp 1713338890
transform 1 0 62054 0 1 57992
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_926
timestamp 1713338890
transform 1 0 61790 0 1 58256
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_927
timestamp 1713338890
transform 1 0 61658 0 1 58388
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_928
timestamp 1713338890
transform 1 0 61526 0 1 58520
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_929
timestamp 1713338890
transform 1 0 61394 0 1 58652
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_930
timestamp 1713338890
transform 1 0 63654 0 1 58655
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_931
timestamp 1713338890
transform 1 0 61262 0 1 58784
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_932
timestamp 1713338890
transform 1 0 63522 0 1 58787
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_933
timestamp 1713338890
transform 1 0 60998 0 1 59048
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_934
timestamp 1713338890
transform 1 0 61130 0 1 58916
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_935
timestamp 1713338890
transform 1 0 63258 0 1 59051
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_936
timestamp 1713338890
transform 1 0 63390 0 1 58919
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_937
timestamp 1713338890
transform 1 0 60866 0 1 59180
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_938
timestamp 1713338890
transform 1 0 60734 0 1 59312
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_939
timestamp 1713338890
transform 1 0 62994 0 1 59315
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_940
timestamp 1713338890
transform 1 0 63126 0 1 59183
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_941
timestamp 1713338890
transform 1 0 60602 0 1 59444
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_942
timestamp 1713338890
transform 1 0 62862 0 1 59447
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_943
timestamp 1713338890
transform 1 0 60470 0 1 59576
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_944
timestamp 1713338890
transform 1 0 60338 0 1 59708
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_945
timestamp 1713338890
transform 1 0 62598 0 1 59711
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_946
timestamp 1713338890
transform 1 0 62730 0 1 59579
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_947
timestamp 1713338890
transform 1 0 62466 0 1 59843
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_948
timestamp 1713338890
transform 1 0 62202 0 1 60107
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_949
timestamp 1713338890
transform 1 0 62334 0 1 59975
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_950
timestamp 1713338890
transform 1 0 62070 0 1 60239
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_951
timestamp 1713338890
transform 1 0 61806 0 1 60503
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_952
timestamp 1713338890
transform 1 0 61938 0 1 60371
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_953
timestamp 1713338890
transform 1 0 64198 0 1 60378
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_954
timestamp 1713338890
transform 1 0 64066 0 1 60510
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_955
timestamp 1713338890
transform 1 0 61674 0 1 60635
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_956
timestamp 1713338890
transform 1 0 63934 0 1 60642
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_957
timestamp 1713338890
transform 1 0 61542 0 1 60767
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_958
timestamp 1713338890
transform 1 0 61410 0 1 60899
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_959
timestamp 1713338890
transform 1 0 61278 0 1 61031
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_960
timestamp 1713338890
transform 1 0 61146 0 1 61163
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_961
timestamp 1713338890
transform 1 0 61014 0 1 61295
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_962
timestamp 1713338890
transform 1 0 63802 0 1 60774
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_963
timestamp 1713338890
transform 1 0 63670 0 1 60906
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_964
timestamp 1713338890
transform 1 0 63538 0 1 61038
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_965
timestamp 1713338890
transform 1 0 63406 0 1 61170
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_966
timestamp 1713338890
transform 1 0 63274 0 1 61302
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_967
timestamp 1713338890
transform 1 0 60882 0 1 61427
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_968
timestamp 1713338890
transform 1 0 60750 0 1 61559
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_969
timestamp 1713338890
transform 1 0 60618 0 1 61691
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_970
timestamp 1713338890
transform 1 0 60486 0 1 61823
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_971
timestamp 1713338890
transform 1 0 60354 0 1 61955
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_972
timestamp 1713338890
transform 1 0 61954 0 1 62622
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_973
timestamp 1713338890
transform 1 0 61822 0 1 62754
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_974
timestamp 1713338890
transform 1 0 61690 0 1 62886
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_975
timestamp 1713338890
transform 1 0 61558 0 1 63018
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_976
timestamp 1713338890
transform 1 0 61426 0 1 63150
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_977
timestamp 1713338890
transform 1 0 61294 0 1 63282
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_978
timestamp 1713338890
transform 1 0 61162 0 1 63414
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_979
timestamp 1713338890
transform 1 0 61030 0 1 63546
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_980
timestamp 1713338890
transform 1 0 60898 0 1 63678
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_981
timestamp 1713338890
transform 1 0 60766 0 1 63810
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_982
timestamp 1713338890
transform 1 0 60634 0 1 63942
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_983
timestamp 1713338890
transform 1 0 60502 0 1 64074
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_984
timestamp 1713338890
transform 1 0 60370 0 1 64206
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_985
timestamp 1713338890
transform 1 0 60238 0 1 64338
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_986
timestamp 1713338890
transform 1 0 61970 0 1 64871
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_987
timestamp 1713338890
transform 1 0 61838 0 1 65003
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_988
timestamp 1713338890
transform 1 0 61706 0 1 65135
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_989
timestamp 1713338890
transform 1 0 61574 0 1 65267
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_990
timestamp 1713338890
transform 1 0 61442 0 1 65399
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_991
timestamp 1713338890
transform 1 0 63010 0 1 61566
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_992
timestamp 1713338890
transform 1 0 63142 0 1 61434
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_993
timestamp 1713338890
transform 1 0 62878 0 1 61698
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_994
timestamp 1713338890
transform 1 0 62746 0 1 61830
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_995
timestamp 1713338890
transform 1 0 62614 0 1 61962
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_996
timestamp 1713338890
transform 1 0 62482 0 1 62094
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_997
timestamp 1713338890
transform 1 0 62350 0 1 62226
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_998
timestamp 1713338890
transform 1 0 62218 0 1 62358
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_999
timestamp 1713338890
transform 1 0 62086 0 1 62490
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1000
timestamp 1713338890
transform 1 0 63818 0 1 63023
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1001
timestamp 1713338890
transform 1 0 63686 0 1 63155
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1002
timestamp 1713338890
transform 1 0 63554 0 1 63287
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1003
timestamp 1713338890
transform 1 0 63290 0 1 63551
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1004
timestamp 1713338890
transform 1 0 63422 0 1 63419
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1005
timestamp 1713338890
transform 1 0 63158 0 1 63683
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1006
timestamp 1713338890
transform 1 0 63026 0 1 63815
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1007
timestamp 1713338890
transform 1 0 62894 0 1 63947
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1008
timestamp 1713338890
transform 1 0 62762 0 1 64079
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1009
timestamp 1713338890
transform 1 0 62630 0 1 64211
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1010
timestamp 1713338890
transform 1 0 62498 0 1 64343
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1011
timestamp 1713338890
transform 1 0 62366 0 1 64475
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1012
timestamp 1713338890
transform 1 0 62234 0 1 64607
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1013
timestamp 1713338890
transform 1 0 62102 0 1 64739
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1014
timestamp 1713338890
transform 1 0 63570 0 1 65534
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1015
timestamp 1713338890
transform 1 0 63702 0 1 65402
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1016
timestamp 1713338890
transform 1 0 63438 0 1 65666
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1017
timestamp 1713338890
transform 1 0 63306 0 1 65798
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1018
timestamp 1713338890
transform 1 0 63174 0 1 65930
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1019
timestamp 1713338890
transform 1 0 63042 0 1 66062
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1020
timestamp 1713338890
transform 1 0 64362 0 1 64742
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1021
timestamp 1713338890
transform 1 0 64230 0 1 64874
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1022
timestamp 1713338890
transform 1 0 64098 0 1 65006
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1023
timestamp 1713338890
transform 1 0 63966 0 1 65138
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1024
timestamp 1713338890
transform 1 0 64346 0 1 62495
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1025
timestamp 1713338890
transform 1 0 63834 0 1 65270
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1026
timestamp 1713338890
transform 1 0 63950 0 1 62891
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1027
timestamp 1713338890
transform 1 0 64082 0 1 62759
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1028
timestamp 1713338890
transform 1 0 64214 0 1 62627
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1029
timestamp 1713338890
transform 1 0 64874 0 1 61967
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1030
timestamp 1713338890
transform 1 0 64742 0 1 62099
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1031
timestamp 1713338890
transform 1 0 64478 0 1 62363
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1032
timestamp 1713338890
transform 1 0 64610 0 1 62231
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1033
timestamp 1713338890
transform 1 0 65550 0 1 63554
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1034
timestamp 1713338890
transform 1 0 65418 0 1 63686
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1035
timestamp 1713338890
transform 1 0 65286 0 1 63818
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1036
timestamp 1713338890
transform 1 0 65154 0 1 63950
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1037
timestamp 1713338890
transform 1 0 65022 0 1 64082
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1038
timestamp 1713338890
transform 1 0 64758 0 1 64346
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1039
timestamp 1713338890
transform 1 0 64890 0 1 64214
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1040
timestamp 1713338890
transform 1 0 64626 0 1 64478
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1041
timestamp 1713338890
transform 1 0 64494 0 1 64610
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1042
timestamp 1713338890
transform 1 0 66094 0 1 65282
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1043
timestamp 1713338890
transform 1 0 66226 0 1 65150
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1044
timestamp 1713338890
transform 1 0 65830 0 1 65546
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1045
timestamp 1713338890
transform 1 0 65962 0 1 65414
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1046
timestamp 1713338890
transform 1 0 65698 0 1 65678
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1047
timestamp 1713338890
transform 1 0 65566 0 1 65810
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1048
timestamp 1713338890
transform 1 0 65434 0 1 65942
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1049
timestamp 1713338890
transform 1 0 65170 0 1 66206
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1050
timestamp 1713338890
transform 1 0 65302 0 1 66074
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1051
timestamp 1713338890
transform 1 0 65038 0 1 66338
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1052
timestamp 1713338890
transform 1 0 64906 0 1 66470
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1053
timestamp 1713338890
transform 1 0 64774 0 1 66602
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1054
timestamp 1713338890
transform 1 0 64642 0 1 66734
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1055
timestamp 1713338890
transform 1 0 66775 0 1 66864
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1056
timestamp 1713338890
transform 1 0 66511 0 1 67128
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1057
timestamp 1713338890
transform 1 0 66643 0 1 66996
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1058
timestamp 1713338890
transform 1 0 66379 0 1 67260
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1059
timestamp 1713338890
transform 1 0 66247 0 1 67392
box -896 -38 896 38
use M4_M3_CDNS_69033583165212  M4_M3_CDNS_69033583165212_1060
timestamp 1713338890
transform 1 0 66907 0 1 66732
box -896 -38 896 38
use M4_M3_CDNS_69033583165213  M4_M3_CDNS_69033583165213_0
timestamp 1713338890
transform 1 0 14032 0 1 46995
box 28 -38 3140 38
use M4_M3_CDNS_69033583165213  M4_M3_CDNS_69033583165213_1
timestamp 1713338890
transform 1 0 17232 0 1 48331
box 28 -38 3140 38
use M4_M3_CDNS_69033583165213  M4_M3_CDNS_69033583165213_2
timestamp 1713338890
transform 1 0 20432 0 1 49657
box 28 -38 3140 38
use M4_M3_CDNS_69033583165213  M4_M3_CDNS_69033583165213_3
timestamp 1713338890
transform 1 0 26832 0 1 52337
box 28 -38 3140 38
use M4_M3_CDNS_69033583165213  M4_M3_CDNS_69033583165213_4
timestamp 1713338890
transform 1 0 30032 0 1 53675
box 28 -38 3140 38
use M4_M3_CDNS_69033583165213  M4_M3_CDNS_69033583165213_5
timestamp 1713338890
transform 1 0 33232 0 1 55007
box 28 -38 3140 38
use M4_M3_CDNS_69033583165213  M4_M3_CDNS_69033583165213_6
timestamp 1713338890
transform 1 0 36432 0 1 56348
box 28 -38 3140 38
use M4_M3_CDNS_69033583165213  M4_M3_CDNS_69033583165213_7
timestamp 1713338890
transform 1 0 42832 0 1 59024
box 28 -38 3140 38
use M4_M3_CDNS_69033583165213  M4_M3_CDNS_69033583165213_8
timestamp 1713338890
transform 1 0 46032 0 1 60391
box 28 -38 3140 38
use M4_M3_CDNS_69033583165214  M4_M3_CDNS_69033583165214_0
timestamp 1713338890
transform 1 0 47259 0 1 16288
box -3338 -38 38 38
use M4_M3_CDNS_69033583165214  M4_M3_CDNS_69033583165214_1
timestamp 1713338890
transform 1 0 48595 0 1 19488
box -3338 -38 38 38
use M4_M3_CDNS_69033583165214  M4_M3_CDNS_69033583165214_2
timestamp 1713338890
transform 1 0 49921 0 1 22688
box -3338 -38 38 38
use M4_M3_CDNS_69033583165214  M4_M3_CDNS_69033583165214_3
timestamp 1713338890
transform 1 0 52601 0 1 29088
box -3338 -38 38 38
use M4_M3_CDNS_69033583165214  M4_M3_CDNS_69033583165214_4
timestamp 1713338890
transform 1 0 53939 0 1 32288
box -3338 -38 38 38
use M4_M3_CDNS_69033583165214  M4_M3_CDNS_69033583165214_5
timestamp 1713338890
transform 1 0 55271 0 1 35488
box -3338 -38 38 38
use M4_M3_CDNS_69033583165214  M4_M3_CDNS_69033583165214_6
timestamp 1713338890
transform 1 0 56612 0 1 38688
box -3338 -38 38 38
use M4_M3_CDNS_69033583165214  M4_M3_CDNS_69033583165214_7
timestamp 1713338890
transform 1 0 59288 0 1 45088
box -3338 -38 38 38
use M4_M3_CDNS_69033583165215  M4_M3_CDNS_69033583165215_0
timestamp 1713338890
transform 1 0 14032 0 1 46731
box 28 -38 3404 38
use M4_M3_CDNS_69033583165215  M4_M3_CDNS_69033583165215_1
timestamp 1713338890
transform 1 0 17232 0 1 48067
box 28 -38 3404 38
use M4_M3_CDNS_69033583165215  M4_M3_CDNS_69033583165215_2
timestamp 1713338890
transform 1 0 20432 0 1 49393
box 28 -38 3404 38
use M4_M3_CDNS_69033583165215  M4_M3_CDNS_69033583165215_3
timestamp 1713338890
transform 1 0 26832 0 1 52073
box 28 -38 3404 38
use M4_M3_CDNS_69033583165215  M4_M3_CDNS_69033583165215_4
timestamp 1713338890
transform 1 0 30032 0 1 53411
box 28 -38 3404 38
use M4_M3_CDNS_69033583165215  M4_M3_CDNS_69033583165215_5
timestamp 1713338890
transform 1 0 33232 0 1 54743
box 28 -38 3404 38
use M4_M3_CDNS_69033583165215  M4_M3_CDNS_69033583165215_6
timestamp 1713338890
transform 1 0 36432 0 1 56084
box 28 -38 3404 38
use M4_M3_CDNS_69033583165215  M4_M3_CDNS_69033583165215_7
timestamp 1713338890
transform 1 0 42832 0 1 58760
box 28 -38 3404 38
use M4_M3_CDNS_69033583165215  M4_M3_CDNS_69033583165215_8
timestamp 1713338890
transform 1 0 46032 0 1 60127
box 28 -38 3404 38
use M4_M3_CDNS_69033583165216  M4_M3_CDNS_69033583165216_0
timestamp 1713338890
transform 1 0 14032 0 1 46599
box 28 -38 3536 38
use M4_M3_CDNS_69033583165216  M4_M3_CDNS_69033583165216_1
timestamp 1713338890
transform 1 0 17232 0 1 47935
box 28 -38 3536 38
use M4_M3_CDNS_69033583165216  M4_M3_CDNS_69033583165216_2
timestamp 1713338890
transform 1 0 20432 0 1 49261
box 28 -38 3536 38
use M4_M3_CDNS_69033583165216  M4_M3_CDNS_69033583165216_3
timestamp 1713338890
transform 1 0 26832 0 1 51941
box 28 -38 3536 38
use M4_M3_CDNS_69033583165216  M4_M3_CDNS_69033583165216_4
timestamp 1713338890
transform 1 0 30032 0 1 53279
box 28 -38 3536 38
use M4_M3_CDNS_69033583165216  M4_M3_CDNS_69033583165216_5
timestamp 1713338890
transform 1 0 33232 0 1 54611
box 28 -38 3536 38
use M4_M3_CDNS_69033583165216  M4_M3_CDNS_69033583165216_6
timestamp 1713338890
transform 1 0 36432 0 1 55952
box 28 -38 3536 38
use M4_M3_CDNS_69033583165216  M4_M3_CDNS_69033583165216_7
timestamp 1713338890
transform 1 0 42832 0 1 58628
box 28 -38 3536 38
use M4_M3_CDNS_69033583165216  M4_M3_CDNS_69033583165216_8
timestamp 1713338890
transform 1 0 46032 0 1 59995
box 28 -38 3536 38
use M4_M3_CDNS_69033583165217  M4_M3_CDNS_69033583165217_0
timestamp 1713338890
transform 1 0 14032 0 1 46467
box 28 -38 3668 38
use M4_M3_CDNS_69033583165217  M4_M3_CDNS_69033583165217_1
timestamp 1713338890
transform 1 0 17232 0 1 47803
box 28 -38 3668 38
use M4_M3_CDNS_69033583165217  M4_M3_CDNS_69033583165217_2
timestamp 1713338890
transform 1 0 20432 0 1 49129
box 28 -38 3668 38
use M4_M3_CDNS_69033583165217  M4_M3_CDNS_69033583165217_3
timestamp 1713338890
transform 1 0 26832 0 1 51809
box 28 -38 3668 38
use M4_M3_CDNS_69033583165217  M4_M3_CDNS_69033583165217_4
timestamp 1713338890
transform 1 0 30032 0 1 53147
box 28 -38 3668 38
use M4_M3_CDNS_69033583165217  M4_M3_CDNS_69033583165217_5
timestamp 1713338890
transform 1 0 33232 0 1 54479
box 28 -38 3668 38
use M4_M3_CDNS_69033583165217  M4_M3_CDNS_69033583165217_6
timestamp 1713338890
transform 1 0 36432 0 1 55820
box 28 -38 3668 38
use M4_M3_CDNS_69033583165217  M4_M3_CDNS_69033583165217_7
timestamp 1713338890
transform 1 0 42832 0 1 58496
box 28 -38 3668 38
use M4_M3_CDNS_69033583165217  M4_M3_CDNS_69033583165217_8
timestamp 1713338890
transform 1 0 46032 0 1 59863
box 28 -38 3668 38
use M4_M3_CDNS_69033583165218  M4_M3_CDNS_69033583165218_0
timestamp 1713338890
transform 1 0 14032 0 1 46335
box 28 -38 3800 38
use M4_M3_CDNS_69033583165218  M4_M3_CDNS_69033583165218_1
timestamp 1713338890
transform 1 0 17232 0 1 47671
box 28 -38 3800 38
use M4_M3_CDNS_69033583165218  M4_M3_CDNS_69033583165218_2
timestamp 1713338890
transform 1 0 20432 0 1 48997
box 28 -38 3800 38
use M4_M3_CDNS_69033583165218  M4_M3_CDNS_69033583165218_3
timestamp 1713338890
transform 1 0 26832 0 1 51677
box 28 -38 3800 38
use M4_M3_CDNS_69033583165218  M4_M3_CDNS_69033583165218_4
timestamp 1713338890
transform 1 0 30032 0 1 53015
box 28 -38 3800 38
use M4_M3_CDNS_69033583165218  M4_M3_CDNS_69033583165218_5
timestamp 1713338890
transform 1 0 33232 0 1 54347
box 28 -38 3800 38
use M4_M3_CDNS_69033583165218  M4_M3_CDNS_69033583165218_6
timestamp 1713338890
transform 1 0 36432 0 1 55688
box 28 -38 3800 38
use M4_M3_CDNS_69033583165218  M4_M3_CDNS_69033583165218_7
timestamp 1713338890
transform 1 0 42832 0 1 58364
box 28 -38 3800 38
use M4_M3_CDNS_69033583165218  M4_M3_CDNS_69033583165218_8
timestamp 1713338890
transform 1 0 46032 0 1 59731
box 28 -38 3800 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_0
timestamp 1713338890
transform 1 0 45081 0 1 17109
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1
timestamp 1713338890
transform 1 0 44949 0 1 17241
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_2
timestamp 1713338890
transform 1 0 44817 0 1 17373
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_3
timestamp 1713338890
transform 1 0 44685 0 1 17505
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_4
timestamp 1713338890
transform 1 0 44421 0 1 17769
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_5
timestamp 1713338890
transform 1 0 44289 0 1 17901
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_6
timestamp 1713338890
transform 1 0 44553 0 1 17637
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_7
timestamp 1713338890
transform 1 0 43893 0 1 18297
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_8
timestamp 1713338890
transform 1 0 44025 0 1 18165
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_9
timestamp 1713338890
transform 1 0 44157 0 1 18033
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_10
timestamp 1713338890
transform 1 0 43497 0 1 18693
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_11
timestamp 1713338890
transform 1 0 43629 0 1 18561
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_12
timestamp 1713338890
transform 1 0 43761 0 1 18429
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_13
timestamp 1713338890
transform 1 0 43101 0 1 19089
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_14
timestamp 1713338890
transform 1 0 43365 0 1 18825
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_15
timestamp 1713338890
transform 1 0 43233 0 1 18957
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_16
timestamp 1713338890
transform 1 0 42705 0 1 19485
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_17
timestamp 1713338890
transform 1 0 42837 0 1 19353
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_18
timestamp 1713338890
transform 1 0 42969 0 1 19221
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_19
timestamp 1713338890
transform 1 0 42441 0 1 19749
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_20
timestamp 1713338890
transform 1 0 42573 0 1 19617
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_21
timestamp 1713338890
transform 1 0 42177 0 1 20013
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_22
timestamp 1713338890
transform 1 0 42309 0 1 19881
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_23
timestamp 1713338890
transform 1 0 41781 0 1 20409
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_24
timestamp 1713338890
transform 1 0 42045 0 1 20145
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_25
timestamp 1713338890
transform 1 0 41649 0 1 20541
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_26
timestamp 1713338890
transform 1 0 41913 0 1 20277
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_27
timestamp 1713338890
transform 1 0 46301 0 1 20425
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_28
timestamp 1713338890
transform 1 0 46169 0 1 20557
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_29
timestamp 1713338890
transform 1 0 46433 0 1 20293
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_30
timestamp 1713338890
transform 1 0 41517 0 1 20673
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_31
timestamp 1713338890
transform 1 0 41385 0 1 20805
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_32
timestamp 1713338890
transform 1 0 46037 0 1 20689
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_33
timestamp 1713338890
transform 1 0 45905 0 1 20821
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_34
timestamp 1713338890
transform 1 0 41121 0 1 21069
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_35
timestamp 1713338890
transform 1 0 41253 0 1 20937
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_36
timestamp 1713338890
transform 1 0 45773 0 1 20953
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_37
timestamp 1713338890
transform 1 0 45641 0 1 21085
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_38
timestamp 1713338890
transform 1 0 40725 0 1 21465
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_39
timestamp 1713338890
transform 1 0 40857 0 1 21333
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_40
timestamp 1713338890
transform 1 0 40989 0 1 21201
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_41
timestamp 1713338890
transform 1 0 45245 0 1 21481
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_42
timestamp 1713338890
transform 1 0 45509 0 1 21217
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_43
timestamp 1713338890
transform 1 0 45377 0 1 21349
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_44
timestamp 1713338890
transform 1 0 40593 0 1 21597
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_45
timestamp 1713338890
transform 1 0 40461 0 1 21729
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_46
timestamp 1713338890
transform 1 0 45113 0 1 21613
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_47
timestamp 1713338890
transform 1 0 44981 0 1 21745
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_48
timestamp 1713338890
transform 1 0 40197 0 1 21993
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_49
timestamp 1713338890
transform 1 0 40329 0 1 21861
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_50
timestamp 1713338890
transform 1 0 44849 0 1 21877
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_51
timestamp 1713338890
transform 1 0 44717 0 1 22009
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_52
timestamp 1713338890
transform 1 0 38613 0 1 23577
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_53
timestamp 1713338890
transform 1 0 38481 0 1 23709
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_54
timestamp 1713338890
transform 1 0 38349 0 1 23841
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_55
timestamp 1713338890
transform 1 0 38217 0 1 23973
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_56
timestamp 1713338890
transform 1 0 38085 0 1 24105
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_57
timestamp 1713338890
transform 1 0 37953 0 1 24237
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_58
timestamp 1713338890
transform 1 0 37821 0 1 24369
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_59
timestamp 1713338890
transform 1 0 37689 0 1 24501
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_60
timestamp 1713338890
transform 1 0 37557 0 1 24633
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_61
timestamp 1713338890
transform 1 0 37425 0 1 24765
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_62
timestamp 1713338890
transform 1 0 37293 0 1 24897
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_63
timestamp 1713338890
transform 1 0 37161 0 1 25029
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_64
timestamp 1713338890
transform 1 0 40065 0 1 22125
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_65
timestamp 1713338890
transform 1 0 39933 0 1 22257
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_66
timestamp 1713338890
transform 1 0 44585 0 1 22141
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_67
timestamp 1713338890
transform 1 0 44453 0 1 22273
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_68
timestamp 1713338890
transform 1 0 39669 0 1 22521
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_69
timestamp 1713338890
transform 1 0 39801 0 1 22389
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_70
timestamp 1713338890
transform 1 0 44321 0 1 22405
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_71
timestamp 1713338890
transform 1 0 44189 0 1 22537
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_72
timestamp 1713338890
transform 1 0 39405 0 1 22785
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_73
timestamp 1713338890
transform 1 0 39537 0 1 22653
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_74
timestamp 1713338890
transform 1 0 43925 0 1 22801
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_75
timestamp 1713338890
transform 1 0 44057 0 1 22669
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_76
timestamp 1713338890
transform 1 0 39009 0 1 23181
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_77
timestamp 1713338890
transform 1 0 39141 0 1 23049
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_78
timestamp 1713338890
transform 1 0 39273 0 1 22917
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_79
timestamp 1713338890
transform 1 0 43793 0 1 22933
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_80
timestamp 1713338890
transform 1 0 43661 0 1 23065
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_81
timestamp 1713338890
transform 1 0 38877 0 1 23313
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_82
timestamp 1713338890
transform 1 0 38745 0 1 23445
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_83
timestamp 1713338890
transform 1 0 43529 0 1 23197
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_84
timestamp 1713338890
transform 1 0 43397 0 1 23329
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_85
timestamp 1713338890
transform 1 0 43265 0 1 23461
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_86
timestamp 1713338890
transform 1 0 47785 0 1 23467
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_87
timestamp 1713338890
transform 1 0 43133 0 1 23593
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_88
timestamp 1713338890
transform 1 0 43001 0 1 23725
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_89
timestamp 1713338890
transform 1 0 47653 0 1 23599
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_90
timestamp 1713338890
transform 1 0 47521 0 1 23731
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_91
timestamp 1713338890
transform 1 0 42605 0 1 24121
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_92
timestamp 1713338890
transform 1 0 42869 0 1 23857
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_93
timestamp 1713338890
transform 1 0 42737 0 1 23989
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_94
timestamp 1713338890
transform 1 0 47389 0 1 23863
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_95
timestamp 1713338890
transform 1 0 47257 0 1 23995
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_96
timestamp 1713338890
transform 1 0 47125 0 1 24127
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_97
timestamp 1713338890
transform 1 0 42473 0 1 24253
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_98
timestamp 1713338890
transform 1 0 42341 0 1 24385
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_99
timestamp 1713338890
transform 1 0 42209 0 1 24517
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_100
timestamp 1713338890
transform 1 0 46729 0 1 24523
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_101
timestamp 1713338890
transform 1 0 46993 0 1 24259
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_102
timestamp 1713338890
transform 1 0 46861 0 1 24391
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_103
timestamp 1713338890
transform 1 0 42077 0 1 24649
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_104
timestamp 1713338890
transform 1 0 41945 0 1 24781
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_105
timestamp 1713338890
transform 1 0 46465 0 1 24787
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_106
timestamp 1713338890
transform 1 0 46597 0 1 24655
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_107
timestamp 1713338890
transform 1 0 46333 0 1 24919
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_108
timestamp 1713338890
transform 1 0 46201 0 1 25051
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_109
timestamp 1713338890
transform 1 0 41813 0 1 24913
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_110
timestamp 1713338890
transform 1 0 41681 0 1 25045
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_111
timestamp 1713338890
transform 1 0 37029 0 1 25161
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_112
timestamp 1713338890
transform 1 0 36633 0 1 25557
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_113
timestamp 1713338890
transform 1 0 36369 0 1 25821
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_114
timestamp 1713338890
transform 1 0 36237 0 1 25953
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_115
timestamp 1713338890
transform 1 0 36501 0 1 25689
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_116
timestamp 1713338890
transform 1 0 36765 0 1 25425
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_117
timestamp 1713338890
transform 1 0 36897 0 1 25293
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_118
timestamp 1713338890
transform 1 0 35181 0 1 27009
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_119
timestamp 1713338890
transform 1 0 35841 0 1 26349
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_120
timestamp 1713338890
transform 1 0 36105 0 1 26085
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_121
timestamp 1713338890
transform 1 0 35445 0 1 26745
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_122
timestamp 1713338890
transform 1 0 35313 0 1 26877
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_123
timestamp 1713338890
transform 1 0 35577 0 1 26613
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_124
timestamp 1713338890
transform 1 0 35709 0 1 26481
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_125
timestamp 1713338890
transform 1 0 35973 0 1 26217
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_126
timestamp 1713338890
transform 1 0 34917 0 1 27273
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_127
timestamp 1713338890
transform 1 0 34653 0 1 27537
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_128
timestamp 1713338890
transform 1 0 34257 0 1 27933
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_129
timestamp 1713338890
transform 1 0 35049 0 1 27141
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_130
timestamp 1713338890
transform 1 0 34389 0 1 27801
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_131
timestamp 1713338890
transform 1 0 34521 0 1 27669
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_132
timestamp 1713338890
transform 1 0 34785 0 1 27405
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_133
timestamp 1713338890
transform 1 0 41549 0 1 25177
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_134
timestamp 1713338890
transform 1 0 46069 0 1 25183
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_135
timestamp 1713338890
transform 1 0 41417 0 1 25309
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_136
timestamp 1713338890
transform 1 0 41285 0 1 25441
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_137
timestamp 1713338890
transform 1 0 45937 0 1 25315
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_138
timestamp 1713338890
transform 1 0 45805 0 1 25447
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_139
timestamp 1713338890
transform 1 0 41021 0 1 25705
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_140
timestamp 1713338890
transform 1 0 41153 0 1 25573
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_141
timestamp 1713338890
transform 1 0 45673 0 1 25579
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_142
timestamp 1713338890
transform 1 0 45541 0 1 25711
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_143
timestamp 1713338890
transform 1 0 40889 0 1 25837
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_144
timestamp 1713338890
transform 1 0 40757 0 1 25969
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_145
timestamp 1713338890
transform 1 0 45277 0 1 25975
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_146
timestamp 1713338890
transform 1 0 45409 0 1 25843
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_147
timestamp 1713338890
transform 1 0 40625 0 1 26101
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_148
timestamp 1713338890
transform 1 0 45145 0 1 26107
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_149
timestamp 1713338890
transform 1 0 40493 0 1 26233
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_150
timestamp 1713338890
transform 1 0 45013 0 1 26239
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_151
timestamp 1713338890
transform 1 0 40361 0 1 26365
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_152
timestamp 1713338890
transform 1 0 40229 0 1 26497
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_153
timestamp 1713338890
transform 1 0 44881 0 1 26371
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_154
timestamp 1713338890
transform 1 0 44749 0 1 26503
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_155
timestamp 1713338890
transform 1 0 40097 0 1 26629
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_156
timestamp 1713338890
transform 1 0 44617 0 1 26635
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_157
timestamp 1713338890
transform 1 0 39965 0 1 26761
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_158
timestamp 1713338890
transform 1 0 39833 0 1 26893
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_159
timestamp 1713338890
transform 1 0 44485 0 1 26767
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_160
timestamp 1713338890
transform 1 0 44353 0 1 26899
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_161
timestamp 1713338890
transform 1 0 39701 0 1 27025
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_162
timestamp 1713338890
transform 1 0 44221 0 1 27031
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_163
timestamp 1713338890
transform 1 0 39569 0 1 27157
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_164
timestamp 1713338890
transform 1 0 39437 0 1 27289
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_165
timestamp 1713338890
transform 1 0 44089 0 1 27163
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_166
timestamp 1713338890
transform 1 0 39305 0 1 27421
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_167
timestamp 1713338890
transform 1 0 43825 0 1 27427
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_168
timestamp 1713338890
transform 1 0 43957 0 1 27295
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_169
timestamp 1713338890
transform 1 0 39173 0 1 27553
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_170
timestamp 1713338890
transform 1 0 43693 0 1 27559
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_171
timestamp 1713338890
transform 1 0 39041 0 1 27685
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_172
timestamp 1713338890
transform 1 0 38909 0 1 27817
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_173
timestamp 1713338890
transform 1 0 43561 0 1 27691
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_174
timestamp 1713338890
transform 1 0 43429 0 1 27823
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_175
timestamp 1713338890
transform 1 0 38777 0 1 27949
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_176
timestamp 1713338890
transform 1 0 43297 0 1 27955
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_177
timestamp 1713338890
transform 1 0 33993 0 1 28197
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_178
timestamp 1713338890
transform 1 0 33729 0 1 28461
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_179
timestamp 1713338890
transform 1 0 33861 0 1 28329
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_180
timestamp 1713338890
transform 1 0 34125 0 1 28065
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_181
timestamp 1713338890
transform 1 0 38645 0 1 28081
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_182
timestamp 1713338890
transform 1 0 38513 0 1 28213
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_183
timestamp 1713338890
transform 1 0 38381 0 1 28345
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_184
timestamp 1713338890
transform 1 0 33597 0 1 28593
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_185
timestamp 1713338890
transform 1 0 33333 0 1 28857
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_186
timestamp 1713338890
transform 1 0 33465 0 1 28725
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_187
timestamp 1713338890
transform 1 0 38117 0 1 28609
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_188
timestamp 1713338890
transform 1 0 37985 0 1 28741
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_189
timestamp 1713338890
transform 1 0 38249 0 1 28477
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_190
timestamp 1713338890
transform 1 0 37853 0 1 28873
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_191
timestamp 1713338890
transform 1 0 33069 0 1 29121
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_192
timestamp 1713338890
transform 1 0 32937 0 1 29253
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_193
timestamp 1713338890
transform 1 0 33201 0 1 28989
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_194
timestamp 1713338890
transform 1 0 37457 0 1 29269
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_195
timestamp 1713338890
transform 1 0 37721 0 1 29005
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_196
timestamp 1713338890
transform 1 0 37589 0 1 29137
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_197
timestamp 1713338890
transform 1 0 32541 0 1 29649
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_198
timestamp 1713338890
transform 1 0 32805 0 1 29385
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_199
timestamp 1713338890
transform 1 0 32673 0 1 29517
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_200
timestamp 1713338890
transform 1 0 37325 0 1 29401
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_201
timestamp 1713338890
transform 1 0 37193 0 1 29533
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_202
timestamp 1713338890
transform 1 0 37061 0 1 29665
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_203
timestamp 1713338890
transform 1 0 32277 0 1 29913
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_204
timestamp 1713338890
transform 1 0 32409 0 1 29781
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_205
timestamp 1713338890
transform 1 0 32145 0 1 30045
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_206
timestamp 1713338890
transform 1 0 36797 0 1 29929
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_207
timestamp 1713338890
transform 1 0 36929 0 1 29797
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_208
timestamp 1713338890
transform 1 0 36665 0 1 30061
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_209
timestamp 1713338890
transform 1 0 31749 0 1 30441
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_210
timestamp 1713338890
transform 1 0 32013 0 1 30177
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_211
timestamp 1713338890
transform 1 0 31881 0 1 30309
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_212
timestamp 1713338890
transform 1 0 31617 0 1 30573
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_213
timestamp 1713338890
transform 1 0 36533 0 1 30193
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_214
timestamp 1713338890
transform 1 0 36401 0 1 30325
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_215
timestamp 1713338890
transform 1 0 36269 0 1 30457
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_216
timestamp 1713338890
transform 1 0 36137 0 1 30589
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_217
timestamp 1713338890
transform 1 0 31221 0 1 30969
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_218
timestamp 1713338890
transform 1 0 31353 0 1 30837
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_219
timestamp 1713338890
transform 1 0 31485 0 1 30705
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_220
timestamp 1713338890
transform 1 0 36005 0 1 30721
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_221
timestamp 1713338890
transform 1 0 35873 0 1 30853
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_222
timestamp 1713338890
transform 1 0 35741 0 1 30985
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_223
timestamp 1713338890
transform 1 0 43165 0 1 28087
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_224
timestamp 1713338890
transform 1 0 43033 0 1 28219
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_225
timestamp 1713338890
transform 1 0 42901 0 1 28351
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_226
timestamp 1713338890
transform 1 0 42637 0 1 28615
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_227
timestamp 1713338890
transform 1 0 42769 0 1 28483
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_228
timestamp 1713338890
transform 1 0 42505 0 1 28747
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_229
timestamp 1713338890
transform 1 0 42373 0 1 28879
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_230
timestamp 1713338890
transform 1 0 42241 0 1 29011
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_231
timestamp 1713338890
transform 1 0 42109 0 1 29143
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_232
timestamp 1713338890
transform 1 0 41977 0 1 29275
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_233
timestamp 1713338890
transform 1 0 41845 0 1 29407
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_234
timestamp 1713338890
transform 1 0 41713 0 1 29539
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_235
timestamp 1713338890
transform 1 0 41581 0 1 29671
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_236
timestamp 1713338890
transform 1 0 41449 0 1 29803
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_237
timestamp 1713338890
transform 1 0 41317 0 1 29935
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_238
timestamp 1713338890
transform 1 0 41185 0 1 30067
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_239
timestamp 1713338890
transform 1 0 50357 0 1 29975
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_240
timestamp 1713338890
transform 1 0 41053 0 1 30199
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_241
timestamp 1713338890
transform 1 0 50093 0 1 30239
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_242
timestamp 1713338890
transform 1 0 50225 0 1 30107
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_243
timestamp 1713338890
transform 1 0 40921 0 1 30331
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_244
timestamp 1713338890
transform 1 0 49961 0 1 30371
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_245
timestamp 1713338890
transform 1 0 40789 0 1 30463
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_246
timestamp 1713338890
transform 1 0 40657 0 1 30595
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_247
timestamp 1713338890
transform 1 0 49829 0 1 30503
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_248
timestamp 1713338890
transform 1 0 49697 0 1 30635
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_249
timestamp 1713338890
transform 1 0 40525 0 1 30727
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_250
timestamp 1713338890
transform 1 0 49565 0 1 30767
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_251
timestamp 1713338890
transform 1 0 40393 0 1 30859
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_252
timestamp 1713338890
transform 1 0 40261 0 1 30991
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_253
timestamp 1713338890
transform 1 0 49433 0 1 30899
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_254
timestamp 1713338890
transform 1 0 31089 0 1 31101
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_255
timestamp 1713338890
transform 1 0 30957 0 1 31233
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_256
timestamp 1713338890
transform 1 0 35609 0 1 31117
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_257
timestamp 1713338890
transform 1 0 35477 0 1 31249
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_258
timestamp 1713338890
transform 1 0 30561 0 1 31629
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_259
timestamp 1713338890
transform 1 0 30825 0 1 31365
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_260
timestamp 1713338890
transform 1 0 30693 0 1 31497
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_261
timestamp 1713338890
transform 1 0 35213 0 1 31513
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_262
timestamp 1713338890
transform 1 0 35081 0 1 31645
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_263
timestamp 1713338890
transform 1 0 35345 0 1 31381
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_264
timestamp 1713338890
transform 1 0 30297 0 1 31893
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_265
timestamp 1713338890
transform 1 0 30429 0 1 31761
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_266
timestamp 1713338890
transform 1 0 34949 0 1 31777
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_267
timestamp 1713338890
transform 1 0 34817 0 1 31909
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_268
timestamp 1713338890
transform 1 0 30165 0 1 32025
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_269
timestamp 1713338890
transform 1 0 29901 0 1 32289
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_270
timestamp 1713338890
transform 1 0 30033 0 1 32157
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_271
timestamp 1713338890
transform 1 0 34685 0 1 32041
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_272
timestamp 1713338890
transform 1 0 34553 0 1 32173
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_273
timestamp 1713338890
transform 1 0 34421 0 1 32305
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_274
timestamp 1713338890
transform 1 0 29637 0 1 32553
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_275
timestamp 1713338890
transform 1 0 29769 0 1 32421
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_276
timestamp 1713338890
transform 1 0 34289 0 1 32437
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_277
timestamp 1713338890
transform 1 0 34157 0 1 32569
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_278
timestamp 1713338890
transform 1 0 38677 0 1 32575
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_279
timestamp 1713338890
transform 1 0 29373 0 1 32817
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_280
timestamp 1713338890
transform 1 0 29505 0 1 32685
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_281
timestamp 1713338890
transform 1 0 29241 0 1 32949
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_282
timestamp 1713338890
transform 1 0 34025 0 1 32701
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_283
timestamp 1713338890
transform 1 0 33893 0 1 32833
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_284
timestamp 1713338890
transform 1 0 33761 0 1 32965
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_285
timestamp 1713338890
transform 1 0 38545 0 1 32707
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_286
timestamp 1713338890
transform 1 0 38413 0 1 32839
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_287
timestamp 1713338890
transform 1 0 38281 0 1 32971
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_288
timestamp 1713338890
transform 1 0 28977 0 1 33213
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_289
timestamp 1713338890
transform 1 0 29109 0 1 33081
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_290
timestamp 1713338890
transform 1 0 33629 0 1 33097
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_291
timestamp 1713338890
transform 1 0 33497 0 1 33229
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_292
timestamp 1713338890
transform 1 0 38149 0 1 33103
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_293
timestamp 1713338890
transform 1 0 38017 0 1 33235
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_294
timestamp 1713338890
transform 1 0 28581 0 1 33609
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_295
timestamp 1713338890
transform 1 0 28713 0 1 33477
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_296
timestamp 1713338890
transform 1 0 28845 0 1 33345
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_297
timestamp 1713338890
transform 1 0 33365 0 1 33361
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_298
timestamp 1713338890
transform 1 0 33233 0 1 33493
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_299
timestamp 1713338890
transform 1 0 33101 0 1 33625
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_300
timestamp 1713338890
transform 1 0 37753 0 1 33499
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_301
timestamp 1713338890
transform 1 0 37621 0 1 33631
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_302
timestamp 1713338890
transform 1 0 37885 0 1 33367
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_303
timestamp 1713338890
transform 1 0 28449 0 1 33741
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_304
timestamp 1713338890
transform 1 0 28317 0 1 33873
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_305
timestamp 1713338890
transform 1 0 32969 0 1 33757
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_306
timestamp 1713338890
transform 1 0 32837 0 1 33889
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_307
timestamp 1713338890
transform 1 0 37489 0 1 33763
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_308
timestamp 1713338890
transform 1 0 37357 0 1 33895
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_309
timestamp 1713338890
transform 1 0 40129 0 1 31123
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_310
timestamp 1713338890
transform 1 0 49301 0 1 31031
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_311
timestamp 1713338890
transform 1 0 49169 0 1 31163
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_312
timestamp 1713338890
transform 1 0 39997 0 1 31255
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_313
timestamp 1713338890
transform 1 0 49037 0 1 31295
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_314
timestamp 1713338890
transform 1 0 39865 0 1 31387
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_315
timestamp 1713338890
transform 1 0 48905 0 1 31427
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_316
timestamp 1713338890
transform 1 0 39601 0 1 31651
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_317
timestamp 1713338890
transform 1 0 39733 0 1 31519
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_318
timestamp 1713338890
transform 1 0 48773 0 1 31559
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_319
timestamp 1713338890
transform 1 0 39469 0 1 31783
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_320
timestamp 1713338890
transform 1 0 48641 0 1 31691
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_321
timestamp 1713338890
transform 1 0 48509 0 1 31823
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_322
timestamp 1713338890
transform 1 0 39337 0 1 31915
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_323
timestamp 1713338890
transform 1 0 48377 0 1 31955
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_324
timestamp 1713338890
transform 1 0 39205 0 1 32047
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_325
timestamp 1713338890
transform 1 0 48245 0 1 32087
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_326
timestamp 1713338890
transform 1 0 39073 0 1 32179
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_327
timestamp 1713338890
transform 1 0 38941 0 1 32311
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_328
timestamp 1713338890
transform 1 0 48113 0 1 32219
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_329
timestamp 1713338890
transform 1 0 38809 0 1 32443
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_330
timestamp 1713338890
transform 1 0 47981 0 1 32351
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_331
timestamp 1713338890
transform 1 0 47849 0 1 32483
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_332
timestamp 1713338890
transform 1 0 47717 0 1 32615
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_333
timestamp 1713338890
transform 1 0 47585 0 1 32747
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_334
timestamp 1713338890
transform 1 0 47453 0 1 32879
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_335
timestamp 1713338890
transform 1 0 47321 0 1 33011
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_336
timestamp 1713338890
transform 1 0 47189 0 1 33143
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_337
timestamp 1713338890
transform 1 0 51709 0 1 33161
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_338
timestamp 1713338890
transform 1 0 47057 0 1 33275
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_339
timestamp 1713338890
transform 1 0 46925 0 1 33407
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_340
timestamp 1713338890
transform 1 0 51577 0 1 33293
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_341
timestamp 1713338890
transform 1 0 51445 0 1 33425
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_342
timestamp 1713338890
transform 1 0 46793 0 1 33539
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_343
timestamp 1713338890
transform 1 0 51313 0 1 33557
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_344
timestamp 1713338890
transform 1 0 46529 0 1 33803
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_345
timestamp 1713338890
transform 1 0 46661 0 1 33671
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_346
timestamp 1713338890
transform 1 0 51181 0 1 33689
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_347
timestamp 1713338890
transform 1 0 46397 0 1 33935
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_348
timestamp 1713338890
transform 1 0 51049 0 1 33821
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_349
timestamp 1713338890
transform 1 0 50917 0 1 33953
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_350
timestamp 1713338890
transform 1 0 28053 0 1 34137
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_351
timestamp 1713338890
transform 1 0 28185 0 1 34005
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_352
timestamp 1713338890
transform 1 0 27921 0 1 34269
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_353
timestamp 1713338890
transform 1 0 32573 0 1 34153
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_354
timestamp 1713338890
transform 1 0 32705 0 1 34021
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_355
timestamp 1713338890
transform 1 0 37225 0 1 34027
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_356
timestamp 1713338890
transform 1 0 37093 0 1 34159
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_357
timestamp 1713338890
transform 1 0 27789 0 1 34401
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_358
timestamp 1713338890
transform 1 0 27657 0 1 34533
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_359
timestamp 1713338890
transform 1 0 32441 0 1 34285
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_360
timestamp 1713338890
transform 1 0 32309 0 1 34417
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_361
timestamp 1713338890
transform 1 0 36829 0 1 34423
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_362
timestamp 1713338890
transform 1 0 36961 0 1 34291
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_363
timestamp 1713338890
transform 1 0 27393 0 1 34797
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_364
timestamp 1713338890
transform 1 0 27525 0 1 34665
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_365
timestamp 1713338890
transform 1 0 32177 0 1 34549
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_366
timestamp 1713338890
transform 1 0 32045 0 1 34681
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_367
timestamp 1713338890
transform 1 0 31913 0 1 34813
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_368
timestamp 1713338890
transform 1 0 36697 0 1 34555
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_369
timestamp 1713338890
transform 1 0 36565 0 1 34687
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_370
timestamp 1713338890
transform 1 0 27129 0 1 35061
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_371
timestamp 1713338890
transform 1 0 27261 0 1 34929
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_372
timestamp 1713338890
transform 1 0 31781 0 1 34945
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_373
timestamp 1713338890
transform 1 0 31649 0 1 35077
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_374
timestamp 1713338890
transform 1 0 36433 0 1 34819
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_375
timestamp 1713338890
transform 1 0 36301 0 1 34951
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_376
timestamp 1713338890
transform 1 0 36169 0 1 35083
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_377
timestamp 1713338890
transform 1 0 26865 0 1 35325
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_378
timestamp 1713338890
transform 1 0 26997 0 1 35193
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_379
timestamp 1713338890
transform 1 0 31517 0 1 35209
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_380
timestamp 1713338890
transform 1 0 31385 0 1 35341
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_381
timestamp 1713338890
transform 1 0 36037 0 1 35215
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_382
timestamp 1713338890
transform 1 0 35905 0 1 35347
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_383
timestamp 1713338890
transform 1 0 26601 0 1 35589
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_384
timestamp 1713338890
transform 1 0 26733 0 1 35457
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_385
timestamp 1713338890
transform 1 0 31121 0 1 35605
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_386
timestamp 1713338890
transform 1 0 31253 0 1 35473
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_387
timestamp 1713338890
transform 1 0 35773 0 1 35479
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_388
timestamp 1713338890
transform 1 0 35641 0 1 35611
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_389
timestamp 1713338890
transform 1 0 26337 0 1 35853
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_390
timestamp 1713338890
transform 1 0 26469 0 1 35721
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_391
timestamp 1713338890
transform 1 0 30989 0 1 35737
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_392
timestamp 1713338890
transform 1 0 30857 0 1 35869
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_393
timestamp 1713338890
transform 1 0 35377 0 1 35875
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_394
timestamp 1713338890
transform 1 0 35509 0 1 35743
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_395
timestamp 1713338890
transform 1 0 26073 0 1 36117
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_396
timestamp 1713338890
transform 1 0 26205 0 1 35985
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_397
timestamp 1713338890
transform 1 0 30725 0 1 36001
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_398
timestamp 1713338890
transform 1 0 30593 0 1 36133
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_399
timestamp 1713338890
transform 1 0 35245 0 1 36007
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_400
timestamp 1713338890
transform 1 0 35113 0 1 36139
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_401
timestamp 1713338890
transform 1 0 25809 0 1 36381
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_402
timestamp 1713338890
transform 1 0 25941 0 1 36249
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_403
timestamp 1713338890
transform 1 0 30461 0 1 36265
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_404
timestamp 1713338890
transform 1 0 30329 0 1 36397
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_405
timestamp 1713338890
transform 1 0 34981 0 1 36271
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_406
timestamp 1713338890
transform 1 0 34849 0 1 36403
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_407
timestamp 1713338890
transform 1 0 25677 0 1 36513
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_408
timestamp 1713338890
transform 1 0 25545 0 1 36645
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_409
timestamp 1713338890
transform 1 0 30197 0 1 36529
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_410
timestamp 1713338890
transform 1 0 30065 0 1 36661
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_411
timestamp 1713338890
transform 1 0 34717 0 1 36535
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_412
timestamp 1713338890
transform 1 0 34585 0 1 36667
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_413
timestamp 1713338890
transform 1 0 25413 0 1 36777
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_414
timestamp 1713338890
transform 1 0 25281 0 1 36909
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_415
timestamp 1713338890
transform 1 0 29933 0 1 36793
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_416
timestamp 1713338890
transform 1 0 29801 0 1 36925
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_417
timestamp 1713338890
transform 1 0 34453 0 1 36799
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_418
timestamp 1713338890
transform 1 0 34321 0 1 36931
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_419
timestamp 1713338890
transform 1 0 46265 0 1 34067
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_420
timestamp 1713338890
transform 1 0 50785 0 1 34085
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_421
timestamp 1713338890
transform 1 0 46001 0 1 34331
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_422
timestamp 1713338890
transform 1 0 46133 0 1 34199
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_423
timestamp 1713338890
transform 1 0 50653 0 1 34217
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_424
timestamp 1713338890
transform 1 0 45869 0 1 34463
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_425
timestamp 1713338890
transform 1 0 50521 0 1 34349
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_426
timestamp 1713338890
transform 1 0 50389 0 1 34481
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_427
timestamp 1713338890
transform 1 0 45737 0 1 34595
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_428
timestamp 1713338890
transform 1 0 50257 0 1 34613
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_429
timestamp 1713338890
transform 1 0 45605 0 1 34727
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_430
timestamp 1713338890
transform 1 0 50125 0 1 34745
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_431
timestamp 1713338890
transform 1 0 45473 0 1 34859
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_432
timestamp 1713338890
transform 1 0 45341 0 1 34991
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_433
timestamp 1713338890
transform 1 0 49993 0 1 34877
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_434
timestamp 1713338890
transform 1 0 45209 0 1 35123
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_435
timestamp 1713338890
transform 1 0 49861 0 1 35009
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_436
timestamp 1713338890
transform 1 0 49729 0 1 35141
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_437
timestamp 1713338890
transform 1 0 45077 0 1 35255
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_438
timestamp 1713338890
transform 1 0 49597 0 1 35273
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_439
timestamp 1713338890
transform 1 0 44945 0 1 35387
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_440
timestamp 1713338890
transform 1 0 49465 0 1 35405
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_441
timestamp 1713338890
transform 1 0 44813 0 1 35519
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_442
timestamp 1713338890
transform 1 0 49333 0 1 35537
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_443
timestamp 1713338890
transform 1 0 44549 0 1 35783
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_444
timestamp 1713338890
transform 1 0 44681 0 1 35651
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_445
timestamp 1713338890
transform 1 0 49201 0 1 35669
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_446
timestamp 1713338890
transform 1 0 44417 0 1 35915
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_447
timestamp 1713338890
transform 1 0 48937 0 1 35933
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_448
timestamp 1713338890
transform 1 0 49069 0 1 35801
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_449
timestamp 1713338890
transform 1 0 44285 0 1 36047
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_450
timestamp 1713338890
transform 1 0 48805 0 1 36065
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_451
timestamp 1713338890
transform 1 0 44153 0 1 36179
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_452
timestamp 1713338890
transform 1 0 48673 0 1 36197
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_453
timestamp 1713338890
transform 1 0 44021 0 1 36311
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_454
timestamp 1713338890
transform 1 0 48541 0 1 36329
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_455
timestamp 1713338890
transform 1 0 53061 0 1 36341
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_456
timestamp 1713338890
transform 1 0 43889 0 1 36443
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_457
timestamp 1713338890
transform 1 0 48409 0 1 36461
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_458
timestamp 1713338890
transform 1 0 52929 0 1 36473
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_459
timestamp 1713338890
transform 1 0 43757 0 1 36575
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_460
timestamp 1713338890
transform 1 0 48277 0 1 36593
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_461
timestamp 1713338890
transform 1 0 52797 0 1 36605
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_462
timestamp 1713338890
transform 1 0 43625 0 1 36707
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_463
timestamp 1713338890
transform 1 0 48145 0 1 36725
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_464
timestamp 1713338890
transform 1 0 52665 0 1 36737
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_465
timestamp 1713338890
transform 1 0 43493 0 1 36839
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_466
timestamp 1713338890
transform 1 0 43361 0 1 36971
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_467
timestamp 1713338890
transform 1 0 48013 0 1 36857
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_468
timestamp 1713338890
transform 1 0 52533 0 1 36869
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_469
timestamp 1713338890
transform 1 0 25149 0 1 37041
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_470
timestamp 1713338890
transform 1 0 25017 0 1 37173
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_471
timestamp 1713338890
transform 1 0 29669 0 1 37057
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_472
timestamp 1713338890
transform 1 0 34189 0 1 37063
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_473
timestamp 1713338890
transform 1 0 24885 0 1 37305
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_474
timestamp 1713338890
transform 1 0 29537 0 1 37189
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_475
timestamp 1713338890
transform 1 0 29405 0 1 37321
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_476
timestamp 1713338890
transform 1 0 34057 0 1 37195
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_477
timestamp 1713338890
transform 1 0 33925 0 1 37327
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_478
timestamp 1713338890
transform 1 0 24753 0 1 37437
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_479
timestamp 1713338890
transform 1 0 24621 0 1 37569
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_480
timestamp 1713338890
transform 1 0 29273 0 1 37453
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_481
timestamp 1713338890
transform 1 0 33793 0 1 37459
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_482
timestamp 1713338890
transform 1 0 24489 0 1 37701
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_483
timestamp 1713338890
transform 1 0 29141 0 1 37585
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_484
timestamp 1713338890
transform 1 0 29009 0 1 37717
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_485
timestamp 1713338890
transform 1 0 33661 0 1 37591
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_486
timestamp 1713338890
transform 1 0 33529 0 1 37723
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_487
timestamp 1713338890
transform 1 0 24225 0 1 37965
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_488
timestamp 1713338890
transform 1 0 24357 0 1 37833
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_489
timestamp 1713338890
transform 1 0 28877 0 1 37849
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_490
timestamp 1713338890
transform 1 0 33397 0 1 37855
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_491
timestamp 1713338890
transform 1 0 24093 0 1 38097
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_492
timestamp 1713338890
transform 1 0 28613 0 1 38113
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_493
timestamp 1713338890
transform 1 0 28745 0 1 37981
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_494
timestamp 1713338890
transform 1 0 33133 0 1 38119
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_495
timestamp 1713338890
transform 1 0 33265 0 1 37987
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_496
timestamp 1713338890
transform 1 0 23961 0 1 38229
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_497
timestamp 1713338890
transform 1 0 23829 0 1 38361
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_498
timestamp 1713338890
transform 1 0 28481 0 1 38245
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_499
timestamp 1713338890
transform 1 0 33001 0 1 38251
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_500
timestamp 1713338890
transform 1 0 23697 0 1 38493
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_501
timestamp 1713338890
transform 1 0 28349 0 1 38377
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_502
timestamp 1713338890
transform 1 0 28217 0 1 38509
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_503
timestamp 1713338890
transform 1 0 32869 0 1 38383
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_504
timestamp 1713338890
transform 1 0 32737 0 1 38515
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_505
timestamp 1713338890
transform 1 0 23565 0 1 38625
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_506
timestamp 1713338890
transform 1 0 23433 0 1 38757
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_507
timestamp 1713338890
transform 1 0 28085 0 1 38641
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_508
timestamp 1713338890
transform 1 0 32605 0 1 38647
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_509
timestamp 1713338890
transform 1 0 23301 0 1 38889
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_510
timestamp 1713338890
transform 1 0 27953 0 1 38773
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_511
timestamp 1713338890
transform 1 0 27821 0 1 38905
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_512
timestamp 1713338890
transform 1 0 32341 0 1 38911
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_513
timestamp 1713338890
transform 1 0 32473 0 1 38779
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_514
timestamp 1713338890
transform 1 0 23169 0 1 39021
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_515
timestamp 1713338890
transform 1 0 23037 0 1 39153
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_516
timestamp 1713338890
transform 1 0 27689 0 1 39037
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_517
timestamp 1713338890
transform 1 0 32209 0 1 39043
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_518
timestamp 1713338890
transform 1 0 22905 0 1 39285
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_519
timestamp 1713338890
transform 1 0 27557 0 1 39169
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_520
timestamp 1713338890
transform 1 0 27425 0 1 39301
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_521
timestamp 1713338890
transform 1 0 32077 0 1 39175
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_522
timestamp 1713338890
transform 1 0 31945 0 1 39307
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_523
timestamp 1713338890
transform 1 0 22641 0 1 39549
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_524
timestamp 1713338890
transform 1 0 22773 0 1 39417
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_525
timestamp 1713338890
transform 1 0 27293 0 1 39433
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_526
timestamp 1713338890
transform 1 0 31813 0 1 39439
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_527
timestamp 1713338890
transform 1 0 22509 0 1 39681
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_528
timestamp 1713338890
transform 1 0 27161 0 1 39565
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_529
timestamp 1713338890
transform 1 0 27029 0 1 39697
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_530
timestamp 1713338890
transform 1 0 31681 0 1 39571
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_531
timestamp 1713338890
transform 1 0 31549 0 1 39703
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_532
timestamp 1713338890
transform 1 0 22245 0 1 39945
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_533
timestamp 1713338890
transform 1 0 22377 0 1 39813
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_534
timestamp 1713338890
transform 1 0 26897 0 1 39829
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_535
timestamp 1713338890
transform 1 0 31417 0 1 39835
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_536
timestamp 1713338890
transform 1 0 26765 0 1 39961
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_537
timestamp 1713338890
transform 1 0 43229 0 1 37103
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_538
timestamp 1713338890
transform 1 0 47881 0 1 36989
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_539
timestamp 1713338890
transform 1 0 47749 0 1 37121
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_540
timestamp 1713338890
transform 1 0 52401 0 1 37001
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_541
timestamp 1713338890
transform 1 0 52269 0 1 37133
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_542
timestamp 1713338890
transform 1 0 43097 0 1 37235
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_543
timestamp 1713338890
transform 1 0 47617 0 1 37253
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_544
timestamp 1713338890
transform 1 0 52137 0 1 37265
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_545
timestamp 1713338890
transform 1 0 42965 0 1 37367
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_546
timestamp 1713338890
transform 1 0 42833 0 1 37499
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_547
timestamp 1713338890
transform 1 0 47485 0 1 37385
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_548
timestamp 1713338890
transform 1 0 52005 0 1 37397
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_549
timestamp 1713338890
transform 1 0 42701 0 1 37631
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_550
timestamp 1713338890
transform 1 0 47353 0 1 37517
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_551
timestamp 1713338890
transform 1 0 47221 0 1 37649
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_552
timestamp 1713338890
transform 1 0 51873 0 1 37529
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_553
timestamp 1713338890
transform 1 0 51741 0 1 37661
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_554
timestamp 1713338890
transform 1 0 42569 0 1 37763
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_555
timestamp 1713338890
transform 1 0 47089 0 1 37781
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_556
timestamp 1713338890
transform 1 0 51609 0 1 37793
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_557
timestamp 1713338890
transform 1 0 42437 0 1 37895
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_558
timestamp 1713338890
transform 1 0 46957 0 1 37913
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_559
timestamp 1713338890
transform 1 0 51477 0 1 37925
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_560
timestamp 1713338890
transform 1 0 42305 0 1 38027
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_561
timestamp 1713338890
transform 1 0 42173 0 1 38159
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_562
timestamp 1713338890
transform 1 0 46693 0 1 38177
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_563
timestamp 1713338890
transform 1 0 46825 0 1 38045
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_564
timestamp 1713338890
transform 1 0 51345 0 1 38057
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_565
timestamp 1713338890
transform 1 0 51213 0 1 38189
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_566
timestamp 1713338890
transform 1 0 42041 0 1 38291
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_567
timestamp 1713338890
transform 1 0 46561 0 1 38309
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_568
timestamp 1713338890
transform 1 0 51081 0 1 38321
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_569
timestamp 1713338890
transform 1 0 41909 0 1 38423
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_570
timestamp 1713338890
transform 1 0 46429 0 1 38441
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_571
timestamp 1713338890
transform 1 0 50949 0 1 38453
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_572
timestamp 1713338890
transform 1 0 41777 0 1 38555
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_573
timestamp 1713338890
transform 1 0 41645 0 1 38687
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_574
timestamp 1713338890
transform 1 0 46297 0 1 38573
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_575
timestamp 1713338890
transform 1 0 46165 0 1 38705
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_576
timestamp 1713338890
transform 1 0 50685 0 1 38717
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_577
timestamp 1713338890
transform 1 0 50817 0 1 38585
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_578
timestamp 1713338890
transform 1 0 41513 0 1 38819
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_579
timestamp 1713338890
transform 1 0 46033 0 1 38837
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_580
timestamp 1713338890
transform 1 0 50553 0 1 38849
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_581
timestamp 1713338890
transform 1 0 41381 0 1 38951
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_582
timestamp 1713338890
transform 1 0 45901 0 1 38969
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_583
timestamp 1713338890
transform 1 0 50421 0 1 38981
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_584
timestamp 1713338890
transform 1 0 41249 0 1 39083
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_585
timestamp 1713338890
transform 1 0 41117 0 1 39215
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_586
timestamp 1713338890
transform 1 0 45637 0 1 39233
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_587
timestamp 1713338890
transform 1 0 45769 0 1 39101
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_588
timestamp 1713338890
transform 1 0 50289 0 1 39113
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_589
timestamp 1713338890
transform 1 0 50157 0 1 39245
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_590
timestamp 1713338890
transform 1 0 40985 0 1 39347
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_591
timestamp 1713338890
transform 1 0 45505 0 1 39365
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_592
timestamp 1713338890
transform 1 0 50025 0 1 39377
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_593
timestamp 1713338890
transform 1 0 40853 0 1 39479
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_594
timestamp 1713338890
transform 1 0 45373 0 1 39497
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_595
timestamp 1713338890
transform 1 0 49893 0 1 39509
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_596
timestamp 1713338890
transform 1 0 54413 0 1 39530
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_597
timestamp 1713338890
transform 1 0 40721 0 1 39611
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_598
timestamp 1713338890
transform 1 0 40589 0 1 39743
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_599
timestamp 1713338890
transform 1 0 45241 0 1 39629
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_600
timestamp 1713338890
transform 1 0 45109 0 1 39761
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_601
timestamp 1713338890
transform 1 0 49761 0 1 39641
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_602
timestamp 1713338890
transform 1 0 49629 0 1 39773
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_603
timestamp 1713338890
transform 1 0 54281 0 1 39662
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_604
timestamp 1713338890
transform 1 0 54149 0 1 39794
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_605
timestamp 1713338890
transform 1 0 54017 0 1 39926
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_606
timestamp 1713338890
transform 1 0 44977 0 1 39893
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_607
timestamp 1713338890
transform 1 0 40457 0 1 39875
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_608
timestamp 1713338890
transform 1 0 49497 0 1 39905
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_609
timestamp 1713338890
transform 1 0 22113 0 1 40077
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_610
timestamp 1713338890
transform 1 0 26633 0 1 40093
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_611
timestamp 1713338890
transform 1 0 31153 0 1 40099
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_612
timestamp 1713338890
transform 1 0 31285 0 1 39967
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_613
timestamp 1713338890
transform 1 0 21981 0 1 40209
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_614
timestamp 1713338890
transform 1 0 21849 0 1 40341
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_615
timestamp 1713338890
transform 1 0 26501 0 1 40225
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_616
timestamp 1713338890
transform 1 0 26369 0 1 40357
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_617
timestamp 1713338890
transform 1 0 30889 0 1 40363
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_618
timestamp 1713338890
transform 1 0 31021 0 1 40231
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_619
timestamp 1713338890
transform 1 0 21717 0 1 40473
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_620
timestamp 1713338890
transform 1 0 26237 0 1 40489
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_621
timestamp 1713338890
transform 1 0 30757 0 1 40495
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_622
timestamp 1713338890
transform 1 0 21453 0 1 40737
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_623
timestamp 1713338890
transform 1 0 21585 0 1 40605
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_624
timestamp 1713338890
transform 1 0 26105 0 1 40621
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_625
timestamp 1713338890
transform 1 0 25973 0 1 40753
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_626
timestamp 1713338890
transform 1 0 30625 0 1 40627
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_627
timestamp 1713338890
transform 1 0 30493 0 1 40759
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_628
timestamp 1713338890
transform 1 0 21189 0 1 41001
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_629
timestamp 1713338890
transform 1 0 21321 0 1 40869
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_630
timestamp 1713338890
transform 1 0 25841 0 1 40885
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_631
timestamp 1713338890
transform 1 0 25709 0 1 41017
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_632
timestamp 1713338890
transform 1 0 30361 0 1 40891
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_633
timestamp 1713338890
transform 1 0 30229 0 1 41023
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_634
timestamp 1713338890
transform 1 0 21057 0 1 41133
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_635
timestamp 1713338890
transform 1 0 25577 0 1 41149
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_636
timestamp 1713338890
transform 1 0 30097 0 1 41155
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_637
timestamp 1713338890
transform 1 0 20793 0 1 41397
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_638
timestamp 1713338890
transform 1 0 20925 0 1 41265
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_639
timestamp 1713338890
transform 1 0 25445 0 1 41281
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_640
timestamp 1713338890
transform 1 0 25313 0 1 41413
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_641
timestamp 1713338890
transform 1 0 29965 0 1 41287
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_642
timestamp 1713338890
transform 1 0 29833 0 1 41419
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_643
timestamp 1713338890
transform 1 0 20661 0 1 41529
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_644
timestamp 1713338890
transform 1 0 20529 0 1 41661
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_645
timestamp 1713338890
transform 1 0 25181 0 1 41545
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_646
timestamp 1713338890
transform 1 0 29701 0 1 41551
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_647
timestamp 1713338890
transform 1 0 20397 0 1 41793
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_648
timestamp 1713338890
transform 1 0 25049 0 1 41677
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_649
timestamp 1713338890
transform 1 0 24917 0 1 41809
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_650
timestamp 1713338890
transform 1 0 29569 0 1 41683
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_651
timestamp 1713338890
transform 1 0 29437 0 1 41815
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_652
timestamp 1713338890
transform 1 0 38609 0 1 41723
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_653
timestamp 1713338890
transform 1 0 38477 0 1 41855
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_654
timestamp 1713338890
transform 1 0 20265 0 1 41925
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_655
timestamp 1713338890
transform 1 0 20133 0 1 42057
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_656
timestamp 1713338890
transform 1 0 24785 0 1 41941
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_657
timestamp 1713338890
transform 1 0 24653 0 1 42073
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_658
timestamp 1713338890
transform 1 0 29305 0 1 41947
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_659
timestamp 1713338890
transform 1 0 29173 0 1 42079
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_660
timestamp 1713338890
transform 1 0 38345 0 1 41987
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_661
timestamp 1713338890
transform 1 0 40325 0 1 40007
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_662
timestamp 1713338890
transform 1 0 44845 0 1 40025
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_663
timestamp 1713338890
transform 1 0 49365 0 1 40037
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_664
timestamp 1713338890
transform 1 0 53885 0 1 40058
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_665
timestamp 1713338890
transform 1 0 40193 0 1 40139
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_666
timestamp 1713338890
transform 1 0 40061 0 1 40271
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_667
timestamp 1713338890
transform 1 0 44713 0 1 40157
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_668
timestamp 1713338890
transform 1 0 44581 0 1 40289
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_669
timestamp 1713338890
transform 1 0 49233 0 1 40169
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_670
timestamp 1713338890
transform 1 0 49101 0 1 40301
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_671
timestamp 1713338890
transform 1 0 53753 0 1 40190
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_672
timestamp 1713338890
transform 1 0 39929 0 1 40403
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_673
timestamp 1713338890
transform 1 0 44449 0 1 40421
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_674
timestamp 1713338890
transform 1 0 48969 0 1 40433
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_675
timestamp 1713338890
transform 1 0 53621 0 1 40322
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_676
timestamp 1713338890
transform 1 0 53489 0 1 40454
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_677
timestamp 1713338890
transform 1 0 39797 0 1 40535
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_678
timestamp 1713338890
transform 1 0 44317 0 1 40553
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_679
timestamp 1713338890
transform 1 0 48837 0 1 40565
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_680
timestamp 1713338890
transform 1 0 53357 0 1 40586
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_681
timestamp 1713338890
transform 1 0 39665 0 1 40667
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_682
timestamp 1713338890
transform 1 0 39533 0 1 40799
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_683
timestamp 1713338890
transform 1 0 44185 0 1 40685
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_684
timestamp 1713338890
transform 1 0 44053 0 1 40817
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_685
timestamp 1713338890
transform 1 0 48705 0 1 40697
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_686
timestamp 1713338890
transform 1 0 48573 0 1 40829
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_687
timestamp 1713338890
transform 1 0 53225 0 1 40718
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_688
timestamp 1713338890
transform 1 0 39401 0 1 40931
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_689
timestamp 1713338890
transform 1 0 43921 0 1 40949
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_690
timestamp 1713338890
transform 1 0 48441 0 1 40961
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_691
timestamp 1713338890
transform 1 0 53093 0 1 40850
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_692
timestamp 1713338890
transform 1 0 52961 0 1 40982
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_693
timestamp 1713338890
transform 1 0 39269 0 1 41063
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_694
timestamp 1713338890
transform 1 0 43789 0 1 41081
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_695
timestamp 1713338890
transform 1 0 48309 0 1 41093
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_696
timestamp 1713338890
transform 1 0 52829 0 1 41114
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_697
timestamp 1713338890
transform 1 0 39005 0 1 41327
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_698
timestamp 1713338890
transform 1 0 39137 0 1 41195
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_699
timestamp 1713338890
transform 1 0 43657 0 1 41213
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_700
timestamp 1713338890
transform 1 0 43525 0 1 41345
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_701
timestamp 1713338890
transform 1 0 48177 0 1 41225
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_702
timestamp 1713338890
transform 1 0 48045 0 1 41357
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_703
timestamp 1713338890
transform 1 0 52697 0 1 41246
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_704
timestamp 1713338890
transform 1 0 38873 0 1 41459
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_705
timestamp 1713338890
transform 1 0 38741 0 1 41591
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_706
timestamp 1713338890
transform 1 0 43393 0 1 41477
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_707
timestamp 1713338890
transform 1 0 43261 0 1 41609
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_708
timestamp 1713338890
transform 1 0 47913 0 1 41489
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_709
timestamp 1713338890
transform 1 0 47781 0 1 41621
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_710
timestamp 1713338890
transform 1 0 52301 0 1 41642
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_711
timestamp 1713338890
transform 1 0 52565 0 1 41378
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_712
timestamp 1713338890
transform 1 0 52433 0 1 41510
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_713
timestamp 1713338890
transform 1 0 42865 0 1 42005
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_714
timestamp 1713338890
transform 1 0 43129 0 1 41741
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_715
timestamp 1713338890
transform 1 0 42997 0 1 41873
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_716
timestamp 1713338890
transform 1 0 47385 0 1 42017
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_717
timestamp 1713338890
transform 1 0 47649 0 1 41753
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_718
timestamp 1713338890
transform 1 0 47517 0 1 41885
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_719
timestamp 1713338890
transform 1 0 52169 0 1 41774
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_720
timestamp 1713338890
transform 1 0 52037 0 1 41906
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_721
timestamp 1713338890
transform 1 0 51905 0 1 42038
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_722
timestamp 1713338890
transform 1 0 19077 0 1 43113
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_723
timestamp 1713338890
transform 1 0 18945 0 1 43245
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_724
timestamp 1713338890
transform 1 0 18813 0 1 43377
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_725
timestamp 1713338890
transform 1 0 18417 0 1 43773
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_726
timestamp 1713338890
transform 1 0 18681 0 1 43509
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_727
timestamp 1713338890
transform 1 0 18549 0 1 43641
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_728
timestamp 1713338890
transform 1 0 18285 0 1 43905
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_729
timestamp 1713338890
transform 1 0 18153 0 1 44037
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_730
timestamp 1713338890
transform 1 0 18021 0 1 44169
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_731
timestamp 1713338890
transform 1 0 17889 0 1 44301
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_732
timestamp 1713338890
transform 1 0 17757 0 1 44433
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_733
timestamp 1713338890
transform 1 0 17625 0 1 44565
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_734
timestamp 1713338890
transform 1 0 17493 0 1 44697
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_735
timestamp 1713338890
transform 1 0 17361 0 1 44829
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_736
timestamp 1713338890
transform 1 0 17229 0 1 44961
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_737
timestamp 1713338890
transform 1 0 17097 0 1 45093
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_738
timestamp 1713338890
transform 1 0 16965 0 1 45225
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_739
timestamp 1713338890
transform 1 0 16833 0 1 45357
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_740
timestamp 1713338890
transform 1 0 16701 0 1 45489
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_741
timestamp 1713338890
transform 1 0 16569 0 1 45621
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_742
timestamp 1713338890
transform 1 0 16437 0 1 45753
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_743
timestamp 1713338890
transform 1 0 16305 0 1 45885
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_744
timestamp 1713338890
transform 1 0 16173 0 1 46017
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_745
timestamp 1713338890
transform 1 0 20001 0 1 42189
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_746
timestamp 1713338890
transform 1 0 19869 0 1 42321
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_747
timestamp 1713338890
transform 1 0 19737 0 1 42453
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_748
timestamp 1713338890
transform 1 0 19605 0 1 42585
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_749
timestamp 1713338890
transform 1 0 19473 0 1 42717
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_750
timestamp 1713338890
transform 1 0 19341 0 1 42849
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_751
timestamp 1713338890
transform 1 0 19209 0 1 42981
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_752
timestamp 1713338890
transform 1 0 23069 0 1 43657
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_753
timestamp 1713338890
transform 1 0 22937 0 1 43789
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_754
timestamp 1713338890
transform 1 0 22805 0 1 43921
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_755
timestamp 1713338890
transform 1 0 22673 0 1 44053
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_756
timestamp 1713338890
transform 1 0 22541 0 1 44185
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_757
timestamp 1713338890
transform 1 0 22277 0 1 44449
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_758
timestamp 1713338890
transform 1 0 22409 0 1 44317
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_759
timestamp 1713338890
transform 1 0 22145 0 1 44581
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_760
timestamp 1713338890
transform 1 0 22013 0 1 44713
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_761
timestamp 1713338890
transform 1 0 21881 0 1 44845
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_762
timestamp 1713338890
transform 1 0 21749 0 1 44977
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_763
timestamp 1713338890
transform 1 0 21485 0 1 45241
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_764
timestamp 1713338890
transform 1 0 21617 0 1 45109
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_765
timestamp 1713338890
transform 1 0 21353 0 1 45373
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_766
timestamp 1713338890
transform 1 0 21221 0 1 45505
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_767
timestamp 1713338890
transform 1 0 21089 0 1 45637
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_768
timestamp 1713338890
transform 1 0 20957 0 1 45769
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_769
timestamp 1713338890
transform 1 0 20825 0 1 45901
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_770
timestamp 1713338890
transform 1 0 20693 0 1 46033
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_771
timestamp 1713338890
transform 1 0 20561 0 1 46165
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_772
timestamp 1713338890
transform 1 0 20429 0 1 46297
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_773
timestamp 1713338890
transform 1 0 20297 0 1 46429
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_774
timestamp 1713338890
transform 1 0 20033 0 1 46693
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_775
timestamp 1713338890
transform 1 0 20165 0 1 46561
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_776
timestamp 1713338890
transform 1 0 19769 0 1 46957
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_777
timestamp 1713338890
transform 1 0 19901 0 1 46825
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_778
timestamp 1713338890
transform 1 0 19637 0 1 47089
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_779
timestamp 1713338890
transform 1 0 19505 0 1 47221
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_780
timestamp 1713338890
transform 1 0 19373 0 1 47353
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_781
timestamp 1713338890
transform 1 0 23101 0 1 48151
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_782
timestamp 1713338890
transform 1 0 22969 0 1 48283
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_783
timestamp 1713338890
transform 1 0 22837 0 1 48415
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_784
timestamp 1713338890
transform 1 0 22705 0 1 48547
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_785
timestamp 1713338890
transform 1 0 22573 0 1 48679
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_786
timestamp 1713338890
transform 1 0 24521 0 1 42205
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_787
timestamp 1713338890
transform 1 0 24389 0 1 42337
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_788
timestamp 1713338890
transform 1 0 24125 0 1 42601
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_789
timestamp 1713338890
transform 1 0 24257 0 1 42469
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_790
timestamp 1713338890
transform 1 0 23993 0 1 42733
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_791
timestamp 1713338890
transform 1 0 23861 0 1 42865
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_792
timestamp 1713338890
transform 1 0 23729 0 1 42997
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_793
timestamp 1713338890
transform 1 0 23597 0 1 43129
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_794
timestamp 1713338890
transform 1 0 23465 0 1 43261
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_795
timestamp 1713338890
transform 1 0 23333 0 1 43393
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_796
timestamp 1713338890
transform 1 0 23201 0 1 43525
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_797
timestamp 1713338890
transform 1 0 26665 0 1 44587
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_798
timestamp 1713338890
transform 1 0 26533 0 1 44719
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_799
timestamp 1713338890
transform 1 0 26401 0 1 44851
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_800
timestamp 1713338890
transform 1 0 26269 0 1 44983
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_801
timestamp 1713338890
transform 1 0 26137 0 1 45115
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_802
timestamp 1713338890
transform 1 0 26005 0 1 45247
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_803
timestamp 1713338890
transform 1 0 25873 0 1 45379
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_804
timestamp 1713338890
transform 1 0 25741 0 1 45511
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_805
timestamp 1713338890
transform 1 0 25345 0 1 45907
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_806
timestamp 1713338890
transform 1 0 25609 0 1 45643
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_807
timestamp 1713338890
transform 1 0 25477 0 1 45775
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_808
timestamp 1713338890
transform 1 0 25213 0 1 46039
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_809
timestamp 1713338890
transform 1 0 25081 0 1 46171
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_810
timestamp 1713338890
transform 1 0 24949 0 1 46303
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_811
timestamp 1713338890
transform 1 0 24817 0 1 46435
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_812
timestamp 1713338890
transform 1 0 24685 0 1 46567
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_813
timestamp 1713338890
transform 1 0 24553 0 1 46699
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_814
timestamp 1713338890
transform 1 0 24421 0 1 46831
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_815
timestamp 1713338890
transform 1 0 24289 0 1 46963
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_816
timestamp 1713338890
transform 1 0 24157 0 1 47095
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_817
timestamp 1713338890
transform 1 0 24025 0 1 47227
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_818
timestamp 1713338890
transform 1 0 23893 0 1 47359
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_819
timestamp 1713338890
transform 1 0 23761 0 1 47491
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_820
timestamp 1713338890
transform 1 0 23629 0 1 47623
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_821
timestamp 1713338890
transform 1 0 23497 0 1 47755
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_822
timestamp 1713338890
transform 1 0 23365 0 1 47887
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_823
timestamp 1713338890
transform 1 0 23233 0 1 48019
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_824
timestamp 1713338890
transform 1 0 29041 0 1 42211
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_825
timestamp 1713338890
transform 1 0 28909 0 1 42343
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_826
timestamp 1713338890
transform 1 0 28777 0 1 42475
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_827
timestamp 1713338890
transform 1 0 28645 0 1 42607
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_828
timestamp 1713338890
transform 1 0 28513 0 1 42739
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_829
timestamp 1713338890
transform 1 0 28381 0 1 42871
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_830
timestamp 1713338890
transform 1 0 28249 0 1 43003
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_831
timestamp 1713338890
transform 1 0 28117 0 1 43135
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_832
timestamp 1713338890
transform 1 0 27985 0 1 43267
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_833
timestamp 1713338890
transform 1 0 27853 0 1 43399
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_834
timestamp 1713338890
transform 1 0 27721 0 1 43531
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_835
timestamp 1713338890
transform 1 0 27589 0 1 43663
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_836
timestamp 1713338890
transform 1 0 27457 0 1 43795
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_837
timestamp 1713338890
transform 1 0 27325 0 1 43927
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_838
timestamp 1713338890
transform 1 0 27193 0 1 44059
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_839
timestamp 1713338890
transform 1 0 27061 0 1 44191
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_840
timestamp 1713338890
transform 1 0 26929 0 1 44323
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_841
timestamp 1713338890
transform 1 0 26797 0 1 44455
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_842
timestamp 1713338890
transform 1 0 30689 0 1 49643
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_843
timestamp 1713338890
transform 1 0 30557 0 1 49775
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_844
timestamp 1713338890
transform 1 0 30425 0 1 49907
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_845
timestamp 1713338890
transform 1 0 30293 0 1 50039
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_846
timestamp 1713338890
transform 1 0 30161 0 1 50171
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_847
timestamp 1713338890
transform 1 0 30029 0 1 50303
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_848
timestamp 1713338890
transform 1 0 29897 0 1 50435
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_849
timestamp 1713338890
transform 1 0 29765 0 1 50567
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_850
timestamp 1713338890
transform 1 0 29633 0 1 50699
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_851
timestamp 1713338890
transform 1 0 29501 0 1 50831
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_852
timestamp 1713338890
transform 1 0 29369 0 1 50963
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_853
timestamp 1713338890
transform 1 0 29237 0 1 51095
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_854
timestamp 1713338890
transform 1 0 29105 0 1 51227
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_855
timestamp 1713338890
transform 1 0 28973 0 1 51359
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_856
timestamp 1713338890
transform 1 0 34649 0 1 45683
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_857
timestamp 1713338890
transform 1 0 34517 0 1 45815
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_858
timestamp 1713338890
transform 1 0 34385 0 1 45947
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_859
timestamp 1713338890
transform 1 0 34253 0 1 46079
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_860
timestamp 1713338890
transform 1 0 34121 0 1 46211
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_861
timestamp 1713338890
transform 1 0 33989 0 1 46343
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_862
timestamp 1713338890
transform 1 0 33857 0 1 46475
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_863
timestamp 1713338890
transform 1 0 33725 0 1 46607
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_864
timestamp 1713338890
transform 1 0 33593 0 1 46739
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_865
timestamp 1713338890
transform 1 0 33461 0 1 46871
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_866
timestamp 1713338890
transform 1 0 33329 0 1 47003
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_867
timestamp 1713338890
transform 1 0 33197 0 1 47135
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_868
timestamp 1713338890
transform 1 0 33065 0 1 47267
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_869
timestamp 1713338890
transform 1 0 32933 0 1 47399
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_870
timestamp 1713338890
transform 1 0 32801 0 1 47531
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_871
timestamp 1713338890
transform 1 0 32669 0 1 47663
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_872
timestamp 1713338890
transform 1 0 32537 0 1 47795
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_873
timestamp 1713338890
transform 1 0 32405 0 1 47927
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_874
timestamp 1713338890
transform 1 0 32273 0 1 48059
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_875
timestamp 1713338890
transform 1 0 32141 0 1 48191
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_876
timestamp 1713338890
transform 1 0 32009 0 1 48323
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_877
timestamp 1713338890
transform 1 0 31877 0 1 48455
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_878
timestamp 1713338890
transform 1 0 31745 0 1 48587
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_879
timestamp 1713338890
transform 1 0 31613 0 1 48719
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_880
timestamp 1713338890
transform 1 0 31481 0 1 48851
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_881
timestamp 1713338890
transform 1 0 31349 0 1 48983
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_882
timestamp 1713338890
transform 1 0 31217 0 1 49115
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_883
timestamp 1713338890
transform 1 0 31085 0 1 49247
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_884
timestamp 1713338890
transform 1 0 30953 0 1 49379
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_885
timestamp 1713338890
transform 1 0 30821 0 1 49511
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_886
timestamp 1713338890
transform 1 0 34681 0 1 50189
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_887
timestamp 1713338890
transform 1 0 34549 0 1 50321
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_888
timestamp 1713338890
transform 1 0 34417 0 1 50453
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_889
timestamp 1713338890
transform 1 0 34285 0 1 50585
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_890
timestamp 1713338890
transform 1 0 34153 0 1 50717
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_891
timestamp 1713338890
transform 1 0 34021 0 1 50849
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_892
timestamp 1713338890
transform 1 0 33889 0 1 50981
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_893
timestamp 1713338890
transform 1 0 33757 0 1 51113
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_894
timestamp 1713338890
transform 1 0 33625 0 1 51245
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_895
timestamp 1713338890
transform 1 0 33493 0 1 51377
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_896
timestamp 1713338890
transform 1 0 33361 0 1 51509
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_897
timestamp 1713338890
transform 1 0 33229 0 1 51641
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_898
timestamp 1713338890
transform 1 0 33097 0 1 51773
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_899
timestamp 1713338890
transform 1 0 32965 0 1 51905
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_900
timestamp 1713338890
transform 1 0 32833 0 1 52037
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_901
timestamp 1713338890
transform 1 0 32701 0 1 52169
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_902
timestamp 1713338890
transform 1 0 32569 0 1 52301
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_903
timestamp 1713338890
transform 1 0 32437 0 1 52433
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_904
timestamp 1713338890
transform 1 0 32305 0 1 52565
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_905
timestamp 1713338890
transform 1 0 32173 0 1 52697
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_906
timestamp 1713338890
transform 1 0 38213 0 1 42119
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_907
timestamp 1713338890
transform 1 0 38081 0 1 42251
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_908
timestamp 1713338890
transform 1 0 37949 0 1 42383
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_909
timestamp 1713338890
transform 1 0 37817 0 1 42515
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_910
timestamp 1713338890
transform 1 0 37685 0 1 42647
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_911
timestamp 1713338890
transform 1 0 37553 0 1 42779
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_912
timestamp 1713338890
transform 1 0 37421 0 1 42911
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_913
timestamp 1713338890
transform 1 0 37289 0 1 43043
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_914
timestamp 1713338890
transform 1 0 37157 0 1 43175
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_915
timestamp 1713338890
transform 1 0 37025 0 1 43307
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_916
timestamp 1713338890
transform 1 0 36893 0 1 43439
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_917
timestamp 1713338890
transform 1 0 36761 0 1 43571
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_918
timestamp 1713338890
transform 1 0 36629 0 1 43703
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_919
timestamp 1713338890
transform 1 0 36497 0 1 43835
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_920
timestamp 1713338890
transform 1 0 36365 0 1 43967
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_921
timestamp 1713338890
transform 1 0 36101 0 1 44231
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_922
timestamp 1713338890
transform 1 0 36233 0 1 44099
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_923
timestamp 1713338890
transform 1 0 35969 0 1 44363
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_924
timestamp 1713338890
transform 1 0 35837 0 1 44495
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_925
timestamp 1713338890
transform 1 0 35705 0 1 44627
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_926
timestamp 1713338890
transform 1 0 35573 0 1 44759
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_927
timestamp 1713338890
transform 1 0 35441 0 1 44891
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_928
timestamp 1713338890
transform 1 0 35309 0 1 45023
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_929
timestamp 1713338890
transform 1 0 35177 0 1 45155
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_930
timestamp 1713338890
transform 1 0 35045 0 1 45287
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_931
timestamp 1713338890
transform 1 0 34913 0 1 45419
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_932
timestamp 1713338890
transform 1 0 34781 0 1 45551
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_933
timestamp 1713338890
transform 1 0 38113 0 1 46757
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_934
timestamp 1713338890
transform 1 0 37981 0 1 46889
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_935
timestamp 1713338890
transform 1 0 37849 0 1 47021
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_936
timestamp 1713338890
transform 1 0 37717 0 1 47153
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_937
timestamp 1713338890
transform 1 0 37585 0 1 47285
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_938
timestamp 1713338890
transform 1 0 37453 0 1 47417
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_939
timestamp 1713338890
transform 1 0 37321 0 1 47549
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_940
timestamp 1713338890
transform 1 0 37189 0 1 47681
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_941
timestamp 1713338890
transform 1 0 37057 0 1 47813
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_942
timestamp 1713338890
transform 1 0 36925 0 1 47945
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_943
timestamp 1713338890
transform 1 0 36793 0 1 48077
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_944
timestamp 1713338890
transform 1 0 36661 0 1 48209
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_945
timestamp 1713338890
transform 1 0 36529 0 1 48341
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_946
timestamp 1713338890
transform 1 0 36397 0 1 48473
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_947
timestamp 1713338890
transform 1 0 36265 0 1 48605
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_948
timestamp 1713338890
transform 1 0 36133 0 1 48737
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_949
timestamp 1713338890
transform 1 0 36001 0 1 48869
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_950
timestamp 1713338890
transform 1 0 35869 0 1 49001
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_951
timestamp 1713338890
transform 1 0 35737 0 1 49133
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_952
timestamp 1713338890
transform 1 0 35605 0 1 49265
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_953
timestamp 1713338890
transform 1 0 35473 0 1 49397
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_954
timestamp 1713338890
transform 1 0 35341 0 1 49529
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_955
timestamp 1713338890
transform 1 0 35209 0 1 49661
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_956
timestamp 1713338890
transform 1 0 35077 0 1 49793
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_957
timestamp 1713338890
transform 1 0 34945 0 1 49925
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_958
timestamp 1713338890
transform 1 0 34813 0 1 50057
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_959
timestamp 1713338890
transform 1 0 38145 0 1 51257
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_960
timestamp 1713338890
transform 1 0 38013 0 1 51389
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_961
timestamp 1713338890
transform 1 0 37881 0 1 51521
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_962
timestamp 1713338890
transform 1 0 37617 0 1 51785
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_963
timestamp 1713338890
transform 1 0 37749 0 1 51653
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_964
timestamp 1713338890
transform 1 0 37485 0 1 51917
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_965
timestamp 1713338890
transform 1 0 37353 0 1 52049
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_966
timestamp 1713338890
transform 1 0 37221 0 1 52181
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_967
timestamp 1713338890
transform 1 0 37089 0 1 52313
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_968
timestamp 1713338890
transform 1 0 36957 0 1 52445
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_969
timestamp 1713338890
transform 1 0 36825 0 1 52577
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_970
timestamp 1713338890
transform 1 0 36693 0 1 52709
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_971
timestamp 1713338890
transform 1 0 36561 0 1 52841
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_972
timestamp 1713338890
transform 1 0 36429 0 1 52973
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_973
timestamp 1713338890
transform 1 0 36297 0 1 53105
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_974
timestamp 1713338890
transform 1 0 36165 0 1 53237
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_975
timestamp 1713338890
transform 1 0 36033 0 1 53369
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_976
timestamp 1713338890
transform 1 0 35901 0 1 53501
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_977
timestamp 1713338890
transform 1 0 35769 0 1 53633
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_978
timestamp 1713338890
transform 1 0 35637 0 1 53765
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_979
timestamp 1713338890
transform 1 0 35505 0 1 53897
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_980
timestamp 1713338890
transform 1 0 35373 0 1 54029
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_981
timestamp 1713338890
transform 1 0 42205 0 1 42665
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_982
timestamp 1713338890
transform 1 0 42073 0 1 42797
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_983
timestamp 1713338890
transform 1 0 41941 0 1 42929
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_984
timestamp 1713338890
transform 1 0 41809 0 1 43061
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_985
timestamp 1713338890
transform 1 0 41677 0 1 43193
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_986
timestamp 1713338890
transform 1 0 41545 0 1 43325
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_987
timestamp 1713338890
transform 1 0 41413 0 1 43457
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_988
timestamp 1713338890
transform 1 0 41281 0 1 43589
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_989
timestamp 1713338890
transform 1 0 41149 0 1 43721
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_990
timestamp 1713338890
transform 1 0 41017 0 1 43853
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_991
timestamp 1713338890
transform 1 0 40885 0 1 43985
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_992
timestamp 1713338890
transform 1 0 40753 0 1 44117
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_993
timestamp 1713338890
transform 1 0 40621 0 1 44249
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_994
timestamp 1713338890
transform 1 0 40489 0 1 44381
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_995
timestamp 1713338890
transform 1 0 40357 0 1 44513
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_996
timestamp 1713338890
transform 1 0 40225 0 1 44645
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_997
timestamp 1713338890
transform 1 0 40093 0 1 44777
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_998
timestamp 1713338890
transform 1 0 39961 0 1 44909
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_999
timestamp 1713338890
transform 1 0 39829 0 1 45041
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1000
timestamp 1713338890
transform 1 0 39697 0 1 45173
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1001
timestamp 1713338890
transform 1 0 39565 0 1 45305
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1002
timestamp 1713338890
transform 1 0 39433 0 1 45437
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1003
timestamp 1713338890
transform 1 0 39301 0 1 45569
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1004
timestamp 1713338890
transform 1 0 39169 0 1 45701
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1005
timestamp 1713338890
transform 1 0 39037 0 1 45833
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1006
timestamp 1713338890
transform 1 0 38905 0 1 45965
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1007
timestamp 1713338890
transform 1 0 38773 0 1 46097
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1008
timestamp 1713338890
transform 1 0 38641 0 1 46229
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1009
timestamp 1713338890
transform 1 0 38509 0 1 46361
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1010
timestamp 1713338890
transform 1 0 38377 0 1 46493
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1011
timestamp 1713338890
transform 1 0 38245 0 1 46625
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1012
timestamp 1713338890
transform 1 0 42237 0 1 47165
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1013
timestamp 1713338890
transform 1 0 42105 0 1 47297
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1014
timestamp 1713338890
transform 1 0 41973 0 1 47429
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1015
timestamp 1713338890
transform 1 0 41841 0 1 47561
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1016
timestamp 1713338890
transform 1 0 41709 0 1 47693
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1017
timestamp 1713338890
transform 1 0 41577 0 1 47825
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1018
timestamp 1713338890
transform 1 0 41445 0 1 47957
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1019
timestamp 1713338890
transform 1 0 41313 0 1 48089
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1020
timestamp 1713338890
transform 1 0 41181 0 1 48221
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1021
timestamp 1713338890
transform 1 0 41049 0 1 48353
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1022
timestamp 1713338890
transform 1 0 40917 0 1 48485
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1023
timestamp 1713338890
transform 1 0 40785 0 1 48617
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1024
timestamp 1713338890
transform 1 0 40653 0 1 48749
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1025
timestamp 1713338890
transform 1 0 40521 0 1 48881
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1026
timestamp 1713338890
transform 1 0 40389 0 1 49013
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1027
timestamp 1713338890
transform 1 0 40257 0 1 49145
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1028
timestamp 1713338890
transform 1 0 40125 0 1 49277
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1029
timestamp 1713338890
transform 1 0 39993 0 1 49409
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1030
timestamp 1713338890
transform 1 0 39861 0 1 49541
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1031
timestamp 1713338890
transform 1 0 39729 0 1 49673
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1032
timestamp 1713338890
transform 1 0 39597 0 1 49805
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1033
timestamp 1713338890
transform 1 0 39465 0 1 49937
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1034
timestamp 1713338890
transform 1 0 39333 0 1 50069
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1035
timestamp 1713338890
transform 1 0 39201 0 1 50201
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1036
timestamp 1713338890
transform 1 0 39069 0 1 50333
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1037
timestamp 1713338890
transform 1 0 38937 0 1 50465
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1038
timestamp 1713338890
transform 1 0 38805 0 1 50597
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1039
timestamp 1713338890
transform 1 0 38673 0 1 50729
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1040
timestamp 1713338890
transform 1 0 38541 0 1 50861
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1041
timestamp 1713338890
transform 1 0 38409 0 1 50993
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1042
timestamp 1713338890
transform 1 0 38277 0 1 51125
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1043
timestamp 1713338890
transform 1 0 42269 0 1 51674
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1044
timestamp 1713338890
transform 1 0 42137 0 1 51806
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1045
timestamp 1713338890
transform 1 0 42005 0 1 51938
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1046
timestamp 1713338890
transform 1 0 41873 0 1 52070
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1047
timestamp 1713338890
transform 1 0 41741 0 1 52202
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1048
timestamp 1713338890
transform 1 0 41609 0 1 52334
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1049
timestamp 1713338890
transform 1 0 41477 0 1 52466
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1050
timestamp 1713338890
transform 1 0 41345 0 1 52598
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1051
timestamp 1713338890
transform 1 0 41213 0 1 52730
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1052
timestamp 1713338890
transform 1 0 41081 0 1 52862
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1053
timestamp 1713338890
transform 1 0 40949 0 1 52994
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1054
timestamp 1713338890
transform 1 0 40817 0 1 53126
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1055
timestamp 1713338890
transform 1 0 40685 0 1 53258
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1056
timestamp 1713338890
transform 1 0 40553 0 1 53390
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1057
timestamp 1713338890
transform 1 0 40421 0 1 53522
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1058
timestamp 1713338890
transform 1 0 40289 0 1 53654
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1059
timestamp 1713338890
transform 1 0 40157 0 1 53786
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1060
timestamp 1713338890
transform 1 0 40025 0 1 53918
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1061
timestamp 1713338890
transform 1 0 39893 0 1 54050
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1062
timestamp 1713338890
transform 1 0 39761 0 1 54182
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1063
timestamp 1713338890
transform 1 0 39629 0 1 54314
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1064
timestamp 1713338890
transform 1 0 39497 0 1 54446
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1065
timestamp 1713338890
transform 1 0 39365 0 1 54578
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1066
timestamp 1713338890
transform 1 0 39233 0 1 54710
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1067
timestamp 1713338890
transform 1 0 39101 0 1 54842
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1068
timestamp 1713338890
transform 1 0 38969 0 1 54974
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1069
timestamp 1713338890
transform 1 0 38837 0 1 55106
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1070
timestamp 1713338890
transform 1 0 38705 0 1 55238
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1071
timestamp 1713338890
transform 1 0 38573 0 1 55370
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1072
timestamp 1713338890
transform 1 0 42733 0 1 42137
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1073
timestamp 1713338890
transform 1 0 42601 0 1 42269
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1074
timestamp 1713338890
transform 1 0 42469 0 1 42401
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1075
timestamp 1713338890
transform 1 0 42337 0 1 42533
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1076
timestamp 1713338890
transform 1 0 46197 0 1 43205
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1077
timestamp 1713338890
transform 1 0 46065 0 1 43337
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1078
timestamp 1713338890
transform 1 0 45933 0 1 43469
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1079
timestamp 1713338890
transform 1 0 45801 0 1 43601
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1080
timestamp 1713338890
transform 1 0 45669 0 1 43733
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1081
timestamp 1713338890
transform 1 0 45537 0 1 43865
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1082
timestamp 1713338890
transform 1 0 45405 0 1 43997
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1083
timestamp 1713338890
transform 1 0 45273 0 1 44129
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1084
timestamp 1713338890
transform 1 0 45141 0 1 44261
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1085
timestamp 1713338890
transform 1 0 45009 0 1 44393
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1086
timestamp 1713338890
transform 1 0 44877 0 1 44525
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1087
timestamp 1713338890
transform 1 0 44745 0 1 44657
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1088
timestamp 1713338890
transform 1 0 44613 0 1 44789
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1089
timestamp 1713338890
transform 1 0 44481 0 1 44921
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1090
timestamp 1713338890
transform 1 0 44349 0 1 45053
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1091
timestamp 1713338890
transform 1 0 44217 0 1 45185
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1092
timestamp 1713338890
transform 1 0 44085 0 1 45317
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1093
timestamp 1713338890
transform 1 0 43953 0 1 45449
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1094
timestamp 1713338890
transform 1 0 43821 0 1 45581
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1095
timestamp 1713338890
transform 1 0 43689 0 1 45713
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1096
timestamp 1713338890
transform 1 0 43557 0 1 45845
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1097
timestamp 1713338890
transform 1 0 43425 0 1 45977
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1098
timestamp 1713338890
transform 1 0 43293 0 1 46109
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1099
timestamp 1713338890
transform 1 0 43161 0 1 46241
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1100
timestamp 1713338890
transform 1 0 43029 0 1 46373
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1101
timestamp 1713338890
transform 1 0 42897 0 1 46505
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1102
timestamp 1713338890
transform 1 0 42765 0 1 46637
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1103
timestamp 1713338890
transform 1 0 42633 0 1 46769
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1104
timestamp 1713338890
transform 1 0 42501 0 1 46901
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1105
timestamp 1713338890
transform 1 0 42369 0 1 47033
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1106
timestamp 1713338890
transform 1 0 46229 0 1 47714
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1107
timestamp 1713338890
transform 1 0 46097 0 1 47846
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1108
timestamp 1713338890
transform 1 0 45965 0 1 47978
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1109
timestamp 1713338890
transform 1 0 45833 0 1 48110
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1110
timestamp 1713338890
transform 1 0 45701 0 1 48242
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1111
timestamp 1713338890
transform 1 0 45569 0 1 48374
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1112
timestamp 1713338890
transform 1 0 45437 0 1 48506
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1113
timestamp 1713338890
transform 1 0 45305 0 1 48638
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1114
timestamp 1713338890
transform 1 0 45173 0 1 48770
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1115
timestamp 1713338890
transform 1 0 45041 0 1 48902
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1116
timestamp 1713338890
transform 1 0 44909 0 1 49034
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1117
timestamp 1713338890
transform 1 0 44777 0 1 49166
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1118
timestamp 1713338890
transform 1 0 44645 0 1 49298
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1119
timestamp 1713338890
transform 1 0 44513 0 1 49430
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1120
timestamp 1713338890
transform 1 0 44381 0 1 49562
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1121
timestamp 1713338890
transform 1 0 44249 0 1 49694
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1122
timestamp 1713338890
transform 1 0 44117 0 1 49826
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1123
timestamp 1713338890
transform 1 0 43985 0 1 49958
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1124
timestamp 1713338890
transform 1 0 43853 0 1 50090
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1125
timestamp 1713338890
transform 1 0 43721 0 1 50222
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1126
timestamp 1713338890
transform 1 0 43589 0 1 50354
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1127
timestamp 1713338890
transform 1 0 43457 0 1 50486
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1128
timestamp 1713338890
transform 1 0 43325 0 1 50618
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1129
timestamp 1713338890
transform 1 0 43193 0 1 50750
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1130
timestamp 1713338890
transform 1 0 43061 0 1 50882
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1131
timestamp 1713338890
transform 1 0 42929 0 1 51014
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1132
timestamp 1713338890
transform 1 0 42797 0 1 51146
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1133
timestamp 1713338890
transform 1 0 42665 0 1 51278
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1134
timestamp 1713338890
transform 1 0 42533 0 1 51410
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1135
timestamp 1713338890
transform 1 0 42401 0 1 51542
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1136
timestamp 1713338890
transform 1 0 47253 0 1 42149
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1137
timestamp 1713338890
transform 1 0 47121 0 1 42281
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1138
timestamp 1713338890
transform 1 0 46989 0 1 42413
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1139
timestamp 1713338890
transform 1 0 46857 0 1 42545
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1140
timestamp 1713338890
transform 1 0 46725 0 1 42677
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1141
timestamp 1713338890
transform 1 0 46593 0 1 42809
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1142
timestamp 1713338890
transform 1 0 46461 0 1 42941
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1143
timestamp 1713338890
transform 1 0 46329 0 1 43073
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1144
timestamp 1713338890
transform 1 0 49793 0 1 44150
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1145
timestamp 1713338890
transform 1 0 49661 0 1 44282
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1146
timestamp 1713338890
transform 1 0 49529 0 1 44414
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1147
timestamp 1713338890
transform 1 0 49397 0 1 44546
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1148
timestamp 1713338890
transform 1 0 49265 0 1 44678
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1149
timestamp 1713338890
transform 1 0 49133 0 1 44810
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1150
timestamp 1713338890
transform 1 0 49001 0 1 44942
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1151
timestamp 1713338890
transform 1 0 48869 0 1 45074
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1152
timestamp 1713338890
transform 1 0 48737 0 1 45206
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1153
timestamp 1713338890
transform 1 0 48605 0 1 45338
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1154
timestamp 1713338890
transform 1 0 48473 0 1 45470
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1155
timestamp 1713338890
transform 1 0 48341 0 1 45602
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1156
timestamp 1713338890
transform 1 0 48209 0 1 45734
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1157
timestamp 1713338890
transform 1 0 48077 0 1 45866
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1158
timestamp 1713338890
transform 1 0 47945 0 1 45998
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1159
timestamp 1713338890
transform 1 0 47813 0 1 46130
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1160
timestamp 1713338890
transform 1 0 47681 0 1 46262
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1161
timestamp 1713338890
transform 1 0 47549 0 1 46394
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1162
timestamp 1713338890
transform 1 0 47417 0 1 46526
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1163
timestamp 1713338890
transform 1 0 47285 0 1 46658
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1164
timestamp 1713338890
transform 1 0 47153 0 1 46790
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1165
timestamp 1713338890
transform 1 0 47021 0 1 46922
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1166
timestamp 1713338890
transform 1 0 46889 0 1 47054
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1167
timestamp 1713338890
transform 1 0 46757 0 1 47186
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1168
timestamp 1713338890
transform 1 0 46625 0 1 47318
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1169
timestamp 1713338890
transform 1 0 46493 0 1 47450
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1170
timestamp 1713338890
transform 1 0 46361 0 1 47582
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1171
timestamp 1713338890
transform 1 0 49725 0 1 53294
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1172
timestamp 1713338890
transform 1 0 49593 0 1 53426
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1173
timestamp 1713338890
transform 1 0 49461 0 1 53558
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1174
timestamp 1713338890
transform 1 0 49329 0 1 53690
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1175
timestamp 1713338890
transform 1 0 49197 0 1 53822
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1176
timestamp 1713338890
transform 1 0 49065 0 1 53954
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1177
timestamp 1713338890
transform 1 0 48933 0 1 54086
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1178
timestamp 1713338890
transform 1 0 48801 0 1 54218
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1179
timestamp 1713338890
transform 1 0 48669 0 1 54350
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1180
timestamp 1713338890
transform 1 0 48537 0 1 54482
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1181
timestamp 1713338890
transform 1 0 48405 0 1 54614
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1182
timestamp 1713338890
transform 1 0 48273 0 1 54746
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1183
timestamp 1713338890
transform 1 0 48141 0 1 54878
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1184
timestamp 1713338890
transform 1 0 48009 0 1 55010
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1185
timestamp 1713338890
transform 1 0 47877 0 1 55142
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1186
timestamp 1713338890
transform 1 0 47745 0 1 55274
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1187
timestamp 1713338890
transform 1 0 47613 0 1 55406
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1188
timestamp 1713338890
transform 1 0 47481 0 1 55538
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1189
timestamp 1713338890
transform 1 0 47349 0 1 55670
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1190
timestamp 1713338890
transform 1 0 47217 0 1 55802
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1191
timestamp 1713338890
transform 1 0 47085 0 1 55934
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1192
timestamp 1713338890
transform 1 0 46953 0 1 56066
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1193
timestamp 1713338890
transform 1 0 46821 0 1 56198
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1194
timestamp 1713338890
transform 1 0 46293 0 1 56726
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1195
timestamp 1713338890
transform 1 0 46161 0 1 56858
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1196
timestamp 1713338890
transform 1 0 46029 0 1 56990
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1197
timestamp 1713338890
transform 1 0 45897 0 1 57122
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1198
timestamp 1713338890
transform 1 0 45765 0 1 57254
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1199
timestamp 1713338890
transform 1 0 45633 0 1 57386
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1200
timestamp 1713338890
transform 1 0 45501 0 1 57518
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1201
timestamp 1713338890
transform 1 0 45369 0 1 57650
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1202
timestamp 1713338890
transform 1 0 45237 0 1 57782
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1203
timestamp 1713338890
transform 1 0 45105 0 1 57914
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1204
timestamp 1713338890
transform 1 0 44973 0 1 58046
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1205
timestamp 1713338890
transform 1 0 46689 0 1 56330
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1206
timestamp 1713338890
transform 1 0 46557 0 1 56462
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1207
timestamp 1713338890
transform 1 0 46425 0 1 56594
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1208
timestamp 1713338890
transform 1 0 49757 0 1 57828
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1209
timestamp 1713338890
transform 1 0 49625 0 1 57960
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1210
timestamp 1713338890
transform 1 0 49493 0 1 58092
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1211
timestamp 1713338890
transform 1 0 49361 0 1 58224
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1212
timestamp 1713338890
transform 1 0 49229 0 1 58356
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1213
timestamp 1713338890
transform 1 0 49097 0 1 58488
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1214
timestamp 1713338890
transform 1 0 48965 0 1 58620
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1215
timestamp 1713338890
transform 1 0 48833 0 1 58752
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1216
timestamp 1713338890
transform 1 0 48701 0 1 58884
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1217
timestamp 1713338890
transform 1 0 48569 0 1 59016
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1218
timestamp 1713338890
transform 1 0 48437 0 1 59148
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1219
timestamp 1713338890
transform 1 0 48305 0 1 59280
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1220
timestamp 1713338890
transform 1 0 48173 0 1 59412
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1221
timestamp 1713338890
transform 1 0 51773 0 1 42170
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1222
timestamp 1713338890
transform 1 0 51641 0 1 42302
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1223
timestamp 1713338890
transform 1 0 51509 0 1 42434
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1224
timestamp 1713338890
transform 1 0 51377 0 1 42566
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1225
timestamp 1713338890
transform 1 0 51245 0 1 42698
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1226
timestamp 1713338890
transform 1 0 51113 0 1 42830
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1227
timestamp 1713338890
transform 1 0 50981 0 1 42962
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1228
timestamp 1713338890
transform 1 0 50849 0 1 43094
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1229
timestamp 1713338890
transform 1 0 50717 0 1 43226
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1230
timestamp 1713338890
transform 1 0 50585 0 1 43358
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1231
timestamp 1713338890
transform 1 0 50453 0 1 43490
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1232
timestamp 1713338890
transform 1 0 50321 0 1 43622
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1233
timestamp 1713338890
transform 1 0 50189 0 1 43754
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1234
timestamp 1713338890
transform 1 0 50057 0 1 43886
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1235
timestamp 1713338890
transform 1 0 49925 0 1 44018
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1236
timestamp 1713338890
transform 1 0 53817 0 1 49202
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1237
timestamp 1713338890
transform 1 0 53685 0 1 49334
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1238
timestamp 1713338890
transform 1 0 53553 0 1 49466
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1239
timestamp 1713338890
transform 1 0 53421 0 1 49598
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1240
timestamp 1713338890
transform 1 0 53289 0 1 49730
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1241
timestamp 1713338890
transform 1 0 53157 0 1 49862
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1242
timestamp 1713338890
transform 1 0 53025 0 1 49994
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1243
timestamp 1713338890
transform 1 0 52893 0 1 50126
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1244
timestamp 1713338890
transform 1 0 52761 0 1 50258
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1245
timestamp 1713338890
transform 1 0 52629 0 1 50390
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1246
timestamp 1713338890
transform 1 0 52497 0 1 50522
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1247
timestamp 1713338890
transform 1 0 52365 0 1 50654
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1248
timestamp 1713338890
transform 1 0 52233 0 1 50786
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1249
timestamp 1713338890
transform 1 0 52101 0 1 50918
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1250
timestamp 1713338890
transform 1 0 51969 0 1 51050
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1251
timestamp 1713338890
transform 1 0 51837 0 1 51182
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1252
timestamp 1713338890
transform 1 0 51705 0 1 51314
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1253
timestamp 1713338890
transform 1 0 51573 0 1 51446
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1254
timestamp 1713338890
transform 1 0 51441 0 1 51578
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1255
timestamp 1713338890
transform 1 0 57117 0 1 45902
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1256
timestamp 1713338890
transform 1 0 56985 0 1 46034
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1257
timestamp 1713338890
transform 1 0 56853 0 1 46166
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1258
timestamp 1713338890
transform 1 0 56721 0 1 46298
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1259
timestamp 1713338890
transform 1 0 56589 0 1 46430
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1260
timestamp 1713338890
transform 1 0 56457 0 1 46562
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1261
timestamp 1713338890
transform 1 0 56325 0 1 46694
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1262
timestamp 1713338890
transform 1 0 56193 0 1 46826
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1263
timestamp 1713338890
transform 1 0 56061 0 1 46958
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1264
timestamp 1713338890
transform 1 0 55929 0 1 47090
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1265
timestamp 1713338890
transform 1 0 55797 0 1 47222
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1266
timestamp 1713338890
transform 1 0 55665 0 1 47354
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1267
timestamp 1713338890
transform 1 0 55533 0 1 47486
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1268
timestamp 1713338890
transform 1 0 55401 0 1 47618
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1269
timestamp 1713338890
transform 1 0 55269 0 1 47750
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1270
timestamp 1713338890
transform 1 0 55137 0 1 47882
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1271
timestamp 1713338890
transform 1 0 55005 0 1 48014
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1272
timestamp 1713338890
transform 1 0 54873 0 1 48146
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1273
timestamp 1713338890
transform 1 0 54741 0 1 48278
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1274
timestamp 1713338890
transform 1 0 54609 0 1 48410
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1275
timestamp 1713338890
transform 1 0 54477 0 1 48542
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1276
timestamp 1713338890
transform 1 0 54345 0 1 48674
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1277
timestamp 1713338890
transform 1 0 54213 0 1 48806
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1278
timestamp 1713338890
transform 1 0 54081 0 1 48938
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1279
timestamp 1713338890
transform 1 0 53949 0 1 49070
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1280
timestamp 1713338890
transform 1 0 57809 0 1 49776
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1281
timestamp 1713338890
transform 1 0 57677 0 1 49908
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1282
timestamp 1713338890
transform 1 0 57545 0 1 50040
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1283
timestamp 1713338890
transform 1 0 57413 0 1 50172
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1284
timestamp 1713338890
transform 1 0 57281 0 1 50304
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1285
timestamp 1713338890
transform 1 0 57149 0 1 50436
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1286
timestamp 1713338890
transform 1 0 57017 0 1 50568
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1287
timestamp 1713338890
transform 1 0 56885 0 1 50700
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1288
timestamp 1713338890
transform 1 0 56753 0 1 50832
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1289
timestamp 1713338890
transform 1 0 56621 0 1 50964
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1290
timestamp 1713338890
transform 1 0 56489 0 1 51096
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1291
timestamp 1713338890
transform 1 0 56357 0 1 51228
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1292
timestamp 1713338890
transform 1 0 56225 0 1 51360
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1293
timestamp 1713338890
transform 1 0 56093 0 1 51492
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1294
timestamp 1713338890
transform 1 0 55961 0 1 51624
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1295
timestamp 1713338890
transform 1 0 58469 0 1 49116
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1296
timestamp 1713338890
transform 1 0 58337 0 1 49248
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1297
timestamp 1713338890
transform 1 0 58205 0 1 49380
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1298
timestamp 1713338890
transform 1 0 58073 0 1 49512
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1299
timestamp 1713338890
transform 1 0 57941 0 1 49644
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1300
timestamp 1713338890
transform 1 0 51309 0 1 51710
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1301
timestamp 1713338890
transform 1 0 51177 0 1 51842
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1302
timestamp 1713338890
transform 1 0 51045 0 1 51974
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1303
timestamp 1713338890
transform 1 0 50913 0 1 52106
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1304
timestamp 1713338890
transform 1 0 50781 0 1 52238
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1305
timestamp 1713338890
transform 1 0 50649 0 1 52370
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1306
timestamp 1713338890
transform 1 0 50517 0 1 52502
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1307
timestamp 1713338890
transform 1 0 50385 0 1 52634
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1308
timestamp 1713338890
transform 1 0 50253 0 1 52766
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1309
timestamp 1713338890
transform 1 0 50121 0 1 52898
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1310
timestamp 1713338890
transform 1 0 49989 0 1 53030
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1311
timestamp 1713338890
transform 1 0 49857 0 1 53162
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1312
timestamp 1713338890
transform 1 0 53717 0 1 53868
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1313
timestamp 1713338890
transform 1 0 53585 0 1 54000
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1314
timestamp 1713338890
transform 1 0 53453 0 1 54132
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1315
timestamp 1713338890
transform 1 0 53321 0 1 54264
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1316
timestamp 1713338890
transform 1 0 53189 0 1 54396
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1317
timestamp 1713338890
transform 1 0 53057 0 1 54528
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1318
timestamp 1713338890
transform 1 0 52925 0 1 54660
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1319
timestamp 1713338890
transform 1 0 52793 0 1 54792
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1320
timestamp 1713338890
transform 1 0 52661 0 1 54924
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1321
timestamp 1713338890
transform 1 0 52529 0 1 55056
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1322
timestamp 1713338890
transform 1 0 52397 0 1 55188
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1323
timestamp 1713338890
transform 1 0 52265 0 1 55320
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1324
timestamp 1713338890
transform 1 0 52133 0 1 55452
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1325
timestamp 1713338890
transform 1 0 52001 0 1 55584
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1326
timestamp 1713338890
transform 1 0 51869 0 1 55716
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1327
timestamp 1713338890
transform 1 0 51737 0 1 55848
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1328
timestamp 1713338890
transform 1 0 51605 0 1 55980
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1329
timestamp 1713338890
transform 1 0 51473 0 1 56112
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1330
timestamp 1713338890
transform 1 0 51341 0 1 56244
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1331
timestamp 1713338890
transform 1 0 51209 0 1 56376
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1332
timestamp 1713338890
transform 1 0 51077 0 1 56508
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1333
timestamp 1713338890
transform 1 0 50945 0 1 56640
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1334
timestamp 1713338890
transform 1 0 50813 0 1 56772
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1335
timestamp 1713338890
transform 1 0 50681 0 1 56904
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1336
timestamp 1713338890
transform 1 0 50549 0 1 57036
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1337
timestamp 1713338890
transform 1 0 50417 0 1 57168
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1338
timestamp 1713338890
transform 1 0 50285 0 1 57300
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1339
timestamp 1713338890
transform 1 0 50153 0 1 57432
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1340
timestamp 1713338890
transform 1 0 50021 0 1 57564
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1341
timestamp 1713338890
transform 1 0 49889 0 1 57696
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1342
timestamp 1713338890
transform 1 0 55829 0 1 51756
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1343
timestamp 1713338890
transform 1 0 55697 0 1 51888
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1344
timestamp 1713338890
transform 1 0 55565 0 1 52020
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1345
timestamp 1713338890
transform 1 0 55433 0 1 52152
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1346
timestamp 1713338890
transform 1 0 55301 0 1 52284
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1347
timestamp 1713338890
transform 1 0 55169 0 1 52416
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1348
timestamp 1713338890
transform 1 0 55037 0 1 52548
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1349
timestamp 1713338890
transform 1 0 54905 0 1 52680
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1350
timestamp 1713338890
transform 1 0 54773 0 1 52812
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1351
timestamp 1713338890
transform 1 0 54641 0 1 52944
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1352
timestamp 1713338890
transform 1 0 54509 0 1 53076
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1353
timestamp 1713338890
transform 1 0 54377 0 1 53208
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1354
timestamp 1713338890
transform 1 0 54245 0 1 53340
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1355
timestamp 1713338890
transform 1 0 54113 0 1 53472
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1356
timestamp 1713338890
transform 1 0 53981 0 1 53604
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165219  M4_M3_CDNS_69033583165219_1357
timestamp 1713338890
transform 1 0 53849 0 1 53736
box -2018 -38 2018 38
use M4_M3_CDNS_69033583165220  M4_M3_CDNS_69033583165220_0
timestamp 1713338890
transform 1 0 14032 0 1 47259
box 28 -38 2876 38
use M4_M3_CDNS_69033583165220  M4_M3_CDNS_69033583165220_1
timestamp 1713338890
transform 1 0 17232 0 1 48595
box 28 -38 2876 38
use M4_M3_CDNS_69033583165220  M4_M3_CDNS_69033583165220_2
timestamp 1713338890
transform 1 0 20432 0 1 49921
box 28 -38 2876 38
use M4_M3_CDNS_69033583165220  M4_M3_CDNS_69033583165220_3
timestamp 1713338890
transform 1 0 26832 0 1 52601
box 28 -38 2876 38
use M4_M3_CDNS_69033583165220  M4_M3_CDNS_69033583165220_4
timestamp 1713338890
transform 1 0 30032 0 1 53939
box 28 -38 2876 38
use M4_M3_CDNS_69033583165220  M4_M3_CDNS_69033583165220_5
timestamp 1713338890
transform 1 0 33232 0 1 55271
box 28 -38 2876 38
use M4_M3_CDNS_69033583165220  M4_M3_CDNS_69033583165220_6
timestamp 1713338890
transform 1 0 36432 0 1 56612
box 28 -38 2876 38
use M4_M3_CDNS_69033583165220  M4_M3_CDNS_69033583165220_7
timestamp 1713338890
transform 1 0 42832 0 1 59288
box 28 -38 2876 38
use M4_M3_CDNS_69033583165220  M4_M3_CDNS_69033583165220_8
timestamp 1713338890
transform 1 0 46032 0 1 60655
box 28 -38 2876 38
use M4_M3_CDNS_69033583165221  M4_M3_CDNS_69033583165221_0
timestamp 1713338890
transform 1 0 47259 0 1 16816
box -3866 -38 38 38
use M4_M3_CDNS_69033583165221  M4_M3_CDNS_69033583165221_1
timestamp 1713338890
transform 1 0 48595 0 1 20016
box -3866 -38 38 38
use M4_M3_CDNS_69033583165221  M4_M3_CDNS_69033583165221_2
timestamp 1713338890
transform 1 0 49921 0 1 23216
box -3866 -38 38 38
use M4_M3_CDNS_69033583165221  M4_M3_CDNS_69033583165221_3
timestamp 1713338890
transform 1 0 52601 0 1 29616
box -3866 -38 38 38
use M4_M3_CDNS_69033583165221  M4_M3_CDNS_69033583165221_4
timestamp 1713338890
transform 1 0 53939 0 1 32816
box -3866 -38 38 38
use M4_M3_CDNS_69033583165221  M4_M3_CDNS_69033583165221_5
timestamp 1713338890
transform 1 0 55271 0 1 36016
box -3866 -38 38 38
use M4_M3_CDNS_69033583165221  M4_M3_CDNS_69033583165221_6
timestamp 1713338890
transform 1 0 56612 0 1 39216
box -3866 -38 38 38
use M4_M3_CDNS_69033583165221  M4_M3_CDNS_69033583165221_7
timestamp 1713338890
transform 1 0 59288 0 1 45616
box -3866 -38 38 38
use M4_M3_CDNS_69033583165222  M4_M3_CDNS_69033583165222_0
timestamp 1713338890
transform 1 0 47259 0 1 16684
box -3734 -38 38 38
use M4_M3_CDNS_69033583165222  M4_M3_CDNS_69033583165222_1
timestamp 1713338890
transform 1 0 48595 0 1 19884
box -3734 -38 38 38
use M4_M3_CDNS_69033583165222  M4_M3_CDNS_69033583165222_2
timestamp 1713338890
transform 1 0 49921 0 1 23084
box -3734 -38 38 38
use M4_M3_CDNS_69033583165222  M4_M3_CDNS_69033583165222_3
timestamp 1713338890
transform 1 0 52601 0 1 29484
box -3734 -38 38 38
use M4_M3_CDNS_69033583165222  M4_M3_CDNS_69033583165222_4
timestamp 1713338890
transform 1 0 53939 0 1 32684
box -3734 -38 38 38
use M4_M3_CDNS_69033583165222  M4_M3_CDNS_69033583165222_5
timestamp 1713338890
transform 1 0 55271 0 1 35884
box -3734 -38 38 38
use M4_M3_CDNS_69033583165222  M4_M3_CDNS_69033583165222_6
timestamp 1713338890
transform 1 0 56612 0 1 39084
box -3734 -38 38 38
use M4_M3_CDNS_69033583165222  M4_M3_CDNS_69033583165222_7
timestamp 1713338890
transform 1 0 59288 0 1 45484
box -3734 -38 38 38
use M4_M3_CDNS_69033583165223  M4_M3_CDNS_69033583165223_0
timestamp 1713338890
transform 1 0 47259 0 1 16552
box -3602 -38 38 38
use M4_M3_CDNS_69033583165223  M4_M3_CDNS_69033583165223_1
timestamp 1713338890
transform 1 0 48595 0 1 19752
box -3602 -38 38 38
use M4_M3_CDNS_69033583165223  M4_M3_CDNS_69033583165223_2
timestamp 1713338890
transform 1 0 49921 0 1 22952
box -3602 -38 38 38
use M4_M3_CDNS_69033583165223  M4_M3_CDNS_69033583165223_3
timestamp 1713338890
transform 1 0 52601 0 1 29352
box -3602 -38 38 38
use M4_M3_CDNS_69033583165223  M4_M3_CDNS_69033583165223_4
timestamp 1713338890
transform 1 0 53939 0 1 32552
box -3602 -38 38 38
use M4_M3_CDNS_69033583165223  M4_M3_CDNS_69033583165223_5
timestamp 1713338890
transform 1 0 55271 0 1 35752
box -3602 -38 38 38
use M4_M3_CDNS_69033583165223  M4_M3_CDNS_69033583165223_6
timestamp 1713338890
transform 1 0 56612 0 1 38952
box -3602 -38 38 38
use M4_M3_CDNS_69033583165223  M4_M3_CDNS_69033583165223_7
timestamp 1713338890
transform 1 0 59288 0 1 45352
box -3602 -38 38 38
use M4_M3_CDNS_69033583165224  M4_M3_CDNS_69033583165224_0
timestamp 1713338890
transform 1 0 47259 0 1 16420
box -3470 -38 38 38
use M4_M3_CDNS_69033583165224  M4_M3_CDNS_69033583165224_1
timestamp 1713338890
transform 1 0 48595 0 1 19620
box -3470 -38 38 38
use M4_M3_CDNS_69033583165224  M4_M3_CDNS_69033583165224_2
timestamp 1713338890
transform 1 0 49921 0 1 22820
box -3470 -38 38 38
use M4_M3_CDNS_69033583165224  M4_M3_CDNS_69033583165224_3
timestamp 1713338890
transform 1 0 52601 0 1 29220
box -3470 -38 38 38
use M4_M3_CDNS_69033583165224  M4_M3_CDNS_69033583165224_4
timestamp 1713338890
transform 1 0 53939 0 1 32420
box -3470 -38 38 38
use M4_M3_CDNS_69033583165224  M4_M3_CDNS_69033583165224_5
timestamp 1713338890
transform 1 0 55271 0 1 35620
box -3470 -38 38 38
use M4_M3_CDNS_69033583165224  M4_M3_CDNS_69033583165224_6
timestamp 1713338890
transform 1 0 56612 0 1 38820
box -3470 -38 38 38
use M4_M3_CDNS_69033583165224  M4_M3_CDNS_69033583165224_7
timestamp 1713338890
transform 1 0 59288 0 1 45220
box -3470 -38 38 38
use M4_M3_CDNS_69033583165225  M4_M3_CDNS_69033583165225_0
timestamp 1713338890
transform 1 0 47259 0 1 16948
box -3998 -38 38 38
use M4_M3_CDNS_69033583165225  M4_M3_CDNS_69033583165225_1
timestamp 1713338890
transform 1 0 48595 0 1 20148
box -3998 -38 38 38
use M4_M3_CDNS_69033583165225  M4_M3_CDNS_69033583165225_2
timestamp 1713338890
transform 1 0 49921 0 1 23348
box -3998 -38 38 38
use M4_M3_CDNS_69033583165225  M4_M3_CDNS_69033583165225_3
timestamp 1713338890
transform 1 0 52601 0 1 29748
box -3998 -38 38 38
use M4_M3_CDNS_69033583165225  M4_M3_CDNS_69033583165225_4
timestamp 1713338890
transform 1 0 53939 0 1 32948
box -3998 -38 38 38
use M4_M3_CDNS_69033583165225  M4_M3_CDNS_69033583165225_5
timestamp 1713338890
transform 1 0 55271 0 1 36148
box -3998 -38 38 38
use M4_M3_CDNS_69033583165225  M4_M3_CDNS_69033583165225_6
timestamp 1713338890
transform 1 0 56612 0 1 39348
box -3998 -38 38 38
use M4_M3_CDNS_69033583165225  M4_M3_CDNS_69033583165225_7
timestamp 1713338890
transform 1 0 59288 0 1 45748
box -3998 -38 38 38
use M4_M3_CDNS_69033583165226  M4_M3_CDNS_69033583165226_0
timestamp 1713338890
transform 1 0 53100 0 1 66854
box -698 -4130 698 4130
use M4_M3_CDNS_69033583165227  M4_M3_CDNS_69033583165227_0
timestamp 1713338890
transform 1 0 66854 0 1 53100
box -4130 -698 4130 698
use M4_M3_CDNS_69033583165228  M4_M3_CDNS_69033583165228_0
timestamp 1713338890
transform 1 0 23632 0 1 50203
box 28 -38 1688 38
use M4_M3_CDNS_69033583165228  M4_M3_CDNS_69033583165228_1
timestamp 1713338890
transform 1 0 25232 0 1 50872
box 28 -38 1688 38
use M4_M3_CDNS_69033583165228  M4_M3_CDNS_69033583165228_2
timestamp 1713338890
transform 1 0 39632 0 1 56890
box 28 -38 1688 38
use M4_M3_CDNS_69033583165228  M4_M3_CDNS_69033583165228_3
timestamp 1713338890
transform 1 0 41232 0 1 57562
box 28 -38 1688 38
use M4_M3_CDNS_69033583165228  M4_M3_CDNS_69033583165228_4
timestamp 1713338890
transform 1 0 49232 0 1 60927
box 28 -38 1688 38
use M4_M3_CDNS_69033583165228  M4_M3_CDNS_69033583165228_5
timestamp 1713338890
transform 1 0 50832 0 1 61591
box 28 -38 1688 38
use M4_M3_CDNS_69033583165228  M4_M3_CDNS_69033583165228_6
timestamp 1713338890
transform 1 0 52432 0 1 62259
box 28 -38 1688 38
use M4_M3_CDNS_69033583165228  M4_M3_CDNS_69033583165228_7
timestamp 1713338890
transform 1 0 54032 0 1 62925
box 28 -38 1688 38
use M4_M3_CDNS_69033583165228  M4_M3_CDNS_69033583165228_8
timestamp 1713338890
transform 1 0 55632 0 1 63588
box 28 -38 1688 38
use M4_M3_CDNS_69033583165228  M4_M3_CDNS_69033583165228_9
timestamp 1713338890
transform 1 0 57232 0 1 64251
box 28 -38 1688 38
use M4_M3_CDNS_69033583165228  M4_M3_CDNS_69033583165228_10
timestamp 1713338890
transform 1 0 58832 0 1 64918
box 28 -38 1688 38
use M4_M3_CDNS_69033583165228  M4_M3_CDNS_69033583165228_11
timestamp 1713338890
transform 1 0 60432 0 1 65583
box 28 -38 1688 38
use M4_M3_CDNS_69033583165228  M4_M3_CDNS_69033583165228_12
timestamp 1713338890
transform 1 0 62032 0 1 66246
box 28 -38 1688 38
use M4_M3_CDNS_69033583165228  M4_M3_CDNS_69033583165228_13
timestamp 1713338890
transform 1 0 63632 0 1 66918
box 28 -38 1688 38
use M4_M3_CDNS_69033583165228  M4_M3_CDNS_69033583165228_14
timestamp 1713338890
transform 1 0 65237 0 1 67576
box 28 -38 1688 38
use M4_M3_CDNS_69033583165229  M4_M3_CDNS_69033583165229_0
timestamp 1713338890
transform 1 0 23632 0 1 50335
box 28 -38 1556 38
use M4_M3_CDNS_69033583165229  M4_M3_CDNS_69033583165229_1
timestamp 1713338890
transform 1 0 25232 0 1 51004
box 28 -38 1556 38
use M4_M3_CDNS_69033583165229  M4_M3_CDNS_69033583165229_2
timestamp 1713338890
transform 1 0 39632 0 1 57022
box 28 -38 1556 38
use M4_M3_CDNS_69033583165229  M4_M3_CDNS_69033583165229_3
timestamp 1713338890
transform 1 0 41232 0 1 57694
box 28 -38 1556 38
use M4_M3_CDNS_69033583165229  M4_M3_CDNS_69033583165229_4
timestamp 1713338890
transform 1 0 49232 0 1 61059
box 28 -38 1556 38
use M4_M3_CDNS_69033583165229  M4_M3_CDNS_69033583165229_5
timestamp 1713338890
transform 1 0 50832 0 1 61723
box 28 -38 1556 38
use M4_M3_CDNS_69033583165229  M4_M3_CDNS_69033583165229_6
timestamp 1713338890
transform 1 0 52432 0 1 62391
box 28 -38 1556 38
use M4_M3_CDNS_69033583165229  M4_M3_CDNS_69033583165229_7
timestamp 1713338890
transform 1 0 54032 0 1 63057
box 28 -38 1556 38
use M4_M3_CDNS_69033583165229  M4_M3_CDNS_69033583165229_8
timestamp 1713338890
transform 1 0 55632 0 1 63720
box 28 -38 1556 38
use M4_M3_CDNS_69033583165229  M4_M3_CDNS_69033583165229_9
timestamp 1713338890
transform 1 0 57232 0 1 64383
box 28 -38 1556 38
use M4_M3_CDNS_69033583165229  M4_M3_CDNS_69033583165229_10
timestamp 1713338890
transform 1 0 58832 0 1 65050
box 28 -38 1556 38
use M4_M3_CDNS_69033583165229  M4_M3_CDNS_69033583165229_11
timestamp 1713338890
transform 1 0 60432 0 1 65715
box 28 -38 1556 38
use M4_M3_CDNS_69033583165229  M4_M3_CDNS_69033583165229_12
timestamp 1713338890
transform 1 0 62032 0 1 66378
box 28 -38 1556 38
use M4_M3_CDNS_69033583165229  M4_M3_CDNS_69033583165229_13
timestamp 1713338890
transform 1 0 63632 0 1 67050
box 28 -38 1556 38
use M4_M3_CDNS_69033583165229  M4_M3_CDNS_69033583165229_14
timestamp 1713338890
transform 1 0 65237 0 1 67708
box 28 -38 1556 38
use M4_M3_CDNS_69033583165229  M4_M3_CDNS_69033583165229_15
timestamp 1713338890
transform 1 0 66832 0 1 68318
box 28 -38 1556 38
use M4_M3_CDNS_69033583165230  M4_M3_CDNS_69033583165230_0
timestamp 1713338890
transform 1 0 23632 0 1 50467
box 28 -38 1424 38
use M4_M3_CDNS_69033583165230  M4_M3_CDNS_69033583165230_1
timestamp 1713338890
transform 1 0 25232 0 1 51136
box 28 -38 1424 38
use M4_M3_CDNS_69033583165230  M4_M3_CDNS_69033583165230_2
timestamp 1713338890
transform 1 0 39632 0 1 57154
box 28 -38 1424 38
use M4_M3_CDNS_69033583165230  M4_M3_CDNS_69033583165230_3
timestamp 1713338890
transform 1 0 41232 0 1 57826
box 28 -38 1424 38
use M4_M3_CDNS_69033583165230  M4_M3_CDNS_69033583165230_4
timestamp 1713338890
transform 1 0 49232 0 1 61191
box 28 -38 1424 38
use M4_M3_CDNS_69033583165230  M4_M3_CDNS_69033583165230_5
timestamp 1713338890
transform 1 0 50832 0 1 61855
box 28 -38 1424 38
use M4_M3_CDNS_69033583165230  M4_M3_CDNS_69033583165230_6
timestamp 1713338890
transform 1 0 52432 0 1 62523
box 28 -38 1424 38
use M4_M3_CDNS_69033583165230  M4_M3_CDNS_69033583165230_7
timestamp 1713338890
transform 1 0 54032 0 1 63189
box 28 -38 1424 38
use M4_M3_CDNS_69033583165230  M4_M3_CDNS_69033583165230_8
timestamp 1713338890
transform 1 0 55632 0 1 63852
box 28 -38 1424 38
use M4_M3_CDNS_69033583165230  M4_M3_CDNS_69033583165230_9
timestamp 1713338890
transform 1 0 57232 0 1 64515
box 28 -38 1424 38
use M4_M3_CDNS_69033583165230  M4_M3_CDNS_69033583165230_10
timestamp 1713338890
transform 1 0 58832 0 1 65182
box 28 -38 1424 38
use M4_M3_CDNS_69033583165230  M4_M3_CDNS_69033583165230_11
timestamp 1713338890
transform 1 0 60432 0 1 65847
box 28 -38 1424 38
use M4_M3_CDNS_69033583165230  M4_M3_CDNS_69033583165230_12
timestamp 1713338890
transform 1 0 62032 0 1 66510
box 28 -38 1424 38
use M4_M3_CDNS_69033583165230  M4_M3_CDNS_69033583165230_13
timestamp 1713338890
transform 1 0 63632 0 1 67182
box 28 -38 1424 38
use M4_M3_CDNS_69033583165230  M4_M3_CDNS_69033583165230_14
timestamp 1713338890
transform 1 0 65237 0 1 67840
box 28 -38 1424 38
use M4_M3_CDNS_69033583165230  M4_M3_CDNS_69033583165230_15
timestamp 1713338890
transform 1 0 66832 0 1 68509
box 28 -38 1424 38
use M4_M3_CDNS_69033583165231  M4_M3_CDNS_69033583165231_0
timestamp 1713338890
transform 1 0 23632 0 1 50599
box 28 -38 1292 38
use M4_M3_CDNS_69033583165231  M4_M3_CDNS_69033583165231_1
timestamp 1713338890
transform 1 0 25232 0 1 51268
box 28 -38 1292 38
use M4_M3_CDNS_69033583165231  M4_M3_CDNS_69033583165231_2
timestamp 1713338890
transform 1 0 39632 0 1 57286
box 28 -38 1292 38
use M4_M3_CDNS_69033583165231  M4_M3_CDNS_69033583165231_3
timestamp 1713338890
transform 1 0 41232 0 1 57958
box 28 -38 1292 38
use M4_M3_CDNS_69033583165231  M4_M3_CDNS_69033583165231_4
timestamp 1713338890
transform 1 0 50832 0 1 61987
box 28 -38 1292 38
use M4_M3_CDNS_69033583165231  M4_M3_CDNS_69033583165231_5
timestamp 1713338890
transform 1 0 49232 0 1 61323
box 28 -38 1292 38
use M4_M3_CDNS_69033583165231  M4_M3_CDNS_69033583165231_6
timestamp 1713338890
transform 1 0 52432 0 1 62655
box 28 -38 1292 38
use M4_M3_CDNS_69033583165231  M4_M3_CDNS_69033583165231_7
timestamp 1713338890
transform 1 0 54032 0 1 63321
box 28 -38 1292 38
use M4_M3_CDNS_69033583165231  M4_M3_CDNS_69033583165231_8
timestamp 1713338890
transform 1 0 55632 0 1 63984
box 28 -38 1292 38
use M4_M3_CDNS_69033583165231  M4_M3_CDNS_69033583165231_9
timestamp 1713338890
transform 1 0 57232 0 1 64647
box 28 -38 1292 38
use M4_M3_CDNS_69033583165231  M4_M3_CDNS_69033583165231_10
timestamp 1713338890
transform 1 0 58832 0 1 65314
box 28 -38 1292 38
use M4_M3_CDNS_69033583165231  M4_M3_CDNS_69033583165231_11
timestamp 1713338890
transform 1 0 60432 0 1 65979
box 28 -38 1292 38
use M4_M3_CDNS_69033583165231  M4_M3_CDNS_69033583165231_12
timestamp 1713338890
transform 1 0 62032 0 1 66642
box 28 -38 1292 38
use M4_M3_CDNS_69033583165231  M4_M3_CDNS_69033583165231_13
timestamp 1713338890
transform 1 0 63632 0 1 67314
box 28 -38 1292 38
use M4_M3_CDNS_69033583165231  M4_M3_CDNS_69033583165231_14
timestamp 1713338890
transform 1 0 65237 0 1 67972
box 28 -38 1292 38
use M4_M3_CDNS_69033583165231  M4_M3_CDNS_69033583165231_15
timestamp 1713338890
transform 1 0 66832 0 1 68641
box 28 -38 1292 38
use M4_M3_CDNS_69033583165232  M4_M3_CDNS_69033583165232_0
timestamp 1713338890
transform 1 0 47259 0 1 14572
box -1622 -38 38 38
use M4_M3_CDNS_69033583165232  M4_M3_CDNS_69033583165232_1
timestamp 1713338890
transform 1 0 48595 0 1 17772
box -1622 -38 38 38
use M4_M3_CDNS_69033583165232  M4_M3_CDNS_69033583165232_2
timestamp 1713338890
transform 1 0 49921 0 1 20972
box -1622 -38 38 38
use M4_M3_CDNS_69033583165232  M4_M3_CDNS_69033583165232_3
timestamp 1713338890
transform 1 0 50599 0 1 24816
box -1622 -38 38 38
use M4_M3_CDNS_69033583165232  M4_M3_CDNS_69033583165232_4
timestamp 1713338890
transform 1 0 51268 0 1 26416
box -1622 -38 38 38
use M4_M3_CDNS_69033583165232  M4_M3_CDNS_69033583165232_5
timestamp 1713338890
transform 1 0 52601 0 1 27372
box -1622 -38 38 38
use M4_M3_CDNS_69033583165232  M4_M3_CDNS_69033583165232_6
timestamp 1713338890
transform 1 0 53939 0 1 30572
box -1622 -38 38 38
use M4_M3_CDNS_69033583165232  M4_M3_CDNS_69033583165232_7
timestamp 1713338890
transform 1 0 55271 0 1 33772
box -1622 -38 38 38
use M4_M3_CDNS_69033583165232  M4_M3_CDNS_69033583165232_8
timestamp 1713338890
transform 1 0 56612 0 1 36972
box -1622 -38 38 38
use M4_M3_CDNS_69033583165232  M4_M3_CDNS_69033583165232_9
timestamp 1713338890
transform 1 0 57286 0 1 40816
box -1622 -38 38 38
use M4_M3_CDNS_69033583165232  M4_M3_CDNS_69033583165232_10
timestamp 1713338890
transform 1 0 57958 0 1 42416
box -1622 -38 38 38
use M4_M3_CDNS_69033583165232  M4_M3_CDNS_69033583165232_11
timestamp 1713338890
transform 1 0 59288 0 1 43372
box -1622 -38 38 38
use M4_M3_CDNS_69033583165232  M4_M3_CDNS_69033583165232_12
timestamp 1713338890
transform 1 0 63321 0 1 55216
box -1622 -38 38 38
use M4_M3_CDNS_69033583165232  M4_M3_CDNS_69033583165232_13
timestamp 1713338890
transform 1 0 63984 0 1 56816
box -1622 -38 38 38
use M4_M3_CDNS_69033583165232  M4_M3_CDNS_69033583165232_14
timestamp 1713338890
transform 1 0 64647 0 1 58416
box -1622 -38 38 38
use M4_M3_CDNS_69033583165232  M4_M3_CDNS_69033583165232_15
timestamp 1713338890
transform 1 0 65314 0 1 60016
box -1622 -38 38 38
use M4_M3_CDNS_69033583165232  M4_M3_CDNS_69033583165232_16
timestamp 1713338890
transform 1 0 65978 0 1 61617
box -1622 -38 38 38
use M4_M3_CDNS_69033583165232  M4_M3_CDNS_69033583165232_17
timestamp 1713338890
transform 1 0 66642 0 1 63216
box -1622 -38 38 38
use M4_M3_CDNS_69033583165232  M4_M3_CDNS_69033583165232_18
timestamp 1713338890
transform 1 0 67314 0 1 64816
box -1622 -38 38 38
use M4_M3_CDNS_69033583165232  M4_M3_CDNS_69033583165232_19
timestamp 1713338890
transform 1 0 67977 0 1 66416
box -1622 -38 38 38
use M4_M3_CDNS_69033583165232  M4_M3_CDNS_69033583165232_20
timestamp 1713338890
transform 1 0 68641 0 1 68016
box -1622 -38 38 38
use M4_M3_CDNS_69033583165233  M4_M3_CDNS_69033583165233_0
timestamp 1713338890
transform 1 0 47259 0 1 14308
box -1358 -38 38 38
use M4_M3_CDNS_69033583165233  M4_M3_CDNS_69033583165233_1
timestamp 1713338890
transform 1 0 48595 0 1 17508
box -1358 -38 38 38
use M4_M3_CDNS_69033583165233  M4_M3_CDNS_69033583165233_2
timestamp 1713338890
transform 1 0 49921 0 1 20708
box -1358 -38 38 38
use M4_M3_CDNS_69033583165233  M4_M3_CDNS_69033583165233_3
timestamp 1713338890
transform 1 0 50599 0 1 24552
box -1358 -38 38 38
use M4_M3_CDNS_69033583165233  M4_M3_CDNS_69033583165233_4
timestamp 1713338890
transform 1 0 51268 0 1 26152
box -1358 -38 38 38
use M4_M3_CDNS_69033583165233  M4_M3_CDNS_69033583165233_5
timestamp 1713338890
transform 1 0 52601 0 1 27108
box -1358 -38 38 38
use M4_M3_CDNS_69033583165233  M4_M3_CDNS_69033583165233_6
timestamp 1713338890
transform 1 0 53939 0 1 30308
box -1358 -38 38 38
use M4_M3_CDNS_69033583165233  M4_M3_CDNS_69033583165233_7
timestamp 1713338890
transform 1 0 55271 0 1 33508
box -1358 -38 38 38
use M4_M3_CDNS_69033583165233  M4_M3_CDNS_69033583165233_8
timestamp 1713338890
transform 1 0 56612 0 1 36708
box -1358 -38 38 38
use M4_M3_CDNS_69033583165233  M4_M3_CDNS_69033583165233_9
timestamp 1713338890
transform 1 0 57286 0 1 40552
box -1358 -38 38 38
use M4_M3_CDNS_69033583165233  M4_M3_CDNS_69033583165233_10
timestamp 1713338890
transform 1 0 57958 0 1 42152
box -1358 -38 38 38
use M4_M3_CDNS_69033583165233  M4_M3_CDNS_69033583165233_11
timestamp 1713338890
transform 1 0 59288 0 1 43108
box -1358 -38 38 38
use M4_M3_CDNS_69033583165233  M4_M3_CDNS_69033583165233_12
timestamp 1713338890
transform 1 0 63321 0 1 54952
box -1358 -38 38 38
use M4_M3_CDNS_69033583165233  M4_M3_CDNS_69033583165233_13
timestamp 1713338890
transform 1 0 63984 0 1 56552
box -1358 -38 38 38
use M4_M3_CDNS_69033583165233  M4_M3_CDNS_69033583165233_14
timestamp 1713338890
transform 1 0 64647 0 1 58152
box -1358 -38 38 38
use M4_M3_CDNS_69033583165233  M4_M3_CDNS_69033583165233_15
timestamp 1713338890
transform 1 0 65314 0 1 59752
box -1358 -38 38 38
use M4_M3_CDNS_69033583165233  M4_M3_CDNS_69033583165233_16
timestamp 1713338890
transform 1 0 65978 0 1 61353
box -1358 -38 38 38
use M4_M3_CDNS_69033583165233  M4_M3_CDNS_69033583165233_17
timestamp 1713338890
transform 1 0 66642 0 1 62952
box -1358 -38 38 38
use M4_M3_CDNS_69033583165233  M4_M3_CDNS_69033583165233_18
timestamp 1713338890
transform 1 0 67314 0 1 64552
box -1358 -38 38 38
use M4_M3_CDNS_69033583165233  M4_M3_CDNS_69033583165233_19
timestamp 1713338890
transform 1 0 67977 0 1 66152
box -1358 -38 38 38
use M4_M3_CDNS_69033583165233  M4_M3_CDNS_69033583165233_20
timestamp 1713338890
transform 1 0 68641 0 1 67752
box -1358 -38 38 38
use M4_M3_CDNS_69033583165234  M4_M3_CDNS_69033583165234_0
timestamp 1713338890
transform 1 0 50599 0 1 23760
box -566 -38 38 38
use M4_M3_CDNS_69033583165234  M4_M3_CDNS_69033583165234_1
timestamp 1713338890
transform 1 0 51268 0 1 25360
box -566 -38 38 38
use M4_M3_CDNS_69033583165234  M4_M3_CDNS_69033583165234_2
timestamp 1713338890
transform 1 0 57286 0 1 39760
box -566 -38 38 38
use M4_M3_CDNS_69033583165234  M4_M3_CDNS_69033583165234_3
timestamp 1713338890
transform 1 0 57958 0 1 41360
box -566 -38 38 38
use M4_M3_CDNS_69033583165234  M4_M3_CDNS_69033583165234_4
timestamp 1713338890
transform 1 0 63321 0 1 54160
box -566 -38 38 38
use M4_M3_CDNS_69033583165234  M4_M3_CDNS_69033583165234_5
timestamp 1713338890
transform 1 0 63984 0 1 55760
box -566 -38 38 38
use M4_M3_CDNS_69033583165234  M4_M3_CDNS_69033583165234_6
timestamp 1713338890
transform 1 0 64647 0 1 57360
box -566 -38 38 38
use M4_M3_CDNS_69033583165234  M4_M3_CDNS_69033583165234_7
timestamp 1713338890
transform 1 0 65314 0 1 58960
box -566 -38 38 38
use M4_M3_CDNS_69033583165234  M4_M3_CDNS_69033583165234_8
timestamp 1713338890
transform 1 0 65978 0 1 60561
box -566 -38 38 38
use M4_M3_CDNS_69033583165234  M4_M3_CDNS_69033583165234_9
timestamp 1713338890
transform 1 0 66642 0 1 62160
box -566 -38 38 38
use M4_M3_CDNS_69033583165234  M4_M3_CDNS_69033583165234_10
timestamp 1713338890
transform 1 0 67314 0 1 63760
box -566 -38 38 38
use M4_M3_CDNS_69033583165234  M4_M3_CDNS_69033583165234_11
timestamp 1713338890
transform 1 0 67977 0 1 65360
box -566 -38 38 38
use M4_M3_CDNS_69033583165234  M4_M3_CDNS_69033583165234_12
timestamp 1713338890
transform 1 0 68641 0 1 66960
box -566 -38 38 38
use M4_M3_CDNS_69033583165235  M4_M3_CDNS_69033583165235_0
timestamp 1713338890
transform 1 0 47259 0 1 14440
box -1490 -38 38 38
use M4_M3_CDNS_69033583165235  M4_M3_CDNS_69033583165235_1
timestamp 1713338890
transform 1 0 48595 0 1 17640
box -1490 -38 38 38
use M4_M3_CDNS_69033583165235  M4_M3_CDNS_69033583165235_2
timestamp 1713338890
transform 1 0 49921 0 1 20840
box -1490 -38 38 38
use M4_M3_CDNS_69033583165235  M4_M3_CDNS_69033583165235_3
timestamp 1713338890
transform 1 0 50599 0 1 24684
box -1490 -38 38 38
use M4_M3_CDNS_69033583165235  M4_M3_CDNS_69033583165235_4
timestamp 1713338890
transform 1 0 51268 0 1 26284
box -1490 -38 38 38
use M4_M3_CDNS_69033583165235  M4_M3_CDNS_69033583165235_5
timestamp 1713338890
transform 1 0 52601 0 1 27240
box -1490 -38 38 38
use M4_M3_CDNS_69033583165235  M4_M3_CDNS_69033583165235_6
timestamp 1713338890
transform 1 0 53939 0 1 30440
box -1490 -38 38 38
use M4_M3_CDNS_69033583165235  M4_M3_CDNS_69033583165235_7
timestamp 1713338890
transform 1 0 55271 0 1 33640
box -1490 -38 38 38
use M4_M3_CDNS_69033583165235  M4_M3_CDNS_69033583165235_8
timestamp 1713338890
transform 1 0 56612 0 1 36840
box -1490 -38 38 38
use M4_M3_CDNS_69033583165235  M4_M3_CDNS_69033583165235_9
timestamp 1713338890
transform 1 0 57286 0 1 40684
box -1490 -38 38 38
use M4_M3_CDNS_69033583165235  M4_M3_CDNS_69033583165235_10
timestamp 1713338890
transform 1 0 57958 0 1 42284
box -1490 -38 38 38
use M4_M3_CDNS_69033583165235  M4_M3_CDNS_69033583165235_11
timestamp 1713338890
transform 1 0 59288 0 1 43240
box -1490 -38 38 38
use M4_M3_CDNS_69033583165235  M4_M3_CDNS_69033583165235_12
timestamp 1713338890
transform 1 0 63321 0 1 55084
box -1490 -38 38 38
use M4_M3_CDNS_69033583165235  M4_M3_CDNS_69033583165235_13
timestamp 1713338890
transform 1 0 63984 0 1 56684
box -1490 -38 38 38
use M4_M3_CDNS_69033583165235  M4_M3_CDNS_69033583165235_14
timestamp 1713338890
transform 1 0 64647 0 1 58284
box -1490 -38 38 38
use M4_M3_CDNS_69033583165235  M4_M3_CDNS_69033583165235_15
timestamp 1713338890
transform 1 0 65314 0 1 59884
box -1490 -38 38 38
use M4_M3_CDNS_69033583165235  M4_M3_CDNS_69033583165235_16
timestamp 1713338890
transform 1 0 65978 0 1 61485
box -1490 -38 38 38
use M4_M3_CDNS_69033583165235  M4_M3_CDNS_69033583165235_17
timestamp 1713338890
transform 1 0 66642 0 1 63084
box -1490 -38 38 38
use M4_M3_CDNS_69033583165235  M4_M3_CDNS_69033583165235_18
timestamp 1713338890
transform 1 0 67314 0 1 64684
box -1490 -38 38 38
use M4_M3_CDNS_69033583165235  M4_M3_CDNS_69033583165235_19
timestamp 1713338890
transform 1 0 67977 0 1 66284
box -1490 -38 38 38
use M4_M3_CDNS_69033583165235  M4_M3_CDNS_69033583165235_20
timestamp 1713338890
transform 1 0 68641 0 1 67884
box -1490 -38 38 38
use M4_M3_CDNS_69033583165236  M4_M3_CDNS_69033583165236_0
timestamp 1713338890
transform 1 0 47259 0 1 14176
box -1226 -38 38 38
use M4_M3_CDNS_69033583165236  M4_M3_CDNS_69033583165236_1
timestamp 1713338890
transform 1 0 48595 0 1 17376
box -1226 -38 38 38
use M4_M3_CDNS_69033583165236  M4_M3_CDNS_69033583165236_2
timestamp 1713338890
transform 1 0 49921 0 1 20576
box -1226 -38 38 38
use M4_M3_CDNS_69033583165236  M4_M3_CDNS_69033583165236_3
timestamp 1713338890
transform 1 0 50599 0 1 24420
box -1226 -38 38 38
use M4_M3_CDNS_69033583165236  M4_M3_CDNS_69033583165236_4
timestamp 1713338890
transform 1 0 51268 0 1 26020
box -1226 -38 38 38
use M4_M3_CDNS_69033583165236  M4_M3_CDNS_69033583165236_5
timestamp 1713338890
transform 1 0 52601 0 1 26976
box -1226 -38 38 38
use M4_M3_CDNS_69033583165236  M4_M3_CDNS_69033583165236_6
timestamp 1713338890
transform 1 0 53939 0 1 30176
box -1226 -38 38 38
use M4_M3_CDNS_69033583165236  M4_M3_CDNS_69033583165236_7
timestamp 1713338890
transform 1 0 55271 0 1 33376
box -1226 -38 38 38
use M4_M3_CDNS_69033583165236  M4_M3_CDNS_69033583165236_8
timestamp 1713338890
transform 1 0 56612 0 1 36576
box -1226 -38 38 38
use M4_M3_CDNS_69033583165236  M4_M3_CDNS_69033583165236_9
timestamp 1713338890
transform 1 0 57286 0 1 40420
box -1226 -38 38 38
use M4_M3_CDNS_69033583165236  M4_M3_CDNS_69033583165236_10
timestamp 1713338890
transform 1 0 57958 0 1 42020
box -1226 -38 38 38
use M4_M3_CDNS_69033583165236  M4_M3_CDNS_69033583165236_11
timestamp 1713338890
transform 1 0 59288 0 1 42976
box -1226 -38 38 38
use M4_M3_CDNS_69033583165236  M4_M3_CDNS_69033583165236_12
timestamp 1713338890
transform 1 0 63321 0 1 54820
box -1226 -38 38 38
use M4_M3_CDNS_69033583165236  M4_M3_CDNS_69033583165236_13
timestamp 1713338890
transform 1 0 63984 0 1 56420
box -1226 -38 38 38
use M4_M3_CDNS_69033583165236  M4_M3_CDNS_69033583165236_14
timestamp 1713338890
transform 1 0 64647 0 1 58020
box -1226 -38 38 38
use M4_M3_CDNS_69033583165236  M4_M3_CDNS_69033583165236_15
timestamp 1713338890
transform 1 0 65314 0 1 59620
box -1226 -38 38 38
use M4_M3_CDNS_69033583165236  M4_M3_CDNS_69033583165236_16
timestamp 1713338890
transform 1 0 65978 0 1 61221
box -1226 -38 38 38
use M4_M3_CDNS_69033583165236  M4_M3_CDNS_69033583165236_17
timestamp 1713338890
transform 1 0 66642 0 1 62820
box -1226 -38 38 38
use M4_M3_CDNS_69033583165236  M4_M3_CDNS_69033583165236_18
timestamp 1713338890
transform 1 0 67314 0 1 64420
box -1226 -38 38 38
use M4_M3_CDNS_69033583165236  M4_M3_CDNS_69033583165236_19
timestamp 1713338890
transform 1 0 67977 0 1 66020
box -1226 -38 38 38
use M4_M3_CDNS_69033583165236  M4_M3_CDNS_69033583165236_20
timestamp 1713338890
transform 1 0 68641 0 1 67620
box -1226 -38 38 38
use M4_M3_CDNS_69033583165237  M4_M3_CDNS_69033583165237_0
timestamp 1713338890
transform 1 0 47259 0 1 14704
box -1754 -38 38 38
use M4_M3_CDNS_69033583165237  M4_M3_CDNS_69033583165237_1
timestamp 1713338890
transform 1 0 48595 0 1 17904
box -1754 -38 38 38
use M4_M3_CDNS_69033583165237  M4_M3_CDNS_69033583165237_2
timestamp 1713338890
transform 1 0 49921 0 1 21104
box -1754 -38 38 38
use M4_M3_CDNS_69033583165237  M4_M3_CDNS_69033583165237_3
timestamp 1713338890
transform 1 0 50599 0 1 24948
box -1754 -38 38 38
use M4_M3_CDNS_69033583165237  M4_M3_CDNS_69033583165237_4
timestamp 1713338890
transform 1 0 51268 0 1 26548
box -1754 -38 38 38
use M4_M3_CDNS_69033583165237  M4_M3_CDNS_69033583165237_5
timestamp 1713338890
transform 1 0 52601 0 1 27504
box -1754 -38 38 38
use M4_M3_CDNS_69033583165237  M4_M3_CDNS_69033583165237_6
timestamp 1713338890
transform 1 0 53939 0 1 30704
box -1754 -38 38 38
use M4_M3_CDNS_69033583165237  M4_M3_CDNS_69033583165237_7
timestamp 1713338890
transform 1 0 55271 0 1 33904
box -1754 -38 38 38
use M4_M3_CDNS_69033583165237  M4_M3_CDNS_69033583165237_8
timestamp 1713338890
transform 1 0 56612 0 1 37104
box -1754 -38 38 38
use M4_M3_CDNS_69033583165237  M4_M3_CDNS_69033583165237_9
timestamp 1713338890
transform 1 0 57286 0 1 40948
box -1754 -38 38 38
use M4_M3_CDNS_69033583165237  M4_M3_CDNS_69033583165237_10
timestamp 1713338890
transform 1 0 57958 0 1 42548
box -1754 -38 38 38
use M4_M3_CDNS_69033583165237  M4_M3_CDNS_69033583165237_11
timestamp 1713338890
transform 1 0 59288 0 1 43504
box -1754 -38 38 38
use M4_M3_CDNS_69033583165237  M4_M3_CDNS_69033583165237_12
timestamp 1713338890
transform 1 0 63321 0 1 55348
box -1754 -38 38 38
use M4_M3_CDNS_69033583165237  M4_M3_CDNS_69033583165237_13
timestamp 1713338890
transform 1 0 63984 0 1 56948
box -1754 -38 38 38
use M4_M3_CDNS_69033583165237  M4_M3_CDNS_69033583165237_14
timestamp 1713338890
transform 1 0 64647 0 1 58548
box -1754 -38 38 38
use M4_M3_CDNS_69033583165237  M4_M3_CDNS_69033583165237_15
timestamp 1713338890
transform 1 0 65314 0 1 60148
box -1754 -38 38 38
use M4_M3_CDNS_69033583165237  M4_M3_CDNS_69033583165237_16
timestamp 1713338890
transform 1 0 65978 0 1 61749
box -1754 -38 38 38
use M4_M3_CDNS_69033583165237  M4_M3_CDNS_69033583165237_17
timestamp 1713338890
transform 1 0 66642 0 1 63348
box -1754 -38 38 38
use M4_M3_CDNS_69033583165237  M4_M3_CDNS_69033583165237_18
timestamp 1713338890
transform 1 0 67314 0 1 64948
box -1754 -38 38 38
use M4_M3_CDNS_69033583165237  M4_M3_CDNS_69033583165237_19
timestamp 1713338890
transform 1 0 67977 0 1 66548
box -1754 -38 38 38
use M4_M3_CDNS_69033583165237  M4_M3_CDNS_69033583165237_20
timestamp 1713338890
transform 1 0 68641 0 1 68148
box -1754 -38 38 38
use M4_M3_CDNS_69033583165238  M4_M3_CDNS_69033583165238_0
timestamp 1713338890
transform 1 0 60655 0 1 46308
box -1292 -38 -28 38
use M4_M3_CDNS_69033583165238  M4_M3_CDNS_69033583165238_1
timestamp 1713338890
transform 1 0 61323 0 1 50152
box -1292 -38 -28 38
use M4_M3_CDNS_69033583165238  M4_M3_CDNS_69033583165238_2
timestamp 1713338890
transform 1 0 61987 0 1 51752
box -1292 -38 -28 38
use M4_M3_CDNS_69033583165238  M4_M3_CDNS_69033583165238_3
timestamp 1713338890
transform 1 0 62655 0 1 53352
box -1292 -38 -28 38
use M4_M3_CDNS_69033583165239  M4_M3_CDNS_69033583165239_0
timestamp 1713338890
transform 1 0 60655 0 1 46440
box -1424 -38 -28 38
use M4_M3_CDNS_69033583165239  M4_M3_CDNS_69033583165239_1
timestamp 1713338890
transform 1 0 61323 0 1 50284
box -1424 -38 -28 38
use M4_M3_CDNS_69033583165239  M4_M3_CDNS_69033583165239_2
timestamp 1713338890
transform 1 0 61987 0 1 51884
box -1424 -38 -28 38
use M4_M3_CDNS_69033583165239  M4_M3_CDNS_69033583165239_3
timestamp 1713338890
transform 1 0 62655 0 1 53484
box -1424 -38 -28 38
use M4_M3_CDNS_69033583165240  M4_M3_CDNS_69033583165240_0
timestamp 1713338890
transform 1 0 60655 0 1 46704
box -1688 -38 -28 38
use M4_M3_CDNS_69033583165240  M4_M3_CDNS_69033583165240_1
timestamp 1713338890
transform 1 0 61323 0 1 50548
box -1688 -38 -28 38
use M4_M3_CDNS_69033583165240  M4_M3_CDNS_69033583165240_2
timestamp 1713338890
transform 1 0 61987 0 1 52148
box -1688 -38 -28 38
use M4_M3_CDNS_69033583165240  M4_M3_CDNS_69033583165240_3
timestamp 1713338890
transform 1 0 62655 0 1 53748
box -1688 -38 -28 38
use M4_M3_CDNS_69033583165241  M4_M3_CDNS_69033583165241_0
timestamp 1713338890
transform 1 0 60655 0 1 46572
box -1556 -38 -28 38
use M4_M3_CDNS_69033583165241  M4_M3_CDNS_69033583165241_1
timestamp 1713338890
transform 1 0 61323 0 1 50416
box -1556 -38 -28 38
use M4_M3_CDNS_69033583165241  M4_M3_CDNS_69033583165241_2
timestamp 1713338890
transform 1 0 61987 0 1 52016
box -1556 -38 -28 38
use M4_M3_CDNS_69033583165241  M4_M3_CDNS_69033583165241_3
timestamp 1713338890
transform 1 0 62655 0 1 53616
box -1556 -38 -28 38
use M4_M3_CDNS_69033583165242  M4_M3_CDNS_69033583165242_0
timestamp 1713338890
transform 1 0 62700 0 1 68847
box -698 -2084 698 2084
use M4_M3_CDNS_69033583165243  M4_M3_CDNS_69033583165243_0
timestamp 1713338890
transform 1 0 68847 0 1 62700
box -2084 -698 2084 698
use M4_M3_CDNS_69033583165244  M4_M3_CDNS_69033583165244_0
timestamp 1713338890
transform 1 0 50599 0 1 24288
box -1094 -38 38 38
use M4_M3_CDNS_69033583165244  M4_M3_CDNS_69033583165244_1
timestamp 1713338890
transform 1 0 51268 0 1 25888
box -1094 -38 38 38
use M4_M3_CDNS_69033583165244  M4_M3_CDNS_69033583165244_2
timestamp 1713338890
transform 1 0 57286 0 1 40288
box -1094 -38 38 38
use M4_M3_CDNS_69033583165244  M4_M3_CDNS_69033583165244_3
timestamp 1713338890
transform 1 0 57958 0 1 41888
box -1094 -38 38 38
use M4_M3_CDNS_69033583165244  M4_M3_CDNS_69033583165244_4
timestamp 1713338890
transform 1 0 63321 0 1 54688
box -1094 -38 38 38
use M4_M3_CDNS_69033583165244  M4_M3_CDNS_69033583165244_5
timestamp 1713338890
transform 1 0 63984 0 1 56288
box -1094 -38 38 38
use M4_M3_CDNS_69033583165244  M4_M3_CDNS_69033583165244_6
timestamp 1713338890
transform 1 0 64647 0 1 57888
box -1094 -38 38 38
use M4_M3_CDNS_69033583165244  M4_M3_CDNS_69033583165244_7
timestamp 1713338890
transform 1 0 65314 0 1 59488
box -1094 -38 38 38
use M4_M3_CDNS_69033583165244  M4_M3_CDNS_69033583165244_8
timestamp 1713338890
transform 1 0 65978 0 1 61089
box -1094 -38 38 38
use M4_M3_CDNS_69033583165244  M4_M3_CDNS_69033583165244_9
timestamp 1713338890
transform 1 0 66642 0 1 62688
box -1094 -38 38 38
use M4_M3_CDNS_69033583165244  M4_M3_CDNS_69033583165244_10
timestamp 1713338890
transform 1 0 67314 0 1 64288
box -1094 -38 38 38
use M4_M3_CDNS_69033583165244  M4_M3_CDNS_69033583165244_11
timestamp 1713338890
transform 1 0 67977 0 1 65888
box -1094 -38 38 38
use M4_M3_CDNS_69033583165244  M4_M3_CDNS_69033583165244_12
timestamp 1713338890
transform 1 0 68641 0 1 67488
box -1094 -38 38 38
use M4_M3_CDNS_69033583165245  M4_M3_CDNS_69033583165245_0
timestamp 1713338890
transform 1 0 50599 0 1 24024
box -830 -38 38 38
use M4_M3_CDNS_69033583165245  M4_M3_CDNS_69033583165245_1
timestamp 1713338890
transform 1 0 51268 0 1 25624
box -830 -38 38 38
use M4_M3_CDNS_69033583165245  M4_M3_CDNS_69033583165245_2
timestamp 1713338890
transform 1 0 57286 0 1 40024
box -830 -38 38 38
use M4_M3_CDNS_69033583165245  M4_M3_CDNS_69033583165245_3
timestamp 1713338890
transform 1 0 57958 0 1 41624
box -830 -38 38 38
use M4_M3_CDNS_69033583165245  M4_M3_CDNS_69033583165245_4
timestamp 1713338890
transform 1 0 63321 0 1 54424
box -830 -38 38 38
use M4_M3_CDNS_69033583165245  M4_M3_CDNS_69033583165245_5
timestamp 1713338890
transform 1 0 63984 0 1 56024
box -830 -38 38 38
use M4_M3_CDNS_69033583165245  M4_M3_CDNS_69033583165245_6
timestamp 1713338890
transform 1 0 64647 0 1 57624
box -830 -38 38 38
use M4_M3_CDNS_69033583165245  M4_M3_CDNS_69033583165245_7
timestamp 1713338890
transform 1 0 65314 0 1 59224
box -830 -38 38 38
use M4_M3_CDNS_69033583165245  M4_M3_CDNS_69033583165245_8
timestamp 1713338890
transform 1 0 65978 0 1 60825
box -830 -38 38 38
use M4_M3_CDNS_69033583165245  M4_M3_CDNS_69033583165245_9
timestamp 1713338890
transform 1 0 66642 0 1 62424
box -830 -38 38 38
use M4_M3_CDNS_69033583165245  M4_M3_CDNS_69033583165245_10
timestamp 1713338890
transform 1 0 67314 0 1 64024
box -830 -38 38 38
use M4_M3_CDNS_69033583165245  M4_M3_CDNS_69033583165245_11
timestamp 1713338890
transform 1 0 67977 0 1 65624
box -830 -38 38 38
use M4_M3_CDNS_69033583165245  M4_M3_CDNS_69033583165245_12
timestamp 1713338890
transform 1 0 68641 0 1 67224
box -830 -38 38 38
use M4_M3_CDNS_69033583165246  M4_M3_CDNS_69033583165246_0
timestamp 1713338890
transform 1 0 50599 0 1 23892
box -698 -38 38 38
use M4_M3_CDNS_69033583165246  M4_M3_CDNS_69033583165246_1
timestamp 1713338890
transform 1 0 51268 0 1 25492
box -698 -38 38 38
use M4_M3_CDNS_69033583165246  M4_M3_CDNS_69033583165246_2
timestamp 1713338890
transform 1 0 57286 0 1 39892
box -698 -38 38 38
use M4_M3_CDNS_69033583165246  M4_M3_CDNS_69033583165246_3
timestamp 1713338890
transform 1 0 57958 0 1 41492
box -698 -38 38 38
use M4_M3_CDNS_69033583165246  M4_M3_CDNS_69033583165246_4
timestamp 1713338890
transform 1 0 63321 0 1 54292
box -698 -38 38 38
use M4_M3_CDNS_69033583165246  M4_M3_CDNS_69033583165246_5
timestamp 1713338890
transform 1 0 63984 0 1 55892
box -698 -38 38 38
use M4_M3_CDNS_69033583165246  M4_M3_CDNS_69033583165246_6
timestamp 1713338890
transform 1 0 64647 0 1 57492
box -698 -38 38 38
use M4_M3_CDNS_69033583165246  M4_M3_CDNS_69033583165246_7
timestamp 1713338890
transform 1 0 65314 0 1 59092
box -698 -38 38 38
use M4_M3_CDNS_69033583165246  M4_M3_CDNS_69033583165246_8
timestamp 1713338890
transform 1 0 65978 0 1 60693
box -698 -38 38 38
use M4_M3_CDNS_69033583165246  M4_M3_CDNS_69033583165246_9
timestamp 1713338890
transform 1 0 66642 0 1 62292
box -698 -38 38 38
use M4_M3_CDNS_69033583165246  M4_M3_CDNS_69033583165246_10
timestamp 1713338890
transform 1 0 67314 0 1 63892
box -698 -38 38 38
use M4_M3_CDNS_69033583165246  M4_M3_CDNS_69033583165246_11
timestamp 1713338890
transform 1 0 67977 0 1 65492
box -698 -38 38 38
use M4_M3_CDNS_69033583165246  M4_M3_CDNS_69033583165246_12
timestamp 1713338890
transform 1 0 68641 0 1 67092
box -698 -38 38 38
use M4_M3_CDNS_69033583165247  M4_M3_CDNS_69033583165247_0
timestamp 1713338890
transform 1 0 50599 0 1 24156
box -962 -38 38 38
use M4_M3_CDNS_69033583165247  M4_M3_CDNS_69033583165247_1
timestamp 1713338890
transform 1 0 51268 0 1 25756
box -962 -38 38 38
use M4_M3_CDNS_69033583165247  M4_M3_CDNS_69033583165247_2
timestamp 1713338890
transform 1 0 57286 0 1 40156
box -962 -38 38 38
use M4_M3_CDNS_69033583165247  M4_M3_CDNS_69033583165247_3
timestamp 1713338890
transform 1 0 57958 0 1 41756
box -962 -38 38 38
use M4_M3_CDNS_69033583165247  M4_M3_CDNS_69033583165247_4
timestamp 1713338890
transform 1 0 63321 0 1 54556
box -962 -38 38 38
use M4_M3_CDNS_69033583165247  M4_M3_CDNS_69033583165247_5
timestamp 1713338890
transform 1 0 63984 0 1 56156
box -962 -38 38 38
use M4_M3_CDNS_69033583165247  M4_M3_CDNS_69033583165247_6
timestamp 1713338890
transform 1 0 64647 0 1 57756
box -962 -38 38 38
use M4_M3_CDNS_69033583165247  M4_M3_CDNS_69033583165247_7
timestamp 1713338890
transform 1 0 65314 0 1 59356
box -962 -38 38 38
use M4_M3_CDNS_69033583165247  M4_M3_CDNS_69033583165247_8
timestamp 1713338890
transform 1 0 65978 0 1 60957
box -962 -38 38 38
use M4_M3_CDNS_69033583165247  M4_M3_CDNS_69033583165247_9
timestamp 1713338890
transform 1 0 66642 0 1 62556
box -962 -38 38 38
use M4_M3_CDNS_69033583165247  M4_M3_CDNS_69033583165247_10
timestamp 1713338890
transform 1 0 67314 0 1 64156
box -962 -38 38 38
use M4_M3_CDNS_69033583165247  M4_M3_CDNS_69033583165247_11
timestamp 1713338890
transform 1 0 67977 0 1 65756
box -962 -38 38 38
use M4_M3_CDNS_69033583165247  M4_M3_CDNS_69033583165247_12
timestamp 1713338890
transform 1 0 68641 0 1 67356
box -962 -38 38 38
use M4_M3_CDNS_69033583165248  M4_M3_CDNS_69033583165248_0
timestamp 1713338890
transform 1 0 65902 0 1 69512
box -698 -1424 698 1424
use M4_M3_CDNS_69033583165249  M4_M3_CDNS_69033583165249_0
timestamp 1713338890
transform 1 0 69514 0 1 65900
box -1424 -698 1424 698
use M4_M3_CDNS_69033583165250  M4_M3_CDNS_69033583165250_0
timestamp 1713338890
transform 1 0 69600 0 1 69230
box -1160 -38 104 38
use M4_M3_CDNS_69033583165251  M4_M3_CDNS_69033583165251_0
timestamp 1713338890
transform 1 0 69550 0 1 69098
box -1094 -38 170 38
use M4_M3_CDNS_69033583165252  M4_M3_CDNS_69033583165252_0
timestamp 1713338890
transform 1 0 67500 0 1 69846
box -698 -1094 698 1094
use M4_M3_CDNS_69033583165253  M4_M3_CDNS_69033583165253_0
timestamp 1713338890
transform 1 0 69846 0 1 67500
box -1094 -698 1094 698
use M4_M3_CDNS_69033583165254  M4_M3_CDNS_69033583165254_0
timestamp 1713338890
transform 1 0 69039 0 1 70154
box -632 -830 632 830
use M4_M3_CDNS_69033583165255  M4_M3_CDNS_69033583165255_0
timestamp 1713338890
transform 1 0 69427 0 1 68570
box -698 -38 302 38
use M4_M3_CDNS_69033583165256  M4_M3_CDNS_69033583165256_0
timestamp 1713338890
transform 1 0 69487 0 1 68966
box -1028 -38 236 38
use M4_M3_CDNS_69033583165257  M4_M3_CDNS_69033583165257_0
timestamp 1713338890
transform 1 0 70367 0 1 69039
box -566 -632 566 632
use M4_M3_CDNS_69033583165258  M4_M3_CDNS_69033583165258_0
timestamp 1713338890
transform 1 0 69427 0 1 68702
box -830 -38 302 38
use M4_M3_CDNS_69033583165259  M4_M3_CDNS_69033583165259_0
timestamp 1713338890
transform 1 0 69427 0 1 68834
box -962 -38 302 38
use M4_M3_CDNS_69033583165260  M4_M3_CDNS_69033583165260_0
timestamp 1713338890
transform 1 0 64300 0 1 69183
box -698 -1754 698 1754
use M4_M3_CDNS_69033583165261  M4_M3_CDNS_69033583165261_0
timestamp 1713338890
transform 1 0 69183 0 1 64300
box -1754 -698 1754 698
use M4_M3_CDNS_69033583165262  M4_M3_CDNS_69033583165262_0
timestamp 1713338890
transform 1 0 54700 0 1 67186
box -698 -3734 698 3734
use M4_M3_CDNS_69033583165263  M4_M3_CDNS_69033583165263_0
timestamp 1713338890
transform 1 0 56300 0 1 67518
box -698 -3404 698 3404
use M4_M3_CDNS_69033583165264  M4_M3_CDNS_69033583165264_0
timestamp 1713338890
transform 1 0 57900 0 1 67850
box -698 -3074 698 3074
use M4_M3_CDNS_69033583165265  M4_M3_CDNS_69033583165265_0
timestamp 1713338890
transform 1 0 59500 0 1 68183
box -698 -2744 698 2744
use M4_M3_CDNS_69033583165266  M4_M3_CDNS_69033583165266_0
timestamp 1713338890
transform 1 0 61100 0 1 68516
box -698 -2414 698 2414
use M4_M3_CDNS_69033583165267  M4_M3_CDNS_69033583165267_0
timestamp 1713338890
transform 1 0 67186 0 1 54700
box -3734 -698 3734 698
use M4_M3_CDNS_69033583165268  M4_M3_CDNS_69033583165268_0
timestamp 1713338890
transform 1 0 67518 0 1 56300
box -3404 -698 3404 698
use M4_M3_CDNS_69033583165269  M4_M3_CDNS_69033583165269_0
timestamp 1713338890
transform 1 0 67850 0 1 57900
box -3074 -698 3074 698
use M4_M3_CDNS_69033583165270  M4_M3_CDNS_69033583165270_0
timestamp 1713338890
transform 1 0 68183 0 1 59500
box -2744 -698 2744 698
use M4_M3_CDNS_69033583165271  M4_M3_CDNS_69033583165271_0
timestamp 1713338890
transform 1 0 68515 0 1 61101
box -2414 -698 2414 698
use M4_M3_CDNS_69033583165272  M4_M3_CDNS_69033583165272_0
timestamp 1713338890
transform 1 0 40300 0 1 64169
box -698 -6770 698 6770
use M4_M3_CDNS_69033583165273  M4_M3_CDNS_69033583165273_0
timestamp 1713338890
transform 1 0 41900 0 1 64505
box -698 -6440 698 6440
use M4_M3_CDNS_69033583165274  M4_M3_CDNS_69033583165274_0
timestamp 1713338890
transform 1 0 47500 0 1 65853
box -1490 -5120 1490 5120
use M4_M3_CDNS_69033583165275  M4_M3_CDNS_69033583165275_0
timestamp 1713338890
transform 1 0 44300 0 1 65170
box -1490 -5780 1490 5780
use M4_M3_CDNS_69033583165276  M4_M3_CDNS_69033583165276_0
timestamp 1713338890
transform 1 0 37900 0 1 63832
box -1490 -7100 1490 7100
use M4_M3_CDNS_69033583165277  M4_M3_CDNS_69033583165277_0
timestamp 1713338890
transform 1 0 49900 0 1 66188
box -698 -4790 698 4790
use M4_M3_CDNS_69033583165278  M4_M3_CDNS_69033583165278_0
timestamp 1713338890
transform 1 0 51500 0 1 66519
box -698 -4460 698 4460
use M4_M3_CDNS_69033583165279  M4_M3_CDNS_69033583165279_0
timestamp 1713338890
transform 1 0 65170 0 1 44300
box -5780 -1490 5780 1490
use M4_M3_CDNS_69033583165280  M4_M3_CDNS_69033583165280_0
timestamp 1713338890
transform 1 0 63832 0 1 37900
box -7100 -1490 7100 1490
use M4_M3_CDNS_69033583165281  M4_M3_CDNS_69033583165281_0
timestamp 1713338890
transform 1 0 64505 0 1 41900
box -6440 -698 6440 698
use M4_M3_CDNS_69033583165282  M4_M3_CDNS_69033583165282_0
timestamp 1713338890
transform 1 0 47259 0 1 15628
box -2678 -38 38 38
use M4_M3_CDNS_69033583165282  M4_M3_CDNS_69033583165282_1
timestamp 1713338890
transform 1 0 48595 0 1 18828
box -2678 -38 38 38
use M4_M3_CDNS_69033583165282  M4_M3_CDNS_69033583165282_2
timestamp 1713338890
transform 1 0 49921 0 1 22028
box -2678 -38 38 38
use M4_M3_CDNS_69033583165282  M4_M3_CDNS_69033583165282_3
timestamp 1713338890
transform 1 0 52601 0 1 28428
box -2678 -38 38 38
use M4_M3_CDNS_69033583165282  M4_M3_CDNS_69033583165282_4
timestamp 1713338890
transform 1 0 53939 0 1 31628
box -2678 -38 38 38
use M4_M3_CDNS_69033583165282  M4_M3_CDNS_69033583165282_5
timestamp 1713338890
transform 1 0 55271 0 1 34828
box -2678 -38 38 38
use M4_M3_CDNS_69033583165282  M4_M3_CDNS_69033583165282_6
timestamp 1713338890
transform 1 0 56612 0 1 38028
box -2678 -38 38 38
use M4_M3_CDNS_69033583165282  M4_M3_CDNS_69033583165282_7
timestamp 1713338890
transform 1 0 59288 0 1 44428
box -2678 -38 38 38
use M4_M3_CDNS_69033583165283  M4_M3_CDNS_69033583165283_0
timestamp 1713338890
transform 1 0 65853 0 1 47500
box -5120 -1490 5120 1490
use M4_M3_CDNS_69033583165284  M4_M3_CDNS_69033583165284_0
timestamp 1713338890
transform 1 0 66188 0 1 49900
box -4790 -698 4790 698
use M4_M3_CDNS_69033583165285  M4_M3_CDNS_69033583165285_0
timestamp 1713338890
transform 1 0 66519 0 1 51500
box -4460 -698 4460 698
use M4_M3_CDNS_69033583165286  M4_M3_CDNS_69033583165286_0
timestamp 1713338890
transform 1 0 61323 0 1 49492
box -632 -38 -28 38
use M4_M3_CDNS_69033583165286  M4_M3_CDNS_69033583165286_1
timestamp 1713338890
transform 1 0 61987 0 1 51092
box -632 -38 -28 38
use M4_M3_CDNS_69033583165286  M4_M3_CDNS_69033583165286_2
timestamp 1713338890
transform 1 0 62655 0 1 52692
box -632 -38 -28 38
use M4_M3_CDNS_69033583165287  M4_M3_CDNS_69033583165287_0
timestamp 1713338890
transform 1 0 61323 0 1 49624
box -764 -38 -28 38
use M4_M3_CDNS_69033583165287  M4_M3_CDNS_69033583165287_1
timestamp 1713338890
transform 1 0 61987 0 1 51224
box -764 -38 -28 38
use M4_M3_CDNS_69033583165287  M4_M3_CDNS_69033583165287_2
timestamp 1713338890
transform 1 0 62655 0 1 52824
box -764 -38 -28 38
use M4_M3_CDNS_69033583165288  M4_M3_CDNS_69033583165288_0
timestamp 1713338890
transform 1 0 61323 0 1 49756
box -896 -38 -28 38
use M4_M3_CDNS_69033583165288  M4_M3_CDNS_69033583165288_1
timestamp 1713338890
transform 1 0 61987 0 1 51356
box -896 -38 -28 38
use M4_M3_CDNS_69033583165288  M4_M3_CDNS_69033583165288_2
timestamp 1713338890
transform 1 0 62655 0 1 52956
box -896 -38 -28 38
use M4_M3_CDNS_69033583165289  M4_M3_CDNS_69033583165289_0
timestamp 1713338890
transform 1 0 61323 0 1 49888
box -1028 -38 -28 38
use M4_M3_CDNS_69033583165289  M4_M3_CDNS_69033583165289_1
timestamp 1713338890
transform 1 0 61987 0 1 51488
box -1028 -38 -28 38
use M4_M3_CDNS_69033583165289  M4_M3_CDNS_69033583165289_2
timestamp 1713338890
transform 1 0 62655 0 1 53088
box -1028 -38 -28 38
use M4_M3_CDNS_69033583165290  M4_M3_CDNS_69033583165290_0
timestamp 1713338890
transform 1 0 60655 0 1 46176
box -1160 -38 -28 38
use M4_M3_CDNS_69033583165290  M4_M3_CDNS_69033583165290_1
timestamp 1713338890
transform 1 0 61323 0 1 50020
box -1160 -38 -28 38
use M4_M3_CDNS_69033583165290  M4_M3_CDNS_69033583165290_2
timestamp 1713338890
transform 1 0 61987 0 1 51620
box -1160 -38 -28 38
use M4_M3_CDNS_69033583165290  M4_M3_CDNS_69033583165290_3
timestamp 1713338890
transform 1 0 62655 0 1 53220
box -1160 -38 -28 38
use M4_M3_CDNS_69033583165291  M4_M3_CDNS_69033583165291_0
timestamp 1713338890
transform 1 0 64169 0 1 40300
box -6770 -698 6770 698
use M4_M3_CDNS_69033583165292  M4_M3_CDNS_69033583165292_0
timestamp 1713338890
transform 1 0 61323 0 1 49360
box -500 -38 -28 38
use M4_M3_CDNS_69033583165292  M4_M3_CDNS_69033583165292_1
timestamp 1713338890
transform 1 0 61987 0 1 50960
box -500 -38 -28 38
use M4_M3_CDNS_69033583165292  M4_M3_CDNS_69033583165292_2
timestamp 1713338890
transform 1 0 62655 0 1 52560
box -500 -38 -28 38
use M4_M3_CDNS_69033583165293  M4_M3_CDNS_69033583165293_0
timestamp 1713338890
transform 1 0 47259 0 1 16156
box -3206 -38 38 38
use M4_M3_CDNS_69033583165293  M4_M3_CDNS_69033583165293_1
timestamp 1713338890
transform 1 0 48595 0 1 19356
box -3206 -38 38 38
use M4_M3_CDNS_69033583165293  M4_M3_CDNS_69033583165293_2
timestamp 1713338890
transform 1 0 49921 0 1 22556
box -3206 -38 38 38
use M4_M3_CDNS_69033583165293  M4_M3_CDNS_69033583165293_3
timestamp 1713338890
transform 1 0 52601 0 1 28956
box -3206 -38 38 38
use M4_M3_CDNS_69033583165293  M4_M3_CDNS_69033583165293_4
timestamp 1713338890
transform 1 0 53939 0 1 32156
box -3206 -38 38 38
use M4_M3_CDNS_69033583165293  M4_M3_CDNS_69033583165293_5
timestamp 1713338890
transform 1 0 55271 0 1 35356
box -3206 -38 38 38
use M4_M3_CDNS_69033583165293  M4_M3_CDNS_69033583165293_6
timestamp 1713338890
transform 1 0 56612 0 1 38556
box -3206 -38 38 38
use M4_M3_CDNS_69033583165293  M4_M3_CDNS_69033583165293_7
timestamp 1713338890
transform 1 0 59288 0 1 44956
box -3206 -38 38 38
use M4_M3_CDNS_69033583165294  M4_M3_CDNS_69033583165294_0
timestamp 1713338890
transform 1 0 47259 0 1 16024
box -3074 -38 38 38
use M4_M3_CDNS_69033583165294  M4_M3_CDNS_69033583165294_1
timestamp 1713338890
transform 1 0 48595 0 1 19224
box -3074 -38 38 38
use M4_M3_CDNS_69033583165294  M4_M3_CDNS_69033583165294_2
timestamp 1713338890
transform 1 0 49921 0 1 22424
box -3074 -38 38 38
use M4_M3_CDNS_69033583165294  M4_M3_CDNS_69033583165294_3
timestamp 1713338890
transform 1 0 52601 0 1 28824
box -3074 -38 38 38
use M4_M3_CDNS_69033583165294  M4_M3_CDNS_69033583165294_4
timestamp 1713338890
transform 1 0 53939 0 1 32024
box -3074 -38 38 38
use M4_M3_CDNS_69033583165294  M4_M3_CDNS_69033583165294_5
timestamp 1713338890
transform 1 0 55271 0 1 35224
box -3074 -38 38 38
use M4_M3_CDNS_69033583165294  M4_M3_CDNS_69033583165294_6
timestamp 1713338890
transform 1 0 56612 0 1 38424
box -3074 -38 38 38
use M4_M3_CDNS_69033583165294  M4_M3_CDNS_69033583165294_7
timestamp 1713338890
transform 1 0 59288 0 1 44824
box -3074 -38 38 38
use M4_M3_CDNS_69033583165295  M4_M3_CDNS_69033583165295_0
timestamp 1713338890
transform 1 0 47259 0 1 15892
box -2942 -38 38 38
use M4_M3_CDNS_69033583165295  M4_M3_CDNS_69033583165295_1
timestamp 1713338890
transform 1 0 48595 0 1 19092
box -2942 -38 38 38
use M4_M3_CDNS_69033583165295  M4_M3_CDNS_69033583165295_2
timestamp 1713338890
transform 1 0 49921 0 1 22292
box -2942 -38 38 38
use M4_M3_CDNS_69033583165295  M4_M3_CDNS_69033583165295_3
timestamp 1713338890
transform 1 0 52601 0 1 28692
box -2942 -38 38 38
use M4_M3_CDNS_69033583165295  M4_M3_CDNS_69033583165295_4
timestamp 1713338890
transform 1 0 53939 0 1 31892
box -2942 -38 38 38
use M4_M3_CDNS_69033583165295  M4_M3_CDNS_69033583165295_5
timestamp 1713338890
transform 1 0 55271 0 1 35092
box -2942 -38 38 38
use M4_M3_CDNS_69033583165295  M4_M3_CDNS_69033583165295_6
timestamp 1713338890
transform 1 0 56612 0 1 38292
box -2942 -38 38 38
use M4_M3_CDNS_69033583165295  M4_M3_CDNS_69033583165295_7
timestamp 1713338890
transform 1 0 59288 0 1 44692
box -2942 -38 38 38
use M4_M3_CDNS_69033583165296  M4_M3_CDNS_69033583165296_0
timestamp 1713338890
transform 1 0 47259 0 1 15760
box -2810 -38 38 38
use M4_M3_CDNS_69033583165296  M4_M3_CDNS_69033583165296_1
timestamp 1713338890
transform 1 0 48595 0 1 18960
box -2810 -38 38 38
use M4_M3_CDNS_69033583165296  M4_M3_CDNS_69033583165296_2
timestamp 1713338890
transform 1 0 49921 0 1 22160
box -2810 -38 38 38
use M4_M3_CDNS_69033583165296  M4_M3_CDNS_69033583165296_3
timestamp 1713338890
transform 1 0 52601 0 1 28560
box -2810 -38 38 38
use M4_M3_CDNS_69033583165296  M4_M3_CDNS_69033583165296_4
timestamp 1713338890
transform 1 0 53939 0 1 31760
box -2810 -38 38 38
use M4_M3_CDNS_69033583165296  M4_M3_CDNS_69033583165296_5
timestamp 1713338890
transform 1 0 55271 0 1 34960
box -2810 -38 38 38
use M4_M3_CDNS_69033583165296  M4_M3_CDNS_69033583165296_6
timestamp 1713338890
transform 1 0 56612 0 1 38160
box -2810 -38 38 38
use M4_M3_CDNS_69033583165296  M4_M3_CDNS_69033583165296_7
timestamp 1713338890
transform 1 0 59288 0 1 44560
box -2810 -38 38 38
use M4_M3_CDNS_69033583165297  M4_M3_CDNS_69033583165297_0
timestamp 1713338890
transform 1 0 60655 0 1 48024
box -3008 -38 -28 38
use M4_M3_CDNS_69033583165298  M4_M3_CDNS_69033583165298_0
timestamp 1713338890
transform 1 0 60655 0 1 48156
box -3140 -38 -28 38
use M4_M3_CDNS_69033583165299  M4_M3_CDNS_69033583165299_0
timestamp 1713338890
transform 1 0 60655 0 1 48288
box -3272 -38 -28 38
use M4_M3_CDNS_69033583165300  M4_M3_CDNS_69033583165300_0
timestamp 1713338890
transform 1 0 60655 0 1 48420
box -3404 -38 -28 38
use M4_M3_CDNS_69033583165301  M4_M3_CDNS_69033583165301_0
timestamp 1713338890
transform 1 0 60655 0 1 48552
box -3536 -38 -28 38
use M4_M3_CDNS_69033583165302  M4_M3_CDNS_69033583165302_0
timestamp 1713338890
transform 1 0 60655 0 1 48684
box -3668 -38 -28 38
use M4_M3_CDNS_69033583165303  M4_M3_CDNS_69033583165303_0
timestamp 1713338890
transform 1 0 60655 0 1 48816
box -3800 -38 -28 38
use M4_M3_CDNS_69033583165304  M4_M3_CDNS_69033583165304_0
timestamp 1713338890
transform 1 0 60655 0 1 48948
box -3932 -38 -28 38
use M4_M3_CDNS_69033583165305  M4_M3_CDNS_69033583165305_0
timestamp 1713338890
transform 1 0 60655 0 1 47628
box -2612 -38 -28 38
use M4_M3_CDNS_69033583165306  M4_M3_CDNS_69033583165306_0
timestamp 1713338890
transform 1 0 60655 0 1 47760
box -2744 -38 -28 38
use M4_M3_CDNS_69033583165307  M4_M3_CDNS_69033583165307_0
timestamp 1713338890
transform 1 0 60655 0 1 47892
box -2876 -38 -28 38
use M4_M3_CDNS_69033583165308  M4_M3_CDNS_69033583165308_0
timestamp 1713338890
transform 1 0 60655 0 1 46836
box -1820 -38 -28 38
use M4_M3_CDNS_69033583165309  M4_M3_CDNS_69033583165309_0
timestamp 1713338890
transform 1 0 60655 0 1 46968
box -1952 -38 -28 38
use M4_M3_CDNS_69033583165310  M4_M3_CDNS_69033583165310_0
timestamp 1713338890
transform 1 0 60655 0 1 47100
box -2084 -38 -28 38
use M4_M3_CDNS_69033583165311  M4_M3_CDNS_69033583165311_0
timestamp 1713338890
transform 1 0 60655 0 1 47232
box -2216 -38 -28 38
use M4_M3_CDNS_69033583165312  M4_M3_CDNS_69033583165312_0
timestamp 1713338890
transform 1 0 60655 0 1 47364
box -2348 -38 -28 38
use M4_M3_CDNS_69033583165313  M4_M3_CDNS_69033583165313_0
timestamp 1713338890
transform 1 0 60655 0 1 47496
box -2480 -38 -28 38
use M4_M3_CDNS_69033583165314  M4_M3_CDNS_69033583165314_0
timestamp 1713338890
transform 1 0 47259 0 1 15496
box -2546 -38 38 38
use M4_M3_CDNS_69033583165314  M4_M3_CDNS_69033583165314_1
timestamp 1713338890
transform 1 0 48595 0 1 18696
box -2546 -38 38 38
use M4_M3_CDNS_69033583165314  M4_M3_CDNS_69033583165314_2
timestamp 1713338890
transform 1 0 49921 0 1 21896
box -2546 -38 38 38
use M4_M3_CDNS_69033583165314  M4_M3_CDNS_69033583165314_3
timestamp 1713338890
transform 1 0 52601 0 1 28296
box -2546 -38 38 38
use M4_M3_CDNS_69033583165314  M4_M3_CDNS_69033583165314_4
timestamp 1713338890
transform 1 0 53939 0 1 31496
box -2546 -38 38 38
use M4_M3_CDNS_69033583165314  M4_M3_CDNS_69033583165314_5
timestamp 1713338890
transform 1 0 55271 0 1 34696
box -2546 -38 38 38
use M4_M3_CDNS_69033583165314  M4_M3_CDNS_69033583165314_6
timestamp 1713338890
transform 1 0 56612 0 1 37896
box -2546 -38 38 38
use M4_M3_CDNS_69033583165314  M4_M3_CDNS_69033583165314_7
timestamp 1713338890
transform 1 0 59288 0 1 44296
box -2546 -38 38 38
use M4_M3_CDNS_69033583165315  M4_M3_CDNS_69033583165315_0
timestamp 1713338890
transform 1 0 47259 0 1 15364
box -2414 -38 38 38
use M4_M3_CDNS_69033583165315  M4_M3_CDNS_69033583165315_1
timestamp 1713338890
transform 1 0 48595 0 1 18564
box -2414 -38 38 38
use M4_M3_CDNS_69033583165315  M4_M3_CDNS_69033583165315_2
timestamp 1713338890
transform 1 0 49921 0 1 21764
box -2414 -38 38 38
use M4_M3_CDNS_69033583165315  M4_M3_CDNS_69033583165315_3
timestamp 1713338890
transform 1 0 52601 0 1 28164
box -2414 -38 38 38
use M4_M3_CDNS_69033583165315  M4_M3_CDNS_69033583165315_4
timestamp 1713338890
transform 1 0 53939 0 1 31364
box -2414 -38 38 38
use M4_M3_CDNS_69033583165315  M4_M3_CDNS_69033583165315_5
timestamp 1713338890
transform 1 0 55271 0 1 34564
box -2414 -38 38 38
use M4_M3_CDNS_69033583165315  M4_M3_CDNS_69033583165315_6
timestamp 1713338890
transform 1 0 56612 0 1 37764
box -2414 -38 38 38
use M4_M3_CDNS_69033583165315  M4_M3_CDNS_69033583165315_7
timestamp 1713338890
transform 1 0 59288 0 1 44164
box -2414 -38 38 38
use M4_M3_CDNS_69033583165316  M4_M3_CDNS_69033583165316_0
timestamp 1713338890
transform 1 0 47259 0 1 15232
box -2282 -38 38 38
use M4_M3_CDNS_69033583165316  M4_M3_CDNS_69033583165316_1
timestamp 1713338890
transform 1 0 48595 0 1 18432
box -2282 -38 38 38
use M4_M3_CDNS_69033583165316  M4_M3_CDNS_69033583165316_2
timestamp 1713338890
transform 1 0 49921 0 1 21632
box -2282 -38 38 38
use M4_M3_CDNS_69033583165316  M4_M3_CDNS_69033583165316_3
timestamp 1713338890
transform 1 0 52601 0 1 28032
box -2282 -38 38 38
use M4_M3_CDNS_69033583165316  M4_M3_CDNS_69033583165316_4
timestamp 1713338890
transform 1 0 53939 0 1 31232
box -2282 -38 38 38
use M4_M3_CDNS_69033583165316  M4_M3_CDNS_69033583165316_5
timestamp 1713338890
transform 1 0 55271 0 1 34432
box -2282 -38 38 38
use M4_M3_CDNS_69033583165316  M4_M3_CDNS_69033583165316_6
timestamp 1713338890
transform 1 0 56612 0 1 37632
box -2282 -38 38 38
use M4_M3_CDNS_69033583165316  M4_M3_CDNS_69033583165316_7
timestamp 1713338890
transform 1 0 59288 0 1 44032
box -2282 -38 38 38
use M4_M3_CDNS_69033583165317  M4_M3_CDNS_69033583165317_0
timestamp 1713338890
transform 1 0 47259 0 1 15100
box -2150 -38 38 38
use M4_M3_CDNS_69033583165317  M4_M3_CDNS_69033583165317_1
timestamp 1713338890
transform 1 0 48595 0 1 18300
box -2150 -38 38 38
use M4_M3_CDNS_69033583165317  M4_M3_CDNS_69033583165317_2
timestamp 1713338890
transform 1 0 49921 0 1 21500
box -2150 -38 38 38
use M4_M3_CDNS_69033583165317  M4_M3_CDNS_69033583165317_3
timestamp 1713338890
transform 1 0 52601 0 1 27900
box -2150 -38 38 38
use M4_M3_CDNS_69033583165317  M4_M3_CDNS_69033583165317_4
timestamp 1713338890
transform 1 0 53939 0 1 31100
box -2150 -38 38 38
use M4_M3_CDNS_69033583165317  M4_M3_CDNS_69033583165317_5
timestamp 1713338890
transform 1 0 55271 0 1 34300
box -2150 -38 38 38
use M4_M3_CDNS_69033583165317  M4_M3_CDNS_69033583165317_6
timestamp 1713338890
transform 1 0 56612 0 1 37500
box -2150 -38 38 38
use M4_M3_CDNS_69033583165317  M4_M3_CDNS_69033583165317_7
timestamp 1713338890
transform 1 0 59288 0 1 43900
box -2150 -38 38 38
use M4_M3_CDNS_69033583165318  M4_M3_CDNS_69033583165318_0
timestamp 1713338890
transform 1 0 47259 0 1 14968
box -2018 -38 38 38
use M4_M3_CDNS_69033583165318  M4_M3_CDNS_69033583165318_1
timestamp 1713338890
transform 1 0 48595 0 1 18168
box -2018 -38 38 38
use M4_M3_CDNS_69033583165318  M4_M3_CDNS_69033583165318_2
timestamp 1713338890
transform 1 0 49921 0 1 21368
box -2018 -38 38 38
use M4_M3_CDNS_69033583165318  M4_M3_CDNS_69033583165318_3
timestamp 1713338890
transform 1 0 52601 0 1 27768
box -2018 -38 38 38
use M4_M3_CDNS_69033583165318  M4_M3_CDNS_69033583165318_4
timestamp 1713338890
transform 1 0 53939 0 1 30968
box -2018 -38 38 38
use M4_M3_CDNS_69033583165318  M4_M3_CDNS_69033583165318_5
timestamp 1713338890
transform 1 0 55271 0 1 34168
box -2018 -38 38 38
use M4_M3_CDNS_69033583165318  M4_M3_CDNS_69033583165318_6
timestamp 1713338890
transform 1 0 56612 0 1 37368
box -2018 -38 38 38
use M4_M3_CDNS_69033583165318  M4_M3_CDNS_69033583165318_7
timestamp 1713338890
transform 1 0 59288 0 1 43768
box -2018 -38 38 38
use M4_M3_CDNS_69033583165319  M4_M3_CDNS_69033583165319_0
timestamp 1713338890
transform 1 0 47259 0 1 14836
box -1886 -38 38 38
use M4_M3_CDNS_69033583165319  M4_M3_CDNS_69033583165319_1
timestamp 1713338890
transform 1 0 48595 0 1 18036
box -1886 -38 38 38
use M4_M3_CDNS_69033583165319  M4_M3_CDNS_69033583165319_2
timestamp 1713338890
transform 1 0 49921 0 1 21236
box -1886 -38 38 38
use M4_M3_CDNS_69033583165319  M4_M3_CDNS_69033583165319_3
timestamp 1713338890
transform 1 0 52601 0 1 27636
box -1886 -38 38 38
use M4_M3_CDNS_69033583165319  M4_M3_CDNS_69033583165319_4
timestamp 1713338890
transform 1 0 53939 0 1 30836
box -1886 -38 38 38
use M4_M3_CDNS_69033583165319  M4_M3_CDNS_69033583165319_5
timestamp 1713338890
transform 1 0 55271 0 1 34036
box -1886 -38 38 38
use M4_M3_CDNS_69033583165319  M4_M3_CDNS_69033583165319_6
timestamp 1713338890
transform 1 0 56612 0 1 37236
box -1886 -38 38 38
use M4_M3_CDNS_69033583165319  M4_M3_CDNS_69033583165319_7
timestamp 1713338890
transform 1 0 59288 0 1 43636
box -1886 -38 38 38
use M4_M3_CDNS_69033583165320  M4_M3_CDNS_69033583165320_0
timestamp 1713338890
transform 1 0 18700 0 1 59824
box -1490 -11126 1490 11126
use M4_M3_CDNS_69033583165321  M4_M3_CDNS_69033583165321_0
timestamp 1713338890
transform 1 0 15500 0 1 59156
box -1490 -11786 1490 11786
use M4_M3_CDNS_69033583165322  M4_M3_CDNS_69033583165322_0
timestamp 1713338890
transform 1 0 25900 0 1 61160
box -698 -9806 698 9806
use M4_M3_CDNS_69033583165323  M4_M3_CDNS_69033583165323_0
timestamp 1713338890
transform 1 0 28300 0 1 61827
box -1490 -9146 1490 9146
use M4_M3_CDNS_69033583165324  M4_M3_CDNS_69033583165324_0
timestamp 1713338890
transform 1 0 21900 0 1 60487
box -1490 -10466 1490 10466
use M4_M3_CDNS_69033583165325  M4_M3_CDNS_69033583165325_0
timestamp 1713338890
transform 1 0 24300 0 1 60826
box -698 -10136 698 10136
use M4_M3_CDNS_69033583165326  M4_M3_CDNS_69033583165326_0
timestamp 1713338890
transform 1 0 31500 0 1 62496
box -1490 -8486 1490 8486
use M4_M3_CDNS_69033583165327  M4_M3_CDNS_69033583165327_0
timestamp 1713338890
transform 1 0 60826 0 1 24300
box -10136 -698 10136 698
use M4_M3_CDNS_69033583165328  M4_M3_CDNS_69033583165328_0
timestamp 1713338890
transform 1 0 61160 0 1 25900
box -9806 -698 9806 698
use M4_M3_CDNS_69033583165329  M4_M3_CDNS_69033583165329_0
timestamp 1713338890
transform 1 0 61827 0 1 28300
box -9146 -1490 9146 1490
use M4_M3_CDNS_69033583165330  M4_M3_CDNS_69033583165330_0
timestamp 1713338890
transform 1 0 59824 0 1 18700
box -11126 -1490 11126 1490
use M4_M3_CDNS_69033583165331  M4_M3_CDNS_69033583165331_0
timestamp 1713338890
transform 1 0 60487 0 1 21900
box -10466 -1490 10466 1490
use M4_M3_CDNS_69033583165332  M4_M3_CDNS_69033583165332_0
timestamp 1713338890
transform 1 0 59156 0 1 15500
box -11786 -1490 11786 1490
use M4_M3_CDNS_69033583165333  M4_M3_CDNS_69033583165333_0
timestamp 1713338890
transform 1 0 62496 0 1 31500
box -8486 -1490 8486 1490
use POWER_RAIL_COR_1  POWER_RAIL_COR_1_0
timestamp 1713338890
transform 1 0 0 0 1 0
box 13097 13097 71000 71000
<< labels >>
rlabel metal3 s 70444 56376 70444 56376 4 DVDD
port 1 nsew
rlabel metal3 s 70444 59576 70444 59576 4 DVDD
port 1 nsew
rlabel metal3 s 70444 67411 70444 67411 4 DVDD
port 1 nsew
rlabel metal3 s 70444 24237 70444 24237 4 DVDD
port 1 nsew
rlabel metal3 s 70444 28347 70444 28347 4 DVDD
port 1 nsew
rlabel metal3 s 70444 31562 70444 31562 4 DVDD
port 1 nsew
rlabel metal3 s 70444 34676 70444 34676 4 DVDD
port 1 nsew
rlabel metal3 s 70444 37912 70444 37912 4 DVDD
port 1 nsew
rlabel metal3 s 70444 41930 70444 41930 4 DVDD
port 1 nsew
rlabel metal3 s 70444 44321 70444 44321 4 DVDD
port 1 nsew
rlabel metal3 s 70444 53176 70444 53176 4 DVDD
port 1 nsew
rlabel metal3 s 70444 54611 70444 54611 4 DVDD
port 1 nsew
rlabel metal3 s 70445 64211 70445 64211 4 VSS
port 2 nsew
rlabel metal3 s 70549 49976 70549 49976 4 VSS
port 2 nsew
rlabel metal3 s 70444 57811 70444 57811 4 DVSS
port 3 nsew
rlabel metal3 s 70444 61011 70444 61011 4 DVSS
port 3 nsew
rlabel metal3 s 70444 65976 70444 65976 4 DVSS
port 3 nsew
rlabel metal3 s 70444 69002 70444 69002 4 DVSS
port 3 nsew
rlabel metal3 s 70422 15703 70422 15703 4 DVSS
port 3 nsew
rlabel metal3 s 70375 18874 70375 18874 4 DVSS
port 3 nsew
rlabel metal3 s 70444 21860 70444 21860 4 DVSS
port 3 nsew
rlabel metal3 s 70444 26053 70444 26053 4 DVSS
port 3 nsew
rlabel metal3 s 70444 40295 70444 40295 4 DVSS
port 3 nsew
rlabel metal3 s 70444 47548 70444 47548 4 DVSS
port 3 nsew
rlabel metal3 s 70549 51411 70549 51411 4 VDD
port 4 nsew
rlabel metal3 s 70444 62776 70444 62776 4 VDD
port 4 nsew
<< end >>
