magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1045 -1305 1045 1305
<< metal1 >>
rect -45 299 45 305
rect -45 -299 -39 299
rect 39 -299 45 299
rect -45 -305 45 -299
<< via1 >>
rect -39 -299 39 299
<< metal2 >>
rect -45 299 45 305
rect -45 -299 -39 299
rect 39 -299 45 299
rect -45 -305 45 -299
<< end >>
