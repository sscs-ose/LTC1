magic
tech gf180mcuC
magscale 1 10
timestamp 1693281404
<< error_p >>
rect -5527 -58 -5481 58
rect -5183 -58 -5137 58
rect -4839 -58 -4793 58
rect -4495 -58 -4449 58
rect -4151 -58 -4105 58
rect -3807 -58 -3761 58
rect -3463 -58 -3417 58
rect -3119 -58 -3073 58
rect -2775 -58 -2729 58
rect -2431 -58 -2385 58
rect -2087 -58 -2041 58
rect -1743 -58 -1697 58
rect -1399 -58 -1353 58
rect -1055 -58 -1009 58
rect -711 -58 -665 58
rect -367 -58 -321 58
rect -23 -58 23 58
rect 321 -58 367 58
rect 665 -58 711 58
rect 1009 -58 1055 58
rect 1353 -58 1399 58
rect 1697 -58 1743 58
rect 2041 -58 2087 58
rect 2385 -58 2431 58
rect 2729 -58 2775 58
rect 3073 -58 3119 58
rect 3417 -58 3463 58
rect 3761 -58 3807 58
rect 4105 -58 4151 58
rect 4449 -58 4495 58
rect 4793 -58 4839 58
rect 5137 -58 5183 58
rect 5481 -58 5527 58
<< pwell >>
rect -5564 -128 5564 128
<< nmos >>
rect -5452 -60 -5212 60
rect -5108 -60 -4868 60
rect -4764 -60 -4524 60
rect -4420 -60 -4180 60
rect -4076 -60 -3836 60
rect -3732 -60 -3492 60
rect -3388 -60 -3148 60
rect -3044 -60 -2804 60
rect -2700 -60 -2460 60
rect -2356 -60 -2116 60
rect -2012 -60 -1772 60
rect -1668 -60 -1428 60
rect -1324 -60 -1084 60
rect -980 -60 -740 60
rect -636 -60 -396 60
rect -292 -60 -52 60
rect 52 -60 292 60
rect 396 -60 636 60
rect 740 -60 980 60
rect 1084 -60 1324 60
rect 1428 -60 1668 60
rect 1772 -60 2012 60
rect 2116 -60 2356 60
rect 2460 -60 2700 60
rect 2804 -60 3044 60
rect 3148 -60 3388 60
rect 3492 -60 3732 60
rect 3836 -60 4076 60
rect 4180 -60 4420 60
rect 4524 -60 4764 60
rect 4868 -60 5108 60
rect 5212 -60 5452 60
<< ndiff >>
rect -5540 47 -5452 60
rect -5540 -47 -5527 47
rect -5481 -47 -5452 47
rect -5540 -60 -5452 -47
rect -5212 47 -5108 60
rect -5212 -47 -5183 47
rect -5137 -47 -5108 47
rect -5212 -60 -5108 -47
rect -4868 47 -4764 60
rect -4868 -47 -4839 47
rect -4793 -47 -4764 47
rect -4868 -60 -4764 -47
rect -4524 47 -4420 60
rect -4524 -47 -4495 47
rect -4449 -47 -4420 47
rect -4524 -60 -4420 -47
rect -4180 47 -4076 60
rect -4180 -47 -4151 47
rect -4105 -47 -4076 47
rect -4180 -60 -4076 -47
rect -3836 47 -3732 60
rect -3836 -47 -3807 47
rect -3761 -47 -3732 47
rect -3836 -60 -3732 -47
rect -3492 47 -3388 60
rect -3492 -47 -3463 47
rect -3417 -47 -3388 47
rect -3492 -60 -3388 -47
rect -3148 47 -3044 60
rect -3148 -47 -3119 47
rect -3073 -47 -3044 47
rect -3148 -60 -3044 -47
rect -2804 47 -2700 60
rect -2804 -47 -2775 47
rect -2729 -47 -2700 47
rect -2804 -60 -2700 -47
rect -2460 47 -2356 60
rect -2460 -47 -2431 47
rect -2385 -47 -2356 47
rect -2460 -60 -2356 -47
rect -2116 47 -2012 60
rect -2116 -47 -2087 47
rect -2041 -47 -2012 47
rect -2116 -60 -2012 -47
rect -1772 47 -1668 60
rect -1772 -47 -1743 47
rect -1697 -47 -1668 47
rect -1772 -60 -1668 -47
rect -1428 47 -1324 60
rect -1428 -47 -1399 47
rect -1353 -47 -1324 47
rect -1428 -60 -1324 -47
rect -1084 47 -980 60
rect -1084 -47 -1055 47
rect -1009 -47 -980 47
rect -1084 -60 -980 -47
rect -740 47 -636 60
rect -740 -47 -711 47
rect -665 -47 -636 47
rect -740 -60 -636 -47
rect -396 47 -292 60
rect -396 -47 -367 47
rect -321 -47 -292 47
rect -396 -60 -292 -47
rect -52 47 52 60
rect -52 -47 -23 47
rect 23 -47 52 47
rect -52 -60 52 -47
rect 292 47 396 60
rect 292 -47 321 47
rect 367 -47 396 47
rect 292 -60 396 -47
rect 636 47 740 60
rect 636 -47 665 47
rect 711 -47 740 47
rect 636 -60 740 -47
rect 980 47 1084 60
rect 980 -47 1009 47
rect 1055 -47 1084 47
rect 980 -60 1084 -47
rect 1324 47 1428 60
rect 1324 -47 1353 47
rect 1399 -47 1428 47
rect 1324 -60 1428 -47
rect 1668 47 1772 60
rect 1668 -47 1697 47
rect 1743 -47 1772 47
rect 1668 -60 1772 -47
rect 2012 47 2116 60
rect 2012 -47 2041 47
rect 2087 -47 2116 47
rect 2012 -60 2116 -47
rect 2356 47 2460 60
rect 2356 -47 2385 47
rect 2431 -47 2460 47
rect 2356 -60 2460 -47
rect 2700 47 2804 60
rect 2700 -47 2729 47
rect 2775 -47 2804 47
rect 2700 -60 2804 -47
rect 3044 47 3148 60
rect 3044 -47 3073 47
rect 3119 -47 3148 47
rect 3044 -60 3148 -47
rect 3388 47 3492 60
rect 3388 -47 3417 47
rect 3463 -47 3492 47
rect 3388 -60 3492 -47
rect 3732 47 3836 60
rect 3732 -47 3761 47
rect 3807 -47 3836 47
rect 3732 -60 3836 -47
rect 4076 47 4180 60
rect 4076 -47 4105 47
rect 4151 -47 4180 47
rect 4076 -60 4180 -47
rect 4420 47 4524 60
rect 4420 -47 4449 47
rect 4495 -47 4524 47
rect 4420 -60 4524 -47
rect 4764 47 4868 60
rect 4764 -47 4793 47
rect 4839 -47 4868 47
rect 4764 -60 4868 -47
rect 5108 47 5212 60
rect 5108 -47 5137 47
rect 5183 -47 5212 47
rect 5108 -60 5212 -47
rect 5452 47 5540 60
rect 5452 -47 5481 47
rect 5527 -47 5540 47
rect 5452 -60 5540 -47
<< ndiffc >>
rect -5527 -47 -5481 47
rect -5183 -47 -5137 47
rect -4839 -47 -4793 47
rect -4495 -47 -4449 47
rect -4151 -47 -4105 47
rect -3807 -47 -3761 47
rect -3463 -47 -3417 47
rect -3119 -47 -3073 47
rect -2775 -47 -2729 47
rect -2431 -47 -2385 47
rect -2087 -47 -2041 47
rect -1743 -47 -1697 47
rect -1399 -47 -1353 47
rect -1055 -47 -1009 47
rect -711 -47 -665 47
rect -367 -47 -321 47
rect -23 -47 23 47
rect 321 -47 367 47
rect 665 -47 711 47
rect 1009 -47 1055 47
rect 1353 -47 1399 47
rect 1697 -47 1743 47
rect 2041 -47 2087 47
rect 2385 -47 2431 47
rect 2729 -47 2775 47
rect 3073 -47 3119 47
rect 3417 -47 3463 47
rect 3761 -47 3807 47
rect 4105 -47 4151 47
rect 4449 -47 4495 47
rect 4793 -47 4839 47
rect 5137 -47 5183 47
rect 5481 -47 5527 47
<< polysilicon >>
rect -5452 60 -5212 104
rect -5108 60 -4868 104
rect -4764 60 -4524 104
rect -4420 60 -4180 104
rect -4076 60 -3836 104
rect -3732 60 -3492 104
rect -3388 60 -3148 104
rect -3044 60 -2804 104
rect -2700 60 -2460 104
rect -2356 60 -2116 104
rect -2012 60 -1772 104
rect -1668 60 -1428 104
rect -1324 60 -1084 104
rect -980 60 -740 104
rect -636 60 -396 104
rect -292 60 -52 104
rect 52 60 292 104
rect 396 60 636 104
rect 740 60 980 104
rect 1084 60 1324 104
rect 1428 60 1668 104
rect 1772 60 2012 104
rect 2116 60 2356 104
rect 2460 60 2700 104
rect 2804 60 3044 104
rect 3148 60 3388 104
rect 3492 60 3732 104
rect 3836 60 4076 104
rect 4180 60 4420 104
rect 4524 60 4764 104
rect 4868 60 5108 104
rect 5212 60 5452 104
rect -5452 -104 -5212 -60
rect -5108 -104 -4868 -60
rect -4764 -104 -4524 -60
rect -4420 -104 -4180 -60
rect -4076 -104 -3836 -60
rect -3732 -104 -3492 -60
rect -3388 -104 -3148 -60
rect -3044 -104 -2804 -60
rect -2700 -104 -2460 -60
rect -2356 -104 -2116 -60
rect -2012 -104 -1772 -60
rect -1668 -104 -1428 -60
rect -1324 -104 -1084 -60
rect -980 -104 -740 -60
rect -636 -104 -396 -60
rect -292 -104 -52 -60
rect 52 -104 292 -60
rect 396 -104 636 -60
rect 740 -104 980 -60
rect 1084 -104 1324 -60
rect 1428 -104 1668 -60
rect 1772 -104 2012 -60
rect 2116 -104 2356 -60
rect 2460 -104 2700 -60
rect 2804 -104 3044 -60
rect 3148 -104 3388 -60
rect 3492 -104 3732 -60
rect 3836 -104 4076 -60
rect 4180 -104 4420 -60
rect 4524 -104 4764 -60
rect 4868 -104 5108 -60
rect 5212 -104 5452 -60
<< metal1 >>
rect -5527 47 -5481 58
rect -5527 -58 -5481 -47
rect -5183 47 -5137 58
rect -5183 -58 -5137 -47
rect -4839 47 -4793 58
rect -4839 -58 -4793 -47
rect -4495 47 -4449 58
rect -4495 -58 -4449 -47
rect -4151 47 -4105 58
rect -4151 -58 -4105 -47
rect -3807 47 -3761 58
rect -3807 -58 -3761 -47
rect -3463 47 -3417 58
rect -3463 -58 -3417 -47
rect -3119 47 -3073 58
rect -3119 -58 -3073 -47
rect -2775 47 -2729 58
rect -2775 -58 -2729 -47
rect -2431 47 -2385 58
rect -2431 -58 -2385 -47
rect -2087 47 -2041 58
rect -2087 -58 -2041 -47
rect -1743 47 -1697 58
rect -1743 -58 -1697 -47
rect -1399 47 -1353 58
rect -1399 -58 -1353 -47
rect -1055 47 -1009 58
rect -1055 -58 -1009 -47
rect -711 47 -665 58
rect -711 -58 -665 -47
rect -367 47 -321 58
rect -367 -58 -321 -47
rect -23 47 23 58
rect -23 -58 23 -47
rect 321 47 367 58
rect 321 -58 367 -47
rect 665 47 711 58
rect 665 -58 711 -47
rect 1009 47 1055 58
rect 1009 -58 1055 -47
rect 1353 47 1399 58
rect 1353 -58 1399 -47
rect 1697 47 1743 58
rect 1697 -58 1743 -47
rect 2041 47 2087 58
rect 2041 -58 2087 -47
rect 2385 47 2431 58
rect 2385 -58 2431 -47
rect 2729 47 2775 58
rect 2729 -58 2775 -47
rect 3073 47 3119 58
rect 3073 -58 3119 -47
rect 3417 47 3463 58
rect 3417 -58 3463 -47
rect 3761 47 3807 58
rect 3761 -58 3807 -47
rect 4105 47 4151 58
rect 4105 -58 4151 -47
rect 4449 47 4495 58
rect 4449 -58 4495 -47
rect 4793 47 4839 58
rect 4793 -58 4839 -47
rect 5137 47 5183 58
rect 5137 -58 5183 -47
rect 5481 47 5527 58
rect 5481 -58 5527 -47
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 0.6 l 1.2 m 1 nf 32 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
