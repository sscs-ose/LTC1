magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2000 -2000 2984 2160
<< polysilicon >>
rect 0 103 102 160
rect 0 57 13 103
rect 59 57 102 103
rect 0 0 102 57
rect 882 103 984 160
rect 882 57 925 103
rect 971 57 984 103
rect 882 0 984 57
<< polycontact >>
rect 13 57 59 103
rect 925 57 971 103
<< ppolyres >>
rect 102 0 882 160
<< metal1 >>
rect 2 103 70 158
rect 2 57 13 103
rect 59 57 70 103
rect 2 2 70 57
rect 914 103 982 158
rect 914 57 925 103
rect 971 57 982 103
rect 914 2 982 57
<< labels >>
rlabel polycontact 948 80 948 80 4 MINUS
rlabel polycontact 36 80 36 80 4 PLUS
<< end >>
