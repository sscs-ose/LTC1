magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1305 -1019 1305 1019
<< metal1 >>
rect -305 13 305 19
rect -305 -13 -299 13
rect 299 -13 305 13
rect -305 -19 305 -13
<< via1 >>
rect -299 -13 299 13
<< metal2 >>
rect -305 13 305 19
rect -305 -13 -299 13
rect 299 -13 305 13
rect -305 -19 305 -13
<< end >>
