* NGSPICE file created from and_2_flat.ext - technology: gf180mcuC

.subckt and_2_flat VDD IN2 OUT IN1 VSS
X0 VDD IN1.t0 nand2_0.OUT VDD.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1 nand2_0.OUT IN2.t0 VDD.t5 VDD.t0 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2 OUT nand2_0.OUT VSS.t2 VSS.t1 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X3 OUT nand2_0.OUT VDD.t4 VDD.t3 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X4 nand2_0.OUT IN1.t1 a_495_1252# VSS.t0 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X5 a_495_1252# IN2.t1 VSS.t4 VSS.t3 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
R0 IN1.n0 IN1.t1 31.528
R1 IN1.n0 IN1.t0 15.3826
R2 IN1 IN1.n0 8.85806
R3 VDD.n5 VDD.n4 213.458
R4 VDD.n5 VDD.n3 52.9326
R5 VDD.n4 VDD.t3 22.7928
R6 VDD VDD.n5 6.3005
R7 VDD VDD.t5 5.21701
R8 VDD.n2 VDD.t4 5.14703
R9 VDD.n1 VDD.n0 5.13287
R10 VDD.n2 VDD.n1 0.136194
R11 VDD VDD.n1 0.106177
R12 VDD.n3 VDD.n2 0.0460556
R13 VDD.n4 VDD.t0 0.00528088
R14 VDD.n3 VDD 0.00105556
R15 IN2.n0 IN2.t0 30.9379
R16 IN2.n0 IN2.t1 21.6422
R17 IN2 IN2.n0 4.00388
R18 VSS.t0 VSS.n1 1242.83
R19 VSS.n1 VSS.t1 1037.75
R20 VSS.n2 VSS.t0 596.558
R21 VSS.n2 VSS.t3 397.707
R22 VSS.n1 VSS 391.339
R23 VSS.n0 VSS.t2 9.34566
R24 VSS VSS.t4 7.30963
R25 VSS VSS.n2 5.2005
R26 VSS.n0 VSS 0.375997
R27 VSS VSS.n0 0.0647857
R28 OUT OUT.n1 9.42932
R29 OUT OUT.n0 5.13104
C0 VDD IN2 0.146f
C1 OUT IN1 0.00888f
C2 nand2_0.OUT OUT 0.125f
C3 a_495_1252# IN1 0.00348f
C4 nand2_0.OUT IN1 0.267f
C5 nand2_0.OUT a_495_1252# 0.0691f
C6 OUT VDD 0.122f
C7 VDD IN1 0.239f
C8 IN2 IN1 0.0466f
C9 VDD a_495_1252# 3.14e-19
C10 a_495_1252# IN2 0.00347f
C11 nand2_0.OUT VDD 0.408f
C12 nand2_0.OUT IN2 0.0956f
C13 a_495_1252# VSS 0.0678f
C14 OUT VSS 0.148f
C15 nand2_0.OUT VSS 0.485f
C16 IN1 VSS 0.219f
C17 IN2 VSS 0.292f
C18 VDD VSS 1.85f
.ends

