magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -7811 -3285 7811 3285
<< psubdiff >>
rect -5811 1263 5811 1285
rect -5811 1217 -5789 1263
rect -5743 1217 -5665 1263
rect -5619 1217 -5541 1263
rect -5495 1217 -5417 1263
rect -5371 1217 -5293 1263
rect -5247 1217 -5169 1263
rect -5123 1217 -5045 1263
rect -4999 1217 -4921 1263
rect -4875 1217 -4797 1263
rect -4751 1217 -4673 1263
rect -4627 1217 -4549 1263
rect -4503 1217 -4425 1263
rect -4379 1217 -4301 1263
rect -4255 1217 -4177 1263
rect -4131 1217 -4053 1263
rect -4007 1217 -3929 1263
rect -3883 1217 -3805 1263
rect -3759 1217 -3681 1263
rect -3635 1217 -3557 1263
rect -3511 1217 -3433 1263
rect -3387 1217 -3309 1263
rect -3263 1217 -3185 1263
rect -3139 1217 -3061 1263
rect -3015 1217 -2937 1263
rect -2891 1217 -2813 1263
rect -2767 1217 -2689 1263
rect -2643 1217 -2565 1263
rect -2519 1217 -2441 1263
rect -2395 1217 -2317 1263
rect -2271 1217 -2193 1263
rect -2147 1217 -2069 1263
rect -2023 1217 -1945 1263
rect -1899 1217 -1821 1263
rect -1775 1217 -1697 1263
rect -1651 1217 -1573 1263
rect -1527 1217 -1449 1263
rect -1403 1217 -1325 1263
rect -1279 1217 -1201 1263
rect -1155 1217 -1077 1263
rect -1031 1217 -953 1263
rect -907 1217 -829 1263
rect -783 1217 -705 1263
rect -659 1217 -581 1263
rect -535 1217 -457 1263
rect -411 1217 -333 1263
rect -287 1217 -209 1263
rect -163 1217 -85 1263
rect -39 1217 39 1263
rect 85 1217 163 1263
rect 209 1217 287 1263
rect 333 1217 411 1263
rect 457 1217 535 1263
rect 581 1217 659 1263
rect 705 1217 783 1263
rect 829 1217 907 1263
rect 953 1217 1031 1263
rect 1077 1217 1155 1263
rect 1201 1217 1279 1263
rect 1325 1217 1403 1263
rect 1449 1217 1527 1263
rect 1573 1217 1651 1263
rect 1697 1217 1775 1263
rect 1821 1217 1899 1263
rect 1945 1217 2023 1263
rect 2069 1217 2147 1263
rect 2193 1217 2271 1263
rect 2317 1217 2395 1263
rect 2441 1217 2519 1263
rect 2565 1217 2643 1263
rect 2689 1217 2767 1263
rect 2813 1217 2891 1263
rect 2937 1217 3015 1263
rect 3061 1217 3139 1263
rect 3185 1217 3263 1263
rect 3309 1217 3387 1263
rect 3433 1217 3511 1263
rect 3557 1217 3635 1263
rect 3681 1217 3759 1263
rect 3805 1217 3883 1263
rect 3929 1217 4007 1263
rect 4053 1217 4131 1263
rect 4177 1217 4255 1263
rect 4301 1217 4379 1263
rect 4425 1217 4503 1263
rect 4549 1217 4627 1263
rect 4673 1217 4751 1263
rect 4797 1217 4875 1263
rect 4921 1217 4999 1263
rect 5045 1217 5123 1263
rect 5169 1217 5247 1263
rect 5293 1217 5371 1263
rect 5417 1217 5495 1263
rect 5541 1217 5619 1263
rect 5665 1217 5743 1263
rect 5789 1217 5811 1263
rect -5811 1139 5811 1217
rect -5811 1093 -5789 1139
rect -5743 1093 -5665 1139
rect -5619 1093 -5541 1139
rect -5495 1093 -5417 1139
rect -5371 1093 -5293 1139
rect -5247 1093 -5169 1139
rect -5123 1093 -5045 1139
rect -4999 1093 -4921 1139
rect -4875 1093 -4797 1139
rect -4751 1093 -4673 1139
rect -4627 1093 -4549 1139
rect -4503 1093 -4425 1139
rect -4379 1093 -4301 1139
rect -4255 1093 -4177 1139
rect -4131 1093 -4053 1139
rect -4007 1093 -3929 1139
rect -3883 1093 -3805 1139
rect -3759 1093 -3681 1139
rect -3635 1093 -3557 1139
rect -3511 1093 -3433 1139
rect -3387 1093 -3309 1139
rect -3263 1093 -3185 1139
rect -3139 1093 -3061 1139
rect -3015 1093 -2937 1139
rect -2891 1093 -2813 1139
rect -2767 1093 -2689 1139
rect -2643 1093 -2565 1139
rect -2519 1093 -2441 1139
rect -2395 1093 -2317 1139
rect -2271 1093 -2193 1139
rect -2147 1093 -2069 1139
rect -2023 1093 -1945 1139
rect -1899 1093 -1821 1139
rect -1775 1093 -1697 1139
rect -1651 1093 -1573 1139
rect -1527 1093 -1449 1139
rect -1403 1093 -1325 1139
rect -1279 1093 -1201 1139
rect -1155 1093 -1077 1139
rect -1031 1093 -953 1139
rect -907 1093 -829 1139
rect -783 1093 -705 1139
rect -659 1093 -581 1139
rect -535 1093 -457 1139
rect -411 1093 -333 1139
rect -287 1093 -209 1139
rect -163 1093 -85 1139
rect -39 1093 39 1139
rect 85 1093 163 1139
rect 209 1093 287 1139
rect 333 1093 411 1139
rect 457 1093 535 1139
rect 581 1093 659 1139
rect 705 1093 783 1139
rect 829 1093 907 1139
rect 953 1093 1031 1139
rect 1077 1093 1155 1139
rect 1201 1093 1279 1139
rect 1325 1093 1403 1139
rect 1449 1093 1527 1139
rect 1573 1093 1651 1139
rect 1697 1093 1775 1139
rect 1821 1093 1899 1139
rect 1945 1093 2023 1139
rect 2069 1093 2147 1139
rect 2193 1093 2271 1139
rect 2317 1093 2395 1139
rect 2441 1093 2519 1139
rect 2565 1093 2643 1139
rect 2689 1093 2767 1139
rect 2813 1093 2891 1139
rect 2937 1093 3015 1139
rect 3061 1093 3139 1139
rect 3185 1093 3263 1139
rect 3309 1093 3387 1139
rect 3433 1093 3511 1139
rect 3557 1093 3635 1139
rect 3681 1093 3759 1139
rect 3805 1093 3883 1139
rect 3929 1093 4007 1139
rect 4053 1093 4131 1139
rect 4177 1093 4255 1139
rect 4301 1093 4379 1139
rect 4425 1093 4503 1139
rect 4549 1093 4627 1139
rect 4673 1093 4751 1139
rect 4797 1093 4875 1139
rect 4921 1093 4999 1139
rect 5045 1093 5123 1139
rect 5169 1093 5247 1139
rect 5293 1093 5371 1139
rect 5417 1093 5495 1139
rect 5541 1093 5619 1139
rect 5665 1093 5743 1139
rect 5789 1093 5811 1139
rect -5811 1015 5811 1093
rect -5811 969 -5789 1015
rect -5743 969 -5665 1015
rect -5619 969 -5541 1015
rect -5495 969 -5417 1015
rect -5371 969 -5293 1015
rect -5247 969 -5169 1015
rect -5123 969 -5045 1015
rect -4999 969 -4921 1015
rect -4875 969 -4797 1015
rect -4751 969 -4673 1015
rect -4627 969 -4549 1015
rect -4503 969 -4425 1015
rect -4379 969 -4301 1015
rect -4255 969 -4177 1015
rect -4131 969 -4053 1015
rect -4007 969 -3929 1015
rect -3883 969 -3805 1015
rect -3759 969 -3681 1015
rect -3635 969 -3557 1015
rect -3511 969 -3433 1015
rect -3387 969 -3309 1015
rect -3263 969 -3185 1015
rect -3139 969 -3061 1015
rect -3015 969 -2937 1015
rect -2891 969 -2813 1015
rect -2767 969 -2689 1015
rect -2643 969 -2565 1015
rect -2519 969 -2441 1015
rect -2395 969 -2317 1015
rect -2271 969 -2193 1015
rect -2147 969 -2069 1015
rect -2023 969 -1945 1015
rect -1899 969 -1821 1015
rect -1775 969 -1697 1015
rect -1651 969 -1573 1015
rect -1527 969 -1449 1015
rect -1403 969 -1325 1015
rect -1279 969 -1201 1015
rect -1155 969 -1077 1015
rect -1031 969 -953 1015
rect -907 969 -829 1015
rect -783 969 -705 1015
rect -659 969 -581 1015
rect -535 969 -457 1015
rect -411 969 -333 1015
rect -287 969 -209 1015
rect -163 969 -85 1015
rect -39 969 39 1015
rect 85 969 163 1015
rect 209 969 287 1015
rect 333 969 411 1015
rect 457 969 535 1015
rect 581 969 659 1015
rect 705 969 783 1015
rect 829 969 907 1015
rect 953 969 1031 1015
rect 1077 969 1155 1015
rect 1201 969 1279 1015
rect 1325 969 1403 1015
rect 1449 969 1527 1015
rect 1573 969 1651 1015
rect 1697 969 1775 1015
rect 1821 969 1899 1015
rect 1945 969 2023 1015
rect 2069 969 2147 1015
rect 2193 969 2271 1015
rect 2317 969 2395 1015
rect 2441 969 2519 1015
rect 2565 969 2643 1015
rect 2689 969 2767 1015
rect 2813 969 2891 1015
rect 2937 969 3015 1015
rect 3061 969 3139 1015
rect 3185 969 3263 1015
rect 3309 969 3387 1015
rect 3433 969 3511 1015
rect 3557 969 3635 1015
rect 3681 969 3759 1015
rect 3805 969 3883 1015
rect 3929 969 4007 1015
rect 4053 969 4131 1015
rect 4177 969 4255 1015
rect 4301 969 4379 1015
rect 4425 969 4503 1015
rect 4549 969 4627 1015
rect 4673 969 4751 1015
rect 4797 969 4875 1015
rect 4921 969 4999 1015
rect 5045 969 5123 1015
rect 5169 969 5247 1015
rect 5293 969 5371 1015
rect 5417 969 5495 1015
rect 5541 969 5619 1015
rect 5665 969 5743 1015
rect 5789 969 5811 1015
rect -5811 891 5811 969
rect -5811 845 -5789 891
rect -5743 845 -5665 891
rect -5619 845 -5541 891
rect -5495 845 -5417 891
rect -5371 845 -5293 891
rect -5247 845 -5169 891
rect -5123 845 -5045 891
rect -4999 845 -4921 891
rect -4875 845 -4797 891
rect -4751 845 -4673 891
rect -4627 845 -4549 891
rect -4503 845 -4425 891
rect -4379 845 -4301 891
rect -4255 845 -4177 891
rect -4131 845 -4053 891
rect -4007 845 -3929 891
rect -3883 845 -3805 891
rect -3759 845 -3681 891
rect -3635 845 -3557 891
rect -3511 845 -3433 891
rect -3387 845 -3309 891
rect -3263 845 -3185 891
rect -3139 845 -3061 891
rect -3015 845 -2937 891
rect -2891 845 -2813 891
rect -2767 845 -2689 891
rect -2643 845 -2565 891
rect -2519 845 -2441 891
rect -2395 845 -2317 891
rect -2271 845 -2193 891
rect -2147 845 -2069 891
rect -2023 845 -1945 891
rect -1899 845 -1821 891
rect -1775 845 -1697 891
rect -1651 845 -1573 891
rect -1527 845 -1449 891
rect -1403 845 -1325 891
rect -1279 845 -1201 891
rect -1155 845 -1077 891
rect -1031 845 -953 891
rect -907 845 -829 891
rect -783 845 -705 891
rect -659 845 -581 891
rect -535 845 -457 891
rect -411 845 -333 891
rect -287 845 -209 891
rect -163 845 -85 891
rect -39 845 39 891
rect 85 845 163 891
rect 209 845 287 891
rect 333 845 411 891
rect 457 845 535 891
rect 581 845 659 891
rect 705 845 783 891
rect 829 845 907 891
rect 953 845 1031 891
rect 1077 845 1155 891
rect 1201 845 1279 891
rect 1325 845 1403 891
rect 1449 845 1527 891
rect 1573 845 1651 891
rect 1697 845 1775 891
rect 1821 845 1899 891
rect 1945 845 2023 891
rect 2069 845 2147 891
rect 2193 845 2271 891
rect 2317 845 2395 891
rect 2441 845 2519 891
rect 2565 845 2643 891
rect 2689 845 2767 891
rect 2813 845 2891 891
rect 2937 845 3015 891
rect 3061 845 3139 891
rect 3185 845 3263 891
rect 3309 845 3387 891
rect 3433 845 3511 891
rect 3557 845 3635 891
rect 3681 845 3759 891
rect 3805 845 3883 891
rect 3929 845 4007 891
rect 4053 845 4131 891
rect 4177 845 4255 891
rect 4301 845 4379 891
rect 4425 845 4503 891
rect 4549 845 4627 891
rect 4673 845 4751 891
rect 4797 845 4875 891
rect 4921 845 4999 891
rect 5045 845 5123 891
rect 5169 845 5247 891
rect 5293 845 5371 891
rect 5417 845 5495 891
rect 5541 845 5619 891
rect 5665 845 5743 891
rect 5789 845 5811 891
rect -5811 767 5811 845
rect -5811 721 -5789 767
rect -5743 721 -5665 767
rect -5619 721 -5541 767
rect -5495 721 -5417 767
rect -5371 721 -5293 767
rect -5247 721 -5169 767
rect -5123 721 -5045 767
rect -4999 721 -4921 767
rect -4875 721 -4797 767
rect -4751 721 -4673 767
rect -4627 721 -4549 767
rect -4503 721 -4425 767
rect -4379 721 -4301 767
rect -4255 721 -4177 767
rect -4131 721 -4053 767
rect -4007 721 -3929 767
rect -3883 721 -3805 767
rect -3759 721 -3681 767
rect -3635 721 -3557 767
rect -3511 721 -3433 767
rect -3387 721 -3309 767
rect -3263 721 -3185 767
rect -3139 721 -3061 767
rect -3015 721 -2937 767
rect -2891 721 -2813 767
rect -2767 721 -2689 767
rect -2643 721 -2565 767
rect -2519 721 -2441 767
rect -2395 721 -2317 767
rect -2271 721 -2193 767
rect -2147 721 -2069 767
rect -2023 721 -1945 767
rect -1899 721 -1821 767
rect -1775 721 -1697 767
rect -1651 721 -1573 767
rect -1527 721 -1449 767
rect -1403 721 -1325 767
rect -1279 721 -1201 767
rect -1155 721 -1077 767
rect -1031 721 -953 767
rect -907 721 -829 767
rect -783 721 -705 767
rect -659 721 -581 767
rect -535 721 -457 767
rect -411 721 -333 767
rect -287 721 -209 767
rect -163 721 -85 767
rect -39 721 39 767
rect 85 721 163 767
rect 209 721 287 767
rect 333 721 411 767
rect 457 721 535 767
rect 581 721 659 767
rect 705 721 783 767
rect 829 721 907 767
rect 953 721 1031 767
rect 1077 721 1155 767
rect 1201 721 1279 767
rect 1325 721 1403 767
rect 1449 721 1527 767
rect 1573 721 1651 767
rect 1697 721 1775 767
rect 1821 721 1899 767
rect 1945 721 2023 767
rect 2069 721 2147 767
rect 2193 721 2271 767
rect 2317 721 2395 767
rect 2441 721 2519 767
rect 2565 721 2643 767
rect 2689 721 2767 767
rect 2813 721 2891 767
rect 2937 721 3015 767
rect 3061 721 3139 767
rect 3185 721 3263 767
rect 3309 721 3387 767
rect 3433 721 3511 767
rect 3557 721 3635 767
rect 3681 721 3759 767
rect 3805 721 3883 767
rect 3929 721 4007 767
rect 4053 721 4131 767
rect 4177 721 4255 767
rect 4301 721 4379 767
rect 4425 721 4503 767
rect 4549 721 4627 767
rect 4673 721 4751 767
rect 4797 721 4875 767
rect 4921 721 4999 767
rect 5045 721 5123 767
rect 5169 721 5247 767
rect 5293 721 5371 767
rect 5417 721 5495 767
rect 5541 721 5619 767
rect 5665 721 5743 767
rect 5789 721 5811 767
rect -5811 643 5811 721
rect -5811 597 -5789 643
rect -5743 597 -5665 643
rect -5619 597 -5541 643
rect -5495 597 -5417 643
rect -5371 597 -5293 643
rect -5247 597 -5169 643
rect -5123 597 -5045 643
rect -4999 597 -4921 643
rect -4875 597 -4797 643
rect -4751 597 -4673 643
rect -4627 597 -4549 643
rect -4503 597 -4425 643
rect -4379 597 -4301 643
rect -4255 597 -4177 643
rect -4131 597 -4053 643
rect -4007 597 -3929 643
rect -3883 597 -3805 643
rect -3759 597 -3681 643
rect -3635 597 -3557 643
rect -3511 597 -3433 643
rect -3387 597 -3309 643
rect -3263 597 -3185 643
rect -3139 597 -3061 643
rect -3015 597 -2937 643
rect -2891 597 -2813 643
rect -2767 597 -2689 643
rect -2643 597 -2565 643
rect -2519 597 -2441 643
rect -2395 597 -2317 643
rect -2271 597 -2193 643
rect -2147 597 -2069 643
rect -2023 597 -1945 643
rect -1899 597 -1821 643
rect -1775 597 -1697 643
rect -1651 597 -1573 643
rect -1527 597 -1449 643
rect -1403 597 -1325 643
rect -1279 597 -1201 643
rect -1155 597 -1077 643
rect -1031 597 -953 643
rect -907 597 -829 643
rect -783 597 -705 643
rect -659 597 -581 643
rect -535 597 -457 643
rect -411 597 -333 643
rect -287 597 -209 643
rect -163 597 -85 643
rect -39 597 39 643
rect 85 597 163 643
rect 209 597 287 643
rect 333 597 411 643
rect 457 597 535 643
rect 581 597 659 643
rect 705 597 783 643
rect 829 597 907 643
rect 953 597 1031 643
rect 1077 597 1155 643
rect 1201 597 1279 643
rect 1325 597 1403 643
rect 1449 597 1527 643
rect 1573 597 1651 643
rect 1697 597 1775 643
rect 1821 597 1899 643
rect 1945 597 2023 643
rect 2069 597 2147 643
rect 2193 597 2271 643
rect 2317 597 2395 643
rect 2441 597 2519 643
rect 2565 597 2643 643
rect 2689 597 2767 643
rect 2813 597 2891 643
rect 2937 597 3015 643
rect 3061 597 3139 643
rect 3185 597 3263 643
rect 3309 597 3387 643
rect 3433 597 3511 643
rect 3557 597 3635 643
rect 3681 597 3759 643
rect 3805 597 3883 643
rect 3929 597 4007 643
rect 4053 597 4131 643
rect 4177 597 4255 643
rect 4301 597 4379 643
rect 4425 597 4503 643
rect 4549 597 4627 643
rect 4673 597 4751 643
rect 4797 597 4875 643
rect 4921 597 4999 643
rect 5045 597 5123 643
rect 5169 597 5247 643
rect 5293 597 5371 643
rect 5417 597 5495 643
rect 5541 597 5619 643
rect 5665 597 5743 643
rect 5789 597 5811 643
rect -5811 519 5811 597
rect -5811 473 -5789 519
rect -5743 473 -5665 519
rect -5619 473 -5541 519
rect -5495 473 -5417 519
rect -5371 473 -5293 519
rect -5247 473 -5169 519
rect -5123 473 -5045 519
rect -4999 473 -4921 519
rect -4875 473 -4797 519
rect -4751 473 -4673 519
rect -4627 473 -4549 519
rect -4503 473 -4425 519
rect -4379 473 -4301 519
rect -4255 473 -4177 519
rect -4131 473 -4053 519
rect -4007 473 -3929 519
rect -3883 473 -3805 519
rect -3759 473 -3681 519
rect -3635 473 -3557 519
rect -3511 473 -3433 519
rect -3387 473 -3309 519
rect -3263 473 -3185 519
rect -3139 473 -3061 519
rect -3015 473 -2937 519
rect -2891 473 -2813 519
rect -2767 473 -2689 519
rect -2643 473 -2565 519
rect -2519 473 -2441 519
rect -2395 473 -2317 519
rect -2271 473 -2193 519
rect -2147 473 -2069 519
rect -2023 473 -1945 519
rect -1899 473 -1821 519
rect -1775 473 -1697 519
rect -1651 473 -1573 519
rect -1527 473 -1449 519
rect -1403 473 -1325 519
rect -1279 473 -1201 519
rect -1155 473 -1077 519
rect -1031 473 -953 519
rect -907 473 -829 519
rect -783 473 -705 519
rect -659 473 -581 519
rect -535 473 -457 519
rect -411 473 -333 519
rect -287 473 -209 519
rect -163 473 -85 519
rect -39 473 39 519
rect 85 473 163 519
rect 209 473 287 519
rect 333 473 411 519
rect 457 473 535 519
rect 581 473 659 519
rect 705 473 783 519
rect 829 473 907 519
rect 953 473 1031 519
rect 1077 473 1155 519
rect 1201 473 1279 519
rect 1325 473 1403 519
rect 1449 473 1527 519
rect 1573 473 1651 519
rect 1697 473 1775 519
rect 1821 473 1899 519
rect 1945 473 2023 519
rect 2069 473 2147 519
rect 2193 473 2271 519
rect 2317 473 2395 519
rect 2441 473 2519 519
rect 2565 473 2643 519
rect 2689 473 2767 519
rect 2813 473 2891 519
rect 2937 473 3015 519
rect 3061 473 3139 519
rect 3185 473 3263 519
rect 3309 473 3387 519
rect 3433 473 3511 519
rect 3557 473 3635 519
rect 3681 473 3759 519
rect 3805 473 3883 519
rect 3929 473 4007 519
rect 4053 473 4131 519
rect 4177 473 4255 519
rect 4301 473 4379 519
rect 4425 473 4503 519
rect 4549 473 4627 519
rect 4673 473 4751 519
rect 4797 473 4875 519
rect 4921 473 4999 519
rect 5045 473 5123 519
rect 5169 473 5247 519
rect 5293 473 5371 519
rect 5417 473 5495 519
rect 5541 473 5619 519
rect 5665 473 5743 519
rect 5789 473 5811 519
rect -5811 395 5811 473
rect -5811 349 -5789 395
rect -5743 349 -5665 395
rect -5619 349 -5541 395
rect -5495 349 -5417 395
rect -5371 349 -5293 395
rect -5247 349 -5169 395
rect -5123 349 -5045 395
rect -4999 349 -4921 395
rect -4875 349 -4797 395
rect -4751 349 -4673 395
rect -4627 349 -4549 395
rect -4503 349 -4425 395
rect -4379 349 -4301 395
rect -4255 349 -4177 395
rect -4131 349 -4053 395
rect -4007 349 -3929 395
rect -3883 349 -3805 395
rect -3759 349 -3681 395
rect -3635 349 -3557 395
rect -3511 349 -3433 395
rect -3387 349 -3309 395
rect -3263 349 -3185 395
rect -3139 349 -3061 395
rect -3015 349 -2937 395
rect -2891 349 -2813 395
rect -2767 349 -2689 395
rect -2643 349 -2565 395
rect -2519 349 -2441 395
rect -2395 349 -2317 395
rect -2271 349 -2193 395
rect -2147 349 -2069 395
rect -2023 349 -1945 395
rect -1899 349 -1821 395
rect -1775 349 -1697 395
rect -1651 349 -1573 395
rect -1527 349 -1449 395
rect -1403 349 -1325 395
rect -1279 349 -1201 395
rect -1155 349 -1077 395
rect -1031 349 -953 395
rect -907 349 -829 395
rect -783 349 -705 395
rect -659 349 -581 395
rect -535 349 -457 395
rect -411 349 -333 395
rect -287 349 -209 395
rect -163 349 -85 395
rect -39 349 39 395
rect 85 349 163 395
rect 209 349 287 395
rect 333 349 411 395
rect 457 349 535 395
rect 581 349 659 395
rect 705 349 783 395
rect 829 349 907 395
rect 953 349 1031 395
rect 1077 349 1155 395
rect 1201 349 1279 395
rect 1325 349 1403 395
rect 1449 349 1527 395
rect 1573 349 1651 395
rect 1697 349 1775 395
rect 1821 349 1899 395
rect 1945 349 2023 395
rect 2069 349 2147 395
rect 2193 349 2271 395
rect 2317 349 2395 395
rect 2441 349 2519 395
rect 2565 349 2643 395
rect 2689 349 2767 395
rect 2813 349 2891 395
rect 2937 349 3015 395
rect 3061 349 3139 395
rect 3185 349 3263 395
rect 3309 349 3387 395
rect 3433 349 3511 395
rect 3557 349 3635 395
rect 3681 349 3759 395
rect 3805 349 3883 395
rect 3929 349 4007 395
rect 4053 349 4131 395
rect 4177 349 4255 395
rect 4301 349 4379 395
rect 4425 349 4503 395
rect 4549 349 4627 395
rect 4673 349 4751 395
rect 4797 349 4875 395
rect 4921 349 4999 395
rect 5045 349 5123 395
rect 5169 349 5247 395
rect 5293 349 5371 395
rect 5417 349 5495 395
rect 5541 349 5619 395
rect 5665 349 5743 395
rect 5789 349 5811 395
rect -5811 271 5811 349
rect -5811 225 -5789 271
rect -5743 225 -5665 271
rect -5619 225 -5541 271
rect -5495 225 -5417 271
rect -5371 225 -5293 271
rect -5247 225 -5169 271
rect -5123 225 -5045 271
rect -4999 225 -4921 271
rect -4875 225 -4797 271
rect -4751 225 -4673 271
rect -4627 225 -4549 271
rect -4503 225 -4425 271
rect -4379 225 -4301 271
rect -4255 225 -4177 271
rect -4131 225 -4053 271
rect -4007 225 -3929 271
rect -3883 225 -3805 271
rect -3759 225 -3681 271
rect -3635 225 -3557 271
rect -3511 225 -3433 271
rect -3387 225 -3309 271
rect -3263 225 -3185 271
rect -3139 225 -3061 271
rect -3015 225 -2937 271
rect -2891 225 -2813 271
rect -2767 225 -2689 271
rect -2643 225 -2565 271
rect -2519 225 -2441 271
rect -2395 225 -2317 271
rect -2271 225 -2193 271
rect -2147 225 -2069 271
rect -2023 225 -1945 271
rect -1899 225 -1821 271
rect -1775 225 -1697 271
rect -1651 225 -1573 271
rect -1527 225 -1449 271
rect -1403 225 -1325 271
rect -1279 225 -1201 271
rect -1155 225 -1077 271
rect -1031 225 -953 271
rect -907 225 -829 271
rect -783 225 -705 271
rect -659 225 -581 271
rect -535 225 -457 271
rect -411 225 -333 271
rect -287 225 -209 271
rect -163 225 -85 271
rect -39 225 39 271
rect 85 225 163 271
rect 209 225 287 271
rect 333 225 411 271
rect 457 225 535 271
rect 581 225 659 271
rect 705 225 783 271
rect 829 225 907 271
rect 953 225 1031 271
rect 1077 225 1155 271
rect 1201 225 1279 271
rect 1325 225 1403 271
rect 1449 225 1527 271
rect 1573 225 1651 271
rect 1697 225 1775 271
rect 1821 225 1899 271
rect 1945 225 2023 271
rect 2069 225 2147 271
rect 2193 225 2271 271
rect 2317 225 2395 271
rect 2441 225 2519 271
rect 2565 225 2643 271
rect 2689 225 2767 271
rect 2813 225 2891 271
rect 2937 225 3015 271
rect 3061 225 3139 271
rect 3185 225 3263 271
rect 3309 225 3387 271
rect 3433 225 3511 271
rect 3557 225 3635 271
rect 3681 225 3759 271
rect 3805 225 3883 271
rect 3929 225 4007 271
rect 4053 225 4131 271
rect 4177 225 4255 271
rect 4301 225 4379 271
rect 4425 225 4503 271
rect 4549 225 4627 271
rect 4673 225 4751 271
rect 4797 225 4875 271
rect 4921 225 4999 271
rect 5045 225 5123 271
rect 5169 225 5247 271
rect 5293 225 5371 271
rect 5417 225 5495 271
rect 5541 225 5619 271
rect 5665 225 5743 271
rect 5789 225 5811 271
rect -5811 147 5811 225
rect -5811 101 -5789 147
rect -5743 101 -5665 147
rect -5619 101 -5541 147
rect -5495 101 -5417 147
rect -5371 101 -5293 147
rect -5247 101 -5169 147
rect -5123 101 -5045 147
rect -4999 101 -4921 147
rect -4875 101 -4797 147
rect -4751 101 -4673 147
rect -4627 101 -4549 147
rect -4503 101 -4425 147
rect -4379 101 -4301 147
rect -4255 101 -4177 147
rect -4131 101 -4053 147
rect -4007 101 -3929 147
rect -3883 101 -3805 147
rect -3759 101 -3681 147
rect -3635 101 -3557 147
rect -3511 101 -3433 147
rect -3387 101 -3309 147
rect -3263 101 -3185 147
rect -3139 101 -3061 147
rect -3015 101 -2937 147
rect -2891 101 -2813 147
rect -2767 101 -2689 147
rect -2643 101 -2565 147
rect -2519 101 -2441 147
rect -2395 101 -2317 147
rect -2271 101 -2193 147
rect -2147 101 -2069 147
rect -2023 101 -1945 147
rect -1899 101 -1821 147
rect -1775 101 -1697 147
rect -1651 101 -1573 147
rect -1527 101 -1449 147
rect -1403 101 -1325 147
rect -1279 101 -1201 147
rect -1155 101 -1077 147
rect -1031 101 -953 147
rect -907 101 -829 147
rect -783 101 -705 147
rect -659 101 -581 147
rect -535 101 -457 147
rect -411 101 -333 147
rect -287 101 -209 147
rect -163 101 -85 147
rect -39 101 39 147
rect 85 101 163 147
rect 209 101 287 147
rect 333 101 411 147
rect 457 101 535 147
rect 581 101 659 147
rect 705 101 783 147
rect 829 101 907 147
rect 953 101 1031 147
rect 1077 101 1155 147
rect 1201 101 1279 147
rect 1325 101 1403 147
rect 1449 101 1527 147
rect 1573 101 1651 147
rect 1697 101 1775 147
rect 1821 101 1899 147
rect 1945 101 2023 147
rect 2069 101 2147 147
rect 2193 101 2271 147
rect 2317 101 2395 147
rect 2441 101 2519 147
rect 2565 101 2643 147
rect 2689 101 2767 147
rect 2813 101 2891 147
rect 2937 101 3015 147
rect 3061 101 3139 147
rect 3185 101 3263 147
rect 3309 101 3387 147
rect 3433 101 3511 147
rect 3557 101 3635 147
rect 3681 101 3759 147
rect 3805 101 3883 147
rect 3929 101 4007 147
rect 4053 101 4131 147
rect 4177 101 4255 147
rect 4301 101 4379 147
rect 4425 101 4503 147
rect 4549 101 4627 147
rect 4673 101 4751 147
rect 4797 101 4875 147
rect 4921 101 4999 147
rect 5045 101 5123 147
rect 5169 101 5247 147
rect 5293 101 5371 147
rect 5417 101 5495 147
rect 5541 101 5619 147
rect 5665 101 5743 147
rect 5789 101 5811 147
rect -5811 23 5811 101
rect -5811 -23 -5789 23
rect -5743 -23 -5665 23
rect -5619 -23 -5541 23
rect -5495 -23 -5417 23
rect -5371 -23 -5293 23
rect -5247 -23 -5169 23
rect -5123 -23 -5045 23
rect -4999 -23 -4921 23
rect -4875 -23 -4797 23
rect -4751 -23 -4673 23
rect -4627 -23 -4549 23
rect -4503 -23 -4425 23
rect -4379 -23 -4301 23
rect -4255 -23 -4177 23
rect -4131 -23 -4053 23
rect -4007 -23 -3929 23
rect -3883 -23 -3805 23
rect -3759 -23 -3681 23
rect -3635 -23 -3557 23
rect -3511 -23 -3433 23
rect -3387 -23 -3309 23
rect -3263 -23 -3185 23
rect -3139 -23 -3061 23
rect -3015 -23 -2937 23
rect -2891 -23 -2813 23
rect -2767 -23 -2689 23
rect -2643 -23 -2565 23
rect -2519 -23 -2441 23
rect -2395 -23 -2317 23
rect -2271 -23 -2193 23
rect -2147 -23 -2069 23
rect -2023 -23 -1945 23
rect -1899 -23 -1821 23
rect -1775 -23 -1697 23
rect -1651 -23 -1573 23
rect -1527 -23 -1449 23
rect -1403 -23 -1325 23
rect -1279 -23 -1201 23
rect -1155 -23 -1077 23
rect -1031 -23 -953 23
rect -907 -23 -829 23
rect -783 -23 -705 23
rect -659 -23 -581 23
rect -535 -23 -457 23
rect -411 -23 -333 23
rect -287 -23 -209 23
rect -163 -23 -85 23
rect -39 -23 39 23
rect 85 -23 163 23
rect 209 -23 287 23
rect 333 -23 411 23
rect 457 -23 535 23
rect 581 -23 659 23
rect 705 -23 783 23
rect 829 -23 907 23
rect 953 -23 1031 23
rect 1077 -23 1155 23
rect 1201 -23 1279 23
rect 1325 -23 1403 23
rect 1449 -23 1527 23
rect 1573 -23 1651 23
rect 1697 -23 1775 23
rect 1821 -23 1899 23
rect 1945 -23 2023 23
rect 2069 -23 2147 23
rect 2193 -23 2271 23
rect 2317 -23 2395 23
rect 2441 -23 2519 23
rect 2565 -23 2643 23
rect 2689 -23 2767 23
rect 2813 -23 2891 23
rect 2937 -23 3015 23
rect 3061 -23 3139 23
rect 3185 -23 3263 23
rect 3309 -23 3387 23
rect 3433 -23 3511 23
rect 3557 -23 3635 23
rect 3681 -23 3759 23
rect 3805 -23 3883 23
rect 3929 -23 4007 23
rect 4053 -23 4131 23
rect 4177 -23 4255 23
rect 4301 -23 4379 23
rect 4425 -23 4503 23
rect 4549 -23 4627 23
rect 4673 -23 4751 23
rect 4797 -23 4875 23
rect 4921 -23 4999 23
rect 5045 -23 5123 23
rect 5169 -23 5247 23
rect 5293 -23 5371 23
rect 5417 -23 5495 23
rect 5541 -23 5619 23
rect 5665 -23 5743 23
rect 5789 -23 5811 23
rect -5811 -101 5811 -23
rect -5811 -147 -5789 -101
rect -5743 -147 -5665 -101
rect -5619 -147 -5541 -101
rect -5495 -147 -5417 -101
rect -5371 -147 -5293 -101
rect -5247 -147 -5169 -101
rect -5123 -147 -5045 -101
rect -4999 -147 -4921 -101
rect -4875 -147 -4797 -101
rect -4751 -147 -4673 -101
rect -4627 -147 -4549 -101
rect -4503 -147 -4425 -101
rect -4379 -147 -4301 -101
rect -4255 -147 -4177 -101
rect -4131 -147 -4053 -101
rect -4007 -147 -3929 -101
rect -3883 -147 -3805 -101
rect -3759 -147 -3681 -101
rect -3635 -147 -3557 -101
rect -3511 -147 -3433 -101
rect -3387 -147 -3309 -101
rect -3263 -147 -3185 -101
rect -3139 -147 -3061 -101
rect -3015 -147 -2937 -101
rect -2891 -147 -2813 -101
rect -2767 -147 -2689 -101
rect -2643 -147 -2565 -101
rect -2519 -147 -2441 -101
rect -2395 -147 -2317 -101
rect -2271 -147 -2193 -101
rect -2147 -147 -2069 -101
rect -2023 -147 -1945 -101
rect -1899 -147 -1821 -101
rect -1775 -147 -1697 -101
rect -1651 -147 -1573 -101
rect -1527 -147 -1449 -101
rect -1403 -147 -1325 -101
rect -1279 -147 -1201 -101
rect -1155 -147 -1077 -101
rect -1031 -147 -953 -101
rect -907 -147 -829 -101
rect -783 -147 -705 -101
rect -659 -147 -581 -101
rect -535 -147 -457 -101
rect -411 -147 -333 -101
rect -287 -147 -209 -101
rect -163 -147 -85 -101
rect -39 -147 39 -101
rect 85 -147 163 -101
rect 209 -147 287 -101
rect 333 -147 411 -101
rect 457 -147 535 -101
rect 581 -147 659 -101
rect 705 -147 783 -101
rect 829 -147 907 -101
rect 953 -147 1031 -101
rect 1077 -147 1155 -101
rect 1201 -147 1279 -101
rect 1325 -147 1403 -101
rect 1449 -147 1527 -101
rect 1573 -147 1651 -101
rect 1697 -147 1775 -101
rect 1821 -147 1899 -101
rect 1945 -147 2023 -101
rect 2069 -147 2147 -101
rect 2193 -147 2271 -101
rect 2317 -147 2395 -101
rect 2441 -147 2519 -101
rect 2565 -147 2643 -101
rect 2689 -147 2767 -101
rect 2813 -147 2891 -101
rect 2937 -147 3015 -101
rect 3061 -147 3139 -101
rect 3185 -147 3263 -101
rect 3309 -147 3387 -101
rect 3433 -147 3511 -101
rect 3557 -147 3635 -101
rect 3681 -147 3759 -101
rect 3805 -147 3883 -101
rect 3929 -147 4007 -101
rect 4053 -147 4131 -101
rect 4177 -147 4255 -101
rect 4301 -147 4379 -101
rect 4425 -147 4503 -101
rect 4549 -147 4627 -101
rect 4673 -147 4751 -101
rect 4797 -147 4875 -101
rect 4921 -147 4999 -101
rect 5045 -147 5123 -101
rect 5169 -147 5247 -101
rect 5293 -147 5371 -101
rect 5417 -147 5495 -101
rect 5541 -147 5619 -101
rect 5665 -147 5743 -101
rect 5789 -147 5811 -101
rect -5811 -225 5811 -147
rect -5811 -271 -5789 -225
rect -5743 -271 -5665 -225
rect -5619 -271 -5541 -225
rect -5495 -271 -5417 -225
rect -5371 -271 -5293 -225
rect -5247 -271 -5169 -225
rect -5123 -271 -5045 -225
rect -4999 -271 -4921 -225
rect -4875 -271 -4797 -225
rect -4751 -271 -4673 -225
rect -4627 -271 -4549 -225
rect -4503 -271 -4425 -225
rect -4379 -271 -4301 -225
rect -4255 -271 -4177 -225
rect -4131 -271 -4053 -225
rect -4007 -271 -3929 -225
rect -3883 -271 -3805 -225
rect -3759 -271 -3681 -225
rect -3635 -271 -3557 -225
rect -3511 -271 -3433 -225
rect -3387 -271 -3309 -225
rect -3263 -271 -3185 -225
rect -3139 -271 -3061 -225
rect -3015 -271 -2937 -225
rect -2891 -271 -2813 -225
rect -2767 -271 -2689 -225
rect -2643 -271 -2565 -225
rect -2519 -271 -2441 -225
rect -2395 -271 -2317 -225
rect -2271 -271 -2193 -225
rect -2147 -271 -2069 -225
rect -2023 -271 -1945 -225
rect -1899 -271 -1821 -225
rect -1775 -271 -1697 -225
rect -1651 -271 -1573 -225
rect -1527 -271 -1449 -225
rect -1403 -271 -1325 -225
rect -1279 -271 -1201 -225
rect -1155 -271 -1077 -225
rect -1031 -271 -953 -225
rect -907 -271 -829 -225
rect -783 -271 -705 -225
rect -659 -271 -581 -225
rect -535 -271 -457 -225
rect -411 -271 -333 -225
rect -287 -271 -209 -225
rect -163 -271 -85 -225
rect -39 -271 39 -225
rect 85 -271 163 -225
rect 209 -271 287 -225
rect 333 -271 411 -225
rect 457 -271 535 -225
rect 581 -271 659 -225
rect 705 -271 783 -225
rect 829 -271 907 -225
rect 953 -271 1031 -225
rect 1077 -271 1155 -225
rect 1201 -271 1279 -225
rect 1325 -271 1403 -225
rect 1449 -271 1527 -225
rect 1573 -271 1651 -225
rect 1697 -271 1775 -225
rect 1821 -271 1899 -225
rect 1945 -271 2023 -225
rect 2069 -271 2147 -225
rect 2193 -271 2271 -225
rect 2317 -271 2395 -225
rect 2441 -271 2519 -225
rect 2565 -271 2643 -225
rect 2689 -271 2767 -225
rect 2813 -271 2891 -225
rect 2937 -271 3015 -225
rect 3061 -271 3139 -225
rect 3185 -271 3263 -225
rect 3309 -271 3387 -225
rect 3433 -271 3511 -225
rect 3557 -271 3635 -225
rect 3681 -271 3759 -225
rect 3805 -271 3883 -225
rect 3929 -271 4007 -225
rect 4053 -271 4131 -225
rect 4177 -271 4255 -225
rect 4301 -271 4379 -225
rect 4425 -271 4503 -225
rect 4549 -271 4627 -225
rect 4673 -271 4751 -225
rect 4797 -271 4875 -225
rect 4921 -271 4999 -225
rect 5045 -271 5123 -225
rect 5169 -271 5247 -225
rect 5293 -271 5371 -225
rect 5417 -271 5495 -225
rect 5541 -271 5619 -225
rect 5665 -271 5743 -225
rect 5789 -271 5811 -225
rect -5811 -349 5811 -271
rect -5811 -395 -5789 -349
rect -5743 -395 -5665 -349
rect -5619 -395 -5541 -349
rect -5495 -395 -5417 -349
rect -5371 -395 -5293 -349
rect -5247 -395 -5169 -349
rect -5123 -395 -5045 -349
rect -4999 -395 -4921 -349
rect -4875 -395 -4797 -349
rect -4751 -395 -4673 -349
rect -4627 -395 -4549 -349
rect -4503 -395 -4425 -349
rect -4379 -395 -4301 -349
rect -4255 -395 -4177 -349
rect -4131 -395 -4053 -349
rect -4007 -395 -3929 -349
rect -3883 -395 -3805 -349
rect -3759 -395 -3681 -349
rect -3635 -395 -3557 -349
rect -3511 -395 -3433 -349
rect -3387 -395 -3309 -349
rect -3263 -395 -3185 -349
rect -3139 -395 -3061 -349
rect -3015 -395 -2937 -349
rect -2891 -395 -2813 -349
rect -2767 -395 -2689 -349
rect -2643 -395 -2565 -349
rect -2519 -395 -2441 -349
rect -2395 -395 -2317 -349
rect -2271 -395 -2193 -349
rect -2147 -395 -2069 -349
rect -2023 -395 -1945 -349
rect -1899 -395 -1821 -349
rect -1775 -395 -1697 -349
rect -1651 -395 -1573 -349
rect -1527 -395 -1449 -349
rect -1403 -395 -1325 -349
rect -1279 -395 -1201 -349
rect -1155 -395 -1077 -349
rect -1031 -395 -953 -349
rect -907 -395 -829 -349
rect -783 -395 -705 -349
rect -659 -395 -581 -349
rect -535 -395 -457 -349
rect -411 -395 -333 -349
rect -287 -395 -209 -349
rect -163 -395 -85 -349
rect -39 -395 39 -349
rect 85 -395 163 -349
rect 209 -395 287 -349
rect 333 -395 411 -349
rect 457 -395 535 -349
rect 581 -395 659 -349
rect 705 -395 783 -349
rect 829 -395 907 -349
rect 953 -395 1031 -349
rect 1077 -395 1155 -349
rect 1201 -395 1279 -349
rect 1325 -395 1403 -349
rect 1449 -395 1527 -349
rect 1573 -395 1651 -349
rect 1697 -395 1775 -349
rect 1821 -395 1899 -349
rect 1945 -395 2023 -349
rect 2069 -395 2147 -349
rect 2193 -395 2271 -349
rect 2317 -395 2395 -349
rect 2441 -395 2519 -349
rect 2565 -395 2643 -349
rect 2689 -395 2767 -349
rect 2813 -395 2891 -349
rect 2937 -395 3015 -349
rect 3061 -395 3139 -349
rect 3185 -395 3263 -349
rect 3309 -395 3387 -349
rect 3433 -395 3511 -349
rect 3557 -395 3635 -349
rect 3681 -395 3759 -349
rect 3805 -395 3883 -349
rect 3929 -395 4007 -349
rect 4053 -395 4131 -349
rect 4177 -395 4255 -349
rect 4301 -395 4379 -349
rect 4425 -395 4503 -349
rect 4549 -395 4627 -349
rect 4673 -395 4751 -349
rect 4797 -395 4875 -349
rect 4921 -395 4999 -349
rect 5045 -395 5123 -349
rect 5169 -395 5247 -349
rect 5293 -395 5371 -349
rect 5417 -395 5495 -349
rect 5541 -395 5619 -349
rect 5665 -395 5743 -349
rect 5789 -395 5811 -349
rect -5811 -473 5811 -395
rect -5811 -519 -5789 -473
rect -5743 -519 -5665 -473
rect -5619 -519 -5541 -473
rect -5495 -519 -5417 -473
rect -5371 -519 -5293 -473
rect -5247 -519 -5169 -473
rect -5123 -519 -5045 -473
rect -4999 -519 -4921 -473
rect -4875 -519 -4797 -473
rect -4751 -519 -4673 -473
rect -4627 -519 -4549 -473
rect -4503 -519 -4425 -473
rect -4379 -519 -4301 -473
rect -4255 -519 -4177 -473
rect -4131 -519 -4053 -473
rect -4007 -519 -3929 -473
rect -3883 -519 -3805 -473
rect -3759 -519 -3681 -473
rect -3635 -519 -3557 -473
rect -3511 -519 -3433 -473
rect -3387 -519 -3309 -473
rect -3263 -519 -3185 -473
rect -3139 -519 -3061 -473
rect -3015 -519 -2937 -473
rect -2891 -519 -2813 -473
rect -2767 -519 -2689 -473
rect -2643 -519 -2565 -473
rect -2519 -519 -2441 -473
rect -2395 -519 -2317 -473
rect -2271 -519 -2193 -473
rect -2147 -519 -2069 -473
rect -2023 -519 -1945 -473
rect -1899 -519 -1821 -473
rect -1775 -519 -1697 -473
rect -1651 -519 -1573 -473
rect -1527 -519 -1449 -473
rect -1403 -519 -1325 -473
rect -1279 -519 -1201 -473
rect -1155 -519 -1077 -473
rect -1031 -519 -953 -473
rect -907 -519 -829 -473
rect -783 -519 -705 -473
rect -659 -519 -581 -473
rect -535 -519 -457 -473
rect -411 -519 -333 -473
rect -287 -519 -209 -473
rect -163 -519 -85 -473
rect -39 -519 39 -473
rect 85 -519 163 -473
rect 209 -519 287 -473
rect 333 -519 411 -473
rect 457 -519 535 -473
rect 581 -519 659 -473
rect 705 -519 783 -473
rect 829 -519 907 -473
rect 953 -519 1031 -473
rect 1077 -519 1155 -473
rect 1201 -519 1279 -473
rect 1325 -519 1403 -473
rect 1449 -519 1527 -473
rect 1573 -519 1651 -473
rect 1697 -519 1775 -473
rect 1821 -519 1899 -473
rect 1945 -519 2023 -473
rect 2069 -519 2147 -473
rect 2193 -519 2271 -473
rect 2317 -519 2395 -473
rect 2441 -519 2519 -473
rect 2565 -519 2643 -473
rect 2689 -519 2767 -473
rect 2813 -519 2891 -473
rect 2937 -519 3015 -473
rect 3061 -519 3139 -473
rect 3185 -519 3263 -473
rect 3309 -519 3387 -473
rect 3433 -519 3511 -473
rect 3557 -519 3635 -473
rect 3681 -519 3759 -473
rect 3805 -519 3883 -473
rect 3929 -519 4007 -473
rect 4053 -519 4131 -473
rect 4177 -519 4255 -473
rect 4301 -519 4379 -473
rect 4425 -519 4503 -473
rect 4549 -519 4627 -473
rect 4673 -519 4751 -473
rect 4797 -519 4875 -473
rect 4921 -519 4999 -473
rect 5045 -519 5123 -473
rect 5169 -519 5247 -473
rect 5293 -519 5371 -473
rect 5417 -519 5495 -473
rect 5541 -519 5619 -473
rect 5665 -519 5743 -473
rect 5789 -519 5811 -473
rect -5811 -597 5811 -519
rect -5811 -643 -5789 -597
rect -5743 -643 -5665 -597
rect -5619 -643 -5541 -597
rect -5495 -643 -5417 -597
rect -5371 -643 -5293 -597
rect -5247 -643 -5169 -597
rect -5123 -643 -5045 -597
rect -4999 -643 -4921 -597
rect -4875 -643 -4797 -597
rect -4751 -643 -4673 -597
rect -4627 -643 -4549 -597
rect -4503 -643 -4425 -597
rect -4379 -643 -4301 -597
rect -4255 -643 -4177 -597
rect -4131 -643 -4053 -597
rect -4007 -643 -3929 -597
rect -3883 -643 -3805 -597
rect -3759 -643 -3681 -597
rect -3635 -643 -3557 -597
rect -3511 -643 -3433 -597
rect -3387 -643 -3309 -597
rect -3263 -643 -3185 -597
rect -3139 -643 -3061 -597
rect -3015 -643 -2937 -597
rect -2891 -643 -2813 -597
rect -2767 -643 -2689 -597
rect -2643 -643 -2565 -597
rect -2519 -643 -2441 -597
rect -2395 -643 -2317 -597
rect -2271 -643 -2193 -597
rect -2147 -643 -2069 -597
rect -2023 -643 -1945 -597
rect -1899 -643 -1821 -597
rect -1775 -643 -1697 -597
rect -1651 -643 -1573 -597
rect -1527 -643 -1449 -597
rect -1403 -643 -1325 -597
rect -1279 -643 -1201 -597
rect -1155 -643 -1077 -597
rect -1031 -643 -953 -597
rect -907 -643 -829 -597
rect -783 -643 -705 -597
rect -659 -643 -581 -597
rect -535 -643 -457 -597
rect -411 -643 -333 -597
rect -287 -643 -209 -597
rect -163 -643 -85 -597
rect -39 -643 39 -597
rect 85 -643 163 -597
rect 209 -643 287 -597
rect 333 -643 411 -597
rect 457 -643 535 -597
rect 581 -643 659 -597
rect 705 -643 783 -597
rect 829 -643 907 -597
rect 953 -643 1031 -597
rect 1077 -643 1155 -597
rect 1201 -643 1279 -597
rect 1325 -643 1403 -597
rect 1449 -643 1527 -597
rect 1573 -643 1651 -597
rect 1697 -643 1775 -597
rect 1821 -643 1899 -597
rect 1945 -643 2023 -597
rect 2069 -643 2147 -597
rect 2193 -643 2271 -597
rect 2317 -643 2395 -597
rect 2441 -643 2519 -597
rect 2565 -643 2643 -597
rect 2689 -643 2767 -597
rect 2813 -643 2891 -597
rect 2937 -643 3015 -597
rect 3061 -643 3139 -597
rect 3185 -643 3263 -597
rect 3309 -643 3387 -597
rect 3433 -643 3511 -597
rect 3557 -643 3635 -597
rect 3681 -643 3759 -597
rect 3805 -643 3883 -597
rect 3929 -643 4007 -597
rect 4053 -643 4131 -597
rect 4177 -643 4255 -597
rect 4301 -643 4379 -597
rect 4425 -643 4503 -597
rect 4549 -643 4627 -597
rect 4673 -643 4751 -597
rect 4797 -643 4875 -597
rect 4921 -643 4999 -597
rect 5045 -643 5123 -597
rect 5169 -643 5247 -597
rect 5293 -643 5371 -597
rect 5417 -643 5495 -597
rect 5541 -643 5619 -597
rect 5665 -643 5743 -597
rect 5789 -643 5811 -597
rect -5811 -721 5811 -643
rect -5811 -767 -5789 -721
rect -5743 -767 -5665 -721
rect -5619 -767 -5541 -721
rect -5495 -767 -5417 -721
rect -5371 -767 -5293 -721
rect -5247 -767 -5169 -721
rect -5123 -767 -5045 -721
rect -4999 -767 -4921 -721
rect -4875 -767 -4797 -721
rect -4751 -767 -4673 -721
rect -4627 -767 -4549 -721
rect -4503 -767 -4425 -721
rect -4379 -767 -4301 -721
rect -4255 -767 -4177 -721
rect -4131 -767 -4053 -721
rect -4007 -767 -3929 -721
rect -3883 -767 -3805 -721
rect -3759 -767 -3681 -721
rect -3635 -767 -3557 -721
rect -3511 -767 -3433 -721
rect -3387 -767 -3309 -721
rect -3263 -767 -3185 -721
rect -3139 -767 -3061 -721
rect -3015 -767 -2937 -721
rect -2891 -767 -2813 -721
rect -2767 -767 -2689 -721
rect -2643 -767 -2565 -721
rect -2519 -767 -2441 -721
rect -2395 -767 -2317 -721
rect -2271 -767 -2193 -721
rect -2147 -767 -2069 -721
rect -2023 -767 -1945 -721
rect -1899 -767 -1821 -721
rect -1775 -767 -1697 -721
rect -1651 -767 -1573 -721
rect -1527 -767 -1449 -721
rect -1403 -767 -1325 -721
rect -1279 -767 -1201 -721
rect -1155 -767 -1077 -721
rect -1031 -767 -953 -721
rect -907 -767 -829 -721
rect -783 -767 -705 -721
rect -659 -767 -581 -721
rect -535 -767 -457 -721
rect -411 -767 -333 -721
rect -287 -767 -209 -721
rect -163 -767 -85 -721
rect -39 -767 39 -721
rect 85 -767 163 -721
rect 209 -767 287 -721
rect 333 -767 411 -721
rect 457 -767 535 -721
rect 581 -767 659 -721
rect 705 -767 783 -721
rect 829 -767 907 -721
rect 953 -767 1031 -721
rect 1077 -767 1155 -721
rect 1201 -767 1279 -721
rect 1325 -767 1403 -721
rect 1449 -767 1527 -721
rect 1573 -767 1651 -721
rect 1697 -767 1775 -721
rect 1821 -767 1899 -721
rect 1945 -767 2023 -721
rect 2069 -767 2147 -721
rect 2193 -767 2271 -721
rect 2317 -767 2395 -721
rect 2441 -767 2519 -721
rect 2565 -767 2643 -721
rect 2689 -767 2767 -721
rect 2813 -767 2891 -721
rect 2937 -767 3015 -721
rect 3061 -767 3139 -721
rect 3185 -767 3263 -721
rect 3309 -767 3387 -721
rect 3433 -767 3511 -721
rect 3557 -767 3635 -721
rect 3681 -767 3759 -721
rect 3805 -767 3883 -721
rect 3929 -767 4007 -721
rect 4053 -767 4131 -721
rect 4177 -767 4255 -721
rect 4301 -767 4379 -721
rect 4425 -767 4503 -721
rect 4549 -767 4627 -721
rect 4673 -767 4751 -721
rect 4797 -767 4875 -721
rect 4921 -767 4999 -721
rect 5045 -767 5123 -721
rect 5169 -767 5247 -721
rect 5293 -767 5371 -721
rect 5417 -767 5495 -721
rect 5541 -767 5619 -721
rect 5665 -767 5743 -721
rect 5789 -767 5811 -721
rect -5811 -845 5811 -767
rect -5811 -891 -5789 -845
rect -5743 -891 -5665 -845
rect -5619 -891 -5541 -845
rect -5495 -891 -5417 -845
rect -5371 -891 -5293 -845
rect -5247 -891 -5169 -845
rect -5123 -891 -5045 -845
rect -4999 -891 -4921 -845
rect -4875 -891 -4797 -845
rect -4751 -891 -4673 -845
rect -4627 -891 -4549 -845
rect -4503 -891 -4425 -845
rect -4379 -891 -4301 -845
rect -4255 -891 -4177 -845
rect -4131 -891 -4053 -845
rect -4007 -891 -3929 -845
rect -3883 -891 -3805 -845
rect -3759 -891 -3681 -845
rect -3635 -891 -3557 -845
rect -3511 -891 -3433 -845
rect -3387 -891 -3309 -845
rect -3263 -891 -3185 -845
rect -3139 -891 -3061 -845
rect -3015 -891 -2937 -845
rect -2891 -891 -2813 -845
rect -2767 -891 -2689 -845
rect -2643 -891 -2565 -845
rect -2519 -891 -2441 -845
rect -2395 -891 -2317 -845
rect -2271 -891 -2193 -845
rect -2147 -891 -2069 -845
rect -2023 -891 -1945 -845
rect -1899 -891 -1821 -845
rect -1775 -891 -1697 -845
rect -1651 -891 -1573 -845
rect -1527 -891 -1449 -845
rect -1403 -891 -1325 -845
rect -1279 -891 -1201 -845
rect -1155 -891 -1077 -845
rect -1031 -891 -953 -845
rect -907 -891 -829 -845
rect -783 -891 -705 -845
rect -659 -891 -581 -845
rect -535 -891 -457 -845
rect -411 -891 -333 -845
rect -287 -891 -209 -845
rect -163 -891 -85 -845
rect -39 -891 39 -845
rect 85 -891 163 -845
rect 209 -891 287 -845
rect 333 -891 411 -845
rect 457 -891 535 -845
rect 581 -891 659 -845
rect 705 -891 783 -845
rect 829 -891 907 -845
rect 953 -891 1031 -845
rect 1077 -891 1155 -845
rect 1201 -891 1279 -845
rect 1325 -891 1403 -845
rect 1449 -891 1527 -845
rect 1573 -891 1651 -845
rect 1697 -891 1775 -845
rect 1821 -891 1899 -845
rect 1945 -891 2023 -845
rect 2069 -891 2147 -845
rect 2193 -891 2271 -845
rect 2317 -891 2395 -845
rect 2441 -891 2519 -845
rect 2565 -891 2643 -845
rect 2689 -891 2767 -845
rect 2813 -891 2891 -845
rect 2937 -891 3015 -845
rect 3061 -891 3139 -845
rect 3185 -891 3263 -845
rect 3309 -891 3387 -845
rect 3433 -891 3511 -845
rect 3557 -891 3635 -845
rect 3681 -891 3759 -845
rect 3805 -891 3883 -845
rect 3929 -891 4007 -845
rect 4053 -891 4131 -845
rect 4177 -891 4255 -845
rect 4301 -891 4379 -845
rect 4425 -891 4503 -845
rect 4549 -891 4627 -845
rect 4673 -891 4751 -845
rect 4797 -891 4875 -845
rect 4921 -891 4999 -845
rect 5045 -891 5123 -845
rect 5169 -891 5247 -845
rect 5293 -891 5371 -845
rect 5417 -891 5495 -845
rect 5541 -891 5619 -845
rect 5665 -891 5743 -845
rect 5789 -891 5811 -845
rect -5811 -969 5811 -891
rect -5811 -1015 -5789 -969
rect -5743 -1015 -5665 -969
rect -5619 -1015 -5541 -969
rect -5495 -1015 -5417 -969
rect -5371 -1015 -5293 -969
rect -5247 -1015 -5169 -969
rect -5123 -1015 -5045 -969
rect -4999 -1015 -4921 -969
rect -4875 -1015 -4797 -969
rect -4751 -1015 -4673 -969
rect -4627 -1015 -4549 -969
rect -4503 -1015 -4425 -969
rect -4379 -1015 -4301 -969
rect -4255 -1015 -4177 -969
rect -4131 -1015 -4053 -969
rect -4007 -1015 -3929 -969
rect -3883 -1015 -3805 -969
rect -3759 -1015 -3681 -969
rect -3635 -1015 -3557 -969
rect -3511 -1015 -3433 -969
rect -3387 -1015 -3309 -969
rect -3263 -1015 -3185 -969
rect -3139 -1015 -3061 -969
rect -3015 -1015 -2937 -969
rect -2891 -1015 -2813 -969
rect -2767 -1015 -2689 -969
rect -2643 -1015 -2565 -969
rect -2519 -1015 -2441 -969
rect -2395 -1015 -2317 -969
rect -2271 -1015 -2193 -969
rect -2147 -1015 -2069 -969
rect -2023 -1015 -1945 -969
rect -1899 -1015 -1821 -969
rect -1775 -1015 -1697 -969
rect -1651 -1015 -1573 -969
rect -1527 -1015 -1449 -969
rect -1403 -1015 -1325 -969
rect -1279 -1015 -1201 -969
rect -1155 -1015 -1077 -969
rect -1031 -1015 -953 -969
rect -907 -1015 -829 -969
rect -783 -1015 -705 -969
rect -659 -1015 -581 -969
rect -535 -1015 -457 -969
rect -411 -1015 -333 -969
rect -287 -1015 -209 -969
rect -163 -1015 -85 -969
rect -39 -1015 39 -969
rect 85 -1015 163 -969
rect 209 -1015 287 -969
rect 333 -1015 411 -969
rect 457 -1015 535 -969
rect 581 -1015 659 -969
rect 705 -1015 783 -969
rect 829 -1015 907 -969
rect 953 -1015 1031 -969
rect 1077 -1015 1155 -969
rect 1201 -1015 1279 -969
rect 1325 -1015 1403 -969
rect 1449 -1015 1527 -969
rect 1573 -1015 1651 -969
rect 1697 -1015 1775 -969
rect 1821 -1015 1899 -969
rect 1945 -1015 2023 -969
rect 2069 -1015 2147 -969
rect 2193 -1015 2271 -969
rect 2317 -1015 2395 -969
rect 2441 -1015 2519 -969
rect 2565 -1015 2643 -969
rect 2689 -1015 2767 -969
rect 2813 -1015 2891 -969
rect 2937 -1015 3015 -969
rect 3061 -1015 3139 -969
rect 3185 -1015 3263 -969
rect 3309 -1015 3387 -969
rect 3433 -1015 3511 -969
rect 3557 -1015 3635 -969
rect 3681 -1015 3759 -969
rect 3805 -1015 3883 -969
rect 3929 -1015 4007 -969
rect 4053 -1015 4131 -969
rect 4177 -1015 4255 -969
rect 4301 -1015 4379 -969
rect 4425 -1015 4503 -969
rect 4549 -1015 4627 -969
rect 4673 -1015 4751 -969
rect 4797 -1015 4875 -969
rect 4921 -1015 4999 -969
rect 5045 -1015 5123 -969
rect 5169 -1015 5247 -969
rect 5293 -1015 5371 -969
rect 5417 -1015 5495 -969
rect 5541 -1015 5619 -969
rect 5665 -1015 5743 -969
rect 5789 -1015 5811 -969
rect -5811 -1093 5811 -1015
rect -5811 -1139 -5789 -1093
rect -5743 -1139 -5665 -1093
rect -5619 -1139 -5541 -1093
rect -5495 -1139 -5417 -1093
rect -5371 -1139 -5293 -1093
rect -5247 -1139 -5169 -1093
rect -5123 -1139 -5045 -1093
rect -4999 -1139 -4921 -1093
rect -4875 -1139 -4797 -1093
rect -4751 -1139 -4673 -1093
rect -4627 -1139 -4549 -1093
rect -4503 -1139 -4425 -1093
rect -4379 -1139 -4301 -1093
rect -4255 -1139 -4177 -1093
rect -4131 -1139 -4053 -1093
rect -4007 -1139 -3929 -1093
rect -3883 -1139 -3805 -1093
rect -3759 -1139 -3681 -1093
rect -3635 -1139 -3557 -1093
rect -3511 -1139 -3433 -1093
rect -3387 -1139 -3309 -1093
rect -3263 -1139 -3185 -1093
rect -3139 -1139 -3061 -1093
rect -3015 -1139 -2937 -1093
rect -2891 -1139 -2813 -1093
rect -2767 -1139 -2689 -1093
rect -2643 -1139 -2565 -1093
rect -2519 -1139 -2441 -1093
rect -2395 -1139 -2317 -1093
rect -2271 -1139 -2193 -1093
rect -2147 -1139 -2069 -1093
rect -2023 -1139 -1945 -1093
rect -1899 -1139 -1821 -1093
rect -1775 -1139 -1697 -1093
rect -1651 -1139 -1573 -1093
rect -1527 -1139 -1449 -1093
rect -1403 -1139 -1325 -1093
rect -1279 -1139 -1201 -1093
rect -1155 -1139 -1077 -1093
rect -1031 -1139 -953 -1093
rect -907 -1139 -829 -1093
rect -783 -1139 -705 -1093
rect -659 -1139 -581 -1093
rect -535 -1139 -457 -1093
rect -411 -1139 -333 -1093
rect -287 -1139 -209 -1093
rect -163 -1139 -85 -1093
rect -39 -1139 39 -1093
rect 85 -1139 163 -1093
rect 209 -1139 287 -1093
rect 333 -1139 411 -1093
rect 457 -1139 535 -1093
rect 581 -1139 659 -1093
rect 705 -1139 783 -1093
rect 829 -1139 907 -1093
rect 953 -1139 1031 -1093
rect 1077 -1139 1155 -1093
rect 1201 -1139 1279 -1093
rect 1325 -1139 1403 -1093
rect 1449 -1139 1527 -1093
rect 1573 -1139 1651 -1093
rect 1697 -1139 1775 -1093
rect 1821 -1139 1899 -1093
rect 1945 -1139 2023 -1093
rect 2069 -1139 2147 -1093
rect 2193 -1139 2271 -1093
rect 2317 -1139 2395 -1093
rect 2441 -1139 2519 -1093
rect 2565 -1139 2643 -1093
rect 2689 -1139 2767 -1093
rect 2813 -1139 2891 -1093
rect 2937 -1139 3015 -1093
rect 3061 -1139 3139 -1093
rect 3185 -1139 3263 -1093
rect 3309 -1139 3387 -1093
rect 3433 -1139 3511 -1093
rect 3557 -1139 3635 -1093
rect 3681 -1139 3759 -1093
rect 3805 -1139 3883 -1093
rect 3929 -1139 4007 -1093
rect 4053 -1139 4131 -1093
rect 4177 -1139 4255 -1093
rect 4301 -1139 4379 -1093
rect 4425 -1139 4503 -1093
rect 4549 -1139 4627 -1093
rect 4673 -1139 4751 -1093
rect 4797 -1139 4875 -1093
rect 4921 -1139 4999 -1093
rect 5045 -1139 5123 -1093
rect 5169 -1139 5247 -1093
rect 5293 -1139 5371 -1093
rect 5417 -1139 5495 -1093
rect 5541 -1139 5619 -1093
rect 5665 -1139 5743 -1093
rect 5789 -1139 5811 -1093
rect -5811 -1217 5811 -1139
rect -5811 -1263 -5789 -1217
rect -5743 -1263 -5665 -1217
rect -5619 -1263 -5541 -1217
rect -5495 -1263 -5417 -1217
rect -5371 -1263 -5293 -1217
rect -5247 -1263 -5169 -1217
rect -5123 -1263 -5045 -1217
rect -4999 -1263 -4921 -1217
rect -4875 -1263 -4797 -1217
rect -4751 -1263 -4673 -1217
rect -4627 -1263 -4549 -1217
rect -4503 -1263 -4425 -1217
rect -4379 -1263 -4301 -1217
rect -4255 -1263 -4177 -1217
rect -4131 -1263 -4053 -1217
rect -4007 -1263 -3929 -1217
rect -3883 -1263 -3805 -1217
rect -3759 -1263 -3681 -1217
rect -3635 -1263 -3557 -1217
rect -3511 -1263 -3433 -1217
rect -3387 -1263 -3309 -1217
rect -3263 -1263 -3185 -1217
rect -3139 -1263 -3061 -1217
rect -3015 -1263 -2937 -1217
rect -2891 -1263 -2813 -1217
rect -2767 -1263 -2689 -1217
rect -2643 -1263 -2565 -1217
rect -2519 -1263 -2441 -1217
rect -2395 -1263 -2317 -1217
rect -2271 -1263 -2193 -1217
rect -2147 -1263 -2069 -1217
rect -2023 -1263 -1945 -1217
rect -1899 -1263 -1821 -1217
rect -1775 -1263 -1697 -1217
rect -1651 -1263 -1573 -1217
rect -1527 -1263 -1449 -1217
rect -1403 -1263 -1325 -1217
rect -1279 -1263 -1201 -1217
rect -1155 -1263 -1077 -1217
rect -1031 -1263 -953 -1217
rect -907 -1263 -829 -1217
rect -783 -1263 -705 -1217
rect -659 -1263 -581 -1217
rect -535 -1263 -457 -1217
rect -411 -1263 -333 -1217
rect -287 -1263 -209 -1217
rect -163 -1263 -85 -1217
rect -39 -1263 39 -1217
rect 85 -1263 163 -1217
rect 209 -1263 287 -1217
rect 333 -1263 411 -1217
rect 457 -1263 535 -1217
rect 581 -1263 659 -1217
rect 705 -1263 783 -1217
rect 829 -1263 907 -1217
rect 953 -1263 1031 -1217
rect 1077 -1263 1155 -1217
rect 1201 -1263 1279 -1217
rect 1325 -1263 1403 -1217
rect 1449 -1263 1527 -1217
rect 1573 -1263 1651 -1217
rect 1697 -1263 1775 -1217
rect 1821 -1263 1899 -1217
rect 1945 -1263 2023 -1217
rect 2069 -1263 2147 -1217
rect 2193 -1263 2271 -1217
rect 2317 -1263 2395 -1217
rect 2441 -1263 2519 -1217
rect 2565 -1263 2643 -1217
rect 2689 -1263 2767 -1217
rect 2813 -1263 2891 -1217
rect 2937 -1263 3015 -1217
rect 3061 -1263 3139 -1217
rect 3185 -1263 3263 -1217
rect 3309 -1263 3387 -1217
rect 3433 -1263 3511 -1217
rect 3557 -1263 3635 -1217
rect 3681 -1263 3759 -1217
rect 3805 -1263 3883 -1217
rect 3929 -1263 4007 -1217
rect 4053 -1263 4131 -1217
rect 4177 -1263 4255 -1217
rect 4301 -1263 4379 -1217
rect 4425 -1263 4503 -1217
rect 4549 -1263 4627 -1217
rect 4673 -1263 4751 -1217
rect 4797 -1263 4875 -1217
rect 4921 -1263 4999 -1217
rect 5045 -1263 5123 -1217
rect 5169 -1263 5247 -1217
rect 5293 -1263 5371 -1217
rect 5417 -1263 5495 -1217
rect 5541 -1263 5619 -1217
rect 5665 -1263 5743 -1217
rect 5789 -1263 5811 -1217
rect -5811 -1285 5811 -1263
<< psubdiffcont >>
rect -5789 1217 -5743 1263
rect -5665 1217 -5619 1263
rect -5541 1217 -5495 1263
rect -5417 1217 -5371 1263
rect -5293 1217 -5247 1263
rect -5169 1217 -5123 1263
rect -5045 1217 -4999 1263
rect -4921 1217 -4875 1263
rect -4797 1217 -4751 1263
rect -4673 1217 -4627 1263
rect -4549 1217 -4503 1263
rect -4425 1217 -4379 1263
rect -4301 1217 -4255 1263
rect -4177 1217 -4131 1263
rect -4053 1217 -4007 1263
rect -3929 1217 -3883 1263
rect -3805 1217 -3759 1263
rect -3681 1217 -3635 1263
rect -3557 1217 -3511 1263
rect -3433 1217 -3387 1263
rect -3309 1217 -3263 1263
rect -3185 1217 -3139 1263
rect -3061 1217 -3015 1263
rect -2937 1217 -2891 1263
rect -2813 1217 -2767 1263
rect -2689 1217 -2643 1263
rect -2565 1217 -2519 1263
rect -2441 1217 -2395 1263
rect -2317 1217 -2271 1263
rect -2193 1217 -2147 1263
rect -2069 1217 -2023 1263
rect -1945 1217 -1899 1263
rect -1821 1217 -1775 1263
rect -1697 1217 -1651 1263
rect -1573 1217 -1527 1263
rect -1449 1217 -1403 1263
rect -1325 1217 -1279 1263
rect -1201 1217 -1155 1263
rect -1077 1217 -1031 1263
rect -953 1217 -907 1263
rect -829 1217 -783 1263
rect -705 1217 -659 1263
rect -581 1217 -535 1263
rect -457 1217 -411 1263
rect -333 1217 -287 1263
rect -209 1217 -163 1263
rect -85 1217 -39 1263
rect 39 1217 85 1263
rect 163 1217 209 1263
rect 287 1217 333 1263
rect 411 1217 457 1263
rect 535 1217 581 1263
rect 659 1217 705 1263
rect 783 1217 829 1263
rect 907 1217 953 1263
rect 1031 1217 1077 1263
rect 1155 1217 1201 1263
rect 1279 1217 1325 1263
rect 1403 1217 1449 1263
rect 1527 1217 1573 1263
rect 1651 1217 1697 1263
rect 1775 1217 1821 1263
rect 1899 1217 1945 1263
rect 2023 1217 2069 1263
rect 2147 1217 2193 1263
rect 2271 1217 2317 1263
rect 2395 1217 2441 1263
rect 2519 1217 2565 1263
rect 2643 1217 2689 1263
rect 2767 1217 2813 1263
rect 2891 1217 2937 1263
rect 3015 1217 3061 1263
rect 3139 1217 3185 1263
rect 3263 1217 3309 1263
rect 3387 1217 3433 1263
rect 3511 1217 3557 1263
rect 3635 1217 3681 1263
rect 3759 1217 3805 1263
rect 3883 1217 3929 1263
rect 4007 1217 4053 1263
rect 4131 1217 4177 1263
rect 4255 1217 4301 1263
rect 4379 1217 4425 1263
rect 4503 1217 4549 1263
rect 4627 1217 4673 1263
rect 4751 1217 4797 1263
rect 4875 1217 4921 1263
rect 4999 1217 5045 1263
rect 5123 1217 5169 1263
rect 5247 1217 5293 1263
rect 5371 1217 5417 1263
rect 5495 1217 5541 1263
rect 5619 1217 5665 1263
rect 5743 1217 5789 1263
rect -5789 1093 -5743 1139
rect -5665 1093 -5619 1139
rect -5541 1093 -5495 1139
rect -5417 1093 -5371 1139
rect -5293 1093 -5247 1139
rect -5169 1093 -5123 1139
rect -5045 1093 -4999 1139
rect -4921 1093 -4875 1139
rect -4797 1093 -4751 1139
rect -4673 1093 -4627 1139
rect -4549 1093 -4503 1139
rect -4425 1093 -4379 1139
rect -4301 1093 -4255 1139
rect -4177 1093 -4131 1139
rect -4053 1093 -4007 1139
rect -3929 1093 -3883 1139
rect -3805 1093 -3759 1139
rect -3681 1093 -3635 1139
rect -3557 1093 -3511 1139
rect -3433 1093 -3387 1139
rect -3309 1093 -3263 1139
rect -3185 1093 -3139 1139
rect -3061 1093 -3015 1139
rect -2937 1093 -2891 1139
rect -2813 1093 -2767 1139
rect -2689 1093 -2643 1139
rect -2565 1093 -2519 1139
rect -2441 1093 -2395 1139
rect -2317 1093 -2271 1139
rect -2193 1093 -2147 1139
rect -2069 1093 -2023 1139
rect -1945 1093 -1899 1139
rect -1821 1093 -1775 1139
rect -1697 1093 -1651 1139
rect -1573 1093 -1527 1139
rect -1449 1093 -1403 1139
rect -1325 1093 -1279 1139
rect -1201 1093 -1155 1139
rect -1077 1093 -1031 1139
rect -953 1093 -907 1139
rect -829 1093 -783 1139
rect -705 1093 -659 1139
rect -581 1093 -535 1139
rect -457 1093 -411 1139
rect -333 1093 -287 1139
rect -209 1093 -163 1139
rect -85 1093 -39 1139
rect 39 1093 85 1139
rect 163 1093 209 1139
rect 287 1093 333 1139
rect 411 1093 457 1139
rect 535 1093 581 1139
rect 659 1093 705 1139
rect 783 1093 829 1139
rect 907 1093 953 1139
rect 1031 1093 1077 1139
rect 1155 1093 1201 1139
rect 1279 1093 1325 1139
rect 1403 1093 1449 1139
rect 1527 1093 1573 1139
rect 1651 1093 1697 1139
rect 1775 1093 1821 1139
rect 1899 1093 1945 1139
rect 2023 1093 2069 1139
rect 2147 1093 2193 1139
rect 2271 1093 2317 1139
rect 2395 1093 2441 1139
rect 2519 1093 2565 1139
rect 2643 1093 2689 1139
rect 2767 1093 2813 1139
rect 2891 1093 2937 1139
rect 3015 1093 3061 1139
rect 3139 1093 3185 1139
rect 3263 1093 3309 1139
rect 3387 1093 3433 1139
rect 3511 1093 3557 1139
rect 3635 1093 3681 1139
rect 3759 1093 3805 1139
rect 3883 1093 3929 1139
rect 4007 1093 4053 1139
rect 4131 1093 4177 1139
rect 4255 1093 4301 1139
rect 4379 1093 4425 1139
rect 4503 1093 4549 1139
rect 4627 1093 4673 1139
rect 4751 1093 4797 1139
rect 4875 1093 4921 1139
rect 4999 1093 5045 1139
rect 5123 1093 5169 1139
rect 5247 1093 5293 1139
rect 5371 1093 5417 1139
rect 5495 1093 5541 1139
rect 5619 1093 5665 1139
rect 5743 1093 5789 1139
rect -5789 969 -5743 1015
rect -5665 969 -5619 1015
rect -5541 969 -5495 1015
rect -5417 969 -5371 1015
rect -5293 969 -5247 1015
rect -5169 969 -5123 1015
rect -5045 969 -4999 1015
rect -4921 969 -4875 1015
rect -4797 969 -4751 1015
rect -4673 969 -4627 1015
rect -4549 969 -4503 1015
rect -4425 969 -4379 1015
rect -4301 969 -4255 1015
rect -4177 969 -4131 1015
rect -4053 969 -4007 1015
rect -3929 969 -3883 1015
rect -3805 969 -3759 1015
rect -3681 969 -3635 1015
rect -3557 969 -3511 1015
rect -3433 969 -3387 1015
rect -3309 969 -3263 1015
rect -3185 969 -3139 1015
rect -3061 969 -3015 1015
rect -2937 969 -2891 1015
rect -2813 969 -2767 1015
rect -2689 969 -2643 1015
rect -2565 969 -2519 1015
rect -2441 969 -2395 1015
rect -2317 969 -2271 1015
rect -2193 969 -2147 1015
rect -2069 969 -2023 1015
rect -1945 969 -1899 1015
rect -1821 969 -1775 1015
rect -1697 969 -1651 1015
rect -1573 969 -1527 1015
rect -1449 969 -1403 1015
rect -1325 969 -1279 1015
rect -1201 969 -1155 1015
rect -1077 969 -1031 1015
rect -953 969 -907 1015
rect -829 969 -783 1015
rect -705 969 -659 1015
rect -581 969 -535 1015
rect -457 969 -411 1015
rect -333 969 -287 1015
rect -209 969 -163 1015
rect -85 969 -39 1015
rect 39 969 85 1015
rect 163 969 209 1015
rect 287 969 333 1015
rect 411 969 457 1015
rect 535 969 581 1015
rect 659 969 705 1015
rect 783 969 829 1015
rect 907 969 953 1015
rect 1031 969 1077 1015
rect 1155 969 1201 1015
rect 1279 969 1325 1015
rect 1403 969 1449 1015
rect 1527 969 1573 1015
rect 1651 969 1697 1015
rect 1775 969 1821 1015
rect 1899 969 1945 1015
rect 2023 969 2069 1015
rect 2147 969 2193 1015
rect 2271 969 2317 1015
rect 2395 969 2441 1015
rect 2519 969 2565 1015
rect 2643 969 2689 1015
rect 2767 969 2813 1015
rect 2891 969 2937 1015
rect 3015 969 3061 1015
rect 3139 969 3185 1015
rect 3263 969 3309 1015
rect 3387 969 3433 1015
rect 3511 969 3557 1015
rect 3635 969 3681 1015
rect 3759 969 3805 1015
rect 3883 969 3929 1015
rect 4007 969 4053 1015
rect 4131 969 4177 1015
rect 4255 969 4301 1015
rect 4379 969 4425 1015
rect 4503 969 4549 1015
rect 4627 969 4673 1015
rect 4751 969 4797 1015
rect 4875 969 4921 1015
rect 4999 969 5045 1015
rect 5123 969 5169 1015
rect 5247 969 5293 1015
rect 5371 969 5417 1015
rect 5495 969 5541 1015
rect 5619 969 5665 1015
rect 5743 969 5789 1015
rect -5789 845 -5743 891
rect -5665 845 -5619 891
rect -5541 845 -5495 891
rect -5417 845 -5371 891
rect -5293 845 -5247 891
rect -5169 845 -5123 891
rect -5045 845 -4999 891
rect -4921 845 -4875 891
rect -4797 845 -4751 891
rect -4673 845 -4627 891
rect -4549 845 -4503 891
rect -4425 845 -4379 891
rect -4301 845 -4255 891
rect -4177 845 -4131 891
rect -4053 845 -4007 891
rect -3929 845 -3883 891
rect -3805 845 -3759 891
rect -3681 845 -3635 891
rect -3557 845 -3511 891
rect -3433 845 -3387 891
rect -3309 845 -3263 891
rect -3185 845 -3139 891
rect -3061 845 -3015 891
rect -2937 845 -2891 891
rect -2813 845 -2767 891
rect -2689 845 -2643 891
rect -2565 845 -2519 891
rect -2441 845 -2395 891
rect -2317 845 -2271 891
rect -2193 845 -2147 891
rect -2069 845 -2023 891
rect -1945 845 -1899 891
rect -1821 845 -1775 891
rect -1697 845 -1651 891
rect -1573 845 -1527 891
rect -1449 845 -1403 891
rect -1325 845 -1279 891
rect -1201 845 -1155 891
rect -1077 845 -1031 891
rect -953 845 -907 891
rect -829 845 -783 891
rect -705 845 -659 891
rect -581 845 -535 891
rect -457 845 -411 891
rect -333 845 -287 891
rect -209 845 -163 891
rect -85 845 -39 891
rect 39 845 85 891
rect 163 845 209 891
rect 287 845 333 891
rect 411 845 457 891
rect 535 845 581 891
rect 659 845 705 891
rect 783 845 829 891
rect 907 845 953 891
rect 1031 845 1077 891
rect 1155 845 1201 891
rect 1279 845 1325 891
rect 1403 845 1449 891
rect 1527 845 1573 891
rect 1651 845 1697 891
rect 1775 845 1821 891
rect 1899 845 1945 891
rect 2023 845 2069 891
rect 2147 845 2193 891
rect 2271 845 2317 891
rect 2395 845 2441 891
rect 2519 845 2565 891
rect 2643 845 2689 891
rect 2767 845 2813 891
rect 2891 845 2937 891
rect 3015 845 3061 891
rect 3139 845 3185 891
rect 3263 845 3309 891
rect 3387 845 3433 891
rect 3511 845 3557 891
rect 3635 845 3681 891
rect 3759 845 3805 891
rect 3883 845 3929 891
rect 4007 845 4053 891
rect 4131 845 4177 891
rect 4255 845 4301 891
rect 4379 845 4425 891
rect 4503 845 4549 891
rect 4627 845 4673 891
rect 4751 845 4797 891
rect 4875 845 4921 891
rect 4999 845 5045 891
rect 5123 845 5169 891
rect 5247 845 5293 891
rect 5371 845 5417 891
rect 5495 845 5541 891
rect 5619 845 5665 891
rect 5743 845 5789 891
rect -5789 721 -5743 767
rect -5665 721 -5619 767
rect -5541 721 -5495 767
rect -5417 721 -5371 767
rect -5293 721 -5247 767
rect -5169 721 -5123 767
rect -5045 721 -4999 767
rect -4921 721 -4875 767
rect -4797 721 -4751 767
rect -4673 721 -4627 767
rect -4549 721 -4503 767
rect -4425 721 -4379 767
rect -4301 721 -4255 767
rect -4177 721 -4131 767
rect -4053 721 -4007 767
rect -3929 721 -3883 767
rect -3805 721 -3759 767
rect -3681 721 -3635 767
rect -3557 721 -3511 767
rect -3433 721 -3387 767
rect -3309 721 -3263 767
rect -3185 721 -3139 767
rect -3061 721 -3015 767
rect -2937 721 -2891 767
rect -2813 721 -2767 767
rect -2689 721 -2643 767
rect -2565 721 -2519 767
rect -2441 721 -2395 767
rect -2317 721 -2271 767
rect -2193 721 -2147 767
rect -2069 721 -2023 767
rect -1945 721 -1899 767
rect -1821 721 -1775 767
rect -1697 721 -1651 767
rect -1573 721 -1527 767
rect -1449 721 -1403 767
rect -1325 721 -1279 767
rect -1201 721 -1155 767
rect -1077 721 -1031 767
rect -953 721 -907 767
rect -829 721 -783 767
rect -705 721 -659 767
rect -581 721 -535 767
rect -457 721 -411 767
rect -333 721 -287 767
rect -209 721 -163 767
rect -85 721 -39 767
rect 39 721 85 767
rect 163 721 209 767
rect 287 721 333 767
rect 411 721 457 767
rect 535 721 581 767
rect 659 721 705 767
rect 783 721 829 767
rect 907 721 953 767
rect 1031 721 1077 767
rect 1155 721 1201 767
rect 1279 721 1325 767
rect 1403 721 1449 767
rect 1527 721 1573 767
rect 1651 721 1697 767
rect 1775 721 1821 767
rect 1899 721 1945 767
rect 2023 721 2069 767
rect 2147 721 2193 767
rect 2271 721 2317 767
rect 2395 721 2441 767
rect 2519 721 2565 767
rect 2643 721 2689 767
rect 2767 721 2813 767
rect 2891 721 2937 767
rect 3015 721 3061 767
rect 3139 721 3185 767
rect 3263 721 3309 767
rect 3387 721 3433 767
rect 3511 721 3557 767
rect 3635 721 3681 767
rect 3759 721 3805 767
rect 3883 721 3929 767
rect 4007 721 4053 767
rect 4131 721 4177 767
rect 4255 721 4301 767
rect 4379 721 4425 767
rect 4503 721 4549 767
rect 4627 721 4673 767
rect 4751 721 4797 767
rect 4875 721 4921 767
rect 4999 721 5045 767
rect 5123 721 5169 767
rect 5247 721 5293 767
rect 5371 721 5417 767
rect 5495 721 5541 767
rect 5619 721 5665 767
rect 5743 721 5789 767
rect -5789 597 -5743 643
rect -5665 597 -5619 643
rect -5541 597 -5495 643
rect -5417 597 -5371 643
rect -5293 597 -5247 643
rect -5169 597 -5123 643
rect -5045 597 -4999 643
rect -4921 597 -4875 643
rect -4797 597 -4751 643
rect -4673 597 -4627 643
rect -4549 597 -4503 643
rect -4425 597 -4379 643
rect -4301 597 -4255 643
rect -4177 597 -4131 643
rect -4053 597 -4007 643
rect -3929 597 -3883 643
rect -3805 597 -3759 643
rect -3681 597 -3635 643
rect -3557 597 -3511 643
rect -3433 597 -3387 643
rect -3309 597 -3263 643
rect -3185 597 -3139 643
rect -3061 597 -3015 643
rect -2937 597 -2891 643
rect -2813 597 -2767 643
rect -2689 597 -2643 643
rect -2565 597 -2519 643
rect -2441 597 -2395 643
rect -2317 597 -2271 643
rect -2193 597 -2147 643
rect -2069 597 -2023 643
rect -1945 597 -1899 643
rect -1821 597 -1775 643
rect -1697 597 -1651 643
rect -1573 597 -1527 643
rect -1449 597 -1403 643
rect -1325 597 -1279 643
rect -1201 597 -1155 643
rect -1077 597 -1031 643
rect -953 597 -907 643
rect -829 597 -783 643
rect -705 597 -659 643
rect -581 597 -535 643
rect -457 597 -411 643
rect -333 597 -287 643
rect -209 597 -163 643
rect -85 597 -39 643
rect 39 597 85 643
rect 163 597 209 643
rect 287 597 333 643
rect 411 597 457 643
rect 535 597 581 643
rect 659 597 705 643
rect 783 597 829 643
rect 907 597 953 643
rect 1031 597 1077 643
rect 1155 597 1201 643
rect 1279 597 1325 643
rect 1403 597 1449 643
rect 1527 597 1573 643
rect 1651 597 1697 643
rect 1775 597 1821 643
rect 1899 597 1945 643
rect 2023 597 2069 643
rect 2147 597 2193 643
rect 2271 597 2317 643
rect 2395 597 2441 643
rect 2519 597 2565 643
rect 2643 597 2689 643
rect 2767 597 2813 643
rect 2891 597 2937 643
rect 3015 597 3061 643
rect 3139 597 3185 643
rect 3263 597 3309 643
rect 3387 597 3433 643
rect 3511 597 3557 643
rect 3635 597 3681 643
rect 3759 597 3805 643
rect 3883 597 3929 643
rect 4007 597 4053 643
rect 4131 597 4177 643
rect 4255 597 4301 643
rect 4379 597 4425 643
rect 4503 597 4549 643
rect 4627 597 4673 643
rect 4751 597 4797 643
rect 4875 597 4921 643
rect 4999 597 5045 643
rect 5123 597 5169 643
rect 5247 597 5293 643
rect 5371 597 5417 643
rect 5495 597 5541 643
rect 5619 597 5665 643
rect 5743 597 5789 643
rect -5789 473 -5743 519
rect -5665 473 -5619 519
rect -5541 473 -5495 519
rect -5417 473 -5371 519
rect -5293 473 -5247 519
rect -5169 473 -5123 519
rect -5045 473 -4999 519
rect -4921 473 -4875 519
rect -4797 473 -4751 519
rect -4673 473 -4627 519
rect -4549 473 -4503 519
rect -4425 473 -4379 519
rect -4301 473 -4255 519
rect -4177 473 -4131 519
rect -4053 473 -4007 519
rect -3929 473 -3883 519
rect -3805 473 -3759 519
rect -3681 473 -3635 519
rect -3557 473 -3511 519
rect -3433 473 -3387 519
rect -3309 473 -3263 519
rect -3185 473 -3139 519
rect -3061 473 -3015 519
rect -2937 473 -2891 519
rect -2813 473 -2767 519
rect -2689 473 -2643 519
rect -2565 473 -2519 519
rect -2441 473 -2395 519
rect -2317 473 -2271 519
rect -2193 473 -2147 519
rect -2069 473 -2023 519
rect -1945 473 -1899 519
rect -1821 473 -1775 519
rect -1697 473 -1651 519
rect -1573 473 -1527 519
rect -1449 473 -1403 519
rect -1325 473 -1279 519
rect -1201 473 -1155 519
rect -1077 473 -1031 519
rect -953 473 -907 519
rect -829 473 -783 519
rect -705 473 -659 519
rect -581 473 -535 519
rect -457 473 -411 519
rect -333 473 -287 519
rect -209 473 -163 519
rect -85 473 -39 519
rect 39 473 85 519
rect 163 473 209 519
rect 287 473 333 519
rect 411 473 457 519
rect 535 473 581 519
rect 659 473 705 519
rect 783 473 829 519
rect 907 473 953 519
rect 1031 473 1077 519
rect 1155 473 1201 519
rect 1279 473 1325 519
rect 1403 473 1449 519
rect 1527 473 1573 519
rect 1651 473 1697 519
rect 1775 473 1821 519
rect 1899 473 1945 519
rect 2023 473 2069 519
rect 2147 473 2193 519
rect 2271 473 2317 519
rect 2395 473 2441 519
rect 2519 473 2565 519
rect 2643 473 2689 519
rect 2767 473 2813 519
rect 2891 473 2937 519
rect 3015 473 3061 519
rect 3139 473 3185 519
rect 3263 473 3309 519
rect 3387 473 3433 519
rect 3511 473 3557 519
rect 3635 473 3681 519
rect 3759 473 3805 519
rect 3883 473 3929 519
rect 4007 473 4053 519
rect 4131 473 4177 519
rect 4255 473 4301 519
rect 4379 473 4425 519
rect 4503 473 4549 519
rect 4627 473 4673 519
rect 4751 473 4797 519
rect 4875 473 4921 519
rect 4999 473 5045 519
rect 5123 473 5169 519
rect 5247 473 5293 519
rect 5371 473 5417 519
rect 5495 473 5541 519
rect 5619 473 5665 519
rect 5743 473 5789 519
rect -5789 349 -5743 395
rect -5665 349 -5619 395
rect -5541 349 -5495 395
rect -5417 349 -5371 395
rect -5293 349 -5247 395
rect -5169 349 -5123 395
rect -5045 349 -4999 395
rect -4921 349 -4875 395
rect -4797 349 -4751 395
rect -4673 349 -4627 395
rect -4549 349 -4503 395
rect -4425 349 -4379 395
rect -4301 349 -4255 395
rect -4177 349 -4131 395
rect -4053 349 -4007 395
rect -3929 349 -3883 395
rect -3805 349 -3759 395
rect -3681 349 -3635 395
rect -3557 349 -3511 395
rect -3433 349 -3387 395
rect -3309 349 -3263 395
rect -3185 349 -3139 395
rect -3061 349 -3015 395
rect -2937 349 -2891 395
rect -2813 349 -2767 395
rect -2689 349 -2643 395
rect -2565 349 -2519 395
rect -2441 349 -2395 395
rect -2317 349 -2271 395
rect -2193 349 -2147 395
rect -2069 349 -2023 395
rect -1945 349 -1899 395
rect -1821 349 -1775 395
rect -1697 349 -1651 395
rect -1573 349 -1527 395
rect -1449 349 -1403 395
rect -1325 349 -1279 395
rect -1201 349 -1155 395
rect -1077 349 -1031 395
rect -953 349 -907 395
rect -829 349 -783 395
rect -705 349 -659 395
rect -581 349 -535 395
rect -457 349 -411 395
rect -333 349 -287 395
rect -209 349 -163 395
rect -85 349 -39 395
rect 39 349 85 395
rect 163 349 209 395
rect 287 349 333 395
rect 411 349 457 395
rect 535 349 581 395
rect 659 349 705 395
rect 783 349 829 395
rect 907 349 953 395
rect 1031 349 1077 395
rect 1155 349 1201 395
rect 1279 349 1325 395
rect 1403 349 1449 395
rect 1527 349 1573 395
rect 1651 349 1697 395
rect 1775 349 1821 395
rect 1899 349 1945 395
rect 2023 349 2069 395
rect 2147 349 2193 395
rect 2271 349 2317 395
rect 2395 349 2441 395
rect 2519 349 2565 395
rect 2643 349 2689 395
rect 2767 349 2813 395
rect 2891 349 2937 395
rect 3015 349 3061 395
rect 3139 349 3185 395
rect 3263 349 3309 395
rect 3387 349 3433 395
rect 3511 349 3557 395
rect 3635 349 3681 395
rect 3759 349 3805 395
rect 3883 349 3929 395
rect 4007 349 4053 395
rect 4131 349 4177 395
rect 4255 349 4301 395
rect 4379 349 4425 395
rect 4503 349 4549 395
rect 4627 349 4673 395
rect 4751 349 4797 395
rect 4875 349 4921 395
rect 4999 349 5045 395
rect 5123 349 5169 395
rect 5247 349 5293 395
rect 5371 349 5417 395
rect 5495 349 5541 395
rect 5619 349 5665 395
rect 5743 349 5789 395
rect -5789 225 -5743 271
rect -5665 225 -5619 271
rect -5541 225 -5495 271
rect -5417 225 -5371 271
rect -5293 225 -5247 271
rect -5169 225 -5123 271
rect -5045 225 -4999 271
rect -4921 225 -4875 271
rect -4797 225 -4751 271
rect -4673 225 -4627 271
rect -4549 225 -4503 271
rect -4425 225 -4379 271
rect -4301 225 -4255 271
rect -4177 225 -4131 271
rect -4053 225 -4007 271
rect -3929 225 -3883 271
rect -3805 225 -3759 271
rect -3681 225 -3635 271
rect -3557 225 -3511 271
rect -3433 225 -3387 271
rect -3309 225 -3263 271
rect -3185 225 -3139 271
rect -3061 225 -3015 271
rect -2937 225 -2891 271
rect -2813 225 -2767 271
rect -2689 225 -2643 271
rect -2565 225 -2519 271
rect -2441 225 -2395 271
rect -2317 225 -2271 271
rect -2193 225 -2147 271
rect -2069 225 -2023 271
rect -1945 225 -1899 271
rect -1821 225 -1775 271
rect -1697 225 -1651 271
rect -1573 225 -1527 271
rect -1449 225 -1403 271
rect -1325 225 -1279 271
rect -1201 225 -1155 271
rect -1077 225 -1031 271
rect -953 225 -907 271
rect -829 225 -783 271
rect -705 225 -659 271
rect -581 225 -535 271
rect -457 225 -411 271
rect -333 225 -287 271
rect -209 225 -163 271
rect -85 225 -39 271
rect 39 225 85 271
rect 163 225 209 271
rect 287 225 333 271
rect 411 225 457 271
rect 535 225 581 271
rect 659 225 705 271
rect 783 225 829 271
rect 907 225 953 271
rect 1031 225 1077 271
rect 1155 225 1201 271
rect 1279 225 1325 271
rect 1403 225 1449 271
rect 1527 225 1573 271
rect 1651 225 1697 271
rect 1775 225 1821 271
rect 1899 225 1945 271
rect 2023 225 2069 271
rect 2147 225 2193 271
rect 2271 225 2317 271
rect 2395 225 2441 271
rect 2519 225 2565 271
rect 2643 225 2689 271
rect 2767 225 2813 271
rect 2891 225 2937 271
rect 3015 225 3061 271
rect 3139 225 3185 271
rect 3263 225 3309 271
rect 3387 225 3433 271
rect 3511 225 3557 271
rect 3635 225 3681 271
rect 3759 225 3805 271
rect 3883 225 3929 271
rect 4007 225 4053 271
rect 4131 225 4177 271
rect 4255 225 4301 271
rect 4379 225 4425 271
rect 4503 225 4549 271
rect 4627 225 4673 271
rect 4751 225 4797 271
rect 4875 225 4921 271
rect 4999 225 5045 271
rect 5123 225 5169 271
rect 5247 225 5293 271
rect 5371 225 5417 271
rect 5495 225 5541 271
rect 5619 225 5665 271
rect 5743 225 5789 271
rect -5789 101 -5743 147
rect -5665 101 -5619 147
rect -5541 101 -5495 147
rect -5417 101 -5371 147
rect -5293 101 -5247 147
rect -5169 101 -5123 147
rect -5045 101 -4999 147
rect -4921 101 -4875 147
rect -4797 101 -4751 147
rect -4673 101 -4627 147
rect -4549 101 -4503 147
rect -4425 101 -4379 147
rect -4301 101 -4255 147
rect -4177 101 -4131 147
rect -4053 101 -4007 147
rect -3929 101 -3883 147
rect -3805 101 -3759 147
rect -3681 101 -3635 147
rect -3557 101 -3511 147
rect -3433 101 -3387 147
rect -3309 101 -3263 147
rect -3185 101 -3139 147
rect -3061 101 -3015 147
rect -2937 101 -2891 147
rect -2813 101 -2767 147
rect -2689 101 -2643 147
rect -2565 101 -2519 147
rect -2441 101 -2395 147
rect -2317 101 -2271 147
rect -2193 101 -2147 147
rect -2069 101 -2023 147
rect -1945 101 -1899 147
rect -1821 101 -1775 147
rect -1697 101 -1651 147
rect -1573 101 -1527 147
rect -1449 101 -1403 147
rect -1325 101 -1279 147
rect -1201 101 -1155 147
rect -1077 101 -1031 147
rect -953 101 -907 147
rect -829 101 -783 147
rect -705 101 -659 147
rect -581 101 -535 147
rect -457 101 -411 147
rect -333 101 -287 147
rect -209 101 -163 147
rect -85 101 -39 147
rect 39 101 85 147
rect 163 101 209 147
rect 287 101 333 147
rect 411 101 457 147
rect 535 101 581 147
rect 659 101 705 147
rect 783 101 829 147
rect 907 101 953 147
rect 1031 101 1077 147
rect 1155 101 1201 147
rect 1279 101 1325 147
rect 1403 101 1449 147
rect 1527 101 1573 147
rect 1651 101 1697 147
rect 1775 101 1821 147
rect 1899 101 1945 147
rect 2023 101 2069 147
rect 2147 101 2193 147
rect 2271 101 2317 147
rect 2395 101 2441 147
rect 2519 101 2565 147
rect 2643 101 2689 147
rect 2767 101 2813 147
rect 2891 101 2937 147
rect 3015 101 3061 147
rect 3139 101 3185 147
rect 3263 101 3309 147
rect 3387 101 3433 147
rect 3511 101 3557 147
rect 3635 101 3681 147
rect 3759 101 3805 147
rect 3883 101 3929 147
rect 4007 101 4053 147
rect 4131 101 4177 147
rect 4255 101 4301 147
rect 4379 101 4425 147
rect 4503 101 4549 147
rect 4627 101 4673 147
rect 4751 101 4797 147
rect 4875 101 4921 147
rect 4999 101 5045 147
rect 5123 101 5169 147
rect 5247 101 5293 147
rect 5371 101 5417 147
rect 5495 101 5541 147
rect 5619 101 5665 147
rect 5743 101 5789 147
rect -5789 -23 -5743 23
rect -5665 -23 -5619 23
rect -5541 -23 -5495 23
rect -5417 -23 -5371 23
rect -5293 -23 -5247 23
rect -5169 -23 -5123 23
rect -5045 -23 -4999 23
rect -4921 -23 -4875 23
rect -4797 -23 -4751 23
rect -4673 -23 -4627 23
rect -4549 -23 -4503 23
rect -4425 -23 -4379 23
rect -4301 -23 -4255 23
rect -4177 -23 -4131 23
rect -4053 -23 -4007 23
rect -3929 -23 -3883 23
rect -3805 -23 -3759 23
rect -3681 -23 -3635 23
rect -3557 -23 -3511 23
rect -3433 -23 -3387 23
rect -3309 -23 -3263 23
rect -3185 -23 -3139 23
rect -3061 -23 -3015 23
rect -2937 -23 -2891 23
rect -2813 -23 -2767 23
rect -2689 -23 -2643 23
rect -2565 -23 -2519 23
rect -2441 -23 -2395 23
rect -2317 -23 -2271 23
rect -2193 -23 -2147 23
rect -2069 -23 -2023 23
rect -1945 -23 -1899 23
rect -1821 -23 -1775 23
rect -1697 -23 -1651 23
rect -1573 -23 -1527 23
rect -1449 -23 -1403 23
rect -1325 -23 -1279 23
rect -1201 -23 -1155 23
rect -1077 -23 -1031 23
rect -953 -23 -907 23
rect -829 -23 -783 23
rect -705 -23 -659 23
rect -581 -23 -535 23
rect -457 -23 -411 23
rect -333 -23 -287 23
rect -209 -23 -163 23
rect -85 -23 -39 23
rect 39 -23 85 23
rect 163 -23 209 23
rect 287 -23 333 23
rect 411 -23 457 23
rect 535 -23 581 23
rect 659 -23 705 23
rect 783 -23 829 23
rect 907 -23 953 23
rect 1031 -23 1077 23
rect 1155 -23 1201 23
rect 1279 -23 1325 23
rect 1403 -23 1449 23
rect 1527 -23 1573 23
rect 1651 -23 1697 23
rect 1775 -23 1821 23
rect 1899 -23 1945 23
rect 2023 -23 2069 23
rect 2147 -23 2193 23
rect 2271 -23 2317 23
rect 2395 -23 2441 23
rect 2519 -23 2565 23
rect 2643 -23 2689 23
rect 2767 -23 2813 23
rect 2891 -23 2937 23
rect 3015 -23 3061 23
rect 3139 -23 3185 23
rect 3263 -23 3309 23
rect 3387 -23 3433 23
rect 3511 -23 3557 23
rect 3635 -23 3681 23
rect 3759 -23 3805 23
rect 3883 -23 3929 23
rect 4007 -23 4053 23
rect 4131 -23 4177 23
rect 4255 -23 4301 23
rect 4379 -23 4425 23
rect 4503 -23 4549 23
rect 4627 -23 4673 23
rect 4751 -23 4797 23
rect 4875 -23 4921 23
rect 4999 -23 5045 23
rect 5123 -23 5169 23
rect 5247 -23 5293 23
rect 5371 -23 5417 23
rect 5495 -23 5541 23
rect 5619 -23 5665 23
rect 5743 -23 5789 23
rect -5789 -147 -5743 -101
rect -5665 -147 -5619 -101
rect -5541 -147 -5495 -101
rect -5417 -147 -5371 -101
rect -5293 -147 -5247 -101
rect -5169 -147 -5123 -101
rect -5045 -147 -4999 -101
rect -4921 -147 -4875 -101
rect -4797 -147 -4751 -101
rect -4673 -147 -4627 -101
rect -4549 -147 -4503 -101
rect -4425 -147 -4379 -101
rect -4301 -147 -4255 -101
rect -4177 -147 -4131 -101
rect -4053 -147 -4007 -101
rect -3929 -147 -3883 -101
rect -3805 -147 -3759 -101
rect -3681 -147 -3635 -101
rect -3557 -147 -3511 -101
rect -3433 -147 -3387 -101
rect -3309 -147 -3263 -101
rect -3185 -147 -3139 -101
rect -3061 -147 -3015 -101
rect -2937 -147 -2891 -101
rect -2813 -147 -2767 -101
rect -2689 -147 -2643 -101
rect -2565 -147 -2519 -101
rect -2441 -147 -2395 -101
rect -2317 -147 -2271 -101
rect -2193 -147 -2147 -101
rect -2069 -147 -2023 -101
rect -1945 -147 -1899 -101
rect -1821 -147 -1775 -101
rect -1697 -147 -1651 -101
rect -1573 -147 -1527 -101
rect -1449 -147 -1403 -101
rect -1325 -147 -1279 -101
rect -1201 -147 -1155 -101
rect -1077 -147 -1031 -101
rect -953 -147 -907 -101
rect -829 -147 -783 -101
rect -705 -147 -659 -101
rect -581 -147 -535 -101
rect -457 -147 -411 -101
rect -333 -147 -287 -101
rect -209 -147 -163 -101
rect -85 -147 -39 -101
rect 39 -147 85 -101
rect 163 -147 209 -101
rect 287 -147 333 -101
rect 411 -147 457 -101
rect 535 -147 581 -101
rect 659 -147 705 -101
rect 783 -147 829 -101
rect 907 -147 953 -101
rect 1031 -147 1077 -101
rect 1155 -147 1201 -101
rect 1279 -147 1325 -101
rect 1403 -147 1449 -101
rect 1527 -147 1573 -101
rect 1651 -147 1697 -101
rect 1775 -147 1821 -101
rect 1899 -147 1945 -101
rect 2023 -147 2069 -101
rect 2147 -147 2193 -101
rect 2271 -147 2317 -101
rect 2395 -147 2441 -101
rect 2519 -147 2565 -101
rect 2643 -147 2689 -101
rect 2767 -147 2813 -101
rect 2891 -147 2937 -101
rect 3015 -147 3061 -101
rect 3139 -147 3185 -101
rect 3263 -147 3309 -101
rect 3387 -147 3433 -101
rect 3511 -147 3557 -101
rect 3635 -147 3681 -101
rect 3759 -147 3805 -101
rect 3883 -147 3929 -101
rect 4007 -147 4053 -101
rect 4131 -147 4177 -101
rect 4255 -147 4301 -101
rect 4379 -147 4425 -101
rect 4503 -147 4549 -101
rect 4627 -147 4673 -101
rect 4751 -147 4797 -101
rect 4875 -147 4921 -101
rect 4999 -147 5045 -101
rect 5123 -147 5169 -101
rect 5247 -147 5293 -101
rect 5371 -147 5417 -101
rect 5495 -147 5541 -101
rect 5619 -147 5665 -101
rect 5743 -147 5789 -101
rect -5789 -271 -5743 -225
rect -5665 -271 -5619 -225
rect -5541 -271 -5495 -225
rect -5417 -271 -5371 -225
rect -5293 -271 -5247 -225
rect -5169 -271 -5123 -225
rect -5045 -271 -4999 -225
rect -4921 -271 -4875 -225
rect -4797 -271 -4751 -225
rect -4673 -271 -4627 -225
rect -4549 -271 -4503 -225
rect -4425 -271 -4379 -225
rect -4301 -271 -4255 -225
rect -4177 -271 -4131 -225
rect -4053 -271 -4007 -225
rect -3929 -271 -3883 -225
rect -3805 -271 -3759 -225
rect -3681 -271 -3635 -225
rect -3557 -271 -3511 -225
rect -3433 -271 -3387 -225
rect -3309 -271 -3263 -225
rect -3185 -271 -3139 -225
rect -3061 -271 -3015 -225
rect -2937 -271 -2891 -225
rect -2813 -271 -2767 -225
rect -2689 -271 -2643 -225
rect -2565 -271 -2519 -225
rect -2441 -271 -2395 -225
rect -2317 -271 -2271 -225
rect -2193 -271 -2147 -225
rect -2069 -271 -2023 -225
rect -1945 -271 -1899 -225
rect -1821 -271 -1775 -225
rect -1697 -271 -1651 -225
rect -1573 -271 -1527 -225
rect -1449 -271 -1403 -225
rect -1325 -271 -1279 -225
rect -1201 -271 -1155 -225
rect -1077 -271 -1031 -225
rect -953 -271 -907 -225
rect -829 -271 -783 -225
rect -705 -271 -659 -225
rect -581 -271 -535 -225
rect -457 -271 -411 -225
rect -333 -271 -287 -225
rect -209 -271 -163 -225
rect -85 -271 -39 -225
rect 39 -271 85 -225
rect 163 -271 209 -225
rect 287 -271 333 -225
rect 411 -271 457 -225
rect 535 -271 581 -225
rect 659 -271 705 -225
rect 783 -271 829 -225
rect 907 -271 953 -225
rect 1031 -271 1077 -225
rect 1155 -271 1201 -225
rect 1279 -271 1325 -225
rect 1403 -271 1449 -225
rect 1527 -271 1573 -225
rect 1651 -271 1697 -225
rect 1775 -271 1821 -225
rect 1899 -271 1945 -225
rect 2023 -271 2069 -225
rect 2147 -271 2193 -225
rect 2271 -271 2317 -225
rect 2395 -271 2441 -225
rect 2519 -271 2565 -225
rect 2643 -271 2689 -225
rect 2767 -271 2813 -225
rect 2891 -271 2937 -225
rect 3015 -271 3061 -225
rect 3139 -271 3185 -225
rect 3263 -271 3309 -225
rect 3387 -271 3433 -225
rect 3511 -271 3557 -225
rect 3635 -271 3681 -225
rect 3759 -271 3805 -225
rect 3883 -271 3929 -225
rect 4007 -271 4053 -225
rect 4131 -271 4177 -225
rect 4255 -271 4301 -225
rect 4379 -271 4425 -225
rect 4503 -271 4549 -225
rect 4627 -271 4673 -225
rect 4751 -271 4797 -225
rect 4875 -271 4921 -225
rect 4999 -271 5045 -225
rect 5123 -271 5169 -225
rect 5247 -271 5293 -225
rect 5371 -271 5417 -225
rect 5495 -271 5541 -225
rect 5619 -271 5665 -225
rect 5743 -271 5789 -225
rect -5789 -395 -5743 -349
rect -5665 -395 -5619 -349
rect -5541 -395 -5495 -349
rect -5417 -395 -5371 -349
rect -5293 -395 -5247 -349
rect -5169 -395 -5123 -349
rect -5045 -395 -4999 -349
rect -4921 -395 -4875 -349
rect -4797 -395 -4751 -349
rect -4673 -395 -4627 -349
rect -4549 -395 -4503 -349
rect -4425 -395 -4379 -349
rect -4301 -395 -4255 -349
rect -4177 -395 -4131 -349
rect -4053 -395 -4007 -349
rect -3929 -395 -3883 -349
rect -3805 -395 -3759 -349
rect -3681 -395 -3635 -349
rect -3557 -395 -3511 -349
rect -3433 -395 -3387 -349
rect -3309 -395 -3263 -349
rect -3185 -395 -3139 -349
rect -3061 -395 -3015 -349
rect -2937 -395 -2891 -349
rect -2813 -395 -2767 -349
rect -2689 -395 -2643 -349
rect -2565 -395 -2519 -349
rect -2441 -395 -2395 -349
rect -2317 -395 -2271 -349
rect -2193 -395 -2147 -349
rect -2069 -395 -2023 -349
rect -1945 -395 -1899 -349
rect -1821 -395 -1775 -349
rect -1697 -395 -1651 -349
rect -1573 -395 -1527 -349
rect -1449 -395 -1403 -349
rect -1325 -395 -1279 -349
rect -1201 -395 -1155 -349
rect -1077 -395 -1031 -349
rect -953 -395 -907 -349
rect -829 -395 -783 -349
rect -705 -395 -659 -349
rect -581 -395 -535 -349
rect -457 -395 -411 -349
rect -333 -395 -287 -349
rect -209 -395 -163 -349
rect -85 -395 -39 -349
rect 39 -395 85 -349
rect 163 -395 209 -349
rect 287 -395 333 -349
rect 411 -395 457 -349
rect 535 -395 581 -349
rect 659 -395 705 -349
rect 783 -395 829 -349
rect 907 -395 953 -349
rect 1031 -395 1077 -349
rect 1155 -395 1201 -349
rect 1279 -395 1325 -349
rect 1403 -395 1449 -349
rect 1527 -395 1573 -349
rect 1651 -395 1697 -349
rect 1775 -395 1821 -349
rect 1899 -395 1945 -349
rect 2023 -395 2069 -349
rect 2147 -395 2193 -349
rect 2271 -395 2317 -349
rect 2395 -395 2441 -349
rect 2519 -395 2565 -349
rect 2643 -395 2689 -349
rect 2767 -395 2813 -349
rect 2891 -395 2937 -349
rect 3015 -395 3061 -349
rect 3139 -395 3185 -349
rect 3263 -395 3309 -349
rect 3387 -395 3433 -349
rect 3511 -395 3557 -349
rect 3635 -395 3681 -349
rect 3759 -395 3805 -349
rect 3883 -395 3929 -349
rect 4007 -395 4053 -349
rect 4131 -395 4177 -349
rect 4255 -395 4301 -349
rect 4379 -395 4425 -349
rect 4503 -395 4549 -349
rect 4627 -395 4673 -349
rect 4751 -395 4797 -349
rect 4875 -395 4921 -349
rect 4999 -395 5045 -349
rect 5123 -395 5169 -349
rect 5247 -395 5293 -349
rect 5371 -395 5417 -349
rect 5495 -395 5541 -349
rect 5619 -395 5665 -349
rect 5743 -395 5789 -349
rect -5789 -519 -5743 -473
rect -5665 -519 -5619 -473
rect -5541 -519 -5495 -473
rect -5417 -519 -5371 -473
rect -5293 -519 -5247 -473
rect -5169 -519 -5123 -473
rect -5045 -519 -4999 -473
rect -4921 -519 -4875 -473
rect -4797 -519 -4751 -473
rect -4673 -519 -4627 -473
rect -4549 -519 -4503 -473
rect -4425 -519 -4379 -473
rect -4301 -519 -4255 -473
rect -4177 -519 -4131 -473
rect -4053 -519 -4007 -473
rect -3929 -519 -3883 -473
rect -3805 -519 -3759 -473
rect -3681 -519 -3635 -473
rect -3557 -519 -3511 -473
rect -3433 -519 -3387 -473
rect -3309 -519 -3263 -473
rect -3185 -519 -3139 -473
rect -3061 -519 -3015 -473
rect -2937 -519 -2891 -473
rect -2813 -519 -2767 -473
rect -2689 -519 -2643 -473
rect -2565 -519 -2519 -473
rect -2441 -519 -2395 -473
rect -2317 -519 -2271 -473
rect -2193 -519 -2147 -473
rect -2069 -519 -2023 -473
rect -1945 -519 -1899 -473
rect -1821 -519 -1775 -473
rect -1697 -519 -1651 -473
rect -1573 -519 -1527 -473
rect -1449 -519 -1403 -473
rect -1325 -519 -1279 -473
rect -1201 -519 -1155 -473
rect -1077 -519 -1031 -473
rect -953 -519 -907 -473
rect -829 -519 -783 -473
rect -705 -519 -659 -473
rect -581 -519 -535 -473
rect -457 -519 -411 -473
rect -333 -519 -287 -473
rect -209 -519 -163 -473
rect -85 -519 -39 -473
rect 39 -519 85 -473
rect 163 -519 209 -473
rect 287 -519 333 -473
rect 411 -519 457 -473
rect 535 -519 581 -473
rect 659 -519 705 -473
rect 783 -519 829 -473
rect 907 -519 953 -473
rect 1031 -519 1077 -473
rect 1155 -519 1201 -473
rect 1279 -519 1325 -473
rect 1403 -519 1449 -473
rect 1527 -519 1573 -473
rect 1651 -519 1697 -473
rect 1775 -519 1821 -473
rect 1899 -519 1945 -473
rect 2023 -519 2069 -473
rect 2147 -519 2193 -473
rect 2271 -519 2317 -473
rect 2395 -519 2441 -473
rect 2519 -519 2565 -473
rect 2643 -519 2689 -473
rect 2767 -519 2813 -473
rect 2891 -519 2937 -473
rect 3015 -519 3061 -473
rect 3139 -519 3185 -473
rect 3263 -519 3309 -473
rect 3387 -519 3433 -473
rect 3511 -519 3557 -473
rect 3635 -519 3681 -473
rect 3759 -519 3805 -473
rect 3883 -519 3929 -473
rect 4007 -519 4053 -473
rect 4131 -519 4177 -473
rect 4255 -519 4301 -473
rect 4379 -519 4425 -473
rect 4503 -519 4549 -473
rect 4627 -519 4673 -473
rect 4751 -519 4797 -473
rect 4875 -519 4921 -473
rect 4999 -519 5045 -473
rect 5123 -519 5169 -473
rect 5247 -519 5293 -473
rect 5371 -519 5417 -473
rect 5495 -519 5541 -473
rect 5619 -519 5665 -473
rect 5743 -519 5789 -473
rect -5789 -643 -5743 -597
rect -5665 -643 -5619 -597
rect -5541 -643 -5495 -597
rect -5417 -643 -5371 -597
rect -5293 -643 -5247 -597
rect -5169 -643 -5123 -597
rect -5045 -643 -4999 -597
rect -4921 -643 -4875 -597
rect -4797 -643 -4751 -597
rect -4673 -643 -4627 -597
rect -4549 -643 -4503 -597
rect -4425 -643 -4379 -597
rect -4301 -643 -4255 -597
rect -4177 -643 -4131 -597
rect -4053 -643 -4007 -597
rect -3929 -643 -3883 -597
rect -3805 -643 -3759 -597
rect -3681 -643 -3635 -597
rect -3557 -643 -3511 -597
rect -3433 -643 -3387 -597
rect -3309 -643 -3263 -597
rect -3185 -643 -3139 -597
rect -3061 -643 -3015 -597
rect -2937 -643 -2891 -597
rect -2813 -643 -2767 -597
rect -2689 -643 -2643 -597
rect -2565 -643 -2519 -597
rect -2441 -643 -2395 -597
rect -2317 -643 -2271 -597
rect -2193 -643 -2147 -597
rect -2069 -643 -2023 -597
rect -1945 -643 -1899 -597
rect -1821 -643 -1775 -597
rect -1697 -643 -1651 -597
rect -1573 -643 -1527 -597
rect -1449 -643 -1403 -597
rect -1325 -643 -1279 -597
rect -1201 -643 -1155 -597
rect -1077 -643 -1031 -597
rect -953 -643 -907 -597
rect -829 -643 -783 -597
rect -705 -643 -659 -597
rect -581 -643 -535 -597
rect -457 -643 -411 -597
rect -333 -643 -287 -597
rect -209 -643 -163 -597
rect -85 -643 -39 -597
rect 39 -643 85 -597
rect 163 -643 209 -597
rect 287 -643 333 -597
rect 411 -643 457 -597
rect 535 -643 581 -597
rect 659 -643 705 -597
rect 783 -643 829 -597
rect 907 -643 953 -597
rect 1031 -643 1077 -597
rect 1155 -643 1201 -597
rect 1279 -643 1325 -597
rect 1403 -643 1449 -597
rect 1527 -643 1573 -597
rect 1651 -643 1697 -597
rect 1775 -643 1821 -597
rect 1899 -643 1945 -597
rect 2023 -643 2069 -597
rect 2147 -643 2193 -597
rect 2271 -643 2317 -597
rect 2395 -643 2441 -597
rect 2519 -643 2565 -597
rect 2643 -643 2689 -597
rect 2767 -643 2813 -597
rect 2891 -643 2937 -597
rect 3015 -643 3061 -597
rect 3139 -643 3185 -597
rect 3263 -643 3309 -597
rect 3387 -643 3433 -597
rect 3511 -643 3557 -597
rect 3635 -643 3681 -597
rect 3759 -643 3805 -597
rect 3883 -643 3929 -597
rect 4007 -643 4053 -597
rect 4131 -643 4177 -597
rect 4255 -643 4301 -597
rect 4379 -643 4425 -597
rect 4503 -643 4549 -597
rect 4627 -643 4673 -597
rect 4751 -643 4797 -597
rect 4875 -643 4921 -597
rect 4999 -643 5045 -597
rect 5123 -643 5169 -597
rect 5247 -643 5293 -597
rect 5371 -643 5417 -597
rect 5495 -643 5541 -597
rect 5619 -643 5665 -597
rect 5743 -643 5789 -597
rect -5789 -767 -5743 -721
rect -5665 -767 -5619 -721
rect -5541 -767 -5495 -721
rect -5417 -767 -5371 -721
rect -5293 -767 -5247 -721
rect -5169 -767 -5123 -721
rect -5045 -767 -4999 -721
rect -4921 -767 -4875 -721
rect -4797 -767 -4751 -721
rect -4673 -767 -4627 -721
rect -4549 -767 -4503 -721
rect -4425 -767 -4379 -721
rect -4301 -767 -4255 -721
rect -4177 -767 -4131 -721
rect -4053 -767 -4007 -721
rect -3929 -767 -3883 -721
rect -3805 -767 -3759 -721
rect -3681 -767 -3635 -721
rect -3557 -767 -3511 -721
rect -3433 -767 -3387 -721
rect -3309 -767 -3263 -721
rect -3185 -767 -3139 -721
rect -3061 -767 -3015 -721
rect -2937 -767 -2891 -721
rect -2813 -767 -2767 -721
rect -2689 -767 -2643 -721
rect -2565 -767 -2519 -721
rect -2441 -767 -2395 -721
rect -2317 -767 -2271 -721
rect -2193 -767 -2147 -721
rect -2069 -767 -2023 -721
rect -1945 -767 -1899 -721
rect -1821 -767 -1775 -721
rect -1697 -767 -1651 -721
rect -1573 -767 -1527 -721
rect -1449 -767 -1403 -721
rect -1325 -767 -1279 -721
rect -1201 -767 -1155 -721
rect -1077 -767 -1031 -721
rect -953 -767 -907 -721
rect -829 -767 -783 -721
rect -705 -767 -659 -721
rect -581 -767 -535 -721
rect -457 -767 -411 -721
rect -333 -767 -287 -721
rect -209 -767 -163 -721
rect -85 -767 -39 -721
rect 39 -767 85 -721
rect 163 -767 209 -721
rect 287 -767 333 -721
rect 411 -767 457 -721
rect 535 -767 581 -721
rect 659 -767 705 -721
rect 783 -767 829 -721
rect 907 -767 953 -721
rect 1031 -767 1077 -721
rect 1155 -767 1201 -721
rect 1279 -767 1325 -721
rect 1403 -767 1449 -721
rect 1527 -767 1573 -721
rect 1651 -767 1697 -721
rect 1775 -767 1821 -721
rect 1899 -767 1945 -721
rect 2023 -767 2069 -721
rect 2147 -767 2193 -721
rect 2271 -767 2317 -721
rect 2395 -767 2441 -721
rect 2519 -767 2565 -721
rect 2643 -767 2689 -721
rect 2767 -767 2813 -721
rect 2891 -767 2937 -721
rect 3015 -767 3061 -721
rect 3139 -767 3185 -721
rect 3263 -767 3309 -721
rect 3387 -767 3433 -721
rect 3511 -767 3557 -721
rect 3635 -767 3681 -721
rect 3759 -767 3805 -721
rect 3883 -767 3929 -721
rect 4007 -767 4053 -721
rect 4131 -767 4177 -721
rect 4255 -767 4301 -721
rect 4379 -767 4425 -721
rect 4503 -767 4549 -721
rect 4627 -767 4673 -721
rect 4751 -767 4797 -721
rect 4875 -767 4921 -721
rect 4999 -767 5045 -721
rect 5123 -767 5169 -721
rect 5247 -767 5293 -721
rect 5371 -767 5417 -721
rect 5495 -767 5541 -721
rect 5619 -767 5665 -721
rect 5743 -767 5789 -721
rect -5789 -891 -5743 -845
rect -5665 -891 -5619 -845
rect -5541 -891 -5495 -845
rect -5417 -891 -5371 -845
rect -5293 -891 -5247 -845
rect -5169 -891 -5123 -845
rect -5045 -891 -4999 -845
rect -4921 -891 -4875 -845
rect -4797 -891 -4751 -845
rect -4673 -891 -4627 -845
rect -4549 -891 -4503 -845
rect -4425 -891 -4379 -845
rect -4301 -891 -4255 -845
rect -4177 -891 -4131 -845
rect -4053 -891 -4007 -845
rect -3929 -891 -3883 -845
rect -3805 -891 -3759 -845
rect -3681 -891 -3635 -845
rect -3557 -891 -3511 -845
rect -3433 -891 -3387 -845
rect -3309 -891 -3263 -845
rect -3185 -891 -3139 -845
rect -3061 -891 -3015 -845
rect -2937 -891 -2891 -845
rect -2813 -891 -2767 -845
rect -2689 -891 -2643 -845
rect -2565 -891 -2519 -845
rect -2441 -891 -2395 -845
rect -2317 -891 -2271 -845
rect -2193 -891 -2147 -845
rect -2069 -891 -2023 -845
rect -1945 -891 -1899 -845
rect -1821 -891 -1775 -845
rect -1697 -891 -1651 -845
rect -1573 -891 -1527 -845
rect -1449 -891 -1403 -845
rect -1325 -891 -1279 -845
rect -1201 -891 -1155 -845
rect -1077 -891 -1031 -845
rect -953 -891 -907 -845
rect -829 -891 -783 -845
rect -705 -891 -659 -845
rect -581 -891 -535 -845
rect -457 -891 -411 -845
rect -333 -891 -287 -845
rect -209 -891 -163 -845
rect -85 -891 -39 -845
rect 39 -891 85 -845
rect 163 -891 209 -845
rect 287 -891 333 -845
rect 411 -891 457 -845
rect 535 -891 581 -845
rect 659 -891 705 -845
rect 783 -891 829 -845
rect 907 -891 953 -845
rect 1031 -891 1077 -845
rect 1155 -891 1201 -845
rect 1279 -891 1325 -845
rect 1403 -891 1449 -845
rect 1527 -891 1573 -845
rect 1651 -891 1697 -845
rect 1775 -891 1821 -845
rect 1899 -891 1945 -845
rect 2023 -891 2069 -845
rect 2147 -891 2193 -845
rect 2271 -891 2317 -845
rect 2395 -891 2441 -845
rect 2519 -891 2565 -845
rect 2643 -891 2689 -845
rect 2767 -891 2813 -845
rect 2891 -891 2937 -845
rect 3015 -891 3061 -845
rect 3139 -891 3185 -845
rect 3263 -891 3309 -845
rect 3387 -891 3433 -845
rect 3511 -891 3557 -845
rect 3635 -891 3681 -845
rect 3759 -891 3805 -845
rect 3883 -891 3929 -845
rect 4007 -891 4053 -845
rect 4131 -891 4177 -845
rect 4255 -891 4301 -845
rect 4379 -891 4425 -845
rect 4503 -891 4549 -845
rect 4627 -891 4673 -845
rect 4751 -891 4797 -845
rect 4875 -891 4921 -845
rect 4999 -891 5045 -845
rect 5123 -891 5169 -845
rect 5247 -891 5293 -845
rect 5371 -891 5417 -845
rect 5495 -891 5541 -845
rect 5619 -891 5665 -845
rect 5743 -891 5789 -845
rect -5789 -1015 -5743 -969
rect -5665 -1015 -5619 -969
rect -5541 -1015 -5495 -969
rect -5417 -1015 -5371 -969
rect -5293 -1015 -5247 -969
rect -5169 -1015 -5123 -969
rect -5045 -1015 -4999 -969
rect -4921 -1015 -4875 -969
rect -4797 -1015 -4751 -969
rect -4673 -1015 -4627 -969
rect -4549 -1015 -4503 -969
rect -4425 -1015 -4379 -969
rect -4301 -1015 -4255 -969
rect -4177 -1015 -4131 -969
rect -4053 -1015 -4007 -969
rect -3929 -1015 -3883 -969
rect -3805 -1015 -3759 -969
rect -3681 -1015 -3635 -969
rect -3557 -1015 -3511 -969
rect -3433 -1015 -3387 -969
rect -3309 -1015 -3263 -969
rect -3185 -1015 -3139 -969
rect -3061 -1015 -3015 -969
rect -2937 -1015 -2891 -969
rect -2813 -1015 -2767 -969
rect -2689 -1015 -2643 -969
rect -2565 -1015 -2519 -969
rect -2441 -1015 -2395 -969
rect -2317 -1015 -2271 -969
rect -2193 -1015 -2147 -969
rect -2069 -1015 -2023 -969
rect -1945 -1015 -1899 -969
rect -1821 -1015 -1775 -969
rect -1697 -1015 -1651 -969
rect -1573 -1015 -1527 -969
rect -1449 -1015 -1403 -969
rect -1325 -1015 -1279 -969
rect -1201 -1015 -1155 -969
rect -1077 -1015 -1031 -969
rect -953 -1015 -907 -969
rect -829 -1015 -783 -969
rect -705 -1015 -659 -969
rect -581 -1015 -535 -969
rect -457 -1015 -411 -969
rect -333 -1015 -287 -969
rect -209 -1015 -163 -969
rect -85 -1015 -39 -969
rect 39 -1015 85 -969
rect 163 -1015 209 -969
rect 287 -1015 333 -969
rect 411 -1015 457 -969
rect 535 -1015 581 -969
rect 659 -1015 705 -969
rect 783 -1015 829 -969
rect 907 -1015 953 -969
rect 1031 -1015 1077 -969
rect 1155 -1015 1201 -969
rect 1279 -1015 1325 -969
rect 1403 -1015 1449 -969
rect 1527 -1015 1573 -969
rect 1651 -1015 1697 -969
rect 1775 -1015 1821 -969
rect 1899 -1015 1945 -969
rect 2023 -1015 2069 -969
rect 2147 -1015 2193 -969
rect 2271 -1015 2317 -969
rect 2395 -1015 2441 -969
rect 2519 -1015 2565 -969
rect 2643 -1015 2689 -969
rect 2767 -1015 2813 -969
rect 2891 -1015 2937 -969
rect 3015 -1015 3061 -969
rect 3139 -1015 3185 -969
rect 3263 -1015 3309 -969
rect 3387 -1015 3433 -969
rect 3511 -1015 3557 -969
rect 3635 -1015 3681 -969
rect 3759 -1015 3805 -969
rect 3883 -1015 3929 -969
rect 4007 -1015 4053 -969
rect 4131 -1015 4177 -969
rect 4255 -1015 4301 -969
rect 4379 -1015 4425 -969
rect 4503 -1015 4549 -969
rect 4627 -1015 4673 -969
rect 4751 -1015 4797 -969
rect 4875 -1015 4921 -969
rect 4999 -1015 5045 -969
rect 5123 -1015 5169 -969
rect 5247 -1015 5293 -969
rect 5371 -1015 5417 -969
rect 5495 -1015 5541 -969
rect 5619 -1015 5665 -969
rect 5743 -1015 5789 -969
rect -5789 -1139 -5743 -1093
rect -5665 -1139 -5619 -1093
rect -5541 -1139 -5495 -1093
rect -5417 -1139 -5371 -1093
rect -5293 -1139 -5247 -1093
rect -5169 -1139 -5123 -1093
rect -5045 -1139 -4999 -1093
rect -4921 -1139 -4875 -1093
rect -4797 -1139 -4751 -1093
rect -4673 -1139 -4627 -1093
rect -4549 -1139 -4503 -1093
rect -4425 -1139 -4379 -1093
rect -4301 -1139 -4255 -1093
rect -4177 -1139 -4131 -1093
rect -4053 -1139 -4007 -1093
rect -3929 -1139 -3883 -1093
rect -3805 -1139 -3759 -1093
rect -3681 -1139 -3635 -1093
rect -3557 -1139 -3511 -1093
rect -3433 -1139 -3387 -1093
rect -3309 -1139 -3263 -1093
rect -3185 -1139 -3139 -1093
rect -3061 -1139 -3015 -1093
rect -2937 -1139 -2891 -1093
rect -2813 -1139 -2767 -1093
rect -2689 -1139 -2643 -1093
rect -2565 -1139 -2519 -1093
rect -2441 -1139 -2395 -1093
rect -2317 -1139 -2271 -1093
rect -2193 -1139 -2147 -1093
rect -2069 -1139 -2023 -1093
rect -1945 -1139 -1899 -1093
rect -1821 -1139 -1775 -1093
rect -1697 -1139 -1651 -1093
rect -1573 -1139 -1527 -1093
rect -1449 -1139 -1403 -1093
rect -1325 -1139 -1279 -1093
rect -1201 -1139 -1155 -1093
rect -1077 -1139 -1031 -1093
rect -953 -1139 -907 -1093
rect -829 -1139 -783 -1093
rect -705 -1139 -659 -1093
rect -581 -1139 -535 -1093
rect -457 -1139 -411 -1093
rect -333 -1139 -287 -1093
rect -209 -1139 -163 -1093
rect -85 -1139 -39 -1093
rect 39 -1139 85 -1093
rect 163 -1139 209 -1093
rect 287 -1139 333 -1093
rect 411 -1139 457 -1093
rect 535 -1139 581 -1093
rect 659 -1139 705 -1093
rect 783 -1139 829 -1093
rect 907 -1139 953 -1093
rect 1031 -1139 1077 -1093
rect 1155 -1139 1201 -1093
rect 1279 -1139 1325 -1093
rect 1403 -1139 1449 -1093
rect 1527 -1139 1573 -1093
rect 1651 -1139 1697 -1093
rect 1775 -1139 1821 -1093
rect 1899 -1139 1945 -1093
rect 2023 -1139 2069 -1093
rect 2147 -1139 2193 -1093
rect 2271 -1139 2317 -1093
rect 2395 -1139 2441 -1093
rect 2519 -1139 2565 -1093
rect 2643 -1139 2689 -1093
rect 2767 -1139 2813 -1093
rect 2891 -1139 2937 -1093
rect 3015 -1139 3061 -1093
rect 3139 -1139 3185 -1093
rect 3263 -1139 3309 -1093
rect 3387 -1139 3433 -1093
rect 3511 -1139 3557 -1093
rect 3635 -1139 3681 -1093
rect 3759 -1139 3805 -1093
rect 3883 -1139 3929 -1093
rect 4007 -1139 4053 -1093
rect 4131 -1139 4177 -1093
rect 4255 -1139 4301 -1093
rect 4379 -1139 4425 -1093
rect 4503 -1139 4549 -1093
rect 4627 -1139 4673 -1093
rect 4751 -1139 4797 -1093
rect 4875 -1139 4921 -1093
rect 4999 -1139 5045 -1093
rect 5123 -1139 5169 -1093
rect 5247 -1139 5293 -1093
rect 5371 -1139 5417 -1093
rect 5495 -1139 5541 -1093
rect 5619 -1139 5665 -1093
rect 5743 -1139 5789 -1093
rect -5789 -1263 -5743 -1217
rect -5665 -1263 -5619 -1217
rect -5541 -1263 -5495 -1217
rect -5417 -1263 -5371 -1217
rect -5293 -1263 -5247 -1217
rect -5169 -1263 -5123 -1217
rect -5045 -1263 -4999 -1217
rect -4921 -1263 -4875 -1217
rect -4797 -1263 -4751 -1217
rect -4673 -1263 -4627 -1217
rect -4549 -1263 -4503 -1217
rect -4425 -1263 -4379 -1217
rect -4301 -1263 -4255 -1217
rect -4177 -1263 -4131 -1217
rect -4053 -1263 -4007 -1217
rect -3929 -1263 -3883 -1217
rect -3805 -1263 -3759 -1217
rect -3681 -1263 -3635 -1217
rect -3557 -1263 -3511 -1217
rect -3433 -1263 -3387 -1217
rect -3309 -1263 -3263 -1217
rect -3185 -1263 -3139 -1217
rect -3061 -1263 -3015 -1217
rect -2937 -1263 -2891 -1217
rect -2813 -1263 -2767 -1217
rect -2689 -1263 -2643 -1217
rect -2565 -1263 -2519 -1217
rect -2441 -1263 -2395 -1217
rect -2317 -1263 -2271 -1217
rect -2193 -1263 -2147 -1217
rect -2069 -1263 -2023 -1217
rect -1945 -1263 -1899 -1217
rect -1821 -1263 -1775 -1217
rect -1697 -1263 -1651 -1217
rect -1573 -1263 -1527 -1217
rect -1449 -1263 -1403 -1217
rect -1325 -1263 -1279 -1217
rect -1201 -1263 -1155 -1217
rect -1077 -1263 -1031 -1217
rect -953 -1263 -907 -1217
rect -829 -1263 -783 -1217
rect -705 -1263 -659 -1217
rect -581 -1263 -535 -1217
rect -457 -1263 -411 -1217
rect -333 -1263 -287 -1217
rect -209 -1263 -163 -1217
rect -85 -1263 -39 -1217
rect 39 -1263 85 -1217
rect 163 -1263 209 -1217
rect 287 -1263 333 -1217
rect 411 -1263 457 -1217
rect 535 -1263 581 -1217
rect 659 -1263 705 -1217
rect 783 -1263 829 -1217
rect 907 -1263 953 -1217
rect 1031 -1263 1077 -1217
rect 1155 -1263 1201 -1217
rect 1279 -1263 1325 -1217
rect 1403 -1263 1449 -1217
rect 1527 -1263 1573 -1217
rect 1651 -1263 1697 -1217
rect 1775 -1263 1821 -1217
rect 1899 -1263 1945 -1217
rect 2023 -1263 2069 -1217
rect 2147 -1263 2193 -1217
rect 2271 -1263 2317 -1217
rect 2395 -1263 2441 -1217
rect 2519 -1263 2565 -1217
rect 2643 -1263 2689 -1217
rect 2767 -1263 2813 -1217
rect 2891 -1263 2937 -1217
rect 3015 -1263 3061 -1217
rect 3139 -1263 3185 -1217
rect 3263 -1263 3309 -1217
rect 3387 -1263 3433 -1217
rect 3511 -1263 3557 -1217
rect 3635 -1263 3681 -1217
rect 3759 -1263 3805 -1217
rect 3883 -1263 3929 -1217
rect 4007 -1263 4053 -1217
rect 4131 -1263 4177 -1217
rect 4255 -1263 4301 -1217
rect 4379 -1263 4425 -1217
rect 4503 -1263 4549 -1217
rect 4627 -1263 4673 -1217
rect 4751 -1263 4797 -1217
rect 4875 -1263 4921 -1217
rect 4999 -1263 5045 -1217
rect 5123 -1263 5169 -1217
rect 5247 -1263 5293 -1217
rect 5371 -1263 5417 -1217
rect 5495 -1263 5541 -1217
rect 5619 -1263 5665 -1217
rect 5743 -1263 5789 -1217
<< metal1 >>
rect -5800 1263 5800 1274
rect -5800 1217 -5789 1263
rect -5743 1217 -5665 1263
rect -5619 1217 -5541 1263
rect -5495 1217 -5417 1263
rect -5371 1217 -5293 1263
rect -5247 1217 -5169 1263
rect -5123 1217 -5045 1263
rect -4999 1217 -4921 1263
rect -4875 1217 -4797 1263
rect -4751 1217 -4673 1263
rect -4627 1217 -4549 1263
rect -4503 1217 -4425 1263
rect -4379 1217 -4301 1263
rect -4255 1217 -4177 1263
rect -4131 1217 -4053 1263
rect -4007 1217 -3929 1263
rect -3883 1217 -3805 1263
rect -3759 1217 -3681 1263
rect -3635 1217 -3557 1263
rect -3511 1217 -3433 1263
rect -3387 1217 -3309 1263
rect -3263 1217 -3185 1263
rect -3139 1217 -3061 1263
rect -3015 1217 -2937 1263
rect -2891 1217 -2813 1263
rect -2767 1217 -2689 1263
rect -2643 1217 -2565 1263
rect -2519 1217 -2441 1263
rect -2395 1217 -2317 1263
rect -2271 1217 -2193 1263
rect -2147 1217 -2069 1263
rect -2023 1217 -1945 1263
rect -1899 1217 -1821 1263
rect -1775 1217 -1697 1263
rect -1651 1217 -1573 1263
rect -1527 1217 -1449 1263
rect -1403 1217 -1325 1263
rect -1279 1217 -1201 1263
rect -1155 1217 -1077 1263
rect -1031 1217 -953 1263
rect -907 1217 -829 1263
rect -783 1217 -705 1263
rect -659 1217 -581 1263
rect -535 1217 -457 1263
rect -411 1217 -333 1263
rect -287 1217 -209 1263
rect -163 1217 -85 1263
rect -39 1217 39 1263
rect 85 1217 163 1263
rect 209 1217 287 1263
rect 333 1217 411 1263
rect 457 1217 535 1263
rect 581 1217 659 1263
rect 705 1217 783 1263
rect 829 1217 907 1263
rect 953 1217 1031 1263
rect 1077 1217 1155 1263
rect 1201 1217 1279 1263
rect 1325 1217 1403 1263
rect 1449 1217 1527 1263
rect 1573 1217 1651 1263
rect 1697 1217 1775 1263
rect 1821 1217 1899 1263
rect 1945 1217 2023 1263
rect 2069 1217 2147 1263
rect 2193 1217 2271 1263
rect 2317 1217 2395 1263
rect 2441 1217 2519 1263
rect 2565 1217 2643 1263
rect 2689 1217 2767 1263
rect 2813 1217 2891 1263
rect 2937 1217 3015 1263
rect 3061 1217 3139 1263
rect 3185 1217 3263 1263
rect 3309 1217 3387 1263
rect 3433 1217 3511 1263
rect 3557 1217 3635 1263
rect 3681 1217 3759 1263
rect 3805 1217 3883 1263
rect 3929 1217 4007 1263
rect 4053 1217 4131 1263
rect 4177 1217 4255 1263
rect 4301 1217 4379 1263
rect 4425 1217 4503 1263
rect 4549 1217 4627 1263
rect 4673 1217 4751 1263
rect 4797 1217 4875 1263
rect 4921 1217 4999 1263
rect 5045 1217 5123 1263
rect 5169 1217 5247 1263
rect 5293 1217 5371 1263
rect 5417 1217 5495 1263
rect 5541 1217 5619 1263
rect 5665 1217 5743 1263
rect 5789 1217 5800 1263
rect -5800 1139 5800 1217
rect -5800 1093 -5789 1139
rect -5743 1093 -5665 1139
rect -5619 1093 -5541 1139
rect -5495 1093 -5417 1139
rect -5371 1093 -5293 1139
rect -5247 1093 -5169 1139
rect -5123 1093 -5045 1139
rect -4999 1093 -4921 1139
rect -4875 1093 -4797 1139
rect -4751 1093 -4673 1139
rect -4627 1093 -4549 1139
rect -4503 1093 -4425 1139
rect -4379 1093 -4301 1139
rect -4255 1093 -4177 1139
rect -4131 1093 -4053 1139
rect -4007 1093 -3929 1139
rect -3883 1093 -3805 1139
rect -3759 1093 -3681 1139
rect -3635 1093 -3557 1139
rect -3511 1093 -3433 1139
rect -3387 1093 -3309 1139
rect -3263 1093 -3185 1139
rect -3139 1093 -3061 1139
rect -3015 1093 -2937 1139
rect -2891 1093 -2813 1139
rect -2767 1093 -2689 1139
rect -2643 1093 -2565 1139
rect -2519 1093 -2441 1139
rect -2395 1093 -2317 1139
rect -2271 1093 -2193 1139
rect -2147 1093 -2069 1139
rect -2023 1093 -1945 1139
rect -1899 1093 -1821 1139
rect -1775 1093 -1697 1139
rect -1651 1093 -1573 1139
rect -1527 1093 -1449 1139
rect -1403 1093 -1325 1139
rect -1279 1093 -1201 1139
rect -1155 1093 -1077 1139
rect -1031 1093 -953 1139
rect -907 1093 -829 1139
rect -783 1093 -705 1139
rect -659 1093 -581 1139
rect -535 1093 -457 1139
rect -411 1093 -333 1139
rect -287 1093 -209 1139
rect -163 1093 -85 1139
rect -39 1093 39 1139
rect 85 1093 163 1139
rect 209 1093 287 1139
rect 333 1093 411 1139
rect 457 1093 535 1139
rect 581 1093 659 1139
rect 705 1093 783 1139
rect 829 1093 907 1139
rect 953 1093 1031 1139
rect 1077 1093 1155 1139
rect 1201 1093 1279 1139
rect 1325 1093 1403 1139
rect 1449 1093 1527 1139
rect 1573 1093 1651 1139
rect 1697 1093 1775 1139
rect 1821 1093 1899 1139
rect 1945 1093 2023 1139
rect 2069 1093 2147 1139
rect 2193 1093 2271 1139
rect 2317 1093 2395 1139
rect 2441 1093 2519 1139
rect 2565 1093 2643 1139
rect 2689 1093 2767 1139
rect 2813 1093 2891 1139
rect 2937 1093 3015 1139
rect 3061 1093 3139 1139
rect 3185 1093 3263 1139
rect 3309 1093 3387 1139
rect 3433 1093 3511 1139
rect 3557 1093 3635 1139
rect 3681 1093 3759 1139
rect 3805 1093 3883 1139
rect 3929 1093 4007 1139
rect 4053 1093 4131 1139
rect 4177 1093 4255 1139
rect 4301 1093 4379 1139
rect 4425 1093 4503 1139
rect 4549 1093 4627 1139
rect 4673 1093 4751 1139
rect 4797 1093 4875 1139
rect 4921 1093 4999 1139
rect 5045 1093 5123 1139
rect 5169 1093 5247 1139
rect 5293 1093 5371 1139
rect 5417 1093 5495 1139
rect 5541 1093 5619 1139
rect 5665 1093 5743 1139
rect 5789 1093 5800 1139
rect -5800 1015 5800 1093
rect -5800 969 -5789 1015
rect -5743 969 -5665 1015
rect -5619 969 -5541 1015
rect -5495 969 -5417 1015
rect -5371 969 -5293 1015
rect -5247 969 -5169 1015
rect -5123 969 -5045 1015
rect -4999 969 -4921 1015
rect -4875 969 -4797 1015
rect -4751 969 -4673 1015
rect -4627 969 -4549 1015
rect -4503 969 -4425 1015
rect -4379 969 -4301 1015
rect -4255 969 -4177 1015
rect -4131 969 -4053 1015
rect -4007 969 -3929 1015
rect -3883 969 -3805 1015
rect -3759 969 -3681 1015
rect -3635 969 -3557 1015
rect -3511 969 -3433 1015
rect -3387 969 -3309 1015
rect -3263 969 -3185 1015
rect -3139 969 -3061 1015
rect -3015 969 -2937 1015
rect -2891 969 -2813 1015
rect -2767 969 -2689 1015
rect -2643 969 -2565 1015
rect -2519 969 -2441 1015
rect -2395 969 -2317 1015
rect -2271 969 -2193 1015
rect -2147 969 -2069 1015
rect -2023 969 -1945 1015
rect -1899 969 -1821 1015
rect -1775 969 -1697 1015
rect -1651 969 -1573 1015
rect -1527 969 -1449 1015
rect -1403 969 -1325 1015
rect -1279 969 -1201 1015
rect -1155 969 -1077 1015
rect -1031 969 -953 1015
rect -907 969 -829 1015
rect -783 969 -705 1015
rect -659 969 -581 1015
rect -535 969 -457 1015
rect -411 969 -333 1015
rect -287 969 -209 1015
rect -163 969 -85 1015
rect -39 969 39 1015
rect 85 969 163 1015
rect 209 969 287 1015
rect 333 969 411 1015
rect 457 969 535 1015
rect 581 969 659 1015
rect 705 969 783 1015
rect 829 969 907 1015
rect 953 969 1031 1015
rect 1077 969 1155 1015
rect 1201 969 1279 1015
rect 1325 969 1403 1015
rect 1449 969 1527 1015
rect 1573 969 1651 1015
rect 1697 969 1775 1015
rect 1821 969 1899 1015
rect 1945 969 2023 1015
rect 2069 969 2147 1015
rect 2193 969 2271 1015
rect 2317 969 2395 1015
rect 2441 969 2519 1015
rect 2565 969 2643 1015
rect 2689 969 2767 1015
rect 2813 969 2891 1015
rect 2937 969 3015 1015
rect 3061 969 3139 1015
rect 3185 969 3263 1015
rect 3309 969 3387 1015
rect 3433 969 3511 1015
rect 3557 969 3635 1015
rect 3681 969 3759 1015
rect 3805 969 3883 1015
rect 3929 969 4007 1015
rect 4053 969 4131 1015
rect 4177 969 4255 1015
rect 4301 969 4379 1015
rect 4425 969 4503 1015
rect 4549 969 4627 1015
rect 4673 969 4751 1015
rect 4797 969 4875 1015
rect 4921 969 4999 1015
rect 5045 969 5123 1015
rect 5169 969 5247 1015
rect 5293 969 5371 1015
rect 5417 969 5495 1015
rect 5541 969 5619 1015
rect 5665 969 5743 1015
rect 5789 969 5800 1015
rect -5800 891 5800 969
rect -5800 845 -5789 891
rect -5743 845 -5665 891
rect -5619 845 -5541 891
rect -5495 845 -5417 891
rect -5371 845 -5293 891
rect -5247 845 -5169 891
rect -5123 845 -5045 891
rect -4999 845 -4921 891
rect -4875 845 -4797 891
rect -4751 845 -4673 891
rect -4627 845 -4549 891
rect -4503 845 -4425 891
rect -4379 845 -4301 891
rect -4255 845 -4177 891
rect -4131 845 -4053 891
rect -4007 845 -3929 891
rect -3883 845 -3805 891
rect -3759 845 -3681 891
rect -3635 845 -3557 891
rect -3511 845 -3433 891
rect -3387 845 -3309 891
rect -3263 845 -3185 891
rect -3139 845 -3061 891
rect -3015 845 -2937 891
rect -2891 845 -2813 891
rect -2767 845 -2689 891
rect -2643 845 -2565 891
rect -2519 845 -2441 891
rect -2395 845 -2317 891
rect -2271 845 -2193 891
rect -2147 845 -2069 891
rect -2023 845 -1945 891
rect -1899 845 -1821 891
rect -1775 845 -1697 891
rect -1651 845 -1573 891
rect -1527 845 -1449 891
rect -1403 845 -1325 891
rect -1279 845 -1201 891
rect -1155 845 -1077 891
rect -1031 845 -953 891
rect -907 845 -829 891
rect -783 845 -705 891
rect -659 845 -581 891
rect -535 845 -457 891
rect -411 845 -333 891
rect -287 845 -209 891
rect -163 845 -85 891
rect -39 845 39 891
rect 85 845 163 891
rect 209 845 287 891
rect 333 845 411 891
rect 457 845 535 891
rect 581 845 659 891
rect 705 845 783 891
rect 829 845 907 891
rect 953 845 1031 891
rect 1077 845 1155 891
rect 1201 845 1279 891
rect 1325 845 1403 891
rect 1449 845 1527 891
rect 1573 845 1651 891
rect 1697 845 1775 891
rect 1821 845 1899 891
rect 1945 845 2023 891
rect 2069 845 2147 891
rect 2193 845 2271 891
rect 2317 845 2395 891
rect 2441 845 2519 891
rect 2565 845 2643 891
rect 2689 845 2767 891
rect 2813 845 2891 891
rect 2937 845 3015 891
rect 3061 845 3139 891
rect 3185 845 3263 891
rect 3309 845 3387 891
rect 3433 845 3511 891
rect 3557 845 3635 891
rect 3681 845 3759 891
rect 3805 845 3883 891
rect 3929 845 4007 891
rect 4053 845 4131 891
rect 4177 845 4255 891
rect 4301 845 4379 891
rect 4425 845 4503 891
rect 4549 845 4627 891
rect 4673 845 4751 891
rect 4797 845 4875 891
rect 4921 845 4999 891
rect 5045 845 5123 891
rect 5169 845 5247 891
rect 5293 845 5371 891
rect 5417 845 5495 891
rect 5541 845 5619 891
rect 5665 845 5743 891
rect 5789 845 5800 891
rect -5800 767 5800 845
rect -5800 721 -5789 767
rect -5743 721 -5665 767
rect -5619 721 -5541 767
rect -5495 721 -5417 767
rect -5371 721 -5293 767
rect -5247 721 -5169 767
rect -5123 721 -5045 767
rect -4999 721 -4921 767
rect -4875 721 -4797 767
rect -4751 721 -4673 767
rect -4627 721 -4549 767
rect -4503 721 -4425 767
rect -4379 721 -4301 767
rect -4255 721 -4177 767
rect -4131 721 -4053 767
rect -4007 721 -3929 767
rect -3883 721 -3805 767
rect -3759 721 -3681 767
rect -3635 721 -3557 767
rect -3511 721 -3433 767
rect -3387 721 -3309 767
rect -3263 721 -3185 767
rect -3139 721 -3061 767
rect -3015 721 -2937 767
rect -2891 721 -2813 767
rect -2767 721 -2689 767
rect -2643 721 -2565 767
rect -2519 721 -2441 767
rect -2395 721 -2317 767
rect -2271 721 -2193 767
rect -2147 721 -2069 767
rect -2023 721 -1945 767
rect -1899 721 -1821 767
rect -1775 721 -1697 767
rect -1651 721 -1573 767
rect -1527 721 -1449 767
rect -1403 721 -1325 767
rect -1279 721 -1201 767
rect -1155 721 -1077 767
rect -1031 721 -953 767
rect -907 721 -829 767
rect -783 721 -705 767
rect -659 721 -581 767
rect -535 721 -457 767
rect -411 721 -333 767
rect -287 721 -209 767
rect -163 721 -85 767
rect -39 721 39 767
rect 85 721 163 767
rect 209 721 287 767
rect 333 721 411 767
rect 457 721 535 767
rect 581 721 659 767
rect 705 721 783 767
rect 829 721 907 767
rect 953 721 1031 767
rect 1077 721 1155 767
rect 1201 721 1279 767
rect 1325 721 1403 767
rect 1449 721 1527 767
rect 1573 721 1651 767
rect 1697 721 1775 767
rect 1821 721 1899 767
rect 1945 721 2023 767
rect 2069 721 2147 767
rect 2193 721 2271 767
rect 2317 721 2395 767
rect 2441 721 2519 767
rect 2565 721 2643 767
rect 2689 721 2767 767
rect 2813 721 2891 767
rect 2937 721 3015 767
rect 3061 721 3139 767
rect 3185 721 3263 767
rect 3309 721 3387 767
rect 3433 721 3511 767
rect 3557 721 3635 767
rect 3681 721 3759 767
rect 3805 721 3883 767
rect 3929 721 4007 767
rect 4053 721 4131 767
rect 4177 721 4255 767
rect 4301 721 4379 767
rect 4425 721 4503 767
rect 4549 721 4627 767
rect 4673 721 4751 767
rect 4797 721 4875 767
rect 4921 721 4999 767
rect 5045 721 5123 767
rect 5169 721 5247 767
rect 5293 721 5371 767
rect 5417 721 5495 767
rect 5541 721 5619 767
rect 5665 721 5743 767
rect 5789 721 5800 767
rect -5800 643 5800 721
rect -5800 597 -5789 643
rect -5743 597 -5665 643
rect -5619 597 -5541 643
rect -5495 597 -5417 643
rect -5371 597 -5293 643
rect -5247 597 -5169 643
rect -5123 597 -5045 643
rect -4999 597 -4921 643
rect -4875 597 -4797 643
rect -4751 597 -4673 643
rect -4627 597 -4549 643
rect -4503 597 -4425 643
rect -4379 597 -4301 643
rect -4255 597 -4177 643
rect -4131 597 -4053 643
rect -4007 597 -3929 643
rect -3883 597 -3805 643
rect -3759 597 -3681 643
rect -3635 597 -3557 643
rect -3511 597 -3433 643
rect -3387 597 -3309 643
rect -3263 597 -3185 643
rect -3139 597 -3061 643
rect -3015 597 -2937 643
rect -2891 597 -2813 643
rect -2767 597 -2689 643
rect -2643 597 -2565 643
rect -2519 597 -2441 643
rect -2395 597 -2317 643
rect -2271 597 -2193 643
rect -2147 597 -2069 643
rect -2023 597 -1945 643
rect -1899 597 -1821 643
rect -1775 597 -1697 643
rect -1651 597 -1573 643
rect -1527 597 -1449 643
rect -1403 597 -1325 643
rect -1279 597 -1201 643
rect -1155 597 -1077 643
rect -1031 597 -953 643
rect -907 597 -829 643
rect -783 597 -705 643
rect -659 597 -581 643
rect -535 597 -457 643
rect -411 597 -333 643
rect -287 597 -209 643
rect -163 597 -85 643
rect -39 597 39 643
rect 85 597 163 643
rect 209 597 287 643
rect 333 597 411 643
rect 457 597 535 643
rect 581 597 659 643
rect 705 597 783 643
rect 829 597 907 643
rect 953 597 1031 643
rect 1077 597 1155 643
rect 1201 597 1279 643
rect 1325 597 1403 643
rect 1449 597 1527 643
rect 1573 597 1651 643
rect 1697 597 1775 643
rect 1821 597 1899 643
rect 1945 597 2023 643
rect 2069 597 2147 643
rect 2193 597 2271 643
rect 2317 597 2395 643
rect 2441 597 2519 643
rect 2565 597 2643 643
rect 2689 597 2767 643
rect 2813 597 2891 643
rect 2937 597 3015 643
rect 3061 597 3139 643
rect 3185 597 3263 643
rect 3309 597 3387 643
rect 3433 597 3511 643
rect 3557 597 3635 643
rect 3681 597 3759 643
rect 3805 597 3883 643
rect 3929 597 4007 643
rect 4053 597 4131 643
rect 4177 597 4255 643
rect 4301 597 4379 643
rect 4425 597 4503 643
rect 4549 597 4627 643
rect 4673 597 4751 643
rect 4797 597 4875 643
rect 4921 597 4999 643
rect 5045 597 5123 643
rect 5169 597 5247 643
rect 5293 597 5371 643
rect 5417 597 5495 643
rect 5541 597 5619 643
rect 5665 597 5743 643
rect 5789 597 5800 643
rect -5800 519 5800 597
rect -5800 473 -5789 519
rect -5743 473 -5665 519
rect -5619 473 -5541 519
rect -5495 473 -5417 519
rect -5371 473 -5293 519
rect -5247 473 -5169 519
rect -5123 473 -5045 519
rect -4999 473 -4921 519
rect -4875 473 -4797 519
rect -4751 473 -4673 519
rect -4627 473 -4549 519
rect -4503 473 -4425 519
rect -4379 473 -4301 519
rect -4255 473 -4177 519
rect -4131 473 -4053 519
rect -4007 473 -3929 519
rect -3883 473 -3805 519
rect -3759 473 -3681 519
rect -3635 473 -3557 519
rect -3511 473 -3433 519
rect -3387 473 -3309 519
rect -3263 473 -3185 519
rect -3139 473 -3061 519
rect -3015 473 -2937 519
rect -2891 473 -2813 519
rect -2767 473 -2689 519
rect -2643 473 -2565 519
rect -2519 473 -2441 519
rect -2395 473 -2317 519
rect -2271 473 -2193 519
rect -2147 473 -2069 519
rect -2023 473 -1945 519
rect -1899 473 -1821 519
rect -1775 473 -1697 519
rect -1651 473 -1573 519
rect -1527 473 -1449 519
rect -1403 473 -1325 519
rect -1279 473 -1201 519
rect -1155 473 -1077 519
rect -1031 473 -953 519
rect -907 473 -829 519
rect -783 473 -705 519
rect -659 473 -581 519
rect -535 473 -457 519
rect -411 473 -333 519
rect -287 473 -209 519
rect -163 473 -85 519
rect -39 473 39 519
rect 85 473 163 519
rect 209 473 287 519
rect 333 473 411 519
rect 457 473 535 519
rect 581 473 659 519
rect 705 473 783 519
rect 829 473 907 519
rect 953 473 1031 519
rect 1077 473 1155 519
rect 1201 473 1279 519
rect 1325 473 1403 519
rect 1449 473 1527 519
rect 1573 473 1651 519
rect 1697 473 1775 519
rect 1821 473 1899 519
rect 1945 473 2023 519
rect 2069 473 2147 519
rect 2193 473 2271 519
rect 2317 473 2395 519
rect 2441 473 2519 519
rect 2565 473 2643 519
rect 2689 473 2767 519
rect 2813 473 2891 519
rect 2937 473 3015 519
rect 3061 473 3139 519
rect 3185 473 3263 519
rect 3309 473 3387 519
rect 3433 473 3511 519
rect 3557 473 3635 519
rect 3681 473 3759 519
rect 3805 473 3883 519
rect 3929 473 4007 519
rect 4053 473 4131 519
rect 4177 473 4255 519
rect 4301 473 4379 519
rect 4425 473 4503 519
rect 4549 473 4627 519
rect 4673 473 4751 519
rect 4797 473 4875 519
rect 4921 473 4999 519
rect 5045 473 5123 519
rect 5169 473 5247 519
rect 5293 473 5371 519
rect 5417 473 5495 519
rect 5541 473 5619 519
rect 5665 473 5743 519
rect 5789 473 5800 519
rect -5800 395 5800 473
rect -5800 349 -5789 395
rect -5743 349 -5665 395
rect -5619 349 -5541 395
rect -5495 349 -5417 395
rect -5371 349 -5293 395
rect -5247 349 -5169 395
rect -5123 349 -5045 395
rect -4999 349 -4921 395
rect -4875 349 -4797 395
rect -4751 349 -4673 395
rect -4627 349 -4549 395
rect -4503 349 -4425 395
rect -4379 349 -4301 395
rect -4255 349 -4177 395
rect -4131 349 -4053 395
rect -4007 349 -3929 395
rect -3883 349 -3805 395
rect -3759 349 -3681 395
rect -3635 349 -3557 395
rect -3511 349 -3433 395
rect -3387 349 -3309 395
rect -3263 349 -3185 395
rect -3139 349 -3061 395
rect -3015 349 -2937 395
rect -2891 349 -2813 395
rect -2767 349 -2689 395
rect -2643 349 -2565 395
rect -2519 349 -2441 395
rect -2395 349 -2317 395
rect -2271 349 -2193 395
rect -2147 349 -2069 395
rect -2023 349 -1945 395
rect -1899 349 -1821 395
rect -1775 349 -1697 395
rect -1651 349 -1573 395
rect -1527 349 -1449 395
rect -1403 349 -1325 395
rect -1279 349 -1201 395
rect -1155 349 -1077 395
rect -1031 349 -953 395
rect -907 349 -829 395
rect -783 349 -705 395
rect -659 349 -581 395
rect -535 349 -457 395
rect -411 349 -333 395
rect -287 349 -209 395
rect -163 349 -85 395
rect -39 349 39 395
rect 85 349 163 395
rect 209 349 287 395
rect 333 349 411 395
rect 457 349 535 395
rect 581 349 659 395
rect 705 349 783 395
rect 829 349 907 395
rect 953 349 1031 395
rect 1077 349 1155 395
rect 1201 349 1279 395
rect 1325 349 1403 395
rect 1449 349 1527 395
rect 1573 349 1651 395
rect 1697 349 1775 395
rect 1821 349 1899 395
rect 1945 349 2023 395
rect 2069 349 2147 395
rect 2193 349 2271 395
rect 2317 349 2395 395
rect 2441 349 2519 395
rect 2565 349 2643 395
rect 2689 349 2767 395
rect 2813 349 2891 395
rect 2937 349 3015 395
rect 3061 349 3139 395
rect 3185 349 3263 395
rect 3309 349 3387 395
rect 3433 349 3511 395
rect 3557 349 3635 395
rect 3681 349 3759 395
rect 3805 349 3883 395
rect 3929 349 4007 395
rect 4053 349 4131 395
rect 4177 349 4255 395
rect 4301 349 4379 395
rect 4425 349 4503 395
rect 4549 349 4627 395
rect 4673 349 4751 395
rect 4797 349 4875 395
rect 4921 349 4999 395
rect 5045 349 5123 395
rect 5169 349 5247 395
rect 5293 349 5371 395
rect 5417 349 5495 395
rect 5541 349 5619 395
rect 5665 349 5743 395
rect 5789 349 5800 395
rect -5800 271 5800 349
rect -5800 225 -5789 271
rect -5743 225 -5665 271
rect -5619 225 -5541 271
rect -5495 225 -5417 271
rect -5371 225 -5293 271
rect -5247 225 -5169 271
rect -5123 225 -5045 271
rect -4999 225 -4921 271
rect -4875 225 -4797 271
rect -4751 225 -4673 271
rect -4627 225 -4549 271
rect -4503 225 -4425 271
rect -4379 225 -4301 271
rect -4255 225 -4177 271
rect -4131 225 -4053 271
rect -4007 225 -3929 271
rect -3883 225 -3805 271
rect -3759 225 -3681 271
rect -3635 225 -3557 271
rect -3511 225 -3433 271
rect -3387 225 -3309 271
rect -3263 225 -3185 271
rect -3139 225 -3061 271
rect -3015 225 -2937 271
rect -2891 225 -2813 271
rect -2767 225 -2689 271
rect -2643 225 -2565 271
rect -2519 225 -2441 271
rect -2395 225 -2317 271
rect -2271 225 -2193 271
rect -2147 225 -2069 271
rect -2023 225 -1945 271
rect -1899 225 -1821 271
rect -1775 225 -1697 271
rect -1651 225 -1573 271
rect -1527 225 -1449 271
rect -1403 225 -1325 271
rect -1279 225 -1201 271
rect -1155 225 -1077 271
rect -1031 225 -953 271
rect -907 225 -829 271
rect -783 225 -705 271
rect -659 225 -581 271
rect -535 225 -457 271
rect -411 225 -333 271
rect -287 225 -209 271
rect -163 225 -85 271
rect -39 225 39 271
rect 85 225 163 271
rect 209 225 287 271
rect 333 225 411 271
rect 457 225 535 271
rect 581 225 659 271
rect 705 225 783 271
rect 829 225 907 271
rect 953 225 1031 271
rect 1077 225 1155 271
rect 1201 225 1279 271
rect 1325 225 1403 271
rect 1449 225 1527 271
rect 1573 225 1651 271
rect 1697 225 1775 271
rect 1821 225 1899 271
rect 1945 225 2023 271
rect 2069 225 2147 271
rect 2193 225 2271 271
rect 2317 225 2395 271
rect 2441 225 2519 271
rect 2565 225 2643 271
rect 2689 225 2767 271
rect 2813 225 2891 271
rect 2937 225 3015 271
rect 3061 225 3139 271
rect 3185 225 3263 271
rect 3309 225 3387 271
rect 3433 225 3511 271
rect 3557 225 3635 271
rect 3681 225 3759 271
rect 3805 225 3883 271
rect 3929 225 4007 271
rect 4053 225 4131 271
rect 4177 225 4255 271
rect 4301 225 4379 271
rect 4425 225 4503 271
rect 4549 225 4627 271
rect 4673 225 4751 271
rect 4797 225 4875 271
rect 4921 225 4999 271
rect 5045 225 5123 271
rect 5169 225 5247 271
rect 5293 225 5371 271
rect 5417 225 5495 271
rect 5541 225 5619 271
rect 5665 225 5743 271
rect 5789 225 5800 271
rect -5800 147 5800 225
rect -5800 101 -5789 147
rect -5743 101 -5665 147
rect -5619 101 -5541 147
rect -5495 101 -5417 147
rect -5371 101 -5293 147
rect -5247 101 -5169 147
rect -5123 101 -5045 147
rect -4999 101 -4921 147
rect -4875 101 -4797 147
rect -4751 101 -4673 147
rect -4627 101 -4549 147
rect -4503 101 -4425 147
rect -4379 101 -4301 147
rect -4255 101 -4177 147
rect -4131 101 -4053 147
rect -4007 101 -3929 147
rect -3883 101 -3805 147
rect -3759 101 -3681 147
rect -3635 101 -3557 147
rect -3511 101 -3433 147
rect -3387 101 -3309 147
rect -3263 101 -3185 147
rect -3139 101 -3061 147
rect -3015 101 -2937 147
rect -2891 101 -2813 147
rect -2767 101 -2689 147
rect -2643 101 -2565 147
rect -2519 101 -2441 147
rect -2395 101 -2317 147
rect -2271 101 -2193 147
rect -2147 101 -2069 147
rect -2023 101 -1945 147
rect -1899 101 -1821 147
rect -1775 101 -1697 147
rect -1651 101 -1573 147
rect -1527 101 -1449 147
rect -1403 101 -1325 147
rect -1279 101 -1201 147
rect -1155 101 -1077 147
rect -1031 101 -953 147
rect -907 101 -829 147
rect -783 101 -705 147
rect -659 101 -581 147
rect -535 101 -457 147
rect -411 101 -333 147
rect -287 101 -209 147
rect -163 101 -85 147
rect -39 101 39 147
rect 85 101 163 147
rect 209 101 287 147
rect 333 101 411 147
rect 457 101 535 147
rect 581 101 659 147
rect 705 101 783 147
rect 829 101 907 147
rect 953 101 1031 147
rect 1077 101 1155 147
rect 1201 101 1279 147
rect 1325 101 1403 147
rect 1449 101 1527 147
rect 1573 101 1651 147
rect 1697 101 1775 147
rect 1821 101 1899 147
rect 1945 101 2023 147
rect 2069 101 2147 147
rect 2193 101 2271 147
rect 2317 101 2395 147
rect 2441 101 2519 147
rect 2565 101 2643 147
rect 2689 101 2767 147
rect 2813 101 2891 147
rect 2937 101 3015 147
rect 3061 101 3139 147
rect 3185 101 3263 147
rect 3309 101 3387 147
rect 3433 101 3511 147
rect 3557 101 3635 147
rect 3681 101 3759 147
rect 3805 101 3883 147
rect 3929 101 4007 147
rect 4053 101 4131 147
rect 4177 101 4255 147
rect 4301 101 4379 147
rect 4425 101 4503 147
rect 4549 101 4627 147
rect 4673 101 4751 147
rect 4797 101 4875 147
rect 4921 101 4999 147
rect 5045 101 5123 147
rect 5169 101 5247 147
rect 5293 101 5371 147
rect 5417 101 5495 147
rect 5541 101 5619 147
rect 5665 101 5743 147
rect 5789 101 5800 147
rect -5800 23 5800 101
rect -5800 -23 -5789 23
rect -5743 -23 -5665 23
rect -5619 -23 -5541 23
rect -5495 -23 -5417 23
rect -5371 -23 -5293 23
rect -5247 -23 -5169 23
rect -5123 -23 -5045 23
rect -4999 -23 -4921 23
rect -4875 -23 -4797 23
rect -4751 -23 -4673 23
rect -4627 -23 -4549 23
rect -4503 -23 -4425 23
rect -4379 -23 -4301 23
rect -4255 -23 -4177 23
rect -4131 -23 -4053 23
rect -4007 -23 -3929 23
rect -3883 -23 -3805 23
rect -3759 -23 -3681 23
rect -3635 -23 -3557 23
rect -3511 -23 -3433 23
rect -3387 -23 -3309 23
rect -3263 -23 -3185 23
rect -3139 -23 -3061 23
rect -3015 -23 -2937 23
rect -2891 -23 -2813 23
rect -2767 -23 -2689 23
rect -2643 -23 -2565 23
rect -2519 -23 -2441 23
rect -2395 -23 -2317 23
rect -2271 -23 -2193 23
rect -2147 -23 -2069 23
rect -2023 -23 -1945 23
rect -1899 -23 -1821 23
rect -1775 -23 -1697 23
rect -1651 -23 -1573 23
rect -1527 -23 -1449 23
rect -1403 -23 -1325 23
rect -1279 -23 -1201 23
rect -1155 -23 -1077 23
rect -1031 -23 -953 23
rect -907 -23 -829 23
rect -783 -23 -705 23
rect -659 -23 -581 23
rect -535 -23 -457 23
rect -411 -23 -333 23
rect -287 -23 -209 23
rect -163 -23 -85 23
rect -39 -23 39 23
rect 85 -23 163 23
rect 209 -23 287 23
rect 333 -23 411 23
rect 457 -23 535 23
rect 581 -23 659 23
rect 705 -23 783 23
rect 829 -23 907 23
rect 953 -23 1031 23
rect 1077 -23 1155 23
rect 1201 -23 1279 23
rect 1325 -23 1403 23
rect 1449 -23 1527 23
rect 1573 -23 1651 23
rect 1697 -23 1775 23
rect 1821 -23 1899 23
rect 1945 -23 2023 23
rect 2069 -23 2147 23
rect 2193 -23 2271 23
rect 2317 -23 2395 23
rect 2441 -23 2519 23
rect 2565 -23 2643 23
rect 2689 -23 2767 23
rect 2813 -23 2891 23
rect 2937 -23 3015 23
rect 3061 -23 3139 23
rect 3185 -23 3263 23
rect 3309 -23 3387 23
rect 3433 -23 3511 23
rect 3557 -23 3635 23
rect 3681 -23 3759 23
rect 3805 -23 3883 23
rect 3929 -23 4007 23
rect 4053 -23 4131 23
rect 4177 -23 4255 23
rect 4301 -23 4379 23
rect 4425 -23 4503 23
rect 4549 -23 4627 23
rect 4673 -23 4751 23
rect 4797 -23 4875 23
rect 4921 -23 4999 23
rect 5045 -23 5123 23
rect 5169 -23 5247 23
rect 5293 -23 5371 23
rect 5417 -23 5495 23
rect 5541 -23 5619 23
rect 5665 -23 5743 23
rect 5789 -23 5800 23
rect -5800 -101 5800 -23
rect -5800 -147 -5789 -101
rect -5743 -147 -5665 -101
rect -5619 -147 -5541 -101
rect -5495 -147 -5417 -101
rect -5371 -147 -5293 -101
rect -5247 -147 -5169 -101
rect -5123 -147 -5045 -101
rect -4999 -147 -4921 -101
rect -4875 -147 -4797 -101
rect -4751 -147 -4673 -101
rect -4627 -147 -4549 -101
rect -4503 -147 -4425 -101
rect -4379 -147 -4301 -101
rect -4255 -147 -4177 -101
rect -4131 -147 -4053 -101
rect -4007 -147 -3929 -101
rect -3883 -147 -3805 -101
rect -3759 -147 -3681 -101
rect -3635 -147 -3557 -101
rect -3511 -147 -3433 -101
rect -3387 -147 -3309 -101
rect -3263 -147 -3185 -101
rect -3139 -147 -3061 -101
rect -3015 -147 -2937 -101
rect -2891 -147 -2813 -101
rect -2767 -147 -2689 -101
rect -2643 -147 -2565 -101
rect -2519 -147 -2441 -101
rect -2395 -147 -2317 -101
rect -2271 -147 -2193 -101
rect -2147 -147 -2069 -101
rect -2023 -147 -1945 -101
rect -1899 -147 -1821 -101
rect -1775 -147 -1697 -101
rect -1651 -147 -1573 -101
rect -1527 -147 -1449 -101
rect -1403 -147 -1325 -101
rect -1279 -147 -1201 -101
rect -1155 -147 -1077 -101
rect -1031 -147 -953 -101
rect -907 -147 -829 -101
rect -783 -147 -705 -101
rect -659 -147 -581 -101
rect -535 -147 -457 -101
rect -411 -147 -333 -101
rect -287 -147 -209 -101
rect -163 -147 -85 -101
rect -39 -147 39 -101
rect 85 -147 163 -101
rect 209 -147 287 -101
rect 333 -147 411 -101
rect 457 -147 535 -101
rect 581 -147 659 -101
rect 705 -147 783 -101
rect 829 -147 907 -101
rect 953 -147 1031 -101
rect 1077 -147 1155 -101
rect 1201 -147 1279 -101
rect 1325 -147 1403 -101
rect 1449 -147 1527 -101
rect 1573 -147 1651 -101
rect 1697 -147 1775 -101
rect 1821 -147 1899 -101
rect 1945 -147 2023 -101
rect 2069 -147 2147 -101
rect 2193 -147 2271 -101
rect 2317 -147 2395 -101
rect 2441 -147 2519 -101
rect 2565 -147 2643 -101
rect 2689 -147 2767 -101
rect 2813 -147 2891 -101
rect 2937 -147 3015 -101
rect 3061 -147 3139 -101
rect 3185 -147 3263 -101
rect 3309 -147 3387 -101
rect 3433 -147 3511 -101
rect 3557 -147 3635 -101
rect 3681 -147 3759 -101
rect 3805 -147 3883 -101
rect 3929 -147 4007 -101
rect 4053 -147 4131 -101
rect 4177 -147 4255 -101
rect 4301 -147 4379 -101
rect 4425 -147 4503 -101
rect 4549 -147 4627 -101
rect 4673 -147 4751 -101
rect 4797 -147 4875 -101
rect 4921 -147 4999 -101
rect 5045 -147 5123 -101
rect 5169 -147 5247 -101
rect 5293 -147 5371 -101
rect 5417 -147 5495 -101
rect 5541 -147 5619 -101
rect 5665 -147 5743 -101
rect 5789 -147 5800 -101
rect -5800 -225 5800 -147
rect -5800 -271 -5789 -225
rect -5743 -271 -5665 -225
rect -5619 -271 -5541 -225
rect -5495 -271 -5417 -225
rect -5371 -271 -5293 -225
rect -5247 -271 -5169 -225
rect -5123 -271 -5045 -225
rect -4999 -271 -4921 -225
rect -4875 -271 -4797 -225
rect -4751 -271 -4673 -225
rect -4627 -271 -4549 -225
rect -4503 -271 -4425 -225
rect -4379 -271 -4301 -225
rect -4255 -271 -4177 -225
rect -4131 -271 -4053 -225
rect -4007 -271 -3929 -225
rect -3883 -271 -3805 -225
rect -3759 -271 -3681 -225
rect -3635 -271 -3557 -225
rect -3511 -271 -3433 -225
rect -3387 -271 -3309 -225
rect -3263 -271 -3185 -225
rect -3139 -271 -3061 -225
rect -3015 -271 -2937 -225
rect -2891 -271 -2813 -225
rect -2767 -271 -2689 -225
rect -2643 -271 -2565 -225
rect -2519 -271 -2441 -225
rect -2395 -271 -2317 -225
rect -2271 -271 -2193 -225
rect -2147 -271 -2069 -225
rect -2023 -271 -1945 -225
rect -1899 -271 -1821 -225
rect -1775 -271 -1697 -225
rect -1651 -271 -1573 -225
rect -1527 -271 -1449 -225
rect -1403 -271 -1325 -225
rect -1279 -271 -1201 -225
rect -1155 -271 -1077 -225
rect -1031 -271 -953 -225
rect -907 -271 -829 -225
rect -783 -271 -705 -225
rect -659 -271 -581 -225
rect -535 -271 -457 -225
rect -411 -271 -333 -225
rect -287 -271 -209 -225
rect -163 -271 -85 -225
rect -39 -271 39 -225
rect 85 -271 163 -225
rect 209 -271 287 -225
rect 333 -271 411 -225
rect 457 -271 535 -225
rect 581 -271 659 -225
rect 705 -271 783 -225
rect 829 -271 907 -225
rect 953 -271 1031 -225
rect 1077 -271 1155 -225
rect 1201 -271 1279 -225
rect 1325 -271 1403 -225
rect 1449 -271 1527 -225
rect 1573 -271 1651 -225
rect 1697 -271 1775 -225
rect 1821 -271 1899 -225
rect 1945 -271 2023 -225
rect 2069 -271 2147 -225
rect 2193 -271 2271 -225
rect 2317 -271 2395 -225
rect 2441 -271 2519 -225
rect 2565 -271 2643 -225
rect 2689 -271 2767 -225
rect 2813 -271 2891 -225
rect 2937 -271 3015 -225
rect 3061 -271 3139 -225
rect 3185 -271 3263 -225
rect 3309 -271 3387 -225
rect 3433 -271 3511 -225
rect 3557 -271 3635 -225
rect 3681 -271 3759 -225
rect 3805 -271 3883 -225
rect 3929 -271 4007 -225
rect 4053 -271 4131 -225
rect 4177 -271 4255 -225
rect 4301 -271 4379 -225
rect 4425 -271 4503 -225
rect 4549 -271 4627 -225
rect 4673 -271 4751 -225
rect 4797 -271 4875 -225
rect 4921 -271 4999 -225
rect 5045 -271 5123 -225
rect 5169 -271 5247 -225
rect 5293 -271 5371 -225
rect 5417 -271 5495 -225
rect 5541 -271 5619 -225
rect 5665 -271 5743 -225
rect 5789 -271 5800 -225
rect -5800 -349 5800 -271
rect -5800 -395 -5789 -349
rect -5743 -395 -5665 -349
rect -5619 -395 -5541 -349
rect -5495 -395 -5417 -349
rect -5371 -395 -5293 -349
rect -5247 -395 -5169 -349
rect -5123 -395 -5045 -349
rect -4999 -395 -4921 -349
rect -4875 -395 -4797 -349
rect -4751 -395 -4673 -349
rect -4627 -395 -4549 -349
rect -4503 -395 -4425 -349
rect -4379 -395 -4301 -349
rect -4255 -395 -4177 -349
rect -4131 -395 -4053 -349
rect -4007 -395 -3929 -349
rect -3883 -395 -3805 -349
rect -3759 -395 -3681 -349
rect -3635 -395 -3557 -349
rect -3511 -395 -3433 -349
rect -3387 -395 -3309 -349
rect -3263 -395 -3185 -349
rect -3139 -395 -3061 -349
rect -3015 -395 -2937 -349
rect -2891 -395 -2813 -349
rect -2767 -395 -2689 -349
rect -2643 -395 -2565 -349
rect -2519 -395 -2441 -349
rect -2395 -395 -2317 -349
rect -2271 -395 -2193 -349
rect -2147 -395 -2069 -349
rect -2023 -395 -1945 -349
rect -1899 -395 -1821 -349
rect -1775 -395 -1697 -349
rect -1651 -395 -1573 -349
rect -1527 -395 -1449 -349
rect -1403 -395 -1325 -349
rect -1279 -395 -1201 -349
rect -1155 -395 -1077 -349
rect -1031 -395 -953 -349
rect -907 -395 -829 -349
rect -783 -395 -705 -349
rect -659 -395 -581 -349
rect -535 -395 -457 -349
rect -411 -395 -333 -349
rect -287 -395 -209 -349
rect -163 -395 -85 -349
rect -39 -395 39 -349
rect 85 -395 163 -349
rect 209 -395 287 -349
rect 333 -395 411 -349
rect 457 -395 535 -349
rect 581 -395 659 -349
rect 705 -395 783 -349
rect 829 -395 907 -349
rect 953 -395 1031 -349
rect 1077 -395 1155 -349
rect 1201 -395 1279 -349
rect 1325 -395 1403 -349
rect 1449 -395 1527 -349
rect 1573 -395 1651 -349
rect 1697 -395 1775 -349
rect 1821 -395 1899 -349
rect 1945 -395 2023 -349
rect 2069 -395 2147 -349
rect 2193 -395 2271 -349
rect 2317 -395 2395 -349
rect 2441 -395 2519 -349
rect 2565 -395 2643 -349
rect 2689 -395 2767 -349
rect 2813 -395 2891 -349
rect 2937 -395 3015 -349
rect 3061 -395 3139 -349
rect 3185 -395 3263 -349
rect 3309 -395 3387 -349
rect 3433 -395 3511 -349
rect 3557 -395 3635 -349
rect 3681 -395 3759 -349
rect 3805 -395 3883 -349
rect 3929 -395 4007 -349
rect 4053 -395 4131 -349
rect 4177 -395 4255 -349
rect 4301 -395 4379 -349
rect 4425 -395 4503 -349
rect 4549 -395 4627 -349
rect 4673 -395 4751 -349
rect 4797 -395 4875 -349
rect 4921 -395 4999 -349
rect 5045 -395 5123 -349
rect 5169 -395 5247 -349
rect 5293 -395 5371 -349
rect 5417 -395 5495 -349
rect 5541 -395 5619 -349
rect 5665 -395 5743 -349
rect 5789 -395 5800 -349
rect -5800 -473 5800 -395
rect -5800 -519 -5789 -473
rect -5743 -519 -5665 -473
rect -5619 -519 -5541 -473
rect -5495 -519 -5417 -473
rect -5371 -519 -5293 -473
rect -5247 -519 -5169 -473
rect -5123 -519 -5045 -473
rect -4999 -519 -4921 -473
rect -4875 -519 -4797 -473
rect -4751 -519 -4673 -473
rect -4627 -519 -4549 -473
rect -4503 -519 -4425 -473
rect -4379 -519 -4301 -473
rect -4255 -519 -4177 -473
rect -4131 -519 -4053 -473
rect -4007 -519 -3929 -473
rect -3883 -519 -3805 -473
rect -3759 -519 -3681 -473
rect -3635 -519 -3557 -473
rect -3511 -519 -3433 -473
rect -3387 -519 -3309 -473
rect -3263 -519 -3185 -473
rect -3139 -519 -3061 -473
rect -3015 -519 -2937 -473
rect -2891 -519 -2813 -473
rect -2767 -519 -2689 -473
rect -2643 -519 -2565 -473
rect -2519 -519 -2441 -473
rect -2395 -519 -2317 -473
rect -2271 -519 -2193 -473
rect -2147 -519 -2069 -473
rect -2023 -519 -1945 -473
rect -1899 -519 -1821 -473
rect -1775 -519 -1697 -473
rect -1651 -519 -1573 -473
rect -1527 -519 -1449 -473
rect -1403 -519 -1325 -473
rect -1279 -519 -1201 -473
rect -1155 -519 -1077 -473
rect -1031 -519 -953 -473
rect -907 -519 -829 -473
rect -783 -519 -705 -473
rect -659 -519 -581 -473
rect -535 -519 -457 -473
rect -411 -519 -333 -473
rect -287 -519 -209 -473
rect -163 -519 -85 -473
rect -39 -519 39 -473
rect 85 -519 163 -473
rect 209 -519 287 -473
rect 333 -519 411 -473
rect 457 -519 535 -473
rect 581 -519 659 -473
rect 705 -519 783 -473
rect 829 -519 907 -473
rect 953 -519 1031 -473
rect 1077 -519 1155 -473
rect 1201 -519 1279 -473
rect 1325 -519 1403 -473
rect 1449 -519 1527 -473
rect 1573 -519 1651 -473
rect 1697 -519 1775 -473
rect 1821 -519 1899 -473
rect 1945 -519 2023 -473
rect 2069 -519 2147 -473
rect 2193 -519 2271 -473
rect 2317 -519 2395 -473
rect 2441 -519 2519 -473
rect 2565 -519 2643 -473
rect 2689 -519 2767 -473
rect 2813 -519 2891 -473
rect 2937 -519 3015 -473
rect 3061 -519 3139 -473
rect 3185 -519 3263 -473
rect 3309 -519 3387 -473
rect 3433 -519 3511 -473
rect 3557 -519 3635 -473
rect 3681 -519 3759 -473
rect 3805 -519 3883 -473
rect 3929 -519 4007 -473
rect 4053 -519 4131 -473
rect 4177 -519 4255 -473
rect 4301 -519 4379 -473
rect 4425 -519 4503 -473
rect 4549 -519 4627 -473
rect 4673 -519 4751 -473
rect 4797 -519 4875 -473
rect 4921 -519 4999 -473
rect 5045 -519 5123 -473
rect 5169 -519 5247 -473
rect 5293 -519 5371 -473
rect 5417 -519 5495 -473
rect 5541 -519 5619 -473
rect 5665 -519 5743 -473
rect 5789 -519 5800 -473
rect -5800 -597 5800 -519
rect -5800 -643 -5789 -597
rect -5743 -643 -5665 -597
rect -5619 -643 -5541 -597
rect -5495 -643 -5417 -597
rect -5371 -643 -5293 -597
rect -5247 -643 -5169 -597
rect -5123 -643 -5045 -597
rect -4999 -643 -4921 -597
rect -4875 -643 -4797 -597
rect -4751 -643 -4673 -597
rect -4627 -643 -4549 -597
rect -4503 -643 -4425 -597
rect -4379 -643 -4301 -597
rect -4255 -643 -4177 -597
rect -4131 -643 -4053 -597
rect -4007 -643 -3929 -597
rect -3883 -643 -3805 -597
rect -3759 -643 -3681 -597
rect -3635 -643 -3557 -597
rect -3511 -643 -3433 -597
rect -3387 -643 -3309 -597
rect -3263 -643 -3185 -597
rect -3139 -643 -3061 -597
rect -3015 -643 -2937 -597
rect -2891 -643 -2813 -597
rect -2767 -643 -2689 -597
rect -2643 -643 -2565 -597
rect -2519 -643 -2441 -597
rect -2395 -643 -2317 -597
rect -2271 -643 -2193 -597
rect -2147 -643 -2069 -597
rect -2023 -643 -1945 -597
rect -1899 -643 -1821 -597
rect -1775 -643 -1697 -597
rect -1651 -643 -1573 -597
rect -1527 -643 -1449 -597
rect -1403 -643 -1325 -597
rect -1279 -643 -1201 -597
rect -1155 -643 -1077 -597
rect -1031 -643 -953 -597
rect -907 -643 -829 -597
rect -783 -643 -705 -597
rect -659 -643 -581 -597
rect -535 -643 -457 -597
rect -411 -643 -333 -597
rect -287 -643 -209 -597
rect -163 -643 -85 -597
rect -39 -643 39 -597
rect 85 -643 163 -597
rect 209 -643 287 -597
rect 333 -643 411 -597
rect 457 -643 535 -597
rect 581 -643 659 -597
rect 705 -643 783 -597
rect 829 -643 907 -597
rect 953 -643 1031 -597
rect 1077 -643 1155 -597
rect 1201 -643 1279 -597
rect 1325 -643 1403 -597
rect 1449 -643 1527 -597
rect 1573 -643 1651 -597
rect 1697 -643 1775 -597
rect 1821 -643 1899 -597
rect 1945 -643 2023 -597
rect 2069 -643 2147 -597
rect 2193 -643 2271 -597
rect 2317 -643 2395 -597
rect 2441 -643 2519 -597
rect 2565 -643 2643 -597
rect 2689 -643 2767 -597
rect 2813 -643 2891 -597
rect 2937 -643 3015 -597
rect 3061 -643 3139 -597
rect 3185 -643 3263 -597
rect 3309 -643 3387 -597
rect 3433 -643 3511 -597
rect 3557 -643 3635 -597
rect 3681 -643 3759 -597
rect 3805 -643 3883 -597
rect 3929 -643 4007 -597
rect 4053 -643 4131 -597
rect 4177 -643 4255 -597
rect 4301 -643 4379 -597
rect 4425 -643 4503 -597
rect 4549 -643 4627 -597
rect 4673 -643 4751 -597
rect 4797 -643 4875 -597
rect 4921 -643 4999 -597
rect 5045 -643 5123 -597
rect 5169 -643 5247 -597
rect 5293 -643 5371 -597
rect 5417 -643 5495 -597
rect 5541 -643 5619 -597
rect 5665 -643 5743 -597
rect 5789 -643 5800 -597
rect -5800 -721 5800 -643
rect -5800 -767 -5789 -721
rect -5743 -767 -5665 -721
rect -5619 -767 -5541 -721
rect -5495 -767 -5417 -721
rect -5371 -767 -5293 -721
rect -5247 -767 -5169 -721
rect -5123 -767 -5045 -721
rect -4999 -767 -4921 -721
rect -4875 -767 -4797 -721
rect -4751 -767 -4673 -721
rect -4627 -767 -4549 -721
rect -4503 -767 -4425 -721
rect -4379 -767 -4301 -721
rect -4255 -767 -4177 -721
rect -4131 -767 -4053 -721
rect -4007 -767 -3929 -721
rect -3883 -767 -3805 -721
rect -3759 -767 -3681 -721
rect -3635 -767 -3557 -721
rect -3511 -767 -3433 -721
rect -3387 -767 -3309 -721
rect -3263 -767 -3185 -721
rect -3139 -767 -3061 -721
rect -3015 -767 -2937 -721
rect -2891 -767 -2813 -721
rect -2767 -767 -2689 -721
rect -2643 -767 -2565 -721
rect -2519 -767 -2441 -721
rect -2395 -767 -2317 -721
rect -2271 -767 -2193 -721
rect -2147 -767 -2069 -721
rect -2023 -767 -1945 -721
rect -1899 -767 -1821 -721
rect -1775 -767 -1697 -721
rect -1651 -767 -1573 -721
rect -1527 -767 -1449 -721
rect -1403 -767 -1325 -721
rect -1279 -767 -1201 -721
rect -1155 -767 -1077 -721
rect -1031 -767 -953 -721
rect -907 -767 -829 -721
rect -783 -767 -705 -721
rect -659 -767 -581 -721
rect -535 -767 -457 -721
rect -411 -767 -333 -721
rect -287 -767 -209 -721
rect -163 -767 -85 -721
rect -39 -767 39 -721
rect 85 -767 163 -721
rect 209 -767 287 -721
rect 333 -767 411 -721
rect 457 -767 535 -721
rect 581 -767 659 -721
rect 705 -767 783 -721
rect 829 -767 907 -721
rect 953 -767 1031 -721
rect 1077 -767 1155 -721
rect 1201 -767 1279 -721
rect 1325 -767 1403 -721
rect 1449 -767 1527 -721
rect 1573 -767 1651 -721
rect 1697 -767 1775 -721
rect 1821 -767 1899 -721
rect 1945 -767 2023 -721
rect 2069 -767 2147 -721
rect 2193 -767 2271 -721
rect 2317 -767 2395 -721
rect 2441 -767 2519 -721
rect 2565 -767 2643 -721
rect 2689 -767 2767 -721
rect 2813 -767 2891 -721
rect 2937 -767 3015 -721
rect 3061 -767 3139 -721
rect 3185 -767 3263 -721
rect 3309 -767 3387 -721
rect 3433 -767 3511 -721
rect 3557 -767 3635 -721
rect 3681 -767 3759 -721
rect 3805 -767 3883 -721
rect 3929 -767 4007 -721
rect 4053 -767 4131 -721
rect 4177 -767 4255 -721
rect 4301 -767 4379 -721
rect 4425 -767 4503 -721
rect 4549 -767 4627 -721
rect 4673 -767 4751 -721
rect 4797 -767 4875 -721
rect 4921 -767 4999 -721
rect 5045 -767 5123 -721
rect 5169 -767 5247 -721
rect 5293 -767 5371 -721
rect 5417 -767 5495 -721
rect 5541 -767 5619 -721
rect 5665 -767 5743 -721
rect 5789 -767 5800 -721
rect -5800 -845 5800 -767
rect -5800 -891 -5789 -845
rect -5743 -891 -5665 -845
rect -5619 -891 -5541 -845
rect -5495 -891 -5417 -845
rect -5371 -891 -5293 -845
rect -5247 -891 -5169 -845
rect -5123 -891 -5045 -845
rect -4999 -891 -4921 -845
rect -4875 -891 -4797 -845
rect -4751 -891 -4673 -845
rect -4627 -891 -4549 -845
rect -4503 -891 -4425 -845
rect -4379 -891 -4301 -845
rect -4255 -891 -4177 -845
rect -4131 -891 -4053 -845
rect -4007 -891 -3929 -845
rect -3883 -891 -3805 -845
rect -3759 -891 -3681 -845
rect -3635 -891 -3557 -845
rect -3511 -891 -3433 -845
rect -3387 -891 -3309 -845
rect -3263 -891 -3185 -845
rect -3139 -891 -3061 -845
rect -3015 -891 -2937 -845
rect -2891 -891 -2813 -845
rect -2767 -891 -2689 -845
rect -2643 -891 -2565 -845
rect -2519 -891 -2441 -845
rect -2395 -891 -2317 -845
rect -2271 -891 -2193 -845
rect -2147 -891 -2069 -845
rect -2023 -891 -1945 -845
rect -1899 -891 -1821 -845
rect -1775 -891 -1697 -845
rect -1651 -891 -1573 -845
rect -1527 -891 -1449 -845
rect -1403 -891 -1325 -845
rect -1279 -891 -1201 -845
rect -1155 -891 -1077 -845
rect -1031 -891 -953 -845
rect -907 -891 -829 -845
rect -783 -891 -705 -845
rect -659 -891 -581 -845
rect -535 -891 -457 -845
rect -411 -891 -333 -845
rect -287 -891 -209 -845
rect -163 -891 -85 -845
rect -39 -891 39 -845
rect 85 -891 163 -845
rect 209 -891 287 -845
rect 333 -891 411 -845
rect 457 -891 535 -845
rect 581 -891 659 -845
rect 705 -891 783 -845
rect 829 -891 907 -845
rect 953 -891 1031 -845
rect 1077 -891 1155 -845
rect 1201 -891 1279 -845
rect 1325 -891 1403 -845
rect 1449 -891 1527 -845
rect 1573 -891 1651 -845
rect 1697 -891 1775 -845
rect 1821 -891 1899 -845
rect 1945 -891 2023 -845
rect 2069 -891 2147 -845
rect 2193 -891 2271 -845
rect 2317 -891 2395 -845
rect 2441 -891 2519 -845
rect 2565 -891 2643 -845
rect 2689 -891 2767 -845
rect 2813 -891 2891 -845
rect 2937 -891 3015 -845
rect 3061 -891 3139 -845
rect 3185 -891 3263 -845
rect 3309 -891 3387 -845
rect 3433 -891 3511 -845
rect 3557 -891 3635 -845
rect 3681 -891 3759 -845
rect 3805 -891 3883 -845
rect 3929 -891 4007 -845
rect 4053 -891 4131 -845
rect 4177 -891 4255 -845
rect 4301 -891 4379 -845
rect 4425 -891 4503 -845
rect 4549 -891 4627 -845
rect 4673 -891 4751 -845
rect 4797 -891 4875 -845
rect 4921 -891 4999 -845
rect 5045 -891 5123 -845
rect 5169 -891 5247 -845
rect 5293 -891 5371 -845
rect 5417 -891 5495 -845
rect 5541 -891 5619 -845
rect 5665 -891 5743 -845
rect 5789 -891 5800 -845
rect -5800 -969 5800 -891
rect -5800 -1015 -5789 -969
rect -5743 -1015 -5665 -969
rect -5619 -1015 -5541 -969
rect -5495 -1015 -5417 -969
rect -5371 -1015 -5293 -969
rect -5247 -1015 -5169 -969
rect -5123 -1015 -5045 -969
rect -4999 -1015 -4921 -969
rect -4875 -1015 -4797 -969
rect -4751 -1015 -4673 -969
rect -4627 -1015 -4549 -969
rect -4503 -1015 -4425 -969
rect -4379 -1015 -4301 -969
rect -4255 -1015 -4177 -969
rect -4131 -1015 -4053 -969
rect -4007 -1015 -3929 -969
rect -3883 -1015 -3805 -969
rect -3759 -1015 -3681 -969
rect -3635 -1015 -3557 -969
rect -3511 -1015 -3433 -969
rect -3387 -1015 -3309 -969
rect -3263 -1015 -3185 -969
rect -3139 -1015 -3061 -969
rect -3015 -1015 -2937 -969
rect -2891 -1015 -2813 -969
rect -2767 -1015 -2689 -969
rect -2643 -1015 -2565 -969
rect -2519 -1015 -2441 -969
rect -2395 -1015 -2317 -969
rect -2271 -1015 -2193 -969
rect -2147 -1015 -2069 -969
rect -2023 -1015 -1945 -969
rect -1899 -1015 -1821 -969
rect -1775 -1015 -1697 -969
rect -1651 -1015 -1573 -969
rect -1527 -1015 -1449 -969
rect -1403 -1015 -1325 -969
rect -1279 -1015 -1201 -969
rect -1155 -1015 -1077 -969
rect -1031 -1015 -953 -969
rect -907 -1015 -829 -969
rect -783 -1015 -705 -969
rect -659 -1015 -581 -969
rect -535 -1015 -457 -969
rect -411 -1015 -333 -969
rect -287 -1015 -209 -969
rect -163 -1015 -85 -969
rect -39 -1015 39 -969
rect 85 -1015 163 -969
rect 209 -1015 287 -969
rect 333 -1015 411 -969
rect 457 -1015 535 -969
rect 581 -1015 659 -969
rect 705 -1015 783 -969
rect 829 -1015 907 -969
rect 953 -1015 1031 -969
rect 1077 -1015 1155 -969
rect 1201 -1015 1279 -969
rect 1325 -1015 1403 -969
rect 1449 -1015 1527 -969
rect 1573 -1015 1651 -969
rect 1697 -1015 1775 -969
rect 1821 -1015 1899 -969
rect 1945 -1015 2023 -969
rect 2069 -1015 2147 -969
rect 2193 -1015 2271 -969
rect 2317 -1015 2395 -969
rect 2441 -1015 2519 -969
rect 2565 -1015 2643 -969
rect 2689 -1015 2767 -969
rect 2813 -1015 2891 -969
rect 2937 -1015 3015 -969
rect 3061 -1015 3139 -969
rect 3185 -1015 3263 -969
rect 3309 -1015 3387 -969
rect 3433 -1015 3511 -969
rect 3557 -1015 3635 -969
rect 3681 -1015 3759 -969
rect 3805 -1015 3883 -969
rect 3929 -1015 4007 -969
rect 4053 -1015 4131 -969
rect 4177 -1015 4255 -969
rect 4301 -1015 4379 -969
rect 4425 -1015 4503 -969
rect 4549 -1015 4627 -969
rect 4673 -1015 4751 -969
rect 4797 -1015 4875 -969
rect 4921 -1015 4999 -969
rect 5045 -1015 5123 -969
rect 5169 -1015 5247 -969
rect 5293 -1015 5371 -969
rect 5417 -1015 5495 -969
rect 5541 -1015 5619 -969
rect 5665 -1015 5743 -969
rect 5789 -1015 5800 -969
rect -5800 -1093 5800 -1015
rect -5800 -1139 -5789 -1093
rect -5743 -1139 -5665 -1093
rect -5619 -1139 -5541 -1093
rect -5495 -1139 -5417 -1093
rect -5371 -1139 -5293 -1093
rect -5247 -1139 -5169 -1093
rect -5123 -1139 -5045 -1093
rect -4999 -1139 -4921 -1093
rect -4875 -1139 -4797 -1093
rect -4751 -1139 -4673 -1093
rect -4627 -1139 -4549 -1093
rect -4503 -1139 -4425 -1093
rect -4379 -1139 -4301 -1093
rect -4255 -1139 -4177 -1093
rect -4131 -1139 -4053 -1093
rect -4007 -1139 -3929 -1093
rect -3883 -1139 -3805 -1093
rect -3759 -1139 -3681 -1093
rect -3635 -1139 -3557 -1093
rect -3511 -1139 -3433 -1093
rect -3387 -1139 -3309 -1093
rect -3263 -1139 -3185 -1093
rect -3139 -1139 -3061 -1093
rect -3015 -1139 -2937 -1093
rect -2891 -1139 -2813 -1093
rect -2767 -1139 -2689 -1093
rect -2643 -1139 -2565 -1093
rect -2519 -1139 -2441 -1093
rect -2395 -1139 -2317 -1093
rect -2271 -1139 -2193 -1093
rect -2147 -1139 -2069 -1093
rect -2023 -1139 -1945 -1093
rect -1899 -1139 -1821 -1093
rect -1775 -1139 -1697 -1093
rect -1651 -1139 -1573 -1093
rect -1527 -1139 -1449 -1093
rect -1403 -1139 -1325 -1093
rect -1279 -1139 -1201 -1093
rect -1155 -1139 -1077 -1093
rect -1031 -1139 -953 -1093
rect -907 -1139 -829 -1093
rect -783 -1139 -705 -1093
rect -659 -1139 -581 -1093
rect -535 -1139 -457 -1093
rect -411 -1139 -333 -1093
rect -287 -1139 -209 -1093
rect -163 -1139 -85 -1093
rect -39 -1139 39 -1093
rect 85 -1139 163 -1093
rect 209 -1139 287 -1093
rect 333 -1139 411 -1093
rect 457 -1139 535 -1093
rect 581 -1139 659 -1093
rect 705 -1139 783 -1093
rect 829 -1139 907 -1093
rect 953 -1139 1031 -1093
rect 1077 -1139 1155 -1093
rect 1201 -1139 1279 -1093
rect 1325 -1139 1403 -1093
rect 1449 -1139 1527 -1093
rect 1573 -1139 1651 -1093
rect 1697 -1139 1775 -1093
rect 1821 -1139 1899 -1093
rect 1945 -1139 2023 -1093
rect 2069 -1139 2147 -1093
rect 2193 -1139 2271 -1093
rect 2317 -1139 2395 -1093
rect 2441 -1139 2519 -1093
rect 2565 -1139 2643 -1093
rect 2689 -1139 2767 -1093
rect 2813 -1139 2891 -1093
rect 2937 -1139 3015 -1093
rect 3061 -1139 3139 -1093
rect 3185 -1139 3263 -1093
rect 3309 -1139 3387 -1093
rect 3433 -1139 3511 -1093
rect 3557 -1139 3635 -1093
rect 3681 -1139 3759 -1093
rect 3805 -1139 3883 -1093
rect 3929 -1139 4007 -1093
rect 4053 -1139 4131 -1093
rect 4177 -1139 4255 -1093
rect 4301 -1139 4379 -1093
rect 4425 -1139 4503 -1093
rect 4549 -1139 4627 -1093
rect 4673 -1139 4751 -1093
rect 4797 -1139 4875 -1093
rect 4921 -1139 4999 -1093
rect 5045 -1139 5123 -1093
rect 5169 -1139 5247 -1093
rect 5293 -1139 5371 -1093
rect 5417 -1139 5495 -1093
rect 5541 -1139 5619 -1093
rect 5665 -1139 5743 -1093
rect 5789 -1139 5800 -1093
rect -5800 -1217 5800 -1139
rect -5800 -1263 -5789 -1217
rect -5743 -1263 -5665 -1217
rect -5619 -1263 -5541 -1217
rect -5495 -1263 -5417 -1217
rect -5371 -1263 -5293 -1217
rect -5247 -1263 -5169 -1217
rect -5123 -1263 -5045 -1217
rect -4999 -1263 -4921 -1217
rect -4875 -1263 -4797 -1217
rect -4751 -1263 -4673 -1217
rect -4627 -1263 -4549 -1217
rect -4503 -1263 -4425 -1217
rect -4379 -1263 -4301 -1217
rect -4255 -1263 -4177 -1217
rect -4131 -1263 -4053 -1217
rect -4007 -1263 -3929 -1217
rect -3883 -1263 -3805 -1217
rect -3759 -1263 -3681 -1217
rect -3635 -1263 -3557 -1217
rect -3511 -1263 -3433 -1217
rect -3387 -1263 -3309 -1217
rect -3263 -1263 -3185 -1217
rect -3139 -1263 -3061 -1217
rect -3015 -1263 -2937 -1217
rect -2891 -1263 -2813 -1217
rect -2767 -1263 -2689 -1217
rect -2643 -1263 -2565 -1217
rect -2519 -1263 -2441 -1217
rect -2395 -1263 -2317 -1217
rect -2271 -1263 -2193 -1217
rect -2147 -1263 -2069 -1217
rect -2023 -1263 -1945 -1217
rect -1899 -1263 -1821 -1217
rect -1775 -1263 -1697 -1217
rect -1651 -1263 -1573 -1217
rect -1527 -1263 -1449 -1217
rect -1403 -1263 -1325 -1217
rect -1279 -1263 -1201 -1217
rect -1155 -1263 -1077 -1217
rect -1031 -1263 -953 -1217
rect -907 -1263 -829 -1217
rect -783 -1263 -705 -1217
rect -659 -1263 -581 -1217
rect -535 -1263 -457 -1217
rect -411 -1263 -333 -1217
rect -287 -1263 -209 -1217
rect -163 -1263 -85 -1217
rect -39 -1263 39 -1217
rect 85 -1263 163 -1217
rect 209 -1263 287 -1217
rect 333 -1263 411 -1217
rect 457 -1263 535 -1217
rect 581 -1263 659 -1217
rect 705 -1263 783 -1217
rect 829 -1263 907 -1217
rect 953 -1263 1031 -1217
rect 1077 -1263 1155 -1217
rect 1201 -1263 1279 -1217
rect 1325 -1263 1403 -1217
rect 1449 -1263 1527 -1217
rect 1573 -1263 1651 -1217
rect 1697 -1263 1775 -1217
rect 1821 -1263 1899 -1217
rect 1945 -1263 2023 -1217
rect 2069 -1263 2147 -1217
rect 2193 -1263 2271 -1217
rect 2317 -1263 2395 -1217
rect 2441 -1263 2519 -1217
rect 2565 -1263 2643 -1217
rect 2689 -1263 2767 -1217
rect 2813 -1263 2891 -1217
rect 2937 -1263 3015 -1217
rect 3061 -1263 3139 -1217
rect 3185 -1263 3263 -1217
rect 3309 -1263 3387 -1217
rect 3433 -1263 3511 -1217
rect 3557 -1263 3635 -1217
rect 3681 -1263 3759 -1217
rect 3805 -1263 3883 -1217
rect 3929 -1263 4007 -1217
rect 4053 -1263 4131 -1217
rect 4177 -1263 4255 -1217
rect 4301 -1263 4379 -1217
rect 4425 -1263 4503 -1217
rect 4549 -1263 4627 -1217
rect 4673 -1263 4751 -1217
rect 4797 -1263 4875 -1217
rect 4921 -1263 4999 -1217
rect 5045 -1263 5123 -1217
rect 5169 -1263 5247 -1217
rect 5293 -1263 5371 -1217
rect 5417 -1263 5495 -1217
rect 5541 -1263 5619 -1217
rect 5665 -1263 5743 -1217
rect 5789 -1263 5800 -1217
rect -5800 -1274 5800 -1263
<< end >>
