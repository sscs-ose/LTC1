magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -3778 -1081 3778 1081
<< metal1 >>
rect -2778 75 2778 81
rect -2778 49 -2772 75
rect -2746 49 -2710 75
rect -2684 49 -2648 75
rect -2622 49 -2586 75
rect -2560 49 -2524 75
rect -2498 49 -2462 75
rect -2436 49 -2400 75
rect -2374 49 -2338 75
rect -2312 49 -2276 75
rect -2250 49 -2214 75
rect -2188 49 -2152 75
rect -2126 49 -2090 75
rect -2064 49 -2028 75
rect -2002 49 -1966 75
rect -1940 49 -1904 75
rect -1878 49 -1842 75
rect -1816 49 -1780 75
rect -1754 49 -1718 75
rect -1692 49 -1656 75
rect -1630 49 -1594 75
rect -1568 49 -1532 75
rect -1506 49 -1470 75
rect -1444 49 -1408 75
rect -1382 49 -1346 75
rect -1320 49 -1284 75
rect -1258 49 -1222 75
rect -1196 49 -1160 75
rect -1134 49 -1098 75
rect -1072 49 -1036 75
rect -1010 49 -974 75
rect -948 49 -912 75
rect -886 49 -850 75
rect -824 49 -788 75
rect -762 49 -726 75
rect -700 49 -664 75
rect -638 49 -602 75
rect -576 49 -540 75
rect -514 49 -478 75
rect -452 49 -416 75
rect -390 49 -354 75
rect -328 49 -292 75
rect -266 49 -230 75
rect -204 49 -168 75
rect -142 49 -106 75
rect -80 49 -44 75
rect -18 49 18 75
rect 44 49 80 75
rect 106 49 142 75
rect 168 49 204 75
rect 230 49 266 75
rect 292 49 328 75
rect 354 49 390 75
rect 416 49 452 75
rect 478 49 514 75
rect 540 49 576 75
rect 602 49 638 75
rect 664 49 700 75
rect 726 49 762 75
rect 788 49 824 75
rect 850 49 886 75
rect 912 49 948 75
rect 974 49 1010 75
rect 1036 49 1072 75
rect 1098 49 1134 75
rect 1160 49 1196 75
rect 1222 49 1258 75
rect 1284 49 1320 75
rect 1346 49 1382 75
rect 1408 49 1444 75
rect 1470 49 1506 75
rect 1532 49 1568 75
rect 1594 49 1630 75
rect 1656 49 1692 75
rect 1718 49 1754 75
rect 1780 49 1816 75
rect 1842 49 1878 75
rect 1904 49 1940 75
rect 1966 49 2002 75
rect 2028 49 2064 75
rect 2090 49 2126 75
rect 2152 49 2188 75
rect 2214 49 2250 75
rect 2276 49 2312 75
rect 2338 49 2374 75
rect 2400 49 2436 75
rect 2462 49 2498 75
rect 2524 49 2560 75
rect 2586 49 2622 75
rect 2648 49 2684 75
rect 2710 49 2746 75
rect 2772 49 2778 75
rect -2778 13 2778 49
rect -2778 -13 -2772 13
rect -2746 -13 -2710 13
rect -2684 -13 -2648 13
rect -2622 -13 -2586 13
rect -2560 -13 -2524 13
rect -2498 -13 -2462 13
rect -2436 -13 -2400 13
rect -2374 -13 -2338 13
rect -2312 -13 -2276 13
rect -2250 -13 -2214 13
rect -2188 -13 -2152 13
rect -2126 -13 -2090 13
rect -2064 -13 -2028 13
rect -2002 -13 -1966 13
rect -1940 -13 -1904 13
rect -1878 -13 -1842 13
rect -1816 -13 -1780 13
rect -1754 -13 -1718 13
rect -1692 -13 -1656 13
rect -1630 -13 -1594 13
rect -1568 -13 -1532 13
rect -1506 -13 -1470 13
rect -1444 -13 -1408 13
rect -1382 -13 -1346 13
rect -1320 -13 -1284 13
rect -1258 -13 -1222 13
rect -1196 -13 -1160 13
rect -1134 -13 -1098 13
rect -1072 -13 -1036 13
rect -1010 -13 -974 13
rect -948 -13 -912 13
rect -886 -13 -850 13
rect -824 -13 -788 13
rect -762 -13 -726 13
rect -700 -13 -664 13
rect -638 -13 -602 13
rect -576 -13 -540 13
rect -514 -13 -478 13
rect -452 -13 -416 13
rect -390 -13 -354 13
rect -328 -13 -292 13
rect -266 -13 -230 13
rect -204 -13 -168 13
rect -142 -13 -106 13
rect -80 -13 -44 13
rect -18 -13 18 13
rect 44 -13 80 13
rect 106 -13 142 13
rect 168 -13 204 13
rect 230 -13 266 13
rect 292 -13 328 13
rect 354 -13 390 13
rect 416 -13 452 13
rect 478 -13 514 13
rect 540 -13 576 13
rect 602 -13 638 13
rect 664 -13 700 13
rect 726 -13 762 13
rect 788 -13 824 13
rect 850 -13 886 13
rect 912 -13 948 13
rect 974 -13 1010 13
rect 1036 -13 1072 13
rect 1098 -13 1134 13
rect 1160 -13 1196 13
rect 1222 -13 1258 13
rect 1284 -13 1320 13
rect 1346 -13 1382 13
rect 1408 -13 1444 13
rect 1470 -13 1506 13
rect 1532 -13 1568 13
rect 1594 -13 1630 13
rect 1656 -13 1692 13
rect 1718 -13 1754 13
rect 1780 -13 1816 13
rect 1842 -13 1878 13
rect 1904 -13 1940 13
rect 1966 -13 2002 13
rect 2028 -13 2064 13
rect 2090 -13 2126 13
rect 2152 -13 2188 13
rect 2214 -13 2250 13
rect 2276 -13 2312 13
rect 2338 -13 2374 13
rect 2400 -13 2436 13
rect 2462 -13 2498 13
rect 2524 -13 2560 13
rect 2586 -13 2622 13
rect 2648 -13 2684 13
rect 2710 -13 2746 13
rect 2772 -13 2778 13
rect -2778 -49 2778 -13
rect -2778 -75 -2772 -49
rect -2746 -75 -2710 -49
rect -2684 -75 -2648 -49
rect -2622 -75 -2586 -49
rect -2560 -75 -2524 -49
rect -2498 -75 -2462 -49
rect -2436 -75 -2400 -49
rect -2374 -75 -2338 -49
rect -2312 -75 -2276 -49
rect -2250 -75 -2214 -49
rect -2188 -75 -2152 -49
rect -2126 -75 -2090 -49
rect -2064 -75 -2028 -49
rect -2002 -75 -1966 -49
rect -1940 -75 -1904 -49
rect -1878 -75 -1842 -49
rect -1816 -75 -1780 -49
rect -1754 -75 -1718 -49
rect -1692 -75 -1656 -49
rect -1630 -75 -1594 -49
rect -1568 -75 -1532 -49
rect -1506 -75 -1470 -49
rect -1444 -75 -1408 -49
rect -1382 -75 -1346 -49
rect -1320 -75 -1284 -49
rect -1258 -75 -1222 -49
rect -1196 -75 -1160 -49
rect -1134 -75 -1098 -49
rect -1072 -75 -1036 -49
rect -1010 -75 -974 -49
rect -948 -75 -912 -49
rect -886 -75 -850 -49
rect -824 -75 -788 -49
rect -762 -75 -726 -49
rect -700 -75 -664 -49
rect -638 -75 -602 -49
rect -576 -75 -540 -49
rect -514 -75 -478 -49
rect -452 -75 -416 -49
rect -390 -75 -354 -49
rect -328 -75 -292 -49
rect -266 -75 -230 -49
rect -204 -75 -168 -49
rect -142 -75 -106 -49
rect -80 -75 -44 -49
rect -18 -75 18 -49
rect 44 -75 80 -49
rect 106 -75 142 -49
rect 168 -75 204 -49
rect 230 -75 266 -49
rect 292 -75 328 -49
rect 354 -75 390 -49
rect 416 -75 452 -49
rect 478 -75 514 -49
rect 540 -75 576 -49
rect 602 -75 638 -49
rect 664 -75 700 -49
rect 726 -75 762 -49
rect 788 -75 824 -49
rect 850 -75 886 -49
rect 912 -75 948 -49
rect 974 -75 1010 -49
rect 1036 -75 1072 -49
rect 1098 -75 1134 -49
rect 1160 -75 1196 -49
rect 1222 -75 1258 -49
rect 1284 -75 1320 -49
rect 1346 -75 1382 -49
rect 1408 -75 1444 -49
rect 1470 -75 1506 -49
rect 1532 -75 1568 -49
rect 1594 -75 1630 -49
rect 1656 -75 1692 -49
rect 1718 -75 1754 -49
rect 1780 -75 1816 -49
rect 1842 -75 1878 -49
rect 1904 -75 1940 -49
rect 1966 -75 2002 -49
rect 2028 -75 2064 -49
rect 2090 -75 2126 -49
rect 2152 -75 2188 -49
rect 2214 -75 2250 -49
rect 2276 -75 2312 -49
rect 2338 -75 2374 -49
rect 2400 -75 2436 -49
rect 2462 -75 2498 -49
rect 2524 -75 2560 -49
rect 2586 -75 2622 -49
rect 2648 -75 2684 -49
rect 2710 -75 2746 -49
rect 2772 -75 2778 -49
rect -2778 -81 2778 -75
<< via1 >>
rect -2772 49 -2746 75
rect -2710 49 -2684 75
rect -2648 49 -2622 75
rect -2586 49 -2560 75
rect -2524 49 -2498 75
rect -2462 49 -2436 75
rect -2400 49 -2374 75
rect -2338 49 -2312 75
rect -2276 49 -2250 75
rect -2214 49 -2188 75
rect -2152 49 -2126 75
rect -2090 49 -2064 75
rect -2028 49 -2002 75
rect -1966 49 -1940 75
rect -1904 49 -1878 75
rect -1842 49 -1816 75
rect -1780 49 -1754 75
rect -1718 49 -1692 75
rect -1656 49 -1630 75
rect -1594 49 -1568 75
rect -1532 49 -1506 75
rect -1470 49 -1444 75
rect -1408 49 -1382 75
rect -1346 49 -1320 75
rect -1284 49 -1258 75
rect -1222 49 -1196 75
rect -1160 49 -1134 75
rect -1098 49 -1072 75
rect -1036 49 -1010 75
rect -974 49 -948 75
rect -912 49 -886 75
rect -850 49 -824 75
rect -788 49 -762 75
rect -726 49 -700 75
rect -664 49 -638 75
rect -602 49 -576 75
rect -540 49 -514 75
rect -478 49 -452 75
rect -416 49 -390 75
rect -354 49 -328 75
rect -292 49 -266 75
rect -230 49 -204 75
rect -168 49 -142 75
rect -106 49 -80 75
rect -44 49 -18 75
rect 18 49 44 75
rect 80 49 106 75
rect 142 49 168 75
rect 204 49 230 75
rect 266 49 292 75
rect 328 49 354 75
rect 390 49 416 75
rect 452 49 478 75
rect 514 49 540 75
rect 576 49 602 75
rect 638 49 664 75
rect 700 49 726 75
rect 762 49 788 75
rect 824 49 850 75
rect 886 49 912 75
rect 948 49 974 75
rect 1010 49 1036 75
rect 1072 49 1098 75
rect 1134 49 1160 75
rect 1196 49 1222 75
rect 1258 49 1284 75
rect 1320 49 1346 75
rect 1382 49 1408 75
rect 1444 49 1470 75
rect 1506 49 1532 75
rect 1568 49 1594 75
rect 1630 49 1656 75
rect 1692 49 1718 75
rect 1754 49 1780 75
rect 1816 49 1842 75
rect 1878 49 1904 75
rect 1940 49 1966 75
rect 2002 49 2028 75
rect 2064 49 2090 75
rect 2126 49 2152 75
rect 2188 49 2214 75
rect 2250 49 2276 75
rect 2312 49 2338 75
rect 2374 49 2400 75
rect 2436 49 2462 75
rect 2498 49 2524 75
rect 2560 49 2586 75
rect 2622 49 2648 75
rect 2684 49 2710 75
rect 2746 49 2772 75
rect -2772 -13 -2746 13
rect -2710 -13 -2684 13
rect -2648 -13 -2622 13
rect -2586 -13 -2560 13
rect -2524 -13 -2498 13
rect -2462 -13 -2436 13
rect -2400 -13 -2374 13
rect -2338 -13 -2312 13
rect -2276 -13 -2250 13
rect -2214 -13 -2188 13
rect -2152 -13 -2126 13
rect -2090 -13 -2064 13
rect -2028 -13 -2002 13
rect -1966 -13 -1940 13
rect -1904 -13 -1878 13
rect -1842 -13 -1816 13
rect -1780 -13 -1754 13
rect -1718 -13 -1692 13
rect -1656 -13 -1630 13
rect -1594 -13 -1568 13
rect -1532 -13 -1506 13
rect -1470 -13 -1444 13
rect -1408 -13 -1382 13
rect -1346 -13 -1320 13
rect -1284 -13 -1258 13
rect -1222 -13 -1196 13
rect -1160 -13 -1134 13
rect -1098 -13 -1072 13
rect -1036 -13 -1010 13
rect -974 -13 -948 13
rect -912 -13 -886 13
rect -850 -13 -824 13
rect -788 -13 -762 13
rect -726 -13 -700 13
rect -664 -13 -638 13
rect -602 -13 -576 13
rect -540 -13 -514 13
rect -478 -13 -452 13
rect -416 -13 -390 13
rect -354 -13 -328 13
rect -292 -13 -266 13
rect -230 -13 -204 13
rect -168 -13 -142 13
rect -106 -13 -80 13
rect -44 -13 -18 13
rect 18 -13 44 13
rect 80 -13 106 13
rect 142 -13 168 13
rect 204 -13 230 13
rect 266 -13 292 13
rect 328 -13 354 13
rect 390 -13 416 13
rect 452 -13 478 13
rect 514 -13 540 13
rect 576 -13 602 13
rect 638 -13 664 13
rect 700 -13 726 13
rect 762 -13 788 13
rect 824 -13 850 13
rect 886 -13 912 13
rect 948 -13 974 13
rect 1010 -13 1036 13
rect 1072 -13 1098 13
rect 1134 -13 1160 13
rect 1196 -13 1222 13
rect 1258 -13 1284 13
rect 1320 -13 1346 13
rect 1382 -13 1408 13
rect 1444 -13 1470 13
rect 1506 -13 1532 13
rect 1568 -13 1594 13
rect 1630 -13 1656 13
rect 1692 -13 1718 13
rect 1754 -13 1780 13
rect 1816 -13 1842 13
rect 1878 -13 1904 13
rect 1940 -13 1966 13
rect 2002 -13 2028 13
rect 2064 -13 2090 13
rect 2126 -13 2152 13
rect 2188 -13 2214 13
rect 2250 -13 2276 13
rect 2312 -13 2338 13
rect 2374 -13 2400 13
rect 2436 -13 2462 13
rect 2498 -13 2524 13
rect 2560 -13 2586 13
rect 2622 -13 2648 13
rect 2684 -13 2710 13
rect 2746 -13 2772 13
rect -2772 -75 -2746 -49
rect -2710 -75 -2684 -49
rect -2648 -75 -2622 -49
rect -2586 -75 -2560 -49
rect -2524 -75 -2498 -49
rect -2462 -75 -2436 -49
rect -2400 -75 -2374 -49
rect -2338 -75 -2312 -49
rect -2276 -75 -2250 -49
rect -2214 -75 -2188 -49
rect -2152 -75 -2126 -49
rect -2090 -75 -2064 -49
rect -2028 -75 -2002 -49
rect -1966 -75 -1940 -49
rect -1904 -75 -1878 -49
rect -1842 -75 -1816 -49
rect -1780 -75 -1754 -49
rect -1718 -75 -1692 -49
rect -1656 -75 -1630 -49
rect -1594 -75 -1568 -49
rect -1532 -75 -1506 -49
rect -1470 -75 -1444 -49
rect -1408 -75 -1382 -49
rect -1346 -75 -1320 -49
rect -1284 -75 -1258 -49
rect -1222 -75 -1196 -49
rect -1160 -75 -1134 -49
rect -1098 -75 -1072 -49
rect -1036 -75 -1010 -49
rect -974 -75 -948 -49
rect -912 -75 -886 -49
rect -850 -75 -824 -49
rect -788 -75 -762 -49
rect -726 -75 -700 -49
rect -664 -75 -638 -49
rect -602 -75 -576 -49
rect -540 -75 -514 -49
rect -478 -75 -452 -49
rect -416 -75 -390 -49
rect -354 -75 -328 -49
rect -292 -75 -266 -49
rect -230 -75 -204 -49
rect -168 -75 -142 -49
rect -106 -75 -80 -49
rect -44 -75 -18 -49
rect 18 -75 44 -49
rect 80 -75 106 -49
rect 142 -75 168 -49
rect 204 -75 230 -49
rect 266 -75 292 -49
rect 328 -75 354 -49
rect 390 -75 416 -49
rect 452 -75 478 -49
rect 514 -75 540 -49
rect 576 -75 602 -49
rect 638 -75 664 -49
rect 700 -75 726 -49
rect 762 -75 788 -49
rect 824 -75 850 -49
rect 886 -75 912 -49
rect 948 -75 974 -49
rect 1010 -75 1036 -49
rect 1072 -75 1098 -49
rect 1134 -75 1160 -49
rect 1196 -75 1222 -49
rect 1258 -75 1284 -49
rect 1320 -75 1346 -49
rect 1382 -75 1408 -49
rect 1444 -75 1470 -49
rect 1506 -75 1532 -49
rect 1568 -75 1594 -49
rect 1630 -75 1656 -49
rect 1692 -75 1718 -49
rect 1754 -75 1780 -49
rect 1816 -75 1842 -49
rect 1878 -75 1904 -49
rect 1940 -75 1966 -49
rect 2002 -75 2028 -49
rect 2064 -75 2090 -49
rect 2126 -75 2152 -49
rect 2188 -75 2214 -49
rect 2250 -75 2276 -49
rect 2312 -75 2338 -49
rect 2374 -75 2400 -49
rect 2436 -75 2462 -49
rect 2498 -75 2524 -49
rect 2560 -75 2586 -49
rect 2622 -75 2648 -49
rect 2684 -75 2710 -49
rect 2746 -75 2772 -49
<< metal2 >>
rect -2778 75 2778 81
rect -2778 49 -2772 75
rect -2746 49 -2710 75
rect -2684 49 -2648 75
rect -2622 49 -2586 75
rect -2560 49 -2524 75
rect -2498 49 -2462 75
rect -2436 49 -2400 75
rect -2374 49 -2338 75
rect -2312 49 -2276 75
rect -2250 49 -2214 75
rect -2188 49 -2152 75
rect -2126 49 -2090 75
rect -2064 49 -2028 75
rect -2002 49 -1966 75
rect -1940 49 -1904 75
rect -1878 49 -1842 75
rect -1816 49 -1780 75
rect -1754 49 -1718 75
rect -1692 49 -1656 75
rect -1630 49 -1594 75
rect -1568 49 -1532 75
rect -1506 49 -1470 75
rect -1444 49 -1408 75
rect -1382 49 -1346 75
rect -1320 49 -1284 75
rect -1258 49 -1222 75
rect -1196 49 -1160 75
rect -1134 49 -1098 75
rect -1072 49 -1036 75
rect -1010 49 -974 75
rect -948 49 -912 75
rect -886 49 -850 75
rect -824 49 -788 75
rect -762 49 -726 75
rect -700 49 -664 75
rect -638 49 -602 75
rect -576 49 -540 75
rect -514 49 -478 75
rect -452 49 -416 75
rect -390 49 -354 75
rect -328 49 -292 75
rect -266 49 -230 75
rect -204 49 -168 75
rect -142 49 -106 75
rect -80 49 -44 75
rect -18 49 18 75
rect 44 49 80 75
rect 106 49 142 75
rect 168 49 204 75
rect 230 49 266 75
rect 292 49 328 75
rect 354 49 390 75
rect 416 49 452 75
rect 478 49 514 75
rect 540 49 576 75
rect 602 49 638 75
rect 664 49 700 75
rect 726 49 762 75
rect 788 49 824 75
rect 850 49 886 75
rect 912 49 948 75
rect 974 49 1010 75
rect 1036 49 1072 75
rect 1098 49 1134 75
rect 1160 49 1196 75
rect 1222 49 1258 75
rect 1284 49 1320 75
rect 1346 49 1382 75
rect 1408 49 1444 75
rect 1470 49 1506 75
rect 1532 49 1568 75
rect 1594 49 1630 75
rect 1656 49 1692 75
rect 1718 49 1754 75
rect 1780 49 1816 75
rect 1842 49 1878 75
rect 1904 49 1940 75
rect 1966 49 2002 75
rect 2028 49 2064 75
rect 2090 49 2126 75
rect 2152 49 2188 75
rect 2214 49 2250 75
rect 2276 49 2312 75
rect 2338 49 2374 75
rect 2400 49 2436 75
rect 2462 49 2498 75
rect 2524 49 2560 75
rect 2586 49 2622 75
rect 2648 49 2684 75
rect 2710 49 2746 75
rect 2772 49 2778 75
rect -2778 13 2778 49
rect -2778 -13 -2772 13
rect -2746 -13 -2710 13
rect -2684 -13 -2648 13
rect -2622 -13 -2586 13
rect -2560 -13 -2524 13
rect -2498 -13 -2462 13
rect -2436 -13 -2400 13
rect -2374 -13 -2338 13
rect -2312 -13 -2276 13
rect -2250 -13 -2214 13
rect -2188 -13 -2152 13
rect -2126 -13 -2090 13
rect -2064 -13 -2028 13
rect -2002 -13 -1966 13
rect -1940 -13 -1904 13
rect -1878 -13 -1842 13
rect -1816 -13 -1780 13
rect -1754 -13 -1718 13
rect -1692 -13 -1656 13
rect -1630 -13 -1594 13
rect -1568 -13 -1532 13
rect -1506 -13 -1470 13
rect -1444 -13 -1408 13
rect -1382 -13 -1346 13
rect -1320 -13 -1284 13
rect -1258 -13 -1222 13
rect -1196 -13 -1160 13
rect -1134 -13 -1098 13
rect -1072 -13 -1036 13
rect -1010 -13 -974 13
rect -948 -13 -912 13
rect -886 -13 -850 13
rect -824 -13 -788 13
rect -762 -13 -726 13
rect -700 -13 -664 13
rect -638 -13 -602 13
rect -576 -13 -540 13
rect -514 -13 -478 13
rect -452 -13 -416 13
rect -390 -13 -354 13
rect -328 -13 -292 13
rect -266 -13 -230 13
rect -204 -13 -168 13
rect -142 -13 -106 13
rect -80 -13 -44 13
rect -18 -13 18 13
rect 44 -13 80 13
rect 106 -13 142 13
rect 168 -13 204 13
rect 230 -13 266 13
rect 292 -13 328 13
rect 354 -13 390 13
rect 416 -13 452 13
rect 478 -13 514 13
rect 540 -13 576 13
rect 602 -13 638 13
rect 664 -13 700 13
rect 726 -13 762 13
rect 788 -13 824 13
rect 850 -13 886 13
rect 912 -13 948 13
rect 974 -13 1010 13
rect 1036 -13 1072 13
rect 1098 -13 1134 13
rect 1160 -13 1196 13
rect 1222 -13 1258 13
rect 1284 -13 1320 13
rect 1346 -13 1382 13
rect 1408 -13 1444 13
rect 1470 -13 1506 13
rect 1532 -13 1568 13
rect 1594 -13 1630 13
rect 1656 -13 1692 13
rect 1718 -13 1754 13
rect 1780 -13 1816 13
rect 1842 -13 1878 13
rect 1904 -13 1940 13
rect 1966 -13 2002 13
rect 2028 -13 2064 13
rect 2090 -13 2126 13
rect 2152 -13 2188 13
rect 2214 -13 2250 13
rect 2276 -13 2312 13
rect 2338 -13 2374 13
rect 2400 -13 2436 13
rect 2462 -13 2498 13
rect 2524 -13 2560 13
rect 2586 -13 2622 13
rect 2648 -13 2684 13
rect 2710 -13 2746 13
rect 2772 -13 2778 13
rect -2778 -49 2778 -13
rect -2778 -75 -2772 -49
rect -2746 -75 -2710 -49
rect -2684 -75 -2648 -49
rect -2622 -75 -2586 -49
rect -2560 -75 -2524 -49
rect -2498 -75 -2462 -49
rect -2436 -75 -2400 -49
rect -2374 -75 -2338 -49
rect -2312 -75 -2276 -49
rect -2250 -75 -2214 -49
rect -2188 -75 -2152 -49
rect -2126 -75 -2090 -49
rect -2064 -75 -2028 -49
rect -2002 -75 -1966 -49
rect -1940 -75 -1904 -49
rect -1878 -75 -1842 -49
rect -1816 -75 -1780 -49
rect -1754 -75 -1718 -49
rect -1692 -75 -1656 -49
rect -1630 -75 -1594 -49
rect -1568 -75 -1532 -49
rect -1506 -75 -1470 -49
rect -1444 -75 -1408 -49
rect -1382 -75 -1346 -49
rect -1320 -75 -1284 -49
rect -1258 -75 -1222 -49
rect -1196 -75 -1160 -49
rect -1134 -75 -1098 -49
rect -1072 -75 -1036 -49
rect -1010 -75 -974 -49
rect -948 -75 -912 -49
rect -886 -75 -850 -49
rect -824 -75 -788 -49
rect -762 -75 -726 -49
rect -700 -75 -664 -49
rect -638 -75 -602 -49
rect -576 -75 -540 -49
rect -514 -75 -478 -49
rect -452 -75 -416 -49
rect -390 -75 -354 -49
rect -328 -75 -292 -49
rect -266 -75 -230 -49
rect -204 -75 -168 -49
rect -142 -75 -106 -49
rect -80 -75 -44 -49
rect -18 -75 18 -49
rect 44 -75 80 -49
rect 106 -75 142 -49
rect 168 -75 204 -49
rect 230 -75 266 -49
rect 292 -75 328 -49
rect 354 -75 390 -49
rect 416 -75 452 -49
rect 478 -75 514 -49
rect 540 -75 576 -49
rect 602 -75 638 -49
rect 664 -75 700 -49
rect 726 -75 762 -49
rect 788 -75 824 -49
rect 850 -75 886 -49
rect 912 -75 948 -49
rect 974 -75 1010 -49
rect 1036 -75 1072 -49
rect 1098 -75 1134 -49
rect 1160 -75 1196 -49
rect 1222 -75 1258 -49
rect 1284 -75 1320 -49
rect 1346 -75 1382 -49
rect 1408 -75 1444 -49
rect 1470 -75 1506 -49
rect 1532 -75 1568 -49
rect 1594 -75 1630 -49
rect 1656 -75 1692 -49
rect 1718 -75 1754 -49
rect 1780 -75 1816 -49
rect 1842 -75 1878 -49
rect 1904 -75 1940 -49
rect 1966 -75 2002 -49
rect 2028 -75 2064 -49
rect 2090 -75 2126 -49
rect 2152 -75 2188 -49
rect 2214 -75 2250 -49
rect 2276 -75 2312 -49
rect 2338 -75 2374 -49
rect 2400 -75 2436 -49
rect 2462 -75 2498 -49
rect 2524 -75 2560 -49
rect 2586 -75 2622 -49
rect 2648 -75 2684 -49
rect 2710 -75 2746 -49
rect 2772 -75 2778 -49
rect -2778 -81 2778 -75
<< end >>
