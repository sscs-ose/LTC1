magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1285 -1285 1285 1285
<< metal2 >>
rect -285 280 285 285
rect -285 252 -280 280
rect -252 252 -204 280
rect -176 252 -128 280
rect -100 252 -52 280
rect -24 252 24 280
rect 52 252 100 280
rect 128 252 176 280
rect 204 252 252 280
rect 280 252 285 280
rect -285 204 285 252
rect -285 176 -280 204
rect -252 176 -204 204
rect -176 176 -128 204
rect -100 176 -52 204
rect -24 176 24 204
rect 52 176 100 204
rect 128 176 176 204
rect 204 176 252 204
rect 280 176 285 204
rect -285 128 285 176
rect -285 100 -280 128
rect -252 100 -204 128
rect -176 100 -128 128
rect -100 100 -52 128
rect -24 100 24 128
rect 52 100 100 128
rect 128 100 176 128
rect 204 100 252 128
rect 280 100 285 128
rect -285 52 285 100
rect -285 24 -280 52
rect -252 24 -204 52
rect -176 24 -128 52
rect -100 24 -52 52
rect -24 24 24 52
rect 52 24 100 52
rect 128 24 176 52
rect 204 24 252 52
rect 280 24 285 52
rect -285 -24 285 24
rect -285 -52 -280 -24
rect -252 -52 -204 -24
rect -176 -52 -128 -24
rect -100 -52 -52 -24
rect -24 -52 24 -24
rect 52 -52 100 -24
rect 128 -52 176 -24
rect 204 -52 252 -24
rect 280 -52 285 -24
rect -285 -100 285 -52
rect -285 -128 -280 -100
rect -252 -128 -204 -100
rect -176 -128 -128 -100
rect -100 -128 -52 -100
rect -24 -128 24 -100
rect 52 -128 100 -100
rect 128 -128 176 -100
rect 204 -128 252 -100
rect 280 -128 285 -100
rect -285 -176 285 -128
rect -285 -204 -280 -176
rect -252 -204 -204 -176
rect -176 -204 -128 -176
rect -100 -204 -52 -176
rect -24 -204 24 -176
rect 52 -204 100 -176
rect 128 -204 176 -176
rect 204 -204 252 -176
rect 280 -204 285 -176
rect -285 -252 285 -204
rect -285 -280 -280 -252
rect -252 -280 -204 -252
rect -176 -280 -128 -252
rect -100 -280 -52 -252
rect -24 -280 24 -252
rect 52 -280 100 -252
rect 128 -280 176 -252
rect 204 -280 252 -252
rect 280 -280 285 -252
rect -285 -285 285 -280
<< via2 >>
rect -280 252 -252 280
rect -204 252 -176 280
rect -128 252 -100 280
rect -52 252 -24 280
rect 24 252 52 280
rect 100 252 128 280
rect 176 252 204 280
rect 252 252 280 280
rect -280 176 -252 204
rect -204 176 -176 204
rect -128 176 -100 204
rect -52 176 -24 204
rect 24 176 52 204
rect 100 176 128 204
rect 176 176 204 204
rect 252 176 280 204
rect -280 100 -252 128
rect -204 100 -176 128
rect -128 100 -100 128
rect -52 100 -24 128
rect 24 100 52 128
rect 100 100 128 128
rect 176 100 204 128
rect 252 100 280 128
rect -280 24 -252 52
rect -204 24 -176 52
rect -128 24 -100 52
rect -52 24 -24 52
rect 24 24 52 52
rect 100 24 128 52
rect 176 24 204 52
rect 252 24 280 52
rect -280 -52 -252 -24
rect -204 -52 -176 -24
rect -128 -52 -100 -24
rect -52 -52 -24 -24
rect 24 -52 52 -24
rect 100 -52 128 -24
rect 176 -52 204 -24
rect 252 -52 280 -24
rect -280 -128 -252 -100
rect -204 -128 -176 -100
rect -128 -128 -100 -100
rect -52 -128 -24 -100
rect 24 -128 52 -100
rect 100 -128 128 -100
rect 176 -128 204 -100
rect 252 -128 280 -100
rect -280 -204 -252 -176
rect -204 -204 -176 -176
rect -128 -204 -100 -176
rect -52 -204 -24 -176
rect 24 -204 52 -176
rect 100 -204 128 -176
rect 176 -204 204 -176
rect 252 -204 280 -176
rect -280 -280 -252 -252
rect -204 -280 -176 -252
rect -128 -280 -100 -252
rect -52 -280 -24 -252
rect 24 -280 52 -252
rect 100 -280 128 -252
rect 176 -280 204 -252
rect 252 -280 280 -252
<< metal3 >>
rect -285 280 285 285
rect -285 252 -280 280
rect -252 252 -204 280
rect -176 252 -128 280
rect -100 252 -52 280
rect -24 252 24 280
rect 52 252 100 280
rect 128 252 176 280
rect 204 252 252 280
rect 280 252 285 280
rect -285 204 285 252
rect -285 176 -280 204
rect -252 176 -204 204
rect -176 176 -128 204
rect -100 176 -52 204
rect -24 176 24 204
rect 52 176 100 204
rect 128 176 176 204
rect 204 176 252 204
rect 280 176 285 204
rect -285 128 285 176
rect -285 100 -280 128
rect -252 100 -204 128
rect -176 100 -128 128
rect -100 100 -52 128
rect -24 100 24 128
rect 52 100 100 128
rect 128 100 176 128
rect 204 100 252 128
rect 280 100 285 128
rect -285 52 285 100
rect -285 24 -280 52
rect -252 24 -204 52
rect -176 24 -128 52
rect -100 24 -52 52
rect -24 24 24 52
rect 52 24 100 52
rect 128 24 176 52
rect 204 24 252 52
rect 280 24 285 52
rect -285 -24 285 24
rect -285 -52 -280 -24
rect -252 -52 -204 -24
rect -176 -52 -128 -24
rect -100 -52 -52 -24
rect -24 -52 24 -24
rect 52 -52 100 -24
rect 128 -52 176 -24
rect 204 -52 252 -24
rect 280 -52 285 -24
rect -285 -100 285 -52
rect -285 -128 -280 -100
rect -252 -128 -204 -100
rect -176 -128 -128 -100
rect -100 -128 -52 -100
rect -24 -128 24 -100
rect 52 -128 100 -100
rect 128 -128 176 -100
rect 204 -128 252 -100
rect 280 -128 285 -100
rect -285 -176 285 -128
rect -285 -204 -280 -176
rect -252 -204 -204 -176
rect -176 -204 -128 -176
rect -100 -204 -52 -176
rect -24 -204 24 -176
rect 52 -204 100 -176
rect 128 -204 176 -176
rect 204 -204 252 -176
rect 280 -204 285 -176
rect -285 -252 285 -204
rect -285 -280 -280 -252
rect -252 -280 -204 -252
rect -176 -280 -128 -252
rect -100 -280 -52 -252
rect -24 -280 24 -252
rect 52 -280 100 -252
rect 128 -280 176 -252
rect 204 -280 252 -252
rect 280 -280 285 -252
rect -285 -285 285 -280
<< end >>
