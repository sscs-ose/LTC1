magic
tech gf180mcuC
magscale 1 10
timestamp 1714490790
<< nwell >>
rect 0 875 434 950
rect 0 820 5956 875
rect 0 770 608 820
rect 673 770 852 820
rect 918 770 1097 820
rect 1162 770 1341 820
rect 1407 770 1586 820
rect 1652 770 1831 820
rect 1896 770 2075 820
rect 2141 770 2320 820
rect 2386 770 2565 820
rect 2630 770 2809 820
rect 2885 785 2886 820
rect 2885 772 3062 785
rect 3313 772 3495 820
rect 3733 772 3915 820
rect 4155 772 4337 820
rect 4577 772 4759 820
rect 5052 772 5234 820
rect 5527 772 5709 820
rect 0 752 434 770
<< pwell >>
rect 2920 -2260 2970 -2254
rect 3327 -2260 3381 -2253
rect 3735 -2260 3791 -2252
rect 4144 -2260 4198 -2253
rect 4551 -2260 4605 -2254
rect 4959 -2260 5014 -2254
rect 5368 -2260 5429 -2254
<< psubdiff >>
rect 68 -3064 244 -3051
rect 68 -3115 91 -3064
rect 228 -3115 244 -3064
rect 68 -3130 244 -3115
rect 368 -3064 544 -3051
rect 368 -3115 391 -3064
rect 528 -3115 544 -3064
rect 368 -3130 544 -3115
rect 668 -3064 844 -3051
rect 668 -3115 691 -3064
rect 828 -3115 844 -3064
rect 668 -3130 844 -3115
rect 968 -3064 1144 -3051
rect 968 -3115 991 -3064
rect 1128 -3115 1144 -3064
rect 968 -3130 1144 -3115
rect 1268 -3064 1444 -3051
rect 1268 -3115 1291 -3064
rect 1428 -3115 1444 -3064
rect 1268 -3130 1444 -3115
rect 1568 -3064 1744 -3051
rect 1568 -3115 1591 -3064
rect 1728 -3115 1744 -3064
rect 1568 -3130 1744 -3115
rect 1868 -3064 2044 -3051
rect 1868 -3115 1891 -3064
rect 2028 -3115 2044 -3064
rect 1868 -3130 2044 -3115
rect 2168 -3064 2344 -3051
rect 2168 -3115 2191 -3064
rect 2328 -3115 2344 -3064
rect 2168 -3130 2344 -3115
rect 2468 -3064 2644 -3051
rect 2468 -3115 2491 -3064
rect 2628 -3115 2644 -3064
rect 2468 -3130 2644 -3115
rect 2768 -3064 2944 -3051
rect 2768 -3115 2791 -3064
rect 2928 -3115 2944 -3064
rect 2768 -3130 2944 -3115
rect 3068 -3064 3244 -3051
rect 3068 -3115 3091 -3064
rect 3228 -3115 3244 -3064
rect 3068 -3130 3244 -3115
rect 3368 -3064 3544 -3051
rect 3368 -3115 3391 -3064
rect 3528 -3115 3544 -3064
rect 3368 -3130 3544 -3115
rect 3668 -3064 3844 -3051
rect 3668 -3115 3691 -3064
rect 3828 -3115 3844 -3064
rect 3668 -3130 3844 -3115
rect 3968 -3064 4144 -3051
rect 3968 -3115 3991 -3064
rect 4128 -3115 4144 -3064
rect 3968 -3130 4144 -3115
rect 4268 -3064 4444 -3051
rect 4268 -3115 4291 -3064
rect 4428 -3115 4444 -3064
rect 4268 -3130 4444 -3115
rect 4568 -3064 4744 -3051
rect 4568 -3115 4591 -3064
rect 4728 -3115 4744 -3064
rect 4568 -3130 4744 -3115
rect 4868 -3064 5044 -3051
rect 4868 -3115 4891 -3064
rect 5028 -3115 5044 -3064
rect 4868 -3130 5044 -3115
rect 5168 -3064 5344 -3051
rect 5168 -3115 5191 -3064
rect 5328 -3115 5344 -3064
rect 5168 -3130 5344 -3115
rect 5468 -3064 5644 -3051
rect 5468 -3115 5491 -3064
rect 5628 -3115 5644 -3064
rect 5468 -3130 5644 -3115
rect 5718 -3064 5894 -3051
rect 5718 -3115 5741 -3064
rect 5878 -3115 5894 -3064
rect 5718 -3130 5894 -3115
<< nsubdiff >>
rect 128 911 296 925
rect 128 850 158 911
rect 251 850 296 911
rect 128 822 296 850
<< psubdiffcont >>
rect 91 -3115 228 -3064
rect 391 -3115 528 -3064
rect 691 -3115 828 -3064
rect 991 -3115 1128 -3064
rect 1291 -3115 1428 -3064
rect 1591 -3115 1728 -3064
rect 1891 -3115 2028 -3064
rect 2191 -3115 2328 -3064
rect 2491 -3115 2628 -3064
rect 2791 -3115 2928 -3064
rect 3091 -3115 3228 -3064
rect 3391 -3115 3528 -3064
rect 3691 -3115 3828 -3064
rect 3991 -3115 4128 -3064
rect 4291 -3115 4428 -3064
rect 4591 -3115 4728 -3064
rect 4891 -3115 5028 -3064
rect 5191 -3115 5328 -3064
rect 5491 -3115 5628 -3064
rect 5741 -3115 5878 -3064
<< nsubdiffcont >>
rect 158 850 251 911
<< polysilicon >>
rect 175 91 273 120
rect 786 91 878 121
rect 173 89 878 91
rect -158 64 878 89
rect -158 -4 -137 64
rect -85 -4 878 64
rect -158 -28 878 -4
rect 988 60 4150 86
rect 988 10 1009 60
rect 1059 10 4150 60
rect -158 -29 185 -28
rect 988 -30 4150 10
rect 4254 66 5782 88
rect 4254 16 4274 66
rect 4327 16 5782 66
rect 4254 -29 5782 16
rect 5681 -99 5782 -29
rect 174 -728 477 -727
rect 174 -776 5781 -728
rect 2620 -1433 2722 -1404
rect 2620 -1479 2640 -1433
rect 2697 -1479 2722 -1433
rect -161 -1492 -66 -1482
rect -161 -1500 451 -1492
rect -161 -1552 -146 -1500
rect -93 -1552 451 -1500
rect -161 -1563 451 -1552
rect 548 -1500 645 -1487
rect 548 -1547 564 -1500
rect 616 -1511 645 -1500
rect 2620 -1505 2722 -1479
rect 2826 -1490 2926 -1424
rect 3438 -1490 3538 -1424
rect 4050 -1490 4150 -1424
rect 4662 -1490 4762 -1424
rect 5274 -1490 5374 -1424
rect 616 -1547 2076 -1511
rect 548 -1560 2076 -1547
rect 2792 -1560 5748 -1490
rect -161 -1568 -66 -1563
rect 2179 -2203 2279 -2200
rect 2179 -2260 2892 -2203
rect 138 -2895 646 -2887
rect 138 -2897 2279 -2895
rect 138 -2984 2891 -2897
rect 2276 -2985 2891 -2984
rect 2996 -2915 5748 -2890
rect 2996 -2961 3226 -2915
rect 3279 -2961 5748 -2915
rect 2996 -3001 5748 -2961
<< polycontact >>
rect -137 -4 -85 64
rect 1009 10 1059 60
rect 4274 16 4327 66
rect 2640 -1479 2697 -1433
rect -146 -1552 -93 -1500
rect 564 -1547 616 -1500
rect 3226 -2961 3279 -2915
<< metal1 >>
rect 143 911 263 924
rect 143 876 158 911
rect 0 850 158 876
rect 251 876 263 911
rect 251 850 5956 876
rect 0 753 5956 850
rect 0 752 434 753
rect 99 677 145 752
rect 507 677 553 753
rect 914 675 961 753
rect 1323 677 1369 753
rect 1731 677 1777 753
rect 2139 677 2185 753
rect 2547 677 2593 753
rect 2955 677 3001 753
rect 3363 677 3409 753
rect 3771 676 3817 753
rect 4178 666 4226 753
rect 4587 675 4633 753
rect 4995 677 5041 753
rect 5403 678 5449 753
rect 5811 678 5857 753
rect 300 86 351 136
rect 709 86 758 147
rect -153 64 -76 78
rect -153 28 -137 64
rect -154 -4 -137 28
rect -85 -4 -76 64
rect 300 73 758 86
rect 1117 82 1166 166
rect 1526 82 1573 155
rect 1934 82 1981 156
rect 2343 82 2390 156
rect 2750 82 2797 154
rect 3158 82 3205 154
rect 3566 82 3613 154
rect 3974 82 4021 155
rect 1117 79 4021 82
rect 4383 80 4430 155
rect 4789 80 4836 155
rect 5198 80 5245 159
rect 5607 80 5654 155
rect 300 60 1070 73
rect 300 54 1009 60
rect -154 -16 -76 -4
rect -24 10 1009 54
rect 1059 10 1070 60
rect -24 9 1070 10
rect -24 8 758 9
rect -154 -73 -80 -16
rect -154 -1500 -85 -73
rect -154 -1552 -146 -1500
rect -93 -1552 -85 -1500
rect -154 -1568 -85 -1552
rect -24 -1508 22 8
rect 987 -5 1070 9
rect 1117 66 4336 79
rect 1117 16 4274 66
rect 4327 16 4336 66
rect 1117 3 4336 16
rect 4383 7 5654 80
rect 5606 -164 5654 7
rect 5811 -136 5857 145
rect 68 -318 169 -304
rect 68 -387 83 -318
rect 157 -387 169 -318
rect 68 -401 169 -387
rect 474 -311 575 -294
rect 474 -380 488 -311
rect 562 -380 575 -311
rect 474 -392 575 -380
rect 879 -310 979 -289
rect 879 -379 893 -310
rect 967 -379 979 -310
rect 1289 -297 1389 -277
rect 1289 -366 1303 -297
rect 1377 -366 1389 -297
rect 1289 -378 1389 -366
rect 1699 -293 1799 -274
rect 1699 -362 1711 -293
rect 1785 -362 1799 -293
rect 1699 -375 1799 -362
rect 2109 -284 2209 -265
rect 2109 -353 2121 -284
rect 2195 -353 2209 -284
rect 2109 -366 2209 -353
rect 2515 -283 2615 -265
rect 2515 -352 2530 -283
rect 2609 -352 2615 -283
rect 2515 -366 2615 -352
rect 2918 -274 3018 -255
rect 2918 -343 2934 -274
rect 3008 -343 3018 -274
rect 2918 -356 3018 -343
rect 3328 -271 3428 -249
rect 3328 -340 3344 -271
rect 3418 -340 3428 -271
rect 3328 -350 3428 -340
rect 3743 -269 3843 -250
rect 3743 -338 3755 -269
rect 3829 -338 3843 -269
rect 3743 -351 3843 -338
rect 4147 -271 4247 -251
rect 4147 -340 4160 -271
rect 4234 -340 4247 -271
rect 4147 -352 4247 -340
rect 4555 -271 4655 -255
rect 4555 -340 4570 -271
rect 4644 -340 4655 -271
rect 4555 -356 4655 -340
rect 4958 -271 5058 -251
rect 4958 -340 4971 -271
rect 5045 -340 5058 -271
rect 4958 -352 5058 -340
rect 5374 -267 5474 -247
rect 5374 -336 5387 -267
rect 5461 -336 5474 -267
rect 5374 -348 5474 -336
rect 5775 -252 5875 -236
rect 5775 -321 5788 -252
rect 5862 -321 5875 -252
rect 5775 -337 5875 -321
rect 879 -390 979 -379
rect 302 -728 349 -658
rect 711 -728 757 -658
rect 1119 -728 1165 -651
rect 1526 -728 1572 -651
rect 1934 -728 1980 -651
rect 2342 -728 2388 -651
rect 2751 -728 2797 -653
rect 3158 -728 3204 -651
rect 3566 -728 3612 -652
rect 3975 -728 4021 -660
rect 4382 -728 4428 -662
rect 4791 -728 4837 -658
rect 5198 -728 5244 -657
rect 5606 -728 5653 -662
rect 302 -775 5653 -728
rect 302 -844 349 -775
rect 710 -836 757 -775
rect 1119 -836 1166 -775
rect 1527 -836 1574 -775
rect 1935 -835 1982 -775
rect 2343 -835 2390 -775
rect 2751 -835 2798 -775
rect 3159 -835 3206 -775
rect 3567 -835 3614 -775
rect 3975 -834 4022 -775
rect 4383 -834 4430 -775
rect 4792 -834 4839 -775
rect 5200 -834 5247 -775
rect 5606 -833 5653 -775
rect 5810 -838 5857 -667
rect 68 -1012 183 -988
rect 68 -1081 87 -1012
rect 166 -1081 183 -1012
rect 68 -1097 183 -1081
rect 471 -1006 586 -977
rect 471 -1075 486 -1006
rect 565 -1075 586 -1006
rect 471 -1086 586 -1075
rect 877 -1010 992 -981
rect 877 -1079 894 -1010
rect 973 -1079 992 -1010
rect 877 -1090 992 -1079
rect 1282 -1004 1397 -981
rect 1282 -1073 1299 -1004
rect 1378 -1073 1397 -1004
rect 1282 -1090 1397 -1073
rect 1692 -1021 1807 -995
rect 1692 -1090 1709 -1021
rect 1788 -1090 1807 -1021
rect 1692 -1104 1807 -1090
rect 2100 -1022 2215 -998
rect 2100 -1091 2117 -1022
rect 2196 -1091 2215 -1022
rect 2100 -1107 2215 -1091
rect 2504 -1033 2619 -1008
rect 2504 -1102 2525 -1033
rect 2604 -1102 2619 -1033
rect 2504 -1117 2619 -1102
rect 2918 -1043 3033 -1018
rect 2918 -1112 2937 -1043
rect 3016 -1112 3033 -1043
rect 3330 -1029 3445 -1003
rect 3330 -1098 3348 -1029
rect 3427 -1098 3445 -1029
rect 3330 -1112 3445 -1098
rect 3737 -1027 3852 -1006
rect 3737 -1096 3755 -1027
rect 3834 -1096 3852 -1027
rect 2918 -1127 3033 -1112
rect 3737 -1115 3852 -1096
rect 4139 -1024 4254 -999
rect 4139 -1093 4162 -1024
rect 4241 -1093 4254 -1024
rect 4550 -1008 4665 -981
rect 4550 -1077 4567 -1008
rect 4646 -1077 4665 -1008
rect 4550 -1090 4665 -1077
rect 4966 -996 5081 -972
rect 4966 -1065 4980 -996
rect 5059 -1065 5081 -996
rect 4966 -1081 5081 -1065
rect 5372 -990 5487 -964
rect 5372 -1059 5388 -990
rect 5467 -1059 5487 -990
rect 5372 -1073 5487 -1059
rect 5769 -982 5884 -959
rect 5769 -1051 5790 -982
rect 5869 -1051 5884 -982
rect 5769 -1068 5884 -1051
rect 4139 -1108 4254 -1093
rect 2621 -1428 2718 -1415
rect 2621 -1483 2635 -1428
rect 2702 -1483 2718 -1428
rect 5607 -1438 5654 -1286
rect 258 -1500 628 -1487
rect 2621 -1495 2718 -1483
rect 258 -1508 564 -1500
rect -24 -1547 564 -1508
rect 616 -1547 628 -1500
rect -24 -1554 628 -1547
rect 269 -1617 315 -1554
rect 548 -1560 628 -1554
rect 5572 -1509 5955 -1438
rect 5572 -1615 5619 -1509
rect 654 -1821 743 -1810
rect 654 -1874 668 -1821
rect 731 -1874 743 -1821
rect 654 -1884 743 -1874
rect 1060 -1812 1149 -1798
rect 1060 -1865 1074 -1812
rect 1137 -1865 1149 -1812
rect 1470 -1800 1559 -1785
rect 1470 -1853 1485 -1800
rect 1548 -1853 1559 -1800
rect 1470 -1863 1559 -1853
rect 1875 -1792 1964 -1778
rect 1875 -1845 1889 -1792
rect 1952 -1845 1964 -1792
rect 1875 -1856 1964 -1845
rect 1060 -1876 1149 -1865
rect 2289 -2042 2379 -2029
rect 2289 -2101 2299 -2042
rect 2368 -2101 2379 -2042
rect 2289 -2114 2379 -2101
rect 2692 -2042 2782 -2029
rect 2692 -2099 2704 -2042
rect 2771 -2099 2782 -2042
rect 2692 -2111 2782 -2099
rect 3098 -2039 3192 -2025
rect 3098 -2094 3111 -2039
rect 3181 -2094 3192 -2039
rect 3098 -2105 3192 -2094
rect 3509 -2029 3596 -2016
rect 3509 -2085 3520 -2029
rect 3586 -2085 3596 -2029
rect 3916 -2018 4006 -2005
rect 3916 -2074 3929 -2018
rect 3995 -2074 4006 -2018
rect 3916 -2085 4006 -2074
rect 4324 -2021 4415 -2006
rect 4324 -2076 4338 -2021
rect 4405 -2076 4415 -2021
rect 3509 -2095 3596 -2085
rect 4324 -2089 4415 -2076
rect 4733 -2018 4826 -2005
rect 4733 -2072 4745 -2018
rect 4814 -2072 4826 -2018
rect 4733 -2085 4826 -2072
rect 5142 -2019 5231 -2005
rect 5142 -2073 5153 -2019
rect 5219 -2073 5231 -2019
rect 5142 -2085 5231 -2073
rect 5552 -2021 5640 -2008
rect 5552 -2074 5563 -2021
rect 5629 -2074 5640 -2021
rect 5552 -2086 5640 -2074
rect 64 -2208 111 -2149
rect 472 -2208 519 -2147
rect 881 -2208 928 -2149
rect 1289 -2208 1336 -2148
rect 1696 -2208 1743 -2148
rect 2104 -2208 2151 -2149
rect 2513 -2208 2560 -2147
rect 2920 -2208 2967 -2149
rect 3328 -2208 3375 -2149
rect 3737 -2208 3784 -2149
rect 4145 -2208 4192 -2149
rect 4553 -2208 4600 -2148
rect 4961 -2208 5008 -2148
rect 5369 -2208 5416 -2147
rect 5776 -2208 5823 -2149
rect 64 -2254 5823 -2208
rect 64 -2313 111 -2254
rect 472 -2313 519 -2254
rect 881 -2313 928 -2254
rect 1289 -2312 1336 -2254
rect 1696 -2312 1743 -2254
rect 2104 -2313 2151 -2254
rect 2513 -2311 2560 -2254
rect 2921 -2553 2997 -2254
rect 248 -2603 334 -2589
rect 248 -2659 261 -2603
rect 323 -2659 334 -2603
rect 248 -2671 334 -2659
rect 657 -2598 743 -2583
rect 657 -2654 669 -2598
rect 731 -2654 743 -2598
rect 657 -2666 743 -2654
rect 1063 -2596 1149 -2582
rect 1063 -2652 1076 -2596
rect 1138 -2652 1149 -2596
rect 1063 -2665 1149 -2652
rect 1473 -2596 1560 -2583
rect 1473 -2652 1486 -2596
rect 1548 -2652 1560 -2596
rect 1473 -2665 1560 -2652
rect 1882 -2596 1969 -2582
rect 1882 -2652 1894 -2596
rect 1956 -2652 1969 -2596
rect 1882 -2664 1969 -2652
rect 2287 -2595 2374 -2581
rect 2287 -2651 2299 -2595
rect 2361 -2651 2374 -2595
rect 2287 -2663 2374 -2651
rect 2695 -2594 2782 -2580
rect 2695 -2650 2707 -2594
rect 2769 -2650 2782 -2594
rect 2921 -2645 5822 -2553
rect 2695 -2662 2782 -2650
rect 65 -3024 111 -2858
rect 881 -3024 927 -2858
rect 1691 -3024 1751 -2832
rect 2503 -3024 2563 -2835
rect 3220 -2915 3282 -2645
rect 3220 -2961 3226 -2915
rect 3279 -2961 3282 -2915
rect 3220 -2973 3282 -2961
rect 3724 -3024 3784 -2833
rect 4954 -3024 5014 -2844
rect 0 -3064 5956 -3024
rect 0 -3115 91 -3064
rect 228 -3115 391 -3064
rect 528 -3115 691 -3064
rect 828 -3115 991 -3064
rect 1128 -3115 1291 -3064
rect 1428 -3115 1591 -3064
rect 1728 -3115 1891 -3064
rect 2028 -3115 2191 -3064
rect 2328 -3115 2491 -3064
rect 2628 -3115 2791 -3064
rect 2928 -3115 3091 -3064
rect 3228 -3115 3391 -3064
rect 3528 -3115 3691 -3064
rect 3828 -3115 3991 -3064
rect 4128 -3115 4291 -3064
rect 4428 -3115 4591 -3064
rect 4728 -3115 4891 -3064
rect 5028 -3115 5191 -3064
rect 5328 -3115 5491 -3064
rect 5628 -3115 5741 -3064
rect 5878 -3115 5956 -3064
rect 0 -3147 5956 -3115
<< via1 >>
rect 83 -387 157 -318
rect 488 -380 562 -311
rect 893 -379 967 -310
rect 1303 -366 1377 -297
rect 1711 -362 1785 -293
rect 2121 -353 2195 -284
rect 2530 -352 2609 -283
rect 2934 -343 3008 -274
rect 3344 -340 3418 -271
rect 3755 -338 3829 -269
rect 4160 -340 4234 -271
rect 4570 -340 4644 -271
rect 4971 -340 5045 -271
rect 5387 -336 5461 -267
rect 5788 -321 5862 -252
rect 87 -1081 166 -1012
rect 486 -1075 565 -1006
rect 894 -1079 973 -1010
rect 1299 -1073 1378 -1004
rect 1709 -1090 1788 -1021
rect 2117 -1091 2196 -1022
rect 2525 -1102 2604 -1033
rect 2937 -1112 3016 -1043
rect 3348 -1098 3427 -1029
rect 3755 -1096 3834 -1027
rect 4162 -1093 4241 -1024
rect 4567 -1077 4646 -1008
rect 4980 -1065 5059 -996
rect 5388 -1059 5467 -990
rect 5790 -1051 5869 -982
rect 2635 -1433 2702 -1428
rect 2635 -1479 2640 -1433
rect 2640 -1479 2697 -1433
rect 2697 -1479 2702 -1433
rect 2635 -1483 2702 -1479
rect 668 -1874 731 -1821
rect 1074 -1865 1137 -1812
rect 1485 -1853 1548 -1800
rect 1889 -1845 1952 -1792
rect 2299 -2101 2368 -2042
rect 2704 -2099 2771 -2042
rect 3111 -2094 3181 -2039
rect 3520 -2085 3586 -2029
rect 3929 -2074 3995 -2018
rect 4338 -2076 4405 -2021
rect 4745 -2072 4814 -2018
rect 5153 -2073 5219 -2019
rect 5563 -2074 5629 -2021
rect 261 -2659 323 -2603
rect 669 -2654 731 -2598
rect 1076 -2652 1138 -2596
rect 1486 -2652 1548 -2596
rect 1894 -2652 1956 -2596
rect 2299 -2651 2361 -2595
rect 2707 -2650 2769 -2594
<< metal2 >>
rect 66 -252 5875 -234
rect 66 -267 5788 -252
rect 66 -269 5387 -267
rect 66 -271 3755 -269
rect 66 -274 3344 -271
rect 66 -283 2934 -274
rect 66 -284 2530 -283
rect 66 -293 2121 -284
rect 66 -297 1711 -293
rect 66 -310 1303 -297
rect 66 -311 893 -310
rect 66 -318 488 -311
rect 66 -387 83 -318
rect 157 -380 488 -318
rect 562 -379 893 -311
rect 967 -366 1303 -310
rect 1377 -362 1711 -297
rect 1785 -353 2121 -293
rect 2195 -352 2530 -284
rect 2609 -343 2934 -283
rect 3008 -340 3344 -274
rect 3418 -338 3755 -271
rect 3829 -271 5387 -269
rect 3829 -338 4160 -271
rect 3418 -340 4160 -338
rect 4234 -340 4570 -271
rect 4644 -340 4971 -271
rect 5045 -336 5387 -271
rect 5461 -321 5788 -267
rect 5862 -321 5875 -252
rect 5461 -336 5875 -321
rect 5045 -340 5875 -336
rect 3008 -343 5875 -340
rect 2609 -352 5875 -343
rect 2195 -353 5875 -352
rect 1785 -362 5875 -353
rect 1377 -366 5875 -362
rect 967 -379 5875 -366
rect 562 -380 5875 -379
rect 157 -387 5875 -380
rect 66 -400 5875 -387
rect 68 -401 169 -400
rect 61 -982 5885 -949
rect 61 -990 5790 -982
rect 61 -996 5388 -990
rect 61 -1004 4980 -996
rect 61 -1006 1299 -1004
rect 61 -1012 486 -1006
rect 61 -1081 87 -1012
rect 166 -1075 486 -1012
rect 565 -1010 1299 -1006
rect 565 -1075 894 -1010
rect 166 -1079 894 -1075
rect 973 -1073 1299 -1010
rect 1378 -1008 4980 -1004
rect 1378 -1021 4567 -1008
rect 1378 -1073 1709 -1021
rect 973 -1079 1709 -1073
rect 166 -1081 1709 -1079
rect 61 -1090 1709 -1081
rect 1788 -1022 4567 -1021
rect 1788 -1090 2117 -1022
rect 61 -1091 2117 -1090
rect 2196 -1024 4567 -1022
rect 2196 -1027 4162 -1024
rect 2196 -1029 3755 -1027
rect 2196 -1033 3348 -1029
rect 2196 -1091 2525 -1033
rect 61 -1102 2525 -1091
rect 2604 -1043 3348 -1033
rect 2604 -1102 2937 -1043
rect 61 -1108 2937 -1102
rect 2504 -1117 2619 -1108
rect 2918 -1112 2937 -1108
rect 3016 -1098 3348 -1043
rect 3427 -1096 3755 -1029
rect 3834 -1093 4162 -1027
rect 4241 -1077 4567 -1024
rect 4646 -1065 4980 -1008
rect 5059 -1059 5388 -996
rect 5467 -1051 5790 -990
rect 5869 -1051 5885 -982
rect 5467 -1059 5885 -1051
rect 5059 -1065 5885 -1059
rect 4646 -1077 5885 -1065
rect 4241 -1093 5885 -1077
rect 3834 -1096 5885 -1093
rect 3427 -1098 5885 -1096
rect 3016 -1108 5885 -1098
rect 3016 -1112 3033 -1108
rect 3330 -1112 3445 -1108
rect 2918 -1127 3033 -1112
rect 3737 -1115 3852 -1108
rect 2619 -1428 2718 -1413
rect 2619 -1483 2635 -1428
rect 2702 -1483 2718 -1428
rect 2619 -1773 2718 -1483
rect 1883 -1775 2718 -1773
rect 653 -1792 2718 -1775
rect 653 -1800 1889 -1792
rect 653 -1812 1485 -1800
rect 653 -1821 1074 -1812
rect 653 -1874 668 -1821
rect 731 -1865 1074 -1821
rect 1137 -1853 1485 -1812
rect 1548 -1845 1889 -1800
rect 1952 -1845 2718 -1792
rect 1548 -1853 2718 -1845
rect 1137 -1865 2718 -1853
rect 731 -1874 2718 -1865
rect 653 -1884 2718 -1874
rect 2289 -2018 5640 -2003
rect 2289 -2029 3929 -2018
rect 2289 -2039 3520 -2029
rect 2289 -2042 3111 -2039
rect 2289 -2101 2299 -2042
rect 2368 -2099 2704 -2042
rect 2771 -2094 3111 -2042
rect 3181 -2085 3520 -2039
rect 3586 -2074 3929 -2029
rect 3995 -2021 4745 -2018
rect 3995 -2074 4338 -2021
rect 3586 -2076 4338 -2074
rect 4405 -2072 4745 -2021
rect 4814 -2019 5640 -2018
rect 4814 -2072 5153 -2019
rect 4405 -2073 5153 -2072
rect 5219 -2021 5640 -2019
rect 5219 -2073 5563 -2021
rect 4405 -2074 5563 -2073
rect 5629 -2074 5640 -2021
rect 4405 -2076 5640 -2074
rect 3586 -2085 5640 -2076
rect 3181 -2094 5640 -2085
rect 2771 -2099 5640 -2094
rect 2368 -2101 5640 -2099
rect 2289 -2114 5640 -2101
rect 2398 -2579 2480 -2114
rect 248 -2594 2791 -2579
rect 248 -2595 2707 -2594
rect 248 -2596 2299 -2595
rect 248 -2598 1076 -2596
rect 248 -2603 669 -2598
rect 248 -2659 261 -2603
rect 323 -2654 669 -2603
rect 731 -2652 1076 -2598
rect 1138 -2652 1486 -2596
rect 1548 -2652 1894 -2596
rect 1956 -2651 2299 -2596
rect 2361 -2650 2707 -2595
rect 2769 -2650 2791 -2594
rect 2361 -2651 2791 -2650
rect 1956 -2652 2791 -2651
rect 731 -2654 2791 -2652
rect 323 -2659 2791 -2654
rect 248 -2671 2791 -2659
use nmos_3p3_7NPLVN  nmos_3p3_7NPLVN_0
timestamp 1714126980
transform 1 0 2944 0 1 -2580
box -2916 -348 2916 348
use nmos_3p3_8FEAMQ  nmos_3p3_8FEAMQ_0
timestamp 1714126980
transform 1 0 292 0 1 -1884
box -264 -348 264 348
use nmos_3p3_JEEAMQ  nmos_3p3_JEEAMQ_0
timestamp 1714126980
transform 1 0 1312 0 1 -1884
box -876 -348 876 348
use nmos_3p3_PLQLVN  nmos_3p3_PLQLVN_0
timestamp 1714126980
transform 1 0 3964 0 1 -1884
box -1896 -348 1896 348
use pmos_3p3_MDMPD7  pmos_3p3_MDMPD7_0
timestamp 1714126980
transform 1 0 2978 0 1 -752
box -2978 -758 2978 758
use pmos_3p3_MV44E7  pmos_3p3_MV44E7_0
timestamp 1714126980
transform 1 0 2570 0 1 410
box -1754 -410 1754 410
use pmos_3p3_PPYSL5  pmos_3p3_PPYSL5_0
timestamp 1714126980
transform 1 0 530 0 1 410
box -530 -410 530 410
use pmos_3p3_PPZSL5  pmos_3p3_PPZSL5_0
timestamp 1714126980
transform 1 0 5018 0 1 410
box -938 -410 938 410
<< labels >>
flabel metal1 -131 -741 -131 -741 0 FreeSans 480 0 0 0 IN
port 2 nsew
flabel metal1 5909 -1469 5909 -1469 0 FreeSans 480 0 0 0 OUT
port 3 nsew
flabel psubdiffcont 2859 -3090 2859 -3090 0 FreeSans 480 0 0 0 VSS
port 4 nsew
flabel metal1 3404 811 3404 811 0 FreeSans 480 0 0 0 VDD
port 1 nsew
<< end >>
