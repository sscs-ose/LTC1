* NGSPICE file created from CLK_div_100_mag_flat.ext - technology: gf180mcuC

.subckt pex_CLK_div_100_mag VSS VDD RST Vdiv100 CLK
X0 a_6311_5223# CLK_div_10_mag_1.Q1.t3 CLK_div_10_mag_1.JK_FF_mag_2.QB VSS.t207 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1 VDD CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t133 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2 VDD VDD.t184 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VDD.t185 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_10_mag_0.Q1 VDD.t24 VDD.t23 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X4 a_8323_5223# CLK_div_10_mag_1.Q0.t3 a_8163_5223# VSS.t216 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X5 VDD CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_10_mag_1.JK_FF_mag_3.QB VDD.t357 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X6 a_5300_4126# CLK_div_10_mag_1.Q1.t4 a_5140_4126# VSS.t206 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X7 a_230_2335# CLK_div_10_mag_1.Q3 Vdiv100.t2 VDD.t72 pfet_03v3 ad=0.624p pd=2.92u as=1.06p ps=5.68u w=2.4u l=0.28u
X8 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 VDD.t320 VDD.t319 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X9 VDD CLK_div_10_mag_1.JK_FF_mag_0.J CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VDD.t297 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X10 a_794_1309# CLK.t0 a_634_1309# VSS.t296 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X11 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_2.QB a_5503_1353# VSS.t213 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X12 VDD VDD.t180 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT VDD.t181 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X13 VDD CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t64 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X14 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD.t90 VDD.t89 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X15 a_4375_1353# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VSS.t87 VSS.t86 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X16 VDD CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t423 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X17 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT RST.t0 VDD.t347 VDD.t346 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X18 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.Q0 VDD.t422 VDD.t421 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X19 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.J.t3 VDD.t93 VDD.t92 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X20 VSS CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT a_3858_5223# VSS.t120 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X21 CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_10_mag_1.Q2.t3 VDD.t194 VDD.t193 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X22 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD.t50 VDD.t49 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X23 VSS CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_1.CLK VSS.t65 nfet_03v3 ad=86.8f pd=0.92u as=86.8f ps=0.92u w=0.22u l=0.28u
X24 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD.t54 VDD.t53 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X25 a_8163_5223# CLK_div_10_mag_1.Q1.t5 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT VSS.t205 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X26 VSS CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_10610_4126# VSS.t68 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X27 a_9510_2450# CLK_div_10_mag_0.Q0 VSS.t276 VSS.t275 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X28 a_2076_256# CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS.t128 VSS.t127 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X29 VSS CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT a_4582_5223# VSS.t83 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X30 VSS CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_1559_4126# VSS.t93 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X31 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_10_mag_1.Q0.t4 VDD.t337 VDD.t336 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X32 CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS.t24 VSS.t23 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X33 VSS CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 a_3294_5223# VSS.t227 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X34 VSS VDD.t476 a_11334_4126# VSS.t109 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X35 VDD CLK_div_10_mag_1.Q0.t5 CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN VDD.t338 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X36 VSS CLK_div_10_mag_1.JK_FF_mag_0.J a_2283_4126# VSS.t196 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X37 VDD CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN CLK_div_10_mag_1.JK_FF_mag_0.J VDD.t43 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X38 a_788_212# CLK.t1 a_628_212# VSS.t297 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X39 a_3858_5223# CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 VSS.t209 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X40 VSS VDD.t477 a_5306_5223# VSS.t112 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X41 VSS CLK_div_10_mag_1.Q1.t6 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 VSS.t202 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X42 VDD CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD.t244 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X43 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD.t322 VDD.t321 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X44 a_9845_1309# CLK_div_10_mag_0.Q0 a_9685_1309# VSS.t274 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X45 VSS CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_995_4126# VSS.t44 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X46 VDD CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_10_mag_1.Q3 VDD.t365 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X47 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VDD.t132 VDD.t131 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X48 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VDD.t354 VDD.t353 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X49 a_4582_5223# RST.t1 a_4422_5223# VSS.t324 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X50 a_1559_4126# CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t33 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X51 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_10_mag_0.Q1 a_3805_212# VSS.t13 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X52 a_3294_5223# CLK_div_10_mag_1.Q2.t4 CLK_div_10_mag_1.JK_FF_mag_3.QB VSS.t103 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X53 VDD CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD.t261 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X54 CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_1.Q2.t5 VDD.t104 VDD.t103 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X55 a_2283_4126# CLK_div_10_mag_1.Q0.t6 a_2123_4126# VSS.t217 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X56 VDD RST.t2 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t323 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X57 CLK_div_10_mag_0.JK_FF_mag_0.J CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VSS.t118 VSS.t117 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X58 VDD CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t75 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X59 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t267 VDD.t266 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X60 a_9839_212# CLK_div_10_mag_0.Q0 a_9679_212# VSS.t273 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X61 a_9685_1309# CLK_div_10_mag_0.JK_FF_mag_0.J VSS.t299 VSS.t298 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X62 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.Q2 a_7574_2450# VSS.t290 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X63 VDD CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t218 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X64 VSS CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN CLK_div_10_mag_1.JK_FF_mag_0.J VSS.t27 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X65 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t215 VDD.t214 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X66 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_7546_212# VSS.t36 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X67 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT RST.t3 VDD.t460 VDD.t459 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X68 VSS CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 a_431_4126# VSS.t235 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X69 Vdiv100 CLK_div_10_mag_1.and2_mag_0.OUT VSS.t42 VSS.t41 nfet_03v3 ad=86.8f pd=0.92u as=86.8f ps=0.92u w=0.22u l=0.28u
X70 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_10_mag_0.Q0 VDD.t420 VDD.t419 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X71 a_995_4126# CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t92 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X72 VDD CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_10_mag_1.Q0.t0 VDD.t126 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X73 VDD CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_10_mag_1.nor_3_mag_0.IN3 VDD.t188 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X74 VSS CLK_div_10_mag_1.Q2.t6 a_3426_3029# VSS.t73 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X75 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.Q0 a_2640_256# VSS.t272 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X76 VDD CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_2.QB VDD.t20 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X77 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD.t177 VDD.t179 VDD.t178 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X78 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_3.QB a_6828_1309# VSS.t22 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X79 VSS CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_1565_5223# VSS.t159 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X80 a_7574_2450# CLK_div_10_mag_0.Q1 VSS.t12 VSS.t11 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X81 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_11127_256# VSS.t80 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X82 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t464 VDD.t463 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X83 VDD RST.t4 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD.t331 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X84 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_1.QB VDD.t235 VDD.t234 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X85 VDD CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t277 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X86 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.JK_FF_mag_1.QB VDD.t240 VDD.t239 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X87 a_1565_5223# RST.t5 a_1405_5223# VSS.t241 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X88 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_7956_1353# VSS.t72 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X89 VSS CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_9482_4126# VSS.t88 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X90 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t469 VDD.t468 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X91 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_10_mag_0.Q2 VDD.t448 VDD.t447 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X92 a_10563_212# RST.t6 a_10403_212# VSS.t316 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X93 a_8520_1353# CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VSS.t26 VSS.t25 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X94 a_5657_256# CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VSS.t135 VSS.t134 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X95 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_2076_256# VSS.t170 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X96 VDD CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT VDD.t28 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X97 VSS CLK_div_10_mag_1.Q3 Vdiv100.t1 VSS.t49 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X98 VDD CLK.t2 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t374 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X99 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_10_mag_0.Q2 VDD.t445 VDD.t444 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X100 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD.t248 VDD.t247 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X101 VDD CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT VDD.t343 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X102 VDD CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD.t442 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X103 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_10_mag_0.Q0 a_788_212# VSS.t271 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X104 a_9482_4126# CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_10_mag_1.Q0.t2 VSS.t142 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X105 VSS CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_10_mag_1.nor_3_mag_0.IN3 VSS.t98 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X106 a_3645_212# VDD.t478 VSS.t172 VSS.t171 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X107 VDD CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_10_mag_1.Q1.t0 VDD.t4 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X108 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.QB a_3811_1309# VSS.t212 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X109 a_4939_1353# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VSS.t64 VSS.t63 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X110 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD.t225 VDD.t224 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X111 VDD CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD.t241 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X112 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_10_mag_0.and2_mag_1.OUT VSS.t105 VSS.t104 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X113 VDD CLK_div_10_mag_1.CLK CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VDD.t273 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X114 a_1512_212# RST.t7 a_1352_212# VSS.t185 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X115 VDD CLK_div_10_mag_1.Q0.t7 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VDD.t136 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X116 VDD CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t84 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X117 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VDD.t402 VDD.t401 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X118 a_7439_5223# CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT VSS.t17 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X119 VDD CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t416 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X120 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t265 VDD.t264 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X121 CLK_div_10_mag_1.Q1 CLK_div_10_mag_1.JK_FF_mag_2.QB VDD.t292 VDD.t291 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X122 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_10_mag_1.CLK VDD.t431 VDD.t430 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X123 a_5140_4126# CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT VSS.t219 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X124 CLK_div_10_mag_1.CLK CLK_div_10_mag_0.Q3 a_11738_2752# VDD.t273 pfet_03v3 ad=1.06p pd=5.68u as=0.624p ps=2.92u w=2.4u l=0.28u
X125 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_4939_1353# VSS.t144 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X126 a_634_1309# VDD.t479 VSS.t174 VSS.t173 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X127 a_5503_1353# CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VSS.t211 VSS.t210 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X128 a_5093_256# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VSS.t224 VSS.t223 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X129 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VDD.t112 VDD.t111 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X130 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_10_mag_1.Q1.t7 VDD.t316 VDD.t315 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X131 VSS CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 a_6465_4126# VSS.t2 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X132 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.Q0 VDD.t415 VDD.t414 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X133 VDD CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT VDD.t285 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X134 VSS CLK_div_10_mag_1.nor_3_mag_0.IN3 Vdiv100.t3 VSS.t106 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X135 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_0.J VDD.t458 VDD.t457 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X136 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_10_mag_0.Q2 a_6822_212# VSS.t289 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X137 a_4369_212# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VSS.t146 VSS.t145 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X138 VSS CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_10046_4126# VSS.t59 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X139 VDD CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VDD.t236 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X140 a_10610_4126# CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t264 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X141 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.Q0 VSS.t270 VSS.t269 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X142 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_10409_1353# VSS.t54 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X143 VDD CLK_div_10_mag_1.JK_FF_mag_2.J.t2 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VDD.t382 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X144 a_10973_1353# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t164 VSS.t163 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X145 VDD CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VDD.t385 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X146 a_6465_4126# CLK_div_10_mag_1.JK_FF_mag_2.QB CLK_div_10_mag_1.Q1.t2 VSS.t191 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X147 a_11334_4126# CLK_div_10_mag_1.CLK a_11174_4126# VSS.t282 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X148 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_3.QB VDD.t38 VDD.t37 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X149 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_1358_1353# VSS.t126 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X150 a_1922_1353# CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t125 VSS.t124 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X151 a_5306_5223# CLK_div_10_mag_1.Q1.t8 a_5146_5223# VSS.t201 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X152 VDD VDD.t173 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VDD.t174 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X153 VDD VDD.t169 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VDD.t170 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X154 CLK_div_10_mag_1.Q3 CLK_div_10_mag_1.JK_FF_mag_2.J.t3 VDD.t427 VDD.t426 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X155 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_10563_212# VSS.t162 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X156 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.Q1 a_5657_256# VSS.t10 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X157 a_4422_5223# CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT VSS.t189 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X158 VDD CLK_div_10_mag_1.Q2.t7 CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN VDD.t105 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X159 a_11174_4126# CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VSS.t141 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X160 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD.t356 VDD.t355 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X161 VDD CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_1.and2_mag_0.OUT VDD.t249 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X162 VDD CLK_div_10_mag_0.JK_FF_mag_2.J.t4 CLK_div_10_mag_0.Q3 VDD.t362 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X163 a_1358_1353# CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS.t303 VSS.t302 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X164 VDD RST.t8 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VDD.t390 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X165 a_2123_4126# CLK_div_10_mag_1.JK_FF_mag_2.J.t4 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VSS.t277 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X166 VSS CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_10616_5223# VSS.t249 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X167 VDD CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.Q0 VDD.t231 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X168 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t281 VDD.t280 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X169 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_1922_1353# VSS.t169 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X170 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_10_mag_1.Q0.t8 VDD.t140 VDD.t139 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X171 CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VDD.t473 VDD.t472 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X172 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.Q1 VDD.t19 VDD.t18 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X173 VDD CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_3.QB VDD.t439 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X174 VSS VDD.t482 a_11340_5223# VSS.t175 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X175 VDD CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t116 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X176 VDD CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD.t61 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X177 a_431_4126# CLK_div_10_mag_1.JK_FF_mag_2.J.t5 CLK_div_10_mag_1.Q3 VSS.t257 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X178 VSS VDD.t483 a_2289_5223# VSS.t178 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X179 a_3426_3029# CLK_div_10_mag_1.Q1.t9 CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN VSS.t73 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X180 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_10_mag_0.Q1 a_8542_2450# VSS.t9 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X181 a_6828_1309# CLK_div_10_mag_0.Q1 a_6668_1309# VSS.t8 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X182 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t389 VDD.t388 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X183 CLK_div_10_mag_0.JK_FF_mag_2.J CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t361 VDD.t360 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X184 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_10_mag_0.Q3 VDD.t272 VDD.t271 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X185 VDD CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t46 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X186 VSS CLK_div_10_mag_1.Q1.t10 a_4394_3029# VSS.t73 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X187 VSS CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_1.and2_mag_0.OUT VSS.t147 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X188 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.QB VDD.t330 VDD.t329 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X189 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD.t120 VDD.t119 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X190 a_10046_4126# CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t323 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X191 a_2289_5223# CLK_div_10_mag_1.Q0.t9 a_2129_5223# VSS.t96 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X192 a_6668_1309# VDD.t484 VSS.t182 VSS.t181 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X193 a_8674_256# CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VSS.t133 VSS.t132 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X194 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_5093_256# VSS.t143 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X195 a_1405_5223# CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VSS.t43 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X196 a_4529_212# RST.t9 a_4369_212# VSS.t97 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X197 a_4394_3029# CLK_div_10_mag_1.Q2.t8 CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN VSS.t73 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X198 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK.t3 VDD.t377 VDD.t72 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X199 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t74 VDD.t73 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X200 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t435 VDD.t434 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X201 VSS CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_841_5223# VSS.t30 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X202 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t166 VDD.t168 VDD.t167 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X203 VDD CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t398 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X204 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 VDD.t3 VDD.t2 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X205 CLK_div_10_mag_0.JK_FF_mag_0.J CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD.t206 VDD.t205 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X206 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.Q0 VDD.t413 VDD.t412 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X207 VDD CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 VDD.t255 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X208 a_8110_256# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VSS.t78 VSS.t77 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X209 a_3811_1309# CLK_div_10_mag_0.Q0 a_3651_1309# VSS.t268 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X210 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_10_mag_0.Q3 a_9839_212# VSS.t168 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X211 VDD CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_10_mag_1.JK_FF_mag_1.QB VDD.t449 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X212 CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VDD.t471 VDD.t470 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X213 a_7386_212# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VSS.t82 VSS.t81 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X214 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t163 VDD.t165 VDD.t164 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X215 VDD CLK_div_10_mag_1.JK_FF_mag_2.J.t6 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT VDD.t395 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X216 VDD CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 VDD.t25 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X217 VDD CLK_div_10_mag_1.Q0.t10 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 VDD.t368 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X218 VSS CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_9892_5223# VSS.t261 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X219 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT VDD.t59 VDD.t58 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X220 a_7029_4126# CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 VSS.t1 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X221 VDD CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD.t409 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X222 a_11738_2752# CLK_div_10_mag_0.and2_mag_0.OUT a_11578_2752# VDD.t91 pfet_03v3 ad=0.624p pd=2.92u as=0.624p ps=2.92u w=2.4u l=0.28u
X223 VSS CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT a_7593_4126# VSS.t153 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X224 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t213 VDD.t212 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X225 VDD CLK_div_10_mag_1.Q2.t9 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT VDD.t202 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X226 VDD CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t436 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X227 VSS CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_9328_5223# VSS.t291 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X228 a_9892_5223# CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t322 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X229 VDD CLK_div_10_mag_0.Q3 CLK_div_10_mag_0.JK_FF_mag_2.J.t0 VDD.t268 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X230 VDD CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 VDD.t55 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X231 VSS CLK_div_10_mag_1.JK_FF_mag_2.J.t7 a_8317_4126# VSS.t258 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X232 VDD CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_10_mag_1.Q2.t0 VDD.t252 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X233 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 VDD.t318 VDD.t317 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X234 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.Q0 VSS.t267 VSS.t266 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X235 VDD RST.t10 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VDD.t141 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X236 CLK_div_10_mag_0.Q3 CLK_div_10_mag_0.JK_FF_mag_2.J.t5 a_11537_1353# VSS.t232 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X237 VSS CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 a_7029_4126# VSS.t14 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X238 a_11578_2752# CLK_div_10_mag_0.nor_3_mag_0.IN3 VDD.t381 VDD.t380 pfet_03v3 ad=0.624p pd=2.92u as=1.06p ps=5.68u w=2.4u l=0.28u
X239 a_10409_1353# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS.t184 VSS.t183 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X240 a_7593_4126# CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 VSS.t40 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X241 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.Q1 VDD.t17 VDD.t16 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X242 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.QB a_2486_1353# VSS.t140 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X243 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD.t160 VDD.t162 VDD.t161 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X244 VDD CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT VDD.t465 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X245 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT RST.t11 VDD.t145 VDD.t144 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X246 VDD CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD.t13 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X247 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.Q2 a_8674_256# VSS.t288 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X248 a_628_212# VDD.t485 VSS.t305 VSS.t304 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X249 VDD CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_10_mag_1.JK_FF_mag_2.QB VDD.t78 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X250 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_10973_1353# VSS.t79 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X251 a_5146_5223# CLK_div_10_mag_1.Q2.t10 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT VSS.t116 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X252 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 VDD.t1 VDD.t0 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X253 VDD VDD.t156 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT VDD.t157 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X254 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_10_mag_1.CLK VDD.t429 VDD.t428 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X255 VDD VDD.t152 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT VDD.t153 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X256 VDD CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD.t108 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X257 VDD CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 VDD.t282 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X258 VDD CLK_div_10_mag_1.Q1.t11 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 VDD.t312 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X259 VDD CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VDD.t81 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X260 VSS CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 a_3448_4126# VSS.t150 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X261 VDD CLK_div_10_mag_1.and2_mag_1.OUT CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VDD.t31 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X262 CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN CLK_div_10_mag_1.Q1.t12 VDD.t311 VDD.t310 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X263 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD.t52 VDD.t51 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X264 a_2486_1353# CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t253 VSS.t252 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X265 a_11691_256# CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t231 VSS.t230 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X266 a_3805_212# CLK_div_10_mag_0.Q0 a_3645_212# VSS.t265 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X267 VSS CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT a_6875_5223# VSS.t37 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X268 a_4012_4126# CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 VSS.t208 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X269 VSS CLK_div_10_mag_1.CLK CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VSS.t279 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X270 VDD CLK_div_10_mag_1.nor_3_mag_0.IN3 a_390_2335# VDD.t197 pfet_03v3 ad=1.06p pd=5.68u as=0.624p ps=2.92u w=2.4u l=0.28u
X271 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD.t149 VDD.t151 VDD.t150 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X272 VSS CLK_div_10_mag_1.Q0.t11 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VSS.t238 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X273 VDD CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.Q2 VDD.t34 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X274 CLK_div_10_mag_0.Q3 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t456 VDD.t455 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X275 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_1512_212# VSS.t123 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X276 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t349 VDD.t348 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X277 a_10616_5223# RST.t12 a_10456_5223# VSS.t192 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X278 VDD CLK_div_10_mag_1.Q0.t12 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VDD.t371 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X279 VDD CLK_div_10_mag_1.Q1.t13 CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN VDD.t307 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X280 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD.t296 VDD.t295 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X281 VSS CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT a_7599_5223# VSS.t317 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X282 VDD CLK_div_10_mag_1.Q3 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VDD.t69 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X283 CLK_div_10_mag_1.CLK CLK_div_10_mag_0.Q3 VSS.t167 VSS.t166 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X284 VSS CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 a_6311_5223# VSS.t55 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X285 a_11340_5223# CLK_div_10_mag_1.CLK a_11180_5223# VSS.t278 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X286 a_7546_212# RST.t13 a_7386_212# VSS.t193 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X287 a_6875_5223# CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 VSS.t0 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X288 VSS VDD.t488 a_8323_5223# VSS.t306 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X289 VSS VDD.t489 a_5300_4126# VSS.t309 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X290 a_390_2335# CLK_div_10_mag_1.and2_mag_0.OUT a_230_2335# VDD.t60 pfet_03v3 ad=0.624p pd=2.92u as=0.624p ps=2.92u w=2.4u l=0.28u
X291 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.Q1 VSS.t7 VSS.t6 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X292 VSS CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 a_4012_4126# VSS.t186 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X293 a_8542_2450# CLK_div_10_mag_0.Q2 VSS.t287 VSS.t286 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X294 a_11127_256# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS.t53 VSS.t52 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X295 a_6662_212# VDD.t490 VSS.t313 VSS.t312 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X296 a_2640_256# CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t284 VSS.t283 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X297 a_10456_5223# CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VSS.t58 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X298 VDD CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_10_mag_1.JK_FF_mag_2.J.t1 VDD.t221 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X299 CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_1.Q2.t11 VDD.t201 VDD.t200 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X300 CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VDD.t40 VDD.t39 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X301 VDD CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD.t100 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X302 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VDD.t130 VDD.t129 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X303 VDD CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VDD.t406 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X304 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t462 VDD.t461 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X305 a_11180_5223# CLK_div_10_mag_1.Q0.t13 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VSS.t254 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X306 VDD CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_1.and2_mag_1.OUT VDD.t228 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X307 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.Q2 a_9510_2450# VSS.t285 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X308 a_2129_5223# CLK_div_10_mag_1.Q3 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VSS.t48 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X309 VSS CLK_div_10_mag_1.and2_mag_1.OUT CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS.t18 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X310 VDD CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD.t350 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X311 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.Q3 VDD.t68 VDD.t67 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X312 a_10403_212# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS.t221 VSS.t220 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X313 VDD CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.Q1 VDD.t326 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X314 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.J.t6 a_9845_1309# VSS.t233 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X315 VSS CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_277_5223# VSS.t129 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X316 a_841_5223# CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t91 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X317 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VDD.t125 VDD.t124 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X318 VDD CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD.t10 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X319 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS.t321 VSS.t320 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X320 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK.t4 VSS.t243 VSS.t242 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X321 VSS CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_1.and2_mag_1.OUT VSS.t136 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X322 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD.t88 VDD.t87 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X323 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD.t217 VDD.t216 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X324 VSS CLK_div_10_mag_1.Q0.t14 a_2458_3029# VSS.t115 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X325 a_3651_1309# CLK_div_10_mag_0.JK_FF_mag_2.J.t7 VSS.t102 VSS.t101 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X326 a_277_5223# CLK_div_10_mag_1.Q3 CLK_div_10_mag_1.JK_FF_mag_2.J VSS.t47 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X327 CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_10_mag_1.Q0.t15 VDD.t394 VDD.t393 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X328 CLK_div_10_mag_0.JK_FF_mag_2.J CLK_div_10_mag_0.Q3 a_11691_256# VSS.t165 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X329 a_1352_212# CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS.t301 VSS.t300 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X330 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_10_mag_1.Q0.t16 VDD.t335 VDD.t334 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X331 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t146 VDD.t148 VDD.t147 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X332 a_2458_3029# CLK_div_10_mag_1.Q2.t12 CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN VSS.t115 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X333 CLK_div_10_mag_1.CLK CLK_div_10_mag_0.nor_3_mag_0.IN3 VSS.t248 VSS.t247 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X334 VDD CLK_div_10_mag_1.JK_FF_mag_2.QB CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT VDD.t288 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X335 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_7392_1353# VSS.t76 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X336 VDD CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 VDD.t258 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X337 a_6822_212# CLK_div_10_mag_0.Q1 a_6662_212# VSS.t5 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X338 a_9328_5223# CLK_div_10_mag_1.Q0.t17 CLK_div_10_mag_1.JK_FF_mag_1.QB VSS.t214 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X339 a_7956_1353# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VSS.t35 VSS.t34 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X340 a_8317_4126# CLK_div_10_mag_1.Q0.t18 a_8157_4126# VSS.t215 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X341 a_11537_1353# CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t295 VSS.t294 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X342 VDD CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD.t7 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X343 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_4529_212# VSS.t62 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X344 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_3.QB a_8520_1353# VSS.t21 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X345 a_7392_1353# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VSS.t195 VSS.t194 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X346 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT RST.t14 VDD.t294 VDD.t293 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X347 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT VDD.t211 VDD.t210 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X348 VDD CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t113 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X349 VDD CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.QB VDD.t403 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X350 CLK_div_10_mag_1.JK_FF_mag_2.QB CLK_div_10_mag_1.Q1.t14 VDD.t306 VDD.t305 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X351 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_10_mag_0.and2_mag_1.OUT VDD.t196 VDD.t195 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X352 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_10_mag_1.Q0.t19 VDD.t379 VDD.t378 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X353 a_8157_4126# CLK_div_10_mag_1.JK_FF_mag_2.QB CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT VSS.t190 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X354 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_10_mag_1.Q1.t15 VDD.t304 VDD.t303 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X355 VSS CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT a_4576_4126# VSS.t156 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X356 a_9679_212# VDD.t491 VSS.t315 VSS.t314 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X357 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_8110_256# VSS.t71 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X358 a_3448_4126# CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_10_mag_1.Q2.t1 VSS.t218 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X359 VSS CLK_div_10_mag_1.Q0.t20 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 VSS.t244 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X360 VDD CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD.t97 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X361 VDD CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 VDD.t207 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X362 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD.t42 VDD.t41 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X363 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_1.QB a_794_1309# VSS.t139 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X364 VDD CLK.t5 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t452 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X365 VDD CLK_div_10_mag_1.Q1.t16 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT VDD.t300 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X366 VDD CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t94 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X367 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_4375_1353# VSS.t222 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X368 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD.t227 VDD.t226 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X369 VDD CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t274 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X370 a_7599_5223# RST.t15 a_7439_5223# VSS.t234 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X371 VDD CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT VDD.t121 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X372 a_4576_4126# CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 VSS.t119 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X373 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VSS.t226 VSS.t225 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X374 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.J.t8 VDD.t192 VDD.t191 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
R0 CLK_div_10_mag_1.Q1.n17 CLK_div_10_mag_1.Q1.t4 36.935
R1 CLK_div_10_mag_1.Q1.n18 CLK_div_10_mag_1.Q1.t8 36.935
R2 CLK_div_10_mag_1.Q1.n12 CLK_div_10_mag_1.Q1.t5 36.935
R3 CLK_div_10_mag_1.Q1.n19 CLK_div_10_mag_1.Q1.t9 31.4332
R4 CLK_div_10_mag_1.Q1.n14 CLK_div_10_mag_1.Q1.t3 31.4332
R5 CLK_div_10_mag_1.Q1.n20 CLK_div_10_mag_1.Q1.t13 30.9379
R6 CLK_div_10_mag_1.Q1.n22 CLK_div_10_mag_1.Q1.t11 25.4744
R7 CLK_div_10_mag_1.Q1.n20 CLK_div_10_mag_1.Q1.t10 21.6422
R8 CLK_div_10_mag_1.Q1.n17 CLK_div_10_mag_1.Q1.t15 18.1962
R9 CLK_div_10_mag_1.Q1.n18 CLK_div_10_mag_1.Q1.t7 18.1962
R10 CLK_div_10_mag_1.Q1.n12 CLK_div_10_mag_1.Q1.t16 18.1962
R11 CLK_div_10_mag_1.Q1.n19 CLK_div_10_mag_1.Q1.t12 15.3826
R12 CLK_div_10_mag_1.Q1.n14 CLK_div_10_mag_1.Q1.t14 15.3826
R13 CLK_div_10_mag_1.Q1.n22 CLK_div_10_mag_1.Q1.t6 14.1417
R14 CLK_div_10_mag_1.Q1.n11 CLK_div_10_mag_1.Q1.t2 7.09905
R15 CLK_div_10_mag_1.Q1.n15 CLK_div_10_mag_1.Q1.n14 6.86029
R16 CLK_div_10_mag_1.Q1.n16 CLK_div_10_mag_1.Q1.n13 5.01077
R17 CLK_div_10_mag_1.Q1.n2 CLK_div_10_mag_1.Q1.n4 0.0219501
R18 CLK_div_10_mag_1.Q1.n1 CLK_div_10_mag_1.Q1.n0 0.0360559
R19 CLK_div_10_mag_1.Q1.n19 CLK_div_10_mag_1.Q1 5.69501
R20 CLK_div_10_mag_1.Q1.n4 CLK_div_10_mag_1.Q1.n1 2.23369
R21 CLK_div_10_mag_1.Q1.n2 CLK_div_10_mag_1.Q1.n0 1.11499
R22 CLK_div_10_mag_1.Q1.n23 CLK_div_10_mag_1.Q1.n8 2.2429
R23 CLK_div_10_mag_1.Q1.n8 CLK_div_10_mag_1.Q1.n7 0.0171915
R24 CLK_div_10_mag_1.Q1.n11 CLK_div_10_mag_1.Q1.n10 3.25053
R25 CLK_div_10_mag_1.Q1.n10 CLK_div_10_mag_1.Q1.t0 2.2755
R26 CLK_div_10_mag_1.Q1.n10 CLK_div_10_mag_1.Q1.n9 2.2755
R27 CLK_div_10_mag_1.Q1.n25 CLK_div_10_mag_1.Q1.n24 2.2505
R28 CLK_div_10_mag_1.Q1.n7 CLK_div_10_mag_1.Q1.n6 2.24196
R29 CLK_div_10_mag_1.Q1.n13 CLK_div_10_mag_1.Q1.n12 2.13459
R30 CLK_div_10_mag_1.Q1.n3 CLK_div_10_mag_1.Q1.n20 2.13074
R31 CLK_div_10_mag_1.Q1.n4 CLK_div_10_mag_1.Q1.n17 2.12093
R32 CLK_div_10_mag_1.Q1.n1 CLK_div_10_mag_1.Q1.n5 2.64237
R33 CLK_div_10_mag_1.Q1.n0 CLK_div_10_mag_1.Q1.n21 4.95192
R34 CLK_div_10_mag_1.Q1.n21 CLK_div_10_mag_1.Q1 4.19069
R35 CLK_div_10_mag_1.Q1.n24 CLK_div_10_mag_1.Q1.n16 1.52773
R36 CLK_div_10_mag_1.Q1.n18 CLK_div_10_mag_1.Q1.n5 2.13281
R37 CLK_div_10_mag_1.Q1.n7 CLK_div_10_mag_1.Q1.n22 1.42118
R38 CLK_div_10_mag_1.Q1.n16 CLK_div_10_mag_1.Q1.n15 1.12067
R39 CLK_div_10_mag_1.Q1.n6 CLK_div_10_mag_1.Q1.n0 0.960138
R40 CLK_div_10_mag_1.Q1 CLK_div_10_mag_1.Q1.n23 0.646487
R41 CLK_div_10_mag_1.Q1.n8 CLK_div_10_mag_1.Q1 0.187192
R42 CLK_div_10_mag_1.Q1.n25 CLK_div_10_mag_1.Q1.n11 0.0905
R43 CLK_div_10_mag_1.Q1.n15 CLK_div_10_mag_1.Q1 0.0857632
R44 CLK_div_10_mag_1.Q1 CLK_div_10_mag_1.Q1.n25 0.0834687
R45 CLK_div_10_mag_1.Q1.n13 CLK_div_10_mag_1.Q1 0.0800273
R46 CLK_div_10_mag_1.Q1.n3 CLK_div_10_mag_1.Q1 0.0980715
R47 CLK_div_10_mag_1.Q1.n2 CLK_div_10_mag_1.Q1 0.0672526
R48 CLK_div_10_mag_1.Q1.n5 CLK_div_10_mag_1.Q1 0.0771461
R49 CLK_div_10_mag_1.Q1.n24 CLK_div_10_mag_1.Q1 0.0322045
R50 CLK_div_10_mag_1.Q1.n23 CLK_div_10_mag_1.Q1.n6 0.0238218
R51 CLK_div_10_mag_1.Q1.n21 CLK_div_10_mag_1.Q1.n3 2.08419
R52 VSS.n245 VSS.n232 36515.7
R53 VSS.n349 VSS.n348 36280.3
R54 VSS.n227 VSS.n226 18801.2
R55 VSS.n258 VSS.n228 18801.2
R56 VSS.t47 VSS.n4 12177.1
R57 VSS.n78 VSS.n77 9589.42
R58 VSS.n266 VSS.n265 9584.01
R59 VSS.n348 VSS.t304 6168.75
R60 VSS.n289 VSS.n288 5257.24
R61 VSS.n349 VSS.n4 5257.24
R62 VSS.n178 VSS.n177 3893.61
R63 VSS.n305 VSS.n304 3893.61
R64 VSS.n15 VSS.t23 3606.54
R65 VSS.t98 VSS.n65 3606.54
R66 VSS.n14 VSS.t247 3112.87
R67 VSS.n67 VSS.t106 3112.87
R68 VSS.n228 VSS.n36 3086.35
R69 VSS.t225 VSS.t104 3055.32
R70 VSS.t214 VSS.n149 2628.58
R71 VSS.n166 VSS.t207 2628.58
R72 VSS.n177 VSS.t103 2628.58
R73 VSS.t314 VSS.n305 2628.58
R74 VSS.t312 VSS.n318 2628.58
R75 VSS.t171 VSS.n331 2628.58
R76 VSS.n149 VSS.t306 2622.37
R77 VSS.t112 VSS.n166 2622.37
R78 VSS.n305 VSS.t288 2622.37
R79 VSS.n318 VSS.t10 2622.37
R80 VSS.n331 VSS.t272 2622.37
R81 VSS.t249 VSS.t254 2510.52
R82 VSS.t291 VSS.t322 2510.52
R83 VSS.t317 VSS.t205 2510.52
R84 VSS.t0 VSS.t55 2510.52
R85 VSS.t83 VSS.t116 2510.52
R86 VSS.t227 VSS.t209 2510.52
R87 VSS.t159 VSS.t48 2510.52
R88 VSS.t129 VSS.t91 2510.52
R89 VSS.t80 VSS.t230 2510.52
R90 VSS.t168 VSS.t220 2510.52
R91 VSS.t71 VSS.t132 2510.52
R92 VSS.t289 VSS.t81 2510.52
R93 VSS.t143 VSS.t134 2510.52
R94 VSS.t13 VSS.t145 2510.52
R95 VSS.t170 VSS.t283 2510.52
R96 VSS.t300 VSS.t271 2510.52
R97 VSS.t320 VSS.t286 2307.56
R98 VSS.t279 VSS.t109 2307.56
R99 VSS.t141 VSS.t68 2307.56
R100 VSS.t264 VSS.t59 2307.56
R101 VSS.t323 VSS.t88 2307.56
R102 VSS.t244 VSS.t258 2307.56
R103 VSS.t190 VSS.t153 2307.56
R104 VSS.t40 VSS.t14 2307.56
R105 VSS.t1 VSS.t2 2307.56
R106 VSS.t156 VSS.t219 2307.56
R107 VSS.t186 VSS.t119 2307.56
R108 VSS.t150 VSS.t208 2307.56
R109 VSS.t238 VSS.t196 2307.56
R110 VSS.t277 VSS.t93 2307.56
R111 VSS.t33 VSS.t44 2307.56
R112 VSS.t92 VSS.t235 2307.56
R113 VSS.t294 VSS.t79 2307.56
R114 VSS.t54 VSS.t163 2307.56
R115 VSS.t183 VSS.t233 2307.56
R116 VSS.t266 VSS.t298 2307.56
R117 VSS.t25 VSS.t72 2307.56
R118 VSS.t34 VSS.t76 2307.56
R119 VSS.t194 VSS.t22 2307.56
R120 VSS.t181 VSS.t6 2307.56
R121 VSS.t144 VSS.t210 2307.56
R122 VSS.t222 VSS.t63 2307.56
R123 VSS.t212 VSS.t86 2307.56
R124 VSS.t101 VSS.t269 2307.56
R125 VSS.t252 VSS.t169 2307.56
R126 VSS.t124 VSS.t126 2307.56
R127 VSS.t302 VSS.t139 2307.56
R128 VSS.t173 VSS.t242 2307.56
R129 VSS.t257 VSS.n4 2084.8
R130 VSS.t232 VSS.n289 2084.8
R131 VSS.t18 VSS.n47 1878.69
R132 VSS.t142 VSS.n131 1719.24
R133 VSS.n226 VSS.t191 1719.24
R134 VSS.t218 VSS.n78 1719.24
R135 VSS.n265 VSS.t21 1713.53
R136 VSS.n258 VSS.t213 1713.53
R137 VSS.n245 VSS.t140 1713.53
R138 VSS.n131 VSS.n130 1565.03
R139 VSS.n226 VSS.n225 1565.03
R140 VSS.n259 VSS.n258 1565.03
R141 VSS.n246 VSS.n245 1565.03
R142 VSS.t65 VSS.t166 1151.9
R143 VSS.t41 VSS.t49 1151.9
R144 VSS.t49 VSS.n349 1007.91
R145 VSS.t254 VSS.t278 994.264
R146 VSS.t192 VSS.t58 994.264
R147 VSS.t205 VSS.t216 994.264
R148 VSS.t234 VSS.t17 994.264
R149 VSS.t116 VSS.t201 994.264
R150 VSS.t324 VSS.t189 994.264
R151 VSS.t48 VSS.t96 994.264
R152 VSS.t241 VSS.t43 994.264
R153 VSS.t316 VSS.t162 994.264
R154 VSS.t273 VSS.t168 994.264
R155 VSS.t193 VSS.t36 994.264
R156 VSS.t5 VSS.t289 994.264
R157 VSS.t97 VSS.t62 994.264
R158 VSS.t265 VSS.t13 994.264
R159 VSS.t185 VSS.t123 994.264
R160 VSS.t271 VSS.t297 994.264
R161 VSS.t282 VSS.t141 913.885
R162 VSS.t215 VSS.t190 913.885
R163 VSS.t219 VSS.t206 913.885
R164 VSS.t217 VSS.t277 913.885
R165 VSS.t233 VSS.t274 913.885
R166 VSS.t22 VSS.t8 913.885
R167 VSS.t268 VSS.t212 913.885
R168 VSS.t139 VSS.t296 913.885
R169 VSS.n46 VSS.t27 838.187
R170 VSS.n267 VSS.t117 838.187
R171 VSS.n13 VSS.t65 671.942
R172 VSS.n350 VSS.t41 671.942
R173 VSS.t278 VSS.n143 596.558
R174 VSS.n144 VSS.t192 596.558
R175 VSS.t322 VSS.n148 596.558
R176 VSS.n150 VSS.t214 596.558
R177 VSS.t216 VSS.n157 596.558
R178 VSS.n158 VSS.t234 596.558
R179 VSS.n161 VSS.t0 596.558
R180 VSS.t207 VSS.n165 596.558
R181 VSS.t201 VSS.n167 596.558
R182 VSS.n169 VSS.t324 596.558
R183 VSS.t209 VSS.n171 596.558
R184 VSS.t103 VSS.n173 596.558
R185 VSS.t96 VSS.n197 596.558
R186 VSS.n199 VSS.t241 596.558
R187 VSS.t91 VSS.n201 596.558
R188 VSS.n203 VSS.t47 596.558
R189 VSS.n282 VSS.t165 596.558
R190 VSS.n283 VSS.t80 596.558
R191 VSS.n287 VSS.t316 596.558
R192 VSS.n306 VSS.t273 596.558
R193 VSS.n312 VSS.t288 596.558
R194 VSS.n313 VSS.t71 596.558
R195 VSS.n317 VSS.t193 596.558
R196 VSS.n319 VSS.t5 596.558
R197 VSS.n325 VSS.t10 596.558
R198 VSS.n326 VSS.t143 596.558
R199 VSS.n330 VSS.t97 596.558
R200 VSS.n332 VSS.t265 596.558
R201 VSS.n338 VSS.t272 596.558
R202 VSS.n339 VSS.t170 596.558
R203 VSS.n342 VSS.t185 596.558
R204 VSS.n347 VSS.t297 596.558
R205 VSS.n18 VSS.t9 548.331
R206 VSS.n20 VSS.t290 548.331
R207 VSS.n17 VSS.t285 548.331
R208 VSS.n135 VSS.t282 548.331
R209 VSS.n134 VSS.t264 548.331
R210 VSS.n133 VSS.t323 548.331
R211 VSS.n132 VSS.t142 548.331
R212 VSS.n128 VSS.t215 548.331
R213 VSS.n127 VSS.t40 548.331
R214 VSS.n126 VSS.t1 548.331
R215 VSS.n125 VSS.t191 548.331
R216 VSS.t206 VSS.n39 548.331
R217 VSS.t119 VSS.n41 548.331
R218 VSS.t208 VSS.n43 548.331
R219 VSS.n79 VSS.t218 548.331
R220 VSS.n192 VSS.t217 548.331
R221 VSS.n191 VSS.t33 548.331
R222 VSS.n190 VSS.t92 548.331
R223 VSS.n189 VSS.t257 548.331
R224 VSS.n290 VSS.t232 548.331
R225 VSS.n295 VSS.t79 548.331
R226 VSS.n296 VSS.t54 548.331
R227 VSS.n301 VSS.t274 548.331
R228 VSS.t21 VSS.n264 548.331
R229 VSS.t72 VSS.n263 548.331
R230 VSS.t76 VSS.n262 548.331
R231 VSS.t8 VSS.n261 548.331
R232 VSS.t213 VSS.n257 548.331
R233 VSS.n229 VSS.t144 548.331
R234 VSS.n230 VSS.t222 548.331
R235 VSS.n248 VSS.t268 548.331
R236 VSS.t140 VSS.n244 548.331
R237 VSS.t169 VSS.n243 548.331
R238 VSS.t126 VSS.n242 548.331
R239 VSS.t296 VSS.n241 548.331
R240 VSS.n228 VSS.n227 508.851
R241 VSS.t247 VSS.n13 479.959
R242 VSS.n350 VSS.t106 479.959
R243 VSS.t115 VSS.t136 398.623
R244 VSS.n143 VSS.t175 397.707
R245 VSS.n144 VSS.t249 397.707
R246 VSS.n148 VSS.t261 397.707
R247 VSS.n150 VSS.t291 397.707
R248 VSS.n157 VSS.t306 397.707
R249 VSS.n158 VSS.t317 397.707
R250 VSS.n161 VSS.t37 397.707
R251 VSS.n165 VSS.t55 397.707
R252 VSS.n167 VSS.t112 397.707
R253 VSS.n169 VSS.t83 397.707
R254 VSS.n171 VSS.t120 397.707
R255 VSS.n173 VSS.t227 397.707
R256 VSS.n197 VSS.t178 397.707
R257 VSS.n199 VSS.t159 397.707
R258 VSS.n201 VSS.t30 397.707
R259 VSS.n203 VSS.t129 397.707
R260 VSS.t230 VSS.n282 397.707
R261 VSS.n283 VSS.t52 397.707
R262 VSS.t220 VSS.n287 397.707
R263 VSS.n306 VSS.t314 397.707
R264 VSS.t132 VSS.n312 397.707
R265 VSS.n313 VSS.t77 397.707
R266 VSS.t81 VSS.n317 397.707
R267 VSS.n319 VSS.t312 397.707
R268 VSS.t134 VSS.n325 397.707
R269 VSS.n326 VSS.t223 397.707
R270 VSS.t145 VSS.n330 397.707
R271 VSS.n332 VSS.t171 397.707
R272 VSS.t283 VSS.n338 397.707
R273 VSS.n339 VSS.t127 397.707
R274 VSS.n342 VSS.t300 397.707
R275 VSS.t304 VSS.n347 397.707
R276 VSS.t286 VSS.n18 365.555
R277 VSS.n20 VSS.t11 365.555
R278 VSS.t275 VSS.n17 365.555
R279 VSS.t109 VSS.n135 365.555
R280 VSS.t68 VSS.n134 365.555
R281 VSS.t59 VSS.n133 365.555
R282 VSS.t88 VSS.n132 365.555
R283 VSS.t258 VSS.n128 365.555
R284 VSS.t153 VSS.n127 365.555
R285 VSS.t14 VSS.n126 365.555
R286 VSS.t2 VSS.n125 365.555
R287 VSS.n39 VSS.t309 365.555
R288 VSS.n41 VSS.t156 365.555
R289 VSS.n43 VSS.t186 365.555
R290 VSS.n79 VSS.t150 365.555
R291 VSS.t196 VSS.n192 365.555
R292 VSS.t93 VSS.n191 365.555
R293 VSS.t44 VSS.n190 365.555
R294 VSS.t235 VSS.n189 365.555
R295 VSS.n290 VSS.t294 365.555
R296 VSS.t163 VSS.n295 365.555
R297 VSS.n296 VSS.t183 365.555
R298 VSS.t298 VSS.n301 365.555
R299 VSS.n264 VSS.t25 365.555
R300 VSS.n263 VSS.t34 365.555
R301 VSS.n262 VSS.t194 365.555
R302 VSS.n261 VSS.t181 365.555
R303 VSS.n257 VSS.t210 365.555
R304 VSS.t63 VSS.n229 365.555
R305 VSS.t86 VSS.n230 365.555
R306 VSS.n248 VSS.t101 365.555
R307 VSS.n244 VSS.t252 365.555
R308 VSS.n243 VSS.t124 365.555
R309 VSS.n242 VSS.t302 365.555
R310 VSS.n241 VSS.t173 365.555
R311 VSS.n348 VSS.n1 348.418
R312 VSS.n136 VSS.n100 342.707
R313 VSS.n76 VSS.t115 231.852
R314 VSS.t73 VSS.t147 211.208
R315 VSS.n77 VSS.n47 195.244
R316 VSS.n266 VSS.t275 165.642
R317 VSS.t23 VSS.n14 150.845
R318 VSS.t104 VSS.n15 150.845
R319 VSS.n65 VSS.t18 150.845
R320 VSS.n67 VSS.t98 150.845
R321 VSS.n45 VSS.t73 122.846
R322 VSS.n304 VSS.n303 119.948
R323 VSS.n260 VSS.n259 119.948
R324 VSS.n247 VSS.n246 119.948
R325 VSS.n130 VSS.n129 114.236
R326 VSS.n225 VSS.n224 114.236
R327 VSS.n193 VSS.n178 114.236
R328 VSS.n19 VSS.t320 34.2711
R329 VSS.n16 VSS.t225 34.2711
R330 VSS.n136 VSS.t279 34.2711
R331 VSS.n129 VSS.t244 34.2711
R332 VSS.n224 VSS.t202 34.2711
R333 VSS.n193 VSS.t238 34.2711
R334 VSS.n303 VSS.t266 34.2711
R335 VSS.t6 VSS.n260 34.2711
R336 VSS.t269 VSS.n247 34.2711
R337 VSS.t242 VSS.n1 34.2711
R338 VSS.n267 VSS.n266 27.0388
R339 VSS.n77 VSS.n46 21.6311
R340 VSS.n77 VSS.n76 16.2708
R341 VSS.n277 VSS.t248 9.37686
R342 VSS.n69 VSS.n68 9.37686
R343 VSS.n231 VSS.t270 9.3736
R344 VSS.n35 VSS.t7 9.3736
R345 VSS.n302 VSS.t267 9.3736
R346 VSS.n194 VSS.n176 9.37275
R347 VSS.n223 VSS.n37 9.37275
R348 VSS.n112 VSS.n111 9.37275
R349 VSS.n137 VSS.n99 9.37275
R350 VSS.n271 VSS.t226 9.30652
R351 VSS.n26 VSS.t118 9.30652
R352 VSS.n22 VSS.t321 9.30652
R353 VSS.n64 VSS.n48 9.30652
R354 VSS.n60 VSS.n50 9.30652
R355 VSS.n56 VSS.n52 9.30652
R356 VSS.n354 VSS.t243 9.30652
R357 VSS.n275 VSS.t24 9.30518
R358 VSS.n71 VSS.n66 9.30518
R359 VSS.n273 VSS.t105 9.25414
R360 VSS.n74 VSS.n73 9.25414
R361 VSS.n77 VSS.n45 8.62119
R362 VSS VSS.n51 7.30633
R363 VSS VSS.t12 7.30633
R364 VSS.n280 VSS.t231 7.19156
R365 VSS.n285 VSS.t53 7.19156
R366 VSS.n310 VSS.t133 7.19156
R367 VSS.n315 VSS.t78 7.19156
R368 VSS.n323 VSS.t135 7.19156
R369 VSS.n328 VSS.t224 7.19156
R370 VSS.n28 VSS.t26 7.19156
R371 VSS.n30 VSS.t35 7.19156
R372 VSS.n32 VSS.t195 7.19156
R373 VSS.n292 VSS.t295 7.19156
R374 VSS.n293 VSS.t164 7.19156
R375 VSS.n298 VSS.t184 7.19156
R376 VSS.n234 VSS.t253 7.19156
R377 VSS.n236 VSS.t125 7.19156
R378 VSS.n238 VSS.t303 7.19156
R379 VSS.n205 VSS.n202 7.19156
R380 VSS.n207 VSS.n200 7.19156
R381 VSS.n187 VSS.n186 7.19156
R382 VSS.n184 VSS.n183 7.19156
R383 VSS.n181 VSS.n180 7.19156
R384 VSS.n214 VSS.n172 7.19156
R385 VSS.n216 VSS.n170 7.19156
R386 VSS.n81 VSS.n44 7.19156
R387 VSS.n83 VSS.n42 7.19156
R388 VSS.n85 VSS.n40 7.19156
R389 VSS.n163 VSS.n89 7.19156
R390 VSS.n160 VSS.n90 7.19156
R391 VSS.n123 VSS.n122 7.19156
R392 VSS.n120 VSS.n119 7.19156
R393 VSS.n117 VSS.n116 7.19156
R394 VSS.n94 VSS.n93 7.19156
R395 VSS.n146 VSS.n95 7.19156
R396 VSS.n109 VSS.n108 7.19156
R397 VSS.n106 VSS.n105 7.19156
R398 VSS.n103 VSS.n102 7.19156
R399 VSS.n255 VSS.t211 7.19156
R400 VSS.n253 VSS.t64 7.19156
R401 VSS.n251 VSS.t87 7.19156
R402 VSS.n336 VSS.t284 7.19156
R403 VSS.n341 VSS.t128 7.19156
R404 VSS.n269 VSS.t276 6.88656
R405 VSS.n24 VSS.t287 6.88656
R406 VSS.n62 VSS.n49 6.88656
R407 VSS.n54 VSS.n53 6.88656
R408 VSS.n12 VSS.n11 6.01414
R409 VSS.n12 VSS.t167 6.01414
R410 VSS.n3 VSS.n2 6.01414
R411 VSS.n3 VSS.t42 6.01414
R412 VSS.n10 VSS.t221 5.91399
R413 VSS.n308 VSS.t315 5.91399
R414 VSS.n8 VSS.t82 5.91399
R415 VSS.n321 VSS.t313 5.91399
R416 VSS.n6 VSS.t146 5.91399
R417 VSS.n334 VSS.t172 5.91399
R418 VSS.n33 VSS.t182 5.91399
R419 VSS.n299 VSS.t299 5.91399
R420 VSS.n239 VSS.t174 5.91399
R421 VSS.n209 VSS.n198 5.91399
R422 VSS.n211 VSS.n196 5.91399
R423 VSS.n175 VSS.n174 5.91399
R424 VSS.n218 VSS.n168 5.91399
R425 VSS.n220 VSS.n88 5.91399
R426 VSS.n87 VSS.n38 5.91399
R427 VSS.n155 VSS.n154 5.91399
R428 VSS.n153 VSS.n91 5.91399
R429 VSS.n114 VSS.n113 5.91399
R430 VSS.n141 VSS.n140 5.91399
R431 VSS.n139 VSS.n96 5.91399
R432 VSS.n98 VSS.n97 5.91399
R433 VSS.n249 VSS.t102 5.91399
R434 VSS.n344 VSS.t301 5.91399
R435 VSS.n345 VSS.t305 5.91399
R436 VSS.n143 VSS.n142 5.2005
R437 VSS.n145 VSS.n144 5.2005
R438 VSS.n148 VSS.n147 5.2005
R439 VSS.n151 VSS.n150 5.2005
R440 VSS.n157 VSS.n156 5.2005
R441 VSS.n159 VSS.n158 5.2005
R442 VSS.n162 VSS.n161 5.2005
R443 VSS.n165 VSS.n164 5.2005
R444 VSS.n219 VSS.n167 5.2005
R445 VSS.n217 VSS.n169 5.2005
R446 VSS.n215 VSS.n171 5.2005
R447 VSS.n213 VSS.n173 5.2005
R448 VSS.n210 VSS.n197 5.2005
R449 VSS.n208 VSS.n199 5.2005
R450 VSS.n206 VSS.n201 5.2005
R451 VSS.n204 VSS.n203 5.2005
R452 VSS.n76 VSS.n75 5.2005
R453 VSS.n59 VSS.n58 5.2005
R454 VSS.n58 VSS.n57 5.2005
R455 VSS.n55 VSS.n45 5.2005
R456 VSS.n21 VSS.n20 5.2005
R457 VSS.n23 VSS.n19 5.2005
R458 VSS.n25 VSS.n18 5.2005
R459 VSS.n268 VSS.n267 5.2005
R460 VSS.n272 VSS.n16 5.2005
R461 VSS.n270 VSS.n17 5.2005
R462 VSS.n278 VSS.n13 5.2005
R463 VSS.n276 VSS.n14 5.2005
R464 VSS.n274 VSS.n15 5.2005
R465 VSS.n189 VSS.n188 5.2005
R466 VSS.n190 VSS.n185 5.2005
R467 VSS.n191 VSS.n182 5.2005
R468 VSS.n192 VSS.n179 5.2005
R469 VSS.n194 VSS.n193 5.2005
R470 VSS.n80 VSS.n79 5.2005
R471 VSS.n82 VSS.n43 5.2005
R472 VSS.n84 VSS.n41 5.2005
R473 VSS.n86 VSS.n39 5.2005
R474 VSS.n224 VSS.n223 5.2005
R475 VSS.n125 VSS.n124 5.2005
R476 VSS.n126 VSS.n121 5.2005
R477 VSS.n127 VSS.n118 5.2005
R478 VSS.n128 VSS.n115 5.2005
R479 VSS.n129 VSS.n112 5.2005
R480 VSS.n132 VSS.n110 5.2005
R481 VSS.n133 VSS.n107 5.2005
R482 VSS.n134 VSS.n104 5.2005
R483 VSS.n135 VSS.n101 5.2005
R484 VSS.n137 VSS.n136 5.2005
R485 VSS.n351 VSS.n350 5.2005
R486 VSS.n70 VSS.n67 5.2005
R487 VSS.n72 VSS.n65 5.2005
R488 VSS.n241 VSS.n240 5.2005
R489 VSS.n242 VSS.n237 5.2005
R490 VSS.n243 VSS.n235 5.2005
R491 VSS.n244 VSS.n233 5.2005
R492 VSS.n291 VSS.n290 5.2005
R493 VSS.n295 VSS.n294 5.2005
R494 VSS.n297 VSS.n296 5.2005
R495 VSS.n301 VSS.n300 5.2005
R496 VSS.n303 VSS.n302 5.2005
R497 VSS.n264 VSS.n27 5.2005
R498 VSS.n263 VSS.n29 5.2005
R499 VSS.n262 VSS.n31 5.2005
R500 VSS.n261 VSS.n34 5.2005
R501 VSS.n260 VSS.n35 5.2005
R502 VSS.n247 VSS.n231 5.2005
R503 VSS.n257 VSS.n256 5.2005
R504 VSS.n254 VSS.n229 5.2005
R505 VSS.n252 VSS.n230 5.2005
R506 VSS.n250 VSS.n248 5.2005
R507 VSS.n347 VSS.n346 5.2005
R508 VSS.n343 VSS.n342 5.2005
R509 VSS.n340 VSS.n339 5.2005
R510 VSS.n338 VSS.n337 5.2005
R511 VSS.n333 VSS.n332 5.2005
R512 VSS.n330 VSS.n329 5.2005
R513 VSS.n327 VSS.n326 5.2005
R514 VSS.n325 VSS.n324 5.2005
R515 VSS.n320 VSS.n319 5.2005
R516 VSS.n317 VSS.n316 5.2005
R517 VSS.n314 VSS.n313 5.2005
R518 VSS.n312 VSS.n311 5.2005
R519 VSS.n307 VSS.n306 5.2005
R520 VSS.n287 VSS.n286 5.2005
R521 VSS.n284 VSS.n283 5.2005
R522 VSS.n282 VSS.n281 5.2005
R523 VSS.n355 VSS.n1 5.2005
R524 VSS.n279 VSS.n12 3.36323
R525 VSS.n352 VSS.n3 3.36323
R526 VSS VSS.n279 2.40845
R527 VSS.n353 VSS 2.1304
R528 VSS.n354 VSS 1.99132
R529 VSS.n345 VSS.n0 1.03335
R530 VSS.n139 VSS.n138 1.03307
R531 VSS.n212 VSS.n195 0.846463
R532 VSS.n222 VSS.n221 0.846463
R533 VSS.n152 VSS.n92 0.846463
R534 VSS.n322 VSS.n7 0.845914
R535 VSS.n309 VSS.n9 0.845914
R536 VSS.n335 VSS.n5 0.845914
R537 VSS.n221 VSS 0.520683
R538 VSS VSS.n212 0.520683
R539 VSS VSS.n309 0.519858
R540 VSS VSS.n322 0.519858
R541 VSS.n142 VSS.n141 0.480225
R542 VSS.n146 VSS.n145 0.480225
R543 VSS.n156 VSS.n155 0.480225
R544 VSS.n160 VSS.n159 0.480225
R545 VSS.n219 VSS.n218 0.480225
R546 VSS.n217 VSS.n216 0.480225
R547 VSS.n210 VSS.n209 0.480225
R548 VSS.n208 VSS.n207 0.480225
R549 VSS.n286 VSS.n285 0.480225
R550 VSS.n307 VSS.n10 0.480225
R551 VSS.n316 VSS.n315 0.480225
R552 VSS.n320 VSS.n8 0.480225
R553 VSS.n329 VSS.n328 0.480225
R554 VSS.n333 VSS.n6 0.480225
R555 VSS.n343 VSS.n341 0.480225
R556 VSS.n346 VSS.n344 0.480225
R557 VSS.n64 VSS.n63 0.396541
R558 VSS.n60 VSS.n59 0.396541
R559 VSS.n57 VSS.n56 0.396541
R560 VSS.n271 VSS.n270 0.396455
R561 VSS.n22 VSS.n21 0.396455
R562 VSS.n26 VSS.n25 0.396455
R563 VSS.n277 VSS 0.379596
R564 VSS VSS.n69 0.378121
R565 VSS VSS.n353 0.357797
R566 VSS VSS.n28 0.343161
R567 VSS VSS.n30 0.343161
R568 VSS VSS.n292 0.343161
R569 VSS.n293 VSS 0.343161
R570 VSS VSS.n234 0.343161
R571 VSS VSS.n236 0.343161
R572 VSS.n184 VSS 0.343161
R573 VSS.n187 VSS 0.343161
R574 VSS VSS.n83 0.343161
R575 VSS VSS.n81 0.343161
R576 VSS.n120 VSS 0.343161
R577 VSS.n123 VSS 0.343161
R578 VSS.n106 VSS 0.343161
R579 VSS.n109 VSS 0.343161
R580 VSS VSS.n94 0.343161
R581 VSS.n163 VSS 0.343161
R582 VSS VSS.n214 0.343161
R583 VSS VSS.n205 0.343161
R584 VSS.n255 VSS 0.343161
R585 VSS.n253 VSS 0.343161
R586 VSS.n280 VSS 0.343161
R587 VSS.n310 VSS 0.343161
R588 VSS.n323 VSS 0.343161
R589 VSS.n336 VSS 0.343161
R590 VSS VSS.n71 0.311509
R591 VSS.n275 VSS 0.310668
R592 VSS.n34 VSS 0.289491
R593 VSS.n300 VSS 0.289491
R594 VSS.n240 VSS 0.289491
R595 VSS VSS.n179 0.289491
R596 VSS.n86 VSS 0.289491
R597 VSS VSS.n115 0.289491
R598 VSS VSS.n101 0.289491
R599 VSS VSS.n250 0.289491
R600 VSS.n353 VSS.n352 0.280231
R601 VSS.n62 VSS 0.27984
R602 VSS VSS.n54 0.27984
R603 VSS.n24 VSS 0.27984
R604 VSS.n269 VSS 0.27984
R605 VSS.n273 VSS 0.250123
R606 VSS VSS.n74 0.250123
R607 VSS.n274 VSS.n273 0.247195
R608 VSS.n74 VSS.n72 0.247195
R609 VSS VSS.n269 0.243604
R610 VSS VSS.n62 0.243604
R611 VSS.n54 VSS 0.243604
R612 VSS VSS.n24 0.243604
R613 VSS.n152 VSS 0.217656
R614 VSS VSS.n335 0.21683
R615 VSS VSS.n32 0.191234
R616 VSS VSS.n298 0.191234
R617 VSS VSS.n238 0.191234
R618 VSS.n181 VSS 0.191234
R619 VSS VSS.n85 0.191234
R620 VSS.n117 VSS 0.191234
R621 VSS.n103 VSS 0.191234
R622 VSS.n251 VSS 0.191234
R623 VSS.n309 VSS.n308 0.187931
R624 VSS.n322 VSS.n321 0.187931
R625 VSS.n335 VSS.n334 0.187931
R626 VSS.n153 VSS.n152 0.187105
R627 VSS.n221 VSS.n220 0.187105
R628 VSS.n212 VSS.n211 0.187105
R629 VSS.n276 VSS.n275 0.152211
R630 VSS.n71 VSS.n70 0.15137
R631 VSS.n279 VSS.n278 0.138903
R632 VSS.n352 VSS.n351 0.138903
R633 VSS VSS.n5 0.137685
R634 VSS VSS.n7 0.137685
R635 VSS VSS.n9 0.137685
R636 VSS VSS.n0 0.137685
R637 VSS.n195 VSS 0.137136
R638 VSS VSS.n222 0.137136
R639 VSS VSS.n92 0.137136
R640 VSS.n138 VSS 0.137136
R641 VSS.n28 VSS.n27 0.118573
R642 VSS.n30 VSS.n29 0.118573
R643 VSS.n32 VSS.n31 0.118573
R644 VSS.n292 VSS.n291 0.118573
R645 VSS.n294 VSS.n293 0.118573
R646 VSS.n298 VSS.n297 0.118573
R647 VSS.n234 VSS.n233 0.118573
R648 VSS.n236 VSS.n235 0.118573
R649 VSS.n238 VSS.n237 0.118573
R650 VSS.n182 VSS.n181 0.118573
R651 VSS.n185 VSS.n184 0.118573
R652 VSS.n188 VSS.n187 0.118573
R653 VSS.n85 VSS.n84 0.118573
R654 VSS.n83 VSS.n82 0.118573
R655 VSS.n81 VSS.n80 0.118573
R656 VSS.n118 VSS.n117 0.118573
R657 VSS.n121 VSS.n120 0.118573
R658 VSS.n124 VSS.n123 0.118573
R659 VSS.n104 VSS.n103 0.118573
R660 VSS.n107 VSS.n106 0.118573
R661 VSS.n110 VSS.n109 0.118573
R662 VSS.n147 VSS.n146 0.118573
R663 VSS.n151 VSS.n94 0.118573
R664 VSS.n162 VSS.n160 0.118573
R665 VSS.n164 VSS.n163 0.118573
R666 VSS.n216 VSS.n215 0.118573
R667 VSS.n214 VSS.n213 0.118573
R668 VSS.n207 VSS.n206 0.118573
R669 VSS.n205 VSS.n204 0.118573
R670 VSS.n256 VSS.n255 0.118573
R671 VSS.n254 VSS.n253 0.118573
R672 VSS.n252 VSS.n251 0.118573
R673 VSS.n281 VSS.n280 0.118573
R674 VSS.n285 VSS.n284 0.118573
R675 VSS.n311 VSS.n310 0.118573
R676 VSS.n315 VSS.n314 0.118573
R677 VSS.n324 VSS.n323 0.118573
R678 VSS.n328 VSS.n327 0.118573
R679 VSS.n337 VSS.n336 0.118573
R680 VSS.n341 VSS.n340 0.118573
R681 VSS VSS.n33 0.115271
R682 VSS VSS.n299 0.115271
R683 VSS VSS.n239 0.115271
R684 VSS VSS.n175 0.115271
R685 VSS.n87 VSS 0.115271
R686 VSS VSS.n114 0.115271
R687 VSS VSS.n98 0.115271
R688 VSS VSS.n139 0.115271
R689 VSS.n141 VSS 0.115271
R690 VSS VSS.n153 0.115271
R691 VSS.n155 VSS 0.115271
R692 VSS.n220 VSS 0.115271
R693 VSS.n218 VSS 0.115271
R694 VSS.n211 VSS 0.115271
R695 VSS.n209 VSS 0.115271
R696 VSS VSS.n249 0.115271
R697 VSS VSS.n10 0.115271
R698 VSS.n308 VSS 0.115271
R699 VSS VSS.n8 0.115271
R700 VSS.n321 VSS 0.115271
R701 VSS VSS.n6 0.115271
R702 VSS.n334 VSS 0.115271
R703 VSS.n344 VSS 0.115271
R704 VSS VSS.n345 0.115271
R705 VSS VSS.n277 0.113945
R706 VSS.n69 VSS 0.113945
R707 VSS.n33 VSS.n7 0.10206
R708 VSS.n299 VSS.n9 0.10206
R709 VSS.n239 VSS.n0 0.10206
R710 VSS.n195 VSS.n175 0.10206
R711 VSS.n222 VSS.n87 0.10206
R712 VSS.n114 VSS.n92 0.10206
R713 VSS.n138 VSS.n98 0.10206
R714 VSS.n249 VSS.n5 0.10206
R715 VSS.n272 VSS.n271 0.0675755
R716 VSS.n23 VSS.n22 0.0675755
R717 VSS.n268 VSS.n26 0.0675755
R718 VSS.n355 VSS.n354 0.0675755
R719 VSS.n75 VSS.n64 0.0667264
R720 VSS.n61 VSS.n60 0.0667264
R721 VSS.n56 VSS.n55 0.0667264
R722 VSS.n27 VSS 0.00545413
R723 VSS.n29 VSS 0.00545413
R724 VSS.n31 VSS 0.00545413
R725 VSS.n291 VSS 0.00545413
R726 VSS.n294 VSS 0.00545413
R727 VSS.n297 VSS 0.00545413
R728 VSS.n233 VSS 0.00545413
R729 VSS.n235 VSS 0.00545413
R730 VSS.n237 VSS 0.00545413
R731 VSS VSS.n182 0.00545413
R732 VSS VSS.n185 0.00545413
R733 VSS.n188 VSS 0.00545413
R734 VSS.n84 VSS 0.00545413
R735 VSS.n82 VSS 0.00545413
R736 VSS.n80 VSS 0.00545413
R737 VSS VSS.n118 0.00545413
R738 VSS VSS.n121 0.00545413
R739 VSS.n124 VSS 0.00545413
R740 VSS VSS.n104 0.00545413
R741 VSS VSS.n107 0.00545413
R742 VSS.n110 VSS 0.00545413
R743 VSS.n147 VSS 0.00545413
R744 VSS VSS.n151 0.00545413
R745 VSS VSS.n162 0.00545413
R746 VSS.n164 VSS 0.00545413
R747 VSS.n215 VSS 0.00545413
R748 VSS.n213 VSS 0.00545413
R749 VSS.n206 VSS 0.00545413
R750 VSS.n204 VSS 0.00545413
R751 VSS.n256 VSS 0.00545413
R752 VSS VSS.n254 0.00545413
R753 VSS VSS.n252 0.00545413
R754 VSS.n281 VSS 0.00545413
R755 VSS.n284 VSS 0.00545413
R756 VSS.n311 VSS 0.00545413
R757 VSS.n314 VSS 0.00545413
R758 VSS.n324 VSS 0.00545413
R759 VSS.n327 VSS 0.00545413
R760 VSS.n337 VSS 0.00545413
R761 VSS.n340 VSS 0.00545413
R762 VSS.n34 VSS 0.00380275
R763 VSS.n300 VSS 0.00380275
R764 VSS.n240 VSS 0.00380275
R765 VSS.n270 VSS 0.00380275
R766 VSS.n179 VSS 0.00380275
R767 VSS VSS.n86 0.00380275
R768 VSS.n115 VSS 0.00380275
R769 VSS.n101 VSS 0.00380275
R770 VSS.n142 VSS 0.00380275
R771 VSS.n145 VSS 0.00380275
R772 VSS.n156 VSS 0.00380275
R773 VSS.n159 VSS 0.00380275
R774 VSS VSS.n219 0.00380275
R775 VSS VSS.n217 0.00380275
R776 VSS VSS.n210 0.00380275
R777 VSS VSS.n208 0.00380275
R778 VSS.n63 VSS 0.00380275
R779 VSS.n57 VSS 0.00380275
R780 VSS.n59 VSS 0.00380275
R781 VSS.n21 VSS 0.00380275
R782 VSS.n25 VSS 0.00380275
R783 VSS.n250 VSS 0.00380275
R784 VSS.n286 VSS 0.00380275
R785 VSS VSS.n307 0.00380275
R786 VSS.n316 VSS 0.00380275
R787 VSS VSS.n320 0.00380275
R788 VSS.n329 VSS 0.00380275
R789 VSS VSS.n333 0.00380275
R790 VSS VSS.n343 0.00380275
R791 VSS.n346 VSS 0.00380275
R792 VSS.n278 VSS 0.00352521
R793 VSS.n351 VSS 0.00352521
R794 VSS.n231 VSS 0.00219811
R795 VSS.n35 VSS 0.00219811
R796 VSS.n302 VSS 0.00219811
R797 VSS VSS.n276 0.00219811
R798 VSS VSS.n274 0.00219811
R799 VSS VSS.n272 0.00219811
R800 VSS VSS.n194 0.00219811
R801 VSS.n223 VSS 0.00219811
R802 VSS.n112 VSS 0.00219811
R803 VSS VSS.n137 0.00219811
R804 VSS.n70 VSS 0.00219811
R805 VSS.n72 VSS 0.00219811
R806 VSS.n75 VSS 0.00219811
R807 VSS VSS.n61 0.00219811
R808 VSS.n55 VSS 0.00219811
R809 VSS VSS.n23 0.00219811
R810 VSS VSS.n268 0.00219811
R811 VSS VSS.n355 0.00219811
R812 VDD.n428 VDD.n139 190685
R813 VDD.n428 VDD.t374 83097.6
R814 VDD.t430 VDD.n243 29077.7
R815 VDD.n119 VDD.n118 11185.2
R816 VDD.n130 VDD.n129 11185.2
R817 VDD.t188 VDD.n426 1105.93
R818 VDD.t39 VDD.n241 1105.93
R819 VDD.t97 VDD.t41 961.905
R820 VDD.t295 VDD.t37 961.905
R821 VDD.t244 VDD.t321 961.905
R822 VDD.t329 VDD.t124 961.905
R823 VDD.t277 VDD.t388 961.905
R824 VDD.t234 VDD.t463 961.905
R825 VDD.t133 VDD.t382 765.152
R826 VDD.t64 VDD.t49 765.152
R827 VDD.t365 VDD.t131 765.152
R828 VDD.t261 VDD.t69 765.152
R829 VDD.t61 VDD.t46 765.152
R830 VDD.t221 VDD.t129 765.152
R831 VDD.t121 VDD.t202 765.152
R832 VDD.t285 VDD.t207 765.152
R833 VDD.t357 VDD.t319 765.152
R834 VDD.t258 VDD.t343 765.152
R835 VDD.t282 VDD.t210 765.152
R836 VDD.t252 VDD.t317 765.152
R837 VDD.t255 VDD.t288 765.152
R838 VDD.t58 VDD.t25 765.152
R839 VDD.t4 VDD.t2 765.152
R840 VDD.t94 VDD.t236 765.152
R841 VDD.t401 VDD.t84 765.152
R842 VDD.t126 VDD.t472 765.152
R843 VDD.t385 VDD.t371 765.152
R844 VDD.t81 VDD.t398 765.152
R845 VDD.t449 VDD.t470 765.152
R846 VDD.t465 VDD.t300 765.152
R847 VDD.t28 VDD.t55 765.152
R848 VDD.t78 VDD.t0 765.152
R849 VDD.t274 VDD.t434 765.152
R850 VDD.t212 VDD.t216 765.152
R851 VDD.t419 VDD.t461 765.152
R852 VDD.t241 VDD.t226 765.152
R853 VDD.t87 VDD.t353 765.152
R854 VDD.t23 VDD.t247 765.152
R855 VDD.t455 VDD.t116 765.152
R856 VDD.t75 VDD.t266 765.152
R857 VDD.t280 VDD.t191 765.152
R858 VDD.t113 VDD.t360 765.152
R859 VDD.t264 VDD.t73 765.152
R860 VDD.t271 VDD.t348 765.152
R861 VDD.t100 VDD.t224 765.152
R862 VDD.t53 VDD.t111 765.152
R863 VDD.t444 VDD.t119 765.152
R864 VDD.n118 VDD.t51 676.191
R865 VDD.n129 VDD.t89 676.191
R866 VDD.n139 VDD.t218 669.048
R867 VDD.t195 VDD.t355 645.307
R868 VDD.t228 VDD.t31 642.843
R869 VDD.n428 VDD.n427 525.424
R870 VDD.n243 VDD.n242 525.424
R871 VDD.n119 VDD.t150 485.714
R872 VDD.n130 VDD.t92 485.714
R873 VDD VDD.n83 429.187
R874 VDD.n236 VDD 427.092
R875 VDD.n238 VDD 427.092
R876 VDD VDD.n294 426.699
R877 VDD VDD.n258 426.699
R878 VDD VDD.n281 426.699
R879 VDD.t18 VDD.n119 426.44
R880 VDD.t421 VDD.n130 426.44
R881 VDD.n240 VDD 425.019
R882 VDD VDD.n416 424.618
R883 VDD VDD.n411 424.618
R884 VDD VDD.n421 422.557
R885 VDD.n416 VDD.t338 386.365
R886 VDD.n411 VDD.t105 386.365
R887 VDD.t297 VDD.n294 386.365
R888 VDD.n281 VDD.t153 386.365
R889 VDD.n258 VDD.t395 386.365
R890 VDD.t412 VDD.n238 386.365
R891 VDD.t447 VDD.n236 386.365
R892 VDD.n83 VDD.t457 386.365
R893 VDD.t37 VDD.t13 380.952
R894 VDD.t406 VDD.t329 380.952
R895 VDD.t374 VDD.t234 380.952
R896 VDD.n421 VDD.t103 378.788
R897 VDD.n416 VDD.t310 378.788
R898 VDD.n411 VDD.t200 378.788
R899 VDD.n240 VDD.t442 378.788
R900 VDD.n238 VDD.t7 378.788
R901 VDD.n236 VDD.t436 378.788
R902 VDD.t382 VDD.t336 303.031
R903 VDD.t69 VDD.t139 303.031
R904 VDD.t459 VDD.t61 303.031
R905 VDD.t202 VDD.t315 303.031
R906 VDD.t346 VDD.t285 303.031
R907 VDD.t343 VDD.t303 303.031
R908 VDD.t288 VDD.t334 303.031
R909 VDD.t236 VDD.t430 303.031
R910 VDD.t371 VDD.t428 303.031
R911 VDD.t144 VDD.t81 303.031
R912 VDD.t300 VDD.t378 303.031
R913 VDD.t293 VDD.t28 303.031
R914 VDD.t331 VDD.t212 303.031
R915 VDD.t452 VDD.t419 303.031
R916 VDD.t390 VDD.t87 303.031
R917 VDD.t409 VDD.t23 303.031
R918 VDD.t191 VDD.t416 303.031
R919 VDD.t323 VDD.t264 303.031
R920 VDD.t423 VDD.t271 303.031
R921 VDD.t141 VDD.t53 303.031
R922 VDD.t10 VDD.t444 303.031
R923 VDD.n139 VDD.t214 292.858
R924 VDD.n118 VDD.t108 285.714
R925 VDD.n129 VDD.t350 285.714
R926 VDD.n110 VDD.t34 242.857
R927 VDD.n111 VDD.t97 242.857
R928 VDD.t108 VDD.n117 242.857
R929 VDD.t13 VDD.n3 242.857
R930 VDD.n121 VDD.t326 242.857
R931 VDD.n123 VDD.t244 242.857
R932 VDD.t350 VDD.n125 242.857
R933 VDD.n128 VDD.t406 242.857
R934 VDD.n132 VDD.t231 242.857
R935 VDD.n134 VDD.t277 242.857
R936 VDD.t218 VDD.n136 242.857
R937 VDD.t442 VDD.n239 193.183
R938 VDD.t7 VDD.n237 193.183
R939 VDD.t436 VDD.n235 193.183
R940 VDD.n448 VDD.t403 193.183
R941 VDD.n450 VDD.t274 193.183
R942 VDD.n453 VDD.t331 193.183
R943 VDD.n456 VDD.t452 193.183
R944 VDD.n483 VDD.t20 193.183
R945 VDD.n485 VDD.t241 193.183
R946 VDD.n488 VDD.t390 193.183
R947 VDD.n491 VDD.t409 193.183
R948 VDD.n70 VDD.t362 193.183
R949 VDD.n76 VDD.t116 193.183
R950 VDD.n77 VDD.t75 193.183
R951 VDD.n82 VDD.t416 193.183
R952 VDD.n16 VDD.t268 193.183
R953 VDD.n18 VDD.t113 193.183
R954 VDD.n21 VDD.t323 193.183
R955 VDD.n24 VDD.t423 193.183
R956 VDD.n86 VDD.t439 193.183
R957 VDD.n88 VDD.t100 193.183
R958 VDD.n91 VDD.t141 193.183
R959 VDD.n94 VDD.t10 193.183
R960 VDD.t103 VDD.n420 191.288
R961 VDD.t310 VDD.n415 191.288
R962 VDD.t200 VDD.n410 191.288
R963 VDD.t336 VDD.n296 191.288
R964 VDD.t49 VDD.n300 191.288
R965 VDD.t131 VDD.n302 191.288
R966 VDD.n304 VDD.t426 191.288
R967 VDD.t139 VDD.n347 191.288
R968 VDD.n348 VDD.t459 191.288
R969 VDD.t129 VDD.n356 191.288
R970 VDD.n357 VDD.t67 191.288
R971 VDD.t315 VDD.n383 191.288
R972 VDD.n384 VDD.t346 191.288
R973 VDD.t319 VDD.n392 191.288
R974 VDD.n393 VDD.t193 191.288
R975 VDD.t303 VDD.n287 191.288
R976 VDD.t210 VDD.n288 191.288
R977 VDD.t317 VDD.n290 191.288
R978 VDD.n292 VDD.t341 191.288
R979 VDD.t334 VDD.n266 191.288
R980 VDD.n267 VDD.t58 191.288
R981 VDD.t2 VDD.n275 191.288
R982 VDD.n276 VDD.t291 191.288
R983 VDD.n244 VDD.t401 191.288
R984 VDD.t472 VDD.n252 191.288
R985 VDD.n253 VDD.t239 191.288
R986 VDD.t428 VDD.n189 191.288
R987 VDD.n190 VDD.t144 191.288
R988 VDD.t470 VDD.n198 191.288
R989 VDD.n199 VDD.t393 191.288
R990 VDD.t378 VDD.n163 191.288
R991 VDD.n164 VDD.t293 191.288
R992 VDD.t0 VDD.n172 191.288
R993 VDD.n173 VDD.t305 191.288
R994 VDD.t41 VDD.n110 138.095
R995 VDD.n111 VDD.t51 138.095
R996 VDD.n117 VDD.t295 138.095
R997 VDD.t150 VDD.n3 138.095
R998 VDD.t321 VDD.n121 138.095
R999 VDD.t89 VDD.n123 138.095
R1000 VDD.t124 VDD.n125 138.095
R1001 VDD.t92 VDD.n128 138.095
R1002 VDD.t388 VDD.n132 138.095
R1003 VDD.t214 VDD.n134 138.095
R1004 VDD.t463 VDD.n136 138.095
R1005 VDD.t72 VDD.t60 120.755
R1006 VDD.t91 VDD.t273 120.755
R1007 VDD.n420 VDD.t338 111.743
R1008 VDD.n415 VDD.t105 111.743
R1009 VDD.n410 VDD.t307 111.743
R1010 VDD.n296 VDD.t297 111.743
R1011 VDD.n300 VDD.t133 111.743
R1012 VDD.n302 VDD.t64 111.743
R1013 VDD.n304 VDD.t365 111.743
R1014 VDD.n347 VDD.t170 111.743
R1015 VDD.n348 VDD.t261 111.743
R1016 VDD.n356 VDD.t46 111.743
R1017 VDD.n357 VDD.t221 111.743
R1018 VDD.n383 VDD.t181 111.743
R1019 VDD.n384 VDD.t121 111.743
R1020 VDD.n392 VDD.t207 111.743
R1021 VDD.n393 VDD.t357 111.743
R1022 VDD.n287 VDD.t153 111.743
R1023 VDD.n288 VDD.t258 111.743
R1024 VDD.n290 VDD.t282 111.743
R1025 VDD.n292 VDD.t252 111.743
R1026 VDD.n266 VDD.t395 111.743
R1027 VDD.n267 VDD.t255 111.743
R1028 VDD.n275 VDD.t25 111.743
R1029 VDD.n276 VDD.t4 111.743
R1030 VDD.n244 VDD.t94 111.743
R1031 VDD.n252 VDD.t84 111.743
R1032 VDD.n253 VDD.t126 111.743
R1033 VDD.n189 VDD.t174 111.743
R1034 VDD.n190 VDD.t385 111.743
R1035 VDD.n198 VDD.t398 111.743
R1036 VDD.n199 VDD.t449 111.743
R1037 VDD.n163 VDD.t157 111.743
R1038 VDD.n164 VDD.t465 111.743
R1039 VDD.n172 VDD.t55 111.743
R1040 VDD.n173 VDD.t78 111.743
R1041 VDD.n239 VDD.t412 109.849
R1042 VDD.n237 VDD.t447 109.849
R1043 VDD.n235 VDD.t16 109.849
R1044 VDD.t434 VDD.n448 109.849
R1045 VDD.t216 VDD.n450 109.849
R1046 VDD.t461 VDD.n453 109.849
R1047 VDD.n456 VDD.t164 109.849
R1048 VDD.t226 VDD.n483 109.849
R1049 VDD.t353 VDD.n485 109.849
R1050 VDD.t247 VDD.n488 109.849
R1051 VDD.n491 VDD.t178 109.849
R1052 VDD.n70 VDD.t455 109.849
R1053 VDD.t266 VDD.n76 109.849
R1054 VDD.n77 VDD.t280 109.849
R1055 VDD.t457 VDD.n82 109.849
R1056 VDD.t360 VDD.n16 109.849
R1057 VDD.t73 VDD.n18 109.849
R1058 VDD.t348 VDD.n21 109.849
R1059 VDD.n24 VDD.t147 109.849
R1060 VDD.t224 VDD.n86 109.849
R1061 VDD.t111 VDD.n88 109.849
R1062 VDD.t119 VDD.n91 109.849
R1063 VDD.n94 VDD.t161 109.849
R1064 VDD.n431 VDD.t197 105.66
R1065 VDD.n206 VDD.t380 105.66
R1066 VDD.t197 VDD.t167 63.3967
R1067 VDD.t380 VDD.t185 63.3967
R1068 VDD.n294 VDD.t136 62.1896
R1069 VDD.n281 VDD.t312 62.1896
R1070 VDD.n258 VDD.t368 62.1896
R1071 VDD.n416 VDD.t43 61.8817
R1072 VDD.n411 VDD.t249 61.8817
R1073 VDD.n421 VDD.t228 61.5769
R1074 VDD.n83 VDD.t414 59.702
R1075 VDD.n238 VDD.t205 59.4064
R1076 VDD.n236 VDD.t468 59.4064
R1077 VDD.t355 VDD.n240 59.1138
R1078 VDD.n426 VDD.t31 55.0852
R1079 VDD.n427 VDD.t188 55.0852
R1080 VDD.n242 VDD.t39 55.0852
R1081 VDD.n241 VDD.t195 55.0852
R1082 VDD.n429 VDD.n428 45.2835
R1083 VDD.t185 VDD.n203 44.5288
R1084 VDD.n243 VDD.n203 44.5288
R1085 VDD.t167 VDD.n429 43.7741
R1086 VDD.n338 VDD.t169 30.9379
R1087 VDD.n312 VDD.t156 30.9379
R1088 VDD.n25 VDD.t146 30.9379
R1089 VDD.n27 VDD.t177 30.9379
R1090 VDD.n48 VDD.t149 30.721
R1091 VDD.n330 VDD.t152 30.7204
R1092 VDD.n318 VDD.t184 30.7203
R1093 VDD.n38 VDD.t166 30.7203
R1094 VDD.n45 VDD.t160 30.3459
R1095 VDD.n324 VDD.t173 30.2877
R1096 VDD.n334 VDD.t180 30.2877
R1097 VDD.n33 VDD.t163 30.0062
R1098 VDD.n334 VDD.t477 24.9141
R1099 VDD.n45 VDD.t490 24.8618
R1100 VDD.n338 VDD.t483 24.5101
R1101 VDD.n323 VDD.t482 24.5101
R1102 VDD.n312 VDD.t488 24.5101
R1103 VDD.n25 VDD.t491 24.5101
R1104 VDD.n27 VDD.t478 24.5101
R1105 VDD.n48 VDD.t484 24.4816
R1106 VDD.n38 VDD.t479 24.4814
R1107 VDD.n318 VDD.t476 24.4814
R1108 VDD.n330 VDD.t489 24.4813
R1109 VDD.n35 VDD.t485 24.4392
R1110 VDD.t60 VDD.n431 15.0948
R1111 VDD.n206 VDD.t91 15.0948
R1112 VDD VDD.t421 10.5649
R1113 VDD VDD.t18 10.5649
R1114 VDD.n323 VDD.n322 8.0005
R1115 VDD.n35 VDD.n34 8.0005
R1116 VDD VDD.t72 7.80993
R1117 VDD.t273 VDD 7.80993
R1118 VDD.n55 VDD.n54 6.39748
R1119 VDD.n339 VDD.n337 6.39705
R1120 VDD.n431 VDD 6.30126
R1121 VDD VDD.n206 6.30126
R1122 VDD.n358 VDD.n357 6.3005
R1123 VDD.n356 VDD.n355 6.3005
R1124 VDD.n349 VDD.n348 6.3005
R1125 VDD.n347 VDD.n346 6.3005
R1126 VDD.n370 VDD.n296 6.3005
R1127 VDD.n367 VDD.n300 6.3005
R1128 VDD.n364 VDD.n302 6.3005
R1129 VDD.n361 VDD.n304 6.3005
R1130 VDD.n383 VDD.n382 6.3005
R1131 VDD.n385 VDD.n384 6.3005
R1132 VDD.n392 VDD.n391 6.3005
R1133 VDD.n394 VDD.n393 6.3005
R1134 VDD.n235 VDD.n234 6.3005
R1135 VDD.n237 VDD.n228 6.3005
R1136 VDD.n239 VDD.n223 6.3005
R1137 VDD.n241 VDD.n218 6.3005
R1138 VDD.n242 VDD 6.3005
R1139 VDD.n210 VDD.n203 6.3005
R1140 VDD.n245 VDD.n244 6.3005
R1141 VDD.n252 VDD.n251 6.3005
R1142 VDD.n254 VDD.n253 6.3005
R1143 VDD.n189 VDD.n188 6.3005
R1144 VDD.n191 VDD.n190 6.3005
R1145 VDD.n198 VDD.n197 6.3005
R1146 VDD.n200 VDD.n199 6.3005
R1147 VDD.n266 VDD.n265 6.3005
R1148 VDD.n268 VDD.n267 6.3005
R1149 VDD.n275 VDD.n274 6.3005
R1150 VDD.n277 VDD.n276 6.3005
R1151 VDD.n163 VDD.n162 6.3005
R1152 VDD.n165 VDD.n164 6.3005
R1153 VDD.n172 VDD.n171 6.3005
R1154 VDD.n174 VDD.n173 6.3005
R1155 VDD.n287 VDD.n286 6.3005
R1156 VDD.n404 VDD.n288 6.3005
R1157 VDD.n401 VDD.n290 6.3005
R1158 VDD.n398 VDD.n292 6.3005
R1159 VDD.n410 VDD.n409 6.3005
R1160 VDD.n415 VDD.n414 6.3005
R1161 VDD.n420 VDD.n419 6.3005
R1162 VDD.n426 VDD.n425 6.3005
R1163 VDD.n427 VDD 6.3005
R1164 VDD.n435 VDD.n429 6.3005
R1165 VDD.n439 VDD.n136 6.3005
R1166 VDD.n442 VDD.n134 6.3005
R1167 VDD.n445 VDD.n132 6.3005
R1168 VDD.n457 VDD.n456 6.3005
R1169 VDD.n460 VDD.n453 6.3005
R1170 VDD.n463 VDD.n450 6.3005
R1171 VDD.n466 VDD.n448 6.3005
R1172 VDD.n471 VDD.n128 6.3005
R1173 VDD.n474 VDD.n125 6.3005
R1174 VDD.n477 VDD.n123 6.3005
R1175 VDD.n480 VDD.n121 6.3005
R1176 VDD.n492 VDD.n491 6.3005
R1177 VDD.n495 VDD.n488 6.3005
R1178 VDD.n498 VDD.n485 6.3005
R1179 VDD.n501 VDD.n483 6.3005
R1180 VDD.n58 VDD.n24 6.3005
R1181 VDD.n61 VDD.n21 6.3005
R1182 VDD.n64 VDD.n18 6.3005
R1183 VDD.n67 VDD.n16 6.3005
R1184 VDD.n82 VDD.n81 6.3005
R1185 VDD.n78 VDD.n77 6.3005
R1186 VDD.n76 VDD.n75 6.3005
R1187 VDD.n71 VDD.n70 6.3005
R1188 VDD.n95 VDD.n94 6.3005
R1189 VDD.n98 VDD.n91 6.3005
R1190 VDD.n101 VDD.n88 6.3005
R1191 VDD.n104 VDD.n86 6.3005
R1192 VDD.n506 VDD.n3 6.3005
R1193 VDD.n117 VDD.n116 6.3005
R1194 VDD.n112 VDD.n111 6.3005
R1195 VDD.n110 VDD.n109 6.3005
R1196 VDD.n327 VDD.n326 5.30733
R1197 VDD.n44 VDD.n43 5.30657
R1198 VDD.n382 VDD.n378 5.213
R1199 VDD.n188 VDD.n184 5.213
R1200 VDD.n162 VDD.n158 5.213
R1201 VDD.n457 VDD.t165 5.213
R1202 VDD.n492 VDD.t179 5.213
R1203 VDD.n95 VDD.t162 5.213
R1204 VDD VDD.t377 5.16454
R1205 VDD VDD.n205 5.16369
R1206 VDD.n219 VDD.t196 5.14212
R1207 VDD.n422 VDD.n140 5.14212
R1208 VDD.n371 VDD.n295 5.13287
R1209 VDD.n368 VDD.n299 5.13287
R1210 VDD.n366 VDD.t50 5.13287
R1211 VDD.n365 VDD.n301 5.13287
R1212 VDD.n363 VDD.t132 5.13287
R1213 VDD.n362 VDD.n303 5.13287
R1214 VDD.n360 VDD.t427 5.13287
R1215 VDD.n309 VDD.n308 5.13287
R1216 VDD.n351 VDD.n305 5.13287
R1217 VDD.n354 VDD.t130 5.13287
R1218 VDD.n353 VDD.n352 5.13287
R1219 VDD.n359 VDD.t68 5.13287
R1220 VDD.n377 VDD.n376 5.13287
R1221 VDD.n387 VDD.n373 5.13287
R1222 VDD.n390 VDD.t320 5.13287
R1223 VDD.n389 VDD.n388 5.13287
R1224 VDD.n395 VDD.t194 5.13287
R1225 VDD.n208 VDD.n204 5.13287
R1226 VDD.n233 VDD.t17 5.13287
R1227 VDD.n232 VDD.n230 5.13287
R1228 VDD.n229 VDD.t448 5.13287
R1229 VDD.n227 VDD.n225 5.13287
R1230 VDD.n224 VDD.t413 5.13287
R1231 VDD.n222 VDD.n220 5.13287
R1232 VDD.n212 VDD.n211 5.13287
R1233 VDD.n246 VDD.t402 5.13287
R1234 VDD.n247 VDD.n202 5.13287
R1235 VDD.n250 VDD.t473 5.13287
R1236 VDD.n249 VDD.n248 5.13287
R1237 VDD.n255 VDD.t240 5.13287
R1238 VDD.n183 VDD.n182 5.13287
R1239 VDD.n193 VDD.n179 5.13287
R1240 VDD.n196 VDD.t471 5.13287
R1241 VDD.n195 VDD.n194 5.13287
R1242 VDD.n201 VDD.t394 5.13287
R1243 VDD.n259 VDD.n177 5.13287
R1244 VDD.n263 VDD.n262 5.13287
R1245 VDD.n269 VDD.t59 5.13287
R1246 VDD.n270 VDD.n176 5.13287
R1247 VDD.n273 VDD.t3 5.13287
R1248 VDD.n272 VDD.n271 5.13287
R1249 VDD.n278 VDD.t292 5.13287
R1250 VDD.n157 VDD.n156 5.13287
R1251 VDD.n167 VDD.n153 5.13287
R1252 VDD.n170 VDD.t1 5.13287
R1253 VDD.n169 VDD.n168 5.13287
R1254 VDD.n175 VDD.t306 5.13287
R1255 VDD.n282 VDD.n151 5.13287
R1256 VDD.n405 VDD.n150 5.13287
R1257 VDD.n403 VDD.t211 5.13287
R1258 VDD.n402 VDD.n289 5.13287
R1259 VDD.n400 VDD.t318 5.13287
R1260 VDD.n399 VDD.n291 5.13287
R1261 VDD.n397 VDD.t342 5.13287
R1262 VDD.n407 VDD.n149 5.13287
R1263 VDD.n408 VDD.t201 5.13287
R1264 VDD.n412 VDD.n146 5.13287
R1265 VDD.n413 VDD.t311 5.13287
R1266 VDD.n417 VDD.n143 5.13287
R1267 VDD.n418 VDD.t104 5.13287
R1268 VDD.n433 VDD.t168 5.13287
R1269 VDD.n438 VDD.t464 5.13287
R1270 VDD.n440 VDD.n135 5.13287
R1271 VDD.n441 VDD.t215 5.13287
R1272 VDD.n443 VDD.n133 5.13287
R1273 VDD.n444 VDD.t389 5.13287
R1274 VDD.n446 VDD.n131 5.13287
R1275 VDD.n459 VDD.t462 5.13287
R1276 VDD.n462 VDD.t217 5.13287
R1277 VDD.n464 VDD.n449 5.13287
R1278 VDD.n465 VDD.t435 5.13287
R1279 VDD.n467 VDD.n447 5.13287
R1280 VDD.n470 VDD.t93 5.13287
R1281 VDD.n473 VDD.t125 5.13287
R1282 VDD.n475 VDD.n124 5.13287
R1283 VDD.n476 VDD.t90 5.13287
R1284 VDD.n478 VDD.n122 5.13287
R1285 VDD.n479 VDD.t322 5.13287
R1286 VDD.n481 VDD.n120 5.13287
R1287 VDD.n494 VDD.t248 5.13287
R1288 VDD.n497 VDD.t354 5.13287
R1289 VDD.n499 VDD.n484 5.13287
R1290 VDD.n500 VDD.t227 5.13287
R1291 VDD.n502 VDD.n482 5.13287
R1292 VDD.n8 VDD.t458 5.13287
R1293 VDD.n79 VDD.t281 5.13287
R1294 VDD.n12 VDD.n11 5.13287
R1295 VDD.n74 VDD.t267 5.13287
R1296 VDD.n73 VDD.n13 5.13287
R1297 VDD.n72 VDD.t456 5.13287
R1298 VDD.n69 VDD.n14 5.13287
R1299 VDD.n60 VDD.t349 5.13287
R1300 VDD.n63 VDD.t74 5.13287
R1301 VDD.n65 VDD.n17 5.13287
R1302 VDD.n66 VDD.t361 5.13287
R1303 VDD.n68 VDD.n15 5.13287
R1304 VDD.n97 VDD.t120 5.13287
R1305 VDD.n100 VDD.t112 5.13287
R1306 VDD.n102 VDD.n87 5.13287
R1307 VDD.n103 VDD.t225 5.13287
R1308 VDD.n105 VDD.n85 5.13287
R1309 VDD.n505 VDD.t151 5.13287
R1310 VDD.n115 VDD.t296 5.13287
R1311 VDD.n114 VDD.n4 5.13287
R1312 VDD.n113 VDD.t52 5.13287
R1313 VDD.n6 VDD.n5 5.13287
R1314 VDD.n108 VDD.t42 5.13287
R1315 VDD.n107 VDD.n7 5.13287
R1316 VDD.n217 VDD.t40 5.09693
R1317 VDD.n424 VDD.n423 5.09693
R1318 VDD.n372 VDD.n293 5.09407
R1319 VDD.n231 VDD.t469 5.09407
R1320 VDD.n226 VDD.t206 5.09407
R1321 VDD.n221 VDD.t356 5.09407
R1322 VDD.n257 VDD.n178 5.09407
R1323 VDD.n280 VDD.n152 5.09407
R1324 VDD.n148 VDD.n147 5.09407
R1325 VDD.n145 VDD.n144 5.09407
R1326 VDD.n142 VDD.n141 5.09407
R1327 VDD.n469 VDD.t422 5.09407
R1328 VDD.n504 VDD.t19 5.09407
R1329 VDD.n84 VDD.t415 5.09407
R1330 VDD.n342 VDD.n341 4.8755
R1331 VDD.n57 VDD.t148 4.8755
R1332 VDD.n337 VDD.n327 4.84121
R1333 VDD.n54 VDD.n44 4.84121
R1334 VDD.n317 VDD.n316 4.5005
R1335 VDD.n319 VDD.n316 4.5005
R1336 VDD.n311 VDD.n310 4.5005
R1337 VDD.n313 VDD.n310 4.5005
R1338 VDD.n329 VDD.n328 4.5005
R1339 VDD.n331 VDD.n328 4.5005
R1340 VDD.n36 VDD.n35 4.5005
R1341 VDD.n39 VDD.n37 4.5005
R1342 VDD.n40 VDD.n37 4.5005
R1343 VDD.n28 VDD.n26 4.5005
R1344 VDD.n29 VDD.n26 4.5005
R1345 VDD.n49 VDD.n47 4.5005
R1346 VDD.n50 VDD.n47 4.5005
R1347 VDD.n432 VDD 4.40201
R1348 VDD.n207 VDD 4.40201
R1349 VDD.n209 VDD.t381 3.94862
R1350 VDD.n434 VDD.n430 3.94862
R1351 VDD.n33 VDD.n32 3.61662
R1352 VDD.n207 VDD 3.52487
R1353 VDD.n432 VDD 3.47987
R1354 VDD.n339 VDD.n338 2.88198
R1355 VDD.n55 VDD.n25 2.88182
R1356 VDD.n215 VDD.n214 2.88011
R1357 VDD.n437 VDD.n138 2.87966
R1358 VDD.n369 VDD.n298 2.85787
R1359 VDD.n345 VDD.n344 2.85787
R1360 VDD.n350 VDD.n307 2.85787
R1361 VDD.n381 VDD.n380 2.85787
R1362 VDD.n386 VDD.n375 2.85787
R1363 VDD.n187 VDD.n186 2.85787
R1364 VDD.n192 VDD.n181 2.85787
R1365 VDD.n264 VDD.n261 2.85787
R1366 VDD.n161 VDD.n160 2.85787
R1367 VDD.n166 VDD.n155 2.85787
R1368 VDD.n285 VDD.n284 2.85787
R1369 VDD.n458 VDD.n455 2.85787
R1370 VDD.n461 VDD.n452 2.85787
R1371 VDD.n472 VDD.n127 2.85787
R1372 VDD.n493 VDD.n490 2.85787
R1373 VDD.n496 VDD.n487 2.85787
R1374 VDD.n80 VDD.n10 2.85787
R1375 VDD.n59 VDD.n23 2.85787
R1376 VDD.n62 VDD.n20 2.85787
R1377 VDD.n96 VDD.n93 2.85787
R1378 VDD.n99 VDD.n90 2.85787
R1379 VDD.n507 VDD.n2 2.85787
R1380 VDD.n138 VDD.t235 2.2755
R1381 VDD.n138 VDD.n137 2.2755
R1382 VDD.n298 VDD.t337 2.2755
R1383 VDD.n298 VDD.n297 2.2755
R1384 VDD.n344 VDD.t140 2.2755
R1385 VDD.n344 VDD.n343 2.2755
R1386 VDD.n307 VDD.t460 2.2755
R1387 VDD.n307 VDD.n306 2.2755
R1388 VDD.n380 VDD.t316 2.2755
R1389 VDD.n380 VDD.n379 2.2755
R1390 VDD.n375 VDD.t347 2.2755
R1391 VDD.n375 VDD.n374 2.2755
R1392 VDD.n214 VDD.t431 2.2755
R1393 VDD.n214 VDD.n213 2.2755
R1394 VDD.n186 VDD.t429 2.2755
R1395 VDD.n186 VDD.n185 2.2755
R1396 VDD.n181 VDD.t145 2.2755
R1397 VDD.n181 VDD.n180 2.2755
R1398 VDD.n261 VDD.t335 2.2755
R1399 VDD.n261 VDD.n260 2.2755
R1400 VDD.n160 VDD.t379 2.2755
R1401 VDD.n160 VDD.n159 2.2755
R1402 VDD.n155 VDD.t294 2.2755
R1403 VDD.n155 VDD.n154 2.2755
R1404 VDD.n284 VDD.t304 2.2755
R1405 VDD.n284 VDD.n283 2.2755
R1406 VDD.n455 VDD.t420 2.2755
R1407 VDD.n455 VDD.n454 2.2755
R1408 VDD.n452 VDD.t213 2.2755
R1409 VDD.n452 VDD.n451 2.2755
R1410 VDD.n127 VDD.t330 2.2755
R1411 VDD.n127 VDD.n126 2.2755
R1412 VDD.n490 VDD.t24 2.2755
R1413 VDD.n490 VDD.n489 2.2755
R1414 VDD.n487 VDD.t88 2.2755
R1415 VDD.n487 VDD.n486 2.2755
R1416 VDD.n10 VDD.t192 2.2755
R1417 VDD.n10 VDD.n9 2.2755
R1418 VDD.n23 VDD.t272 2.2755
R1419 VDD.n23 VDD.n22 2.2755
R1420 VDD.n20 VDD.t265 2.2755
R1421 VDD.n20 VDD.n19 2.2755
R1422 VDD.n93 VDD.t445 2.2755
R1423 VDD.n93 VDD.n92 2.2755
R1424 VDD.n90 VDD.t54 2.2755
R1425 VDD.n90 VDD.n89 2.2755
R1426 VDD.n2 VDD.t38 2.2755
R1427 VDD.n2 VDD.n1 2.2755
R1428 VDD.n321 VDD.n320 2.2439
R1429 VDD.n333 VDD.n332 2.2439
R1430 VDD.n42 VDD.n41 2.2439
R1431 VDD.n52 VDD.n51 2.2439
R1432 VDD.n315 VDD.n314 2.24362
R1433 VDD.n31 VDD.n30 2.24362
R1434 VDD.n313 VDD.n312 2.12269
R1435 VDD.n28 VDD.n27 2.12257
R1436 VDD.n325 VDD.n324 1.82213
R1437 VDD.n335 VDD.n334 1.82213
R1438 VDD VDD.n371 1.81843
R1439 VDD.n259 VDD 1.81843
R1440 VDD.n282 VDD 1.81843
R1441 VDD.n412 VDD 1.81843
R1442 VDD.n417 VDD 1.81843
R1443 VDD.n46 VDD.n45 1.81789
R1444 VDD VDD.n229 1.77285
R1445 VDD VDD.n224 1.77285
R1446 VDD.n470 VDD 1.77285
R1447 VDD.n505 VDD 1.77285
R1448 VDD VDD.n8 1.77285
R1449 VDD.n43 VDD.n42 1.62565
R1450 VDD.n53 VDD.n52 1.62565
R1451 VDD.n336 VDD.n333 1.6239
R1452 VDD.n326 VDD.n321 1.6239
R1453 VDD.n331 VDD.n330 1.39892
R1454 VDD.n319 VDD.n318 1.3985
R1455 VDD.n49 VDD.n48 1.39782
R1456 VDD.n39 VDD.n38 1.39728
R1457 VDD.n69 VDD.n68 1.16167
R1458 VDD.n360 VDD.n359 1.16051
R1459 VDD.n326 VDD.n325 1.12224
R1460 VDD.n43 VDD.n36 1.12171
R1461 VDD.n53 VDD.n46 1.12171
R1462 VDD.n336 VDD.n335 1.12167
R1463 VDD.n468 VDD.n467 1.07428
R1464 VDD.n503 VDD.n502 1.07428
R1465 VDD.n106 VDD.n105 1.07428
R1466 VDD.n396 VDD.n395 1.0737
R1467 VDD.n256 VDD.n201 1.0737
R1468 VDD.n279 VDD.n175 1.0737
R1469 VDD.n35 VDD.n33 0.840632
R1470 VDD.n407 VDD.n406 0.715235
R1471 VDD.n342 VDD.n340 0.603658
R1472 VDD.n337 VDD.n336 0.523557
R1473 VDD.n54 VDD.n53 0.5228
R1474 VDD.n327 VDD.n315 0.497812
R1475 VDD.n44 VDD.n31 0.497812
R1476 VDD.n233 VDD 0.434967
R1477 VDD.n324 VDD.n323 0.404541
R1478 VDD.n436 VDD 0.339236
R1479 VDD VDD.n216 0.338387
R1480 VDD.n346 VDD.n342 0.337997
R1481 VDD.n58 VDD.n57 0.337997
R1482 VDD VDD.n219 0.334577
R1483 VDD.n422 VDD 0.334577
R1484 VDD.n57 VDD.n56 0.333658
R1485 VDD.n425 VDD.n424 0.318198
R1486 VDD.n218 VDD.n217 0.317357
R1487 VDD VDD.n0 0.280768
R1488 VDD.n345 VDD.n309 0.233919
R1489 VDD.n351 VDD.n350 0.233919
R1490 VDD.n381 VDD.n377 0.233919
R1491 VDD.n387 VDD.n386 0.233919
R1492 VDD.n187 VDD.n183 0.233919
R1493 VDD.n193 VDD.n192 0.233919
R1494 VDD.n161 VDD.n157 0.233919
R1495 VDD.n167 VDD.n166 0.233919
R1496 VDD.n462 VDD.n461 0.233919
R1497 VDD.n459 VDD.n458 0.233919
R1498 VDD.n497 VDD.n496 0.233919
R1499 VDD.n494 VDD.n493 0.233919
R1500 VDD.n63 VDD.n62 0.233919
R1501 VDD.n60 VDD.n59 0.233919
R1502 VDD.n100 VDD.n99 0.233919
R1503 VDD.n97 VDD.n96 0.233919
R1504 VDD.n408 VDD.n148 0.170499
R1505 VDD.n413 VDD.n145 0.170499
R1506 VDD.n418 VDD.n142 0.170499
R1507 VDD.n232 VDD.n231 0.170231
R1508 VDD.n227 VDD.n226 0.170231
R1509 VDD.n222 VDD.n221 0.170231
R1510 VDD.n217 VDD 0.147133
R1511 VDD.n424 VDD 0.146292
R1512 VDD.n397 VDD.n396 0.143967
R1513 VDD.n256 VDD.n255 0.143967
R1514 VDD.n279 VDD.n278 0.143967
R1515 VDD.n468 VDD.n446 0.143501
R1516 VDD.n503 VDD.n481 0.143501
R1517 VDD.n107 VDD.n106 0.143501
R1518 VDD.n354 VDD.n353 0.141016
R1519 VDD.n366 VDD.n365 0.141016
R1520 VDD.n363 VDD.n362 0.141016
R1521 VDD.n390 VDD.n389 0.141016
R1522 VDD.n247 VDD.n246 0.141016
R1523 VDD.n250 VDD.n249 0.141016
R1524 VDD.n196 VDD.n195 0.141016
R1525 VDD.n270 VDD.n269 0.141016
R1526 VDD.n273 VDD.n272 0.141016
R1527 VDD.n170 VDD.n169 0.141016
R1528 VDD.n403 VDD.n402 0.141016
R1529 VDD.n400 VDD.n399 0.141016
R1530 VDD.n444 VDD.n443 0.141016
R1531 VDD.n441 VDD.n440 0.141016
R1532 VDD.n465 VDD.n464 0.141016
R1533 VDD.n479 VDD.n478 0.141016
R1534 VDD.n476 VDD.n475 0.141016
R1535 VDD.n500 VDD.n499 0.141016
R1536 VDD.n66 VDD.n65 0.141016
R1537 VDD.n73 VDD.n72 0.141016
R1538 VDD.n74 VDD.n12 0.141016
R1539 VDD.n103 VDD.n102 0.141016
R1540 VDD.n108 VDD.n6 0.141016
R1541 VDD.n114 VDD.n113 0.141016
R1542 VDD.n396 VDD.n372 0.139745
R1543 VDD.n280 VDD.n279 0.139745
R1544 VDD.n504 VDD.n503 0.138896
R1545 VDD.n106 VDD.n84 0.138896
R1546 VDD.n257 VDD 0.128708
R1547 VDD.n469 VDD 0.127858
R1548 VDD VDD.n368 0.123016
R1549 VDD VDD.n212 0.123016
R1550 VDD VDD.n263 0.123016
R1551 VDD.n438 VDD 0.122435
R1552 VDD.n473 VDD 0.122435
R1553 VDD VDD.n79 0.122435
R1554 VDD.n335 VDD 0.112066
R1555 VDD VDD.n472 0.111984
R1556 VDD.n80 VDD 0.111984
R1557 VDD VDD.n507 0.111984
R1558 VDD.n340 VDD 0.111564
R1559 VDD.n369 VDD 0.111403
R1560 VDD.n264 VDD 0.111403
R1561 VDD.n285 VDD 0.111403
R1562 VDD.n46 VDD 0.110941
R1563 VDD VDD.n437 0.108832
R1564 VDD.n215 VDD 0.108613
R1565 VDD.n355 VDD.n354 0.107339
R1566 VDD.n359 VDD.n358 0.107339
R1567 VDD.n367 VDD.n366 0.107339
R1568 VDD.n364 VDD.n363 0.107339
R1569 VDD.n361 VDD.n360 0.107339
R1570 VDD.n391 VDD.n390 0.107339
R1571 VDD.n395 VDD.n394 0.107339
R1572 VDD.n234 VDD.n232 0.107339
R1573 VDD.n228 VDD.n227 0.107339
R1574 VDD.n223 VDD.n222 0.107339
R1575 VDD.n246 VDD.n245 0.107339
R1576 VDD.n251 VDD.n250 0.107339
R1577 VDD.n255 VDD.n254 0.107339
R1578 VDD.n197 VDD.n196 0.107339
R1579 VDD.n201 VDD.n200 0.107339
R1580 VDD.n269 VDD.n268 0.107339
R1581 VDD.n274 VDD.n273 0.107339
R1582 VDD.n278 VDD.n277 0.107339
R1583 VDD.n171 VDD.n170 0.107339
R1584 VDD.n175 VDD.n174 0.107339
R1585 VDD.n404 VDD.n403 0.107339
R1586 VDD.n401 VDD.n400 0.107339
R1587 VDD.n398 VDD.n397 0.107339
R1588 VDD.n409 VDD.n408 0.107339
R1589 VDD.n414 VDD.n413 0.107339
R1590 VDD.n419 VDD.n418 0.107339
R1591 VDD.n446 VDD.n445 0.107339
R1592 VDD.n443 VDD.n442 0.107339
R1593 VDD.n440 VDD.n439 0.107339
R1594 VDD.n467 VDD.n466 0.107339
R1595 VDD.n464 VDD.n463 0.107339
R1596 VDD.n481 VDD.n480 0.107339
R1597 VDD.n478 VDD.n477 0.107339
R1598 VDD.n475 VDD.n474 0.107339
R1599 VDD.n502 VDD.n501 0.107339
R1600 VDD.n499 VDD.n498 0.107339
R1601 VDD.n68 VDD.n67 0.107339
R1602 VDD.n65 VDD.n64 0.107339
R1603 VDD.n71 VDD.n69 0.107339
R1604 VDD.n75 VDD.n73 0.107339
R1605 VDD.n78 VDD.n12 0.107339
R1606 VDD.n105 VDD.n104 0.107339
R1607 VDD.n102 VDD.n101 0.107339
R1608 VDD.n109 VDD.n107 0.107339
R1609 VDD.n112 VDD.n6 0.107339
R1610 VDD.n116 VDD.n114 0.107339
R1611 VDD VDD.n345 0.106758
R1612 VDD.n350 VDD 0.106758
R1613 VDD VDD.n369 0.106758
R1614 VDD VDD.n381 0.106758
R1615 VDD.n386 VDD 0.106758
R1616 VDD VDD.n187 0.106758
R1617 VDD.n192 VDD 0.106758
R1618 VDD VDD.n264 0.106758
R1619 VDD VDD.n161 0.106758
R1620 VDD.n166 VDD 0.106758
R1621 VDD VDD.n285 0.106758
R1622 VDD.n461 VDD 0.106177
R1623 VDD.n458 VDD 0.106177
R1624 VDD.n472 VDD 0.106177
R1625 VDD.n496 VDD 0.106177
R1626 VDD.n493 VDD 0.106177
R1627 VDD.n62 VDD 0.106177
R1628 VDD.n59 VDD 0.106177
R1629 VDD VDD.n80 0.106177
R1630 VDD.n99 VDD 0.106177
R1631 VDD.n96 VDD 0.106177
R1632 VDD.n507 VDD 0.106177
R1633 VDD.n322 VDD 0.0850665
R1634 VDD.n34 VDD 0.0839415
R1635 VDD.n406 VDD 0.0829516
R1636 VDD VDD.n0 0.082371
R1637 VDD.n317 VDD 0.0816915
R1638 VDD.n40 VDD 0.0816915
R1639 VDD.n349 VDD.n309 0.080629
R1640 VDD.n371 VDD.n370 0.080629
R1641 VDD.n385 VDD.n377 0.080629
R1642 VDD.n191 VDD.n183 0.080629
R1643 VDD.n265 VDD.n259 0.080629
R1644 VDD.n165 VDD.n157 0.080629
R1645 VDD.n286 VDD.n282 0.080629
R1646 VDD.n460 VDD.n459 0.080629
R1647 VDD.n471 VDD.n470 0.080629
R1648 VDD.n495 VDD.n494 0.080629
R1649 VDD.n61 VDD.n60 0.080629
R1650 VDD.n81 VDD.n8 0.080629
R1651 VDD.n98 VDD.n97 0.080629
R1652 VDD.n506 VDD.n505 0.080629
R1653 VDD.n329 VDD 0.0805665
R1654 VDD.n50 VDD 0.0805665
R1655 VDD VDD.n444 0.0794677
R1656 VDD VDD.n441 0.0794677
R1657 VDD VDD.n438 0.0794677
R1658 VDD VDD.n465 0.0794677
R1659 VDD VDD.n462 0.0794677
R1660 VDD VDD.n479 0.0794677
R1661 VDD VDD.n476 0.0794677
R1662 VDD VDD.n473 0.0794677
R1663 VDD VDD.n500 0.0794677
R1664 VDD VDD.n497 0.0794677
R1665 VDD VDD.n66 0.0794677
R1666 VDD VDD.n63 0.0794677
R1667 VDD.n72 VDD 0.0794677
R1668 VDD VDD.n74 0.0794677
R1669 VDD.n79 VDD 0.0794677
R1670 VDD VDD.n103 0.0794677
R1671 VDD VDD.n100 0.0794677
R1672 VDD VDD.n108 0.0794677
R1673 VDD.n113 VDD 0.0794677
R1674 VDD VDD.n115 0.0794677
R1675 VDD.n219 VDD 0.0794623
R1676 VDD VDD.n422 0.0794623
R1677 VDD VDD.n351 0.0788871
R1678 VDD.n353 VDD 0.0788871
R1679 VDD.n368 VDD 0.0788871
R1680 VDD.n365 VDD 0.0788871
R1681 VDD.n362 VDD 0.0788871
R1682 VDD VDD.n387 0.0788871
R1683 VDD.n389 VDD 0.0788871
R1684 VDD.n212 VDD 0.0788871
R1685 VDD VDD.n247 0.0788871
R1686 VDD.n249 VDD 0.0788871
R1687 VDD VDD.n193 0.0788871
R1688 VDD.n195 VDD 0.0788871
R1689 VDD.n263 VDD 0.0788871
R1690 VDD VDD.n270 0.0788871
R1691 VDD.n272 VDD 0.0788871
R1692 VDD VDD.n167 0.0788871
R1693 VDD.n169 VDD 0.0788871
R1694 VDD.n405 VDD 0.0788871
R1695 VDD.n402 VDD 0.0788871
R1696 VDD.n399 VDD 0.0788871
R1697 VDD VDD.n233 0.0759839
R1698 VDD.n229 VDD 0.0759839
R1699 VDD.n224 VDD 0.0759839
R1700 VDD VDD.n407 0.0754032
R1701 VDD VDD.n412 0.0754032
R1702 VDD VDD.n417 0.0754032
R1703 VDD.n311 VDD 0.0749415
R1704 VDD.n29 VDD 0.0738165
R1705 VDD.n56 VDD.n55 0.0725
R1706 VDD.n231 VDD 0.0709717
R1707 VDD.n226 VDD 0.0709717
R1708 VDD.n221 VDD 0.0709717
R1709 VDD VDD.n469 0.0709717
R1710 VDD VDD.n504 0.0709717
R1711 VDD.n84 VDD 0.0709717
R1712 VDD.n372 VDD 0.0701226
R1713 VDD VDD.n257 0.0701226
R1714 VDD VDD.n280 0.0701226
R1715 VDD VDD.n148 0.0701226
R1716 VDD VDD.n145 0.0701226
R1717 VDD VDD.n142 0.0701226
R1718 VDD.n56 VDD 0.0493298
R1719 VDD.n216 VDD 0.0491131
R1720 VDD.n436 VDD 0.0487847
R1721 VDD.n208 VDD.n207 0.0409015
R1722 VDD.n433 VDD.n432 0.040573
R1723 VDD.n406 VDD.n405 0.0405645
R1724 VDD.n115 VDD.n0 0.0405645
R1725 VDD.n340 VDD.n339 0.0344894
R1726 VDD.n320 VDD.n317 0.0275
R1727 VDD.n325 VDD.n322 0.0275
R1728 VDD.n41 VDD.n40 0.0275
R1729 VDD.n34 VDD.n32 0.0275
R1730 VDD.n332 VDD.n329 0.026375
R1731 VDD.n51 VDD.n50 0.026375
R1732 VDD.n321 VDD.n316 0.025705
R1733 VDD.n333 VDD.n328 0.025705
R1734 VDD.n42 VDD.n37 0.025705
R1735 VDD.n52 VDD.n47 0.025705
R1736 VDD.n209 VDD.n208 0.025135
R1737 VDD.n434 VDD.n433 0.025135
R1738 VDD.n210 VDD.n209 0.0211934
R1739 VDD.n435 VDD.n434 0.0211934
R1740 VDD.n30 VDD.n29 0.02075
R1741 VDD.n314 VDD.n311 0.019625
R1742 VDD.n315 VDD.n310 0.0169383
R1743 VDD.n31 VDD.n26 0.0169383
R1744 VDD.n437 VDD.n436 0.0132147
R1745 VDD.n216 VDD.n215 0.0131133
R1746 VDD VDD.n256 0.0115377
R1747 VDD VDD.n468 0.0115377
R1748 VDD.n314 VDD.n313 0.010625
R1749 VDD.n30 VDD.n28 0.0095
R1750 VDD.n409 VDD 0.00572581
R1751 VDD.n414 VDD 0.00572581
R1752 VDD.n419 VDD 0.00572581
R1753 VDD.n234 VDD 0.00514516
R1754 VDD VDD.n228 0.00514516
R1755 VDD VDD.n223 0.00514516
R1756 VDD.n332 VDD.n331 0.003875
R1757 VDD.n51 VDD.n49 0.003875
R1758 VDD.n320 VDD.n319 0.00275
R1759 VDD.n41 VDD.n39 0.00275
R1760 VDD.n355 VDD 0.00224194
R1761 VDD.n358 VDD 0.00224194
R1762 VDD VDD.n367 0.00224194
R1763 VDD VDD.n364 0.00224194
R1764 VDD VDD.n361 0.00224194
R1765 VDD.n391 VDD 0.00224194
R1766 VDD.n394 VDD 0.00224194
R1767 VDD.n245 VDD 0.00224194
R1768 VDD.n251 VDD 0.00224194
R1769 VDD.n254 VDD 0.00224194
R1770 VDD.n197 VDD 0.00224194
R1771 VDD.n200 VDD 0.00224194
R1772 VDD.n268 VDD 0.00224194
R1773 VDD.n274 VDD 0.00224194
R1774 VDD.n277 VDD 0.00224194
R1775 VDD.n171 VDD 0.00224194
R1776 VDD.n174 VDD 0.00224194
R1777 VDD VDD.n404 0.00224194
R1778 VDD VDD.n401 0.00224194
R1779 VDD VDD.n398 0.00224194
R1780 VDD VDD.n218 0.00219811
R1781 VDD.n425 VDD 0.00219811
R1782 VDD.n445 VDD 0.00166129
R1783 VDD.n442 VDD 0.00166129
R1784 VDD.n439 VDD 0.00166129
R1785 VDD.n466 VDD 0.00166129
R1786 VDD.n463 VDD 0.00166129
R1787 VDD VDD.n460 0.00166129
R1788 VDD VDD.n457 0.00166129
R1789 VDD.n480 VDD 0.00166129
R1790 VDD.n477 VDD 0.00166129
R1791 VDD.n474 VDD 0.00166129
R1792 VDD VDD.n471 0.00166129
R1793 VDD.n501 VDD 0.00166129
R1794 VDD.n498 VDD 0.00166129
R1795 VDD VDD.n495 0.00166129
R1796 VDD VDD.n492 0.00166129
R1797 VDD.n67 VDD 0.00166129
R1798 VDD.n64 VDD 0.00166129
R1799 VDD VDD.n61 0.00166129
R1800 VDD VDD.n58 0.00166129
R1801 VDD VDD.n71 0.00166129
R1802 VDD.n75 VDD 0.00166129
R1803 VDD VDD.n78 0.00166129
R1804 VDD.n81 VDD 0.00166129
R1805 VDD.n104 VDD 0.00166129
R1806 VDD.n101 VDD 0.00166129
R1807 VDD VDD.n98 0.00166129
R1808 VDD VDD.n95 0.00166129
R1809 VDD.n109 VDD 0.00166129
R1810 VDD VDD.n112 0.00166129
R1811 VDD.n116 VDD 0.00166129
R1812 VDD VDD.n506 0.00166129
R1813 VDD.n36 VDD.n32 0.001625
R1814 VDD VDD.n435 0.00115693
R1815 VDD.n346 VDD 0.00108064
R1816 VDD VDD.n349 0.00108064
R1817 VDD.n370 VDD 0.00108064
R1818 VDD.n382 VDD 0.00108064
R1819 VDD VDD.n385 0.00108064
R1820 VDD.n188 VDD 0.00108064
R1821 VDD VDD.n191 0.00108064
R1822 VDD.n265 VDD 0.00108064
R1823 VDD.n162 VDD 0.00108064
R1824 VDD VDD.n165 0.00108064
R1825 VDD.n286 VDD 0.00108064
R1826 VDD VDD.n210 0.000828467
R1827 CLK_div_10_mag_1.Q0.n19 CLK_div_10_mag_1.Q0.t18 36.935
R1828 CLK_div_10_mag_1.Q0.n18 CLK_div_10_mag_1.Q0.t3 36.935
R1829 CLK_div_10_mag_1.Q0.n22 CLK_div_10_mag_1.Q0.t6 36.935
R1830 CLK_div_10_mag_1.Q0.n21 CLK_div_10_mag_1.Q0.t9 36.935
R1831 CLK_div_10_mag_1.Q0.n13 CLK_div_10_mag_1.Q0.t13 36.935
R1832 CLK_div_10_mag_1.Q0.n15 CLK_div_10_mag_1.Q0.t17 31.4332
R1833 CLK_div_10_mag_1.Q0.n24 CLK_div_10_mag_1.Q0.t5 30.6613
R1834 CLK_div_10_mag_1.Q0.n20 CLK_div_10_mag_1.Q0.t7 25.4744
R1835 CLK_div_10_mag_1.Q0.n26 CLK_div_10_mag_1.Q0.t10 25.4744
R1836 CLK_div_10_mag_1.Q0.n24 CLK_div_10_mag_1.Q0.t14 21.6718
R1837 CLK_div_10_mag_1.Q0.n19 CLK_div_10_mag_1.Q0.t16 18.1962
R1838 CLK_div_10_mag_1.Q0.n18 CLK_div_10_mag_1.Q0.t19 18.1962
R1839 CLK_div_10_mag_1.Q0.n22 CLK_div_10_mag_1.Q0.t4 18.1962
R1840 CLK_div_10_mag_1.Q0.n21 CLK_div_10_mag_1.Q0.t8 18.1962
R1841 CLK_div_10_mag_1.Q0.n13 CLK_div_10_mag_1.Q0.t12 18.1962
R1842 CLK_div_10_mag_1.Q0.n15 CLK_div_10_mag_1.Q0.t15 15.3826
R1843 CLK_div_10_mag_1.Q0.n26 CLK_div_10_mag_1.Q0.t20 14.1417
R1844 CLK_div_10_mag_1.Q0.n20 CLK_div_10_mag_1.Q0.t11 14.1417
R1845 CLK_div_10_mag_1.Q0.n0 CLK_div_10_mag_1.Q0.n25 9.9005
R1846 CLK_div_10_mag_1.Q0.n12 CLK_div_10_mag_1.Q0.t2 7.09905
R1847 CLK_div_10_mag_1.Q0.n16 CLK_div_10_mag_1.Q0.n15 6.86029
R1848 CLK_div_10_mag_1.Q0.n17 CLK_div_10_mag_1.Q0.n14 5.01077
R1849 CLK_div_10_mag_1.Q0.n2 CLK_div_10_mag_1.Q0.n3 1.11863
R1850 CLK_div_10_mag_1.Q0.n4 CLK_div_10_mag_1.Q0.n5 1.11863
R1851 CLK_div_10_mag_1.Q0.n20 CLK_div_10_mag_1.Q0.n9 1.42995
R1852 CLK_div_10_mag_1.Q0.n0 CLK_div_10_mag_1.Q0.n1 1.11781
R1853 CLK_div_10_mag_1.Q0.n12 CLK_div_10_mag_1.Q0.n11 3.25053
R1854 CLK_div_10_mag_1.Q0.n11 CLK_div_10_mag_1.Q0.t0 2.2755
R1855 CLK_div_10_mag_1.Q0.n11 CLK_div_10_mag_1.Q0.n10 2.2755
R1856 CLK_div_10_mag_1.Q0.n28 CLK_div_10_mag_1.Q0.n27 2.2505
R1857 CLK_div_10_mag_1.Q0.n23 CLK_div_10_mag_1.Q0.n9 1.16587
R1858 CLK_div_10_mag_1.Q0.n14 CLK_div_10_mag_1.Q0.n13 2.13459
R1859 CLK_div_10_mag_1.Q0.n3 CLK_div_10_mag_1.Q0.n19 2.13265
R1860 CLK_div_10_mag_1.Q0.n5 CLK_div_10_mag_1.Q0.n22 2.13265
R1861 CLK_div_10_mag_1.Q0.n2 CLK_div_10_mag_1.Q0.n7 2.63776
R1862 CLK_div_10_mag_1.Q0.n4 CLK_div_10_mag_1.Q0.n8 2.63776
R1863 CLK_div_10_mag_1.Q0.n27 CLK_div_10_mag_1.Q0.n17 1.52773
R1864 CLK_div_10_mag_1.Q0.n18 CLK_div_10_mag_1.Q0.n7 2.13261
R1865 CLK_div_10_mag_1.Q0.n21 CLK_div_10_mag_1.Q0.n8 2.13281
R1866 CLK_div_10_mag_1.Q0.n1 CLK_div_10_mag_1.Q0.n26 1.42999
R1867 CLK_div_10_mag_1.Q0.n6 CLK_div_10_mag_1.Q0.n24 1.41101
R1868 CLK_div_10_mag_1.Q0.n17 CLK_div_10_mag_1.Q0.n16 1.12067
R1869 CLK_div_10_mag_1.Q0.n25 CLK_div_10_mag_1.Q0.n23 0.286289
R1870 CLK_div_10_mag_1.Q0.n1 CLK_div_10_mag_1.Q0 0.196008
R1871 CLK_div_10_mag_1.Q0.n9 CLK_div_10_mag_1.Q0 0.196051
R1872 CLK_div_10_mag_1.Q0.n28 CLK_div_10_mag_1.Q0.n12 0.0905
R1873 CLK_div_10_mag_1.Q0.n16 CLK_div_10_mag_1.Q0 0.0857632
R1874 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.Q0.n28 0.0834687
R1875 CLK_div_10_mag_1.Q0.n6 CLK_div_10_mag_1.Q0 0.104828
R1876 CLK_div_10_mag_1.Q0.n14 CLK_div_10_mag_1.Q0 0.0800273
R1877 CLK_div_10_mag_1.Q0.n8 CLK_div_10_mag_1.Q0 0.0771461
R1878 CLK_div_10_mag_1.Q0.n7 CLK_div_10_mag_1.Q0 0.0771461
R1879 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.Q0.n5 0.077103
R1880 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.Q0.n3 0.077103
R1881 CLK_div_10_mag_1.Q0.n27 CLK_div_10_mag_1.Q0 0.0289903
R1882 CLK_div_10_mag_1.Q0.n25 CLK_div_10_mag_1.Q0.n6 7.13895
R1883 CLK_div_10_mag_1.Q0.n0 CLK_div_10_mag_1.Q0.n2 1.18681
R1884 CLK_div_10_mag_1.Q0.n23 CLK_div_10_mag_1.Q0.n4 0.938524
R1885 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.Q0.n0 0.680217
R1886 Vdiv100.n2 Vdiv100.t1 9.28805
R1887 Vdiv100.n1 Vdiv100.n0 6.01414
R1888 Vdiv100.n1 Vdiv100.t3 6.01414
R1889 Vdiv100.n3 Vdiv100.t2 3.87536
R1890 Vdiv100.n2 Vdiv100.n1 3.74829
R1891 Vdiv100.n3 Vdiv100.n2 0.0409348
R1892 Vdiv100 Vdiv100.n3 0.0031087
R1893 CLK.n9 CLK.t0 36.935
R1894 CLK.n3 CLK.t1 36.935
R1895 CLK.n14 CLK.t3 25.5361
R1896 CLK.n9 CLK.t2 18.1962
R1897 CLK.n3 CLK.t5 18.1962
R1898 CLK.n14 CLK.t4 14.0734
R1899 CLK.n5 CLK.n2 4.5005
R1900 CLK.n5 CLK.n4 4.5005
R1901 CLK.n8 CLK.n7 4.5005
R1902 CLK.n10 CLK.n7 4.5005
R1903 CLK.n16 CLK.n15 4.5005
R1904 CLK.n17 CLK.n16 4.5005
R1905 CLK.n12 CLK.n11 2.25107
R1906 CLK.n13 CLK.n0 2.24235
R1907 CLK.n4 CLK.n3 2.12175
R1908 CLK.n10 CLK.n9 2.12075
R1909 CLK.n7 CLK.n6 1.74297
R1910 CLK.n6 CLK.n1 1.49778
R1911 CLK.n15 CLK.n14 1.42775
R1912 CLK.n13 CLK.n12 0.97145
R1913 CLK CLK.n17 0.1355
R1914 CLK.n8 CLK 0.0473512
R1915 CLK.n2 CLK 0.0473512
R1916 CLK.n11 CLK.n8 0.0361897
R1917 CLK.n2 CLK.n1 0.0361897
R1918 CLK.n17 CLK.n0 0.03175
R1919 CLK.n16 CLK.n13 0.0246174
R1920 CLK.n6 CLK.n5 0.0131772
R1921 CLK.n12 CLK.n7 0.0122182
R1922 CLK.n11 CLK.n10 0.00515517
R1923 CLK.n4 CLK.n1 0.00515517
R1924 CLK.n15 CLK.n0 0.00175
R1925 RST.n27 RST.t15 37.2596
R1926 RST.n0 RST.t5 36.935
R1927 RST.n22 RST.t1 36.935
R1928 RST.n29 RST.t12 36.935
R1929 RST.n15 RST.t6 36.935
R1930 RST.n13 RST.t13 36.935
R1931 RST.n2 RST.t7 36.935
R1932 RST.n8 RST.t9 36.859
R1933 RST.n0 RST.t3 18.1962
R1934 RST.n22 RST.t0 18.1962
R1935 RST.n29 RST.t11 18.1962
R1936 RST.n15 RST.t2 18.1962
R1937 RST.n13 RST.t10 18.1962
R1938 RST.n2 RST.t4 18.1962
R1939 RST.n27 RST.t14 17.5947
R1940 RST.n7 RST.t8 17.236
R1941 RST.n33 RST.n19 6.72677
R1942 RST.n17 RST.n16 5.39891
R1943 RST.n12 RST.n11 4.5005
R1944 RST.n6 RST.n5 4.5005
R1945 RST.n12 RST.n4 4.5005
R1946 RST.n7 RST.n4 3.60685
R1947 RST.n18 RST.n17 3.52872
R1948 RST.n33 RST.n32 3.52871
R1949 RST.n32 RST.n31 3.52813
R1950 RST.n31 RST 3.47503
R1951 RST RST.n18 3.47443
R1952 RST.n9 RST.n8 2.88526
R1953 RST.n16 RST.n15 2.13713
R1954 RST.n14 RST.n13 2.13713
R1955 RST.n30 RST.n29 2.13592
R1956 RST.n3 RST.n2 2.1349
R1957 RST.n23 RST.n22 2.12075
R1958 RST.n1 RST.n0 2.12075
R1959 RST.n17 RST.n14 1.87041
R1960 RST.n31 RST.n28 1.8703
R1961 RST RST.n30 1.81628
R1962 RST.n19 RST.n3 1.76851
R1963 RST.n36 RST.n35 1.51229
R1964 RST.n10 RST.n5 1.51223
R1965 RST.n25 RST.n24 1.51214
R1966 RST.n28 RST.n27 1.43806
R1967 RST.n34 RST.n33 1.12379
R1968 RST.n18 RST.n12 1.12371
R1969 RST.n32 RST.n26 1.1235
R1970 RST.n8 RST.n7 0.865351
R1971 RST.n30 RST 0.0704961
R1972 RST.n3 RST 0.0687763
R1973 RST.n14 RST 0.06755
R1974 RST.n16 RST 0.0675495
R1975 RST.n28 RST 0.0659998
R1976 RST.n19 RST 0.0484016
R1977 RST.n20 RST 0.0394837
R1978 RST.n6 RST 0.0394837
R1979 RST RST.n39 0.0383947
R1980 RST.n37 RST.n36 0.0377319
R1981 RST.n24 RST.n21 0.0377318
R1982 RST.n11 RST.n10 0.0367013
R1983 RST.n39 RST.n38 0.028431
R1984 RST.n39 RST 0.0194474
R1985 RST.n10 RST.n9 0.0051456
R1986 RST.n24 RST.n23 0.00438036
R1987 RST.n36 RST.n1 0.00438025
R1988 RST.n35 RST.n34 0.00391772
R1989 RST.n26 RST.n25 0.003875
R1990 RST.n12 RST.n5 0.003875
R1991 RST.n21 RST.n20 0.00205172
R1992 RST.n11 RST.n6 0.00205172
R1993 RST.n38 RST.n37 0.00205172
R1994 RST.n9 RST.n4 0.00199457
R1995 CLK_div_10_mag_0.JK_FF_mag_2.J.n2 CLK_div_10_mag_0.JK_FF_mag_2.J.t6 37.1986
R1996 CLK_div_10_mag_0.JK_FF_mag_2.J.n1 CLK_div_10_mag_0.JK_FF_mag_2.J.t5 31.528
R1997 CLK_div_10_mag_0.JK_FF_mag_2.J.n3 CLK_div_10_mag_0.JK_FF_mag_2.J.t3 30.6315
R1998 CLK_div_10_mag_0.JK_FF_mag_2.J.n3 CLK_div_10_mag_0.JK_FF_mag_2.J.t7 24.5953
R1999 CLK_div_10_mag_0.JK_FF_mag_2.J.n2 CLK_div_10_mag_0.JK_FF_mag_2.J.t8 17.6614
R2000 CLK_div_10_mag_0.JK_FF_mag_2.J.n4 CLK_div_10_mag_0.JK_FF_mag_2.J 17.0516
R2001 CLK_div_10_mag_0.JK_FF_mag_2.J.n1 CLK_div_10_mag_0.JK_FF_mag_2.J.t4 15.3826
R2002 CLK_div_10_mag_0.JK_FF_mag_2.J CLK_div_10_mag_0.JK_FF_mag_2.J.n1 7.62751
R2003 CLK_div_10_mag_0.JK_FF_mag_2.J.n5 CLK_div_10_mag_0.JK_FF_mag_2.J.n4 3.28711
R2004 CLK_div_10_mag_0.JK_FF_mag_2.J.n0 CLK_div_10_mag_0.JK_FF_mag_2.J.n7 2.99416
R2005 CLK_div_10_mag_0.JK_FF_mag_2.J.n4 CLK_div_10_mag_0.JK_FF_mag_2.J 2.81128
R2006 CLK_div_10_mag_0.JK_FF_mag_2.J.n5 CLK_div_10_mag_0.JK_FF_mag_2.J 2.67866
R2007 CLK_div_10_mag_0.JK_FF_mag_2.J.n7 CLK_div_10_mag_0.JK_FF_mag_2.J.t0 2.2755
R2008 CLK_div_10_mag_0.JK_FF_mag_2.J.n7 CLK_div_10_mag_0.JK_FF_mag_2.J.n6 2.2755
R2009 CLK_div_10_mag_0.JK_FF_mag_2.J.n0 CLK_div_10_mag_0.JK_FF_mag_2.J.n5 2.2505
R2010 CLK_div_10_mag_0.JK_FF_mag_2.J CLK_div_10_mag_0.JK_FF_mag_2.J.n3 1.80496
R2011 CLK_div_10_mag_0.JK_FF_mag_2.J CLK_div_10_mag_0.JK_FF_mag_2.J.n2 1.43709
R2012 CLK_div_10_mag_0.JK_FF_mag_2.J CLK_div_10_mag_0.JK_FF_mag_2.J.n0 0.281955
R2013 CLK_div_10_mag_1.Q2.n2 CLK_div_10_mag_1.Q2.t10 36.935
R2014 CLK_div_10_mag_1.Q2.n6 CLK_div_10_mag_1.Q2.t8 31.4332
R2015 CLK_div_10_mag_1.Q2.n8 CLK_div_10_mag_1.Q2.t12 31.4332
R2016 CLK_div_10_mag_1.Q2.n3 CLK_div_10_mag_1.Q2.t4 31.4332
R2017 CLK_div_10_mag_1.Q2.n5 CLK_div_10_mag_1.Q2.t7 30.5752
R2018 CLK_div_10_mag_1.Q2.n5 CLK_div_10_mag_1.Q2.t6 21.7814
R2019 CLK_div_10_mag_1.Q2.n2 CLK_div_10_mag_1.Q2.t9 18.1962
R2020 CLK_div_10_mag_1.Q2.n6 CLK_div_10_mag_1.Q2.t11 15.3826
R2021 CLK_div_10_mag_1.Q2.n8 CLK_div_10_mag_1.Q2.t5 15.3826
R2022 CLK_div_10_mag_1.Q2.n3 CLK_div_10_mag_1.Q2.t3 15.3826
R2023 CLK_div_10_mag_1.Q2 CLK_div_10_mag_1.Q2.t1 7.09905
R2024 CLK_div_10_mag_1.Q2 CLK_div_10_mag_1.Q2.n8 6.86658
R2025 CLK_div_10_mag_1.Q2 CLK_div_10_mag_1.Q2.n6 6.86658
R2026 CLK_div_10_mag_1.Q2 CLK_div_10_mag_1.Q2.n3 6.86029
R2027 CLK_div_10_mag_1.Q2.n9 CLK_div_10_mag_1.Q2 5.61266
R2028 CLK_div_10_mag_1.Q2.n4 CLK_div_10_mag_1.Q2 5.01077
R2029 CLK_div_10_mag_1.Q2 CLK_div_10_mag_1.Q2.n1 3.25053
R2030 CLK_div_10_mag_1.Q2.n7 CLK_div_10_mag_1.Q2 3.01024
R2031 CLK_div_10_mag_1.Q2.n9 CLK_div_10_mag_1.Q2.n7 2.84996
R2032 CLK_div_10_mag_1.Q2 CLK_div_10_mag_1.Q2.n10 2.34645
R2033 CLK_div_10_mag_1.Q2.n1 CLK_div_10_mag_1.Q2.t0 2.2755
R2034 CLK_div_10_mag_1.Q2.n1 CLK_div_10_mag_1.Q2.n0 2.2755
R2035 CLK_div_10_mag_1.Q2 CLK_div_10_mag_1.Q2.n2 2.13459
R2036 CLK_div_10_mag_1.Q2 CLK_div_10_mag_1.Q2.n5 1.80883
R2037 CLK_div_10_mag_1.Q2.n7 CLK_div_10_mag_1.Q2 1.67882
R2038 CLK_div_10_mag_1.Q2.n10 CLK_div_10_mag_1.Q2.n4 1.5246
R2039 CLK_div_10_mag_1.Q2.n10 CLK_div_10_mag_1.Q2.n9 1.44585
R2040 CLK_div_10_mag_1.Q2.n4 CLK_div_10_mag_1.Q2 1.12067
R2041 CLK_div_10_mag_1.JK_FF_mag_2.J.n3 CLK_div_10_mag_1.JK_FF_mag_2.J.t4 37.1981
R2042 CLK_div_10_mag_1.JK_FF_mag_2.J.n5 CLK_div_10_mag_1.JK_FF_mag_2.J.t5 31.4332
R2043 CLK_div_10_mag_1.JK_FF_mag_2.J.n2 CLK_div_10_mag_1.JK_FF_mag_2.J.t6 30.5752
R2044 CLK_div_10_mag_1.JK_FF_mag_2.J.n2 CLK_div_10_mag_1.JK_FF_mag_2.J.t7 24.6493
R2045 CLK_div_10_mag_1.JK_FF_mag_2.J.n3 CLK_div_10_mag_1.JK_FF_mag_2.J.t2 17.6611
R2046 CLK_div_10_mag_1.JK_FF_mag_2.J.n4 CLK_div_10_mag_1.JK_FF_mag_2.J 17.0516
R2047 CLK_div_10_mag_1.JK_FF_mag_2.J.n5 CLK_div_10_mag_1.JK_FF_mag_2.J.t3 15.3826
R2048 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.JK_FF_mag_2.J.n5 7.62776
R2049 CLK_div_10_mag_1.JK_FF_mag_2.J.n6 CLK_div_10_mag_1.JK_FF_mag_2.J.n4 3.28711
R2050 CLK_div_10_mag_1.JK_FF_mag_2.J.n7 CLK_div_10_mag_1.JK_FF_mag_2.J.n1 2.99416
R2051 CLK_div_10_mag_1.JK_FF_mag_2.J.n4 CLK_div_10_mag_1.JK_FF_mag_2.J 2.81128
R2052 CLK_div_10_mag_1.JK_FF_mag_2.J.n6 CLK_div_10_mag_1.JK_FF_mag_2.J 2.67895
R2053 CLK_div_10_mag_1.JK_FF_mag_2.J.n1 CLK_div_10_mag_1.JK_FF_mag_2.J.t1 2.2755
R2054 CLK_div_10_mag_1.JK_FF_mag_2.J.n1 CLK_div_10_mag_1.JK_FF_mag_2.J.n0 2.2755
R2055 CLK_div_10_mag_1.JK_FF_mag_2.J.n7 CLK_div_10_mag_1.JK_FF_mag_2.J.n6 2.2505
R2056 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.JK_FF_mag_2.J.n2 1.80883
R2057 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.JK_FF_mag_2.J.n3 1.43706
R2058 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.JK_FF_mag_2.J.n7 0.4325
C0 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_3645_212# 1.17e-20
C1 RST CLK 0.00772f
C2 a_11691_256# CLK_div_10_mag_0.JK_FF_mag_2.J 0.0811f
C3 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_1559_4126# 0.0697f
C4 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_1.JK_FF_mag_2.J 0.25f
C5 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 0.109f
C6 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_0.and2_mag_0.OUT 5.05e-20
C7 RST a_7546_212# 0.00186f
C8 a_230_2335# CLK_div_10_mag_1.nor_3_mag_0.IN3 2.44e-20
C9 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_1512_212# 8.64e-19
C10 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT 0.00395f
C11 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.00335f
C12 CLK_div_10_mag_1.Q0 a_7593_4126# 6.43e-21
C13 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C14 a_9482_4126# CLK_div_10_mag_0.and2_mag_0.OUT 2.05e-19
C15 a_4422_5223# a_4582_5223# 0.0504f
C16 CLK_div_10_mag_1.JK_FF_mag_2.J a_1559_4126# 3.25e-19
C17 CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_10_mag_1.JK_FF_mag_2.QB 2.59e-21
C18 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_1.nor_3_mag_0.IN3 4.39e-19
C19 CLK_div_10_mag_0.JK_FF_mag_1.QB a_1512_212# 0.00696f
C20 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_10_mag_1.JK_FF_mag_2.QB 0.343f
C21 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 1.29e-19
C22 CLK_div_10_mag_1.JK_FF_mag_1.QB a_10616_5223# 0.00695f
C23 CLK_div_10_mag_0.Q0 a_9510_2450# 0.01f
C24 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_3805_212# 1.46e-19
C25 a_10456_5223# CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 8.64e-19
C26 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT a_5306_5223# 0.0202f
C27 a_11180_5223# CLK_div_10_mag_1.CLK 0.00164f
C28 a_7029_4126# CLK_div_10_mag_1.Q1 6.06e-21
C29 CLK a_628_212# 0.00117f
C30 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 7.24e-19
C31 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_10_mag_1.Q3 0.338f
C32 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 9.64e-19
C33 CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.198f
C34 RST CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 0.0568f
C35 a_11127_256# CLK_div_10_mag_0.JK_FF_mag_2.J 0.00964f
C36 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_2.J 1.54e-19
C37 a_8157_4126# CLK_div_10_mag_1.JK_FF_mag_2.QB 0.00392f
C38 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 2.89e-19
C39 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD 0.994f
C40 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.0126f
C41 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_10_mag_1.Q3 0.00393f
C42 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00118f
C43 VDD CLK_div_10_mag_0.and2_mag_0.OUT 0.977f
C44 a_230_2335# CLK 4.82e-19
C45 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.and2_mag_1.OUT 0.124f
C46 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 6.82e-19
C47 VDD a_1559_4126# 3.14e-19
C48 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 8.27e-19
C49 a_9892_5223# CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.0036f
C50 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.Q3 2f
C51 CLK_div_10_mag_1.JK_FF_mag_1.QB a_10456_5223# 0.00696f
C52 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_2.J 9.73e-19
C53 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_1.Q1 0.00145f
C54 a_7956_1353# CLK_div_10_mag_0.JK_FF_mag_2.J 7.4e-19
C55 CLK_div_10_mag_0.JK_FF_mag_2.QB a_4369_212# 0.00695f
C56 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 RST 0.177f
C57 CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.16f
C58 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT a_5146_5223# 0.0731f
C59 a_6465_4126# CLK_div_10_mag_1.Q1 0.069f
C60 CLK_div_10_mag_0.Q1 a_5093_256# 0.00859f
C61 RST CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.0172f
C62 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_2.QB 2.59e-21
C63 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_1.JK_FF_mag_2.QB 0.00123f
C64 CLK_div_10_mag_0.Q2 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 3.85e-20
C65 VDD a_6822_212# 0.00891f
C66 CLK_div_10_mag_1.JK_FF_mag_0.J CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.106f
C67 CLK_div_10_mag_0.JK_FF_mag_0.J CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.106f
C68 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.00118f
C69 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.768f
C70 CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 3.38e-19
C71 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 9.9e-19
C72 a_10563_212# CLK_div_10_mag_0.JK_FF_mag_2.J 0.00696f
C73 CLK_div_10_mag_1.Q0 CLK_div_10_mag_0.JK_FF_mag_1.QB 0.00158f
C74 VDD a_9839_212# 0.00299f
C75 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.00164f
C76 RST Vdiv100 0.00303f
C77 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN a_8542_2450# 0.069f
C78 CLK_div_10_mag_1.Q0 a_6465_4126# 9.26e-19
C79 RST CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.255f
C80 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 0.00233f
C81 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.Q3 9.83e-19
C82 VDD CLK_div_10_mag_1.Q3 1.18f
C83 CLK_div_10_mag_1.JK_FF_mag_0.J CLK_div_10_mag_0.Q0 4.2e-19
C84 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0209f
C85 CLK_div_10_mag_1.JK_FF_mag_1.QB a_9892_5223# 0.00964f
C86 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 6.88e-21
C87 a_7392_1353# CLK_div_10_mag_0.JK_FF_mag_2.J 3.12e-19
C88 a_1922_1353# CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 4.52e-20
C89 RST CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.00434f
C90 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT a_4582_5223# 9.1e-19
C91 a_5140_4126# a_5300_4126# 0.0504f
C92 CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.25f
C93 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_10_mag_1.JK_FF_mag_2.QB 0.103f
C94 CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 2.81e-20
C95 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 a_995_4126# 0.069f
C96 a_10403_212# CLK_div_10_mag_0.JK_FF_mag_2.J 0.00695f
C97 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_2.QB 1.96f
C98 CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 5.98e-20
C99 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.00233f
C100 CLK_div_10_mag_1.JK_FF_mag_0.J RST 0.0484f
C101 CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.103f
C102 CLK CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 6.64e-19
C103 a_1358_1353# CLK 6.43e-21
C104 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.103f
C105 CLK_div_10_mag_0.JK_FF_mag_0.J CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 1.41e-20
C106 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 8.16e-20
C107 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_4369_212# 0.0203f
C108 CLK_div_10_mag_1.CLK CLK_div_10_mag_0.JK_FF_mag_2.J 4.19e-19
C109 CLK_div_10_mag_0.Q2 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 1.49e-21
C110 RST a_8674_256# 9.66e-19
C111 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.298f
C112 a_230_2335# Vdiv100 0.198f
C113 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT 0.122f
C114 CLK_div_10_mag_1.JK_FF_mag_1.QB a_9328_5223# 0.0811f
C115 a_6828_1309# CLK_div_10_mag_0.JK_FF_mag_2.J 9.32e-19
C116 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00311f
C117 a_4394_3029# CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT 3.38e-20
C118 CLK_div_10_mag_0.JK_FF_mag_1.QB a_2640_256# 0.0811f
C119 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 2.86e-19
C120 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT a_4422_5223# 2.88e-20
C121 VDD CLK_div_10_mag_1.nor_3_mag_0.IN3 0.399f
C122 CLK_div_10_mag_1.CLK CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 6.64e-19
C123 a_4375_1353# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.00378f
C124 CLK_div_10_mag_0.JK_FF_mag_0.J CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00264f
C125 RST CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 3.84e-20
C126 a_841_5223# CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.069f
C127 RST CLK_div_10_mag_1.JK_FF_mag_3.QB 0.179f
C128 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_10_mag_1.JK_FF_mag_2.QB 2.81e-20
C129 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT RST 3.84e-20
C130 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_10_mag_1.CLK 0.235f
C131 CLK_div_10_mag_0.nor_3_mag_0.IN3 a_11738_2752# 2.44e-20
C132 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.235f
C133 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.0228f
C134 VDD CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.792f
C135 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_10_mag_0.and2_mag_0.OUT 8.94e-19
C136 VDD a_1922_1353# 3.14e-19
C137 CLK_div_10_mag_1.JK_FF_mag_0.J CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 1.41e-20
C138 CLK_div_10_mag_0.Q0 a_794_1309# 2.79e-20
C139 a_6668_1309# CLK_div_10_mag_0.JK_FF_mag_2.J 0.00111f
C140 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0343f
C141 CLK_div_10_mag_1.JK_FF_mag_0.J CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.0823f
C142 VDD CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.741f
C143 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.00356f
C144 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_10_mag_1.and2_mag_0.OUT 8.94e-19
C145 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_2.J 0.00488f
C146 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.121f
C147 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 0.0905f
C148 a_3811_1309# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.0732f
C149 a_634_1309# a_794_1309# 0.0504f
C150 a_4939_1353# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0059f
C151 CLK_div_10_mag_0.JK_FF_mag_2.QB a_5093_256# 0.00964f
C152 VDD CLK 1.1f
C153 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 4.36e-20
C154 RST a_794_1309# 9.5e-19
C155 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_11537_1353# 0.00118f
C156 CLK_div_10_mag_0.Q1 a_6662_212# 0.00119f
C157 VDD a_7546_212# 0.00101f
C158 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00718f
C159 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0228f
C160 CLK_div_10_mag_0.nor_3_mag_0.IN3 a_11578_2752# 9.02e-19
C161 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 RST 0.177f
C162 CLK_div_10_mag_0.Q0 CLK_div_10_mag_1.and2_mag_0.OUT 0.0635f
C163 CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_10_mag_1.Q0 1.96f
C164 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.J 0.283f
C165 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0129f
C166 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_1.JK_FF_mag_3.QB 0.28f
C167 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.Q3 0.124f
C168 a_5503_1353# CLK_div_10_mag_0.JK_FF_mag_2.J 7.4e-19
C169 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_6662_212# 1.17e-20
C170 a_4394_3029# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 7.43e-22
C171 a_7599_5223# CLK_div_10_mag_1.JK_FF_mag_2.QB 0.00695f
C172 CLK_div_10_mag_0.Q0 a_788_212# 0.00789f
C173 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.and2_mag_0.OUT 6.22e-20
C174 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_1.JK_FF_mag_3.QB 7.08e-20
C175 RST CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.118f
C176 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.338f
C177 CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_10046_4126# 0.069f
C178 CLK_div_10_mag_1.and2_mag_1.OUT CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 1.29e-19
C179 RST CLK_div_10_mag_1.and2_mag_0.OUT 0.0507f
C180 a_3651_1309# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.0203f
C181 VDD CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 1.03f
C182 a_4375_1353# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0697f
C183 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_2640_256# 0.00372f
C184 VDD a_9510_2450# 3.14e-19
C185 a_11691_256# CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.00372f
C186 RST CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.177f
C187 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_10973_1353# 0.011f
C188 a_10616_5223# RST 8.64e-19
C189 RST CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.0543f
C190 CLK_div_10_mag_1.JK_FF_mag_2.J Vdiv100 4.19e-19
C191 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_6822_212# 1.46e-19
C192 CLK_div_10_mag_0.JK_FF_mag_3.QB a_7956_1353# 2.96e-19
C193 RST CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.019f
C194 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_10_mag_0.and2_mag_0.OUT 6.69e-19
C195 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT RST 0.0763f
C196 a_9839_212# CLK_div_10_mag_0.Q3 0.00789f
C197 a_390_2335# RST 0.00198f
C198 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_5093_256# 0.00378f
C199 a_4939_1353# CLK_div_10_mag_0.JK_FF_mag_2.J 7.4e-19
C200 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.CLK 0.149f
C201 a_7439_5223# CLK_div_10_mag_1.JK_FF_mag_2.QB 0.00696f
C202 VDD CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.652f
C203 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.0654f
C204 CLK_div_10_mag_1.JK_FF_mag_0.J CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.00102f
C205 CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_9482_4126# 0.00372f
C206 CLK_div_10_mag_1.Q1 CLK_div_10_mag_1.JK_FF_mag_2.QB 1.96f
C207 VDD CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.395f
C208 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.122f
C209 CLK_div_10_mag_1.and2_mag_1.OUT RST 0.0284f
C210 a_628_212# a_788_212# 0.0504f
C211 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 0.231f
C212 a_11127_256# CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.069f
C213 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.and2_mag_1.OUT 2.11e-20
C214 VDD a_11738_2752# 0.0407f
C215 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.JK_FF_mag_0.J 0.0156f
C216 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_628_212# 0.0202f
C217 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_10409_1353# 1.43e-19
C218 CLK_div_10_mag_0.JK_FF_mag_0.J CLK_div_10_mag_0.Q2 0.289f
C219 a_230_2335# CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00261f
C220 a_10456_5223# RST 0.00186f
C221 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C222 a_230_2335# CLK_div_10_mag_1.and2_mag_0.OUT 0.00894f
C223 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.J 0.783f
C224 VDD Vdiv100 0.0814f
C225 CLK_div_10_mag_0.JK_FF_mag_3.QB a_7392_1353# 3.25e-19
C226 RST a_8323_5223# 0.00186f
C227 CLK_div_10_mag_0.JK_FF_mag_3.QB a_7386_212# 0.00695f
C228 a_4012_4126# CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 0.069f
C229 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.109f
C230 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.Q1 1.17e-19
C231 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.JK_FF_mag_2.QB 0.348f
C232 CLK_div_10_mag_0.and2_mag_1.OUT RST 4.25e-20
C233 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_1.and2_mag_0.OUT 6.22e-20
C234 VDD CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.994f
C235 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_1.and2_mag_0.OUT 0.065f
C236 a_4375_1353# CLK_div_10_mag_0.JK_FF_mag_2.J 3.12e-19
C237 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00183f
C238 CLK_div_10_mag_1.JK_FF_mag_2.J a_8317_4126# 0.00876f
C239 CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 8.02e-20
C240 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 0.321f
C241 VDD CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.399f
C242 a_6875_5223# CLK_div_10_mag_1.JK_FF_mag_2.QB 0.00964f
C243 RST CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 3.84e-20
C244 RST CLK_div_10_mag_0.JK_FF_mag_2.J 3.04f
C245 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.JK_FF_mag_1.QB 2.59e-21
C246 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.25f
C247 a_230_2335# a_390_2335# 0.186f
C248 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_7956_1353# 4.52e-20
C249 VDD a_11578_2752# 0.234f
C250 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.JK_FF_mag_3.QB 0.0835f
C251 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_9845_1309# 0.00119f
C252 CLK_div_10_mag_1.JK_FF_mag_0.J VDD 0.487f
C253 a_9892_5223# RST 9.41e-19
C254 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT 0.1f
C255 CLK_div_10_mag_0.Q0 CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN 0.00116f
C256 CLK_div_10_mag_0.JK_FF_mag_3.QB a_6828_1309# 0.00392f
C257 RST CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.261f
C258 a_3448_4126# CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 0.00372f
C259 RST a_8163_5223# 0.00186f
C260 CLK_div_10_mag_0.Q1 a_7392_1353# 1.25e-20
C261 CLK_div_10_mag_0.Q0 a_3645_212# 0.001f
C262 CLK_div_10_mag_0.Q1 a_7386_212# 3.6e-22
C263 VDD a_8674_256# 0.00152f
C264 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_1.and2_mag_1.OUT 0.00718f
C265 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT RST 0.0495f
C266 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 4.25e-20
C267 CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_1.nor_3_mag_0.IN3 4.85e-20
C268 CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN RST 9.43e-19
C269 CLK_div_10_mag_1.JK_FF_mag_2.J a_8157_4126# 9.32e-19
C270 a_3811_1309# CLK_div_10_mag_0.JK_FF_mag_2.J 9.32e-19
C271 a_2486_1353# CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00118f
C272 a_3426_3029# CLK_div_10_mag_1.JK_FF_mag_3.QB 1.45e-20
C273 VDD a_8317_4126# 3.78e-19
C274 a_6311_5223# CLK_div_10_mag_1.JK_FF_mag_2.QB 0.0811f
C275 a_8674_256# CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.00372f
C276 CLK_div_10_mag_0.Q0 a_10409_1353# 6.43e-21
C277 a_1405_5223# a_1565_5223# 0.0504f
C278 CLK_div_10_mag_0.Q3 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.338f
C279 a_2486_1353# CLK_div_10_mag_1.and2_mag_0.OUT 2.05e-19
C280 RST a_3645_212# 0.00186f
C281 a_1358_1353# CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.43e-19
C282 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_7392_1353# 0.0202f
C283 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.16f
C284 CLK_div_10_mag_0.Q0 a_1512_212# 0.0101f
C285 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_7386_212# 0.0203f
C286 VDD a_8542_2450# 3.14e-19
C287 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN 1.36e-19
C288 VDD CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.649f
C289 a_9328_5223# RST 9.66e-19
C290 a_11340_5223# VDD 0.0132f
C291 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0854f
C292 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_2129_5223# 1.5e-20
C293 VDD CLK_div_10_mag_1.JK_FF_mag_3.QB 0.911f
C294 CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 4.84e-19
C295 a_277_5223# CLK_div_10_mag_1.Q3 0.0157f
C296 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0384f
C297 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_2.J 0.00488f
C298 VDD CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT 0.649f
C299 a_8542_2450# CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 1.29e-22
C300 a_1922_1353# CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 8.17e-21
C301 RST a_10409_1353# 2.78e-19
C302 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 0.0854f
C303 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 a_8520_1353# 0.00372f
C304 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_788_212# 1.5e-20
C305 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_10_mag_1.Q0 0.00116f
C306 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 0.0432f
C307 RST a_7599_5223# 0.00169f
C308 CLK_div_10_mag_1.CLK CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 3.1e-22
C309 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.121f
C310 RST a_1512_212# 0.00186f
C311 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.0591f
C312 CLK_div_10_mag_0.Q1 a_6828_1309# 0.00939f
C313 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.and2_mag_0.OUT 0.179f
C314 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_10_mag_1.and2_mag_0.OUT 6.69e-19
C315 CLK_div_10_mag_0.nor_3_mag_0.IN3 a_11537_1353# 2.1e-20
C316 CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_1.and2_mag_0.OUT 0.125f
C317 a_2458_3029# RST 4.48e-19
C318 a_3651_1309# CLK_div_10_mag_0.JK_FF_mag_2.J 0.00876f
C319 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00157f
C320 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 0.159f
C321 a_6662_212# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.0202f
C322 VDD a_8157_4126# 2.66e-19
C323 CLK_div_10_mag_0.Q0 a_9845_1309# 0.00939f
C324 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.and2_mag_0.OUT 0.00656f
C325 a_2123_4126# a_2283_4126# 0.0504f
C326 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.27f
C327 CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_10_mag_1.Q3 0.00357f
C328 VDD a_7574_2450# 6e-19
C329 CLK_div_10_mag_0.Q0 CLK_div_10_mag_1.Q1 0.0314f
C330 CLK_div_10_mag_1.and2_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0018f
C331 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_1565_5223# 0.0203f
C332 VDD a_794_1309# 2.66e-19
C333 a_11180_5223# VDD 0.00892f
C334 CLK_div_10_mag_0.JK_FF_mag_0.J CLK_div_10_mag_0.and2_mag_0.OUT 0.0659f
C335 CLK_div_10_mag_0.Q2 a_6822_212# 0.00789f
C336 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 7.08e-20
C337 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 1.54e-19
C338 RST a_7439_5223# 0.00186f
C339 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_1352_212# 9.1e-19
C340 VDD CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 0.652f
C341 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.0894f
C342 a_10610_4126# CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.0202f
C343 a_9482_4126# CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 4.52e-20
C344 a_2129_5223# CLK_div_10_mag_1.Q3 0.00789f
C345 CLK_div_10_mag_0.Q1 a_6668_1309# 0.0101f
C346 CLK_div_10_mag_0.Q2 a_9839_212# 1.86e-20
C347 CLK_div_10_mag_1.JK_FF_mag_2.J a_390_2335# 9.21e-20
C348 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT 0.0286f
C349 RST CLK_div_10_mag_1.Q1 0.133f
C350 VDD CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.457f
C351 a_3426_3029# CLK_div_10_mag_1.and2_mag_0.OUT 0.00138f
C352 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_10_mag_1.and2_mag_1.OUT 4.42e-19
C353 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_3.QB 1e-19
C354 CLK_div_10_mag_0.Q0 CLK_div_10_mag_1.Q0 5.98e-20
C355 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C356 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 5.37e-19
C357 CLK_div_10_mag_0.JK_FF_mag_3.QB a_8110_256# 0.00964f
C358 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0622f
C359 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.122f
C360 CLK_div_10_mag_1.Q3 a_431_4126# 0.069f
C361 VDD CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.22f
C362 CLK_div_10_mag_0.Q0 a_9685_1309# 0.0101f
C363 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.J 4.24e-20
C364 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 0.359f
C365 VDD CLK_div_10_mag_1.and2_mag_0.OUT 0.977f
C366 VDD CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.653f
C367 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.00975f
C368 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.231f
C369 a_10616_5223# VDD 0.00123f
C370 CLK_div_10_mag_1.Q0 RST 0.169f
C371 VDD a_788_212# 0.00892f
C372 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_1405_5223# 0.0733f
C373 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 0.231f
C374 VDD CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.768f
C375 CLK_div_10_mag_1.JK_FF_mag_2.J a_8323_5223# 2.81e-19
C376 CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_10_mag_1.nor_3_mag_0.IN3 0.11f
C377 CLK_div_10_mag_0.Q3 a_11738_2752# 0.019f
C378 RST a_6875_5223# 9.41e-19
C379 VDD CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.395f
C380 a_10046_4126# CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 4.52e-20
C381 a_1565_5223# CLK_div_10_mag_1.Q3 0.0102f
C382 CLK_div_10_mag_0.Q1 a_5503_1353# 0.069f
C383 CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C384 VDD a_390_2335# 0.234f
C385 VDD CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT 0.748f
C386 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.198f
C387 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.321f
C388 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00183f
C389 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 0.00602f
C390 CLK_div_10_mag_0.Q0 a_8520_1353# 9.45e-19
C391 RST CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.00739f
C392 CLK_div_10_mag_0.Q0 a_4369_212# 3.6e-22
C393 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.303f
C394 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.Q3 0.0345f
C395 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_3.QB 0.0615f
C396 VDD CLK_div_10_mag_1.and2_mag_1.OUT 0.58f
C397 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_1.Q1 0.447f
C398 a_431_4126# CLK_div_10_mag_1.nor_3_mag_0.IN3 2.1e-20
C399 a_10456_5223# VDD 0.00101f
C400 CLK_div_10_mag_1.Q0 a_11174_4126# 2.79e-20
C401 VDD a_11537_1353# 3.56e-19
C402 RST a_4369_212# 0.00169f
C403 CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN 2.86e-19
C404 CLK_div_10_mag_0.Q0 a_2640_256# 0.0157f
C405 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 4.24e-20
C406 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_8110_256# 0.00378f
C407 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 5.08e-20
C408 CLK_div_10_mag_0.JK_FF_mag_3.QB RST 0.179f
C409 VDD a_8323_5223# 0.0123f
C410 RST a_6311_5223# 9.66e-19
C411 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_11738_2752# 5.39e-20
C412 CLK_div_10_mag_0.Q1 a_4939_1353# 6.06e-21
C413 CLK_div_10_mag_0.and2_mag_1.OUT VDD 0.58f
C414 a_1405_5223# CLK_div_10_mag_1.Q3 0.0101f
C415 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 0.857f
C416 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_1512_212# 0.0733f
C417 a_6828_1309# CLK_div_10_mag_0.JK_FF_mag_2.QB 1.41e-20
C418 CLK_div_10_mag_1.CLK CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.267f
C419 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C420 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_1559_4126# 0.0202f
C421 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 9.98e-19
C422 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.529f
C423 CLK_div_10_mag_1.JK_FF_mag_0.J CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 0.0275f
C424 RST a_2640_256# 9.66e-19
C425 VDD CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 0.741f
C426 VDD CLK_div_10_mag_0.JK_FF_mag_2.J 1.65f
C427 a_7593_4126# CLK_div_10_mag_1.JK_FF_mag_2.QB 3.25e-19
C428 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 0.0622f
C429 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 4.25e-20
C430 CLK_div_10_mag_0.JK_FF_mag_2.J CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.00586f
C431 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.00125f
C432 a_1922_1353# CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.069f
C433 CLK_div_10_mag_1.Q3 a_2123_4126# 2.79e-20
C434 a_7386_212# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 9.1e-19
C435 a_9892_5223# VDD 0.00152f
C436 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.Q1 1.16f
C437 VDD a_10973_1353# 3.14e-19
C438 CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN a_3426_3029# 0.069f
C439 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_2076_256# 0.0036f
C440 VDD a_8163_5223# 0.00863f
C441 VDD CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 1f
C442 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C443 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 4.27e-20
C444 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_11578_2752# 9.16e-20
C445 CLK_div_10_mag_0.Q2 a_7546_212# 0.0101f
C446 CLK CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 1.48e-20
C447 VDD CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.768f
C448 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.00395f
C449 CLK_div_10_mag_0.Q1 RST 0.133f
C450 a_1352_212# a_1512_212# 0.0504f
C451 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00157f
C452 VDD CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN 0.431f
C453 a_6668_1309# CLK_div_10_mag_0.JK_FF_mag_2.QB 1.86e-20
C454 a_7574_2450# CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 7.43e-22
C455 RST CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 2.96e-19
C456 CLK_div_10_mag_1.JK_FF_mag_3.QB a_4582_5223# 0.00695f
C457 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_1.Q3 0.0345f
C458 a_7029_4126# CLK_div_10_mag_1.JK_FF_mag_2.QB 2.96e-19
C459 VDD a_3645_212# 0.0123f
C460 CLK_div_10_mag_1.Q0 a_2486_1353# 8.17e-21
C461 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT RST 0.266f
C462 CLK_div_10_mag_0.Q0 a_4394_3029# 2.48e-19
C463 a_9328_5223# VDD 0.00152f
C464 CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_1.Q1 0.0995f
C465 CLK_div_10_mag_1.Q0 a_10046_4126# 6.06e-21
C466 CLK_div_10_mag_0.Q2 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 2.64e-19
C467 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 1.49e-21
C468 VDD a_10409_1353# 3.14e-19
C469 CLK_div_10_mag_0.Q2 a_9510_2450# 0.0096f
C470 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.233f
C471 VDD a_7599_5223# 0.00123f
C472 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.235f
C473 VDD a_1512_212# 0.00101f
C474 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.Q1 0.0871f
C475 RST CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 0.0172f
C476 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 0.122f
C477 CLK_div_10_mag_0.Q1 a_3811_1309# 2.79e-20
C478 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 RST 0.00143f
C479 CLK_div_10_mag_1.JK_FF_mag_3.QB a_3858_5223# 0.00964f
C480 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.00163f
C481 CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN Vdiv100 1.82e-19
C482 a_5503_1353# CLK_div_10_mag_0.JK_FF_mag_2.QB 0.0114f
C483 VDD a_2458_3029# 3.14e-19
C484 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN 4.36e-20
C485 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 5.11e-19
C486 CLK_div_10_mag_1.JK_FF_mag_3.QB a_4422_5223# 0.00696f
C487 a_6465_4126# CLK_div_10_mag_1.JK_FF_mag_2.QB 0.0114f
C488 CLK_div_10_mag_0.JK_FF_mag_0.J a_9510_2450# 0.0027f
C489 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00545f
C490 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00137f
C491 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.108f
C492 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.Q0 0.783f
C493 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_10_mag_0.nor_3_mag_0.IN3 7.14e-19
C494 CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.28f
C495 a_3426_3029# CLK_div_10_mag_1.Q1 0.0084f
C496 CLK_div_10_mag_1.Q0 a_9482_4126# 0.069f
C497 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 0.121f
C498 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_10_mag_0.JK_FF_mag_2.J 0.0286f
C499 VDD a_7439_5223# 0.00101f
C500 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 1.54e-21
C501 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C502 CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00163f
C503 CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.0384f
C504 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 a_5657_256# 0.00372f
C505 RST a_2289_5223# 0.00186f
C506 RST a_5093_256# 9.41e-19
C507 VDD CLK_div_10_mag_1.Q1 4.08f
C508 CLK_div_10_mag_1.JK_FF_mag_3.QB a_3294_5223# 0.0811f
C509 a_4939_1353# CLK_div_10_mag_0.JK_FF_mag_2.QB 2.96e-19
C510 CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_1.and2_mag_0.OUT 0.0496f
C511 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.321f
C512 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 1.29e-19
C513 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 7.24e-19
C514 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.0592f
C515 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 2.45e-22
C516 a_3645_212# a_3805_212# 0.0504f
C517 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.J 0.346f
C518 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 0.321f
C519 a_634_1309# CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0203f
C520 CLK_div_10_mag_0.Q2 CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.00114f
C521 a_8323_5223# CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 1.17e-20
C522 a_5140_4126# CLK_div_10_mag_1.JK_FF_mag_3.QB 0.00392f
C523 VDD CLK_div_10_mag_1.Q0 5.05f
C524 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 a_4422_5223# 8.64e-19
C525 RST CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0134f
C526 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.321f
C527 VDD a_9685_1309# 2.21e-19
C528 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.QB 0.348f
C529 CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN a_390_2335# 2.85e-20
C530 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_4529_212# 8.64e-19
C531 CLK_div_10_mag_0.JK_FF_mag_0.J CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00174f
C532 CLK_div_10_mag_1.CLK CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.42f
C533 VDD a_6875_5223# 0.00152f
C534 RST CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT 0.266f
C535 a_7593_4126# RST 1.23e-20
C536 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_3645_212# 0.0202f
C537 CLK_div_10_mag_0.Q3 a_11537_1353# 0.069f
C538 CLK_div_10_mag_1.Q3 CLK_div_10_mag_1.nor_3_mag_0.IN3 0.00442f
C539 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_10_mag_1.CLK 9.71e-20
C540 CLK_div_10_mag_1.JK_FF_mag_0.J CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 2.61e-19
C541 CLK_div_10_mag_0.JK_FF_mag_0.J CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 2.61e-19
C542 a_4375_1353# CLK_div_10_mag_0.JK_FF_mag_2.QB 3.25e-19
C543 CLK_div_10_mag_1.and2_mag_1.OUT CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 0.124f
C544 a_9839_212# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0731f
C545 RST CLK_div_10_mag_0.JK_FF_mag_2.QB 0.179f
C546 a_10403_212# a_10563_212# 0.0504f
C547 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_0.Q3 0.00132f
C548 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 0.00157f
C549 VDD CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.398f
C550 CLK_div_10_mag_0.Q2 a_8674_256# 0.0157f
C551 a_4576_4126# CLK_div_10_mag_1.JK_FF_mag_3.QB 3.25e-19
C552 a_8163_5223# CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 1.5e-20
C553 CLK_div_10_mag_0.Q3 CLK_div_10_mag_0.JK_FF_mag_2.J 2f
C554 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_11334_4126# 0.0203f
C555 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.J 0.0501f
C556 CLK_div_10_mag_1.Q1 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 0.0635f
C557 VDD a_4369_212# 0.00123f
C558 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_10_mag_1.JK_FF_mag_3.QB 0.103f
C559 VDD a_8520_1353# 3.56e-19
C560 a_4939_1353# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 4.52e-20
C561 CLK_div_10_mag_0.Q2 a_8542_2450# 0.0112f
C562 VDD CLK_div_10_mag_0.JK_FF_mag_3.QB 0.911f
C563 CLK_div_10_mag_0.and2_mag_0.OUT a_9510_2450# 0.00138f
C564 VDD a_6311_5223# 0.00152f
C565 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_10409_1353# 0.00378f
C566 CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_10_mag_1.CLK 0.307f
C567 a_8520_1353# CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 4.52e-20
C568 CLK_div_10_mag_0.Q2 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT 0.00146f
C569 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.198f
C570 CLK_div_10_mag_1.JK_FF_mag_0.J a_2283_4126# 8.64e-19
C571 CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 0.0591f
C572 CLK_div_10_mag_1.Q3 CLK 0.00639f
C573 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 4.42e-19
C574 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00356f
C575 a_3811_1309# CLK_div_10_mag_0.JK_FF_mag_2.QB 0.00392f
C576 VDD a_2640_256# 0.00152f
C577 VDD CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.398f
C578 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 6.82e-19
C579 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0854f
C580 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.QB 1.96f
C581 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.11f
C582 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_2.J 0.038f
C583 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT 0.159f
C584 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.00481f
C585 a_7599_5223# CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 0.0203f
C586 a_4012_4126# CLK_div_10_mag_1.JK_FF_mag_3.QB 2.96e-19
C587 a_6875_5223# CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 0.069f
C588 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_11174_4126# 0.0732f
C589 RST CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.0758f
C590 CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 5.13e-19
C591 RST CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.257f
C592 CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_10_mag_1.JK_FF_mag_2.QB 2.59e-21
C593 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.0591f
C594 a_4394_3029# CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.069f
C595 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 a_7956_1353# 0.069f
C596 CLK_div_10_mag_1.Q1 a_5306_5223# 0.00119f
C597 CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN 2.86e-19
C598 CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_10_mag_1.and2_mag_0.OUT 0.0654f
C599 a_4375_1353# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0202f
C600 CLK_div_10_mag_0.Q2 a_7574_2450# 0.00929f
C601 CLK_div_10_mag_0.and2_mag_0.OUT a_11738_2752# 0.00894f
C602 RST CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.266f
C603 RST CLK_div_10_mag_0.JK_FF_mag_1.QB 0.16f
C604 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 a_4576_4126# 0.0697f
C605 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 0.00586f
C606 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_10973_1353# 0.0059f
C607 a_11127_256# CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0036f
C608 RST a_995_4126# 0.0011f
C609 a_841_5223# CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.0036f
C610 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_9845_1309# 0.0732f
C611 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.198f
C612 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT 0.00157f
C613 CLK_div_10_mag_1.JK_FF_mag_3.QB a_2283_4126# 1.86e-20
C614 VDD CLK_div_10_mag_0.Q1 4.08f
C615 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_10973_1353# 5.94e-20
C616 a_5300_4126# CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 0.0203f
C617 CLK_div_10_mag_0.Q0 a_9679_212# 0.00117f
C618 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_2289_5223# 0.0202f
C619 VDD CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.391f
C620 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.and2_mag_0.OUT 3.38e-19
C621 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.322f
C622 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 0.109f
C623 RST a_6662_212# 0.00186f
C624 CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_390_2335# 9.16e-20
C625 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00213f
C626 CLK_div_10_mag_1.nor_3_mag_0.IN3 CLK 2.42e-19
C627 CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_10_mag_0.and2_mag_0.OUT 0.00252f
C628 a_3448_4126# CLK_div_10_mag_1.JK_FF_mag_3.QB 0.0114f
C629 a_7439_5223# CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 0.0733f
C630 VDD CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.999f
C631 a_6311_5223# CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 0.00372f
C632 a_3426_3029# CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 1.29e-22
C633 a_431_4126# CLK_div_10_mag_1.and2_mag_0.OUT 1.54e-19
C634 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_10610_4126# 0.00378f
C635 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.122f
C636 a_9679_212# RST 0.00186f
C637 CLK_div_10_mag_1.Q1 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 0.0343f
C638 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.36f
C639 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0622f
C640 a_3811_1309# CLK_div_10_mag_0.JK_FF_mag_1.QB 1.41e-20
C641 CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN a_2458_3029# 0.069f
C642 a_1358_1353# CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.00378f
C643 CLK_div_10_mag_1.Q1 a_5146_5223# 0.00166f
C644 CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_10_mag_1.and2_mag_1.OUT 0.11f
C645 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 a_4012_4126# 0.0059f
C646 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_1.JK_FF_mag_0.J 9.55e-19
C647 CLK_div_10_mag_0.and2_mag_0.OUT a_11578_2752# 0.0294f
C648 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_10409_1353# 0.0697f
C649 CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00252f
C650 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 2.86e-19
C651 VDD CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 0.395f
C652 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_9685_1309# 0.0203f
C653 VDD CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.391f
C654 CLK_div_10_mag_0.Q3 a_9845_1309# 2.79e-20
C655 VDD a_4394_3029# 6e-19
C656 CLK_div_10_mag_1.JK_FF_mag_3.QB a_2123_4126# 1.41e-20
C657 a_5140_4126# CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 0.0732f
C658 a_9839_212# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 1.5e-20
C659 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 0.00481f
C660 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.231f
C661 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.00975f
C662 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_4369_212# 9.1e-19
C663 CLK_div_10_mag_1.Q3 Vdiv100 0.242f
C664 a_6875_5223# CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 0.00378f
C665 a_6668_1309# a_6828_1309# 0.0504f
C666 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_995_4126# 0.011f
C667 CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT 5.7e-20
C668 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0635f
C669 a_3651_1309# CLK_div_10_mag_0.JK_FF_mag_1.QB 1.86e-20
C670 CLK_div_10_mag_1.Q1 a_4582_5223# 3.6e-22
C671 CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_1.Q1 1.17e-19
C672 CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_2.QB 0.00123f
C673 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT 0.0334f
C674 CLK_div_10_mag_0.and2_mag_0.OUT a_8542_2450# 0.00138f
C675 CLK_div_10_mag_1.JK_FF_mag_2.J a_7593_4126# 3.12e-19
C676 VDD a_2289_5223# 0.00727f
C677 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_10_mag_1.Q1 0.108f
C678 CLK_div_10_mag_0.Q1 a_3805_212# 0.00789f
C679 RST CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0201f
C680 VDD a_5093_256# 0.00152f
C681 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 2.81e-20
C682 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 a_7439_5223# 8.64e-19
C683 RST CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.0675f
C684 a_4576_4126# CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 0.00378f
C685 CLK_div_10_mag_0.Q0 a_7956_1353# 6.06e-21
C686 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.0979f
C687 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 0.0979f
C688 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_0.Q2 0.0165f
C689 CLK_div_10_mag_1.Q1 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 0.00335f
C690 CLK_div_10_mag_1.JK_FF_mag_2.J a_841_5223# 0.00964f
C691 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 RST 0.189f
C692 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 0.00183f
C693 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 0.0205f
C694 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_2.J 0.0626f
C695 VDD CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.742f
C696 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.338f
C697 a_2486_1353# CLK_div_10_mag_0.JK_FF_mag_1.QB 0.0114f
C698 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.768f
C699 a_1358_1353# CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0697f
C700 Vdiv100 CLK_div_10_mag_1.nor_3_mag_0.IN3 0.0263f
C701 CLK_div_10_mag_0.JK_FF_mag_0.J CLK_div_10_mag_0.and2_mag_1.OUT 2.57e-20
C702 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 0.0129f
C703 CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_10_mag_0.Q0 0.00158f
C704 CLK_div_10_mag_1.JK_FF_mag_2.J a_7029_4126# 7.4e-19
C705 VDD CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT 0.999f
C706 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.122f
C707 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.25f
C708 a_1358_1353# CLK_div_10_mag_0.JK_FF_mag_1.QB 3.33e-19
C709 a_5300_4126# CLK_div_10_mag_1.Q1 0.0101f
C710 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.J 0.0905f
C711 a_10563_212# RST 0.00127f
C712 VDD a_7593_4126# 3.14e-19
C713 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_8520_1353# 0.00118f
C714 CLK_div_10_mag_0.JK_FF_mag_0.J CLK_div_10_mag_0.JK_FF_mag_2.J 0.0156f
C715 VDD CLK_div_10_mag_0.JK_FF_mag_2.QB 0.913f
C716 CLK_div_10_mag_1.JK_FF_mag_1.QB RST 0.144f
C717 a_11174_4126# CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.00119f
C718 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.28f
C719 a_841_5223# VDD 3.14e-19
C720 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.and2_mag_0.OUT 0.125f
C721 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_7546_212# 8.64e-19
C722 CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 1.49e-21
C723 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.121f
C724 VDD CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.742f
C725 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_995_4126# 0.0059f
C726 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_10_mag_0.Q3 0.11f
C727 a_7392_1353# RST 1.23e-20
C728 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_1.and2_mag_0.OUT 3.38e-19
C729 CLK_div_10_mag_0.Q1 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 0.00145f
C730 RST a_7386_212# 0.00169f
C731 Vdiv100 CLK 0.00102f
C732 CLK_div_10_mag_1.JK_FF_mag_2.J a_995_4126# 2.96e-19
C733 CLK_div_10_mag_1.JK_FF_mag_2.J a_6465_4126# 7.4e-19
C734 a_5140_4126# CLK_div_10_mag_1.Q1 0.00939f
C735 CLK_div_10_mag_0.JK_FF_mag_1.QB a_1352_212# 0.00695f
C736 VDD a_7029_4126# 3.14e-19
C737 a_4369_212# a_4529_212# 0.0504f
C738 a_10403_212# RST 0.00169f
C739 a_10610_4126# CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 1.43e-19
C740 CLK_div_10_mag_1.CLK RST 5.44e-19
C741 CLK_div_10_mag_1.JK_FF_mag_1.QB a_11174_4126# 0.00392f
C742 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_10610_4126# 0.0697f
C743 CLK_div_10_mag_1.CLK a_11334_4126# 0.0101f
C744 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C745 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.447f
C746 CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.00182f
C747 CLK_div_10_mag_0.Q3 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C748 VDD CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.654f
C749 a_2458_3029# CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 8.17e-21
C750 VDD CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.768f
C751 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 4.42e-19
C752 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_1.and2_mag_1.OUT 0.00243f
C753 VDD CLK_div_10_mag_0.JK_FF_mag_1.QB 0.92f
C754 CLK_div_10_mag_1.Q3 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 6.63e-19
C755 VDD CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 1f
C756 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.159f
C757 VDD a_995_4126# 3.14e-19
C758 CLK_div_10_mag_1.and2_mag_1.OUT a_1559_4126# 5.94e-20
C759 a_4576_4126# CLK_div_10_mag_1.Q1 1.25e-20
C760 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.nor_3_mag_0.IN3 4.85e-20
C761 a_2486_1353# CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 4.52e-20
C762 VDD a_6465_4126# 3.56e-19
C763 CLK_div_10_mag_0.and2_mag_0.OUT a_11537_1353# 1.54e-19
C764 CLK_div_10_mag_1.Q3 CLK_div_10_mag_1.and2_mag_0.OUT 0.124f
C765 RST CLK_div_10_mag_1.JK_FF_mag_2.QB 0.179f
C766 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_10_mag_1.Q1 0.235f
C767 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.122f
C768 a_10046_4126# CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.011f
C769 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_0.and2_mag_0.OUT 0.0693f
C770 CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_9510_2450# 8.17e-21
C771 CLK_div_10_mag_0.Q1 a_4529_212# 0.0101f
C772 CLK_div_10_mag_0.Q1 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 1.58e-20
C773 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.0215f
C774 VDD a_6662_212# 0.0132f
C775 CLK_div_10_mag_1.JK_FF_mag_1.QB a_10610_4126# 3.33e-19
C776 CLK_div_10_mag_1.CLK a_11174_4126# 0.00939f
C777 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_10046_4126# 0.0059f
C778 a_2129_5223# CLK_div_10_mag_1.Q0 0.00164f
C779 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_10_mag_1.Q1 5.37e-19
C780 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.J 0.00656f
C781 CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 4.42e-19
C782 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT a_5306_5223# 1.17e-20
C783 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN a_10046_4126# 8.17e-21
C784 VDD a_9679_212# 0.00727f
C785 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.103f
C786 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_1.Q1 2.96e-19
C787 CLK_div_10_mag_0.Q2 CLK_div_10_mag_1.Q0 0.0204f
C788 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 RST 9.24e-20
C789 CLK_div_10_mag_0.Q2 a_9685_1309# 6.36e-19
C790 VDD a_11691_256# 3.14e-19
C791 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 0.0215f
C792 CLK_div_10_mag_1.and2_mag_1.OUT CLK_div_10_mag_1.Q3 0.00132f
C793 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 1.48e-19
C794 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 4.84e-19
C795 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.529f
C796 CLK_div_10_mag_0.Q0 a_5503_1353# 9.26e-19
C797 CLK_div_10_mag_1.nor_3_mag_0.IN3 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00182f
C798 a_9482_4126# CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.00118f
C799 CLK_div_10_mag_1.JK_FF_mag_1.QB a_10046_4126# 2.96e-19
C800 CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_10_mag_1.nor_3_mag_0.IN3 0.144f
C801 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 a_3858_5223# 0.069f
C802 CLK_div_10_mag_1.CLK a_10610_4126# 6.43e-21
C803 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 a_431_4126# 0.00372f
C804 CLK_div_10_mag_0.JK_FF_mag_0.J CLK_div_10_mag_1.Q0 4.2e-19
C805 CLK_div_10_mag_1.Q0 a_4012_4126# 6.06e-21
C806 a_11578_2752# a_11738_2752# 0.186f
C807 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.0116f
C808 CLK_div_10_mag_0.JK_FF_mag_0.J a_9685_1309# 8.64e-19
C809 RST CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00237f
C810 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT a_5146_5223# 1.5e-20
C811 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_1.JK_FF_mag_2.QB 3.49e-19
C812 a_6465_4126# CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 4.52e-20
C813 a_794_1309# CLK 0.00939f
C814 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 0.0854f
C815 a_7593_4126# CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 0.0202f
C816 CLK_div_10_mag_1.CLK CLK_div_10_mag_0.nor_3_mag_0.IN3 0.0267f
C817 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_3805_212# 1.5e-20
C818 a_1922_1353# CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.011f
C819 CLK_div_10_mag_0.Q2 a_8520_1353# 0.069f
C820 VDD a_11127_256# 3.14e-19
C821 a_390_2335# CLK_div_10_mag_1.nor_3_mag_0.IN3 9.02e-19
C822 RST a_8110_256# 9.41e-19
C823 VDD CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.395f
C824 CLK_div_10_mag_1.Q0 a_2283_4126# 0.0101f
C825 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_3.QB 1.96f
C826 VDD CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 1.22f
C827 a_8157_4126# CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 0.00119f
C828 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.JK_FF_mag_1.QB 9.14e-19
C829 CLK CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.407f
C830 CLK_div_10_mag_0.JK_FF_mag_1.QB a_2076_256# 0.00964f
C831 CLK_div_10_mag_1.JK_FF_mag_1.QB a_9482_4126# 0.0114f
C832 VDD CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.654f
C833 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 a_3294_5223# 0.00372f
C834 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.121f
C835 CLK_div_10_mag_1.and2_mag_0.OUT CLK 6.39e-19
C836 CLK_div_10_mag_1.Q0 a_3448_4126# 9.45e-19
C837 RST CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.0152f
C838 a_277_5223# CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.00372f
C839 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.QB 3.49e-19
C840 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT a_4582_5223# 0.0203f
C841 CLK a_788_212# 0.00164f
C842 VDD a_7956_1353# 3.14e-19
C843 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD 0.442f
C844 a_7029_4126# CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 4.52e-20
C845 CLK_div_10_mag_0.JK_FF_mag_0.J CLK_div_10_mag_0.JK_FF_mag_3.QB 5.7e-19
C846 CLK CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.235f
C847 CLK_div_10_mag_1.Q0 a_2123_4126# 0.00939f
C848 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 2.48e-20
C849 a_5503_1353# CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.00372f
C850 CLK_div_10_mag_0.JK_FF_mag_0.J CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 8.2e-19
C851 CLK_div_10_mag_0.Q0 a_4375_1353# 6.43e-21
C852 a_7593_4126# CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 0.0697f
C853 CLK_div_10_mag_1.JK_FF_mag_1.QB VDD 0.92f
C854 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_7574_2450# 2.36e-22
C855 CLK_div_10_mag_0.Q0 RST 0.158f
C856 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.Q2 0.98f
C857 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT a_3858_5223# 0.00378f
C858 CLK_div_10_mag_0.JK_FF_mag_2.QB a_4529_212# 0.00696f
C859 RST a_634_1309# 8.88e-19
C860 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT a_4422_5223# 0.0733f
C861 VDD a_7392_1353# 3.14e-19
C862 CLK_div_10_mag_0.Q1 a_5657_256# 0.0157f
C863 a_4375_1353# RST 1.23e-20
C864 VDD a_7386_212# 0.00123f
C865 CLK_div_10_mag_1.JK_FF_mag_0.J CLK_div_10_mag_1.JK_FF_mag_3.QB 5.7e-19
C866 CLK_div_10_mag_0.JK_FF_mag_2.J CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.11f
C867 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.018f
C868 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 1.36e-19
C869 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0352f
C870 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_1.Q0 9.9e-19
C871 CLK_div_10_mag_0.JK_FF_mag_0.J CLK_div_10_mag_0.Q1 0.0685f
C872 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 a_7029_4126# 0.069f
C873 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 6.89e-19
C874 CLK_div_10_mag_1.Q0 CLK_div_10_mag_0.and2_mag_0.OUT 0.0635f
C875 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.J 0.00602f
C876 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.nor_3_mag_0.IN3 4.39e-19
C877 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.JK_FF_mag_2.QB 0.0838f
C878 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00118f
C879 VDD a_10403_212# 2.21e-19
C880 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 0.00118f
C881 CLK_div_10_mag_1.Q0 a_1559_4126# 6.43e-21
C882 a_4939_1353# CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.069f
C883 CLK_div_10_mag_0.Q0 a_628_212# 0.00335f
C884 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_431_4126# 4.52e-20
C885 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.0894f
C886 CLK_div_10_mag_0.Q0 a_3811_1309# 0.00939f
C887 a_7029_4126# CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 0.0059f
C888 VDD CLK_div_10_mag_1.CLK 1.47f
C889 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT a_8317_4126# 0.0203f
C890 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 8.16e-20
C891 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_2076_256# 0.069f
C892 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C893 Vdiv100 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 8.11e-20
C894 VDD a_6828_1309# 2.66e-19
C895 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.0205f
C896 Vdiv100 CLK_div_10_mag_1.and2_mag_0.OUT 0.119f
C897 a_2129_5223# a_2289_5223# 0.0504f
C898 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 a_6465_4126# 0.00372f
C899 a_11174_4126# a_11334_4126# 0.0504f
C900 CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 6.89e-19
C901 a_8157_4126# a_8317_4126# 0.0504f
C902 CLK_div_10_mag_0.and2_mag_1.OUT a_9510_2450# 3.92e-20
C903 a_9679_212# CLK_div_10_mag_0.Q3 0.00335f
C904 a_230_2335# RST 0.00189f
C905 VDD CLK_div_10_mag_1.JK_FF_mag_2.QB 0.913f
C906 RST CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 9.24e-20
C907 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_4529_212# 0.0733f
C908 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.Q3 0.149f
C909 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.and2_mag_0.OUT 1.33e-20
C910 CLK_div_10_mag_0.Q0 a_3651_1309# 0.0101f
C911 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 4.27e-20
C912 RST CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 0.055f
C913 a_11691_256# CLK_div_10_mag_0.Q3 0.0157f
C914 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 RST 0.0521f
C915 a_390_2335# Vdiv100 0.0132f
C916 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT a_8157_4126# 0.0732f
C917 CLK_div_10_mag_1.JK_FF_mag_0.J CLK_div_10_mag_1.and2_mag_0.OUT 0.0659f
C918 CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 8.16e-20
C919 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_10_mag_0.and2_mag_0.OUT 0.00178f
C920 VDD a_6668_1309# 0.00746f
C921 a_11180_5223# a_11340_5223# 0.0504f
C922 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_5093_256# 0.0036f
C923 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 1.98e-19
C924 VDD CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.397f
C925 a_8163_5223# CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 1.46e-19
C926 a_4576_4126# CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT 0.0202f
C927 a_3448_4126# CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 4.52e-20
C928 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.00183f
C929 CLK_div_10_mag_1.Q3 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.11f
C930 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_2.J 0.0432f
C931 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 8.16e-20
C932 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_3.QB 0.0378f
C933 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT 0.121f
C934 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_8542_2450# 5.1e-20
C935 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_2.J 0.00586f
C936 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT 8.02e-20
C937 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.122f
C938 CLK_div_10_mag_0.Q0 a_2486_1353# 0.069f
C939 CLK_div_10_mag_0.Q2 a_7593_4126# 7.43e-22
C940 a_11738_2752# CLK_div_10_mag_0.JK_FF_mag_2.J 3.02e-19
C941 a_11127_256# CLK_div_10_mag_0.Q3 0.00859f
C942 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.and2_mag_0.OUT 0.0529f
C943 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 0.00975f
C944 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00243f
C945 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0343f
C946 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.346f
C947 CLK_div_10_mag_0.Q3 CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 6.63e-19
C948 CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_10_mag_1.and2_mag_0.OUT 1.33e-20
C949 CLK_div_10_mag_1.JK_FF_mag_0.J CLK_div_10_mag_1.and2_mag_1.OUT 2.57e-20
C950 a_3651_1309# a_3811_1309# 0.0504f
C951 VDD CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.14f
C952 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.122f
C953 a_2486_1353# RST 0.00104f
C954 VDD a_5503_1353# 3.56e-19
C955 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.J 0.251f
C956 CLK_div_10_mag_0.JK_FF_mag_2.QB a_5657_256# 0.0811f
C957 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_10_mag_1.JK_FF_mag_2.QB 0.198f
C958 a_4012_4126# CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT 4.52e-20
C959 RST a_10046_4126# 6.14e-19
C960 RST a_1358_1353# 0.0012f
C961 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.28f
C962 CLK_div_10_mag_0.Q0 CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.0042f
C963 RST CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.374f
C964 CLK_div_10_mag_0.Q1 a_6822_212# 0.00166f
C965 VDD CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.431f
C966 VDD a_8110_256# 0.00152f
C967 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_7956_1353# 0.011f
C968 RST CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.0795f
C969 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_7574_2450# 0.069f
C970 CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_10_mag_0.JK_FF_mag_1.QB 0.00154f
C971 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_10973_1353# 4.52e-20
C972 a_8110_256# CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.069f
C973 CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_995_4126# 5.94e-20
C974 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_10_mag_1.nor_3_mag_0.IN3 7.14e-19
C975 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT 0.00183f
C976 a_11578_2752# CLK_div_10_mag_0.JK_FF_mag_2.J 9.21e-20
C977 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.122f
C978 a_10563_212# CLK_div_10_mag_0.Q3 0.0101f
C979 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 RST 0.225f
C980 CLK_div_10_mag_0.Q0 a_9482_4126# 8.17e-21
C981 a_794_1309# CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00119f
C982 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_6822_212# 1.5e-20
C983 CLK_div_10_mag_0.Q0 a_1352_212# 0.0102f
C984 CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.00975f
C985 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 5.13e-19
C986 VDD CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.648f
C987 CLK_div_10_mag_1.JK_FF_mag_2.J RST 3.06f
C988 VDD a_4939_1353# 3.14e-19
C989 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_628_212# 1.17e-20
C990 RST a_9482_4126# 6.14e-19
C991 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.338f
C992 RST a_1352_212# 8.64e-19
C993 CLK_div_10_mag_1.Q1 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 0.018f
C994 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_7392_1353# 1.43e-19
C995 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 3.38e-19
C996 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C997 a_10563_212# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 8.64e-19
C998 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_10409_1353# 0.0202f
C999 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_2289_5223# 1.17e-20
C1000 CLK_div_10_mag_1.JK_FF_mag_0.J CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN 0.125f
C1001 CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.101f
C1002 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0592f
C1003 CLK_div_10_mag_0.Q0 VDD 5.05f
C1004 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.J 0.1f
C1005 CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 0.343f
C1006 a_10403_212# CLK_div_10_mag_0.Q3 0.0102f
C1007 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_788_212# 1.46e-19
C1008 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00118f
C1009 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 6.82e-19
C1010 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_1.QB 7.08e-20
C1011 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.159f
C1012 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 1.3f
C1013 VDD a_634_1309# 0.00752f
C1014 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.00118f
C1015 CLK_div_10_mag_0.Q2 a_6662_212# 0.00335f
C1016 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_10_mag_1.Q3 0.0635f
C1017 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.343f
C1018 VDD a_4375_1353# 3.14e-19
C1019 CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00154f
C1020 CLK_div_10_mag_1.CLK CLK_div_10_mag_0.Q3 0.256f
C1021 VDD RST 2.73f
C1022 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_1.JK_FF_mag_2.QB 0.25f
C1023 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_788_212# 0.0731f
C1024 VDD a_11334_4126# 0.00752f
C1025 a_6875_5223# CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 0.0036f
C1026 a_390_2335# CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00239f
C1027 CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 0.00137f
C1028 RST CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.0172f
C1029 a_11340_5223# CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 1.17e-20
C1030 CLK_div_10_mag_0.Q2 a_9679_212# 2.55e-20
C1031 CLK_div_10_mag_1.JK_FF_mag_2.J a_230_2335# 3.02e-19
C1032 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.233f
C1033 a_390_2335# CLK_div_10_mag_1.and2_mag_0.OUT 0.0294f
C1034 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_6828_1309# 0.00119f
C1035 CLK_div_10_mag_0.JK_FF_mag_3.QB a_7546_212# 0.00696f
C1036 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 0.0501f
C1037 a_11340_5223# CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.0202f
C1038 CLK_div_10_mag_1.JK_FF_mag_0.J a_2458_3029# 0.0027f
C1039 CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN CLK_div_10_mag_1.JK_FF_mag_3.QB 1e-19
C1040 CLK_div_10_mag_1.and2_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 9.64e-19
C1041 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.283f
C1042 CLK_div_10_mag_1.and2_mag_1.OUT CLK_div_10_mag_1.and2_mag_0.OUT 0.0693f
C1043 CLK_div_10_mag_1.Q3 a_2289_5223# 0.00335f
C1044 VDD a_628_212# 0.0132f
C1045 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_841_5223# 0.00378f
C1046 VDD a_3811_1309# 2.66e-19
C1047 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 0.122f
C1048 a_10456_5223# a_10616_5223# 0.0504f
C1049 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.273f
C1050 CLK_div_10_mag_1.CLK CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 2.16e-19
C1051 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0894f
C1052 VDD a_11174_4126# 2.66e-19
C1053 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_10_mag_0.and2_mag_0.OUT 0.00157f
C1054 a_11180_5223# CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 1.5e-20
C1055 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_10_mag_1.JK_FF_mag_2.QB 0.0591f
C1056 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.J 1.48e-19
C1057 VDD a_230_2335# 0.0407f
C1058 a_1358_1353# CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0202f
C1059 CLK_div_10_mag_1.JK_FF_mag_0.J CLK_div_10_mag_1.Q1 0.0685f
C1060 VDD CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.397f
C1061 CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.J 5.05e-20
C1062 a_11180_5223# CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.0731f
C1063 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.359f
C1064 VDD CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 1.07f
C1065 CLK_div_10_mag_0.Q0 a_3805_212# 0.00166f
C1066 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0622f
C1067 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_2.J 0.0432f
C1068 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_2.QB 0.0378f
C1069 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.108f
C1070 VDD CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 1.14f
C1071 RST CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 0.0172f
C1072 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT a_8323_5223# 0.0202f
C1073 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 8.16e-20
C1074 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.0378f
C1075 VDD a_3651_1309# 3.78e-19
C1076 RST a_3805_212# 0.00186f
C1077 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.00157f
C1078 CLK_div_10_mag_1.JK_FF_mag_0.J CLK_div_10_mag_1.Q0 0.487f
C1079 CLK_div_10_mag_0.Q0 a_2076_256# 0.00859f
C1080 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_7546_212# 0.0733f
C1081 VDD a_10610_4126# 3.14e-19
C1082 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.233f
C1083 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.Q2 0.305f
C1084 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.Q3 0.0263f
C1085 a_10616_5223# CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.0203f
C1086 a_841_5223# CLK_div_10_mag_1.Q3 0.00859f
C1087 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.11f
C1088 a_9892_5223# CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.069f
C1089 a_5300_4126# CLK_div_10_mag_1.JK_FF_mag_2.QB 1.86e-20
C1090 CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN CLK_div_10_mag_1.and2_mag_0.OUT 0.0758f
C1091 CLK_div_10_mag_0.Q1 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 2.96e-19
C1092 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_1352_212# 0.0203f
C1093 VDD CLK_div_10_mag_0.nor_3_mag_0.IN3 0.399f
C1094 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_10_mag_1.Q1 4.66e-21
C1095 CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_10_mag_1.Q1 0.311f
C1096 a_10616_5223# CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 9.1e-19
C1097 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_995_4126# 4.52e-20
C1098 RST a_2076_256# 9.41e-19
C1099 CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.122f
C1100 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_10_mag_1.Q1 7.24e-19
C1101 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.0376f
C1102 CLK_div_10_mag_1.Q0 a_8317_4126# 0.0101f
C1103 RST CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.0763f
C1104 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_8110_256# 0.0036f
C1105 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_0.J 0.0275f
C1106 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT a_8163_5223# 0.0731f
C1107 RST a_5306_5223# 0.00186f
C1108 a_11537_1353# CLK_div_10_mag_0.JK_FF_mag_2.J 0.0114f
C1109 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.27f
C1110 a_6822_212# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.0731f
C1111 VDD a_2486_1353# 3.56e-19
C1112 a_11340_5223# CLK_div_10_mag_1.Q0 0.00335f
C1113 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.JK_FF_mag_3.QB 0.0615f
C1114 a_8157_4126# CLK_div_10_mag_1.Q1 2.79e-20
C1115 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00152f
C1116 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C1117 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C1118 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT 0.298f
C1119 VDD a_10046_4126# 3.14e-19
C1120 VDD CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1f
C1121 VDD a_1358_1353# 3.14e-19
C1122 RST CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00229f
C1123 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.0635f
C1124 CLK_div_10_mag_0.Q2 a_7386_212# 0.0102f
C1125 a_10456_5223# CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.0733f
C1126 a_5140_4126# CLK_div_10_mag_1.JK_FF_mag_2.QB 1.41e-20
C1127 a_9328_5223# CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.00372f
C1128 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00943f
C1129 a_3426_3029# CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN 5.1e-20
C1130 a_2458_3029# CLK_div_10_mag_1.and2_mag_0.OUT 0.00138f
C1131 VDD CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.792f
C1132 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_1512_212# 2.88e-20
C1133 a_10456_5223# CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 2.88e-20
C1134 a_8163_5223# a_8323_5223# 0.0504f
C1135 CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 1.98e-19
C1136 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.768f
C1137 CLK_div_10_mag_0.Q2 a_10403_212# 3.6e-22
C1138 a_6662_212# a_6822_212# 0.0504f
C1139 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.0018f
C1140 CLK_div_10_mag_1.Q0 a_8157_4126# 0.00939f
C1141 VDD CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.457f
C1142 VDD CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.652f
C1143 RST CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 0.266f
C1144 RST a_5146_5223# 0.00186f
C1145 a_10973_1353# CLK_div_10_mag_0.JK_FF_mag_2.J 2.96e-19
C1146 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT a_7599_5223# 9.1e-19
C1147 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_10_mag_1.Q1 0.00152f
C1148 CLK_div_10_mag_0.JK_FF_mag_3.QB a_8674_256# 0.0811f
C1149 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.Q3 0.149f
C1150 CLK_div_10_mag_1.Q0 a_7574_2450# 2.48e-19
C1151 CLK CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.267f
C1152 CLK_div_10_mag_1.JK_FF_mag_2.J VDD 1.65f
C1153 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.857f
C1154 a_11180_5223# CLK_div_10_mag_1.Q0 0.00789f
C1155 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.122f
C1156 VDD a_9482_4126# 3.56e-19
C1157 VDD a_1352_212# 0.00123f
C1158 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.QB 2.81e-20
C1159 CLK_div_10_mag_0.Q2 a_6828_1309# 2.79e-20
C1160 CLK_div_10_mag_0.JK_FF_mag_3.QB a_8542_2450# 1.45e-20
C1161 a_9679_212# a_9839_212# 0.0504f
C1162 CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_10_mag_1.Q1 0.0529f
C1163 a_9892_5223# CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.00378f
C1164 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 0.0126f
C1165 RST CLK_div_10_mag_0.Q3 0.0395f
C1166 CLK_div_10_mag_1.and2_mag_1.OUT a_2458_3029# 3.92e-20
C1167 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_10_mag_1.Q1 1.58e-20
C1168 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 RST 0.055f
C1169 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_1.Q0 0.0042f
C1170 CLK_div_10_mag_0.and2_mag_1.OUT a_10409_1353# 5.94e-20
C1171 CLK_div_10_mag_0.JK_FF_mag_2.J a_3645_212# 2.81e-19
C1172 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 Vdiv100 3.1e-22
C1173 CLK_div_10_mag_0.Q2 CLK_div_10_mag_1.JK_FF_mag_2.QB 1.28e-20
C1174 CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN RST 0.00594f
C1175 VDD a_3426_3029# 3.14e-19
C1176 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.121f
C1177 RST a_4582_5223# 0.00169f
C1178 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT a_7439_5223# 2.88e-20
C1179 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.101f
C1180 a_10409_1353# CLK_div_10_mag_0.JK_FF_mag_2.J 3.25e-19
C1181 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 5.11e-19
C1182 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.and2_mag_0.OUT 0.026f
C1183 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 RST 9.24e-20
C1184 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_10_mag_1.Q1 0.338f
C1185 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_10_mag_0.and2_mag_0.OUT 0.00101f
C1186 a_10616_5223# CLK_div_10_mag_1.Q0 0.0102f
C1187 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 a_5093_256# 0.069f
C1188 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 a_5146_5223# 1.46e-19
C1189 RST CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.152f
C1190 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.0635f
C1191 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.and2_mag_0.OUT 0.0496f
C1192 VDD CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.395f
C1193 RST CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 0.177f
C1194 a_7593_4126# CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 1.43e-19
C1195 RST a_4529_212# 0.00186f
C1196 CLK_div_10_mag_1.and2_mag_1.OUT CLK_div_10_mag_1.Q1 8.51e-22
C1197 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.113f
C1198 CLK_div_10_mag_0.Q1 a_8542_2450# 0.0084f
C1199 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 7.24e-19
C1200 a_1922_1353# CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0059f
C1201 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT 0.233f
C1202 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_10_mag_1.and2_mag_0.OUT 0.00178f
C1203 RST a_3858_5223# 9.41e-19
C1204 CLK_div_10_mag_0.Q1 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT 4.66e-21
C1205 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 0.00586f
C1206 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00183f
C1207 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_2076_256# 0.00378f
C1208 CLK_div_10_mag_1.Q1 a_8323_5223# 0.00335f
C1209 a_1922_1353# CLK_div_10_mag_0.JK_FF_mag_1.QB 2.96e-19
C1210 RST a_4422_5223# 0.00186f
C1211 a_9845_1309# CLK_div_10_mag_0.JK_FF_mag_2.J 0.00486f
C1212 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.and2_mag_1.OUT 2.11e-20
C1213 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 2.11e-19
C1214 CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_10_mag_0.and2_mag_0.OUT 0.0063f
C1215 CLK CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 9.71e-20
C1216 a_2458_3029# CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN 5.1e-20
C1217 a_10456_5223# CLK_div_10_mag_1.Q0 0.0101f
C1218 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_10_mag_1.Q1 0.273f
C1219 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0569f
C1220 a_7546_212# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 2.88e-20
C1221 CLK CLK_div_10_mag_0.JK_FF_mag_1.QB 0.307f
C1222 CLK_div_10_mag_1.Q0 a_8323_5223# 0.001f
C1223 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 0.00213f
C1224 a_7029_4126# CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 0.011f
C1225 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_10_mag_1.JK_FF_mag_3.QB 0.198f
C1226 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.198f
C1227 CLK_div_10_mag_0.Q1 a_7574_2450# 0.0105f
C1228 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 2.11e-19
C1229 a_9679_212# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0202f
C1230 RST a_3294_5223# 9.66e-19
C1231 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.103f
C1232 CLK_div_10_mag_0.Q2 a_8110_256# 0.00859f
C1233 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 0.0285f
C1234 a_5503_1353# CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.00118f
C1235 CLK_div_10_mag_1.Q1 a_8163_5223# 0.00789f
C1236 VDD CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 0.395f
C1237 CLK_div_10_mag_0.JK_FF_mag_0.J CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0836f
C1238 CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_10_mag_0.Q3 0.00442f
C1239 a_9685_1309# CLK_div_10_mag_0.JK_FF_mag_2.J 0.00111f
C1240 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 1.54e-21
C1241 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_7574_2450# 3.38e-20
C1242 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0995f
C1243 CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN CLK_div_10_mag_1.Q1 0.303f
C1244 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 a_3858_5223# 0.0036f
C1245 a_9892_5223# CLK_div_10_mag_1.Q0 0.00859f
C1246 VDD a_3805_212# 0.00863f
C1247 CLK_div_10_mag_1.CLK CLK_div_10_mag_0.and2_mag_0.OUT 0.122f
C1248 CLK_div_10_mag_0.JK_FF_mag_0.J CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.125f
C1249 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.0343f
C1250 a_6465_4126# CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 0.00118f
C1251 CLK_div_10_mag_1.Q0 a_8163_5223# 0.00166f
C1252 CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN RST 0.021f
C1253 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 5.7e-20
C1254 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.00335f
C1255 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.338f
C1256 VDD a_2076_256# 0.00152f
C1257 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN 0.0116f
C1258 a_7439_5223# a_7599_5223# 0.0504f
C1259 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00157f
C1260 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 0.0334f
C1261 VDD CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.748f
C1262 a_4939_1353# CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.011f
C1263 CLK_div_10_mag_1.Q1 a_7599_5223# 0.0102f
C1264 VDD a_5306_5223# 0.0132f
C1265 a_8520_1353# CLK_div_10_mag_0.JK_FF_mag_2.J 7.4e-19
C1266 a_4394_3029# CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 2.36e-22
C1267 CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.11f
C1268 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_11537_1353# 0.00372f
C1269 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.Q2 0.622f
C1270 a_2129_5223# RST 0.00186f
C1271 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_2.J 0.0835f
C1272 a_4576_4126# RST 1.23e-20
C1273 a_9328_5223# CLK_div_10_mag_1.Q0 0.0157f
C1274 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.108f
C1275 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.122f
C1276 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT RST 0.0758f
C1277 RST a_431_4126# 4.42e-19
C1278 VDD CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.648f
C1279 CLK_div_10_mag_0.Q2 RST 0.105f
C1280 CLK_div_10_mag_1.Q0 a_7599_5223# 3.6e-22
C1281 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_2.J 0.0592f
C1282 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_1.JK_FF_mag_3.QB 0.25f
C1283 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 1.3f
C1284 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_2283_4126# 0.0203f
C1285 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.J 0.487f
C1286 a_5140_4126# CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 0.00119f
C1287 CLK_div_10_mag_1.Q0 a_2458_3029# 0.01f
C1288 RST CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 9.24e-20
C1289 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT a_7593_4126# 0.00378f
C1290 RST CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0115f
C1291 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.343f
C1292 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 9.73e-19
C1293 RST a_5657_256# 9.66e-19
C1294 CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_230_2335# 5.39e-20
C1295 VDD CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 1f
C1296 a_4375_1353# CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 1.43e-19
C1297 CLK_div_10_mag_1.Q1 a_7439_5223# 0.0101f
C1298 RST CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0568f
C1299 VDD a_5146_5223# 0.00891f
C1300 a_11537_1353# CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 4.52e-20
C1301 a_10563_212# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 2.88e-20
C1302 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_10973_1353# 0.069f
C1303 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_0.Q1 8.51e-22
C1304 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 0.00488f
C1305 CLK_div_10_mag_0.JK_FF_mag_0.J RST 1.55e-19
C1306 a_1565_5223# RST 0.00169f
C1307 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00943f
C1308 a_794_1309# CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0732f
C1309 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_2.J 0.0871f
C1310 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 0.0432f
C1311 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.and2_mag_0.OUT 0.065f
C1312 a_9685_1309# a_9845_1309# 0.0504f
C1313 CLK_div_10_mag_0.JK_FF_mag_2.J CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.199f
C1314 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_2123_4126# 0.0732f
C1315 VDD CLK_div_10_mag_0.Q3 1.18f
C1316 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.Q1 1.16f
C1317 VDD CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 1.07f
C1318 a_4576_4126# CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 1.43e-19
C1319 a_9679_212# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 1.17e-20
C1320 a_2129_5223# CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 1.46e-19
C1321 RST a_2283_4126# 8.64e-19
C1322 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_3805_212# 0.0731f
C1323 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.J 0.0334f
C1324 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.321f
C1325 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_10_mag_0.and2_mag_0.OUT 0.0758f
C1326 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT 0.768f
C1327 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 0.00118f
C1328 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT a_7392_1353# 0.00378f
C1329 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0894f
C1330 a_3811_1309# CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.00119f
C1331 VDD CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 0.442f
C1332 VDD a_4582_5223# 0.00123f
C1333 CLK_div_10_mag_1.Q1 a_6875_5223# 0.00859f
C1334 a_10403_212# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 9.1e-19
C1335 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_431_4126# 0.00118f
C1336 CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.00157f
C1337 CLK_div_10_mag_1.JK_FF_mag_2.J a_5300_4126# 0.00111f
C1338 VDD CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 0.397f
C1339 a_1405_5223# RST 0.00128f
C1340 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN a_9510_2450# 0.069f
C1341 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 0.359f
C1342 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.00183f
C1343 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.0622f
C1344 a_9839_212# CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.46e-19
C1345 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.359f
C1346 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_1.QB 2.81e-20
C1347 VDD CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.652f
C1348 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0622f
C1349 a_7386_212# a_7546_212# 0.0504f
C1350 VDD CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 0.653f
C1351 CLK_div_10_mag_0.Q1 a_3645_212# 0.00335f
C1352 VDD a_4529_212# 0.00101f
C1353 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_1559_4126# 0.00378f
C1354 CLK_div_10_mag_0.JK_FF_mag_3.QB a_9845_1309# 1.41e-20
C1355 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 0.122f
C1356 VDD CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.514f
C1357 a_4012_4126# CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 0.011f
C1358 a_11738_2752# CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.00261f
C1359 RST a_2123_4126# 9.22e-19
C1360 VDD a_3858_5223# 0.00152f
C1361 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0378f
C1362 CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 7.08e-20
C1363 CLK_div_10_mag_1.JK_FF_mag_2.J a_277_5223# 0.0811f
C1364 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.nor_3_mag_0.IN3 3.87e-19
C1365 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT a_6828_1309# 0.0732f
C1366 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 5.08e-20
C1367 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_7956_1353# 0.0059f
C1368 CLK_div_10_mag_1.Q1 a_6311_5223# 0.0157f
C1369 VDD a_4422_5223# 0.00101f
C1370 a_11127_256# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00378f
C1371 CLK_div_10_mag_1.JK_FF_mag_2.J a_5140_4126# 9.32e-19
C1372 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.and2_mag_0.OUT 0.026f
C1373 VDD a_5300_4126# 0.00746f
C1374 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 1.29e-19
C1375 CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.36f
C1376 a_2129_5223# CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.0731f
C1377 a_794_1309# CLK_div_10_mag_0.JK_FF_mag_1.QB 0.00392f
C1378 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT RST 0.361f
C1379 a_2486_1353# CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00372f
C1380 CLK_div_10_mag_0.JK_FF_mag_3.QB a_9685_1309# 1.86e-20
C1381 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C1382 a_5146_5223# a_5306_5223# 0.0504f
C1383 a_3448_4126# CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 0.00118f
C1384 RST a_1559_4126# 0.0014f
C1385 a_11578_2752# CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.00239f
C1386 CLK_div_10_mag_1.Q3 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 8.98e-19
C1387 VDD a_3294_5223# 0.00152f
C1388 a_277_5223# VDD 3.14e-19
C1389 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C1390 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_7392_1353# 0.0697f
C1391 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.233f
C1392 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 5.98e-20
C1393 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 8.16e-20
C1394 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT a_6668_1309# 0.0203f
C1395 a_10563_212# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0733f
C1396 CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00101f
C1397 CLK_div_10_mag_0.Q0 a_9839_212# 0.00164f
C1398 CLK_div_10_mag_1.JK_FF_mag_2.J a_4576_4126# 3.12e-19
C1399 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.28f
C1400 RST a_6822_212# 0.00186f
C1401 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 0.0622f
C1402 VDD a_5140_4126# 2.66e-19
C1403 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN a_11578_2752# 2.85e-20
C1404 CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_1.QB 0.0063f
C1405 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT 0.0151f
C1406 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_2123_4126# 0.00119f
C1407 CLK_div_10_mag_1.JK_FF_mag_2.J a_431_4126# 0.0114f
C1408 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00164f
C1409 CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 6.88e-21
C1410 a_1565_5223# CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 9.1e-19
C1411 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_0.Q2 0.0011f
C1412 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.768f
C1413 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.JK_FF_mag_2.J 0.0838f
C1414 a_9839_212# RST 0.00186f
C1415 CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.0592f
C1416 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.103f
C1417 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_1.JK_FF_mag_2.QB 0.28f
C1418 VDD CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.514f
C1419 CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 2.48e-20
C1420 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00118f
C1421 CLK_div_10_mag_0.JK_FF_mag_3.QB a_8520_1353# 0.0114f
C1422 CLK_div_10_mag_1.JK_FF_mag_2.J CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 0.00488f
C1423 CLK_div_10_mag_0.Q1 CLK_div_10_mag_1.Q0 0.0314f
C1424 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_10_mag_0.Q3 8.98e-19
C1425 RST CLK_div_10_mag_1.Q3 0.0465f
C1426 CLK_div_10_mag_1.CLK a_11738_2752# 0.198f
C1427 a_10403_212# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0203f
C1428 CLK_div_10_mag_1.and2_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 2.89e-19
C1429 CLK_div_10_mag_1.JK_FF_mag_2.J a_1565_5223# 0.00695f
C1430 CLK_div_10_mag_1.JK_FF_mag_2.J a_4012_4126# 7.4e-19
C1431 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_4529_212# 2.88e-20
C1432 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C1433 a_4394_3029# CLK_div_10_mag_1.Q1 0.0105f
C1434 VDD a_4576_4126# 3.14e-19
C1435 a_2129_5223# VDD 0.00299f
C1436 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_1559_4126# 1.43e-19
C1437 VDD CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT 0.768f
C1438 VDD a_431_4126# 3.56e-19
C1439 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.0622f
C1440 a_1405_5223# CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 2.88e-20
C1441 VDD CLK_div_10_mag_0.Q2 2.86f
C1442 CLK_div_10_mag_1.JK_FF_mag_1.QB a_8317_4126# 1.86e-20
C1443 CLK_div_10_mag_1.Q0 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 6.82e-19
C1444 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.122f
C1445 CLK_div_10_mag_1.CLK CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 1.48e-20
C1446 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.00183f
C1447 CLK_div_10_mag_1.JK_FF_mag_2.J a_2283_4126# 0.00111f
C1448 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.0635f
C1449 VDD CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 0.397f
C1450 VDD CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.399f
C1451 a_1405_5223# CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 8.64e-19
C1452 CLK_div_10_mag_0.Q1 a_4369_212# 0.0102f
C1453 a_11180_5223# CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 1.46e-19
C1454 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 0.00975f
C1455 VDD a_5657_256# 0.00152f
C1456 CLK_div_10_mag_0.JK_FF_mag_2.J CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.0151f
C1457 CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_10_mag_0.and2_mag_0.OUT 0.144f
C1458 CLK_div_10_mag_1.CLK a_11578_2752# 0.0133f
C1459 VDD CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 1.03f
C1460 CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT 2.81e-20
C1461 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_3.QB 0.311f
C1462 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.109f
C1463 CLK_div_10_mag_1.JK_FF_mag_2.J a_1405_5223# 0.00696f
C1464 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.JK_FF_mag_2.J 9.14e-19
C1465 CLK_div_10_mag_0.JK_FF_mag_0.J VDD 0.496f
C1466 CLK_div_10_mag_1.JK_FF_mag_2.J a_3448_4126# 7.4e-19
C1467 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.J 0.0334f
C1468 a_1565_5223# VDD 2.21e-19
C1469 VDD a_4012_4126# 3.14e-19
C1470 a_230_2335# CLK_div_10_mag_1.Q3 0.019f
C1471 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 0.768f
C1472 RST CLK_div_10_mag_1.nor_3_mag_0.IN3 0.00649f
C1473 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.321f
C1474 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.235f
C1475 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 8.16e-20
C1476 CLK_div_10_mag_0.Q0 a_1922_1353# 6.06e-21
C1477 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_1.Q3 0.0263f
C1478 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.25f
C1479 CLK_div_10_mag_1.JK_FF_mag_1.QB a_8157_4126# 1.41e-20
C1480 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN a_9510_2450# 5.1e-20
C1481 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.0285f
C1482 CLK_div_10_mag_1.Q0 a_2289_5223# 0.00117f
C1483 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 8.16e-20
C1484 CLK_div_10_mag_1.JK_FF_mag_2.J a_2123_4126# 0.00486f
C1485 VDD a_2283_4126# 2.21e-19
C1486 RST CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0759f
C1487 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_10_mag_0.Q3 0.00393f
C1488 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.121f
C1489 a_1922_1353# RST 0.00167f
C1490 CLK_div_10_mag_0.Q0 CLK 0.149f
C1491 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT RST 3.84e-20
C1492 a_11340_5223# CLK_div_10_mag_1.CLK 0.00117f
C1493 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_1.Q1 0.00335f
C1494 CLK_div_10_mag_0.Q3 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00357f
C1495 CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.321f
C1496 a_5503_1353# CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 4.52e-20
C1497 a_634_1309# CLK 0.0101f
C1498 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C1499 VDD a_3448_4126# 3.56e-19
C1500 a_11691_256# VSS 0.0675f
C1501 a_11127_256# VSS 0.0676f
C1502 a_10563_212# VSS 0.0343f
C1503 a_10403_212# VSS 0.0881f
C1504 a_9839_212# VSS 0.0343f
C1505 a_9679_212# VSS 0.0881f
C1506 a_8674_256# VSS 0.0675f
C1507 a_8110_256# VSS 0.0676f
C1508 a_7546_212# VSS 0.0343f
C1509 a_7386_212# VSS 0.0881f
C1510 a_6822_212# VSS 0.0343f
C1511 a_6662_212# VSS 0.0881f
C1512 a_5657_256# VSS 0.0675f
C1513 a_5093_256# VSS 0.0676f
C1514 a_4529_212# VSS 0.0343f
C1515 a_4369_212# VSS 0.0881f
C1516 a_3805_212# VSS 0.0343f
C1517 a_3645_212# VSS 0.0881f
C1518 a_2640_256# VSS 0.0675f
C1519 a_2076_256# VSS 0.0676f
C1520 a_1512_212# VSS 0.0343f
C1521 a_1352_212# VSS 0.0881f
C1522 a_788_212# VSS 0.0343f
C1523 a_628_212# VSS 0.0881f
C1524 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.415f
C1525 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.519f
C1526 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VSS 0.415f
C1527 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VSS 0.539f
C1528 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VSS 0.415f
C1529 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VSS 0.539f
C1530 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.415f
C1531 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.539f
C1532 a_11537_1353# VSS 0.0676f
C1533 a_10973_1353# VSS 0.0676f
C1534 a_10409_1353# VSS 0.0676f
C1535 a_9845_1309# VSS 0.0343f
C1536 a_9685_1309# VSS 0.0881f
C1537 a_8520_1353# VSS 0.0676f
C1538 a_7956_1353# VSS 0.0676f
C1539 a_7392_1353# VSS 0.0676f
C1540 a_6828_1309# VSS 0.0343f
C1541 a_6668_1309# VSS 0.0881f
C1542 a_5503_1353# VSS 0.0676f
C1543 a_4939_1353# VSS 0.0676f
C1544 a_4375_1353# VSS 0.0676f
C1545 a_3811_1309# VSS 0.0343f
C1546 a_3651_1309# VSS 0.0881f
C1547 a_2486_1353# VSS 0.0676f
C1548 a_1922_1353# VSS 0.0676f
C1549 a_1358_1353# VSS 0.0676f
C1550 a_794_1309# VSS 0.0343f
C1551 a_634_1309# VSS 0.0881f
C1552 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.414f
C1553 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.753f
C1554 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.724f
C1555 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.807f
C1556 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C1557 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VSS 0.413f
C1558 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 VSS 0.692f
C1559 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VSS 0.724f
C1560 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VSS 0.808f
C1561 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VSS 0.509f
C1562 CLK_div_10_mag_0.JK_FF_mag_3.QB VSS 0.877f
C1563 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VSS 0.415f
C1564 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 VSS 0.695f
C1565 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VSS 0.724f
C1566 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VSS 0.806f
C1567 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VSS 0.506f
C1568 CLK_div_10_mag_0.JK_FF_mag_2.QB VSS 0.876f
C1569 CLK_div_10_mag_0.JK_FF_mag_2.J VSS 3.11f
C1570 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.412f
C1571 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.772f
C1572 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.723f
C1573 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.806f
C1574 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.508f
C1575 CLK_div_10_mag_0.JK_FF_mag_1.QB VSS 0.888f
C1576 CLK VSS 0.913f
C1577 a_9510_2450# VSS 0.0679f
C1578 a_11738_2752# VSS 0.0371f
C1579 a_11578_2752# VSS 0.038f
C1580 a_8542_2450# VSS 0.0679f
C1581 a_7574_2450# VSS 0.0676f
C1582 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS 0.664f
C1583 CLK_div_10_mag_0.and2_mag_1.OUT VSS 0.701f
C1584 CLK_div_10_mag_0.JK_FF_mag_0.J VSS 0.633f
C1585 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VSS 0.432f
C1586 CLK_div_10_mag_0.Q0 VSS 3.36f
C1587 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VSS 0.438f
C1588 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS 0.433f
C1589 CLK_div_10_mag_0.Q2 VSS 2.2f
C1590 CLK_div_10_mag_0.Q1 VSS 2.59f
C1591 a_4394_3029# VSS 0.0676f
C1592 CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN VSS 0.433f
C1593 a_3426_3029# VSS 0.0679f
C1594 a_390_2335# VSS 0.038f
C1595 a_230_2335# VSS 0.0371f
C1596 CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN VSS 0.438f
C1597 a_2458_3029# VSS 0.0679f
C1598 CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN VSS 0.432f
C1599 CLK_div_10_mag_1.and2_mag_1.OUT VSS 0.701f
C1600 CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS 0.664f
C1601 CLK_div_10_mag_1.nor_3_mag_0.IN3 VSS 0.335f
C1602 CLK_div_10_mag_1.and2_mag_0.OUT VSS 0.601f
C1603 Vdiv100 VSS 0.634f
C1604 CLK_div_10_mag_0.Q3 VSS 1.92f
C1605 CLK_div_10_mag_0.and2_mag_0.OUT VSS 0.599f
C1606 CLK_div_10_mag_0.nor_3_mag_0.IN3 VSS 0.335f
C1607 a_11334_4126# VSS 0.0881f
C1608 a_11174_4126# VSS 0.0343f
C1609 a_10610_4126# VSS 0.0676f
C1610 a_10046_4126# VSS 0.0676f
C1611 a_9482_4126# VSS 0.0676f
C1612 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.508f
C1613 CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.412f
C1614 a_8317_4126# VSS 0.0881f
C1615 a_8157_4126# VSS 0.0343f
C1616 a_7593_4126# VSS 0.0676f
C1617 a_7029_4126# VSS 0.0676f
C1618 a_6465_4126# VSS 0.0676f
C1619 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT VSS 0.506f
C1620 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 VSS 0.415f
C1621 a_5300_4126# VSS 0.0881f
C1622 a_5140_4126# VSS 0.0343f
C1623 a_4576_4126# VSS 0.0676f
C1624 a_4012_4126# VSS 0.0676f
C1625 a_3448_4126# VSS 0.0676f
C1626 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT VSS 0.509f
C1627 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 VSS 0.413f
C1628 a_2283_4126# VSS 0.0881f
C1629 a_2123_4126# VSS 0.0343f
C1630 a_1559_4126# VSS 0.0676f
C1631 a_995_4126# VSS 0.0676f
C1632 a_431_4126# VSS 0.0676f
C1633 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C1634 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.414f
C1635 CLK_div_10_mag_1.JK_FF_mag_0.J VSS 0.598f
C1636 a_11340_5223# VSS 0.0881f
C1637 a_11180_5223# VSS 0.0343f
C1638 a_10616_5223# VSS 0.0881f
C1639 a_10456_5223# VSS 0.0343f
C1640 a_9892_5223# VSS 0.0676f
C1641 a_9328_5223# VSS 0.0675f
C1642 CLK_div_10_mag_1.JK_FF_mag_1.QB VSS 0.888f
C1643 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.806f
C1644 CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.757f
C1645 CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.415f
C1646 a_8323_5223# VSS 0.0881f
C1647 a_8163_5223# VSS 0.0343f
C1648 a_7599_5223# VSS 0.0881f
C1649 a_7439_5223# VSS 0.0343f
C1650 a_6875_5223# VSS 0.0676f
C1651 a_6311_5223# VSS 0.0675f
C1652 CLK_div_10_mag_1.JK_FF_mag_2.QB VSS 0.876f
C1653 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT VSS 0.806f
C1654 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 VSS 0.695f
C1655 CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 VSS 0.415f
C1656 a_5306_5223# VSS 0.0881f
C1657 a_5146_5223# VSS 0.0343f
C1658 a_4582_5223# VSS 0.0881f
C1659 a_4422_5223# VSS 0.0343f
C1660 a_3858_5223# VSS 0.0676f
C1661 a_3294_5223# VSS 0.0675f
C1662 CLK_div_10_mag_1.JK_FF_mag_3.QB VSS 0.877f
C1663 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT VSS 0.808f
C1664 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 VSS 0.692f
C1665 CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 VSS 0.415f
C1666 a_2289_5223# VSS 0.0881f
C1667 a_2129_5223# VSS 0.0343f
C1668 a_1565_5223# VSS 0.0881f
C1669 a_1405_5223# VSS 0.0343f
C1670 a_841_5223# VSS 0.0676f
C1671 a_277_5223# VSS 0.0675f
C1672 CLK_div_10_mag_1.JK_FF_mag_2.J VSS 3.12f
C1673 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.807f
C1674 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.753f
C1675 CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.415f
C1676 CLK_div_10_mag_1.CLK VSS 1.63f
C1677 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.539f
C1678 CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.723f
C1679 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT VSS 0.539f
C1680 CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 VSS 0.724f
C1681 CLK_div_10_mag_1.Q1 VSS 2.99f
C1682 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT VSS 0.539f
C1683 CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 VSS 0.724f
C1684 CLK_div_10_mag_1.Q0 VSS 3.52f
C1685 CLK_div_10_mag_1.Q3 VSS 1.93f
C1686 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.519f
C1687 RST VSS 6.42f
C1688 CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.724f
C1689 VDD VSS 0.135p
C1690 CLK_div_10_mag_1.JK_FF_mag_2.J.t1 VSS 0.0149f
C1691 CLK_div_10_mag_1.JK_FF_mag_2.J.n0 VSS 0.0149f
C1692 CLK_div_10_mag_1.JK_FF_mag_2.J.n1 VSS 0.0318f
C1693 CLK_div_10_mag_1.JK_FF_mag_2.J.t7 VSS 0.0238f
C1694 CLK_div_10_mag_1.JK_FF_mag_2.J.t6 VSS 0.0308f
C1695 CLK_div_10_mag_1.JK_FF_mag_2.J.n2 VSS 0.0609f
C1696 CLK_div_10_mag_1.JK_FF_mag_2.J.t4 VSS 0.0335f
C1697 CLK_div_10_mag_1.JK_FF_mag_2.J.t2 VSS 0.0214f
C1698 CLK_div_10_mag_1.JK_FF_mag_2.J.n3 VSS 0.0593f
C1699 CLK_div_10_mag_1.JK_FF_mag_2.J.n4 VSS 1.14f
C1700 CLK_div_10_mag_1.JK_FF_mag_2.J.t5 VSS 0.0238f
C1701 CLK_div_10_mag_1.JK_FF_mag_2.J.t3 VSS 0.0191f
C1702 CLK_div_10_mag_1.JK_FF_mag_2.J.n5 VSS 0.0566f
C1703 CLK_div_10_mag_1.JK_FF_mag_2.J.n6 VSS 0.381f
C1704 CLK_div_10_mag_1.JK_FF_mag_2.J.n7 VSS 0.0932f
C1705 CLK_div_10_mag_1.Q2.t1 VSS 0.02f
C1706 CLK_div_10_mag_1.Q2.t0 VSS 0.0165f
C1707 CLK_div_10_mag_1.Q2.n0 VSS 0.0165f
C1708 CLK_div_10_mag_1.Q2.n1 VSS 0.0396f
C1709 CLK_div_10_mag_1.Q2.t10 VSS 0.0367f
C1710 CLK_div_10_mag_1.Q2.t9 VSS 0.0242f
C1711 CLK_div_10_mag_1.Q2.n2 VSS 0.0652f
C1712 CLK_div_10_mag_1.Q2.t4 VSS 0.0263f
C1713 CLK_div_10_mag_1.Q2.t3 VSS 0.0211f
C1714 CLK_div_10_mag_1.Q2.n3 VSS 0.0612f
C1715 CLK_div_10_mag_1.Q2.n4 VSS 0.486f
C1716 CLK_div_10_mag_1.Q2.t6 VSS 0.019f
C1717 CLK_div_10_mag_1.Q2.t7 VSS 0.034f
C1718 CLK_div_10_mag_1.Q2.n5 VSS 0.0648f
C1719 CLK_div_10_mag_1.Q2.t8 VSS 0.0263f
C1720 CLK_div_10_mag_1.Q2.t11 VSS 0.0211f
C1721 CLK_div_10_mag_1.Q2.n6 VSS 0.0612f
C1722 CLK_div_10_mag_1.Q2.n7 VSS 0.325f
C1723 CLK_div_10_mag_1.Q2.t12 VSS 0.0263f
C1724 CLK_div_10_mag_1.Q2.t5 VSS 0.0211f
C1725 CLK_div_10_mag_1.Q2.n8 VSS 0.0612f
C1726 CLK_div_10_mag_1.Q2.n9 VSS 0.308f
C1727 CLK_div_10_mag_1.Q2.n10 VSS 0.15f
C1728 CLK_div_10_mag_0.JK_FF_mag_2.J.n0 VSS 0.0848f
C1729 CLK_div_10_mag_0.JK_FF_mag_2.J.t4 VSS 0.0183f
C1730 CLK_div_10_mag_0.JK_FF_mag_2.J.t5 VSS 0.0229f
C1731 CLK_div_10_mag_0.JK_FF_mag_2.J.n1 VSS 0.0543f
C1732 CLK_div_10_mag_0.JK_FF_mag_2.J.t6 VSS 0.0322f
C1733 CLK_div_10_mag_0.JK_FF_mag_2.J.t8 VSS 0.0205f
C1734 CLK_div_10_mag_0.JK_FF_mag_2.J.n2 VSS 0.0569f
C1735 CLK_div_10_mag_0.JK_FF_mag_2.J.t3 VSS 0.0296f
C1736 CLK_div_10_mag_0.JK_FF_mag_2.J.t7 VSS 0.0228f
C1737 CLK_div_10_mag_0.JK_FF_mag_2.J.n3 VSS 0.0585f
C1738 CLK_div_10_mag_0.JK_FF_mag_2.J.n4 VSS 1.1f
C1739 CLK_div_10_mag_0.JK_FF_mag_2.J.n5 VSS 0.366f
C1740 CLK_div_10_mag_0.JK_FF_mag_2.J.t0 VSS 0.0143f
C1741 CLK_div_10_mag_0.JK_FF_mag_2.J.n6 VSS 0.0143f
C1742 CLK_div_10_mag_0.JK_FF_mag_2.J.n7 VSS 0.0338f
C1743 RST.t5 VSS 0.0404f
C1744 RST.t3 VSS 0.0266f
C1745 RST.n0 VSS 0.0713f
C1746 RST.n1 VSS 0.00918f
C1747 RST.t4 VSS 0.0266f
C1748 RST.t7 VSS 0.0404f
C1749 RST.n2 VSS 0.0714f
C1750 RST.n3 VSS 0.0364f
C1751 RST.n4 VSS 0.00894f
C1752 RST.n5 VSS 0.0205f
C1753 RST.n6 VSS 0.00329f
C1754 RST.t8 VSS 0.0254f
C1755 RST.n7 VSS 0.0232f
C1756 RST.t9 VSS 0.0403f
C1757 RST.n8 VSS 0.0494f
C1758 RST.n9 VSS 3.9e-19
C1759 RST.n10 VSS 0.00328f
C1760 RST.n11 VSS 0.00309f
C1761 RST.n12 VSS 0.0164f
C1762 RST.t10 VSS 0.0266f
C1763 RST.t13 VSS 0.0404f
C1764 RST.n13 VSS 0.0714f
C1765 RST.n14 VSS 0.0384f
C1766 RST.t2 VSS 0.0266f
C1767 RST.t6 VSS 0.0404f
C1768 RST.n15 VSS 0.0714f
C1769 RST.n16 VSS 0.389f
C1770 RST.n17 VSS 1.21f
C1771 RST.n18 VSS 1f
C1772 RST.n19 VSS 0.575f
C1773 RST.n20 VSS 0.00329f
C1774 RST.n21 VSS 0.00317f
C1775 RST.t1 VSS 0.0404f
C1776 RST.t0 VSS 0.0266f
C1777 RST.n22 VSS 0.0713f
C1778 RST.n23 VSS 0.00918f
C1779 RST.n24 VSS 0.00334f
C1780 RST.n25 VSS 0.0209f
C1781 RST.n26 VSS 0.0161f
C1782 RST.t15 VSS 0.0408f
C1783 RST.t14 VSS 0.0258f
C1784 RST.n27 VSS 0.0717f
C1785 RST.n28 VSS 0.0385f
C1786 RST.t12 VSS 0.0404f
C1787 RST.t11 VSS 0.0266f
C1788 RST.n29 VSS 0.0714f
C1789 RST.n30 VSS 0.0371f
C1790 RST.n31 VSS 1.02f
C1791 RST.n32 VSS 1.01f
C1792 RST.n33 VSS 1.07f
C1793 RST.n34 VSS 0.0159f
C1794 RST.n35 VSS 0.0206f
C1795 RST.n36 VSS 0.00334f
C1796 RST.n37 VSS 0.00317f
C1797 RST.n38 VSS 0.0024f
C1798 RST.n39 VSS 0.00277f
C1799 CLK_div_10_mag_1.Q0.n0 VSS 0.826f
C1800 CLK_div_10_mag_1.Q0.n1 VSS 0.0344f
C1801 CLK_div_10_mag_1.Q0.n2 VSS 0.254f
C1802 CLK_div_10_mag_1.Q0.n3 VSS 0.0151f
C1803 CLK_div_10_mag_1.Q0.n4 VSS 0.241f
C1804 CLK_div_10_mag_1.Q0.n5 VSS 0.0151f
C1805 CLK_div_10_mag_1.Q0.n6 VSS 0.15f
C1806 CLK_div_10_mag_1.Q0.n7 VSS 0.103f
C1807 CLK_div_10_mag_1.Q0.n8 VSS 0.103f
C1808 CLK_div_10_mag_1.Q0.n9 VSS 0.035f
C1809 CLK_div_10_mag_1.Q0.t2 VSS 0.0201f
C1810 CLK_div_10_mag_1.Q0.t0 VSS 0.0165f
C1811 CLK_div_10_mag_1.Q0.n10 VSS 0.0165f
C1812 CLK_div_10_mag_1.Q0.n11 VSS 0.0397f
C1813 CLK_div_10_mag_1.Q0.n12 VSS 0.124f
C1814 CLK_div_10_mag_1.Q0.t13 VSS 0.0368f
C1815 CLK_div_10_mag_1.Q0.t12 VSS 0.0243f
C1816 CLK_div_10_mag_1.Q0.n13 VSS 0.0654f
C1817 CLK_div_10_mag_1.Q0.n14 VSS 0.257f
C1818 CLK_div_10_mag_1.Q0.t17 VSS 0.0264f
C1819 CLK_div_10_mag_1.Q0.t15 VSS 0.0211f
C1820 CLK_div_10_mag_1.Q0.n15 VSS 0.0614f
C1821 CLK_div_10_mag_1.Q0.n16 VSS 0.0381f
C1822 CLK_div_10_mag_1.Q0.n17 VSS 0.488f
C1823 CLK_div_10_mag_1.Q0.t3 VSS 0.0368f
C1824 CLK_div_10_mag_1.Q0.t19 VSS 0.0243f
C1825 CLK_div_10_mag_1.Q0.n18 VSS 0.0651f
C1826 CLK_div_10_mag_1.Q0.t18 VSS 0.0368f
C1827 CLK_div_10_mag_1.Q0.t16 VSS 0.0243f
C1828 CLK_div_10_mag_1.Q0.n19 VSS 0.0651f
C1829 CLK_div_10_mag_1.Q0.t7 VSS 0.0304f
C1830 CLK_div_10_mag_1.Q0.t11 VSS 0.00786f
C1831 CLK_div_10_mag_1.Q0.n20 VSS 0.0504f
C1832 CLK_div_10_mag_1.Q0.t9 VSS 0.0368f
C1833 CLK_div_10_mag_1.Q0.t8 VSS 0.0243f
C1834 CLK_div_10_mag_1.Q0.n21 VSS 0.0651f
C1835 CLK_div_10_mag_1.Q0.t6 VSS 0.0368f
C1836 CLK_div_10_mag_1.Q0.t4 VSS 0.0243f
C1837 CLK_div_10_mag_1.Q0.n22 VSS 0.0651f
C1838 CLK_div_10_mag_1.Q0.n23 VSS 0.11f
C1839 CLK_div_10_mag_1.Q0.t5 VSS 0.0342f
C1840 CLK_div_10_mag_1.Q0.t14 VSS 0.0189f
C1841 CLK_div_10_mag_1.Q0.n24 VSS 0.0652f
C1842 CLK_div_10_mag_1.Q0.n25 VSS 0.869f
C1843 CLK_div_10_mag_1.Q0.t10 VSS 0.0304f
C1844 CLK_div_10_mag_1.Q0.t20 VSS 0.00786f
C1845 CLK_div_10_mag_1.Q0.n26 VSS 0.0504f
C1846 CLK_div_10_mag_1.Q0.n27 VSS 0.124f
C1847 CLK_div_10_mag_1.Q0.n28 VSS 0.0156f
C1848 VDD.n0 VSS 0.0293f
C1849 VDD.t38 VSS 0.0024f
C1850 VDD.n1 VSS 0.0024f
C1851 VDD.n2 VSS 0.00524f
C1852 VDD.n3 VSS 0.0312f
C1853 VDD.t151 VSS 0.00583f
C1854 VDD.t51 VSS 0.0414f
C1855 VDD.n4 VSS 0.00583f
C1856 VDD.t52 VSS 0.00583f
C1857 VDD.n5 VSS 0.00583f
C1858 VDD.n6 VSS 0.0289f
C1859 VDD.t34 VSS 0.0613f
C1860 VDD.n7 VSS 0.00583f
C1861 VDD.t415 VSS 0.00581f
C1862 VDD.t458 VSS 0.00583f
C1863 VDD.n8 VSS 0.0275f
C1864 VDD.t414 VSS 0.0515f
C1865 VDD.t416 VSS 0.0399f
C1866 VDD.t192 VSS 0.0024f
C1867 VDD.n9 VSS 0.0024f
C1868 VDD.n10 VSS 0.00524f
C1869 VDD.t281 VSS 0.00583f
C1870 VDD.n11 VSS 0.00583f
C1871 VDD.n12 VSS 0.0289f
C1872 VDD.t116 VSS 0.077f
C1873 VDD.n13 VSS 0.00583f
C1874 VDD.t456 VSS 0.00583f
C1875 VDD.n14 VSS 0.00583f
C1876 VDD.n15 VSS 0.00583f
C1877 VDD.t268 VSS 0.0759f
C1878 VDD.n16 VSS 0.0362f
C1879 VDD.t361 VSS 0.00583f
C1880 VDD.n17 VSS 0.00583f
C1881 VDD.t360 VSS 0.0703f
C1882 VDD.t113 VSS 0.077f
C1883 VDD.n18 VSS 0.0362f
C1884 VDD.t74 VSS 0.00583f
C1885 VDD.t265 VSS 0.0024f
C1886 VDD.n19 VSS 0.0024f
C1887 VDD.n20 VSS 0.00524f
C1888 VDD.t73 VSS 0.0703f
C1889 VDD.t264 VSS 0.0859f
C1890 VDD.t323 VSS 0.0399f
C1891 VDD.n21 VSS 0.0362f
C1892 VDD.t349 VSS 0.00583f
C1893 VDD.t272 VSS 0.0024f
C1894 VDD.n22 VSS 0.0024f
C1895 VDD.n23 VSS 0.00524f
C1896 VDD.t348 VSS 0.0703f
C1897 VDD.t271 VSS 0.0859f
C1898 VDD.t423 VSS 0.0399f
C1899 VDD.t147 VSS 0.0701f
C1900 VDD.n24 VSS 0.0362f
C1901 VDD.t148 VSS 0.00545f
C1902 VDD.t146 VSS 0.005f
C1903 VDD.t491 VSS 0.00379f
C1904 VDD.n25 VSS 0.00977f
C1905 VDD.n26 VSS 0.00173f
C1906 VDD.t177 VSS 0.005f
C1907 VDD.t478 VSS 0.00379f
C1908 VDD.n27 VSS 0.00978f
C1909 VDD.n28 VSS 0.0023f
C1910 VDD.n29 VSS 0.00119f
C1911 VDD.n30 VSS 6e-19
C1912 VDD.n31 VSS 0.00534f
C1913 VDD.n32 VSS 5.77e-19
C1914 VDD.t163 VSS 0.00486f
C1915 VDD.n33 VSS 0.0048f
C1916 VDD.t485 VSS 0.00378f
C1917 VDD.n34 VSS 0.00162f
C1918 VDD.n35 VSS 0.00513f
C1919 VDD.n36 VSS 0.00177f
C1920 VDD.n37 VSS 0.00146f
C1921 VDD.t166 VSS 0.00498f
C1922 VDD.t479 VSS 0.0038f
C1923 VDD.n38 VSS 0.0098f
C1924 VDD.n39 VSS 0.00184f
C1925 VDD.n40 VSS 0.00156f
C1926 VDD.n41 VSS 6e-19
C1927 VDD.n42 VSS 0.0189f
C1928 VDD.n43 VSS 0.0733f
C1929 VDD.n44 VSS 0.107f
C1930 VDD.t490 VSS 0.00387f
C1931 VDD.t160 VSS 0.00491f
C1932 VDD.n45 VSS 0.00979f
C1933 VDD.n46 VSS 0.00357f
C1934 VDD.n47 VSS 0.00146f
C1935 VDD.t484 VSS 0.0038f
C1936 VDD.t149 VSS 0.00498f
C1937 VDD.n48 VSS 0.0098f
C1938 VDD.n49 VSS 0.00191f
C1939 VDD.n50 VSS 0.0015f
C1940 VDD.n51 VSS 6e-19
C1941 VDD.n52 VSS 0.0189f
C1942 VDD.n53 VSS 0.0247f
C1943 VDD.n54 VSS 0.119f
C1944 VDD.n55 VSS 0.0499f
C1945 VDD.n56 VSS 0.00472f
C1946 VDD.n57 VSS 0.0135f
C1947 VDD.n58 VSS 0.0333f
C1948 VDD.n59 VSS 0.0332f
C1949 VDD.n60 VSS 0.0341f
C1950 VDD.n61 VSS 0.0181f
C1951 VDD.n62 VSS 0.0332f
C1952 VDD.n63 VSS 0.034f
C1953 VDD.n64 VSS 0.0201f
C1954 VDD.n65 VSS 0.0289f
C1955 VDD.n66 VSS 0.0269f
C1956 VDD.n67 VSS 0.0201f
C1957 VDD.n68 VSS 0.055f
C1958 VDD.n69 VSS 0.0625f
C1959 VDD.t362 VSS 0.0759f
C1960 VDD.t455 VSS 0.0703f
C1961 VDD.n70 VSS 0.0362f
C1962 VDD.n71 VSS 0.0201f
C1963 VDD.n72 VSS 0.0269f
C1964 VDD.n73 VSS 0.0289f
C1965 VDD.t267 VSS 0.00583f
C1966 VDD.n74 VSS 0.0269f
C1967 VDD.n75 VSS 0.0201f
C1968 VDD.n76 VSS 0.0362f
C1969 VDD.t266 VSS 0.0703f
C1970 VDD.t75 VSS 0.077f
C1971 VDD.t191 VSS 0.0859f
C1972 VDD.t280 VSS 0.0703f
C1973 VDD.n77 VSS 0.0362f
C1974 VDD.n78 VSS 0.0201f
C1975 VDD.n79 VSS 0.0254f
C1976 VDD.n80 VSS 0.0238f
C1977 VDD.n81 VSS 0.0181f
C1978 VDD.n82 VSS 0.0362f
C1979 VDD.t457 VSS 0.0399f
C1980 VDD.n83 VSS 0.0542f
C1981 VDD.n84 VSS 0.0183f
C1982 VDD.n85 VSS 0.00583f
C1983 VDD.t439 VSS 0.0759f
C1984 VDD.n86 VSS 0.0362f
C1985 VDD.t225 VSS 0.00583f
C1986 VDD.n87 VSS 0.00583f
C1987 VDD.t224 VSS 0.0703f
C1988 VDD.t100 VSS 0.077f
C1989 VDD.n88 VSS 0.0362f
C1990 VDD.t112 VSS 0.00583f
C1991 VDD.t54 VSS 0.0024f
C1992 VDD.n89 VSS 0.0024f
C1993 VDD.n90 VSS 0.00524f
C1994 VDD.t111 VSS 0.0703f
C1995 VDD.t53 VSS 0.0859f
C1996 VDD.t141 VSS 0.0399f
C1997 VDD.n91 VSS 0.0362f
C1998 VDD.t120 VSS 0.00583f
C1999 VDD.t445 VSS 0.0024f
C2000 VDD.n92 VSS 0.0024f
C2001 VDD.n93 VSS 0.00524f
C2002 VDD.t119 VSS 0.0703f
C2003 VDD.t444 VSS 0.0859f
C2004 VDD.t10 VSS 0.0399f
C2005 VDD.t161 VSS 0.0701f
C2006 VDD.n94 VSS 0.0362f
C2007 VDD.t162 VSS 0.00625f
C2008 VDD.n95 VSS 0.0449f
C2009 VDD.n96 VSS 0.0332f
C2010 VDD.n97 VSS 0.0341f
C2011 VDD.n98 VSS 0.0181f
C2012 VDD.n99 VSS 0.0332f
C2013 VDD.n100 VSS 0.034f
C2014 VDD.n101 VSS 0.0201f
C2015 VDD.n102 VSS 0.0289f
C2016 VDD.n103 VSS 0.0269f
C2017 VDD.n104 VSS 0.0201f
C2018 VDD.n105 VSS 0.0517f
C2019 VDD.n106 VSS 0.0413f
C2020 VDD.n107 VSS 0.0296f
C2021 VDD.t42 VSS 0.00583f
C2022 VDD.n108 VSS 0.0269f
C2023 VDD.n109 VSS 0.0201f
C2024 VDD.n110 VSS 0.0312f
C2025 VDD.t41 VSS 0.0559f
C2026 VDD.t97 VSS 0.0613f
C2027 VDD.n111 VSS 0.0312f
C2028 VDD.n112 VSS 0.0201f
C2029 VDD.n113 VSS 0.0269f
C2030 VDD.n114 VSS 0.0289f
C2031 VDD.t296 VSS 0.00583f
C2032 VDD.n115 VSS 0.0191f
C2033 VDD.n116 VSS 0.0201f
C2034 VDD.t13 VSS 0.0317f
C2035 VDD.t37 VSS 0.0683f
C2036 VDD.t295 VSS 0.0559f
C2037 VDD.n117 VSS 0.0312f
C2038 VDD.t108 VSS 0.0269f
C2039 VDD.n118 VSS 0.162f
C2040 VDD.t150 VSS 0.0317f
C2041 VDD.n119 VSS 0.0894f
C2042 VDD.t18 VSS 0.0643f
C2043 VDD.t19 VSS 0.00581f
C2044 VDD.n120 VSS 0.00583f
C2045 VDD.t326 VSS 0.0613f
C2046 VDD.n121 VSS 0.0312f
C2047 VDD.t322 VSS 0.00583f
C2048 VDD.n122 VSS 0.00583f
C2049 VDD.t321 VSS 0.0559f
C2050 VDD.t244 VSS 0.0613f
C2051 VDD.n123 VSS 0.0312f
C2052 VDD.t90 VSS 0.00583f
C2053 VDD.n124 VSS 0.00583f
C2054 VDD.n125 VSS 0.0312f
C2055 VDD.t125 VSS 0.00583f
C2056 VDD.t330 VSS 0.0024f
C2057 VDD.n126 VSS 0.0024f
C2058 VDD.n127 VSS 0.00524f
C2059 VDD.t124 VSS 0.0559f
C2060 VDD.t329 VSS 0.0683f
C2061 VDD.t406 VSS 0.0317f
C2062 VDD.n128 VSS 0.0312f
C2063 VDD.t93 VSS 0.00583f
C2064 VDD.t89 VSS 0.0414f
C2065 VDD.t350 VSS 0.0269f
C2066 VDD.n129 VSS 0.162f
C2067 VDD.t92 VSS 0.0317f
C2068 VDD.n130 VSS 0.0894f
C2069 VDD.t421 VSS 0.0643f
C2070 VDD.t422 VSS 0.00581f
C2071 VDD.n131 VSS 0.00583f
C2072 VDD.t231 VSS 0.0613f
C2073 VDD.n132 VSS 0.0312f
C2074 VDD.t389 VSS 0.00583f
C2075 VDD.n133 VSS 0.00583f
C2076 VDD.t388 VSS 0.0559f
C2077 VDD.t277 VSS 0.0613f
C2078 VDD.n134 VSS 0.0312f
C2079 VDD.t215 VSS 0.00583f
C2080 VDD.n135 VSS 0.00583f
C2081 VDD.n136 VSS 0.0312f
C2082 VDD.t464 VSS 0.00583f
C2083 VDD.t235 VSS 0.0024f
C2084 VDD.n137 VSS 0.0024f
C2085 VDD.n138 VSS 0.00526f
C2086 VDD.t214 VSS 0.0219f
C2087 VDD.t218 VSS 0.0464f
C2088 VDD.n139 VSS 0.178f
C2089 VDD.t463 VSS 0.0559f
C2090 VDD.t234 VSS 0.0683f
C2091 VDD.t374 VSS 0.0294f
C2092 VDD.t31 VSS 0.0483f
C2093 VDD.n140 VSS 0.00592f
C2094 VDD.n141 VSS 0.00581f
C2095 VDD.n142 VSS 0.0205f
C2096 VDD.t228 VSS 0.0828f
C2097 VDD.t338 VSS 0.04f
C2098 VDD.n143 VSS 0.00583f
C2099 VDD.n144 VSS 0.00581f
C2100 VDD.n145 VSS 0.0205f
C2101 VDD.t43 VSS 0.0518f
C2102 VDD.t105 VSS 0.04f
C2103 VDD.n146 VSS 0.00583f
C2104 VDD.n147 VSS 0.00581f
C2105 VDD.n148 VSS 0.0205f
C2106 VDD.t249 VSS 0.0518f
C2107 VDD.t307 VSS 0.0703f
C2108 VDD.n149 VSS 0.00583f
C2109 VDD.n150 VSS 0.00583f
C2110 VDD.t153 VSS 0.04f
C2111 VDD.n151 VSS 0.00583f
C2112 VDD.n152 VSS 0.00581f
C2113 VDD.t306 VSS 0.00583f
C2114 VDD.t55 VSS 0.0705f
C2115 VDD.n153 VSS 0.00583f
C2116 VDD.t294 VSS 0.0024f
C2117 VDD.n154 VSS 0.0024f
C2118 VDD.n155 VSS 0.00524f
C2119 VDD.n156 VSS 0.00583f
C2120 VDD.n157 VSS 0.0341f
C2121 VDD.t157 VSS 0.0703f
C2122 VDD.n158 VSS 0.00625f
C2123 VDD.t379 VSS 0.0024f
C2124 VDD.n159 VSS 0.0024f
C2125 VDD.n160 VSS 0.00524f
C2126 VDD.n161 VSS 0.0333f
C2127 VDD.n162 VSS 0.0449f
C2128 VDD.n163 VSS 0.0362f
C2129 VDD.t378 VSS 0.0397f
C2130 VDD.t300 VSS 0.0859f
C2131 VDD.t465 VSS 0.0705f
C2132 VDD.t28 VSS 0.0859f
C2133 VDD.t293 VSS 0.0397f
C2134 VDD.n164 VSS 0.0362f
C2135 VDD.n165 VSS 0.018f
C2136 VDD.n166 VSS 0.0333f
C2137 VDD.n167 VSS 0.034f
C2138 VDD.t1 VSS 0.00583f
C2139 VDD.n168 VSS 0.00583f
C2140 VDD.n169 VSS 0.0268f
C2141 VDD.n170 VSS 0.0289f
C2142 VDD.n171 VSS 0.0202f
C2143 VDD.n172 VSS 0.0362f
C2144 VDD.t0 VSS 0.0769f
C2145 VDD.t78 VSS 0.0705f
C2146 VDD.t305 VSS 0.0758f
C2147 VDD.n173 VSS 0.0362f
C2148 VDD.n174 VSS 0.0202f
C2149 VDD.n175 VSS 0.0516f
C2150 VDD.t292 VSS 0.00583f
C2151 VDD.t25 VSS 0.0705f
C2152 VDD.n176 VSS 0.00583f
C2153 VDD.t59 VSS 0.00583f
C2154 VDD.t395 VSS 0.04f
C2155 VDD.n177 VSS 0.00583f
C2156 VDD.n178 VSS 0.00581f
C2157 VDD.t394 VSS 0.00583f
C2158 VDD.t398 VSS 0.0705f
C2159 VDD.n179 VSS 0.00583f
C2160 VDD.t145 VSS 0.0024f
C2161 VDD.n180 VSS 0.0024f
C2162 VDD.n181 VSS 0.00524f
C2163 VDD.n182 VSS 0.00583f
C2164 VDD.n183 VSS 0.0341f
C2165 VDD.t174 VSS 0.0703f
C2166 VDD.n184 VSS 0.00625f
C2167 VDD.t429 VSS 0.0024f
C2168 VDD.n185 VSS 0.0024f
C2169 VDD.n186 VSS 0.00524f
C2170 VDD.n187 VSS 0.0333f
C2171 VDD.n188 VSS 0.0449f
C2172 VDD.n189 VSS 0.0362f
C2173 VDD.t428 VSS 0.0397f
C2174 VDD.t371 VSS 0.0859f
C2175 VDD.t385 VSS 0.0705f
C2176 VDD.t81 VSS 0.0859f
C2177 VDD.t144 VSS 0.0397f
C2178 VDD.n190 VSS 0.0362f
C2179 VDD.n191 VSS 0.018f
C2180 VDD.n192 VSS 0.0333f
C2181 VDD.n193 VSS 0.034f
C2182 VDD.t471 VSS 0.00583f
C2183 VDD.n194 VSS 0.00583f
C2184 VDD.n195 VSS 0.0268f
C2185 VDD.n196 VSS 0.0289f
C2186 VDD.n197 VSS 0.0202f
C2187 VDD.n198 VSS 0.0362f
C2188 VDD.t470 VSS 0.0769f
C2189 VDD.t449 VSS 0.0705f
C2190 VDD.t393 VSS 0.0758f
C2191 VDD.n199 VSS 0.0362f
C2192 VDD.n200 VSS 0.0202f
C2193 VDD.n201 VSS 0.0516f
C2194 VDD.t240 VSS 0.00583f
C2195 VDD.t84 VSS 0.0705f
C2196 VDD.n202 VSS 0.00583f
C2197 VDD.t402 VSS 0.00583f
C2198 VDD.n203 VSS 0.0569f
C2199 VDD.t381 VSS 0.0226f
C2200 VDD.n204 VSS 0.00583f
C2201 VDD.n205 VSS 0.00608f
C2202 VDD.t273 VSS 0.192f
C2203 VDD.t91 VSS 0.0688f
C2204 VDD.t185 VSS 0.0546f
C2205 VDD.t380 VSS 0.0856f
C2206 VDD.n206 VSS 0.0739f
C2207 VDD.n207 VSS 0.0101f
C2208 VDD.n208 VSS 0.0256f
C2209 VDD.n209 VSS 0.0274f
C2210 VDD.n210 VSS 0.0169f
C2211 VDD.n211 VSS 0.00583f
C2212 VDD.n212 VSS 0.0254f
C2213 VDD.t431 VSS 0.0024f
C2214 VDD.n213 VSS 0.0024f
C2215 VDD.n214 VSS 0.00526f
C2216 VDD.n215 VSS 0.0184f
C2217 VDD.n216 VSS 0.0262f
C2218 VDD.t40 VSS 0.00581f
C2219 VDD.n217 VSS 0.0276f
C2220 VDD.n218 VSS 0.0192f
C2221 VDD.t196 VSS 0.00592f
C2222 VDD.n219 VSS 0.0317f
C2223 VDD.n220 VSS 0.00583f
C2224 VDD.t356 VSS 0.00581f
C2225 VDD.n221 VSS 0.0205f
C2226 VDD.n222 VSS 0.0287f
C2227 VDD.n223 VSS 0.0204f
C2228 VDD.t413 VSS 0.00583f
C2229 VDD.n224 VSS 0.0272f
C2230 VDD.t205 VSS 0.0517f
C2231 VDD.n225 VSS 0.00583f
C2232 VDD.t206 VSS 0.00581f
C2233 VDD.n226 VSS 0.0205f
C2234 VDD.n227 VSS 0.0287f
C2235 VDD.n228 VSS 0.0204f
C2236 VDD.t448 VSS 0.00583f
C2237 VDD.n229 VSS 0.0272f
C2238 VDD.t468 VSS 0.0517f
C2239 VDD.t16 VSS 0.0701f
C2240 VDD.n230 VSS 0.00583f
C2241 VDD.t469 VSS 0.00581f
C2242 VDD.n231 VSS 0.0205f
C2243 VDD.n232 VSS 0.0287f
C2244 VDD.t17 VSS 0.00583f
C2245 VDD.n233 VSS 0.0525f
C2246 VDD.n234 VSS 0.0204f
C2247 VDD.n235 VSS 0.0362f
C2248 VDD.t436 VSS 0.046f
C2249 VDD.n236 VSS 0.0847f
C2250 VDD.t447 VSS 0.0399f
C2251 VDD.n237 VSS 0.0362f
C2252 VDD.t7 VSS 0.046f
C2253 VDD.n238 VSS 0.0847f
C2254 VDD.t412 VSS 0.0399f
C2255 VDD.n239 VSS 0.0362f
C2256 VDD.t442 VSS 0.046f
C2257 VDD.n240 VSS 0.0538f
C2258 VDD.t355 VSS 0.0824f
C2259 VDD.t195 VSS 0.0486f
C2260 VDD.n241 VSS 0.0822f
C2261 VDD.t39 VSS 0.0746f
C2262 VDD.n242 VSS 0.0449f
C2263 VDD.n243 VSS 0.0565f
C2264 VDD.t430 VSS 0.037f
C2265 VDD.t236 VSS 0.0859f
C2266 VDD.t94 VSS 0.0705f
C2267 VDD.t401 VSS 0.0769f
C2268 VDD.n244 VSS 0.0362f
C2269 VDD.n245 VSS 0.0202f
C2270 VDD.n246 VSS 0.0289f
C2271 VDD.n247 VSS 0.0268f
C2272 VDD.t473 VSS 0.00583f
C2273 VDD.n248 VSS 0.00583f
C2274 VDD.n249 VSS 0.0268f
C2275 VDD.n250 VSS 0.0289f
C2276 VDD.n251 VSS 0.0202f
C2277 VDD.n252 VSS 0.0362f
C2278 VDD.t472 VSS 0.0769f
C2279 VDD.t126 VSS 0.0705f
C2280 VDD.t239 VSS 0.0758f
C2281 VDD.n253 VSS 0.0362f
C2282 VDD.n254 VSS 0.0202f
C2283 VDD.n255 VSS 0.0296f
C2284 VDD.n256 VSS 0.0365f
C2285 VDD.n257 VSS 0.0179f
C2286 VDD.t368 VSS 0.0516f
C2287 VDD.n258 VSS 0.0542f
C2288 VDD.n259 VSS 0.0276f
C2289 VDD.t335 VSS 0.0024f
C2290 VDD.n260 VSS 0.0024f
C2291 VDD.n261 VSS 0.00524f
C2292 VDD.n262 VSS 0.00583f
C2293 VDD.n263 VSS 0.0254f
C2294 VDD.n264 VSS 0.0238f
C2295 VDD.n265 VSS 0.018f
C2296 VDD.n266 VSS 0.0362f
C2297 VDD.t334 VSS 0.0397f
C2298 VDD.t288 VSS 0.0859f
C2299 VDD.t255 VSS 0.0705f
C2300 VDD.t58 VSS 0.0769f
C2301 VDD.n267 VSS 0.0362f
C2302 VDD.n268 VSS 0.0202f
C2303 VDD.n269 VSS 0.0289f
C2304 VDD.n270 VSS 0.0268f
C2305 VDD.t3 VSS 0.00583f
C2306 VDD.n271 VSS 0.00583f
C2307 VDD.n272 VSS 0.0268f
C2308 VDD.n273 VSS 0.0289f
C2309 VDD.n274 VSS 0.0202f
C2310 VDD.n275 VSS 0.0362f
C2311 VDD.t2 VSS 0.0769f
C2312 VDD.t4 VSS 0.0705f
C2313 VDD.t291 VSS 0.0758f
C2314 VDD.n276 VSS 0.0362f
C2315 VDD.n277 VSS 0.0202f
C2316 VDD.n278 VSS 0.0296f
C2317 VDD.n279 VSS 0.0412f
C2318 VDD.n280 VSS 0.0183f
C2319 VDD.t312 VSS 0.0516f
C2320 VDD.n281 VSS 0.0542f
C2321 VDD.n282 VSS 0.0276f
C2322 VDD.t304 VSS 0.0024f
C2323 VDD.n283 VSS 0.0024f
C2324 VDD.n284 VSS 0.00524f
C2325 VDD.n285 VSS 0.0238f
C2326 VDD.n286 VSS 0.018f
C2327 VDD.n287 VSS 0.0362f
C2328 VDD.t303 VSS 0.0397f
C2329 VDD.t343 VSS 0.0859f
C2330 VDD.t258 VSS 0.0705f
C2331 VDD.n288 VSS 0.0362f
C2332 VDD.t211 VSS 0.00583f
C2333 VDD.n289 VSS 0.00583f
C2334 VDD.t210 VSS 0.0769f
C2335 VDD.t282 VSS 0.0705f
C2336 VDD.n290 VSS 0.0362f
C2337 VDD.t318 VSS 0.00583f
C2338 VDD.n291 VSS 0.00583f
C2339 VDD.t317 VSS 0.0769f
C2340 VDD.t252 VSS 0.0705f
C2341 VDD.t341 VSS 0.0758f
C2342 VDD.n292 VSS 0.0362f
C2343 VDD.t342 VSS 0.00583f
C2344 VDD.n293 VSS 0.00581f
C2345 VDD.t136 VSS 0.0516f
C2346 VDD.n294 VSS 0.0542f
C2347 VDD.n295 VSS 0.00583f
C2348 VDD.t297 VSS 0.04f
C2349 VDD.n296 VSS 0.0362f
C2350 VDD.t337 VSS 0.0024f
C2351 VDD.n297 VSS 0.0024f
C2352 VDD.n298 VSS 0.00524f
C2353 VDD.n299 VSS 0.00583f
C2354 VDD.t336 VSS 0.0397f
C2355 VDD.t382 VSS 0.0859f
C2356 VDD.t133 VSS 0.0705f
C2357 VDD.n300 VSS 0.0362f
C2358 VDD.t50 VSS 0.00583f
C2359 VDD.n301 VSS 0.00583f
C2360 VDD.t49 VSS 0.0769f
C2361 VDD.t64 VSS 0.0705f
C2362 VDD.n302 VSS 0.0362f
C2363 VDD.t132 VSS 0.00583f
C2364 VDD.n303 VSS 0.00583f
C2365 VDD.t131 VSS 0.0769f
C2366 VDD.t365 VSS 0.0705f
C2367 VDD.t426 VSS 0.0758f
C2368 VDD.n304 VSS 0.0362f
C2369 VDD.t427 VSS 0.00583f
C2370 VDD.t68 VSS 0.00583f
C2371 VDD.t46 VSS 0.0705f
C2372 VDD.n305 VSS 0.00583f
C2373 VDD.t460 VSS 0.0024f
C2374 VDD.n306 VSS 0.0024f
C2375 VDD.n307 VSS 0.00524f
C2376 VDD.n308 VSS 0.00583f
C2377 VDD.n309 VSS 0.0341f
C2378 VDD.t170 VSS 0.0703f
C2379 VDD.n310 VSS 0.00173f
C2380 VDD.n311 VSS 0.0012f
C2381 VDD.t488 VSS 0.00379f
C2382 VDD.t156 VSS 0.005f
C2383 VDD.n312 VSS 0.00978f
C2384 VDD.n313 VSS 0.00228f
C2385 VDD.n314 VSS 6e-19
C2386 VDD.n315 VSS 0.00534f
C2387 VDD.n316 VSS 0.00146f
C2388 VDD.n317 VSS 0.00156f
C2389 VDD.t184 VSS 0.00498f
C2390 VDD.t476 VSS 0.0038f
C2391 VDD.n318 VSS 0.0098f
C2392 VDD.n319 VSS 0.00184f
C2393 VDD.n320 VSS 6e-19
C2394 VDD.n321 VSS 0.0189f
C2395 VDD.n322 VSS 0.00165f
C2396 VDD.t482 VSS 0.00379f
C2397 VDD.n323 VSS 0.00521f
C2398 VDD.t173 VSS 0.00491f
C2399 VDD.n324 VSS 0.00466f
C2400 VDD.n325 VSS 0.0023f
C2401 VDD.n326 VSS 0.0733f
C2402 VDD.n327 VSS 0.107f
C2403 VDD.n328 VSS 0.00146f
C2404 VDD.n329 VSS 0.0015f
C2405 VDD.t152 VSS 0.00498f
C2406 VDD.t489 VSS 0.0038f
C2407 VDD.n330 VSS 0.0098f
C2408 VDD.n331 VSS 0.00191f
C2409 VDD.n332 VSS 6e-19
C2410 VDD.n333 VSS 0.0189f
C2411 VDD.t477 VSS 0.00388f
C2412 VDD.t180 VSS 0.00491f
C2413 VDD.n334 VSS 0.00978f
C2414 VDD.n335 VSS 0.00355f
C2415 VDD.n336 VSS 0.0247f
C2416 VDD.n337 VSS 0.119f
C2417 VDD.t483 VSS 0.00379f
C2418 VDD.t169 VSS 0.005f
C2419 VDD.n338 VSS 0.00977f
C2420 VDD.n339 VSS 0.0492f
C2421 VDD.n340 VSS 0.00353f
C2422 VDD.n341 VSS 0.00545f
C2423 VDD.n342 VSS 0.0152f
C2424 VDD.t140 VSS 0.0024f
C2425 VDD.n343 VSS 0.0024f
C2426 VDD.n344 VSS 0.00524f
C2427 VDD.n345 VSS 0.0333f
C2428 VDD.n346 VSS 0.0333f
C2429 VDD.n347 VSS 0.0362f
C2430 VDD.t139 VSS 0.0397f
C2431 VDD.t69 VSS 0.0859f
C2432 VDD.t261 VSS 0.0705f
C2433 VDD.t61 VSS 0.0859f
C2434 VDD.t459 VSS 0.0397f
C2435 VDD.n348 VSS 0.0362f
C2436 VDD.n349 VSS 0.018f
C2437 VDD.n350 VSS 0.0333f
C2438 VDD.n351 VSS 0.034f
C2439 VDD.t130 VSS 0.00583f
C2440 VDD.n352 VSS 0.00583f
C2441 VDD.n353 VSS 0.0268f
C2442 VDD.n354 VSS 0.0289f
C2443 VDD.n355 VSS 0.0202f
C2444 VDD.n356 VSS 0.0362f
C2445 VDD.t129 VSS 0.0769f
C2446 VDD.t221 VSS 0.0705f
C2447 VDD.t67 VSS 0.0758f
C2448 VDD.n357 VSS 0.0362f
C2449 VDD.n358 VSS 0.0202f
C2450 VDD.n359 VSS 0.0549f
C2451 VDD.n360 VSS 0.0624f
C2452 VDD.n361 VSS 0.0202f
C2453 VDD.n362 VSS 0.0268f
C2454 VDD.n363 VSS 0.0289f
C2455 VDD.n364 VSS 0.0202f
C2456 VDD.n365 VSS 0.0268f
C2457 VDD.n366 VSS 0.0289f
C2458 VDD.n367 VSS 0.0202f
C2459 VDD.n368 VSS 0.0254f
C2460 VDD.n369 VSS 0.0238f
C2461 VDD.n370 VSS 0.018f
C2462 VDD.n371 VSS 0.0276f
C2463 VDD.n372 VSS 0.0183f
C2464 VDD.t194 VSS 0.00583f
C2465 VDD.t207 VSS 0.0705f
C2466 VDD.n373 VSS 0.00583f
C2467 VDD.t347 VSS 0.0024f
C2468 VDD.n374 VSS 0.0024f
C2469 VDD.n375 VSS 0.00524f
C2470 VDD.n376 VSS 0.00583f
C2471 VDD.n377 VSS 0.0341f
C2472 VDD.t181 VSS 0.0703f
C2473 VDD.n378 VSS 0.00625f
C2474 VDD.t316 VSS 0.0024f
C2475 VDD.n379 VSS 0.0024f
C2476 VDD.n380 VSS 0.00524f
C2477 VDD.n381 VSS 0.0333f
C2478 VDD.n382 VSS 0.0449f
C2479 VDD.n383 VSS 0.0362f
C2480 VDD.t315 VSS 0.0397f
C2481 VDD.t202 VSS 0.0859f
C2482 VDD.t121 VSS 0.0705f
C2483 VDD.t285 VSS 0.0859f
C2484 VDD.t346 VSS 0.0397f
C2485 VDD.n384 VSS 0.0362f
C2486 VDD.n385 VSS 0.018f
C2487 VDD.n386 VSS 0.0333f
C2488 VDD.n387 VSS 0.034f
C2489 VDD.t320 VSS 0.00583f
C2490 VDD.n388 VSS 0.00583f
C2491 VDD.n389 VSS 0.0268f
C2492 VDD.n390 VSS 0.0289f
C2493 VDD.n391 VSS 0.0202f
C2494 VDD.n392 VSS 0.0362f
C2495 VDD.t319 VSS 0.0769f
C2496 VDD.t357 VSS 0.0705f
C2497 VDD.t193 VSS 0.0758f
C2498 VDD.n393 VSS 0.0362f
C2499 VDD.n394 VSS 0.0202f
C2500 VDD.n395 VSS 0.0516f
C2501 VDD.n396 VSS 0.0412f
C2502 VDD.n397 VSS 0.0296f
C2503 VDD.n398 VSS 0.0202f
C2504 VDD.n399 VSS 0.0268f
C2505 VDD.n400 VSS 0.0289f
C2506 VDD.n401 VSS 0.0202f
C2507 VDD.n402 VSS 0.0268f
C2508 VDD.n403 VSS 0.0289f
C2509 VDD.n404 VSS 0.0202f
C2510 VDD.n405 VSS 0.0191f
C2511 VDD.n406 VSS 0.0618f
C2512 VDD.n407 VSS 0.0734f
C2513 VDD.t201 VSS 0.00583f
C2514 VDD.n408 VSS 0.0286f
C2515 VDD.n409 VSS 0.0205f
C2516 VDD.n410 VSS 0.0362f
C2517 VDD.t200 VSS 0.0458f
C2518 VDD.n411 VSS 0.0847f
C2519 VDD.n412 VSS 0.0272f
C2520 VDD.t311 VSS 0.00583f
C2521 VDD.n413 VSS 0.0286f
C2522 VDD.n414 VSS 0.0205f
C2523 VDD.n415 VSS 0.0362f
C2524 VDD.t310 VSS 0.0458f
C2525 VDD.n416 VSS 0.0847f
C2526 VDD.n417 VSS 0.0272f
C2527 VDD.t104 VSS 0.00583f
C2528 VDD.n418 VSS 0.0286f
C2529 VDD.n419 VSS 0.0205f
C2530 VDD.n420 VSS 0.0362f
C2531 VDD.t103 VSS 0.0458f
C2532 VDD.n421 VSS 0.0538f
C2533 VDD.n422 VSS 0.0317f
C2534 VDD.n423 VSS 0.00581f
C2535 VDD.n424 VSS 0.0276f
C2536 VDD.n425 VSS 0.0192f
C2537 VDD.n426 VSS 0.0822f
C2538 VDD.t188 VSS 0.0746f
C2539 VDD.n427 VSS 0.0449f
C2540 VDD.n428 VSS 0.0584f
C2541 VDD.n429 VSS 0.0569f
C2542 VDD.n430 VSS 0.0226f
C2543 VDD.t168 VSS 0.00583f
C2544 VDD.t167 VSS 0.0542f
C2545 VDD.t197 VSS 0.0856f
C2546 VDD.n431 VSS 0.0739f
C2547 VDD.t60 VSS 0.0688f
C2548 VDD.t72 VSS 0.192f
C2549 VDD.t377 VSS 0.00609f
C2550 VDD.n432 VSS 0.00998f
C2551 VDD.n433 VSS 0.0255f
C2552 VDD.n434 VSS 0.0274f
C2553 VDD.n435 VSS 0.017f
C2554 VDD.n436 VSS 0.0262f
C2555 VDD.n437 VSS 0.0184f
C2556 VDD.n438 VSS 0.0254f
C2557 VDD.n439 VSS 0.0201f
C2558 VDD.n440 VSS 0.0289f
C2559 VDD.n441 VSS 0.0269f
C2560 VDD.n442 VSS 0.0201f
C2561 VDD.n443 VSS 0.0289f
C2562 VDD.n444 VSS 0.0269f
C2563 VDD.n445 VSS 0.0201f
C2564 VDD.n446 VSS 0.0296f
C2565 VDD.n447 VSS 0.00583f
C2566 VDD.t403 VSS 0.0759f
C2567 VDD.n448 VSS 0.0362f
C2568 VDD.t435 VSS 0.00583f
C2569 VDD.n449 VSS 0.00583f
C2570 VDD.t434 VSS 0.0703f
C2571 VDD.t274 VSS 0.077f
C2572 VDD.n450 VSS 0.0362f
C2573 VDD.t217 VSS 0.00583f
C2574 VDD.t213 VSS 0.0024f
C2575 VDD.n451 VSS 0.0024f
C2576 VDD.n452 VSS 0.00524f
C2577 VDD.t216 VSS 0.0703f
C2578 VDD.t212 VSS 0.0859f
C2579 VDD.t331 VSS 0.0399f
C2580 VDD.n453 VSS 0.0362f
C2581 VDD.t462 VSS 0.00583f
C2582 VDD.t420 VSS 0.0024f
C2583 VDD.n454 VSS 0.0024f
C2584 VDD.n455 VSS 0.00524f
C2585 VDD.t461 VSS 0.0703f
C2586 VDD.t419 VSS 0.0859f
C2587 VDD.t452 VSS 0.0399f
C2588 VDD.t164 VSS 0.0701f
C2589 VDD.n456 VSS 0.0362f
C2590 VDD.t165 VSS 0.00625f
C2591 VDD.n457 VSS 0.0449f
C2592 VDD.n458 VSS 0.0332f
C2593 VDD.n459 VSS 0.0341f
C2594 VDD.n460 VSS 0.0181f
C2595 VDD.n461 VSS 0.0332f
C2596 VDD.n462 VSS 0.034f
C2597 VDD.n463 VSS 0.0201f
C2598 VDD.n464 VSS 0.0289f
C2599 VDD.n465 VSS 0.0269f
C2600 VDD.n466 VSS 0.0201f
C2601 VDD.n467 VSS 0.0517f
C2602 VDD.n468 VSS 0.0367f
C2603 VDD.n469 VSS 0.0179f
C2604 VDD.n470 VSS 0.0275f
C2605 VDD.n471 VSS 0.0181f
C2606 VDD.n472 VSS 0.0238f
C2607 VDD.n473 VSS 0.0254f
C2608 VDD.n474 VSS 0.0201f
C2609 VDD.n475 VSS 0.0289f
C2610 VDD.n476 VSS 0.0269f
C2611 VDD.n477 VSS 0.0201f
C2612 VDD.n478 VSS 0.0289f
C2613 VDD.n479 VSS 0.0269f
C2614 VDD.n480 VSS 0.0201f
C2615 VDD.n481 VSS 0.0296f
C2616 VDD.n482 VSS 0.00583f
C2617 VDD.t20 VSS 0.0759f
C2618 VDD.n483 VSS 0.0362f
C2619 VDD.t227 VSS 0.00583f
C2620 VDD.n484 VSS 0.00583f
C2621 VDD.t226 VSS 0.0703f
C2622 VDD.t241 VSS 0.077f
C2623 VDD.n485 VSS 0.0362f
C2624 VDD.t354 VSS 0.00583f
C2625 VDD.t88 VSS 0.0024f
C2626 VDD.n486 VSS 0.0024f
C2627 VDD.n487 VSS 0.00524f
C2628 VDD.t353 VSS 0.0703f
C2629 VDD.t87 VSS 0.0859f
C2630 VDD.t390 VSS 0.0399f
C2631 VDD.n488 VSS 0.0362f
C2632 VDD.t248 VSS 0.00583f
C2633 VDD.t24 VSS 0.0024f
C2634 VDD.n489 VSS 0.0024f
C2635 VDD.n490 VSS 0.00524f
C2636 VDD.t247 VSS 0.0703f
C2637 VDD.t23 VSS 0.0859f
C2638 VDD.t409 VSS 0.0399f
C2639 VDD.t178 VSS 0.0701f
C2640 VDD.n491 VSS 0.0362f
C2641 VDD.t179 VSS 0.00625f
C2642 VDD.n492 VSS 0.0449f
C2643 VDD.n493 VSS 0.0332f
C2644 VDD.n494 VSS 0.0341f
C2645 VDD.n495 VSS 0.0181f
C2646 VDD.n496 VSS 0.0332f
C2647 VDD.n497 VSS 0.034f
C2648 VDD.n498 VSS 0.0201f
C2649 VDD.n499 VSS 0.0289f
C2650 VDD.n500 VSS 0.0269f
C2651 VDD.n501 VSS 0.0201f
C2652 VDD.n502 VSS 0.0517f
C2653 VDD.n503 VSS 0.0413f
C2654 VDD.n504 VSS 0.0183f
C2655 VDD.n505 VSS 0.0275f
C2656 VDD.n506 VSS 0.0181f
C2657 VDD.n507 VSS 0.0238f
C2658 CLK_div_10_mag_1.Q1.n0 VSS 0.196f
C2659 CLK_div_10_mag_1.Q1.n1 VSS 0.191f
C2660 CLK_div_10_mag_1.Q1.n2 VSS 0.00491f
C2661 CLK_div_10_mag_1.Q1.n3 VSS 0.0761f
C2662 CLK_div_10_mag_1.Q1.n4 VSS 0.0132f
C2663 CLK_div_10_mag_1.Q1.n5 VSS 0.119f
C2664 CLK_div_10_mag_1.Q1.n6 VSS 0.0879f
C2665 CLK_div_10_mag_1.Q1.n7 VSS 0.0167f
C2666 CLK_div_10_mag_1.Q1.n8 VSS 0.0244f
C2667 CLK_div_10_mag_1.Q1.t2 VSS 0.0233f
C2668 CLK_div_10_mag_1.Q1.t0 VSS 0.0192f
C2669 CLK_div_10_mag_1.Q1.n9 VSS 0.0192f
C2670 CLK_div_10_mag_1.Q1.n10 VSS 0.0462f
C2671 CLK_div_10_mag_1.Q1.n11 VSS 0.144f
C2672 CLK_div_10_mag_1.Q1.t5 VSS 0.0428f
C2673 CLK_div_10_mag_1.Q1.t16 VSS 0.0282f
C2674 CLK_div_10_mag_1.Q1.n12 VSS 0.076f
C2675 CLK_div_10_mag_1.Q1.n13 VSS 0.298f
C2676 CLK_div_10_mag_1.Q1.t3 VSS 0.0307f
C2677 CLK_div_10_mag_1.Q1.t14 VSS 0.0246f
C2678 CLK_div_10_mag_1.Q1.n14 VSS 0.0713f
C2679 CLK_div_10_mag_1.Q1.n15 VSS 0.0442f
C2680 CLK_div_10_mag_1.Q1.n16 VSS 0.567f
C2681 CLK_div_10_mag_1.Q1.t4 VSS 0.0428f
C2682 CLK_div_10_mag_1.Q1.t15 VSS 0.0282f
C2683 CLK_div_10_mag_1.Q1.n17 VSS 0.0756f
C2684 CLK_div_10_mag_1.Q1.t8 VSS 0.0428f
C2685 CLK_div_10_mag_1.Q1.t7 VSS 0.0282f
C2686 CLK_div_10_mag_1.Q1.n18 VSS 0.0757f
C2687 CLK_div_10_mag_1.Q1.t9 VSS 0.0307f
C2688 CLK_div_10_mag_1.Q1.t12 VSS 0.0246f
C2689 CLK_div_10_mag_1.Q1.n19 VSS 0.0695f
C2690 CLK_div_10_mag_1.Q1.t10 VSS 0.0219f
C2691 CLK_div_10_mag_1.Q1.t13 VSS 0.0401f
C2692 CLK_div_10_mag_1.Q1.n20 VSS 0.0755f
C2693 CLK_div_10_mag_1.Q1.n21 VSS 0.66f
C2694 CLK_div_10_mag_1.Q1.t11 VSS 0.0353f
C2695 CLK_div_10_mag_1.Q1.t6 VSS 0.00913f
C2696 CLK_div_10_mag_1.Q1.n22 VSS 0.0585f
C2697 CLK_div_10_mag_1.Q1.n23 VSS 0.0619f
C2698 CLK_div_10_mag_1.Q1.n24 VSS 0.144f
C2699 CLK_div_10_mag_1.Q1.n25 VSS 0.0182f
.ends

