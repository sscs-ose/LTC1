magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -4254 -2045 4254 2045
<< ndiff >>
rect -2254 23 2254 45
rect -2254 -23 -2232 23
rect 2232 -23 2254 23
rect -2254 -45 2254 -23
<< ndiffc >>
rect -2232 -23 2232 23
<< metal1 >>
rect -2243 23 2243 34
rect -2243 -23 -2232 23
rect 2232 -23 2243 23
rect -2243 -34 2243 -23
<< end >>
