magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2445 -8095 2445 8095
<< psubdiff >>
rect -445 6073 445 6095
rect -445 -6073 -423 6073
rect 423 -6073 445 6073
rect -445 -6095 445 -6073
<< psubdiffcont >>
rect -423 -6073 423 6073
<< metal1 >>
rect -434 6073 434 6084
rect -434 -6073 -423 6073
rect 423 -6073 434 6073
rect -434 -6084 434 -6073
<< end >>
