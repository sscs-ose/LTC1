* NGSPICE file created from nmos_3p3_GGGST2_flat.ext - technology: gf180mcuC

.subckt nmos_3p3_GGGST2_flat OUT VDD VSS A B
X0 VDD A.t0 a_86_440.t1 VDD.t3 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X1 VDD a_390_68.t4 OUT.t0 VDD.t7 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X2 OUT a_390_68.t5 VSS.t6 VSS.t5 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X3 VSS B.t2 a_390_68.t1 VSS.t2 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
R0 A.n0 A.t0 36.5005
R1 A.n2 A.n1 18.2505
R2 A.n1 A.t1 16.0344
R3 A.n0 A.t2 15.6434
R4 A.n1 A.n0 8.73443
R5 A A.n2 8.0005
R6 A A.n2 8.0005
R7 a_86_440.n2 a_86_440.t1 5.61007
R8 a_86_440.n3 a_86_440.n2 5.61007
R9 a_86_440.n2 a_86_440.n1 2.6005
R10 a_86_440.n1 a_86_440.t3 1.8205
R11 a_86_440.n1 a_86_440.n0 1.8205
R12 VDD.n11 VDD.t0 82.9108
R13 VDD.n19 VDD.t3 77.8347
R14 VDD.n2 VDD.t7 75.7026
R15 VDD.n23 VDD.t1 33.8415
R16 VDD.n29 VDD.t6 13.5369
R17 VDD.n1 VDD.n0 4.88224
R18 VDD.n4 VDD.n3 3.1505
R19 VDD.n7 VDD.n6 3.1505
R20 VDD.n6 VDD.n5 3.1505
R21 VDD.n10 VDD.n9 3.1505
R22 VDD.n9 VDD.n8 3.1505
R23 VDD.n13 VDD.n12 3.1505
R24 VDD.n12 VDD.n11 3.1505
R25 VDD.n16 VDD.n15 3.1505
R26 VDD.n15 VDD.n14 3.1505
R27 VDD.n31 VDD.n30 3.1505
R28 VDD.n30 VDD.n29 3.1505
R29 VDD.n28 VDD.n27 3.1505
R30 VDD.n27 VDD.n26 3.1505
R31 VDD.n25 VDD.n24 3.1505
R32 VDD.n24 VDD.n23 3.1505
R33 VDD.n20 VDD.n19 3.1505
R34 VDD.n22 VDD.n18 3.06224
R35 VDD.n21 VDD.n20 1.87197
R36 VDD.n18 VDD.t2 1.8205
R37 VDD.n18 VDD.n17 1.8205
R38 VDD.n22 VDD.n21 0.593718
R39 VDD.n3 VDD.n2 0.150506
R40 VDD.n16 VDD.n13 0.0864821
R41 VDD.n7 VDD.n4 0.0760357
R42 VDD.n10 VDD.n7 0.0760357
R43 VDD.n13 VDD.n10 0.0760357
R44 VDD.n31 VDD.n28 0.0760357
R45 VDD.n28 VDD.n25 0.0760357
R46 VDD.n25 VDD.n22 0.0487143
R47 VDD VDD.n16 0.0382679
R48 VDD VDD.n31 0.0382679
R49 VDD.n4 VDD.n1 0.0302321
R50 B.n1 B.t2 63.6148
R51 B.n0 B.t0 36.5005
R52 B.t2 B.n0 32.0684
R53 B.n0 B.t1 15.6434
R54 B B.n1 8.0005
R55 B B.n1 8.0005
R56 a_390_68.n0 a_390_68.t4 68.3076
R57 a_390_68.n0 a_390_68.t5 15.2404
R58 a_390_68.n3 a_390_68.n0 4.04418
R59 a_390_68.n3 a_390_68.n2 3.62789
R60 a_390_68.n2 a_390_68.t1 3.2765
R61 a_390_68.n2 a_390_68.n1 3.2765
R62 a_390_68.n5 a_390_68.n3 3.1718
R63 a_390_68.t3 a_390_68.n5 1.8205
R64 a_390_68.n5 a_390_68.n4 1.8205
R65 OUT.n1 OUT.n0 6.93911
R66 OUT.n1 OUT.t0 4.80398
R67 OUT OUT.n1 0.340935
R68 VSS.n6 VSS.t2 277.728
R69 VSS.n2 VSS.t5 112.273
R70 VSS.n11 VSS.t0 112.273
R71 VSS.n10 VSS.t1 6.91182
R72 VSS.n5 VSS.n1 3.6318
R73 VSS.n1 VSS.t6 3.2765
R74 VSS.n1 VSS.n0 3.2765
R75 VSS.n10 VSS.n9 2.6005
R76 VSS.n3 VSS.n2 2.6005
R77 VSS.n8 VSS.n7 2.6005
R78 VSS.n7 VSS.n6 2.6005
R79 VSS.n16 VSS.n15 2.6005
R80 VSS.n15 VSS.n14 2.6005
R81 VSS.n13 VSS.n12 2.6005
R82 VSS.n12 VSS.n11 2.6005
R83 VSS.n4 VSS.n3 1.64943
R84 VSS.n5 VSS.n4 0.532617
R85 VSS.n16 VSS.n13 0.0760357
R86 VSS.n13 VSS.n10 0.0760357
R87 VSS VSS.n16 0.0446964
R88 VSS VSS.n8 0.0318393
R89 VSS.n8 VSS.n5 0.0270179
C0 B VDD 0.204f
C1 OUT VDD 0.177f
C2 B OUT 0.00407f
C3 A VDD 0.234f
C4 A B 0.0839f
.ends

