* NGSPICE file created from JK_FF_mag_flat.ext - technology: gf180mcuC

.subckt pex_JK_FF_mag CLK VSS VDD Q J QB RST K
X0 nand2_mag_3.IN1 CLK.t0 VSS.t23 VSS.t22 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1 nand3_mag_1.IN1 nand3_mag_1.OUT a_968_1353# VSS.t12 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2 nand2_mag_4.IN2 nand3_mag_1.OUT VDD.t20 VDD.t19 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X3 a_398_212# CLK.t1 a_238_212# VSS.t21 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X4 a_1532_1353# nand3_mag_1.IN1 VSS.t15 VSS.t14 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X5 Q QB.t3 a_2096_1353# VSS.t9 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X6 a_968_1353# nand3_mag_0.OUT VSS.t1 VSS.t0 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X7 Q nand2_mag_1.IN2 VDD.t45 VDD.t44 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X8 VDD RST.t0 nand3_mag_1.OUT VDD.t4 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X9 QB Q.t3 a_2250_256# VSS.t6 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X10 nand3_mag_0.OUT J.t0 VDD.t13 VDD.t12 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X11 VDD nand2_mag_3.IN1 nand2_mag_4.IN2 VDD.t28 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X12 a_1122_212# RST.t1 a_962_212# VSS.t4 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X13 a_1686_256# nand3_mag_1.OUT VSS.t11 VSS.t10 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X14 a_2096_1353# nand2_mag_1.IN2 VSS.t25 VSS.t24 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X15 nand3_mag_2.OUT Q.t4 VDD.t11 VDD.t10 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X16 nand3_mag_0.OUT QB.t4 a_404_1309# VSS.t26 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X17 nand2_mag_4.IN2 nand2_mag_3.IN1 a_1686_256# VSS.t17 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X18 QB nand2_mag_4.IN2 VDD.t3 VDD.t2 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X19 nand3_mag_2.OUT Q.t5 a_398_212# VSS.t5 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X20 nand3_mag_2.OUT K.t0 VDD.t40 VDD.t39 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X21 VDD nand2_mag_3.IN1 nand2_mag_1.IN2 VDD.t25 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X22 nand3_mag_1.OUT nand3_mag_1.IN1 VDD.t24 VDD.t23 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X23 a_238_212# K.t1 VSS.t8 VSS.t7 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X24 nand3_mag_0.OUT QB.t5 VDD.t15 VDD.t14 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X25 nand3_mag_1.OUT nand3_mag_1.IN1 a_1122_212# VSS.t13 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X26 a_2250_256# nand2_mag_4.IN2 VSS.t3 VSS.t2 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X27 nand2_mag_3.IN1 CLK.t2 VDD.t38 VDD.t37 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X28 a_404_1309# CLK.t3 a_244_1309# VSS.t20 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X29 nand2_mag_1.IN2 nand2_mag_3.IN1 a_1532_1353# VSS.t16 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X30 VDD nand3_mag_1.OUT nand3_mag_1.IN1 VDD.t16 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X31 nand2_mag_1.IN2 nand3_mag_1.IN1 VDD.t22 VDD.t21 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X32 VDD QB.t6 Q.t0 VDD.t41 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X33 nand3_mag_1.IN1 nand3_mag_0.OUT VDD.t1 VDD.t0 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X34 nand3_mag_1.OUT nand3_mag_2.OUT VDD.t47 VDD.t46 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X35 VDD Q.t6 QB.t1 VDD.t7 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X36 VDD CLK.t4 nand3_mag_0.OUT VDD.t34 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X37 VDD CLK.t5 nand3_mag_2.OUT VDD.t31 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X38 a_962_212# nand3_mag_2.OUT VSS.t28 VSS.t27 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X39 a_244_1309# J.t1 VSS.t19 VSS.t18 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
R0 CLK.n9 CLK.t3 36.935
R1 CLK.n3 CLK.t1 36.935
R2 CLK.n14 CLK.t2 25.5361
R3 CLK.n9 CLK.t4 18.1962
R4 CLK.n3 CLK.t5 18.1962
R5 CLK.n14 CLK.t0 14.0734
R6 CLK.n5 CLK.n2 4.5005
R7 CLK.n5 CLK.n4 4.5005
R8 CLK.n8 CLK.n7 4.5005
R9 CLK.n10 CLK.n7 4.5005
R10 CLK.n16 CLK.n15 4.5005
R11 CLK.n17 CLK.n16 4.5005
R12 CLK.n12 CLK.n11 2.25107
R13 CLK.n13 CLK.n0 2.24235
R14 CLK.n4 CLK.n3 2.12175
R15 CLK.n10 CLK.n9 2.12075
R16 CLK.n7 CLK.n6 1.74297
R17 CLK.n6 CLK.n1 1.49778
R18 CLK.n15 CLK.n14 1.42775
R19 CLK.n13 CLK.n12 0.97145
R20 CLK CLK.n17 0.1605
R21 CLK.n8 CLK 0.0473512
R22 CLK.n2 CLK 0.0473512
R23 CLK.n11 CLK.n8 0.0361897
R24 CLK.n2 CLK.n1 0.0361897
R25 CLK.n17 CLK.n0 0.03175
R26 CLK.n16 CLK.n13 0.0246174
R27 CLK.n6 CLK.n5 0.0131772
R28 CLK.n12 CLK.n7 0.0122182
R29 CLK.n11 CLK.n10 0.00515517
R30 CLK.n4 CLK.n1 0.00515517
R31 CLK.n15 CLK.n0 0.00175
R32 VSS.t7 VSS.n21 6810.9
R33 VSS.t17 VSS.t2 2510.52
R34 VSS.t5 VSS.t27 2510.52
R35 VSS.t16 VSS.t24 2307.56
R36 VSS.t14 VSS.t12 2307.56
R37 VSS.t26 VSS.t0 2307.56
R38 VSS.t22 VSS.t18 2307.56
R39 VSS.t4 VSS.t13 994.264
R40 VSS.t21 VSS.t5 994.264
R41 VSS.t20 VSS.t26 913.885
R42 VSS.n4 VSS.t6 596.558
R43 VSS.n5 VSS.t17 596.558
R44 VSS.n9 VSS.t4 596.558
R45 VSS.n22 VSS.t21 596.558
R46 VSS.n12 VSS.t9 548.331
R47 VSS.n13 VSS.t16 548.331
R48 VSS.n18 VSS.t12 548.331
R49 VSS.n19 VSS.t20 548.331
R50 VSS.t2 VSS.n4 397.707
R51 VSS.n5 VSS.t10 397.707
R52 VSS.t27 VSS.n9 397.707
R53 VSS.n22 VSS.t7 397.707
R54 VSS.t24 VSS.n12 365.555
R55 VSS.n13 VSS.t14 365.555
R56 VSS.t0 VSS.n18 365.555
R57 VSS.t18 VSS.n19 365.555
R58 VSS.n21 VSS.t22 22.8476
R59 VSS.n21 VSS.n20 16.6241
R60 VSS.n20 VSS.t23 9.3736
R61 VSS.n2 VSS.t3 7.19156
R62 VSS.n7 VSS.t11 7.19156
R63 VSS.n10 VSS.t25 7.19156
R64 VSS.n15 VSS.t15 7.19156
R65 VSS.n16 VSS.t1 7.19156
R66 VSS.n1 VSS.t28 5.91399
R67 VSS.n24 VSS.t8 5.91399
R68 VSS.n26 VSS.t19 5.91399
R69 VSS.n23 VSS.n22 5.2005
R70 VSS.n9 VSS.n8 5.2005
R71 VSS.n6 VSS.n5 5.2005
R72 VSS.n4 VSS.n3 5.2005
R73 VSS.n19 VSS.n0 5.2005
R74 VSS.n18 VSS.n17 5.2005
R75 VSS.n14 VSS.n13 5.2005
R76 VSS.n12 VSS.n11 5.2005
R77 VSS.n25 VSS.n24 1.03335
R78 VSS.n8 VSS.n7 0.480225
R79 VSS.n23 VSS.n1 0.480225
R80 VSS.n2 VSS 0.343161
R81 VSS.n10 VSS 0.343161
R82 VSS VSS.n15 0.343161
R83 VSS VSS.n0 0.289491
R84 VSS.n16 VSS 0.191234
R85 VSS.n25 VSS 0.137685
R86 VSS.n3 VSS.n2 0.118573
R87 VSS.n7 VSS.n6 0.118573
R88 VSS.n11 VSS.n10 0.118573
R89 VSS.n15 VSS.n14 0.118573
R90 VSS.n17 VSS.n16 0.118573
R91 VSS VSS.n1 0.115271
R92 VSS.n24 VSS 0.115271
R93 VSS VSS.n26 0.115271
R94 VSS.n26 VSS.n25 0.10206
R95 VSS.n3 VSS 0.00545413
R96 VSS.n6 VSS 0.00545413
R97 VSS.n11 VSS 0.00545413
R98 VSS.n14 VSS 0.00545413
R99 VSS.n17 VSS 0.00545413
R100 VSS.n8 VSS 0.00380275
R101 VSS VSS.n23 0.00380275
R102 VSS VSS.n0 0.00380275
R103 VSS.n20 VSS 0.00219811
R104 VDD.t16 VDD.t21 765.152
R105 VDD.t14 VDD.t0 765.152
R106 VDD.t28 VDD.t2 765.152
R107 VDD.t23 VDD.t19 765.152
R108 VDD.t10 VDD.t46 765.152
R109 VDD VDD.n32 429.187
R110 VDD.n32 VDD.t12 386.365
R111 VDD.t34 VDD.t14 303.031
R112 VDD.t4 VDD.t23 303.031
R113 VDD.t31 VDD.t10 303.031
R114 VDD.n23 VDD.t41 193.183
R115 VDD.n26 VDD.t25 193.183
R116 VDD.n28 VDD.t16 193.183
R117 VDD.n31 VDD.t34 193.183
R118 VDD.n2 VDD.t7 193.183
R119 VDD.n4 VDD.t28 193.183
R120 VDD.n7 VDD.t4 193.183
R121 VDD.n10 VDD.t31 193.183
R122 VDD.n23 VDD.t44 109.849
R123 VDD.t21 VDD.n26 109.849
R124 VDD.t0 VDD.n28 109.849
R125 VDD.t12 VDD.n31 109.849
R126 VDD.t2 VDD.n2 109.849
R127 VDD.t19 VDD.n4 109.849
R128 VDD.t46 VDD.n7 109.849
R129 VDD.n10 VDD.t39 109.849
R130 VDD.n32 VDD.t37 59.702
R131 VDD.n11 VDD.n10 6.3005
R132 VDD.n14 VDD.n7 6.3005
R133 VDD.n17 VDD.n4 6.3005
R134 VDD.n20 VDD.n2 6.3005
R135 VDD.n24 VDD.n23 6.3005
R136 VDD.n40 VDD.n26 6.3005
R137 VDD.n37 VDD.n28 6.3005
R138 VDD.n34 VDD.n31 6.3005
R139 VDD.n11 VDD.t40 5.213
R140 VDD VDD.t38 5.16454
R141 VDD.n33 VDD.t13 5.13287
R142 VDD.n36 VDD.t1 5.13287
R143 VDD.n38 VDD.n27 5.13287
R144 VDD.n39 VDD.t22 5.13287
R145 VDD.n41 VDD.n25 5.13287
R146 VDD.n42 VDD.t45 5.13287
R147 VDD.n22 VDD.n0 5.13287
R148 VDD.n13 VDD.t47 5.13287
R149 VDD.n16 VDD.t20 5.13287
R150 VDD.n18 VDD.n3 5.13287
R151 VDD.n19 VDD.t3 5.13287
R152 VDD.n21 VDD.n1 5.13287
R153 VDD.n35 VDD.n30 2.85787
R154 VDD.n12 VDD.n9 2.85787
R155 VDD.n15 VDD.n6 2.85787
R156 VDD.n30 VDD.t15 2.2755
R157 VDD.n30 VDD.n29 2.2755
R158 VDD.n9 VDD.t11 2.2755
R159 VDD.n9 VDD.n8 2.2755
R160 VDD.n6 VDD.t24 2.2755
R161 VDD.n6 VDD.n5 2.2755
R162 VDD.n33 VDD 1.77285
R163 VDD.n22 VDD.n21 1.16167
R164 VDD.n16 VDD.n15 0.233919
R165 VDD.n13 VDD.n12 0.233919
R166 VDD.n19 VDD.n18 0.141016
R167 VDD.n42 VDD.n41 0.141016
R168 VDD.n39 VDD.n38 0.141016
R169 VDD.n36 VDD 0.122435
R170 VDD VDD.n35 0.111984
R171 VDD.n21 VDD.n20 0.107339
R172 VDD.n18 VDD.n17 0.107339
R173 VDD.n24 VDD.n22 0.107339
R174 VDD.n41 VDD.n40 0.107339
R175 VDD.n38 VDD.n37 0.107339
R176 VDD.n15 VDD 0.106177
R177 VDD.n12 VDD 0.106177
R178 VDD.n35 VDD 0.106177
R179 VDD.n14 VDD.n13 0.080629
R180 VDD.n34 VDD.n33 0.080629
R181 VDD VDD.n19 0.0794677
R182 VDD VDD.n16 0.0794677
R183 VDD VDD.n42 0.0794677
R184 VDD VDD.n39 0.0794677
R185 VDD VDD.n36 0.0794677
R186 VDD.n20 VDD 0.00166129
R187 VDD.n17 VDD 0.00166129
R188 VDD VDD.n14 0.00166129
R189 VDD VDD.n11 0.00166129
R190 VDD VDD.n24 0.00166129
R191 VDD.n40 VDD 0.00166129
R192 VDD.n37 VDD 0.00166129
R193 VDD VDD.n34 0.00166129
R194 QB.n3 QB.t4 37.1981
R195 QB.n1 QB.t3 31.528
R196 QB.n3 QB.t5 17.6611
R197 QB.n1 QB.t6 15.3826
R198 QB.n2 QB.n1 7.62751
R199 QB.n9 QB.n0 7.11377
R200 QB.n5 QB.n4 6.09789
R201 QB.n8 QB.n7 2.99416
R202 QB.n5 QB.n2 2.67866
R203 QB.n7 QB.t1 2.2755
R204 QB.n7 QB.n6 2.2755
R205 QB.n8 QB.n5 2.2505
R206 QB.n4 QB.n3 1.43706
R207 QB.n9 QB.n8 0.241045
R208 QB.n2 QB 0.144374
R209 QB.n4 QB 0.0670696
R210 QB QB.n9 0.0414091
R211 Q.n0 Q.t5 36.935
R212 Q.n2 Q.t3 31.528
R213 Q.n0 Q.t4 18.1962
R214 Q.n2 Q.t6 15.3826
R215 Q.n8 Q.n5 7.09905
R216 Q.n3 Q.n2 6.86134
R217 Q.n4 Q.n1 5.01116
R218 Q.n9 Q.n4 3.7789
R219 Q.n8 Q.n7 3.25085
R220 Q.n7 Q.t0 2.2755
R221 Q.n7 Q.n6 2.2755
R222 Q.n1 Q.n0 2.13398
R223 Q.n4 Q.n3 1.12056
R224 Q.n9 Q.n8 0.0919062
R225 Q.n3 Q 0.0857632
R226 Q.n1 Q 0.0810725
R227 Q Q.n9 0.073625
R228 RST.n0 RST.t1 36.935
R229 RST.n0 RST.t0 18.1962
R230 RST RST.n0 4.08138
R231 J.n0 J.t0 30.9379
R232 J.n0 J.t1 24.5101
R233 J J.n0 4.11094
R234 K.n0 K.t0 30.9379
R235 K.n0 K.t1 24.5101
R236 K K.n0 4.11094
C0 nand2_mag_3.IN1 Q 0.0168f
C1 a_968_1353# nand3_mag_1.IN1 0.0697f
C2 CLK nand3_mag_0.OUT 0.268f
C3 a_2096_1353# nand2_mag_3.IN1 0.00118f
C4 nand3_mag_2.OUT Q 0.338f
C5 K nand3_mag_2.OUT 0.0904f
C6 nand2_mag_3.IN1 J 0.0393f
C7 VDD CLK 0.695f
C8 a_1122_212# nand3_mag_1.IN1 8.64e-19
C9 a_238_212# Q 0.00335f
C10 RST nand3_mag_1.IN1 0.123f
C11 nand2_mag_3.IN1 nand3_mag_1.OUT 0.16f
C12 a_2250_256# Q 0.0157f
C13 K a_238_212# 8.64e-19
C14 a_398_212# nand2_mag_3.IN1 1.46e-19
C15 nand3_mag_2.OUT nand3_mag_1.OUT 0.121f
C16 nand2_mag_4.IN2 nand2_mag_1.IN2 8.16e-20
C17 a_404_1309# Q 2.79e-20
C18 a_1686_256# Q 0.00859f
C19 a_238_212# nand3_mag_1.OUT 1.17e-20
C20 QB nand2_mag_1.IN2 0.0592f
C21 a_1122_212# Q 0.0101f
C22 a_398_212# nand3_mag_2.OUT 0.0731f
C23 RST Q 0.00332f
C24 nand2_mag_4.IN2 QB 0.199f
C25 a_968_1353# nand3_mag_1.OUT 0.0202f
C26 a_398_212# a_238_212# 0.0504f
C27 a_1532_1353# nand2_mag_1.IN2 0.069f
C28 a_1686_256# nand3_mag_1.OUT 0.00378f
C29 QB nand3_mag_0.OUT 0.343f
C30 VDD nand2_mag_1.IN2 0.397f
C31 a_1122_212# nand3_mag_1.OUT 0.0733f
C32 RST nand3_mag_1.OUT 0.216f
C33 a_1532_1353# QB 2.96e-19
C34 a_404_1309# a_244_1309# 0.0504f
C35 VDD nand2_mag_4.IN2 0.391f
C36 VDD QB 0.909f
C37 nand3_mag_2.OUT nand2_mag_3.IN1 0.00119f
C38 VDD nand3_mag_0.OUT 0.647f
C39 a_962_212# Q 0.0102f
C40 VDD a_1532_1353# 3.14e-19
C41 CLK nand3_mag_1.IN1 9.71e-20
C42 a_968_1353# nand2_mag_3.IN1 1.43e-19
C43 a_238_212# nand3_mag_2.OUT 0.0202f
C44 a_404_1309# nand2_mag_3.IN1 0.00119f
C45 a_962_212# nand3_mag_1.OUT 0.0203f
C46 a_1686_256# nand2_mag_3.IN1 0.0036f
C47 RST nand2_mag_3.IN1 1.35e-20
C48 CLK Q 0.149f
C49 K CLK 0.0518f
C50 a_1122_212# nand3_mag_2.OUT 2.88e-20
C51 RST nand3_mag_2.OUT 0.0475f
C52 CLK J 0.0832f
C53 nand3_mag_1.IN1 nand2_mag_1.IN2 0.109f
C54 CLK nand3_mag_1.OUT 6.64e-19
C55 nand3_mag_1.IN1 QB 0.0445f
C56 CLK a_244_1309# 0.0101f
C57 a_398_212# CLK 0.00164f
C58 nand3_mag_1.IN1 nand3_mag_0.OUT 0.122f
C59 a_1122_212# RST 0.00103f
C60 Q nand2_mag_1.IN2 0.107f
C61 a_1532_1353# nand3_mag_1.IN1 0.0059f
C62 a_962_212# nand3_mag_2.OUT 9.1e-19
C63 nand2_mag_4.IN2 Q 0.0635f
C64 VDD nand3_mag_1.IN1 0.653f
C65 a_2096_1353# nand2_mag_1.IN2 0.00372f
C66 QB Q 1.94f
C67 a_2096_1353# nand2_mag_4.IN2 4.52e-20
C68 nand2_mag_1.IN2 nand3_mag_1.OUT 0.00975f
C69 Q nand3_mag_0.OUT 7.24e-19
C70 a_2096_1353# QB 0.0114f
C71 CLK nand2_mag_3.IN1 0.408f
C72 nand2_mag_4.IN2 nand3_mag_1.OUT 0.122f
C73 QB J 1.3e-19
C74 QB nand3_mag_1.OUT 0.254f
C75 VDD Q 0.858f
C76 a_1122_212# a_962_212# 0.0504f
C77 CLK nand3_mag_2.OUT 0.235f
C78 nand3_mag_0.OUT J 0.0904f
C79 RST a_962_212# 8.64e-19
C80 VDD K 0.158f
C81 nand3_mag_1.OUT nand3_mag_0.OUT 0.0622f
C82 a_238_212# CLK 0.00117f
C83 VDD a_2096_1353# 3.56e-19
C84 a_1532_1353# nand3_mag_1.OUT 4.52e-20
C85 VDD J 0.168f
C86 CLK a_968_1353# 6.43e-21
C87 a_244_1309# nand3_mag_0.OUT 0.0203f
C88 VDD nand3_mag_1.OUT 0.994f
C89 CLK a_404_1309# 0.00939f
C90 VDD a_244_1309# 2.21e-19
C91 nand2_mag_3.IN1 nand2_mag_1.IN2 0.36f
C92 nand2_mag_4.IN2 nand2_mag_3.IN1 0.321f
C93 nand2_mag_3.IN1 QB 0.281f
C94 nand2_mag_3.IN1 nand3_mag_0.OUT 0.0894f
C95 nand3_mag_2.OUT QB 0.103f
C96 a_1532_1353# nand2_mag_3.IN1 0.011f
C97 a_2250_256# nand2_mag_4.IN2 0.00372f
C98 nand3_mag_2.OUT nand3_mag_0.OUT 0.00183f
C99 VDD nand2_mag_3.IN1 1.14f
C100 a_2250_256# QB 0.0811f
C101 nand3_mag_1.IN1 Q 0.00335f
C102 a_968_1353# QB 3.33e-19
C103 a_1686_256# nand2_mag_4.IN2 0.069f
C104 VDD nand3_mag_2.OUT 0.642f
C105 a_404_1309# QB 0.00392f
C106 a_968_1353# nand3_mag_0.OUT 0.00378f
C107 a_1686_256# QB 0.00964f
C108 VDD a_238_212# 2.21e-19
C109 a_2250_256# VDD 3.14e-19
C110 a_404_1309# nand3_mag_0.OUT 0.0732f
C111 a_1122_212# QB 0.00696f
C112 RST QB 0.0121f
C113 nand3_mag_1.IN1 nand3_mag_1.OUT 0.769f
C114 VDD a_968_1353# 3.14e-19
C115 K Q 0.00438f
C116 a_1686_256# VDD 3.14e-19
C117 a_2096_1353# Q 0.069f
C118 VDD RST 0.171f
C119 Q nand3_mag_1.OUT 0.0343f
C120 K J 0.00197f
C121 a_962_212# QB 0.00695f
C122 a_398_212# Q 0.00789f
C123 nand2_mag_3.IN1 nand3_mag_1.IN1 0.233f
C124 a_244_1309# J 8.64e-19
C125 CLK nand2_mag_1.IN2 1.48e-20
C126 a_398_212# nand3_mag_1.OUT 1.5e-20
C127 VDD a_962_212# 2.21e-19
C128 nand3_mag_2.OUT nand3_mag_1.IN1 0.00224f
C129 CLK QB 0.307f
C130 a_2250_256# VSS 0.0675f
C131 a_1686_256# VSS 0.0676f
C132 a_1122_212# VSS 0.0343f
C133 a_962_212# VSS 0.0881f
C134 a_398_212# VSS 0.0343f
C135 a_238_212# VSS 0.0881f
C136 nand2_mag_4.IN2 VSS 0.415f
C137 RST VSS 0.19f
C138 nand3_mag_2.OUT VSS 0.539f
C139 K VSS 0.33f
C140 a_2096_1353# VSS 0.0676f
C141 a_1532_1353# VSS 0.0676f
C142 a_968_1353# VSS 0.0676f
C143 a_404_1309# VSS 0.0343f
C144 a_244_1309# VSS 0.0881f
C145 Q VSS 1.4f
C146 nand2_mag_1.IN2 VSS 0.415f
C147 nand2_mag_3.IN1 VSS 0.963f
C148 nand3_mag_1.IN1 VSS 0.724f
C149 nand3_mag_1.OUT VSS 0.809f
C150 nand3_mag_0.OUT VSS 0.509f
C151 QB VSS 0.92f
C152 J VSS 0.275f
C153 CLK VSS 1.01f
C154 VDD VSS 12.4f
.ends

