magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1073 -7310 1073 7310
<< metal1 >>
rect -73 6304 73 6310
rect -73 6278 -67 6304
rect -41 6278 -13 6304
rect 13 6278 41 6304
rect 67 6278 73 6304
rect -73 6250 73 6278
rect -73 6224 -67 6250
rect -41 6224 -13 6250
rect 13 6224 41 6250
rect 67 6224 73 6250
rect -73 6196 73 6224
rect -73 6170 -67 6196
rect -41 6170 -13 6196
rect 13 6170 41 6196
rect 67 6170 73 6196
rect -73 6142 73 6170
rect -73 6116 -67 6142
rect -41 6116 -13 6142
rect 13 6116 41 6142
rect 67 6116 73 6142
rect -73 6088 73 6116
rect -73 6062 -67 6088
rect -41 6062 -13 6088
rect 13 6062 41 6088
rect 67 6062 73 6088
rect -73 6034 73 6062
rect -73 6008 -67 6034
rect -41 6008 -13 6034
rect 13 6008 41 6034
rect 67 6008 73 6034
rect -73 5980 73 6008
rect -73 5954 -67 5980
rect -41 5954 -13 5980
rect 13 5954 41 5980
rect 67 5954 73 5980
rect -73 5926 73 5954
rect -73 5900 -67 5926
rect -41 5900 -13 5926
rect 13 5900 41 5926
rect 67 5900 73 5926
rect -73 5872 73 5900
rect -73 5846 -67 5872
rect -41 5846 -13 5872
rect 13 5846 41 5872
rect 67 5846 73 5872
rect -73 5818 73 5846
rect -73 5792 -67 5818
rect -41 5792 -13 5818
rect 13 5792 41 5818
rect 67 5792 73 5818
rect -73 5764 73 5792
rect -73 5738 -67 5764
rect -41 5738 -13 5764
rect 13 5738 41 5764
rect 67 5738 73 5764
rect -73 5710 73 5738
rect -73 5684 -67 5710
rect -41 5684 -13 5710
rect 13 5684 41 5710
rect 67 5684 73 5710
rect -73 5656 73 5684
rect -73 5630 -67 5656
rect -41 5630 -13 5656
rect 13 5630 41 5656
rect 67 5630 73 5656
rect -73 5602 73 5630
rect -73 5576 -67 5602
rect -41 5576 -13 5602
rect 13 5576 41 5602
rect 67 5576 73 5602
rect -73 5548 73 5576
rect -73 5522 -67 5548
rect -41 5522 -13 5548
rect 13 5522 41 5548
rect 67 5522 73 5548
rect -73 5494 73 5522
rect -73 5468 -67 5494
rect -41 5468 -13 5494
rect 13 5468 41 5494
rect 67 5468 73 5494
rect -73 5440 73 5468
rect -73 5414 -67 5440
rect -41 5414 -13 5440
rect 13 5414 41 5440
rect 67 5414 73 5440
rect -73 5386 73 5414
rect -73 5360 -67 5386
rect -41 5360 -13 5386
rect 13 5360 41 5386
rect 67 5360 73 5386
rect -73 5332 73 5360
rect -73 5306 -67 5332
rect -41 5306 -13 5332
rect 13 5306 41 5332
rect 67 5306 73 5332
rect -73 5278 73 5306
rect -73 5252 -67 5278
rect -41 5252 -13 5278
rect 13 5252 41 5278
rect 67 5252 73 5278
rect -73 5224 73 5252
rect -73 5198 -67 5224
rect -41 5198 -13 5224
rect 13 5198 41 5224
rect 67 5198 73 5224
rect -73 5170 73 5198
rect -73 5144 -67 5170
rect -41 5144 -13 5170
rect 13 5144 41 5170
rect 67 5144 73 5170
rect -73 5116 73 5144
rect -73 5090 -67 5116
rect -41 5090 -13 5116
rect 13 5090 41 5116
rect 67 5090 73 5116
rect -73 5062 73 5090
rect -73 5036 -67 5062
rect -41 5036 -13 5062
rect 13 5036 41 5062
rect 67 5036 73 5062
rect -73 5008 73 5036
rect -73 4982 -67 5008
rect -41 4982 -13 5008
rect 13 4982 41 5008
rect 67 4982 73 5008
rect -73 4954 73 4982
rect -73 4928 -67 4954
rect -41 4928 -13 4954
rect 13 4928 41 4954
rect 67 4928 73 4954
rect -73 4900 73 4928
rect -73 4874 -67 4900
rect -41 4874 -13 4900
rect 13 4874 41 4900
rect 67 4874 73 4900
rect -73 4846 73 4874
rect -73 4820 -67 4846
rect -41 4820 -13 4846
rect 13 4820 41 4846
rect 67 4820 73 4846
rect -73 4792 73 4820
rect -73 4766 -67 4792
rect -41 4766 -13 4792
rect 13 4766 41 4792
rect 67 4766 73 4792
rect -73 4738 73 4766
rect -73 4712 -67 4738
rect -41 4712 -13 4738
rect 13 4712 41 4738
rect 67 4712 73 4738
rect -73 4684 73 4712
rect -73 4658 -67 4684
rect -41 4658 -13 4684
rect 13 4658 41 4684
rect 67 4658 73 4684
rect -73 4630 73 4658
rect -73 4604 -67 4630
rect -41 4604 -13 4630
rect 13 4604 41 4630
rect 67 4604 73 4630
rect -73 4576 73 4604
rect -73 4550 -67 4576
rect -41 4550 -13 4576
rect 13 4550 41 4576
rect 67 4550 73 4576
rect -73 4522 73 4550
rect -73 4496 -67 4522
rect -41 4496 -13 4522
rect 13 4496 41 4522
rect 67 4496 73 4522
rect -73 4468 73 4496
rect -73 4442 -67 4468
rect -41 4442 -13 4468
rect 13 4442 41 4468
rect 67 4442 73 4468
rect -73 4414 73 4442
rect -73 4388 -67 4414
rect -41 4388 -13 4414
rect 13 4388 41 4414
rect 67 4388 73 4414
rect -73 4360 73 4388
rect -73 4334 -67 4360
rect -41 4334 -13 4360
rect 13 4334 41 4360
rect 67 4334 73 4360
rect -73 4306 73 4334
rect -73 4280 -67 4306
rect -41 4280 -13 4306
rect 13 4280 41 4306
rect 67 4280 73 4306
rect -73 4252 73 4280
rect -73 4226 -67 4252
rect -41 4226 -13 4252
rect 13 4226 41 4252
rect 67 4226 73 4252
rect -73 4198 73 4226
rect -73 4172 -67 4198
rect -41 4172 -13 4198
rect 13 4172 41 4198
rect 67 4172 73 4198
rect -73 4144 73 4172
rect -73 4118 -67 4144
rect -41 4118 -13 4144
rect 13 4118 41 4144
rect 67 4118 73 4144
rect -73 4090 73 4118
rect -73 4064 -67 4090
rect -41 4064 -13 4090
rect 13 4064 41 4090
rect 67 4064 73 4090
rect -73 4036 73 4064
rect -73 4010 -67 4036
rect -41 4010 -13 4036
rect 13 4010 41 4036
rect 67 4010 73 4036
rect -73 3982 73 4010
rect -73 3956 -67 3982
rect -41 3956 -13 3982
rect 13 3956 41 3982
rect 67 3956 73 3982
rect -73 3928 73 3956
rect -73 3902 -67 3928
rect -41 3902 -13 3928
rect 13 3902 41 3928
rect 67 3902 73 3928
rect -73 3874 73 3902
rect -73 3848 -67 3874
rect -41 3848 -13 3874
rect 13 3848 41 3874
rect 67 3848 73 3874
rect -73 3820 73 3848
rect -73 3794 -67 3820
rect -41 3794 -13 3820
rect 13 3794 41 3820
rect 67 3794 73 3820
rect -73 3766 73 3794
rect -73 3740 -67 3766
rect -41 3740 -13 3766
rect 13 3740 41 3766
rect 67 3740 73 3766
rect -73 3712 73 3740
rect -73 3686 -67 3712
rect -41 3686 -13 3712
rect 13 3686 41 3712
rect 67 3686 73 3712
rect -73 3658 73 3686
rect -73 3632 -67 3658
rect -41 3632 -13 3658
rect 13 3632 41 3658
rect 67 3632 73 3658
rect -73 3604 73 3632
rect -73 3578 -67 3604
rect -41 3578 -13 3604
rect 13 3578 41 3604
rect 67 3578 73 3604
rect -73 3550 73 3578
rect -73 3524 -67 3550
rect -41 3524 -13 3550
rect 13 3524 41 3550
rect 67 3524 73 3550
rect -73 3496 73 3524
rect -73 3470 -67 3496
rect -41 3470 -13 3496
rect 13 3470 41 3496
rect 67 3470 73 3496
rect -73 3442 73 3470
rect -73 3416 -67 3442
rect -41 3416 -13 3442
rect 13 3416 41 3442
rect 67 3416 73 3442
rect -73 3388 73 3416
rect -73 3362 -67 3388
rect -41 3362 -13 3388
rect 13 3362 41 3388
rect 67 3362 73 3388
rect -73 3334 73 3362
rect -73 3308 -67 3334
rect -41 3308 -13 3334
rect 13 3308 41 3334
rect 67 3308 73 3334
rect -73 3280 73 3308
rect -73 3254 -67 3280
rect -41 3254 -13 3280
rect 13 3254 41 3280
rect 67 3254 73 3280
rect -73 3226 73 3254
rect -73 3200 -67 3226
rect -41 3200 -13 3226
rect 13 3200 41 3226
rect 67 3200 73 3226
rect -73 3172 73 3200
rect -73 3146 -67 3172
rect -41 3146 -13 3172
rect 13 3146 41 3172
rect 67 3146 73 3172
rect -73 3118 73 3146
rect -73 3092 -67 3118
rect -41 3092 -13 3118
rect 13 3092 41 3118
rect 67 3092 73 3118
rect -73 3064 73 3092
rect -73 3038 -67 3064
rect -41 3038 -13 3064
rect 13 3038 41 3064
rect 67 3038 73 3064
rect -73 3010 73 3038
rect -73 2984 -67 3010
rect -41 2984 -13 3010
rect 13 2984 41 3010
rect 67 2984 73 3010
rect -73 2956 73 2984
rect -73 2930 -67 2956
rect -41 2930 -13 2956
rect 13 2930 41 2956
rect 67 2930 73 2956
rect -73 2902 73 2930
rect -73 2876 -67 2902
rect -41 2876 -13 2902
rect 13 2876 41 2902
rect 67 2876 73 2902
rect -73 2848 73 2876
rect -73 2822 -67 2848
rect -41 2822 -13 2848
rect 13 2822 41 2848
rect 67 2822 73 2848
rect -73 2794 73 2822
rect -73 2768 -67 2794
rect -41 2768 -13 2794
rect 13 2768 41 2794
rect 67 2768 73 2794
rect -73 2740 73 2768
rect -73 2714 -67 2740
rect -41 2714 -13 2740
rect 13 2714 41 2740
rect 67 2714 73 2740
rect -73 2686 73 2714
rect -73 2660 -67 2686
rect -41 2660 -13 2686
rect 13 2660 41 2686
rect 67 2660 73 2686
rect -73 2632 73 2660
rect -73 2606 -67 2632
rect -41 2606 -13 2632
rect 13 2606 41 2632
rect 67 2606 73 2632
rect -73 2578 73 2606
rect -73 2552 -67 2578
rect -41 2552 -13 2578
rect 13 2552 41 2578
rect 67 2552 73 2578
rect -73 2524 73 2552
rect -73 2498 -67 2524
rect -41 2498 -13 2524
rect 13 2498 41 2524
rect 67 2498 73 2524
rect -73 2470 73 2498
rect -73 2444 -67 2470
rect -41 2444 -13 2470
rect 13 2444 41 2470
rect 67 2444 73 2470
rect -73 2416 73 2444
rect -73 2390 -67 2416
rect -41 2390 -13 2416
rect 13 2390 41 2416
rect 67 2390 73 2416
rect -73 2362 73 2390
rect -73 2336 -67 2362
rect -41 2336 -13 2362
rect 13 2336 41 2362
rect 67 2336 73 2362
rect -73 2308 73 2336
rect -73 2282 -67 2308
rect -41 2282 -13 2308
rect 13 2282 41 2308
rect 67 2282 73 2308
rect -73 2254 73 2282
rect -73 2228 -67 2254
rect -41 2228 -13 2254
rect 13 2228 41 2254
rect 67 2228 73 2254
rect -73 2200 73 2228
rect -73 2174 -67 2200
rect -41 2174 -13 2200
rect 13 2174 41 2200
rect 67 2174 73 2200
rect -73 2146 73 2174
rect -73 2120 -67 2146
rect -41 2120 -13 2146
rect 13 2120 41 2146
rect 67 2120 73 2146
rect -73 2092 73 2120
rect -73 2066 -67 2092
rect -41 2066 -13 2092
rect 13 2066 41 2092
rect 67 2066 73 2092
rect -73 2038 73 2066
rect -73 2012 -67 2038
rect -41 2012 -13 2038
rect 13 2012 41 2038
rect 67 2012 73 2038
rect -73 1984 73 2012
rect -73 1958 -67 1984
rect -41 1958 -13 1984
rect 13 1958 41 1984
rect 67 1958 73 1984
rect -73 1930 73 1958
rect -73 1904 -67 1930
rect -41 1904 -13 1930
rect 13 1904 41 1930
rect 67 1904 73 1930
rect -73 1876 73 1904
rect -73 1850 -67 1876
rect -41 1850 -13 1876
rect 13 1850 41 1876
rect 67 1850 73 1876
rect -73 1822 73 1850
rect -73 1796 -67 1822
rect -41 1796 -13 1822
rect 13 1796 41 1822
rect 67 1796 73 1822
rect -73 1768 73 1796
rect -73 1742 -67 1768
rect -41 1742 -13 1768
rect 13 1742 41 1768
rect 67 1742 73 1768
rect -73 1714 73 1742
rect -73 1688 -67 1714
rect -41 1688 -13 1714
rect 13 1688 41 1714
rect 67 1688 73 1714
rect -73 1660 73 1688
rect -73 1634 -67 1660
rect -41 1634 -13 1660
rect 13 1634 41 1660
rect 67 1634 73 1660
rect -73 1606 73 1634
rect -73 1580 -67 1606
rect -41 1580 -13 1606
rect 13 1580 41 1606
rect 67 1580 73 1606
rect -73 1552 73 1580
rect -73 1526 -67 1552
rect -41 1526 -13 1552
rect 13 1526 41 1552
rect 67 1526 73 1552
rect -73 1498 73 1526
rect -73 1472 -67 1498
rect -41 1472 -13 1498
rect 13 1472 41 1498
rect 67 1472 73 1498
rect -73 1444 73 1472
rect -73 1418 -67 1444
rect -41 1418 -13 1444
rect 13 1418 41 1444
rect 67 1418 73 1444
rect -73 1390 73 1418
rect -73 1364 -67 1390
rect -41 1364 -13 1390
rect 13 1364 41 1390
rect 67 1364 73 1390
rect -73 1336 73 1364
rect -73 1310 -67 1336
rect -41 1310 -13 1336
rect 13 1310 41 1336
rect 67 1310 73 1336
rect -73 1282 73 1310
rect -73 1256 -67 1282
rect -41 1256 -13 1282
rect 13 1256 41 1282
rect 67 1256 73 1282
rect -73 1228 73 1256
rect -73 1202 -67 1228
rect -41 1202 -13 1228
rect 13 1202 41 1228
rect 67 1202 73 1228
rect -73 1174 73 1202
rect -73 1148 -67 1174
rect -41 1148 -13 1174
rect 13 1148 41 1174
rect 67 1148 73 1174
rect -73 1120 73 1148
rect -73 1094 -67 1120
rect -41 1094 -13 1120
rect 13 1094 41 1120
rect 67 1094 73 1120
rect -73 1066 73 1094
rect -73 1040 -67 1066
rect -41 1040 -13 1066
rect 13 1040 41 1066
rect 67 1040 73 1066
rect -73 1012 73 1040
rect -73 986 -67 1012
rect -41 986 -13 1012
rect 13 986 41 1012
rect 67 986 73 1012
rect -73 958 73 986
rect -73 932 -67 958
rect -41 932 -13 958
rect 13 932 41 958
rect 67 932 73 958
rect -73 904 73 932
rect -73 878 -67 904
rect -41 878 -13 904
rect 13 878 41 904
rect 67 878 73 904
rect -73 850 73 878
rect -73 824 -67 850
rect -41 824 -13 850
rect 13 824 41 850
rect 67 824 73 850
rect -73 796 73 824
rect -73 770 -67 796
rect -41 770 -13 796
rect 13 770 41 796
rect 67 770 73 796
rect -73 742 73 770
rect -73 716 -67 742
rect -41 716 -13 742
rect 13 716 41 742
rect 67 716 73 742
rect -73 688 73 716
rect -73 662 -67 688
rect -41 662 -13 688
rect 13 662 41 688
rect 67 662 73 688
rect -73 634 73 662
rect -73 608 -67 634
rect -41 608 -13 634
rect 13 608 41 634
rect 67 608 73 634
rect -73 580 73 608
rect -73 554 -67 580
rect -41 554 -13 580
rect 13 554 41 580
rect 67 554 73 580
rect -73 526 73 554
rect -73 500 -67 526
rect -41 500 -13 526
rect 13 500 41 526
rect 67 500 73 526
rect -73 472 73 500
rect -73 446 -67 472
rect -41 446 -13 472
rect 13 446 41 472
rect 67 446 73 472
rect -73 418 73 446
rect -73 392 -67 418
rect -41 392 -13 418
rect 13 392 41 418
rect 67 392 73 418
rect -73 364 73 392
rect -73 338 -67 364
rect -41 338 -13 364
rect 13 338 41 364
rect 67 338 73 364
rect -73 310 73 338
rect -73 284 -67 310
rect -41 284 -13 310
rect 13 284 41 310
rect 67 284 73 310
rect -73 256 73 284
rect -73 230 -67 256
rect -41 230 -13 256
rect 13 230 41 256
rect 67 230 73 256
rect -73 202 73 230
rect -73 176 -67 202
rect -41 176 -13 202
rect 13 176 41 202
rect 67 176 73 202
rect -73 148 73 176
rect -73 122 -67 148
rect -41 122 -13 148
rect 13 122 41 148
rect 67 122 73 148
rect -73 94 73 122
rect -73 68 -67 94
rect -41 68 -13 94
rect 13 68 41 94
rect 67 68 73 94
rect -73 40 73 68
rect -73 14 -67 40
rect -41 14 -13 40
rect 13 14 41 40
rect 67 14 73 40
rect -73 -14 73 14
rect -73 -40 -67 -14
rect -41 -40 -13 -14
rect 13 -40 41 -14
rect 67 -40 73 -14
rect -73 -68 73 -40
rect -73 -94 -67 -68
rect -41 -94 -13 -68
rect 13 -94 41 -68
rect 67 -94 73 -68
rect -73 -122 73 -94
rect -73 -148 -67 -122
rect -41 -148 -13 -122
rect 13 -148 41 -122
rect 67 -148 73 -122
rect -73 -176 73 -148
rect -73 -202 -67 -176
rect -41 -202 -13 -176
rect 13 -202 41 -176
rect 67 -202 73 -176
rect -73 -230 73 -202
rect -73 -256 -67 -230
rect -41 -256 -13 -230
rect 13 -256 41 -230
rect 67 -256 73 -230
rect -73 -284 73 -256
rect -73 -310 -67 -284
rect -41 -310 -13 -284
rect 13 -310 41 -284
rect 67 -310 73 -284
rect -73 -338 73 -310
rect -73 -364 -67 -338
rect -41 -364 -13 -338
rect 13 -364 41 -338
rect 67 -364 73 -338
rect -73 -392 73 -364
rect -73 -418 -67 -392
rect -41 -418 -13 -392
rect 13 -418 41 -392
rect 67 -418 73 -392
rect -73 -446 73 -418
rect -73 -472 -67 -446
rect -41 -472 -13 -446
rect 13 -472 41 -446
rect 67 -472 73 -446
rect -73 -500 73 -472
rect -73 -526 -67 -500
rect -41 -526 -13 -500
rect 13 -526 41 -500
rect 67 -526 73 -500
rect -73 -554 73 -526
rect -73 -580 -67 -554
rect -41 -580 -13 -554
rect 13 -580 41 -554
rect 67 -580 73 -554
rect -73 -608 73 -580
rect -73 -634 -67 -608
rect -41 -634 -13 -608
rect 13 -634 41 -608
rect 67 -634 73 -608
rect -73 -662 73 -634
rect -73 -688 -67 -662
rect -41 -688 -13 -662
rect 13 -688 41 -662
rect 67 -688 73 -662
rect -73 -716 73 -688
rect -73 -742 -67 -716
rect -41 -742 -13 -716
rect 13 -742 41 -716
rect 67 -742 73 -716
rect -73 -770 73 -742
rect -73 -796 -67 -770
rect -41 -796 -13 -770
rect 13 -796 41 -770
rect 67 -796 73 -770
rect -73 -824 73 -796
rect -73 -850 -67 -824
rect -41 -850 -13 -824
rect 13 -850 41 -824
rect 67 -850 73 -824
rect -73 -878 73 -850
rect -73 -904 -67 -878
rect -41 -904 -13 -878
rect 13 -904 41 -878
rect 67 -904 73 -878
rect -73 -932 73 -904
rect -73 -958 -67 -932
rect -41 -958 -13 -932
rect 13 -958 41 -932
rect 67 -958 73 -932
rect -73 -986 73 -958
rect -73 -1012 -67 -986
rect -41 -1012 -13 -986
rect 13 -1012 41 -986
rect 67 -1012 73 -986
rect -73 -1040 73 -1012
rect -73 -1066 -67 -1040
rect -41 -1066 -13 -1040
rect 13 -1066 41 -1040
rect 67 -1066 73 -1040
rect -73 -1094 73 -1066
rect -73 -1120 -67 -1094
rect -41 -1120 -13 -1094
rect 13 -1120 41 -1094
rect 67 -1120 73 -1094
rect -73 -1148 73 -1120
rect -73 -1174 -67 -1148
rect -41 -1174 -13 -1148
rect 13 -1174 41 -1148
rect 67 -1174 73 -1148
rect -73 -1202 73 -1174
rect -73 -1228 -67 -1202
rect -41 -1228 -13 -1202
rect 13 -1228 41 -1202
rect 67 -1228 73 -1202
rect -73 -1256 73 -1228
rect -73 -1282 -67 -1256
rect -41 -1282 -13 -1256
rect 13 -1282 41 -1256
rect 67 -1282 73 -1256
rect -73 -1310 73 -1282
rect -73 -1336 -67 -1310
rect -41 -1336 -13 -1310
rect 13 -1336 41 -1310
rect 67 -1336 73 -1310
rect -73 -1364 73 -1336
rect -73 -1390 -67 -1364
rect -41 -1390 -13 -1364
rect 13 -1390 41 -1364
rect 67 -1390 73 -1364
rect -73 -1418 73 -1390
rect -73 -1444 -67 -1418
rect -41 -1444 -13 -1418
rect 13 -1444 41 -1418
rect 67 -1444 73 -1418
rect -73 -1472 73 -1444
rect -73 -1498 -67 -1472
rect -41 -1498 -13 -1472
rect 13 -1498 41 -1472
rect 67 -1498 73 -1472
rect -73 -1526 73 -1498
rect -73 -1552 -67 -1526
rect -41 -1552 -13 -1526
rect 13 -1552 41 -1526
rect 67 -1552 73 -1526
rect -73 -1580 73 -1552
rect -73 -1606 -67 -1580
rect -41 -1606 -13 -1580
rect 13 -1606 41 -1580
rect 67 -1606 73 -1580
rect -73 -1634 73 -1606
rect -73 -1660 -67 -1634
rect -41 -1660 -13 -1634
rect 13 -1660 41 -1634
rect 67 -1660 73 -1634
rect -73 -1688 73 -1660
rect -73 -1714 -67 -1688
rect -41 -1714 -13 -1688
rect 13 -1714 41 -1688
rect 67 -1714 73 -1688
rect -73 -1742 73 -1714
rect -73 -1768 -67 -1742
rect -41 -1768 -13 -1742
rect 13 -1768 41 -1742
rect 67 -1768 73 -1742
rect -73 -1796 73 -1768
rect -73 -1822 -67 -1796
rect -41 -1822 -13 -1796
rect 13 -1822 41 -1796
rect 67 -1822 73 -1796
rect -73 -1850 73 -1822
rect -73 -1876 -67 -1850
rect -41 -1876 -13 -1850
rect 13 -1876 41 -1850
rect 67 -1876 73 -1850
rect -73 -1904 73 -1876
rect -73 -1930 -67 -1904
rect -41 -1930 -13 -1904
rect 13 -1930 41 -1904
rect 67 -1930 73 -1904
rect -73 -1958 73 -1930
rect -73 -1984 -67 -1958
rect -41 -1984 -13 -1958
rect 13 -1984 41 -1958
rect 67 -1984 73 -1958
rect -73 -2012 73 -1984
rect -73 -2038 -67 -2012
rect -41 -2038 -13 -2012
rect 13 -2038 41 -2012
rect 67 -2038 73 -2012
rect -73 -2066 73 -2038
rect -73 -2092 -67 -2066
rect -41 -2092 -13 -2066
rect 13 -2092 41 -2066
rect 67 -2092 73 -2066
rect -73 -2120 73 -2092
rect -73 -2146 -67 -2120
rect -41 -2146 -13 -2120
rect 13 -2146 41 -2120
rect 67 -2146 73 -2120
rect -73 -2174 73 -2146
rect -73 -2200 -67 -2174
rect -41 -2200 -13 -2174
rect 13 -2200 41 -2174
rect 67 -2200 73 -2174
rect -73 -2228 73 -2200
rect -73 -2254 -67 -2228
rect -41 -2254 -13 -2228
rect 13 -2254 41 -2228
rect 67 -2254 73 -2228
rect -73 -2282 73 -2254
rect -73 -2308 -67 -2282
rect -41 -2308 -13 -2282
rect 13 -2308 41 -2282
rect 67 -2308 73 -2282
rect -73 -2336 73 -2308
rect -73 -2362 -67 -2336
rect -41 -2362 -13 -2336
rect 13 -2362 41 -2336
rect 67 -2362 73 -2336
rect -73 -2390 73 -2362
rect -73 -2416 -67 -2390
rect -41 -2416 -13 -2390
rect 13 -2416 41 -2390
rect 67 -2416 73 -2390
rect -73 -2444 73 -2416
rect -73 -2470 -67 -2444
rect -41 -2470 -13 -2444
rect 13 -2470 41 -2444
rect 67 -2470 73 -2444
rect -73 -2498 73 -2470
rect -73 -2524 -67 -2498
rect -41 -2524 -13 -2498
rect 13 -2524 41 -2498
rect 67 -2524 73 -2498
rect -73 -2552 73 -2524
rect -73 -2578 -67 -2552
rect -41 -2578 -13 -2552
rect 13 -2578 41 -2552
rect 67 -2578 73 -2552
rect -73 -2606 73 -2578
rect -73 -2632 -67 -2606
rect -41 -2632 -13 -2606
rect 13 -2632 41 -2606
rect 67 -2632 73 -2606
rect -73 -2660 73 -2632
rect -73 -2686 -67 -2660
rect -41 -2686 -13 -2660
rect 13 -2686 41 -2660
rect 67 -2686 73 -2660
rect -73 -2714 73 -2686
rect -73 -2740 -67 -2714
rect -41 -2740 -13 -2714
rect 13 -2740 41 -2714
rect 67 -2740 73 -2714
rect -73 -2768 73 -2740
rect -73 -2794 -67 -2768
rect -41 -2794 -13 -2768
rect 13 -2794 41 -2768
rect 67 -2794 73 -2768
rect -73 -2822 73 -2794
rect -73 -2848 -67 -2822
rect -41 -2848 -13 -2822
rect 13 -2848 41 -2822
rect 67 -2848 73 -2822
rect -73 -2876 73 -2848
rect -73 -2902 -67 -2876
rect -41 -2902 -13 -2876
rect 13 -2902 41 -2876
rect 67 -2902 73 -2876
rect -73 -2930 73 -2902
rect -73 -2956 -67 -2930
rect -41 -2956 -13 -2930
rect 13 -2956 41 -2930
rect 67 -2956 73 -2930
rect -73 -2984 73 -2956
rect -73 -3010 -67 -2984
rect -41 -3010 -13 -2984
rect 13 -3010 41 -2984
rect 67 -3010 73 -2984
rect -73 -3038 73 -3010
rect -73 -3064 -67 -3038
rect -41 -3064 -13 -3038
rect 13 -3064 41 -3038
rect 67 -3064 73 -3038
rect -73 -3092 73 -3064
rect -73 -3118 -67 -3092
rect -41 -3118 -13 -3092
rect 13 -3118 41 -3092
rect 67 -3118 73 -3092
rect -73 -3146 73 -3118
rect -73 -3172 -67 -3146
rect -41 -3172 -13 -3146
rect 13 -3172 41 -3146
rect 67 -3172 73 -3146
rect -73 -3200 73 -3172
rect -73 -3226 -67 -3200
rect -41 -3226 -13 -3200
rect 13 -3226 41 -3200
rect 67 -3226 73 -3200
rect -73 -3254 73 -3226
rect -73 -3280 -67 -3254
rect -41 -3280 -13 -3254
rect 13 -3280 41 -3254
rect 67 -3280 73 -3254
rect -73 -3308 73 -3280
rect -73 -3334 -67 -3308
rect -41 -3334 -13 -3308
rect 13 -3334 41 -3308
rect 67 -3334 73 -3308
rect -73 -3362 73 -3334
rect -73 -3388 -67 -3362
rect -41 -3388 -13 -3362
rect 13 -3388 41 -3362
rect 67 -3388 73 -3362
rect -73 -3416 73 -3388
rect -73 -3442 -67 -3416
rect -41 -3442 -13 -3416
rect 13 -3442 41 -3416
rect 67 -3442 73 -3416
rect -73 -3470 73 -3442
rect -73 -3496 -67 -3470
rect -41 -3496 -13 -3470
rect 13 -3496 41 -3470
rect 67 -3496 73 -3470
rect -73 -3524 73 -3496
rect -73 -3550 -67 -3524
rect -41 -3550 -13 -3524
rect 13 -3550 41 -3524
rect 67 -3550 73 -3524
rect -73 -3578 73 -3550
rect -73 -3604 -67 -3578
rect -41 -3604 -13 -3578
rect 13 -3604 41 -3578
rect 67 -3604 73 -3578
rect -73 -3632 73 -3604
rect -73 -3658 -67 -3632
rect -41 -3658 -13 -3632
rect 13 -3658 41 -3632
rect 67 -3658 73 -3632
rect -73 -3686 73 -3658
rect -73 -3712 -67 -3686
rect -41 -3712 -13 -3686
rect 13 -3712 41 -3686
rect 67 -3712 73 -3686
rect -73 -3740 73 -3712
rect -73 -3766 -67 -3740
rect -41 -3766 -13 -3740
rect 13 -3766 41 -3740
rect 67 -3766 73 -3740
rect -73 -3794 73 -3766
rect -73 -3820 -67 -3794
rect -41 -3820 -13 -3794
rect 13 -3820 41 -3794
rect 67 -3820 73 -3794
rect -73 -3848 73 -3820
rect -73 -3874 -67 -3848
rect -41 -3874 -13 -3848
rect 13 -3874 41 -3848
rect 67 -3874 73 -3848
rect -73 -3902 73 -3874
rect -73 -3928 -67 -3902
rect -41 -3928 -13 -3902
rect 13 -3928 41 -3902
rect 67 -3928 73 -3902
rect -73 -3956 73 -3928
rect -73 -3982 -67 -3956
rect -41 -3982 -13 -3956
rect 13 -3982 41 -3956
rect 67 -3982 73 -3956
rect -73 -4010 73 -3982
rect -73 -4036 -67 -4010
rect -41 -4036 -13 -4010
rect 13 -4036 41 -4010
rect 67 -4036 73 -4010
rect -73 -4064 73 -4036
rect -73 -4090 -67 -4064
rect -41 -4090 -13 -4064
rect 13 -4090 41 -4064
rect 67 -4090 73 -4064
rect -73 -4118 73 -4090
rect -73 -4144 -67 -4118
rect -41 -4144 -13 -4118
rect 13 -4144 41 -4118
rect 67 -4144 73 -4118
rect -73 -4172 73 -4144
rect -73 -4198 -67 -4172
rect -41 -4198 -13 -4172
rect 13 -4198 41 -4172
rect 67 -4198 73 -4172
rect -73 -4226 73 -4198
rect -73 -4252 -67 -4226
rect -41 -4252 -13 -4226
rect 13 -4252 41 -4226
rect 67 -4252 73 -4226
rect -73 -4280 73 -4252
rect -73 -4306 -67 -4280
rect -41 -4306 -13 -4280
rect 13 -4306 41 -4280
rect 67 -4306 73 -4280
rect -73 -4334 73 -4306
rect -73 -4360 -67 -4334
rect -41 -4360 -13 -4334
rect 13 -4360 41 -4334
rect 67 -4360 73 -4334
rect -73 -4388 73 -4360
rect -73 -4414 -67 -4388
rect -41 -4414 -13 -4388
rect 13 -4414 41 -4388
rect 67 -4414 73 -4388
rect -73 -4442 73 -4414
rect -73 -4468 -67 -4442
rect -41 -4468 -13 -4442
rect 13 -4468 41 -4442
rect 67 -4468 73 -4442
rect -73 -4496 73 -4468
rect -73 -4522 -67 -4496
rect -41 -4522 -13 -4496
rect 13 -4522 41 -4496
rect 67 -4522 73 -4496
rect -73 -4550 73 -4522
rect -73 -4576 -67 -4550
rect -41 -4576 -13 -4550
rect 13 -4576 41 -4550
rect 67 -4576 73 -4550
rect -73 -4604 73 -4576
rect -73 -4630 -67 -4604
rect -41 -4630 -13 -4604
rect 13 -4630 41 -4604
rect 67 -4630 73 -4604
rect -73 -4658 73 -4630
rect -73 -4684 -67 -4658
rect -41 -4684 -13 -4658
rect 13 -4684 41 -4658
rect 67 -4684 73 -4658
rect -73 -4712 73 -4684
rect -73 -4738 -67 -4712
rect -41 -4738 -13 -4712
rect 13 -4738 41 -4712
rect 67 -4738 73 -4712
rect -73 -4766 73 -4738
rect -73 -4792 -67 -4766
rect -41 -4792 -13 -4766
rect 13 -4792 41 -4766
rect 67 -4792 73 -4766
rect -73 -4820 73 -4792
rect -73 -4846 -67 -4820
rect -41 -4846 -13 -4820
rect 13 -4846 41 -4820
rect 67 -4846 73 -4820
rect -73 -4874 73 -4846
rect -73 -4900 -67 -4874
rect -41 -4900 -13 -4874
rect 13 -4900 41 -4874
rect 67 -4900 73 -4874
rect -73 -4928 73 -4900
rect -73 -4954 -67 -4928
rect -41 -4954 -13 -4928
rect 13 -4954 41 -4928
rect 67 -4954 73 -4928
rect -73 -4982 73 -4954
rect -73 -5008 -67 -4982
rect -41 -5008 -13 -4982
rect 13 -5008 41 -4982
rect 67 -5008 73 -4982
rect -73 -5036 73 -5008
rect -73 -5062 -67 -5036
rect -41 -5062 -13 -5036
rect 13 -5062 41 -5036
rect 67 -5062 73 -5036
rect -73 -5090 73 -5062
rect -73 -5116 -67 -5090
rect -41 -5116 -13 -5090
rect 13 -5116 41 -5090
rect 67 -5116 73 -5090
rect -73 -5144 73 -5116
rect -73 -5170 -67 -5144
rect -41 -5170 -13 -5144
rect 13 -5170 41 -5144
rect 67 -5170 73 -5144
rect -73 -5198 73 -5170
rect -73 -5224 -67 -5198
rect -41 -5224 -13 -5198
rect 13 -5224 41 -5198
rect 67 -5224 73 -5198
rect -73 -5252 73 -5224
rect -73 -5278 -67 -5252
rect -41 -5278 -13 -5252
rect 13 -5278 41 -5252
rect 67 -5278 73 -5252
rect -73 -5306 73 -5278
rect -73 -5332 -67 -5306
rect -41 -5332 -13 -5306
rect 13 -5332 41 -5306
rect 67 -5332 73 -5306
rect -73 -5360 73 -5332
rect -73 -5386 -67 -5360
rect -41 -5386 -13 -5360
rect 13 -5386 41 -5360
rect 67 -5386 73 -5360
rect -73 -5414 73 -5386
rect -73 -5440 -67 -5414
rect -41 -5440 -13 -5414
rect 13 -5440 41 -5414
rect 67 -5440 73 -5414
rect -73 -5468 73 -5440
rect -73 -5494 -67 -5468
rect -41 -5494 -13 -5468
rect 13 -5494 41 -5468
rect 67 -5494 73 -5468
rect -73 -5522 73 -5494
rect -73 -5548 -67 -5522
rect -41 -5548 -13 -5522
rect 13 -5548 41 -5522
rect 67 -5548 73 -5522
rect -73 -5576 73 -5548
rect -73 -5602 -67 -5576
rect -41 -5602 -13 -5576
rect 13 -5602 41 -5576
rect 67 -5602 73 -5576
rect -73 -5630 73 -5602
rect -73 -5656 -67 -5630
rect -41 -5656 -13 -5630
rect 13 -5656 41 -5630
rect 67 -5656 73 -5630
rect -73 -5684 73 -5656
rect -73 -5710 -67 -5684
rect -41 -5710 -13 -5684
rect 13 -5710 41 -5684
rect 67 -5710 73 -5684
rect -73 -5738 73 -5710
rect -73 -5764 -67 -5738
rect -41 -5764 -13 -5738
rect 13 -5764 41 -5738
rect 67 -5764 73 -5738
rect -73 -5792 73 -5764
rect -73 -5818 -67 -5792
rect -41 -5818 -13 -5792
rect 13 -5818 41 -5792
rect 67 -5818 73 -5792
rect -73 -5846 73 -5818
rect -73 -5872 -67 -5846
rect -41 -5872 -13 -5846
rect 13 -5872 41 -5846
rect 67 -5872 73 -5846
rect -73 -5900 73 -5872
rect -73 -5926 -67 -5900
rect -41 -5926 -13 -5900
rect 13 -5926 41 -5900
rect 67 -5926 73 -5900
rect -73 -5954 73 -5926
rect -73 -5980 -67 -5954
rect -41 -5980 -13 -5954
rect 13 -5980 41 -5954
rect 67 -5980 73 -5954
rect -73 -6008 73 -5980
rect -73 -6034 -67 -6008
rect -41 -6034 -13 -6008
rect 13 -6034 41 -6008
rect 67 -6034 73 -6008
rect -73 -6062 73 -6034
rect -73 -6088 -67 -6062
rect -41 -6088 -13 -6062
rect 13 -6088 41 -6062
rect 67 -6088 73 -6062
rect -73 -6116 73 -6088
rect -73 -6142 -67 -6116
rect -41 -6142 -13 -6116
rect 13 -6142 41 -6116
rect 67 -6142 73 -6116
rect -73 -6170 73 -6142
rect -73 -6196 -67 -6170
rect -41 -6196 -13 -6170
rect 13 -6196 41 -6170
rect 67 -6196 73 -6170
rect -73 -6224 73 -6196
rect -73 -6250 -67 -6224
rect -41 -6250 -13 -6224
rect 13 -6250 41 -6224
rect 67 -6250 73 -6224
rect -73 -6278 73 -6250
rect -73 -6304 -67 -6278
rect -41 -6304 -13 -6278
rect 13 -6304 41 -6278
rect 67 -6304 73 -6278
rect -73 -6310 73 -6304
<< via1 >>
rect -67 6278 -41 6304
rect -13 6278 13 6304
rect 41 6278 67 6304
rect -67 6224 -41 6250
rect -13 6224 13 6250
rect 41 6224 67 6250
rect -67 6170 -41 6196
rect -13 6170 13 6196
rect 41 6170 67 6196
rect -67 6116 -41 6142
rect -13 6116 13 6142
rect 41 6116 67 6142
rect -67 6062 -41 6088
rect -13 6062 13 6088
rect 41 6062 67 6088
rect -67 6008 -41 6034
rect -13 6008 13 6034
rect 41 6008 67 6034
rect -67 5954 -41 5980
rect -13 5954 13 5980
rect 41 5954 67 5980
rect -67 5900 -41 5926
rect -13 5900 13 5926
rect 41 5900 67 5926
rect -67 5846 -41 5872
rect -13 5846 13 5872
rect 41 5846 67 5872
rect -67 5792 -41 5818
rect -13 5792 13 5818
rect 41 5792 67 5818
rect -67 5738 -41 5764
rect -13 5738 13 5764
rect 41 5738 67 5764
rect -67 5684 -41 5710
rect -13 5684 13 5710
rect 41 5684 67 5710
rect -67 5630 -41 5656
rect -13 5630 13 5656
rect 41 5630 67 5656
rect -67 5576 -41 5602
rect -13 5576 13 5602
rect 41 5576 67 5602
rect -67 5522 -41 5548
rect -13 5522 13 5548
rect 41 5522 67 5548
rect -67 5468 -41 5494
rect -13 5468 13 5494
rect 41 5468 67 5494
rect -67 5414 -41 5440
rect -13 5414 13 5440
rect 41 5414 67 5440
rect -67 5360 -41 5386
rect -13 5360 13 5386
rect 41 5360 67 5386
rect -67 5306 -41 5332
rect -13 5306 13 5332
rect 41 5306 67 5332
rect -67 5252 -41 5278
rect -13 5252 13 5278
rect 41 5252 67 5278
rect -67 5198 -41 5224
rect -13 5198 13 5224
rect 41 5198 67 5224
rect -67 5144 -41 5170
rect -13 5144 13 5170
rect 41 5144 67 5170
rect -67 5090 -41 5116
rect -13 5090 13 5116
rect 41 5090 67 5116
rect -67 5036 -41 5062
rect -13 5036 13 5062
rect 41 5036 67 5062
rect -67 4982 -41 5008
rect -13 4982 13 5008
rect 41 4982 67 5008
rect -67 4928 -41 4954
rect -13 4928 13 4954
rect 41 4928 67 4954
rect -67 4874 -41 4900
rect -13 4874 13 4900
rect 41 4874 67 4900
rect -67 4820 -41 4846
rect -13 4820 13 4846
rect 41 4820 67 4846
rect -67 4766 -41 4792
rect -13 4766 13 4792
rect 41 4766 67 4792
rect -67 4712 -41 4738
rect -13 4712 13 4738
rect 41 4712 67 4738
rect -67 4658 -41 4684
rect -13 4658 13 4684
rect 41 4658 67 4684
rect -67 4604 -41 4630
rect -13 4604 13 4630
rect 41 4604 67 4630
rect -67 4550 -41 4576
rect -13 4550 13 4576
rect 41 4550 67 4576
rect -67 4496 -41 4522
rect -13 4496 13 4522
rect 41 4496 67 4522
rect -67 4442 -41 4468
rect -13 4442 13 4468
rect 41 4442 67 4468
rect -67 4388 -41 4414
rect -13 4388 13 4414
rect 41 4388 67 4414
rect -67 4334 -41 4360
rect -13 4334 13 4360
rect 41 4334 67 4360
rect -67 4280 -41 4306
rect -13 4280 13 4306
rect 41 4280 67 4306
rect -67 4226 -41 4252
rect -13 4226 13 4252
rect 41 4226 67 4252
rect -67 4172 -41 4198
rect -13 4172 13 4198
rect 41 4172 67 4198
rect -67 4118 -41 4144
rect -13 4118 13 4144
rect 41 4118 67 4144
rect -67 4064 -41 4090
rect -13 4064 13 4090
rect 41 4064 67 4090
rect -67 4010 -41 4036
rect -13 4010 13 4036
rect 41 4010 67 4036
rect -67 3956 -41 3982
rect -13 3956 13 3982
rect 41 3956 67 3982
rect -67 3902 -41 3928
rect -13 3902 13 3928
rect 41 3902 67 3928
rect -67 3848 -41 3874
rect -13 3848 13 3874
rect 41 3848 67 3874
rect -67 3794 -41 3820
rect -13 3794 13 3820
rect 41 3794 67 3820
rect -67 3740 -41 3766
rect -13 3740 13 3766
rect 41 3740 67 3766
rect -67 3686 -41 3712
rect -13 3686 13 3712
rect 41 3686 67 3712
rect -67 3632 -41 3658
rect -13 3632 13 3658
rect 41 3632 67 3658
rect -67 3578 -41 3604
rect -13 3578 13 3604
rect 41 3578 67 3604
rect -67 3524 -41 3550
rect -13 3524 13 3550
rect 41 3524 67 3550
rect -67 3470 -41 3496
rect -13 3470 13 3496
rect 41 3470 67 3496
rect -67 3416 -41 3442
rect -13 3416 13 3442
rect 41 3416 67 3442
rect -67 3362 -41 3388
rect -13 3362 13 3388
rect 41 3362 67 3388
rect -67 3308 -41 3334
rect -13 3308 13 3334
rect 41 3308 67 3334
rect -67 3254 -41 3280
rect -13 3254 13 3280
rect 41 3254 67 3280
rect -67 3200 -41 3226
rect -13 3200 13 3226
rect 41 3200 67 3226
rect -67 3146 -41 3172
rect -13 3146 13 3172
rect 41 3146 67 3172
rect -67 3092 -41 3118
rect -13 3092 13 3118
rect 41 3092 67 3118
rect -67 3038 -41 3064
rect -13 3038 13 3064
rect 41 3038 67 3064
rect -67 2984 -41 3010
rect -13 2984 13 3010
rect 41 2984 67 3010
rect -67 2930 -41 2956
rect -13 2930 13 2956
rect 41 2930 67 2956
rect -67 2876 -41 2902
rect -13 2876 13 2902
rect 41 2876 67 2902
rect -67 2822 -41 2848
rect -13 2822 13 2848
rect 41 2822 67 2848
rect -67 2768 -41 2794
rect -13 2768 13 2794
rect 41 2768 67 2794
rect -67 2714 -41 2740
rect -13 2714 13 2740
rect 41 2714 67 2740
rect -67 2660 -41 2686
rect -13 2660 13 2686
rect 41 2660 67 2686
rect -67 2606 -41 2632
rect -13 2606 13 2632
rect 41 2606 67 2632
rect -67 2552 -41 2578
rect -13 2552 13 2578
rect 41 2552 67 2578
rect -67 2498 -41 2524
rect -13 2498 13 2524
rect 41 2498 67 2524
rect -67 2444 -41 2470
rect -13 2444 13 2470
rect 41 2444 67 2470
rect -67 2390 -41 2416
rect -13 2390 13 2416
rect 41 2390 67 2416
rect -67 2336 -41 2362
rect -13 2336 13 2362
rect 41 2336 67 2362
rect -67 2282 -41 2308
rect -13 2282 13 2308
rect 41 2282 67 2308
rect -67 2228 -41 2254
rect -13 2228 13 2254
rect 41 2228 67 2254
rect -67 2174 -41 2200
rect -13 2174 13 2200
rect 41 2174 67 2200
rect -67 2120 -41 2146
rect -13 2120 13 2146
rect 41 2120 67 2146
rect -67 2066 -41 2092
rect -13 2066 13 2092
rect 41 2066 67 2092
rect -67 2012 -41 2038
rect -13 2012 13 2038
rect 41 2012 67 2038
rect -67 1958 -41 1984
rect -13 1958 13 1984
rect 41 1958 67 1984
rect -67 1904 -41 1930
rect -13 1904 13 1930
rect 41 1904 67 1930
rect -67 1850 -41 1876
rect -13 1850 13 1876
rect 41 1850 67 1876
rect -67 1796 -41 1822
rect -13 1796 13 1822
rect 41 1796 67 1822
rect -67 1742 -41 1768
rect -13 1742 13 1768
rect 41 1742 67 1768
rect -67 1688 -41 1714
rect -13 1688 13 1714
rect 41 1688 67 1714
rect -67 1634 -41 1660
rect -13 1634 13 1660
rect 41 1634 67 1660
rect -67 1580 -41 1606
rect -13 1580 13 1606
rect 41 1580 67 1606
rect -67 1526 -41 1552
rect -13 1526 13 1552
rect 41 1526 67 1552
rect -67 1472 -41 1498
rect -13 1472 13 1498
rect 41 1472 67 1498
rect -67 1418 -41 1444
rect -13 1418 13 1444
rect 41 1418 67 1444
rect -67 1364 -41 1390
rect -13 1364 13 1390
rect 41 1364 67 1390
rect -67 1310 -41 1336
rect -13 1310 13 1336
rect 41 1310 67 1336
rect -67 1256 -41 1282
rect -13 1256 13 1282
rect 41 1256 67 1282
rect -67 1202 -41 1228
rect -13 1202 13 1228
rect 41 1202 67 1228
rect -67 1148 -41 1174
rect -13 1148 13 1174
rect 41 1148 67 1174
rect -67 1094 -41 1120
rect -13 1094 13 1120
rect 41 1094 67 1120
rect -67 1040 -41 1066
rect -13 1040 13 1066
rect 41 1040 67 1066
rect -67 986 -41 1012
rect -13 986 13 1012
rect 41 986 67 1012
rect -67 932 -41 958
rect -13 932 13 958
rect 41 932 67 958
rect -67 878 -41 904
rect -13 878 13 904
rect 41 878 67 904
rect -67 824 -41 850
rect -13 824 13 850
rect 41 824 67 850
rect -67 770 -41 796
rect -13 770 13 796
rect 41 770 67 796
rect -67 716 -41 742
rect -13 716 13 742
rect 41 716 67 742
rect -67 662 -41 688
rect -13 662 13 688
rect 41 662 67 688
rect -67 608 -41 634
rect -13 608 13 634
rect 41 608 67 634
rect -67 554 -41 580
rect -13 554 13 580
rect 41 554 67 580
rect -67 500 -41 526
rect -13 500 13 526
rect 41 500 67 526
rect -67 446 -41 472
rect -13 446 13 472
rect 41 446 67 472
rect -67 392 -41 418
rect -13 392 13 418
rect 41 392 67 418
rect -67 338 -41 364
rect -13 338 13 364
rect 41 338 67 364
rect -67 284 -41 310
rect -13 284 13 310
rect 41 284 67 310
rect -67 230 -41 256
rect -13 230 13 256
rect 41 230 67 256
rect -67 176 -41 202
rect -13 176 13 202
rect 41 176 67 202
rect -67 122 -41 148
rect -13 122 13 148
rect 41 122 67 148
rect -67 68 -41 94
rect -13 68 13 94
rect 41 68 67 94
rect -67 14 -41 40
rect -13 14 13 40
rect 41 14 67 40
rect -67 -40 -41 -14
rect -13 -40 13 -14
rect 41 -40 67 -14
rect -67 -94 -41 -68
rect -13 -94 13 -68
rect 41 -94 67 -68
rect -67 -148 -41 -122
rect -13 -148 13 -122
rect 41 -148 67 -122
rect -67 -202 -41 -176
rect -13 -202 13 -176
rect 41 -202 67 -176
rect -67 -256 -41 -230
rect -13 -256 13 -230
rect 41 -256 67 -230
rect -67 -310 -41 -284
rect -13 -310 13 -284
rect 41 -310 67 -284
rect -67 -364 -41 -338
rect -13 -364 13 -338
rect 41 -364 67 -338
rect -67 -418 -41 -392
rect -13 -418 13 -392
rect 41 -418 67 -392
rect -67 -472 -41 -446
rect -13 -472 13 -446
rect 41 -472 67 -446
rect -67 -526 -41 -500
rect -13 -526 13 -500
rect 41 -526 67 -500
rect -67 -580 -41 -554
rect -13 -580 13 -554
rect 41 -580 67 -554
rect -67 -634 -41 -608
rect -13 -634 13 -608
rect 41 -634 67 -608
rect -67 -688 -41 -662
rect -13 -688 13 -662
rect 41 -688 67 -662
rect -67 -742 -41 -716
rect -13 -742 13 -716
rect 41 -742 67 -716
rect -67 -796 -41 -770
rect -13 -796 13 -770
rect 41 -796 67 -770
rect -67 -850 -41 -824
rect -13 -850 13 -824
rect 41 -850 67 -824
rect -67 -904 -41 -878
rect -13 -904 13 -878
rect 41 -904 67 -878
rect -67 -958 -41 -932
rect -13 -958 13 -932
rect 41 -958 67 -932
rect -67 -1012 -41 -986
rect -13 -1012 13 -986
rect 41 -1012 67 -986
rect -67 -1066 -41 -1040
rect -13 -1066 13 -1040
rect 41 -1066 67 -1040
rect -67 -1120 -41 -1094
rect -13 -1120 13 -1094
rect 41 -1120 67 -1094
rect -67 -1174 -41 -1148
rect -13 -1174 13 -1148
rect 41 -1174 67 -1148
rect -67 -1228 -41 -1202
rect -13 -1228 13 -1202
rect 41 -1228 67 -1202
rect -67 -1282 -41 -1256
rect -13 -1282 13 -1256
rect 41 -1282 67 -1256
rect -67 -1336 -41 -1310
rect -13 -1336 13 -1310
rect 41 -1336 67 -1310
rect -67 -1390 -41 -1364
rect -13 -1390 13 -1364
rect 41 -1390 67 -1364
rect -67 -1444 -41 -1418
rect -13 -1444 13 -1418
rect 41 -1444 67 -1418
rect -67 -1498 -41 -1472
rect -13 -1498 13 -1472
rect 41 -1498 67 -1472
rect -67 -1552 -41 -1526
rect -13 -1552 13 -1526
rect 41 -1552 67 -1526
rect -67 -1606 -41 -1580
rect -13 -1606 13 -1580
rect 41 -1606 67 -1580
rect -67 -1660 -41 -1634
rect -13 -1660 13 -1634
rect 41 -1660 67 -1634
rect -67 -1714 -41 -1688
rect -13 -1714 13 -1688
rect 41 -1714 67 -1688
rect -67 -1768 -41 -1742
rect -13 -1768 13 -1742
rect 41 -1768 67 -1742
rect -67 -1822 -41 -1796
rect -13 -1822 13 -1796
rect 41 -1822 67 -1796
rect -67 -1876 -41 -1850
rect -13 -1876 13 -1850
rect 41 -1876 67 -1850
rect -67 -1930 -41 -1904
rect -13 -1930 13 -1904
rect 41 -1930 67 -1904
rect -67 -1984 -41 -1958
rect -13 -1984 13 -1958
rect 41 -1984 67 -1958
rect -67 -2038 -41 -2012
rect -13 -2038 13 -2012
rect 41 -2038 67 -2012
rect -67 -2092 -41 -2066
rect -13 -2092 13 -2066
rect 41 -2092 67 -2066
rect -67 -2146 -41 -2120
rect -13 -2146 13 -2120
rect 41 -2146 67 -2120
rect -67 -2200 -41 -2174
rect -13 -2200 13 -2174
rect 41 -2200 67 -2174
rect -67 -2254 -41 -2228
rect -13 -2254 13 -2228
rect 41 -2254 67 -2228
rect -67 -2308 -41 -2282
rect -13 -2308 13 -2282
rect 41 -2308 67 -2282
rect -67 -2362 -41 -2336
rect -13 -2362 13 -2336
rect 41 -2362 67 -2336
rect -67 -2416 -41 -2390
rect -13 -2416 13 -2390
rect 41 -2416 67 -2390
rect -67 -2470 -41 -2444
rect -13 -2470 13 -2444
rect 41 -2470 67 -2444
rect -67 -2524 -41 -2498
rect -13 -2524 13 -2498
rect 41 -2524 67 -2498
rect -67 -2578 -41 -2552
rect -13 -2578 13 -2552
rect 41 -2578 67 -2552
rect -67 -2632 -41 -2606
rect -13 -2632 13 -2606
rect 41 -2632 67 -2606
rect -67 -2686 -41 -2660
rect -13 -2686 13 -2660
rect 41 -2686 67 -2660
rect -67 -2740 -41 -2714
rect -13 -2740 13 -2714
rect 41 -2740 67 -2714
rect -67 -2794 -41 -2768
rect -13 -2794 13 -2768
rect 41 -2794 67 -2768
rect -67 -2848 -41 -2822
rect -13 -2848 13 -2822
rect 41 -2848 67 -2822
rect -67 -2902 -41 -2876
rect -13 -2902 13 -2876
rect 41 -2902 67 -2876
rect -67 -2956 -41 -2930
rect -13 -2956 13 -2930
rect 41 -2956 67 -2930
rect -67 -3010 -41 -2984
rect -13 -3010 13 -2984
rect 41 -3010 67 -2984
rect -67 -3064 -41 -3038
rect -13 -3064 13 -3038
rect 41 -3064 67 -3038
rect -67 -3118 -41 -3092
rect -13 -3118 13 -3092
rect 41 -3118 67 -3092
rect -67 -3172 -41 -3146
rect -13 -3172 13 -3146
rect 41 -3172 67 -3146
rect -67 -3226 -41 -3200
rect -13 -3226 13 -3200
rect 41 -3226 67 -3200
rect -67 -3280 -41 -3254
rect -13 -3280 13 -3254
rect 41 -3280 67 -3254
rect -67 -3334 -41 -3308
rect -13 -3334 13 -3308
rect 41 -3334 67 -3308
rect -67 -3388 -41 -3362
rect -13 -3388 13 -3362
rect 41 -3388 67 -3362
rect -67 -3442 -41 -3416
rect -13 -3442 13 -3416
rect 41 -3442 67 -3416
rect -67 -3496 -41 -3470
rect -13 -3496 13 -3470
rect 41 -3496 67 -3470
rect -67 -3550 -41 -3524
rect -13 -3550 13 -3524
rect 41 -3550 67 -3524
rect -67 -3604 -41 -3578
rect -13 -3604 13 -3578
rect 41 -3604 67 -3578
rect -67 -3658 -41 -3632
rect -13 -3658 13 -3632
rect 41 -3658 67 -3632
rect -67 -3712 -41 -3686
rect -13 -3712 13 -3686
rect 41 -3712 67 -3686
rect -67 -3766 -41 -3740
rect -13 -3766 13 -3740
rect 41 -3766 67 -3740
rect -67 -3820 -41 -3794
rect -13 -3820 13 -3794
rect 41 -3820 67 -3794
rect -67 -3874 -41 -3848
rect -13 -3874 13 -3848
rect 41 -3874 67 -3848
rect -67 -3928 -41 -3902
rect -13 -3928 13 -3902
rect 41 -3928 67 -3902
rect -67 -3982 -41 -3956
rect -13 -3982 13 -3956
rect 41 -3982 67 -3956
rect -67 -4036 -41 -4010
rect -13 -4036 13 -4010
rect 41 -4036 67 -4010
rect -67 -4090 -41 -4064
rect -13 -4090 13 -4064
rect 41 -4090 67 -4064
rect -67 -4144 -41 -4118
rect -13 -4144 13 -4118
rect 41 -4144 67 -4118
rect -67 -4198 -41 -4172
rect -13 -4198 13 -4172
rect 41 -4198 67 -4172
rect -67 -4252 -41 -4226
rect -13 -4252 13 -4226
rect 41 -4252 67 -4226
rect -67 -4306 -41 -4280
rect -13 -4306 13 -4280
rect 41 -4306 67 -4280
rect -67 -4360 -41 -4334
rect -13 -4360 13 -4334
rect 41 -4360 67 -4334
rect -67 -4414 -41 -4388
rect -13 -4414 13 -4388
rect 41 -4414 67 -4388
rect -67 -4468 -41 -4442
rect -13 -4468 13 -4442
rect 41 -4468 67 -4442
rect -67 -4522 -41 -4496
rect -13 -4522 13 -4496
rect 41 -4522 67 -4496
rect -67 -4576 -41 -4550
rect -13 -4576 13 -4550
rect 41 -4576 67 -4550
rect -67 -4630 -41 -4604
rect -13 -4630 13 -4604
rect 41 -4630 67 -4604
rect -67 -4684 -41 -4658
rect -13 -4684 13 -4658
rect 41 -4684 67 -4658
rect -67 -4738 -41 -4712
rect -13 -4738 13 -4712
rect 41 -4738 67 -4712
rect -67 -4792 -41 -4766
rect -13 -4792 13 -4766
rect 41 -4792 67 -4766
rect -67 -4846 -41 -4820
rect -13 -4846 13 -4820
rect 41 -4846 67 -4820
rect -67 -4900 -41 -4874
rect -13 -4900 13 -4874
rect 41 -4900 67 -4874
rect -67 -4954 -41 -4928
rect -13 -4954 13 -4928
rect 41 -4954 67 -4928
rect -67 -5008 -41 -4982
rect -13 -5008 13 -4982
rect 41 -5008 67 -4982
rect -67 -5062 -41 -5036
rect -13 -5062 13 -5036
rect 41 -5062 67 -5036
rect -67 -5116 -41 -5090
rect -13 -5116 13 -5090
rect 41 -5116 67 -5090
rect -67 -5170 -41 -5144
rect -13 -5170 13 -5144
rect 41 -5170 67 -5144
rect -67 -5224 -41 -5198
rect -13 -5224 13 -5198
rect 41 -5224 67 -5198
rect -67 -5278 -41 -5252
rect -13 -5278 13 -5252
rect 41 -5278 67 -5252
rect -67 -5332 -41 -5306
rect -13 -5332 13 -5306
rect 41 -5332 67 -5306
rect -67 -5386 -41 -5360
rect -13 -5386 13 -5360
rect 41 -5386 67 -5360
rect -67 -5440 -41 -5414
rect -13 -5440 13 -5414
rect 41 -5440 67 -5414
rect -67 -5494 -41 -5468
rect -13 -5494 13 -5468
rect 41 -5494 67 -5468
rect -67 -5548 -41 -5522
rect -13 -5548 13 -5522
rect 41 -5548 67 -5522
rect -67 -5602 -41 -5576
rect -13 -5602 13 -5576
rect 41 -5602 67 -5576
rect -67 -5656 -41 -5630
rect -13 -5656 13 -5630
rect 41 -5656 67 -5630
rect -67 -5710 -41 -5684
rect -13 -5710 13 -5684
rect 41 -5710 67 -5684
rect -67 -5764 -41 -5738
rect -13 -5764 13 -5738
rect 41 -5764 67 -5738
rect -67 -5818 -41 -5792
rect -13 -5818 13 -5792
rect 41 -5818 67 -5792
rect -67 -5872 -41 -5846
rect -13 -5872 13 -5846
rect 41 -5872 67 -5846
rect -67 -5926 -41 -5900
rect -13 -5926 13 -5900
rect 41 -5926 67 -5900
rect -67 -5980 -41 -5954
rect -13 -5980 13 -5954
rect 41 -5980 67 -5954
rect -67 -6034 -41 -6008
rect -13 -6034 13 -6008
rect 41 -6034 67 -6008
rect -67 -6088 -41 -6062
rect -13 -6088 13 -6062
rect 41 -6088 67 -6062
rect -67 -6142 -41 -6116
rect -13 -6142 13 -6116
rect 41 -6142 67 -6116
rect -67 -6196 -41 -6170
rect -13 -6196 13 -6170
rect 41 -6196 67 -6170
rect -67 -6250 -41 -6224
rect -13 -6250 13 -6224
rect 41 -6250 67 -6224
rect -67 -6304 -41 -6278
rect -13 -6304 13 -6278
rect 41 -6304 67 -6278
<< metal2 >>
rect -73 6304 73 6310
rect -73 6278 -67 6304
rect -41 6278 -13 6304
rect 13 6278 41 6304
rect 67 6278 73 6304
rect -73 6250 73 6278
rect -73 6224 -67 6250
rect -41 6224 -13 6250
rect 13 6224 41 6250
rect 67 6224 73 6250
rect -73 6196 73 6224
rect -73 6170 -67 6196
rect -41 6170 -13 6196
rect 13 6170 41 6196
rect 67 6170 73 6196
rect -73 6142 73 6170
rect -73 6116 -67 6142
rect -41 6116 -13 6142
rect 13 6116 41 6142
rect 67 6116 73 6142
rect -73 6088 73 6116
rect -73 6062 -67 6088
rect -41 6062 -13 6088
rect 13 6062 41 6088
rect 67 6062 73 6088
rect -73 6034 73 6062
rect -73 6008 -67 6034
rect -41 6008 -13 6034
rect 13 6008 41 6034
rect 67 6008 73 6034
rect -73 5980 73 6008
rect -73 5954 -67 5980
rect -41 5954 -13 5980
rect 13 5954 41 5980
rect 67 5954 73 5980
rect -73 5926 73 5954
rect -73 5900 -67 5926
rect -41 5900 -13 5926
rect 13 5900 41 5926
rect 67 5900 73 5926
rect -73 5872 73 5900
rect -73 5846 -67 5872
rect -41 5846 -13 5872
rect 13 5846 41 5872
rect 67 5846 73 5872
rect -73 5818 73 5846
rect -73 5792 -67 5818
rect -41 5792 -13 5818
rect 13 5792 41 5818
rect 67 5792 73 5818
rect -73 5764 73 5792
rect -73 5738 -67 5764
rect -41 5738 -13 5764
rect 13 5738 41 5764
rect 67 5738 73 5764
rect -73 5710 73 5738
rect -73 5684 -67 5710
rect -41 5684 -13 5710
rect 13 5684 41 5710
rect 67 5684 73 5710
rect -73 5656 73 5684
rect -73 5630 -67 5656
rect -41 5630 -13 5656
rect 13 5630 41 5656
rect 67 5630 73 5656
rect -73 5602 73 5630
rect -73 5576 -67 5602
rect -41 5576 -13 5602
rect 13 5576 41 5602
rect 67 5576 73 5602
rect -73 5548 73 5576
rect -73 5522 -67 5548
rect -41 5522 -13 5548
rect 13 5522 41 5548
rect 67 5522 73 5548
rect -73 5494 73 5522
rect -73 5468 -67 5494
rect -41 5468 -13 5494
rect 13 5468 41 5494
rect 67 5468 73 5494
rect -73 5440 73 5468
rect -73 5414 -67 5440
rect -41 5414 -13 5440
rect 13 5414 41 5440
rect 67 5414 73 5440
rect -73 5386 73 5414
rect -73 5360 -67 5386
rect -41 5360 -13 5386
rect 13 5360 41 5386
rect 67 5360 73 5386
rect -73 5332 73 5360
rect -73 5306 -67 5332
rect -41 5306 -13 5332
rect 13 5306 41 5332
rect 67 5306 73 5332
rect -73 5278 73 5306
rect -73 5252 -67 5278
rect -41 5252 -13 5278
rect 13 5252 41 5278
rect 67 5252 73 5278
rect -73 5224 73 5252
rect -73 5198 -67 5224
rect -41 5198 -13 5224
rect 13 5198 41 5224
rect 67 5198 73 5224
rect -73 5170 73 5198
rect -73 5144 -67 5170
rect -41 5144 -13 5170
rect 13 5144 41 5170
rect 67 5144 73 5170
rect -73 5116 73 5144
rect -73 5090 -67 5116
rect -41 5090 -13 5116
rect 13 5090 41 5116
rect 67 5090 73 5116
rect -73 5062 73 5090
rect -73 5036 -67 5062
rect -41 5036 -13 5062
rect 13 5036 41 5062
rect 67 5036 73 5062
rect -73 5008 73 5036
rect -73 4982 -67 5008
rect -41 4982 -13 5008
rect 13 4982 41 5008
rect 67 4982 73 5008
rect -73 4954 73 4982
rect -73 4928 -67 4954
rect -41 4928 -13 4954
rect 13 4928 41 4954
rect 67 4928 73 4954
rect -73 4900 73 4928
rect -73 4874 -67 4900
rect -41 4874 -13 4900
rect 13 4874 41 4900
rect 67 4874 73 4900
rect -73 4846 73 4874
rect -73 4820 -67 4846
rect -41 4820 -13 4846
rect 13 4820 41 4846
rect 67 4820 73 4846
rect -73 4792 73 4820
rect -73 4766 -67 4792
rect -41 4766 -13 4792
rect 13 4766 41 4792
rect 67 4766 73 4792
rect -73 4738 73 4766
rect -73 4712 -67 4738
rect -41 4712 -13 4738
rect 13 4712 41 4738
rect 67 4712 73 4738
rect -73 4684 73 4712
rect -73 4658 -67 4684
rect -41 4658 -13 4684
rect 13 4658 41 4684
rect 67 4658 73 4684
rect -73 4630 73 4658
rect -73 4604 -67 4630
rect -41 4604 -13 4630
rect 13 4604 41 4630
rect 67 4604 73 4630
rect -73 4576 73 4604
rect -73 4550 -67 4576
rect -41 4550 -13 4576
rect 13 4550 41 4576
rect 67 4550 73 4576
rect -73 4522 73 4550
rect -73 4496 -67 4522
rect -41 4496 -13 4522
rect 13 4496 41 4522
rect 67 4496 73 4522
rect -73 4468 73 4496
rect -73 4442 -67 4468
rect -41 4442 -13 4468
rect 13 4442 41 4468
rect 67 4442 73 4468
rect -73 4414 73 4442
rect -73 4388 -67 4414
rect -41 4388 -13 4414
rect 13 4388 41 4414
rect 67 4388 73 4414
rect -73 4360 73 4388
rect -73 4334 -67 4360
rect -41 4334 -13 4360
rect 13 4334 41 4360
rect 67 4334 73 4360
rect -73 4306 73 4334
rect -73 4280 -67 4306
rect -41 4280 -13 4306
rect 13 4280 41 4306
rect 67 4280 73 4306
rect -73 4252 73 4280
rect -73 4226 -67 4252
rect -41 4226 -13 4252
rect 13 4226 41 4252
rect 67 4226 73 4252
rect -73 4198 73 4226
rect -73 4172 -67 4198
rect -41 4172 -13 4198
rect 13 4172 41 4198
rect 67 4172 73 4198
rect -73 4144 73 4172
rect -73 4118 -67 4144
rect -41 4118 -13 4144
rect 13 4118 41 4144
rect 67 4118 73 4144
rect -73 4090 73 4118
rect -73 4064 -67 4090
rect -41 4064 -13 4090
rect 13 4064 41 4090
rect 67 4064 73 4090
rect -73 4036 73 4064
rect -73 4010 -67 4036
rect -41 4010 -13 4036
rect 13 4010 41 4036
rect 67 4010 73 4036
rect -73 3982 73 4010
rect -73 3956 -67 3982
rect -41 3956 -13 3982
rect 13 3956 41 3982
rect 67 3956 73 3982
rect -73 3928 73 3956
rect -73 3902 -67 3928
rect -41 3902 -13 3928
rect 13 3902 41 3928
rect 67 3902 73 3928
rect -73 3874 73 3902
rect -73 3848 -67 3874
rect -41 3848 -13 3874
rect 13 3848 41 3874
rect 67 3848 73 3874
rect -73 3820 73 3848
rect -73 3794 -67 3820
rect -41 3794 -13 3820
rect 13 3794 41 3820
rect 67 3794 73 3820
rect -73 3766 73 3794
rect -73 3740 -67 3766
rect -41 3740 -13 3766
rect 13 3740 41 3766
rect 67 3740 73 3766
rect -73 3712 73 3740
rect -73 3686 -67 3712
rect -41 3686 -13 3712
rect 13 3686 41 3712
rect 67 3686 73 3712
rect -73 3658 73 3686
rect -73 3632 -67 3658
rect -41 3632 -13 3658
rect 13 3632 41 3658
rect 67 3632 73 3658
rect -73 3604 73 3632
rect -73 3578 -67 3604
rect -41 3578 -13 3604
rect 13 3578 41 3604
rect 67 3578 73 3604
rect -73 3550 73 3578
rect -73 3524 -67 3550
rect -41 3524 -13 3550
rect 13 3524 41 3550
rect 67 3524 73 3550
rect -73 3496 73 3524
rect -73 3470 -67 3496
rect -41 3470 -13 3496
rect 13 3470 41 3496
rect 67 3470 73 3496
rect -73 3442 73 3470
rect -73 3416 -67 3442
rect -41 3416 -13 3442
rect 13 3416 41 3442
rect 67 3416 73 3442
rect -73 3388 73 3416
rect -73 3362 -67 3388
rect -41 3362 -13 3388
rect 13 3362 41 3388
rect 67 3362 73 3388
rect -73 3334 73 3362
rect -73 3308 -67 3334
rect -41 3308 -13 3334
rect 13 3308 41 3334
rect 67 3308 73 3334
rect -73 3280 73 3308
rect -73 3254 -67 3280
rect -41 3254 -13 3280
rect 13 3254 41 3280
rect 67 3254 73 3280
rect -73 3226 73 3254
rect -73 3200 -67 3226
rect -41 3200 -13 3226
rect 13 3200 41 3226
rect 67 3200 73 3226
rect -73 3172 73 3200
rect -73 3146 -67 3172
rect -41 3146 -13 3172
rect 13 3146 41 3172
rect 67 3146 73 3172
rect -73 3118 73 3146
rect -73 3092 -67 3118
rect -41 3092 -13 3118
rect 13 3092 41 3118
rect 67 3092 73 3118
rect -73 3064 73 3092
rect -73 3038 -67 3064
rect -41 3038 -13 3064
rect 13 3038 41 3064
rect 67 3038 73 3064
rect -73 3010 73 3038
rect -73 2984 -67 3010
rect -41 2984 -13 3010
rect 13 2984 41 3010
rect 67 2984 73 3010
rect -73 2956 73 2984
rect -73 2930 -67 2956
rect -41 2930 -13 2956
rect 13 2930 41 2956
rect 67 2930 73 2956
rect -73 2902 73 2930
rect -73 2876 -67 2902
rect -41 2876 -13 2902
rect 13 2876 41 2902
rect 67 2876 73 2902
rect -73 2848 73 2876
rect -73 2822 -67 2848
rect -41 2822 -13 2848
rect 13 2822 41 2848
rect 67 2822 73 2848
rect -73 2794 73 2822
rect -73 2768 -67 2794
rect -41 2768 -13 2794
rect 13 2768 41 2794
rect 67 2768 73 2794
rect -73 2740 73 2768
rect -73 2714 -67 2740
rect -41 2714 -13 2740
rect 13 2714 41 2740
rect 67 2714 73 2740
rect -73 2686 73 2714
rect -73 2660 -67 2686
rect -41 2660 -13 2686
rect 13 2660 41 2686
rect 67 2660 73 2686
rect -73 2632 73 2660
rect -73 2606 -67 2632
rect -41 2606 -13 2632
rect 13 2606 41 2632
rect 67 2606 73 2632
rect -73 2578 73 2606
rect -73 2552 -67 2578
rect -41 2552 -13 2578
rect 13 2552 41 2578
rect 67 2552 73 2578
rect -73 2524 73 2552
rect -73 2498 -67 2524
rect -41 2498 -13 2524
rect 13 2498 41 2524
rect 67 2498 73 2524
rect -73 2470 73 2498
rect -73 2444 -67 2470
rect -41 2444 -13 2470
rect 13 2444 41 2470
rect 67 2444 73 2470
rect -73 2416 73 2444
rect -73 2390 -67 2416
rect -41 2390 -13 2416
rect 13 2390 41 2416
rect 67 2390 73 2416
rect -73 2362 73 2390
rect -73 2336 -67 2362
rect -41 2336 -13 2362
rect 13 2336 41 2362
rect 67 2336 73 2362
rect -73 2308 73 2336
rect -73 2282 -67 2308
rect -41 2282 -13 2308
rect 13 2282 41 2308
rect 67 2282 73 2308
rect -73 2254 73 2282
rect -73 2228 -67 2254
rect -41 2228 -13 2254
rect 13 2228 41 2254
rect 67 2228 73 2254
rect -73 2200 73 2228
rect -73 2174 -67 2200
rect -41 2174 -13 2200
rect 13 2174 41 2200
rect 67 2174 73 2200
rect -73 2146 73 2174
rect -73 2120 -67 2146
rect -41 2120 -13 2146
rect 13 2120 41 2146
rect 67 2120 73 2146
rect -73 2092 73 2120
rect -73 2066 -67 2092
rect -41 2066 -13 2092
rect 13 2066 41 2092
rect 67 2066 73 2092
rect -73 2038 73 2066
rect -73 2012 -67 2038
rect -41 2012 -13 2038
rect 13 2012 41 2038
rect 67 2012 73 2038
rect -73 1984 73 2012
rect -73 1958 -67 1984
rect -41 1958 -13 1984
rect 13 1958 41 1984
rect 67 1958 73 1984
rect -73 1930 73 1958
rect -73 1904 -67 1930
rect -41 1904 -13 1930
rect 13 1904 41 1930
rect 67 1904 73 1930
rect -73 1876 73 1904
rect -73 1850 -67 1876
rect -41 1850 -13 1876
rect 13 1850 41 1876
rect 67 1850 73 1876
rect -73 1822 73 1850
rect -73 1796 -67 1822
rect -41 1796 -13 1822
rect 13 1796 41 1822
rect 67 1796 73 1822
rect -73 1768 73 1796
rect -73 1742 -67 1768
rect -41 1742 -13 1768
rect 13 1742 41 1768
rect 67 1742 73 1768
rect -73 1714 73 1742
rect -73 1688 -67 1714
rect -41 1688 -13 1714
rect 13 1688 41 1714
rect 67 1688 73 1714
rect -73 1660 73 1688
rect -73 1634 -67 1660
rect -41 1634 -13 1660
rect 13 1634 41 1660
rect 67 1634 73 1660
rect -73 1606 73 1634
rect -73 1580 -67 1606
rect -41 1580 -13 1606
rect 13 1580 41 1606
rect 67 1580 73 1606
rect -73 1552 73 1580
rect -73 1526 -67 1552
rect -41 1526 -13 1552
rect 13 1526 41 1552
rect 67 1526 73 1552
rect -73 1498 73 1526
rect -73 1472 -67 1498
rect -41 1472 -13 1498
rect 13 1472 41 1498
rect 67 1472 73 1498
rect -73 1444 73 1472
rect -73 1418 -67 1444
rect -41 1418 -13 1444
rect 13 1418 41 1444
rect 67 1418 73 1444
rect -73 1390 73 1418
rect -73 1364 -67 1390
rect -41 1364 -13 1390
rect 13 1364 41 1390
rect 67 1364 73 1390
rect -73 1336 73 1364
rect -73 1310 -67 1336
rect -41 1310 -13 1336
rect 13 1310 41 1336
rect 67 1310 73 1336
rect -73 1282 73 1310
rect -73 1256 -67 1282
rect -41 1256 -13 1282
rect 13 1256 41 1282
rect 67 1256 73 1282
rect -73 1228 73 1256
rect -73 1202 -67 1228
rect -41 1202 -13 1228
rect 13 1202 41 1228
rect 67 1202 73 1228
rect -73 1174 73 1202
rect -73 1148 -67 1174
rect -41 1148 -13 1174
rect 13 1148 41 1174
rect 67 1148 73 1174
rect -73 1120 73 1148
rect -73 1094 -67 1120
rect -41 1094 -13 1120
rect 13 1094 41 1120
rect 67 1094 73 1120
rect -73 1066 73 1094
rect -73 1040 -67 1066
rect -41 1040 -13 1066
rect 13 1040 41 1066
rect 67 1040 73 1066
rect -73 1012 73 1040
rect -73 986 -67 1012
rect -41 986 -13 1012
rect 13 986 41 1012
rect 67 986 73 1012
rect -73 958 73 986
rect -73 932 -67 958
rect -41 932 -13 958
rect 13 932 41 958
rect 67 932 73 958
rect -73 904 73 932
rect -73 878 -67 904
rect -41 878 -13 904
rect 13 878 41 904
rect 67 878 73 904
rect -73 850 73 878
rect -73 824 -67 850
rect -41 824 -13 850
rect 13 824 41 850
rect 67 824 73 850
rect -73 796 73 824
rect -73 770 -67 796
rect -41 770 -13 796
rect 13 770 41 796
rect 67 770 73 796
rect -73 742 73 770
rect -73 716 -67 742
rect -41 716 -13 742
rect 13 716 41 742
rect 67 716 73 742
rect -73 688 73 716
rect -73 662 -67 688
rect -41 662 -13 688
rect 13 662 41 688
rect 67 662 73 688
rect -73 634 73 662
rect -73 608 -67 634
rect -41 608 -13 634
rect 13 608 41 634
rect 67 608 73 634
rect -73 580 73 608
rect -73 554 -67 580
rect -41 554 -13 580
rect 13 554 41 580
rect 67 554 73 580
rect -73 526 73 554
rect -73 500 -67 526
rect -41 500 -13 526
rect 13 500 41 526
rect 67 500 73 526
rect -73 472 73 500
rect -73 446 -67 472
rect -41 446 -13 472
rect 13 446 41 472
rect 67 446 73 472
rect -73 418 73 446
rect -73 392 -67 418
rect -41 392 -13 418
rect 13 392 41 418
rect 67 392 73 418
rect -73 364 73 392
rect -73 338 -67 364
rect -41 338 -13 364
rect 13 338 41 364
rect 67 338 73 364
rect -73 310 73 338
rect -73 284 -67 310
rect -41 284 -13 310
rect 13 284 41 310
rect 67 284 73 310
rect -73 256 73 284
rect -73 230 -67 256
rect -41 230 -13 256
rect 13 230 41 256
rect 67 230 73 256
rect -73 202 73 230
rect -73 176 -67 202
rect -41 176 -13 202
rect 13 176 41 202
rect 67 176 73 202
rect -73 148 73 176
rect -73 122 -67 148
rect -41 122 -13 148
rect 13 122 41 148
rect 67 122 73 148
rect -73 94 73 122
rect -73 68 -67 94
rect -41 68 -13 94
rect 13 68 41 94
rect 67 68 73 94
rect -73 40 73 68
rect -73 14 -67 40
rect -41 14 -13 40
rect 13 14 41 40
rect 67 14 73 40
rect -73 -14 73 14
rect -73 -40 -67 -14
rect -41 -40 -13 -14
rect 13 -40 41 -14
rect 67 -40 73 -14
rect -73 -68 73 -40
rect -73 -94 -67 -68
rect -41 -94 -13 -68
rect 13 -94 41 -68
rect 67 -94 73 -68
rect -73 -122 73 -94
rect -73 -148 -67 -122
rect -41 -148 -13 -122
rect 13 -148 41 -122
rect 67 -148 73 -122
rect -73 -176 73 -148
rect -73 -202 -67 -176
rect -41 -202 -13 -176
rect 13 -202 41 -176
rect 67 -202 73 -176
rect -73 -230 73 -202
rect -73 -256 -67 -230
rect -41 -256 -13 -230
rect 13 -256 41 -230
rect 67 -256 73 -230
rect -73 -284 73 -256
rect -73 -310 -67 -284
rect -41 -310 -13 -284
rect 13 -310 41 -284
rect 67 -310 73 -284
rect -73 -338 73 -310
rect -73 -364 -67 -338
rect -41 -364 -13 -338
rect 13 -364 41 -338
rect 67 -364 73 -338
rect -73 -392 73 -364
rect -73 -418 -67 -392
rect -41 -418 -13 -392
rect 13 -418 41 -392
rect 67 -418 73 -392
rect -73 -446 73 -418
rect -73 -472 -67 -446
rect -41 -472 -13 -446
rect 13 -472 41 -446
rect 67 -472 73 -446
rect -73 -500 73 -472
rect -73 -526 -67 -500
rect -41 -526 -13 -500
rect 13 -526 41 -500
rect 67 -526 73 -500
rect -73 -554 73 -526
rect -73 -580 -67 -554
rect -41 -580 -13 -554
rect 13 -580 41 -554
rect 67 -580 73 -554
rect -73 -608 73 -580
rect -73 -634 -67 -608
rect -41 -634 -13 -608
rect 13 -634 41 -608
rect 67 -634 73 -608
rect -73 -662 73 -634
rect -73 -688 -67 -662
rect -41 -688 -13 -662
rect 13 -688 41 -662
rect 67 -688 73 -662
rect -73 -716 73 -688
rect -73 -742 -67 -716
rect -41 -742 -13 -716
rect 13 -742 41 -716
rect 67 -742 73 -716
rect -73 -770 73 -742
rect -73 -796 -67 -770
rect -41 -796 -13 -770
rect 13 -796 41 -770
rect 67 -796 73 -770
rect -73 -824 73 -796
rect -73 -850 -67 -824
rect -41 -850 -13 -824
rect 13 -850 41 -824
rect 67 -850 73 -824
rect -73 -878 73 -850
rect -73 -904 -67 -878
rect -41 -904 -13 -878
rect 13 -904 41 -878
rect 67 -904 73 -878
rect -73 -932 73 -904
rect -73 -958 -67 -932
rect -41 -958 -13 -932
rect 13 -958 41 -932
rect 67 -958 73 -932
rect -73 -986 73 -958
rect -73 -1012 -67 -986
rect -41 -1012 -13 -986
rect 13 -1012 41 -986
rect 67 -1012 73 -986
rect -73 -1040 73 -1012
rect -73 -1066 -67 -1040
rect -41 -1066 -13 -1040
rect 13 -1066 41 -1040
rect 67 -1066 73 -1040
rect -73 -1094 73 -1066
rect -73 -1120 -67 -1094
rect -41 -1120 -13 -1094
rect 13 -1120 41 -1094
rect 67 -1120 73 -1094
rect -73 -1148 73 -1120
rect -73 -1174 -67 -1148
rect -41 -1174 -13 -1148
rect 13 -1174 41 -1148
rect 67 -1174 73 -1148
rect -73 -1202 73 -1174
rect -73 -1228 -67 -1202
rect -41 -1228 -13 -1202
rect 13 -1228 41 -1202
rect 67 -1228 73 -1202
rect -73 -1256 73 -1228
rect -73 -1282 -67 -1256
rect -41 -1282 -13 -1256
rect 13 -1282 41 -1256
rect 67 -1282 73 -1256
rect -73 -1310 73 -1282
rect -73 -1336 -67 -1310
rect -41 -1336 -13 -1310
rect 13 -1336 41 -1310
rect 67 -1336 73 -1310
rect -73 -1364 73 -1336
rect -73 -1390 -67 -1364
rect -41 -1390 -13 -1364
rect 13 -1390 41 -1364
rect 67 -1390 73 -1364
rect -73 -1418 73 -1390
rect -73 -1444 -67 -1418
rect -41 -1444 -13 -1418
rect 13 -1444 41 -1418
rect 67 -1444 73 -1418
rect -73 -1472 73 -1444
rect -73 -1498 -67 -1472
rect -41 -1498 -13 -1472
rect 13 -1498 41 -1472
rect 67 -1498 73 -1472
rect -73 -1526 73 -1498
rect -73 -1552 -67 -1526
rect -41 -1552 -13 -1526
rect 13 -1552 41 -1526
rect 67 -1552 73 -1526
rect -73 -1580 73 -1552
rect -73 -1606 -67 -1580
rect -41 -1606 -13 -1580
rect 13 -1606 41 -1580
rect 67 -1606 73 -1580
rect -73 -1634 73 -1606
rect -73 -1660 -67 -1634
rect -41 -1660 -13 -1634
rect 13 -1660 41 -1634
rect 67 -1660 73 -1634
rect -73 -1688 73 -1660
rect -73 -1714 -67 -1688
rect -41 -1714 -13 -1688
rect 13 -1714 41 -1688
rect 67 -1714 73 -1688
rect -73 -1742 73 -1714
rect -73 -1768 -67 -1742
rect -41 -1768 -13 -1742
rect 13 -1768 41 -1742
rect 67 -1768 73 -1742
rect -73 -1796 73 -1768
rect -73 -1822 -67 -1796
rect -41 -1822 -13 -1796
rect 13 -1822 41 -1796
rect 67 -1822 73 -1796
rect -73 -1850 73 -1822
rect -73 -1876 -67 -1850
rect -41 -1876 -13 -1850
rect 13 -1876 41 -1850
rect 67 -1876 73 -1850
rect -73 -1904 73 -1876
rect -73 -1930 -67 -1904
rect -41 -1930 -13 -1904
rect 13 -1930 41 -1904
rect 67 -1930 73 -1904
rect -73 -1958 73 -1930
rect -73 -1984 -67 -1958
rect -41 -1984 -13 -1958
rect 13 -1984 41 -1958
rect 67 -1984 73 -1958
rect -73 -2012 73 -1984
rect -73 -2038 -67 -2012
rect -41 -2038 -13 -2012
rect 13 -2038 41 -2012
rect 67 -2038 73 -2012
rect -73 -2066 73 -2038
rect -73 -2092 -67 -2066
rect -41 -2092 -13 -2066
rect 13 -2092 41 -2066
rect 67 -2092 73 -2066
rect -73 -2120 73 -2092
rect -73 -2146 -67 -2120
rect -41 -2146 -13 -2120
rect 13 -2146 41 -2120
rect 67 -2146 73 -2120
rect -73 -2174 73 -2146
rect -73 -2200 -67 -2174
rect -41 -2200 -13 -2174
rect 13 -2200 41 -2174
rect 67 -2200 73 -2174
rect -73 -2228 73 -2200
rect -73 -2254 -67 -2228
rect -41 -2254 -13 -2228
rect 13 -2254 41 -2228
rect 67 -2254 73 -2228
rect -73 -2282 73 -2254
rect -73 -2308 -67 -2282
rect -41 -2308 -13 -2282
rect 13 -2308 41 -2282
rect 67 -2308 73 -2282
rect -73 -2336 73 -2308
rect -73 -2362 -67 -2336
rect -41 -2362 -13 -2336
rect 13 -2362 41 -2336
rect 67 -2362 73 -2336
rect -73 -2390 73 -2362
rect -73 -2416 -67 -2390
rect -41 -2416 -13 -2390
rect 13 -2416 41 -2390
rect 67 -2416 73 -2390
rect -73 -2444 73 -2416
rect -73 -2470 -67 -2444
rect -41 -2470 -13 -2444
rect 13 -2470 41 -2444
rect 67 -2470 73 -2444
rect -73 -2498 73 -2470
rect -73 -2524 -67 -2498
rect -41 -2524 -13 -2498
rect 13 -2524 41 -2498
rect 67 -2524 73 -2498
rect -73 -2552 73 -2524
rect -73 -2578 -67 -2552
rect -41 -2578 -13 -2552
rect 13 -2578 41 -2552
rect 67 -2578 73 -2552
rect -73 -2606 73 -2578
rect -73 -2632 -67 -2606
rect -41 -2632 -13 -2606
rect 13 -2632 41 -2606
rect 67 -2632 73 -2606
rect -73 -2660 73 -2632
rect -73 -2686 -67 -2660
rect -41 -2686 -13 -2660
rect 13 -2686 41 -2660
rect 67 -2686 73 -2660
rect -73 -2714 73 -2686
rect -73 -2740 -67 -2714
rect -41 -2740 -13 -2714
rect 13 -2740 41 -2714
rect 67 -2740 73 -2714
rect -73 -2768 73 -2740
rect -73 -2794 -67 -2768
rect -41 -2794 -13 -2768
rect 13 -2794 41 -2768
rect 67 -2794 73 -2768
rect -73 -2822 73 -2794
rect -73 -2848 -67 -2822
rect -41 -2848 -13 -2822
rect 13 -2848 41 -2822
rect 67 -2848 73 -2822
rect -73 -2876 73 -2848
rect -73 -2902 -67 -2876
rect -41 -2902 -13 -2876
rect 13 -2902 41 -2876
rect 67 -2902 73 -2876
rect -73 -2930 73 -2902
rect -73 -2956 -67 -2930
rect -41 -2956 -13 -2930
rect 13 -2956 41 -2930
rect 67 -2956 73 -2930
rect -73 -2984 73 -2956
rect -73 -3010 -67 -2984
rect -41 -3010 -13 -2984
rect 13 -3010 41 -2984
rect 67 -3010 73 -2984
rect -73 -3038 73 -3010
rect -73 -3064 -67 -3038
rect -41 -3064 -13 -3038
rect 13 -3064 41 -3038
rect 67 -3064 73 -3038
rect -73 -3092 73 -3064
rect -73 -3118 -67 -3092
rect -41 -3118 -13 -3092
rect 13 -3118 41 -3092
rect 67 -3118 73 -3092
rect -73 -3146 73 -3118
rect -73 -3172 -67 -3146
rect -41 -3172 -13 -3146
rect 13 -3172 41 -3146
rect 67 -3172 73 -3146
rect -73 -3200 73 -3172
rect -73 -3226 -67 -3200
rect -41 -3226 -13 -3200
rect 13 -3226 41 -3200
rect 67 -3226 73 -3200
rect -73 -3254 73 -3226
rect -73 -3280 -67 -3254
rect -41 -3280 -13 -3254
rect 13 -3280 41 -3254
rect 67 -3280 73 -3254
rect -73 -3308 73 -3280
rect -73 -3334 -67 -3308
rect -41 -3334 -13 -3308
rect 13 -3334 41 -3308
rect 67 -3334 73 -3308
rect -73 -3362 73 -3334
rect -73 -3388 -67 -3362
rect -41 -3388 -13 -3362
rect 13 -3388 41 -3362
rect 67 -3388 73 -3362
rect -73 -3416 73 -3388
rect -73 -3442 -67 -3416
rect -41 -3442 -13 -3416
rect 13 -3442 41 -3416
rect 67 -3442 73 -3416
rect -73 -3470 73 -3442
rect -73 -3496 -67 -3470
rect -41 -3496 -13 -3470
rect 13 -3496 41 -3470
rect 67 -3496 73 -3470
rect -73 -3524 73 -3496
rect -73 -3550 -67 -3524
rect -41 -3550 -13 -3524
rect 13 -3550 41 -3524
rect 67 -3550 73 -3524
rect -73 -3578 73 -3550
rect -73 -3604 -67 -3578
rect -41 -3604 -13 -3578
rect 13 -3604 41 -3578
rect 67 -3604 73 -3578
rect -73 -3632 73 -3604
rect -73 -3658 -67 -3632
rect -41 -3658 -13 -3632
rect 13 -3658 41 -3632
rect 67 -3658 73 -3632
rect -73 -3686 73 -3658
rect -73 -3712 -67 -3686
rect -41 -3712 -13 -3686
rect 13 -3712 41 -3686
rect 67 -3712 73 -3686
rect -73 -3740 73 -3712
rect -73 -3766 -67 -3740
rect -41 -3766 -13 -3740
rect 13 -3766 41 -3740
rect 67 -3766 73 -3740
rect -73 -3794 73 -3766
rect -73 -3820 -67 -3794
rect -41 -3820 -13 -3794
rect 13 -3820 41 -3794
rect 67 -3820 73 -3794
rect -73 -3848 73 -3820
rect -73 -3874 -67 -3848
rect -41 -3874 -13 -3848
rect 13 -3874 41 -3848
rect 67 -3874 73 -3848
rect -73 -3902 73 -3874
rect -73 -3928 -67 -3902
rect -41 -3928 -13 -3902
rect 13 -3928 41 -3902
rect 67 -3928 73 -3902
rect -73 -3956 73 -3928
rect -73 -3982 -67 -3956
rect -41 -3982 -13 -3956
rect 13 -3982 41 -3956
rect 67 -3982 73 -3956
rect -73 -4010 73 -3982
rect -73 -4036 -67 -4010
rect -41 -4036 -13 -4010
rect 13 -4036 41 -4010
rect 67 -4036 73 -4010
rect -73 -4064 73 -4036
rect -73 -4090 -67 -4064
rect -41 -4090 -13 -4064
rect 13 -4090 41 -4064
rect 67 -4090 73 -4064
rect -73 -4118 73 -4090
rect -73 -4144 -67 -4118
rect -41 -4144 -13 -4118
rect 13 -4144 41 -4118
rect 67 -4144 73 -4118
rect -73 -4172 73 -4144
rect -73 -4198 -67 -4172
rect -41 -4198 -13 -4172
rect 13 -4198 41 -4172
rect 67 -4198 73 -4172
rect -73 -4226 73 -4198
rect -73 -4252 -67 -4226
rect -41 -4252 -13 -4226
rect 13 -4252 41 -4226
rect 67 -4252 73 -4226
rect -73 -4280 73 -4252
rect -73 -4306 -67 -4280
rect -41 -4306 -13 -4280
rect 13 -4306 41 -4280
rect 67 -4306 73 -4280
rect -73 -4334 73 -4306
rect -73 -4360 -67 -4334
rect -41 -4360 -13 -4334
rect 13 -4360 41 -4334
rect 67 -4360 73 -4334
rect -73 -4388 73 -4360
rect -73 -4414 -67 -4388
rect -41 -4414 -13 -4388
rect 13 -4414 41 -4388
rect 67 -4414 73 -4388
rect -73 -4442 73 -4414
rect -73 -4468 -67 -4442
rect -41 -4468 -13 -4442
rect 13 -4468 41 -4442
rect 67 -4468 73 -4442
rect -73 -4496 73 -4468
rect -73 -4522 -67 -4496
rect -41 -4522 -13 -4496
rect 13 -4522 41 -4496
rect 67 -4522 73 -4496
rect -73 -4550 73 -4522
rect -73 -4576 -67 -4550
rect -41 -4576 -13 -4550
rect 13 -4576 41 -4550
rect 67 -4576 73 -4550
rect -73 -4604 73 -4576
rect -73 -4630 -67 -4604
rect -41 -4630 -13 -4604
rect 13 -4630 41 -4604
rect 67 -4630 73 -4604
rect -73 -4658 73 -4630
rect -73 -4684 -67 -4658
rect -41 -4684 -13 -4658
rect 13 -4684 41 -4658
rect 67 -4684 73 -4658
rect -73 -4712 73 -4684
rect -73 -4738 -67 -4712
rect -41 -4738 -13 -4712
rect 13 -4738 41 -4712
rect 67 -4738 73 -4712
rect -73 -4766 73 -4738
rect -73 -4792 -67 -4766
rect -41 -4792 -13 -4766
rect 13 -4792 41 -4766
rect 67 -4792 73 -4766
rect -73 -4820 73 -4792
rect -73 -4846 -67 -4820
rect -41 -4846 -13 -4820
rect 13 -4846 41 -4820
rect 67 -4846 73 -4820
rect -73 -4874 73 -4846
rect -73 -4900 -67 -4874
rect -41 -4900 -13 -4874
rect 13 -4900 41 -4874
rect 67 -4900 73 -4874
rect -73 -4928 73 -4900
rect -73 -4954 -67 -4928
rect -41 -4954 -13 -4928
rect 13 -4954 41 -4928
rect 67 -4954 73 -4928
rect -73 -4982 73 -4954
rect -73 -5008 -67 -4982
rect -41 -5008 -13 -4982
rect 13 -5008 41 -4982
rect 67 -5008 73 -4982
rect -73 -5036 73 -5008
rect -73 -5062 -67 -5036
rect -41 -5062 -13 -5036
rect 13 -5062 41 -5036
rect 67 -5062 73 -5036
rect -73 -5090 73 -5062
rect -73 -5116 -67 -5090
rect -41 -5116 -13 -5090
rect 13 -5116 41 -5090
rect 67 -5116 73 -5090
rect -73 -5144 73 -5116
rect -73 -5170 -67 -5144
rect -41 -5170 -13 -5144
rect 13 -5170 41 -5144
rect 67 -5170 73 -5144
rect -73 -5198 73 -5170
rect -73 -5224 -67 -5198
rect -41 -5224 -13 -5198
rect 13 -5224 41 -5198
rect 67 -5224 73 -5198
rect -73 -5252 73 -5224
rect -73 -5278 -67 -5252
rect -41 -5278 -13 -5252
rect 13 -5278 41 -5252
rect 67 -5278 73 -5252
rect -73 -5306 73 -5278
rect -73 -5332 -67 -5306
rect -41 -5332 -13 -5306
rect 13 -5332 41 -5306
rect 67 -5332 73 -5306
rect -73 -5360 73 -5332
rect -73 -5386 -67 -5360
rect -41 -5386 -13 -5360
rect 13 -5386 41 -5360
rect 67 -5386 73 -5360
rect -73 -5414 73 -5386
rect -73 -5440 -67 -5414
rect -41 -5440 -13 -5414
rect 13 -5440 41 -5414
rect 67 -5440 73 -5414
rect -73 -5468 73 -5440
rect -73 -5494 -67 -5468
rect -41 -5494 -13 -5468
rect 13 -5494 41 -5468
rect 67 -5494 73 -5468
rect -73 -5522 73 -5494
rect -73 -5548 -67 -5522
rect -41 -5548 -13 -5522
rect 13 -5548 41 -5522
rect 67 -5548 73 -5522
rect -73 -5576 73 -5548
rect -73 -5602 -67 -5576
rect -41 -5602 -13 -5576
rect 13 -5602 41 -5576
rect 67 -5602 73 -5576
rect -73 -5630 73 -5602
rect -73 -5656 -67 -5630
rect -41 -5656 -13 -5630
rect 13 -5656 41 -5630
rect 67 -5656 73 -5630
rect -73 -5684 73 -5656
rect -73 -5710 -67 -5684
rect -41 -5710 -13 -5684
rect 13 -5710 41 -5684
rect 67 -5710 73 -5684
rect -73 -5738 73 -5710
rect -73 -5764 -67 -5738
rect -41 -5764 -13 -5738
rect 13 -5764 41 -5738
rect 67 -5764 73 -5738
rect -73 -5792 73 -5764
rect -73 -5818 -67 -5792
rect -41 -5818 -13 -5792
rect 13 -5818 41 -5792
rect 67 -5818 73 -5792
rect -73 -5846 73 -5818
rect -73 -5872 -67 -5846
rect -41 -5872 -13 -5846
rect 13 -5872 41 -5846
rect 67 -5872 73 -5846
rect -73 -5900 73 -5872
rect -73 -5926 -67 -5900
rect -41 -5926 -13 -5900
rect 13 -5926 41 -5900
rect 67 -5926 73 -5900
rect -73 -5954 73 -5926
rect -73 -5980 -67 -5954
rect -41 -5980 -13 -5954
rect 13 -5980 41 -5954
rect 67 -5980 73 -5954
rect -73 -6008 73 -5980
rect -73 -6034 -67 -6008
rect -41 -6034 -13 -6008
rect 13 -6034 41 -6008
rect 67 -6034 73 -6008
rect -73 -6062 73 -6034
rect -73 -6088 -67 -6062
rect -41 -6088 -13 -6062
rect 13 -6088 41 -6062
rect 67 -6088 73 -6062
rect -73 -6116 73 -6088
rect -73 -6142 -67 -6116
rect -41 -6142 -13 -6116
rect 13 -6142 41 -6116
rect 67 -6142 73 -6116
rect -73 -6170 73 -6142
rect -73 -6196 -67 -6170
rect -41 -6196 -13 -6170
rect 13 -6196 41 -6170
rect 67 -6196 73 -6170
rect -73 -6224 73 -6196
rect -73 -6250 -67 -6224
rect -41 -6250 -13 -6224
rect 13 -6250 41 -6224
rect 67 -6250 73 -6224
rect -73 -6278 73 -6250
rect -73 -6304 -67 -6278
rect -41 -6304 -13 -6278
rect 13 -6304 41 -6278
rect 67 -6304 73 -6278
rect -73 -6310 73 -6304
<< end >>
