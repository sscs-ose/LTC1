magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1349 -2537 1349 2537
<< metal3 >>
rect -349 1532 349 1537
rect -349 1504 -344 1532
rect -316 1504 -278 1532
rect -250 1504 -212 1532
rect -184 1504 -146 1532
rect -118 1504 -80 1532
rect -52 1504 -14 1532
rect 14 1504 52 1532
rect 80 1504 118 1532
rect 146 1504 184 1532
rect 212 1504 250 1532
rect 278 1504 316 1532
rect 344 1504 349 1532
rect -349 1466 349 1504
rect -349 1438 -344 1466
rect -316 1438 -278 1466
rect -250 1438 -212 1466
rect -184 1438 -146 1466
rect -118 1438 -80 1466
rect -52 1438 -14 1466
rect 14 1438 52 1466
rect 80 1438 118 1466
rect 146 1438 184 1466
rect 212 1438 250 1466
rect 278 1438 316 1466
rect 344 1438 349 1466
rect -349 1400 349 1438
rect -349 1372 -344 1400
rect -316 1372 -278 1400
rect -250 1372 -212 1400
rect -184 1372 -146 1400
rect -118 1372 -80 1400
rect -52 1372 -14 1400
rect 14 1372 52 1400
rect 80 1372 118 1400
rect 146 1372 184 1400
rect 212 1372 250 1400
rect 278 1372 316 1400
rect 344 1372 349 1400
rect -349 1334 349 1372
rect -349 1306 -344 1334
rect -316 1306 -278 1334
rect -250 1306 -212 1334
rect -184 1306 -146 1334
rect -118 1306 -80 1334
rect -52 1306 -14 1334
rect 14 1306 52 1334
rect 80 1306 118 1334
rect 146 1306 184 1334
rect 212 1306 250 1334
rect 278 1306 316 1334
rect 344 1306 349 1334
rect -349 1268 349 1306
rect -349 1240 -344 1268
rect -316 1240 -278 1268
rect -250 1240 -212 1268
rect -184 1240 -146 1268
rect -118 1240 -80 1268
rect -52 1240 -14 1268
rect 14 1240 52 1268
rect 80 1240 118 1268
rect 146 1240 184 1268
rect 212 1240 250 1268
rect 278 1240 316 1268
rect 344 1240 349 1268
rect -349 1202 349 1240
rect -349 1174 -344 1202
rect -316 1174 -278 1202
rect -250 1174 -212 1202
rect -184 1174 -146 1202
rect -118 1174 -80 1202
rect -52 1174 -14 1202
rect 14 1174 52 1202
rect 80 1174 118 1202
rect 146 1174 184 1202
rect 212 1174 250 1202
rect 278 1174 316 1202
rect 344 1174 349 1202
rect -349 1136 349 1174
rect -349 1108 -344 1136
rect -316 1108 -278 1136
rect -250 1108 -212 1136
rect -184 1108 -146 1136
rect -118 1108 -80 1136
rect -52 1108 -14 1136
rect 14 1108 52 1136
rect 80 1108 118 1136
rect 146 1108 184 1136
rect 212 1108 250 1136
rect 278 1108 316 1136
rect 344 1108 349 1136
rect -349 1070 349 1108
rect -349 1042 -344 1070
rect -316 1042 -278 1070
rect -250 1042 -212 1070
rect -184 1042 -146 1070
rect -118 1042 -80 1070
rect -52 1042 -14 1070
rect 14 1042 52 1070
rect 80 1042 118 1070
rect 146 1042 184 1070
rect 212 1042 250 1070
rect 278 1042 316 1070
rect 344 1042 349 1070
rect -349 1004 349 1042
rect -349 976 -344 1004
rect -316 976 -278 1004
rect -250 976 -212 1004
rect -184 976 -146 1004
rect -118 976 -80 1004
rect -52 976 -14 1004
rect 14 976 52 1004
rect 80 976 118 1004
rect 146 976 184 1004
rect 212 976 250 1004
rect 278 976 316 1004
rect 344 976 349 1004
rect -349 938 349 976
rect -349 910 -344 938
rect -316 910 -278 938
rect -250 910 -212 938
rect -184 910 -146 938
rect -118 910 -80 938
rect -52 910 -14 938
rect 14 910 52 938
rect 80 910 118 938
rect 146 910 184 938
rect 212 910 250 938
rect 278 910 316 938
rect 344 910 349 938
rect -349 872 349 910
rect -349 844 -344 872
rect -316 844 -278 872
rect -250 844 -212 872
rect -184 844 -146 872
rect -118 844 -80 872
rect -52 844 -14 872
rect 14 844 52 872
rect 80 844 118 872
rect 146 844 184 872
rect 212 844 250 872
rect 278 844 316 872
rect 344 844 349 872
rect -349 806 349 844
rect -349 778 -344 806
rect -316 778 -278 806
rect -250 778 -212 806
rect -184 778 -146 806
rect -118 778 -80 806
rect -52 778 -14 806
rect 14 778 52 806
rect 80 778 118 806
rect 146 778 184 806
rect 212 778 250 806
rect 278 778 316 806
rect 344 778 349 806
rect -349 740 349 778
rect -349 712 -344 740
rect -316 712 -278 740
rect -250 712 -212 740
rect -184 712 -146 740
rect -118 712 -80 740
rect -52 712 -14 740
rect 14 712 52 740
rect 80 712 118 740
rect 146 712 184 740
rect 212 712 250 740
rect 278 712 316 740
rect 344 712 349 740
rect -349 674 349 712
rect -349 646 -344 674
rect -316 646 -278 674
rect -250 646 -212 674
rect -184 646 -146 674
rect -118 646 -80 674
rect -52 646 -14 674
rect 14 646 52 674
rect 80 646 118 674
rect 146 646 184 674
rect 212 646 250 674
rect 278 646 316 674
rect 344 646 349 674
rect -349 608 349 646
rect -349 580 -344 608
rect -316 580 -278 608
rect -250 580 -212 608
rect -184 580 -146 608
rect -118 580 -80 608
rect -52 580 -14 608
rect 14 580 52 608
rect 80 580 118 608
rect 146 580 184 608
rect 212 580 250 608
rect 278 580 316 608
rect 344 580 349 608
rect -349 542 349 580
rect -349 514 -344 542
rect -316 514 -278 542
rect -250 514 -212 542
rect -184 514 -146 542
rect -118 514 -80 542
rect -52 514 -14 542
rect 14 514 52 542
rect 80 514 118 542
rect 146 514 184 542
rect 212 514 250 542
rect 278 514 316 542
rect 344 514 349 542
rect -349 476 349 514
rect -349 448 -344 476
rect -316 448 -278 476
rect -250 448 -212 476
rect -184 448 -146 476
rect -118 448 -80 476
rect -52 448 -14 476
rect 14 448 52 476
rect 80 448 118 476
rect 146 448 184 476
rect 212 448 250 476
rect 278 448 316 476
rect 344 448 349 476
rect -349 410 349 448
rect -349 382 -344 410
rect -316 382 -278 410
rect -250 382 -212 410
rect -184 382 -146 410
rect -118 382 -80 410
rect -52 382 -14 410
rect 14 382 52 410
rect 80 382 118 410
rect 146 382 184 410
rect 212 382 250 410
rect 278 382 316 410
rect 344 382 349 410
rect -349 344 349 382
rect -349 316 -344 344
rect -316 316 -278 344
rect -250 316 -212 344
rect -184 316 -146 344
rect -118 316 -80 344
rect -52 316 -14 344
rect 14 316 52 344
rect 80 316 118 344
rect 146 316 184 344
rect 212 316 250 344
rect 278 316 316 344
rect 344 316 349 344
rect -349 278 349 316
rect -349 250 -344 278
rect -316 250 -278 278
rect -250 250 -212 278
rect -184 250 -146 278
rect -118 250 -80 278
rect -52 250 -14 278
rect 14 250 52 278
rect 80 250 118 278
rect 146 250 184 278
rect 212 250 250 278
rect 278 250 316 278
rect 344 250 349 278
rect -349 212 349 250
rect -349 184 -344 212
rect -316 184 -278 212
rect -250 184 -212 212
rect -184 184 -146 212
rect -118 184 -80 212
rect -52 184 -14 212
rect 14 184 52 212
rect 80 184 118 212
rect 146 184 184 212
rect 212 184 250 212
rect 278 184 316 212
rect 344 184 349 212
rect -349 146 349 184
rect -349 118 -344 146
rect -316 118 -278 146
rect -250 118 -212 146
rect -184 118 -146 146
rect -118 118 -80 146
rect -52 118 -14 146
rect 14 118 52 146
rect 80 118 118 146
rect 146 118 184 146
rect 212 118 250 146
rect 278 118 316 146
rect 344 118 349 146
rect -349 80 349 118
rect -349 52 -344 80
rect -316 52 -278 80
rect -250 52 -212 80
rect -184 52 -146 80
rect -118 52 -80 80
rect -52 52 -14 80
rect 14 52 52 80
rect 80 52 118 80
rect 146 52 184 80
rect 212 52 250 80
rect 278 52 316 80
rect 344 52 349 80
rect -349 14 349 52
rect -349 -14 -344 14
rect -316 -14 -278 14
rect -250 -14 -212 14
rect -184 -14 -146 14
rect -118 -14 -80 14
rect -52 -14 -14 14
rect 14 -14 52 14
rect 80 -14 118 14
rect 146 -14 184 14
rect 212 -14 250 14
rect 278 -14 316 14
rect 344 -14 349 14
rect -349 -52 349 -14
rect -349 -80 -344 -52
rect -316 -80 -278 -52
rect -250 -80 -212 -52
rect -184 -80 -146 -52
rect -118 -80 -80 -52
rect -52 -80 -14 -52
rect 14 -80 52 -52
rect 80 -80 118 -52
rect 146 -80 184 -52
rect 212 -80 250 -52
rect 278 -80 316 -52
rect 344 -80 349 -52
rect -349 -118 349 -80
rect -349 -146 -344 -118
rect -316 -146 -278 -118
rect -250 -146 -212 -118
rect -184 -146 -146 -118
rect -118 -146 -80 -118
rect -52 -146 -14 -118
rect 14 -146 52 -118
rect 80 -146 118 -118
rect 146 -146 184 -118
rect 212 -146 250 -118
rect 278 -146 316 -118
rect 344 -146 349 -118
rect -349 -184 349 -146
rect -349 -212 -344 -184
rect -316 -212 -278 -184
rect -250 -212 -212 -184
rect -184 -212 -146 -184
rect -118 -212 -80 -184
rect -52 -212 -14 -184
rect 14 -212 52 -184
rect 80 -212 118 -184
rect 146 -212 184 -184
rect 212 -212 250 -184
rect 278 -212 316 -184
rect 344 -212 349 -184
rect -349 -250 349 -212
rect -349 -278 -344 -250
rect -316 -278 -278 -250
rect -250 -278 -212 -250
rect -184 -278 -146 -250
rect -118 -278 -80 -250
rect -52 -278 -14 -250
rect 14 -278 52 -250
rect 80 -278 118 -250
rect 146 -278 184 -250
rect 212 -278 250 -250
rect 278 -278 316 -250
rect 344 -278 349 -250
rect -349 -316 349 -278
rect -349 -344 -344 -316
rect -316 -344 -278 -316
rect -250 -344 -212 -316
rect -184 -344 -146 -316
rect -118 -344 -80 -316
rect -52 -344 -14 -316
rect 14 -344 52 -316
rect 80 -344 118 -316
rect 146 -344 184 -316
rect 212 -344 250 -316
rect 278 -344 316 -316
rect 344 -344 349 -316
rect -349 -382 349 -344
rect -349 -410 -344 -382
rect -316 -410 -278 -382
rect -250 -410 -212 -382
rect -184 -410 -146 -382
rect -118 -410 -80 -382
rect -52 -410 -14 -382
rect 14 -410 52 -382
rect 80 -410 118 -382
rect 146 -410 184 -382
rect 212 -410 250 -382
rect 278 -410 316 -382
rect 344 -410 349 -382
rect -349 -448 349 -410
rect -349 -476 -344 -448
rect -316 -476 -278 -448
rect -250 -476 -212 -448
rect -184 -476 -146 -448
rect -118 -476 -80 -448
rect -52 -476 -14 -448
rect 14 -476 52 -448
rect 80 -476 118 -448
rect 146 -476 184 -448
rect 212 -476 250 -448
rect 278 -476 316 -448
rect 344 -476 349 -448
rect -349 -514 349 -476
rect -349 -542 -344 -514
rect -316 -542 -278 -514
rect -250 -542 -212 -514
rect -184 -542 -146 -514
rect -118 -542 -80 -514
rect -52 -542 -14 -514
rect 14 -542 52 -514
rect 80 -542 118 -514
rect 146 -542 184 -514
rect 212 -542 250 -514
rect 278 -542 316 -514
rect 344 -542 349 -514
rect -349 -580 349 -542
rect -349 -608 -344 -580
rect -316 -608 -278 -580
rect -250 -608 -212 -580
rect -184 -608 -146 -580
rect -118 -608 -80 -580
rect -52 -608 -14 -580
rect 14 -608 52 -580
rect 80 -608 118 -580
rect 146 -608 184 -580
rect 212 -608 250 -580
rect 278 -608 316 -580
rect 344 -608 349 -580
rect -349 -646 349 -608
rect -349 -674 -344 -646
rect -316 -674 -278 -646
rect -250 -674 -212 -646
rect -184 -674 -146 -646
rect -118 -674 -80 -646
rect -52 -674 -14 -646
rect 14 -674 52 -646
rect 80 -674 118 -646
rect 146 -674 184 -646
rect 212 -674 250 -646
rect 278 -674 316 -646
rect 344 -674 349 -646
rect -349 -712 349 -674
rect -349 -740 -344 -712
rect -316 -740 -278 -712
rect -250 -740 -212 -712
rect -184 -740 -146 -712
rect -118 -740 -80 -712
rect -52 -740 -14 -712
rect 14 -740 52 -712
rect 80 -740 118 -712
rect 146 -740 184 -712
rect 212 -740 250 -712
rect 278 -740 316 -712
rect 344 -740 349 -712
rect -349 -778 349 -740
rect -349 -806 -344 -778
rect -316 -806 -278 -778
rect -250 -806 -212 -778
rect -184 -806 -146 -778
rect -118 -806 -80 -778
rect -52 -806 -14 -778
rect 14 -806 52 -778
rect 80 -806 118 -778
rect 146 -806 184 -778
rect 212 -806 250 -778
rect 278 -806 316 -778
rect 344 -806 349 -778
rect -349 -844 349 -806
rect -349 -872 -344 -844
rect -316 -872 -278 -844
rect -250 -872 -212 -844
rect -184 -872 -146 -844
rect -118 -872 -80 -844
rect -52 -872 -14 -844
rect 14 -872 52 -844
rect 80 -872 118 -844
rect 146 -872 184 -844
rect 212 -872 250 -844
rect 278 -872 316 -844
rect 344 -872 349 -844
rect -349 -910 349 -872
rect -349 -938 -344 -910
rect -316 -938 -278 -910
rect -250 -938 -212 -910
rect -184 -938 -146 -910
rect -118 -938 -80 -910
rect -52 -938 -14 -910
rect 14 -938 52 -910
rect 80 -938 118 -910
rect 146 -938 184 -910
rect 212 -938 250 -910
rect 278 -938 316 -910
rect 344 -938 349 -910
rect -349 -976 349 -938
rect -349 -1004 -344 -976
rect -316 -1004 -278 -976
rect -250 -1004 -212 -976
rect -184 -1004 -146 -976
rect -118 -1004 -80 -976
rect -52 -1004 -14 -976
rect 14 -1004 52 -976
rect 80 -1004 118 -976
rect 146 -1004 184 -976
rect 212 -1004 250 -976
rect 278 -1004 316 -976
rect 344 -1004 349 -976
rect -349 -1042 349 -1004
rect -349 -1070 -344 -1042
rect -316 -1070 -278 -1042
rect -250 -1070 -212 -1042
rect -184 -1070 -146 -1042
rect -118 -1070 -80 -1042
rect -52 -1070 -14 -1042
rect 14 -1070 52 -1042
rect 80 -1070 118 -1042
rect 146 -1070 184 -1042
rect 212 -1070 250 -1042
rect 278 -1070 316 -1042
rect 344 -1070 349 -1042
rect -349 -1108 349 -1070
rect -349 -1136 -344 -1108
rect -316 -1136 -278 -1108
rect -250 -1136 -212 -1108
rect -184 -1136 -146 -1108
rect -118 -1136 -80 -1108
rect -52 -1136 -14 -1108
rect 14 -1136 52 -1108
rect 80 -1136 118 -1108
rect 146 -1136 184 -1108
rect 212 -1136 250 -1108
rect 278 -1136 316 -1108
rect 344 -1136 349 -1108
rect -349 -1174 349 -1136
rect -349 -1202 -344 -1174
rect -316 -1202 -278 -1174
rect -250 -1202 -212 -1174
rect -184 -1202 -146 -1174
rect -118 -1202 -80 -1174
rect -52 -1202 -14 -1174
rect 14 -1202 52 -1174
rect 80 -1202 118 -1174
rect 146 -1202 184 -1174
rect 212 -1202 250 -1174
rect 278 -1202 316 -1174
rect 344 -1202 349 -1174
rect -349 -1240 349 -1202
rect -349 -1268 -344 -1240
rect -316 -1268 -278 -1240
rect -250 -1268 -212 -1240
rect -184 -1268 -146 -1240
rect -118 -1268 -80 -1240
rect -52 -1268 -14 -1240
rect 14 -1268 52 -1240
rect 80 -1268 118 -1240
rect 146 -1268 184 -1240
rect 212 -1268 250 -1240
rect 278 -1268 316 -1240
rect 344 -1268 349 -1240
rect -349 -1306 349 -1268
rect -349 -1334 -344 -1306
rect -316 -1334 -278 -1306
rect -250 -1334 -212 -1306
rect -184 -1334 -146 -1306
rect -118 -1334 -80 -1306
rect -52 -1334 -14 -1306
rect 14 -1334 52 -1306
rect 80 -1334 118 -1306
rect 146 -1334 184 -1306
rect 212 -1334 250 -1306
rect 278 -1334 316 -1306
rect 344 -1334 349 -1306
rect -349 -1372 349 -1334
rect -349 -1400 -344 -1372
rect -316 -1400 -278 -1372
rect -250 -1400 -212 -1372
rect -184 -1400 -146 -1372
rect -118 -1400 -80 -1372
rect -52 -1400 -14 -1372
rect 14 -1400 52 -1372
rect 80 -1400 118 -1372
rect 146 -1400 184 -1372
rect 212 -1400 250 -1372
rect 278 -1400 316 -1372
rect 344 -1400 349 -1372
rect -349 -1438 349 -1400
rect -349 -1466 -344 -1438
rect -316 -1466 -278 -1438
rect -250 -1466 -212 -1438
rect -184 -1466 -146 -1438
rect -118 -1466 -80 -1438
rect -52 -1466 -14 -1438
rect 14 -1466 52 -1438
rect 80 -1466 118 -1438
rect 146 -1466 184 -1438
rect 212 -1466 250 -1438
rect 278 -1466 316 -1438
rect 344 -1466 349 -1438
rect -349 -1504 349 -1466
rect -349 -1532 -344 -1504
rect -316 -1532 -278 -1504
rect -250 -1532 -212 -1504
rect -184 -1532 -146 -1504
rect -118 -1532 -80 -1504
rect -52 -1532 -14 -1504
rect 14 -1532 52 -1504
rect 80 -1532 118 -1504
rect 146 -1532 184 -1504
rect 212 -1532 250 -1504
rect 278 -1532 316 -1504
rect 344 -1532 349 -1504
rect -349 -1537 349 -1532
<< via3 >>
rect -344 1504 -316 1532
rect -278 1504 -250 1532
rect -212 1504 -184 1532
rect -146 1504 -118 1532
rect -80 1504 -52 1532
rect -14 1504 14 1532
rect 52 1504 80 1532
rect 118 1504 146 1532
rect 184 1504 212 1532
rect 250 1504 278 1532
rect 316 1504 344 1532
rect -344 1438 -316 1466
rect -278 1438 -250 1466
rect -212 1438 -184 1466
rect -146 1438 -118 1466
rect -80 1438 -52 1466
rect -14 1438 14 1466
rect 52 1438 80 1466
rect 118 1438 146 1466
rect 184 1438 212 1466
rect 250 1438 278 1466
rect 316 1438 344 1466
rect -344 1372 -316 1400
rect -278 1372 -250 1400
rect -212 1372 -184 1400
rect -146 1372 -118 1400
rect -80 1372 -52 1400
rect -14 1372 14 1400
rect 52 1372 80 1400
rect 118 1372 146 1400
rect 184 1372 212 1400
rect 250 1372 278 1400
rect 316 1372 344 1400
rect -344 1306 -316 1334
rect -278 1306 -250 1334
rect -212 1306 -184 1334
rect -146 1306 -118 1334
rect -80 1306 -52 1334
rect -14 1306 14 1334
rect 52 1306 80 1334
rect 118 1306 146 1334
rect 184 1306 212 1334
rect 250 1306 278 1334
rect 316 1306 344 1334
rect -344 1240 -316 1268
rect -278 1240 -250 1268
rect -212 1240 -184 1268
rect -146 1240 -118 1268
rect -80 1240 -52 1268
rect -14 1240 14 1268
rect 52 1240 80 1268
rect 118 1240 146 1268
rect 184 1240 212 1268
rect 250 1240 278 1268
rect 316 1240 344 1268
rect -344 1174 -316 1202
rect -278 1174 -250 1202
rect -212 1174 -184 1202
rect -146 1174 -118 1202
rect -80 1174 -52 1202
rect -14 1174 14 1202
rect 52 1174 80 1202
rect 118 1174 146 1202
rect 184 1174 212 1202
rect 250 1174 278 1202
rect 316 1174 344 1202
rect -344 1108 -316 1136
rect -278 1108 -250 1136
rect -212 1108 -184 1136
rect -146 1108 -118 1136
rect -80 1108 -52 1136
rect -14 1108 14 1136
rect 52 1108 80 1136
rect 118 1108 146 1136
rect 184 1108 212 1136
rect 250 1108 278 1136
rect 316 1108 344 1136
rect -344 1042 -316 1070
rect -278 1042 -250 1070
rect -212 1042 -184 1070
rect -146 1042 -118 1070
rect -80 1042 -52 1070
rect -14 1042 14 1070
rect 52 1042 80 1070
rect 118 1042 146 1070
rect 184 1042 212 1070
rect 250 1042 278 1070
rect 316 1042 344 1070
rect -344 976 -316 1004
rect -278 976 -250 1004
rect -212 976 -184 1004
rect -146 976 -118 1004
rect -80 976 -52 1004
rect -14 976 14 1004
rect 52 976 80 1004
rect 118 976 146 1004
rect 184 976 212 1004
rect 250 976 278 1004
rect 316 976 344 1004
rect -344 910 -316 938
rect -278 910 -250 938
rect -212 910 -184 938
rect -146 910 -118 938
rect -80 910 -52 938
rect -14 910 14 938
rect 52 910 80 938
rect 118 910 146 938
rect 184 910 212 938
rect 250 910 278 938
rect 316 910 344 938
rect -344 844 -316 872
rect -278 844 -250 872
rect -212 844 -184 872
rect -146 844 -118 872
rect -80 844 -52 872
rect -14 844 14 872
rect 52 844 80 872
rect 118 844 146 872
rect 184 844 212 872
rect 250 844 278 872
rect 316 844 344 872
rect -344 778 -316 806
rect -278 778 -250 806
rect -212 778 -184 806
rect -146 778 -118 806
rect -80 778 -52 806
rect -14 778 14 806
rect 52 778 80 806
rect 118 778 146 806
rect 184 778 212 806
rect 250 778 278 806
rect 316 778 344 806
rect -344 712 -316 740
rect -278 712 -250 740
rect -212 712 -184 740
rect -146 712 -118 740
rect -80 712 -52 740
rect -14 712 14 740
rect 52 712 80 740
rect 118 712 146 740
rect 184 712 212 740
rect 250 712 278 740
rect 316 712 344 740
rect -344 646 -316 674
rect -278 646 -250 674
rect -212 646 -184 674
rect -146 646 -118 674
rect -80 646 -52 674
rect -14 646 14 674
rect 52 646 80 674
rect 118 646 146 674
rect 184 646 212 674
rect 250 646 278 674
rect 316 646 344 674
rect -344 580 -316 608
rect -278 580 -250 608
rect -212 580 -184 608
rect -146 580 -118 608
rect -80 580 -52 608
rect -14 580 14 608
rect 52 580 80 608
rect 118 580 146 608
rect 184 580 212 608
rect 250 580 278 608
rect 316 580 344 608
rect -344 514 -316 542
rect -278 514 -250 542
rect -212 514 -184 542
rect -146 514 -118 542
rect -80 514 -52 542
rect -14 514 14 542
rect 52 514 80 542
rect 118 514 146 542
rect 184 514 212 542
rect 250 514 278 542
rect 316 514 344 542
rect -344 448 -316 476
rect -278 448 -250 476
rect -212 448 -184 476
rect -146 448 -118 476
rect -80 448 -52 476
rect -14 448 14 476
rect 52 448 80 476
rect 118 448 146 476
rect 184 448 212 476
rect 250 448 278 476
rect 316 448 344 476
rect -344 382 -316 410
rect -278 382 -250 410
rect -212 382 -184 410
rect -146 382 -118 410
rect -80 382 -52 410
rect -14 382 14 410
rect 52 382 80 410
rect 118 382 146 410
rect 184 382 212 410
rect 250 382 278 410
rect 316 382 344 410
rect -344 316 -316 344
rect -278 316 -250 344
rect -212 316 -184 344
rect -146 316 -118 344
rect -80 316 -52 344
rect -14 316 14 344
rect 52 316 80 344
rect 118 316 146 344
rect 184 316 212 344
rect 250 316 278 344
rect 316 316 344 344
rect -344 250 -316 278
rect -278 250 -250 278
rect -212 250 -184 278
rect -146 250 -118 278
rect -80 250 -52 278
rect -14 250 14 278
rect 52 250 80 278
rect 118 250 146 278
rect 184 250 212 278
rect 250 250 278 278
rect 316 250 344 278
rect -344 184 -316 212
rect -278 184 -250 212
rect -212 184 -184 212
rect -146 184 -118 212
rect -80 184 -52 212
rect -14 184 14 212
rect 52 184 80 212
rect 118 184 146 212
rect 184 184 212 212
rect 250 184 278 212
rect 316 184 344 212
rect -344 118 -316 146
rect -278 118 -250 146
rect -212 118 -184 146
rect -146 118 -118 146
rect -80 118 -52 146
rect -14 118 14 146
rect 52 118 80 146
rect 118 118 146 146
rect 184 118 212 146
rect 250 118 278 146
rect 316 118 344 146
rect -344 52 -316 80
rect -278 52 -250 80
rect -212 52 -184 80
rect -146 52 -118 80
rect -80 52 -52 80
rect -14 52 14 80
rect 52 52 80 80
rect 118 52 146 80
rect 184 52 212 80
rect 250 52 278 80
rect 316 52 344 80
rect -344 -14 -316 14
rect -278 -14 -250 14
rect -212 -14 -184 14
rect -146 -14 -118 14
rect -80 -14 -52 14
rect -14 -14 14 14
rect 52 -14 80 14
rect 118 -14 146 14
rect 184 -14 212 14
rect 250 -14 278 14
rect 316 -14 344 14
rect -344 -80 -316 -52
rect -278 -80 -250 -52
rect -212 -80 -184 -52
rect -146 -80 -118 -52
rect -80 -80 -52 -52
rect -14 -80 14 -52
rect 52 -80 80 -52
rect 118 -80 146 -52
rect 184 -80 212 -52
rect 250 -80 278 -52
rect 316 -80 344 -52
rect -344 -146 -316 -118
rect -278 -146 -250 -118
rect -212 -146 -184 -118
rect -146 -146 -118 -118
rect -80 -146 -52 -118
rect -14 -146 14 -118
rect 52 -146 80 -118
rect 118 -146 146 -118
rect 184 -146 212 -118
rect 250 -146 278 -118
rect 316 -146 344 -118
rect -344 -212 -316 -184
rect -278 -212 -250 -184
rect -212 -212 -184 -184
rect -146 -212 -118 -184
rect -80 -212 -52 -184
rect -14 -212 14 -184
rect 52 -212 80 -184
rect 118 -212 146 -184
rect 184 -212 212 -184
rect 250 -212 278 -184
rect 316 -212 344 -184
rect -344 -278 -316 -250
rect -278 -278 -250 -250
rect -212 -278 -184 -250
rect -146 -278 -118 -250
rect -80 -278 -52 -250
rect -14 -278 14 -250
rect 52 -278 80 -250
rect 118 -278 146 -250
rect 184 -278 212 -250
rect 250 -278 278 -250
rect 316 -278 344 -250
rect -344 -344 -316 -316
rect -278 -344 -250 -316
rect -212 -344 -184 -316
rect -146 -344 -118 -316
rect -80 -344 -52 -316
rect -14 -344 14 -316
rect 52 -344 80 -316
rect 118 -344 146 -316
rect 184 -344 212 -316
rect 250 -344 278 -316
rect 316 -344 344 -316
rect -344 -410 -316 -382
rect -278 -410 -250 -382
rect -212 -410 -184 -382
rect -146 -410 -118 -382
rect -80 -410 -52 -382
rect -14 -410 14 -382
rect 52 -410 80 -382
rect 118 -410 146 -382
rect 184 -410 212 -382
rect 250 -410 278 -382
rect 316 -410 344 -382
rect -344 -476 -316 -448
rect -278 -476 -250 -448
rect -212 -476 -184 -448
rect -146 -476 -118 -448
rect -80 -476 -52 -448
rect -14 -476 14 -448
rect 52 -476 80 -448
rect 118 -476 146 -448
rect 184 -476 212 -448
rect 250 -476 278 -448
rect 316 -476 344 -448
rect -344 -542 -316 -514
rect -278 -542 -250 -514
rect -212 -542 -184 -514
rect -146 -542 -118 -514
rect -80 -542 -52 -514
rect -14 -542 14 -514
rect 52 -542 80 -514
rect 118 -542 146 -514
rect 184 -542 212 -514
rect 250 -542 278 -514
rect 316 -542 344 -514
rect -344 -608 -316 -580
rect -278 -608 -250 -580
rect -212 -608 -184 -580
rect -146 -608 -118 -580
rect -80 -608 -52 -580
rect -14 -608 14 -580
rect 52 -608 80 -580
rect 118 -608 146 -580
rect 184 -608 212 -580
rect 250 -608 278 -580
rect 316 -608 344 -580
rect -344 -674 -316 -646
rect -278 -674 -250 -646
rect -212 -674 -184 -646
rect -146 -674 -118 -646
rect -80 -674 -52 -646
rect -14 -674 14 -646
rect 52 -674 80 -646
rect 118 -674 146 -646
rect 184 -674 212 -646
rect 250 -674 278 -646
rect 316 -674 344 -646
rect -344 -740 -316 -712
rect -278 -740 -250 -712
rect -212 -740 -184 -712
rect -146 -740 -118 -712
rect -80 -740 -52 -712
rect -14 -740 14 -712
rect 52 -740 80 -712
rect 118 -740 146 -712
rect 184 -740 212 -712
rect 250 -740 278 -712
rect 316 -740 344 -712
rect -344 -806 -316 -778
rect -278 -806 -250 -778
rect -212 -806 -184 -778
rect -146 -806 -118 -778
rect -80 -806 -52 -778
rect -14 -806 14 -778
rect 52 -806 80 -778
rect 118 -806 146 -778
rect 184 -806 212 -778
rect 250 -806 278 -778
rect 316 -806 344 -778
rect -344 -872 -316 -844
rect -278 -872 -250 -844
rect -212 -872 -184 -844
rect -146 -872 -118 -844
rect -80 -872 -52 -844
rect -14 -872 14 -844
rect 52 -872 80 -844
rect 118 -872 146 -844
rect 184 -872 212 -844
rect 250 -872 278 -844
rect 316 -872 344 -844
rect -344 -938 -316 -910
rect -278 -938 -250 -910
rect -212 -938 -184 -910
rect -146 -938 -118 -910
rect -80 -938 -52 -910
rect -14 -938 14 -910
rect 52 -938 80 -910
rect 118 -938 146 -910
rect 184 -938 212 -910
rect 250 -938 278 -910
rect 316 -938 344 -910
rect -344 -1004 -316 -976
rect -278 -1004 -250 -976
rect -212 -1004 -184 -976
rect -146 -1004 -118 -976
rect -80 -1004 -52 -976
rect -14 -1004 14 -976
rect 52 -1004 80 -976
rect 118 -1004 146 -976
rect 184 -1004 212 -976
rect 250 -1004 278 -976
rect 316 -1004 344 -976
rect -344 -1070 -316 -1042
rect -278 -1070 -250 -1042
rect -212 -1070 -184 -1042
rect -146 -1070 -118 -1042
rect -80 -1070 -52 -1042
rect -14 -1070 14 -1042
rect 52 -1070 80 -1042
rect 118 -1070 146 -1042
rect 184 -1070 212 -1042
rect 250 -1070 278 -1042
rect 316 -1070 344 -1042
rect -344 -1136 -316 -1108
rect -278 -1136 -250 -1108
rect -212 -1136 -184 -1108
rect -146 -1136 -118 -1108
rect -80 -1136 -52 -1108
rect -14 -1136 14 -1108
rect 52 -1136 80 -1108
rect 118 -1136 146 -1108
rect 184 -1136 212 -1108
rect 250 -1136 278 -1108
rect 316 -1136 344 -1108
rect -344 -1202 -316 -1174
rect -278 -1202 -250 -1174
rect -212 -1202 -184 -1174
rect -146 -1202 -118 -1174
rect -80 -1202 -52 -1174
rect -14 -1202 14 -1174
rect 52 -1202 80 -1174
rect 118 -1202 146 -1174
rect 184 -1202 212 -1174
rect 250 -1202 278 -1174
rect 316 -1202 344 -1174
rect -344 -1268 -316 -1240
rect -278 -1268 -250 -1240
rect -212 -1268 -184 -1240
rect -146 -1268 -118 -1240
rect -80 -1268 -52 -1240
rect -14 -1268 14 -1240
rect 52 -1268 80 -1240
rect 118 -1268 146 -1240
rect 184 -1268 212 -1240
rect 250 -1268 278 -1240
rect 316 -1268 344 -1240
rect -344 -1334 -316 -1306
rect -278 -1334 -250 -1306
rect -212 -1334 -184 -1306
rect -146 -1334 -118 -1306
rect -80 -1334 -52 -1306
rect -14 -1334 14 -1306
rect 52 -1334 80 -1306
rect 118 -1334 146 -1306
rect 184 -1334 212 -1306
rect 250 -1334 278 -1306
rect 316 -1334 344 -1306
rect -344 -1400 -316 -1372
rect -278 -1400 -250 -1372
rect -212 -1400 -184 -1372
rect -146 -1400 -118 -1372
rect -80 -1400 -52 -1372
rect -14 -1400 14 -1372
rect 52 -1400 80 -1372
rect 118 -1400 146 -1372
rect 184 -1400 212 -1372
rect 250 -1400 278 -1372
rect 316 -1400 344 -1372
rect -344 -1466 -316 -1438
rect -278 -1466 -250 -1438
rect -212 -1466 -184 -1438
rect -146 -1466 -118 -1438
rect -80 -1466 -52 -1438
rect -14 -1466 14 -1438
rect 52 -1466 80 -1438
rect 118 -1466 146 -1438
rect 184 -1466 212 -1438
rect 250 -1466 278 -1438
rect 316 -1466 344 -1438
rect -344 -1532 -316 -1504
rect -278 -1532 -250 -1504
rect -212 -1532 -184 -1504
rect -146 -1532 -118 -1504
rect -80 -1532 -52 -1504
rect -14 -1532 14 -1504
rect 52 -1532 80 -1504
rect 118 -1532 146 -1504
rect 184 -1532 212 -1504
rect 250 -1532 278 -1504
rect 316 -1532 344 -1504
<< metal4 >>
rect -349 1532 349 1537
rect -349 1504 -344 1532
rect -316 1504 -278 1532
rect -250 1504 -212 1532
rect -184 1504 -146 1532
rect -118 1504 -80 1532
rect -52 1504 -14 1532
rect 14 1504 52 1532
rect 80 1504 118 1532
rect 146 1504 184 1532
rect 212 1504 250 1532
rect 278 1504 316 1532
rect 344 1504 349 1532
rect -349 1466 349 1504
rect -349 1438 -344 1466
rect -316 1438 -278 1466
rect -250 1438 -212 1466
rect -184 1438 -146 1466
rect -118 1438 -80 1466
rect -52 1438 -14 1466
rect 14 1438 52 1466
rect 80 1438 118 1466
rect 146 1438 184 1466
rect 212 1438 250 1466
rect 278 1438 316 1466
rect 344 1438 349 1466
rect -349 1400 349 1438
rect -349 1372 -344 1400
rect -316 1372 -278 1400
rect -250 1372 -212 1400
rect -184 1372 -146 1400
rect -118 1372 -80 1400
rect -52 1372 -14 1400
rect 14 1372 52 1400
rect 80 1372 118 1400
rect 146 1372 184 1400
rect 212 1372 250 1400
rect 278 1372 316 1400
rect 344 1372 349 1400
rect -349 1334 349 1372
rect -349 1306 -344 1334
rect -316 1306 -278 1334
rect -250 1306 -212 1334
rect -184 1306 -146 1334
rect -118 1306 -80 1334
rect -52 1306 -14 1334
rect 14 1306 52 1334
rect 80 1306 118 1334
rect 146 1306 184 1334
rect 212 1306 250 1334
rect 278 1306 316 1334
rect 344 1306 349 1334
rect -349 1268 349 1306
rect -349 1240 -344 1268
rect -316 1240 -278 1268
rect -250 1240 -212 1268
rect -184 1240 -146 1268
rect -118 1240 -80 1268
rect -52 1240 -14 1268
rect 14 1240 52 1268
rect 80 1240 118 1268
rect 146 1240 184 1268
rect 212 1240 250 1268
rect 278 1240 316 1268
rect 344 1240 349 1268
rect -349 1202 349 1240
rect -349 1174 -344 1202
rect -316 1174 -278 1202
rect -250 1174 -212 1202
rect -184 1174 -146 1202
rect -118 1174 -80 1202
rect -52 1174 -14 1202
rect 14 1174 52 1202
rect 80 1174 118 1202
rect 146 1174 184 1202
rect 212 1174 250 1202
rect 278 1174 316 1202
rect 344 1174 349 1202
rect -349 1136 349 1174
rect -349 1108 -344 1136
rect -316 1108 -278 1136
rect -250 1108 -212 1136
rect -184 1108 -146 1136
rect -118 1108 -80 1136
rect -52 1108 -14 1136
rect 14 1108 52 1136
rect 80 1108 118 1136
rect 146 1108 184 1136
rect 212 1108 250 1136
rect 278 1108 316 1136
rect 344 1108 349 1136
rect -349 1070 349 1108
rect -349 1042 -344 1070
rect -316 1042 -278 1070
rect -250 1042 -212 1070
rect -184 1042 -146 1070
rect -118 1042 -80 1070
rect -52 1042 -14 1070
rect 14 1042 52 1070
rect 80 1042 118 1070
rect 146 1042 184 1070
rect 212 1042 250 1070
rect 278 1042 316 1070
rect 344 1042 349 1070
rect -349 1004 349 1042
rect -349 976 -344 1004
rect -316 976 -278 1004
rect -250 976 -212 1004
rect -184 976 -146 1004
rect -118 976 -80 1004
rect -52 976 -14 1004
rect 14 976 52 1004
rect 80 976 118 1004
rect 146 976 184 1004
rect 212 976 250 1004
rect 278 976 316 1004
rect 344 976 349 1004
rect -349 938 349 976
rect -349 910 -344 938
rect -316 910 -278 938
rect -250 910 -212 938
rect -184 910 -146 938
rect -118 910 -80 938
rect -52 910 -14 938
rect 14 910 52 938
rect 80 910 118 938
rect 146 910 184 938
rect 212 910 250 938
rect 278 910 316 938
rect 344 910 349 938
rect -349 872 349 910
rect -349 844 -344 872
rect -316 844 -278 872
rect -250 844 -212 872
rect -184 844 -146 872
rect -118 844 -80 872
rect -52 844 -14 872
rect 14 844 52 872
rect 80 844 118 872
rect 146 844 184 872
rect 212 844 250 872
rect 278 844 316 872
rect 344 844 349 872
rect -349 806 349 844
rect -349 778 -344 806
rect -316 778 -278 806
rect -250 778 -212 806
rect -184 778 -146 806
rect -118 778 -80 806
rect -52 778 -14 806
rect 14 778 52 806
rect 80 778 118 806
rect 146 778 184 806
rect 212 778 250 806
rect 278 778 316 806
rect 344 778 349 806
rect -349 740 349 778
rect -349 712 -344 740
rect -316 712 -278 740
rect -250 712 -212 740
rect -184 712 -146 740
rect -118 712 -80 740
rect -52 712 -14 740
rect 14 712 52 740
rect 80 712 118 740
rect 146 712 184 740
rect 212 712 250 740
rect 278 712 316 740
rect 344 712 349 740
rect -349 674 349 712
rect -349 646 -344 674
rect -316 646 -278 674
rect -250 646 -212 674
rect -184 646 -146 674
rect -118 646 -80 674
rect -52 646 -14 674
rect 14 646 52 674
rect 80 646 118 674
rect 146 646 184 674
rect 212 646 250 674
rect 278 646 316 674
rect 344 646 349 674
rect -349 608 349 646
rect -349 580 -344 608
rect -316 580 -278 608
rect -250 580 -212 608
rect -184 580 -146 608
rect -118 580 -80 608
rect -52 580 -14 608
rect 14 580 52 608
rect 80 580 118 608
rect 146 580 184 608
rect 212 580 250 608
rect 278 580 316 608
rect 344 580 349 608
rect -349 542 349 580
rect -349 514 -344 542
rect -316 514 -278 542
rect -250 514 -212 542
rect -184 514 -146 542
rect -118 514 -80 542
rect -52 514 -14 542
rect 14 514 52 542
rect 80 514 118 542
rect 146 514 184 542
rect 212 514 250 542
rect 278 514 316 542
rect 344 514 349 542
rect -349 476 349 514
rect -349 448 -344 476
rect -316 448 -278 476
rect -250 448 -212 476
rect -184 448 -146 476
rect -118 448 -80 476
rect -52 448 -14 476
rect 14 448 52 476
rect 80 448 118 476
rect 146 448 184 476
rect 212 448 250 476
rect 278 448 316 476
rect 344 448 349 476
rect -349 410 349 448
rect -349 382 -344 410
rect -316 382 -278 410
rect -250 382 -212 410
rect -184 382 -146 410
rect -118 382 -80 410
rect -52 382 -14 410
rect 14 382 52 410
rect 80 382 118 410
rect 146 382 184 410
rect 212 382 250 410
rect 278 382 316 410
rect 344 382 349 410
rect -349 344 349 382
rect -349 316 -344 344
rect -316 316 -278 344
rect -250 316 -212 344
rect -184 316 -146 344
rect -118 316 -80 344
rect -52 316 -14 344
rect 14 316 52 344
rect 80 316 118 344
rect 146 316 184 344
rect 212 316 250 344
rect 278 316 316 344
rect 344 316 349 344
rect -349 278 349 316
rect -349 250 -344 278
rect -316 250 -278 278
rect -250 250 -212 278
rect -184 250 -146 278
rect -118 250 -80 278
rect -52 250 -14 278
rect 14 250 52 278
rect 80 250 118 278
rect 146 250 184 278
rect 212 250 250 278
rect 278 250 316 278
rect 344 250 349 278
rect -349 212 349 250
rect -349 184 -344 212
rect -316 184 -278 212
rect -250 184 -212 212
rect -184 184 -146 212
rect -118 184 -80 212
rect -52 184 -14 212
rect 14 184 52 212
rect 80 184 118 212
rect 146 184 184 212
rect 212 184 250 212
rect 278 184 316 212
rect 344 184 349 212
rect -349 146 349 184
rect -349 118 -344 146
rect -316 118 -278 146
rect -250 118 -212 146
rect -184 118 -146 146
rect -118 118 -80 146
rect -52 118 -14 146
rect 14 118 52 146
rect 80 118 118 146
rect 146 118 184 146
rect 212 118 250 146
rect 278 118 316 146
rect 344 118 349 146
rect -349 80 349 118
rect -349 52 -344 80
rect -316 52 -278 80
rect -250 52 -212 80
rect -184 52 -146 80
rect -118 52 -80 80
rect -52 52 -14 80
rect 14 52 52 80
rect 80 52 118 80
rect 146 52 184 80
rect 212 52 250 80
rect 278 52 316 80
rect 344 52 349 80
rect -349 14 349 52
rect -349 -14 -344 14
rect -316 -14 -278 14
rect -250 -14 -212 14
rect -184 -14 -146 14
rect -118 -14 -80 14
rect -52 -14 -14 14
rect 14 -14 52 14
rect 80 -14 118 14
rect 146 -14 184 14
rect 212 -14 250 14
rect 278 -14 316 14
rect 344 -14 349 14
rect -349 -52 349 -14
rect -349 -80 -344 -52
rect -316 -80 -278 -52
rect -250 -80 -212 -52
rect -184 -80 -146 -52
rect -118 -80 -80 -52
rect -52 -80 -14 -52
rect 14 -80 52 -52
rect 80 -80 118 -52
rect 146 -80 184 -52
rect 212 -80 250 -52
rect 278 -80 316 -52
rect 344 -80 349 -52
rect -349 -118 349 -80
rect -349 -146 -344 -118
rect -316 -146 -278 -118
rect -250 -146 -212 -118
rect -184 -146 -146 -118
rect -118 -146 -80 -118
rect -52 -146 -14 -118
rect 14 -146 52 -118
rect 80 -146 118 -118
rect 146 -146 184 -118
rect 212 -146 250 -118
rect 278 -146 316 -118
rect 344 -146 349 -118
rect -349 -184 349 -146
rect -349 -212 -344 -184
rect -316 -212 -278 -184
rect -250 -212 -212 -184
rect -184 -212 -146 -184
rect -118 -212 -80 -184
rect -52 -212 -14 -184
rect 14 -212 52 -184
rect 80 -212 118 -184
rect 146 -212 184 -184
rect 212 -212 250 -184
rect 278 -212 316 -184
rect 344 -212 349 -184
rect -349 -250 349 -212
rect -349 -278 -344 -250
rect -316 -278 -278 -250
rect -250 -278 -212 -250
rect -184 -278 -146 -250
rect -118 -278 -80 -250
rect -52 -278 -14 -250
rect 14 -278 52 -250
rect 80 -278 118 -250
rect 146 -278 184 -250
rect 212 -278 250 -250
rect 278 -278 316 -250
rect 344 -278 349 -250
rect -349 -316 349 -278
rect -349 -344 -344 -316
rect -316 -344 -278 -316
rect -250 -344 -212 -316
rect -184 -344 -146 -316
rect -118 -344 -80 -316
rect -52 -344 -14 -316
rect 14 -344 52 -316
rect 80 -344 118 -316
rect 146 -344 184 -316
rect 212 -344 250 -316
rect 278 -344 316 -316
rect 344 -344 349 -316
rect -349 -382 349 -344
rect -349 -410 -344 -382
rect -316 -410 -278 -382
rect -250 -410 -212 -382
rect -184 -410 -146 -382
rect -118 -410 -80 -382
rect -52 -410 -14 -382
rect 14 -410 52 -382
rect 80 -410 118 -382
rect 146 -410 184 -382
rect 212 -410 250 -382
rect 278 -410 316 -382
rect 344 -410 349 -382
rect -349 -448 349 -410
rect -349 -476 -344 -448
rect -316 -476 -278 -448
rect -250 -476 -212 -448
rect -184 -476 -146 -448
rect -118 -476 -80 -448
rect -52 -476 -14 -448
rect 14 -476 52 -448
rect 80 -476 118 -448
rect 146 -476 184 -448
rect 212 -476 250 -448
rect 278 -476 316 -448
rect 344 -476 349 -448
rect -349 -514 349 -476
rect -349 -542 -344 -514
rect -316 -542 -278 -514
rect -250 -542 -212 -514
rect -184 -542 -146 -514
rect -118 -542 -80 -514
rect -52 -542 -14 -514
rect 14 -542 52 -514
rect 80 -542 118 -514
rect 146 -542 184 -514
rect 212 -542 250 -514
rect 278 -542 316 -514
rect 344 -542 349 -514
rect -349 -580 349 -542
rect -349 -608 -344 -580
rect -316 -608 -278 -580
rect -250 -608 -212 -580
rect -184 -608 -146 -580
rect -118 -608 -80 -580
rect -52 -608 -14 -580
rect 14 -608 52 -580
rect 80 -608 118 -580
rect 146 -608 184 -580
rect 212 -608 250 -580
rect 278 -608 316 -580
rect 344 -608 349 -580
rect -349 -646 349 -608
rect -349 -674 -344 -646
rect -316 -674 -278 -646
rect -250 -674 -212 -646
rect -184 -674 -146 -646
rect -118 -674 -80 -646
rect -52 -674 -14 -646
rect 14 -674 52 -646
rect 80 -674 118 -646
rect 146 -674 184 -646
rect 212 -674 250 -646
rect 278 -674 316 -646
rect 344 -674 349 -646
rect -349 -712 349 -674
rect -349 -740 -344 -712
rect -316 -740 -278 -712
rect -250 -740 -212 -712
rect -184 -740 -146 -712
rect -118 -740 -80 -712
rect -52 -740 -14 -712
rect 14 -740 52 -712
rect 80 -740 118 -712
rect 146 -740 184 -712
rect 212 -740 250 -712
rect 278 -740 316 -712
rect 344 -740 349 -712
rect -349 -778 349 -740
rect -349 -806 -344 -778
rect -316 -806 -278 -778
rect -250 -806 -212 -778
rect -184 -806 -146 -778
rect -118 -806 -80 -778
rect -52 -806 -14 -778
rect 14 -806 52 -778
rect 80 -806 118 -778
rect 146 -806 184 -778
rect 212 -806 250 -778
rect 278 -806 316 -778
rect 344 -806 349 -778
rect -349 -844 349 -806
rect -349 -872 -344 -844
rect -316 -872 -278 -844
rect -250 -872 -212 -844
rect -184 -872 -146 -844
rect -118 -872 -80 -844
rect -52 -872 -14 -844
rect 14 -872 52 -844
rect 80 -872 118 -844
rect 146 -872 184 -844
rect 212 -872 250 -844
rect 278 -872 316 -844
rect 344 -872 349 -844
rect -349 -910 349 -872
rect -349 -938 -344 -910
rect -316 -938 -278 -910
rect -250 -938 -212 -910
rect -184 -938 -146 -910
rect -118 -938 -80 -910
rect -52 -938 -14 -910
rect 14 -938 52 -910
rect 80 -938 118 -910
rect 146 -938 184 -910
rect 212 -938 250 -910
rect 278 -938 316 -910
rect 344 -938 349 -910
rect -349 -976 349 -938
rect -349 -1004 -344 -976
rect -316 -1004 -278 -976
rect -250 -1004 -212 -976
rect -184 -1004 -146 -976
rect -118 -1004 -80 -976
rect -52 -1004 -14 -976
rect 14 -1004 52 -976
rect 80 -1004 118 -976
rect 146 -1004 184 -976
rect 212 -1004 250 -976
rect 278 -1004 316 -976
rect 344 -1004 349 -976
rect -349 -1042 349 -1004
rect -349 -1070 -344 -1042
rect -316 -1070 -278 -1042
rect -250 -1070 -212 -1042
rect -184 -1070 -146 -1042
rect -118 -1070 -80 -1042
rect -52 -1070 -14 -1042
rect 14 -1070 52 -1042
rect 80 -1070 118 -1042
rect 146 -1070 184 -1042
rect 212 -1070 250 -1042
rect 278 -1070 316 -1042
rect 344 -1070 349 -1042
rect -349 -1108 349 -1070
rect -349 -1136 -344 -1108
rect -316 -1136 -278 -1108
rect -250 -1136 -212 -1108
rect -184 -1136 -146 -1108
rect -118 -1136 -80 -1108
rect -52 -1136 -14 -1108
rect 14 -1136 52 -1108
rect 80 -1136 118 -1108
rect 146 -1136 184 -1108
rect 212 -1136 250 -1108
rect 278 -1136 316 -1108
rect 344 -1136 349 -1108
rect -349 -1174 349 -1136
rect -349 -1202 -344 -1174
rect -316 -1202 -278 -1174
rect -250 -1202 -212 -1174
rect -184 -1202 -146 -1174
rect -118 -1202 -80 -1174
rect -52 -1202 -14 -1174
rect 14 -1202 52 -1174
rect 80 -1202 118 -1174
rect 146 -1202 184 -1174
rect 212 -1202 250 -1174
rect 278 -1202 316 -1174
rect 344 -1202 349 -1174
rect -349 -1240 349 -1202
rect -349 -1268 -344 -1240
rect -316 -1268 -278 -1240
rect -250 -1268 -212 -1240
rect -184 -1268 -146 -1240
rect -118 -1268 -80 -1240
rect -52 -1268 -14 -1240
rect 14 -1268 52 -1240
rect 80 -1268 118 -1240
rect 146 -1268 184 -1240
rect 212 -1268 250 -1240
rect 278 -1268 316 -1240
rect 344 -1268 349 -1240
rect -349 -1306 349 -1268
rect -349 -1334 -344 -1306
rect -316 -1334 -278 -1306
rect -250 -1334 -212 -1306
rect -184 -1334 -146 -1306
rect -118 -1334 -80 -1306
rect -52 -1334 -14 -1306
rect 14 -1334 52 -1306
rect 80 -1334 118 -1306
rect 146 -1334 184 -1306
rect 212 -1334 250 -1306
rect 278 -1334 316 -1306
rect 344 -1334 349 -1306
rect -349 -1372 349 -1334
rect -349 -1400 -344 -1372
rect -316 -1400 -278 -1372
rect -250 -1400 -212 -1372
rect -184 -1400 -146 -1372
rect -118 -1400 -80 -1372
rect -52 -1400 -14 -1372
rect 14 -1400 52 -1372
rect 80 -1400 118 -1372
rect 146 -1400 184 -1372
rect 212 -1400 250 -1372
rect 278 -1400 316 -1372
rect 344 -1400 349 -1372
rect -349 -1438 349 -1400
rect -349 -1466 -344 -1438
rect -316 -1466 -278 -1438
rect -250 -1466 -212 -1438
rect -184 -1466 -146 -1438
rect -118 -1466 -80 -1438
rect -52 -1466 -14 -1438
rect 14 -1466 52 -1438
rect 80 -1466 118 -1438
rect 146 -1466 184 -1438
rect 212 -1466 250 -1438
rect 278 -1466 316 -1438
rect 344 -1466 349 -1438
rect -349 -1504 349 -1466
rect -349 -1532 -344 -1504
rect -316 -1532 -278 -1504
rect -250 -1532 -212 -1504
rect -184 -1532 -146 -1504
rect -118 -1532 -80 -1504
rect -52 -1532 -14 -1504
rect 14 -1532 52 -1504
rect 80 -1532 118 -1504
rect 146 -1532 184 -1504
rect 212 -1532 250 -1504
rect 278 -1532 316 -1504
rect 344 -1532 349 -1504
rect -349 -1537 349 -1532
<< end >>
