magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2045 -3784 2045 3784
<< psubdiff >>
rect -45 1762 45 1784
rect -45 -1762 -23 1762
rect 23 -1762 45 1762
rect -45 -1784 45 -1762
<< psubdiffcont >>
rect -23 -1762 23 1762
<< metal1 >>
rect -34 1762 34 1773
rect -34 -1762 -23 1762
rect 23 -1762 34 1762
rect -34 -1773 34 -1762
<< end >>
