magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -2053 -3233 3187 2569
<< nwell >>
rect 0 428 1060 569
rect 815 342 870 380
rect 397 -180 398 -151
rect 600 -242 725 -89
rect 145 -341 916 -337
<< pwell >>
rect 205 -475 206 -466
rect 217 -480 269 -442
rect 609 -1050 620 -442
<< pmos >>
rect 662 -180 663 -151
<< psubdiff >>
rect 58 -1162 787 -1141
rect 58 -1208 97 -1162
rect 143 -1208 297 -1162
rect 343 -1208 497 -1162
rect 543 -1208 697 -1162
rect 743 -1208 787 -1162
rect 58 -1223 787 -1208
<< nsubdiff >>
rect 58 529 816 545
rect 58 483 89 529
rect 135 483 289 529
rect 335 483 509 529
rect 555 483 729 529
rect 775 483 816 529
rect 58 469 816 483
rect 898 529 1016 545
rect 898 483 929 529
rect 975 483 1016 529
rect 898 469 1016 483
<< psubdiffcont >>
rect 97 -1208 143 -1162
rect 297 -1208 343 -1162
rect 497 -1208 543 -1162
rect 697 -1208 743 -1162
<< nsubdiffcont >>
rect 89 483 135 529
rect 289 483 335 529
rect 509 483 555 529
rect 729 483 775 529
rect 929 483 975 529
<< polysilicon >>
rect 174 342 886 394
rect 113 89 174 97
rect 113 83 274 89
rect 113 37 127 83
rect 173 37 274 83
rect 113 21 274 37
rect 786 -26 886 4
rect 786 -28 811 -26
rect 174 -72 811 -28
rect 857 -72 886 -26
rect 174 -81 886 -72
rect 192 -431 498 -418
rect 192 -466 220 -431
rect 205 -477 220 -466
rect 266 -466 498 -431
rect 266 -477 478 -466
rect 204 -490 478 -477
rect 490 -490 498 -466
rect 732 -770 832 -722
rect 212 -1017 264 -1016
rect 212 -1025 215 -1017
rect 192 -1063 215 -1025
rect 261 -1025 264 -1017
rect 261 -1063 832 -1025
rect 192 -1081 832 -1063
<< polycontact >>
rect 127 37 173 83
rect 811 -72 857 -26
rect 220 -477 266 -431
rect 215 -1063 261 -1017
<< metal1 >>
rect 0 529 1060 569
rect 0 483 89 529
rect 135 483 289 529
rect 335 483 509 529
rect 555 483 729 529
rect 775 483 929 529
rect 975 483 1060 529
rect 0 455 1060 483
rect 885 405 961 455
rect 99 355 961 405
rect 99 285 145 355
rect 507 285 553 355
rect 915 285 961 355
rect 270 246 369 265
rect 270 194 295 246
rect 347 194 369 246
rect 270 178 369 194
rect -52 83 185 85
rect -52 37 127 83
rect 173 37 185 83
rect -52 30 185 37
rect 303 84 349 132
rect 711 86 757 132
rect 711 84 886 86
rect 303 36 886 84
rect -52 -722 3 30
rect 786 -26 886 36
rect 302 -75 648 -26
rect 302 -288 351 -75
rect 599 -127 648 -75
rect 786 -72 811 -26
rect 857 -72 886 -26
rect 786 -80 886 -72
rect 599 -180 771 -127
rect 599 -226 701 -180
rect 663 -232 701 -226
rect 753 -195 771 -180
rect 1011 -178 1187 -155
rect 753 -232 770 -195
rect 663 -263 770 -232
rect 1011 -230 1030 -178
rect 1082 -230 1187 -178
rect 1011 -252 1187 -230
rect 99 -336 145 -290
rect 507 -336 553 -290
rect 915 -336 961 -290
rect 99 -382 961 -336
rect 205 -431 280 -429
rect 205 -477 220 -431
rect 266 -477 280 -431
rect 205 -490 280 -477
rect 81 -571 154 -558
rect 81 -623 98 -571
rect 150 -623 154 -571
rect 81 -635 154 -623
rect 211 -722 269 -490
rect 657 -540 703 -509
rect 329 -560 409 -542
rect 329 -612 338 -560
rect 390 -612 409 -560
rect 329 -629 409 -612
rect 494 -562 567 -549
rect 494 -614 510 -562
rect 562 -614 567 -562
rect 494 -626 567 -614
rect 657 -554 743 -540
rect 657 -606 675 -554
rect 727 -606 743 -554
rect 657 -620 743 -606
rect -52 -762 269 -722
rect -53 -770 269 -762
rect -53 -1026 -6 -770
rect 106 -860 212 -833
rect 657 -834 703 -620
rect 859 -665 906 -382
rect 859 -667 907 -665
rect 106 -912 127 -860
rect 179 -912 212 -860
rect 106 -932 212 -912
rect 510 -863 703 -834
rect 510 -915 535 -863
rect 587 -915 703 -863
rect 510 -927 703 -915
rect 205 -1017 273 -1003
rect 205 -1026 215 -1017
rect -53 -1063 215 -1026
rect 261 -1063 273 -1017
rect -53 -1073 273 -1063
rect 321 -1027 368 -953
rect 657 -977 703 -927
rect 860 -717 907 -667
rect 860 -763 1001 -717
rect 860 -953 906 -763
rect 861 -1027 908 -954
rect 321 -1067 908 -1027
rect 321 -1072 907 -1067
rect 321 -1075 906 -1072
rect 38 -1148 957 -1121
rect 38 -1162 770 -1148
rect 38 -1208 97 -1162
rect 143 -1208 297 -1162
rect 343 -1208 497 -1162
rect 543 -1208 697 -1162
rect 743 -1200 770 -1162
rect 822 -1200 957 -1148
rect 743 -1208 957 -1200
rect 38 -1233 957 -1208
<< via1 >>
rect 295 194 347 246
rect 701 -232 753 -180
rect 1030 -230 1082 -178
rect 98 -623 150 -571
rect 338 -612 390 -560
rect 510 -614 562 -562
rect 675 -606 727 -554
rect 127 -912 179 -860
rect 535 -915 587 -863
rect 770 -1200 822 -1148
<< metal2 >>
rect 270 265 375 270
rect 270 246 376 265
rect 270 194 295 246
rect 347 194 376 246
rect 270 191 376 194
rect 270 -298 375 191
rect 663 -178 1111 -151
rect 663 -180 1030 -178
rect 663 -232 701 -180
rect 753 -230 1030 -180
rect 1082 -230 1111 -178
rect 753 -232 1111 -230
rect 663 -264 1111 -232
rect 80 -404 583 -298
rect 80 -550 190 -404
rect 373 -405 583 -404
rect 81 -571 190 -550
rect 81 -623 98 -571
rect 150 -623 190 -571
rect 81 -635 190 -623
rect 327 -542 408 -535
rect 327 -560 409 -542
rect 327 -612 338 -560
rect 390 -612 409 -560
rect 327 -629 409 -612
rect 490 -562 583 -405
rect 490 -614 510 -562
rect 562 -614 583 -562
rect 327 -682 408 -629
rect 490 -635 583 -614
rect 666 -554 757 -264
rect 1015 -265 1111 -264
rect 666 -606 675 -554
rect 727 -606 757 -554
rect 666 -620 757 -606
rect 325 -707 408 -682
rect 325 -708 807 -707
rect 325 -763 828 -708
rect 106 -860 703 -834
rect 106 -912 127 -860
rect 179 -863 703 -860
rect 179 -912 535 -863
rect 106 -915 535 -912
rect 587 -915 703 -863
rect 106 -932 703 -915
rect 772 -1126 828 -763
rect 731 -1148 867 -1126
rect 731 -1200 770 -1148
rect 822 -1200 867 -1148
rect 731 -1223 867 -1200
use nmos_3p3_UKFAHE  nmos_3p3_UKFAHE_0
timestamp 1713185578
transform 1 0 243 0 1 -898
box -162 -152 162 152
use nmos_3p3_UKFAHE  nmos_3p3_UKFAHE_1
timestamp 1713185578
transform 1 0 447 0 1 -898
box -162 -152 162 152
use nmos_3p3_UKFAHE  nmos_3p3_UKFAHE_2
timestamp 1713185578
transform 1 0 782 0 1 -594
box -162 -152 162 152
use nmos_3p3_UKFAHE  nmos_3p3_UKFAHE_3
timestamp 1713185578
transform 1 0 782 0 1 -898
box -162 -152 162 152
use nmos_3p3_UKFAHE  nmos_3p3_UKFAHE_4
timestamp 1713185578
transform 1 0 447 0 1 -594
box -162 -152 162 152
use nmos_3p3_UKFAHE  nmos_3p3_UKFAHE_5
timestamp 1713185578
transform 1 0 243 0 1 -594
box -162 -152 162 152
use pmos_3p3_YMKZL5  pmos_3p3_YMKZL5_0
timestamp 1713185578
transform 1 0 428 0 1 -208
box -224 -214 224 214
use pmos_3p3_YMKZL5  pmos_3p3_YMKZL5_1
timestamp 1713185578
transform 1 0 632 0 1 -208
box -224 -214 224 214
use pmos_3p3_YMKZL5  pmos_3p3_YMKZL5_2
timestamp 1713185578
transform 1 0 836 0 1 -208
box -224 -214 224 214
use pmos_3p3_YMKZL5  pmos_3p3_YMKZL5_3
timestamp 1713185578
transform 1 0 224 0 1 -208
box -224 -214 224 214
use pmos_3p3_YMKZL5  pmos_3p3_YMKZL5_4
timestamp 1713185578
transform 1 0 836 0 1 214
box -224 -214 224 214
use pmos_3p3_YMKZL5  pmos_3p3_YMKZL5_5
timestamp 1713185578
transform 1 0 632 0 1 214
box -224 -214 224 214
use pmos_3p3_YMKZL5  pmos_3p3_YMKZL5_6
timestamp 1713185578
transform 1 0 428 0 1 214
box -224 -214 224 214
use pmos_3p3_YMKZL5  pmos_3p3_YMKZL5_7
timestamp 1713185578
transform 1 0 224 0 1 214
box -224 -214 224 214
<< labels >>
flabel psubdiffcont 514 -1187 514 -1187 0 FreeSans 750 0 0 0 VSS
flabel nsubdiffcont 533 506 533 506 0 FreeSans 1000 0 0 0 VDD
flabel metal1 s 1133 -218 1133 -218 0 FreeSans 750 0 0 0 OUT
port 1 nsew
flabel metal1 s 966 -741 966 -741 0 FreeSans 750 0 0 0 IN
port 2 nsew
flabel metal1 s -37 -344 -37 -344 0 FreeSans 750 0 0 0 CLK
port 3 nsew
<< end >>
