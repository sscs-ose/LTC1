magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2109 -2322 2109 2322
<< metal2 >>
rect -109 312 109 322
rect -109 256 -99 312
rect -43 256 43 312
rect 99 256 109 312
rect -109 170 109 256
rect -109 114 -99 170
rect -43 114 43 170
rect 99 114 109 170
rect -109 28 109 114
rect -109 -28 -99 28
rect -43 -28 43 28
rect 99 -28 109 28
rect -109 -114 109 -28
rect -109 -170 -99 -114
rect -43 -170 43 -114
rect 99 -170 109 -114
rect -109 -256 109 -170
rect -109 -312 -99 -256
rect -43 -312 43 -256
rect 99 -312 109 -256
rect -109 -322 109 -312
<< via2 >>
rect -99 256 -43 312
rect 43 256 99 312
rect -99 114 -43 170
rect 43 114 99 170
rect -99 -28 -43 28
rect 43 -28 99 28
rect -99 -170 -43 -114
rect 43 -170 99 -114
rect -99 -312 -43 -256
rect 43 -312 99 -256
<< metal3 >>
rect -109 312 109 322
rect -109 256 -99 312
rect -43 256 43 312
rect 99 256 109 312
rect -109 170 109 256
rect -109 114 -99 170
rect -43 114 43 170
rect 99 114 109 170
rect -109 28 109 114
rect -109 -28 -99 28
rect -43 -28 43 28
rect 99 -28 109 28
rect -109 -114 109 -28
rect -109 -170 -99 -114
rect -43 -170 43 -114
rect 99 -170 109 -114
rect -109 -256 109 -170
rect -109 -312 -99 -256
rect -43 -312 43 -256
rect 99 -312 109 -256
rect -109 -322 109 -312
<< end >>
