magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -4978 -2758 4978 2758
<< nwell >>
rect -2978 -758 2978 758
<< pmos >>
rect -2804 68 -2704 628
rect -2600 68 -2500 628
rect -2396 68 -2296 628
rect -2192 68 -2092 628
rect -1988 68 -1888 628
rect -1784 68 -1684 628
rect -1580 68 -1480 628
rect -1376 68 -1276 628
rect -1172 68 -1072 628
rect -968 68 -868 628
rect -764 68 -664 628
rect -560 68 -460 628
rect -356 68 -256 628
rect -152 68 -52 628
rect 52 68 152 628
rect 256 68 356 628
rect 460 68 560 628
rect 664 68 764 628
rect 868 68 968 628
rect 1072 68 1172 628
rect 1276 68 1376 628
rect 1480 68 1580 628
rect 1684 68 1784 628
rect 1888 68 1988 628
rect 2092 68 2192 628
rect 2296 68 2396 628
rect 2500 68 2600 628
rect 2704 68 2804 628
rect -2804 -628 -2704 -68
rect -2600 -628 -2500 -68
rect -2396 -628 -2296 -68
rect -2192 -628 -2092 -68
rect -1988 -628 -1888 -68
rect -1784 -628 -1684 -68
rect -1580 -628 -1480 -68
rect -1376 -628 -1276 -68
rect -1172 -628 -1072 -68
rect -968 -628 -868 -68
rect -764 -628 -664 -68
rect -560 -628 -460 -68
rect -356 -628 -256 -68
rect -152 -628 -52 -68
rect 52 -628 152 -68
rect 256 -628 356 -68
rect 460 -628 560 -68
rect 664 -628 764 -68
rect 868 -628 968 -68
rect 1072 -628 1172 -68
rect 1276 -628 1376 -68
rect 1480 -628 1580 -68
rect 1684 -628 1784 -68
rect 1888 -628 1988 -68
rect 2092 -628 2192 -68
rect 2296 -628 2396 -68
rect 2500 -628 2600 -68
rect 2704 -628 2804 -68
<< pdiff >>
rect -2892 606 -2804 628
rect -2892 90 -2879 606
rect -2833 90 -2804 606
rect -2892 68 -2804 90
rect -2704 606 -2600 628
rect -2704 90 -2675 606
rect -2629 90 -2600 606
rect -2704 68 -2600 90
rect -2500 606 -2396 628
rect -2500 90 -2471 606
rect -2425 90 -2396 606
rect -2500 68 -2396 90
rect -2296 606 -2192 628
rect -2296 90 -2267 606
rect -2221 90 -2192 606
rect -2296 68 -2192 90
rect -2092 606 -1988 628
rect -2092 90 -2063 606
rect -2017 90 -1988 606
rect -2092 68 -1988 90
rect -1888 606 -1784 628
rect -1888 90 -1859 606
rect -1813 90 -1784 606
rect -1888 68 -1784 90
rect -1684 606 -1580 628
rect -1684 90 -1655 606
rect -1609 90 -1580 606
rect -1684 68 -1580 90
rect -1480 606 -1376 628
rect -1480 90 -1451 606
rect -1405 90 -1376 606
rect -1480 68 -1376 90
rect -1276 606 -1172 628
rect -1276 90 -1247 606
rect -1201 90 -1172 606
rect -1276 68 -1172 90
rect -1072 606 -968 628
rect -1072 90 -1043 606
rect -997 90 -968 606
rect -1072 68 -968 90
rect -868 606 -764 628
rect -868 90 -839 606
rect -793 90 -764 606
rect -868 68 -764 90
rect -664 606 -560 628
rect -664 90 -635 606
rect -589 90 -560 606
rect -664 68 -560 90
rect -460 606 -356 628
rect -460 90 -431 606
rect -385 90 -356 606
rect -460 68 -356 90
rect -256 606 -152 628
rect -256 90 -227 606
rect -181 90 -152 606
rect -256 68 -152 90
rect -52 606 52 628
rect -52 90 -23 606
rect 23 90 52 606
rect -52 68 52 90
rect 152 606 256 628
rect 152 90 181 606
rect 227 90 256 606
rect 152 68 256 90
rect 356 606 460 628
rect 356 90 385 606
rect 431 90 460 606
rect 356 68 460 90
rect 560 606 664 628
rect 560 90 589 606
rect 635 90 664 606
rect 560 68 664 90
rect 764 606 868 628
rect 764 90 793 606
rect 839 90 868 606
rect 764 68 868 90
rect 968 606 1072 628
rect 968 90 997 606
rect 1043 90 1072 606
rect 968 68 1072 90
rect 1172 606 1276 628
rect 1172 90 1201 606
rect 1247 90 1276 606
rect 1172 68 1276 90
rect 1376 606 1480 628
rect 1376 90 1405 606
rect 1451 90 1480 606
rect 1376 68 1480 90
rect 1580 606 1684 628
rect 1580 90 1609 606
rect 1655 90 1684 606
rect 1580 68 1684 90
rect 1784 606 1888 628
rect 1784 90 1813 606
rect 1859 90 1888 606
rect 1784 68 1888 90
rect 1988 606 2092 628
rect 1988 90 2017 606
rect 2063 90 2092 606
rect 1988 68 2092 90
rect 2192 606 2296 628
rect 2192 90 2221 606
rect 2267 90 2296 606
rect 2192 68 2296 90
rect 2396 606 2500 628
rect 2396 90 2425 606
rect 2471 90 2500 606
rect 2396 68 2500 90
rect 2600 606 2704 628
rect 2600 90 2629 606
rect 2675 90 2704 606
rect 2600 68 2704 90
rect 2804 606 2892 628
rect 2804 90 2833 606
rect 2879 90 2892 606
rect 2804 68 2892 90
rect -2892 -90 -2804 -68
rect -2892 -606 -2879 -90
rect -2833 -606 -2804 -90
rect -2892 -628 -2804 -606
rect -2704 -90 -2600 -68
rect -2704 -606 -2675 -90
rect -2629 -606 -2600 -90
rect -2704 -628 -2600 -606
rect -2500 -90 -2396 -68
rect -2500 -606 -2471 -90
rect -2425 -606 -2396 -90
rect -2500 -628 -2396 -606
rect -2296 -90 -2192 -68
rect -2296 -606 -2267 -90
rect -2221 -606 -2192 -90
rect -2296 -628 -2192 -606
rect -2092 -90 -1988 -68
rect -2092 -606 -2063 -90
rect -2017 -606 -1988 -90
rect -2092 -628 -1988 -606
rect -1888 -90 -1784 -68
rect -1888 -606 -1859 -90
rect -1813 -606 -1784 -90
rect -1888 -628 -1784 -606
rect -1684 -90 -1580 -68
rect -1684 -606 -1655 -90
rect -1609 -606 -1580 -90
rect -1684 -628 -1580 -606
rect -1480 -90 -1376 -68
rect -1480 -606 -1451 -90
rect -1405 -606 -1376 -90
rect -1480 -628 -1376 -606
rect -1276 -90 -1172 -68
rect -1276 -606 -1247 -90
rect -1201 -606 -1172 -90
rect -1276 -628 -1172 -606
rect -1072 -90 -968 -68
rect -1072 -606 -1043 -90
rect -997 -606 -968 -90
rect -1072 -628 -968 -606
rect -868 -90 -764 -68
rect -868 -606 -839 -90
rect -793 -606 -764 -90
rect -868 -628 -764 -606
rect -664 -90 -560 -68
rect -664 -606 -635 -90
rect -589 -606 -560 -90
rect -664 -628 -560 -606
rect -460 -90 -356 -68
rect -460 -606 -431 -90
rect -385 -606 -356 -90
rect -460 -628 -356 -606
rect -256 -90 -152 -68
rect -256 -606 -227 -90
rect -181 -606 -152 -90
rect -256 -628 -152 -606
rect -52 -90 52 -68
rect -52 -606 -23 -90
rect 23 -606 52 -90
rect -52 -628 52 -606
rect 152 -90 256 -68
rect 152 -606 181 -90
rect 227 -606 256 -90
rect 152 -628 256 -606
rect 356 -90 460 -68
rect 356 -606 385 -90
rect 431 -606 460 -90
rect 356 -628 460 -606
rect 560 -90 664 -68
rect 560 -606 589 -90
rect 635 -606 664 -90
rect 560 -628 664 -606
rect 764 -90 868 -68
rect 764 -606 793 -90
rect 839 -606 868 -90
rect 764 -628 868 -606
rect 968 -90 1072 -68
rect 968 -606 997 -90
rect 1043 -606 1072 -90
rect 968 -628 1072 -606
rect 1172 -90 1276 -68
rect 1172 -606 1201 -90
rect 1247 -606 1276 -90
rect 1172 -628 1276 -606
rect 1376 -90 1480 -68
rect 1376 -606 1405 -90
rect 1451 -606 1480 -90
rect 1376 -628 1480 -606
rect 1580 -90 1684 -68
rect 1580 -606 1609 -90
rect 1655 -606 1684 -90
rect 1580 -628 1684 -606
rect 1784 -90 1888 -68
rect 1784 -606 1813 -90
rect 1859 -606 1888 -90
rect 1784 -628 1888 -606
rect 1988 -90 2092 -68
rect 1988 -606 2017 -90
rect 2063 -606 2092 -90
rect 1988 -628 2092 -606
rect 2192 -90 2296 -68
rect 2192 -606 2221 -90
rect 2267 -606 2296 -90
rect 2192 -628 2296 -606
rect 2396 -90 2500 -68
rect 2396 -606 2425 -90
rect 2471 -606 2500 -90
rect 2396 -628 2500 -606
rect 2600 -90 2704 -68
rect 2600 -606 2629 -90
rect 2675 -606 2704 -90
rect 2600 -628 2704 -606
rect 2804 -90 2892 -68
rect 2804 -606 2833 -90
rect 2879 -606 2892 -90
rect 2804 -628 2892 -606
<< pdiffc >>
rect -2879 90 -2833 606
rect -2675 90 -2629 606
rect -2471 90 -2425 606
rect -2267 90 -2221 606
rect -2063 90 -2017 606
rect -1859 90 -1813 606
rect -1655 90 -1609 606
rect -1451 90 -1405 606
rect -1247 90 -1201 606
rect -1043 90 -997 606
rect -839 90 -793 606
rect -635 90 -589 606
rect -431 90 -385 606
rect -227 90 -181 606
rect -23 90 23 606
rect 181 90 227 606
rect 385 90 431 606
rect 589 90 635 606
rect 793 90 839 606
rect 997 90 1043 606
rect 1201 90 1247 606
rect 1405 90 1451 606
rect 1609 90 1655 606
rect 1813 90 1859 606
rect 2017 90 2063 606
rect 2221 90 2267 606
rect 2425 90 2471 606
rect 2629 90 2675 606
rect 2833 90 2879 606
rect -2879 -606 -2833 -90
rect -2675 -606 -2629 -90
rect -2471 -606 -2425 -90
rect -2267 -606 -2221 -90
rect -2063 -606 -2017 -90
rect -1859 -606 -1813 -90
rect -1655 -606 -1609 -90
rect -1451 -606 -1405 -90
rect -1247 -606 -1201 -90
rect -1043 -606 -997 -90
rect -839 -606 -793 -90
rect -635 -606 -589 -90
rect -431 -606 -385 -90
rect -227 -606 -181 -90
rect -23 -606 23 -90
rect 181 -606 227 -90
rect 385 -606 431 -90
rect 589 -606 635 -90
rect 793 -606 839 -90
rect 997 -606 1043 -90
rect 1201 -606 1247 -90
rect 1405 -606 1451 -90
rect 1609 -606 1655 -90
rect 1813 -606 1859 -90
rect 2017 -606 2063 -90
rect 2221 -606 2267 -90
rect 2425 -606 2471 -90
rect 2629 -606 2675 -90
rect 2833 -606 2879 -90
<< polysilicon >>
rect -2804 628 -2704 672
rect -2600 628 -2500 672
rect -2396 628 -2296 672
rect -2192 628 -2092 672
rect -1988 628 -1888 672
rect -1784 628 -1684 672
rect -1580 628 -1480 672
rect -1376 628 -1276 672
rect -1172 628 -1072 672
rect -968 628 -868 672
rect -764 628 -664 672
rect -560 628 -460 672
rect -356 628 -256 672
rect -152 628 -52 672
rect 52 628 152 672
rect 256 628 356 672
rect 460 628 560 672
rect 664 628 764 672
rect 868 628 968 672
rect 1072 628 1172 672
rect 1276 628 1376 672
rect 1480 628 1580 672
rect 1684 628 1784 672
rect 1888 628 1988 672
rect 2092 628 2192 672
rect 2296 628 2396 672
rect 2500 628 2600 672
rect 2704 628 2804 672
rect -2804 24 -2704 68
rect -2600 24 -2500 68
rect -2396 24 -2296 68
rect -2192 24 -2092 68
rect -1988 24 -1888 68
rect -1784 24 -1684 68
rect -1580 24 -1480 68
rect -1376 24 -1276 68
rect -1172 24 -1072 68
rect -968 24 -868 68
rect -764 24 -664 68
rect -560 24 -460 68
rect -356 24 -256 68
rect -152 24 -52 68
rect 52 24 152 68
rect 256 24 356 68
rect 460 24 560 68
rect 664 24 764 68
rect 868 24 968 68
rect 1072 24 1172 68
rect 1276 24 1376 68
rect 1480 24 1580 68
rect 1684 24 1784 68
rect 1888 24 1988 68
rect 2092 24 2192 68
rect 2296 24 2396 68
rect 2500 24 2600 68
rect 2704 24 2804 68
rect -2804 -68 -2704 -24
rect -2600 -68 -2500 -24
rect -2396 -68 -2296 -24
rect -2192 -68 -2092 -24
rect -1988 -68 -1888 -24
rect -1784 -68 -1684 -24
rect -1580 -68 -1480 -24
rect -1376 -68 -1276 -24
rect -1172 -68 -1072 -24
rect -968 -68 -868 -24
rect -764 -68 -664 -24
rect -560 -68 -460 -24
rect -356 -68 -256 -24
rect -152 -68 -52 -24
rect 52 -68 152 -24
rect 256 -68 356 -24
rect 460 -68 560 -24
rect 664 -68 764 -24
rect 868 -68 968 -24
rect 1072 -68 1172 -24
rect 1276 -68 1376 -24
rect 1480 -68 1580 -24
rect 1684 -68 1784 -24
rect 1888 -68 1988 -24
rect 2092 -68 2192 -24
rect 2296 -68 2396 -24
rect 2500 -68 2600 -24
rect 2704 -68 2804 -24
rect -2804 -672 -2704 -628
rect -2600 -672 -2500 -628
rect -2396 -672 -2296 -628
rect -2192 -672 -2092 -628
rect -1988 -672 -1888 -628
rect -1784 -672 -1684 -628
rect -1580 -672 -1480 -628
rect -1376 -672 -1276 -628
rect -1172 -672 -1072 -628
rect -968 -672 -868 -628
rect -764 -672 -664 -628
rect -560 -672 -460 -628
rect -356 -672 -256 -628
rect -152 -672 -52 -628
rect 52 -672 152 -628
rect 256 -672 356 -628
rect 460 -672 560 -628
rect 664 -672 764 -628
rect 868 -672 968 -628
rect 1072 -672 1172 -628
rect 1276 -672 1376 -628
rect 1480 -672 1580 -628
rect 1684 -672 1784 -628
rect 1888 -672 1988 -628
rect 2092 -672 2192 -628
rect 2296 -672 2396 -628
rect 2500 -672 2600 -628
rect 2704 -672 2804 -628
<< metal1 >>
rect -2879 606 -2833 626
rect -2879 70 -2833 90
rect -2675 606 -2629 626
rect -2675 70 -2629 90
rect -2471 606 -2425 626
rect -2471 70 -2425 90
rect -2267 606 -2221 626
rect -2267 70 -2221 90
rect -2063 606 -2017 626
rect -2063 70 -2017 90
rect -1859 606 -1813 626
rect -1859 70 -1813 90
rect -1655 606 -1609 626
rect -1655 70 -1609 90
rect -1451 606 -1405 626
rect -1451 70 -1405 90
rect -1247 606 -1201 626
rect -1247 70 -1201 90
rect -1043 606 -997 626
rect -1043 70 -997 90
rect -839 606 -793 626
rect -839 70 -793 90
rect -635 606 -589 626
rect -635 70 -589 90
rect -431 606 -385 626
rect -431 70 -385 90
rect -227 606 -181 626
rect -227 70 -181 90
rect -23 606 23 626
rect -23 70 23 90
rect 181 606 227 626
rect 181 70 227 90
rect 385 606 431 626
rect 385 70 431 90
rect 589 606 635 626
rect 589 70 635 90
rect 793 606 839 626
rect 793 70 839 90
rect 997 606 1043 626
rect 997 70 1043 90
rect 1201 606 1247 626
rect 1201 70 1247 90
rect 1405 606 1451 626
rect 1405 70 1451 90
rect 1609 606 1655 626
rect 1609 70 1655 90
rect 1813 606 1859 626
rect 1813 70 1859 90
rect 2017 606 2063 626
rect 2017 70 2063 90
rect 2221 606 2267 626
rect 2221 70 2267 90
rect 2425 606 2471 626
rect 2425 70 2471 90
rect 2629 606 2675 626
rect 2629 70 2675 90
rect 2833 606 2879 626
rect 2833 70 2879 90
rect -2879 -90 -2833 -70
rect -2879 -626 -2833 -606
rect -2675 -90 -2629 -70
rect -2675 -626 -2629 -606
rect -2471 -90 -2425 -70
rect -2471 -626 -2425 -606
rect -2267 -90 -2221 -70
rect -2267 -626 -2221 -606
rect -2063 -90 -2017 -70
rect -2063 -626 -2017 -606
rect -1859 -90 -1813 -70
rect -1859 -626 -1813 -606
rect -1655 -90 -1609 -70
rect -1655 -626 -1609 -606
rect -1451 -90 -1405 -70
rect -1451 -626 -1405 -606
rect -1247 -90 -1201 -70
rect -1247 -626 -1201 -606
rect -1043 -90 -997 -70
rect -1043 -626 -997 -606
rect -839 -90 -793 -70
rect -839 -626 -793 -606
rect -635 -90 -589 -70
rect -635 -626 -589 -606
rect -431 -90 -385 -70
rect -431 -626 -385 -606
rect -227 -90 -181 -70
rect -227 -626 -181 -606
rect -23 -90 23 -70
rect -23 -626 23 -606
rect 181 -90 227 -70
rect 181 -626 227 -606
rect 385 -90 431 -70
rect 385 -626 431 -606
rect 589 -90 635 -70
rect 589 -626 635 -606
rect 793 -90 839 -70
rect 793 -626 839 -606
rect 997 -90 1043 -70
rect 997 -626 1043 -606
rect 1201 -90 1247 -70
rect 1201 -626 1247 -606
rect 1405 -90 1451 -70
rect 1405 -626 1451 -606
rect 1609 -90 1655 -70
rect 1609 -626 1655 -606
rect 1813 -90 1859 -70
rect 1813 -626 1859 -606
rect 2017 -90 2063 -70
rect 2017 -626 2063 -606
rect 2221 -90 2267 -70
rect 2221 -626 2267 -606
rect 2425 -90 2471 -70
rect 2425 -626 2471 -606
rect 2629 -90 2675 -70
rect 2629 -626 2675 -606
rect 2833 -90 2879 -70
rect 2833 -626 2879 -606
<< end >>
