magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1451 -1019 1451 1019
<< metal1 >>
rect -451 13 451 19
rect -451 -13 -445 13
rect -419 -13 -391 13
rect -365 -13 -337 13
rect -311 -13 -283 13
rect -257 -13 -229 13
rect -203 -13 -175 13
rect -149 -13 -121 13
rect -95 -13 -67 13
rect -41 -13 -13 13
rect 13 -13 41 13
rect 67 -13 95 13
rect 121 -13 149 13
rect 175 -13 203 13
rect 229 -13 257 13
rect 283 -13 311 13
rect 337 -13 365 13
rect 391 -13 419 13
rect 445 -13 451 13
rect -451 -19 451 -13
<< via1 >>
rect -445 -13 -419 13
rect -391 -13 -365 13
rect -337 -13 -311 13
rect -283 -13 -257 13
rect -229 -13 -203 13
rect -175 -13 -149 13
rect -121 -13 -95 13
rect -67 -13 -41 13
rect -13 -13 13 13
rect 41 -13 67 13
rect 95 -13 121 13
rect 149 -13 175 13
rect 203 -13 229 13
rect 257 -13 283 13
rect 311 -13 337 13
rect 365 -13 391 13
rect 419 -13 445 13
<< metal2 >>
rect -451 13 451 19
rect -451 -13 -445 13
rect -419 -13 -391 13
rect -365 -13 -337 13
rect -311 -13 -283 13
rect -257 -13 -229 13
rect -203 -13 -175 13
rect -149 -13 -121 13
rect -95 -13 -67 13
rect -41 -13 -13 13
rect 13 -13 41 13
rect 67 -13 95 13
rect 121 -13 149 13
rect 175 -13 203 13
rect 229 -13 257 13
rect 283 -13 311 13
rect 337 -13 365 13
rect 391 -13 419 13
rect 445 -13 451 13
rect -451 -19 451 -13
<< end >>
