magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2088 -2044 2960 2574
<< mvnmos >>
rect 0 0 140 530
rect 244 0 384 530
rect 488 0 628 530
rect 732 0 872 530
<< mvndiff >>
rect -88 517 0 530
rect -88 471 -75 517
rect -29 471 0 517
rect -88 403 0 471
rect -88 357 -75 403
rect -29 357 0 403
rect -88 289 0 357
rect -88 243 -75 289
rect -29 243 0 289
rect -88 174 0 243
rect -88 128 -75 174
rect -29 128 0 174
rect -88 59 0 128
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 140 517 244 530
rect 140 471 169 517
rect 215 471 244 517
rect 140 403 244 471
rect 140 357 169 403
rect 215 357 244 403
rect 140 289 244 357
rect 140 243 169 289
rect 215 243 244 289
rect 140 174 244 243
rect 140 128 169 174
rect 215 128 244 174
rect 140 59 244 128
rect 140 13 169 59
rect 215 13 244 59
rect 140 0 244 13
rect 384 517 488 530
rect 384 471 413 517
rect 459 471 488 517
rect 384 403 488 471
rect 384 357 413 403
rect 459 357 488 403
rect 384 289 488 357
rect 384 243 413 289
rect 459 243 488 289
rect 384 174 488 243
rect 384 128 413 174
rect 459 128 488 174
rect 384 59 488 128
rect 384 13 413 59
rect 459 13 488 59
rect 384 0 488 13
rect 628 517 732 530
rect 628 471 657 517
rect 703 471 732 517
rect 628 403 732 471
rect 628 357 657 403
rect 703 357 732 403
rect 628 289 732 357
rect 628 243 657 289
rect 703 243 732 289
rect 628 174 732 243
rect 628 128 657 174
rect 703 128 732 174
rect 628 59 732 128
rect 628 13 657 59
rect 703 13 732 59
rect 628 0 732 13
rect 872 517 960 530
rect 872 471 901 517
rect 947 471 960 517
rect 872 403 960 471
rect 872 357 901 403
rect 947 357 960 403
rect 872 289 960 357
rect 872 243 901 289
rect 947 243 960 289
rect 872 174 960 243
rect 872 128 901 174
rect 947 128 960 174
rect 872 59 960 128
rect 872 13 901 59
rect 947 13 960 59
rect 872 0 960 13
<< mvndiffc >>
rect -75 471 -29 517
rect -75 357 -29 403
rect -75 243 -29 289
rect -75 128 -29 174
rect -75 13 -29 59
rect 169 471 215 517
rect 169 357 215 403
rect 169 243 215 289
rect 169 128 215 174
rect 169 13 215 59
rect 413 471 459 517
rect 413 357 459 403
rect 413 243 459 289
rect 413 128 459 174
rect 413 13 459 59
rect 657 471 703 517
rect 657 357 703 403
rect 657 243 703 289
rect 657 128 703 174
rect 657 13 703 59
rect 901 471 947 517
rect 901 357 947 403
rect 901 243 947 289
rect 901 128 947 174
rect 901 13 947 59
<< polysilicon >>
rect 0 530 140 574
rect 244 530 384 574
rect 488 530 628 574
rect 732 530 872 574
rect 0 -44 140 0
rect 244 -44 384 0
rect 488 -44 628 0
rect 732 -44 872 0
<< metal1 >>
rect -75 517 -29 530
rect -75 403 -29 471
rect -75 289 -29 357
rect -75 174 -29 243
rect -75 59 -29 128
rect -75 0 -29 13
rect 169 517 215 530
rect 169 403 215 471
rect 169 289 215 357
rect 169 174 215 243
rect 169 59 215 128
rect 169 0 215 13
rect 413 517 459 530
rect 413 403 459 471
rect 413 289 459 357
rect 413 174 459 243
rect 413 59 459 128
rect 413 0 459 13
rect 657 517 703 530
rect 657 403 703 471
rect 657 289 703 357
rect 657 174 703 243
rect 657 59 703 128
rect 657 0 703 13
rect 901 517 947 530
rect 901 403 947 471
rect 901 289 947 357
rect 901 174 947 243
rect 901 59 947 128
rect 901 0 947 13
<< labels >>
rlabel mvndiffc 680 265 680 265 4 D
rlabel mvndiffc 436 265 436 265 4 S
rlabel mvndiffc 192 265 192 265 4 D
rlabel mvndiffc 924 265 924 265 4 S
rlabel mvndiffc -52 265 -52 265 4 S
<< end >>
