* NGSPICE file created from CM_64_flat.ext - technology: gf180mcuC

.subckt pex_CM_64 OUT IM_T IM VSS
X0 VSS IM.t1 a_424_490.t111 VSS.t11 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X1 OUT IM_T.t4 a_424_490.t19 VSS.t11 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X2 OUT IM_T.t5 a_424_490.t20 VSS.t12 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X3 VSS IM.t7 a_424_490.t105 VSS.t2 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=1u
X4 OUT IM_T.t8 a_424_490.t24 VSS.t13 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X5 VSS IM.t10 a_424_490.t102 VSS.t12 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X6 OUT IM_T.t11 a_424_490.t27 VSS.t2 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=1u
X7 OUT IM_T.t12 a_424_490.t13 VSS.t0 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X8 OUT IM_T.t14 a_424_490.t45 VSS.t1 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X9 VSS IM.t13 a_424_490.t99 VSS.t7 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X10 VSS IM.t14 a_424_490.t98 VSS.t1 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X11 VSS IM.t15 a_424_490.t97 VSS.t0 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X12 VSS IM.t16 a_424_490.t96 VSS.t1 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X13 OUT IM_T.t17 a_424_490.t41 VSS.t12 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X14 OUT IM_T.t18 a_424_490.t42 VSS.t12 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X15 OUT IM_T.t19 a_424_490.t0 VSS.t0 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X16 VSS IM.t19 a_424_490.t93 VSS.t2 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=1u
X17 VSS IM.t20 a_424_490.t92 VSS.t12 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X18 VSS IM.t22 a_424_490.t90 VSS.t6 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X19 OUT IM_T.t20 a_424_490.t1 VSS.t1 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X20 VSS IM.t23 a_424_490.t89 VSS.t12 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X21 OUT IM_T.t21 a_424_490.t47 VSS.t2 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=1u
X22 VSS IM.t24 a_424_490.t88 VSS.t11 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X23 VSS IM.t26 a_424_490.t86 VSS.t1 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X24 OUT IM_T.t25 a_424_490.t6 VSS.t6 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X25 VSS IM.t29 a_424_490.t83 VSS.t0 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X26 OUT IM_T.t26 a_424_490.t7 VSS.t6 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X27 VSS IM.t31 a_424_490.t81 VSS.t6 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X28 VSS IM.t32 a_424_490.t80 VSS.t13 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X29 OUT IM_T.t28 a_424_490.t43 VSS.t0 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X30 VSS IM.t34 a_424_490.t78 VSS.t6 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X31 OUT IM_T.t29 a_424_490.t44 VSS.t13 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X32 OUT IM_T.t30 a_424_490.t37 VSS.t1 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X33 OUT IM_T.t32 a_424_490.t28 VSS.t13 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X34 OUT IM_T.t33 a_424_490.t29 VSS.t7 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X35 VSS IM.t36 a_424_490.t76 VSS.t13 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X36 VSS IM.t37 a_424_490.t75 VSS.t1 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X37 OUT IM_T.t36 a_424_490.t116 VSS.t6 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X38 VSS IM.t39 a_424_490.t73 VSS.t13 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X39 OUT IM_T.t37 a_424_490.t117 VSS.t12 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X40 VSS IM.t41 a_424_490.t71 VSS.t2 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=1u
X41 VSS IM.t42 a_424_490.t70 VSS.t7 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X42 VSS IM.t43 a_424_490.t69 VSS.t6 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X43 OUT IM_T.t41 a_424_490.t35 VSS.t7 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X44 OUT IM_T.t42 a_424_490.t36 VSS.t11 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X45 VSS IM.t48 a_424_490.t64 VSS.t2 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=1u
X46 OUT IM_T.t46 a_424_490.t22 VSS.t13 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X47 VSS IM.t49 a_424_490.t63 VSS.t0 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X48 VSS IM.t50 a_424_490.t62 VSS.t11 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X49 VSS IM.t51 a_424_490.t61 VSS.t13 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X50 OUT IM_T.t50 a_424_490.t2 VSS.t2 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=1u
X51 VSS IM.t53 a_424_490.t59 VSS.t0 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X52 VSS IM.t55 a_424_490.t57 VSS.t7 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X53 OUT IM_T.t52 a_424_490.t31 VSS.t11 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X54 VSS IM.t56 a_424_490.t56 VSS.t7 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X55 OUT IM_T.t53 a_424_490.t113 VSS.t0 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X56 OUT IM_T.t55 a_424_490.t12 VSS.t1 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X57 OUT IM_T.t56 a_424_490.t9 VSS.t7 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X58 OUT IM_T.t57 a_424_490.t124 VSS.t7 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X59 VSS IM.t61 a_424_490.t51 VSS.t11 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X60 OUT IM_T.t60 a_424_490.t8 VSS.t6 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X61 OUT IM_T.t61 a_424_490.t125 VSS.t11 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X62 VSS IM.t63 a_424_490.t49 VSS.t12 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X63 OUT IM_T.t63 a_424_490.t34 VSS.t2 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=1u
R0 IM IM.n60 39.4161
R1 IM.n15 IM.n14 39.4095
R2 IM.n62 IM.n30 39.4095
R3 IM.n61 IM.n45 39.4095
R4 IM.n0 IM.t19 32.6004
R5 IM.n16 IM.t41 32.6004
R6 IM.n31 IM.t7 32.6004
R7 IM.n46 IM.t48 32.6004
R8 IM.n1 IM.n0 30.5194
R9 IM.n5 IM.n4 30.5194
R10 IM.n9 IM.n8 30.5194
R11 IM.n13 IM.n12 30.5194
R12 IM.n17 IM.n16 30.5194
R13 IM.n21 IM.n20 30.5194
R14 IM.n25 IM.n24 30.5194
R15 IM.n29 IM.n28 30.5194
R16 IM.n32 IM.n31 30.5194
R17 IM.n36 IM.n35 30.5194
R18 IM.n40 IM.n39 30.5194
R19 IM.n44 IM.n43 30.5194
R20 IM.n47 IM.n46 30.5194
R21 IM.n51 IM.n50 30.5194
R22 IM.n55 IM.n54 30.5194
R23 IM.n59 IM.n58 30.5194
R24 IM.n2 IM.n1 30.2907
R25 IM.n4 IM.n3 30.2907
R26 IM.n6 IM.n5 30.2907
R27 IM.n8 IM.n7 30.2907
R28 IM.n10 IM.n9 30.2907
R29 IM.n12 IM.n11 30.2907
R30 IM.n14 IM.n13 30.2907
R31 IM.n18 IM.n17 30.2907
R32 IM.n20 IM.n19 30.2907
R33 IM.n22 IM.n21 30.2907
R34 IM.n24 IM.n23 30.2907
R35 IM.n26 IM.n25 30.2907
R36 IM.n28 IM.n27 30.2907
R37 IM.n30 IM.n29 30.2907
R38 IM.n33 IM.n32 30.2907
R39 IM.n35 IM.n34 30.2907
R40 IM.n37 IM.n36 30.2907
R41 IM.n39 IM.n38 30.2907
R42 IM.n41 IM.n40 30.2907
R43 IM.n43 IM.n42 30.2907
R44 IM.n45 IM.n44 30.2907
R45 IM.n48 IM.n47 30.2907
R46 IM.n50 IM.n49 30.2907
R47 IM.n52 IM.n51 30.2907
R48 IM.n54 IM.n53 30.2907
R49 IM.n56 IM.n55 30.2907
R50 IM.n58 IM.n57 30.2907
R51 IM.n60 IM.n59 30.2907
R52 IM.n3 IM.n2 30.0619
R53 IM.n7 IM.n6 30.0619
R54 IM.n11 IM.n10 30.0619
R55 IM.n19 IM.n18 30.0619
R56 IM.n23 IM.n22 30.0619
R57 IM.n27 IM.n26 30.0619
R58 IM.n34 IM.n33 30.0619
R59 IM.n38 IM.n37 30.0619
R60 IM.n42 IM.n41 30.0619
R61 IM.n49 IM.n48 30.0619
R62 IM.n53 IM.n52 30.0619
R63 IM.n57 IM.n56 30.0619
R64 IM.n0 IM.t8 2.1905
R65 IM.n1 IM.t37 2.1905
R66 IM.n2 IM.t62 2.1905
R67 IM.n3 IM.t29 2.1905
R68 IM.n4 IM.t17 2.1905
R69 IM.n5 IM.t43 2.1905
R70 IM.n6 IM.t9 2.1905
R71 IM.n7 IM.t56 2.1905
R72 IM.n8 IM.t27 2.1905
R73 IM.n9 IM.t51 2.1905
R74 IM.n10 IM.t35 2.1905
R75 IM.n11 IM.t1 2.1905
R76 IM.n12 IM.t54 2.1905
R77 IM.n13 IM.t23 2.1905
R78 IM.n14 IM.t2 2.1905
R79 IM.n16 IM.t47 2.1905
R80 IM.n17 IM.t16 2.1905
R81 IM.n18 IM.t18 2.1905
R82 IM.n19 IM.t49 2.1905
R83 IM.n20 IM.t60 2.1905
R84 IM.n21 IM.t22 2.1905
R85 IM.n22 IM.t30 2.1905
R86 IM.n23 IM.t13 2.1905
R87 IM.n24 IM.t4 2.1905
R88 IM.n25 IM.t32 2.1905
R89 IM.n26 IM.t57 2.1905
R90 IM.n27 IM.t24 2.1905
R91 IM.n28 IM.t33 2.1905
R92 IM.n29 IM.t63 2.1905
R93 IM.n30 IM.t25 2.1905
R94 IM.n31 IM.t59 2.1905
R95 IM.n32 IM.t26 2.1905
R96 IM.n33 IM.t46 2.1905
R97 IM.n34 IM.t15 2.1905
R98 IM.n35 IM.t3 2.1905
R99 IM.n36 IM.t31 2.1905
R100 IM.n37 IM.t58 2.1905
R101 IM.n38 IM.t42 2.1905
R102 IM.n39 IM.t12 2.1905
R103 IM.n40 IM.t39 2.1905
R104 IM.n41 IM.t21 2.1905
R105 IM.n42 IM.t50 2.1905
R106 IM.n43 IM.t40 2.1905
R107 IM.n44 IM.t10 2.1905
R108 IM.n45 IM.t52 2.1905
R109 IM.n46 IM.t0 2.1905
R110 IM.n47 IM.t14 2.1905
R111 IM.n48 IM.t38 2.1905
R112 IM.n49 IM.t53 2.1905
R113 IM.n50 IM.t5 2.1905
R114 IM.n51 IM.t34 2.1905
R115 IM.n52 IM.t44 2.1905
R116 IM.n53 IM.t55 2.1905
R117 IM.n54 IM.t11 2.1905
R118 IM.n55 IM.t36 2.1905
R119 IM.n56 IM.t45 2.1905
R120 IM.n57 IM.t61 2.1905
R121 IM.n58 IM.t6 2.1905
R122 IM.n59 IM.t20 2.1905
R123 IM.n60 IM.t28 2.1905
R124 IM.n61 IM 1.61818
R125 IM.n62 IM 1.61818
R126 IM IM.n15 0.0659954
R127 IM.n15 IM 0.00703226
R128 IM IM.n61 0.00703226
R129 IM IM.n62 0.00703226
R130 VSS.n174 VSS.t2 73.1772
R131 VSS.n217 VSS.t13 51.4363
R132 VSS.n240 VSS.t1 41.8915
R133 VSS.n187 VSS.t10 39.2402
R134 VSS.n207 VSS.t12 36.5889
R135 VSS.n1 VSS.t6 33.9375
R136 VSS.n17 VSS.t8 29.6954
R137 VSS.n220 VSS.t14 27.0441
R138 VSS.n227 VSS.t5 21.7414
R139 VSS.n9 VSS.t9 19.0901
R140 VSS.n243 VSS.t3 17.4993
R141 VSS.n184 VSS.t0 14.8479
R142 VSS.n204 VSS.t15 12.1966
R143 VSS.n326 VSS.n25 11.6672
R144 VSS.n181 VSS.t4 9.54529
R145 VSS.n125 VSS.t26 6.55042
R146 VSS.n261 VSS.t75 6.55042
R147 VSS.n206 VSS.t108 6.55042
R148 VSS.n56 VSS.t72 6.55042
R149 VSS.n83 VSS.n47 6.52684
R150 VSS.n156 VSS.n155 6.50224
R151 VSS.n252 VSS.n251 6.50224
R152 VSS.n196 VSS.n195 6.50224
R153 VSS.n14 VSS.t11 5.30316
R154 VSS.n93 VSS.n91 3.85174
R155 VSS.n312 VSS.n311 3.85174
R156 VSS.n35 VSS.n33 3.85174
R157 VSS.n11 VSS.n7 3.85174
R158 VSS.n100 VSS.n89 3.80202
R159 VSS.n103 VSS.n87 3.80202
R160 VSS.n112 VSS.n85 3.80202
R161 VSS.n318 VSS.n309 3.80202
R162 VSS.n305 VSS.n44 3.80202
R163 VSS.n296 VSS.n46 3.80202
R164 VSS.n41 VSS.n31 3.80202
R165 VSS.n162 VSS.n161 3.80202
R166 VSS.n171 VSS.n159 3.80202
R167 VSS.n23 VSS.n5 3.80202
R168 VSS.n180 VSS.n179 3.80202
R169 VSS.n193 VSS.n177 3.80202
R170 VSS.n146 VSS.n119 3.75507
R171 VSS.n139 VSS.n121 3.75507
R172 VSS.n130 VSS.n123 3.75507
R173 VSS.n282 VSS.n255 3.75507
R174 VSS.n275 VSS.n257 3.75507
R175 VSS.n266 VSS.n259 3.75507
R176 VSS.n236 VSS.n199 3.75507
R177 VSS.n226 VSS.n201 3.75507
R178 VSS.n213 VSS.n203 3.75507
R179 VSS.n77 VSS.n50 3.75507
R180 VSS.n70 VSS.n52 3.75507
R181 VSS.n61 VSS.n54 3.75507
R182 VSS.n91 VSS.t104 2.7305
R183 VSS.n91 VSS.n90 2.7305
R184 VSS.n89 VSS.t97 2.7305
R185 VSS.n89 VSS.n88 2.7305
R186 VSS.n87 VSS.t105 2.7305
R187 VSS.n87 VSS.n86 2.7305
R188 VSS.n85 VSS.t111 2.7305
R189 VSS.n85 VSS.n84 2.7305
R190 VSS.n119 VSS.t40 2.7305
R191 VSS.n119 VSS.n118 2.7305
R192 VSS.n121 VSS.t24 2.7305
R193 VSS.n121 VSS.n120 2.7305
R194 VSS.n123 VSS.t81 2.7305
R195 VSS.n123 VSS.n122 2.7305
R196 VSS.n311 VSS.t51 2.7305
R197 VSS.n311 VSS.n310 2.7305
R198 VSS.n309 VSS.t96 2.7305
R199 VSS.n309 VSS.n308 2.7305
R200 VSS.n44 VSS.t107 2.7305
R201 VSS.n44 VSS.n43 2.7305
R202 VSS.n46 VSS.t23 2.7305
R203 VSS.n46 VSS.n45 2.7305
R204 VSS.n255 VSS.t86 2.7305
R205 VSS.n255 VSS.n254 2.7305
R206 VSS.n257 VSS.t69 2.7305
R207 VSS.n257 VSS.n256 2.7305
R208 VSS.n259 VSS.t17 2.7305
R209 VSS.n259 VSS.n258 2.7305
R210 VSS.n33 VSS.t62 2.7305
R211 VSS.n33 VSS.n32 2.7305
R212 VSS.n31 VSS.t106 2.7305
R213 VSS.n31 VSS.n30 2.7305
R214 VSS.n161 VSS.t22 2.7305
R215 VSS.n161 VSS.n160 2.7305
R216 VSS.n159 VSS.t43 2.7305
R217 VSS.n159 VSS.n158 2.7305
R218 VSS.n199 VSS.t19 2.7305
R219 VSS.n199 VSS.n198 2.7305
R220 VSS.n201 VSS.t99 2.7305
R221 VSS.n201 VSS.n200 2.7305
R222 VSS.n203 VSS.t59 2.7305
R223 VSS.n203 VSS.n202 2.7305
R224 VSS.n50 VSS.t54 2.7305
R225 VSS.n50 VSS.n49 2.7305
R226 VSS.n52 VSS.t44 2.7305
R227 VSS.n52 VSS.n51 2.7305
R228 VSS.n54 VSS.t41 2.7305
R229 VSS.n54 VSS.n53 2.7305
R230 VSS.n7 VSS.t30 2.7305
R231 VSS.n7 VSS.n6 2.7305
R232 VSS.n5 VSS.t73 2.7305
R233 VSS.n5 VSS.n4 2.7305
R234 VSS.n179 VSS.t88 2.7305
R235 VSS.n179 VSS.n178 2.7305
R236 VSS.n177 VSS.t101 2.7305
R237 VSS.n177 VSS.n176 2.7305
R238 VSS.n223 VSS.t7 2.65183
R239 VSS.n242 VSS.n241 2.6005
R240 VSS.n241 VSS.n240 2.6005
R241 VSS.n239 VSS.n238 2.6005
R242 VSS.n238 VSS.n237 2.6005
R243 VSS.n235 VSS.n234 2.6005
R244 VSS.n234 VSS.n233 2.6005
R245 VSS.n232 VSS.n231 2.6005
R246 VSS.n231 VSS.n230 2.6005
R247 VSS.n229 VSS.n228 2.6005
R248 VSS.n228 VSS.n227 2.6005
R249 VSS.n225 VSS.n224 2.6005
R250 VSS.n224 VSS.n223 2.6005
R251 VSS.n222 VSS.n221 2.6005
R252 VSS.n221 VSS.n220 2.6005
R253 VSS.n219 VSS.n218 2.6005
R254 VSS.n218 VSS.n217 2.6005
R255 VSS.n216 VSS.n215 2.6005
R256 VSS.n215 VSS.n214 2.6005
R257 VSS.n212 VSS.n211 2.6005
R258 VSS.n211 VSS.n210 2.6005
R259 VSS.n209 VSS.n208 2.6005
R260 VSS.n208 VSS.n207 2.6005
R261 VSS.n206 VSS.n205 2.6005
R262 VSS.n205 VSS.n204 2.6005
R263 VSS.n245 VSS.n244 2.6005
R264 VSS.n244 VSS.n243 2.6005
R265 VSS.n173 VSS.n172 2.6005
R266 VSS.n170 VSS.n169 2.6005
R267 VSS.n168 VSS.n167 2.6005
R268 VSS.n166 VSS.n165 2.6005
R269 VSS.n164 VSS.n163 2.6005
R270 VSS.n29 VSS.n28 2.6005
R271 VSS.n324 VSS 2.6005
R272 VSS.n325 VSS.n324 2.6005
R273 VSS.n323 VSS.n322 2.6005
R274 VSS.n322 VSS.n321 2.6005
R275 VSS.n40 VSS.n39 2.6005
R276 VSS.n38 VSS.n37 2.6005
R277 VSS.n14 VSS.n13 2.6005
R278 VSS.n35 VSS.n34 2.6005
R279 VSS.n286 VSS.n285 2.6005
R280 VSS.n284 VSS.n283 2.6005
R281 VSS.n281 VSS.n280 2.6005
R282 VSS.n279 VSS.n278 2.6005
R283 VSS.n277 VSS.n276 2.6005
R284 VSS.n274 VSS.n273 2.6005
R285 VSS.n272 VSS.n271 2.6005
R286 VSS.n270 VSS.n269 2.6005
R287 VSS.n268 VSS.n267 2.6005
R288 VSS.n265 VSS.n264 2.6005
R289 VSS.n263 VSS.n262 2.6005
R290 VSS.n261 VSS.n260 2.6005
R291 VSS.n288 VSS.n287 2.6005
R292 VSS.n295 VSS.n294 2.6005
R293 VSS.n298 VSS.n297 2.6005
R294 VSS.n300 VSS.n299 2.6005
R295 VSS.n302 VSS.n301 2.6005
R296 VSS.n304 VSS.n303 2.6005
R297 VSS.n307 VSS.n306 2.6005
R298 VSS VSS.n27 2.6005
R299 VSS.n325 VSS.n27 2.6005
R300 VSS.n320 VSS.n319 2.6005
R301 VSS.n321 VSS.n320 2.6005
R302 VSS.n317 VSS.n316 2.6005
R303 VSS.n315 VSS.n314 2.6005
R304 VSS.n14 VSS.n12 2.6005
R305 VSS.n9 VSS.n8 2.6005
R306 VSS.n150 VSS.n149 2.6005
R307 VSS.n148 VSS.n147 2.6005
R308 VSS.n145 VSS.n144 2.6005
R309 VSS.n143 VSS.n142 2.6005
R310 VSS.n141 VSS.n140 2.6005
R311 VSS.n138 VSS.n137 2.6005
R312 VSS.n136 VSS.n135 2.6005
R313 VSS.n134 VSS.n133 2.6005
R314 VSS.n132 VSS.n131 2.6005
R315 VSS.n129 VSS.n128 2.6005
R316 VSS.n127 VSS.n126 2.6005
R317 VSS.n125 VSS.n124 2.6005
R318 VSS.n152 VSS.n151 2.6005
R319 VSS.n114 VSS.n113 2.6005
R320 VSS.n111 VSS.n110 2.6005
R321 VSS.n109 VSS.n108 2.6005
R322 VSS.n107 VSS.n106 2.6005
R323 VSS.n105 VSS.n104 2.6005
R324 VSS.n1 VSS.n0 2.6005
R325 VSS VSS.n26 2.6005
R326 VSS.n325 VSS.n26 2.6005
R327 VSS.n101 VSS.n42 2.6005
R328 VSS.n321 VSS.n42 2.6005
R329 VSS.n99 VSS.n98 2.6005
R330 VSS.n97 VSS.n96 2.6005
R331 VSS.n95 VSS.n94 2.6005
R332 VSS.n93 VSS.n92 2.6005
R333 VSS.n80 VSS.n48 2.6005
R334 VSS.n79 VSS.n78 2.6005
R335 VSS.n76 VSS.n75 2.6005
R336 VSS.n74 VSS.n73 2.6005
R337 VSS.n72 VSS.n71 2.6005
R338 VSS.n69 VSS.n68 2.6005
R339 VSS.n67 VSS.n66 2.6005
R340 VSS.n65 VSS.n64 2.6005
R341 VSS.n63 VSS.n62 2.6005
R342 VSS.n60 VSS.n59 2.6005
R343 VSS.n58 VSS.n57 2.6005
R344 VSS.n56 VSS.n55 2.6005
R345 VSS.n82 VSS.n81 2.6005
R346 VSS.n194 VSS.n175 2.6005
R347 VSS.n175 VSS.n174 2.6005
R348 VSS.n192 VSS.n191 2.6005
R349 VSS.n191 VSS.n190 2.6005
R350 VSS.n189 VSS.n188 2.6005
R351 VSS.n188 VSS.n187 2.6005
R352 VSS.n186 VSS.n185 2.6005
R353 VSS.n185 VSS.n184 2.6005
R354 VSS.n183 VSS.n182 2.6005
R355 VSS.n182 VSS.n181 2.6005
R356 VSS.n3 VSS.n2 2.6005
R357 VSS.n2 VSS.n1 2.6005
R358 VSS VSS.n326 2.6005
R359 VSS.n326 VSS.n325 2.6005
R360 VSS.n25 VSS.n24 2.6005
R361 VSS.n321 VSS.n25 2.6005
R362 VSS.n22 VSS.n21 2.6005
R363 VSS.n21 VSS.n20 2.6005
R364 VSS.n19 VSS.n18 2.6005
R365 VSS.n18 VSS.n17 2.6005
R366 VSS.n16 VSS.n15 2.6005
R367 VSS.n15 VSS.n14 2.6005
R368 VSS.n11 VSS.n10 2.6005
R369 VSS.n10 VSS.n9 2.6005
R370 VSS.n154 VSS.n153 2.2505
R371 VSS.n157 VSS.n156 2.2505
R372 VSS.n290 VSS.n289 2.2505
R373 VSS.n253 VSS.n252 2.2505
R374 VSS.n247 VSS.n246 2.2505
R375 VSS.n197 VSS.n196 2.2505
R376 VSS.n197 VSS.n194 1.33855
R377 VSS.n115 VSS.n83 1.2659
R378 VSS.n293 VSS.n157 0.703183
R379 VSS.n253 VSS.n250 0.703183
R380 VSS.n115 VSS.n114 0.635926
R381 VSS.n295 VSS.n293 0.635926
R382 VSS.n250 VSS.n173 0.635926
R383 VSS.n111 VSS.n109 0.1505
R384 VSS.n109 VSS.n107 0.1505
R385 VSS.n107 VSS.n105 0.1505
R386 VSS.n102 VSS 0.1505
R387 VSS VSS.n101 0.1505
R388 VSS.n99 VSS.n97 0.1505
R389 VSS.n97 VSS.n95 0.1505
R390 VSS.n95 VSS.n93 0.1505
R391 VSS.n300 VSS.n298 0.1505
R392 VSS.n302 VSS.n300 0.1505
R393 VSS.n304 VSS.n302 0.1505
R394 VSS VSS.n307 0.1505
R395 VSS.n319 VSS 0.1505
R396 VSS.n317 VSS.n315 0.1505
R397 VSS.n315 VSS.n313 0.1505
R398 VSS.n313 VSS.n312 0.1505
R399 VSS.n170 VSS.n168 0.1505
R400 VSS.n168 VSS.n166 0.1505
R401 VSS.n166 VSS.n164 0.1505
R402 VSS VSS.n29 0.1505
R403 VSS VSS.n323 0.1505
R404 VSS.n40 VSS.n38 0.1505
R405 VSS.n38 VSS.n36 0.1505
R406 VSS.n36 VSS.n35 0.1505
R407 VSS.n192 VSS.n189 0.1505
R408 VSS.n189 VSS.n186 0.1505
R409 VSS.n186 VSS.n183 0.1505
R410 VSS VSS.n3 0.1505
R411 VSS.n22 VSS.n19 0.1505
R412 VSS.n19 VSS.n16 0.1505
R413 VSS.n16 VSS.n11 0.1505
R414 VSS.n24 VSS 0.150071
R415 VSS.n83 VSS.n82 0.142302
R416 VSS.n114 VSS.n112 0.136786
R417 VSS.n296 VSS.n295 0.136786
R418 VSS.n173 VSS.n171 0.136786
R419 VSS.n194 VSS.n193 0.136786
R420 VSS.n152 VSS.n150 0.131205
R421 VSS.n150 VSS.n148 0.131205
R422 VSS.n145 VSS.n143 0.131205
R423 VSS.n143 VSS.n141 0.131205
R424 VSS.n138 VSS.n136 0.131205
R425 VSS.n136 VSS.n134 0.131205
R426 VSS.n134 VSS.n132 0.131205
R427 VSS.n129 VSS.n127 0.131205
R428 VSS.n127 VSS.n125 0.131205
R429 VSS.n288 VSS.n286 0.131205
R430 VSS.n286 VSS.n284 0.131205
R431 VSS.n281 VSS.n279 0.131205
R432 VSS.n279 VSS.n277 0.131205
R433 VSS.n274 VSS.n272 0.131205
R434 VSS.n272 VSS.n270 0.131205
R435 VSS.n270 VSS.n268 0.131205
R436 VSS.n265 VSS.n263 0.131205
R437 VSS.n263 VSS.n261 0.131205
R438 VSS.n245 VSS.n242 0.131205
R439 VSS.n242 VSS.n239 0.131205
R440 VSS.n235 VSS.n232 0.131205
R441 VSS.n232 VSS.n229 0.131205
R442 VSS.n225 VSS.n222 0.131205
R443 VSS.n222 VSS.n219 0.131205
R444 VSS.n219 VSS.n216 0.131205
R445 VSS.n212 VSS.n209 0.131205
R446 VSS.n209 VSS.n206 0.131205
R447 VSS.n82 VSS.n80 0.131205
R448 VSS.n80 VSS.n79 0.131205
R449 VSS.n76 VSS.n74 0.131205
R450 VSS.n74 VSS.n72 0.131205
R451 VSS.n69 VSS.n67 0.131205
R452 VSS.n67 VSS.n65 0.131205
R453 VSS.n65 VSS.n63 0.131205
R454 VSS.n60 VSS.n58 0.131205
R455 VSS.n58 VSS.n56 0.131205
R456 VSS.n101 VSS.n100 0.129071
R457 VSS.n319 VSS.n318 0.129071
R458 VSS.n323 VSS.n41 0.129071
R459 VSS.n24 VSS.n23 0.129071
R460 VSS.n130 VSS.n129 0.127844
R461 VSS.n266 VSS.n265 0.127844
R462 VSS.n213 VSS.n212 0.127844
R463 VSS.n61 VSS.n60 0.127844
R464 VSS.n146 VSS.n145 0.121122
R465 VSS.n282 VSS.n281 0.121122
R466 VSS.n236 VSS.n235 0.121122
R467 VSS.n77 VSS.n76 0.121122
R468 VSS.n153 VSS.n152 0.117388
R469 VSS.n289 VSS.n288 0.117388
R470 VSS.n246 VSS.n245 0.117388
R471 VSS.n116 VSS.n115 0.106138
R472 VSS.n293 VSS.n292 0.106138
R473 VSS.n250 VSS.n249 0.106138
R474 VSS.n103 VSS.n102 0.0930714
R475 VSS.n307 VSS.n305 0.0930714
R476 VSS.n162 VSS.n29 0.0930714
R477 VSS.n180 VSS.n3 0.0930714
R478 VSS.n141 VSS.n139 0.0725747
R479 VSS.n277 VSS.n275 0.0725747
R480 VSS.n229 VSS.n226 0.0725747
R481 VSS.n72 VSS.n70 0.0725747
R482 VSS.n139 VSS.n138 0.0591307
R483 VSS.n275 VSS.n274 0.0591307
R484 VSS.n226 VSS.n225 0.0591307
R485 VSS.n70 VSS.n69 0.0591307
R486 VSS.n105 VSS.n103 0.0579286
R487 VSS.n305 VSS.n304 0.0579286
R488 VSS.n164 VSS.n162 0.0579286
R489 VSS.n183 VSS.n180 0.0579286
R490 VSS.n154 VSS.n117 0.0419226
R491 VSS.n291 VSS.n290 0.0419226
R492 VSS.n248 VSS.n247 0.0419226
R493 VSS.n100 VSS.n99 0.0219286
R494 VSS.n318 VSS.n317 0.0219286
R495 VSS.n41 VSS.n40 0.0219286
R496 VSS.n23 VSS.n22 0.0219286
R497 VSS.n112 VSS.n111 0.0142143
R498 VSS.n298 VSS.n296 0.0142143
R499 VSS.n171 VSS.n170 0.0142143
R500 VSS.n193 VSS.n192 0.0142143
R501 VSS.n148 VSS.n146 0.010583
R502 VSS.n284 VSS.n282 0.010583
R503 VSS.n239 VSS.n236 0.010583
R504 VSS.n79 VSS.n77 0.010583
R505 VSS.n132 VSS.n130 0.003861
R506 VSS.n268 VSS.n266 0.003861
R507 VSS.n216 VSS.n213 0.003861
R508 VSS.n63 VSS.n61 0.003861
R509 VSS.n117 VSS.n116 0.00351255
R510 VSS.n292 VSS.n291 0.00351255
R511 VSS.n249 VSS.n248 0.00351255
R512 VSS.n157 VSS.n154 0.00162971
R513 VSS.n290 VSS.n253 0.00162971
R514 VSS.n247 VSS.n197 0.00162971
R515 a_424_490.n26 a_424_490.n20 3.22004
R516 a_424_490.n193 a_424_490.n1 3.07769
R517 a_424_490.n82 a_424_490.n81 3.07769
R518 a_424_490.n42 a_424_490.n41 3.07769
R519 a_424_490.n10 a_424_490.n9 3.07769
R520 a_424_490.n179 a_424_490.n178 2.93817
R521 a_424_490.n151 a_424_490.n150 2.93817
R522 a_424_490.n139 a_424_490.n138 2.93817
R523 a_424_490.n24 a_424_490.n23 2.87833
R524 a_424_490.n143 a_424_490.n142 2.87833
R525 a_424_490.n155 a_424_490.n154 2.87833
R526 a_424_490.n185 a_424_490.n184 2.87833
R527 a_424_490.n194 a_424_490.n193 2.80003
R528 a_424_490.n82 a_424_490.n79 2.79937
R529 a_424_490.n42 a_424_490.n39 2.79937
R530 a_424_490.n10 a_424_490.n7 2.79937
R531 a_424_490.n29 a_424_490.n14 2.79724
R532 a_424_490.n28 a_424_490.n16 2.79662
R533 a_424_490.n30 a_424_490.n12 2.79463
R534 a_424_490.n25 a_424_490.n22 2.79421
R535 a_424_490.n144 a_424_490.n141 2.79377
R536 a_424_490.n156 a_424_490.n153 2.79377
R537 a_424_490.n186 a_424_490.n183 2.79377
R538 a_424_490.n31 a_424_490.n5 2.79336
R539 a_424_490.n27 a_424_490.n18 2.79324
R540 a_424_490.n1 a_424_490.t64 2.7305
R541 a_424_490.n1 a_424_490.n0 2.7305
R542 a_424_490.n3 a_424_490.t45 2.7305
R543 a_424_490.n3 a_424_490.n2 2.7305
R544 a_424_490.n105 a_424_490.t59 2.7305
R545 a_424_490.n105 a_424_490.n104 2.7305
R546 a_424_490.n113 a_424_490.t7 2.7305
R547 a_424_490.n113 a_424_490.n112 2.7305
R548 a_424_490.n121 a_424_490.t57 2.7305
R549 a_424_490.n121 a_424_490.n120 2.7305
R550 a_424_490.n167 a_424_490.t44 2.7305
R551 a_424_490.n167 a_424_490.n166 2.7305
R552 a_424_490.n181 a_424_490.t51 2.7305
R553 a_424_490.n181 a_424_490.n180 2.7305
R554 a_424_490.n178 a_424_490.t125 2.7305
R555 a_424_490.n178 a_424_490.n177 2.7305
R556 a_424_490.n175 a_424_490.t62 2.7305
R557 a_424_490.n175 a_424_490.n174 2.7305
R558 a_424_490.n81 a_424_490.t105 2.7305
R559 a_424_490.n81 a_424_490.n80 2.7305
R560 a_424_490.n79 a_424_490.t27 2.7305
R561 a_424_490.n79 a_424_490.n78 2.7305
R562 a_424_490.n99 a_424_490.t1 2.7305
R563 a_424_490.n99 a_424_490.n98 2.7305
R564 a_424_490.n102 a_424_490.t98 2.7305
R565 a_424_490.n102 a_424_490.n101 2.7305
R566 a_424_490.n107 a_424_490.t97 2.7305
R567 a_424_490.n107 a_424_490.n106 2.7305
R568 a_424_490.n110 a_424_490.t113 2.7305
R569 a_424_490.n110 a_424_490.n109 2.7305
R570 a_424_490.n115 a_424_490.t6 2.7305
R571 a_424_490.n115 a_424_490.n114 2.7305
R572 a_424_490.n118 a_424_490.t78 2.7305
R573 a_424_490.n118 a_424_490.n117 2.7305
R574 a_424_490.n161 a_424_490.t70 2.7305
R575 a_424_490.n161 a_424_490.n160 2.7305
R576 a_424_490.n164 a_424_490.t124 2.7305
R577 a_424_490.n164 a_424_490.n163 2.7305
R578 a_424_490.n169 a_424_490.t28 2.7305
R579 a_424_490.n169 a_424_490.n168 2.7305
R580 a_424_490.n172 a_424_490.t76 2.7305
R581 a_424_490.n172 a_424_490.n171 2.7305
R582 a_424_490.n132 a_424_490.t73 2.7305
R583 a_424_490.n132 a_424_490.n131 2.7305
R584 a_424_490.n129 a_424_490.t24 2.7305
R585 a_424_490.n129 a_424_490.n128 2.7305
R586 a_424_490.n41 a_424_490.t71 2.7305
R587 a_424_490.n41 a_424_490.n40 2.7305
R588 a_424_490.n39 a_424_490.t34 2.7305
R589 a_424_490.n39 a_424_490.n38 2.7305
R590 a_424_490.n73 a_424_490.t12 2.7305
R591 a_424_490.n73 a_424_490.n72 2.7305
R592 a_424_490.n76 a_424_490.t86 2.7305
R593 a_424_490.n76 a_424_490.n75 2.7305
R594 a_424_490.n84 a_424_490.t63 2.7305
R595 a_424_490.n84 a_424_490.n83 2.7305
R596 a_424_490.n87 a_424_490.t0 2.7305
R597 a_424_490.n87 a_424_490.n86 2.7305
R598 a_424_490.n90 a_424_490.t8 2.7305
R599 a_424_490.n90 a_424_490.n89 2.7305
R600 a_424_490.n93 a_424_490.t81 2.7305
R601 a_424_490.n93 a_424_490.n92 2.7305
R602 a_424_490.n123 a_424_490.t99 2.7305
R603 a_424_490.n123 a_424_490.n122 2.7305
R604 a_424_490.n126 a_424_490.t35 2.7305
R605 a_424_490.n126 a_424_490.n125 2.7305
R606 a_424_490.n147 a_424_490.t88 2.7305
R607 a_424_490.n147 a_424_490.n146 2.7305
R608 a_424_490.n150 a_424_490.t31 2.7305
R609 a_424_490.n150 a_424_490.n149 2.7305
R610 a_424_490.n138 a_424_490.t36 2.7305
R611 a_424_490.n138 a_424_490.n137 2.7305
R612 a_424_490.n135 a_424_490.t111 2.7305
R613 a_424_490.n135 a_424_490.n134 2.7305
R614 a_424_490.n20 a_424_490.t19 2.7305
R615 a_424_490.n20 a_424_490.n19 2.7305
R616 a_424_490.n9 a_424_490.t93 2.7305
R617 a_424_490.n9 a_424_490.n8 2.7305
R618 a_424_490.n7 a_424_490.t47 2.7305
R619 a_424_490.n7 a_424_490.n6 2.7305
R620 a_424_490.n33 a_424_490.t37 2.7305
R621 a_424_490.n33 a_424_490.n32 2.7305
R622 a_424_490.n36 a_424_490.t96 2.7305
R623 a_424_490.n36 a_424_490.n35 2.7305
R624 a_424_490.n5 a_424_490.t75 2.7305
R625 a_424_490.n5 a_424_490.n4 2.7305
R626 a_424_490.n44 a_424_490.t83 2.7305
R627 a_424_490.n44 a_424_490.n43 2.7305
R628 a_424_490.n47 a_424_490.t13 2.7305
R629 a_424_490.n47 a_424_490.n46 2.7305
R630 a_424_490.n12 a_424_490.t43 2.7305
R631 a_424_490.n12 a_424_490.n11 2.7305
R632 a_424_490.n50 a_424_490.t116 2.7305
R633 a_424_490.n50 a_424_490.n49 2.7305
R634 a_424_490.n53 a_424_490.t90 2.7305
R635 a_424_490.n53 a_424_490.n52 2.7305
R636 a_424_490.n14 a_424_490.t69 2.7305
R637 a_424_490.n14 a_424_490.n13 2.7305
R638 a_424_490.n56 a_424_490.t56 2.7305
R639 a_424_490.n56 a_424_490.n55 2.7305
R640 a_424_490.n59 a_424_490.t29 2.7305
R641 a_424_490.n59 a_424_490.n58 2.7305
R642 a_424_490.n16 a_424_490.t9 2.7305
R643 a_424_490.n16 a_424_490.n15 2.7305
R644 a_424_490.n62 a_424_490.t22 2.7305
R645 a_424_490.n62 a_424_490.n61 2.7305
R646 a_424_490.n65 a_424_490.t80 2.7305
R647 a_424_490.n65 a_424_490.n64 2.7305
R648 a_424_490.n18 a_424_490.t61 2.7305
R649 a_424_490.n18 a_424_490.n17 2.7305
R650 a_424_490.n22 a_424_490.t89 2.7305
R651 a_424_490.n22 a_424_490.n21 2.7305
R652 a_424_490.n141 a_424_490.t49 2.7305
R653 a_424_490.n141 a_424_490.n140 2.7305
R654 a_424_490.n153 a_424_490.t102 2.7305
R655 a_424_490.n153 a_424_490.n152 2.7305
R656 a_424_490.n183 a_424_490.t92 2.7305
R657 a_424_490.n183 a_424_490.n182 2.7305
R658 a_424_490.n194 a_424_490.t2 2.7305
R659 a_424_490.n195 a_424_490.n194 2.7305
R660 a_424_490.n190 a_424_490.n113 2.68248
R661 a_424_490.n191 a_424_490.n105 2.68235
R662 a_424_490.n189 a_424_490.n121 2.67583
R663 a_424_490.n192 a_424_490.n3 2.67342
R664 a_424_490.n187 a_424_490.n181 2.67239
R665 a_424_490.n188 a_424_490.n167 2.67214
R666 a_424_490.n25 a_424_490.n24 2.66766
R667 a_424_490.n144 a_424_490.n143 2.66766
R668 a_424_490.n156 a_424_490.n155 2.66766
R669 a_424_490.n186 a_424_490.n185 2.66766
R670 a_424_490.n176 a_424_490.n175 2.56335
R671 a_424_490.n148 a_424_490.n147 2.56335
R672 a_424_490.n136 a_424_490.n135 2.56335
R673 a_424_490.n170 a_424_490.n169 2.56317
R674 a_424_490.n130 a_424_490.n129 2.56317
R675 a_424_490.n63 a_424_490.n62 2.56317
R676 a_424_490.n100 a_424_490.n99 2.56299
R677 a_424_490.n74 a_424_490.n73 2.56299
R678 a_424_490.n34 a_424_490.n33 2.56299
R679 a_424_490.n119 a_424_490.n118 2.56281
R680 a_424_490.n165 a_424_490.n164 2.56281
R681 a_424_490.n94 a_424_490.n93 2.56281
R682 a_424_490.n127 a_424_490.n126 2.56281
R683 a_424_490.n54 a_424_490.n53 2.56281
R684 a_424_490.n60 a_424_490.n59 2.56281
R685 a_424_490.n108 a_424_490.n107 2.56272
R686 a_424_490.n116 a_424_490.n115 2.56272
R687 a_424_490.n85 a_424_490.n84 2.56272
R688 a_424_490.n91 a_424_490.n90 2.56272
R689 a_424_490.n45 a_424_490.n44 2.56272
R690 a_424_490.n51 a_424_490.n50 2.56272
R691 a_424_490.n162 a_424_490.n161 2.56263
R692 a_424_490.n124 a_424_490.n123 2.56263
R693 a_424_490.n57 a_424_490.n56 2.56263
R694 a_424_490.n103 a_424_490.n102 2.56245
R695 a_424_490.n111 a_424_490.n110 2.56245
R696 a_424_490.n173 a_424_490.n172 2.56245
R697 a_424_490.n133 a_424_490.n132 2.56245
R698 a_424_490.n77 a_424_490.n76 2.56245
R699 a_424_490.n88 a_424_490.n87 2.56245
R700 a_424_490.n37 a_424_490.n36 2.56245
R701 a_424_490.n48 a_424_490.n47 2.56245
R702 a_424_490.n66 a_424_490.n65 2.56245
R703 a_424_490.n24 a_424_490.t42 2.4382
R704 a_424_490.n143 a_424_490.t117 2.4382
R705 a_424_490.n155 a_424_490.t20 2.4382
R706 a_424_490.n185 a_424_490.t41 2.4382
R707 a_424_490.n173 a_424_490.n170 1.66688
R708 a_424_490.n66 a_424_490.n63 1.66688
R709 a_424_490.n133 a_424_490.n130 1.66688
R710 a_424_490.n103 a_424_490.n100 1.66543
R711 a_424_490.n77 a_424_490.n74 1.66543
R712 a_424_490.n37 a_424_490.n34 1.66543
R713 a_424_490.n151 a_424_490.n148 1.66252
R714 a_424_490.n139 a_424_490.n136 1.66252
R715 a_424_490.n179 a_424_490.n176 1.66252
R716 a_424_490.n165 a_424_490.n162 1.65962
R717 a_424_490.n127 a_424_490.n124 1.65962
R718 a_424_490.n60 a_424_490.n57 1.65962
R719 a_424_490.n111 a_424_490.n108 1.65672
R720 a_424_490.n88 a_424_490.n85 1.65672
R721 a_424_490.n48 a_424_490.n45 1.65672
R722 a_424_490.n119 a_424_490.n116 1.65381
R723 a_424_490.n94 a_424_490.n91 1.65381
R724 a_424_490.n54 a_424_490.n51 1.65381
R725 a_424_490.n26 a_424_490.n25 0.890339
R726 a_424_490.n145 a_424_490.n144 0.890339
R727 a_424_490.n157 a_424_490.n156 0.890339
R728 a_424_490.n187 a_424_490.n186 0.890339
R729 a_424_490.n30 a_424_490.n29 0.888887
R730 a_424_490.n70 a_424_490.n69 0.888887
R731 a_424_490.n96 a_424_490.n95 0.888887
R732 a_424_490.n191 a_424_490.n190 0.888887
R733 a_424_490.n28 a_424_490.n27 0.887435
R734 a_424_490.n68 a_424_490.n67 0.887435
R735 a_424_490.n159 a_424_490.n158 0.887435
R736 a_424_490.n189 a_424_490.n188 0.887435
R737 a_424_490.n31 a_424_490.n10 0.883081
R738 a_424_490.n71 a_424_490.n42 0.883081
R739 a_424_490.n97 a_424_490.n82 0.883081
R740 a_424_490.n193 a_424_490.n192 0.883081
R741 a_424_490.n31 a_424_490.n30 0.880177
R742 a_424_490.n71 a_424_490.n70 0.880177
R743 a_424_490.n97 a_424_490.n96 0.880177
R744 a_424_490.n192 a_424_490.n191 0.880177
R745 a_424_490.n29 a_424_490.n28 0.878726
R746 a_424_490.n69 a_424_490.n68 0.878726
R747 a_424_490.n190 a_424_490.n189 0.878726
R748 a_424_490.n27 a_424_490.n26 0.874371
R749 a_424_490.n158 a_424_490.n157 0.874371
R750 a_424_490.n188 a_424_490.n187 0.874371
R751 a_424_490.n157 a_424_490.n151 0.282373
R752 a_424_490.n145 a_424_490.n139 0.282373
R753 a_424_490.n187 a_424_490.n179 0.282373
R754 a_424_490.n190 a_424_490.n119 0.27947
R755 a_424_490.n189 a_424_490.n165 0.27947
R756 a_424_490.n95 a_424_490.n94 0.27947
R757 a_424_490.n159 a_424_490.n127 0.27947
R758 a_424_490.n69 a_424_490.n54 0.27947
R759 a_424_490.n68 a_424_490.n60 0.27947
R760 a_424_490.n192 a_424_490.n103 0.276567
R761 a_424_490.n191 a_424_490.n111 0.276567
R762 a_424_490.n188 a_424_490.n173 0.276567
R763 a_424_490.n97 a_424_490.n77 0.276567
R764 a_424_490.n96 a_424_490.n88 0.276567
R765 a_424_490.n71 a_424_490.n37 0.276567
R766 a_424_490.n70 a_424_490.n48 0.276567
R767 a_424_490.n67 a_424_490.n66 0.276567
R768 a_424_490.n158 a_424_490.n133 0.276567
R769 a_424_490.n162 a_424_490.n159 0.161294
R770 a_424_490.n100 a_424_490.n97 0.158391
R771 a_424_490.n74 a_424_490.n71 0.158391
R772 a_424_490.n34 a_424_490.n31 0.158391
R773 a_424_490.n148 a_424_490.n145 0.155488
R774 IM_T.n8 IM_T.n7 147.633
R775 IM_T.n10 IM_T.n9 147.633
R776 IM_T.n12 IM_T.n11 147.633
R777 IM_T.n23 IM_T.n22 147.633
R778 IM_T.n25 IM_T.n24 147.633
R779 IM_T.n27 IM_T.n26 147.633
R780 IM_T.n37 IM_T.n36 147.633
R781 IM_T.n39 IM_T.n38 147.633
R782 IM_T.n41 IM_T.n40 147.633
R783 IM_T.n51 IM_T.n50 147.633
R784 IM_T.n53 IM_T.n52 147.633
R785 IM_T.n55 IM_T.n54 147.633
R786 IM_T.n0 IM_T.t21 60.7907
R787 IM_T.n15 IM_T.t63 60.7907
R788 IM_T.n29 IM_T.t11 60.7907
R789 IM_T.n43 IM_T.t50 60.7907
R790 IM_T.n2 IM_T.n1 54.4633
R791 IM_T.n4 IM_T.n3 54.4633
R792 IM_T.n17 IM_T.n16 54.4633
R793 IM_T.n19 IM_T.n18 54.4633
R794 IM_T.n31 IM_T.n30 54.4633
R795 IM_T.n33 IM_T.n32 54.4633
R796 IM_T.n45 IM_T.n44 54.4633
R797 IM_T.n47 IM_T.n46 54.4633
R798 IM_T.n21 IM_T.n20 51.6858
R799 IM_T.n35 IM_T.n34 51.6858
R800 IM_T.n49 IM_T.n48 51.6858
R801 IM_T.n6 IM_T.n5 51.6849
R802 IM_T IM_T.n56 44.1559
R803 IM_T.n14 IM_T.n13 43.3679
R804 IM_T.n58 IM_T.n28 43.3679
R805 IM_T.n57 IM_T.n42 43.3679
R806 IM_T.n7 IM_T.t3 33.0769
R807 IM_T.n22 IM_T.t24 33.0769
R808 IM_T.n36 IM_T.t51 33.0769
R809 IM_T.n50 IM_T.t58 33.0769
R810 IM_T.n9 IM_T.n8 27.6763
R811 IM_T.n11 IM_T.n10 27.6763
R812 IM_T.n13 IM_T.n12 27.6763
R813 IM_T.n24 IM_T.n23 27.6763
R814 IM_T.n26 IM_T.n25 27.6763
R815 IM_T.n28 IM_T.n27 27.6763
R816 IM_T.n38 IM_T.n37 27.6763
R817 IM_T.n40 IM_T.n39 27.6763
R818 IM_T.n42 IM_T.n41 27.6763
R819 IM_T.n52 IM_T.n51 27.6763
R820 IM_T.n54 IM_T.n53 27.6763
R821 IM_T.n56 IM_T.n55 27.6763
R822 IM_T.n1 IM_T.n0 12.9829
R823 IM_T.n3 IM_T.n2 12.9829
R824 IM_T.n5 IM_T.n4 12.9829
R825 IM_T.n16 IM_T.n15 12.9829
R826 IM_T.n18 IM_T.n17 12.9829
R827 IM_T.n20 IM_T.n19 12.9829
R828 IM_T.n30 IM_T.n29 12.9829
R829 IM_T.n32 IM_T.n31 12.9829
R830 IM_T.n34 IM_T.n33 12.9829
R831 IM_T.n44 IM_T.n43 12.9829
R832 IM_T.n46 IM_T.n45 12.9829
R833 IM_T.n48 IM_T.n47 12.9829
R834 IM_T.n21 IM_T.t44 8.96618
R835 IM_T.n35 IM_T.t54 8.96618
R836 IM_T.n49 IM_T.t27 8.96618
R837 IM_T.n6 IM_T.t7 8.96331
R838 IM_T IM_T.n21 3.31674
R839 IM_T IM_T.n35 3.31674
R840 IM_T IM_T.n49 3.31674
R841 IM_T IM_T.n6 3.31651
R842 IM_T.n0 IM_T.t0 2.1905
R843 IM_T.n1 IM_T.t28 2.1905
R844 IM_T.n2 IM_T.t13 2.1905
R845 IM_T.n3 IM_T.t56 2.1905
R846 IM_T.n4 IM_T.t34 2.1905
R847 IM_T.n5 IM_T.t4 2.1905
R848 IM_T.n7 IM_T.t30 2.1905
R849 IM_T.n8 IM_T.t15 2.1905
R850 IM_T.n9 IM_T.t36 2.1905
R851 IM_T.n10 IM_T.t22 2.1905
R852 IM_T.n11 IM_T.t46 2.1905
R853 IM_T.n12 IM_T.t47 2.1905
R854 IM_T.n13 IM_T.t18 2.1905
R855 IM_T.n15 IM_T.t38 2.1905
R856 IM_T.n16 IM_T.t12 2.1905
R857 IM_T.n17 IM_T.t49 2.1905
R858 IM_T.n18 IM_T.t33 2.1905
R859 IM_T.n19 IM_T.t16 2.1905
R860 IM_T.n20 IM_T.t42 2.1905
R861 IM_T.n22 IM_T.t55 2.1905
R862 IM_T.n23 IM_T.t31 2.1905
R863 IM_T.n24 IM_T.t60 2.1905
R864 IM_T.n25 IM_T.t40 2.1905
R865 IM_T.n26 IM_T.t8 2.1905
R866 IM_T.n27 IM_T.t9 2.1905
R867 IM_T.n28 IM_T.t37 2.1905
R868 IM_T.n29 IM_T.t48 2.1905
R869 IM_T.n30 IM_T.t19 2.1905
R870 IM_T.n31 IM_T.t59 2.1905
R871 IM_T.n32 IM_T.t41 2.1905
R872 IM_T.n33 IM_T.t23 2.1905
R873 IM_T.n34 IM_T.t52 2.1905
R874 IM_T.n36 IM_T.t20 2.1905
R875 IM_T.n37 IM_T.t62 2.1905
R876 IM_T.n38 IM_T.t25 2.1905
R877 IM_T.n39 IM_T.t10 2.1905
R878 IM_T.n40 IM_T.t32 2.1905
R879 IM_T.n41 IM_T.t35 2.1905
R880 IM_T.n42 IM_T.t5 2.1905
R881 IM_T.n43 IM_T.t39 2.1905
R882 IM_T.n44 IM_T.t53 2.1905
R883 IM_T.n45 IM_T.t43 2.1905
R884 IM_T.n46 IM_T.t57 2.1905
R885 IM_T.n47 IM_T.t45 2.1905
R886 IM_T.n48 IM_T.t61 2.1905
R887 IM_T.n50 IM_T.t14 2.1905
R888 IM_T.n51 IM_T.t1 2.1905
R889 IM_T.n52 IM_T.t26 2.1905
R890 IM_T.n53 IM_T.t6 2.1905
R891 IM_T.n54 IM_T.t29 2.1905
R892 IM_T.n55 IM_T.t2 2.1905
R893 IM_T.n56 IM_T.t17 2.1905
R894 IM_T IM_T.n58 0.790466
R895 IM_T.n14 IM_T 0.790466
R896 IM_T IM_T.n57 0.783502
R897 IM_T.n58 IM_T 0.642327
R898 IM_T IM_T.n14 0.642327
R899 IM_T.n57 IM_T 0.636351
R900 OUT.n61 OUT.t36 6.79341
R901 OUT.n38 OUT.t9 6.79341
R902 OUT.n15 OUT.t19 6.79341
R903 OUT.n86 OUT.t56 6.79341
R904 OUT.n68 OUT.n46 6.10941
R905 OUT.n45 OUT.n23 6.10941
R906 OUT.n22 OUT.n0 6.10941
R907 OUT.n93 OUT.n71 6.10941
R908 OUT.n61 OUT.n60 3.51246
R909 OUT.n63 OUT.n56 3.51246
R910 OUT.n65 OUT.n52 3.51246
R911 OUT.n67 OUT.n48 3.51246
R912 OUT.n38 OUT.n37 3.51246
R913 OUT.n40 OUT.n33 3.51246
R914 OUT.n42 OUT.n29 3.51246
R915 OUT.n44 OUT.n25 3.51246
R916 OUT.n15 OUT.n14 3.51246
R917 OUT.n17 OUT.n10 3.51246
R918 OUT.n19 OUT.n6 3.51246
R919 OUT.n21 OUT.n2 3.51246
R920 OUT.n86 OUT.n85 3.51246
R921 OUT.n88 OUT.n81 3.51246
R922 OUT.n90 OUT.n77 3.51246
R923 OUT.n92 OUT.n73 3.51246
R924 OUT.n66 OUT.n50 3.37941
R925 OUT.n64 OUT.n54 3.37941
R926 OUT.n62 OUT.n58 3.37941
R927 OUT.n43 OUT.n27 3.37941
R928 OUT.n41 OUT.n31 3.37941
R929 OUT.n39 OUT.n35 3.37941
R930 OUT.n20 OUT.n4 3.37941
R931 OUT.n18 OUT.n8 3.37941
R932 OUT.n16 OUT.n12 3.37941
R933 OUT.n91 OUT.n75 3.37941
R934 OUT.n89 OUT.n79 3.37941
R935 OUT.n87 OUT.n83 3.37941
R936 OUT.n50 OUT.t24 2.7305
R937 OUT.n50 OUT.n49 2.7305
R938 OUT.n54 OUT.t20 2.7305
R939 OUT.n54 OUT.n53 2.7305
R940 OUT.n58 OUT.t18 2.7305
R941 OUT.n58 OUT.n57 2.7305
R942 OUT.n60 OUT.t61 2.7305
R943 OUT.n60 OUT.n59 2.7305
R944 OUT.n56 OUT.t57 2.7305
R945 OUT.n56 OUT.n55 2.7305
R946 OUT.n52 OUT.t62 2.7305
R947 OUT.n52 OUT.n51 2.7305
R948 OUT.n48 OUT.t5 2.7305
R949 OUT.n48 OUT.n47 2.7305
R950 OUT.n27 OUT.t15 2.7305
R951 OUT.n27 OUT.n26 2.7305
R952 OUT.n31 OUT.t4 2.7305
R953 OUT.n31 OUT.n30 2.7305
R954 OUT.n35 OUT.t40 2.7305
R955 OUT.n35 OUT.n34 2.7305
R956 OUT.n37 OUT.t28 2.7305
R957 OUT.n37 OUT.n36 2.7305
R958 OUT.n33 OUT.t53 2.7305
R959 OUT.n33 OUT.n32 2.7305
R960 OUT.n29 OUT.t1 2.7305
R961 OUT.n29 OUT.n28 2.7305
R962 OUT.n25 OUT.t12 2.7305
R963 OUT.n25 OUT.n24 2.7305
R964 OUT.n4 OUT.t25 2.7305
R965 OUT.n4 OUT.n3 2.7305
R966 OUT.n8 OUT.t14 2.7305
R967 OUT.n8 OUT.n7 2.7305
R968 OUT.n12 OUT.t47 2.7305
R969 OUT.n12 OUT.n11 2.7305
R970 OUT.n14 OUT.t54 2.7305
R971 OUT.n14 OUT.n13 2.7305
R972 OUT.n10 OUT.t23 2.7305
R973 OUT.n10 OUT.n9 2.7305
R974 OUT.n6 OUT.t32 2.7305
R975 OUT.n6 OUT.n5 2.7305
R976 OUT.n2 OUT.t39 2.7305
R977 OUT.n2 OUT.n1 2.7305
R978 OUT.n75 OUT.t63 2.7305
R979 OUT.n75 OUT.n74 2.7305
R980 OUT.n79 OUT.t50 2.7305
R981 OUT.n79 OUT.n78 2.7305
R982 OUT.n83 OUT.t29 2.7305
R983 OUT.n83 OUT.n82 2.7305
R984 OUT.n85 OUT.t16 2.7305
R985 OUT.n85 OUT.n84 2.7305
R986 OUT.n81 OUT.t41 2.7305
R987 OUT.n81 OUT.n80 2.7305
R988 OUT.n77 OUT.t48 2.7305
R989 OUT.n77 OUT.n76 2.7305
R990 OUT.n73 OUT.t60 2.7305
R991 OUT.n73 OUT.n72 2.7305
R992 OUT.n69 OUT 0.9359
R993 OUT.n70 OUT.n69 0.9269
R994 OUT OUT.n70 0.8093
R995 OUT.n68 OUT.n67 0.6845
R996 OUT.n67 OUT.n66 0.6845
R997 OUT.n66 OUT.n65 0.6845
R998 OUT.n65 OUT.n64 0.6845
R999 OUT.n64 OUT.n63 0.6845
R1000 OUT.n63 OUT.n62 0.6845
R1001 OUT.n62 OUT.n61 0.6845
R1002 OUT.n45 OUT.n44 0.6845
R1003 OUT.n44 OUT.n43 0.6845
R1004 OUT.n43 OUT.n42 0.6845
R1005 OUT.n42 OUT.n41 0.6845
R1006 OUT.n41 OUT.n40 0.6845
R1007 OUT.n40 OUT.n39 0.6845
R1008 OUT.n39 OUT.n38 0.6845
R1009 OUT.n22 OUT.n21 0.6845
R1010 OUT.n21 OUT.n20 0.6845
R1011 OUT.n20 OUT.n19 0.6845
R1012 OUT.n19 OUT.n18 0.6845
R1013 OUT.n18 OUT.n17 0.6845
R1014 OUT.n17 OUT.n16 0.6845
R1015 OUT.n16 OUT.n15 0.6845
R1016 OUT.n93 OUT.n92 0.6845
R1017 OUT.n92 OUT.n91 0.6845
R1018 OUT.n91 OUT.n90 0.6845
R1019 OUT.n90 OUT.n89 0.6845
R1020 OUT.n89 OUT.n88 0.6845
R1021 OUT.n88 OUT.n87 0.6845
R1022 OUT.n87 OUT.n86 0.6845
R1023 OUT OUT.n68 0.27275
R1024 OUT OUT.n45 0.27275
R1025 OUT OUT.n22 0.27275
R1026 OUT OUT.n93 0.27275
R1027 OUT.n69 OUT 0.0095
R1028 OUT.n70 OUT 0.0095
C0 OUT IM_T 3.01f
C1 IM_T IM 5.3f
C2 OUT IM 4.14f
C3 OUT VSS 11.7f
C4 IM VSS 28.7f
C5 IM_T VSS 49.5f
C6 OUT.n0 VSS 0.0355f
C7 OUT.t39 VSS 0.0149f
C8 OUT.n1 VSS 0.0149f
C9 OUT.n2 VSS 0.0332f
C10 OUT.t25 VSS 0.0149f
C11 OUT.n3 VSS 0.0149f
C12 OUT.n4 VSS 0.0315f
C13 OUT.t32 VSS 0.0149f
C14 OUT.n5 VSS 0.0149f
C15 OUT.n6 VSS 0.0332f
C16 OUT.t14 VSS 0.0149f
C17 OUT.n7 VSS 0.0149f
C18 OUT.n8 VSS 0.0315f
C19 OUT.t23 VSS 0.0149f
C20 OUT.n9 VSS 0.0149f
C21 OUT.n10 VSS 0.0332f
C22 OUT.t47 VSS 0.0149f
C23 OUT.n11 VSS 0.0149f
C24 OUT.n12 VSS 0.0315f
C25 OUT.t54 VSS 0.0149f
C26 OUT.n13 VSS 0.0149f
C27 OUT.n14 VSS 0.0332f
C28 OUT.t19 VSS 0.0534f
C29 OUT.n15 VSS 0.442f
C30 OUT.n16 VSS 0.269f
C31 OUT.n17 VSS 0.282f
C32 OUT.n18 VSS 0.269f
C33 OUT.n19 VSS 0.282f
C34 OUT.n20 VSS 0.269f
C35 OUT.n21 VSS 0.282f
C36 OUT.n22 VSS 0.215f
C37 OUT.n23 VSS 0.0355f
C38 OUT.t12 VSS 0.0149f
C39 OUT.n24 VSS 0.0149f
C40 OUT.n25 VSS 0.0332f
C41 OUT.t15 VSS 0.0149f
C42 OUT.n26 VSS 0.0149f
C43 OUT.n27 VSS 0.0315f
C44 OUT.t1 VSS 0.0149f
C45 OUT.n28 VSS 0.0149f
C46 OUT.n29 VSS 0.0332f
C47 OUT.t4 VSS 0.0149f
C48 OUT.n30 VSS 0.0149f
C49 OUT.n31 VSS 0.0315f
C50 OUT.t53 VSS 0.0149f
C51 OUT.n32 VSS 0.0149f
C52 OUT.n33 VSS 0.0332f
C53 OUT.t40 VSS 0.0149f
C54 OUT.n34 VSS 0.0149f
C55 OUT.n35 VSS 0.0315f
C56 OUT.t28 VSS 0.0149f
C57 OUT.n36 VSS 0.0149f
C58 OUT.n37 VSS 0.0332f
C59 OUT.t9 VSS 0.0534f
C60 OUT.n38 VSS 0.442f
C61 OUT.n39 VSS 0.269f
C62 OUT.n40 VSS 0.282f
C63 OUT.n41 VSS 0.269f
C64 OUT.n42 VSS 0.282f
C65 OUT.n43 VSS 0.269f
C66 OUT.n44 VSS 0.282f
C67 OUT.n45 VSS 0.215f
C68 OUT.n46 VSS 0.0355f
C69 OUT.t5 VSS 0.0149f
C70 OUT.n47 VSS 0.0149f
C71 OUT.n48 VSS 0.0332f
C72 OUT.t24 VSS 0.0149f
C73 OUT.n49 VSS 0.0149f
C74 OUT.n50 VSS 0.0315f
C75 OUT.t62 VSS 0.0149f
C76 OUT.n51 VSS 0.0149f
C77 OUT.n52 VSS 0.0332f
C78 OUT.t20 VSS 0.0149f
C79 OUT.n53 VSS 0.0149f
C80 OUT.n54 VSS 0.0315f
C81 OUT.t57 VSS 0.0149f
C82 OUT.n55 VSS 0.0149f
C83 OUT.n56 VSS 0.0332f
C84 OUT.t18 VSS 0.0149f
C85 OUT.n57 VSS 0.0149f
C86 OUT.n58 VSS 0.0315f
C87 OUT.t61 VSS 0.0149f
C88 OUT.n59 VSS 0.0149f
C89 OUT.n60 VSS 0.0332f
C90 OUT.t36 VSS 0.0534f
C91 OUT.n61 VSS 0.442f
C92 OUT.n62 VSS 0.269f
C93 OUT.n63 VSS 0.282f
C94 OUT.n64 VSS 0.269f
C95 OUT.n65 VSS 0.282f
C96 OUT.n66 VSS 0.269f
C97 OUT.n67 VSS 0.282f
C98 OUT.n68 VSS 0.215f
C99 OUT.n69 VSS 1.11f
C100 OUT.n70 VSS 1.04f
C101 OUT.n71 VSS 0.0355f
C102 OUT.t60 VSS 0.0149f
C103 OUT.n72 VSS 0.0149f
C104 OUT.n73 VSS 0.0332f
C105 OUT.t63 VSS 0.0149f
C106 OUT.n74 VSS 0.0149f
C107 OUT.n75 VSS 0.0315f
C108 OUT.t48 VSS 0.0149f
C109 OUT.n76 VSS 0.0149f
C110 OUT.n77 VSS 0.0332f
C111 OUT.t50 VSS 0.0149f
C112 OUT.n78 VSS 0.0149f
C113 OUT.n79 VSS 0.0315f
C114 OUT.t41 VSS 0.0149f
C115 OUT.n80 VSS 0.0149f
C116 OUT.n81 VSS 0.0332f
C117 OUT.t29 VSS 0.0149f
C118 OUT.n82 VSS 0.0149f
C119 OUT.n83 VSS 0.0315f
C120 OUT.t16 VSS 0.0149f
C121 OUT.n84 VSS 0.0149f
C122 OUT.n85 VSS 0.0332f
C123 OUT.t56 VSS 0.0534f
C124 OUT.n86 VSS 0.442f
C125 OUT.n87 VSS 0.269f
C126 OUT.n88 VSS 0.282f
C127 OUT.n89 VSS 0.269f
C128 OUT.n90 VSS 0.282f
C129 OUT.n91 VSS 0.269f
C130 OUT.n92 VSS 0.282f
C131 OUT.n93 VSS 0.215f
C132 IM_T.t4 VSS 0.0191f
C133 IM_T.t34 VSS 0.0191f
C134 IM_T.t56 VSS 0.0191f
C135 IM_T.t13 VSS 0.0191f
C136 IM_T.t28 VSS 0.0191f
C137 IM_T.t0 VSS 0.0191f
C138 IM_T.t21 VSS 0.195f
C139 IM_T.n0 VSS 0.224f
C140 IM_T.n1 VSS 0.206f
C141 IM_T.n2 VSS 0.206f
C142 IM_T.n3 VSS 0.206f
C143 IM_T.n4 VSS 0.206f
C144 IM_T.n5 VSS 0.2f
C145 IM_T.t7 VSS 0.0577f
C146 IM_T.n6 VSS 0.174f
C147 IM_T.t18 VSS 0.0191f
C148 IM_T.t47 VSS 0.0191f
C149 IM_T.t46 VSS 0.0191f
C150 IM_T.t22 VSS 0.0191f
C151 IM_T.t36 VSS 0.0191f
C152 IM_T.t15 VSS 0.0191f
C153 IM_T.t30 VSS 0.0191f
C154 IM_T.t3 VSS 0.106f
C155 IM_T.n7 VSS 0.142f
C156 IM_T.n8 VSS 0.128f
C157 IM_T.n9 VSS 0.128f
C158 IM_T.n10 VSS 0.128f
C159 IM_T.n11 VSS 0.128f
C160 IM_T.n12 VSS 0.128f
C161 IM_T.n13 VSS 0.109f
C162 IM_T.n14 VSS 0.195f
C163 IM_T.t42 VSS 0.0191f
C164 IM_T.t16 VSS 0.0191f
C165 IM_T.t33 VSS 0.0191f
C166 IM_T.t49 VSS 0.0191f
C167 IM_T.t12 VSS 0.0191f
C168 IM_T.t38 VSS 0.0191f
C169 IM_T.t63 VSS 0.195f
C170 IM_T.n15 VSS 0.224f
C171 IM_T.n16 VSS 0.206f
C172 IM_T.n17 VSS 0.206f
C173 IM_T.n18 VSS 0.206f
C174 IM_T.n19 VSS 0.206f
C175 IM_T.n20 VSS 0.2f
C176 IM_T.t44 VSS 0.0577f
C177 IM_T.n21 VSS 0.174f
C178 IM_T.t37 VSS 0.0191f
C179 IM_T.t9 VSS 0.0191f
C180 IM_T.t8 VSS 0.0191f
C181 IM_T.t40 VSS 0.0191f
C182 IM_T.t60 VSS 0.0191f
C183 IM_T.t31 VSS 0.0191f
C184 IM_T.t55 VSS 0.0191f
C185 IM_T.t24 VSS 0.106f
C186 IM_T.n22 VSS 0.142f
C187 IM_T.n23 VSS 0.128f
C188 IM_T.n24 VSS 0.128f
C189 IM_T.n25 VSS 0.128f
C190 IM_T.n26 VSS 0.128f
C191 IM_T.n27 VSS 0.128f
C192 IM_T.n28 VSS 0.109f
C193 IM_T.t52 VSS 0.0191f
C194 IM_T.t23 VSS 0.0191f
C195 IM_T.t41 VSS 0.0191f
C196 IM_T.t59 VSS 0.0191f
C197 IM_T.t19 VSS 0.0191f
C198 IM_T.t48 VSS 0.0191f
C199 IM_T.t11 VSS 0.195f
C200 IM_T.n29 VSS 0.224f
C201 IM_T.n30 VSS 0.206f
C202 IM_T.n31 VSS 0.206f
C203 IM_T.n32 VSS 0.206f
C204 IM_T.n33 VSS 0.206f
C205 IM_T.n34 VSS 0.2f
C206 IM_T.t54 VSS 0.0577f
C207 IM_T.n35 VSS 0.174f
C208 IM_T.t5 VSS 0.0191f
C209 IM_T.t35 VSS 0.0191f
C210 IM_T.t32 VSS 0.0191f
C211 IM_T.t10 VSS 0.0191f
C212 IM_T.t25 VSS 0.0191f
C213 IM_T.t62 VSS 0.0191f
C214 IM_T.t20 VSS 0.0191f
C215 IM_T.t51 VSS 0.106f
C216 IM_T.n36 VSS 0.142f
C217 IM_T.n37 VSS 0.128f
C218 IM_T.n38 VSS 0.128f
C219 IM_T.n39 VSS 0.128f
C220 IM_T.n40 VSS 0.128f
C221 IM_T.n41 VSS 0.128f
C222 IM_T.n42 VSS 0.109f
C223 IM_T.t61 VSS 0.0191f
C224 IM_T.t45 VSS 0.0191f
C225 IM_T.t57 VSS 0.0191f
C226 IM_T.t43 VSS 0.0191f
C227 IM_T.t53 VSS 0.0191f
C228 IM_T.t39 VSS 0.0191f
C229 IM_T.t50 VSS 0.195f
C230 IM_T.n43 VSS 0.224f
C231 IM_T.n44 VSS 0.206f
C232 IM_T.n45 VSS 0.206f
C233 IM_T.n46 VSS 0.206f
C234 IM_T.n47 VSS 0.206f
C235 IM_T.n48 VSS 0.2f
C236 IM_T.t27 VSS 0.0577f
C237 IM_T.n49 VSS 0.174f
C238 IM_T.t17 VSS 0.0191f
C239 IM_T.t2 VSS 0.0191f
C240 IM_T.t29 VSS 0.0191f
C241 IM_T.t6 VSS 0.0191f
C242 IM_T.t26 VSS 0.0191f
C243 IM_T.t1 VSS 0.0191f
C244 IM_T.t14 VSS 0.0191f
C245 IM_T.t58 VSS 0.106f
C246 IM_T.n50 VSS 0.142f
C247 IM_T.n51 VSS 0.128f
C248 IM_T.n52 VSS 0.128f
C249 IM_T.n53 VSS 0.128f
C250 IM_T.n54 VSS 0.128f
C251 IM_T.n55 VSS 0.128f
C252 IM_T.n56 VSS 0.111f
C253 IM_T.n57 VSS 0.197f
C254 IM_T.n58 VSS 0.195f
C255 a_424_490.t2 VSS 0.0109f
C256 a_424_490.t64 VSS 0.0109f
C257 a_424_490.n0 VSS 0.0109f
C258 a_424_490.n1 VSS 0.034f
C259 a_424_490.t45 VSS 0.0109f
C260 a_424_490.n2 VSS 0.0109f
C261 a_424_490.n3 VSS 0.0321f
C262 a_424_490.t75 VSS 0.0109f
C263 a_424_490.n4 VSS 0.0109f
C264 a_424_490.n5 VSS 0.0346f
C265 a_424_490.t47 VSS 0.0109f
C266 a_424_490.n6 VSS 0.0109f
C267 a_424_490.n7 VSS 0.0347f
C268 a_424_490.t93 VSS 0.0109f
C269 a_424_490.n8 VSS 0.0109f
C270 a_424_490.n9 VSS 0.034f
C271 a_424_490.n10 VSS 0.191f
C272 a_424_490.t43 VSS 0.0109f
C273 a_424_490.n11 VSS 0.0109f
C274 a_424_490.n12 VSS 0.0346f
C275 a_424_490.t69 VSS 0.0109f
C276 a_424_490.n13 VSS 0.0109f
C277 a_424_490.n14 VSS 0.0346f
C278 a_424_490.t9 VSS 0.0109f
C279 a_424_490.n15 VSS 0.0109f
C280 a_424_490.n16 VSS 0.0346f
C281 a_424_490.t61 VSS 0.0109f
C282 a_424_490.n17 VSS 0.0109f
C283 a_424_490.n18 VSS 0.0346f
C284 a_424_490.t19 VSS 0.0109f
C285 a_424_490.n19 VSS 0.0109f
C286 a_424_490.n20 VSS 0.0358f
C287 a_424_490.t89 VSS 0.0109f
C288 a_424_490.n21 VSS 0.0109f
C289 a_424_490.n22 VSS 0.0345f
C290 a_424_490.n23 VSS 0.0117f
C291 a_424_490.t42 VSS 0.0101f
C292 a_424_490.n24 VSS 0.0354f
C293 a_424_490.n25 VSS 0.183f
C294 a_424_490.n26 VSS 0.207f
C295 a_424_490.n27 VSS 0.208f
C296 a_424_490.n28 VSS 0.209f
C297 a_424_490.n29 VSS 0.209f
C298 a_424_490.n30 VSS 0.209f
C299 a_424_490.n31 VSS 0.208f
C300 a_424_490.t37 VSS 0.0109f
C301 a_424_490.n32 VSS 0.0109f
C302 a_424_490.n33 VSS 0.0303f
C303 a_424_490.n34 VSS 0.155f
C304 a_424_490.t96 VSS 0.0109f
C305 a_424_490.n35 VSS 0.0109f
C306 a_424_490.n36 VSS 0.0303f
C307 a_424_490.n37 VSS 0.164f
C308 a_424_490.t34 VSS 0.0109f
C309 a_424_490.n38 VSS 0.0109f
C310 a_424_490.n39 VSS 0.0347f
C311 a_424_490.t71 VSS 0.0109f
C312 a_424_490.n40 VSS 0.0109f
C313 a_424_490.n41 VSS 0.034f
C314 a_424_490.n42 VSS 0.191f
C315 a_424_490.t83 VSS 0.0109f
C316 a_424_490.n43 VSS 0.0109f
C317 a_424_490.n44 VSS 0.0303f
C318 a_424_490.n45 VSS 0.155f
C319 a_424_490.t13 VSS 0.0109f
C320 a_424_490.n46 VSS 0.0109f
C321 a_424_490.n47 VSS 0.0303f
C322 a_424_490.n48 VSS 0.163f
C323 a_424_490.t116 VSS 0.0109f
C324 a_424_490.n49 VSS 0.0109f
C325 a_424_490.n50 VSS 0.0303f
C326 a_424_490.n51 VSS 0.154f
C327 a_424_490.t90 VSS 0.0109f
C328 a_424_490.n52 VSS 0.0109f
C329 a_424_490.n53 VSS 0.0303f
C330 a_424_490.n54 VSS 0.163f
C331 a_424_490.t56 VSS 0.0109f
C332 a_424_490.n55 VSS 0.0109f
C333 a_424_490.n56 VSS 0.0303f
C334 a_424_490.n57 VSS 0.154f
C335 a_424_490.t29 VSS 0.0109f
C336 a_424_490.n58 VSS 0.0109f
C337 a_424_490.n59 VSS 0.0303f
C338 a_424_490.n60 VSS 0.164f
C339 a_424_490.t22 VSS 0.0109f
C340 a_424_490.n61 VSS 0.0109f
C341 a_424_490.n62 VSS 0.0303f
C342 a_424_490.n63 VSS 0.155f
C343 a_424_490.t80 VSS 0.0109f
C344 a_424_490.n64 VSS 0.0109f
C345 a_424_490.n65 VSS 0.0303f
C346 a_424_490.n66 VSS 0.164f
C347 a_424_490.n67 VSS 0.164f
C348 a_424_490.n68 VSS 0.165f
C349 a_424_490.n69 VSS 0.166f
C350 a_424_490.n70 VSS 0.166f
C351 a_424_490.n71 VSS 0.165f
C352 a_424_490.t12 VSS 0.0109f
C353 a_424_490.n72 VSS 0.0109f
C354 a_424_490.n73 VSS 0.0303f
C355 a_424_490.n74 VSS 0.155f
C356 a_424_490.t86 VSS 0.0109f
C357 a_424_490.n75 VSS 0.0109f
C358 a_424_490.n76 VSS 0.0303f
C359 a_424_490.n77 VSS 0.164f
C360 a_424_490.t27 VSS 0.0109f
C361 a_424_490.n78 VSS 0.0109f
C362 a_424_490.n79 VSS 0.0347f
C363 a_424_490.t105 VSS 0.0109f
C364 a_424_490.n80 VSS 0.0109f
C365 a_424_490.n81 VSS 0.034f
C366 a_424_490.n82 VSS 0.191f
C367 a_424_490.t63 VSS 0.0109f
C368 a_424_490.n83 VSS 0.0109f
C369 a_424_490.n84 VSS 0.0303f
C370 a_424_490.n85 VSS 0.155f
C371 a_424_490.t0 VSS 0.0109f
C372 a_424_490.n86 VSS 0.0109f
C373 a_424_490.n87 VSS 0.0303f
C374 a_424_490.n88 VSS 0.163f
C375 a_424_490.t8 VSS 0.0109f
C376 a_424_490.n89 VSS 0.0109f
C377 a_424_490.n90 VSS 0.0303f
C378 a_424_490.n91 VSS 0.154f
C379 a_424_490.t81 VSS 0.0109f
C380 a_424_490.n92 VSS 0.0109f
C381 a_424_490.n93 VSS 0.0303f
C382 a_424_490.n94 VSS 0.163f
C383 a_424_490.n95 VSS 0.166f
C384 a_424_490.n96 VSS 0.166f
C385 a_424_490.n97 VSS 0.165f
C386 a_424_490.t1 VSS 0.0109f
C387 a_424_490.n98 VSS 0.0109f
C388 a_424_490.n99 VSS 0.0303f
C389 a_424_490.n100 VSS 0.155f
C390 a_424_490.t98 VSS 0.0109f
C391 a_424_490.n101 VSS 0.0109f
C392 a_424_490.n102 VSS 0.0303f
C393 a_424_490.n103 VSS 0.164f
C394 a_424_490.t59 VSS 0.0109f
C395 a_424_490.n104 VSS 0.0109f
C396 a_424_490.n105 VSS 0.0322f
C397 a_424_490.t97 VSS 0.0109f
C398 a_424_490.n106 VSS 0.0109f
C399 a_424_490.n107 VSS 0.0303f
C400 a_424_490.n108 VSS 0.155f
C401 a_424_490.t113 VSS 0.0109f
C402 a_424_490.n109 VSS 0.0109f
C403 a_424_490.n110 VSS 0.0303f
C404 a_424_490.n111 VSS 0.163f
C405 a_424_490.t7 VSS 0.0109f
C406 a_424_490.n112 VSS 0.0109f
C407 a_424_490.n113 VSS 0.0322f
C408 a_424_490.t6 VSS 0.0109f
C409 a_424_490.n114 VSS 0.0109f
C410 a_424_490.n115 VSS 0.0303f
C411 a_424_490.n116 VSS 0.154f
C412 a_424_490.t78 VSS 0.0109f
C413 a_424_490.n117 VSS 0.0109f
C414 a_424_490.n118 VSS 0.0303f
C415 a_424_490.n119 VSS 0.163f
C416 a_424_490.t57 VSS 0.0109f
C417 a_424_490.n120 VSS 0.0109f
C418 a_424_490.n121 VSS 0.0321f
C419 a_424_490.t99 VSS 0.0109f
C420 a_424_490.n122 VSS 0.0109f
C421 a_424_490.n123 VSS 0.0303f
C422 a_424_490.n124 VSS 0.154f
C423 a_424_490.t35 VSS 0.0109f
C424 a_424_490.n125 VSS 0.0109f
C425 a_424_490.n126 VSS 0.0303f
C426 a_424_490.n127 VSS 0.164f
C427 a_424_490.t24 VSS 0.0109f
C428 a_424_490.n128 VSS 0.0109f
C429 a_424_490.n129 VSS 0.0303f
C430 a_424_490.n130 VSS 0.155f
C431 a_424_490.t73 VSS 0.0109f
C432 a_424_490.n131 VSS 0.0109f
C433 a_424_490.n132 VSS 0.0303f
C434 a_424_490.n133 VSS 0.164f
C435 a_424_490.t111 VSS 0.0109f
C436 a_424_490.n134 VSS 0.0109f
C437 a_424_490.n135 VSS 0.0303f
C438 a_424_490.n136 VSS 0.154f
C439 a_424_490.t36 VSS 0.0109f
C440 a_424_490.n137 VSS 0.0109f
C441 a_424_490.n138 VSS 0.0317f
C442 a_424_490.n139 VSS 0.163f
C443 a_424_490.t49 VSS 0.0109f
C444 a_424_490.n140 VSS 0.0109f
C445 a_424_490.n141 VSS 0.0345f
C446 a_424_490.n142 VSS 0.0117f
C447 a_424_490.t117 VSS 0.0101f
C448 a_424_490.n143 VSS 0.0354f
C449 a_424_490.n144 VSS 0.183f
C450 a_424_490.n145 VSS 0.165f
C451 a_424_490.t88 VSS 0.0109f
C452 a_424_490.n146 VSS 0.0109f
C453 a_424_490.n147 VSS 0.0303f
C454 a_424_490.n148 VSS 0.154f
C455 a_424_490.t31 VSS 0.0109f
C456 a_424_490.n149 VSS 0.0109f
C457 a_424_490.n150 VSS 0.0317f
C458 a_424_490.n151 VSS 0.163f
C459 a_424_490.t102 VSS 0.0109f
C460 a_424_490.n152 VSS 0.0109f
C461 a_424_490.n153 VSS 0.0345f
C462 a_424_490.n154 VSS 0.0117f
C463 a_424_490.t20 VSS 0.0101f
C464 a_424_490.n155 VSS 0.0354f
C465 a_424_490.n156 VSS 0.183f
C466 a_424_490.n157 VSS 0.165f
C467 a_424_490.n158 VSS 0.164f
C468 a_424_490.n159 VSS 0.165f
C469 a_424_490.t70 VSS 0.0109f
C470 a_424_490.n160 VSS 0.0109f
C471 a_424_490.n161 VSS 0.0303f
C472 a_424_490.n162 VSS 0.154f
C473 a_424_490.t124 VSS 0.0109f
C474 a_424_490.n163 VSS 0.0109f
C475 a_424_490.n164 VSS 0.0303f
C476 a_424_490.n165 VSS 0.164f
C477 a_424_490.t44 VSS 0.0109f
C478 a_424_490.n166 VSS 0.0109f
C479 a_424_490.n167 VSS 0.032f
C480 a_424_490.t28 VSS 0.0109f
C481 a_424_490.n168 VSS 0.0109f
C482 a_424_490.n169 VSS 0.0303f
C483 a_424_490.n170 VSS 0.155f
C484 a_424_490.t76 VSS 0.0109f
C485 a_424_490.n171 VSS 0.0109f
C486 a_424_490.n172 VSS 0.0303f
C487 a_424_490.n173 VSS 0.164f
C488 a_424_490.t62 VSS 0.0109f
C489 a_424_490.n174 VSS 0.0109f
C490 a_424_490.n175 VSS 0.0303f
C491 a_424_490.n176 VSS 0.154f
C492 a_424_490.t125 VSS 0.0109f
C493 a_424_490.n177 VSS 0.0109f
C494 a_424_490.n178 VSS 0.0317f
C495 a_424_490.n179 VSS 0.163f
C496 a_424_490.t51 VSS 0.0109f
C497 a_424_490.n180 VSS 0.0109f
C498 a_424_490.n181 VSS 0.032f
C499 a_424_490.t92 VSS 0.0109f
C500 a_424_490.n182 VSS 0.0109f
C501 a_424_490.n183 VSS 0.0345f
C502 a_424_490.n184 VSS 0.0117f
C503 a_424_490.t41 VSS 0.0101f
C504 a_424_490.n185 VSS 0.0354f
C505 a_424_490.n186 VSS 0.183f
C506 a_424_490.n187 VSS 0.201f
C507 a_424_490.n188 VSS 0.201f
C508 a_424_490.n189 VSS 0.202f
C509 a_424_490.n190 VSS 0.203f
C510 a_424_490.n191 VSS 0.202f
C511 a_424_490.n192 VSS 0.201f
C512 a_424_490.n193 VSS 0.191f
C513 a_424_490.n194 VSS 0.0347f
C514 a_424_490.n195 VSS 0.0109f
C515 IM.t2 VSS 0.0309f
C516 IM.t23 VSS 0.0309f
C517 IM.t54 VSS 0.0309f
C518 IM.t1 VSS 0.0309f
C519 IM.t35 VSS 0.0309f
C520 IM.t51 VSS 0.0309f
C521 IM.t27 VSS 0.0309f
C522 IM.t56 VSS 0.0309f
C523 IM.t9 VSS 0.0309f
C524 IM.t43 VSS 0.0309f
C525 IM.t17 VSS 0.0309f
C526 IM.t29 VSS 0.0309f
C527 IM.t62 VSS 0.0309f
C528 IM.t37 VSS 0.0309f
C529 IM.t8 VSS 0.0309f
C530 IM.t19 VSS 0.147f
C531 IM.n0 VSS 0.145f
C532 IM.n1 VSS 0.131f
C533 IM.n2 VSS 0.136f
C534 IM.n3 VSS 0.136f
C535 IM.n4 VSS 0.131f
C536 IM.n5 VSS 0.131f
C537 IM.n6 VSS 0.136f
C538 IM.n7 VSS 0.136f
C539 IM.n8 VSS 0.131f
C540 IM.n9 VSS 0.131f
C541 IM.n10 VSS 0.136f
C542 IM.n11 VSS 0.136f
C543 IM.n12 VSS 0.131f
C544 IM.n13 VSS 0.131f
C545 IM.n14 VSS 0.139f
C546 IM.n15 VSS 0.0511f
C547 IM.t25 VSS 0.0309f
C548 IM.t63 VSS 0.0309f
C549 IM.t33 VSS 0.0309f
C550 IM.t24 VSS 0.0309f
C551 IM.t57 VSS 0.0309f
C552 IM.t32 VSS 0.0309f
C553 IM.t4 VSS 0.0309f
C554 IM.t13 VSS 0.0309f
C555 IM.t30 VSS 0.0309f
C556 IM.t22 VSS 0.0309f
C557 IM.t60 VSS 0.0309f
C558 IM.t49 VSS 0.0309f
C559 IM.t18 VSS 0.0309f
C560 IM.t16 VSS 0.0309f
C561 IM.t47 VSS 0.0309f
C562 IM.t41 VSS 0.147f
C563 IM.n16 VSS 0.145f
C564 IM.n17 VSS 0.131f
C565 IM.n18 VSS 0.136f
C566 IM.n19 VSS 0.136f
C567 IM.n20 VSS 0.131f
C568 IM.n21 VSS 0.131f
C569 IM.n22 VSS 0.136f
C570 IM.n23 VSS 0.136f
C571 IM.n24 VSS 0.131f
C572 IM.n25 VSS 0.131f
C573 IM.n26 VSS 0.136f
C574 IM.n27 VSS 0.136f
C575 IM.n28 VSS 0.131f
C576 IM.n29 VSS 0.131f
C577 IM.n30 VSS 0.139f
C578 IM.t52 VSS 0.0309f
C579 IM.t10 VSS 0.0309f
C580 IM.t40 VSS 0.0309f
C581 IM.t50 VSS 0.0309f
C582 IM.t21 VSS 0.0309f
C583 IM.t39 VSS 0.0309f
C584 IM.t12 VSS 0.0309f
C585 IM.t42 VSS 0.0309f
C586 IM.t58 VSS 0.0309f
C587 IM.t31 VSS 0.0309f
C588 IM.t3 VSS 0.0309f
C589 IM.t15 VSS 0.0309f
C590 IM.t46 VSS 0.0309f
C591 IM.t26 VSS 0.0309f
C592 IM.t59 VSS 0.0309f
C593 IM.t7 VSS 0.147f
C594 IM.n31 VSS 0.145f
C595 IM.n32 VSS 0.131f
C596 IM.n33 VSS 0.136f
C597 IM.n34 VSS 0.136f
C598 IM.n35 VSS 0.131f
C599 IM.n36 VSS 0.131f
C600 IM.n37 VSS 0.136f
C601 IM.n38 VSS 0.136f
C602 IM.n39 VSS 0.131f
C603 IM.n40 VSS 0.131f
C604 IM.n41 VSS 0.136f
C605 IM.n42 VSS 0.136f
C606 IM.n43 VSS 0.131f
C607 IM.n44 VSS 0.131f
C608 IM.n45 VSS 0.139f
C609 IM.t28 VSS 0.0309f
C610 IM.t20 VSS 0.0309f
C611 IM.t6 VSS 0.0309f
C612 IM.t61 VSS 0.0309f
C613 IM.t45 VSS 0.0309f
C614 IM.t36 VSS 0.0309f
C615 IM.t11 VSS 0.0309f
C616 IM.t55 VSS 0.0309f
C617 IM.t44 VSS 0.0309f
C618 IM.t34 VSS 0.0309f
C619 IM.t5 VSS 0.0309f
C620 IM.t53 VSS 0.0309f
C621 IM.t38 VSS 0.0309f
C622 IM.t14 VSS 0.0309f
C623 IM.t0 VSS 0.0309f
C624 IM.t48 VSS 0.147f
C625 IM.n46 VSS 0.145f
C626 IM.n47 VSS 0.131f
C627 IM.n48 VSS 0.136f
C628 IM.n49 VSS 0.136f
C629 IM.n50 VSS 0.131f
C630 IM.n51 VSS 0.131f
C631 IM.n52 VSS 0.136f
C632 IM.n53 VSS 0.136f
C633 IM.n54 VSS 0.131f
C634 IM.n55 VSS 0.131f
C635 IM.n56 VSS 0.136f
C636 IM.n57 VSS 0.136f
C637 IM.n58 VSS 0.131f
C638 IM.n59 VSS 0.131f
C639 IM.n60 VSS 0.139f
C640 IM.n61 VSS 0.258f
C641 IM.n62 VSS 0.258f
.ends

