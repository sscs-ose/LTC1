magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -1968 -1968 12576 14320
<< psubdiff >>
rect 32 12298 368 12320
rect 32 12252 54 12298
rect 100 12252 168 12298
rect 214 12252 368 12298
rect 32 12184 368 12252
rect 32 12138 54 12184
rect 100 12138 168 12184
rect 214 12138 368 12184
rect 32 12116 368 12138
rect 32 12070 236 12116
rect 32 12024 54 12070
rect 100 12024 168 12070
rect 214 12024 236 12070
rect 32 11500 236 12024
rect 32 11454 54 11500
rect 100 11454 168 11500
rect 214 11454 236 11500
rect 32 11386 236 11454
rect 32 11340 54 11386
rect 100 11340 168 11386
rect 214 11340 236 11386
rect 32 11272 236 11340
rect 32 11226 54 11272
rect 100 11226 168 11272
rect 214 11226 236 11272
rect 32 11158 236 11226
rect 32 11112 54 11158
rect 100 11112 168 11158
rect 214 11112 236 11158
rect 32 11044 236 11112
rect 32 10998 54 11044
rect 100 10998 168 11044
rect 214 10998 236 11044
rect 32 10930 236 10998
rect 32 10884 54 10930
rect 100 10884 168 10930
rect 214 10884 236 10930
rect 32 10816 236 10884
rect 32 10770 54 10816
rect 100 10770 168 10816
rect 214 10770 236 10816
rect 32 10702 236 10770
rect 32 10656 54 10702
rect 100 10656 168 10702
rect 214 10656 236 10702
rect 32 10588 236 10656
rect 32 10542 54 10588
rect 100 10542 168 10588
rect 214 10542 236 10588
rect 32 10474 236 10542
rect 32 10428 54 10474
rect 100 10428 168 10474
rect 214 10428 236 10474
rect 32 10360 236 10428
rect 32 10314 54 10360
rect 100 10314 168 10360
rect 214 10314 236 10360
rect 32 10246 236 10314
rect 32 10200 54 10246
rect 100 10200 168 10246
rect 214 10200 236 10246
rect 32 10132 236 10200
rect 32 10086 54 10132
rect 100 10086 168 10132
rect 214 10086 236 10132
rect 32 10018 236 10086
rect 32 9972 54 10018
rect 100 9972 168 10018
rect 214 9972 236 10018
rect 32 9904 236 9972
rect 32 9858 54 9904
rect 100 9858 168 9904
rect 214 9858 236 9904
rect 32 9790 236 9858
rect 32 9744 54 9790
rect 100 9744 168 9790
rect 214 9744 236 9790
rect 32 9676 236 9744
rect 32 9630 54 9676
rect 100 9630 168 9676
rect 214 9630 236 9676
rect 32 9562 236 9630
rect 32 9516 54 9562
rect 100 9516 168 9562
rect 214 9516 236 9562
rect 32 9448 236 9516
rect 32 9402 54 9448
rect 100 9402 168 9448
rect 214 9402 236 9448
rect 32 9334 236 9402
rect 32 9288 54 9334
rect 100 9288 168 9334
rect 214 9288 236 9334
rect 32 9220 236 9288
rect 32 9174 54 9220
rect 100 9174 168 9220
rect 214 9174 236 9220
rect 32 9106 236 9174
rect 32 9060 54 9106
rect 100 9060 168 9106
rect 214 9060 236 9106
rect 32 8992 236 9060
rect 32 8946 54 8992
rect 100 8946 168 8992
rect 214 8946 236 8992
rect 32 8878 236 8946
rect 32 8832 54 8878
rect 100 8832 168 8878
rect 214 8832 236 8878
rect 32 8764 236 8832
rect 32 8718 54 8764
rect 100 8718 168 8764
rect 214 8718 236 8764
rect 32 8650 236 8718
rect 32 8604 54 8650
rect 100 8604 168 8650
rect 214 8604 236 8650
rect 32 8536 236 8604
rect 32 8490 54 8536
rect 100 8490 168 8536
rect 214 8490 236 8536
rect 32 8422 236 8490
rect 32 8376 54 8422
rect 100 8376 168 8422
rect 214 8376 236 8422
rect 32 8308 236 8376
rect 32 8262 54 8308
rect 100 8262 168 8308
rect 214 8262 236 8308
rect 32 8194 236 8262
rect 32 8148 54 8194
rect 100 8148 168 8194
rect 214 8148 236 8194
rect 32 8080 236 8148
rect 32 8034 54 8080
rect 100 8034 168 8080
rect 214 8034 236 8080
rect 32 7966 236 8034
rect 32 7920 54 7966
rect 100 7920 168 7966
rect 214 7920 236 7966
rect 32 7852 236 7920
rect 32 7806 54 7852
rect 100 7806 168 7852
rect 214 7806 236 7852
rect 32 7738 236 7806
rect 32 7692 54 7738
rect 100 7692 168 7738
rect 214 7692 236 7738
rect 32 7624 236 7692
rect 32 7578 54 7624
rect 100 7578 168 7624
rect 214 7578 236 7624
rect 32 7510 236 7578
rect 32 7464 54 7510
rect 100 7464 168 7510
rect 214 7464 236 7510
rect 32 7396 236 7464
rect 32 7350 54 7396
rect 100 7350 168 7396
rect 214 7350 236 7396
rect 32 7282 236 7350
rect 32 7236 54 7282
rect 100 7236 168 7282
rect 214 7236 236 7282
rect 32 7168 236 7236
rect 32 7122 54 7168
rect 100 7122 168 7168
rect 214 7122 236 7168
rect 32 7054 236 7122
rect 32 7008 54 7054
rect 100 7008 168 7054
rect 214 7008 236 7054
rect 32 6940 236 7008
rect 32 6894 54 6940
rect 100 6894 168 6940
rect 214 6894 236 6940
rect 32 6826 236 6894
rect 32 6780 54 6826
rect 100 6780 168 6826
rect 214 6780 236 6826
rect 32 6712 236 6780
rect 32 6666 54 6712
rect 100 6666 168 6712
rect 214 6666 236 6712
rect 32 6598 236 6666
rect 32 6552 54 6598
rect 100 6552 168 6598
rect 214 6552 236 6598
rect 32 6484 236 6552
rect 32 6438 54 6484
rect 100 6438 168 6484
rect 214 6438 236 6484
rect 32 6370 236 6438
rect 32 6324 54 6370
rect 100 6324 168 6370
rect 214 6324 236 6370
rect 32 6229 236 6324
rect 32 6025 300 6229
rect 4998 32 5400 236
<< psubdiffcont >>
rect 54 12252 100 12298
rect 168 12252 214 12298
rect 54 12138 100 12184
rect 168 12138 214 12184
rect 54 12024 100 12070
rect 168 12024 214 12070
rect 54 11454 100 11500
rect 168 11454 214 11500
rect 54 11340 100 11386
rect 168 11340 214 11386
rect 54 11226 100 11272
rect 168 11226 214 11272
rect 54 11112 100 11158
rect 168 11112 214 11158
rect 54 10998 100 11044
rect 168 10998 214 11044
rect 54 10884 100 10930
rect 168 10884 214 10930
rect 54 10770 100 10816
rect 168 10770 214 10816
rect 54 10656 100 10702
rect 168 10656 214 10702
rect 54 10542 100 10588
rect 168 10542 214 10588
rect 54 10428 100 10474
rect 168 10428 214 10474
rect 54 10314 100 10360
rect 168 10314 214 10360
rect 54 10200 100 10246
rect 168 10200 214 10246
rect 54 10086 100 10132
rect 168 10086 214 10132
rect 54 9972 100 10018
rect 168 9972 214 10018
rect 54 9858 100 9904
rect 168 9858 214 9904
rect 54 9744 100 9790
rect 168 9744 214 9790
rect 54 9630 100 9676
rect 168 9630 214 9676
rect 54 9516 100 9562
rect 168 9516 214 9562
rect 54 9402 100 9448
rect 168 9402 214 9448
rect 54 9288 100 9334
rect 168 9288 214 9334
rect 54 9174 100 9220
rect 168 9174 214 9220
rect 54 9060 100 9106
rect 168 9060 214 9106
rect 54 8946 100 8992
rect 168 8946 214 8992
rect 54 8832 100 8878
rect 168 8832 214 8878
rect 54 8718 100 8764
rect 168 8718 214 8764
rect 54 8604 100 8650
rect 168 8604 214 8650
rect 54 8490 100 8536
rect 168 8490 214 8536
rect 54 8376 100 8422
rect 168 8376 214 8422
rect 54 8262 100 8308
rect 168 8262 214 8308
rect 54 8148 100 8194
rect 168 8148 214 8194
rect 54 8034 100 8080
rect 168 8034 214 8080
rect 54 7920 100 7966
rect 168 7920 214 7966
rect 54 7806 100 7852
rect 168 7806 214 7852
rect 54 7692 100 7738
rect 168 7692 214 7738
rect 54 7578 100 7624
rect 168 7578 214 7624
rect 54 7464 100 7510
rect 168 7464 214 7510
rect 54 7350 100 7396
rect 168 7350 214 7396
rect 54 7236 100 7282
rect 168 7236 214 7282
rect 54 7122 100 7168
rect 168 7122 214 7168
rect 54 7008 100 7054
rect 168 7008 214 7054
rect 54 6894 100 6940
rect 168 6894 214 6940
rect 54 6780 100 6826
rect 168 6780 214 6826
rect 54 6666 100 6712
rect 168 6666 214 6712
rect 54 6552 100 6598
rect 168 6552 214 6598
rect 54 6438 100 6484
rect 168 6438 214 6484
rect 54 6324 100 6370
rect 168 6324 214 6370
<< metal1 >>
rect 43 12298 10565 12310
rect 43 12252 54 12298
rect 100 12252 168 12298
rect 214 12252 10565 12298
rect 43 12184 10565 12252
rect 43 12138 54 12184
rect 100 12138 168 12184
rect 214 12138 10565 12184
rect 43 12126 10565 12138
rect 43 12070 225 12126
rect 43 12024 54 12070
rect 100 12024 168 12070
rect 214 12024 225 12070
rect 43 11633 225 12024
rect 689 11723 9913 11855
rect 689 11655 2605 11723
rect 3125 11655 5041 11723
rect 5561 11655 7477 11723
rect 7997 11655 9913 11723
rect 43 11500 429 11633
rect 43 11454 54 11500
rect 100 11454 168 11500
rect 214 11454 429 11500
rect 43 11386 429 11454
rect 43 11340 54 11386
rect 100 11340 168 11386
rect 214 11340 429 11386
rect 43 11272 429 11340
rect 43 11226 54 11272
rect 100 11226 168 11272
rect 214 11226 429 11272
rect 43 11158 429 11226
rect 43 11112 54 11158
rect 100 11112 168 11158
rect 214 11112 429 11158
rect 43 11044 429 11112
rect 43 10998 54 11044
rect 100 10998 168 11044
rect 214 10998 429 11044
rect 43 10930 429 10998
rect 43 10884 54 10930
rect 100 10884 168 10930
rect 214 10884 429 10930
rect 43 10816 429 10884
rect 43 10770 54 10816
rect 100 10770 168 10816
rect 214 10770 429 10816
rect 43 10702 429 10770
rect 43 10656 54 10702
rect 100 10656 168 10702
rect 214 10656 429 10702
rect 43 10588 429 10656
rect 43 10542 54 10588
rect 100 10542 168 10588
rect 214 10542 429 10588
rect 43 10474 429 10542
rect 43 10428 54 10474
rect 100 10428 168 10474
rect 214 10428 429 10474
rect 43 10360 429 10428
rect 43 10314 54 10360
rect 100 10314 168 10360
rect 214 10314 429 10360
rect 43 10246 429 10314
rect 43 10200 54 10246
rect 100 10200 168 10246
rect 214 10200 429 10246
rect 43 10132 429 10200
rect 43 10086 54 10132
rect 100 10086 168 10132
rect 214 10086 429 10132
rect 43 10018 429 10086
rect 43 9972 54 10018
rect 100 9972 168 10018
rect 214 9972 429 10018
rect 43 9904 429 9972
rect 43 9858 54 9904
rect 100 9858 168 9904
rect 214 9858 429 9904
rect 43 9790 429 9858
rect 43 9744 54 9790
rect 100 9744 168 9790
rect 214 9744 429 9790
rect 43 9676 429 9744
rect 43 9630 54 9676
rect 100 9630 168 9676
rect 214 9630 429 9676
rect 43 9562 429 9630
rect 43 9516 54 9562
rect 100 9516 168 9562
rect 214 9516 429 9562
rect 43 9448 429 9516
rect 43 9402 54 9448
rect 100 9402 168 9448
rect 214 9402 429 9448
rect 43 9334 429 9402
rect 43 9288 54 9334
rect 100 9288 168 9334
rect 214 9288 429 9334
rect 43 9220 429 9288
rect 43 9174 54 9220
rect 100 9174 168 9220
rect 214 9174 429 9220
rect 43 9106 429 9174
rect 43 9060 54 9106
rect 100 9060 168 9106
rect 214 9060 429 9106
rect 43 8992 429 9060
rect 43 8946 54 8992
rect 100 8946 168 8992
rect 214 8946 429 8992
rect 43 8878 429 8946
rect 43 8832 54 8878
rect 100 8832 168 8878
rect 214 8832 429 8878
rect 43 8764 429 8832
rect 43 8718 54 8764
rect 100 8718 168 8764
rect 214 8718 429 8764
rect 43 8650 429 8718
rect 43 8604 54 8650
rect 100 8604 168 8650
rect 214 8604 429 8650
rect 43 8536 429 8604
rect 43 8490 54 8536
rect 100 8490 168 8536
rect 214 8490 429 8536
rect 43 8422 429 8490
rect 43 8376 54 8422
rect 100 8376 168 8422
rect 214 8376 429 8422
rect 43 8308 429 8376
rect 43 8262 54 8308
rect 100 8262 168 8308
rect 214 8262 429 8308
rect 43 8194 429 8262
rect 43 8148 54 8194
rect 100 8148 168 8194
rect 214 8148 429 8194
rect 43 8080 429 8148
rect 43 8034 54 8080
rect 100 8034 168 8080
rect 214 8034 429 8080
rect 43 7966 429 8034
rect 43 7920 54 7966
rect 100 7920 168 7966
rect 214 7920 429 7966
rect 43 7852 429 7920
rect 43 7806 54 7852
rect 100 7806 168 7852
rect 214 7806 429 7852
rect 43 7738 429 7806
rect 43 7692 54 7738
rect 100 7692 168 7738
rect 214 7692 429 7738
rect 43 7624 429 7692
rect 43 7578 54 7624
rect 100 7578 168 7624
rect 214 7578 429 7624
rect 43 7510 429 7578
rect 43 7464 54 7510
rect 100 7464 168 7510
rect 214 7464 429 7510
rect 43 7396 429 7464
rect 43 7350 54 7396
rect 100 7350 168 7396
rect 214 7350 429 7396
rect 43 7282 429 7350
rect 43 7236 54 7282
rect 100 7236 168 7282
rect 214 7236 429 7282
rect 43 7168 429 7236
rect 43 7122 54 7168
rect 100 7122 168 7168
rect 214 7122 429 7168
rect 43 7054 429 7122
rect 43 7008 54 7054
rect 100 7008 168 7054
rect 214 7008 429 7054
rect 43 6940 429 7008
rect 43 6894 54 6940
rect 100 6894 168 6940
rect 214 6894 429 6940
rect 43 6826 429 6894
rect 43 6780 54 6826
rect 100 6780 168 6826
rect 214 6780 429 6826
rect 43 6712 429 6780
rect 43 6666 54 6712
rect 100 6666 168 6712
rect 214 6666 429 6712
rect 43 6598 429 6666
rect 43 6552 54 6598
rect 100 6552 168 6598
rect 214 6552 429 6598
rect 43 6484 429 6552
rect 43 6438 54 6484
rect 100 6438 168 6484
rect 214 6483 429 6484
rect 10173 6483 10383 11633
rect 214 6438 10383 6483
rect 43 6370 10383 6438
rect 43 6324 54 6370
rect 100 6324 168 6370
rect 214 6324 10383 6370
rect 43 5771 10383 6324
rect 5058 226 5301 5771
rect 10173 621 10383 5771
rect 5561 531 7477 599
rect 7997 531 9913 599
rect 5561 399 9913 531
rect 5009 42 10565 226
use M1_PSUB_CDNS_69033583165350  M1_PSUB_CDNS_69033583165350_0
timestamp 1713338890
transform 0 -1 5304 1 0 6127
box -102 -5004 102 5004
use M1_PSUB_CDNS_69033583165350  M1_PSUB_CDNS_69033583165350_1
timestamp 1713338890
transform 0 -1 5304 1 0 12218
box -102 -5004 102 5004
use M1_PSUB_CDNS_69033583165351  M1_PSUB_CDNS_69033583165351_0
timestamp 1713338890
transform 1 0 10474 0 1 6176
box -102 -6144 102 6144
use M1_PSUB_CDNS_69033583165484  M1_PSUB_CDNS_69033583165484_0
timestamp 1713338890
transform 0 -1 7828 1 0 134
box -102 -2496 102 2496
use M1_PSUB_CDNS_69033583165485  M1_PSUB_CDNS_69033583165485_0
timestamp 1713338890
transform 1 0 5043 0 1 3014
box -45 -2959 45 2959
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_0
timestamp 1713338890
transform 1 0 5519 0 -1 5621
box -218 -350 2218 5092
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_1
timestamp 1713338890
transform 1 0 7955 0 -1 5621
box -218 -350 2218 5092
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_2
timestamp 1713338890
transform 1 0 647 0 1 6633
box -218 -350 2218 5092
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_3
timestamp 1713338890
transform 1 0 3083 0 1 6633
box -218 -350 2218 5092
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_4
timestamp 1713338890
transform 1 0 5519 0 1 6633
box -218 -350 2218 5092
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_5
timestamp 1713338890
transform 1 0 7955 0 1 6633
box -218 -350 2218 5092
<< labels >>
rlabel metal1 s 5302 6126 5302 6126 4 VMINUS
port 1 nsew
<< end >>
