magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1045 -2879 1045 2879
<< metal1 >>
rect -45 1873 45 1879
rect -45 1847 -39 1873
rect 39 1847 45 1873
rect -45 1811 45 1847
rect -45 1785 -39 1811
rect 39 1785 45 1811
rect -45 1749 45 1785
rect -45 1723 -39 1749
rect 39 1723 45 1749
rect -45 1687 45 1723
rect -45 1661 -39 1687
rect 39 1661 45 1687
rect -45 1625 45 1661
rect -45 1599 -39 1625
rect 39 1599 45 1625
rect -45 1563 45 1599
rect -45 1537 -39 1563
rect 39 1537 45 1563
rect -45 1501 45 1537
rect -45 1475 -39 1501
rect 39 1475 45 1501
rect -45 1439 45 1475
rect -45 1413 -39 1439
rect 39 1413 45 1439
rect -45 1377 45 1413
rect -45 1351 -39 1377
rect 39 1351 45 1377
rect -45 1315 45 1351
rect -45 1289 -39 1315
rect 39 1289 45 1315
rect -45 1253 45 1289
rect -45 1227 -39 1253
rect 39 1227 45 1253
rect -45 1191 45 1227
rect -45 1165 -39 1191
rect 39 1165 45 1191
rect -45 1129 45 1165
rect -45 1103 -39 1129
rect 39 1103 45 1129
rect -45 1067 45 1103
rect -45 1041 -39 1067
rect 39 1041 45 1067
rect -45 1005 45 1041
rect -45 979 -39 1005
rect 39 979 45 1005
rect -45 943 45 979
rect -45 917 -39 943
rect 39 917 45 943
rect -45 881 45 917
rect -45 855 -39 881
rect 39 855 45 881
rect -45 819 45 855
rect -45 793 -39 819
rect 39 793 45 819
rect -45 757 45 793
rect -45 731 -39 757
rect 39 731 45 757
rect -45 695 45 731
rect -45 669 -39 695
rect 39 669 45 695
rect -45 633 45 669
rect -45 607 -39 633
rect 39 607 45 633
rect -45 571 45 607
rect -45 545 -39 571
rect 39 545 45 571
rect -45 509 45 545
rect -45 483 -39 509
rect 39 483 45 509
rect -45 447 45 483
rect -45 421 -39 447
rect 39 421 45 447
rect -45 385 45 421
rect -45 359 -39 385
rect 39 359 45 385
rect -45 323 45 359
rect -45 297 -39 323
rect 39 297 45 323
rect -45 261 45 297
rect -45 235 -39 261
rect 39 235 45 261
rect -45 199 45 235
rect -45 173 -39 199
rect 39 173 45 199
rect -45 137 45 173
rect -45 111 -39 137
rect 39 111 45 137
rect -45 75 45 111
rect -45 49 -39 75
rect 39 49 45 75
rect -45 13 45 49
rect -45 -13 -39 13
rect 39 -13 45 13
rect -45 -49 45 -13
rect -45 -75 -39 -49
rect 39 -75 45 -49
rect -45 -111 45 -75
rect -45 -137 -39 -111
rect 39 -137 45 -111
rect -45 -173 45 -137
rect -45 -199 -39 -173
rect 39 -199 45 -173
rect -45 -235 45 -199
rect -45 -261 -39 -235
rect 39 -261 45 -235
rect -45 -297 45 -261
rect -45 -323 -39 -297
rect 39 -323 45 -297
rect -45 -359 45 -323
rect -45 -385 -39 -359
rect 39 -385 45 -359
rect -45 -421 45 -385
rect -45 -447 -39 -421
rect 39 -447 45 -421
rect -45 -483 45 -447
rect -45 -509 -39 -483
rect 39 -509 45 -483
rect -45 -545 45 -509
rect -45 -571 -39 -545
rect 39 -571 45 -545
rect -45 -607 45 -571
rect -45 -633 -39 -607
rect 39 -633 45 -607
rect -45 -669 45 -633
rect -45 -695 -39 -669
rect 39 -695 45 -669
rect -45 -731 45 -695
rect -45 -757 -39 -731
rect 39 -757 45 -731
rect -45 -793 45 -757
rect -45 -819 -39 -793
rect 39 -819 45 -793
rect -45 -855 45 -819
rect -45 -881 -39 -855
rect 39 -881 45 -855
rect -45 -917 45 -881
rect -45 -943 -39 -917
rect 39 -943 45 -917
rect -45 -979 45 -943
rect -45 -1005 -39 -979
rect 39 -1005 45 -979
rect -45 -1041 45 -1005
rect -45 -1067 -39 -1041
rect 39 -1067 45 -1041
rect -45 -1103 45 -1067
rect -45 -1129 -39 -1103
rect 39 -1129 45 -1103
rect -45 -1165 45 -1129
rect -45 -1191 -39 -1165
rect 39 -1191 45 -1165
rect -45 -1227 45 -1191
rect -45 -1253 -39 -1227
rect 39 -1253 45 -1227
rect -45 -1289 45 -1253
rect -45 -1315 -39 -1289
rect 39 -1315 45 -1289
rect -45 -1351 45 -1315
rect -45 -1377 -39 -1351
rect 39 -1377 45 -1351
rect -45 -1413 45 -1377
rect -45 -1439 -39 -1413
rect 39 -1439 45 -1413
rect -45 -1475 45 -1439
rect -45 -1501 -39 -1475
rect 39 -1501 45 -1475
rect -45 -1537 45 -1501
rect -45 -1563 -39 -1537
rect 39 -1563 45 -1537
rect -45 -1599 45 -1563
rect -45 -1625 -39 -1599
rect 39 -1625 45 -1599
rect -45 -1661 45 -1625
rect -45 -1687 -39 -1661
rect 39 -1687 45 -1661
rect -45 -1723 45 -1687
rect -45 -1749 -39 -1723
rect 39 -1749 45 -1723
rect -45 -1785 45 -1749
rect -45 -1811 -39 -1785
rect 39 -1811 45 -1785
rect -45 -1847 45 -1811
rect -45 -1873 -39 -1847
rect 39 -1873 45 -1847
rect -45 -1879 45 -1873
<< via1 >>
rect -39 1847 39 1873
rect -39 1785 39 1811
rect -39 1723 39 1749
rect -39 1661 39 1687
rect -39 1599 39 1625
rect -39 1537 39 1563
rect -39 1475 39 1501
rect -39 1413 39 1439
rect -39 1351 39 1377
rect -39 1289 39 1315
rect -39 1227 39 1253
rect -39 1165 39 1191
rect -39 1103 39 1129
rect -39 1041 39 1067
rect -39 979 39 1005
rect -39 917 39 943
rect -39 855 39 881
rect -39 793 39 819
rect -39 731 39 757
rect -39 669 39 695
rect -39 607 39 633
rect -39 545 39 571
rect -39 483 39 509
rect -39 421 39 447
rect -39 359 39 385
rect -39 297 39 323
rect -39 235 39 261
rect -39 173 39 199
rect -39 111 39 137
rect -39 49 39 75
rect -39 -13 39 13
rect -39 -75 39 -49
rect -39 -137 39 -111
rect -39 -199 39 -173
rect -39 -261 39 -235
rect -39 -323 39 -297
rect -39 -385 39 -359
rect -39 -447 39 -421
rect -39 -509 39 -483
rect -39 -571 39 -545
rect -39 -633 39 -607
rect -39 -695 39 -669
rect -39 -757 39 -731
rect -39 -819 39 -793
rect -39 -881 39 -855
rect -39 -943 39 -917
rect -39 -1005 39 -979
rect -39 -1067 39 -1041
rect -39 -1129 39 -1103
rect -39 -1191 39 -1165
rect -39 -1253 39 -1227
rect -39 -1315 39 -1289
rect -39 -1377 39 -1351
rect -39 -1439 39 -1413
rect -39 -1501 39 -1475
rect -39 -1563 39 -1537
rect -39 -1625 39 -1599
rect -39 -1687 39 -1661
rect -39 -1749 39 -1723
rect -39 -1811 39 -1785
rect -39 -1873 39 -1847
<< metal2 >>
rect -45 1873 45 1879
rect -45 1847 -39 1873
rect 39 1847 45 1873
rect -45 1811 45 1847
rect -45 1785 -39 1811
rect 39 1785 45 1811
rect -45 1749 45 1785
rect -45 1723 -39 1749
rect 39 1723 45 1749
rect -45 1687 45 1723
rect -45 1661 -39 1687
rect 39 1661 45 1687
rect -45 1625 45 1661
rect -45 1599 -39 1625
rect 39 1599 45 1625
rect -45 1563 45 1599
rect -45 1537 -39 1563
rect 39 1537 45 1563
rect -45 1501 45 1537
rect -45 1475 -39 1501
rect 39 1475 45 1501
rect -45 1439 45 1475
rect -45 1413 -39 1439
rect 39 1413 45 1439
rect -45 1377 45 1413
rect -45 1351 -39 1377
rect 39 1351 45 1377
rect -45 1315 45 1351
rect -45 1289 -39 1315
rect 39 1289 45 1315
rect -45 1253 45 1289
rect -45 1227 -39 1253
rect 39 1227 45 1253
rect -45 1191 45 1227
rect -45 1165 -39 1191
rect 39 1165 45 1191
rect -45 1129 45 1165
rect -45 1103 -39 1129
rect 39 1103 45 1129
rect -45 1067 45 1103
rect -45 1041 -39 1067
rect 39 1041 45 1067
rect -45 1005 45 1041
rect -45 979 -39 1005
rect 39 979 45 1005
rect -45 943 45 979
rect -45 917 -39 943
rect 39 917 45 943
rect -45 881 45 917
rect -45 855 -39 881
rect 39 855 45 881
rect -45 819 45 855
rect -45 793 -39 819
rect 39 793 45 819
rect -45 757 45 793
rect -45 731 -39 757
rect 39 731 45 757
rect -45 695 45 731
rect -45 669 -39 695
rect 39 669 45 695
rect -45 633 45 669
rect -45 607 -39 633
rect 39 607 45 633
rect -45 571 45 607
rect -45 545 -39 571
rect 39 545 45 571
rect -45 509 45 545
rect -45 483 -39 509
rect 39 483 45 509
rect -45 447 45 483
rect -45 421 -39 447
rect 39 421 45 447
rect -45 385 45 421
rect -45 359 -39 385
rect 39 359 45 385
rect -45 323 45 359
rect -45 297 -39 323
rect 39 297 45 323
rect -45 261 45 297
rect -45 235 -39 261
rect 39 235 45 261
rect -45 199 45 235
rect -45 173 -39 199
rect 39 173 45 199
rect -45 137 45 173
rect -45 111 -39 137
rect 39 111 45 137
rect -45 75 45 111
rect -45 49 -39 75
rect 39 49 45 75
rect -45 13 45 49
rect -45 -13 -39 13
rect 39 -13 45 13
rect -45 -49 45 -13
rect -45 -75 -39 -49
rect 39 -75 45 -49
rect -45 -111 45 -75
rect -45 -137 -39 -111
rect 39 -137 45 -111
rect -45 -173 45 -137
rect -45 -199 -39 -173
rect 39 -199 45 -173
rect -45 -235 45 -199
rect -45 -261 -39 -235
rect 39 -261 45 -235
rect -45 -297 45 -261
rect -45 -323 -39 -297
rect 39 -323 45 -297
rect -45 -359 45 -323
rect -45 -385 -39 -359
rect 39 -385 45 -359
rect -45 -421 45 -385
rect -45 -447 -39 -421
rect 39 -447 45 -421
rect -45 -483 45 -447
rect -45 -509 -39 -483
rect 39 -509 45 -483
rect -45 -545 45 -509
rect -45 -571 -39 -545
rect 39 -571 45 -545
rect -45 -607 45 -571
rect -45 -633 -39 -607
rect 39 -633 45 -607
rect -45 -669 45 -633
rect -45 -695 -39 -669
rect 39 -695 45 -669
rect -45 -731 45 -695
rect -45 -757 -39 -731
rect 39 -757 45 -731
rect -45 -793 45 -757
rect -45 -819 -39 -793
rect 39 -819 45 -793
rect -45 -855 45 -819
rect -45 -881 -39 -855
rect 39 -881 45 -855
rect -45 -917 45 -881
rect -45 -943 -39 -917
rect 39 -943 45 -917
rect -45 -979 45 -943
rect -45 -1005 -39 -979
rect 39 -1005 45 -979
rect -45 -1041 45 -1005
rect -45 -1067 -39 -1041
rect 39 -1067 45 -1041
rect -45 -1103 45 -1067
rect -45 -1129 -39 -1103
rect 39 -1129 45 -1103
rect -45 -1165 45 -1129
rect -45 -1191 -39 -1165
rect 39 -1191 45 -1165
rect -45 -1227 45 -1191
rect -45 -1253 -39 -1227
rect 39 -1253 45 -1227
rect -45 -1289 45 -1253
rect -45 -1315 -39 -1289
rect 39 -1315 45 -1289
rect -45 -1351 45 -1315
rect -45 -1377 -39 -1351
rect 39 -1377 45 -1351
rect -45 -1413 45 -1377
rect -45 -1439 -39 -1413
rect 39 -1439 45 -1413
rect -45 -1475 45 -1439
rect -45 -1501 -39 -1475
rect 39 -1501 45 -1475
rect -45 -1537 45 -1501
rect -45 -1563 -39 -1537
rect 39 -1563 45 -1537
rect -45 -1599 45 -1563
rect -45 -1625 -39 -1599
rect 39 -1625 45 -1599
rect -45 -1661 45 -1625
rect -45 -1687 -39 -1661
rect 39 -1687 45 -1661
rect -45 -1723 45 -1687
rect -45 -1749 -39 -1723
rect 39 -1749 45 -1723
rect -45 -1785 45 -1749
rect -45 -1811 -39 -1785
rect 39 -1811 45 -1785
rect -45 -1847 45 -1811
rect -45 -1873 -39 -1847
rect 39 -1873 45 -1847
rect -45 -1879 45 -1873
<< end >>
