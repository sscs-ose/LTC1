magic
tech gf180mcuC
magscale 1 10
timestamp 1694501647
<< nwell >>
rect -1104 -386 1104 386
<< nsubdiff >>
rect -1080 290 1080 362
rect -1080 -290 -1008 290
rect 1008 -290 1080 290
rect -1080 -362 1080 -290
<< polysilicon >>
rect -920 189 -680 202
rect -920 143 -907 189
rect -693 143 -680 189
rect -920 100 -680 143
rect -920 -143 -680 -100
rect -920 -189 -907 -143
rect -693 -189 -680 -143
rect -920 -202 -680 -189
rect -600 189 -360 202
rect -600 143 -587 189
rect -373 143 -360 189
rect -600 100 -360 143
rect -600 -143 -360 -100
rect -600 -189 -587 -143
rect -373 -189 -360 -143
rect -600 -202 -360 -189
rect -280 189 -40 202
rect -280 143 -267 189
rect -53 143 -40 189
rect -280 100 -40 143
rect -280 -143 -40 -100
rect -280 -189 -267 -143
rect -53 -189 -40 -143
rect -280 -202 -40 -189
rect 40 189 280 202
rect 40 143 53 189
rect 267 143 280 189
rect 40 100 280 143
rect 40 -143 280 -100
rect 40 -189 53 -143
rect 267 -189 280 -143
rect 40 -202 280 -189
rect 360 189 600 202
rect 360 143 373 189
rect 587 143 600 189
rect 360 100 600 143
rect 360 -143 600 -100
rect 360 -189 373 -143
rect 587 -189 600 -143
rect 360 -202 600 -189
rect 680 189 920 202
rect 680 143 693 189
rect 907 143 920 189
rect 680 100 920 143
rect 680 -143 920 -100
rect 680 -189 693 -143
rect 907 -189 920 -143
rect 680 -202 920 -189
<< polycontact >>
rect -907 143 -693 189
rect -907 -189 -693 -143
rect -587 143 -373 189
rect -587 -189 -373 -143
rect -267 143 -53 189
rect -267 -189 -53 -143
rect 53 143 267 189
rect 53 -189 267 -143
rect 373 143 587 189
rect 373 -189 587 -143
rect 693 143 907 189
rect 693 -189 907 -143
<< ppolyres >>
rect -920 -100 -680 100
rect -600 -100 -360 100
rect -280 -100 -40 100
rect 40 -100 280 100
rect 360 -100 600 100
rect 680 -100 920 100
<< metal1 >>
rect -918 143 -907 189
rect -693 143 -682 189
rect -598 143 -587 189
rect -373 143 -362 189
rect -278 143 -267 189
rect -53 143 -42 189
rect 42 143 53 189
rect 267 143 278 189
rect 362 143 373 189
rect 587 143 598 189
rect 682 143 693 189
rect 907 143 918 189
rect -918 -189 -907 -143
rect -693 -189 -682 -143
rect -598 -189 -587 -143
rect -373 -189 -362 -143
rect -278 -189 -267 -143
rect -53 -189 -42 -143
rect 42 -189 53 -143
rect 267 -189 278 -143
rect 362 -189 373 -143
rect 587 -189 598 -143
rect 682 -189 693 -143
rect 907 -189 918 -143
<< properties >>
string FIXED_BBOX -1044 -326 1044 326
string gencell ppolyf_u
string library gf180mcu
string parameters w 1.2 l 1.0 m 1 nx 6 wmin 0.80 lmin 1.00 rho 315 val 278.761 dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 0 grc 0 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 0
<< end >>
