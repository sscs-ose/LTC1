magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -3148 -2118 3148 2118
<< pwell >>
rect -1148 -118 1148 118
<< nmos >>
rect -1036 -50 -868 50
rect -764 -50 -596 50
rect -492 -50 -324 50
rect -220 -50 -52 50
rect 52 -50 220 50
rect 324 -50 492 50
rect 596 -50 764 50
rect 868 -50 1036 50
<< ndiff >>
rect -1124 23 -1036 50
rect -1124 -23 -1111 23
rect -1065 -23 -1036 23
rect -1124 -50 -1036 -23
rect -868 23 -764 50
rect -868 -23 -839 23
rect -793 -23 -764 23
rect -868 -50 -764 -23
rect -596 23 -492 50
rect -596 -23 -567 23
rect -521 -23 -492 23
rect -596 -50 -492 -23
rect -324 23 -220 50
rect -324 -23 -295 23
rect -249 -23 -220 23
rect -324 -50 -220 -23
rect -52 23 52 50
rect -52 -23 -23 23
rect 23 -23 52 23
rect -52 -50 52 -23
rect 220 23 324 50
rect 220 -23 249 23
rect 295 -23 324 23
rect 220 -50 324 -23
rect 492 23 596 50
rect 492 -23 521 23
rect 567 -23 596 23
rect 492 -50 596 -23
rect 764 23 868 50
rect 764 -23 793 23
rect 839 -23 868 23
rect 764 -50 868 -23
rect 1036 23 1124 50
rect 1036 -23 1065 23
rect 1111 -23 1124 23
rect 1036 -50 1124 -23
<< ndiffc >>
rect -1111 -23 -1065 23
rect -839 -23 -793 23
rect -567 -23 -521 23
rect -295 -23 -249 23
rect -23 -23 23 23
rect 249 -23 295 23
rect 521 -23 567 23
rect 793 -23 839 23
rect 1065 -23 1111 23
<< polysilicon >>
rect -1036 50 -868 94
rect -764 50 -596 94
rect -492 50 -324 94
rect -220 50 -52 94
rect 52 50 220 94
rect 324 50 492 94
rect 596 50 764 94
rect 868 50 1036 94
rect -1036 -94 -868 -50
rect -764 -94 -596 -50
rect -492 -94 -324 -50
rect -220 -94 -52 -50
rect 52 -94 220 -50
rect 324 -94 492 -50
rect 596 -94 764 -50
rect 868 -94 1036 -50
<< metal1 >>
rect -1111 23 -1065 48
rect -1111 -48 -1065 -23
rect -839 23 -793 48
rect -839 -48 -793 -23
rect -567 23 -521 48
rect -567 -48 -521 -23
rect -295 23 -249 48
rect -295 -48 -249 -23
rect -23 23 23 48
rect -23 -48 23 -23
rect 249 23 295 48
rect 249 -48 295 -23
rect 521 23 567 48
rect 521 -48 567 -23
rect 793 23 839 48
rect 793 -48 839 -23
rect 1065 23 1111 48
rect 1065 -48 1111 -23
<< end >>
