magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -4862 -2042 4862 2042
<< polysilicon >>
rect -2862 23 2862 42
rect -2862 -23 -2843 23
rect 2843 -23 2862 23
rect -2862 -42 2862 -23
<< polycontact >>
rect -2843 -23 2843 23
<< metal1 >>
rect -2854 23 2854 34
rect -2854 -23 -2843 23
rect 2843 -23 2854 23
rect -2854 -34 2854 -23
<< end >>
