magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1453 -1329 1453 1329
<< metal2 >>
rect -453 324 453 329
rect -453 296 -448 324
rect -420 296 -386 324
rect -358 296 -324 324
rect -296 296 -262 324
rect -234 296 -200 324
rect -172 296 -138 324
rect -110 296 -76 324
rect -48 296 -14 324
rect 14 296 48 324
rect 76 296 110 324
rect 138 296 172 324
rect 200 296 234 324
rect 262 296 296 324
rect 324 296 358 324
rect 386 296 420 324
rect 448 296 453 324
rect -453 262 453 296
rect -453 234 -448 262
rect -420 234 -386 262
rect -358 234 -324 262
rect -296 234 -262 262
rect -234 234 -200 262
rect -172 234 -138 262
rect -110 234 -76 262
rect -48 234 -14 262
rect 14 234 48 262
rect 76 234 110 262
rect 138 234 172 262
rect 200 234 234 262
rect 262 234 296 262
rect 324 234 358 262
rect 386 234 420 262
rect 448 234 453 262
rect -453 200 453 234
rect -453 172 -448 200
rect -420 172 -386 200
rect -358 172 -324 200
rect -296 172 -262 200
rect -234 172 -200 200
rect -172 172 -138 200
rect -110 172 -76 200
rect -48 172 -14 200
rect 14 172 48 200
rect 76 172 110 200
rect 138 172 172 200
rect 200 172 234 200
rect 262 172 296 200
rect 324 172 358 200
rect 386 172 420 200
rect 448 172 453 200
rect -453 138 453 172
rect -453 110 -448 138
rect -420 110 -386 138
rect -358 110 -324 138
rect -296 110 -262 138
rect -234 110 -200 138
rect -172 110 -138 138
rect -110 110 -76 138
rect -48 110 -14 138
rect 14 110 48 138
rect 76 110 110 138
rect 138 110 172 138
rect 200 110 234 138
rect 262 110 296 138
rect 324 110 358 138
rect 386 110 420 138
rect 448 110 453 138
rect -453 76 453 110
rect -453 48 -448 76
rect -420 48 -386 76
rect -358 48 -324 76
rect -296 48 -262 76
rect -234 48 -200 76
rect -172 48 -138 76
rect -110 48 -76 76
rect -48 48 -14 76
rect 14 48 48 76
rect 76 48 110 76
rect 138 48 172 76
rect 200 48 234 76
rect 262 48 296 76
rect 324 48 358 76
rect 386 48 420 76
rect 448 48 453 76
rect -453 14 453 48
rect -453 -14 -448 14
rect -420 -14 -386 14
rect -358 -14 -324 14
rect -296 -14 -262 14
rect -234 -14 -200 14
rect -172 -14 -138 14
rect -110 -14 -76 14
rect -48 -14 -14 14
rect 14 -14 48 14
rect 76 -14 110 14
rect 138 -14 172 14
rect 200 -14 234 14
rect 262 -14 296 14
rect 324 -14 358 14
rect 386 -14 420 14
rect 448 -14 453 14
rect -453 -48 453 -14
rect -453 -76 -448 -48
rect -420 -76 -386 -48
rect -358 -76 -324 -48
rect -296 -76 -262 -48
rect -234 -76 -200 -48
rect -172 -76 -138 -48
rect -110 -76 -76 -48
rect -48 -76 -14 -48
rect 14 -76 48 -48
rect 76 -76 110 -48
rect 138 -76 172 -48
rect 200 -76 234 -48
rect 262 -76 296 -48
rect 324 -76 358 -48
rect 386 -76 420 -48
rect 448 -76 453 -48
rect -453 -110 453 -76
rect -453 -138 -448 -110
rect -420 -138 -386 -110
rect -358 -138 -324 -110
rect -296 -138 -262 -110
rect -234 -138 -200 -110
rect -172 -138 -138 -110
rect -110 -138 -76 -110
rect -48 -138 -14 -110
rect 14 -138 48 -110
rect 76 -138 110 -110
rect 138 -138 172 -110
rect 200 -138 234 -110
rect 262 -138 296 -110
rect 324 -138 358 -110
rect 386 -138 420 -110
rect 448 -138 453 -110
rect -453 -172 453 -138
rect -453 -200 -448 -172
rect -420 -200 -386 -172
rect -358 -200 -324 -172
rect -296 -200 -262 -172
rect -234 -200 -200 -172
rect -172 -200 -138 -172
rect -110 -200 -76 -172
rect -48 -200 -14 -172
rect 14 -200 48 -172
rect 76 -200 110 -172
rect 138 -200 172 -172
rect 200 -200 234 -172
rect 262 -200 296 -172
rect 324 -200 358 -172
rect 386 -200 420 -172
rect 448 -200 453 -172
rect -453 -234 453 -200
rect -453 -262 -448 -234
rect -420 -262 -386 -234
rect -358 -262 -324 -234
rect -296 -262 -262 -234
rect -234 -262 -200 -234
rect -172 -262 -138 -234
rect -110 -262 -76 -234
rect -48 -262 -14 -234
rect 14 -262 48 -234
rect 76 -262 110 -234
rect 138 -262 172 -234
rect 200 -262 234 -234
rect 262 -262 296 -234
rect 324 -262 358 -234
rect 386 -262 420 -234
rect 448 -262 453 -234
rect -453 -296 453 -262
rect -453 -324 -448 -296
rect -420 -324 -386 -296
rect -358 -324 -324 -296
rect -296 -324 -262 -296
rect -234 -324 -200 -296
rect -172 -324 -138 -296
rect -110 -324 -76 -296
rect -48 -324 -14 -296
rect 14 -324 48 -296
rect 76 -324 110 -296
rect 138 -324 172 -296
rect 200 -324 234 -296
rect 262 -324 296 -296
rect 324 -324 358 -296
rect 386 -324 420 -296
rect 448 -324 453 -296
rect -453 -329 453 -324
<< via2 >>
rect -448 296 -420 324
rect -386 296 -358 324
rect -324 296 -296 324
rect -262 296 -234 324
rect -200 296 -172 324
rect -138 296 -110 324
rect -76 296 -48 324
rect -14 296 14 324
rect 48 296 76 324
rect 110 296 138 324
rect 172 296 200 324
rect 234 296 262 324
rect 296 296 324 324
rect 358 296 386 324
rect 420 296 448 324
rect -448 234 -420 262
rect -386 234 -358 262
rect -324 234 -296 262
rect -262 234 -234 262
rect -200 234 -172 262
rect -138 234 -110 262
rect -76 234 -48 262
rect -14 234 14 262
rect 48 234 76 262
rect 110 234 138 262
rect 172 234 200 262
rect 234 234 262 262
rect 296 234 324 262
rect 358 234 386 262
rect 420 234 448 262
rect -448 172 -420 200
rect -386 172 -358 200
rect -324 172 -296 200
rect -262 172 -234 200
rect -200 172 -172 200
rect -138 172 -110 200
rect -76 172 -48 200
rect -14 172 14 200
rect 48 172 76 200
rect 110 172 138 200
rect 172 172 200 200
rect 234 172 262 200
rect 296 172 324 200
rect 358 172 386 200
rect 420 172 448 200
rect -448 110 -420 138
rect -386 110 -358 138
rect -324 110 -296 138
rect -262 110 -234 138
rect -200 110 -172 138
rect -138 110 -110 138
rect -76 110 -48 138
rect -14 110 14 138
rect 48 110 76 138
rect 110 110 138 138
rect 172 110 200 138
rect 234 110 262 138
rect 296 110 324 138
rect 358 110 386 138
rect 420 110 448 138
rect -448 48 -420 76
rect -386 48 -358 76
rect -324 48 -296 76
rect -262 48 -234 76
rect -200 48 -172 76
rect -138 48 -110 76
rect -76 48 -48 76
rect -14 48 14 76
rect 48 48 76 76
rect 110 48 138 76
rect 172 48 200 76
rect 234 48 262 76
rect 296 48 324 76
rect 358 48 386 76
rect 420 48 448 76
rect -448 -14 -420 14
rect -386 -14 -358 14
rect -324 -14 -296 14
rect -262 -14 -234 14
rect -200 -14 -172 14
rect -138 -14 -110 14
rect -76 -14 -48 14
rect -14 -14 14 14
rect 48 -14 76 14
rect 110 -14 138 14
rect 172 -14 200 14
rect 234 -14 262 14
rect 296 -14 324 14
rect 358 -14 386 14
rect 420 -14 448 14
rect -448 -76 -420 -48
rect -386 -76 -358 -48
rect -324 -76 -296 -48
rect -262 -76 -234 -48
rect -200 -76 -172 -48
rect -138 -76 -110 -48
rect -76 -76 -48 -48
rect -14 -76 14 -48
rect 48 -76 76 -48
rect 110 -76 138 -48
rect 172 -76 200 -48
rect 234 -76 262 -48
rect 296 -76 324 -48
rect 358 -76 386 -48
rect 420 -76 448 -48
rect -448 -138 -420 -110
rect -386 -138 -358 -110
rect -324 -138 -296 -110
rect -262 -138 -234 -110
rect -200 -138 -172 -110
rect -138 -138 -110 -110
rect -76 -138 -48 -110
rect -14 -138 14 -110
rect 48 -138 76 -110
rect 110 -138 138 -110
rect 172 -138 200 -110
rect 234 -138 262 -110
rect 296 -138 324 -110
rect 358 -138 386 -110
rect 420 -138 448 -110
rect -448 -200 -420 -172
rect -386 -200 -358 -172
rect -324 -200 -296 -172
rect -262 -200 -234 -172
rect -200 -200 -172 -172
rect -138 -200 -110 -172
rect -76 -200 -48 -172
rect -14 -200 14 -172
rect 48 -200 76 -172
rect 110 -200 138 -172
rect 172 -200 200 -172
rect 234 -200 262 -172
rect 296 -200 324 -172
rect 358 -200 386 -172
rect 420 -200 448 -172
rect -448 -262 -420 -234
rect -386 -262 -358 -234
rect -324 -262 -296 -234
rect -262 -262 -234 -234
rect -200 -262 -172 -234
rect -138 -262 -110 -234
rect -76 -262 -48 -234
rect -14 -262 14 -234
rect 48 -262 76 -234
rect 110 -262 138 -234
rect 172 -262 200 -234
rect 234 -262 262 -234
rect 296 -262 324 -234
rect 358 -262 386 -234
rect 420 -262 448 -234
rect -448 -324 -420 -296
rect -386 -324 -358 -296
rect -324 -324 -296 -296
rect -262 -324 -234 -296
rect -200 -324 -172 -296
rect -138 -324 -110 -296
rect -76 -324 -48 -296
rect -14 -324 14 -296
rect 48 -324 76 -296
rect 110 -324 138 -296
rect 172 -324 200 -296
rect 234 -324 262 -296
rect 296 -324 324 -296
rect 358 -324 386 -296
rect 420 -324 448 -296
<< metal3 >>
rect -453 324 453 329
rect -453 296 -448 324
rect -420 296 -386 324
rect -358 296 -324 324
rect -296 296 -262 324
rect -234 296 -200 324
rect -172 296 -138 324
rect -110 296 -76 324
rect -48 296 -14 324
rect 14 296 48 324
rect 76 296 110 324
rect 138 296 172 324
rect 200 296 234 324
rect 262 296 296 324
rect 324 296 358 324
rect 386 296 420 324
rect 448 296 453 324
rect -453 262 453 296
rect -453 234 -448 262
rect -420 234 -386 262
rect -358 234 -324 262
rect -296 234 -262 262
rect -234 234 -200 262
rect -172 234 -138 262
rect -110 234 -76 262
rect -48 234 -14 262
rect 14 234 48 262
rect 76 234 110 262
rect 138 234 172 262
rect 200 234 234 262
rect 262 234 296 262
rect 324 234 358 262
rect 386 234 420 262
rect 448 234 453 262
rect -453 200 453 234
rect -453 172 -448 200
rect -420 172 -386 200
rect -358 172 -324 200
rect -296 172 -262 200
rect -234 172 -200 200
rect -172 172 -138 200
rect -110 172 -76 200
rect -48 172 -14 200
rect 14 172 48 200
rect 76 172 110 200
rect 138 172 172 200
rect 200 172 234 200
rect 262 172 296 200
rect 324 172 358 200
rect 386 172 420 200
rect 448 172 453 200
rect -453 138 453 172
rect -453 110 -448 138
rect -420 110 -386 138
rect -358 110 -324 138
rect -296 110 -262 138
rect -234 110 -200 138
rect -172 110 -138 138
rect -110 110 -76 138
rect -48 110 -14 138
rect 14 110 48 138
rect 76 110 110 138
rect 138 110 172 138
rect 200 110 234 138
rect 262 110 296 138
rect 324 110 358 138
rect 386 110 420 138
rect 448 110 453 138
rect -453 76 453 110
rect -453 48 -448 76
rect -420 48 -386 76
rect -358 48 -324 76
rect -296 48 -262 76
rect -234 48 -200 76
rect -172 48 -138 76
rect -110 48 -76 76
rect -48 48 -14 76
rect 14 48 48 76
rect 76 48 110 76
rect 138 48 172 76
rect 200 48 234 76
rect 262 48 296 76
rect 324 48 358 76
rect 386 48 420 76
rect 448 48 453 76
rect -453 14 453 48
rect -453 -14 -448 14
rect -420 -14 -386 14
rect -358 -14 -324 14
rect -296 -14 -262 14
rect -234 -14 -200 14
rect -172 -14 -138 14
rect -110 -14 -76 14
rect -48 -14 -14 14
rect 14 -14 48 14
rect 76 -14 110 14
rect 138 -14 172 14
rect 200 -14 234 14
rect 262 -14 296 14
rect 324 -14 358 14
rect 386 -14 420 14
rect 448 -14 453 14
rect -453 -48 453 -14
rect -453 -76 -448 -48
rect -420 -76 -386 -48
rect -358 -76 -324 -48
rect -296 -76 -262 -48
rect -234 -76 -200 -48
rect -172 -76 -138 -48
rect -110 -76 -76 -48
rect -48 -76 -14 -48
rect 14 -76 48 -48
rect 76 -76 110 -48
rect 138 -76 172 -48
rect 200 -76 234 -48
rect 262 -76 296 -48
rect 324 -76 358 -48
rect 386 -76 420 -48
rect 448 -76 453 -48
rect -453 -110 453 -76
rect -453 -138 -448 -110
rect -420 -138 -386 -110
rect -358 -138 -324 -110
rect -296 -138 -262 -110
rect -234 -138 -200 -110
rect -172 -138 -138 -110
rect -110 -138 -76 -110
rect -48 -138 -14 -110
rect 14 -138 48 -110
rect 76 -138 110 -110
rect 138 -138 172 -110
rect 200 -138 234 -110
rect 262 -138 296 -110
rect 324 -138 358 -110
rect 386 -138 420 -110
rect 448 -138 453 -110
rect -453 -172 453 -138
rect -453 -200 -448 -172
rect -420 -200 -386 -172
rect -358 -200 -324 -172
rect -296 -200 -262 -172
rect -234 -200 -200 -172
rect -172 -200 -138 -172
rect -110 -200 -76 -172
rect -48 -200 -14 -172
rect 14 -200 48 -172
rect 76 -200 110 -172
rect 138 -200 172 -172
rect 200 -200 234 -172
rect 262 -200 296 -172
rect 324 -200 358 -172
rect 386 -200 420 -172
rect 448 -200 453 -172
rect -453 -234 453 -200
rect -453 -262 -448 -234
rect -420 -262 -386 -234
rect -358 -262 -324 -234
rect -296 -262 -262 -234
rect -234 -262 -200 -234
rect -172 -262 -138 -234
rect -110 -262 -76 -234
rect -48 -262 -14 -234
rect 14 -262 48 -234
rect 76 -262 110 -234
rect 138 -262 172 -234
rect 200 -262 234 -234
rect 262 -262 296 -234
rect 324 -262 358 -234
rect 386 -262 420 -234
rect 448 -262 453 -234
rect -453 -296 453 -262
rect -453 -324 -448 -296
rect -420 -324 -386 -296
rect -358 -324 -324 -296
rect -296 -324 -262 -296
rect -234 -324 -200 -296
rect -172 -324 -138 -296
rect -110 -324 -76 -296
rect -48 -324 -14 -296
rect 14 -324 48 -296
rect 76 -324 110 -296
rect 138 -324 172 -296
rect 200 -324 234 -296
rect 262 -324 296 -296
rect 324 -324 358 -296
rect 386 -324 420 -296
rect 448 -324 453 -296
rect -453 -329 453 -324
<< end >>
