magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2083 -2000 4361 4575
<< nwell >>
rect -83 1281 2361 2575
<< polysilicon >>
rect 462 698 602 1442
rect 878 1142 1018 1442
rect 1294 1142 1434 1442
rect 1710 995 1850 1442
rect 878 698 1018 995
rect 1294 817 1850 995
rect 1294 698 1434 817
rect 1710 698 1850 817
<< metal1 >>
rect 79 2413 165 2481
rect 372 1486 448 2468
rect 616 2186 1524 2262
rect 616 1486 692 2186
rect 788 1090 864 2086
rect 1032 1486 1280 2086
rect 1448 1486 1524 2186
rect 498 928 864 1090
rect 1326 987 1402 1312
rect 1620 987 1696 2086
rect 1864 1486 1940 2468
rect 2113 2413 2199 2481
rect 79 11 165 79
rect 372 25 448 654
rect 616 254 692 654
rect 788 354 864 928
rect 914 825 1696 987
rect 1032 354 1280 654
rect 1448 254 1524 654
rect 1620 354 1696 825
rect 616 178 1524 254
rect 1864 25 1940 654
rect 2113 11 2199 79
<< metal2 >>
rect 616 474 692 1666
rect 752 1486 1108 1666
rect 752 654 828 1486
rect 914 1141 1822 1321
rect 752 474 1108 654
use M1_NWELL_CDNS_40661953145315  M1_NWELL_CDNS_40661953145315_0
timestamp 1713338890
transform 1 0 2233 0 1 1977
box -128 -598 128 598
use M1_NWELL_CDNS_40661953145315  M1_NWELL_CDNS_40661953145315_1
timestamp 1713338890
transform 1 0 45 0 1 1977
box -128 -598 128 598
use M1_NWELL_CDNS_40661953145323  M1_NWELL_CDNS_40661953145323_0
timestamp 1713338890
transform 1 0 1139 0 1 2447
box -1068 -128 1068 128
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_0
timestamp 1713338890
transform 1 0 532 0 1 1009
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_1
timestamp 1713338890
transform 1 0 1780 0 1 1231
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_2
timestamp 1713338890
transform 1 0 948 0 1 1231
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_3
timestamp 1713338890
transform 1 0 1364 0 1 1231
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_4
timestamp 1713338890
transform 1 0 948 0 1 906
box -42 -89 42 89
use M1_PSUB_CDNS_69033583165609  M1_PSUB_CDNS_69033583165609_0
timestamp 1713338890
transform 1 0 2233 0 -1 515
box -45 -515 45 515
use M1_PSUB_CDNS_69033583165609  M1_PSUB_CDNS_69033583165609_1
timestamp 1713338890
transform 1 0 45 0 -1 515
box -45 -515 45 515
use M1_PSUB_CDNS_69033583165622  M1_PSUB_CDNS_69033583165622_0
timestamp 1713338890
transform 1 0 1139 0 -1 45
box -985 -45 985 45
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_0
timestamp 1713338890
transform 1 0 1784 0 1 1231
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_1
timestamp 1713338890
transform 1 0 952 0 1 1231
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_2
timestamp 1713338890
transform 1 0 1070 0 1 1576
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_3
timestamp 1713338890
transform 1 0 1070 0 1 564
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_4
timestamp 1713338890
transform 1 0 654 0 1 564
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_5
timestamp 1713338890
transform 1 0 654 0 1 1576
box -38 -90 38 90
use nmos_6p0_CDNS_4066195314530  nmos_6p0_CDNS_4066195314530_0
timestamp 1713338890
transform 1 0 462 0 1 354
box -88 -44 228 344
use nmos_6p0_CDNS_4066195314530  nmos_6p0_CDNS_4066195314530_1
timestamp 1713338890
transform 1 0 1294 0 1 354
box -88 -44 228 344
use nmos_6p0_CDNS_4066195314530  nmos_6p0_CDNS_4066195314530_2
timestamp 1713338890
transform -1 0 1018 0 -1 654
box -88 -44 228 344
use nmos_6p0_CDNS_4066195314530  nmos_6p0_CDNS_4066195314530_3
timestamp 1713338890
transform -1 0 1850 0 -1 654
box -88 -44 228 344
use pmos_6p0_CDNS_4066195314512  pmos_6p0_CDNS_4066195314512_0
timestamp 1713338890
transform 1 0 462 0 1 1486
box -208 -120 348 720
use pmos_6p0_CDNS_4066195314512  pmos_6p0_CDNS_4066195314512_1
timestamp 1713338890
transform -1 0 1850 0 -1 2086
box -208 -120 348 720
use pmos_6p0_CDNS_4066195314512  pmos_6p0_CDNS_4066195314512_2
timestamp 1713338890
transform 1 0 1294 0 -1 2086
box -208 -120 348 720
use pmos_6p0_CDNS_4066195314512  pmos_6p0_CDNS_4066195314512_3
timestamp 1713338890
transform -1 0 1018 0 1 1486
box -208 -120 348 720
<< labels >>
rlabel metal2 s 1507 1222 1507 1222 4 B
port 1 nsew
rlabel metal1 s 1781 1234 1781 1234 4 B
port 1 nsew
rlabel metal1 s 533 1012 533 1012 4 A
port 2 nsew
rlabel metal1 s 244 45 244 45 4 VSS
port 3 nsew
rlabel metal1 s 270 2452 270 2452 4 VDD
port 4 nsew
rlabel metal2 s 783 1222 783 1222 4 Z
port 5 nsew
<< end >>
