* NGSPICE file created from CLK_div_99_mag_flat.ext - technology: gf180mcuC

.subckt pex_CLK_div_99_mag VSS VDD Vdiv99 RST CLK
X0 a_4437_8231# CLK_div_3_mag_0.Q0.t3 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VDD.t315 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X1 CLK_DIV_11_mag_new_0.Q2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t386 VDD.t385 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t498 VDD.t497 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X3 VSS CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 a_10363_9798# VSS.t313 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X4 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 a_12501_11889# VSS.t22 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X5 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_1.K.t2 VDD.t129 VDD.t128 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X6 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.Q0.t3 VDD.t142 VDD.t141 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X7 a_11337_10895# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VSS.t228 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X8 VDD CLK_div_3_mag_1.Q1.t3 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VDD.t285 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X9 a_9951_11931# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT VSS.t190 VSS.t189 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X10 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VDD.t39 VDD.t38 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X11 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD.t32 VDD.t31 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X12 a_4002_14308# CLK_DIV_11_mag_new_0.Q0 VSS.t148 VSS.t84 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X13 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t183 VDD.t182 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X14 a_3556_12901# CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 VDD.t195 VDD.t194 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X15 VDD CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VDD.t104 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X16 VDD CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.CLK.t0 VDD.t72 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X17 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 a_3994_15139# VDD.t384 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X18 a_2597_12515# CLK_DIV_11_mag_new_0.Q1 VSS.t89 VSS.t88 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X19 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t196 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X20 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t79 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X21 CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT VSS.t192 VSS.t191 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X22 VDD CLK_div_3_mag_1.JK_FF_mag_1.K.t2 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VDD.t378 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X23 CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT CLK_DIV_11_mag_new_0.nand3_mag_1.OUT VDD.t500 VDD.t499 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X24 a_10363_9798# CLK_div_3_mag_1.JK_FF_mag_1.K.t3 CLK_div_3_mag_1.Q0.t1 VSS.t263 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X25 CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 VSS.t285 VSS.t284 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X26 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_12347_13030# VSS.t187 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X27 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD.t264 VDD.t263 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X28 a_7226_13030# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t230 VSS.t229 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X29 VSS CLK_div_3_mag_1.Q1.t4 a_12215_9798# VSS.t195 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X30 VSS CLK.t0 a_11779_8699# VSS.t28 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X31 VSS CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_10209_10895# VSS.t155 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X32 CLK_DIV_11_mag_new_0.Q1 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t3 a_13475_13030# VSS.t253 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X33 VDD CLK_div_3_mag_0.Q0.t4 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t312 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X34 VDD CLK.t1 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VDD.t40 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X35 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t332 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X36 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD.t296 VDD.t295 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X37 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.Q2 a_8663_11887# VSS.t279 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X38 CLK_DIV_11_mag_new_0.Q1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD.t471 VDD.t470 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X39 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.Q1.t3 VDD.t137 VDD.t136 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X40 a_5128_10895# RST.t0 a_4968_10895# VSS.t257 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X41 a_6816_11933# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT VSS.t118 VSS.t117 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X42 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.K VDD.t494 VDD.t493 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X43 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_6098_13030# VSS.t116 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X44 VSS CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.CLK.t1 VSS.t51 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X45 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD.t53 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X46 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK.t2 VDD.t44 VDD.t43 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X47 a_11779_8699# CLK_div_3_mag_1.Q1.t5 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN VSS.t28 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X48 a_15500_11885# CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT VSS.t72 VSS.t71 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X49 CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT CLK_DIV_11_mag_new_0.Q3 a_13858_15251# VDD.t309 pfet_03v3 ad=1.06p pd=5.68u as=0.624p ps=2.92u w=2.4u l=0.28u
X50 VDD CLK.t3 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN VDD.t45 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X51 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.Q1 a_11777_11889# VSS.t87 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X52 CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.and2_mag_3.IN1 VDD.t251 VDD.t250 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X53 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN VSS.t1 VSS.t0 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X54 CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT CLK_DIV_11_mag_new_0.nand3_mag_1.OUT VSS.t338 VSS.t337 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X55 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t260 VDD.t259 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X56 a_7421_10895# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t243 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X57 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN VSS.t165 VSS.t164 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X58 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN VSS.t99 VSS.t98 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X59 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.Q1 VDD.t124 VDD.t123 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X60 CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 VSS.t242 VSS.t241 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X61 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.Q2 a_10515_11931# VSS.t278 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X62 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.Q1 VDD.t122 VDD.t110 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X63 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK.t4 VDD.t49 VDD.t48 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X64 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.Vdiv3.t2 VDD.t414 VDD.t413 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X65 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_1.Q1.t6 VDD.t289 VDD.t288 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X66 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.Q3 a_5528_11889# VSS.t212 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X67 a_10096_15189# CLK_DIV_11_mag_new_0.and2_mag_3.IN1 VSS.t168 VSS.t167 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X68 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t2 VDD.t244 VDD.t243 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X69 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_1.QB VDD.t8 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X70 VDD CLK_div_3_mag_1.or_2_mag_0.IN2 a_10806_8231# VDD.t184 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X71 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT RST.t1 VDD.t371 VDD.t370 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X72 a_9227_11887# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT VSS.t47 VSS.t46 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X73 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.Q3 VDD.t308 VDD.t307 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X74 a_7011_9798# CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.Q1.t2 VSS.t2 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X75 CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS.t326 VSS.t325 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X76 a_13629_11933# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 VSS.t200 VSS.t199 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X77 VSS CLK_div_3_mag_0.JK_FF_mag_1.K.t3 a_8863_9798# VSS.t11 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X78 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_12911_13030# VSS.t270 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X79 VSS VDD.t507 a_12221_10895# VSS.t111 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X80 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD.t475 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X81 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 VSS.t133 VSS.t132 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X82 VSS CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_7575_9798# VSS.t2 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X83 VSS CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t4 CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN VSS.t254 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X84 a_2597_14017# CLK_DIV_11_mag_new_0.Q1 VSS.t86 VSS.t85 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X85 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.K.t0 VDD.t16 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X86 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD.t189 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X87 a_5534_12986# CLK_div_3_mag_0.Vdiv3.t3 a_5374_12986# VSS.t301 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X88 VSS CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT VSS.t304 nfet_03v3 ad=86.8f pd=0.92u as=86.8f ps=0.92u w=0.22u l=0.28u
X89 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_16070_13026# VSS.t321 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X90 VSS CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_14514_10895# VSS.t48 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X91 VDD CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN VDD.t304 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X92 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.CLK.t2 VDD.t12 VDD.t11 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X93 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_DIV_11_mag_new_0.Q0 VDD.t176 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X94 a_7380_11933# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t125 VSS.t124 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X95 a_8863_9798# CLK_div_3_mag_0.CLK.t3 a_8703_9798# VSS.t11 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X96 VSS CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_7011_9798# VSS.t2 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X97 VDD CLK_div_3_mag_0.Vdiv3.t4 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT VDD.t442 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X98 a_7575_9798# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t2 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X99 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB VDD.t175 VDD.t174 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X100 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD.t222 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X101 a_8669_12984# CLK_div_3_mag_0.Vdiv3.t5 a_8509_12984# VSS.t302 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X102 a_12501_11889# RST.t2 a_12341_11889# VSS.t258 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X103 CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN VDD.t193 VDD.t192 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X104 a_14508_9798# CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t59 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X105 VSS CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN VSS.t316 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X106 VSS CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN VSS.t96 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X107 a_10361_13028# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t268 VSS.t267 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X108 CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN VSS.t184 VSS.t183 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X109 VDD RST.t3 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT VDD.t372 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X110 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t125 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X111 a_15232_9798# CLK.t5 a_15072_9798# VSS.t37 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X112 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN VSS.t249 VSS.t248 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X113 VDD CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t424 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X114 VDD CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.Vdiv3.t0 VDD.t341 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X115 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VDD.t37 VDD.t36 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X116 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.K VDD.t492 VDD.t491 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X117 CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT CLK_DIV_11_mag_new_0.Q3 VSS.t211 VSS.t210 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X118 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.Vdiv3.t6 VSS.t300 VSS.t299 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X119 a_12347_13030# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT VSS.t55 VSS.t54 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X120 a_3994_9798# CLK_div_3_mag_0.JK_FF_mag_1.K.t4 CLK_div_3_mag_0.Q0.t2 VSS.t2 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X121 VDD VDD.t163 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VDD.t164 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X122 a_10209_10895# CLK_div_3_mag_1.Q0.t4 CLK_div_3_mag_1.JK_FF_mag_1.K VSS.t95 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X123 a_15078_10895# CLK_div_3_mag_1.Q1.t7 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VSS.t198 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X124 a_10927_9798# CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t27 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X125 VDD CLK_div_3_mag_0.Q1.t4 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t138 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X126 a_15072_9798# CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VSS.t76 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X127 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t481 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X128 VSS CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_11491_9798# VSS.t134 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X129 VSS CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_13790_10895# VSS.t56 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X130 a_12055_9798# CLK_div_3_mag_1.JK_FF_mag_1.K.t4 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VSS.t264 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X131 a_6098_13030# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT VSS.t170 VSS.t169 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X132 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_1.Q0.t5 VSS.t97 VSS.t96 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X133 VSS CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.Vdiv3.t1 VSS.t235 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X134 VDD VDD.t159 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t160 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X135 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t488 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X136 CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.and2_mag_3.IN1 a_10961_15230# VSS.t166 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X137 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.Q0.t0 VDD.t62 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X138 a_5692_10895# CLK_div_3_mag_0.Q0.t5 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS.t215 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X139 VDD CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.Q3 VDD.t348 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X140 VSS CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_10927_9798# VSS.t225 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X141 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VDD.t450 VDD.t449 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X142 VSS CLK.t6 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VSS.t38 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X143 a_11491_9798# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t204 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X144 a_6857_10895# CLK_div_3_mag_0.Q1.t5 CLK_div_3_mag_0.JK_FF_mag_1.QB VSS.t94 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X145 a_10515_11931# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t234 VSS.t233 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X146 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 a_15660_11885# VSS.t178 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X147 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t2 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X148 a_7985_10895# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS.t31 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X149 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_16224_11929# VSS.t73 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X150 VDD CLK_div_3_mag_0.Vdiv3.t7 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t437 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X151 a_12215_9798# CLK.t7 a_12055_9798# VSS.t41 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X152 CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_3_mag_0.Vdiv3.t8 VDD.t441 VDD.t440 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X153 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_DIV_11_mag_new_0.Q2 VSS.t277 VSS.t276 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X154 VDD CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.or_2_mag_0.IN2 VDD.t375 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X155 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD.t5 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X156 a_5528_11889# CLK_div_3_mag_0.Vdiv3.t9 a_5368_11889# VSS.t171 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X157 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT VDD.t275 VDD.t274 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X158 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD.t101 VDD.t100 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X159 VSS CLK_div_3_mag_0.CLK.t4 a_5410_8699# VSS.t12 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X160 CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.Q1.t8 VDD.t325 VDD.t324 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X161 CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN VDD.t88 VDD.t87 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X162 VDD CLK_div_3_mag_0.Vdiv3.t10 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t254 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X163 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VDD.t92 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X164 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.Q2 VDD.t408 VDD.t407 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X165 a_14782_12982# CLK_DIV_11_mag_new_0.JK_FF_mag_3.K VSS.t333 VSS.t332 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X166 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.Q0 VDD.t221 VDD.t220 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X167 a_12221_10895# CLK.t8 a_12061_10895# VSS.t42 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X168 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT VDD.t188 VDD.t187 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X169 CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_3_mag_0.Vdiv3.t11 a_10256_15189# VSS.t172 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X170 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB VDD.t431 VDD.t430 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X171 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 a_9387_11887# VSS.t175 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X172 VSS CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_13226_10895# VSS.t8 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X173 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.Q0.t6 VDD.t311 VDD.t310 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X174 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT VDD.t206 VDD.t205 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X175 VDD CLK_div_3_mag_0.CLK.t5 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t13 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X176 a_14514_10895# RST.t4 a_14354_10895# VSS.t259 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X177 VDD CLK_div_3_mag_0.Q1.t6 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t359 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X178 CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD.t168 VDD.t167 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X179 VSS CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.or_2_mag_0.IN2 VSS.t260 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X180 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_15506_13026# VSS.t129 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X181 CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t5 a_5466_15136# VDD.t369 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X182 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.K VDD.t412 VDD.t411 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X183 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t504 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X184 CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_16634_13026# VSS.t120 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X185 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.Q2 a_2757_14017# VSS.t275 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X186 a_8509_12984# CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t3 VSS.t163 VSS.t162 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X187 VSS CLK.t9 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VSS.t43 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X188 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT RST.t5 VDD.t20 VDD.t19 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X189 a_12341_11889# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT VSS.t140 VSS.t139 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X190 CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q3 a_2590_14702# VSS.t209 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X191 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT VDD.t356 VDD.t355 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X192 a_10806_8231# CLK_div_3_mag_1.Q0.t6 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN VDD.t143 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X193 VSS CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_3840_10895# VSS.t16 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X194 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT VDD.t204 VDD.t203 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X195 CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN VSS.t62 VSS.t61 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X196 CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q1 VDD.t121 VDD.t120 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X197 a_8869_10895# CLK_div_3_mag_0.CLK.t6 a_8709_10895# VSS.t15 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X198 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.Q2 VDD.t427 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X199 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t319 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X200 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.K VDD.t268 VDD.t267 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X201 a_6092_11889# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT VSS.t272 VSS.t271 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X202 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK.t10 VDD.t66 VDD.t65 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X203 VSS CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_8145_10895# VSS.t149 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X204 VDD CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 VDD.t301 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X205 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 a_3556_12901# VDD.t469 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X206 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t501 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X207 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t394 VDD.t393 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X208 VSS CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_8139_9798# VSS.t2 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X209 a_12911_13030# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 VSS.t21 VSS.t20 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X210 a_8703_9798# CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS.t11 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X211 a_10773_10895# CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t26 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X212 a_11783_12986# CLK_div_3_mag_0.Vdiv3.t12 a_11623_12986# VSS.t308 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X213 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t478 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X214 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_14942_12982# VSS.t119 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X215 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t278 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X216 VSS VDD.t510 a_15238_10895# VSS.t108 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X217 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.CLK.t7 VDD.t234 VDD.t233 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X218 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT VSS.t244 VSS.t61 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X219 VDD CLK_div_3_mag_0.CLK.t8 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VDD.t235 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X220 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VDD.t448 VDD.t447 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X221 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD.t262 VDD.t261 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X222 CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN VDD.t284 VDD.t283 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X223 a_13065_11933# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT VSS.t186 VSS.t185 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X224 a_6662_13030# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t336 VSS.t335 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X225 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD.t368 VDD.t367 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X226 a_14776_11885# CLK_DIV_11_mag_new_0.JK_FF_mag_3.K VSS.t331 VSS.t330 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X227 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD.t271 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X228 VSS CLK_div_3_mag_0.Q1.t7 a_5846_9798# VSS.t11 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X229 CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t336 VDD.t335 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X230 a_16788_11929# CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 VSS.t74 VSS.t73 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X231 VDD CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t6 CLK_DIV_11_mag_new_0.Q1 VDD.t452 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X232 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.QB VDD.t95 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X233 VDD CLK_div_3_mag_0.Vdiv3.t13 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT VDD.t457 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X234 VSS CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_4558_9798# VSS.t2 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X235 CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VDD.t485 VDD.t484 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X236 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT VDD.t277 VDD.t276 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X237 a_16224_11929# CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT VSS.t128 VSS.t73 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X238 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t4 VDD.t298 VDD.t297 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X239 VSS VDD.t511 a_5852_10895# VSS.t105 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X240 VSS CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_4404_10895# VSS.t327 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X241 Vdiv99 CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT VDD.t150 VDD.t149 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X242 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT RST.t6 VDD.t22 VDD.t21 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X243 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN VDD.t148 VDD.t147 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X244 VSS CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_3994_9798# VSS.t2 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X245 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t171 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X246 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.CLK.t9 VDD.t239 VDD.t238 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X247 a_4558_9798# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t2 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X248 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_3_mag_0.Vdiv3.t14 VSS.t310 VSS.t309 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X249 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VDD.t202 VDD.t201 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X250 VSS CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_5122_9798# VSS.t2 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X251 VSS CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_11497_10895# VSS.t5 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X252 VDD RST.t7 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT VDD.t23 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X253 VDD CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t209 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X254 VDD CLK_div_3_mag_0.JK_FF_mag_1.K.t5 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t130 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X255 a_13475_13030# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 VSS.t320 VSS.t319 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X256 a_13226_10895# CLK_div_3_mag_1.Q1.t9 CLK_div_3_mag_1.JK_FF_mag_1.QB VSS.t224 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X257 a_14354_10895# CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VSS.t66 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X258 VDD CLK_div_3_mag_0.CLK.t10 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VDD.t240 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X259 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t419 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X260 a_15506_13026# CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT VSS.t142 VSS.t141 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X261 a_8663_11887# CLK_div_3_mag_0.Vdiv3.t15 a_8503_11887# VSS.t297 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X262 CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT VDD.t282 VDD.t281 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X263 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t487 VDD.t486 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X264 a_16634_13026# CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 VSS.t115 VSS.t114 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X265 VDD CLK_DIV_11_mag_new_0.Q1 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN VDD.t117 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X266 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD.t390 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X267 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_3_mag_0.Vdiv3.t16 VDD.t436 VDD.t435 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X268 a_13858_15251# CLK_DIV_11_mag_new_0.and2_mag_3.OUT a_13698_15251# VDD.t451 pfet_03v3 ad=0.624p pd=2.92u as=0.624p ps=2.92u w=2.4u l=0.28u
X269 a_5410_8699# CLK_div_3_mag_0.Q1.t8 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS.t12 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X270 VDD VDD.t155 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t156 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X271 a_3840_10895# CLK_div_3_mag_0.Q0.t7 CLK_div_3_mag_0.JK_FF_mag_1.K VSS.t214 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X272 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t364 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X273 a_11777_11889# CLK_div_3_mag_0.Vdiv3.t17 a_11617_11889# VSS.t298 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X274 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.Q3 a_7380_11933# VSS.t208 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X275 VDD CLK_DIV_11_mag_new_0.Q2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB VDD.t404 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X276 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_1.Q1.t2 VDD.t432 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X277 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.Q0 a_14936_11885# VSS.t147 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X278 a_8709_10895# CLK_div_3_mag_0.Q1.t9 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS.t247 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X279 VDD RST.t8 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT VDD.t26 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X280 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VDD.t200 VDD.t199 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X281 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t7 VDD.t456 VDD.t455 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X282 VDD CLK_div_3_mag_0.Vdiv3.t18 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT VDD.t460 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X283 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_8669_12984# VSS.t293 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X284 VDD CLK_div_3_mag_1.Q0.t7 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VDD.t144 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X285 CLK_DIV_11_mag_new_0.Q2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_10361_13028# VSS.t292 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X286 a_8145_10895# RST.t9 a_7985_10895# VSS.t19 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X287 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t179 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X288 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t258 VDD.t257 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X289 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.Q1.t10 VDD.t358 VDD.t357 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X290 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t292 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X291 VDD CLK_div_3_mag_0.Vdiv3.t19 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT VDD.t463 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X292 a_3994_15139# CLK_DIV_11_mag_new_0.Q0 VDD.t219 VDD.t218 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X293 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 VDD.t347 VDD.t346 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X294 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t316 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X295 VDD CLK_div_3_mag_1.JK_FF_mag_1.K.t5 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VDD.t381 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X296 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q1 a_4002_14308# VSS.t84 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X297 VDD CLK_div_3_mag_0.or_2_mag_0.IN2 a_4437_8231# VDD.t225 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X298 a_11623_12986# CLK_DIV_11_mag_new_0.JK_FF_mag_2.K VSS.t283 VSS.t282 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X299 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_9797_13028# VSS.t340 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X300 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 a_6252_11889# VSS.t334 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X301 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t89 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X302 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t338 VDD.t337 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X303 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t496 VDD.t495 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X304 a_15238_10895# CLK.t11 a_15078_10895# VSS.t60 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X305 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_9233_13028# VSS.t188 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X306 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_DIV_11_mag_new_0.Q2 VDD.t403 VDD.t402 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X307 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.Vdiv3.t20 VSS.t312 VSS.t311 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X308 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT VDD.t76 VDD.t75 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X309 a_5374_12986# CLK_DIV_11_mag_new_0.JK_FF_mag_0.K VSS.t182 VSS.t181 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X310 a_16070_13026# CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 VSS.t177 VSS.t176 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X311 CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q1 VDD.t116 VDD.t115 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X312 a_4968_10895# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS.t322 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X313 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_1.Q0.t2 VDD.t466 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X314 a_5852_10895# CLK_div_3_mag_0.CLK.t11 a_5692_10895# VSS.t161 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X315 a_4404_10895# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t303 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X316 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD.t329 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X317 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t253 VDD.t252 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X318 a_8139_9798# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t2 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X319 VSS CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS.t152 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X320 VDD CLK_DIV_11_mag_new_0.Q1 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t0 VDD.t112 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X321 VDD CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN VDD.t247 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X322 VSS CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_6857_10895# VSS.t67 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X323 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.Q2 VDD.t401 VDD.t400 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X324 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.JK_FF_mag_1.K.t6 VDD.t232 VDD.t231 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X325 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD.t387 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X326 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_1.K.t0 VDD.t228 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X327 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN VDD.t1 VDD.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X328 VDD CLK_div_3_mag_1.Q1.t10 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VDD.t326 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X329 VDD CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB VDD.t215 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X330 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q1 VDD.t111 VDD.t110 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X331 a_11497_10895# RST.t10 a_11337_10895# VSS.t273 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X332 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT VDD.t99 VDD.t98 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X333 a_5846_9798# CLK_div_3_mag_0.CLK.t12 a_5686_9798# VSS.t11 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X334 a_14942_12982# CLK_div_3_mag_0.Vdiv3.t21 a_14782_12982# VSS.t34 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X335 CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN VSS.t131 VSS.t130 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X336 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q3 a_2597_12515# VSS.t207 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X337 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN VDD.t363 VDD.t362 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X338 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT RST.t11 VDD.t396 VDD.t395 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X339 CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN VSS.t194 VSS.t193 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X340 a_8503_11887# CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t5 VSS.t206 VSS.t205 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X341 a_13790_10895# CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t138 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X342 CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_7226_13030# VSS.t240 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X343 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.Q0 VSS.t146 VSS.t145 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X344 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.Q0.t8 VSS.t213 VSS.t152 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X345 a_5686_9798# CLK_div_3_mag_0.JK_FF_mag_1.K.t6 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS.t11 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X346 a_13698_15251# CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 VDD.t416 VDD.t415 pfet_03v3 ad=0.624p pd=2.92u as=1.06p ps=5.68u w=2.4u l=0.28u
X347 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN VDD.t246 VDD.t245 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X348 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VDD.t354 VDD.t353 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X349 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t340 VDD.t339 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X350 a_11617_11889# CLK_DIV_11_mag_new_0.JK_FF_mag_2.K VSS.t281 VSS.t280 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X351 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t68 VDD.t67 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X352 VSS CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_5128_10895# VSS.t289 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X353 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_6816_11933# VSS.t217 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X354 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.K VDD.t410 VDD.t409 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X355 VDD CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_1.or_2_mag_0.IN2 VDD.t33 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X356 VSS CLK_div_3_mag_0.CLK.t13 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VSS.t218 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X357 VSS CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN VSS.t145 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X358 a_5122_9798# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t2 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X359 a_15660_11885# RST.t12 a_15500_11885# VSS.t178 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X360 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_9951_11931# VSS.t339 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X361 VDD CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.nand3_mag_1.OUT VDD.t212 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X362 VSS VDD.t513 a_8869_10895# VSS.t102 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X363 a_5368_11889# CLK_DIV_11_mag_new_0.JK_FF_mag_0.K VSS.t180 VSS.t179 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X364 VSS CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_7421_10895# VSS.t250 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X365 VSS CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_13380_9798# VSS.t294 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X366 VDD CLK_div_3_mag_0.Vdiv3.t22 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t56 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X367 a_13944_9798# CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t137 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X368 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t170 VDD.t169 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X369 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.K VDD.t266 VDD.t265 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X370 VDD CLK_div_3_mag_0.JK_FF_mag_1.K.t7 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t133 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X371 a_9797_13028# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t174 VSS.t173 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X372 VDD CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT VDD.t209 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X373 VDD VDD.t151 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VDD.t152 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X374 a_6252_11889# RST.t13 a_6092_11889# VSS.t274 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X375 Vdiv99 CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT VSS.t101 VSS.t100 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X376 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t50 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X377 CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t270 VDD.t269 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X378 a_12061_10895# CLK_div_3_mag_1.Q0.t8 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VSS.t70 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X379 VDD RST.t14 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t397 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X380 a_10256_15189# CLK_DIV_11_mag_new_0.Q0 a_10096_15189# VSS.t144 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X381 VDD CLK_div_3_mag_0.Vdiv3.t23 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t59 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X382 VSS CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_14508_9798# VSS.t121 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X383 a_9233_13028# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT VSS.t232 VSS.t231 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X384 VSS CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_1.or_2_mag_0.IN2 VSS.t23 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X385 a_13380_9798# CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.Q1.t1 VSS.t75 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X386 a_9387_11887# RST.t15 a_9227_11887# VSS.t238 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X387 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VDD.t69 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X388 VSS CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_10773_10895# VSS.t201 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X389 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t8 a_11783_12986# VSS.t307 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X390 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_3_mag_0.Vdiv3.t24 VSS.t287 VSS.t286 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X391 VSS CLK_div_3_mag_1.JK_FF_mag_1.K.t7 a_15232_9798# VSS.t158 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X392 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.CLK.t14 VDD.t323 VDD.t322 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X393 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.Q1 a_13629_11933# VSS.t83 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X394 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.Vdiv3.t25 VDD.t418 VDD.t417 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X395 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_0.Q1.t0 VDD.t107 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X396 VSS CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_13944_9798# VSS.t63 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X397 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VDD.t352 VDD.t351 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X398 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q0 VDD.t208 VDD.t207 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X399 VDD CLK.t12 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VDD.t82 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X400 a_5466_15136# CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 VDD.t345 VDD.t344 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X401 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD.t30 VDD.t29 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X402 a_10961_15230# CLK_DIV_11_mag_new_0.Q1 VSS.t82 VSS.t81 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X403 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD.t472 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X404 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VDD.t78 VDD.t77 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X405 a_2757_14017# CLK_DIV_11_mag_new_0.Q0 a_2597_14017# VSS.t143 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X406 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_13065_11933# VSS.t269 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X407 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_6662_13030# VSS.t216 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X408 a_14936_11885# CLK_div_3_mag_0.Vdiv3.t26 a_14776_11885# VSS.t288 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X409 a_2590_14702# CLK_DIV_11_mag_new_0.Q1 VSS.t80 VSS.t79 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X410 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_3_mag_0.Vdiv3.t27 VDD.t446 VDD.t445 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X411 VSS CLK_div_3_mag_0.CLK.t15 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VSS.t221 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X412 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_DIV_11_mag_new_0.Q0 a_16788_11929# VSS.t73 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X413 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_5534_12986# VSS.t239 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X414 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK.t13 VDD.t86 VDD.t85 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X415 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD.t291 VDD.t290 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
R0 CLK_div_3_mag_0.Q0.n2 CLK_div_3_mag_0.Q0.t5 36.935
R1 CLK_div_3_mag_0.Q0.n3 CLK_div_3_mag_0.Q0.t7 31.4332
R2 CLK_div_3_mag_0.Q0.n5 CLK_div_3_mag_0.Q0.t3 29.8135
R3 CLK_div_3_mag_0.Q0.n5 CLK_div_3_mag_0.Q0.t8 27.8352
R4 CLK_div_3_mag_0.Q0.n2 CLK_div_3_mag_0.Q0.t4 18.1962
R5 CLK_div_3_mag_0.Q0.n3 CLK_div_3_mag_0.Q0.t6 15.3826
R6 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.Q0.t2 7.09905
R7 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.Q0.n3 6.86029
R8 CLK_div_3_mag_0.Q0.n4 CLK_div_3_mag_0.Q0 5.01077
R9 CLK_div_3_mag_0.Q0.n6 CLK_div_3_mag_0.Q0 3.41843
R10 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.Q0.n1 3.25053
R11 CLK_div_3_mag_0.Q0.n1 CLK_div_3_mag_0.Q0.t0 2.2755
R12 CLK_div_3_mag_0.Q0.n1 CLK_div_3_mag_0.Q0.n0 2.2755
R13 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.Q0.n6 2.2505
R14 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.Q0.n2 2.13459
R15 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.Q0.n5 1.74998
R16 CLK_div_3_mag_0.Q0.n6 CLK_div_3_mag_0.Q0.n4 1.50381
R17 CLK_div_3_mag_0.Q0.n4 CLK_div_3_mag_0.Q0 1.12067
R18 VDD.n229 VDD.t415 2529.02
R19 VDD.n235 VDD 2301.38
R20 VDD.n208 VDD 2301.38
R21 VDD.n236 VDD.n235 1842.37
R22 VDD.n209 VDD.n208 1842.37
R23 VDD.n239 VDD.t212 1403.56
R24 VDD.n241 VDD.t484 1242.86
R25 VDD.n232 VDD.t87 1105.93
R26 VDD.t309 VDD.n226 1011.51
R27 VDD.t384 VDD.n212 857.144
R28 VDD.t369 VDD.n216 857.144
R29 VDD.n235 VDD.t192 812.681
R30 VDD.n208 VDD.t283 812.681
R31 VDD.t179 VDD.t104 765.152
R32 VDD.t77 VDD.t89 765.152
R33 VDD.t432 VDD.t199 765.152
R34 VDD.t69 VDD.t285 765.152
R35 VDD.t92 VDD.t79 765.152
R36 VDD.t8 VDD.t201 765.152
R37 VDD.t378 VDD.t196 765.152
R38 VDD.t332 VDD.t295 765.152
R39 VDD.t466 VDD.t38 765.152
R40 VDD.t5 VDD.t144 765.152
R41 VDD.t329 VDD.t292 765.152
R42 VDD.t228 VDD.t36 765.152
R43 VDD.t419 VDD.t312 765.152
R44 VDD.t478 VDD.t488 765.152
R45 VDD.t16 VDD.t447 765.152
R46 VDD.t130 VDD.t2 765.152
R47 VDD.t486 VDD.t481 765.152
R48 VDD.t449 VDD.t62 765.152
R49 VDD.t501 VDD.t385 765.152
R50 VDD.t257 VDD.t278 765.152
R51 VDD.t430 VDD.t337 765.152
R52 VDD.t319 VDD.t335 765.152
R53 VDD.t171 VDD.t497 765.152
R54 VDD.t346 VDD.t252 765.152
R55 VDD.t316 VDD.t182 765.152
R56 VDD.t495 VDD.t169 765.152
R57 VDD.t307 VDD.t393 765.152
R58 VDD.t470 VDD.t390 765.152
R59 VDD.t271 VDD.t29 765.152
R60 VDD.t75 VDD.t455 765.152
R61 VDD.t167 VDD.t472 765.152
R62 VDD.t189 VDD.t261 765.152
R63 VDD.t205 VDD.t174 765.152
R64 VDD.t475 VDD.t100 765.152
R65 VDD.t263 VDD.t187 765.152
R66 VDD.t220 VDD.t98 765.152
R67 VDD.t387 VDD.t290 765.152
R68 VDD.t31 VDD.t274 765.152
R69 VDD.t123 VDD.t203 765.152
R70 VDD.t504 VDD.t339 765.152
R71 VDD.t259 VDD.t276 765.152
R72 VDD.t400 VDD.t67 765.152
R73 VDD.t222 VDD.t359 765.152
R74 VDD.t53 VDD.t364 765.152
R75 VDD.t95 VDD.t353 765.152
R76 VDD.n233 VDD.t355 581.375
R77 VDD VDD.n233 572.967
R78 VDD.n428 VDD.t281 480.199
R79 VDD.t212 VDD.t440 461.096
R80 VDD.t212 VDD.t250 461.096
R81 VDD.t247 VDD.t120 461.096
R82 VDD.t304 VDD.t115 461.096
R83 VDD VDD.n374 429.187
R84 VDD VDD.n342 429.187
R85 VDD VDD.n359 429.187
R86 VDD.n421 VDD 427.092
R87 VDD VDD.n25 426.699
R88 VDD VDD.n129 426.699
R89 VDD VDD.n511 426.699
R90 VDD VDD.n14 426.699
R91 VDD.n144 VDD 424.618
R92 VDD VDD.n203 424.618
R93 VDD.n226 VDD.t149 420.793
R94 VDD.n143 VDD 418.495
R95 VDD VDD.n198 418.495
R96 VDD.n25 VDD.t381 386.365
R97 VDD.n129 VDD.t326 386.365
R98 VDD.n511 VDD.t138 386.365
R99 VDD.n374 VDD.t243 386.365
R100 VDD.n405 VDD.t267 386.365
R101 VDD.n359 VDD.t411 386.365
R102 VDD.n342 VDD.t493 386.365
R103 VDD.n14 VDD.t133 386.365
R104 VDD.n143 VDD.t288 378.788
R105 VDD.n198 VDD.t357 378.788
R106 VDD.t117 VDD.n409 375
R107 VDD.n406 VDD.n405 368.159
R108 VDD.n235 VDD.t247 351.586
R109 VDD.n208 VDD.t304 351.586
R110 VDD.n409 VDD.n407 343.137
R111 VDD.t184 VDD.n143 322.223
R112 VDD.t225 VDD.n198 322.223
R113 VDD.t143 VDD.n144 320.635
R114 VDD.n203 VDD.t315 320.635
R115 VDD.t469 VDD.n421 306.118
R116 VDD.t104 VDD.t85 303.031
R117 VDD.t285 VDD.t65 303.031
R118 VDD.t370 VDD.t92 303.031
R119 VDD.t43 VDD.t378 303.031
R120 VDD.t144 VDD.t48 303.031
R121 VDD.t21 VDD.t329 303.031
R122 VDD.t312 VDD.t233 303.031
R123 VDD.t395 VDD.t478 303.031
R124 VDD.t238 VDD.t130 303.031
R125 VDD.t59 VDD.t430 303.031
R126 VDD.t56 VDD.t346 303.031
R127 VDD.t397 VDD.t495 303.031
R128 VDD.t254 VDD.t307 303.031
R129 VDD.t455 VDD.t442 303.031
R130 VDD.t174 VDD.t457 303.031
R131 VDD.t23 VDD.t263 303.031
R132 VDD.t463 VDD.t220 303.031
R133 VDD.t372 VDD.t31 303.031
R134 VDD.t460 VDD.t123 303.031
R135 VDD.t26 VDD.t259 303.031
R136 VDD.t437 VDD.t400 303.031
R137 VDD.t359 VDD.t11 303.031
R138 VDD.t19 VDD.t53 303.031
R139 VDD.t322 VDD.t424 303.031
R140 VDD.n424 VDD.n412 298.536
R141 VDD.n428 VDD.n412 288
R142 VDD.n214 VDD.n213 199.562
R143 VDD.n218 VDD.n217 199.562
R144 VDD.n365 VDD.t427 193.183
R145 VDD.n366 VDD.t501 193.183
R146 VDD.n372 VDD.t278 193.183
R147 VDD.n373 VDD.t59 193.183
R148 VDD.n397 VDD.t348 193.183
R149 VDD.n399 VDD.t319 193.183
R150 VDD.n401 VDD.t171 193.183
R151 VDD.n404 VDD.t56 193.183
R152 VDD.n410 VDD.t117 193.183
R153 VDD.n376 VDD.t301 193.183
R154 VDD.n378 VDD.t316 193.183
R155 VDD.n381 VDD.t397 193.183
R156 VDD.n384 VDD.t254 193.183
R157 VDD.n346 VDD.t452 193.183
R158 VDD.n352 VDD.t390 193.183
R159 VDD.n353 VDD.t271 193.183
R160 VDD.n358 VDD.t442 193.183
R161 VDD.n329 VDD.t176 193.183
R162 VDD.n335 VDD.t472 193.183
R163 VDD.n336 VDD.t189 193.183
R164 VDD.n341 VDD.t457 193.183
R165 VDD.n308 VDD.t215 193.183
R166 VDD.n310 VDD.t475 193.183
R167 VDD.n313 VDD.t23 193.183
R168 VDD.n316 VDD.t463 193.183
R169 VDD.n280 VDD.t112 193.183
R170 VDD.n282 VDD.t387 193.183
R171 VDD.n285 VDD.t372 193.183
R172 VDD.n288 VDD.t460 193.183
R173 VDD.n252 VDD.t404 193.183
R174 VDD.n254 VDD.t504 193.183
R175 VDD.n257 VDD.t26 193.183
R176 VDD.n260 VDD.t437 193.183
R177 VDD.t85 VDD.n35 191.288
R178 VDD.n36 VDD.t77 191.288
R179 VDD.t199 VDD.n46 191.288
R180 VDD.n47 VDD.t102 191.288
R181 VDD.t65 VDD.n69 191.288
R182 VDD.n70 VDD.t370 191.288
R183 VDD.t201 VDD.n78 191.288
R184 VDD.n79 VDD.t324 191.288
R185 VDD.n128 VDD.t43 191.288
R186 VDD.n127 VDD.t295 191.288
R187 VDD.t38 VDD.n93 191.288
R188 VDD.n95 VDD.t231 191.288
R189 VDD.t48 VDD.n106 191.288
R190 VDD.n107 VDD.t21 191.288
R191 VDD.t36 VDD.n115 191.288
R192 VDD.n116 VDD.t141 191.288
R193 VDD.n136 VDD.t288 191.288
R194 VDD.t233 VDD.n492 191.288
R195 VDD.n493 VDD.t395 191.288
R196 VDD.t447 VDD.n501 191.288
R197 VDD.n502 VDD.t310 191.288
R198 VDD.n510 VDD.t238 191.288
R199 VDD.n509 VDD.t486 191.288
R200 VDD.n508 VDD.t449 191.288
R201 VDD.n507 VDD.t128 191.288
R202 VDD.n423 VDD.t407 191.288
R203 VDD.t357 VDD.n197 191.288
R204 VDD.t11 VDD.n182 191.288
R205 VDD.n183 VDD.t19 191.288
R206 VDD.t353 VDD.n191 191.288
R207 VDD.n192 VDD.t136 191.288
R208 VDD.n13 VDD.t322 191.288
R209 VDD.n153 VDD.t367 191.288
R210 VDD.n158 VDD.t351 191.288
R211 VDD.n163 VDD.t422 191.288
R212 VDD.t451 VDD.t309 175.631
R213 VDD.n213 VDD.t384 170.577
R214 VDD.n213 VDD.t218 170.577
R215 VDD.n217 VDD.t369 170.577
R216 VDD.n217 VDD.t344 170.577
R217 VDD.t415 VDD.n228 153.678
R218 VDD.t407 VDD.t209 151.516
R219 VDD.n145 VDD.t143 142.857
R220 VDD.t315 VDD.n201 142.857
R221 VDD.n409 VDD.t362 132.353
R222 VDD.n420 VDD.t269 124.511
R223 VDD.n424 VDD.n423 117.216
R224 VDD.n407 VDD.n406 112.746
R225 VDD.n35 VDD.t381 111.743
R226 VDD.n36 VDD.t179 111.743
R227 VDD.n46 VDD.t89 111.743
R228 VDD.n47 VDD.t432 111.743
R229 VDD.n69 VDD.t164 111.743
R230 VDD.n70 VDD.t69 111.743
R231 VDD.n78 VDD.t79 111.743
R232 VDD.n79 VDD.t8 111.743
R233 VDD.t326 VDD.n128 111.743
R234 VDD.t196 VDD.n127 111.743
R235 VDD.n93 VDD.t332 111.743
R236 VDD.n95 VDD.t466 111.743
R237 VDD.n106 VDD.t152 111.743
R238 VDD.n107 VDD.t5 111.743
R239 VDD.n115 VDD.t292 111.743
R240 VDD.n116 VDD.t228 111.743
R241 VDD.n136 VDD.t45 111.743
R242 VDD.n492 VDD.t160 111.743
R243 VDD.n493 VDD.t419 111.743
R244 VDD.n501 VDD.t488 111.743
R245 VDD.n502 VDD.t16 111.743
R246 VDD.t138 VDD.n510 111.743
R247 VDD.t2 VDD.n509 111.743
R248 VDD.t481 VDD.n508 111.743
R249 VDD.t62 VDD.n507 111.743
R250 VDD.n197 VDD.t13 111.743
R251 VDD.n182 VDD.t156 111.743
R252 VDD.n183 VDD.t222 111.743
R253 VDD.n191 VDD.t364 111.743
R254 VDD.n192 VDD.t95 111.743
R255 VDD.t133 VDD.n13 111.743
R256 VDD.n153 VDD.t125 111.743
R257 VDD.n158 VDD.t50 111.743
R258 VDD.n163 VDD.t107 111.743
R259 VDD.n145 VDD.t184 111.112
R260 VDD.n201 VDD.t225 111.112
R261 VDD.t385 VDD.n365 109.849
R262 VDD.n366 VDD.t257 109.849
R263 VDD.t337 VDD.n372 109.849
R264 VDD.t243 VDD.n373 109.849
R265 VDD.t335 VDD.n397 109.849
R266 VDD.t497 VDD.n399 109.849
R267 VDD.t252 VDD.n401 109.849
R268 VDD.t267 VDD.n404 109.849
R269 VDD.n410 VDD.t207 109.849
R270 VDD.t182 VDD.n376 109.849
R271 VDD.t169 VDD.n378 109.849
R272 VDD.t393 VDD.n381 109.849
R273 VDD.n384 VDD.t265 109.849
R274 VDD.n346 VDD.t470 109.849
R275 VDD.t29 VDD.n352 109.849
R276 VDD.n353 VDD.t75 109.849
R277 VDD.t411 VDD.n358 109.849
R278 VDD.n329 VDD.t167 109.849
R279 VDD.t261 VDD.n335 109.849
R280 VDD.n336 VDD.t205 109.849
R281 VDD.t493 VDD.n341 109.849
R282 VDD.t100 VDD.n308 109.849
R283 VDD.t187 VDD.n310 109.849
R284 VDD.t98 VDD.n313 109.849
R285 VDD.n316 VDD.t491 109.849
R286 VDD.t290 VDD.n280 109.849
R287 VDD.t274 VDD.n282 109.849
R288 VDD.t203 VDD.n285 109.849
R289 VDD.n288 VDD.t409 109.849
R290 VDD.t339 VDD.n252 109.849
R291 VDD.t276 VDD.n254 109.849
R292 VDD.t67 VDD.n257 109.849
R293 VDD.n260 VDD.t297 109.849
R294 VDD.t209 VDD.n419 96.5914
R295 VDD.n422 VDD.n420 90.2261
R296 VDD.n233 VDD.t499 80.0005
R297 VDD.n422 VDD.t469 76.2337
R298 VDD.t484 VDD 68.2053
R299 VDD.n226 VDD 65.7064
R300 VDD.n25 VDD.t82 62.1896
R301 VDD.n129 VDD.t40 62.1896
R302 VDD.n511 VDD.t240 62.1896
R303 VDD.n14 VDD.t235 62.1896
R304 VDD.n241 VDD.t402 61.9053
R305 VDD.n144 VDD.t72 61.8817
R306 VDD.n203 VDD.t341 61.8817
R307 VDD VDD.n406 61.0269
R308 VDD.n143 VDD.t33 60.9761
R309 VDD.n198 VDD.t375 60.9761
R310 VDD.n374 VDD.t417 59.702
R311 VDD.n405 VDD.t413 59.702
R312 VDD.n359 VDD.t445 59.702
R313 VDD.n342 VDD.t435 59.702
R314 VDD.n421 VDD.t0 59.4064
R315 VDD.n229 VDD.t87 55.0852
R316 VDD.t355 VDD.n232 55.0852
R317 VDD.n419 VDD.t110 54.9247
R318 VDD.n56 VDD.t151 30.9379
R319 VDD.n170 VDD.t159 30.9379
R320 VDD.n59 VDD.t163 30.2877
R321 VDD.n173 VDD.t155 30.2877
R322 VDD.n60 VDD.t510 24.5101
R323 VDD.n56 VDD.t507 24.5101
R324 VDD.n172 VDD.t513 24.5101
R325 VDD.n170 VDD.t511 24.5101
R326 VDD.n228 VDD.t451 21.9544
R327 VDD.n423 VDD.n422 20.147
R328 VDD.n224 VDD.t356 14.0055
R329 VDD.n227 VDD.t416 13.2223
R330 VDD.n230 VDD.t88 12.3869
R331 VDD.n219 VDD.t485 12.3869
R332 VDD.n224 VDD.t500 10.1341
R333 VDD.n426 VDD.n425 9.64171
R334 VDD.n174 VDD.n171 8.14131
R335 VDD.n58 VDD.n57 8.14083
R336 VDD.n61 VDD.n60 8.0005
R337 VDD.n427 VDD.n426 6.69176
R338 VDD.n35 VDD.n34 6.3005
R339 VDD.n37 VDD.n36 6.3005
R340 VDD.n46 VDD.n45 6.3005
R341 VDD.n48 VDD.n47 6.3005
R342 VDD.n69 VDD.n68 6.3005
R343 VDD.n71 VDD.n70 6.3005
R344 VDD.n78 VDD.n77 6.3005
R345 VDD.n80 VDD.n79 6.3005
R346 VDD.n106 VDD.n105 6.3005
R347 VDD.n108 VDD.n107 6.3005
R348 VDD.n115 VDD.n114 6.3005
R349 VDD.n117 VDD.n116 6.3005
R350 VDD.n127 VDD.n126 6.3005
R351 VDD.n123 VDD.n93 6.3005
R352 VDD.n120 VDD.n95 6.3005
R353 VDD.n128 VDD.n85 6.3005
R354 VDD.n137 VDD.n136 6.3005
R355 VDD.n146 VDD.n145 6.3005
R356 VDD.n492 VDD.n491 6.3005
R357 VDD.n494 VDD.n493 6.3005
R358 VDD.n501 VDD.n500 6.3005
R359 VDD.n503 VDD.n502 6.3005
R360 VDD.n509 VDD.n474 6.3005
R361 VDD.n508 VDD.n478 6.3005
R362 VDD.n507 VDD.n506 6.3005
R363 VDD VDD.n428 6.3005
R364 VDD.n430 VDD.n412 6.3005
R365 VDD VDD.n424 6.3005
R366 VDD.n433 VDD.n410 6.3005
R367 VDD VDD.n407 6.3005
R368 VDD.n385 VDD.n384 6.3005
R369 VDD.n388 VDD.n381 6.3005
R370 VDD.n391 VDD.n378 6.3005
R371 VDD.n394 VDD.n376 6.3005
R372 VDD.n447 VDD.n397 6.3005
R373 VDD.n444 VDD.n399 6.3005
R374 VDD.n441 VDD.n401 6.3005
R375 VDD.n438 VDD.n404 6.3005
R376 VDD.n317 VDD.n316 6.3005
R377 VDD.n320 VDD.n313 6.3005
R378 VDD.n323 VDD.n310 6.3005
R379 VDD.n326 VDD.n308 6.3005
R380 VDD.n330 VDD.n329 6.3005
R381 VDD.n335 VDD.n334 6.3005
R382 VDD.n337 VDD.n336 6.3005
R383 VDD.n341 VDD.n340 6.3005
R384 VDD.n289 VDD.n288 6.3005
R385 VDD.n292 VDD.n285 6.3005
R386 VDD.n295 VDD.n282 6.3005
R387 VDD.n298 VDD.n280 6.3005
R388 VDD.n347 VDD.n346 6.3005
R389 VDD.n352 VDD.n351 6.3005
R390 VDD.n354 VDD.n353 6.3005
R391 VDD.n358 VDD.n357 6.3005
R392 VDD.n261 VDD.n260 6.3005
R393 VDD.n264 VDD.n257 6.3005
R394 VDD.n267 VDD.n254 6.3005
R395 VDD.n270 VDD.n252 6.3005
R396 VDD.n365 VDD.n364 6.3005
R397 VDD.n367 VDD.n366 6.3005
R398 VDD.n372 VDD.n371 6.3005
R399 VDD.n452 VDD.n373 6.3005
R400 VDD.n228 VDD.n227 6.3005
R401 VDD VDD.n229 6.3005
R402 VDD.n232 VDD.n231 6.3005
R403 VDD.n242 VDD.n241 6.3005
R404 VDD.n212 VDD 6.3005
R405 VDD.n216 VDD 6.3005
R406 VDD.n463 VDD.n197 6.3005
R407 VDD.n459 VDD.n201 6.3005
R408 VDD.n510 VDD.n468 6.3005
R409 VDD.n182 VDD.n181 6.3005
R410 VDD.n184 VDD.n183 6.3005
R411 VDD.n191 VDD.n190 6.3005
R412 VDD.n193 VDD.n192 6.3005
R413 VDD.n13 VDD.n12 6.3005
R414 VDD.n154 VDD.n153 6.3005
R415 VDD.n159 VDD.n158 6.3005
R416 VDD.n518 VDD.n163 6.3005
R417 VDD.n234 VDD.t193 5.85907
R418 VDD.n142 VDD.n139 5.85007
R419 VDD.n461 VDD.n199 5.85007
R420 VDD.n454 VDD.n453 5.69603
R421 VDD.n105 VDD.n101 5.213
R422 VDD.n491 VDD.n487 5.213
R423 VDD.n385 VDD.t266 5.213
R424 VDD.n317 VDD.t492 5.213
R425 VDD.n289 VDD.t410 5.213
R426 VDD.n261 VDD.t298 5.213
R427 VDD.n26 VDD.n23 5.17567
R428 VDD.n43 VDD.n42 5.17567
R429 VDD VDD.n24 5.16369
R430 VDD.n432 VDD.t208 5.15377
R431 VDD.n84 VDD.n83 5.13287
R432 VDD.n44 VDD.t200 5.13287
R433 VDD.n39 VDD.t78 5.13287
R434 VDD.n40 VDD.n21 5.13287
R435 VDD.n30 VDD.n29 5.13287
R436 VDD.n49 VDD.t103 5.13287
R437 VDD.n54 VDD.n53 5.13287
R438 VDD.n73 VDD.n50 5.13287
R439 VDD.n76 VDD.t202 5.13287
R440 VDD.n75 VDD.n74 5.13287
R441 VDD.n81 VDD.t325 5.13287
R442 VDD.n91 VDD.n86 5.13287
R443 VDD.n125 VDD.t296 5.13287
R444 VDD.n124 VDD.n92 5.13287
R445 VDD.n122 VDD.t39 5.13287
R446 VDD.n121 VDD.n94 5.13287
R447 VDD.n119 VDD.t232 5.13287
R448 VDD.n100 VDD.n99 5.13287
R449 VDD.n110 VDD.n96 5.13287
R450 VDD.n113 VDD.t37 5.13287
R451 VDD.n112 VDD.n111 5.13287
R452 VDD.n118 VDD.t142 5.13287
R453 VDD.n135 VDD.n18 5.13287
R454 VDD.n138 VDD.t289 5.13287
R455 VDD.n473 VDD.n472 5.13287
R456 VDD.n476 VDD.t487 5.13287
R457 VDD.n477 VDD.n475 5.13287
R458 VDD.n480 VDD.t450 5.13287
R459 VDD.n481 VDD.n479 5.13287
R460 VDD.n505 VDD.t129 5.13287
R461 VDD.n486 VDD.n485 5.13287
R462 VDD.n496 VDD.n482 5.13287
R463 VDD.n499 VDD.t448 5.13287
R464 VDD.n498 VDD.n497 5.13287
R465 VDD.n504 VDD.t311 5.13287
R466 VDD.n434 VDD.n408 5.13287
R467 VDD.n416 VDD.n415 5.13287
R468 VDD.n417 VDD.t122 5.13287
R469 VDD.n417 VDD.t111 5.13287
R470 VDD.n437 VDD.t268 5.13287
R471 VDD.n440 VDD.t253 5.13287
R472 VDD.n442 VDD.n400 5.13287
R473 VDD.n443 VDD.t498 5.13287
R474 VDD.n445 VDD.n398 5.13287
R475 VDD.n446 VDD.t336 5.13287
R476 VDD.n448 VDD.n396 5.13287
R477 VDD.n387 VDD.t394 5.13287
R478 VDD.n390 VDD.t170 5.13287
R479 VDD.n392 VDD.n377 5.13287
R480 VDD.n393 VDD.t183 5.13287
R481 VDD.n395 VDD.n375 5.13287
R482 VDD.n300 VDD.t494 5.13287
R483 VDD.n338 VDD.t206 5.13287
R484 VDD.n304 VDD.n303 5.13287
R485 VDD.n333 VDD.t262 5.13287
R486 VDD.n332 VDD.n305 5.13287
R487 VDD.n331 VDD.t168 5.13287
R488 VDD.n328 VDD.n306 5.13287
R489 VDD.n319 VDD.t99 5.13287
R490 VDD.n322 VDD.t188 5.13287
R491 VDD.n324 VDD.n309 5.13287
R492 VDD.n325 VDD.t101 5.13287
R493 VDD.n327 VDD.n307 5.13287
R494 VDD.n291 VDD.t204 5.13287
R495 VDD.n294 VDD.t275 5.13287
R496 VDD.n296 VDD.n281 5.13287
R497 VDD.n297 VDD.t291 5.13287
R498 VDD.n299 VDD.n279 5.13287
R499 VDD.n272 VDD.t412 5.13287
R500 VDD.n355 VDD.t76 5.13287
R501 VDD.n276 VDD.n275 5.13287
R502 VDD.n350 VDD.t30 5.13287
R503 VDD.n349 VDD.n277 5.13287
R504 VDD.n348 VDD.t471 5.13287
R505 VDD.n345 VDD.n278 5.13287
R506 VDD.n451 VDD.t244 5.13287
R507 VDD.n370 VDD.t338 5.13287
R508 VDD.n369 VDD.n247 5.13287
R509 VDD.n368 VDD.t258 5.13287
R510 VDD.n249 VDD.n248 5.13287
R511 VDD.n363 VDD.t386 5.13287
R512 VDD.n362 VDD.n250 5.13287
R513 VDD.n263 VDD.t68 5.13287
R514 VDD.n266 VDD.t277 5.13287
R515 VDD.n268 VDD.n253 5.13287
R516 VDD.n269 VDD.t340 5.13287
R517 VDD.n271 VDD.n251 5.13287
R518 VDD.n237 VDD.t121 5.13287
R519 VDD.n223 VDD.n222 5.13287
R520 VDD.n240 VDD.t251 5.13287
R521 VDD.n210 VDD.t116 5.13287
R522 VDD.n206 VDD.n205 5.13287
R523 VDD.n464 VDD.n196 5.13287
R524 VDD.n462 VDD.t358 5.13287
R525 VDD.n512 VDD.n469 5.13287
R526 VDD.n168 VDD.n167 5.13287
R527 VDD.n186 VDD.n164 5.13287
R528 VDD.n189 VDD.t354 5.13287
R529 VDD.n188 VDD.n187 5.13287
R530 VDD.n194 VDD.t137 5.13287
R531 VDD.n6 VDD.n5 5.13287
R532 VDD.n152 VDD.n4 5.13287
R533 VDD.n155 VDD.t368 5.13287
R534 VDD.n157 VDD.n2 5.13287
R535 VDD.n160 VDD.t352 5.13287
R536 VDD.n162 VDD.n0 5.13287
R537 VDD.n517 VDD.t423 5.13287
R538 VDD.n15 VDD.n11 5.12213
R539 VDD VDD.t150 5.10424
R540 VDD.n130 VDD.n82 5.09407
R541 VDD.n17 VDD.n16 5.09407
R542 VDD.n425 VDD.t270 5.09407
R543 VDD.n427 VDD.t282 5.09407
R544 VDD.n411 VDD.t1 5.09407
R545 VDD.n435 VDD.t363 5.09407
R546 VDD.n436 VDD.t414 5.09407
R547 VDD.n450 VDD.t418 5.09407
R548 VDD.n343 VDD.t436 5.09407
R549 VDD.n360 VDD.t446 5.09407
R550 VDD.n207 VDD.t284 5.09407
R551 VDD.n211 VDD.t148 5.09407
R552 VDD.n215 VDD.t246 5.09407
R553 VDD.n204 VDD.n202 5.09407
R554 VDD.n471 VDD.n470 5.09407
R555 VDD.n243 VDD.t403 4.9655
R556 VDD.n64 VDD.n63 4.8755
R557 VDD.n177 VDD.n176 4.8755
R558 VDD.n214 VDD.t219 4.40826
R559 VDD.n218 VDD.t345 4.3915
R560 VDD.n212 VDD.t147 4.26489
R561 VDD.n216 VDD.t245 4.26489
R562 VDD.n141 VDD.n140 4.12326
R563 VDD.n460 VDD.n200 4.12326
R564 VDD.n429 VDD.t195 4.11379
R565 VDD.n344 VDD.n299 3.90405
R566 VDD.n458 VDD.n457 3.33671
R567 VDD.n419 VDD.n418 3.1505
R568 VDD.n33 VDD.n28 2.85787
R569 VDD.n67 VDD.n66 2.85787
R570 VDD.n72 VDD.n52 2.85787
R571 VDD.n90 VDD.n88 2.85787
R572 VDD.n104 VDD.n103 2.85787
R573 VDD.n109 VDD.n98 2.85787
R574 VDD.n467 VDD.n466 2.85787
R575 VDD.n490 VDD.n489 2.85787
R576 VDD.n495 VDD.n484 2.85787
R577 VDD.n416 VDD.n414 2.85787
R578 VDD.n439 VDD.n403 2.85787
R579 VDD.n386 VDD.n383 2.85787
R580 VDD.n389 VDD.n380 2.85787
R581 VDD.n339 VDD.n302 2.85787
R582 VDD.n318 VDD.n315 2.85787
R583 VDD.n321 VDD.n312 2.85787
R584 VDD.n290 VDD.n287 2.85787
R585 VDD.n293 VDD.n284 2.85787
R586 VDD.n356 VDD.n274 2.85787
R587 VDD.n246 VDD.n245 2.85787
R588 VDD.n262 VDD.n259 2.85787
R589 VDD.n265 VDD.n256 2.85787
R590 VDD.n238 VDD.n221 2.85787
R591 VDD.n180 VDD.n179 2.85787
R592 VDD.n185 VDD.n166 2.85787
R593 VDD.n9 VDD.n8 2.85787
R594 VDD.n28 VDD.t86 2.2755
R595 VDD.n28 VDD.n27 2.2755
R596 VDD.n66 VDD.t66 2.2755
R597 VDD.n66 VDD.n65 2.2755
R598 VDD.n52 VDD.t371 2.2755
R599 VDD.n52 VDD.n51 2.2755
R600 VDD.n88 VDD.t44 2.2755
R601 VDD.n88 VDD.n87 2.2755
R602 VDD.n103 VDD.t49 2.2755
R603 VDD.n103 VDD.n102 2.2755
R604 VDD.n98 VDD.t22 2.2755
R605 VDD.n98 VDD.n97 2.2755
R606 VDD.n466 VDD.t239 2.2755
R607 VDD.n466 VDD.n465 2.2755
R608 VDD.n489 VDD.t234 2.2755
R609 VDD.n489 VDD.n488 2.2755
R610 VDD.n484 VDD.t396 2.2755
R611 VDD.n484 VDD.n483 2.2755
R612 VDD.n414 VDD.t408 2.2755
R613 VDD.n414 VDD.n413 2.2755
R614 VDD.n403 VDD.t347 2.2755
R615 VDD.n403 VDD.n402 2.2755
R616 VDD.n383 VDD.t308 2.2755
R617 VDD.n383 VDD.n382 2.2755
R618 VDD.n380 VDD.t496 2.2755
R619 VDD.n380 VDD.n379 2.2755
R620 VDD.n302 VDD.t175 2.2755
R621 VDD.n302 VDD.n301 2.2755
R622 VDD.n315 VDD.t221 2.2755
R623 VDD.n315 VDD.n314 2.2755
R624 VDD.n312 VDD.t264 2.2755
R625 VDD.n312 VDD.n311 2.2755
R626 VDD.n287 VDD.t124 2.2755
R627 VDD.n287 VDD.n286 2.2755
R628 VDD.n284 VDD.t32 2.2755
R629 VDD.n284 VDD.n283 2.2755
R630 VDD.n274 VDD.t456 2.2755
R631 VDD.n274 VDD.n273 2.2755
R632 VDD.n245 VDD.t431 2.2755
R633 VDD.n245 VDD.n244 2.2755
R634 VDD.n259 VDD.t401 2.2755
R635 VDD.n259 VDD.n258 2.2755
R636 VDD.n256 VDD.t260 2.2755
R637 VDD.n256 VDD.n255 2.2755
R638 VDD.n221 VDD.t441 2.2755
R639 VDD.n221 VDD.n220 2.2755
R640 VDD.n179 VDD.t12 2.2755
R641 VDD.n179 VDD.n178 2.2755
R642 VDD.n166 VDD.t20 2.2755
R643 VDD.n166 VDD.n165 2.2755
R644 VDD.n8 VDD.t323 2.2755
R645 VDD.n8 VDD.n7 2.2755
R646 VDD.n437 VDD 2.25904
R647 VDD.n57 VDD.n56 2.11346
R648 VDD.n171 VDD.n170 2.11346
R649 VDD.n174 VDD.n173 1.8236
R650 VDD.n59 VDD.n58 1.82345
R651 VDD VDD.n84 1.81843
R652 VDD.n512 VDD 1.81843
R653 VDD.n26 VDD 1.79694
R654 VDD.n119 VDD.n118 1.16051
R655 VDD.n505 VDD.n504 1.16051
R656 VDD.n195 VDD.n194 1.0737
R657 VDD.n449 VDD.n395 1.02928
R658 VDD.n361 VDD.n271 1.02928
R659 VDD.n131 VDD.n81 1.02347
R660 VDD.n328 VDD.n327 0.881662
R661 VDD VDD.n240 0.786716
R662 VDD.n420 VDD.t194 0.783764
R663 VDD.n31 VDD.n26 0.682778
R664 VDD.n456 VDD.n211 0.66512
R665 VDD.n455 VDD.n215 0.634017
R666 VDD.n177 VDD.n175 0.608132
R667 VDD.n148 VDD.n15 0.601963
R668 VDD.n32 VDD.n31 0.582756
R669 VDD.n43 VDD.n19 0.582756
R670 VDD.n149 VDD.n10 0.582756
R671 VDD.n151 VDD.n150 0.582756
R672 VDD.n41 VDD.n20 0.5405
R673 VDD.n38 VDD.n22 0.5405
R674 VDD.n133 VDD.n132 0.5405
R675 VDD.n156 VDD.n3 0.5405
R676 VDD.n161 VDD.n1 0.5405
R677 VDD.n516 VDD.n515 0.5405
R678 VDD.n89 VDD 0.468385
R679 VDD VDD.n513 0.468385
R680 VDD.n60 VDD.n59 0.404541
R681 VDD.n173 VDD.n172 0.404541
R682 VDD.n68 VDD.n64 0.337997
R683 VDD.n181 VDD.n177 0.337997
R684 VDD.n64 VDD.n62 0.328132
R685 VDD.n67 VDD.n54 0.233919
R686 VDD.n73 VDD.n72 0.233919
R687 VDD.n104 VDD.n100 0.233919
R688 VDD.n110 VDD.n109 0.233919
R689 VDD.n490 VDD.n486 0.233919
R690 VDD.n496 VDD.n495 0.233919
R691 VDD.n390 VDD.n389 0.233919
R692 VDD.n387 VDD.n386 0.233919
R693 VDD.n322 VDD.n321 0.233919
R694 VDD.n319 VDD.n318 0.233919
R695 VDD.n294 VDD.n293 0.233919
R696 VDD.n291 VDD.n290 0.233919
R697 VDD.n266 VDD.n265 0.233919
R698 VDD.n263 VDD.n262 0.233919
R699 VDD.n180 VDD.n168 0.233919
R700 VDD.n186 VDD.n185 0.233919
R701 VDD VDD.n454 0.227487
R702 VDD.n431 VDD.n430 0.224447
R703 VDD.n134 VDD 0.223897
R704 VDD.n514 VDD 0.223897
R705 VDD.n436 VDD 0.205357
R706 VDD.n432 VDD.n431 0.202146
R707 VDD.n515 VDD.n514 0.178009
R708 VDD.n207 VDD.n206 0.170231
R709 VDD.n450 VDD.n449 0.167533
R710 VDD VDD.n272 0.160716
R711 VDD.n134 VDD.n133 0.159769
R712 VDD.n451 VDD 0.158984
R713 VDD VDD.n300 0.157289
R714 VDD.n361 VDD.n360 0.155496
R715 VDD VDD.n225 0.154766
R716 VDD.n344 VDD.n343 0.154581
R717 VDD.n40 VDD.n39 0.141016
R718 VDD.n76 VDD.n75 0.141016
R719 VDD.n113 VDD.n112 0.141016
R720 VDD.n125 VDD.n124 0.141016
R721 VDD.n122 VDD.n121 0.141016
R722 VDD.n499 VDD.n498 0.141016
R723 VDD.n477 VDD.n476 0.141016
R724 VDD.n481 VDD.n480 0.141016
R725 VDD.n393 VDD.n392 0.141016
R726 VDD.n325 VDD.n324 0.141016
R727 VDD.n297 VDD.n296 0.141016
R728 VDD.n269 VDD.n268 0.141016
R729 VDD.n189 VDD.n188 0.141016
R730 VDD.n131 VDD.n130 0.139745
R731 VDD.n471 VDD.n195 0.139745
R732 VDD VDD.n147 0.138536
R733 VDD.n147 VDD.n17 0.137219
R734 VDD.n458 VDD.n204 0.137219
R735 VDD.n431 VDD.n411 0.137126
R736 VDD.n345 VDD.n344 0.131861
R737 VDD.n435 VDD.n434 0.130567
R738 VDD.n457 VDD.n210 0.129503
R739 VDD.n457 VDD 0.12689
R740 VDD.n446 VDD.n445 0.123551
R741 VDD.n443 VDD.n442 0.123551
R742 VDD.n349 VDD.n348 0.123551
R743 VDD.n350 VDD.n276 0.123551
R744 VDD.n91 VDD 0.123016
R745 VDD.n473 VDD 0.123016
R746 VDD.n363 VDD.n249 0.122176
R747 VDD.n369 VDD.n368 0.122176
R748 VDD.n332 VDD.n331 0.120831
R749 VDD.n333 VDD.n304 0.120831
R750 VDD.n3 VDD.n1 0.119765
R751 VDD.n449 VDD.n448 0.116432
R752 VDD.n456 VDD.n455 0.115201
R753 VDD.n362 VDD.n361 0.115137
R754 VDD VDD.n90 0.111403
R755 VDD VDD.n467 0.111403
R756 VDD.n9 VDD 0.111403
R757 VDD.n44 VDD.n43 0.109081
R758 VDD.n132 VDD.n49 0.107919
R759 VDD.n57 VDD 0.107393
R760 VDD.n171 VDD 0.107393
R761 VDD.n45 VDD.n44 0.107339
R762 VDD.n49 VDD.n48 0.107339
R763 VDD.n77 VDD.n76 0.107339
R764 VDD.n81 VDD.n80 0.107339
R765 VDD.n114 VDD.n113 0.107339
R766 VDD.n118 VDD.n117 0.107339
R767 VDD.n126 VDD.n125 0.107339
R768 VDD.n123 VDD.n122 0.107339
R769 VDD.n120 VDD.n119 0.107339
R770 VDD.n500 VDD.n499 0.107339
R771 VDD.n504 VDD.n503 0.107339
R772 VDD.n476 VDD.n474 0.107339
R773 VDD.n480 VDD.n478 0.107339
R774 VDD.n506 VDD.n505 0.107339
R775 VDD.n434 VDD.n433 0.107339
R776 VDD.n395 VDD.n394 0.107339
R777 VDD.n392 VDD.n391 0.107339
R778 VDD.n327 VDD.n326 0.107339
R779 VDD.n324 VDD.n323 0.107339
R780 VDD.n299 VDD.n298 0.107339
R781 VDD.n296 VDD.n295 0.107339
R782 VDD.n271 VDD.n270 0.107339
R783 VDD.n268 VDD.n267 0.107339
R784 VDD.n209 VDD.n206 0.107339
R785 VDD.n190 VDD.n189 0.107339
R786 VDD.n194 VDD.n193 0.107339
R787 VDD.n155 VDD.n154 0.107339
R788 VDD.n160 VDD.n159 0.107339
R789 VDD.n518 VDD.n517 0.107339
R790 VDD.n20 VDD.n19 0.107337
R791 VDD.n440 VDD 0.10728
R792 VDD VDD.n355 0.10728
R793 VDD VDD.n33 0.106758
R794 VDD VDD.n67 0.106758
R795 VDD.n72 VDD 0.106758
R796 VDD VDD.n104 0.106758
R797 VDD.n109 VDD 0.106758
R798 VDD VDD.n490 0.106758
R799 VDD.n495 VDD 0.106758
R800 VDD VDD.n180 0.106758
R801 VDD.n185 VDD 0.106758
R802 VDD.n389 VDD 0.106177
R803 VDD.n386 VDD 0.106177
R804 VDD.n321 VDD 0.106177
R805 VDD.n318 VDD 0.106177
R806 VDD.n293 VDD 0.106177
R807 VDD.n290 VDD 0.106177
R808 VDD.n265 VDD 0.106177
R809 VDD.n262 VDD 0.106177
R810 VDD.n370 VDD 0.106087
R811 VDD VDD.n338 0.10492
R812 VDD.n150 VDD.n3 0.10413
R813 VDD.n157 VDD.n156 0.100371
R814 VDD.n169 VDD 0.100075
R815 VDD.n148 VDD 0.09952
R816 VDD VDD.n439 0.0981271
R817 VDD.n356 VDD 0.0981271
R818 VDD VDD.n246 0.0970363
R819 VDD.n133 VDD.n19 0.0967138
R820 VDD.n456 VDD.n214 0.096125
R821 VDD.n339 VDD 0.0959696
R822 VDD.n150 VDD.n149 0.0947094
R823 VDD.n448 VDD.n447 0.0940593
R824 VDD.n445 VDD.n444 0.0940593
R825 VDD.n442 VDD.n441 0.0940593
R826 VDD.n347 VDD.n345 0.0940593
R827 VDD.n351 VDD.n349 0.0940593
R828 VDD.n354 VDD.n276 0.0940593
R829 VDD.n439 VDD 0.0930424
R830 VDD VDD.n356 0.0930424
R831 VDD.n364 VDD.n362 0.093014
R832 VDD.n367 VDD.n249 0.093014
R833 VDD.n371 VDD.n369 0.093014
R834 VDD.n330 VDD.n328 0.0919917
R835 VDD.n334 VDD.n332 0.0919917
R836 VDD.n337 VDD.n304 0.0919917
R837 VDD VDD.n339 0.0909972
R838 VDD.n455 VDD.n218 0.0905
R839 VDD.n516 VDD.n195 0.089386
R840 VDD.n162 VDD.n161 0.082371
R841 VDD.n33 VDD.n32 0.0817903
R842 VDD.n149 VDD.n148 0.08148
R843 VDD.n31 VDD.n22 0.0808786
R844 VDD.n22 VDD.n20 0.0808786
R845 VDD.n71 VDD.n54 0.080629
R846 VDD.n108 VDD.n100 0.080629
R847 VDD.n494 VDD.n486 0.080629
R848 VDD.n388 VDD.n387 0.080629
R849 VDD.n320 VDD.n319 0.080629
R850 VDD.n292 VDD.n291 0.080629
R851 VDD.n264 VDD.n263 0.080629
R852 VDD.n184 VDD.n168 0.080629
R853 VDD VDD.n393 0.0794677
R854 VDD VDD.n390 0.0794677
R855 VDD VDD.n325 0.0794677
R856 VDD VDD.n322 0.0794677
R857 VDD VDD.n297 0.0794677
R858 VDD VDD.n294 0.0794677
R859 VDD VDD.n269 0.0794677
R860 VDD VDD.n266 0.0794677
R861 VDD.n30 VDD 0.0788871
R862 VDD VDD.n73 0.0788871
R863 VDD.n75 VDD 0.0788871
R864 VDD VDD.n110 0.0788871
R865 VDD.n112 VDD 0.0788871
R866 VDD VDD.n91 0.0788871
R867 VDD.n124 VDD 0.0788871
R868 VDD.n121 VDD 0.0788871
R869 VDD VDD.n496 0.0788871
R870 VDD.n498 VDD 0.0788871
R871 VDD VDD.n473 0.0788871
R872 VDD VDD.n477 0.0788871
R873 VDD VDD.n481 0.0788871
R874 VDD VDD.n186 0.0788871
R875 VDD.n188 VDD 0.0788871
R876 VDD VDD.n152 0.0788871
R877 VDD VDD.n157 0.0788871
R878 VDD VDD.n162 0.0788871
R879 VDD VDD.n225 0.0786971
R880 VDD.n210 VDD 0.0759839
R881 VDD.n425 VDD 0.0709717
R882 VDD VDD.n411 0.0709717
R883 VDD VDD.n436 0.0709717
R884 VDD VDD.n207 0.0709717
R885 VDD VDD.n211 0.0709717
R886 VDD VDD.n215 0.0709717
R887 VDD.n438 VDD.n437 0.0706695
R888 VDD.n357 VDD.n272 0.0706695
R889 VDD.n130 VDD 0.0701226
R890 VDD VDD.n17 0.0701226
R891 VDD.n204 VDD 0.0701226
R892 VDD VDD.n471 0.0701226
R893 VDD.n234 VDD 0.0700788
R894 VDD.n452 VDD.n451 0.0698855
R895 VDD VDD.n446 0.0696525
R896 VDD VDD.n443 0.0696525
R897 VDD VDD.n440 0.0696525
R898 VDD.n348 VDD 0.0696525
R899 VDD VDD.n350 0.0696525
R900 VDD.n355 VDD 0.0696525
R901 VDD.n340 VDD.n300 0.0691188
R902 VDD.n55 VDD 0.0690714
R903 VDD VDD.n363 0.0688799
R904 VDD.n368 VDD 0.0688799
R905 VDD VDD.n370 0.0688799
R906 VDD.n331 VDD 0.0681243
R907 VDD VDD.n333 0.0681243
R908 VDD.n338 VDD 0.0681243
R909 VDD.n10 VDD.n9 0.0649516
R910 VDD.n147 VDD.n146 0.0617883
R911 VDD.n459 VDD.n458 0.0617883
R912 VDD.n142 VDD.n141 0.0608681
R913 VDD.n461 VDD.n460 0.0608681
R914 VDD.n238 VDD.n237 0.0598378
R915 VDD VDD.n138 0.0592117
R916 VDD.n462 VDD 0.0592117
R917 VDD.n39 VDD.n38 0.0591452
R918 VDD.n161 VDD.n160 0.0591452
R919 VDD.n32 VDD.n30 0.0574032
R920 VDD.n89 VDD.n84 0.0556613
R921 VDD.n513 VDD.n512 0.0556613
R922 VDD VDD.n429 0.0555633
R923 VDD VDD.n432 0.0550806
R924 VDD.n517 VDD.n516 0.0550806
R925 VDD VDD.n416 0.0533387
R926 VDD.n453 VDD.n246 0.0532933
R927 VDD.n38 VDD.n37 0.0486936
R928 VDD.n62 VDD.n55 0.0471071
R929 VDD VDD.n41 0.0452097
R930 VDD VDD.n435 0.043431
R931 VDD.n90 VDD.n89 0.0417258
R932 VDD.n513 VDD.n467 0.0417258
R933 VDD.n156 VDD.n155 0.0411452
R934 VDD VDD.n224 0.041
R935 VDD.n360 VDD 0.0404465
R936 VDD VDD.n450 0.0400238
R937 VDD.n343 VDD 0.0396099
R938 VDD.n453 VDD 0.0392151
R939 VDD.n61 VDD.n58 0.0387493
R940 VDD VDD.n417 0.0382419
R941 VDD.n62 VDD.n61 0.0358571
R942 VDD.n175 VDD.n174 0.0344878
R943 VDD.n426 VDD.n416 0.0344677
R944 VDD.n138 VDD.n137 0.034365
R945 VDD.n463 VDD.n462 0.034365
R946 VDD.n41 VDD.n40 0.0341774
R947 VDD VDD.n223 0.0333767
R948 VDD.n231 VDD.n230 0.0327683
R949 VDD VDD.n427 0.032019
R950 VDD.n132 VDD.n131 0.0292131
R951 VDD.n230 VDD 0.028378
R952 VDD.n10 VDD.n6 0.0277903
R953 VDD.n141 VDD 0.0270031
R954 VDD.n460 VDD 0.0270031
R955 VDD.n152 VDD.n151 0.0254677
R956 VDD.n242 VDD.n219 0.0254153
R957 VDD VDD.n135 0.0242423
R958 VDD.n464 VDD 0.0242423
R959 VDD.n135 VDD.n134 0.0235061
R960 VDD.n514 VDD.n464 0.0235061
R961 VDD VDD.n219 0.0220254
R962 VDD.n89 VDD.n85 0.0206923
R963 VDD.n513 VDD.n468 0.0206923
R964 VDD.n12 VDD.n10 0.0197073
R965 VDD.n236 VDD.n223 0.0194041
R966 VDD VDD.n238 0.0192629
R967 VDD.n43 VDD 0.0155968
R968 VDD.n243 VDD 0.0147732
R969 VDD.n240 VDD.n239 0.0147268
R970 VDD.n237 VDD 0.0138562
R971 VDD VDD.n225 0.0127264
R972 VDD.n455 VDD 0.0120325
R973 VDD.n175 VDD.n169 0.0119894
R974 VDD.n454 VDD.n243 0.0112532
R975 VDD.n55 VDD 0.00907143
R976 VDD.n15 VDD 0.00708537
R977 VDD.n34 VDD.n26 0.0068871
R978 VDD.n32 VDD 0.00653659
R979 VDD.n429 VDD 0.00543671
R980 VDD.n433 VDD 0.00514516
R981 VDD VDD.n209 0.00514516
R982 VDD VDD.n456 0.00501948
R983 VDD VDD.n224 0.00368293
R984 VDD.n430 VDD 0.00315823
R985 VDD.n418 VDD 0.00282258
R986 VDD.n151 VDD 0.00282258
R987 VDD.n45 VDD 0.00224194
R988 VDD.n37 VDD 0.00224194
R989 VDD.n48 VDD 0.00224194
R990 VDD.n77 VDD 0.00224194
R991 VDD.n80 VDD 0.00224194
R992 VDD.n114 VDD 0.00224194
R993 VDD.n117 VDD 0.00224194
R994 VDD.n126 VDD 0.00224194
R995 VDD VDD.n123 0.00224194
R996 VDD VDD.n120 0.00224194
R997 VDD.n500 VDD 0.00224194
R998 VDD.n503 VDD 0.00224194
R999 VDD.n474 VDD 0.00224194
R1000 VDD.n478 VDD 0.00224194
R1001 VDD.n506 VDD 0.00224194
R1002 VDD.n190 VDD 0.00224194
R1003 VDD.n193 VDD 0.00224194
R1004 VDD.n154 VDD 0.00224194
R1005 VDD.n159 VDD 0.00224194
R1006 VDD VDD.n518 0.00224194
R1007 VDD.n137 VDD 0.00215644
R1008 VDD VDD.n463 0.00215644
R1009 VDD.n146 VDD 0.00178834
R1010 VDD VDD.n459 0.00178834
R1011 VDD.n394 VDD 0.00166129
R1012 VDD.n391 VDD 0.00166129
R1013 VDD VDD.n388 0.00166129
R1014 VDD VDD.n385 0.00166129
R1015 VDD.n326 VDD 0.00166129
R1016 VDD.n323 VDD 0.00166129
R1017 VDD VDD.n320 0.00166129
R1018 VDD VDD.n317 0.00166129
R1019 VDD.n298 VDD 0.00166129
R1020 VDD.n295 VDD 0.00166129
R1021 VDD VDD.n292 0.00166129
R1022 VDD VDD.n289 0.00166129
R1023 VDD.n270 VDD 0.00166129
R1024 VDD.n267 VDD 0.00166129
R1025 VDD VDD.n264 0.00166129
R1026 VDD VDD.n261 0.00166129
R1027 VDD.n447 VDD 0.00151695
R1028 VDD.n444 VDD 0.00151695
R1029 VDD.n441 VDD 0.00151695
R1030 VDD VDD.n438 0.00151695
R1031 VDD VDD.n347 0.00151695
R1032 VDD.n351 VDD 0.00151695
R1033 VDD VDD.n354 0.00151695
R1034 VDD.n357 VDD 0.00151695
R1035 VDD.n364 VDD 0.00150559
R1036 VDD VDD.n367 0.00150559
R1037 VDD.n371 VDD 0.00150559
R1038 VDD VDD.n452 0.00150559
R1039 VDD VDD.n330 0.00149448
R1040 VDD.n334 VDD 0.00149448
R1041 VDD VDD.n337 0.00149448
R1042 VDD.n340 VDD 0.00149448
R1043 VDD VDD.n236 0.00132192
R1044 VDD.n34 VDD 0.00108064
R1045 VDD.n68 VDD 0.00108064
R1046 VDD VDD.n71 0.00108064
R1047 VDD.n105 VDD 0.00108064
R1048 VDD VDD.n108 0.00108064
R1049 VDD.n491 VDD 0.00108064
R1050 VDD VDD.n494 0.00108064
R1051 VDD.n418 VDD 0.00108064
R1052 VDD.n181 VDD 0.00108064
R1053 VDD VDD.n184 0.00108064
R1054 VDD.n85 VDD 0.00107692
R1055 VDD.n468 VDD 0.00107692
R1056 VDD.n12 VDD 0.00104878
R1057 VDD.n227 VDD 0.00100943
R1058 VDD VDD.n142 0.000868098
R1059 VDD VDD.n461 0.000868098
R1060 VDD.n231 VDD 0.000719512
R1061 VDD.n239 VDD 0.000706186
R1062 VDD VDD.n234 0.000705479
R1063 VDD VDD.n242 0.000669492
R1064 VSS.n374 VSS.n373 76606.4
R1065 VSS.n375 VSS.n374 44973
R1066 VSS.n253 VSS.n252 19895.3
R1067 VSS.n244 VSS.t309 17230
R1068 VSS.n354 VSS.n353 16982.4
R1069 VSS.n2 VSS.n1 14181.9
R1070 VSS.n174 VSS.t304 10467.5
R1071 VSS.n353 VSS.t38 9497.33
R1072 VSS.n425 VSS.n19 9415.54
R1073 VSS.n18 VSS.t210 7006.49
R1074 VSS.n260 VSS.n172 6768.84
R1075 VSS.n260 VSS.n171 5510.82
R1076 VSS.n1 VSS.n0 4665.4
R1077 VSS.n92 VSS.t73 4499.58
R1078 VSS.n373 VSS.n372 4367.83
R1079 VSS.n373 VSS.n371 3873.69
R1080 VSS.n3 VSS.n2 3525.32
R1081 VSS.n171 VSS.n169 3387.22
R1082 VSS.n254 VSS.n253 2682.86
R1083 VSS.t263 VSS.n334 2673.11
R1084 VSS.t164 VSS.n260 2644.14
R1085 VSS.n180 VSS.n174 2588.5
R1086 VSS.n171 VSS.n170 2553.84
R1087 VSS.t188 VSS.t173 2307.56
R1088 VSS.t299 VSS.t162 2307.56
R1089 VSS.t319 VSS.t270 2307.56
R1090 VSS.t20 VSS.t187 2307.56
R1091 VSS.t54 VSS.t307 2307.56
R1092 VSS.t229 VSS.t216 2307.56
R1093 VSS.t335 VSS.t116 2307.56
R1094 VSS.t239 VSS.t169 2307.56
R1095 VSS.t114 VSS.t321 2307.56
R1096 VSS.t129 VSS.t176 2307.56
R1097 VSS.t141 VSS.t119 2307.56
R1098 VSS.t76 VSS.t121 2307.56
R1099 VSS.t59 VSS.t63 2307.56
R1100 VSS.t137 VSS.t294 2307.56
R1101 VSS.t43 VSS.t195 2307.56
R1102 VSS.t264 VSS.t134 2307.56
R1103 VSS.t204 VSS.t225 2307.56
R1104 VSS.n333 VSS.n145 2212.13
R1105 VSS.n180 VSS.t284 2166.67
R1106 VSS.n260 VSS.n259 2165.66
R1107 VSS.n349 VSS.n74 2098.2
R1108 VSS.n427 VSS.n426 2091.23
R1109 VSS.t79 VSS.n295 2068.97
R1110 VSS.n226 VSS.t240 2050.53
R1111 VSS.n425 VSS.t253 1731.96
R1112 VSS.t75 VSS.n344 1719.24
R1113 VSS.n191 VSS.t130 1635.55
R1114 VSS.n344 VSS.n343 1565.03
R1115 VSS.n334 VSS.n333 1565.03
R1116 VSS.n289 VSS.t241 1564.96
R1117 VSS.n105 VSS.t286 1272.1
R1118 VSS.n426 VSS.n425 1249.34
R1119 VSS.n242 VSS.t282 1199.47
R1120 VSS.n209 VSS.t181 1199.47
R1121 VSS.t332 VSS.n17 1199.47
R1122 VSS.n349 VSS.t158 1199.47
R1123 VSS.n241 VSS.t292 1153.78
R1124 VSS.t120 VSS.n92 1153.78
R1125 VSS.n371 VSS.n370 1145.32
R1126 VSS.n258 VSS.t325 1143.48
R1127 VSS.n196 VSS.n195 1139.06
R1128 VSS.n161 VSS.t191 1134.57
R1129 VSS.n228 VSS.n227 1119.51
R1130 VSS.t218 VSS.n331 1108.08
R1131 VSS.n227 VSS.n203 1076.69
R1132 VSS.n333 VSS.n332 1073.81
R1133 VSS.t81 VSS.t172 1058.09
R1134 VSS.n290 VSS.n289 988.177
R1135 VSS.n3 VSS.t100 927.716
R1136 VSS.t302 VSS.t293 913.885
R1137 VSS.t301 VSS.t239 913.885
R1138 VSS.t37 VSS.t76 913.885
R1139 VSS.t41 VSS.t264 913.885
R1140 VSS.n51 VSS.t117 836.591
R1141 VSS.t67 VSS.t124 794.981
R1142 VSS.n174 VSS.n19 791.109
R1143 VSS.t309 VSS.n243 730.073
R1144 VSS.n74 VSS.n7 686.213
R1145 VSS.n291 VSS.t275 663.793
R1146 VSS.t193 VSS.n290 596.024
R1147 VSS.n259 VSS.t276 595.653
R1148 VSS.t166 VSS.n196 578.554
R1149 VSS.t185 VSS.n118 573.788
R1150 VSS.t292 VSS.n240 548.331
R1151 VSS.n198 VSS.t340 548.331
R1152 VSS.n199 VSS.t188 548.331
R1153 VSS.n200 VSS.t302 548.331
R1154 VSS.t253 VSS.n424 548.331
R1155 VSS.t270 VSS.n423 548.331
R1156 VSS.t187 VSS.n422 548.331
R1157 VSS.n23 VSS.t308 548.331
R1158 VSS.t240 VSS.n225 548.331
R1159 VSS.t216 VSS.n224 548.331
R1160 VSS.t116 VSS.n223 548.331
R1161 VSS.n208 VSS.t301 548.331
R1162 VSS.n93 VSS.t120 548.331
R1163 VSS.n98 VSS.t321 548.331
R1164 VSS.n99 VSS.t129 548.331
R1165 VSS.n102 VSS.t34 548.331
R1166 VSS.n348 VSS.t37 548.331
R1167 VSS.n347 VSS.t59 548.331
R1168 VSS.n346 VSS.t137 548.331
R1169 VSS.n345 VSS.t75 548.331
R1170 VSS.n341 VSS.t41 548.331
R1171 VSS.n340 VSS.t204 548.331
R1172 VSS.n339 VSS.t27 548.331
R1173 VSS.n335 VSS.t263 548.331
R1174 VSS.n331 VSS.n302 531.466
R1175 VSS.t183 VSS.t132 518.688
R1176 VSS.n211 VSS.t327 503.682
R1177 VSS.t201 VSS.n28 466.476
R1178 VSS.n227 VSS.n226 453.219
R1179 VSS.t102 VSS.t46 434.212
R1180 VSS.t149 VSS.t205 434.212
R1181 VSS.n426 VSS.n17 426.769
R1182 VSS.n265 VSS.t145 426.396
R1183 VSS.n253 VSS.t167 396.058
R1184 VSS.n240 VSS.t267 365.555
R1185 VSS.t173 VSS.n198 365.555
R1186 VSS.n199 VSS.t231 365.555
R1187 VSS.t162 VSS.n200 365.555
R1188 VSS.n424 VSS.t319 365.555
R1189 VSS.n423 VSS.t20 365.555
R1190 VSS.n422 VSS.t54 365.555
R1191 VSS.t282 VSS.n23 365.555
R1192 VSS.n225 VSS.t229 365.555
R1193 VSS.n224 VSS.t335 365.555
R1194 VSS.t181 VSS.n208 365.555
R1195 VSS.n93 VSS.t114 365.555
R1196 VSS.t176 VSS.n98 365.555
R1197 VSS.n99 VSS.t141 365.555
R1198 VSS.n102 VSS.t332 365.555
R1199 VSS.t158 VSS.n348 365.555
R1200 VSS.t121 VSS.n347 365.555
R1201 VSS.t63 VSS.n346 365.555
R1202 VSS.t294 VSS.n345 365.555
R1203 VSS.t195 VSS.n341 365.555
R1204 VSS.t134 VSS.n340 365.555
R1205 VSS.t225 VSS.n339 365.555
R1206 VSS.n335 VSS.t313 365.555
R1207 VSS.t175 VSS.t238 350.877
R1208 VSS.t274 VSS.t334 350.404
R1209 VSS.t215 VSS.t161 350.404
R1210 VSS.t171 VSS.t212 350.404
R1211 VSS.t42 VSS.t70 350.404
R1212 VSS.t298 VSS.t87 350.404
R1213 VSS.t273 VSS.t228 350.404
R1214 VSS.n196 VSS.n174 345.394
R1215 VSS.t178 VSS.n7 331.695
R1216 VSS.t84 VSS.t248 329.029
R1217 VSS.t12 VSS.t260 327.675
R1218 VSS.t28 VSS.t23 327.675
R1219 VSS.t0 VSS.n148 319.466
R1220 VSS.t66 VSS.n16 316.639
R1221 VSS.n428 VSS.n427 311.87
R1222 VSS.t60 VSS.t147 311.825
R1223 VSS.t288 VSS.t198 311.825
R1224 VSS.n118 VSS.t22 310.985
R1225 VSS.n19 VSS.n18 297.363
R1226 VSS.n175 VSS.t337 281.091
R1227 VSS.n360 VSS.n354 272.553
R1228 VSS.n375 VSS.n73 270.834
R1229 VSS.n288 VSS.t254 269.688
R1230 VSS.n164 VSS.t209 255.748
R1231 VSS.n376 VSS.n375 251.548
R1232 VSS.n370 VSS.n369 251.548
R1233 VSS.t259 VSS.n428 249.042
R1234 VSS.t38 VSS.n352 235.839
R1235 VSS.t108 VSS.t71 223.987
R1236 VSS.t330 VSS.t48 223.987
R1237 VSS.t278 VSS.t26 214.912
R1238 VSS.t339 VSS.t95 214.912
R1239 VSS.n11 VSS.t60 210.811
R1240 VSS.n430 VSS.t288 210.811
R1241 VSS.t26 VSS.n29 210.526
R1242 VSS.n30 VSS.t278 210.526
R1243 VSS.t95 VSS.n32 210.526
R1244 VSS.n33 VSS.t339 210.526
R1245 VSS.t238 VSS.n35 210.526
R1246 VSS.n37 VSS.t15 210.526
R1247 VSS.n38 VSS.t297 210.526
R1248 VSS.n52 VSS.t274 210.244
R1249 VSS.t161 VSS.n53 210.244
R1250 VSS.n214 VSS.t171 210.244
R1251 VSS.t138 VSS.n111 210.244
R1252 VSS.n112 VSS.t83 210.244
R1253 VSS.t224 VSS.n117 210.244
R1254 VSS.n119 VSS.t269 210.244
R1255 VSS.n123 VSS.t258 210.244
R1256 VSS.n124 VSS.t42 210.244
R1257 VSS.n126 VSS.t298 210.244
R1258 VSS.n127 VSS.t273 210.244
R1259 VSS.n202 VSS.t31 206.125
R1260 VSS.t311 VSS.t257 198.954
R1261 VSS.t241 VSS.n288 192.633
R1262 VSS.n280 VSS.t84 191.375
R1263 VSS.n72 VSS.t12 190.587
R1264 VSS.n360 VSS.t28 190.587
R1265 VSS.n251 VSS.t144 186.381
R1266 VSS.n429 VSS.t259 185.786
R1267 VSS.t316 VSS.t214 183.456
R1268 VSS.n149 VSS.t16 180.292
R1269 VSS.t172 VSS.n245 176.673
R1270 VSS.t105 VSS.t271 175.202
R1271 VSS.t179 VSS.t289 175.202
R1272 VSS.n375 VSS.t152 174.407
R1273 VSS.n370 VSS.t96 174.407
R1274 VSS.t19 VSS.n40 170.585
R1275 VSS.n296 VSS.t85 163.793
R1276 VSS.n44 VSS.n43 159.873
R1277 VSS.n47 VSS.n46 159.873
R1278 VSS.n145 VSS.t175 157.895
R1279 VSS.n153 VSS.t316 151.768
R1280 VSS.t31 VSS.n201 145.708
R1281 VSS.t71 VSS.n9 140.542
R1282 VSS.n11 VSS.t108 140.542
R1283 VSS.n430 VSS.t330 140.542
R1284 VSS.t48 VSS.n429 140.542
R1285 VSS.n30 VSS.t233 140.351
R1286 VSS.n32 VSS.t155 140.351
R1287 VSS.n33 VSS.t189 140.351
R1288 VSS.t46 VSS.n35 140.351
R1289 VSS.n37 VSS.t102 140.351
R1290 VSS.t205 VSS.n38 140.351
R1291 VSS.n29 VSS.t201 140.185
R1292 VSS.t271 VSS.n52 140.162
R1293 VSS.n53 VSS.t105 140.162
R1294 VSS.n214 VSS.t179 140.162
R1295 VSS.t289 VSS.n55 140.162
R1296 VSS.n111 VSS.t56 140.162
R1297 VSS.n112 VSS.t199 140.162
R1298 VSS.n117 VSS.t8 140.162
R1299 VSS.n119 VSS.t185 140.162
R1300 VSS.n302 VSS.t88 139.192
R1301 VSS.n245 VSS.t144 133.962
R1302 VSS.n301 VSS.t207 126.061
R1303 VSS.n246 VSS.t81 124.254
R1304 VSS.t167 VSS.n251 124.254
R1305 VSS.n343 VSS.n342 114.236
R1306 VSS.n40 VSS.t149 110.543
R1307 VSS.n331 VSS.n327 106.921
R1308 VSS.n148 VSS.t303 103.255
R1309 VSS.t16 VSS.n59 101.218
R1310 VSS.t15 VSS.t279 100.877
R1311 VSS.t297 VSS.t247 100.877
R1312 VSS.n244 VSS.t166 99.0148
R1313 VSS.t145 VSS.t98 94.0088
R1314 VSS.t152 VSS.t235 93.9117
R1315 VSS.t96 VSS.t51 93.9117
R1316 VSS.t132 VSS.n153 91.9197
R1317 VSS.t208 VSS.t250 89.7916
R1318 VSS.t124 VSS.t243 89.7916
R1319 VSS.t217 VSS.t67 89.7916
R1320 VSS.t117 VSS.t94 89.7916
R1321 VSS.t139 VSS.t111 87.6016
R1322 VSS.t280 VSS.t5 87.6016
R1323 VSS.n246 VSS.n244 87.3661
R1324 VSS.t88 VSS.n301 84.0409
R1325 VSS.n202 VSS.t19 78.1853
R1326 VSS.n289 VSS.n167 77.2216
R1327 VSS.t2 VSS.t221 58.5375
R1328 VSS.n210 VSS.n57 56.6646
R1329 VSS.n416 VSS.n25 54.1355
R1330 VSS.t111 VSS.n123 52.5611
R1331 VSS.n124 VSS.t139 52.5611
R1332 VSS.t5 VSS.n126 52.5611
R1333 VSS.n127 VSS.t280 52.5611
R1334 VSS.n43 VSS.t208 50.3711
R1335 VSS.t243 VSS.n44 50.3711
R1336 VSS.n46 VSS.t217 50.3711
R1337 VSS.t94 VSS.n47 50.3711
R1338 VSS.t334 VSS.n51 48.1811
R1339 VSS.n254 VSS.t325 47.8266
R1340 VSS.t276 VSS.n258 47.8266
R1341 VSS.t257 VSS.n209 45.3318
R1342 VSS.n105 VSS.n17 41.0359
R1343 VSS.n428 VSS.t66 35.5779
R1344 VSS.n342 VSS.t43 34.2711
R1345 VSS.n332 VSS.t218 34.2711
R1346 VSS.t73 VSS.t178 33.4743
R1347 VSS.n235 VSS.n41 27.068
R1348 VSS.t327 VSS.n210 23.9253
R1349 VSS.n243 VSS.n242 23.5512
R1350 VSS.n202 VSS.t299 22.8476
R1351 VSS.n330 VSS.t11 20.9066
R1352 VSS.t209 VSS.t143 20.1154
R1353 VSS.t85 VSS.t79 20.1154
R1354 VSS.n291 VSS.t193 17.2419
R1355 VSS.n73 VSS.n72 16.7186
R1356 VSS.n261 VSS.t164 16.5119
R1357 VSS.n370 VSS.n354 14.7536
R1358 VSS.n217 VSS.n160 13.2511
R1359 VSS.t11 VSS.t2 13.1415
R1360 VSS.n228 VSS.n202 11.424
R1361 VSS.n155 VSS.t184 10.2623
R1362 VSS.n149 VSS.t0 9.48955
R1363 VSS.n242 VSS.n241 9.42079
R1364 VSS.n257 VSS.t277 9.40866
R1365 VSS.n106 VSS.t287 9.3736
R1366 VSS.n212 VSS.t312 9.3736
R1367 VSS.n197 VSS.t310 9.3736
R1368 VSS.n229 VSS.t300 9.3736
R1369 VSS.n147 VSS.n146 9.37275
R1370 VSS.n329 VSS.n328 9.37275
R1371 VSS.n88 VSS.n87 9.37275
R1372 VSS.n351 VSS.n350 9.37275
R1373 VSS.n284 VSS.t99 9.3645
R1374 VSS.n279 VSS.n266 9.3221
R1375 VSS.n272 VSS.t146 9.3221
R1376 VSS.n264 VSS.n168 9.3221
R1377 VSS.n286 VSS.t242 9.3221
R1378 VSS.n66 VSS.t213 9.3221
R1379 VSS.n68 VSS.n65 9.3221
R1380 VSS.n366 VSS.t97 9.3221
R1381 VSS.n364 VSS.n356 9.3221
R1382 VSS.n293 VSS.t194 9.30652
R1383 VSS.n163 VSS.t192 9.30652
R1384 VSS.n282 VSS.t249 9.30652
R1385 VSS.n263 VSS.t165 9.30652
R1386 VSS.n190 VSS.t244 9.30652
R1387 VSS.n173 VSS.t131 9.30652
R1388 VSS.n61 VSS.n60 9.30652
R1389 VSS.n70 VSS.n62 9.30652
R1390 VSS.n362 VSS.n359 9.30652
R1391 VSS.n367 VSS.n355 9.30652
R1392 VSS.n5 VSS.t101 9.30652
R1393 VSS.n188 VSS.t62 9.30518
R1394 VSS.n193 VSS.t338 9.30518
R1395 VSS.n182 VSS.t285 9.30323
R1396 VSS.n151 VSS.t1 9.30204
R1397 VSS.n256 VSS.t326 9.29981
R1398 VSS.n158 VSS.n152 9.29009
R1399 VSS.n156 VSS.t133 9.29009
R1400 VSS.t212 VSS.t215 8.76061
R1401 VSS.n154 VSS.t183 7.87929
R1402 VSS.n275 VSS.n274 7.39136
R1403 VSS VSS.n357 7.30633
R1404 VSS VSS.n63 7.30633
R1405 VSS.n391 VSS.n45 7.19156
R1406 VSS.n395 VSS.n42 7.19156
R1407 VSS.n379 VSS.n58 7.19156
R1408 VSS.n381 VSS.n56 7.19156
R1409 VSS.n313 VSS.n312 7.19156
R1410 VSS.n310 VSS.n309 7.19156
R1411 VSS.n307 VSS.n306 7.19156
R1412 VSS.n325 VSS.n324 7.19156
R1413 VSS.n322 VSS.n321 7.19156
R1414 VSS.n319 VSS.n318 7.19156
R1415 VSS.n271 VSS.t148 7.19156
R1416 VSS.n411 VSS.n31 7.19156
R1417 VSS.n414 VSS.n27 7.19156
R1418 VSS.n337 VSS.n144 7.19156
R1419 VSS.n143 VSS.n142 7.19156
R1420 VSS.n140 VSS.n139 7.19156
R1421 VSS.n115 VSS.n90 7.19156
R1422 VSS.n109 VSS.n91 7.19156
R1423 VSS.n85 VSS.n84 7.19156
R1424 VSS.n82 VSS.n81 7.19156
R1425 VSS.n79 VSS.n78 7.19156
R1426 VSS.n114 VSS.t200 7.17323
R1427 VSS.n121 VSS.t186 7.17323
R1428 VSS.n392 VSS.t125 7.17323
R1429 VSS.n388 VSS.t118 7.17323
R1430 VSS.n248 VSS.t82 7.17156
R1431 VSS.n410 VSS.t234 7.16989
R1432 VSS.n406 VSS.t190 7.16989
R1433 VSS.n439 VSS.t74 7.16656
R1434 VSS.n437 VSS.t128 7.16656
R1435 VSS.n298 VSS.t80 7.16085
R1436 VSS.n299 VSS.t89 7.15156
R1437 VSS.n21 VSS.t320 7.13489
R1438 VSS.n24 VSS.t21 7.13489
R1439 VSS.n420 VSS.t55 7.13489
R1440 VSS.n205 VSS.t230 7.13323
R1441 VSS.n207 VSS.t336 7.13323
R1442 VSS.n221 VSS.t170 7.13323
R1443 VSS.n238 VSS.t268 7.13156
R1444 VSS.n236 VSS.t174 7.13156
R1445 VSS.n233 VSS.t232 7.13156
R1446 VSS.n184 VSS.n183 7.1285
R1447 VSS.n95 VSS.t115 7.12823
R1448 VSS.n96 VSS.t177 7.12823
R1449 VSS.n101 VSS.t142 7.12823
R1450 VSS.n299 VSS.n298 6.41993
R1451 VSS.n352 VSS.n349 6.08664
R1452 VSS VSS.t86 6.02876
R1453 VSS.n178 VSS.n177 6.01414
R1454 VSS.n178 VSS.t211 6.01414
R1455 VSS.n398 VSS.n39 5.91399
R1456 VSS.n402 VSS.n36 5.91399
R1457 VSS.n383 VSS.n54 5.91399
R1458 VSS.n385 VSS.n50 5.91399
R1459 VSS.n304 VSS.n303 5.91399
R1460 VSS.n316 VSS.n315 5.91399
R1461 VSS.n130 VSS.n125 5.91399
R1462 VSS.n134 VSS.n122 5.91399
R1463 VSS.n137 VSS.n89 5.91399
R1464 VSS.n13 VSS.n12 5.91399
R1465 VSS.n434 VSS.n10 5.91399
R1466 VSS.n76 VSS.n75 5.91399
R1467 VSS.n249 VSS.t168 5.89898
R1468 VSS.n131 VSS.t140 5.89565
R1469 VSS.n26 VSS.t281 5.89565
R1470 VSS.n213 VSS.t272 5.89565
R1471 VSS.n216 VSS.t180 5.89565
R1472 VSS.n403 VSS.t47 5.89232
R1473 VSS.n399 VSS.t206 5.89232
R1474 VSS.n433 VSS.t72 5.88898
R1475 VSS.n14 VSS.t331 5.88898
R1476 VSS.n418 VSS.t283 5.85732
R1477 VSS.n219 VSS.t182 5.85565
R1478 VSS.n231 VSS.t163 5.85398
R1479 VSS.n104 VSS.t333 5.85065
R1480 VSS VSS.n154 5.20234
R1481 VSS VSS.n228 5.20137
R1482 VSS.n150 VSS.n149 5.2005
R1483 VSS.n157 VSS.n153 5.2005
R1484 VSS.n292 VSS.n291 5.2005
R1485 VSS.n165 VSS.n164 5.2005
R1486 VSS.n297 VSS.n296 5.2005
R1487 VSS.n301 VSS.n300 5.2005
R1488 VSS.n212 VSS.n211 5.2005
R1489 VSS.n162 VSS.n161 5.2005
R1490 VSS.n269 VSS.n268 5.2005
R1491 VSS.n281 VSS.n280 5.2005
R1492 VSS.n285 VSS.n265 5.2005
R1493 VSS.n262 VSS.n261 5.2005
R1494 VSS.n288 VSS.n287 5.2005
R1495 VSS.n240 VSS.n239 5.2005
R1496 VSS.n237 VSS.n198 5.2005
R1497 VSS.n234 VSS.n199 5.2005
R1498 VSS.n232 VSS.n200 5.2005
R1499 VSS.n192 VSS.n191 5.2005
R1500 VSS.n251 VSS.n250 5.2005
R1501 VSS.n247 VSS.n246 5.2005
R1502 VSS.n243 VSS.n197 5.2005
R1503 VSS.n424 VSS.n20 5.2005
R1504 VSS.n423 VSS.n22 5.2005
R1505 VSS.n422 VSS.n421 5.2005
R1506 VSS.n419 VSS.n23 5.2005
R1507 VSS.n195 VSS.n194 5.2005
R1508 VSS.n186 VSS.n185 5.2005
R1509 VSS.n189 VSS.n175 5.2005
R1510 VSS.n258 VSS.n257 5.2005
R1511 VSS.n255 VSS.n254 5.2005
R1512 VSS.n225 VSS.n204 5.2005
R1513 VSS.n224 VSS.n206 5.2005
R1514 VSS.n223 VSS.n222 5.2005
R1515 VSS.n220 VSS.n208 5.2005
R1516 VSS.n215 VSS.n214 5.2005
R1517 VSS.n52 VSS.n48 5.2005
R1518 VSS.n327 VSS.n326 5.2005
R1519 VSS.n327 VSS.n323 5.2005
R1520 VSS.n327 VSS.n320 5.2005
R1521 VSS.n327 VSS.n317 5.2005
R1522 VSS.n327 VSS.n314 5.2005
R1523 VSS.n327 VSS.n311 5.2005
R1524 VSS.n327 VSS.n308 5.2005
R1525 VSS.n327 VSS.n305 5.2005
R1526 VSS.n330 VSS.n329 5.2005
R1527 VSS.n378 VSS.n59 5.2005
R1528 VSS.n380 VSS.n57 5.2005
R1529 VSS.n382 VSS.n55 5.2005
R1530 VSS.n384 VSS.n53 5.2005
R1531 VSS.n72 VSS.n71 5.2005
R1532 VSS.n377 VSS.n376 5.2005
R1533 VSS.n361 VSS.n360 5.2005
R1534 VSS.n369 VSS.n368 5.2005
R1535 VSS.n389 VSS.n47 5.2005
R1536 VSS.n393 VSS.n44 5.2005
R1537 VSS.n412 VSS.n30 5.2005
R1538 VSS.n408 VSS.n33 5.2005
R1539 VSS.n404 VSS.n35 5.2005
R1540 VSS.n400 VSS.n38 5.2005
R1541 VSS.n390 VSS.n46 5.2005
R1542 VSS.n394 VSS.n43 5.2005
R1543 VSS.n397 VSS.n40 5.2005
R1544 VSS.n401 VSS.n37 5.2005
R1545 VSS.n409 VSS.n32 5.2005
R1546 VSS.n413 VSS.n29 5.2005
R1547 VSS.n431 VSS.n430 5.2005
R1548 VSS.n435 VSS.n9 5.2005
R1549 VSS.n429 VSS.n15 5.2005
R1550 VSS.n432 VSS.n11 5.2005
R1551 VSS.n106 VSS.n105 5.2005
R1552 VSS.n94 VSS.n93 5.2005
R1553 VSS.n98 VSS.n97 5.2005
R1554 VSS.n100 VSS.n99 5.2005
R1555 VSS.n103 VSS.n102 5.2005
R1556 VSS.n352 VSS.n351 5.2005
R1557 VSS.n332 VSS.n147 5.2005
R1558 VSS.n336 VSS.n335 5.2005
R1559 VSS.n339 VSS.n338 5.2005
R1560 VSS.n340 VSS.n141 5.2005
R1561 VSS.n341 VSS.n138 5.2005
R1562 VSS.n342 VSS.n88 5.2005
R1563 VSS.n345 VSS.n86 5.2005
R1564 VSS.n346 VSS.n83 5.2005
R1565 VSS.n347 VSS.n80 5.2005
R1566 VSS.n348 VSS.n77 5.2005
R1567 VSS.n129 VSS.n126 5.2005
R1568 VSS.n133 VSS.n123 5.2005
R1569 VSS.n120 VSS.n119 5.2005
R1570 VSS.n113 VSS.n112 5.2005
R1571 VSS.n128 VSS.n127 5.2005
R1572 VSS.n132 VSS.n124 5.2005
R1573 VSS.n117 VSS.n116 5.2005
R1574 VSS.n111 VSS.n110 5.2005
R1575 VSS.n4 VSS.n3 5.2005
R1576 VSS.n181 VSS.n180 5.2005
R1577 VSS.n438 VSS.n7 5.2005
R1578 VSS.n440 VSS.n7 5.2005
R1579 VSS.n211 VSS.t322 5.03731
R1580 VSS.n274 VSS.n273 4.5005
R1581 VSS.n273 VSS 4.12455
R1582 VSS.t337 VSS.t61 3.67489
R1583 VSS.n195 VSS.n175 3.67489
R1584 VSS.n179 VSS.n178 3.28959
R1585 VSS.n185 VSS.n184 3.03722
R1586 VSS.n277 VSS.n276 2.6005
R1587 VSS.n276 VSS.n167 2.6005
R1588 VSS.t322 VSS.t311 2.5189
R1589 VSS.n331 VSS.n330 2.38977
R1590 VSS.n407 VSS 2.24014
R1591 VSS.t83 VSS.t138 2.19053
R1592 VSS.t269 VSS.t224 2.19053
R1593 VSS.n183 VSS.n182 2.13762
R1594 VSS VSS.n6 1.98772
R1595 VSS.n286 VSS 1.09141
R1596 VSS.n184 VSS.n175 1.00481
R1597 VSS.n405 VSS.n34 0.846463
R1598 VSS.n386 VSS.n49 0.846463
R1599 VSS.n136 VSS.n135 0.846463
R1600 VSS.n436 VSS.n8 0.846463
R1601 VSS.n108 VSS.n107 0.843955
R1602 VSS.n300 VSS.n160 0.734346
R1603 VSS.n416 VSS.n415 0.70444
R1604 VSS.n193 VSS 0.676801
R1605 VSS.n218 VSS.n217 0.623774
R1606 VSS.n6 VSS.n5 0.616742
R1607 VSS.n396 VSS.n41 0.574895
R1608 VSS.n185 VSS.n176 0.486611
R1609 VSS.n250 VSS.n248 0.439554
R1610 VSS.n275 VSS.n270 0.365463
R1611 VSS.n310 VSS 0.343161
R1612 VSS.n313 VSS 0.343161
R1613 VSS.n322 VSS 0.343161
R1614 VSS.n325 VSS 0.343161
R1615 VSS.n143 VSS 0.343161
R1616 VSS VSS.n337 0.343161
R1617 VSS.n82 VSS 0.343161
R1618 VSS.n85 VSS 0.343161
R1619 VSS.n166 VSS.n163 0.338437
R1620 VSS.n247 VSS.n173 0.316175
R1621 VSS.n249 VSS 0.311851
R1622 VSS.n69 VSS.n68 0.310174
R1623 VSS.n364 VSS.n363 0.310174
R1624 VSS VSS.n305 0.289491
R1625 VSS VSS.n317 0.289491
R1626 VSS VSS.n138 0.289491
R1627 VSS VSS.n77 0.289491
R1628 VSS.n156 VSS.n155 0.284276
R1629 VSS.n297 VSS.n294 0.277931
R1630 VSS.n166 VSS.n165 0.272151
R1631 VSS VSS.n21 0.265394
R1632 VSS.n238 VSS 0.265394
R1633 VSS VSS.n205 0.259875
R1634 VSS VSS.n207 0.259875
R1635 VSS VSS.n95 0.254582
R1636 VSS.n96 VSS 0.254582
R1637 VSS.n363 VSS.n358 0.254245
R1638 VSS.n69 VSS.n64 0.254245
R1639 VSS.n217 VSS.n216 0.241304
R1640 VSS VSS.n419 0.223904
R1641 VSS VSS.n232 0.223904
R1642 VSS VSS.n256 0.223676
R1643 VSS VSS.n220 0.21925
R1644 VSS.n103 VSS 0.214786
R1645 VSS.n387 VSS.n48 0.203
R1646 VSS.n384 VSS.n383 0.202392
R1647 VSS.n382 VSS.n381 0.202392
R1648 VSS.n159 VSS.n151 0.19152
R1649 VSS.n307 VSS 0.191234
R1650 VSS.n319 VSS 0.191234
R1651 VSS.n140 VSS 0.191234
R1652 VSS.n79 VSS 0.191234
R1653 VSS.n283 VSS.n282 0.187704
R1654 VSS.n264 VSS.n263 0.184546
R1655 VSS VSS.n188 0.182492
R1656 VSS.n179 VSS.n6 0.180913
R1657 VSS.n66 VSS.n61 0.168072
R1658 VSS.n367 VSS.n366 0.168072
R1659 VSS.n158 VSS.n157 0.165806
R1660 VSS.n298 VSS 0.158206
R1661 VSS.n215 VSS.n213 0.156125
R1662 VSS.n420 VSS 0.147947
R1663 VSS.n233 VSS 0.147947
R1664 VSS.n221 VSS 0.144875
R1665 VSS VSS.n379 0.144708
R1666 VSS.n70 VSS.n69 0.142796
R1667 VSS.n363 VSS.n362 0.142796
R1668 VSS VSS.n101 0.141929
R1669 VSS VSS.n156 0.140092
R1670 VSS.n67 VSS.n66 0.137391
R1671 VSS.n366 VSS.n365 0.137391
R1672 VSS VSS.n34 0.137136
R1673 VSS VSS.n49 0.137136
R1674 VSS.n136 VSS 0.137136
R1675 VSS VSS.n8 0.137136
R1676 VSS.n287 VSS.n264 0.136634
R1677 VSS.n25 VSS.n24 0.133266
R1678 VSS.n236 VSS.n235 0.133266
R1679 VSS.n25 VSS 0.132628
R1680 VSS.n235 VSS 0.132628
R1681 VSS.n218 VSS 0.127807
R1682 VSS.n107 VSS 0.127258
R1683 VSS.n294 VSS.n293 0.12579
R1684 VSS.n308 VSS.n307 0.118573
R1685 VSS.n311 VSS.n310 0.118573
R1686 VSS.n314 VSS.n313 0.118573
R1687 VSS.n320 VSS.n319 0.118573
R1688 VSS.n323 VSS.n322 0.118573
R1689 VSS.n326 VSS.n325 0.118573
R1690 VSS.n141 VSS.n140 0.118573
R1691 VSS.n338 VSS.n143 0.118573
R1692 VSS.n337 VSS.n336 0.118573
R1693 VSS.n80 VSS.n79 0.118573
R1694 VSS.n83 VSS.n82 0.118573
R1695 VSS.n86 VSS.n85 0.118573
R1696 VSS VSS.n286 0.115458
R1697 VSS VSS.n304 0.115271
R1698 VSS VSS.n316 0.115271
R1699 VSS VSS.n137 0.115271
R1700 VSS VSS.n76 0.115271
R1701 VSS.n68 VSS 0.114702
R1702 VSS VSS.n364 0.114702
R1703 VSS VSS.n190 0.109909
R1704 VSS.n256 VSS.n255 0.109351
R1705 VSS.n417 VSS 0.106075
R1706 VSS.n304 VSS.n34 0.10206
R1707 VSS.n316 VSS.n49 0.10206
R1708 VSS.n137 VSS.n136 0.10206
R1709 VSS.n76 VSS.n8 0.10206
R1710 VSS.n21 VSS.n20 0.0917766
R1711 VSS.n24 VSS.n22 0.0917766
R1712 VSS.n421 VSS.n420 0.0917766
R1713 VSS.n239 VSS.n238 0.0917766
R1714 VSS.n237 VSS.n236 0.0917766
R1715 VSS.n234 VSS.n233 0.0917766
R1716 VSS.n205 VSS.n204 0.089875
R1717 VSS.n207 VSS.n206 0.089875
R1718 VSS.n222 VSS.n221 0.089875
R1719 VSS.n190 VSS.n189 0.0895055
R1720 VSS VSS.n418 0.0892234
R1721 VSS VSS.n231 0.0892234
R1722 VSS.n95 VSS.n94 0.088051
R1723 VSS.n97 VSS.n96 0.088051
R1724 VSS.n101 VSS.n100 0.088051
R1725 VSS VSS.n299 0.0879825
R1726 VSS VSS.n219 0.087375
R1727 VSS.n188 VSS.n187 0.0869264
R1728 VSS.n104 VSS 0.085602
R1729 VSS.n248 VSS 0.085027
R1730 VSS VSS.n249 0.085027
R1731 VSS.n386 VSS.n385 0.0790328
R1732 VSS.n418 VSS.n417 0.0790106
R1733 VSS.n231 VSS.n230 0.0790106
R1734 VSS.n294 VSS.n166 0.0777727
R1735 VSS.n219 VSS.n218 0.077375
R1736 VSS.n181 VSS.n179 0.0760505
R1737 VSS.n107 VSS.n104 0.0758061
R1738 VSS.n406 VSS.n405 0.0730937
R1739 VSS.n151 VSS.n150 0.073051
R1740 VSS.n230 VSS.n229 0.0718942
R1741 VSS.n276 VSS.n275 0.071566
R1742 VSS.n131 VSS.n130 0.0714745
R1743 VSS.n279 VSS.n278 0.0706762
R1744 VSS.n396 VSS.n395 0.0699903
R1745 VSS.n439 VSS 0.0695388
R1746 VSS.n183 VSS 0.0691188
R1747 VSS.n293 VSS.n292 0.0675755
R1748 VSS.n163 VSS.n162 0.0675755
R1749 VSS.n282 VSS.n281 0.0675755
R1750 VSS.n263 VSS.n262 0.0675755
R1751 VSS.n192 VSS.n173 0.0675755
R1752 VSS.n5 VSS.n4 0.0675755
R1753 VSS.n432 VSS.n431 0.0671567
R1754 VSS.n71 VSS.n70 0.0667264
R1755 VSS.n362 VSS.n361 0.0667264
R1756 VSS.n213 VSS 0.0666607
R1757 VSS.n182 VSS 0.0624266
R1758 VSS.n109 VSS.n108 0.0600053
R1759 VSS.n377 VSS.n61 0.0557756
R1760 VSS.n368 VSS.n367 0.0557756
R1761 VSS.n271 VSS 0.0548172
R1762 VSS.n401 VSS.n400 0.0542031
R1763 VSS VSS.n436 0.0535035
R1764 VSS.n381 VSS.n380 0.0501911
R1765 VSS.n379 VSS.n378 0.0501911
R1766 VSS.n385 VSS 0.0488012
R1767 VSS.n383 VSS 0.0488012
R1768 VSS.n283 VSS.n279 0.0449053
R1769 VSS.n194 VSS.n193 0.04
R1770 VSS.n415 VSS.n414 0.0397654
R1771 VSS.n387 VSS.n386 0.0383764
R1772 VSS.n216 VSS 0.0377321
R1773 VSS.n276 VSS.n269 0.036033
R1774 VSS.n417 VSS.n416 0.036
R1775 VSS.n415 VSS.n26 0.0322091
R1776 VSS.n230 VSS.n41 0.0316538
R1777 VSS.n135 VSS.n134 0.0309948
R1778 VSS.n135 VSS 0.03059
R1779 VSS.n388 VSS 0.0270817
R1780 VSS.n285 VSS.n284 0.0263107
R1781 VSS.n440 VSS.n439 0.0242893
R1782 VSS.n438 VSS.n437 0.0242893
R1783 VSS.n273 VSS.n272 0.0211167
R1784 VSS VSS.n391 0.0206049
R1785 VSS.n110 VSS.n109 0.0197954
R1786 VSS.n114 VSS.n113 0.0197954
R1787 VSS.n116 VSS.n115 0.0197954
R1788 VSS.n121 VSS.n120 0.0197954
R1789 VSS.n414 VSS.n413 0.0197954
R1790 VSS.n395 VSS.n394 0.0197954
R1791 VSS.n393 VSS.n392 0.0197954
R1792 VSS.n391 VSS.n390 0.0197954
R1793 VSS.n389 VSS.n388 0.0197954
R1794 VSS.n159 VSS.n158 0.0197857
R1795 VSS.n108 VSS.n15 0.0193906
R1796 VSS.n437 VSS 0.0192985
R1797 VSS.n436 VSS.n435 0.0192556
R1798 VSS VSS.n403 0.0192556
R1799 VSS.n402 VSS 0.0192556
R1800 VSS VSS.n399 0.0192556
R1801 VSS.n398 VSS 0.0192556
R1802 VSS.n412 VSS.n411 0.0181762
R1803 VSS.n410 VSS.n409 0.0181762
R1804 VSS.n408 VSS.n407 0.0175015
R1805 VSS VSS.n387 0.0158823
R1806 VSS.n115 VSS.n114 0.0119693
R1807 VSS VSS.n434 0.0116994
R1808 VSS.n433 VSS 0.0116994
R1809 VSS.n13 VSS 0.0116994
R1810 VSS VSS.n14 0.0116994
R1811 VSS VSS.n121 0.0108898
R1812 VSS.n284 VSS.n283 0.00961702
R1813 VSS.n397 VSS.n396 0.00940555
R1814 VSS.n434 VSS.n433 0.00805622
R1815 VSS.n14 VSS.n13 0.00805622
R1816 VSS.n392 VSS 0.00805622
R1817 VSS.n134 VSS.n133 0.00792129
R1818 VSS.n132 VSS.n131 0.00792129
R1819 VSS.n130 VSS.n129 0.00792129
R1820 VSS.n128 VSS.n26 0.00792129
R1821 VSS.n272 VSS.n271 0.00644714
R1822 VSS.n405 VSS.n404 0.0063021
R1823 VSS.n403 VSS.n402 0.0058973
R1824 VSS.n399 VSS.n398 0.0058973
R1825 VSS VSS.n308 0.00545413
R1826 VSS VSS.n311 0.00545413
R1827 VSS.n314 VSS 0.00545413
R1828 VSS VSS.n320 0.00545413
R1829 VSS VSS.n323 0.00545413
R1830 VSS.n326 VSS 0.00545413
R1831 VSS VSS.n141 0.00545413
R1832 VSS.n338 VSS 0.00545413
R1833 VSS.n336 VSS 0.00545413
R1834 VSS VSS.n80 0.00545413
R1835 VSS VSS.n83 0.00545413
R1836 VSS.n86 VSS 0.00545413
R1837 VSS.n20 VSS 0.00432979
R1838 VSS.n22 VSS 0.00432979
R1839 VSS.n421 VSS 0.00432979
R1840 VSS.n239 VSS 0.00432979
R1841 VSS VSS.n237 0.00432979
R1842 VSS VSS.n234 0.00432979
R1843 VSS.n204 VSS 0.00425
R1844 VSS.n206 VSS 0.00425
R1845 VSS.n222 VSS 0.00425
R1846 VSS.n94 VSS 0.00417347
R1847 VSS.n97 VSS 0.00417347
R1848 VSS.n100 VSS 0.00417347
R1849 VSS.n157 VSS 0.00417347
R1850 VSS.n155 VSS 0.00417347
R1851 VSS.n358 VSS 0.00380275
R1852 VSS.n305 VSS 0.00380275
R1853 VSS.n317 VSS 0.00380275
R1854 VSS.n165 VSS 0.00380275
R1855 VSS VSS.n297 0.00380275
R1856 VSS.n64 VSS 0.00380275
R1857 VSS.n138 VSS 0.00380275
R1858 VSS.n77 VSS 0.00380275
R1859 VSS.n287 VSS 0.00352521
R1860 VSS VSS.n67 0.00352521
R1861 VSS.n365 VSS 0.00352521
R1862 VSS VSS.n48 0.0035
R1863 VSS.n160 VSS.n159 0.00324928
R1864 VSS.n419 VSS 0.00305319
R1865 VSS.n232 VSS 0.00305319
R1866 VSS.n300 VSS 0.00301748
R1867 VSS.n220 VSS 0.003
R1868 VSS.n187 VSS.n186 0.00298619
R1869 VSS VSS.n103 0.00294898
R1870 VSS VSS.n247 0.00293243
R1871 VSS.n250 VSS 0.00293243
R1872 VSS.n407 VSS.n406 0.00279385
R1873 VSS.n380 VSS 0.00258494
R1874 VSS.n378 VSS 0.00258494
R1875 VSS.n150 VSS 0.00233673
R1876 VSS VSS.n106 0.00219811
R1877 VSS.n147 VSS 0.00219811
R1878 VSS.n292 VSS 0.00219811
R1879 VSS.n162 VSS 0.00219811
R1880 VSS VSS.n212 0.00219811
R1881 VSS.n281 VSS 0.00219811
R1882 VSS.n262 VSS 0.00219811
R1883 VSS.n197 VSS 0.00219811
R1884 VSS VSS.n192 0.00219811
R1885 VSS.n329 VSS 0.00219811
R1886 VSS.n71 VSS 0.00219811
R1887 VSS.n361 VSS 0.00219811
R1888 VSS VSS.n88 0.00219811
R1889 VSS.n351 VSS 0.00219811
R1890 VSS.n4 VSS 0.00219811
R1891 VSS VSS.n181 0.00215138
R1892 VSS.n411 VSS.n410 0.00211919
R1893 VSS VSS.n377 0.00191732
R1894 VSS.n368 VSS 0.00191732
R1895 VSS VSS.n384 0.00188996
R1896 VSS VSS.n382 0.00188996
R1897 VSS.n255 VSS 0.00171622
R1898 VSS.n257 VSS 0.00171622
R1899 VSS VSS.n215 0.00157143
R1900 VSS.n194 VSS 0.0015
R1901 VSS VSS.n440 0.00149815
R1902 VSS VSS.n438 0.00149815
R1903 VSS.n186 VSS 0.00149448
R1904 VSS.n189 VSS 0.00149448
R1905 VSS.n229 VSS 0.00136539
R1906 VSS.n110 VSS 0.00130959
R1907 VSS.n113 VSS 0.00130959
R1908 VSS.n116 VSS 0.00130959
R1909 VSS.n120 VSS 0.00130959
R1910 VSS.n413 VSS 0.00130959
R1911 VSS VSS.n412 0.00130959
R1912 VSS.n409 VSS 0.00130959
R1913 VSS VSS.n408 0.00130959
R1914 VSS.n394 VSS 0.00130959
R1915 VSS VSS.n393 0.00130959
R1916 VSS.n390 VSS 0.00130959
R1917 VSS VSS.n389 0.00130959
R1918 VSS VSS.n285 0.0013
R1919 VSS.n277 VSS.n267 0.00129295
R1920 VSS VSS.n267 0.00129295
R1921 VSS.n435 VSS 0.00103973
R1922 VSS VSS.n432 0.00103973
R1923 VSS.n431 VSS 0.00103973
R1924 VSS.n15 VSS 0.00103973
R1925 VSS.n133 VSS 0.00103973
R1926 VSS VSS.n132 0.00103973
R1927 VSS.n129 VSS 0.00103973
R1928 VSS VSS.n128 0.00103973
R1929 VSS.n404 VSS 0.00103973
R1930 VSS VSS.n401 0.00103973
R1931 VSS.n400 VSS 0.00103973
R1932 VSS VSS.n397 0.00103973
R1933 VSS.n278 VSS.n277 0.000896476
R1934 CLK_div_3_mag_0.JK_FF_mag_1.K.n3 CLK_div_3_mag_0.JK_FF_mag_1.K.t6 37.1981
R1935 CLK_div_3_mag_0.JK_FF_mag_1.K.n5 CLK_div_3_mag_0.JK_FF_mag_1.K.t4 31.4332
R1936 CLK_div_3_mag_0.JK_FF_mag_1.K.n4 CLK_div_3_mag_0.JK_FF_mag_1.K.t7 30.4613
R1937 CLK_div_3_mag_0.JK_FF_mag_1.K.n4 CLK_div_3_mag_0.JK_FF_mag_1.K.t3 24.7562
R1938 CLK_div_3_mag_0.JK_FF_mag_1.K.n3 CLK_div_3_mag_0.JK_FF_mag_1.K.t5 17.6611
R1939 CLK_div_3_mag_0.JK_FF_mag_1.K.n5 CLK_div_3_mag_0.JK_FF_mag_1.K.t2 15.3826
R1940 CLK_div_3_mag_0.JK_FF_mag_1.K.n0 CLK_div_3_mag_0.JK_FF_mag_1.K 12.0716
R1941 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.K.n5 7.62076
R1942 CLK_div_3_mag_0.JK_FF_mag_1.K.n6 CLK_div_3_mag_0.JK_FF_mag_1.K 6.09789
R1943 CLK_div_3_mag_0.JK_FF_mag_1.K.n7 CLK_div_3_mag_0.JK_FF_mag_1.K.n2 2.99416
R1944 CLK_div_3_mag_0.JK_FF_mag_1.K.n2 CLK_div_3_mag_0.JK_FF_mag_1.K.t0 2.2755
R1945 CLK_div_3_mag_0.JK_FF_mag_1.K.n2 CLK_div_3_mag_0.JK_FF_mag_1.K.n1 2.2755
R1946 CLK_div_3_mag_0.JK_FF_mag_1.K.n7 CLK_div_3_mag_0.JK_FF_mag_1.K.n6 2.2505
R1947 CLK_div_3_mag_0.JK_FF_mag_1.K.n0 CLK_div_3_mag_0.JK_FF_mag_1.K 2.24788
R1948 CLK_div_3_mag_0.JK_FF_mag_1.K.n6 CLK_div_3_mag_0.JK_FF_mag_1.K.n0 1.94903
R1949 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.K.n4 1.81638
R1950 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.K.n3 1.43706
R1951 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.K.n7 0.4325
R1952 CLK_div_3_mag_1.Q0.n2 CLK_div_3_mag_1.Q0.t8 36.935
R1953 CLK_div_3_mag_1.Q0.n3 CLK_div_3_mag_1.Q0.t4 31.4332
R1954 CLK_div_3_mag_1.Q0.n5 CLK_div_3_mag_1.Q0.t6 29.8135
R1955 CLK_div_3_mag_1.Q0.n5 CLK_div_3_mag_1.Q0.t5 27.8352
R1956 CLK_div_3_mag_1.Q0.n2 CLK_div_3_mag_1.Q0.t7 18.1962
R1957 CLK_div_3_mag_1.Q0.n3 CLK_div_3_mag_1.Q0.t3 15.3826
R1958 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.Q0.t1 7.09905
R1959 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.Q0.n3 6.86029
R1960 CLK_div_3_mag_1.Q0.n4 CLK_div_3_mag_1.Q0 5.01077
R1961 CLK_div_3_mag_1.Q0.n6 CLK_div_3_mag_1.Q0 3.41843
R1962 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.Q0.n1 3.25053
R1963 CLK_div_3_mag_1.Q0.n1 CLK_div_3_mag_1.Q0.t2 2.2755
R1964 CLK_div_3_mag_1.Q0.n1 CLK_div_3_mag_1.Q0.n0 2.2755
R1965 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.Q0.n6 2.2505
R1966 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.Q0.n2 2.13459
R1967 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.Q0.n5 1.74998
R1968 CLK_div_3_mag_1.Q0.n6 CLK_div_3_mag_1.Q0.n4 1.50381
R1969 CLK_div_3_mag_1.Q0.n4 CLK_div_3_mag_1.Q0 1.12067
R1970 CLK_div_3_mag_1.JK_FF_mag_1.K.n3 CLK_div_3_mag_1.JK_FF_mag_1.K.t4 37.1981
R1971 CLK_div_3_mag_1.JK_FF_mag_1.K.n5 CLK_div_3_mag_1.JK_FF_mag_1.K.t3 31.4332
R1972 CLK_div_3_mag_1.JK_FF_mag_1.K.n4 CLK_div_3_mag_1.JK_FF_mag_1.K.t5 30.4613
R1973 CLK_div_3_mag_1.JK_FF_mag_1.K.n4 CLK_div_3_mag_1.JK_FF_mag_1.K.t7 24.7562
R1974 CLK_div_3_mag_1.JK_FF_mag_1.K.n3 CLK_div_3_mag_1.JK_FF_mag_1.K.t2 17.6611
R1975 CLK_div_3_mag_1.JK_FF_mag_1.K.n5 CLK_div_3_mag_1.JK_FF_mag_1.K.t6 15.3826
R1976 CLK_div_3_mag_1.JK_FF_mag_1.K.n0 CLK_div_3_mag_1.JK_FF_mag_1.K 12.0716
R1977 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.K.n5 7.62076
R1978 CLK_div_3_mag_1.JK_FF_mag_1.K.n6 CLK_div_3_mag_1.JK_FF_mag_1.K 6.09789
R1979 CLK_div_3_mag_1.JK_FF_mag_1.K.n7 CLK_div_3_mag_1.JK_FF_mag_1.K.n2 2.99416
R1980 CLK_div_3_mag_1.JK_FF_mag_1.K.n2 CLK_div_3_mag_1.JK_FF_mag_1.K.t0 2.2755
R1981 CLK_div_3_mag_1.JK_FF_mag_1.K.n2 CLK_div_3_mag_1.JK_FF_mag_1.K.n1 2.2755
R1982 CLK_div_3_mag_1.JK_FF_mag_1.K.n7 CLK_div_3_mag_1.JK_FF_mag_1.K.n6 2.2505
R1983 CLK_div_3_mag_1.JK_FF_mag_1.K.n0 CLK_div_3_mag_1.JK_FF_mag_1.K 2.24788
R1984 CLK_div_3_mag_1.JK_FF_mag_1.K.n6 CLK_div_3_mag_1.JK_FF_mag_1.K.n0 1.94903
R1985 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.K.n4 1.81638
R1986 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.K.n3 1.43706
R1987 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.K.n7 0.4325
R1988 CLK_div_3_mag_1.Q1.n5 CLK_div_3_mag_1.Q1.t7 36.935
R1989 CLK_div_3_mag_1.Q1.n2 CLK_div_3_mag_1.Q1.t5 31.4332
R1990 CLK_div_3_mag_1.Q1.n6 CLK_div_3_mag_1.Q1.t9 31.4332
R1991 CLK_div_3_mag_1.Q1.n3 CLK_div_3_mag_1.Q1.t10 30.4613
R1992 CLK_div_3_mag_1.Q1.n3 CLK_div_3_mag_1.Q1.t4 24.7562
R1993 CLK_div_3_mag_1.Q1.n5 CLK_div_3_mag_1.Q1.t3 18.1962
R1994 CLK_div_3_mag_1.Q1.n2 CLK_div_3_mag_1.Q1.t6 15.3826
R1995 CLK_div_3_mag_1.Q1.n6 CLK_div_3_mag_1.Q1.t8 15.3826
R1996 CLK_div_3_mag_1.Q1.n4 CLK_div_3_mag_1.Q1 8.5575
R1997 CLK_div_3_mag_1.Q1 CLK_div_3_mag_1.Q1.t1 7.09905
R1998 CLK_div_3_mag_1.Q1 CLK_div_3_mag_1.Q1.n6 6.86029
R1999 CLK_div_3_mag_1.Q1.n2 CLK_div_3_mag_1.Q1 5.69501
R2000 CLK_div_3_mag_1.Q1.n7 CLK_div_3_mag_1.Q1 5.01077
R2001 CLK_div_3_mag_1.Q1 CLK_div_3_mag_1.Q1.n1 3.25053
R2002 CLK_div_3_mag_1.Q1 CLK_div_3_mag_1.Q1.n8 2.43532
R2003 CLK_div_3_mag_1.Q1.n1 CLK_div_3_mag_1.Q1.t2 2.2755
R2004 CLK_div_3_mag_1.Q1.n1 CLK_div_3_mag_1.Q1.n0 2.2755
R2005 CLK_div_3_mag_1.Q1 CLK_div_3_mag_1.Q1.n5 2.13459
R2006 CLK_div_3_mag_1.Q1 CLK_div_3_mag_1.Q1.n3 1.81638
R2007 CLK_div_3_mag_1.Q1.n8 CLK_div_3_mag_1.Q1.n7 1.45395
R2008 CLK_div_3_mag_1.Q1.n8 CLK_div_3_mag_1.Q1.n4 1.23718
R2009 CLK_div_3_mag_1.Q1.n7 CLK_div_3_mag_1.Q1 1.12067
R2010 CLK_div_3_mag_1.Q1.n4 CLK_div_3_mag_1.Q1 0.976433
R2011 CLK_div_3_mag_0.CLK.n8 CLK_div_3_mag_0.CLK.t3 36.935
R2012 CLK_div_3_mag_0.CLK.n7 CLK_div_3_mag_0.CLK.t6 36.935
R2013 CLK_div_3_mag_0.CLK.n12 CLK_div_3_mag_0.CLK.t12 36.935
R2014 CLK_div_3_mag_0.CLK.n9 CLK_div_3_mag_0.CLK.t11 36.935
R2015 CLK_div_3_mag_0.CLK.n10 CLK_div_3_mag_0.CLK.t5 30.5752
R2016 CLK_div_3_mag_0.CLK.n13 CLK_div_3_mag_0.CLK.t10 25.4744
R2017 CLK_div_3_mag_0.CLK.n6 CLK_div_3_mag_0.CLK.t8 25.4742
R2018 CLK_div_3_mag_0.CLK.n10 CLK_div_3_mag_0.CLK.t4 21.7814
R2019 CLK_div_3_mag_0.CLK.n8 CLK_div_3_mag_0.CLK.t14 18.1962
R2020 CLK_div_3_mag_0.CLK.n7 CLK_div_3_mag_0.CLK.t2 18.1962
R2021 CLK_div_3_mag_0.CLK.n12 CLK_div_3_mag_0.CLK.t9 18.1962
R2022 CLK_div_3_mag_0.CLK.n9 CLK_div_3_mag_0.CLK.t7 18.1962
R2023 CLK_div_3_mag_0.CLK.n6 CLK_div_3_mag_0.CLK.t13 14.142
R2024 CLK_div_3_mag_0.CLK.n13 CLK_div_3_mag_0.CLK.t15 14.1417
R2025 CLK_div_3_mag_0.CLK.n5 CLK_div_3_mag_0.CLK.t1 9.33985
R2026 CLK_div_3_mag_0.CLK.n0 CLK_div_3_mag_0.CLK.n11 7.41483
R2027 CLK_div_3_mag_0.CLK.n15 CLK_div_3_mag_0.CLK.n14 5.37091
R2028 CLK_div_3_mag_0.CLK.n5 CLK_div_3_mag_0.CLK.t0 5.17836
R2029 CLK_div_3_mag_0.CLK.n2 CLK_div_3_mag_0.CLK.n12 2.13265
R2030 CLK_div_3_mag_0.CLK.n2 CLK_div_3_mag_0.CLK 0.077103
R2031 CLK_div_3_mag_0.CLK.n13 CLK_div_3_mag_0.CLK.n3 1.42996
R2032 CLK_div_3_mag_0.CLK.n0 CLK_div_3_mag_0.CLK.n2 1.11863
R2033 CLK_div_3_mag_0.CLK.n14 CLK_div_3_mag_0.CLK.n3 1.19586
R2034 CLK_div_3_mag_0.CLK CLK_div_3_mag_0.CLK.n8 2.13265
R2035 CLK_div_3_mag_0.CLK.n11 CLK_div_3_mag_0.CLK.n10 1.80883
R2036 CLK_div_3_mag_0.CLK.n1 CLK_div_3_mag_0.CLK 2.63776
R2037 CLK_div_3_mag_0.CLK.n0 CLK_div_3_mag_0.CLK 2.51943
R2038 CLK_div_3_mag_0.CLK.n9 CLK_div_3_mag_0.CLK 2.13281
R2039 CLK_div_3_mag_0.CLK.n7 CLK_div_3_mag_0.CLK 2.13261
R2040 CLK_div_3_mag_0.CLK.n4 CLK_div_3_mag_0.CLK.n6 1.43004
R2041 CLK_div_3_mag_0.CLK.n3 CLK_div_3_mag_0.CLK 0.196041
R2042 CLK_div_3_mag_0.CLK CLK_div_3_mag_0.CLK.n4 0.196041
R2043 CLK_div_3_mag_0.CLK CLK_div_3_mag_0.CLK.n5 0.115328
R2044 CLK_div_3_mag_0.CLK.n11 CLK_div_3_mag_0.CLK 0.108371
R2045 CLK_div_3_mag_0.CLK.n4 CLK_div_3_mag_0.CLK.n15 1.19586
R2046 CLK_div_3_mag_0.CLK.n1 CLK_div_3_mag_0.CLK 1.11863
R2047 CLK_div_3_mag_0.CLK.n14 CLK_div_3_mag_0.CLK.n0 1.01264
R2048 CLK_div_3_mag_0.CLK.n15 CLK_div_3_mag_0.CLK.n1 0.894314
R2049 CLK.n1 CLK.t5 36.935
R2050 CLK.n7 CLK.t11 36.935
R2051 CLK.n13 CLK.t7 36.935
R2052 CLK.n17 CLK.t8 36.935
R2053 CLK.n23 CLK.t3 30.5752
R2054 CLK.n30 CLK.t1 25.4744
R2055 CLK.n37 CLK.t12 25.4742
R2056 CLK.n23 CLK.t0 21.7814
R2057 CLK.n1 CLK.t13 18.1962
R2058 CLK.n7 CLK.t10 18.1962
R2059 CLK.n13 CLK.t2 18.1962
R2060 CLK.n17 CLK.t4 18.1962
R2061 CLK.n37 CLK.t6 14.142
R2062 CLK.n30 CLK.t9 14.1417
R2063 CLK.n25 CLK.n24 7.41483
R2064 CLK.n35 CLK.n34 5.37091
R2065 CLK.n12 CLK.n4 2.25107
R2066 CLK.n27 CLK.n16 2.25107
R2067 CLK.n33 CLK.n32 2.24352
R2068 CLK.n39 CLK.n36 2.24352
R2069 CLK.n20 CLK.n17 2.12464
R2070 CLK.n8 CLK.n7 2.12444
R2071 CLK.n2 CLK.n1 2.12188
R2072 CLK.n14 CLK.n13 2.12188
R2073 CLK.n24 CLK.n23 1.80883
R2074 CLK.n11 CLK.n10 1.71671
R2075 CLK.n25 CLK.n22 1.59838
R2076 CLK.n9 CLK.n8 1.50503
R2077 CLK.n21 CLK.n20 1.50503
R2078 CLK.n38 CLK.n37 1.42126
R2079 CLK.n31 CLK.n30 1.42118
R2080 CLK.n35 CLK.n12 0.882596
R2081 CLK.n34 CLK.n27 0.882596
R2082 CLK.n29 CLK 0.1605
R2083 CLK.n26 CLK.n25 0.118826
R2084 CLK.n24 CLK 0.108371
R2085 CLK.n34 CLK.n33 0.0733415
R2086 CLK.n36 CLK.n35 0.0733415
R2087 CLK CLK.n40 0.05925
R2088 CLK.n3 CLK 0.0457995
R2089 CLK.n5 CLK 0.0457995
R2090 CLK.n15 CLK 0.0457995
R2091 CLK.n18 CLK 0.0457995
R2092 CLK.n10 CLK.n9 0.0386356
R2093 CLK.n22 CLK.n21 0.0386356
R2094 CLK.n4 CLK.n3 0.0377414
R2095 CLK.n6 CLK.n5 0.0377414
R2096 CLK.n16 CLK.n15 0.0377414
R2097 CLK.n19 CLK.n18 0.0377414
R2098 CLK.n32 CLK.n29 0.03175
R2099 CLK.n40 CLK.n39 0.03175
R2100 CLK.n33 CLK.n28 0.0198632
R2101 CLK.n36 CLK.n0 0.0198632
R2102 CLK.n12 CLK.n11 0.0122182
R2103 CLK.n27 CLK.n26 0.0122182
R2104 CLK.n4 CLK.n2 0.00360345
R2105 CLK.n16 CLK.n14 0.00360345
R2106 CLK.n8 CLK.n6 0.00203726
R2107 CLK.n20 CLK.n19 0.00203726
R2108 CLK.n32 CLK.n31 0.00175
R2109 CLK.n39 CLK.n38 0.00175
R2110 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n2 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t8 37.1986
R2111 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n1 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t3 31.528
R2112 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n0 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t5 30.6344
R2113 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n0 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t4 27.3855
R2114 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n2 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t7 17.6614
R2115 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n1 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t6 15.3826
R2116 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n1 7.62751
R2117 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n3 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 6.09789
R2118 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n0 2.8877
R2119 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n3 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 2.67866
R2120 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t0 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n3 2.2505
R2121 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n2 1.43709
R2122 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t0 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.4325
R2123 CLK_div_3_mag_0.Q1.n5 CLK_div_3_mag_0.Q1.t9 36.935
R2124 CLK_div_3_mag_0.Q1.n2 CLK_div_3_mag_0.Q1.t8 31.4332
R2125 CLK_div_3_mag_0.Q1.n6 CLK_div_3_mag_0.Q1.t5 31.4332
R2126 CLK_div_3_mag_0.Q1.n3 CLK_div_3_mag_0.Q1.t4 30.4613
R2127 CLK_div_3_mag_0.Q1.n3 CLK_div_3_mag_0.Q1.t7 24.7562
R2128 CLK_div_3_mag_0.Q1.n5 CLK_div_3_mag_0.Q1.t6 18.1962
R2129 CLK_div_3_mag_0.Q1.n2 CLK_div_3_mag_0.Q1.t10 15.3826
R2130 CLK_div_3_mag_0.Q1.n6 CLK_div_3_mag_0.Q1.t3 15.3826
R2131 CLK_div_3_mag_0.Q1.n4 CLK_div_3_mag_0.Q1 8.5575
R2132 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.Q1.t2 7.09905
R2133 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.Q1.n6 6.86029
R2134 CLK_div_3_mag_0.Q1.n2 CLK_div_3_mag_0.Q1 5.69501
R2135 CLK_div_3_mag_0.Q1.n7 CLK_div_3_mag_0.Q1 5.01077
R2136 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.Q1.n1 3.25053
R2137 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.Q1.n8 2.43532
R2138 CLK_div_3_mag_0.Q1.n1 CLK_div_3_mag_0.Q1.t0 2.2755
R2139 CLK_div_3_mag_0.Q1.n1 CLK_div_3_mag_0.Q1.n0 2.2755
R2140 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.Q1.n5 2.13459
R2141 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.Q1.n3 1.81638
R2142 CLK_div_3_mag_0.Q1.n8 CLK_div_3_mag_0.Q1.n7 1.45395
R2143 CLK_div_3_mag_0.Q1.n8 CLK_div_3_mag_0.Q1.n4 1.23718
R2144 CLK_div_3_mag_0.Q1.n7 CLK_div_3_mag_0.Q1 1.12067
R2145 CLK_div_3_mag_0.Q1.n4 CLK_div_3_mag_0.Q1 0.976433
R2146 RST.n56 RST.t10 37.2596
R2147 RST.n44 RST.t0 37.2596
R2148 RST.n64 RST.t9 36.935
R2149 RST.n51 RST.t4 36.935
R2150 RST.n7 RST.t12 36.935
R2151 RST.n0 RST.t2 36.935
R2152 RST.n20 RST.t15 36.935
R2153 RST.n34 RST.t13 36.935
R2154 RST.n64 RST.t5 18.1962
R2155 RST.n51 RST.t1 18.1962
R2156 RST.n7 RST.t7 18.1962
R2157 RST.n0 RST.t3 18.1962
R2158 RST.n20 RST.t8 18.1962
R2159 RST.n34 RST.t14 18.1962
R2160 RST.n56 RST.t6 17.5947
R2161 RST.n44 RST.t11 17.5947
R2162 RST.n68 RST.n61 6.06869
R2163 RST.n61 RST.n54 4.82595
R2164 RST.n68 RST.n67 4.82279
R2165 RST.n61 RST.n60 4.5933
R2166 RST.n27 RST.n26 4.51211
R2167 RST.n67 RST.n66 4.5005
R2168 RST.n54 RST.n53 4.5005
R2169 RST.n22 RST.n19 4.5005
R2170 RST.n22 RST.n21 4.5005
R2171 RST.n25 RST.n23 4.5005
R2172 RST.n25 RST.n24 4.5005
R2173 RST.n69 RST.n48 4.15909
R2174 RST.n72 RST.n70 3.36603
R2175 RST.n72 RST.n71 2.25598
R2176 RST.n10 RST.n9 2.2505
R2177 RST.n65 RST.n63 2.25022
R2178 RST.n52 RST.n50 2.25022
R2179 RST.n28 RST.n27 2.24707
R2180 RST.n60 RST.n59 2.24196
R2181 RST.n48 RST.n47 2.24196
R2182 RST.n65 RST.n64 2.12393
R2183 RST.n52 RST.n51 2.12393
R2184 RST.n1 RST.n0 2.12318
R2185 RST.n21 RST.n20 2.12318
R2186 RST.n35 RST.n34 2.1224
R2187 RST.n8 RST.n7 2.12188
R2188 RST.n15 RST.n14 1.90023
R2189 RST.n17 RST.n16 1.88263
R2190 RST.n30 RST.n29 1.86678
R2191 RST.n37 RST.n36 1.5005
R2192 RST.n39 RST.n38 1.5005
R2193 RST.n13 RST.n12 1.5005
R2194 RST.n57 RST.n56 1.42168
R2195 RST.n45 RST.n44 1.42168
R2196 RST.n16 RST.n4 1.13307
R2197 RST.n3 RST.n2 0.898107
R2198 RST.n70 RST.n69 0.668278
R2199 RST.n42 RST.n41 0.643971
R2200 RST.n69 RST.n68 0.309974
R2201 RST.n70 RST.n42 0.136193
R2202 RST.n62 RST 0.0584663
R2203 RST.n49 RST 0.0584663
R2204 RST.n2 RST 0.0518307
R2205 RST.n58 RST 0.0394837
R2206 RST.n46 RST 0.0394837
R2207 RST.n59 RST.n58 0.0377414
R2208 RST.n47 RST.n46 0.0377414
R2209 RST.n33 RST 0.0363802
R2210 RST.n9 RST.n6 0.0361897
R2211 RST.n36 RST.n33 0.0346379
R2212 RST.n6 RST 0.031725
R2213 RST.n67 RST 0.0293
R2214 RST.n54 RST 0.0293
R2215 RST.n2 RST.n1 0.0249551
R2216 RST.n23 RST 0.0239664
R2217 RST.n60 RST.n55 0.0238218
R2218 RST.n48 RST.n43 0.0238218
R2219 RST.n22 RST.n18 0.0236959
R2220 RST.n14 RST.n13 0.0205676
R2221 RST.n66 RST.n62 0.0196058
R2222 RST.n53 RST.n49 0.0196058
R2223 RST.n39 RST.n30 0.0193514
R2224 RST.n38 RST.n31 0.0181289
R2225 RST.n29 RST.n28 0.0144865
R2226 RST.n27 RST.n25 0.0130264
R2227 RST.n9 RST.n8 0.0129138
R2228 RST.n16 RST.n15 0.0117735
R2229 RST.n10 RST.n5 0.0116103
R2230 RST.n36 RST.n35 0.00825862
R2231 RST.n28 RST.n17 0.0077973
R2232 RST RST.n72 0.00597826
R2233 RST.n12 RST.n11 0.00513918
R2234 RST.n37 RST.n32 0.00513918
R2235 RST.n59 RST.n57 0.00360345
R2236 RST.n47 RST.n45 0.00360345
R2237 RST.n12 RST.n10 0.00328351
R2238 RST.n4 RST.n3 0.00328351
R2239 RST.n38 RST.n37 0.00328351
R2240 RST.n66 RST.n65 0.00255119
R2241 RST.n53 RST.n52 0.00255119
R2242 RST.n40 RST.n39 0.00232432
R2243 RST.n41 RST.n40 0.00232432
R2244 RST.n63 RST 0.0017
R2245 RST.n50 RST 0.0017
R2246 RST.n25 RST.n22 0.00142783
R2247 RST.n42 RST 0.00104528
R2248 CLK_div_3_mag_0.Vdiv3.n20 CLK_div_3_mag_0.Vdiv3.t3 36.935
R2249 CLK_div_3_mag_0.Vdiv3.n19 CLK_div_3_mag_0.Vdiv3.t9 36.935
R2250 CLK_div_3_mag_0.Vdiv3.n30 CLK_div_3_mag_0.Vdiv3.t12 36.935
R2251 CLK_div_3_mag_0.Vdiv3.n29 CLK_div_3_mag_0.Vdiv3.t17 36.935
R2252 CLK_div_3_mag_0.Vdiv3.n28 CLK_div_3_mag_0.Vdiv3.t11 36.935
R2253 CLK_div_3_mag_0.Vdiv3.n26 CLK_div_3_mag_0.Vdiv3.t21 36.935
R2254 CLK_div_3_mag_0.Vdiv3.n25 CLK_div_3_mag_0.Vdiv3.t26 36.935
R2255 CLK_div_3_mag_0.Vdiv3.n23 CLK_div_3_mag_0.Vdiv3.t5 36.935
R2256 CLK_div_3_mag_0.Vdiv3.n22 CLK_div_3_mag_0.Vdiv3.t15 36.935
R2257 CLK_div_3_mag_0.Vdiv3.n21 CLK_div_3_mag_0.Vdiv3.t2 25.5364
R2258 CLK_div_3_mag_0.Vdiv3.n27 CLK_div_3_mag_0.Vdiv3.t16 25.5364
R2259 CLK_div_3_mag_0.Vdiv3.n24 CLK_div_3_mag_0.Vdiv3.t25 25.5364
R2260 CLK_div_3_mag_0.Vdiv3.n31 CLK_div_3_mag_0.Vdiv3.t27 25.5361
R2261 CLK_div_3_mag_0.Vdiv3.n20 CLK_div_3_mag_0.Vdiv3.t22 18.1962
R2262 CLK_div_3_mag_0.Vdiv3.n19 CLK_div_3_mag_0.Vdiv3.t10 18.1962
R2263 CLK_div_3_mag_0.Vdiv3.n30 CLK_div_3_mag_0.Vdiv3.t4 18.1962
R2264 CLK_div_3_mag_0.Vdiv3.n29 CLK_div_3_mag_0.Vdiv3.t18 18.1962
R2265 CLK_div_3_mag_0.Vdiv3.n28 CLK_div_3_mag_0.Vdiv3.t8 18.1962
R2266 CLK_div_3_mag_0.Vdiv3.n26 CLK_div_3_mag_0.Vdiv3.t13 18.1962
R2267 CLK_div_3_mag_0.Vdiv3.n25 CLK_div_3_mag_0.Vdiv3.t19 18.1962
R2268 CLK_div_3_mag_0.Vdiv3.n23 CLK_div_3_mag_0.Vdiv3.t23 18.1962
R2269 CLK_div_3_mag_0.Vdiv3.n22 CLK_div_3_mag_0.Vdiv3.t7 18.1962
R2270 CLK_div_3_mag_0.Vdiv3.n27 CLK_div_3_mag_0.Vdiv3.t24 14.0749
R2271 CLK_div_3_mag_0.Vdiv3.n24 CLK_div_3_mag_0.Vdiv3.t6 14.0749
R2272 CLK_div_3_mag_0.Vdiv3.n21 CLK_div_3_mag_0.Vdiv3.t20 14.0749
R2273 CLK_div_3_mag_0.Vdiv3.n31 CLK_div_3_mag_0.Vdiv3.t14 14.0734
R2274 CLK_div_3_mag_0.Vdiv3.n18 CLK_div_3_mag_0.Vdiv3.t1 9.33985
R2275 CLK_div_3_mag_0.Vdiv3.n33 CLK_div_3_mag_0.Vdiv3 5.77906
R2276 CLK_div_3_mag_0.Vdiv3.n18 CLK_div_3_mag_0.Vdiv3.t0 5.17836
R2277 CLK_div_3_mag_0.Vdiv3.n35 CLK_div_3_mag_0.Vdiv3.n34 5.11659
R2278 CLK_div_3_mag_0.Vdiv3.n10 CLK_div_3_mag_0.Vdiv3.n19 2.13042
R2279 CLK_div_3_mag_0.Vdiv3.n3 CLK_div_3_mag_0.Vdiv3.n2 1.11863
R2280 CLK_div_3_mag_0.Vdiv3.n11 CLK_div_3_mag_0.Vdiv3.n29 2.13042
R2281 CLK_div_3_mag_0.Vdiv3.n5 CLK_div_3_mag_0.Vdiv3.n4 1.11863
R2282 CLK_div_3_mag_0.Vdiv3.n14 CLK_div_3_mag_0.Vdiv3.n31 1.43628
R2283 CLK_div_3_mag_0.Vdiv3.n0 CLK_div_3_mag_0.Vdiv3.n32 4.94724
R2284 CLK_div_3_mag_0.Vdiv3.n12 CLK_div_3_mag_0.Vdiv3.n25 2.13042
R2285 CLK_div_3_mag_0.Vdiv3.n7 CLK_div_3_mag_0.Vdiv3.n6 1.11863
R2286 CLK_div_3_mag_0.Vdiv3.n15 CLK_div_3_mag_0.Vdiv3.n27 1.43559
R2287 CLK_div_3_mag_0.Vdiv3.n13 CLK_div_3_mag_0.Vdiv3.n22 2.13042
R2288 CLK_div_3_mag_0.Vdiv3.n9 CLK_div_3_mag_0.Vdiv3.n8 1.11863
R2289 CLK_div_3_mag_0.Vdiv3.n16 CLK_div_3_mag_0.Vdiv3.n24 1.43559
R2290 CLK_div_3_mag_0.Vdiv3.n1 CLK_div_3_mag_0.Vdiv3.n17 1.49204
R2291 CLK_div_3_mag_0.Vdiv3.n36 CLK_div_3_mag_0.Vdiv3.n35 4.5005
R2292 CLK_div_3_mag_0.Vdiv3.n34 CLK_div_3_mag_0.Vdiv3 4.43149
R2293 CLK_div_3_mag_0.Vdiv3.n33 CLK_div_3_mag_0.Vdiv3.n32 3.5258
R2294 CLK_div_3_mag_0.Vdiv3.n32 CLK_div_3_mag_0.Vdiv3 2.3355
R2295 CLK_div_3_mag_0.Vdiv3.n3 CLK_div_3_mag_0.Vdiv3.n20 2.13151
R2296 CLK_div_3_mag_0.Vdiv3.n5 CLK_div_3_mag_0.Vdiv3.n30 2.13151
R2297 CLK_div_3_mag_0.Vdiv3.n7 CLK_div_3_mag_0.Vdiv3.n26 2.13151
R2298 CLK_div_3_mag_0.Vdiv3.n9 CLK_div_3_mag_0.Vdiv3.n23 2.13151
R2299 CLK_div_3_mag_0.Vdiv3.n2 CLK_div_3_mag_0.Vdiv3.n10 2.63808
R2300 CLK_div_3_mag_0.Vdiv3.n4 CLK_div_3_mag_0.Vdiv3.n11 2.63808
R2301 CLK_div_3_mag_0.Vdiv3.n6 CLK_div_3_mag_0.Vdiv3.n12 2.63808
R2302 CLK_div_3_mag_0.Vdiv3.n8 CLK_div_3_mag_0.Vdiv3.n13 2.63808
R2303 CLK_div_3_mag_0.Vdiv3.n16 CLK_div_3_mag_0.Vdiv3.n8 2.10738
R2304 CLK_div_3_mag_0.Vdiv3.n15 CLK_div_3_mag_0.Vdiv3.n6 2.10738
R2305 CLK_div_3_mag_0.Vdiv3.n14 CLK_div_3_mag_0.Vdiv3.n4 2.10738
R2306 CLK_div_3_mag_0.Vdiv3.n34 CLK_div_3_mag_0.Vdiv3.n33 1.62556
R2307 CLK_div_3_mag_0.Vdiv3.n17 CLK_div_3_mag_0.Vdiv3.n21 1.42706
R2308 CLK_div_3_mag_0.Vdiv3.n2 CLK_div_3_mag_0.Vdiv3.n1 0.991659
R2309 CLK_div_3_mag_0.Vdiv3 CLK_div_3_mag_0.Vdiv3.n36 0.1705
R2310 CLK_div_3_mag_0.Vdiv3 CLK_div_3_mag_0.Vdiv3.n18 0.115328
R2311 CLK_div_3_mag_0.Vdiv3.n0 CLK_div_3_mag_0.Vdiv3 0.0684998
R2312 CLK_div_3_mag_0.Vdiv3.n3 CLK_div_3_mag_0.Vdiv3 0.0786548
R2313 CLK_div_3_mag_0.Vdiv3.n10 CLK_div_3_mag_0.Vdiv3 0.0807313
R2314 CLK_div_3_mag_0.Vdiv3.n5 CLK_div_3_mag_0.Vdiv3 0.0786548
R2315 CLK_div_3_mag_0.Vdiv3.n11 CLK_div_3_mag_0.Vdiv3 0.0807313
R2316 CLK_div_3_mag_0.Vdiv3.n7 CLK_div_3_mag_0.Vdiv3 0.0786548
R2317 CLK_div_3_mag_0.Vdiv3.n12 CLK_div_3_mag_0.Vdiv3 0.0807313
R2318 CLK_div_3_mag_0.Vdiv3.n9 CLK_div_3_mag_0.Vdiv3 0.0786548
R2319 CLK_div_3_mag_0.Vdiv3.n13 CLK_div_3_mag_0.Vdiv3 0.0807313
R2320 CLK_div_3_mag_0.Vdiv3.n36 CLK_div_3_mag_0.Vdiv3.n17 0.033
R2321 CLK_div_3_mag_0.Vdiv3 CLK_div_3_mag_0.Vdiv3.n16 0.1953
R2322 CLK_div_3_mag_0.Vdiv3 CLK_div_3_mag_0.Vdiv3.n15 0.1953
R2323 CLK_div_3_mag_0.Vdiv3 CLK_div_3_mag_0.Vdiv3.n14 0.1953
R2324 CLK_div_3_mag_0.Vdiv3.n35 CLK_div_3_mag_0.Vdiv3.n1 0.0170403
R2325 CLK_div_3_mag_0.Vdiv3.n0 CLK_div_3_mag_0.Vdiv3.n28 2.14709
R2326 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t4 30.9379
R2327 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n0 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t2 30.664
R2328 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n0 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t3 24.5385
R2329 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t5 24.5101
R2330 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n2 7.46763
R2331 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n3 5.28703
R2332 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n1 4.09208
R2333 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 3.12156
R2334 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 1.86016
R2335 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n0 1.4252
R2336 Vdiv99.n2 Vdiv99.n1 9.33985
R2337 Vdiv99.n2 Vdiv99.n0 5.17836
R2338 Vdiv99 Vdiv99.n2 0.115328
C0 a_5466_15136# CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.132f
C1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT RST 0.0834f
C2 a_14508_9798# VDD 3.14e-19
C3 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 2.56e-19
C4 a_10927_9798# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.0059f
C5 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 7.07e-19
C6 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.Q3 0.349f
C7 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.Q1 0.00825f
C8 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.198f
C9 a_5852_10895# VDD 0.00743f
C10 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.Q3 9.48e-20
C11 a_12221_10895# CLK_DIV_11_mag_new_0.Q1 5.98e-19
C12 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT a_6252_11889# 2.88e-20
C13 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 RST 0.0134f
C14 a_10961_15230# CLK_DIV_11_mag_new_0.nand3_mag_1.OUT 2.05e-19
C15 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.00975f
C16 CLK_div_3_mag_1.or_2_mag_0.IN2 a_10806_8231# 8.64e-19
C17 a_4968_10895# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 8.64e-19
C18 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 a_13629_11933# 0.00372f
C19 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_12501_11889# 0.0733f
C20 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.Q0 0.0709f
C21 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT VDD 0.643f
C22 a_12911_13030# CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 2.96e-19
C23 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_10515_11931# 0.0811f
C24 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 7.63e-19
C25 a_9951_11931# CLK_DIV_11_mag_new_0.Q2 0.00859f
C26 a_12347_13030# VDD 3.14e-19
C27 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 0.198f
C28 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.00183f
C29 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_1.Q0 0.107f
C30 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0894f
C31 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK 0.0983f
C32 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.0052f
C33 a_7985_10895# VDD 9.82e-19
C34 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.103f
C35 CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 0.294f
C36 a_4968_10895# a_5128_10895# 0.0504f
C37 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K VDD 0.593f
C38 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 0.129f
C39 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.Q2 6.13e-20
C40 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00158f
C41 a_13944_9798# VDD 3.14e-19
C42 a_2597_12515# CLK_DIV_11_mag_new_0.Q3 0.0111f
C43 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK 0.00481f
C44 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.Q0 1.65e-21
C45 CLK_div_3_mag_1.JK_FF_mag_1.K VDD 2.4f
C46 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.nand3_mag_0.OUT 4.36e-19
C47 a_5692_10895# VDD 0.00305f
C48 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0718f
C49 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.QB 7.08e-20
C50 CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_div_3_mag_0.JK_FF_mag_1.K 2.14e-21
C51 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT a_6092_11889# 9.1e-19
C52 a_12061_10895# CLK_DIV_11_mag_new_0.Q1 5.98e-19
C53 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.Q2 8.04e-19
C54 a_10256_15189# CLK_DIV_11_mag_new_0.nand3_mag_1.OUT 0.0731f
C55 CLK_div_3_mag_1.or_2_mag_0.IN2 a_11779_8699# 7.48e-20
C56 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 a_13065_11933# 0.069f
C57 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 RST 0.00289f
C58 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_12341_11889# 0.0203f
C59 RST CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 0.16f
C60 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_9951_11931# 0.00964f
C61 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.342f
C62 a_12347_13030# CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 3.08e-19
C63 a_9387_11887# CLK_DIV_11_mag_new_0.Q2 0.0101f
C64 a_11617_11889# CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 8.64e-19
C65 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD 0.653f
C66 a_8863_9798# CLK_div_3_mag_1.Q0 3.69e-19
C67 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 RST 1.36e-19
C68 a_6816_11933# CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.00964f
C69 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_15506_13026# 1.43e-19
C70 a_7421_10895# VDD 0.00149f
C71 a_13790_10895# CLK_DIV_11_mag_new_0.Q1 2.58e-20
C72 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT VDD 0.994f
C73 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_12215_9798# 0.0203f
C74 CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 0.0108f
C75 CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN VDD 0.425f
C76 a_13380_9798# VDD 3.56e-19
C77 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.765f
C78 a_10961_15230# CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 3.04e-20
C79 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD 0.652f
C80 a_5122_9798# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0202f
C81 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 1.57f
C82 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 1.33e-19
C83 a_5128_10895# VDD 2.21e-19
C84 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 2.62e-20
C85 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT a_5528_11889# 0.0731f
C86 a_10096_15189# CLK_DIV_11_mag_new_0.nand3_mag_1.OUT 0.0202f
C87 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_11777_11889# 1.5e-20
C88 a_8863_9798# RST 6.26e-19
C89 a_16070_13026# CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 4.52e-20
C90 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.233f
C91 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 a_9387_11887# 8.64e-19
C92 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_9387_11887# 0.00696f
C93 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 a_7380_11933# 0.00372f
C94 a_11783_12986# CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.00392f
C95 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.Q3 2.92f
C96 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN 1.01e-19
C97 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT VDD 0.994f
C98 a_9227_11887# CLK_DIV_11_mag_new_0.Q2 0.0102f
C99 a_11623_12986# VDD 2.21e-19
C100 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 5.48e-20
C101 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.Q1 0.0309f
C102 a_16788_11929# VDD 3.14e-19
C103 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_9797_13028# 4.52e-20
C104 CLK CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.013f
C105 a_2597_12515# CLK_DIV_11_mag_new_0.Q1 0.00347f
C106 a_6252_11889# CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.00696f
C107 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_14942_12982# 0.00119f
C108 a_6857_10895# VDD 0.00149f
C109 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 4.67e-22
C110 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 7.17e-19
C111 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 4.69e-20
C112 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 5.73e-20
C113 a_8663_11887# CLK_DIV_11_mag_new_0.Q3 4.52e-19
C114 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_1.Q0 8.04e-19
C115 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_12055_9798# 0.0732f
C116 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 RST 0.0698f
C117 CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_DIV_11_mag_new_0.Q3 0.00935f
C118 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.Q3 1.04e-19
C119 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 3.81e-19
C120 a_3994_9798# VDD 3.56e-19
C121 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 6.11e-19
C122 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.Q0 0.0143f
C123 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.359f
C124 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 8.64e-20
C125 a_10256_15189# CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 8.5e-20
C126 CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_DIV_11_mag_new_0.Q3 0.161f
C127 a_4558_9798# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 4.52e-20
C128 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.Q2 0.0661f
C129 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT a_5368_11889# 0.0202f
C130 RST CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 0.00146f
C131 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0881f
C132 CLK_DIV_11_mag_new_0.and2_mag_3.IN1 VDD 0.798f
C133 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_11617_11889# 1.17e-20
C134 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_1.Q0 8.04e-19
C135 a_11337_10895# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 8.64e-19
C136 a_8703_9798# RST 5.13e-19
C137 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.0379f
C138 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 7.11e-19
C139 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_9227_11887# 0.00695f
C140 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 1.53e-19
C141 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_1.JK_FF_mag_1.QB 0.0576f
C142 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 0.00165f
C143 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 2.47e-19
C144 a_8663_11887# CLK_DIV_11_mag_new_0.Q2 0.00789f
C145 a_10361_13028# VDD 3.56e-19
C146 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 RST 0.0706f
C147 CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_DIV_11_mag_new_0.Q2 0.0814f
C148 a_16224_11929# VDD 3.14e-19
C149 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_9233_13028# 0.0195f
C150 a_6092_11889# CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.00695f
C151 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.Q0 0.0343f
C152 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 8.26e-20
C153 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_11491_9798# 0.00378f
C154 a_8503_11887# CLK_DIV_11_mag_new_0.Q3 5.83e-19
C155 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.QB 1.45e-19
C156 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.0622f
C157 CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_3_mag_1.JK_FF_mag_1.K 0.00761f
C158 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK 0.00302f
C159 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.Q3 0.076f
C160 a_16634_13026# CLK_DIV_11_mag_new_0.Q0 0.069f
C161 a_10096_15189# CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 1.32e-19
C162 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 2.25e-21
C163 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.103f
C164 CLK CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 4.05e-20
C165 a_4404_10895# VDD 3.14e-19
C166 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.Q1 0.0161f
C167 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_DIV_11_mag_new_0.and2_mag_3.IN1 2.29e-19
C168 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.and2_mag_3.IN1 2.11e-19
C169 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.28f
C170 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.K 0.69f
C171 a_11497_10895# CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 5.54e-20
C172 a_8703_9798# CLK_div_3_mag_0.JK_FF_mag_1.QB 0.00392f
C173 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN VDD 0.411f
C174 a_8139_9798# RST 1.8e-19
C175 CLK_div_3_mag_1.Q0 CLK 0.149f
C176 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT RST 0.313f
C177 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD 0.397f
C178 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.122f
C179 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00183f
C180 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 0.36f
C181 a_12215_9798# CLK_div_3_mag_1.JK_FF_mag_1.QB 1.86e-20
C182 a_8503_11887# CLK_DIV_11_mag_new_0.Q2 0.00335f
C183 a_9797_13028# VDD 3.14e-19
C184 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0622f
C185 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK 0.298f
C186 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.Q0 8.04e-19
C187 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.Q0 0.0485f
C188 CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_DIV_11_mag_new_0.Q1 3.8e-20
C189 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.Q0 1.09e-20
C190 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.0707f
C191 CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_DIV_11_mag_new_0.Q1 0.209f
C192 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.Q2 4.54f
C193 a_7380_11933# CLK_DIV_11_mag_new_0.Q3 0.0157f
C194 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_0.Q0 0.0635f
C195 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 8.16e-20
C196 CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_DIV_11_mag_new_0.Q0 0.0128f
C197 CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 6.36e-20
C198 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 8.28e-20
C199 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 9.07e-20
C200 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_8869_10895# 1.17e-20
C201 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.Q3 8.83e-19
C202 CLK RST 0.0349f
C203 a_3840_10895# VDD 3.14e-19
C204 CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.Q3 0.299f
C205 CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_DIV_11_mag_new_0.Q0 0.00187f
C206 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN VDD 0.517f
C207 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 VDD 9.72f
C208 a_8139_9798# CLK_div_3_mag_0.JK_FF_mag_1.QB 3.33e-19
C209 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.0598f
C210 a_3556_12901# VDD 0.167f
C211 a_3556_12901# CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 0.132f
C212 a_7575_9798# RST 7.58e-19
C213 a_12055_9798# CLK_div_3_mag_1.JK_FF_mag_1.QB 1.41e-20
C214 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.122f
C215 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT RST 5.36e-20
C216 a_9233_13028# VDD 3.14e-19
C217 a_15500_11885# VDD 2.21e-19
C218 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 8.26e-20
C219 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 3.18e-19
C220 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.Q1 3.7f
C221 a_15500_11885# a_15660_11885# 0.0504f
C222 CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN a_3994_15139# 2.7e-20
C223 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 1.53e-19
C224 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.Q3 9.8e-20
C225 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.122f
C226 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_8709_10895# 1.5e-20
C227 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 RST 0.194f
C228 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.Q0 2.42f
C229 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 0.321f
C230 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 1.2e-19
C231 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.Q2 2.07e-20
C232 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 1.93f
C233 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.0881f
C234 a_8863_9798# CLK_div_3_mag_0.JK_FF_mag_1.K 8.64e-19
C235 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.Q3 0.00154f
C236 a_7011_9798# RST 7.24e-19
C237 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.16f
C238 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.122f
C239 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00158f
C240 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_13944_9798# 0.069f
C241 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 0.777f
C242 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_1.JK_FF_mag_1.K 8.58e-20
C243 a_14936_11885# VDD 7.37e-19
C244 CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 VDD 0.515f
C245 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 1.89e-20
C246 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.Q2 1.5e-19
C247 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_1.Q0 0.0343f
C248 CLK_div_3_mag_1.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00101f
C249 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 4.52e-20
C250 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.nand3_mag_1.OUT 9.75e-21
C251 CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.Q1 0.0409f
C252 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_1.QB 0.175f
C253 CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 a_2597_12515# 4.44e-20
C254 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_6662_13030# 4.52e-20
C255 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.Q2 0.306f
C256 a_13698_15251# a_13858_15251# 0.186f
C257 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_DIV_11_mag_new_0.Q3 0.0127f
C258 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_8145_10895# 0.0203f
C259 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 1.49e-19
C260 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.Q0 0.00123f
C261 a_10363_9798# CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 4.52e-20
C262 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.0894f
C263 a_15238_10895# CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.0202f
C264 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.159f
C265 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.Q3 0.11f
C266 CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.Q0 0.242f
C267 a_2757_14017# CLK_DIV_11_mag_new_0.Q3 6.63e-20
C268 CLK_div_3_mag_1.or_2_mag_0.IN2 VDD 0.492f
C269 a_7011_9798# CLK_div_3_mag_0.JK_FF_mag_1.QB 0.0112f
C270 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_13380_9798# 0.00372f
C271 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT RST 0.306f
C272 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 0.104f
C273 RST CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.0917f
C274 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 6.71e-19
C275 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 RST 0.186f
C276 a_8509_12984# VDD 2.21e-19
C277 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0894f
C278 CLK_div_3_mag_1.JK_FF_mag_1.QB a_14514_10895# 0.00695f
C279 a_14776_11885# VDD 9.58e-19
C280 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.124f
C281 CLK_DIV_11_mag_new_0.Q2 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.101f
C282 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_6816_11933# 0.0036f
C283 CLK_div_3_mag_1.Q0 RST 0.354f
C284 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.195f
C285 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK 1.31f
C286 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.Q2 6.62e-20
C287 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.Q1 0.117f
C288 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_6098_13030# 0.0195f
C289 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_7985_10895# 0.0733f
C290 a_2757_14017# CLK_DIV_11_mag_new_0.Q2 8.95e-19
C291 a_5686_9798# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00119f
C292 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.109f
C293 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 1.5e-20
C294 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 3.34e-19
C295 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C296 a_15078_10895# CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.0731f
C297 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD 0.647f
C298 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 0.122f
C299 a_2597_14017# CLK_DIV_11_mag_new_0.Q3 4.15e-19
C300 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 2.76e-19
C301 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 0.321f
C302 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.Q0 0.305f
C303 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 4.44e-20
C304 a_7226_13030# VDD 3.56e-19
C305 CLK_div_3_mag_1.JK_FF_mag_1.QB a_14354_10895# 0.00696f
C306 a_12055_9798# CLK_div_3_mag_1.JK_FF_mag_1.K 0.00392f
C307 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.Q3 0.0281f
C308 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 3.34e-19
C309 a_13629_11933# VDD 3.14e-19
C310 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.321f
C311 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.and2_mag_3.OUT 2.6e-20
C312 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_DIV_11_mag_new_0.Q1 7.38e-19
C313 CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT 0.163f
C314 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.Q3 1.4e-20
C315 CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 0.209f
C316 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0894f
C317 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.231f
C318 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.109f
C319 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.Q1 1.32e-19
C320 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.nand3_mag_1.OUT 1.32e-19
C321 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT RST 0.00437f
C322 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K a_5374_12986# 0.00472f
C323 a_2757_14017# CLK_DIV_11_mag_new_0.Q1 1.75e-19
C324 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_7421_10895# 0.00378f
C325 a_4437_8231# CLK_div_3_mag_0.JK_FF_mag_1.K 0.00168f
C326 a_5122_9798# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.43e-19
C327 CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00776f
C328 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.Q0 0.00425f
C329 a_14514_10895# CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 9.1e-19
C330 a_10806_8231# CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 1.4e-19
C331 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.Q2 0.00952f
C332 CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.Q3 1.34e-19
C333 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.Q0 2.13e-20
C334 CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 1.48e-19
C335 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 9.8e-19
C336 a_2757_14017# CLK_DIV_11_mag_new_0.Q0 0.0177f
C337 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.765f
C338 CLK_div_3_mag_0.JK_FF_mag_1.QB RST 0.761f
C339 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.Q2 0.0766f
C340 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_3994_9798# 0.00372f
C341 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C342 a_6662_13030# VDD 3.14e-19
C343 a_13629_11933# CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.0811f
C344 CLK_div_3_mag_1.JK_FF_mag_1.QB a_13790_10895# 0.00964f
C345 a_11491_9798# CLK_div_3_mag_1.JK_FF_mag_1.K 1.75e-19
C346 a_13065_11933# VDD 3.14e-19
C347 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 2.12e-19
C348 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK 7.03e-21
C349 a_8509_12984# a_8669_12984# 0.0504f
C350 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VDD 0.739f
C351 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.Q0 0.338f
C352 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT 0.00134f
C353 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_16224_11929# 0.0036f
C354 a_14776_11885# a_14936_11885# 0.0504f
C355 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 VDD 0.4f
C356 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.Q2 0.0274f
C357 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.QB 2.81e-20
C358 CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 7.08e-20
C359 a_2597_14017# CLK_DIV_11_mag_new_0.Q1 0.00369f
C360 a_4558_9798# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.011f
C361 CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.Q2 0.0515f
C362 a_14354_10895# CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 2.88e-20
C363 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.105f
C364 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.Q1 0.00367f
C365 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.QB 7.49e-20
C366 a_4002_14308# CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN 0.069f
C367 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT VDD 0.644f
C368 a_2597_14017# CLK_DIV_11_mag_new_0.Q0 0.00765f
C369 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.Q1 0.0365f
C370 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_5852_10895# 1.17e-20
C371 a_3994_15139# CLK_DIV_11_mag_new_0.Q2 0.00186f
C372 a_6098_13030# VDD 3.14e-19
C373 a_10927_9798# CLK_div_3_mag_1.JK_FF_mag_1.K 2.96e-19
C374 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 VDD 1.16f
C375 a_13065_11933# CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.00964f
C376 CLK_div_3_mag_1.JK_FF_mag_1.QB a_13226_10895# 0.0811f
C377 a_10773_10895# CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.069f
C378 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.Q0 0.0175f
C379 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT a_15660_11885# 2.88e-20
C380 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 3.43e-19
C381 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_5528_11889# 8.66e-20
C382 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 4.04e-19
C383 CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT CLK_DIV_11_mag_new_0.and2_mag_3.IN1 0.00147f
C384 a_13380_9798# CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 4.52e-20
C385 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.0854f
C386 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.Q0 0.0582f
C387 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.233f
C388 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.28f
C389 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_13475_13030# 0.00118f
C390 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C391 a_12215_9798# VDD 2.21e-19
C392 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD 0.398f
C393 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.Q0 0.0635f
C394 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.Q1 0.00917f
C395 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 2.01e-19
C396 CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.Q1 0.0248f
C397 a_5466_15136# CLK_DIV_11_mag_new_0.Q2 0.0115f
C398 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_7575_9798# 0.069f
C399 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 1.47e-20
C400 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.Q0 0.0187f
C401 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 RST 0.132f
C402 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 5.25e-20
C403 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_16634_13026# 0.0114f
C404 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_5692_10895# 1.5e-20
C405 a_3994_15139# CLK_DIV_11_mag_new_0.Q1 0.0186f
C406 CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.Q0 0.0072f
C407 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 1.1e-19
C408 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN a_5534_12986# 1.03e-20
C409 a_10363_9798# CLK_div_3_mag_1.JK_FF_mag_1.K 0.012f
C410 a_12501_11889# CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.00696f
C411 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 3.98e-19
C412 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 1.32e-21
C413 a_12341_11889# VDD 2.77e-19
C414 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT a_15500_11885# 9.1e-19
C415 a_10209_10895# CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.00372f
C416 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 6.02e-20
C417 a_16634_13026# CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 0.00372f
C418 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD 1f
C419 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN VDD 0.434f
C420 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 7.55e-19
C421 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_1.Q0 0.0463f
C422 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.Q1 1.31e-20
C423 RST CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0319f
C424 a_3994_15139# CLK_DIV_11_mag_new_0.Q0 0.00718f
C425 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_12911_13030# 0.011f
C426 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 a_10361_13028# 0.00372f
C427 a_15238_10895# VDD 0.0132f
C428 CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT VDD 0.573f
C429 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C430 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT a_15506_13026# 0.00378f
C431 Vdiv99 CLK_DIV_11_mag_new_0.Q3 0.00382f
C432 a_5466_15136# CLK_DIV_11_mag_new_0.Q1 0.015f
C433 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_7011_9798# 0.00372f
C434 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.105f
C435 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 2.51e-19
C436 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 0.139f
C437 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_1.Q0 0.209f
C438 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.00808f
C439 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_5128_10895# 0.0203f
C440 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_16070_13026# 2.96e-19
C441 a_12341_11889# CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.00695f
C442 a_5466_15136# CLK_DIV_11_mag_new_0.Q0 0.00589f
C443 CLK CLK_DIV_11_mag_new_0.Q1 0.00343f
C444 CLK_div_3_mag_0.JK_FF_mag_1.K RST 0.272f
C445 a_5374_12986# VDD 2.21e-19
C446 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN a_5374_12986# 1.29e-20
C447 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.133f
C448 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT a_14936_11885# 0.0731f
C449 a_16070_13026# CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 0.069f
C450 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK 0.00254f
C451 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN a_3556_12901# 1.14e-19
C452 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT a_9387_11887# 2.88e-20
C453 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD 0.397f
C454 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 1.99e-20
C455 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_14936_11885# 1.46e-19
C456 CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 0.116f
C457 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT 1.2e-19
C458 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_12347_13030# 1.43e-19
C459 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 0.122f
C460 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 2.46e-20
C461 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.Q1 0.00101f
C462 a_15078_10895# VDD 0.00888f
C463 CLK CLK_DIV_11_mag_new_0.Q0 6.19e-21
C464 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 a_9797_13028# 0.069f
C465 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 6.02e-20
C466 a_11491_9798# VDD 3.14e-19
C467 CLK_div_3_mag_1.JK_FF_mag_1.K a_11497_10895# 0.00695f
C468 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.69f
C469 a_13858_15251# CLK_DIV_11_mag_new_0.Q3 0.0504f
C470 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.K 0.352f
C471 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 1.99e-20
C472 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT a_14942_12982# 0.0732f
C473 a_14782_12982# CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.00472f
C474 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.0106f
C475 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_8709_10895# 1.46e-19
C476 a_10096_15189# a_10256_15189# 0.0504f
C477 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.00584f
C478 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.121f
C479 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT RST 1.99e-21
C480 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 1.74e-19
C481 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.Q0 3.4e-19
C482 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 VDD 0.395f
C483 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.313f
C484 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.QB 3.28e-19
C485 RST a_6816_11933# 0.00192f
C486 CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 4.95e-20
C487 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_4968_10895# 0.0733f
C488 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 6.93e-19
C489 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT a_14776_11885# 0.0202f
C490 a_11617_11889# VDD 2.21e-19
C491 RST CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 0.265f
C492 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 6.18e-19
C493 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT a_9227_11887# 9.1e-19
C494 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_9951_11931# 0.00378f
C495 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 5.32e-19
C496 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_11783_12986# 0.00119f
C497 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT RST 5.45e-20
C498 a_10927_9798# VDD 3.14e-19
C499 a_14514_10895# VDD 0.0012f
C500 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.Q2 4.01e-20
C501 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 a_10361_13028# 4.52e-20
C502 CLK_div_3_mag_1.JK_FF_mag_1.K a_11337_10895# 0.00696f
C503 a_13698_15251# CLK_DIV_11_mag_new_0.Q3 0.0186f
C504 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 a_15506_13026# 0.0697f
C505 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT a_14782_12982# 0.0203f
C506 CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 1.5e-20
C507 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K VDD 0.9f
C508 CLK_div_3_mag_1.Q0 CLK_DIV_11_mag_new_0.Q2 0.0327f
C509 a_2590_14702# CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN 0.069f
C510 RST CLK_DIV_11_mag_new_0.Q3 0.22f
C511 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 5.74e-20
C512 a_12221_10895# VDD 0.00743f
C513 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.99e-19
C514 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 7.36e-21
C515 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 RST 0.00218f
C516 RST a_6252_11889# 0.00341f
C517 a_3994_9798# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 4.52e-20
C518 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_4404_10895# 0.00378f
C519 a_10515_11931# VDD 3.14e-19
C520 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT 0.342f
C521 a_8869_10895# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.0202f
C522 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT a_8663_11887# 0.0731f
C523 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD 0.392f
C524 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 2.8e-19
C525 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD 0.995f
C526 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_9387_11887# 0.0733f
C527 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.Q1 0.00403f
C528 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.Q1 0.338f
C529 a_10363_9798# VDD 3.56e-19
C530 a_14354_10895# VDD 9.82e-19
C531 RST CLK_DIV_11_mag_new_0.Q2 0.187f
C532 CLK_div_3_mag_1.JK_FF_mag_1.K a_10773_10895# 0.00964f
C533 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.0998f
C534 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C535 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 2.19f
C536 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_3_mag_1.Q0 3.45e-19
C537 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.Q3 2.95e-20
C538 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 0.00265f
C539 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 RST 0.188f
C540 CLK_div_3_mag_1.Q0 CLK_DIV_11_mag_new_0.Q1 0.00948f
C541 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 5.87e-19
C542 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 8.16e-20
C543 a_12061_10895# VDD 0.00305f
C544 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.Q0 3.56e-19
C545 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.QB 0.0576f
C546 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.Q0 0.00335f
C547 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q2 0.0549f
C548 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 3.25e-20
C549 a_5846_9798# RST 7.78e-19
C550 RST a_6092_11889# 0.0024f
C551 a_4437_8231# CLK_div_3_mag_0.Q0 0.0134f
C552 a_9951_11931# VDD 3.14e-19
C553 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0622f
C554 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD 0.468f
C555 a_4404_10895# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.069f
C556 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 3.6e-21
C557 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT a_8503_11887# 0.0202f
C558 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.25f
C559 a_8709_10895# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.0731f
C560 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_9227_11887# 0.0203f
C561 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT VDD 0.643f
C562 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 0.205f
C563 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 RST 0.187f
C564 a_5846_9798# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0203f
C565 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB RST 0.296f
C566 RST CLK_DIV_11_mag_new_0.Q1 0.164f
C567 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD 0.391f
C568 a_13790_10895# VDD 0.00149f
C569 CLK_div_3_mag_1.JK_FF_mag_1.K a_10209_10895# 0.0811f
C570 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_7421_10895# 0.0036f
C571 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 RST 0.155f
C572 CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q3 0.299f
C573 a_5846_9798# CLK_div_3_mag_0.JK_FF_mag_1.QB 1.86e-20
C574 a_11497_10895# VDD 2.21e-19
C575 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VDD 1.08f
C576 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q1 0.316f
C577 RST CLK_DIV_11_mag_new_0.Q0 0.0664f
C578 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.231f
C579 CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 0.129f
C580 a_5686_9798# RST 6.43e-19
C581 RST a_5528_11889# 0.00139f
C582 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 2.34e-19
C583 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 0.0404f
C584 a_5852_10895# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0202f
C585 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00118f
C586 a_3840_10895# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.00372f
C587 a_8145_10895# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 9.1e-19
C588 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 VDD 1.17f
C589 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 0.36f
C590 a_10961_15230# CLK_DIV_11_mag_new_0.Q1 0.015f
C591 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_8663_11887# 1.5e-20
C592 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 a_6816_11933# 0.069f
C593 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0622f
C594 a_3994_15139# CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 0.0202f
C595 a_2597_12515# VDD 3.14e-19
C596 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 0.109f
C597 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q0 0.107f
C598 CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q2 9.25e-19
C599 CLK_div_3_mag_1.or_2_mag_0.IN2 a_10927_9798# 4.9e-20
C600 a_5686_9798# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0732f
C601 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 1.14e-19
C602 a_13226_10895# VDD 0.00149f
C603 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.105f
C604 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.00154f
C605 CLK_div_3_mag_1.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.00477f
C606 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K a_8509_12984# 0.00472f
C607 a_5686_9798# CLK_div_3_mag_0.JK_FF_mag_1.QB 1.41e-20
C608 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 5.2e-20
C609 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 7.86e-19
C610 a_4002_14308# CLK_DIV_11_mag_new_0.Q1 0.0205f
C611 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 4.11e-19
C612 a_5122_9798# RST 2.97e-19
C613 RST a_5368_11889# 0.00125f
C614 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.Q3 0.0635f
C615 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK 0.272f
C616 a_5692_10895# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0731f
C617 a_9227_11887# VDD 2.21e-19
C618 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.306f
C619 a_7985_10895# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 2.88e-20
C620 a_10256_15189# CLK_DIV_11_mag_new_0.Q1 5.19e-20
C621 Vdiv99 CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT 0.121f
C622 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_8503_11887# 1.17e-20
C623 a_4002_14308# CLK_DIV_11_mag_new_0.Q0 0.00379f
C624 a_16634_13026# VDD 3.56e-19
C625 CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q1 0.146f
C626 CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_DIV_11_mag_new_0.and2_mag_3.IN1 0.012f
C627 a_5122_9798# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00378f
C628 a_12341_11889# a_12501_11889# 0.0504f
C629 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 9.58e-20
C630 a_2590_14702# CLK_DIV_11_mag_new_0.Q3 0.00572f
C631 RST CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.0794f
C632 a_10256_15189# CLK_DIV_11_mag_new_0.Q0 0.0121f
C633 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00169f
C634 CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q0 0.00525f
C635 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 VDD 1.32f
C636 a_10773_10895# VDD 3.14e-19
C637 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.K 8.58e-20
C638 a_4558_9798# RST 2.24e-19
C639 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 0.198f
C640 a_12055_9798# a_12215_9798# 0.0504f
C641 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.00253f
C642 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_5692_10895# 1.46e-19
C643 CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 0.048f
C644 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 8.16e-20
C645 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN a_10806_8231# 3.25e-19
C646 a_8663_11887# VDD 7.34e-19
C647 CLK_div_3_mag_0.or_2_mag_0.IN2 a_4437_8231# 8.64e-19
C648 a_5128_10895# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 9.1e-19
C649 a_13858_15251# CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT 0.198f
C650 CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 VDD 0.378f
C651 CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 0.226f
C652 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VDD 1f
C653 a_10096_15189# CLK_DIV_11_mag_new_0.Q1 3.35e-20
C654 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.121f
C655 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.768f
C656 a_10961_15230# CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 2.5e-19
C657 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.and2_mag_3.IN1 0.00243f
C658 a_16070_13026# VDD 3.14e-19
C659 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.Q1 7.75e-19
C660 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 8.59e-20
C661 CLK_DIV_11_mag_new_0.and2_mag_3.OUT VDD 0.304f
C662 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.and2_mag_3.OUT 3.83e-19
C663 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.Q3 0.00107f
C664 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_11617_11889# 5.54e-20
C665 RST CLK_div_3_mag_0.Q0 0.0893f
C666 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.233f
C667 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00166f
C668 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 7.63e-19
C669 a_4437_8231# CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.132f
C670 a_10096_15189# CLK_DIV_11_mag_new_0.Q0 0.00747f
C671 a_6816_11933# CLK_DIV_11_mag_new_0.Q3 0.00859f
C672 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.211f
C673 CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 5.32e-19
C674 a_10209_10895# VDD 3.14e-19
C675 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.Q0 7.24e-19
C676 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_1.QB 0.215f
C677 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_1.JK_FF_mag_1.K 0.0725f
C678 a_4968_10895# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 2.88e-20
C679 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN a_11779_8699# 0.069f
C680 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.Q2 8.93e-19
C681 a_12221_10895# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.0202f
C682 a_8503_11887# VDD 9.56e-19
C683 a_2590_14702# CLK_DIV_11_mag_new_0.Q1 0.00544f
C684 a_5374_12986# a_5534_12986# 0.0504f
C685 a_13698_15251# CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT 0.0135f
C686 CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 a_3556_12901# 0.0178f
C687 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT RST 0.285f
C688 CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 0.0022f
C689 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K VDD 0.833f
C690 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 0.122f
C691 CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 1.64e-20
C692 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.00165f
C693 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.0622f
C694 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 1.83e-19
C695 CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.and2_mag_3.IN1 0.407f
C696 a_6252_11889# CLK_DIV_11_mag_new_0.Q3 0.0101f
C697 a_15232_9798# CLK 0.0101f
C698 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_1.Q0 7.24e-19
C699 CLK_div_3_mag_1.JK_FF_mag_1.QB CLK 0.362f
C700 CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 RST 7.55e-19
C701 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.Q2 9.75e-19
C702 a_3994_9798# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00118f
C703 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 1.05e-20
C704 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK 1.69e-20
C705 a_5686_9798# CLK_div_3_mag_0.JK_FF_mag_1.K 0.00392f
C706 a_8669_12984# CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 1.24e-20
C707 a_15078_10895# a_15238_10895# 0.0504f
C708 a_8863_9798# CLK_div_3_mag_1.JK_FF_mag_1.K 1.09e-20
C709 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C710 a_11779_8699# CLK 0.0103f
C711 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 0.00574f
C712 a_7380_11933# VDD 3.14e-19
C713 CLK_DIV_11_mag_new_0.Q2 CLK_DIV_11_mag_new_0.Q3 1.19f
C714 a_12061_10895# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.0731f
C715 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 1.89e-19
C716 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.507f
C717 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT VDD 0.647f
C718 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0502f
C719 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD 0.739f
C720 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.Q3 0.00397f
C721 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 2.98e-19
C722 CLK_DIV_11_mag_new_0.nand3_mag_1.OUT VDD 1.19f
C723 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT RST 0.00543f
C724 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 a_6252_11889# 8.64e-19
C725 CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 0.191f
C726 a_15072_9798# CLK 0.00939f
C727 a_6092_11889# CLK_DIV_11_mag_new_0.Q3 0.0102f
C728 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00118f
C729 RST a_15506_13026# 2.67e-19
C730 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.122f
C731 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 0.342f
C732 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.121f
C733 CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.0147f
C734 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.122f
C735 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00975f
C736 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.Q1 1.17e-19
C737 a_6092_11889# a_6252_11889# 0.0504f
C738 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD 0.802f
C739 a_5122_9798# CLK_div_3_mag_0.JK_FF_mag_1.K 1.75e-19
C740 a_8509_12984# CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 1.59e-20
C741 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.Q0 0.0349f
C742 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_4404_10895# 0.0036f
C743 a_14508_9798# CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.0202f
C744 a_8703_9798# CLK_div_3_mag_1.JK_FF_mag_1.K 8.77e-21
C745 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.Q3 9.05e-22
C746 a_11497_10895# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 9.1e-19
C747 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.Q2 1.12e-19
C748 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 2.39e-20
C749 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 9.52e-19
C750 CLK_DIV_11_mag_new_0.Q1 CLK_DIV_11_mag_new_0.Q3 1.83f
C751 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_1.Q0 0.0635f
C752 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.Q0 3.38e-19
C753 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.K 1.33e-19
C754 CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.111f
C755 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VDD 1.08f
C756 RST CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 0.0294f
C757 a_11617_11889# a_11777_11889# 0.0504f
C758 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 2.67e-20
C759 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C760 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_DIV_11_mag_new_0.nand3_mag_1.OUT 9.5e-19
C761 CLK CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.235f
C762 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.nand3_mag_1.OUT 4.78e-20
C763 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_13065_11933# 0.0036f
C764 CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.Q3 0.128f
C765 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 1.82e-19
C766 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT VDD 0.664f
C767 a_14508_9798# CLK 6.43e-21
C768 a_5528_11889# CLK_DIV_11_mag_new_0.Q3 0.0152f
C769 RST a_14942_12982# 7.84e-19
C770 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_1.JK_FF_mag_1.K 0.00384f
C771 a_10806_8231# CLK_div_3_mag_1.Q0 0.0134f
C772 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.Q2 0.00391f
C773 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.Q2 1.97f
C774 CLK_DIV_11_mag_new_0.Q2 CLK_DIV_11_mag_new_0.Q1 2.34f
C775 a_4558_9798# CLK_div_3_mag_0.JK_FF_mag_1.K 2.96e-19
C776 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 RST 0.0222f
C777 a_13944_9798# CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 4.52e-20
C778 a_7226_13030# CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.0114f
C779 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 8.16e-20
C780 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 9.62e-20
C781 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.Q1 1.86e-19
C782 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0854f
C783 a_4002_14308# CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 1.78e-20
C784 a_8869_10895# CLK_div_3_mag_1.Q0 1.38e-20
C785 a_11337_10895# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 2.88e-20
C786 a_7011_9798# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 4.52e-20
C787 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 2.01e-19
C788 CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.Q2 0.888f
C789 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_6857_10895# 2.34e-20
C790 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VDD 0.523f
C791 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD 0.66f
C792 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 a_16788_11929# 0.00372f
C793 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.00166f
C794 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VDD 0.398f
C795 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.Q0 2.37f
C796 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_15232_9798# 0.0203f
C797 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD 0.397f
C798 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 a_15660_11885# 8.64e-19
C799 CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 0.124f
C800 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 8.16e-20
C801 a_14776_11885# CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 8.64e-19
C802 a_14508_9798# CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.0697f
C803 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_1.JK_FF_mag_1.QB 0.343f
C804 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT a_12347_13030# 0.00378f
C805 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.16f
C806 a_13944_9798# CLK 6.06e-21
C807 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0377f
C808 a_5368_11889# CLK_DIV_11_mag_new_0.Q3 0.0124f
C809 a_5686_9798# a_5846_9798# 0.0504f
C810 RST a_14782_12982# 9.41e-19
C811 CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 CLK_DIV_11_mag_new_0.nand3_mag_1.OUT 1.03e-19
C812 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.Q1 6.01e-19
C813 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.Q1 1.17e-19
C814 CLK_div_3_mag_1.JK_FF_mag_1.K CLK 2.11f
C815 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 2e-19
C816 a_8869_10895# RST 0.00466f
C817 a_6662_13030# CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 2.96e-19
C818 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.Q0 3.53e-19
C819 a_8139_9798# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0697f
C820 a_8709_10895# CLK_div_3_mag_1.Q0 1.09e-20
C821 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.Q0 0.00121f
C822 CLK_div_3_mag_1.JK_FF_mag_1.QB RST 0.592f
C823 CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.Q1 3.23f
C824 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.Q3 0.0683f
C825 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB RST 0.141f
C826 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 1.74e-19
C827 a_12055_9798# CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.00119f
C828 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 a_16224_11929# 0.069f
C829 a_8863_9798# VDD 5.99e-19
C830 a_16634_13026# CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00118f
C831 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 6.23e-19
C832 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_15072_9798# 0.0732f
C833 a_13629_11933# CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 2.75e-21
C834 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN a_2597_12515# 0.069f
C835 a_13944_9798# CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.0059f
C836 a_2597_14017# VDD 2.21e-19
C837 a_13380_9798# CLK 9.45e-19
C838 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 a_12911_13030# 0.0059f
C839 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT a_11783_12986# 0.0732f
C840 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_10361_13028# 0.00118f
C841 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 8.58e-20
C842 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.Q2 0.291f
C843 a_8709_10895# RST 0.00464f
C844 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 VDD 1.15f
C845 a_14354_10895# a_14514_10895# 0.0504f
C846 a_6098_13030# CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 3.33e-19
C847 a_7575_9798# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0059f
C848 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN VDD 0.409f
C849 CLK_div_3_mag_0.Q0 CLK_DIV_11_mag_new_0.Q3 0.0506f
C850 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 1.31e-20
C851 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 2.01e-19
C852 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD 0.391f
C853 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 RST 0.067f
C854 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_13790_10895# 0.069f
C855 a_11491_9798# CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 1.43e-19
C856 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.00183f
C857 a_8703_9798# VDD 2.65e-19
C858 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_11777_11889# 1.46e-19
C859 a_16070_13026# CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.011f
C860 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 a_10515_11931# 0.00372f
C861 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_14508_9798# 0.00378f
C862 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 VDD 1.18f
C863 a_13065_11933# CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 5.58e-22
C864 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 a_12347_13030# 0.0697f
C865 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT a_11623_12986# 0.0203f
C866 CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN VDD 0.41f
C867 a_12061_10895# a_12221_10895# 0.0504f
C868 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_9797_13028# 0.011f
C869 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00183f
C870 a_5368_11889# a_5528_11889# 0.0504f
C871 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.0306f
C872 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.00254f
C873 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.00916f
C874 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT RST 0.0568f
C875 a_8145_10895# RST 0.00311f
C876 CLK_div_3_mag_0.Q0 CLK_DIV_11_mag_new_0.Q2 6.41e-20
C877 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.Q1 1.93f
C878 a_5534_12986# CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.00392f
C879 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 9.22e-20
C880 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 2.15e-20
C881 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 1.31e-20
C882 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 1.21e-19
C883 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN VDD 0.468f
C884 a_3994_15139# VDD 0.165f
C885 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_1.K 0.23f
C886 CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT CLK_DIV_11_mag_new_0.Q3 0.257f
C887 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.QB 0.175f
C888 a_5852_10895# RST 0.00549f
C889 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.Q0 1.76f
C890 a_10927_9798# CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.011f
C891 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_13226_10895# 0.00372f
C892 CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 3.81e-19
C893 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.105f
C894 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VDD 1f
C895 a_8139_9798# VDD 3.14e-19
C896 CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 CLK_DIV_11_mag_new_0.Q3 8.02e-19
C897 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.0231f
C898 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 a_9951_11931# 0.069f
C899 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.Q0 2.37f
C900 CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 0.126f
C901 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.JK_FF_mag_1.K 0.00761f
C902 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.159f
C903 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 6.11e-19
C904 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.0715f
C905 RST CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.092f
C906 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_1.JK_FF_mag_1.K 0.0948f
C907 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.211f
C908 RST a_12347_13030# 3.68e-20
C909 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_9233_13028# 1.43e-19
C910 a_5466_15136# VDD 0.165f
C911 CLK_div_3_mag_0.JK_FF_mag_1.QB a_8145_10895# 0.00695f
C912 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_15506_13026# 0.0195f
C913 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.122f
C914 a_7985_10895# RST 0.00359f
C915 CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT 0.00982f
C916 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.QB 0.21f
C917 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K RST 0.0105f
C918 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.JK_FF_mag_1.K 0.00205f
C919 a_4437_8231# VDD 0.165f
C920 a_13944_9798# RST 3.62e-19
C921 CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 CLK_DIV_11_mag_new_0.Q2 0.149f
C922 CLK VDD 2.4f
C923 CLK_div_3_mag_1.JK_FF_mag_1.K RST 0.432f
C924 a_5692_10895# RST 0.00513f
C925 a_5686_9798# CLK_div_3_mag_0.Q0 2.79e-20
C926 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 4.23e-20
C927 a_10363_9798# CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.00118f
C928 a_5528_11889# CLK_div_3_mag_0.Q0 6.19e-21
C929 a_7575_9798# VDD 3.14e-19
C930 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT 0.00183f
C931 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 4.68e-20
C932 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 4.44e-20
C933 CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_DIV_11_mag_new_0.Q3 0.0145f
C934 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT VDD 0.647f
C935 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0894f
C936 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_5466_15136# 0.0131f
C937 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.Q1 0.0346f
C938 a_12061_10895# CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 1.46e-19
C939 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_8669_12984# 0.00119f
C940 RST CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.147f
C941 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 a_7226_13030# 0.00372f
C942 CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT CLK_DIV_11_mag_new_0.Q1 3.11e-19
C943 CLK_div_3_mag_0.JK_FF_mag_1.QB a_7985_10895# 0.00696f
C944 a_7421_10895# RST 0.00439f
C945 a_15072_9798# CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.00119f
C946 CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 1.89e-19
C947 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT RST 0.281f
C948 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN a_10806_8231# 0.132f
C949 CLK CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 5.14e-20
C950 CLK_div_3_mag_0.or_2_mag_0.IN2 a_5410_8699# 7.48e-20
C951 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.Q0 3.94e-19
C952 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 VDD 0.655f
C953 a_13380_9798# RST 7.24e-19
C954 CLK_DIV_11_mag_new_0.Q2 CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 0.026f
C955 CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 CLK_DIV_11_mag_new_0.Q1 0.00103f
C956 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.122f
C957 CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT CLK_DIV_11_mag_new_0.Q0 6.99e-20
C958 a_5128_10895# RST 0.00211f
C959 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 RST 0.205f
C960 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_8863_9798# 0.0203f
C961 Vdiv99 VDD 0.189f
C962 a_7011_9798# VDD 3.56e-19
C963 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.343f
C964 CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 CLK_DIV_11_mag_new_0.Q0 0.0444f
C965 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.412f
C966 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 2.39e-19
C967 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT RST 0.286f
C968 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.00118f
C969 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 8.26e-20
C970 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 a_6662_13030# 0.069f
C971 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.36f
C972 a_10961_15230# CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 0.069f
C973 CLK_div_3_mag_0.JK_FF_mag_1.QB a_7421_10895# 0.00964f
C974 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.QB 1.21e-19
C975 a_14508_9798# CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 1.43e-19
C976 a_6857_10895# RST 0.00379f
C977 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 1.9e-20
C978 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_7226_13030# 0.00118f
C979 CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.124f
C980 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.122f
C981 CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT CLK_DIV_11_mag_new_0.nand3_mag_1.OUT 0.131f
C982 a_3994_9798# RST 2.24e-19
C983 CLK_DIV_11_mag_new_0.Q1 CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 0.203f
C984 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0147f
C985 Vdiv99 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 1.71e-21
C986 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.121f
C987 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.Q2 1.83e-19
C988 a_4968_10895# RST 0.0019f
C989 a_13858_15251# VDD 0.0418f
C990 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_8703_9798# 0.0732f
C991 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 0.249f
C992 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00156f
C993 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD 0.995f
C994 CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 0.205f
C995 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD 0.651f
C996 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 0.109f
C997 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT VDD 0.642f
C998 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.24f
C999 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 0.00975f
C1000 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.Q1 0.0635f
C1001 a_11337_10895# a_11497_10895# 0.0504f
C1002 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.00188f
C1003 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_13226_10895# 2.58e-20
C1004 CLK_div_3_mag_1.Q0 VDD 1.3f
C1005 a_10256_15189# CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 4.43e-21
C1006 CLK_div_3_mag_0.JK_FF_mag_1.QB a_6857_10895# 0.0811f
C1007 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K a_8503_11887# 8.64e-19
C1008 a_13944_9798# CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.011f
C1009 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 9.87e-20
C1010 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VDD 0.647f
C1011 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.Q0 1.71e-21
C1012 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.0718f
C1013 CLK_div_3_mag_1.or_2_mag_0.IN2 CLK 6.62e-20
C1014 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_6662_13030# 0.011f
C1015 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.00238f
C1016 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.103f
C1017 a_13858_15251# CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 2.31e-19
C1018 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 5.25e-20
C1019 a_10961_15230# CLK_DIV_11_mag_new_0.and2_mag_3.IN1 0.00476f
C1020 a_13858_15251# CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 1.9e-19
C1021 a_13698_15251# VDD 0.235f
C1022 a_4404_10895# RST 7.06e-19
C1023 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_8139_9798# 0.00378f
C1024 a_9227_11887# a_9387_11887# 0.0504f
C1025 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.0385f
C1026 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.103f
C1027 a_14942_12982# CLK_DIV_11_mag_new_0.Q0 2.79e-20
C1028 RST VDD 2.62f
C1029 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 RST 1.36e-19
C1030 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN RST 0.00236f
C1031 a_10773_10895# CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.0036f
C1032 CLK_div_3_mag_1.Q0 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 8.39e-21
C1033 RST a_15660_11885# 0.00162f
C1034 a_10096_15189# CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 3.44e-21
C1035 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K a_7380_11933# 1.44e-21
C1036 a_13380_9798# CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.00118f
C1037 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN VDD 0.423f
C1038 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 1.84e-19
C1039 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD 0.647f
C1040 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_div_3_mag_0.JK_FF_mag_1.K 3.78e-20
C1041 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.Q3 9.8e-20
C1042 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_6098_13030# 1.43e-19
C1043 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 8.59e-20
C1044 a_13698_15251# CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 3.59e-19
C1045 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.K 8.36e-19
C1046 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 2.75e-19
C1047 a_10256_15189# CLK_DIV_11_mag_new_0.and2_mag_3.IN1 0.00107f
C1048 a_3840_10895# RST 7.28e-19
C1049 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 0.122f
C1050 a_10961_15230# VDD 3.14e-19
C1051 a_8709_10895# CLK_DIV_11_mag_new_0.Q2 2.98e-20
C1052 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.321f
C1053 CLK_div_3_mag_0.JK_FF_mag_1.QB VDD 0.875f
C1054 a_13858_15251# CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 2.84e-20
C1055 RST CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.378f
C1056 CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.Q1 1.9e-20
C1057 a_3556_12901# RST 4.17e-19
C1058 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 9.82e-20
C1059 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_DIV_11_mag_new_0.Q1 1.76e-21
C1060 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0934f
C1061 RST a_9233_13028# 3.08e-20
C1062 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.0435f
C1063 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_1.JK_FF_mag_1.K 0.00205f
C1064 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.121f
C1065 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.00359f
C1066 RST a_15500_11885# 0.00176f
C1067 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.00126f
C1068 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.00975f
C1069 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00183f
C1070 a_5852_10895# CLK_DIV_11_mag_new_0.Q3 5.98e-19
C1071 a_4002_14308# VDD 3.14e-19
C1072 a_4002_14308# CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 3.01e-20
C1073 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_DIV_11_mag_new_0.Q0 1.99f
C1074 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_5534_12986# 0.00119f
C1075 a_13475_13030# CLK_DIV_11_mag_new_0.Q1 0.069f
C1076 CLK_div_3_mag_0.JK_FF_mag_1.K a_5128_10895# 0.00695f
C1077 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 8.58e-20
C1078 a_10096_15189# CLK_DIV_11_mag_new_0.and2_mag_3.IN1 0.00271f
C1079 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.Q0 0.11f
C1080 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.Q3 3.26e-20
C1081 CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 4.52e-20
C1082 CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN VDD 0.423f
C1083 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 7.98e-20
C1084 CLK_div_3_mag_0.or_2_mag_0.IN2 a_4558_9798# 4.9e-20
C1085 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK 0.235f
C1086 a_13698_15251# CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 9.09e-19
C1087 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.16f
C1088 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK 0.0215f
C1089 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0622f
C1090 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_DIV_11_mag_new_0.Q3 0.133f
C1091 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.0129f
C1092 CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_3_mag_1.Q0 0.0655f
C1093 RST a_14936_11885# 0.00201f
C1094 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_6816_11933# 0.00378f
C1095 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 a_10927_9798# 0.069f
C1096 a_5692_10895# CLK_DIV_11_mag_new_0.Q3 6.04e-19
C1097 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.Q0 0.0655f
C1098 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.Q2 0.338f
C1099 a_3994_9798# CLK_div_3_mag_0.JK_FF_mag_1.K 0.012f
C1100 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 1.45e-19
C1101 CLK CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 3.43e-19
C1102 CLK_div_3_mag_0.JK_FF_mag_1.K a_4968_10895# 0.00696f
C1103 a_10096_15189# VDD 5.08e-19
C1104 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 3.43e-19
C1105 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VDD 1f
C1106 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_DIV_11_mag_new_0.Q2 0.0579f
C1107 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.Q3 2.12e-19
C1108 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.Q0 0.209f
C1109 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 0.122f
C1110 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 3.67e-20
C1111 a_7421_10895# CLK_DIV_11_mag_new_0.Q3 2.34e-20
C1112 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.109f
C1113 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.Q2 3.45e-19
C1114 a_12215_9798# CLK 0.0101f
C1115 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.Q0 1.83e-20
C1116 a_8139_9798# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0202f
C1117 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.Q3 0.0346f
C1118 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.321f
C1119 RST a_14776_11885# 0.00201f
C1120 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD 0.391f
C1121 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_6252_11889# 0.0733f
C1122 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 a_10363_9798# 0.00372f
C1123 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.103f
C1124 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.36f
C1125 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_15238_10895# 1.17e-20
C1126 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00156f
C1127 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0622f
C1128 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.109f
C1129 CLK_div_3_mag_0.JK_FF_mag_1.K a_4404_10895# 0.00964f
C1130 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 1.08f
C1131 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 7.49e-20
C1132 a_2590_14702# VDD 3.14e-19
C1133 a_8503_11887# a_8663_11887# 0.0504f
C1134 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_DIV_11_mag_new_0.Q1 9.69e-19
C1135 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.Q2 1.05e-19
C1136 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT RST 0.00337f
C1137 CLK_div_3_mag_0.JK_FF_mag_1.K VDD 2.41f
C1138 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.Q1 8.39e-21
C1139 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C1140 a_12055_9798# CLK 0.00939f
C1141 a_15238_10895# CLK 0.00117f
C1142 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0135f
C1143 a_7575_9798# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 4.52e-20
C1144 RST a_13629_11933# 0.00106f
C1145 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.0435f
C1146 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 3.61e-21
C1147 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.121f
C1148 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 1.96e-19
C1149 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_6092_11889# 0.0203f
C1150 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_16224_11929# 0.00378f
C1151 CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.00252f
C1152 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_15078_10895# 1.5e-20
C1153 a_7380_11933# CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.0811f
C1154 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_11783_12986# 1.16e-20
C1155 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.Q2 0.0345f
C1156 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN VDD 0.415f
C1157 a_11783_12986# CLK_DIV_11_mag_new_0.Q1 2.79e-20
C1158 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_1.Q0 0.338f
C1159 CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_DIV_11_mag_new_0.Q3 0.119f
C1160 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT VDD 0.647f
C1161 CLK_div_3_mag_0.JK_FF_mag_1.K a_3840_10895# 0.0811f
C1162 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0702f
C1163 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.36f
C1164 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.122f
C1165 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.QB 0.343f
C1166 CLK_DIV_11_mag_new_0.Q1 CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 0.111f
C1167 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_1.QB 3.67e-20
C1168 a_6816_11933# VDD 3.14e-19
C1169 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_7380_11933# 2.34e-20
C1170 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 2.04e-19
C1171 a_15078_10895# CLK 0.00164f
C1172 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT VDD 0.994f
C1173 a_11491_9798# CLK 6.43e-21
C1174 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 a_12501_11889# 8.64e-19
C1175 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT a_12501_11889# 2.88e-20
C1176 RST a_13065_11933# 0.00129f
C1177 CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 8.33e-20
C1178 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT RST 0.11f
C1179 CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_DIV_11_mag_new_0.Q2 0.00392f
C1180 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT VDD 0.648f
C1181 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_15660_11885# 0.0733f
C1182 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_5528_11889# 1.5e-20
C1183 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K a_5368_11889# 8.64e-19
C1184 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 0.321f
C1185 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_14514_10895# 0.0203f
C1186 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.768f
C1187 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 0.25f
C1188 CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_DIV_11_mag_new_0.nand3_mag_1.OUT 0.109f
C1189 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_11623_12986# 1.49e-20
C1190 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.Q1 1.36e-19
C1191 a_5410_8699# VDD 5.92e-19
C1192 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 RST 6.71e-19
C1193 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK 5.57e-19
C1194 a_10361_13028# CLK_DIV_11_mag_new_0.Q2 0.069f
C1195 a_12347_13030# CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 1.39e-19
C1196 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00118f
C1197 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 6.36e-19
C1198 CLK_DIV_11_mag_new_0.Q3 VDD 5.7f
C1199 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.Q3 1.51e-19
C1200 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00118f
C1201 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD 0.397f
C1202 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.Q0 3.92e-19
C1203 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 2.21e-19
C1204 a_16788_11929# CLK_DIV_11_mag_new_0.Q0 0.0157f
C1205 RST CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.0957f
C1206 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_1.JK_FF_mag_1.QB 2.81e-20
C1207 a_5122_9798# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.0697f
C1208 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.0445f
C1209 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 4.19e-20
C1210 a_5852_10895# CLK_div_3_mag_0.Q0 0.00335f
C1211 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT a_12341_11889# 9.1e-19
C1212 RST CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00535f
C1213 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_9951_11931# 0.0036f
C1214 RST a_12501_11889# 0.00222f
C1215 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 6.18e-19
C1216 CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_DIV_11_mag_new_0.Q1 0.106f
C1217 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.0951f
C1218 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_15506_13026# 3.33e-19
C1219 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_5368_11889# 1.17e-20
C1220 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_15500_11885# 0.0203f
C1221 CLK_DIV_11_mag_new_0.Q2 VDD 2.61f
C1222 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 0.00125f
C1223 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_14354_10895# 0.0733f
C1224 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_12911_13030# 4.52e-20
C1225 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.Q2 0.0131f
C1226 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.nand3_mag_1.OUT 0.00452f
C1227 a_12221_10895# CLK 0.00117f
C1228 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT a_9233_13028# 0.00378f
C1229 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_10361_13028# 0.0114f
C1230 a_12215_9798# RST 7.78e-19
C1231 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 RST 3.79e-19
C1232 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_DIV_11_mag_new_0.Q3 0.029f
C1233 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.Q3 0.0631f
C1234 a_11783_12986# CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 8.21e-19
C1235 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD 0.651f
C1236 CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_DIV_11_mag_new_0.Q0 0.104f
C1237 a_12055_9798# CLK_div_3_mag_1.Q0 2.79e-20
C1238 a_14782_12982# a_14942_12982# 0.0504f
C1239 CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 5.74e-20
C1240 a_5846_9798# VDD 2.21e-19
C1241 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_div_3_mag_0.Q0 1.6e-19
C1242 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 2.33e-19
C1243 a_6092_11889# VDD 2.21e-19
C1244 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.0593f
C1245 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 0.00118f
C1246 a_16224_11929# CLK_DIV_11_mag_new_0.Q0 0.00859f
C1247 a_4558_9798# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.0059f
C1248 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_13629_11933# 2.58e-20
C1249 a_5692_10895# CLK_div_3_mag_0.Q0 0.00789f
C1250 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT a_11777_11889# 0.0731f
C1251 a_16070_13026# CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00605f
C1252 RST a_12341_11889# 0.00206f
C1253 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD 0.651f
C1254 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB VDD 0.904f
C1255 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN RST 0.00222f
C1256 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.Q2 0.109f
C1257 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_14942_12982# 0.00392f
C1258 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT RST 0.336f
C1259 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_14936_11885# 1.5e-20
C1260 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 a_13475_13030# 4.52e-20
C1261 CLK_DIV_11_mag_new_0.Q1 VDD 3.59f
C1262 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.Q1 0.11f
C1263 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_12347_13030# 0.0195f
C1264 a_3556_12901# CLK_DIV_11_mag_new_0.Q2 0.00208f
C1265 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.Q1 8.19e-19
C1266 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_13790_10895# 0.00378f
C1267 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 a_7226_13030# 4.52e-20
C1268 a_11491_9798# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.0202f
C1269 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 a_9797_13028# 0.0059f
C1270 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_9797_13028# 2.96e-19
C1271 CLK_div_3_mag_1.Q0 a_11777_11889# 5.98e-19
C1272 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_1.or_2_mag_0.IN2 0.0445f
C1273 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT a_8669_12984# 0.0732f
C1274 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 3.67e-20
C1275 a_12061_10895# CLK 0.00164f
C1276 a_12055_9798# RST 6.43e-19
C1277 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VDD 0.653f
C1278 a_15238_10895# RST 5.2e-19
C1279 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 6.57e-19
C1280 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 3.72e-19
C1281 a_11623_12986# CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.00598f
C1282 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.Q0 0.00335f
C1283 CLK_DIV_11_mag_new_0.Q0 VDD 3.9f
C1284 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.Q0 3.4e-19
C1285 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.Q0 0.00129f
C1286 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_4437_8231# 3.25e-19
C1287 CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 CLK_DIV_11_mag_new_0.Q3 0.0224f
C1288 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.K 0.0948f
C1289 a_16634_13026# CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 4.52e-20
C1290 a_15660_11885# CLK_DIV_11_mag_new_0.Q0 0.0101f
C1291 a_14354_10895# CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 8.64e-19
C1292 CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 0.00121f
C1293 a_5128_10895# CLK_div_3_mag_0.Q0 0.0102f
C1294 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 9.52e-19
C1295 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT a_11617_11889# 0.0202f
C1296 RST a_11777_11889# 0.00273f
C1297 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.289f
C1298 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 6.51e-19
C1299 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.QB 0.215f
C1300 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_DIV_11_mag_new_0.Q1 3.09e-19
C1301 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.00209f
C1302 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 9.58e-19
C1303 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 2.51e-19
C1304 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.Q1 2.57f
C1305 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 RST 1.38e-19
C1306 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.359f
C1307 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_14776_11885# 1.17e-20
C1308 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.and2_mag_3.IN1 0.00441f
C1309 a_10927_9798# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 4.52e-20
C1310 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.00388f
C1311 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 a_9233_13028# 0.0697f
C1312 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_9233_13028# 3.12e-19
C1313 CLK_div_3_mag_1.Q0 a_11617_11889# 5.98e-19
C1314 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT a_8509_12984# 0.0203f
C1315 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK 0.471f
C1316 a_11491_9798# RST 3.71e-19
C1317 a_15078_10895# RST 5.2e-19
C1318 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 8.28e-20
C1319 a_8669_12984# CLK_DIV_11_mag_new_0.Q2 2.79e-20
C1320 a_10361_13028# CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 8.11e-19
C1321 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_DIV_11_mag_new_0.Q0 1.61e-19
C1322 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.Q0 4.75f
C1323 a_3556_12901# CLK_DIV_11_mag_new_0.Q0 3.17e-19
C1324 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_12221_10895# 1.17e-20
C1325 a_5122_9798# VDD 3.14e-19
C1326 a_12221_10895# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 5.54e-20
C1327 a_5368_11889# VDD 2.21e-19
C1328 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 RST 0.0581f
C1329 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 5.42e-20
C1330 a_3994_9798# CLK_div_3_mag_0.Q0 0.069f
C1331 a_15500_11885# CLK_DIV_11_mag_new_0.Q0 0.0102f
C1332 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 0.0592f
C1333 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.0432f
C1334 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_1.JK_FF_mag_1.K 0.352f
C1335 a_12221_10895# CLK_div_3_mag_1.Q0 0.00335f
C1336 a_4968_10895# CLK_div_3_mag_0.Q0 0.0101f
C1337 a_8703_9798# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00119f
C1338 a_8709_10895# a_8869_10895# 0.0504f
C1339 RST a_11617_11889# 0.00273f
C1340 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_8663_11887# 1.46e-19
C1341 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0899f
C1342 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 0.122f
C1343 CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 2.25e-19
C1344 a_3994_15139# CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 2.69e-22
C1345 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K VDD 0.866f
C1346 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_8669_12984# 0.00392f
C1347 a_10927_9798# RST 3.96e-19
C1348 a_14514_10895# RST 0.00108f
C1349 CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 CLK_DIV_11_mag_new_0.Q1 4.07e-19
C1350 a_15072_9798# a_15232_9798# 0.0504f
C1351 a_14936_11885# CLK_DIV_11_mag_new_0.Q1 4.28e-19
C1352 CLK_div_3_mag_1.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 1.83e-19
C1353 a_9797_13028# CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 3.47e-19
C1354 a_15072_9798# CLK_div_3_mag_1.JK_FF_mag_1.QB 0.00392f
C1355 a_10363_9798# CLK_div_3_mag_1.Q0 0.069f
C1356 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K RST 0.0777f
C1357 a_4558_9798# VDD 3.14e-19
C1358 a_7226_13030# CLK_DIV_11_mag_new_0.Q3 0.069f
C1359 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.00544f
C1360 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_12061_10895# 1.5e-20
C1361 a_12221_10895# RST 0.00498f
C1362 CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 CLK_DIV_11_mag_new_0.Q0 1.32e-19
C1363 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 1.84e-21
C1364 a_14936_11885# CLK_DIV_11_mag_new_0.Q0 0.00789f
C1365 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_5466_15136# 8.64e-19
C1366 a_4404_10895# CLK_div_3_mag_0.Q0 0.00859f
C1367 a_10256_15189# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 4.33e-21
C1368 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 0.121f
C1369 a_8139_9798# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.43e-19
C1370 a_12061_10895# CLK_div_3_mag_1.Q0 0.00789f
C1371 RST a_10515_11931# 0.00137f
C1372 RST CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0301f
C1373 CLK_div_3_mag_0.Q0 VDD 1.24f
C1374 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.Q0 1.08e-20
C1375 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.161f
C1376 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT RST 0.286f
C1377 CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.103f
C1378 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.K 0.0725f
C1379 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.198f
C1380 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.00301f
C1381 a_10363_9798# RST 3.96e-19
C1382 CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 1.82e-19
C1383 a_14354_10895# RST 0.00173f
C1384 a_14776_11885# CLK_DIV_11_mag_new_0.Q1 5.5e-19
C1385 a_14508_9798# CLK_div_3_mag_1.JK_FF_mag_1.QB 3.33e-19
C1386 CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.132f
C1387 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.QB 1.04e-19
C1388 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 1.82e-19
C1389 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_11497_10895# 0.0203f
C1390 a_2757_14017# CLK_DIV_11_mag_new_0.nand3_mag_0.OUT 0.0732f
C1391 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C1392 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT a_6098_13030# 0.00378f
C1393 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0622f
C1394 a_12061_10895# RST 0.00495f
C1395 a_14776_11885# CLK_DIV_11_mag_new_0.Q0 0.00335f
C1396 a_10806_8231# CLK_div_3_mag_1.JK_FF_mag_1.K 0.00168f
C1397 a_3840_10895# CLK_div_3_mag_0.Q0 0.0157f
C1398 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 0.121f
C1399 a_7575_9798# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.011f
C1400 a_11497_10895# CLK_div_3_mag_1.Q0 0.0102f
C1401 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_1.Q0 0.0175f
C1402 RST a_9951_11931# 0.00136f
C1403 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.233f
C1404 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00118f
C1405 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT VDD 0.994f
C1406 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 0.00975f
C1407 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.16f
C1408 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 9.62e-20
C1409 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_15078_10895# 1.46e-19
C1410 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT RST 0.0634f
C1411 CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT VDD 0.345f
C1412 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.and2_mag_3.OUT 1.39e-19
C1413 a_13790_10895# RST 0.00108f
C1414 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 RST 0.00825f
C1415 a_13629_11933# CLK_DIV_11_mag_new_0.Q1 0.0157f
C1416 CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 VDD 0.657f
C1417 CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 0.0512f
C1418 a_15232_9798# CLK_div_3_mag_1.JK_FF_mag_1.K 8.64e-19
C1419 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 2.34e-19
C1420 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.313f
C1421 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.QB 3.28e-19
C1422 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 a_6662_13030# 0.0059f
C1423 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_11337_10895# 0.0733f
C1424 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT a_5534_12986# 0.0732f
C1425 a_2597_14017# CLK_DIV_11_mag_new_0.nand3_mag_0.OUT 0.0202f
C1426 a_11497_10895# RST 0.00343f
C1427 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 RST 0.0238f
C1428 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 5.63e-21
C1429 a_7011_9798# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00118f
C1430 a_11337_10895# CLK_div_3_mag_1.Q0 0.0101f
C1431 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.25f
C1432 RST a_9387_11887# 0.00222f
C1433 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT 0.00296f
C1434 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT 1.2e-19
C1435 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 RST 0.0698f
C1436 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VDD 0.647f
C1437 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 1.83e-19
C1438 a_13226_10895# RST 0.00214f
C1439 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN a_3994_9798# 4.94e-20
C1440 a_13065_11933# CLK_DIV_11_mag_new_0.Q1 0.00859f
C1441 a_13380_9798# CLK_div_3_mag_1.JK_FF_mag_1.QB 0.0112f
C1442 a_15506_13026# VDD 3.14e-19
C1443 CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 a_3556_12901# 0.0177f
C1444 CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 VDD 0.339f
C1445 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.Q1 0.00101f
C1446 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 a_6098_13030# 0.0697f
C1447 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT a_5374_12986# 0.0203f
C1448 a_2597_14017# a_2757_14017# 0.0504f
C1449 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_10773_10895# 0.00378f
C1450 a_5534_12986# CLK_DIV_11_mag_new_0.Q3 3.43e-19
C1451 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.00169f
C1452 a_11337_10895# RST 0.00327f
C1453 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.Q3 8.62e-19
C1454 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q3 0.329f
C1455 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C1456 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 2.39e-21
C1457 a_10773_10895# CLK_div_3_mag_1.Q0 0.00859f
C1458 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.00975f
C1459 a_7985_10895# a_8145_10895# 0.0504f
C1460 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD 0.392f
C1461 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 8.16e-20
C1462 RST a_9227_11887# 0.00206f
C1463 CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT CLK_DIV_11_mag_new_0.Q3 0.0238f
C1464 a_13858_15251# CLK_DIV_11_mag_new_0.and2_mag_3.OUT 8.64e-19
C1465 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.Q1 3.39e-20
C1466 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_16788_11929# 0.0811f
C1467 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.and2_mag_3.OUT 2.22e-20
C1468 CLK_div_3_mag_0.or_2_mag_0.IN2 VDD 0.492f
C1469 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_7421_10895# 0.069f
C1470 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_1.Q0 6.11e-20
C1471 a_12501_11889# CLK_DIV_11_mag_new_0.Q1 0.0101f
C1472 CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT 0.0121f
C1473 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q2 0.0609f
C1474 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.Q0 0.338f
C1475 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VDD 0.392f
C1476 a_5374_12986# CLK_DIV_11_mag_new_0.Q3 4.47e-19
C1477 a_4437_8231# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.4e-19
C1478 RST CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.303f
C1479 a_5692_10895# a_5852_10895# 0.0504f
C1480 a_10773_10895# RST 0.00382f
C1481 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.Q0 0.0399f
C1482 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VDD 0.414f
C1483 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.198f
C1484 a_10209_10895# CLK_div_3_mag_1.Q0 0.0157f
C1485 RST a_8663_11887# 0.00273f
C1486 a_13698_15251# CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.0105f
C1487 CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 RST 0.00591f
C1488 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 RST 0.145f
C1489 a_8703_9798# a_8863_9798# 0.0504f
C1490 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.K 0.23f
C1491 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_13790_10895# 0.0036f
C1492 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_16224_11929# 0.00964f
C1493 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 1.83e-19
C1494 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 3.43e-19
C1495 a_10806_8231# VDD 0.165f
C1496 a_14942_12982# CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 1.19e-20
C1497 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_6857_10895# 0.00372f
C1498 a_12341_11889# CLK_DIV_11_mag_new_0.Q1 0.0102f
C1499 a_14782_12982# VDD 2.21e-19
C1500 a_11777_11889# CLK_DIV_11_mag_new_0.Q2 4.66e-19
C1501 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K a_6816_11933# 4.96e-22
C1502 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q1 0.116f
C1503 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 2.32e-19
C1504 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.Q2 0.109f
C1505 a_8869_10895# VDD 0.0132f
C1506 a_10209_10895# RST 0.00373f
C1507 CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT CLK_DIV_11_mag_new_0.Q1 3.09e-19
C1508 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN a_10363_9798# 4.94e-20
C1509 a_15232_9798# VDD 5.99e-19
C1510 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0951f
C1511 CLK_div_3_mag_1.JK_FF_mag_1.QB VDD 0.875f
C1512 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK 7.81e-19
C1513 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q0 0.00115f
C1514 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 6.3e-20
C1515 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 7.97e-19
C1516 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB VDD 0.904f
C1517 RST a_8503_11887# 0.00273f
C1518 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.QB 0.21f
C1519 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.JK_FF_mag_1.K 0.00384f
C1520 a_10961_15230# CLK_DIV_11_mag_new_0.and2_mag_3.OUT 6.43e-19
C1521 CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT CLK_DIV_11_mag_new_0.Q0 1.61e-19
C1522 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 4.26e-19
C1523 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD 0.397f
C1524 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_15660_11885# 0.00696f
C1525 a_11779_8699# VDD 5.92e-19
C1526 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.Q3 0.0703f
C1527 RST CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.0864f
C1528 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.198f
C1529 a_7985_10895# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 8.64e-19
C1530 a_14782_12982# CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 1.52e-20
C1531 a_13475_13030# VDD 3.56e-19
C1532 a_11617_11889# CLK_DIV_11_mag_new_0.Q2 6.02e-19
C1533 a_11777_11889# CLK_DIV_11_mag_new_0.Q1 0.00789f
C1534 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C1535 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0592f
C1536 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 a_13475_13030# 0.00372f
C1537 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.121f
C1538 a_3994_15139# CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 0.132f
C1539 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.Q1 1.17e-19
C1540 a_8709_10895# VDD 0.00888f
C1541 a_15072_9798# VDD 2.65e-19
C1542 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.Q3 9.67e-20
C1543 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00183f
C1544 a_11491_9798# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.0697f
C1545 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.Q0 6.35e-19
C1546 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_1.Q0 4.76e-19
C1547 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD 0.394f
C1548 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.Q2 0.0398f
C1549 RST a_7380_11933# 0.00161f
C1550 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.Q1 1.06e-19
C1551 a_15078_10895# CLK_DIV_11_mag_new_0.Q0 2.58e-20
C1552 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN a_5466_15136# 2.4e-20
C1553 a_4558_9798# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.069f
C1554 a_13698_15251# CLK_DIV_11_mag_new_0.nand3_mag_1.OUT 8.09e-22
C1555 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 3.6e-19
C1556 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_15500_11885# 0.00695f
C1557 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 1.99e-19
C1558 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_13065_11933# 0.00378f
C1559 RST CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.103f
C1560 RST CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT 0.00543f
C1561 a_13475_13030# CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.0114f
C1562 a_11617_11889# CLK_DIV_11_mag_new_0.Q1 0.00335f
C1563 a_12911_13030# VDD 3.14e-19
C1564 a_10515_11931# CLK_DIV_11_mag_new_0.Q2 0.0157f
C1565 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 a_12911_13030# 0.069f
C1566 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.Q2 0.0635f
C1567 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VDD 0.802f
C1568 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_5410_8699# 0.069f
C1569 a_11623_12986# a_11783_12986# 0.0504f
C1570 a_8145_10895# VDD 0.0012f
C1571 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00183f
C1572 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.Q0 0.107f
C1573 a_10806_8231# VSS 0.0247f
C1574 a_11779_8699# VSS 0.0676f
C1575 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN VSS 0.435f
C1576 a_4437_8231# VSS 0.0247f
C1577 CLK_div_3_mag_1.or_2_mag_0.IN2 VSS 0.418f
C1578 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN VSS 0.6f
C1579 a_5410_8699# VSS 0.0676f
C1580 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS 0.435f
C1581 CLK_div_3_mag_0.or_2_mag_0.IN2 VSS 0.418f
C1582 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS 0.6f
C1583 a_15232_9798# VSS 0.0881f
C1584 a_15072_9798# VSS 0.0343f
C1585 a_14508_9798# VSS 0.0676f
C1586 a_13944_9798# VSS 0.0676f
C1587 a_13380_9798# VSS 0.0676f
C1588 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.509f
C1589 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.415f
C1590 a_12215_9798# VSS 0.0881f
C1591 a_12055_9798# VSS 0.0343f
C1592 a_11491_9798# VSS 0.0676f
C1593 a_10927_9798# VSS 0.0676f
C1594 a_10363_9798# VSS 0.0676f
C1595 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C1596 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.415f
C1597 a_8863_9798# VSS 0.0881f
C1598 a_8703_9798# VSS 0.0343f
C1599 a_8139_9798# VSS 0.0676f
C1600 a_7575_9798# VSS 0.0676f
C1601 a_7011_9798# VSS 0.0676f
C1602 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.509f
C1603 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.415f
C1604 a_5846_9798# VSS 0.0881f
C1605 a_5686_9798# VSS 0.0343f
C1606 a_5122_9798# VSS 0.0676f
C1607 a_4558_9798# VSS 0.0676f
C1608 a_3994_9798# VSS 0.0676f
C1609 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C1610 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.415f
C1611 a_15238_10895# VSS 0.0881f
C1612 a_15078_10895# VSS 0.0343f
C1613 a_14514_10895# VSS 0.0881f
C1614 a_14354_10895# VSS 0.0343f
C1615 a_13790_10895# VSS 0.0676f
C1616 a_13226_10895# VSS 0.0675f
C1617 CLK_div_3_mag_1.JK_FF_mag_1.QB VSS 0.859f
C1618 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.811f
C1619 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.695f
C1620 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.418f
C1621 a_12221_10895# VSS 0.0881f
C1622 a_12061_10895# VSS 0.0343f
C1623 a_11497_10895# VSS 0.0881f
C1624 a_11337_10895# VSS 0.0343f
C1625 a_10773_10895# VSS 0.0676f
C1626 a_10209_10895# VSS 0.0675f
C1627 CLK_div_3_mag_1.JK_FF_mag_1.K VSS 4.56f
C1628 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.811f
C1629 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.691f
C1630 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.417f
C1631 a_8869_10895# VSS 0.0881f
C1632 a_8709_10895# VSS 0.0343f
C1633 a_8145_10895# VSS 0.0881f
C1634 a_7985_10895# VSS 0.0343f
C1635 a_7421_10895# VSS 0.0676f
C1636 a_6857_10895# VSS 0.0675f
C1637 CLK_div_3_mag_0.JK_FF_mag_1.QB VSS 0.859f
C1638 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.81f
C1639 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.7f
C1640 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.417f
C1641 a_5852_10895# VSS 0.0881f
C1642 a_5692_10895# VSS 0.0343f
C1643 a_5128_10895# VSS 0.0881f
C1644 a_4968_10895# VSS 0.0343f
C1645 a_4404_10895# VSS 0.0676f
C1646 a_3840_10895# VSS 0.0675f
C1647 CLK_div_3_mag_0.JK_FF_mag_1.K VSS 4.51f
C1648 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.81f
C1649 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.691f
C1650 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.417f
C1651 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.521f
C1652 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.726f
C1653 CLK VSS 2.9f
C1654 CLK_div_3_mag_1.Q0 VSS 2.54f
C1655 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.541f
C1656 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.727f
C1657 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.522f
C1658 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.726f
C1659 CLK_div_3_mag_0.Q0 VSS 2.3f
C1660 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.54f
C1661 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.726f
C1662 a_16788_11929# VSS 0.0696f
C1663 a_16224_11929# VSS 0.0698f
C1664 a_15660_11885# VSS 0.0378f
C1665 a_15500_11885# VSS 0.0916f
C1666 a_14936_11885# VSS 0.0378f
C1667 a_14776_11885# VSS 0.0917f
C1668 a_13629_11933# VSS 0.069f
C1669 a_13065_11933# VSS 0.0691f
C1670 a_12501_11889# VSS 0.0367f
C1671 a_12341_11889# VSS 0.0905f
C1672 a_11777_11889# VSS 0.0368f
C1673 a_11617_11889# VSS 0.0906f
C1674 a_10515_11931# VSS 0.0693f
C1675 a_9951_11931# VSS 0.0694f
C1676 a_9387_11887# VSS 0.0372f
C1677 a_9227_11887# VSS 0.0911f
C1678 a_8663_11887# VSS 0.0373f
C1679 a_8503_11887# VSS 0.0911f
C1680 a_7380_11933# VSS 0.069f
C1681 a_6816_11933# VSS 0.0691f
C1682 a_6252_11889# VSS 0.0367f
C1683 a_6092_11889# VSS 0.0905f
C1684 a_5528_11889# VSS 0.0368f
C1685 a_5368_11889# VSS 0.0906f
C1686 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 VSS 0.421f
C1687 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT VSS 0.553f
C1688 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 VSS 0.42f
C1689 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT VSS 0.549f
C1690 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.42f
C1691 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.551f
C1692 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.419f
C1693 RST VSS 6.79f
C1694 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.548f
C1695 a_2597_12515# VSS 0.0716f
C1696 a_16634_13026# VSS 0.0744f
C1697 a_16070_13026# VSS 0.0745f
C1698 a_15506_13026# VSS 0.0744f
C1699 a_14942_12982# VSS 0.047f
C1700 a_14782_12982# VSS 0.101f
C1701 a_13475_13030# VSS 0.0734f
C1702 a_12911_13030# VSS 0.0735f
C1703 a_12347_13030# VSS 0.0735f
C1704 a_11783_12986# VSS 0.0449f
C1705 a_11623_12986# VSS 0.0987f
C1706 a_10361_13028# VSS 0.0739f
C1707 a_9797_13028# VSS 0.074f
C1708 a_9233_13028# VSS 0.0739f
C1709 a_8669_12984# VSS 0.0459f
C1710 a_8509_12984# VSS 0.0997f
C1711 a_7226_13030# VSS 0.0737f
C1712 a_6662_13030# VSS 0.0737f
C1713 a_6098_13030# VSS 0.0737f
C1714 a_5534_12986# VSS 0.0454f
C1715 a_5374_12986# VSS 0.0992f
C1716 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 VSS 0.425f
C1717 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 VSS 0.908f
C1718 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 VSS 0.756f
C1719 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT VSS 0.832f
C1720 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT VSS 0.549f
C1721 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB VSS 0.954f
C1722 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN VSS 0.612f
C1723 a_3556_12901# VSS 0.0247f
C1724 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN VSS 0.45f
C1725 CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 VSS 0.491f
C1726 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 VSS 0.424f
C1727 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 VSS 0.86f
C1728 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 VSS 0.744f
C1729 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT VSS 0.828f
C1730 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT VSS 0.543f
C1731 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.424f
C1732 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.832f
C1733 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.745f
C1734 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.83f
C1735 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.546f
C1736 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB VSS 0.912f
C1737 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.424f
C1738 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.844f
C1739 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.743f
C1740 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.827f
C1741 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.544f
C1742 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K VSS 1.92f
C1743 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K VSS 3.11f
C1744 CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 VSS 0.403f
C1745 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT VSS 0.585f
C1746 a_2757_14017# VSS 0.0343f
C1747 a_2597_14017# VSS 0.0881f
C1748 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN VSS 0.464f
C1749 a_4002_14308# VSS 0.0676f
C1750 Vdiv99 VSS 0.36f
C1751 a_13858_15251# VSS 0.0376f
C1752 a_13698_15251# VSS 0.0391f
C1753 a_10961_15230# VSS 0.0693f
C1754 a_10256_15189# VSS 0.0362f
C1755 a_10096_15189# VSS 0.0901f
C1756 a_2590_14702# VSS 0.0678f
C1757 CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT VSS 1.03f
C1758 CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 VSS 0.555f
C1759 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K VSS 2.9f
C1760 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN VSS 0.676f
C1761 CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT VSS 0.678f
C1762 CLK_DIV_11_mag_new_0.and2_mag_3.OUT VSS 1.93f
C1763 CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN VSS 0.597f
C1764 a_5466_15136# VSS 0.0247f
C1765 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K VSS 2.89f
C1766 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 VSS 18.6f
C1767 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 VSS 2.52f
C1768 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN VSS 0.589f
C1769 a_3994_15139# VSS 0.0247f
C1770 CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN VSS 0.453f
C1771 CLK_DIV_11_mag_new_0.Q3 VSS 6.57f
C1772 CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 VSS 0.532f
C1773 CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN VSS 0.457f
C1774 CLK_DIV_11_mag_new_0.Q1 VSS 6.69f
C1775 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS 0.701f
C1776 CLK_DIV_11_mag_new_0.Q2 VSS 6.76f
C1777 CLK_DIV_11_mag_new_0.Q0 VSS 6.43f
C1778 CLK_DIV_11_mag_new_0.and2_mag_3.IN1 VSS 0.834f
C1779 CLK_DIV_11_mag_new_0.nand3_mag_1.OUT VSS 0.741f
C1780 VDD VSS 0.173p
C1781 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t3 VSS 0.0207f
C1782 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t2 VSS 0.0271f
C1783 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n0 VSS 0.0537f
C1784 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t4 VSS 0.0273f
C1785 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t5 VSS 0.0207f
C1786 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n1 VSS 0.0537f
C1787 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n2 VSS 0.675f
C1788 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n3 VSS 0.0327f
C1789 CLK_div_3_mag_0.Vdiv3.n0 VSS 0.192f
C1790 CLK_div_3_mag_0.Vdiv3.n1 VSS 0.0484f
C1791 CLK_div_3_mag_0.Vdiv3.n2 VSS 0.156f
C1792 CLK_div_3_mag_0.Vdiv3.n3 VSS 0.00958f
C1793 CLK_div_3_mag_0.Vdiv3.n4 VSS 0.186f
C1794 CLK_div_3_mag_0.Vdiv3.n5 VSS 0.00958f
C1795 CLK_div_3_mag_0.Vdiv3.n6 VSS 0.186f
C1796 CLK_div_3_mag_0.Vdiv3.n7 VSS 0.00958f
C1797 CLK_div_3_mag_0.Vdiv3.n8 VSS 0.186f
C1798 CLK_div_3_mag_0.Vdiv3.n9 VSS 0.00958f
C1799 CLK_div_3_mag_0.Vdiv3.n10 VSS 0.0653f
C1800 CLK_div_3_mag_0.Vdiv3.n11 VSS 0.0653f
C1801 CLK_div_3_mag_0.Vdiv3.n12 VSS 0.0653f
C1802 CLK_div_3_mag_0.Vdiv3.n13 VSS 0.0653f
C1803 CLK_div_3_mag_0.Vdiv3.n14 VSS 0.0478f
C1804 CLK_div_3_mag_0.Vdiv3.n15 VSS 0.0478f
C1805 CLK_div_3_mag_0.Vdiv3.n16 VSS 0.0478f
C1806 CLK_div_3_mag_0.Vdiv3.n17 VSS 0.0092f
C1807 CLK_div_3_mag_0.Vdiv3.t1 VSS 0.00793f
C1808 CLK_div_3_mag_0.Vdiv3.t0 VSS 0.0264f
C1809 CLK_div_3_mag_0.Vdiv3.n18 VSS 0.0913f
C1810 CLK_div_3_mag_0.Vdiv3.t10 VSS 0.0155f
C1811 CLK_div_3_mag_0.Vdiv3.t9 VSS 0.0235f
C1812 CLK_div_3_mag_0.Vdiv3.n19 VSS 0.0416f
C1813 CLK_div_3_mag_0.Vdiv3.t22 VSS 0.0155f
C1814 CLK_div_3_mag_0.Vdiv3.t3 VSS 0.0235f
C1815 CLK_div_3_mag_0.Vdiv3.n20 VSS 0.0416f
C1816 CLK_div_3_mag_0.Vdiv3.t2 VSS 0.0194f
C1817 CLK_div_3_mag_0.Vdiv3.t20 VSS 0.00496f
C1818 CLK_div_3_mag_0.Vdiv3.n21 VSS 0.0321f
C1819 CLK_div_3_mag_0.Vdiv3.t7 VSS 0.0155f
C1820 CLK_div_3_mag_0.Vdiv3.t15 VSS 0.0235f
C1821 CLK_div_3_mag_0.Vdiv3.n22 VSS 0.0416f
C1822 CLK_div_3_mag_0.Vdiv3.t23 VSS 0.0155f
C1823 CLK_div_3_mag_0.Vdiv3.t5 VSS 0.0235f
C1824 CLK_div_3_mag_0.Vdiv3.n23 VSS 0.0416f
C1825 CLK_div_3_mag_0.Vdiv3.t25 VSS 0.0194f
C1826 CLK_div_3_mag_0.Vdiv3.t6 VSS 0.00496f
C1827 CLK_div_3_mag_0.Vdiv3.n24 VSS 0.0322f
C1828 CLK_div_3_mag_0.Vdiv3.t19 VSS 0.0155f
C1829 CLK_div_3_mag_0.Vdiv3.t26 VSS 0.0235f
C1830 CLK_div_3_mag_0.Vdiv3.n25 VSS 0.0416f
C1831 CLK_div_3_mag_0.Vdiv3.t13 VSS 0.0155f
C1832 CLK_div_3_mag_0.Vdiv3.t21 VSS 0.0235f
C1833 CLK_div_3_mag_0.Vdiv3.n26 VSS 0.0416f
C1834 CLK_div_3_mag_0.Vdiv3.t16 VSS 0.0194f
C1835 CLK_div_3_mag_0.Vdiv3.t24 VSS 0.00496f
C1836 CLK_div_3_mag_0.Vdiv3.n27 VSS 0.0322f
C1837 CLK_div_3_mag_0.Vdiv3.t8 VSS 0.0155f
C1838 CLK_div_3_mag_0.Vdiv3.t11 VSS 0.0235f
C1839 CLK_div_3_mag_0.Vdiv3.n28 VSS 0.0418f
C1840 CLK_div_3_mag_0.Vdiv3.t18 VSS 0.0155f
C1841 CLK_div_3_mag_0.Vdiv3.t17 VSS 0.0235f
C1842 CLK_div_3_mag_0.Vdiv3.n29 VSS 0.0416f
C1843 CLK_div_3_mag_0.Vdiv3.t4 VSS 0.0155f
C1844 CLK_div_3_mag_0.Vdiv3.t12 VSS 0.0235f
C1845 CLK_div_3_mag_0.Vdiv3.n30 VSS 0.0416f
C1846 CLK_div_3_mag_0.Vdiv3.t14 VSS 0.00496f
C1847 CLK_div_3_mag_0.Vdiv3.t27 VSS 0.0194f
C1848 CLK_div_3_mag_0.Vdiv3.n31 VSS 0.0322f
C1849 CLK_div_3_mag_0.Vdiv3.n32 VSS 0.368f
C1850 CLK_div_3_mag_0.Vdiv3.n33 VSS 1.93f
C1851 CLK_div_3_mag_0.Vdiv3.n34 VSS 1.85f
C1852 CLK_div_3_mag_0.Vdiv3.n35 VSS 0.321f
C1853 CLK_div_3_mag_0.Vdiv3.n36 VSS 0.0147f
C1854 RST.t3 VSS 0.0116f
C1855 RST.t2 VSS 0.0176f
C1856 RST.n0 VSS 0.031f
C1857 RST.n1 VSS 0.00568f
C1858 RST.n2 VSS 0.00192f
C1859 RST.n3 VSS 0.00701f
C1860 RST.n4 VSS 0.0106f
C1861 RST.n5 VSS 0.00639f
C1862 RST.n6 VSS 0.00238f
C1863 RST.t7 VSS 0.0116f
C1864 RST.t12 VSS 0.0176f
C1865 RST.n7 VSS 0.031f
C1866 RST.n8 VSS 0.00438f
C1867 RST.n9 VSS 0.0017f
C1868 RST.n10 VSS 0.00239f
C1869 RST.n11 VSS 0.00833f
C1870 RST.n12 VSS 7.34e-19
C1871 RST.n13 VSS 0.022f
C1872 RST.n14 VSS 0.443f
C1873 RST.n15 VSS 0.442f
C1874 RST.n16 VSS 0.436f
C1875 RST.n17 VSS 0.436f
C1876 RST.n18 VSS 0.0067f
C1877 RST.n19 VSS 0.00126f
C1878 RST.t8 VSS 0.0116f
C1879 RST.t15 VSS 0.0176f
C1880 RST.n20 VSS 0.031f
C1881 RST.n21 VSS 0.00465f
C1882 RST.n22 VSS 0.00239f
C1883 RST.n23 VSS 0.0011f
C1884 RST.n24 VSS 4.95e-19
C1885 RST.n25 VSS 0.00231f
C1886 RST.n26 VSS 0.00123f
C1887 RST.n27 VSS 0.00676f
C1888 RST.n28 VSS 0.00492f
C1889 RST.n29 VSS 0.434f
C1890 RST.n30 VSS 0.435f
C1891 RST.n31 VSS 0.00652f
C1892 RST.n32 VSS 0.00745f
C1893 RST.n33 VSS 0.00248f
C1894 RST.t14 VSS 0.0116f
C1895 RST.t13 VSS 0.0176f
C1896 RST.n34 VSS 0.031f
C1897 RST.n35 VSS 0.00433f
C1898 RST.n36 VSS 0.00148f
C1899 RST.n37 VSS 7.34e-19
C1900 RST.n38 VSS 0.00202f
C1901 RST.n39 VSS 0.00477f
C1902 RST.n40 VSS 8.42e-19
C1903 RST.n41 VSS 0.0564f
C1904 RST.n42 VSS 0.0761f
C1905 RST.n43 VSS 0.00506f
C1906 RST.t0 VSS 0.0178f
C1907 RST.t11 VSS 0.0113f
C1908 RST.n44 VSS 0.0312f
C1909 RST.n45 VSS 0.00405f
C1910 RST.n46 VSS 0.0027f
C1911 RST.n47 VSS 0.00143f
C1912 RST.n48 VSS 0.06f
C1913 RST.n49 VSS 0.00181f
C1914 RST.n50 VSS 0.00545f
C1915 RST.t4 VSS 0.0176f
C1916 RST.t1 VSS 0.0116f
C1917 RST.n51 VSS 0.031f
C1918 RST.n52 VSS 0.00405f
C1919 RST.n53 VSS 0.00145f
C1920 RST.n54 VSS 0.115f
C1921 RST.n55 VSS 0.00506f
C1922 RST.t10 VSS 0.0178f
C1923 RST.t6 VSS 0.0113f
C1924 RST.n56 VSS 0.0312f
C1925 RST.n57 VSS 0.00405f
C1926 RST.n58 VSS 0.0027f
C1927 RST.n59 VSS 0.00143f
C1928 RST.n60 VSS 0.0692f
C1929 RST.n61 VSS 0.866f
C1930 RST.n62 VSS 0.00181f
C1931 RST.n63 VSS 0.00545f
C1932 RST.t9 VSS 0.0176f
C1933 RST.t5 VSS 0.0116f
C1934 RST.n64 VSS 0.031f
C1935 RST.n65 VSS 0.00405f
C1936 RST.n66 VSS 0.00145f
C1937 RST.n67 VSS 0.115f
C1938 RST.n68 VSS 0.777f
C1939 RST.n69 VSS 0.143f
C1940 RST.n70 VSS 0.296f
C1941 RST.n71 VSS 0.183f
C1942 RST.n72 VSS 0.276f
C1943 CLK_div_3_mag_0.Q1.t2 VSS 0.021f
C1944 CLK_div_3_mag_0.Q1.t0 VSS 0.0173f
C1945 CLK_div_3_mag_0.Q1.n0 VSS 0.0173f
C1946 CLK_div_3_mag_0.Q1.n1 VSS 0.0415f
C1947 CLK_div_3_mag_0.Q1.t8 VSS 0.0276f
C1948 CLK_div_3_mag_0.Q1.t10 VSS 0.0221f
C1949 CLK_div_3_mag_0.Q1.n2 VSS 0.0625f
C1950 CLK_div_3_mag_0.Q1.t7 VSS 0.0277f
C1951 CLK_div_3_mag_0.Q1.t4 VSS 0.0355f
C1952 CLK_div_3_mag_0.Q1.n3 VSS 0.0706f
C1953 CLK_div_3_mag_0.Q1.n4 VSS 0.321f
C1954 CLK_div_3_mag_0.Q1.t9 VSS 0.0385f
C1955 CLK_div_3_mag_0.Q1.t6 VSS 0.0254f
C1956 CLK_div_3_mag_0.Q1.n5 VSS 0.0684f
C1957 CLK_div_3_mag_0.Q1.t5 VSS 0.0276f
C1958 CLK_div_3_mag_0.Q1.t3 VSS 0.0221f
C1959 CLK_div_3_mag_0.Q1.n6 VSS 0.0642f
C1960 CLK_div_3_mag_0.Q1.n7 VSS 0.505f
C1961 CLK_div_3_mag_0.Q1.n8 VSS 0.209f
C1962 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t5 VSS 0.154f
C1963 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t4 VSS 0.0457f
C1964 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n0 VSS 0.158f
C1965 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t6 VSS 0.0621f
C1966 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t3 VSS 0.0779f
C1967 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n1 VSS 0.184f
C1968 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t8 VSS 0.109f
C1969 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t7 VSS 0.0696f
C1970 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n2 VSS 0.193f
C1971 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n3 VSS 1.79f
C1972 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t0 VSS 0.589f
C1973 CLK.n0 VSS 0.0185f
C1974 CLK.t5 VSS 0.0521f
C1975 CLK.t13 VSS 0.0343f
C1976 CLK.n1 VSS 0.0919f
C1977 CLK.n2 VSS 0.012f
C1978 CLK.n3 VSS 0.00864f
C1979 CLK.n4 VSS 0.00427f
C1980 CLK.n5 VSS 0.00864f
C1981 CLK.n6 VSS 0.00431f
C1982 CLK.t11 VSS 0.0521f
C1983 CLK.t10 VSS 0.0343f
C1984 CLK.n7 VSS 0.092f
C1985 CLK.n8 VSS 0.012f
C1986 CLK.n9 VSS 0.017f
C1987 CLK.n10 VSS 0.173f
C1988 CLK.n11 VSS 0.17f
C1989 CLK.n12 VSS 0.0995f
C1990 CLK.t7 VSS 0.0521f
C1991 CLK.t2 VSS 0.0343f
C1992 CLK.n13 VSS 0.0919f
C1993 CLK.n14 VSS 0.012f
C1994 CLK.n15 VSS 0.00864f
C1995 CLK.n16 VSS 0.00427f
C1996 CLK.t8 VSS 0.0521f
C1997 CLK.t4 VSS 0.0343f
C1998 CLK.n17 VSS 0.092f
C1999 CLK.n18 VSS 0.00864f
C2000 CLK.n19 VSS 0.00431f
C2001 CLK.n20 VSS 0.012f
C2002 CLK.n21 VSS 0.017f
C2003 CLK.n22 VSS 0.161f
C2004 CLK.t0 VSS 0.027f
C2005 CLK.t3 VSS 0.0482f
C2006 CLK.n23 VSS 0.0919f
C2007 CLK.n24 VSS 0.295f
C2008 CLK.n25 VSS 0.354f
C2009 CLK.n26 VSS 0.0133f
C2010 CLK.n27 VSS 0.0995f
C2011 CLK.n28 VSS 0.0185f
C2012 CLK.n29 VSS 0.0309f
C2013 CLK.t1 VSS 0.0429f
C2014 CLK.t9 VSS 0.0111f
C2015 CLK.n30 VSS 0.0711f
C2016 CLK.n31 VSS 0.0151f
C2017 CLK.n32 VSS 0.00526f
C2018 CLK.n33 VSS 0.0112f
C2019 CLK.n34 VSS 0.658f
C2020 CLK.n35 VSS 0.658f
C2021 CLK.n36 VSS 0.0112f
C2022 CLK.t6 VSS 0.0111f
C2023 CLK.t12 VSS 0.0429f
C2024 CLK.n37 VSS 0.0711f
C2025 CLK.n38 VSS 0.0151f
C2026 CLK.n39 VSS 0.00526f
C2027 CLK.n40 VSS 0.0146f
C2028 CLK_div_3_mag_0.CLK.n0 VSS 0.52f
C2029 CLK_div_3_mag_0.CLK.n1 VSS 0.328f
C2030 CLK_div_3_mag_0.CLK.n2 VSS 0.0208f
C2031 CLK_div_3_mag_0.CLK.n3 VSS 0.0494f
C2032 CLK_div_3_mag_0.CLK.n4 VSS 0.0494f
C2033 CLK_div_3_mag_0.CLK.t1 VSS 0.0172f
C2034 CLK_div_3_mag_0.CLK.t0 VSS 0.0571f
C2035 CLK_div_3_mag_0.CLK.n5 VSS 0.198f
C2036 CLK_div_3_mag_0.CLK.t13 VSS 0.0109f
C2037 CLK_div_3_mag_0.CLK.t8 VSS 0.042f
C2038 CLK_div_3_mag_0.CLK.n6 VSS 0.0697f
C2039 CLK_div_3_mag_0.CLK.t6 VSS 0.0509f
C2040 CLK_div_3_mag_0.CLK.t2 VSS 0.0335f
C2041 CLK_div_3_mag_0.CLK.n7 VSS 0.09f
C2042 CLK_div_3_mag_0.CLK.t3 VSS 0.0509f
C2043 CLK_div_3_mag_0.CLK.t14 VSS 0.0335f
C2044 CLK_div_3_mag_0.CLK.n8 VSS 0.09f
C2045 CLK_div_3_mag_0.CLK.t11 VSS 0.0509f
C2046 CLK_div_3_mag_0.CLK.t7 VSS 0.0335f
C2047 CLK_div_3_mag_0.CLK.n9 VSS 0.09f
C2048 CLK_div_3_mag_0.CLK.t4 VSS 0.0264f
C2049 CLK_div_3_mag_0.CLK.t5 VSS 0.0472f
C2050 CLK_div_3_mag_0.CLK.n10 VSS 0.0899f
C2051 CLK_div_3_mag_0.CLK.n11 VSS 0.288f
C2052 CLK_div_3_mag_0.CLK.t12 VSS 0.0509f
C2053 CLK_div_3_mag_0.CLK.t9 VSS 0.0335f
C2054 CLK_div_3_mag_0.CLK.n12 VSS 0.09f
C2055 CLK_div_3_mag_0.CLK.t10 VSS 0.042f
C2056 CLK_div_3_mag_0.CLK.t15 VSS 0.0109f
C2057 CLK_div_3_mag_0.CLK.n13 VSS 0.0697f
C2058 CLK_div_3_mag_0.CLK.n14 VSS 0.67f
C2059 CLK_div_3_mag_0.CLK.n15 VSS 0.671f
C2060 CLK_div_3_mag_1.Q1.t1 VSS 0.021f
C2061 CLK_div_3_mag_1.Q1.t2 VSS 0.0173f
C2062 CLK_div_3_mag_1.Q1.n0 VSS 0.0173f
C2063 CLK_div_3_mag_1.Q1.n1 VSS 0.0415f
C2064 CLK_div_3_mag_1.Q1.t5 VSS 0.0276f
C2065 CLK_div_3_mag_1.Q1.t6 VSS 0.0221f
C2066 CLK_div_3_mag_1.Q1.n2 VSS 0.0625f
C2067 CLK_div_3_mag_1.Q1.t4 VSS 0.0277f
C2068 CLK_div_3_mag_1.Q1.t10 VSS 0.0355f
C2069 CLK_div_3_mag_1.Q1.n3 VSS 0.0706f
C2070 CLK_div_3_mag_1.Q1.n4 VSS 0.321f
C2071 CLK_div_3_mag_1.Q1.t7 VSS 0.0385f
C2072 CLK_div_3_mag_1.Q1.t3 VSS 0.0254f
C2073 CLK_div_3_mag_1.Q1.n5 VSS 0.0684f
C2074 CLK_div_3_mag_1.Q1.t9 VSS 0.0276f
C2075 CLK_div_3_mag_1.Q1.t8 VSS 0.0221f
C2076 CLK_div_3_mag_1.Q1.n6 VSS 0.0642f
C2077 CLK_div_3_mag_1.Q1.n7 VSS 0.505f
C2078 CLK_div_3_mag_1.Q1.n8 VSS 0.209f
C2079 CLK_div_3_mag_1.JK_FF_mag_1.K.n0 VSS 2.07f
C2080 CLK_div_3_mag_1.JK_FF_mag_1.K.t0 VSS 0.0344f
C2081 CLK_div_3_mag_1.JK_FF_mag_1.K.n1 VSS 0.0344f
C2082 CLK_div_3_mag_1.JK_FF_mag_1.K.n2 VSS 0.0734f
C2083 CLK_div_3_mag_1.JK_FF_mag_1.K.t4 VSS 0.0774f
C2084 CLK_div_3_mag_1.JK_FF_mag_1.K.t2 VSS 0.0493f
C2085 CLK_div_3_mag_1.JK_FF_mag_1.K.n3 VSS 0.137f
C2086 CLK_div_3_mag_1.JK_FF_mag_1.K.t7 VSS 0.0552f
C2087 CLK_div_3_mag_1.JK_FF_mag_1.K.t5 VSS 0.0708f
C2088 CLK_div_3_mag_1.JK_FF_mag_1.K.n4 VSS 0.141f
C2089 CLK_div_3_mag_1.JK_FF_mag_1.K.t3 VSS 0.055f
C2090 CLK_div_3_mag_1.JK_FF_mag_1.K.t6 VSS 0.044f
C2091 CLK_div_3_mag_1.JK_FF_mag_1.K.n5 VSS 0.131f
C2092 CLK_div_3_mag_1.JK_FF_mag_1.K.n6 VSS 1.18f
C2093 CLK_div_3_mag_1.JK_FF_mag_1.K.n7 VSS 0.215f
C2094 CLK_div_3_mag_1.Q0.t1 VSS 0.025f
C2095 CLK_div_3_mag_1.Q0.t2 VSS 0.0206f
C2096 CLK_div_3_mag_1.Q0.n0 VSS 0.0206f
C2097 CLK_div_3_mag_1.Q0.n1 VSS 0.0494f
C2098 CLK_div_3_mag_1.Q0.t8 VSS 0.0459f
C2099 CLK_div_3_mag_1.Q0.t7 VSS 0.0302f
C2100 CLK_div_3_mag_1.Q0.n2 VSS 0.0814f
C2101 CLK_div_3_mag_1.Q0.t4 VSS 0.0329f
C2102 CLK_div_3_mag_1.Q0.t3 VSS 0.0263f
C2103 CLK_div_3_mag_1.Q0.n3 VSS 0.0764f
C2104 CLK_div_3_mag_1.Q0.n4 VSS 0.606f
C2105 CLK_div_3_mag_1.Q0.t6 VSS 0.0641f
C2106 CLK_div_3_mag_1.Q0.t5 VSS 0.0199f
C2107 CLK_div_3_mag_1.Q0.n5 VSS 0.0675f
C2108 CLK_div_3_mag_1.Q0.n6 VSS 0.447f
C2109 CLK_div_3_mag_0.JK_FF_mag_1.K.n0 VSS 2.07f
C2110 CLK_div_3_mag_0.JK_FF_mag_1.K.t0 VSS 0.0344f
C2111 CLK_div_3_mag_0.JK_FF_mag_1.K.n1 VSS 0.0344f
C2112 CLK_div_3_mag_0.JK_FF_mag_1.K.n2 VSS 0.0734f
C2113 CLK_div_3_mag_0.JK_FF_mag_1.K.t6 VSS 0.0774f
C2114 CLK_div_3_mag_0.JK_FF_mag_1.K.t5 VSS 0.0493f
C2115 CLK_div_3_mag_0.JK_FF_mag_1.K.n3 VSS 0.137f
C2116 CLK_div_3_mag_0.JK_FF_mag_1.K.t3 VSS 0.0552f
C2117 CLK_div_3_mag_0.JK_FF_mag_1.K.t7 VSS 0.0708f
C2118 CLK_div_3_mag_0.JK_FF_mag_1.K.n4 VSS 0.141f
C2119 CLK_div_3_mag_0.JK_FF_mag_1.K.t4 VSS 0.055f
C2120 CLK_div_3_mag_0.JK_FF_mag_1.K.t2 VSS 0.044f
C2121 CLK_div_3_mag_0.JK_FF_mag_1.K.n5 VSS 0.131f
C2122 CLK_div_3_mag_0.JK_FF_mag_1.K.n6 VSS 1.18f
C2123 CLK_div_3_mag_0.JK_FF_mag_1.K.n7 VSS 0.215f
C2124 VDD.n0 VSS 0.0068f
C2125 VDD.n1 VSS 0.228f
C2126 VDD.t352 VSS 0.00679f
C2127 VDD.n2 VSS 0.0068f
C2128 VDD.n3 VSS 0.222f
C2129 VDD.t368 VSS 0.00679f
C2130 VDD.n4 VSS 0.0068f
C2131 VDD.n5 VSS 0.0068f
C2132 VDD.n6 VSS 0.0268f
C2133 VDD.t323 VSS 0.00279f
C2134 VDD.n7 VSS 0.00279f
C2135 VDD.n8 VSS 0.0061f
C2136 VDD.n9 VSS 0.024f
C2137 VDD.n10 VSS 0.0686f
C2138 VDD.n11 VSS 0.00685f
C2139 VDD.t235 VSS 0.0601f
C2140 VDD.t424 VSS 0.1f
C2141 VDD.t322 VSS 0.0463f
C2142 VDD.n12 VSS 0.0158f
C2143 VDD.n13 VSS 0.0422f
C2144 VDD.t133 VSS 0.0466f
C2145 VDD.n14 VSS 0.0631f
C2146 VDD.n15 VSS 0.0907f
C2147 VDD.n16 VSS 0.00677f
C2148 VDD.n17 VSS 0.0221f
C2149 VDD.t288 VSS 0.0534f
C2150 VDD.t33 VSS 0.0613f
C2151 VDD.t289 VSS 0.00679f
C2152 VDD.n18 VSS 0.0068f
C2153 VDD.n19 VSS 0.211f
C2154 VDD.t103 VSS 0.00679f
C2155 VDD.t89 VSS 0.0821f
C2156 VDD.n20 VSS 0.195f
C2157 VDD.n21 VSS 0.0068f
C2158 VDD.t78 VSS 0.00679f
C2159 VDD.n22 VSS 0.175f
C2160 VDD.t381 VSS 0.0466f
C2161 VDD.n23 VSS 0.00693f
C2162 VDD.n24 VSS 0.00709f
C2163 VDD.t82 VSS 0.0601f
C2164 VDD.n25 VSS 0.0631f
C2165 VDD.n26 VSS 0.211f
C2166 VDD.t86 VSS 0.00279f
C2167 VDD.n27 VSS 0.00279f
C2168 VDD.n28 VSS 0.0061f
C2169 VDD.n29 VSS 0.0068f
C2170 VDD.n30 VSS 0.0237f
C2171 VDD.n31 VSS 0.903f
C2172 VDD.n32 VSS 0.0714f
C2173 VDD.n33 VSS 0.0251f
C2174 VDD.n34 VSS 0.0144f
C2175 VDD.n35 VSS 0.0422f
C2176 VDD.t85 VSS 0.0463f
C2177 VDD.t104 VSS 0.1f
C2178 VDD.t179 VSS 0.0821f
C2179 VDD.t77 VSS 0.0896f
C2180 VDD.n36 VSS 0.0422f
C2181 VDD.n37 VSS 0.0183f
C2182 VDD.n38 VSS 0.0638f
C2183 VDD.n39 VSS 0.0293f
C2184 VDD.n40 VSS 0.0272f
C2185 VDD.n41 VSS 0.0612f
C2186 VDD.t200 VSS 0.00679f
C2187 VDD.n42 VSS 0.00693f
C2188 VDD.n43 VSS 0.0896f
C2189 VDD.n44 VSS 0.0308f
C2190 VDD.n45 VSS 0.0235f
C2191 VDD.n46 VSS 0.0422f
C2192 VDD.t199 VSS 0.0896f
C2193 VDD.t432 VSS 0.0821f
C2194 VDD.t102 VSS 0.0883f
C2195 VDD.n47 VSS 0.0422f
C2196 VDD.n48 VSS 0.0235f
C2197 VDD.n49 VSS 0.0307f
C2198 VDD.t325 VSS 0.00679f
C2199 VDD.t79 VSS 0.0821f
C2200 VDD.n50 VSS 0.0068f
C2201 VDD.t371 VSS 0.00279f
C2202 VDD.n51 VSS 0.00279f
C2203 VDD.n52 VSS 0.0061f
C2204 VDD.n53 VSS 0.0068f
C2205 VDD.n54 VSS 0.0397f
C2206 VDD.t164 VSS 0.0819f
C2207 VDD.n55 VSS 6.72e-19
C2208 VDD.t507 VSS 0.00442f
C2209 VDD.t151 VSS 0.00583f
C2210 VDD.n56 VSS 0.0114f
C2211 VDD.n57 VSS 0.0757f
C2212 VDD.n58 VSS 0.0748f
C2213 VDD.t510 VSS 0.00442f
C2214 VDD.t163 VSS 0.00572f
C2215 VDD.n59 VSS 0.00543f
C2216 VDD.n60 VSS 0.00607f
C2217 VDD.n61 VSS 9.6e-19
C2218 VDD.n62 VSS 0.00507f
C2219 VDD.n63 VSS 0.00635f
C2220 VDD.n64 VSS 0.0159f
C2221 VDD.t66 VSS 0.00279f
C2222 VDD.n65 VSS 0.00279f
C2223 VDD.n66 VSS 0.0061f
C2224 VDD.n67 VSS 0.0388f
C2225 VDD.n68 VSS 0.0388f
C2226 VDD.n69 VSS 0.0422f
C2227 VDD.t65 VSS 0.0463f
C2228 VDD.t285 VSS 0.1f
C2229 VDD.t69 VSS 0.0821f
C2230 VDD.t92 VSS 0.1f
C2231 VDD.t370 VSS 0.0463f
C2232 VDD.n70 VSS 0.0422f
C2233 VDD.n71 VSS 0.021f
C2234 VDD.n72 VSS 0.0388f
C2235 VDD.n73 VSS 0.0396f
C2236 VDD.t202 VSS 0.00679f
C2237 VDD.n74 VSS 0.0068f
C2238 VDD.n75 VSS 0.0312f
C2239 VDD.n76 VSS 0.0337f
C2240 VDD.n77 VSS 0.0235f
C2241 VDD.n78 VSS 0.0422f
C2242 VDD.t201 VSS 0.0896f
C2243 VDD.t8 VSS 0.0821f
C2244 VDD.t324 VSS 0.0883f
C2245 VDD.n79 VSS 0.0422f
C2246 VDD.n80 VSS 0.0235f
C2247 VDD.n81 VSS 0.0587f
C2248 VDD.n82 VSS 0.00677f
C2249 VDD.n83 VSS 0.0068f
C2250 VDD.n84 VSS 0.0299f
C2251 VDD.t40 VSS 0.0601f
C2252 VDD.n85 VSS 0.0157f
C2253 VDD.t295 VSS 0.0896f
C2254 VDD.n86 VSS 0.0068f
C2255 VDD.t44 VSS 0.00279f
C2256 VDD.n87 VSS 0.00279f
C2257 VDD.n88 VSS 0.0061f
C2258 VDD.n89 VSS 0.053f
C2259 VDD.n90 VSS 0.0219f
C2260 VDD.n91 VSS 0.0296f
C2261 VDD.t296 VSS 0.00679f
C2262 VDD.n92 VSS 0.0068f
C2263 VDD.t332 VSS 0.0821f
C2264 VDD.n93 VSS 0.0422f
C2265 VDD.t39 VSS 0.00679f
C2266 VDD.n94 VSS 0.0068f
C2267 VDD.t38 VSS 0.0896f
C2268 VDD.t466 VSS 0.0821f
C2269 VDD.t231 VSS 0.0883f
C2270 VDD.n95 VSS 0.0422f
C2271 VDD.t232 VSS 0.00679f
C2272 VDD.t142 VSS 0.00679f
C2273 VDD.t292 VSS 0.0821f
C2274 VDD.n96 VSS 0.0068f
C2275 VDD.t22 VSS 0.00279f
C2276 VDD.n97 VSS 0.00279f
C2277 VDD.n98 VSS 0.0061f
C2278 VDD.n99 VSS 0.0068f
C2279 VDD.n100 VSS 0.0397f
C2280 VDD.t152 VSS 0.0819f
C2281 VDD.n101 VSS 0.00729f
C2282 VDD.t49 VSS 0.00279f
C2283 VDD.n102 VSS 0.00279f
C2284 VDD.n103 VSS 0.0061f
C2285 VDD.n104 VSS 0.0388f
C2286 VDD.n105 VSS 0.0523f
C2287 VDD.n106 VSS 0.0422f
C2288 VDD.t48 VSS 0.0463f
C2289 VDD.t144 VSS 0.1f
C2290 VDD.t5 VSS 0.0821f
C2291 VDD.t329 VSS 0.1f
C2292 VDD.t21 VSS 0.0463f
C2293 VDD.n107 VSS 0.0422f
C2294 VDD.n108 VSS 0.021f
C2295 VDD.n109 VSS 0.0388f
C2296 VDD.n110 VSS 0.0396f
C2297 VDD.t37 VSS 0.00679f
C2298 VDD.n111 VSS 0.0068f
C2299 VDD.n112 VSS 0.0312f
C2300 VDD.n113 VSS 0.0337f
C2301 VDD.n114 VSS 0.0235f
C2302 VDD.n115 VSS 0.0422f
C2303 VDD.t36 VSS 0.0896f
C2304 VDD.t228 VSS 0.0821f
C2305 VDD.t141 VSS 0.0883f
C2306 VDD.n116 VSS 0.0422f
C2307 VDD.n117 VSS 0.0235f
C2308 VDD.n118 VSS 0.064f
C2309 VDD.n119 VSS 0.0727f
C2310 VDD.n120 VSS 0.0235f
C2311 VDD.n121 VSS 0.0312f
C2312 VDD.n122 VSS 0.0337f
C2313 VDD.n123 VSS 0.0235f
C2314 VDD.n124 VSS 0.0312f
C2315 VDD.n125 VSS 0.0337f
C2316 VDD.n126 VSS 0.0235f
C2317 VDD.n127 VSS 0.0422f
C2318 VDD.t196 VSS 0.0821f
C2319 VDD.t378 VSS 0.1f
C2320 VDD.t43 VSS 0.0463f
C2321 VDD.n128 VSS 0.0422f
C2322 VDD.t326 VSS 0.0466f
C2323 VDD.n129 VSS 0.0631f
C2324 VDD.n130 VSS 0.0213f
C2325 VDD.n131 VSS 0.0406f
C2326 VDD.n132 VSS 0.0667f
C2327 VDD.n133 VSS 0.248f
C2328 VDD.n134 VSS 0.195f
C2329 VDD.n135 VSS 0.0533f
C2330 VDD.t45 VSS 0.0819f
C2331 VDD.n136 VSS 0.0422f
C2332 VDD.n137 VSS 0.0455f
C2333 VDD.n138 VSS 0.0941f
C2334 VDD.n139 VSS 0.00853f
C2335 VDD.n140 VSS 0.0162f
C2336 VDD.n141 VSS 0.0957f
C2337 VDD.n142 VSS 0.0677f
C2338 VDD.n143 VSS 0.106f
C2339 VDD.t184 VSS 0.0578f
C2340 VDD.t72 VSS 0.0604f
C2341 VDD.n144 VSS 0.0698f
C2342 VDD.t143 VSS 0.0608f
C2343 VDD.n145 VSS 0.041f
C2344 VDD.n146 VSS 0.0707f
C2345 VDD.n147 VSS 0.166f
C2346 VDD.n148 VSS 0.196f
C2347 VDD.n149 VSS 0.19f
C2348 VDD.n150 VSS 0.207f
C2349 VDD.n151 VSS 0.0695f
C2350 VDD.n152 VSS 0.0209f
C2351 VDD.t125 VSS 0.0821f
C2352 VDD.t367 VSS 0.0896f
C2353 VDD.n153 VSS 0.0422f
C2354 VDD.n154 VSS 0.0235f
C2355 VDD.n155 VSS 0.0247f
C2356 VDD.n156 VSS 0.0668f
C2357 VDD.n157 VSS 0.0276f
C2358 VDD.t50 VSS 0.0821f
C2359 VDD.t351 VSS 0.0896f
C2360 VDD.n158 VSS 0.0422f
C2361 VDD.n159 VSS 0.0235f
C2362 VDD.n160 VSS 0.0263f
C2363 VDD.n161 VSS 0.0668f
C2364 VDD.n162 VSS 0.026f
C2365 VDD.t107 VSS 0.0821f
C2366 VDD.t422 VSS 0.0883f
C2367 VDD.n163 VSS 0.0422f
C2368 VDD.t423 VSS 0.00679f
C2369 VDD.t137 VSS 0.00679f
C2370 VDD.t364 VSS 0.0821f
C2371 VDD.n164 VSS 0.0068f
C2372 VDD.t20 VSS 0.00279f
C2373 VDD.n165 VSS 0.00279f
C2374 VDD.n166 VSS 0.0061f
C2375 VDD.n167 VSS 0.0068f
C2376 VDD.n168 VSS 0.0397f
C2377 VDD.t156 VSS 0.0819f
C2378 VDD.n169 VSS 9.16e-19
C2379 VDD.t511 VSS 0.00442f
C2380 VDD.t159 VSS 0.00583f
C2381 VDD.n170 VSS 0.0114f
C2382 VDD.n171 VSS 0.0757f
C2383 VDD.t513 VSS 0.00442f
C2384 VDD.n172 VSS 0.00607f
C2385 VDD.t155 VSS 0.00572f
C2386 VDD.n173 VSS 0.00543f
C2387 VDD.n174 VSS 0.0743f
C2388 VDD.n175 VSS 0.00328f
C2389 VDD.n176 VSS 0.00635f
C2390 VDD.n177 VSS 0.0179f
C2391 VDD.t12 VSS 0.00279f
C2392 VDD.n178 VSS 0.00279f
C2393 VDD.n179 VSS 0.0061f
C2394 VDD.n180 VSS 0.0388f
C2395 VDD.n181 VSS 0.0388f
C2396 VDD.n182 VSS 0.0422f
C2397 VDD.t11 VSS 0.0463f
C2398 VDD.t359 VSS 0.1f
C2399 VDD.t222 VSS 0.0821f
C2400 VDD.t53 VSS 0.1f
C2401 VDD.t19 VSS 0.0463f
C2402 VDD.n183 VSS 0.0422f
C2403 VDD.n184 VSS 0.021f
C2404 VDD.n185 VSS 0.0388f
C2405 VDD.n186 VSS 0.0396f
C2406 VDD.t354 VSS 0.00679f
C2407 VDD.n187 VSS 0.0068f
C2408 VDD.n188 VSS 0.0312f
C2409 VDD.n189 VSS 0.0337f
C2410 VDD.n190 VSS 0.0235f
C2411 VDD.n191 VSS 0.0422f
C2412 VDD.t353 VSS 0.0896f
C2413 VDD.t95 VSS 0.0821f
C2414 VDD.t136 VSS 0.0883f
C2415 VDD.n192 VSS 0.0422f
C2416 VDD.n193 VSS 0.0235f
C2417 VDD.n194 VSS 0.0601f
C2418 VDD.n195 VSS 0.0427f
C2419 VDD.n196 VSS 0.0068f
C2420 VDD.t13 VSS 0.0819f
C2421 VDD.n197 VSS 0.0422f
C2422 VDD.t358 VSS 0.00679f
C2423 VDD.t357 VSS 0.0534f
C2424 VDD.t375 VSS 0.0613f
C2425 VDD.n198 VSS 0.106f
C2426 VDD.n199 VSS 0.00853f
C2427 VDD.n200 VSS 0.0162f
C2428 VDD.t225 VSS 0.0578f
C2429 VDD.n201 VSS 0.041f
C2430 VDD.n202 VSS 0.00677f
C2431 VDD.t315 VSS 0.0608f
C2432 VDD.t341 VSS 0.0604f
C2433 VDD.n203 VSS 0.0698f
C2434 VDD.n204 VSS 0.0221f
C2435 VDD.t116 VSS 0.0068f
C2436 VDD.n205 VSS 0.00679f
C2437 VDD.n206 VSS 0.0334f
C2438 VDD.t283 VSS 0.0799f
C2439 VDD.t115 VSS 0.0657f
C2440 VDD.t304 VSS 0.0329f
C2441 VDD.t284 VSS 0.00677f
C2442 VDD.n207 VSS 0.0239f
C2443 VDD.n208 VSS 0.0659f
C2444 VDD.n209 VSS 0.0478f
C2445 VDD.n210 VSS 0.0303f
C2446 VDD.t148 VSS 0.00677f
C2447 VDD.n211 VSS 0.031f
C2448 VDD.t147 VSS 0.064f
C2449 VDD.n212 VSS 0.0725f
C2450 VDD.t384 VSS 0.0759f
C2451 VDD.t218 VSS 0.0762f
C2452 VDD.n213 VSS 0.0479f
C2453 VDD.t219 VSS 0.0178f
C2454 VDD.n214 VSS 0.103f
C2455 VDD.t246 VSS 0.00677f
C2456 VDD.n215 VSS 0.0312f
C2457 VDD.t245 VSS 0.064f
C2458 VDD.n216 VSS 0.0725f
C2459 VDD.t369 VSS 0.0759f
C2460 VDD.t344 VSS 0.0762f
C2461 VDD.n217 VSS 0.0479f
C2462 VDD.t345 VSS 0.0178f
C2463 VDD.n218 VSS 0.104f
C2464 VDD.t403 VSS 0.00649f
C2465 VDD.t485 VSS 0.0141f
C2466 VDD.n219 VSS 0.201f
C2467 VDD.t251 VSS 0.0068f
C2468 VDD.t441 VSS 0.00279f
C2469 VDD.n220 VSS 0.00279f
C2470 VDD.n221 VSS 0.0061f
C2471 VDD.t121 VSS 0.0068f
C2472 VDD.n222 VSS 0.00679f
C2473 VDD.n223 VSS 0.16f
C2474 VDD.t192 VSS 0.0799f
C2475 VDD.t120 VSS 0.0657f
C2476 VDD.t247 VSS 0.0329f
C2477 VDD.t193 VSS 0.00854f
C2478 VDD.t356 VSS 0.0148f
C2479 VDD.t500 VSS 0.0131f
C2480 VDD.n224 VSS 0.121f
C2481 VDD.t499 VSS 0.0447f
C2482 VDD.t87 VSS 0.0869f
C2483 VDD.t88 VSS 0.0141f
C2484 VDD.n225 VSS -0.207f
C2485 VDD.t150 VSS 0.0068f
C2486 VDD.t149 VSS 0.0801f
C2487 VDD.n226 VSS 0.0527f
C2488 VDD.t309 VSS 0.165f
C2489 VDD.t451 VSS 0.0551f
C2490 VDD.t416 VSS 0.04f
C2491 VDD.n227 VSS 0.0374f
C2492 VDD.n228 VSS 0.0639f
C2493 VDD.t415 VSS 0.175f
C2494 VDD.n229 VSS 0.0991f
C2495 VDD.n230 VSS 0.156f
C2496 VDD.n231 VSS 0.0904f
C2497 VDD.n232 VSS 0.0958f
C2498 VDD.t355 VSS 0.0476f
C2499 VDD.n233 VSS 0.0633f
C2500 VDD.n234 VSS 0.196f
C2501 VDD.n235 VSS 0.0659f
C2502 VDD.n236 VSS 0.0943f
C2503 VDD.n237 VSS 0.201f
C2504 VDD.n238 VSS 0.212f
C2505 VDD.t440 VSS 0.0657f
C2506 VDD.t250 VSS 0.0657f
C2507 VDD.t212 VSS 0.0495f
C2508 VDD.n239 VSS 0.0511f
C2509 VDD.n240 VSS 0.228f
C2510 VDD.t484 VSS 0.0674f
C2511 VDD.t402 VSS 0.081f
C2512 VDD.n241 VSS 0.0703f
C2513 VDD.n242 VSS 0.114f
C2514 VDD.n243 VSS 0.126f
C2515 VDD.t431 VSS 0.00279f
C2516 VDD.n244 VSS 0.00279f
C2517 VDD.n245 VSS 0.0061f
C2518 VDD.n246 VSS 0.0262f
C2519 VDD.t278 VSS 0.0897f
C2520 VDD.n247 VSS 0.00679f
C2521 VDD.t258 VSS 0.0068f
C2522 VDD.n248 VSS 0.00679f
C2523 VDD.n249 VSS 0.0371f
C2524 VDD.t427 VSS 0.0885f
C2525 VDD.n250 VSS 0.00679f
C2526 VDD.n251 VSS 0.00679f
C2527 VDD.t404 VSS 0.0885f
C2528 VDD.n252 VSS 0.0422f
C2529 VDD.t340 VSS 0.0068f
C2530 VDD.n253 VSS 0.00679f
C2531 VDD.t339 VSS 0.0819f
C2532 VDD.t504 VSS 0.0897f
C2533 VDD.n254 VSS 0.0422f
C2534 VDD.t277 VSS 0.0068f
C2535 VDD.t260 VSS 0.00279f
C2536 VDD.n255 VSS 0.00279f
C2537 VDD.n256 VSS 0.0061f
C2538 VDD.t276 VSS 0.0819f
C2539 VDD.t259 VSS 0.1f
C2540 VDD.t26 VSS 0.0465f
C2541 VDD.n257 VSS 0.0422f
C2542 VDD.t68 VSS 0.0068f
C2543 VDD.t401 VSS 0.00279f
C2544 VDD.n258 VSS 0.00279f
C2545 VDD.n259 VSS 0.0061f
C2546 VDD.t67 VSS 0.0819f
C2547 VDD.t400 VSS 0.1f
C2548 VDD.t437 VSS 0.0465f
C2549 VDD.t297 VSS 0.0817f
C2550 VDD.n260 VSS 0.0422f
C2551 VDD.t298 VSS 0.00728f
C2552 VDD.n261 VSS 0.0523f
C2553 VDD.n262 VSS 0.0387f
C2554 VDD.n263 VSS 0.0397f
C2555 VDD.n264 VSS 0.0211f
C2556 VDD.n265 VSS 0.0387f
C2557 VDD.n266 VSS 0.0396f
C2558 VDD.n267 VSS 0.0235f
C2559 VDD.n268 VSS 0.0337f
C2560 VDD.n269 VSS 0.0313f
C2561 VDD.n270 VSS 0.0235f
C2562 VDD.n271 VSS 0.0589f
C2563 VDD.t446 VSS 0.00677f
C2564 VDD.t412 VSS 0.0068f
C2565 VDD.n272 VSS 0.0394f
C2566 VDD.t445 VSS 0.0599f
C2567 VDD.t442 VSS 0.0465f
C2568 VDD.t456 VSS 0.00279f
C2569 VDD.n273 VSS 0.00279f
C2570 VDD.n274 VSS 0.0061f
C2571 VDD.t76 VSS 0.0068f
C2572 VDD.n275 VSS 0.00679f
C2573 VDD.n276 VSS 0.0368f
C2574 VDD.t390 VSS 0.0897f
C2575 VDD.n277 VSS 0.00679f
C2576 VDD.t471 VSS 0.0068f
C2577 VDD.n278 VSS 0.00679f
C2578 VDD.n279 VSS 0.00679f
C2579 VDD.t112 VSS 0.0885f
C2580 VDD.n280 VSS 0.0422f
C2581 VDD.t291 VSS 0.0068f
C2582 VDD.n281 VSS 0.00679f
C2583 VDD.t290 VSS 0.0819f
C2584 VDD.t387 VSS 0.0897f
C2585 VDD.n282 VSS 0.0422f
C2586 VDD.t275 VSS 0.0068f
C2587 VDD.t32 VSS 0.00279f
C2588 VDD.n283 VSS 0.00279f
C2589 VDD.n284 VSS 0.0061f
C2590 VDD.t274 VSS 0.0819f
C2591 VDD.t31 VSS 0.1f
C2592 VDD.t372 VSS 0.0465f
C2593 VDD.n285 VSS 0.0422f
C2594 VDD.t204 VSS 0.0068f
C2595 VDD.t124 VSS 0.00279f
C2596 VDD.n286 VSS 0.00279f
C2597 VDD.n287 VSS 0.0061f
C2598 VDD.t203 VSS 0.0819f
C2599 VDD.t123 VSS 0.1f
C2600 VDD.t460 VSS 0.0465f
C2601 VDD.t409 VSS 0.0817f
C2602 VDD.n288 VSS 0.0422f
C2603 VDD.t410 VSS 0.00728f
C2604 VDD.n289 VSS 0.0523f
C2605 VDD.n290 VSS 0.0387f
C2606 VDD.n291 VSS 0.0397f
C2607 VDD.n292 VSS 0.0211f
C2608 VDD.n293 VSS 0.0387f
C2609 VDD.n294 VSS 0.0396f
C2610 VDD.n295 VSS 0.0235f
C2611 VDD.n296 VSS 0.0337f
C2612 VDD.n297 VSS 0.0313f
C2613 VDD.n298 VSS 0.0235f
C2614 VDD.n299 VSS 0.0799f
C2615 VDD.t436 VSS 0.00677f
C2616 VDD.t494 VSS 0.0068f
C2617 VDD.n300 VSS 0.04f
C2618 VDD.t435 VSS 0.0599f
C2619 VDD.t457 VSS 0.0465f
C2620 VDD.t175 VSS 0.00279f
C2621 VDD.n301 VSS 0.00279f
C2622 VDD.n302 VSS 0.0061f
C2623 VDD.t206 VSS 0.0068f
C2624 VDD.n303 VSS 0.00679f
C2625 VDD.n304 VSS 0.0374f
C2626 VDD.t472 VSS 0.0897f
C2627 VDD.n305 VSS 0.00679f
C2628 VDD.t168 VSS 0.0068f
C2629 VDD.n306 VSS 0.00679f
C2630 VDD.n307 VSS 0.00679f
C2631 VDD.t215 VSS 0.0885f
C2632 VDD.n308 VSS 0.0422f
C2633 VDD.t101 VSS 0.0068f
C2634 VDD.n309 VSS 0.00679f
C2635 VDD.t100 VSS 0.0819f
C2636 VDD.t475 VSS 0.0897f
C2637 VDD.n310 VSS 0.0422f
C2638 VDD.t188 VSS 0.0068f
C2639 VDD.t264 VSS 0.00279f
C2640 VDD.n311 VSS 0.00279f
C2641 VDD.n312 VSS 0.0061f
C2642 VDD.t187 VSS 0.0819f
C2643 VDD.t263 VSS 0.1f
C2644 VDD.t23 VSS 0.0465f
C2645 VDD.n313 VSS 0.0422f
C2646 VDD.t99 VSS 0.0068f
C2647 VDD.t221 VSS 0.00279f
C2648 VDD.n314 VSS 0.00279f
C2649 VDD.n315 VSS 0.0061f
C2650 VDD.t98 VSS 0.0819f
C2651 VDD.t220 VSS 0.1f
C2652 VDD.t463 VSS 0.0465f
C2653 VDD.t491 VSS 0.0817f
C2654 VDD.n316 VSS 0.0422f
C2655 VDD.t492 VSS 0.00728f
C2656 VDD.n317 VSS 0.0523f
C2657 VDD.n318 VSS 0.0387f
C2658 VDD.n319 VSS 0.0397f
C2659 VDD.n320 VSS 0.0211f
C2660 VDD.n321 VSS 0.0387f
C2661 VDD.n322 VSS 0.0396f
C2662 VDD.n323 VSS 0.0235f
C2663 VDD.n324 VSS 0.0337f
C2664 VDD.n325 VSS 0.0313f
C2665 VDD.n326 VSS 0.0235f
C2666 VDD.n327 VSS 0.0801f
C2667 VDD.n328 VSS 0.0923f
C2668 VDD.t176 VSS 0.0885f
C2669 VDD.t167 VSS 0.0819f
C2670 VDD.n329 VSS 0.0422f
C2671 VDD.n330 VSS 0.0251f
C2672 VDD.n331 VSS 0.0346f
C2673 VDD.n332 VSS 0.0374f
C2674 VDD.t262 VSS 0.0068f
C2675 VDD.n333 VSS 0.0346f
C2676 VDD.n334 VSS 0.0251f
C2677 VDD.n335 VSS 0.0422f
C2678 VDD.t261 VSS 0.0819f
C2679 VDD.t189 VSS 0.0897f
C2680 VDD.t174 VSS 0.1f
C2681 VDD.t205 VSS 0.0819f
C2682 VDD.n336 VSS 0.0422f
C2683 VDD.n337 VSS 0.0251f
C2684 VDD.n338 VSS 0.0326f
C2685 VDD.n339 VSS 0.031f
C2686 VDD.n340 VSS 0.0223f
C2687 VDD.n341 VSS 0.0422f
C2688 VDD.t493 VSS 0.0465f
C2689 VDD.n342 VSS 0.0631f
C2690 VDD.n343 VSS 0.038f
C2691 VDD.n344 VSS 0.0424f
C2692 VDD.n345 VSS 0.0378f
C2693 VDD.t452 VSS 0.0885f
C2694 VDD.t470 VSS 0.0819f
C2695 VDD.n346 VSS 0.0422f
C2696 VDD.n347 VSS 0.0248f
C2697 VDD.n348 VSS 0.0341f
C2698 VDD.n349 VSS 0.0368f
C2699 VDD.t30 VSS 0.0068f
C2700 VDD.n350 VSS 0.0341f
C2701 VDD.n351 VSS 0.0248f
C2702 VDD.n352 VSS 0.0422f
C2703 VDD.t29 VSS 0.0819f
C2704 VDD.t271 VSS 0.0897f
C2705 VDD.t455 VSS 0.1f
C2706 VDD.t75 VSS 0.0819f
C2707 VDD.n353 VSS 0.0422f
C2708 VDD.n354 VSS 0.0248f
C2709 VDD.n355 VSS 0.0322f
C2710 VDD.n356 VSS 0.0305f
C2711 VDD.n357 VSS 0.0221f
C2712 VDD.n358 VSS 0.0422f
C2713 VDD.t411 VSS 0.0465f
C2714 VDD.n359 VSS 0.0631f
C2715 VDD.n360 VSS 0.0364f
C2716 VDD.n361 VSS 0.0597f
C2717 VDD.n362 VSS 0.0362f
C2718 VDD.t386 VSS 0.0068f
C2719 VDD.n363 VSS 0.0343f
C2720 VDD.n364 VSS 0.025f
C2721 VDD.n365 VSS 0.0422f
C2722 VDD.t385 VSS 0.0819f
C2723 VDD.t501 VSS 0.0897f
C2724 VDD.t257 VSS 0.0819f
C2725 VDD.n366 VSS 0.0422f
C2726 VDD.n367 VSS 0.025f
C2727 VDD.n368 VSS 0.0343f
C2728 VDD.n369 VSS 0.0371f
C2729 VDD.t338 VSS 0.0068f
C2730 VDD.n370 VSS 0.0324f
C2731 VDD.n371 VSS 0.025f
C2732 VDD.n372 VSS 0.0422f
C2733 VDD.t337 VSS 0.0819f
C2734 VDD.t430 VSS 0.1f
C2735 VDD.t59 VSS 0.0465f
C2736 VDD.n373 VSS 0.0422f
C2737 VDD.t244 VSS 0.0068f
C2738 VDD.t243 VSS 0.0465f
C2739 VDD.t417 VSS 0.0599f
C2740 VDD.n374 VSS 0.0631f
C2741 VDD.t418 VSS 0.00677f
C2742 VDD.n375 VSS 0.00679f
C2743 VDD.t301 VSS 0.0885f
C2744 VDD.n376 VSS 0.0422f
C2745 VDD.t183 VSS 0.0068f
C2746 VDD.n377 VSS 0.00679f
C2747 VDD.t182 VSS 0.0819f
C2748 VDD.t316 VSS 0.0897f
C2749 VDD.n378 VSS 0.0422f
C2750 VDD.t170 VSS 0.0068f
C2751 VDD.t496 VSS 0.00279f
C2752 VDD.n379 VSS 0.00279f
C2753 VDD.n380 VSS 0.0061f
C2754 VDD.t169 VSS 0.0819f
C2755 VDD.t495 VSS 0.1f
C2756 VDD.t397 VSS 0.0465f
C2757 VDD.n381 VSS 0.0422f
C2758 VDD.t394 VSS 0.0068f
C2759 VDD.t308 VSS 0.00279f
C2760 VDD.n382 VSS 0.00279f
C2761 VDD.n383 VSS 0.0061f
C2762 VDD.t393 VSS 0.0819f
C2763 VDD.t307 VSS 0.1f
C2764 VDD.t254 VSS 0.0465f
C2765 VDD.t265 VSS 0.0817f
C2766 VDD.n384 VSS 0.0422f
C2767 VDD.t266 VSS 0.00728f
C2768 VDD.n385 VSS 0.0523f
C2769 VDD.n386 VSS 0.0387f
C2770 VDD.n387 VSS 0.0397f
C2771 VDD.n388 VSS 0.0211f
C2772 VDD.n389 VSS 0.0387f
C2773 VDD.n390 VSS 0.0396f
C2774 VDD.n391 VSS 0.0235f
C2775 VDD.n392 VSS 0.0337f
C2776 VDD.n393 VSS 0.0313f
C2777 VDD.n394 VSS 0.0235f
C2778 VDD.n395 VSS 0.0589f
C2779 VDD.n396 VSS 0.00679f
C2780 VDD.t348 VSS 0.0885f
C2781 VDD.n397 VSS 0.0422f
C2782 VDD.t336 VSS 0.0068f
C2783 VDD.n398 VSS 0.00679f
C2784 VDD.t335 VSS 0.0819f
C2785 VDD.t319 VSS 0.0897f
C2786 VDD.n399 VSS 0.0422f
C2787 VDD.t498 VSS 0.0068f
C2788 VDD.n400 VSS 0.00679f
C2789 VDD.t497 VSS 0.0819f
C2790 VDD.t171 VSS 0.0897f
C2791 VDD.n401 VSS 0.0422f
C2792 VDD.t253 VSS 0.0068f
C2793 VDD.t347 VSS 0.00279f
C2794 VDD.n402 VSS 0.00279f
C2795 VDD.n403 VSS 0.0061f
C2796 VDD.t252 VSS 0.0819f
C2797 VDD.t346 VSS 0.1f
C2798 VDD.t56 VSS 0.0465f
C2799 VDD.n404 VSS 0.0422f
C2800 VDD.t268 VSS 0.0068f
C2801 VDD.t267 VSS 0.0465f
C2802 VDD.t413 VSS 0.0599f
C2803 VDD.n405 VSS 0.0594f
C2804 VDD.n406 VSS 0.0561f
C2805 VDD.t414 VSS 0.00677f
C2806 VDD.n407 VSS 0.0344f
C2807 VDD.t363 VSS 0.00677f
C2808 VDD.n408 VSS 0.00679f
C2809 VDD.t362 VSS 0.065f
C2810 VDD.n409 VSS 0.0617f
C2811 VDD.t117 VSS 0.0532f
C2812 VDD.t207 VSS 0.0817f
C2813 VDD.n410 VSS 0.0422f
C2814 VDD.t1 VSS 0.00677f
C2815 VDD.n411 VSS 0.0222f
C2816 VDD.n412 VSS 0.0726f
C2817 VDD.t195 VSS 0.0162f
C2818 VDD.t282 VSS 0.00677f
C2819 VDD.t408 VSS 0.00279f
C2820 VDD.n413 VSS 0.00279f
C2821 VDD.n414 VSS 0.0061f
C2822 VDD.n415 VSS 0.00679f
C2823 VDD.n416 VSS 0.0509f
C2824 VDD.t270 VSS 0.00677f
C2825 VDD.t110 VSS 0.163f
C2826 VDD.t122 VSS 0.0068f
C2827 VDD.t111 VSS 0.0068f
C2828 VDD.n417 VSS 0.0626f
C2829 VDD.n418 VSS 0.0286f
C2830 VDD.n419 VSS 0.0843f
C2831 VDD.t209 VSS 0.0929f
C2832 VDD.t407 VSS 0.128f
C2833 VDD.t194 VSS 0.0218f
C2834 VDD.t269 VSS 0.0903f
C2835 VDD.t0 VSS 0.0602f
C2836 VDD.n421 VSS 0.0713f
C2837 VDD.t469 VSS 0.0568f
C2838 VDD.n422 VSS 0.0243f
C2839 VDD.n423 VSS 0.0854f
C2840 VDD.n424 VSS 0.0505f
C2841 VDD.n425 VSS 0.024f
C2842 VDD.n426 VSS 0.013f
C2843 VDD.n427 VSS 0.0706f
C2844 VDD.t281 VSS 0.0833f
C2845 VDD.n428 VSS 0.0579f
C2846 VDD.n429 VSS 0.0305f
C2847 VDD.n430 VSS 0.0338f
C2848 VDD.n431 VSS 0.0261f
C2849 VDD.t208 VSS 0.0069f
C2850 VDD.n432 VSS 0.0378f
C2851 VDD.n433 VSS 0.0238f
C2852 VDD.n434 VSS 0.0334f
C2853 VDD.n435 VSS 0.0313f
C2854 VDD.n436 VSS 0.028f
C2855 VDD.n437 VSS 0.0348f
C2856 VDD.n438 VSS 0.0221f
C2857 VDD.n439 VSS 0.0305f
C2858 VDD.n440 VSS 0.0322f
C2859 VDD.n441 VSS 0.0248f
C2860 VDD.n442 VSS 0.0368f
C2861 VDD.n443 VSS 0.0341f
C2862 VDD.n444 VSS 0.0248f
C2863 VDD.n445 VSS 0.0368f
C2864 VDD.n446 VSS 0.0341f
C2865 VDD.n447 VSS 0.0248f
C2866 VDD.n448 VSS 0.036f
C2867 VDD.n449 VSS 0.0604f
C2868 VDD.n450 VSS 0.0378f
C2869 VDD.n451 VSS 0.0397f
C2870 VDD.n452 VSS 0.0222f
C2871 VDD.n453 VSS 0.104f
C2872 VDD.n454 VSS 1.28f
C2873 VDD.n455 VSS 0.637f
C2874 VDD.n456 VSS 0.601f
C2875 VDD.n457 VSS 2.22f
C2876 VDD.n458 VSS 1.4f
C2877 VDD.n459 VSS 0.0707f
C2878 VDD.n460 VSS 0.0957f
C2879 VDD.n461 VSS 0.0677f
C2880 VDD.n462 VSS 0.0941f
C2881 VDD.n463 VSS 0.0455f
C2882 VDD.n464 VSS 0.0533f
C2883 VDD.t239 VSS 0.00279f
C2884 VDD.n465 VSS 0.00279f
C2885 VDD.n466 VSS 0.0061f
C2886 VDD.n467 VSS 0.0219f
C2887 VDD.n468 VSS 0.0157f
C2888 VDD.n469 VSS 0.0068f
C2889 VDD.n470 VSS 0.00677f
C2890 VDD.n471 VSS 0.0213f
C2891 VDD.t240 VSS 0.0601f
C2892 VDD.n472 VSS 0.0068f
C2893 VDD.n473 VSS 0.0296f
C2894 VDD.n474 VSS 0.0235f
C2895 VDD.n475 VSS 0.0068f
C2896 VDD.t487 VSS 0.00679f
C2897 VDD.n476 VSS 0.0337f
C2898 VDD.n477 VSS 0.0312f
C2899 VDD.n478 VSS 0.0235f
C2900 VDD.n479 VSS 0.0068f
C2901 VDD.t450 VSS 0.00679f
C2902 VDD.n480 VSS 0.0337f
C2903 VDD.n481 VSS 0.0312f
C2904 VDD.t129 VSS 0.00679f
C2905 VDD.t311 VSS 0.00679f
C2906 VDD.t488 VSS 0.0821f
C2907 VDD.n482 VSS 0.0068f
C2908 VDD.t396 VSS 0.00279f
C2909 VDD.n483 VSS 0.00279f
C2910 VDD.n484 VSS 0.0061f
C2911 VDD.n485 VSS 0.0068f
C2912 VDD.n486 VSS 0.0397f
C2913 VDD.t160 VSS 0.0819f
C2914 VDD.n487 VSS 0.00729f
C2915 VDD.t234 VSS 0.00279f
C2916 VDD.n488 VSS 0.00279f
C2917 VDD.n489 VSS 0.0061f
C2918 VDD.n490 VSS 0.0388f
C2919 VDD.n491 VSS 0.0523f
C2920 VDD.n492 VSS 0.0422f
C2921 VDD.t233 VSS 0.0463f
C2922 VDD.t312 VSS 0.1f
C2923 VDD.t419 VSS 0.0821f
C2924 VDD.t478 VSS 0.1f
C2925 VDD.t395 VSS 0.0463f
C2926 VDD.n493 VSS 0.0422f
C2927 VDD.n494 VSS 0.021f
C2928 VDD.n495 VSS 0.0388f
C2929 VDD.n496 VSS 0.0396f
C2930 VDD.t448 VSS 0.00679f
C2931 VDD.n497 VSS 0.0068f
C2932 VDD.n498 VSS 0.0312f
C2933 VDD.n499 VSS 0.0337f
C2934 VDD.n500 VSS 0.0235f
C2935 VDD.n501 VSS 0.0422f
C2936 VDD.t447 VSS 0.0896f
C2937 VDD.t16 VSS 0.0821f
C2938 VDD.t310 VSS 0.0883f
C2939 VDD.n502 VSS 0.0422f
C2940 VDD.n503 VSS 0.0235f
C2941 VDD.n504 VSS 0.064f
C2942 VDD.n505 VSS 0.0727f
C2943 VDD.n506 VSS 0.0235f
C2944 VDD.t128 VSS 0.0883f
C2945 VDD.n507 VSS 0.0422f
C2946 VDD.t62 VSS 0.0821f
C2947 VDD.t449 VSS 0.0896f
C2948 VDD.n508 VSS 0.0422f
C2949 VDD.t481 VSS 0.0821f
C2950 VDD.t486 VSS 0.0896f
C2951 VDD.n509 VSS 0.0422f
C2952 VDD.t2 VSS 0.0821f
C2953 VDD.t130 VSS 0.1f
C2954 VDD.t238 VSS 0.0463f
C2955 VDD.n510 VSS 0.0422f
C2956 VDD.t138 VSS 0.0466f
C2957 VDD.n511 VSS 0.0631f
C2958 VDD.n512 VSS 0.0299f
C2959 VDD.n513 VSS 0.053f
C2960 VDD.n514 VSS 0.209f
C2961 VDD.n515 VSS 0.273f
C2962 VDD.n516 VSS 0.068f
C2963 VDD.n517 VSS 0.026f
C2964 VDD.n518 VSS 0.0235f
C2965 CLK_div_3_mag_0.Q0.t2 VSS 0.025f
C2966 CLK_div_3_mag_0.Q0.t0 VSS 0.0206f
C2967 CLK_div_3_mag_0.Q0.n0 VSS 0.0206f
C2968 CLK_div_3_mag_0.Q0.n1 VSS 0.0494f
C2969 CLK_div_3_mag_0.Q0.t5 VSS 0.0459f
C2970 CLK_div_3_mag_0.Q0.t4 VSS 0.0302f
C2971 CLK_div_3_mag_0.Q0.n2 VSS 0.0814f
C2972 CLK_div_3_mag_0.Q0.t7 VSS 0.0329f
C2973 CLK_div_3_mag_0.Q0.t6 VSS 0.0263f
C2974 CLK_div_3_mag_0.Q0.n3 VSS 0.0764f
C2975 CLK_div_3_mag_0.Q0.n4 VSS 0.606f
C2976 CLK_div_3_mag_0.Q0.t3 VSS 0.0641f
C2977 CLK_div_3_mag_0.Q0.t8 VSS 0.0199f
C2978 CLK_div_3_mag_0.Q0.n5 VSS 0.0675f
C2979 CLK_div_3_mag_0.Q0.n6 VSS 0.447f
.ends

