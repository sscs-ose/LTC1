magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -9351 -3458 9351 3458
<< metal3 >>
rect -7351 1448 7351 1458
rect -7351 1392 -7341 1448
rect -7285 1392 -7199 1448
rect -7143 1392 -7057 1448
rect -7001 1392 -6915 1448
rect -6859 1392 -6773 1448
rect -6717 1392 -6631 1448
rect -6575 1392 -6489 1448
rect -6433 1392 -6347 1448
rect -6291 1392 -6205 1448
rect -6149 1392 -6063 1448
rect -6007 1392 -5921 1448
rect -5865 1392 -5779 1448
rect -5723 1392 -5637 1448
rect -5581 1392 -5495 1448
rect -5439 1392 -5353 1448
rect -5297 1392 -5211 1448
rect -5155 1392 -5069 1448
rect -5013 1392 -4927 1448
rect -4871 1392 -4785 1448
rect -4729 1392 -4643 1448
rect -4587 1392 -4501 1448
rect -4445 1392 -4359 1448
rect -4303 1392 -4217 1448
rect -4161 1392 -4075 1448
rect -4019 1392 -3933 1448
rect -3877 1392 -3791 1448
rect -3735 1392 -3649 1448
rect -3593 1392 -3507 1448
rect -3451 1392 -3365 1448
rect -3309 1392 -3223 1448
rect -3167 1392 -3081 1448
rect -3025 1392 -2939 1448
rect -2883 1392 -2797 1448
rect -2741 1392 -2655 1448
rect -2599 1392 -2513 1448
rect -2457 1392 -2371 1448
rect -2315 1392 -2229 1448
rect -2173 1392 -2087 1448
rect -2031 1392 -1945 1448
rect -1889 1392 -1803 1448
rect -1747 1392 -1661 1448
rect -1605 1392 -1519 1448
rect -1463 1392 -1377 1448
rect -1321 1392 -1235 1448
rect -1179 1392 -1093 1448
rect -1037 1392 -951 1448
rect -895 1392 -809 1448
rect -753 1392 -667 1448
rect -611 1392 -525 1448
rect -469 1392 -383 1448
rect -327 1392 -241 1448
rect -185 1392 -99 1448
rect -43 1392 43 1448
rect 99 1392 185 1448
rect 241 1392 327 1448
rect 383 1392 469 1448
rect 525 1392 611 1448
rect 667 1392 753 1448
rect 809 1392 895 1448
rect 951 1392 1037 1448
rect 1093 1392 1179 1448
rect 1235 1392 1321 1448
rect 1377 1392 1463 1448
rect 1519 1392 1605 1448
rect 1661 1392 1747 1448
rect 1803 1392 1889 1448
rect 1945 1392 2031 1448
rect 2087 1392 2173 1448
rect 2229 1392 2315 1448
rect 2371 1392 2457 1448
rect 2513 1392 2599 1448
rect 2655 1392 2741 1448
rect 2797 1392 2883 1448
rect 2939 1392 3025 1448
rect 3081 1392 3167 1448
rect 3223 1392 3309 1448
rect 3365 1392 3451 1448
rect 3507 1392 3593 1448
rect 3649 1392 3735 1448
rect 3791 1392 3877 1448
rect 3933 1392 4019 1448
rect 4075 1392 4161 1448
rect 4217 1392 4303 1448
rect 4359 1392 4445 1448
rect 4501 1392 4587 1448
rect 4643 1392 4729 1448
rect 4785 1392 4871 1448
rect 4927 1392 5013 1448
rect 5069 1392 5155 1448
rect 5211 1392 5297 1448
rect 5353 1392 5439 1448
rect 5495 1392 5581 1448
rect 5637 1392 5723 1448
rect 5779 1392 5865 1448
rect 5921 1392 6007 1448
rect 6063 1392 6149 1448
rect 6205 1392 6291 1448
rect 6347 1392 6433 1448
rect 6489 1392 6575 1448
rect 6631 1392 6717 1448
rect 6773 1392 6859 1448
rect 6915 1392 7001 1448
rect 7057 1392 7143 1448
rect 7199 1392 7285 1448
rect 7341 1392 7351 1448
rect -7351 1306 7351 1392
rect -7351 1250 -7341 1306
rect -7285 1250 -7199 1306
rect -7143 1250 -7057 1306
rect -7001 1250 -6915 1306
rect -6859 1250 -6773 1306
rect -6717 1250 -6631 1306
rect -6575 1250 -6489 1306
rect -6433 1250 -6347 1306
rect -6291 1250 -6205 1306
rect -6149 1250 -6063 1306
rect -6007 1250 -5921 1306
rect -5865 1250 -5779 1306
rect -5723 1250 -5637 1306
rect -5581 1250 -5495 1306
rect -5439 1250 -5353 1306
rect -5297 1250 -5211 1306
rect -5155 1250 -5069 1306
rect -5013 1250 -4927 1306
rect -4871 1250 -4785 1306
rect -4729 1250 -4643 1306
rect -4587 1250 -4501 1306
rect -4445 1250 -4359 1306
rect -4303 1250 -4217 1306
rect -4161 1250 -4075 1306
rect -4019 1250 -3933 1306
rect -3877 1250 -3791 1306
rect -3735 1250 -3649 1306
rect -3593 1250 -3507 1306
rect -3451 1250 -3365 1306
rect -3309 1250 -3223 1306
rect -3167 1250 -3081 1306
rect -3025 1250 -2939 1306
rect -2883 1250 -2797 1306
rect -2741 1250 -2655 1306
rect -2599 1250 -2513 1306
rect -2457 1250 -2371 1306
rect -2315 1250 -2229 1306
rect -2173 1250 -2087 1306
rect -2031 1250 -1945 1306
rect -1889 1250 -1803 1306
rect -1747 1250 -1661 1306
rect -1605 1250 -1519 1306
rect -1463 1250 -1377 1306
rect -1321 1250 -1235 1306
rect -1179 1250 -1093 1306
rect -1037 1250 -951 1306
rect -895 1250 -809 1306
rect -753 1250 -667 1306
rect -611 1250 -525 1306
rect -469 1250 -383 1306
rect -327 1250 -241 1306
rect -185 1250 -99 1306
rect -43 1250 43 1306
rect 99 1250 185 1306
rect 241 1250 327 1306
rect 383 1250 469 1306
rect 525 1250 611 1306
rect 667 1250 753 1306
rect 809 1250 895 1306
rect 951 1250 1037 1306
rect 1093 1250 1179 1306
rect 1235 1250 1321 1306
rect 1377 1250 1463 1306
rect 1519 1250 1605 1306
rect 1661 1250 1747 1306
rect 1803 1250 1889 1306
rect 1945 1250 2031 1306
rect 2087 1250 2173 1306
rect 2229 1250 2315 1306
rect 2371 1250 2457 1306
rect 2513 1250 2599 1306
rect 2655 1250 2741 1306
rect 2797 1250 2883 1306
rect 2939 1250 3025 1306
rect 3081 1250 3167 1306
rect 3223 1250 3309 1306
rect 3365 1250 3451 1306
rect 3507 1250 3593 1306
rect 3649 1250 3735 1306
rect 3791 1250 3877 1306
rect 3933 1250 4019 1306
rect 4075 1250 4161 1306
rect 4217 1250 4303 1306
rect 4359 1250 4445 1306
rect 4501 1250 4587 1306
rect 4643 1250 4729 1306
rect 4785 1250 4871 1306
rect 4927 1250 5013 1306
rect 5069 1250 5155 1306
rect 5211 1250 5297 1306
rect 5353 1250 5439 1306
rect 5495 1250 5581 1306
rect 5637 1250 5723 1306
rect 5779 1250 5865 1306
rect 5921 1250 6007 1306
rect 6063 1250 6149 1306
rect 6205 1250 6291 1306
rect 6347 1250 6433 1306
rect 6489 1250 6575 1306
rect 6631 1250 6717 1306
rect 6773 1250 6859 1306
rect 6915 1250 7001 1306
rect 7057 1250 7143 1306
rect 7199 1250 7285 1306
rect 7341 1250 7351 1306
rect -7351 1164 7351 1250
rect -7351 1108 -7341 1164
rect -7285 1108 -7199 1164
rect -7143 1108 -7057 1164
rect -7001 1108 -6915 1164
rect -6859 1108 -6773 1164
rect -6717 1108 -6631 1164
rect -6575 1108 -6489 1164
rect -6433 1108 -6347 1164
rect -6291 1108 -6205 1164
rect -6149 1108 -6063 1164
rect -6007 1108 -5921 1164
rect -5865 1108 -5779 1164
rect -5723 1108 -5637 1164
rect -5581 1108 -5495 1164
rect -5439 1108 -5353 1164
rect -5297 1108 -5211 1164
rect -5155 1108 -5069 1164
rect -5013 1108 -4927 1164
rect -4871 1108 -4785 1164
rect -4729 1108 -4643 1164
rect -4587 1108 -4501 1164
rect -4445 1108 -4359 1164
rect -4303 1108 -4217 1164
rect -4161 1108 -4075 1164
rect -4019 1108 -3933 1164
rect -3877 1108 -3791 1164
rect -3735 1108 -3649 1164
rect -3593 1108 -3507 1164
rect -3451 1108 -3365 1164
rect -3309 1108 -3223 1164
rect -3167 1108 -3081 1164
rect -3025 1108 -2939 1164
rect -2883 1108 -2797 1164
rect -2741 1108 -2655 1164
rect -2599 1108 -2513 1164
rect -2457 1108 -2371 1164
rect -2315 1108 -2229 1164
rect -2173 1108 -2087 1164
rect -2031 1108 -1945 1164
rect -1889 1108 -1803 1164
rect -1747 1108 -1661 1164
rect -1605 1108 -1519 1164
rect -1463 1108 -1377 1164
rect -1321 1108 -1235 1164
rect -1179 1108 -1093 1164
rect -1037 1108 -951 1164
rect -895 1108 -809 1164
rect -753 1108 -667 1164
rect -611 1108 -525 1164
rect -469 1108 -383 1164
rect -327 1108 -241 1164
rect -185 1108 -99 1164
rect -43 1108 43 1164
rect 99 1108 185 1164
rect 241 1108 327 1164
rect 383 1108 469 1164
rect 525 1108 611 1164
rect 667 1108 753 1164
rect 809 1108 895 1164
rect 951 1108 1037 1164
rect 1093 1108 1179 1164
rect 1235 1108 1321 1164
rect 1377 1108 1463 1164
rect 1519 1108 1605 1164
rect 1661 1108 1747 1164
rect 1803 1108 1889 1164
rect 1945 1108 2031 1164
rect 2087 1108 2173 1164
rect 2229 1108 2315 1164
rect 2371 1108 2457 1164
rect 2513 1108 2599 1164
rect 2655 1108 2741 1164
rect 2797 1108 2883 1164
rect 2939 1108 3025 1164
rect 3081 1108 3167 1164
rect 3223 1108 3309 1164
rect 3365 1108 3451 1164
rect 3507 1108 3593 1164
rect 3649 1108 3735 1164
rect 3791 1108 3877 1164
rect 3933 1108 4019 1164
rect 4075 1108 4161 1164
rect 4217 1108 4303 1164
rect 4359 1108 4445 1164
rect 4501 1108 4587 1164
rect 4643 1108 4729 1164
rect 4785 1108 4871 1164
rect 4927 1108 5013 1164
rect 5069 1108 5155 1164
rect 5211 1108 5297 1164
rect 5353 1108 5439 1164
rect 5495 1108 5581 1164
rect 5637 1108 5723 1164
rect 5779 1108 5865 1164
rect 5921 1108 6007 1164
rect 6063 1108 6149 1164
rect 6205 1108 6291 1164
rect 6347 1108 6433 1164
rect 6489 1108 6575 1164
rect 6631 1108 6717 1164
rect 6773 1108 6859 1164
rect 6915 1108 7001 1164
rect 7057 1108 7143 1164
rect 7199 1108 7285 1164
rect 7341 1108 7351 1164
rect -7351 1022 7351 1108
rect -7351 966 -7341 1022
rect -7285 966 -7199 1022
rect -7143 966 -7057 1022
rect -7001 966 -6915 1022
rect -6859 966 -6773 1022
rect -6717 966 -6631 1022
rect -6575 966 -6489 1022
rect -6433 966 -6347 1022
rect -6291 966 -6205 1022
rect -6149 966 -6063 1022
rect -6007 966 -5921 1022
rect -5865 966 -5779 1022
rect -5723 966 -5637 1022
rect -5581 966 -5495 1022
rect -5439 966 -5353 1022
rect -5297 966 -5211 1022
rect -5155 966 -5069 1022
rect -5013 966 -4927 1022
rect -4871 966 -4785 1022
rect -4729 966 -4643 1022
rect -4587 966 -4501 1022
rect -4445 966 -4359 1022
rect -4303 966 -4217 1022
rect -4161 966 -4075 1022
rect -4019 966 -3933 1022
rect -3877 966 -3791 1022
rect -3735 966 -3649 1022
rect -3593 966 -3507 1022
rect -3451 966 -3365 1022
rect -3309 966 -3223 1022
rect -3167 966 -3081 1022
rect -3025 966 -2939 1022
rect -2883 966 -2797 1022
rect -2741 966 -2655 1022
rect -2599 966 -2513 1022
rect -2457 966 -2371 1022
rect -2315 966 -2229 1022
rect -2173 966 -2087 1022
rect -2031 966 -1945 1022
rect -1889 966 -1803 1022
rect -1747 966 -1661 1022
rect -1605 966 -1519 1022
rect -1463 966 -1377 1022
rect -1321 966 -1235 1022
rect -1179 966 -1093 1022
rect -1037 966 -951 1022
rect -895 966 -809 1022
rect -753 966 -667 1022
rect -611 966 -525 1022
rect -469 966 -383 1022
rect -327 966 -241 1022
rect -185 966 -99 1022
rect -43 966 43 1022
rect 99 966 185 1022
rect 241 966 327 1022
rect 383 966 469 1022
rect 525 966 611 1022
rect 667 966 753 1022
rect 809 966 895 1022
rect 951 966 1037 1022
rect 1093 966 1179 1022
rect 1235 966 1321 1022
rect 1377 966 1463 1022
rect 1519 966 1605 1022
rect 1661 966 1747 1022
rect 1803 966 1889 1022
rect 1945 966 2031 1022
rect 2087 966 2173 1022
rect 2229 966 2315 1022
rect 2371 966 2457 1022
rect 2513 966 2599 1022
rect 2655 966 2741 1022
rect 2797 966 2883 1022
rect 2939 966 3025 1022
rect 3081 966 3167 1022
rect 3223 966 3309 1022
rect 3365 966 3451 1022
rect 3507 966 3593 1022
rect 3649 966 3735 1022
rect 3791 966 3877 1022
rect 3933 966 4019 1022
rect 4075 966 4161 1022
rect 4217 966 4303 1022
rect 4359 966 4445 1022
rect 4501 966 4587 1022
rect 4643 966 4729 1022
rect 4785 966 4871 1022
rect 4927 966 5013 1022
rect 5069 966 5155 1022
rect 5211 966 5297 1022
rect 5353 966 5439 1022
rect 5495 966 5581 1022
rect 5637 966 5723 1022
rect 5779 966 5865 1022
rect 5921 966 6007 1022
rect 6063 966 6149 1022
rect 6205 966 6291 1022
rect 6347 966 6433 1022
rect 6489 966 6575 1022
rect 6631 966 6717 1022
rect 6773 966 6859 1022
rect 6915 966 7001 1022
rect 7057 966 7143 1022
rect 7199 966 7285 1022
rect 7341 966 7351 1022
rect -7351 880 7351 966
rect -7351 824 -7341 880
rect -7285 824 -7199 880
rect -7143 824 -7057 880
rect -7001 824 -6915 880
rect -6859 824 -6773 880
rect -6717 824 -6631 880
rect -6575 824 -6489 880
rect -6433 824 -6347 880
rect -6291 824 -6205 880
rect -6149 824 -6063 880
rect -6007 824 -5921 880
rect -5865 824 -5779 880
rect -5723 824 -5637 880
rect -5581 824 -5495 880
rect -5439 824 -5353 880
rect -5297 824 -5211 880
rect -5155 824 -5069 880
rect -5013 824 -4927 880
rect -4871 824 -4785 880
rect -4729 824 -4643 880
rect -4587 824 -4501 880
rect -4445 824 -4359 880
rect -4303 824 -4217 880
rect -4161 824 -4075 880
rect -4019 824 -3933 880
rect -3877 824 -3791 880
rect -3735 824 -3649 880
rect -3593 824 -3507 880
rect -3451 824 -3365 880
rect -3309 824 -3223 880
rect -3167 824 -3081 880
rect -3025 824 -2939 880
rect -2883 824 -2797 880
rect -2741 824 -2655 880
rect -2599 824 -2513 880
rect -2457 824 -2371 880
rect -2315 824 -2229 880
rect -2173 824 -2087 880
rect -2031 824 -1945 880
rect -1889 824 -1803 880
rect -1747 824 -1661 880
rect -1605 824 -1519 880
rect -1463 824 -1377 880
rect -1321 824 -1235 880
rect -1179 824 -1093 880
rect -1037 824 -951 880
rect -895 824 -809 880
rect -753 824 -667 880
rect -611 824 -525 880
rect -469 824 -383 880
rect -327 824 -241 880
rect -185 824 -99 880
rect -43 824 43 880
rect 99 824 185 880
rect 241 824 327 880
rect 383 824 469 880
rect 525 824 611 880
rect 667 824 753 880
rect 809 824 895 880
rect 951 824 1037 880
rect 1093 824 1179 880
rect 1235 824 1321 880
rect 1377 824 1463 880
rect 1519 824 1605 880
rect 1661 824 1747 880
rect 1803 824 1889 880
rect 1945 824 2031 880
rect 2087 824 2173 880
rect 2229 824 2315 880
rect 2371 824 2457 880
rect 2513 824 2599 880
rect 2655 824 2741 880
rect 2797 824 2883 880
rect 2939 824 3025 880
rect 3081 824 3167 880
rect 3223 824 3309 880
rect 3365 824 3451 880
rect 3507 824 3593 880
rect 3649 824 3735 880
rect 3791 824 3877 880
rect 3933 824 4019 880
rect 4075 824 4161 880
rect 4217 824 4303 880
rect 4359 824 4445 880
rect 4501 824 4587 880
rect 4643 824 4729 880
rect 4785 824 4871 880
rect 4927 824 5013 880
rect 5069 824 5155 880
rect 5211 824 5297 880
rect 5353 824 5439 880
rect 5495 824 5581 880
rect 5637 824 5723 880
rect 5779 824 5865 880
rect 5921 824 6007 880
rect 6063 824 6149 880
rect 6205 824 6291 880
rect 6347 824 6433 880
rect 6489 824 6575 880
rect 6631 824 6717 880
rect 6773 824 6859 880
rect 6915 824 7001 880
rect 7057 824 7143 880
rect 7199 824 7285 880
rect 7341 824 7351 880
rect -7351 738 7351 824
rect -7351 682 -7341 738
rect -7285 682 -7199 738
rect -7143 682 -7057 738
rect -7001 682 -6915 738
rect -6859 682 -6773 738
rect -6717 682 -6631 738
rect -6575 682 -6489 738
rect -6433 682 -6347 738
rect -6291 682 -6205 738
rect -6149 682 -6063 738
rect -6007 682 -5921 738
rect -5865 682 -5779 738
rect -5723 682 -5637 738
rect -5581 682 -5495 738
rect -5439 682 -5353 738
rect -5297 682 -5211 738
rect -5155 682 -5069 738
rect -5013 682 -4927 738
rect -4871 682 -4785 738
rect -4729 682 -4643 738
rect -4587 682 -4501 738
rect -4445 682 -4359 738
rect -4303 682 -4217 738
rect -4161 682 -4075 738
rect -4019 682 -3933 738
rect -3877 682 -3791 738
rect -3735 682 -3649 738
rect -3593 682 -3507 738
rect -3451 682 -3365 738
rect -3309 682 -3223 738
rect -3167 682 -3081 738
rect -3025 682 -2939 738
rect -2883 682 -2797 738
rect -2741 682 -2655 738
rect -2599 682 -2513 738
rect -2457 682 -2371 738
rect -2315 682 -2229 738
rect -2173 682 -2087 738
rect -2031 682 -1945 738
rect -1889 682 -1803 738
rect -1747 682 -1661 738
rect -1605 682 -1519 738
rect -1463 682 -1377 738
rect -1321 682 -1235 738
rect -1179 682 -1093 738
rect -1037 682 -951 738
rect -895 682 -809 738
rect -753 682 -667 738
rect -611 682 -525 738
rect -469 682 -383 738
rect -327 682 -241 738
rect -185 682 -99 738
rect -43 682 43 738
rect 99 682 185 738
rect 241 682 327 738
rect 383 682 469 738
rect 525 682 611 738
rect 667 682 753 738
rect 809 682 895 738
rect 951 682 1037 738
rect 1093 682 1179 738
rect 1235 682 1321 738
rect 1377 682 1463 738
rect 1519 682 1605 738
rect 1661 682 1747 738
rect 1803 682 1889 738
rect 1945 682 2031 738
rect 2087 682 2173 738
rect 2229 682 2315 738
rect 2371 682 2457 738
rect 2513 682 2599 738
rect 2655 682 2741 738
rect 2797 682 2883 738
rect 2939 682 3025 738
rect 3081 682 3167 738
rect 3223 682 3309 738
rect 3365 682 3451 738
rect 3507 682 3593 738
rect 3649 682 3735 738
rect 3791 682 3877 738
rect 3933 682 4019 738
rect 4075 682 4161 738
rect 4217 682 4303 738
rect 4359 682 4445 738
rect 4501 682 4587 738
rect 4643 682 4729 738
rect 4785 682 4871 738
rect 4927 682 5013 738
rect 5069 682 5155 738
rect 5211 682 5297 738
rect 5353 682 5439 738
rect 5495 682 5581 738
rect 5637 682 5723 738
rect 5779 682 5865 738
rect 5921 682 6007 738
rect 6063 682 6149 738
rect 6205 682 6291 738
rect 6347 682 6433 738
rect 6489 682 6575 738
rect 6631 682 6717 738
rect 6773 682 6859 738
rect 6915 682 7001 738
rect 7057 682 7143 738
rect 7199 682 7285 738
rect 7341 682 7351 738
rect -7351 596 7351 682
rect -7351 540 -7341 596
rect -7285 540 -7199 596
rect -7143 540 -7057 596
rect -7001 540 -6915 596
rect -6859 540 -6773 596
rect -6717 540 -6631 596
rect -6575 540 -6489 596
rect -6433 540 -6347 596
rect -6291 540 -6205 596
rect -6149 540 -6063 596
rect -6007 540 -5921 596
rect -5865 540 -5779 596
rect -5723 540 -5637 596
rect -5581 540 -5495 596
rect -5439 540 -5353 596
rect -5297 540 -5211 596
rect -5155 540 -5069 596
rect -5013 540 -4927 596
rect -4871 540 -4785 596
rect -4729 540 -4643 596
rect -4587 540 -4501 596
rect -4445 540 -4359 596
rect -4303 540 -4217 596
rect -4161 540 -4075 596
rect -4019 540 -3933 596
rect -3877 540 -3791 596
rect -3735 540 -3649 596
rect -3593 540 -3507 596
rect -3451 540 -3365 596
rect -3309 540 -3223 596
rect -3167 540 -3081 596
rect -3025 540 -2939 596
rect -2883 540 -2797 596
rect -2741 540 -2655 596
rect -2599 540 -2513 596
rect -2457 540 -2371 596
rect -2315 540 -2229 596
rect -2173 540 -2087 596
rect -2031 540 -1945 596
rect -1889 540 -1803 596
rect -1747 540 -1661 596
rect -1605 540 -1519 596
rect -1463 540 -1377 596
rect -1321 540 -1235 596
rect -1179 540 -1093 596
rect -1037 540 -951 596
rect -895 540 -809 596
rect -753 540 -667 596
rect -611 540 -525 596
rect -469 540 -383 596
rect -327 540 -241 596
rect -185 540 -99 596
rect -43 540 43 596
rect 99 540 185 596
rect 241 540 327 596
rect 383 540 469 596
rect 525 540 611 596
rect 667 540 753 596
rect 809 540 895 596
rect 951 540 1037 596
rect 1093 540 1179 596
rect 1235 540 1321 596
rect 1377 540 1463 596
rect 1519 540 1605 596
rect 1661 540 1747 596
rect 1803 540 1889 596
rect 1945 540 2031 596
rect 2087 540 2173 596
rect 2229 540 2315 596
rect 2371 540 2457 596
rect 2513 540 2599 596
rect 2655 540 2741 596
rect 2797 540 2883 596
rect 2939 540 3025 596
rect 3081 540 3167 596
rect 3223 540 3309 596
rect 3365 540 3451 596
rect 3507 540 3593 596
rect 3649 540 3735 596
rect 3791 540 3877 596
rect 3933 540 4019 596
rect 4075 540 4161 596
rect 4217 540 4303 596
rect 4359 540 4445 596
rect 4501 540 4587 596
rect 4643 540 4729 596
rect 4785 540 4871 596
rect 4927 540 5013 596
rect 5069 540 5155 596
rect 5211 540 5297 596
rect 5353 540 5439 596
rect 5495 540 5581 596
rect 5637 540 5723 596
rect 5779 540 5865 596
rect 5921 540 6007 596
rect 6063 540 6149 596
rect 6205 540 6291 596
rect 6347 540 6433 596
rect 6489 540 6575 596
rect 6631 540 6717 596
rect 6773 540 6859 596
rect 6915 540 7001 596
rect 7057 540 7143 596
rect 7199 540 7285 596
rect 7341 540 7351 596
rect -7351 454 7351 540
rect -7351 398 -7341 454
rect -7285 398 -7199 454
rect -7143 398 -7057 454
rect -7001 398 -6915 454
rect -6859 398 -6773 454
rect -6717 398 -6631 454
rect -6575 398 -6489 454
rect -6433 398 -6347 454
rect -6291 398 -6205 454
rect -6149 398 -6063 454
rect -6007 398 -5921 454
rect -5865 398 -5779 454
rect -5723 398 -5637 454
rect -5581 398 -5495 454
rect -5439 398 -5353 454
rect -5297 398 -5211 454
rect -5155 398 -5069 454
rect -5013 398 -4927 454
rect -4871 398 -4785 454
rect -4729 398 -4643 454
rect -4587 398 -4501 454
rect -4445 398 -4359 454
rect -4303 398 -4217 454
rect -4161 398 -4075 454
rect -4019 398 -3933 454
rect -3877 398 -3791 454
rect -3735 398 -3649 454
rect -3593 398 -3507 454
rect -3451 398 -3365 454
rect -3309 398 -3223 454
rect -3167 398 -3081 454
rect -3025 398 -2939 454
rect -2883 398 -2797 454
rect -2741 398 -2655 454
rect -2599 398 -2513 454
rect -2457 398 -2371 454
rect -2315 398 -2229 454
rect -2173 398 -2087 454
rect -2031 398 -1945 454
rect -1889 398 -1803 454
rect -1747 398 -1661 454
rect -1605 398 -1519 454
rect -1463 398 -1377 454
rect -1321 398 -1235 454
rect -1179 398 -1093 454
rect -1037 398 -951 454
rect -895 398 -809 454
rect -753 398 -667 454
rect -611 398 -525 454
rect -469 398 -383 454
rect -327 398 -241 454
rect -185 398 -99 454
rect -43 398 43 454
rect 99 398 185 454
rect 241 398 327 454
rect 383 398 469 454
rect 525 398 611 454
rect 667 398 753 454
rect 809 398 895 454
rect 951 398 1037 454
rect 1093 398 1179 454
rect 1235 398 1321 454
rect 1377 398 1463 454
rect 1519 398 1605 454
rect 1661 398 1747 454
rect 1803 398 1889 454
rect 1945 398 2031 454
rect 2087 398 2173 454
rect 2229 398 2315 454
rect 2371 398 2457 454
rect 2513 398 2599 454
rect 2655 398 2741 454
rect 2797 398 2883 454
rect 2939 398 3025 454
rect 3081 398 3167 454
rect 3223 398 3309 454
rect 3365 398 3451 454
rect 3507 398 3593 454
rect 3649 398 3735 454
rect 3791 398 3877 454
rect 3933 398 4019 454
rect 4075 398 4161 454
rect 4217 398 4303 454
rect 4359 398 4445 454
rect 4501 398 4587 454
rect 4643 398 4729 454
rect 4785 398 4871 454
rect 4927 398 5013 454
rect 5069 398 5155 454
rect 5211 398 5297 454
rect 5353 398 5439 454
rect 5495 398 5581 454
rect 5637 398 5723 454
rect 5779 398 5865 454
rect 5921 398 6007 454
rect 6063 398 6149 454
rect 6205 398 6291 454
rect 6347 398 6433 454
rect 6489 398 6575 454
rect 6631 398 6717 454
rect 6773 398 6859 454
rect 6915 398 7001 454
rect 7057 398 7143 454
rect 7199 398 7285 454
rect 7341 398 7351 454
rect -7351 312 7351 398
rect -7351 256 -7341 312
rect -7285 256 -7199 312
rect -7143 256 -7057 312
rect -7001 256 -6915 312
rect -6859 256 -6773 312
rect -6717 256 -6631 312
rect -6575 256 -6489 312
rect -6433 256 -6347 312
rect -6291 256 -6205 312
rect -6149 256 -6063 312
rect -6007 256 -5921 312
rect -5865 256 -5779 312
rect -5723 256 -5637 312
rect -5581 256 -5495 312
rect -5439 256 -5353 312
rect -5297 256 -5211 312
rect -5155 256 -5069 312
rect -5013 256 -4927 312
rect -4871 256 -4785 312
rect -4729 256 -4643 312
rect -4587 256 -4501 312
rect -4445 256 -4359 312
rect -4303 256 -4217 312
rect -4161 256 -4075 312
rect -4019 256 -3933 312
rect -3877 256 -3791 312
rect -3735 256 -3649 312
rect -3593 256 -3507 312
rect -3451 256 -3365 312
rect -3309 256 -3223 312
rect -3167 256 -3081 312
rect -3025 256 -2939 312
rect -2883 256 -2797 312
rect -2741 256 -2655 312
rect -2599 256 -2513 312
rect -2457 256 -2371 312
rect -2315 256 -2229 312
rect -2173 256 -2087 312
rect -2031 256 -1945 312
rect -1889 256 -1803 312
rect -1747 256 -1661 312
rect -1605 256 -1519 312
rect -1463 256 -1377 312
rect -1321 256 -1235 312
rect -1179 256 -1093 312
rect -1037 256 -951 312
rect -895 256 -809 312
rect -753 256 -667 312
rect -611 256 -525 312
rect -469 256 -383 312
rect -327 256 -241 312
rect -185 256 -99 312
rect -43 256 43 312
rect 99 256 185 312
rect 241 256 327 312
rect 383 256 469 312
rect 525 256 611 312
rect 667 256 753 312
rect 809 256 895 312
rect 951 256 1037 312
rect 1093 256 1179 312
rect 1235 256 1321 312
rect 1377 256 1463 312
rect 1519 256 1605 312
rect 1661 256 1747 312
rect 1803 256 1889 312
rect 1945 256 2031 312
rect 2087 256 2173 312
rect 2229 256 2315 312
rect 2371 256 2457 312
rect 2513 256 2599 312
rect 2655 256 2741 312
rect 2797 256 2883 312
rect 2939 256 3025 312
rect 3081 256 3167 312
rect 3223 256 3309 312
rect 3365 256 3451 312
rect 3507 256 3593 312
rect 3649 256 3735 312
rect 3791 256 3877 312
rect 3933 256 4019 312
rect 4075 256 4161 312
rect 4217 256 4303 312
rect 4359 256 4445 312
rect 4501 256 4587 312
rect 4643 256 4729 312
rect 4785 256 4871 312
rect 4927 256 5013 312
rect 5069 256 5155 312
rect 5211 256 5297 312
rect 5353 256 5439 312
rect 5495 256 5581 312
rect 5637 256 5723 312
rect 5779 256 5865 312
rect 5921 256 6007 312
rect 6063 256 6149 312
rect 6205 256 6291 312
rect 6347 256 6433 312
rect 6489 256 6575 312
rect 6631 256 6717 312
rect 6773 256 6859 312
rect 6915 256 7001 312
rect 7057 256 7143 312
rect 7199 256 7285 312
rect 7341 256 7351 312
rect -7351 170 7351 256
rect -7351 114 -7341 170
rect -7285 114 -7199 170
rect -7143 114 -7057 170
rect -7001 114 -6915 170
rect -6859 114 -6773 170
rect -6717 114 -6631 170
rect -6575 114 -6489 170
rect -6433 114 -6347 170
rect -6291 114 -6205 170
rect -6149 114 -6063 170
rect -6007 114 -5921 170
rect -5865 114 -5779 170
rect -5723 114 -5637 170
rect -5581 114 -5495 170
rect -5439 114 -5353 170
rect -5297 114 -5211 170
rect -5155 114 -5069 170
rect -5013 114 -4927 170
rect -4871 114 -4785 170
rect -4729 114 -4643 170
rect -4587 114 -4501 170
rect -4445 114 -4359 170
rect -4303 114 -4217 170
rect -4161 114 -4075 170
rect -4019 114 -3933 170
rect -3877 114 -3791 170
rect -3735 114 -3649 170
rect -3593 114 -3507 170
rect -3451 114 -3365 170
rect -3309 114 -3223 170
rect -3167 114 -3081 170
rect -3025 114 -2939 170
rect -2883 114 -2797 170
rect -2741 114 -2655 170
rect -2599 114 -2513 170
rect -2457 114 -2371 170
rect -2315 114 -2229 170
rect -2173 114 -2087 170
rect -2031 114 -1945 170
rect -1889 114 -1803 170
rect -1747 114 -1661 170
rect -1605 114 -1519 170
rect -1463 114 -1377 170
rect -1321 114 -1235 170
rect -1179 114 -1093 170
rect -1037 114 -951 170
rect -895 114 -809 170
rect -753 114 -667 170
rect -611 114 -525 170
rect -469 114 -383 170
rect -327 114 -241 170
rect -185 114 -99 170
rect -43 114 43 170
rect 99 114 185 170
rect 241 114 327 170
rect 383 114 469 170
rect 525 114 611 170
rect 667 114 753 170
rect 809 114 895 170
rect 951 114 1037 170
rect 1093 114 1179 170
rect 1235 114 1321 170
rect 1377 114 1463 170
rect 1519 114 1605 170
rect 1661 114 1747 170
rect 1803 114 1889 170
rect 1945 114 2031 170
rect 2087 114 2173 170
rect 2229 114 2315 170
rect 2371 114 2457 170
rect 2513 114 2599 170
rect 2655 114 2741 170
rect 2797 114 2883 170
rect 2939 114 3025 170
rect 3081 114 3167 170
rect 3223 114 3309 170
rect 3365 114 3451 170
rect 3507 114 3593 170
rect 3649 114 3735 170
rect 3791 114 3877 170
rect 3933 114 4019 170
rect 4075 114 4161 170
rect 4217 114 4303 170
rect 4359 114 4445 170
rect 4501 114 4587 170
rect 4643 114 4729 170
rect 4785 114 4871 170
rect 4927 114 5013 170
rect 5069 114 5155 170
rect 5211 114 5297 170
rect 5353 114 5439 170
rect 5495 114 5581 170
rect 5637 114 5723 170
rect 5779 114 5865 170
rect 5921 114 6007 170
rect 6063 114 6149 170
rect 6205 114 6291 170
rect 6347 114 6433 170
rect 6489 114 6575 170
rect 6631 114 6717 170
rect 6773 114 6859 170
rect 6915 114 7001 170
rect 7057 114 7143 170
rect 7199 114 7285 170
rect 7341 114 7351 170
rect -7351 28 7351 114
rect -7351 -28 -7341 28
rect -7285 -28 -7199 28
rect -7143 -28 -7057 28
rect -7001 -28 -6915 28
rect -6859 -28 -6773 28
rect -6717 -28 -6631 28
rect -6575 -28 -6489 28
rect -6433 -28 -6347 28
rect -6291 -28 -6205 28
rect -6149 -28 -6063 28
rect -6007 -28 -5921 28
rect -5865 -28 -5779 28
rect -5723 -28 -5637 28
rect -5581 -28 -5495 28
rect -5439 -28 -5353 28
rect -5297 -28 -5211 28
rect -5155 -28 -5069 28
rect -5013 -28 -4927 28
rect -4871 -28 -4785 28
rect -4729 -28 -4643 28
rect -4587 -28 -4501 28
rect -4445 -28 -4359 28
rect -4303 -28 -4217 28
rect -4161 -28 -4075 28
rect -4019 -28 -3933 28
rect -3877 -28 -3791 28
rect -3735 -28 -3649 28
rect -3593 -28 -3507 28
rect -3451 -28 -3365 28
rect -3309 -28 -3223 28
rect -3167 -28 -3081 28
rect -3025 -28 -2939 28
rect -2883 -28 -2797 28
rect -2741 -28 -2655 28
rect -2599 -28 -2513 28
rect -2457 -28 -2371 28
rect -2315 -28 -2229 28
rect -2173 -28 -2087 28
rect -2031 -28 -1945 28
rect -1889 -28 -1803 28
rect -1747 -28 -1661 28
rect -1605 -28 -1519 28
rect -1463 -28 -1377 28
rect -1321 -28 -1235 28
rect -1179 -28 -1093 28
rect -1037 -28 -951 28
rect -895 -28 -809 28
rect -753 -28 -667 28
rect -611 -28 -525 28
rect -469 -28 -383 28
rect -327 -28 -241 28
rect -185 -28 -99 28
rect -43 -28 43 28
rect 99 -28 185 28
rect 241 -28 327 28
rect 383 -28 469 28
rect 525 -28 611 28
rect 667 -28 753 28
rect 809 -28 895 28
rect 951 -28 1037 28
rect 1093 -28 1179 28
rect 1235 -28 1321 28
rect 1377 -28 1463 28
rect 1519 -28 1605 28
rect 1661 -28 1747 28
rect 1803 -28 1889 28
rect 1945 -28 2031 28
rect 2087 -28 2173 28
rect 2229 -28 2315 28
rect 2371 -28 2457 28
rect 2513 -28 2599 28
rect 2655 -28 2741 28
rect 2797 -28 2883 28
rect 2939 -28 3025 28
rect 3081 -28 3167 28
rect 3223 -28 3309 28
rect 3365 -28 3451 28
rect 3507 -28 3593 28
rect 3649 -28 3735 28
rect 3791 -28 3877 28
rect 3933 -28 4019 28
rect 4075 -28 4161 28
rect 4217 -28 4303 28
rect 4359 -28 4445 28
rect 4501 -28 4587 28
rect 4643 -28 4729 28
rect 4785 -28 4871 28
rect 4927 -28 5013 28
rect 5069 -28 5155 28
rect 5211 -28 5297 28
rect 5353 -28 5439 28
rect 5495 -28 5581 28
rect 5637 -28 5723 28
rect 5779 -28 5865 28
rect 5921 -28 6007 28
rect 6063 -28 6149 28
rect 6205 -28 6291 28
rect 6347 -28 6433 28
rect 6489 -28 6575 28
rect 6631 -28 6717 28
rect 6773 -28 6859 28
rect 6915 -28 7001 28
rect 7057 -28 7143 28
rect 7199 -28 7285 28
rect 7341 -28 7351 28
rect -7351 -114 7351 -28
rect -7351 -170 -7341 -114
rect -7285 -170 -7199 -114
rect -7143 -170 -7057 -114
rect -7001 -170 -6915 -114
rect -6859 -170 -6773 -114
rect -6717 -170 -6631 -114
rect -6575 -170 -6489 -114
rect -6433 -170 -6347 -114
rect -6291 -170 -6205 -114
rect -6149 -170 -6063 -114
rect -6007 -170 -5921 -114
rect -5865 -170 -5779 -114
rect -5723 -170 -5637 -114
rect -5581 -170 -5495 -114
rect -5439 -170 -5353 -114
rect -5297 -170 -5211 -114
rect -5155 -170 -5069 -114
rect -5013 -170 -4927 -114
rect -4871 -170 -4785 -114
rect -4729 -170 -4643 -114
rect -4587 -170 -4501 -114
rect -4445 -170 -4359 -114
rect -4303 -170 -4217 -114
rect -4161 -170 -4075 -114
rect -4019 -170 -3933 -114
rect -3877 -170 -3791 -114
rect -3735 -170 -3649 -114
rect -3593 -170 -3507 -114
rect -3451 -170 -3365 -114
rect -3309 -170 -3223 -114
rect -3167 -170 -3081 -114
rect -3025 -170 -2939 -114
rect -2883 -170 -2797 -114
rect -2741 -170 -2655 -114
rect -2599 -170 -2513 -114
rect -2457 -170 -2371 -114
rect -2315 -170 -2229 -114
rect -2173 -170 -2087 -114
rect -2031 -170 -1945 -114
rect -1889 -170 -1803 -114
rect -1747 -170 -1661 -114
rect -1605 -170 -1519 -114
rect -1463 -170 -1377 -114
rect -1321 -170 -1235 -114
rect -1179 -170 -1093 -114
rect -1037 -170 -951 -114
rect -895 -170 -809 -114
rect -753 -170 -667 -114
rect -611 -170 -525 -114
rect -469 -170 -383 -114
rect -327 -170 -241 -114
rect -185 -170 -99 -114
rect -43 -170 43 -114
rect 99 -170 185 -114
rect 241 -170 327 -114
rect 383 -170 469 -114
rect 525 -170 611 -114
rect 667 -170 753 -114
rect 809 -170 895 -114
rect 951 -170 1037 -114
rect 1093 -170 1179 -114
rect 1235 -170 1321 -114
rect 1377 -170 1463 -114
rect 1519 -170 1605 -114
rect 1661 -170 1747 -114
rect 1803 -170 1889 -114
rect 1945 -170 2031 -114
rect 2087 -170 2173 -114
rect 2229 -170 2315 -114
rect 2371 -170 2457 -114
rect 2513 -170 2599 -114
rect 2655 -170 2741 -114
rect 2797 -170 2883 -114
rect 2939 -170 3025 -114
rect 3081 -170 3167 -114
rect 3223 -170 3309 -114
rect 3365 -170 3451 -114
rect 3507 -170 3593 -114
rect 3649 -170 3735 -114
rect 3791 -170 3877 -114
rect 3933 -170 4019 -114
rect 4075 -170 4161 -114
rect 4217 -170 4303 -114
rect 4359 -170 4445 -114
rect 4501 -170 4587 -114
rect 4643 -170 4729 -114
rect 4785 -170 4871 -114
rect 4927 -170 5013 -114
rect 5069 -170 5155 -114
rect 5211 -170 5297 -114
rect 5353 -170 5439 -114
rect 5495 -170 5581 -114
rect 5637 -170 5723 -114
rect 5779 -170 5865 -114
rect 5921 -170 6007 -114
rect 6063 -170 6149 -114
rect 6205 -170 6291 -114
rect 6347 -170 6433 -114
rect 6489 -170 6575 -114
rect 6631 -170 6717 -114
rect 6773 -170 6859 -114
rect 6915 -170 7001 -114
rect 7057 -170 7143 -114
rect 7199 -170 7285 -114
rect 7341 -170 7351 -114
rect -7351 -256 7351 -170
rect -7351 -312 -7341 -256
rect -7285 -312 -7199 -256
rect -7143 -312 -7057 -256
rect -7001 -312 -6915 -256
rect -6859 -312 -6773 -256
rect -6717 -312 -6631 -256
rect -6575 -312 -6489 -256
rect -6433 -312 -6347 -256
rect -6291 -312 -6205 -256
rect -6149 -312 -6063 -256
rect -6007 -312 -5921 -256
rect -5865 -312 -5779 -256
rect -5723 -312 -5637 -256
rect -5581 -312 -5495 -256
rect -5439 -312 -5353 -256
rect -5297 -312 -5211 -256
rect -5155 -312 -5069 -256
rect -5013 -312 -4927 -256
rect -4871 -312 -4785 -256
rect -4729 -312 -4643 -256
rect -4587 -312 -4501 -256
rect -4445 -312 -4359 -256
rect -4303 -312 -4217 -256
rect -4161 -312 -4075 -256
rect -4019 -312 -3933 -256
rect -3877 -312 -3791 -256
rect -3735 -312 -3649 -256
rect -3593 -312 -3507 -256
rect -3451 -312 -3365 -256
rect -3309 -312 -3223 -256
rect -3167 -312 -3081 -256
rect -3025 -312 -2939 -256
rect -2883 -312 -2797 -256
rect -2741 -312 -2655 -256
rect -2599 -312 -2513 -256
rect -2457 -312 -2371 -256
rect -2315 -312 -2229 -256
rect -2173 -312 -2087 -256
rect -2031 -312 -1945 -256
rect -1889 -312 -1803 -256
rect -1747 -312 -1661 -256
rect -1605 -312 -1519 -256
rect -1463 -312 -1377 -256
rect -1321 -312 -1235 -256
rect -1179 -312 -1093 -256
rect -1037 -312 -951 -256
rect -895 -312 -809 -256
rect -753 -312 -667 -256
rect -611 -312 -525 -256
rect -469 -312 -383 -256
rect -327 -312 -241 -256
rect -185 -312 -99 -256
rect -43 -312 43 -256
rect 99 -312 185 -256
rect 241 -312 327 -256
rect 383 -312 469 -256
rect 525 -312 611 -256
rect 667 -312 753 -256
rect 809 -312 895 -256
rect 951 -312 1037 -256
rect 1093 -312 1179 -256
rect 1235 -312 1321 -256
rect 1377 -312 1463 -256
rect 1519 -312 1605 -256
rect 1661 -312 1747 -256
rect 1803 -312 1889 -256
rect 1945 -312 2031 -256
rect 2087 -312 2173 -256
rect 2229 -312 2315 -256
rect 2371 -312 2457 -256
rect 2513 -312 2599 -256
rect 2655 -312 2741 -256
rect 2797 -312 2883 -256
rect 2939 -312 3025 -256
rect 3081 -312 3167 -256
rect 3223 -312 3309 -256
rect 3365 -312 3451 -256
rect 3507 -312 3593 -256
rect 3649 -312 3735 -256
rect 3791 -312 3877 -256
rect 3933 -312 4019 -256
rect 4075 -312 4161 -256
rect 4217 -312 4303 -256
rect 4359 -312 4445 -256
rect 4501 -312 4587 -256
rect 4643 -312 4729 -256
rect 4785 -312 4871 -256
rect 4927 -312 5013 -256
rect 5069 -312 5155 -256
rect 5211 -312 5297 -256
rect 5353 -312 5439 -256
rect 5495 -312 5581 -256
rect 5637 -312 5723 -256
rect 5779 -312 5865 -256
rect 5921 -312 6007 -256
rect 6063 -312 6149 -256
rect 6205 -312 6291 -256
rect 6347 -312 6433 -256
rect 6489 -312 6575 -256
rect 6631 -312 6717 -256
rect 6773 -312 6859 -256
rect 6915 -312 7001 -256
rect 7057 -312 7143 -256
rect 7199 -312 7285 -256
rect 7341 -312 7351 -256
rect -7351 -398 7351 -312
rect -7351 -454 -7341 -398
rect -7285 -454 -7199 -398
rect -7143 -454 -7057 -398
rect -7001 -454 -6915 -398
rect -6859 -454 -6773 -398
rect -6717 -454 -6631 -398
rect -6575 -454 -6489 -398
rect -6433 -454 -6347 -398
rect -6291 -454 -6205 -398
rect -6149 -454 -6063 -398
rect -6007 -454 -5921 -398
rect -5865 -454 -5779 -398
rect -5723 -454 -5637 -398
rect -5581 -454 -5495 -398
rect -5439 -454 -5353 -398
rect -5297 -454 -5211 -398
rect -5155 -454 -5069 -398
rect -5013 -454 -4927 -398
rect -4871 -454 -4785 -398
rect -4729 -454 -4643 -398
rect -4587 -454 -4501 -398
rect -4445 -454 -4359 -398
rect -4303 -454 -4217 -398
rect -4161 -454 -4075 -398
rect -4019 -454 -3933 -398
rect -3877 -454 -3791 -398
rect -3735 -454 -3649 -398
rect -3593 -454 -3507 -398
rect -3451 -454 -3365 -398
rect -3309 -454 -3223 -398
rect -3167 -454 -3081 -398
rect -3025 -454 -2939 -398
rect -2883 -454 -2797 -398
rect -2741 -454 -2655 -398
rect -2599 -454 -2513 -398
rect -2457 -454 -2371 -398
rect -2315 -454 -2229 -398
rect -2173 -454 -2087 -398
rect -2031 -454 -1945 -398
rect -1889 -454 -1803 -398
rect -1747 -454 -1661 -398
rect -1605 -454 -1519 -398
rect -1463 -454 -1377 -398
rect -1321 -454 -1235 -398
rect -1179 -454 -1093 -398
rect -1037 -454 -951 -398
rect -895 -454 -809 -398
rect -753 -454 -667 -398
rect -611 -454 -525 -398
rect -469 -454 -383 -398
rect -327 -454 -241 -398
rect -185 -454 -99 -398
rect -43 -454 43 -398
rect 99 -454 185 -398
rect 241 -454 327 -398
rect 383 -454 469 -398
rect 525 -454 611 -398
rect 667 -454 753 -398
rect 809 -454 895 -398
rect 951 -454 1037 -398
rect 1093 -454 1179 -398
rect 1235 -454 1321 -398
rect 1377 -454 1463 -398
rect 1519 -454 1605 -398
rect 1661 -454 1747 -398
rect 1803 -454 1889 -398
rect 1945 -454 2031 -398
rect 2087 -454 2173 -398
rect 2229 -454 2315 -398
rect 2371 -454 2457 -398
rect 2513 -454 2599 -398
rect 2655 -454 2741 -398
rect 2797 -454 2883 -398
rect 2939 -454 3025 -398
rect 3081 -454 3167 -398
rect 3223 -454 3309 -398
rect 3365 -454 3451 -398
rect 3507 -454 3593 -398
rect 3649 -454 3735 -398
rect 3791 -454 3877 -398
rect 3933 -454 4019 -398
rect 4075 -454 4161 -398
rect 4217 -454 4303 -398
rect 4359 -454 4445 -398
rect 4501 -454 4587 -398
rect 4643 -454 4729 -398
rect 4785 -454 4871 -398
rect 4927 -454 5013 -398
rect 5069 -454 5155 -398
rect 5211 -454 5297 -398
rect 5353 -454 5439 -398
rect 5495 -454 5581 -398
rect 5637 -454 5723 -398
rect 5779 -454 5865 -398
rect 5921 -454 6007 -398
rect 6063 -454 6149 -398
rect 6205 -454 6291 -398
rect 6347 -454 6433 -398
rect 6489 -454 6575 -398
rect 6631 -454 6717 -398
rect 6773 -454 6859 -398
rect 6915 -454 7001 -398
rect 7057 -454 7143 -398
rect 7199 -454 7285 -398
rect 7341 -454 7351 -398
rect -7351 -540 7351 -454
rect -7351 -596 -7341 -540
rect -7285 -596 -7199 -540
rect -7143 -596 -7057 -540
rect -7001 -596 -6915 -540
rect -6859 -596 -6773 -540
rect -6717 -596 -6631 -540
rect -6575 -596 -6489 -540
rect -6433 -596 -6347 -540
rect -6291 -596 -6205 -540
rect -6149 -596 -6063 -540
rect -6007 -596 -5921 -540
rect -5865 -596 -5779 -540
rect -5723 -596 -5637 -540
rect -5581 -596 -5495 -540
rect -5439 -596 -5353 -540
rect -5297 -596 -5211 -540
rect -5155 -596 -5069 -540
rect -5013 -596 -4927 -540
rect -4871 -596 -4785 -540
rect -4729 -596 -4643 -540
rect -4587 -596 -4501 -540
rect -4445 -596 -4359 -540
rect -4303 -596 -4217 -540
rect -4161 -596 -4075 -540
rect -4019 -596 -3933 -540
rect -3877 -596 -3791 -540
rect -3735 -596 -3649 -540
rect -3593 -596 -3507 -540
rect -3451 -596 -3365 -540
rect -3309 -596 -3223 -540
rect -3167 -596 -3081 -540
rect -3025 -596 -2939 -540
rect -2883 -596 -2797 -540
rect -2741 -596 -2655 -540
rect -2599 -596 -2513 -540
rect -2457 -596 -2371 -540
rect -2315 -596 -2229 -540
rect -2173 -596 -2087 -540
rect -2031 -596 -1945 -540
rect -1889 -596 -1803 -540
rect -1747 -596 -1661 -540
rect -1605 -596 -1519 -540
rect -1463 -596 -1377 -540
rect -1321 -596 -1235 -540
rect -1179 -596 -1093 -540
rect -1037 -596 -951 -540
rect -895 -596 -809 -540
rect -753 -596 -667 -540
rect -611 -596 -525 -540
rect -469 -596 -383 -540
rect -327 -596 -241 -540
rect -185 -596 -99 -540
rect -43 -596 43 -540
rect 99 -596 185 -540
rect 241 -596 327 -540
rect 383 -596 469 -540
rect 525 -596 611 -540
rect 667 -596 753 -540
rect 809 -596 895 -540
rect 951 -596 1037 -540
rect 1093 -596 1179 -540
rect 1235 -596 1321 -540
rect 1377 -596 1463 -540
rect 1519 -596 1605 -540
rect 1661 -596 1747 -540
rect 1803 -596 1889 -540
rect 1945 -596 2031 -540
rect 2087 -596 2173 -540
rect 2229 -596 2315 -540
rect 2371 -596 2457 -540
rect 2513 -596 2599 -540
rect 2655 -596 2741 -540
rect 2797 -596 2883 -540
rect 2939 -596 3025 -540
rect 3081 -596 3167 -540
rect 3223 -596 3309 -540
rect 3365 -596 3451 -540
rect 3507 -596 3593 -540
rect 3649 -596 3735 -540
rect 3791 -596 3877 -540
rect 3933 -596 4019 -540
rect 4075 -596 4161 -540
rect 4217 -596 4303 -540
rect 4359 -596 4445 -540
rect 4501 -596 4587 -540
rect 4643 -596 4729 -540
rect 4785 -596 4871 -540
rect 4927 -596 5013 -540
rect 5069 -596 5155 -540
rect 5211 -596 5297 -540
rect 5353 -596 5439 -540
rect 5495 -596 5581 -540
rect 5637 -596 5723 -540
rect 5779 -596 5865 -540
rect 5921 -596 6007 -540
rect 6063 -596 6149 -540
rect 6205 -596 6291 -540
rect 6347 -596 6433 -540
rect 6489 -596 6575 -540
rect 6631 -596 6717 -540
rect 6773 -596 6859 -540
rect 6915 -596 7001 -540
rect 7057 -596 7143 -540
rect 7199 -596 7285 -540
rect 7341 -596 7351 -540
rect -7351 -682 7351 -596
rect -7351 -738 -7341 -682
rect -7285 -738 -7199 -682
rect -7143 -738 -7057 -682
rect -7001 -738 -6915 -682
rect -6859 -738 -6773 -682
rect -6717 -738 -6631 -682
rect -6575 -738 -6489 -682
rect -6433 -738 -6347 -682
rect -6291 -738 -6205 -682
rect -6149 -738 -6063 -682
rect -6007 -738 -5921 -682
rect -5865 -738 -5779 -682
rect -5723 -738 -5637 -682
rect -5581 -738 -5495 -682
rect -5439 -738 -5353 -682
rect -5297 -738 -5211 -682
rect -5155 -738 -5069 -682
rect -5013 -738 -4927 -682
rect -4871 -738 -4785 -682
rect -4729 -738 -4643 -682
rect -4587 -738 -4501 -682
rect -4445 -738 -4359 -682
rect -4303 -738 -4217 -682
rect -4161 -738 -4075 -682
rect -4019 -738 -3933 -682
rect -3877 -738 -3791 -682
rect -3735 -738 -3649 -682
rect -3593 -738 -3507 -682
rect -3451 -738 -3365 -682
rect -3309 -738 -3223 -682
rect -3167 -738 -3081 -682
rect -3025 -738 -2939 -682
rect -2883 -738 -2797 -682
rect -2741 -738 -2655 -682
rect -2599 -738 -2513 -682
rect -2457 -738 -2371 -682
rect -2315 -738 -2229 -682
rect -2173 -738 -2087 -682
rect -2031 -738 -1945 -682
rect -1889 -738 -1803 -682
rect -1747 -738 -1661 -682
rect -1605 -738 -1519 -682
rect -1463 -738 -1377 -682
rect -1321 -738 -1235 -682
rect -1179 -738 -1093 -682
rect -1037 -738 -951 -682
rect -895 -738 -809 -682
rect -753 -738 -667 -682
rect -611 -738 -525 -682
rect -469 -738 -383 -682
rect -327 -738 -241 -682
rect -185 -738 -99 -682
rect -43 -738 43 -682
rect 99 -738 185 -682
rect 241 -738 327 -682
rect 383 -738 469 -682
rect 525 -738 611 -682
rect 667 -738 753 -682
rect 809 -738 895 -682
rect 951 -738 1037 -682
rect 1093 -738 1179 -682
rect 1235 -738 1321 -682
rect 1377 -738 1463 -682
rect 1519 -738 1605 -682
rect 1661 -738 1747 -682
rect 1803 -738 1889 -682
rect 1945 -738 2031 -682
rect 2087 -738 2173 -682
rect 2229 -738 2315 -682
rect 2371 -738 2457 -682
rect 2513 -738 2599 -682
rect 2655 -738 2741 -682
rect 2797 -738 2883 -682
rect 2939 -738 3025 -682
rect 3081 -738 3167 -682
rect 3223 -738 3309 -682
rect 3365 -738 3451 -682
rect 3507 -738 3593 -682
rect 3649 -738 3735 -682
rect 3791 -738 3877 -682
rect 3933 -738 4019 -682
rect 4075 -738 4161 -682
rect 4217 -738 4303 -682
rect 4359 -738 4445 -682
rect 4501 -738 4587 -682
rect 4643 -738 4729 -682
rect 4785 -738 4871 -682
rect 4927 -738 5013 -682
rect 5069 -738 5155 -682
rect 5211 -738 5297 -682
rect 5353 -738 5439 -682
rect 5495 -738 5581 -682
rect 5637 -738 5723 -682
rect 5779 -738 5865 -682
rect 5921 -738 6007 -682
rect 6063 -738 6149 -682
rect 6205 -738 6291 -682
rect 6347 -738 6433 -682
rect 6489 -738 6575 -682
rect 6631 -738 6717 -682
rect 6773 -738 6859 -682
rect 6915 -738 7001 -682
rect 7057 -738 7143 -682
rect 7199 -738 7285 -682
rect 7341 -738 7351 -682
rect -7351 -824 7351 -738
rect -7351 -880 -7341 -824
rect -7285 -880 -7199 -824
rect -7143 -880 -7057 -824
rect -7001 -880 -6915 -824
rect -6859 -880 -6773 -824
rect -6717 -880 -6631 -824
rect -6575 -880 -6489 -824
rect -6433 -880 -6347 -824
rect -6291 -880 -6205 -824
rect -6149 -880 -6063 -824
rect -6007 -880 -5921 -824
rect -5865 -880 -5779 -824
rect -5723 -880 -5637 -824
rect -5581 -880 -5495 -824
rect -5439 -880 -5353 -824
rect -5297 -880 -5211 -824
rect -5155 -880 -5069 -824
rect -5013 -880 -4927 -824
rect -4871 -880 -4785 -824
rect -4729 -880 -4643 -824
rect -4587 -880 -4501 -824
rect -4445 -880 -4359 -824
rect -4303 -880 -4217 -824
rect -4161 -880 -4075 -824
rect -4019 -880 -3933 -824
rect -3877 -880 -3791 -824
rect -3735 -880 -3649 -824
rect -3593 -880 -3507 -824
rect -3451 -880 -3365 -824
rect -3309 -880 -3223 -824
rect -3167 -880 -3081 -824
rect -3025 -880 -2939 -824
rect -2883 -880 -2797 -824
rect -2741 -880 -2655 -824
rect -2599 -880 -2513 -824
rect -2457 -880 -2371 -824
rect -2315 -880 -2229 -824
rect -2173 -880 -2087 -824
rect -2031 -880 -1945 -824
rect -1889 -880 -1803 -824
rect -1747 -880 -1661 -824
rect -1605 -880 -1519 -824
rect -1463 -880 -1377 -824
rect -1321 -880 -1235 -824
rect -1179 -880 -1093 -824
rect -1037 -880 -951 -824
rect -895 -880 -809 -824
rect -753 -880 -667 -824
rect -611 -880 -525 -824
rect -469 -880 -383 -824
rect -327 -880 -241 -824
rect -185 -880 -99 -824
rect -43 -880 43 -824
rect 99 -880 185 -824
rect 241 -880 327 -824
rect 383 -880 469 -824
rect 525 -880 611 -824
rect 667 -880 753 -824
rect 809 -880 895 -824
rect 951 -880 1037 -824
rect 1093 -880 1179 -824
rect 1235 -880 1321 -824
rect 1377 -880 1463 -824
rect 1519 -880 1605 -824
rect 1661 -880 1747 -824
rect 1803 -880 1889 -824
rect 1945 -880 2031 -824
rect 2087 -880 2173 -824
rect 2229 -880 2315 -824
rect 2371 -880 2457 -824
rect 2513 -880 2599 -824
rect 2655 -880 2741 -824
rect 2797 -880 2883 -824
rect 2939 -880 3025 -824
rect 3081 -880 3167 -824
rect 3223 -880 3309 -824
rect 3365 -880 3451 -824
rect 3507 -880 3593 -824
rect 3649 -880 3735 -824
rect 3791 -880 3877 -824
rect 3933 -880 4019 -824
rect 4075 -880 4161 -824
rect 4217 -880 4303 -824
rect 4359 -880 4445 -824
rect 4501 -880 4587 -824
rect 4643 -880 4729 -824
rect 4785 -880 4871 -824
rect 4927 -880 5013 -824
rect 5069 -880 5155 -824
rect 5211 -880 5297 -824
rect 5353 -880 5439 -824
rect 5495 -880 5581 -824
rect 5637 -880 5723 -824
rect 5779 -880 5865 -824
rect 5921 -880 6007 -824
rect 6063 -880 6149 -824
rect 6205 -880 6291 -824
rect 6347 -880 6433 -824
rect 6489 -880 6575 -824
rect 6631 -880 6717 -824
rect 6773 -880 6859 -824
rect 6915 -880 7001 -824
rect 7057 -880 7143 -824
rect 7199 -880 7285 -824
rect 7341 -880 7351 -824
rect -7351 -966 7351 -880
rect -7351 -1022 -7341 -966
rect -7285 -1022 -7199 -966
rect -7143 -1022 -7057 -966
rect -7001 -1022 -6915 -966
rect -6859 -1022 -6773 -966
rect -6717 -1022 -6631 -966
rect -6575 -1022 -6489 -966
rect -6433 -1022 -6347 -966
rect -6291 -1022 -6205 -966
rect -6149 -1022 -6063 -966
rect -6007 -1022 -5921 -966
rect -5865 -1022 -5779 -966
rect -5723 -1022 -5637 -966
rect -5581 -1022 -5495 -966
rect -5439 -1022 -5353 -966
rect -5297 -1022 -5211 -966
rect -5155 -1022 -5069 -966
rect -5013 -1022 -4927 -966
rect -4871 -1022 -4785 -966
rect -4729 -1022 -4643 -966
rect -4587 -1022 -4501 -966
rect -4445 -1022 -4359 -966
rect -4303 -1022 -4217 -966
rect -4161 -1022 -4075 -966
rect -4019 -1022 -3933 -966
rect -3877 -1022 -3791 -966
rect -3735 -1022 -3649 -966
rect -3593 -1022 -3507 -966
rect -3451 -1022 -3365 -966
rect -3309 -1022 -3223 -966
rect -3167 -1022 -3081 -966
rect -3025 -1022 -2939 -966
rect -2883 -1022 -2797 -966
rect -2741 -1022 -2655 -966
rect -2599 -1022 -2513 -966
rect -2457 -1022 -2371 -966
rect -2315 -1022 -2229 -966
rect -2173 -1022 -2087 -966
rect -2031 -1022 -1945 -966
rect -1889 -1022 -1803 -966
rect -1747 -1022 -1661 -966
rect -1605 -1022 -1519 -966
rect -1463 -1022 -1377 -966
rect -1321 -1022 -1235 -966
rect -1179 -1022 -1093 -966
rect -1037 -1022 -951 -966
rect -895 -1022 -809 -966
rect -753 -1022 -667 -966
rect -611 -1022 -525 -966
rect -469 -1022 -383 -966
rect -327 -1022 -241 -966
rect -185 -1022 -99 -966
rect -43 -1022 43 -966
rect 99 -1022 185 -966
rect 241 -1022 327 -966
rect 383 -1022 469 -966
rect 525 -1022 611 -966
rect 667 -1022 753 -966
rect 809 -1022 895 -966
rect 951 -1022 1037 -966
rect 1093 -1022 1179 -966
rect 1235 -1022 1321 -966
rect 1377 -1022 1463 -966
rect 1519 -1022 1605 -966
rect 1661 -1022 1747 -966
rect 1803 -1022 1889 -966
rect 1945 -1022 2031 -966
rect 2087 -1022 2173 -966
rect 2229 -1022 2315 -966
rect 2371 -1022 2457 -966
rect 2513 -1022 2599 -966
rect 2655 -1022 2741 -966
rect 2797 -1022 2883 -966
rect 2939 -1022 3025 -966
rect 3081 -1022 3167 -966
rect 3223 -1022 3309 -966
rect 3365 -1022 3451 -966
rect 3507 -1022 3593 -966
rect 3649 -1022 3735 -966
rect 3791 -1022 3877 -966
rect 3933 -1022 4019 -966
rect 4075 -1022 4161 -966
rect 4217 -1022 4303 -966
rect 4359 -1022 4445 -966
rect 4501 -1022 4587 -966
rect 4643 -1022 4729 -966
rect 4785 -1022 4871 -966
rect 4927 -1022 5013 -966
rect 5069 -1022 5155 -966
rect 5211 -1022 5297 -966
rect 5353 -1022 5439 -966
rect 5495 -1022 5581 -966
rect 5637 -1022 5723 -966
rect 5779 -1022 5865 -966
rect 5921 -1022 6007 -966
rect 6063 -1022 6149 -966
rect 6205 -1022 6291 -966
rect 6347 -1022 6433 -966
rect 6489 -1022 6575 -966
rect 6631 -1022 6717 -966
rect 6773 -1022 6859 -966
rect 6915 -1022 7001 -966
rect 7057 -1022 7143 -966
rect 7199 -1022 7285 -966
rect 7341 -1022 7351 -966
rect -7351 -1108 7351 -1022
rect -7351 -1164 -7341 -1108
rect -7285 -1164 -7199 -1108
rect -7143 -1164 -7057 -1108
rect -7001 -1164 -6915 -1108
rect -6859 -1164 -6773 -1108
rect -6717 -1164 -6631 -1108
rect -6575 -1164 -6489 -1108
rect -6433 -1164 -6347 -1108
rect -6291 -1164 -6205 -1108
rect -6149 -1164 -6063 -1108
rect -6007 -1164 -5921 -1108
rect -5865 -1164 -5779 -1108
rect -5723 -1164 -5637 -1108
rect -5581 -1164 -5495 -1108
rect -5439 -1164 -5353 -1108
rect -5297 -1164 -5211 -1108
rect -5155 -1164 -5069 -1108
rect -5013 -1164 -4927 -1108
rect -4871 -1164 -4785 -1108
rect -4729 -1164 -4643 -1108
rect -4587 -1164 -4501 -1108
rect -4445 -1164 -4359 -1108
rect -4303 -1164 -4217 -1108
rect -4161 -1164 -4075 -1108
rect -4019 -1164 -3933 -1108
rect -3877 -1164 -3791 -1108
rect -3735 -1164 -3649 -1108
rect -3593 -1164 -3507 -1108
rect -3451 -1164 -3365 -1108
rect -3309 -1164 -3223 -1108
rect -3167 -1164 -3081 -1108
rect -3025 -1164 -2939 -1108
rect -2883 -1164 -2797 -1108
rect -2741 -1164 -2655 -1108
rect -2599 -1164 -2513 -1108
rect -2457 -1164 -2371 -1108
rect -2315 -1164 -2229 -1108
rect -2173 -1164 -2087 -1108
rect -2031 -1164 -1945 -1108
rect -1889 -1164 -1803 -1108
rect -1747 -1164 -1661 -1108
rect -1605 -1164 -1519 -1108
rect -1463 -1164 -1377 -1108
rect -1321 -1164 -1235 -1108
rect -1179 -1164 -1093 -1108
rect -1037 -1164 -951 -1108
rect -895 -1164 -809 -1108
rect -753 -1164 -667 -1108
rect -611 -1164 -525 -1108
rect -469 -1164 -383 -1108
rect -327 -1164 -241 -1108
rect -185 -1164 -99 -1108
rect -43 -1164 43 -1108
rect 99 -1164 185 -1108
rect 241 -1164 327 -1108
rect 383 -1164 469 -1108
rect 525 -1164 611 -1108
rect 667 -1164 753 -1108
rect 809 -1164 895 -1108
rect 951 -1164 1037 -1108
rect 1093 -1164 1179 -1108
rect 1235 -1164 1321 -1108
rect 1377 -1164 1463 -1108
rect 1519 -1164 1605 -1108
rect 1661 -1164 1747 -1108
rect 1803 -1164 1889 -1108
rect 1945 -1164 2031 -1108
rect 2087 -1164 2173 -1108
rect 2229 -1164 2315 -1108
rect 2371 -1164 2457 -1108
rect 2513 -1164 2599 -1108
rect 2655 -1164 2741 -1108
rect 2797 -1164 2883 -1108
rect 2939 -1164 3025 -1108
rect 3081 -1164 3167 -1108
rect 3223 -1164 3309 -1108
rect 3365 -1164 3451 -1108
rect 3507 -1164 3593 -1108
rect 3649 -1164 3735 -1108
rect 3791 -1164 3877 -1108
rect 3933 -1164 4019 -1108
rect 4075 -1164 4161 -1108
rect 4217 -1164 4303 -1108
rect 4359 -1164 4445 -1108
rect 4501 -1164 4587 -1108
rect 4643 -1164 4729 -1108
rect 4785 -1164 4871 -1108
rect 4927 -1164 5013 -1108
rect 5069 -1164 5155 -1108
rect 5211 -1164 5297 -1108
rect 5353 -1164 5439 -1108
rect 5495 -1164 5581 -1108
rect 5637 -1164 5723 -1108
rect 5779 -1164 5865 -1108
rect 5921 -1164 6007 -1108
rect 6063 -1164 6149 -1108
rect 6205 -1164 6291 -1108
rect 6347 -1164 6433 -1108
rect 6489 -1164 6575 -1108
rect 6631 -1164 6717 -1108
rect 6773 -1164 6859 -1108
rect 6915 -1164 7001 -1108
rect 7057 -1164 7143 -1108
rect 7199 -1164 7285 -1108
rect 7341 -1164 7351 -1108
rect -7351 -1250 7351 -1164
rect -7351 -1306 -7341 -1250
rect -7285 -1306 -7199 -1250
rect -7143 -1306 -7057 -1250
rect -7001 -1306 -6915 -1250
rect -6859 -1306 -6773 -1250
rect -6717 -1306 -6631 -1250
rect -6575 -1306 -6489 -1250
rect -6433 -1306 -6347 -1250
rect -6291 -1306 -6205 -1250
rect -6149 -1306 -6063 -1250
rect -6007 -1306 -5921 -1250
rect -5865 -1306 -5779 -1250
rect -5723 -1306 -5637 -1250
rect -5581 -1306 -5495 -1250
rect -5439 -1306 -5353 -1250
rect -5297 -1306 -5211 -1250
rect -5155 -1306 -5069 -1250
rect -5013 -1306 -4927 -1250
rect -4871 -1306 -4785 -1250
rect -4729 -1306 -4643 -1250
rect -4587 -1306 -4501 -1250
rect -4445 -1306 -4359 -1250
rect -4303 -1306 -4217 -1250
rect -4161 -1306 -4075 -1250
rect -4019 -1306 -3933 -1250
rect -3877 -1306 -3791 -1250
rect -3735 -1306 -3649 -1250
rect -3593 -1306 -3507 -1250
rect -3451 -1306 -3365 -1250
rect -3309 -1306 -3223 -1250
rect -3167 -1306 -3081 -1250
rect -3025 -1306 -2939 -1250
rect -2883 -1306 -2797 -1250
rect -2741 -1306 -2655 -1250
rect -2599 -1306 -2513 -1250
rect -2457 -1306 -2371 -1250
rect -2315 -1306 -2229 -1250
rect -2173 -1306 -2087 -1250
rect -2031 -1306 -1945 -1250
rect -1889 -1306 -1803 -1250
rect -1747 -1306 -1661 -1250
rect -1605 -1306 -1519 -1250
rect -1463 -1306 -1377 -1250
rect -1321 -1306 -1235 -1250
rect -1179 -1306 -1093 -1250
rect -1037 -1306 -951 -1250
rect -895 -1306 -809 -1250
rect -753 -1306 -667 -1250
rect -611 -1306 -525 -1250
rect -469 -1306 -383 -1250
rect -327 -1306 -241 -1250
rect -185 -1306 -99 -1250
rect -43 -1306 43 -1250
rect 99 -1306 185 -1250
rect 241 -1306 327 -1250
rect 383 -1306 469 -1250
rect 525 -1306 611 -1250
rect 667 -1306 753 -1250
rect 809 -1306 895 -1250
rect 951 -1306 1037 -1250
rect 1093 -1306 1179 -1250
rect 1235 -1306 1321 -1250
rect 1377 -1306 1463 -1250
rect 1519 -1306 1605 -1250
rect 1661 -1306 1747 -1250
rect 1803 -1306 1889 -1250
rect 1945 -1306 2031 -1250
rect 2087 -1306 2173 -1250
rect 2229 -1306 2315 -1250
rect 2371 -1306 2457 -1250
rect 2513 -1306 2599 -1250
rect 2655 -1306 2741 -1250
rect 2797 -1306 2883 -1250
rect 2939 -1306 3025 -1250
rect 3081 -1306 3167 -1250
rect 3223 -1306 3309 -1250
rect 3365 -1306 3451 -1250
rect 3507 -1306 3593 -1250
rect 3649 -1306 3735 -1250
rect 3791 -1306 3877 -1250
rect 3933 -1306 4019 -1250
rect 4075 -1306 4161 -1250
rect 4217 -1306 4303 -1250
rect 4359 -1306 4445 -1250
rect 4501 -1306 4587 -1250
rect 4643 -1306 4729 -1250
rect 4785 -1306 4871 -1250
rect 4927 -1306 5013 -1250
rect 5069 -1306 5155 -1250
rect 5211 -1306 5297 -1250
rect 5353 -1306 5439 -1250
rect 5495 -1306 5581 -1250
rect 5637 -1306 5723 -1250
rect 5779 -1306 5865 -1250
rect 5921 -1306 6007 -1250
rect 6063 -1306 6149 -1250
rect 6205 -1306 6291 -1250
rect 6347 -1306 6433 -1250
rect 6489 -1306 6575 -1250
rect 6631 -1306 6717 -1250
rect 6773 -1306 6859 -1250
rect 6915 -1306 7001 -1250
rect 7057 -1306 7143 -1250
rect 7199 -1306 7285 -1250
rect 7341 -1306 7351 -1250
rect -7351 -1392 7351 -1306
rect -7351 -1448 -7341 -1392
rect -7285 -1448 -7199 -1392
rect -7143 -1448 -7057 -1392
rect -7001 -1448 -6915 -1392
rect -6859 -1448 -6773 -1392
rect -6717 -1448 -6631 -1392
rect -6575 -1448 -6489 -1392
rect -6433 -1448 -6347 -1392
rect -6291 -1448 -6205 -1392
rect -6149 -1448 -6063 -1392
rect -6007 -1448 -5921 -1392
rect -5865 -1448 -5779 -1392
rect -5723 -1448 -5637 -1392
rect -5581 -1448 -5495 -1392
rect -5439 -1448 -5353 -1392
rect -5297 -1448 -5211 -1392
rect -5155 -1448 -5069 -1392
rect -5013 -1448 -4927 -1392
rect -4871 -1448 -4785 -1392
rect -4729 -1448 -4643 -1392
rect -4587 -1448 -4501 -1392
rect -4445 -1448 -4359 -1392
rect -4303 -1448 -4217 -1392
rect -4161 -1448 -4075 -1392
rect -4019 -1448 -3933 -1392
rect -3877 -1448 -3791 -1392
rect -3735 -1448 -3649 -1392
rect -3593 -1448 -3507 -1392
rect -3451 -1448 -3365 -1392
rect -3309 -1448 -3223 -1392
rect -3167 -1448 -3081 -1392
rect -3025 -1448 -2939 -1392
rect -2883 -1448 -2797 -1392
rect -2741 -1448 -2655 -1392
rect -2599 -1448 -2513 -1392
rect -2457 -1448 -2371 -1392
rect -2315 -1448 -2229 -1392
rect -2173 -1448 -2087 -1392
rect -2031 -1448 -1945 -1392
rect -1889 -1448 -1803 -1392
rect -1747 -1448 -1661 -1392
rect -1605 -1448 -1519 -1392
rect -1463 -1448 -1377 -1392
rect -1321 -1448 -1235 -1392
rect -1179 -1448 -1093 -1392
rect -1037 -1448 -951 -1392
rect -895 -1448 -809 -1392
rect -753 -1448 -667 -1392
rect -611 -1448 -525 -1392
rect -469 -1448 -383 -1392
rect -327 -1448 -241 -1392
rect -185 -1448 -99 -1392
rect -43 -1448 43 -1392
rect 99 -1448 185 -1392
rect 241 -1448 327 -1392
rect 383 -1448 469 -1392
rect 525 -1448 611 -1392
rect 667 -1448 753 -1392
rect 809 -1448 895 -1392
rect 951 -1448 1037 -1392
rect 1093 -1448 1179 -1392
rect 1235 -1448 1321 -1392
rect 1377 -1448 1463 -1392
rect 1519 -1448 1605 -1392
rect 1661 -1448 1747 -1392
rect 1803 -1448 1889 -1392
rect 1945 -1448 2031 -1392
rect 2087 -1448 2173 -1392
rect 2229 -1448 2315 -1392
rect 2371 -1448 2457 -1392
rect 2513 -1448 2599 -1392
rect 2655 -1448 2741 -1392
rect 2797 -1448 2883 -1392
rect 2939 -1448 3025 -1392
rect 3081 -1448 3167 -1392
rect 3223 -1448 3309 -1392
rect 3365 -1448 3451 -1392
rect 3507 -1448 3593 -1392
rect 3649 -1448 3735 -1392
rect 3791 -1448 3877 -1392
rect 3933 -1448 4019 -1392
rect 4075 -1448 4161 -1392
rect 4217 -1448 4303 -1392
rect 4359 -1448 4445 -1392
rect 4501 -1448 4587 -1392
rect 4643 -1448 4729 -1392
rect 4785 -1448 4871 -1392
rect 4927 -1448 5013 -1392
rect 5069 -1448 5155 -1392
rect 5211 -1448 5297 -1392
rect 5353 -1448 5439 -1392
rect 5495 -1448 5581 -1392
rect 5637 -1448 5723 -1392
rect 5779 -1448 5865 -1392
rect 5921 -1448 6007 -1392
rect 6063 -1448 6149 -1392
rect 6205 -1448 6291 -1392
rect 6347 -1448 6433 -1392
rect 6489 -1448 6575 -1392
rect 6631 -1448 6717 -1392
rect 6773 -1448 6859 -1392
rect 6915 -1448 7001 -1392
rect 7057 -1448 7143 -1392
rect 7199 -1448 7285 -1392
rect 7341 -1448 7351 -1392
rect -7351 -1458 7351 -1448
<< via3 >>
rect -7341 1392 -7285 1448
rect -7199 1392 -7143 1448
rect -7057 1392 -7001 1448
rect -6915 1392 -6859 1448
rect -6773 1392 -6717 1448
rect -6631 1392 -6575 1448
rect -6489 1392 -6433 1448
rect -6347 1392 -6291 1448
rect -6205 1392 -6149 1448
rect -6063 1392 -6007 1448
rect -5921 1392 -5865 1448
rect -5779 1392 -5723 1448
rect -5637 1392 -5581 1448
rect -5495 1392 -5439 1448
rect -5353 1392 -5297 1448
rect -5211 1392 -5155 1448
rect -5069 1392 -5013 1448
rect -4927 1392 -4871 1448
rect -4785 1392 -4729 1448
rect -4643 1392 -4587 1448
rect -4501 1392 -4445 1448
rect -4359 1392 -4303 1448
rect -4217 1392 -4161 1448
rect -4075 1392 -4019 1448
rect -3933 1392 -3877 1448
rect -3791 1392 -3735 1448
rect -3649 1392 -3593 1448
rect -3507 1392 -3451 1448
rect -3365 1392 -3309 1448
rect -3223 1392 -3167 1448
rect -3081 1392 -3025 1448
rect -2939 1392 -2883 1448
rect -2797 1392 -2741 1448
rect -2655 1392 -2599 1448
rect -2513 1392 -2457 1448
rect -2371 1392 -2315 1448
rect -2229 1392 -2173 1448
rect -2087 1392 -2031 1448
rect -1945 1392 -1889 1448
rect -1803 1392 -1747 1448
rect -1661 1392 -1605 1448
rect -1519 1392 -1463 1448
rect -1377 1392 -1321 1448
rect -1235 1392 -1179 1448
rect -1093 1392 -1037 1448
rect -951 1392 -895 1448
rect -809 1392 -753 1448
rect -667 1392 -611 1448
rect -525 1392 -469 1448
rect -383 1392 -327 1448
rect -241 1392 -185 1448
rect -99 1392 -43 1448
rect 43 1392 99 1448
rect 185 1392 241 1448
rect 327 1392 383 1448
rect 469 1392 525 1448
rect 611 1392 667 1448
rect 753 1392 809 1448
rect 895 1392 951 1448
rect 1037 1392 1093 1448
rect 1179 1392 1235 1448
rect 1321 1392 1377 1448
rect 1463 1392 1519 1448
rect 1605 1392 1661 1448
rect 1747 1392 1803 1448
rect 1889 1392 1945 1448
rect 2031 1392 2087 1448
rect 2173 1392 2229 1448
rect 2315 1392 2371 1448
rect 2457 1392 2513 1448
rect 2599 1392 2655 1448
rect 2741 1392 2797 1448
rect 2883 1392 2939 1448
rect 3025 1392 3081 1448
rect 3167 1392 3223 1448
rect 3309 1392 3365 1448
rect 3451 1392 3507 1448
rect 3593 1392 3649 1448
rect 3735 1392 3791 1448
rect 3877 1392 3933 1448
rect 4019 1392 4075 1448
rect 4161 1392 4217 1448
rect 4303 1392 4359 1448
rect 4445 1392 4501 1448
rect 4587 1392 4643 1448
rect 4729 1392 4785 1448
rect 4871 1392 4927 1448
rect 5013 1392 5069 1448
rect 5155 1392 5211 1448
rect 5297 1392 5353 1448
rect 5439 1392 5495 1448
rect 5581 1392 5637 1448
rect 5723 1392 5779 1448
rect 5865 1392 5921 1448
rect 6007 1392 6063 1448
rect 6149 1392 6205 1448
rect 6291 1392 6347 1448
rect 6433 1392 6489 1448
rect 6575 1392 6631 1448
rect 6717 1392 6773 1448
rect 6859 1392 6915 1448
rect 7001 1392 7057 1448
rect 7143 1392 7199 1448
rect 7285 1392 7341 1448
rect -7341 1250 -7285 1306
rect -7199 1250 -7143 1306
rect -7057 1250 -7001 1306
rect -6915 1250 -6859 1306
rect -6773 1250 -6717 1306
rect -6631 1250 -6575 1306
rect -6489 1250 -6433 1306
rect -6347 1250 -6291 1306
rect -6205 1250 -6149 1306
rect -6063 1250 -6007 1306
rect -5921 1250 -5865 1306
rect -5779 1250 -5723 1306
rect -5637 1250 -5581 1306
rect -5495 1250 -5439 1306
rect -5353 1250 -5297 1306
rect -5211 1250 -5155 1306
rect -5069 1250 -5013 1306
rect -4927 1250 -4871 1306
rect -4785 1250 -4729 1306
rect -4643 1250 -4587 1306
rect -4501 1250 -4445 1306
rect -4359 1250 -4303 1306
rect -4217 1250 -4161 1306
rect -4075 1250 -4019 1306
rect -3933 1250 -3877 1306
rect -3791 1250 -3735 1306
rect -3649 1250 -3593 1306
rect -3507 1250 -3451 1306
rect -3365 1250 -3309 1306
rect -3223 1250 -3167 1306
rect -3081 1250 -3025 1306
rect -2939 1250 -2883 1306
rect -2797 1250 -2741 1306
rect -2655 1250 -2599 1306
rect -2513 1250 -2457 1306
rect -2371 1250 -2315 1306
rect -2229 1250 -2173 1306
rect -2087 1250 -2031 1306
rect -1945 1250 -1889 1306
rect -1803 1250 -1747 1306
rect -1661 1250 -1605 1306
rect -1519 1250 -1463 1306
rect -1377 1250 -1321 1306
rect -1235 1250 -1179 1306
rect -1093 1250 -1037 1306
rect -951 1250 -895 1306
rect -809 1250 -753 1306
rect -667 1250 -611 1306
rect -525 1250 -469 1306
rect -383 1250 -327 1306
rect -241 1250 -185 1306
rect -99 1250 -43 1306
rect 43 1250 99 1306
rect 185 1250 241 1306
rect 327 1250 383 1306
rect 469 1250 525 1306
rect 611 1250 667 1306
rect 753 1250 809 1306
rect 895 1250 951 1306
rect 1037 1250 1093 1306
rect 1179 1250 1235 1306
rect 1321 1250 1377 1306
rect 1463 1250 1519 1306
rect 1605 1250 1661 1306
rect 1747 1250 1803 1306
rect 1889 1250 1945 1306
rect 2031 1250 2087 1306
rect 2173 1250 2229 1306
rect 2315 1250 2371 1306
rect 2457 1250 2513 1306
rect 2599 1250 2655 1306
rect 2741 1250 2797 1306
rect 2883 1250 2939 1306
rect 3025 1250 3081 1306
rect 3167 1250 3223 1306
rect 3309 1250 3365 1306
rect 3451 1250 3507 1306
rect 3593 1250 3649 1306
rect 3735 1250 3791 1306
rect 3877 1250 3933 1306
rect 4019 1250 4075 1306
rect 4161 1250 4217 1306
rect 4303 1250 4359 1306
rect 4445 1250 4501 1306
rect 4587 1250 4643 1306
rect 4729 1250 4785 1306
rect 4871 1250 4927 1306
rect 5013 1250 5069 1306
rect 5155 1250 5211 1306
rect 5297 1250 5353 1306
rect 5439 1250 5495 1306
rect 5581 1250 5637 1306
rect 5723 1250 5779 1306
rect 5865 1250 5921 1306
rect 6007 1250 6063 1306
rect 6149 1250 6205 1306
rect 6291 1250 6347 1306
rect 6433 1250 6489 1306
rect 6575 1250 6631 1306
rect 6717 1250 6773 1306
rect 6859 1250 6915 1306
rect 7001 1250 7057 1306
rect 7143 1250 7199 1306
rect 7285 1250 7341 1306
rect -7341 1108 -7285 1164
rect -7199 1108 -7143 1164
rect -7057 1108 -7001 1164
rect -6915 1108 -6859 1164
rect -6773 1108 -6717 1164
rect -6631 1108 -6575 1164
rect -6489 1108 -6433 1164
rect -6347 1108 -6291 1164
rect -6205 1108 -6149 1164
rect -6063 1108 -6007 1164
rect -5921 1108 -5865 1164
rect -5779 1108 -5723 1164
rect -5637 1108 -5581 1164
rect -5495 1108 -5439 1164
rect -5353 1108 -5297 1164
rect -5211 1108 -5155 1164
rect -5069 1108 -5013 1164
rect -4927 1108 -4871 1164
rect -4785 1108 -4729 1164
rect -4643 1108 -4587 1164
rect -4501 1108 -4445 1164
rect -4359 1108 -4303 1164
rect -4217 1108 -4161 1164
rect -4075 1108 -4019 1164
rect -3933 1108 -3877 1164
rect -3791 1108 -3735 1164
rect -3649 1108 -3593 1164
rect -3507 1108 -3451 1164
rect -3365 1108 -3309 1164
rect -3223 1108 -3167 1164
rect -3081 1108 -3025 1164
rect -2939 1108 -2883 1164
rect -2797 1108 -2741 1164
rect -2655 1108 -2599 1164
rect -2513 1108 -2457 1164
rect -2371 1108 -2315 1164
rect -2229 1108 -2173 1164
rect -2087 1108 -2031 1164
rect -1945 1108 -1889 1164
rect -1803 1108 -1747 1164
rect -1661 1108 -1605 1164
rect -1519 1108 -1463 1164
rect -1377 1108 -1321 1164
rect -1235 1108 -1179 1164
rect -1093 1108 -1037 1164
rect -951 1108 -895 1164
rect -809 1108 -753 1164
rect -667 1108 -611 1164
rect -525 1108 -469 1164
rect -383 1108 -327 1164
rect -241 1108 -185 1164
rect -99 1108 -43 1164
rect 43 1108 99 1164
rect 185 1108 241 1164
rect 327 1108 383 1164
rect 469 1108 525 1164
rect 611 1108 667 1164
rect 753 1108 809 1164
rect 895 1108 951 1164
rect 1037 1108 1093 1164
rect 1179 1108 1235 1164
rect 1321 1108 1377 1164
rect 1463 1108 1519 1164
rect 1605 1108 1661 1164
rect 1747 1108 1803 1164
rect 1889 1108 1945 1164
rect 2031 1108 2087 1164
rect 2173 1108 2229 1164
rect 2315 1108 2371 1164
rect 2457 1108 2513 1164
rect 2599 1108 2655 1164
rect 2741 1108 2797 1164
rect 2883 1108 2939 1164
rect 3025 1108 3081 1164
rect 3167 1108 3223 1164
rect 3309 1108 3365 1164
rect 3451 1108 3507 1164
rect 3593 1108 3649 1164
rect 3735 1108 3791 1164
rect 3877 1108 3933 1164
rect 4019 1108 4075 1164
rect 4161 1108 4217 1164
rect 4303 1108 4359 1164
rect 4445 1108 4501 1164
rect 4587 1108 4643 1164
rect 4729 1108 4785 1164
rect 4871 1108 4927 1164
rect 5013 1108 5069 1164
rect 5155 1108 5211 1164
rect 5297 1108 5353 1164
rect 5439 1108 5495 1164
rect 5581 1108 5637 1164
rect 5723 1108 5779 1164
rect 5865 1108 5921 1164
rect 6007 1108 6063 1164
rect 6149 1108 6205 1164
rect 6291 1108 6347 1164
rect 6433 1108 6489 1164
rect 6575 1108 6631 1164
rect 6717 1108 6773 1164
rect 6859 1108 6915 1164
rect 7001 1108 7057 1164
rect 7143 1108 7199 1164
rect 7285 1108 7341 1164
rect -7341 966 -7285 1022
rect -7199 966 -7143 1022
rect -7057 966 -7001 1022
rect -6915 966 -6859 1022
rect -6773 966 -6717 1022
rect -6631 966 -6575 1022
rect -6489 966 -6433 1022
rect -6347 966 -6291 1022
rect -6205 966 -6149 1022
rect -6063 966 -6007 1022
rect -5921 966 -5865 1022
rect -5779 966 -5723 1022
rect -5637 966 -5581 1022
rect -5495 966 -5439 1022
rect -5353 966 -5297 1022
rect -5211 966 -5155 1022
rect -5069 966 -5013 1022
rect -4927 966 -4871 1022
rect -4785 966 -4729 1022
rect -4643 966 -4587 1022
rect -4501 966 -4445 1022
rect -4359 966 -4303 1022
rect -4217 966 -4161 1022
rect -4075 966 -4019 1022
rect -3933 966 -3877 1022
rect -3791 966 -3735 1022
rect -3649 966 -3593 1022
rect -3507 966 -3451 1022
rect -3365 966 -3309 1022
rect -3223 966 -3167 1022
rect -3081 966 -3025 1022
rect -2939 966 -2883 1022
rect -2797 966 -2741 1022
rect -2655 966 -2599 1022
rect -2513 966 -2457 1022
rect -2371 966 -2315 1022
rect -2229 966 -2173 1022
rect -2087 966 -2031 1022
rect -1945 966 -1889 1022
rect -1803 966 -1747 1022
rect -1661 966 -1605 1022
rect -1519 966 -1463 1022
rect -1377 966 -1321 1022
rect -1235 966 -1179 1022
rect -1093 966 -1037 1022
rect -951 966 -895 1022
rect -809 966 -753 1022
rect -667 966 -611 1022
rect -525 966 -469 1022
rect -383 966 -327 1022
rect -241 966 -185 1022
rect -99 966 -43 1022
rect 43 966 99 1022
rect 185 966 241 1022
rect 327 966 383 1022
rect 469 966 525 1022
rect 611 966 667 1022
rect 753 966 809 1022
rect 895 966 951 1022
rect 1037 966 1093 1022
rect 1179 966 1235 1022
rect 1321 966 1377 1022
rect 1463 966 1519 1022
rect 1605 966 1661 1022
rect 1747 966 1803 1022
rect 1889 966 1945 1022
rect 2031 966 2087 1022
rect 2173 966 2229 1022
rect 2315 966 2371 1022
rect 2457 966 2513 1022
rect 2599 966 2655 1022
rect 2741 966 2797 1022
rect 2883 966 2939 1022
rect 3025 966 3081 1022
rect 3167 966 3223 1022
rect 3309 966 3365 1022
rect 3451 966 3507 1022
rect 3593 966 3649 1022
rect 3735 966 3791 1022
rect 3877 966 3933 1022
rect 4019 966 4075 1022
rect 4161 966 4217 1022
rect 4303 966 4359 1022
rect 4445 966 4501 1022
rect 4587 966 4643 1022
rect 4729 966 4785 1022
rect 4871 966 4927 1022
rect 5013 966 5069 1022
rect 5155 966 5211 1022
rect 5297 966 5353 1022
rect 5439 966 5495 1022
rect 5581 966 5637 1022
rect 5723 966 5779 1022
rect 5865 966 5921 1022
rect 6007 966 6063 1022
rect 6149 966 6205 1022
rect 6291 966 6347 1022
rect 6433 966 6489 1022
rect 6575 966 6631 1022
rect 6717 966 6773 1022
rect 6859 966 6915 1022
rect 7001 966 7057 1022
rect 7143 966 7199 1022
rect 7285 966 7341 1022
rect -7341 824 -7285 880
rect -7199 824 -7143 880
rect -7057 824 -7001 880
rect -6915 824 -6859 880
rect -6773 824 -6717 880
rect -6631 824 -6575 880
rect -6489 824 -6433 880
rect -6347 824 -6291 880
rect -6205 824 -6149 880
rect -6063 824 -6007 880
rect -5921 824 -5865 880
rect -5779 824 -5723 880
rect -5637 824 -5581 880
rect -5495 824 -5439 880
rect -5353 824 -5297 880
rect -5211 824 -5155 880
rect -5069 824 -5013 880
rect -4927 824 -4871 880
rect -4785 824 -4729 880
rect -4643 824 -4587 880
rect -4501 824 -4445 880
rect -4359 824 -4303 880
rect -4217 824 -4161 880
rect -4075 824 -4019 880
rect -3933 824 -3877 880
rect -3791 824 -3735 880
rect -3649 824 -3593 880
rect -3507 824 -3451 880
rect -3365 824 -3309 880
rect -3223 824 -3167 880
rect -3081 824 -3025 880
rect -2939 824 -2883 880
rect -2797 824 -2741 880
rect -2655 824 -2599 880
rect -2513 824 -2457 880
rect -2371 824 -2315 880
rect -2229 824 -2173 880
rect -2087 824 -2031 880
rect -1945 824 -1889 880
rect -1803 824 -1747 880
rect -1661 824 -1605 880
rect -1519 824 -1463 880
rect -1377 824 -1321 880
rect -1235 824 -1179 880
rect -1093 824 -1037 880
rect -951 824 -895 880
rect -809 824 -753 880
rect -667 824 -611 880
rect -525 824 -469 880
rect -383 824 -327 880
rect -241 824 -185 880
rect -99 824 -43 880
rect 43 824 99 880
rect 185 824 241 880
rect 327 824 383 880
rect 469 824 525 880
rect 611 824 667 880
rect 753 824 809 880
rect 895 824 951 880
rect 1037 824 1093 880
rect 1179 824 1235 880
rect 1321 824 1377 880
rect 1463 824 1519 880
rect 1605 824 1661 880
rect 1747 824 1803 880
rect 1889 824 1945 880
rect 2031 824 2087 880
rect 2173 824 2229 880
rect 2315 824 2371 880
rect 2457 824 2513 880
rect 2599 824 2655 880
rect 2741 824 2797 880
rect 2883 824 2939 880
rect 3025 824 3081 880
rect 3167 824 3223 880
rect 3309 824 3365 880
rect 3451 824 3507 880
rect 3593 824 3649 880
rect 3735 824 3791 880
rect 3877 824 3933 880
rect 4019 824 4075 880
rect 4161 824 4217 880
rect 4303 824 4359 880
rect 4445 824 4501 880
rect 4587 824 4643 880
rect 4729 824 4785 880
rect 4871 824 4927 880
rect 5013 824 5069 880
rect 5155 824 5211 880
rect 5297 824 5353 880
rect 5439 824 5495 880
rect 5581 824 5637 880
rect 5723 824 5779 880
rect 5865 824 5921 880
rect 6007 824 6063 880
rect 6149 824 6205 880
rect 6291 824 6347 880
rect 6433 824 6489 880
rect 6575 824 6631 880
rect 6717 824 6773 880
rect 6859 824 6915 880
rect 7001 824 7057 880
rect 7143 824 7199 880
rect 7285 824 7341 880
rect -7341 682 -7285 738
rect -7199 682 -7143 738
rect -7057 682 -7001 738
rect -6915 682 -6859 738
rect -6773 682 -6717 738
rect -6631 682 -6575 738
rect -6489 682 -6433 738
rect -6347 682 -6291 738
rect -6205 682 -6149 738
rect -6063 682 -6007 738
rect -5921 682 -5865 738
rect -5779 682 -5723 738
rect -5637 682 -5581 738
rect -5495 682 -5439 738
rect -5353 682 -5297 738
rect -5211 682 -5155 738
rect -5069 682 -5013 738
rect -4927 682 -4871 738
rect -4785 682 -4729 738
rect -4643 682 -4587 738
rect -4501 682 -4445 738
rect -4359 682 -4303 738
rect -4217 682 -4161 738
rect -4075 682 -4019 738
rect -3933 682 -3877 738
rect -3791 682 -3735 738
rect -3649 682 -3593 738
rect -3507 682 -3451 738
rect -3365 682 -3309 738
rect -3223 682 -3167 738
rect -3081 682 -3025 738
rect -2939 682 -2883 738
rect -2797 682 -2741 738
rect -2655 682 -2599 738
rect -2513 682 -2457 738
rect -2371 682 -2315 738
rect -2229 682 -2173 738
rect -2087 682 -2031 738
rect -1945 682 -1889 738
rect -1803 682 -1747 738
rect -1661 682 -1605 738
rect -1519 682 -1463 738
rect -1377 682 -1321 738
rect -1235 682 -1179 738
rect -1093 682 -1037 738
rect -951 682 -895 738
rect -809 682 -753 738
rect -667 682 -611 738
rect -525 682 -469 738
rect -383 682 -327 738
rect -241 682 -185 738
rect -99 682 -43 738
rect 43 682 99 738
rect 185 682 241 738
rect 327 682 383 738
rect 469 682 525 738
rect 611 682 667 738
rect 753 682 809 738
rect 895 682 951 738
rect 1037 682 1093 738
rect 1179 682 1235 738
rect 1321 682 1377 738
rect 1463 682 1519 738
rect 1605 682 1661 738
rect 1747 682 1803 738
rect 1889 682 1945 738
rect 2031 682 2087 738
rect 2173 682 2229 738
rect 2315 682 2371 738
rect 2457 682 2513 738
rect 2599 682 2655 738
rect 2741 682 2797 738
rect 2883 682 2939 738
rect 3025 682 3081 738
rect 3167 682 3223 738
rect 3309 682 3365 738
rect 3451 682 3507 738
rect 3593 682 3649 738
rect 3735 682 3791 738
rect 3877 682 3933 738
rect 4019 682 4075 738
rect 4161 682 4217 738
rect 4303 682 4359 738
rect 4445 682 4501 738
rect 4587 682 4643 738
rect 4729 682 4785 738
rect 4871 682 4927 738
rect 5013 682 5069 738
rect 5155 682 5211 738
rect 5297 682 5353 738
rect 5439 682 5495 738
rect 5581 682 5637 738
rect 5723 682 5779 738
rect 5865 682 5921 738
rect 6007 682 6063 738
rect 6149 682 6205 738
rect 6291 682 6347 738
rect 6433 682 6489 738
rect 6575 682 6631 738
rect 6717 682 6773 738
rect 6859 682 6915 738
rect 7001 682 7057 738
rect 7143 682 7199 738
rect 7285 682 7341 738
rect -7341 540 -7285 596
rect -7199 540 -7143 596
rect -7057 540 -7001 596
rect -6915 540 -6859 596
rect -6773 540 -6717 596
rect -6631 540 -6575 596
rect -6489 540 -6433 596
rect -6347 540 -6291 596
rect -6205 540 -6149 596
rect -6063 540 -6007 596
rect -5921 540 -5865 596
rect -5779 540 -5723 596
rect -5637 540 -5581 596
rect -5495 540 -5439 596
rect -5353 540 -5297 596
rect -5211 540 -5155 596
rect -5069 540 -5013 596
rect -4927 540 -4871 596
rect -4785 540 -4729 596
rect -4643 540 -4587 596
rect -4501 540 -4445 596
rect -4359 540 -4303 596
rect -4217 540 -4161 596
rect -4075 540 -4019 596
rect -3933 540 -3877 596
rect -3791 540 -3735 596
rect -3649 540 -3593 596
rect -3507 540 -3451 596
rect -3365 540 -3309 596
rect -3223 540 -3167 596
rect -3081 540 -3025 596
rect -2939 540 -2883 596
rect -2797 540 -2741 596
rect -2655 540 -2599 596
rect -2513 540 -2457 596
rect -2371 540 -2315 596
rect -2229 540 -2173 596
rect -2087 540 -2031 596
rect -1945 540 -1889 596
rect -1803 540 -1747 596
rect -1661 540 -1605 596
rect -1519 540 -1463 596
rect -1377 540 -1321 596
rect -1235 540 -1179 596
rect -1093 540 -1037 596
rect -951 540 -895 596
rect -809 540 -753 596
rect -667 540 -611 596
rect -525 540 -469 596
rect -383 540 -327 596
rect -241 540 -185 596
rect -99 540 -43 596
rect 43 540 99 596
rect 185 540 241 596
rect 327 540 383 596
rect 469 540 525 596
rect 611 540 667 596
rect 753 540 809 596
rect 895 540 951 596
rect 1037 540 1093 596
rect 1179 540 1235 596
rect 1321 540 1377 596
rect 1463 540 1519 596
rect 1605 540 1661 596
rect 1747 540 1803 596
rect 1889 540 1945 596
rect 2031 540 2087 596
rect 2173 540 2229 596
rect 2315 540 2371 596
rect 2457 540 2513 596
rect 2599 540 2655 596
rect 2741 540 2797 596
rect 2883 540 2939 596
rect 3025 540 3081 596
rect 3167 540 3223 596
rect 3309 540 3365 596
rect 3451 540 3507 596
rect 3593 540 3649 596
rect 3735 540 3791 596
rect 3877 540 3933 596
rect 4019 540 4075 596
rect 4161 540 4217 596
rect 4303 540 4359 596
rect 4445 540 4501 596
rect 4587 540 4643 596
rect 4729 540 4785 596
rect 4871 540 4927 596
rect 5013 540 5069 596
rect 5155 540 5211 596
rect 5297 540 5353 596
rect 5439 540 5495 596
rect 5581 540 5637 596
rect 5723 540 5779 596
rect 5865 540 5921 596
rect 6007 540 6063 596
rect 6149 540 6205 596
rect 6291 540 6347 596
rect 6433 540 6489 596
rect 6575 540 6631 596
rect 6717 540 6773 596
rect 6859 540 6915 596
rect 7001 540 7057 596
rect 7143 540 7199 596
rect 7285 540 7341 596
rect -7341 398 -7285 454
rect -7199 398 -7143 454
rect -7057 398 -7001 454
rect -6915 398 -6859 454
rect -6773 398 -6717 454
rect -6631 398 -6575 454
rect -6489 398 -6433 454
rect -6347 398 -6291 454
rect -6205 398 -6149 454
rect -6063 398 -6007 454
rect -5921 398 -5865 454
rect -5779 398 -5723 454
rect -5637 398 -5581 454
rect -5495 398 -5439 454
rect -5353 398 -5297 454
rect -5211 398 -5155 454
rect -5069 398 -5013 454
rect -4927 398 -4871 454
rect -4785 398 -4729 454
rect -4643 398 -4587 454
rect -4501 398 -4445 454
rect -4359 398 -4303 454
rect -4217 398 -4161 454
rect -4075 398 -4019 454
rect -3933 398 -3877 454
rect -3791 398 -3735 454
rect -3649 398 -3593 454
rect -3507 398 -3451 454
rect -3365 398 -3309 454
rect -3223 398 -3167 454
rect -3081 398 -3025 454
rect -2939 398 -2883 454
rect -2797 398 -2741 454
rect -2655 398 -2599 454
rect -2513 398 -2457 454
rect -2371 398 -2315 454
rect -2229 398 -2173 454
rect -2087 398 -2031 454
rect -1945 398 -1889 454
rect -1803 398 -1747 454
rect -1661 398 -1605 454
rect -1519 398 -1463 454
rect -1377 398 -1321 454
rect -1235 398 -1179 454
rect -1093 398 -1037 454
rect -951 398 -895 454
rect -809 398 -753 454
rect -667 398 -611 454
rect -525 398 -469 454
rect -383 398 -327 454
rect -241 398 -185 454
rect -99 398 -43 454
rect 43 398 99 454
rect 185 398 241 454
rect 327 398 383 454
rect 469 398 525 454
rect 611 398 667 454
rect 753 398 809 454
rect 895 398 951 454
rect 1037 398 1093 454
rect 1179 398 1235 454
rect 1321 398 1377 454
rect 1463 398 1519 454
rect 1605 398 1661 454
rect 1747 398 1803 454
rect 1889 398 1945 454
rect 2031 398 2087 454
rect 2173 398 2229 454
rect 2315 398 2371 454
rect 2457 398 2513 454
rect 2599 398 2655 454
rect 2741 398 2797 454
rect 2883 398 2939 454
rect 3025 398 3081 454
rect 3167 398 3223 454
rect 3309 398 3365 454
rect 3451 398 3507 454
rect 3593 398 3649 454
rect 3735 398 3791 454
rect 3877 398 3933 454
rect 4019 398 4075 454
rect 4161 398 4217 454
rect 4303 398 4359 454
rect 4445 398 4501 454
rect 4587 398 4643 454
rect 4729 398 4785 454
rect 4871 398 4927 454
rect 5013 398 5069 454
rect 5155 398 5211 454
rect 5297 398 5353 454
rect 5439 398 5495 454
rect 5581 398 5637 454
rect 5723 398 5779 454
rect 5865 398 5921 454
rect 6007 398 6063 454
rect 6149 398 6205 454
rect 6291 398 6347 454
rect 6433 398 6489 454
rect 6575 398 6631 454
rect 6717 398 6773 454
rect 6859 398 6915 454
rect 7001 398 7057 454
rect 7143 398 7199 454
rect 7285 398 7341 454
rect -7341 256 -7285 312
rect -7199 256 -7143 312
rect -7057 256 -7001 312
rect -6915 256 -6859 312
rect -6773 256 -6717 312
rect -6631 256 -6575 312
rect -6489 256 -6433 312
rect -6347 256 -6291 312
rect -6205 256 -6149 312
rect -6063 256 -6007 312
rect -5921 256 -5865 312
rect -5779 256 -5723 312
rect -5637 256 -5581 312
rect -5495 256 -5439 312
rect -5353 256 -5297 312
rect -5211 256 -5155 312
rect -5069 256 -5013 312
rect -4927 256 -4871 312
rect -4785 256 -4729 312
rect -4643 256 -4587 312
rect -4501 256 -4445 312
rect -4359 256 -4303 312
rect -4217 256 -4161 312
rect -4075 256 -4019 312
rect -3933 256 -3877 312
rect -3791 256 -3735 312
rect -3649 256 -3593 312
rect -3507 256 -3451 312
rect -3365 256 -3309 312
rect -3223 256 -3167 312
rect -3081 256 -3025 312
rect -2939 256 -2883 312
rect -2797 256 -2741 312
rect -2655 256 -2599 312
rect -2513 256 -2457 312
rect -2371 256 -2315 312
rect -2229 256 -2173 312
rect -2087 256 -2031 312
rect -1945 256 -1889 312
rect -1803 256 -1747 312
rect -1661 256 -1605 312
rect -1519 256 -1463 312
rect -1377 256 -1321 312
rect -1235 256 -1179 312
rect -1093 256 -1037 312
rect -951 256 -895 312
rect -809 256 -753 312
rect -667 256 -611 312
rect -525 256 -469 312
rect -383 256 -327 312
rect -241 256 -185 312
rect -99 256 -43 312
rect 43 256 99 312
rect 185 256 241 312
rect 327 256 383 312
rect 469 256 525 312
rect 611 256 667 312
rect 753 256 809 312
rect 895 256 951 312
rect 1037 256 1093 312
rect 1179 256 1235 312
rect 1321 256 1377 312
rect 1463 256 1519 312
rect 1605 256 1661 312
rect 1747 256 1803 312
rect 1889 256 1945 312
rect 2031 256 2087 312
rect 2173 256 2229 312
rect 2315 256 2371 312
rect 2457 256 2513 312
rect 2599 256 2655 312
rect 2741 256 2797 312
rect 2883 256 2939 312
rect 3025 256 3081 312
rect 3167 256 3223 312
rect 3309 256 3365 312
rect 3451 256 3507 312
rect 3593 256 3649 312
rect 3735 256 3791 312
rect 3877 256 3933 312
rect 4019 256 4075 312
rect 4161 256 4217 312
rect 4303 256 4359 312
rect 4445 256 4501 312
rect 4587 256 4643 312
rect 4729 256 4785 312
rect 4871 256 4927 312
rect 5013 256 5069 312
rect 5155 256 5211 312
rect 5297 256 5353 312
rect 5439 256 5495 312
rect 5581 256 5637 312
rect 5723 256 5779 312
rect 5865 256 5921 312
rect 6007 256 6063 312
rect 6149 256 6205 312
rect 6291 256 6347 312
rect 6433 256 6489 312
rect 6575 256 6631 312
rect 6717 256 6773 312
rect 6859 256 6915 312
rect 7001 256 7057 312
rect 7143 256 7199 312
rect 7285 256 7341 312
rect -7341 114 -7285 170
rect -7199 114 -7143 170
rect -7057 114 -7001 170
rect -6915 114 -6859 170
rect -6773 114 -6717 170
rect -6631 114 -6575 170
rect -6489 114 -6433 170
rect -6347 114 -6291 170
rect -6205 114 -6149 170
rect -6063 114 -6007 170
rect -5921 114 -5865 170
rect -5779 114 -5723 170
rect -5637 114 -5581 170
rect -5495 114 -5439 170
rect -5353 114 -5297 170
rect -5211 114 -5155 170
rect -5069 114 -5013 170
rect -4927 114 -4871 170
rect -4785 114 -4729 170
rect -4643 114 -4587 170
rect -4501 114 -4445 170
rect -4359 114 -4303 170
rect -4217 114 -4161 170
rect -4075 114 -4019 170
rect -3933 114 -3877 170
rect -3791 114 -3735 170
rect -3649 114 -3593 170
rect -3507 114 -3451 170
rect -3365 114 -3309 170
rect -3223 114 -3167 170
rect -3081 114 -3025 170
rect -2939 114 -2883 170
rect -2797 114 -2741 170
rect -2655 114 -2599 170
rect -2513 114 -2457 170
rect -2371 114 -2315 170
rect -2229 114 -2173 170
rect -2087 114 -2031 170
rect -1945 114 -1889 170
rect -1803 114 -1747 170
rect -1661 114 -1605 170
rect -1519 114 -1463 170
rect -1377 114 -1321 170
rect -1235 114 -1179 170
rect -1093 114 -1037 170
rect -951 114 -895 170
rect -809 114 -753 170
rect -667 114 -611 170
rect -525 114 -469 170
rect -383 114 -327 170
rect -241 114 -185 170
rect -99 114 -43 170
rect 43 114 99 170
rect 185 114 241 170
rect 327 114 383 170
rect 469 114 525 170
rect 611 114 667 170
rect 753 114 809 170
rect 895 114 951 170
rect 1037 114 1093 170
rect 1179 114 1235 170
rect 1321 114 1377 170
rect 1463 114 1519 170
rect 1605 114 1661 170
rect 1747 114 1803 170
rect 1889 114 1945 170
rect 2031 114 2087 170
rect 2173 114 2229 170
rect 2315 114 2371 170
rect 2457 114 2513 170
rect 2599 114 2655 170
rect 2741 114 2797 170
rect 2883 114 2939 170
rect 3025 114 3081 170
rect 3167 114 3223 170
rect 3309 114 3365 170
rect 3451 114 3507 170
rect 3593 114 3649 170
rect 3735 114 3791 170
rect 3877 114 3933 170
rect 4019 114 4075 170
rect 4161 114 4217 170
rect 4303 114 4359 170
rect 4445 114 4501 170
rect 4587 114 4643 170
rect 4729 114 4785 170
rect 4871 114 4927 170
rect 5013 114 5069 170
rect 5155 114 5211 170
rect 5297 114 5353 170
rect 5439 114 5495 170
rect 5581 114 5637 170
rect 5723 114 5779 170
rect 5865 114 5921 170
rect 6007 114 6063 170
rect 6149 114 6205 170
rect 6291 114 6347 170
rect 6433 114 6489 170
rect 6575 114 6631 170
rect 6717 114 6773 170
rect 6859 114 6915 170
rect 7001 114 7057 170
rect 7143 114 7199 170
rect 7285 114 7341 170
rect -7341 -28 -7285 28
rect -7199 -28 -7143 28
rect -7057 -28 -7001 28
rect -6915 -28 -6859 28
rect -6773 -28 -6717 28
rect -6631 -28 -6575 28
rect -6489 -28 -6433 28
rect -6347 -28 -6291 28
rect -6205 -28 -6149 28
rect -6063 -28 -6007 28
rect -5921 -28 -5865 28
rect -5779 -28 -5723 28
rect -5637 -28 -5581 28
rect -5495 -28 -5439 28
rect -5353 -28 -5297 28
rect -5211 -28 -5155 28
rect -5069 -28 -5013 28
rect -4927 -28 -4871 28
rect -4785 -28 -4729 28
rect -4643 -28 -4587 28
rect -4501 -28 -4445 28
rect -4359 -28 -4303 28
rect -4217 -28 -4161 28
rect -4075 -28 -4019 28
rect -3933 -28 -3877 28
rect -3791 -28 -3735 28
rect -3649 -28 -3593 28
rect -3507 -28 -3451 28
rect -3365 -28 -3309 28
rect -3223 -28 -3167 28
rect -3081 -28 -3025 28
rect -2939 -28 -2883 28
rect -2797 -28 -2741 28
rect -2655 -28 -2599 28
rect -2513 -28 -2457 28
rect -2371 -28 -2315 28
rect -2229 -28 -2173 28
rect -2087 -28 -2031 28
rect -1945 -28 -1889 28
rect -1803 -28 -1747 28
rect -1661 -28 -1605 28
rect -1519 -28 -1463 28
rect -1377 -28 -1321 28
rect -1235 -28 -1179 28
rect -1093 -28 -1037 28
rect -951 -28 -895 28
rect -809 -28 -753 28
rect -667 -28 -611 28
rect -525 -28 -469 28
rect -383 -28 -327 28
rect -241 -28 -185 28
rect -99 -28 -43 28
rect 43 -28 99 28
rect 185 -28 241 28
rect 327 -28 383 28
rect 469 -28 525 28
rect 611 -28 667 28
rect 753 -28 809 28
rect 895 -28 951 28
rect 1037 -28 1093 28
rect 1179 -28 1235 28
rect 1321 -28 1377 28
rect 1463 -28 1519 28
rect 1605 -28 1661 28
rect 1747 -28 1803 28
rect 1889 -28 1945 28
rect 2031 -28 2087 28
rect 2173 -28 2229 28
rect 2315 -28 2371 28
rect 2457 -28 2513 28
rect 2599 -28 2655 28
rect 2741 -28 2797 28
rect 2883 -28 2939 28
rect 3025 -28 3081 28
rect 3167 -28 3223 28
rect 3309 -28 3365 28
rect 3451 -28 3507 28
rect 3593 -28 3649 28
rect 3735 -28 3791 28
rect 3877 -28 3933 28
rect 4019 -28 4075 28
rect 4161 -28 4217 28
rect 4303 -28 4359 28
rect 4445 -28 4501 28
rect 4587 -28 4643 28
rect 4729 -28 4785 28
rect 4871 -28 4927 28
rect 5013 -28 5069 28
rect 5155 -28 5211 28
rect 5297 -28 5353 28
rect 5439 -28 5495 28
rect 5581 -28 5637 28
rect 5723 -28 5779 28
rect 5865 -28 5921 28
rect 6007 -28 6063 28
rect 6149 -28 6205 28
rect 6291 -28 6347 28
rect 6433 -28 6489 28
rect 6575 -28 6631 28
rect 6717 -28 6773 28
rect 6859 -28 6915 28
rect 7001 -28 7057 28
rect 7143 -28 7199 28
rect 7285 -28 7341 28
rect -7341 -170 -7285 -114
rect -7199 -170 -7143 -114
rect -7057 -170 -7001 -114
rect -6915 -170 -6859 -114
rect -6773 -170 -6717 -114
rect -6631 -170 -6575 -114
rect -6489 -170 -6433 -114
rect -6347 -170 -6291 -114
rect -6205 -170 -6149 -114
rect -6063 -170 -6007 -114
rect -5921 -170 -5865 -114
rect -5779 -170 -5723 -114
rect -5637 -170 -5581 -114
rect -5495 -170 -5439 -114
rect -5353 -170 -5297 -114
rect -5211 -170 -5155 -114
rect -5069 -170 -5013 -114
rect -4927 -170 -4871 -114
rect -4785 -170 -4729 -114
rect -4643 -170 -4587 -114
rect -4501 -170 -4445 -114
rect -4359 -170 -4303 -114
rect -4217 -170 -4161 -114
rect -4075 -170 -4019 -114
rect -3933 -170 -3877 -114
rect -3791 -170 -3735 -114
rect -3649 -170 -3593 -114
rect -3507 -170 -3451 -114
rect -3365 -170 -3309 -114
rect -3223 -170 -3167 -114
rect -3081 -170 -3025 -114
rect -2939 -170 -2883 -114
rect -2797 -170 -2741 -114
rect -2655 -170 -2599 -114
rect -2513 -170 -2457 -114
rect -2371 -170 -2315 -114
rect -2229 -170 -2173 -114
rect -2087 -170 -2031 -114
rect -1945 -170 -1889 -114
rect -1803 -170 -1747 -114
rect -1661 -170 -1605 -114
rect -1519 -170 -1463 -114
rect -1377 -170 -1321 -114
rect -1235 -170 -1179 -114
rect -1093 -170 -1037 -114
rect -951 -170 -895 -114
rect -809 -170 -753 -114
rect -667 -170 -611 -114
rect -525 -170 -469 -114
rect -383 -170 -327 -114
rect -241 -170 -185 -114
rect -99 -170 -43 -114
rect 43 -170 99 -114
rect 185 -170 241 -114
rect 327 -170 383 -114
rect 469 -170 525 -114
rect 611 -170 667 -114
rect 753 -170 809 -114
rect 895 -170 951 -114
rect 1037 -170 1093 -114
rect 1179 -170 1235 -114
rect 1321 -170 1377 -114
rect 1463 -170 1519 -114
rect 1605 -170 1661 -114
rect 1747 -170 1803 -114
rect 1889 -170 1945 -114
rect 2031 -170 2087 -114
rect 2173 -170 2229 -114
rect 2315 -170 2371 -114
rect 2457 -170 2513 -114
rect 2599 -170 2655 -114
rect 2741 -170 2797 -114
rect 2883 -170 2939 -114
rect 3025 -170 3081 -114
rect 3167 -170 3223 -114
rect 3309 -170 3365 -114
rect 3451 -170 3507 -114
rect 3593 -170 3649 -114
rect 3735 -170 3791 -114
rect 3877 -170 3933 -114
rect 4019 -170 4075 -114
rect 4161 -170 4217 -114
rect 4303 -170 4359 -114
rect 4445 -170 4501 -114
rect 4587 -170 4643 -114
rect 4729 -170 4785 -114
rect 4871 -170 4927 -114
rect 5013 -170 5069 -114
rect 5155 -170 5211 -114
rect 5297 -170 5353 -114
rect 5439 -170 5495 -114
rect 5581 -170 5637 -114
rect 5723 -170 5779 -114
rect 5865 -170 5921 -114
rect 6007 -170 6063 -114
rect 6149 -170 6205 -114
rect 6291 -170 6347 -114
rect 6433 -170 6489 -114
rect 6575 -170 6631 -114
rect 6717 -170 6773 -114
rect 6859 -170 6915 -114
rect 7001 -170 7057 -114
rect 7143 -170 7199 -114
rect 7285 -170 7341 -114
rect -7341 -312 -7285 -256
rect -7199 -312 -7143 -256
rect -7057 -312 -7001 -256
rect -6915 -312 -6859 -256
rect -6773 -312 -6717 -256
rect -6631 -312 -6575 -256
rect -6489 -312 -6433 -256
rect -6347 -312 -6291 -256
rect -6205 -312 -6149 -256
rect -6063 -312 -6007 -256
rect -5921 -312 -5865 -256
rect -5779 -312 -5723 -256
rect -5637 -312 -5581 -256
rect -5495 -312 -5439 -256
rect -5353 -312 -5297 -256
rect -5211 -312 -5155 -256
rect -5069 -312 -5013 -256
rect -4927 -312 -4871 -256
rect -4785 -312 -4729 -256
rect -4643 -312 -4587 -256
rect -4501 -312 -4445 -256
rect -4359 -312 -4303 -256
rect -4217 -312 -4161 -256
rect -4075 -312 -4019 -256
rect -3933 -312 -3877 -256
rect -3791 -312 -3735 -256
rect -3649 -312 -3593 -256
rect -3507 -312 -3451 -256
rect -3365 -312 -3309 -256
rect -3223 -312 -3167 -256
rect -3081 -312 -3025 -256
rect -2939 -312 -2883 -256
rect -2797 -312 -2741 -256
rect -2655 -312 -2599 -256
rect -2513 -312 -2457 -256
rect -2371 -312 -2315 -256
rect -2229 -312 -2173 -256
rect -2087 -312 -2031 -256
rect -1945 -312 -1889 -256
rect -1803 -312 -1747 -256
rect -1661 -312 -1605 -256
rect -1519 -312 -1463 -256
rect -1377 -312 -1321 -256
rect -1235 -312 -1179 -256
rect -1093 -312 -1037 -256
rect -951 -312 -895 -256
rect -809 -312 -753 -256
rect -667 -312 -611 -256
rect -525 -312 -469 -256
rect -383 -312 -327 -256
rect -241 -312 -185 -256
rect -99 -312 -43 -256
rect 43 -312 99 -256
rect 185 -312 241 -256
rect 327 -312 383 -256
rect 469 -312 525 -256
rect 611 -312 667 -256
rect 753 -312 809 -256
rect 895 -312 951 -256
rect 1037 -312 1093 -256
rect 1179 -312 1235 -256
rect 1321 -312 1377 -256
rect 1463 -312 1519 -256
rect 1605 -312 1661 -256
rect 1747 -312 1803 -256
rect 1889 -312 1945 -256
rect 2031 -312 2087 -256
rect 2173 -312 2229 -256
rect 2315 -312 2371 -256
rect 2457 -312 2513 -256
rect 2599 -312 2655 -256
rect 2741 -312 2797 -256
rect 2883 -312 2939 -256
rect 3025 -312 3081 -256
rect 3167 -312 3223 -256
rect 3309 -312 3365 -256
rect 3451 -312 3507 -256
rect 3593 -312 3649 -256
rect 3735 -312 3791 -256
rect 3877 -312 3933 -256
rect 4019 -312 4075 -256
rect 4161 -312 4217 -256
rect 4303 -312 4359 -256
rect 4445 -312 4501 -256
rect 4587 -312 4643 -256
rect 4729 -312 4785 -256
rect 4871 -312 4927 -256
rect 5013 -312 5069 -256
rect 5155 -312 5211 -256
rect 5297 -312 5353 -256
rect 5439 -312 5495 -256
rect 5581 -312 5637 -256
rect 5723 -312 5779 -256
rect 5865 -312 5921 -256
rect 6007 -312 6063 -256
rect 6149 -312 6205 -256
rect 6291 -312 6347 -256
rect 6433 -312 6489 -256
rect 6575 -312 6631 -256
rect 6717 -312 6773 -256
rect 6859 -312 6915 -256
rect 7001 -312 7057 -256
rect 7143 -312 7199 -256
rect 7285 -312 7341 -256
rect -7341 -454 -7285 -398
rect -7199 -454 -7143 -398
rect -7057 -454 -7001 -398
rect -6915 -454 -6859 -398
rect -6773 -454 -6717 -398
rect -6631 -454 -6575 -398
rect -6489 -454 -6433 -398
rect -6347 -454 -6291 -398
rect -6205 -454 -6149 -398
rect -6063 -454 -6007 -398
rect -5921 -454 -5865 -398
rect -5779 -454 -5723 -398
rect -5637 -454 -5581 -398
rect -5495 -454 -5439 -398
rect -5353 -454 -5297 -398
rect -5211 -454 -5155 -398
rect -5069 -454 -5013 -398
rect -4927 -454 -4871 -398
rect -4785 -454 -4729 -398
rect -4643 -454 -4587 -398
rect -4501 -454 -4445 -398
rect -4359 -454 -4303 -398
rect -4217 -454 -4161 -398
rect -4075 -454 -4019 -398
rect -3933 -454 -3877 -398
rect -3791 -454 -3735 -398
rect -3649 -454 -3593 -398
rect -3507 -454 -3451 -398
rect -3365 -454 -3309 -398
rect -3223 -454 -3167 -398
rect -3081 -454 -3025 -398
rect -2939 -454 -2883 -398
rect -2797 -454 -2741 -398
rect -2655 -454 -2599 -398
rect -2513 -454 -2457 -398
rect -2371 -454 -2315 -398
rect -2229 -454 -2173 -398
rect -2087 -454 -2031 -398
rect -1945 -454 -1889 -398
rect -1803 -454 -1747 -398
rect -1661 -454 -1605 -398
rect -1519 -454 -1463 -398
rect -1377 -454 -1321 -398
rect -1235 -454 -1179 -398
rect -1093 -454 -1037 -398
rect -951 -454 -895 -398
rect -809 -454 -753 -398
rect -667 -454 -611 -398
rect -525 -454 -469 -398
rect -383 -454 -327 -398
rect -241 -454 -185 -398
rect -99 -454 -43 -398
rect 43 -454 99 -398
rect 185 -454 241 -398
rect 327 -454 383 -398
rect 469 -454 525 -398
rect 611 -454 667 -398
rect 753 -454 809 -398
rect 895 -454 951 -398
rect 1037 -454 1093 -398
rect 1179 -454 1235 -398
rect 1321 -454 1377 -398
rect 1463 -454 1519 -398
rect 1605 -454 1661 -398
rect 1747 -454 1803 -398
rect 1889 -454 1945 -398
rect 2031 -454 2087 -398
rect 2173 -454 2229 -398
rect 2315 -454 2371 -398
rect 2457 -454 2513 -398
rect 2599 -454 2655 -398
rect 2741 -454 2797 -398
rect 2883 -454 2939 -398
rect 3025 -454 3081 -398
rect 3167 -454 3223 -398
rect 3309 -454 3365 -398
rect 3451 -454 3507 -398
rect 3593 -454 3649 -398
rect 3735 -454 3791 -398
rect 3877 -454 3933 -398
rect 4019 -454 4075 -398
rect 4161 -454 4217 -398
rect 4303 -454 4359 -398
rect 4445 -454 4501 -398
rect 4587 -454 4643 -398
rect 4729 -454 4785 -398
rect 4871 -454 4927 -398
rect 5013 -454 5069 -398
rect 5155 -454 5211 -398
rect 5297 -454 5353 -398
rect 5439 -454 5495 -398
rect 5581 -454 5637 -398
rect 5723 -454 5779 -398
rect 5865 -454 5921 -398
rect 6007 -454 6063 -398
rect 6149 -454 6205 -398
rect 6291 -454 6347 -398
rect 6433 -454 6489 -398
rect 6575 -454 6631 -398
rect 6717 -454 6773 -398
rect 6859 -454 6915 -398
rect 7001 -454 7057 -398
rect 7143 -454 7199 -398
rect 7285 -454 7341 -398
rect -7341 -596 -7285 -540
rect -7199 -596 -7143 -540
rect -7057 -596 -7001 -540
rect -6915 -596 -6859 -540
rect -6773 -596 -6717 -540
rect -6631 -596 -6575 -540
rect -6489 -596 -6433 -540
rect -6347 -596 -6291 -540
rect -6205 -596 -6149 -540
rect -6063 -596 -6007 -540
rect -5921 -596 -5865 -540
rect -5779 -596 -5723 -540
rect -5637 -596 -5581 -540
rect -5495 -596 -5439 -540
rect -5353 -596 -5297 -540
rect -5211 -596 -5155 -540
rect -5069 -596 -5013 -540
rect -4927 -596 -4871 -540
rect -4785 -596 -4729 -540
rect -4643 -596 -4587 -540
rect -4501 -596 -4445 -540
rect -4359 -596 -4303 -540
rect -4217 -596 -4161 -540
rect -4075 -596 -4019 -540
rect -3933 -596 -3877 -540
rect -3791 -596 -3735 -540
rect -3649 -596 -3593 -540
rect -3507 -596 -3451 -540
rect -3365 -596 -3309 -540
rect -3223 -596 -3167 -540
rect -3081 -596 -3025 -540
rect -2939 -596 -2883 -540
rect -2797 -596 -2741 -540
rect -2655 -596 -2599 -540
rect -2513 -596 -2457 -540
rect -2371 -596 -2315 -540
rect -2229 -596 -2173 -540
rect -2087 -596 -2031 -540
rect -1945 -596 -1889 -540
rect -1803 -596 -1747 -540
rect -1661 -596 -1605 -540
rect -1519 -596 -1463 -540
rect -1377 -596 -1321 -540
rect -1235 -596 -1179 -540
rect -1093 -596 -1037 -540
rect -951 -596 -895 -540
rect -809 -596 -753 -540
rect -667 -596 -611 -540
rect -525 -596 -469 -540
rect -383 -596 -327 -540
rect -241 -596 -185 -540
rect -99 -596 -43 -540
rect 43 -596 99 -540
rect 185 -596 241 -540
rect 327 -596 383 -540
rect 469 -596 525 -540
rect 611 -596 667 -540
rect 753 -596 809 -540
rect 895 -596 951 -540
rect 1037 -596 1093 -540
rect 1179 -596 1235 -540
rect 1321 -596 1377 -540
rect 1463 -596 1519 -540
rect 1605 -596 1661 -540
rect 1747 -596 1803 -540
rect 1889 -596 1945 -540
rect 2031 -596 2087 -540
rect 2173 -596 2229 -540
rect 2315 -596 2371 -540
rect 2457 -596 2513 -540
rect 2599 -596 2655 -540
rect 2741 -596 2797 -540
rect 2883 -596 2939 -540
rect 3025 -596 3081 -540
rect 3167 -596 3223 -540
rect 3309 -596 3365 -540
rect 3451 -596 3507 -540
rect 3593 -596 3649 -540
rect 3735 -596 3791 -540
rect 3877 -596 3933 -540
rect 4019 -596 4075 -540
rect 4161 -596 4217 -540
rect 4303 -596 4359 -540
rect 4445 -596 4501 -540
rect 4587 -596 4643 -540
rect 4729 -596 4785 -540
rect 4871 -596 4927 -540
rect 5013 -596 5069 -540
rect 5155 -596 5211 -540
rect 5297 -596 5353 -540
rect 5439 -596 5495 -540
rect 5581 -596 5637 -540
rect 5723 -596 5779 -540
rect 5865 -596 5921 -540
rect 6007 -596 6063 -540
rect 6149 -596 6205 -540
rect 6291 -596 6347 -540
rect 6433 -596 6489 -540
rect 6575 -596 6631 -540
rect 6717 -596 6773 -540
rect 6859 -596 6915 -540
rect 7001 -596 7057 -540
rect 7143 -596 7199 -540
rect 7285 -596 7341 -540
rect -7341 -738 -7285 -682
rect -7199 -738 -7143 -682
rect -7057 -738 -7001 -682
rect -6915 -738 -6859 -682
rect -6773 -738 -6717 -682
rect -6631 -738 -6575 -682
rect -6489 -738 -6433 -682
rect -6347 -738 -6291 -682
rect -6205 -738 -6149 -682
rect -6063 -738 -6007 -682
rect -5921 -738 -5865 -682
rect -5779 -738 -5723 -682
rect -5637 -738 -5581 -682
rect -5495 -738 -5439 -682
rect -5353 -738 -5297 -682
rect -5211 -738 -5155 -682
rect -5069 -738 -5013 -682
rect -4927 -738 -4871 -682
rect -4785 -738 -4729 -682
rect -4643 -738 -4587 -682
rect -4501 -738 -4445 -682
rect -4359 -738 -4303 -682
rect -4217 -738 -4161 -682
rect -4075 -738 -4019 -682
rect -3933 -738 -3877 -682
rect -3791 -738 -3735 -682
rect -3649 -738 -3593 -682
rect -3507 -738 -3451 -682
rect -3365 -738 -3309 -682
rect -3223 -738 -3167 -682
rect -3081 -738 -3025 -682
rect -2939 -738 -2883 -682
rect -2797 -738 -2741 -682
rect -2655 -738 -2599 -682
rect -2513 -738 -2457 -682
rect -2371 -738 -2315 -682
rect -2229 -738 -2173 -682
rect -2087 -738 -2031 -682
rect -1945 -738 -1889 -682
rect -1803 -738 -1747 -682
rect -1661 -738 -1605 -682
rect -1519 -738 -1463 -682
rect -1377 -738 -1321 -682
rect -1235 -738 -1179 -682
rect -1093 -738 -1037 -682
rect -951 -738 -895 -682
rect -809 -738 -753 -682
rect -667 -738 -611 -682
rect -525 -738 -469 -682
rect -383 -738 -327 -682
rect -241 -738 -185 -682
rect -99 -738 -43 -682
rect 43 -738 99 -682
rect 185 -738 241 -682
rect 327 -738 383 -682
rect 469 -738 525 -682
rect 611 -738 667 -682
rect 753 -738 809 -682
rect 895 -738 951 -682
rect 1037 -738 1093 -682
rect 1179 -738 1235 -682
rect 1321 -738 1377 -682
rect 1463 -738 1519 -682
rect 1605 -738 1661 -682
rect 1747 -738 1803 -682
rect 1889 -738 1945 -682
rect 2031 -738 2087 -682
rect 2173 -738 2229 -682
rect 2315 -738 2371 -682
rect 2457 -738 2513 -682
rect 2599 -738 2655 -682
rect 2741 -738 2797 -682
rect 2883 -738 2939 -682
rect 3025 -738 3081 -682
rect 3167 -738 3223 -682
rect 3309 -738 3365 -682
rect 3451 -738 3507 -682
rect 3593 -738 3649 -682
rect 3735 -738 3791 -682
rect 3877 -738 3933 -682
rect 4019 -738 4075 -682
rect 4161 -738 4217 -682
rect 4303 -738 4359 -682
rect 4445 -738 4501 -682
rect 4587 -738 4643 -682
rect 4729 -738 4785 -682
rect 4871 -738 4927 -682
rect 5013 -738 5069 -682
rect 5155 -738 5211 -682
rect 5297 -738 5353 -682
rect 5439 -738 5495 -682
rect 5581 -738 5637 -682
rect 5723 -738 5779 -682
rect 5865 -738 5921 -682
rect 6007 -738 6063 -682
rect 6149 -738 6205 -682
rect 6291 -738 6347 -682
rect 6433 -738 6489 -682
rect 6575 -738 6631 -682
rect 6717 -738 6773 -682
rect 6859 -738 6915 -682
rect 7001 -738 7057 -682
rect 7143 -738 7199 -682
rect 7285 -738 7341 -682
rect -7341 -880 -7285 -824
rect -7199 -880 -7143 -824
rect -7057 -880 -7001 -824
rect -6915 -880 -6859 -824
rect -6773 -880 -6717 -824
rect -6631 -880 -6575 -824
rect -6489 -880 -6433 -824
rect -6347 -880 -6291 -824
rect -6205 -880 -6149 -824
rect -6063 -880 -6007 -824
rect -5921 -880 -5865 -824
rect -5779 -880 -5723 -824
rect -5637 -880 -5581 -824
rect -5495 -880 -5439 -824
rect -5353 -880 -5297 -824
rect -5211 -880 -5155 -824
rect -5069 -880 -5013 -824
rect -4927 -880 -4871 -824
rect -4785 -880 -4729 -824
rect -4643 -880 -4587 -824
rect -4501 -880 -4445 -824
rect -4359 -880 -4303 -824
rect -4217 -880 -4161 -824
rect -4075 -880 -4019 -824
rect -3933 -880 -3877 -824
rect -3791 -880 -3735 -824
rect -3649 -880 -3593 -824
rect -3507 -880 -3451 -824
rect -3365 -880 -3309 -824
rect -3223 -880 -3167 -824
rect -3081 -880 -3025 -824
rect -2939 -880 -2883 -824
rect -2797 -880 -2741 -824
rect -2655 -880 -2599 -824
rect -2513 -880 -2457 -824
rect -2371 -880 -2315 -824
rect -2229 -880 -2173 -824
rect -2087 -880 -2031 -824
rect -1945 -880 -1889 -824
rect -1803 -880 -1747 -824
rect -1661 -880 -1605 -824
rect -1519 -880 -1463 -824
rect -1377 -880 -1321 -824
rect -1235 -880 -1179 -824
rect -1093 -880 -1037 -824
rect -951 -880 -895 -824
rect -809 -880 -753 -824
rect -667 -880 -611 -824
rect -525 -880 -469 -824
rect -383 -880 -327 -824
rect -241 -880 -185 -824
rect -99 -880 -43 -824
rect 43 -880 99 -824
rect 185 -880 241 -824
rect 327 -880 383 -824
rect 469 -880 525 -824
rect 611 -880 667 -824
rect 753 -880 809 -824
rect 895 -880 951 -824
rect 1037 -880 1093 -824
rect 1179 -880 1235 -824
rect 1321 -880 1377 -824
rect 1463 -880 1519 -824
rect 1605 -880 1661 -824
rect 1747 -880 1803 -824
rect 1889 -880 1945 -824
rect 2031 -880 2087 -824
rect 2173 -880 2229 -824
rect 2315 -880 2371 -824
rect 2457 -880 2513 -824
rect 2599 -880 2655 -824
rect 2741 -880 2797 -824
rect 2883 -880 2939 -824
rect 3025 -880 3081 -824
rect 3167 -880 3223 -824
rect 3309 -880 3365 -824
rect 3451 -880 3507 -824
rect 3593 -880 3649 -824
rect 3735 -880 3791 -824
rect 3877 -880 3933 -824
rect 4019 -880 4075 -824
rect 4161 -880 4217 -824
rect 4303 -880 4359 -824
rect 4445 -880 4501 -824
rect 4587 -880 4643 -824
rect 4729 -880 4785 -824
rect 4871 -880 4927 -824
rect 5013 -880 5069 -824
rect 5155 -880 5211 -824
rect 5297 -880 5353 -824
rect 5439 -880 5495 -824
rect 5581 -880 5637 -824
rect 5723 -880 5779 -824
rect 5865 -880 5921 -824
rect 6007 -880 6063 -824
rect 6149 -880 6205 -824
rect 6291 -880 6347 -824
rect 6433 -880 6489 -824
rect 6575 -880 6631 -824
rect 6717 -880 6773 -824
rect 6859 -880 6915 -824
rect 7001 -880 7057 -824
rect 7143 -880 7199 -824
rect 7285 -880 7341 -824
rect -7341 -1022 -7285 -966
rect -7199 -1022 -7143 -966
rect -7057 -1022 -7001 -966
rect -6915 -1022 -6859 -966
rect -6773 -1022 -6717 -966
rect -6631 -1022 -6575 -966
rect -6489 -1022 -6433 -966
rect -6347 -1022 -6291 -966
rect -6205 -1022 -6149 -966
rect -6063 -1022 -6007 -966
rect -5921 -1022 -5865 -966
rect -5779 -1022 -5723 -966
rect -5637 -1022 -5581 -966
rect -5495 -1022 -5439 -966
rect -5353 -1022 -5297 -966
rect -5211 -1022 -5155 -966
rect -5069 -1022 -5013 -966
rect -4927 -1022 -4871 -966
rect -4785 -1022 -4729 -966
rect -4643 -1022 -4587 -966
rect -4501 -1022 -4445 -966
rect -4359 -1022 -4303 -966
rect -4217 -1022 -4161 -966
rect -4075 -1022 -4019 -966
rect -3933 -1022 -3877 -966
rect -3791 -1022 -3735 -966
rect -3649 -1022 -3593 -966
rect -3507 -1022 -3451 -966
rect -3365 -1022 -3309 -966
rect -3223 -1022 -3167 -966
rect -3081 -1022 -3025 -966
rect -2939 -1022 -2883 -966
rect -2797 -1022 -2741 -966
rect -2655 -1022 -2599 -966
rect -2513 -1022 -2457 -966
rect -2371 -1022 -2315 -966
rect -2229 -1022 -2173 -966
rect -2087 -1022 -2031 -966
rect -1945 -1022 -1889 -966
rect -1803 -1022 -1747 -966
rect -1661 -1022 -1605 -966
rect -1519 -1022 -1463 -966
rect -1377 -1022 -1321 -966
rect -1235 -1022 -1179 -966
rect -1093 -1022 -1037 -966
rect -951 -1022 -895 -966
rect -809 -1022 -753 -966
rect -667 -1022 -611 -966
rect -525 -1022 -469 -966
rect -383 -1022 -327 -966
rect -241 -1022 -185 -966
rect -99 -1022 -43 -966
rect 43 -1022 99 -966
rect 185 -1022 241 -966
rect 327 -1022 383 -966
rect 469 -1022 525 -966
rect 611 -1022 667 -966
rect 753 -1022 809 -966
rect 895 -1022 951 -966
rect 1037 -1022 1093 -966
rect 1179 -1022 1235 -966
rect 1321 -1022 1377 -966
rect 1463 -1022 1519 -966
rect 1605 -1022 1661 -966
rect 1747 -1022 1803 -966
rect 1889 -1022 1945 -966
rect 2031 -1022 2087 -966
rect 2173 -1022 2229 -966
rect 2315 -1022 2371 -966
rect 2457 -1022 2513 -966
rect 2599 -1022 2655 -966
rect 2741 -1022 2797 -966
rect 2883 -1022 2939 -966
rect 3025 -1022 3081 -966
rect 3167 -1022 3223 -966
rect 3309 -1022 3365 -966
rect 3451 -1022 3507 -966
rect 3593 -1022 3649 -966
rect 3735 -1022 3791 -966
rect 3877 -1022 3933 -966
rect 4019 -1022 4075 -966
rect 4161 -1022 4217 -966
rect 4303 -1022 4359 -966
rect 4445 -1022 4501 -966
rect 4587 -1022 4643 -966
rect 4729 -1022 4785 -966
rect 4871 -1022 4927 -966
rect 5013 -1022 5069 -966
rect 5155 -1022 5211 -966
rect 5297 -1022 5353 -966
rect 5439 -1022 5495 -966
rect 5581 -1022 5637 -966
rect 5723 -1022 5779 -966
rect 5865 -1022 5921 -966
rect 6007 -1022 6063 -966
rect 6149 -1022 6205 -966
rect 6291 -1022 6347 -966
rect 6433 -1022 6489 -966
rect 6575 -1022 6631 -966
rect 6717 -1022 6773 -966
rect 6859 -1022 6915 -966
rect 7001 -1022 7057 -966
rect 7143 -1022 7199 -966
rect 7285 -1022 7341 -966
rect -7341 -1164 -7285 -1108
rect -7199 -1164 -7143 -1108
rect -7057 -1164 -7001 -1108
rect -6915 -1164 -6859 -1108
rect -6773 -1164 -6717 -1108
rect -6631 -1164 -6575 -1108
rect -6489 -1164 -6433 -1108
rect -6347 -1164 -6291 -1108
rect -6205 -1164 -6149 -1108
rect -6063 -1164 -6007 -1108
rect -5921 -1164 -5865 -1108
rect -5779 -1164 -5723 -1108
rect -5637 -1164 -5581 -1108
rect -5495 -1164 -5439 -1108
rect -5353 -1164 -5297 -1108
rect -5211 -1164 -5155 -1108
rect -5069 -1164 -5013 -1108
rect -4927 -1164 -4871 -1108
rect -4785 -1164 -4729 -1108
rect -4643 -1164 -4587 -1108
rect -4501 -1164 -4445 -1108
rect -4359 -1164 -4303 -1108
rect -4217 -1164 -4161 -1108
rect -4075 -1164 -4019 -1108
rect -3933 -1164 -3877 -1108
rect -3791 -1164 -3735 -1108
rect -3649 -1164 -3593 -1108
rect -3507 -1164 -3451 -1108
rect -3365 -1164 -3309 -1108
rect -3223 -1164 -3167 -1108
rect -3081 -1164 -3025 -1108
rect -2939 -1164 -2883 -1108
rect -2797 -1164 -2741 -1108
rect -2655 -1164 -2599 -1108
rect -2513 -1164 -2457 -1108
rect -2371 -1164 -2315 -1108
rect -2229 -1164 -2173 -1108
rect -2087 -1164 -2031 -1108
rect -1945 -1164 -1889 -1108
rect -1803 -1164 -1747 -1108
rect -1661 -1164 -1605 -1108
rect -1519 -1164 -1463 -1108
rect -1377 -1164 -1321 -1108
rect -1235 -1164 -1179 -1108
rect -1093 -1164 -1037 -1108
rect -951 -1164 -895 -1108
rect -809 -1164 -753 -1108
rect -667 -1164 -611 -1108
rect -525 -1164 -469 -1108
rect -383 -1164 -327 -1108
rect -241 -1164 -185 -1108
rect -99 -1164 -43 -1108
rect 43 -1164 99 -1108
rect 185 -1164 241 -1108
rect 327 -1164 383 -1108
rect 469 -1164 525 -1108
rect 611 -1164 667 -1108
rect 753 -1164 809 -1108
rect 895 -1164 951 -1108
rect 1037 -1164 1093 -1108
rect 1179 -1164 1235 -1108
rect 1321 -1164 1377 -1108
rect 1463 -1164 1519 -1108
rect 1605 -1164 1661 -1108
rect 1747 -1164 1803 -1108
rect 1889 -1164 1945 -1108
rect 2031 -1164 2087 -1108
rect 2173 -1164 2229 -1108
rect 2315 -1164 2371 -1108
rect 2457 -1164 2513 -1108
rect 2599 -1164 2655 -1108
rect 2741 -1164 2797 -1108
rect 2883 -1164 2939 -1108
rect 3025 -1164 3081 -1108
rect 3167 -1164 3223 -1108
rect 3309 -1164 3365 -1108
rect 3451 -1164 3507 -1108
rect 3593 -1164 3649 -1108
rect 3735 -1164 3791 -1108
rect 3877 -1164 3933 -1108
rect 4019 -1164 4075 -1108
rect 4161 -1164 4217 -1108
rect 4303 -1164 4359 -1108
rect 4445 -1164 4501 -1108
rect 4587 -1164 4643 -1108
rect 4729 -1164 4785 -1108
rect 4871 -1164 4927 -1108
rect 5013 -1164 5069 -1108
rect 5155 -1164 5211 -1108
rect 5297 -1164 5353 -1108
rect 5439 -1164 5495 -1108
rect 5581 -1164 5637 -1108
rect 5723 -1164 5779 -1108
rect 5865 -1164 5921 -1108
rect 6007 -1164 6063 -1108
rect 6149 -1164 6205 -1108
rect 6291 -1164 6347 -1108
rect 6433 -1164 6489 -1108
rect 6575 -1164 6631 -1108
rect 6717 -1164 6773 -1108
rect 6859 -1164 6915 -1108
rect 7001 -1164 7057 -1108
rect 7143 -1164 7199 -1108
rect 7285 -1164 7341 -1108
rect -7341 -1306 -7285 -1250
rect -7199 -1306 -7143 -1250
rect -7057 -1306 -7001 -1250
rect -6915 -1306 -6859 -1250
rect -6773 -1306 -6717 -1250
rect -6631 -1306 -6575 -1250
rect -6489 -1306 -6433 -1250
rect -6347 -1306 -6291 -1250
rect -6205 -1306 -6149 -1250
rect -6063 -1306 -6007 -1250
rect -5921 -1306 -5865 -1250
rect -5779 -1306 -5723 -1250
rect -5637 -1306 -5581 -1250
rect -5495 -1306 -5439 -1250
rect -5353 -1306 -5297 -1250
rect -5211 -1306 -5155 -1250
rect -5069 -1306 -5013 -1250
rect -4927 -1306 -4871 -1250
rect -4785 -1306 -4729 -1250
rect -4643 -1306 -4587 -1250
rect -4501 -1306 -4445 -1250
rect -4359 -1306 -4303 -1250
rect -4217 -1306 -4161 -1250
rect -4075 -1306 -4019 -1250
rect -3933 -1306 -3877 -1250
rect -3791 -1306 -3735 -1250
rect -3649 -1306 -3593 -1250
rect -3507 -1306 -3451 -1250
rect -3365 -1306 -3309 -1250
rect -3223 -1306 -3167 -1250
rect -3081 -1306 -3025 -1250
rect -2939 -1306 -2883 -1250
rect -2797 -1306 -2741 -1250
rect -2655 -1306 -2599 -1250
rect -2513 -1306 -2457 -1250
rect -2371 -1306 -2315 -1250
rect -2229 -1306 -2173 -1250
rect -2087 -1306 -2031 -1250
rect -1945 -1306 -1889 -1250
rect -1803 -1306 -1747 -1250
rect -1661 -1306 -1605 -1250
rect -1519 -1306 -1463 -1250
rect -1377 -1306 -1321 -1250
rect -1235 -1306 -1179 -1250
rect -1093 -1306 -1037 -1250
rect -951 -1306 -895 -1250
rect -809 -1306 -753 -1250
rect -667 -1306 -611 -1250
rect -525 -1306 -469 -1250
rect -383 -1306 -327 -1250
rect -241 -1306 -185 -1250
rect -99 -1306 -43 -1250
rect 43 -1306 99 -1250
rect 185 -1306 241 -1250
rect 327 -1306 383 -1250
rect 469 -1306 525 -1250
rect 611 -1306 667 -1250
rect 753 -1306 809 -1250
rect 895 -1306 951 -1250
rect 1037 -1306 1093 -1250
rect 1179 -1306 1235 -1250
rect 1321 -1306 1377 -1250
rect 1463 -1306 1519 -1250
rect 1605 -1306 1661 -1250
rect 1747 -1306 1803 -1250
rect 1889 -1306 1945 -1250
rect 2031 -1306 2087 -1250
rect 2173 -1306 2229 -1250
rect 2315 -1306 2371 -1250
rect 2457 -1306 2513 -1250
rect 2599 -1306 2655 -1250
rect 2741 -1306 2797 -1250
rect 2883 -1306 2939 -1250
rect 3025 -1306 3081 -1250
rect 3167 -1306 3223 -1250
rect 3309 -1306 3365 -1250
rect 3451 -1306 3507 -1250
rect 3593 -1306 3649 -1250
rect 3735 -1306 3791 -1250
rect 3877 -1306 3933 -1250
rect 4019 -1306 4075 -1250
rect 4161 -1306 4217 -1250
rect 4303 -1306 4359 -1250
rect 4445 -1306 4501 -1250
rect 4587 -1306 4643 -1250
rect 4729 -1306 4785 -1250
rect 4871 -1306 4927 -1250
rect 5013 -1306 5069 -1250
rect 5155 -1306 5211 -1250
rect 5297 -1306 5353 -1250
rect 5439 -1306 5495 -1250
rect 5581 -1306 5637 -1250
rect 5723 -1306 5779 -1250
rect 5865 -1306 5921 -1250
rect 6007 -1306 6063 -1250
rect 6149 -1306 6205 -1250
rect 6291 -1306 6347 -1250
rect 6433 -1306 6489 -1250
rect 6575 -1306 6631 -1250
rect 6717 -1306 6773 -1250
rect 6859 -1306 6915 -1250
rect 7001 -1306 7057 -1250
rect 7143 -1306 7199 -1250
rect 7285 -1306 7341 -1250
rect -7341 -1448 -7285 -1392
rect -7199 -1448 -7143 -1392
rect -7057 -1448 -7001 -1392
rect -6915 -1448 -6859 -1392
rect -6773 -1448 -6717 -1392
rect -6631 -1448 -6575 -1392
rect -6489 -1448 -6433 -1392
rect -6347 -1448 -6291 -1392
rect -6205 -1448 -6149 -1392
rect -6063 -1448 -6007 -1392
rect -5921 -1448 -5865 -1392
rect -5779 -1448 -5723 -1392
rect -5637 -1448 -5581 -1392
rect -5495 -1448 -5439 -1392
rect -5353 -1448 -5297 -1392
rect -5211 -1448 -5155 -1392
rect -5069 -1448 -5013 -1392
rect -4927 -1448 -4871 -1392
rect -4785 -1448 -4729 -1392
rect -4643 -1448 -4587 -1392
rect -4501 -1448 -4445 -1392
rect -4359 -1448 -4303 -1392
rect -4217 -1448 -4161 -1392
rect -4075 -1448 -4019 -1392
rect -3933 -1448 -3877 -1392
rect -3791 -1448 -3735 -1392
rect -3649 -1448 -3593 -1392
rect -3507 -1448 -3451 -1392
rect -3365 -1448 -3309 -1392
rect -3223 -1448 -3167 -1392
rect -3081 -1448 -3025 -1392
rect -2939 -1448 -2883 -1392
rect -2797 -1448 -2741 -1392
rect -2655 -1448 -2599 -1392
rect -2513 -1448 -2457 -1392
rect -2371 -1448 -2315 -1392
rect -2229 -1448 -2173 -1392
rect -2087 -1448 -2031 -1392
rect -1945 -1448 -1889 -1392
rect -1803 -1448 -1747 -1392
rect -1661 -1448 -1605 -1392
rect -1519 -1448 -1463 -1392
rect -1377 -1448 -1321 -1392
rect -1235 -1448 -1179 -1392
rect -1093 -1448 -1037 -1392
rect -951 -1448 -895 -1392
rect -809 -1448 -753 -1392
rect -667 -1448 -611 -1392
rect -525 -1448 -469 -1392
rect -383 -1448 -327 -1392
rect -241 -1448 -185 -1392
rect -99 -1448 -43 -1392
rect 43 -1448 99 -1392
rect 185 -1448 241 -1392
rect 327 -1448 383 -1392
rect 469 -1448 525 -1392
rect 611 -1448 667 -1392
rect 753 -1448 809 -1392
rect 895 -1448 951 -1392
rect 1037 -1448 1093 -1392
rect 1179 -1448 1235 -1392
rect 1321 -1448 1377 -1392
rect 1463 -1448 1519 -1392
rect 1605 -1448 1661 -1392
rect 1747 -1448 1803 -1392
rect 1889 -1448 1945 -1392
rect 2031 -1448 2087 -1392
rect 2173 -1448 2229 -1392
rect 2315 -1448 2371 -1392
rect 2457 -1448 2513 -1392
rect 2599 -1448 2655 -1392
rect 2741 -1448 2797 -1392
rect 2883 -1448 2939 -1392
rect 3025 -1448 3081 -1392
rect 3167 -1448 3223 -1392
rect 3309 -1448 3365 -1392
rect 3451 -1448 3507 -1392
rect 3593 -1448 3649 -1392
rect 3735 -1448 3791 -1392
rect 3877 -1448 3933 -1392
rect 4019 -1448 4075 -1392
rect 4161 -1448 4217 -1392
rect 4303 -1448 4359 -1392
rect 4445 -1448 4501 -1392
rect 4587 -1448 4643 -1392
rect 4729 -1448 4785 -1392
rect 4871 -1448 4927 -1392
rect 5013 -1448 5069 -1392
rect 5155 -1448 5211 -1392
rect 5297 -1448 5353 -1392
rect 5439 -1448 5495 -1392
rect 5581 -1448 5637 -1392
rect 5723 -1448 5779 -1392
rect 5865 -1448 5921 -1392
rect 6007 -1448 6063 -1392
rect 6149 -1448 6205 -1392
rect 6291 -1448 6347 -1392
rect 6433 -1448 6489 -1392
rect 6575 -1448 6631 -1392
rect 6717 -1448 6773 -1392
rect 6859 -1448 6915 -1392
rect 7001 -1448 7057 -1392
rect 7143 -1448 7199 -1392
rect 7285 -1448 7341 -1392
<< metal4 >>
rect -7351 1448 7351 1458
rect -7351 1392 -7341 1448
rect -7285 1392 -7199 1448
rect -7143 1392 -7057 1448
rect -7001 1392 -6915 1448
rect -6859 1392 -6773 1448
rect -6717 1392 -6631 1448
rect -6575 1392 -6489 1448
rect -6433 1392 -6347 1448
rect -6291 1392 -6205 1448
rect -6149 1392 -6063 1448
rect -6007 1392 -5921 1448
rect -5865 1392 -5779 1448
rect -5723 1392 -5637 1448
rect -5581 1392 -5495 1448
rect -5439 1392 -5353 1448
rect -5297 1392 -5211 1448
rect -5155 1392 -5069 1448
rect -5013 1392 -4927 1448
rect -4871 1392 -4785 1448
rect -4729 1392 -4643 1448
rect -4587 1392 -4501 1448
rect -4445 1392 -4359 1448
rect -4303 1392 -4217 1448
rect -4161 1392 -4075 1448
rect -4019 1392 -3933 1448
rect -3877 1392 -3791 1448
rect -3735 1392 -3649 1448
rect -3593 1392 -3507 1448
rect -3451 1392 -3365 1448
rect -3309 1392 -3223 1448
rect -3167 1392 -3081 1448
rect -3025 1392 -2939 1448
rect -2883 1392 -2797 1448
rect -2741 1392 -2655 1448
rect -2599 1392 -2513 1448
rect -2457 1392 -2371 1448
rect -2315 1392 -2229 1448
rect -2173 1392 -2087 1448
rect -2031 1392 -1945 1448
rect -1889 1392 -1803 1448
rect -1747 1392 -1661 1448
rect -1605 1392 -1519 1448
rect -1463 1392 -1377 1448
rect -1321 1392 -1235 1448
rect -1179 1392 -1093 1448
rect -1037 1392 -951 1448
rect -895 1392 -809 1448
rect -753 1392 -667 1448
rect -611 1392 -525 1448
rect -469 1392 -383 1448
rect -327 1392 -241 1448
rect -185 1392 -99 1448
rect -43 1392 43 1448
rect 99 1392 185 1448
rect 241 1392 327 1448
rect 383 1392 469 1448
rect 525 1392 611 1448
rect 667 1392 753 1448
rect 809 1392 895 1448
rect 951 1392 1037 1448
rect 1093 1392 1179 1448
rect 1235 1392 1321 1448
rect 1377 1392 1463 1448
rect 1519 1392 1605 1448
rect 1661 1392 1747 1448
rect 1803 1392 1889 1448
rect 1945 1392 2031 1448
rect 2087 1392 2173 1448
rect 2229 1392 2315 1448
rect 2371 1392 2457 1448
rect 2513 1392 2599 1448
rect 2655 1392 2741 1448
rect 2797 1392 2883 1448
rect 2939 1392 3025 1448
rect 3081 1392 3167 1448
rect 3223 1392 3309 1448
rect 3365 1392 3451 1448
rect 3507 1392 3593 1448
rect 3649 1392 3735 1448
rect 3791 1392 3877 1448
rect 3933 1392 4019 1448
rect 4075 1392 4161 1448
rect 4217 1392 4303 1448
rect 4359 1392 4445 1448
rect 4501 1392 4587 1448
rect 4643 1392 4729 1448
rect 4785 1392 4871 1448
rect 4927 1392 5013 1448
rect 5069 1392 5155 1448
rect 5211 1392 5297 1448
rect 5353 1392 5439 1448
rect 5495 1392 5581 1448
rect 5637 1392 5723 1448
rect 5779 1392 5865 1448
rect 5921 1392 6007 1448
rect 6063 1392 6149 1448
rect 6205 1392 6291 1448
rect 6347 1392 6433 1448
rect 6489 1392 6575 1448
rect 6631 1392 6717 1448
rect 6773 1392 6859 1448
rect 6915 1392 7001 1448
rect 7057 1392 7143 1448
rect 7199 1392 7285 1448
rect 7341 1392 7351 1448
rect -7351 1306 7351 1392
rect -7351 1250 -7341 1306
rect -7285 1250 -7199 1306
rect -7143 1250 -7057 1306
rect -7001 1250 -6915 1306
rect -6859 1250 -6773 1306
rect -6717 1250 -6631 1306
rect -6575 1250 -6489 1306
rect -6433 1250 -6347 1306
rect -6291 1250 -6205 1306
rect -6149 1250 -6063 1306
rect -6007 1250 -5921 1306
rect -5865 1250 -5779 1306
rect -5723 1250 -5637 1306
rect -5581 1250 -5495 1306
rect -5439 1250 -5353 1306
rect -5297 1250 -5211 1306
rect -5155 1250 -5069 1306
rect -5013 1250 -4927 1306
rect -4871 1250 -4785 1306
rect -4729 1250 -4643 1306
rect -4587 1250 -4501 1306
rect -4445 1250 -4359 1306
rect -4303 1250 -4217 1306
rect -4161 1250 -4075 1306
rect -4019 1250 -3933 1306
rect -3877 1250 -3791 1306
rect -3735 1250 -3649 1306
rect -3593 1250 -3507 1306
rect -3451 1250 -3365 1306
rect -3309 1250 -3223 1306
rect -3167 1250 -3081 1306
rect -3025 1250 -2939 1306
rect -2883 1250 -2797 1306
rect -2741 1250 -2655 1306
rect -2599 1250 -2513 1306
rect -2457 1250 -2371 1306
rect -2315 1250 -2229 1306
rect -2173 1250 -2087 1306
rect -2031 1250 -1945 1306
rect -1889 1250 -1803 1306
rect -1747 1250 -1661 1306
rect -1605 1250 -1519 1306
rect -1463 1250 -1377 1306
rect -1321 1250 -1235 1306
rect -1179 1250 -1093 1306
rect -1037 1250 -951 1306
rect -895 1250 -809 1306
rect -753 1250 -667 1306
rect -611 1250 -525 1306
rect -469 1250 -383 1306
rect -327 1250 -241 1306
rect -185 1250 -99 1306
rect -43 1250 43 1306
rect 99 1250 185 1306
rect 241 1250 327 1306
rect 383 1250 469 1306
rect 525 1250 611 1306
rect 667 1250 753 1306
rect 809 1250 895 1306
rect 951 1250 1037 1306
rect 1093 1250 1179 1306
rect 1235 1250 1321 1306
rect 1377 1250 1463 1306
rect 1519 1250 1605 1306
rect 1661 1250 1747 1306
rect 1803 1250 1889 1306
rect 1945 1250 2031 1306
rect 2087 1250 2173 1306
rect 2229 1250 2315 1306
rect 2371 1250 2457 1306
rect 2513 1250 2599 1306
rect 2655 1250 2741 1306
rect 2797 1250 2883 1306
rect 2939 1250 3025 1306
rect 3081 1250 3167 1306
rect 3223 1250 3309 1306
rect 3365 1250 3451 1306
rect 3507 1250 3593 1306
rect 3649 1250 3735 1306
rect 3791 1250 3877 1306
rect 3933 1250 4019 1306
rect 4075 1250 4161 1306
rect 4217 1250 4303 1306
rect 4359 1250 4445 1306
rect 4501 1250 4587 1306
rect 4643 1250 4729 1306
rect 4785 1250 4871 1306
rect 4927 1250 5013 1306
rect 5069 1250 5155 1306
rect 5211 1250 5297 1306
rect 5353 1250 5439 1306
rect 5495 1250 5581 1306
rect 5637 1250 5723 1306
rect 5779 1250 5865 1306
rect 5921 1250 6007 1306
rect 6063 1250 6149 1306
rect 6205 1250 6291 1306
rect 6347 1250 6433 1306
rect 6489 1250 6575 1306
rect 6631 1250 6717 1306
rect 6773 1250 6859 1306
rect 6915 1250 7001 1306
rect 7057 1250 7143 1306
rect 7199 1250 7285 1306
rect 7341 1250 7351 1306
rect -7351 1164 7351 1250
rect -7351 1108 -7341 1164
rect -7285 1108 -7199 1164
rect -7143 1108 -7057 1164
rect -7001 1108 -6915 1164
rect -6859 1108 -6773 1164
rect -6717 1108 -6631 1164
rect -6575 1108 -6489 1164
rect -6433 1108 -6347 1164
rect -6291 1108 -6205 1164
rect -6149 1108 -6063 1164
rect -6007 1108 -5921 1164
rect -5865 1108 -5779 1164
rect -5723 1108 -5637 1164
rect -5581 1108 -5495 1164
rect -5439 1108 -5353 1164
rect -5297 1108 -5211 1164
rect -5155 1108 -5069 1164
rect -5013 1108 -4927 1164
rect -4871 1108 -4785 1164
rect -4729 1108 -4643 1164
rect -4587 1108 -4501 1164
rect -4445 1108 -4359 1164
rect -4303 1108 -4217 1164
rect -4161 1108 -4075 1164
rect -4019 1108 -3933 1164
rect -3877 1108 -3791 1164
rect -3735 1108 -3649 1164
rect -3593 1108 -3507 1164
rect -3451 1108 -3365 1164
rect -3309 1108 -3223 1164
rect -3167 1108 -3081 1164
rect -3025 1108 -2939 1164
rect -2883 1108 -2797 1164
rect -2741 1108 -2655 1164
rect -2599 1108 -2513 1164
rect -2457 1108 -2371 1164
rect -2315 1108 -2229 1164
rect -2173 1108 -2087 1164
rect -2031 1108 -1945 1164
rect -1889 1108 -1803 1164
rect -1747 1108 -1661 1164
rect -1605 1108 -1519 1164
rect -1463 1108 -1377 1164
rect -1321 1108 -1235 1164
rect -1179 1108 -1093 1164
rect -1037 1108 -951 1164
rect -895 1108 -809 1164
rect -753 1108 -667 1164
rect -611 1108 -525 1164
rect -469 1108 -383 1164
rect -327 1108 -241 1164
rect -185 1108 -99 1164
rect -43 1108 43 1164
rect 99 1108 185 1164
rect 241 1108 327 1164
rect 383 1108 469 1164
rect 525 1108 611 1164
rect 667 1108 753 1164
rect 809 1108 895 1164
rect 951 1108 1037 1164
rect 1093 1108 1179 1164
rect 1235 1108 1321 1164
rect 1377 1108 1463 1164
rect 1519 1108 1605 1164
rect 1661 1108 1747 1164
rect 1803 1108 1889 1164
rect 1945 1108 2031 1164
rect 2087 1108 2173 1164
rect 2229 1108 2315 1164
rect 2371 1108 2457 1164
rect 2513 1108 2599 1164
rect 2655 1108 2741 1164
rect 2797 1108 2883 1164
rect 2939 1108 3025 1164
rect 3081 1108 3167 1164
rect 3223 1108 3309 1164
rect 3365 1108 3451 1164
rect 3507 1108 3593 1164
rect 3649 1108 3735 1164
rect 3791 1108 3877 1164
rect 3933 1108 4019 1164
rect 4075 1108 4161 1164
rect 4217 1108 4303 1164
rect 4359 1108 4445 1164
rect 4501 1108 4587 1164
rect 4643 1108 4729 1164
rect 4785 1108 4871 1164
rect 4927 1108 5013 1164
rect 5069 1108 5155 1164
rect 5211 1108 5297 1164
rect 5353 1108 5439 1164
rect 5495 1108 5581 1164
rect 5637 1108 5723 1164
rect 5779 1108 5865 1164
rect 5921 1108 6007 1164
rect 6063 1108 6149 1164
rect 6205 1108 6291 1164
rect 6347 1108 6433 1164
rect 6489 1108 6575 1164
rect 6631 1108 6717 1164
rect 6773 1108 6859 1164
rect 6915 1108 7001 1164
rect 7057 1108 7143 1164
rect 7199 1108 7285 1164
rect 7341 1108 7351 1164
rect -7351 1022 7351 1108
rect -7351 966 -7341 1022
rect -7285 966 -7199 1022
rect -7143 966 -7057 1022
rect -7001 966 -6915 1022
rect -6859 966 -6773 1022
rect -6717 966 -6631 1022
rect -6575 966 -6489 1022
rect -6433 966 -6347 1022
rect -6291 966 -6205 1022
rect -6149 966 -6063 1022
rect -6007 966 -5921 1022
rect -5865 966 -5779 1022
rect -5723 966 -5637 1022
rect -5581 966 -5495 1022
rect -5439 966 -5353 1022
rect -5297 966 -5211 1022
rect -5155 966 -5069 1022
rect -5013 966 -4927 1022
rect -4871 966 -4785 1022
rect -4729 966 -4643 1022
rect -4587 966 -4501 1022
rect -4445 966 -4359 1022
rect -4303 966 -4217 1022
rect -4161 966 -4075 1022
rect -4019 966 -3933 1022
rect -3877 966 -3791 1022
rect -3735 966 -3649 1022
rect -3593 966 -3507 1022
rect -3451 966 -3365 1022
rect -3309 966 -3223 1022
rect -3167 966 -3081 1022
rect -3025 966 -2939 1022
rect -2883 966 -2797 1022
rect -2741 966 -2655 1022
rect -2599 966 -2513 1022
rect -2457 966 -2371 1022
rect -2315 966 -2229 1022
rect -2173 966 -2087 1022
rect -2031 966 -1945 1022
rect -1889 966 -1803 1022
rect -1747 966 -1661 1022
rect -1605 966 -1519 1022
rect -1463 966 -1377 1022
rect -1321 966 -1235 1022
rect -1179 966 -1093 1022
rect -1037 966 -951 1022
rect -895 966 -809 1022
rect -753 966 -667 1022
rect -611 966 -525 1022
rect -469 966 -383 1022
rect -327 966 -241 1022
rect -185 966 -99 1022
rect -43 966 43 1022
rect 99 966 185 1022
rect 241 966 327 1022
rect 383 966 469 1022
rect 525 966 611 1022
rect 667 966 753 1022
rect 809 966 895 1022
rect 951 966 1037 1022
rect 1093 966 1179 1022
rect 1235 966 1321 1022
rect 1377 966 1463 1022
rect 1519 966 1605 1022
rect 1661 966 1747 1022
rect 1803 966 1889 1022
rect 1945 966 2031 1022
rect 2087 966 2173 1022
rect 2229 966 2315 1022
rect 2371 966 2457 1022
rect 2513 966 2599 1022
rect 2655 966 2741 1022
rect 2797 966 2883 1022
rect 2939 966 3025 1022
rect 3081 966 3167 1022
rect 3223 966 3309 1022
rect 3365 966 3451 1022
rect 3507 966 3593 1022
rect 3649 966 3735 1022
rect 3791 966 3877 1022
rect 3933 966 4019 1022
rect 4075 966 4161 1022
rect 4217 966 4303 1022
rect 4359 966 4445 1022
rect 4501 966 4587 1022
rect 4643 966 4729 1022
rect 4785 966 4871 1022
rect 4927 966 5013 1022
rect 5069 966 5155 1022
rect 5211 966 5297 1022
rect 5353 966 5439 1022
rect 5495 966 5581 1022
rect 5637 966 5723 1022
rect 5779 966 5865 1022
rect 5921 966 6007 1022
rect 6063 966 6149 1022
rect 6205 966 6291 1022
rect 6347 966 6433 1022
rect 6489 966 6575 1022
rect 6631 966 6717 1022
rect 6773 966 6859 1022
rect 6915 966 7001 1022
rect 7057 966 7143 1022
rect 7199 966 7285 1022
rect 7341 966 7351 1022
rect -7351 880 7351 966
rect -7351 824 -7341 880
rect -7285 824 -7199 880
rect -7143 824 -7057 880
rect -7001 824 -6915 880
rect -6859 824 -6773 880
rect -6717 824 -6631 880
rect -6575 824 -6489 880
rect -6433 824 -6347 880
rect -6291 824 -6205 880
rect -6149 824 -6063 880
rect -6007 824 -5921 880
rect -5865 824 -5779 880
rect -5723 824 -5637 880
rect -5581 824 -5495 880
rect -5439 824 -5353 880
rect -5297 824 -5211 880
rect -5155 824 -5069 880
rect -5013 824 -4927 880
rect -4871 824 -4785 880
rect -4729 824 -4643 880
rect -4587 824 -4501 880
rect -4445 824 -4359 880
rect -4303 824 -4217 880
rect -4161 824 -4075 880
rect -4019 824 -3933 880
rect -3877 824 -3791 880
rect -3735 824 -3649 880
rect -3593 824 -3507 880
rect -3451 824 -3365 880
rect -3309 824 -3223 880
rect -3167 824 -3081 880
rect -3025 824 -2939 880
rect -2883 824 -2797 880
rect -2741 824 -2655 880
rect -2599 824 -2513 880
rect -2457 824 -2371 880
rect -2315 824 -2229 880
rect -2173 824 -2087 880
rect -2031 824 -1945 880
rect -1889 824 -1803 880
rect -1747 824 -1661 880
rect -1605 824 -1519 880
rect -1463 824 -1377 880
rect -1321 824 -1235 880
rect -1179 824 -1093 880
rect -1037 824 -951 880
rect -895 824 -809 880
rect -753 824 -667 880
rect -611 824 -525 880
rect -469 824 -383 880
rect -327 824 -241 880
rect -185 824 -99 880
rect -43 824 43 880
rect 99 824 185 880
rect 241 824 327 880
rect 383 824 469 880
rect 525 824 611 880
rect 667 824 753 880
rect 809 824 895 880
rect 951 824 1037 880
rect 1093 824 1179 880
rect 1235 824 1321 880
rect 1377 824 1463 880
rect 1519 824 1605 880
rect 1661 824 1747 880
rect 1803 824 1889 880
rect 1945 824 2031 880
rect 2087 824 2173 880
rect 2229 824 2315 880
rect 2371 824 2457 880
rect 2513 824 2599 880
rect 2655 824 2741 880
rect 2797 824 2883 880
rect 2939 824 3025 880
rect 3081 824 3167 880
rect 3223 824 3309 880
rect 3365 824 3451 880
rect 3507 824 3593 880
rect 3649 824 3735 880
rect 3791 824 3877 880
rect 3933 824 4019 880
rect 4075 824 4161 880
rect 4217 824 4303 880
rect 4359 824 4445 880
rect 4501 824 4587 880
rect 4643 824 4729 880
rect 4785 824 4871 880
rect 4927 824 5013 880
rect 5069 824 5155 880
rect 5211 824 5297 880
rect 5353 824 5439 880
rect 5495 824 5581 880
rect 5637 824 5723 880
rect 5779 824 5865 880
rect 5921 824 6007 880
rect 6063 824 6149 880
rect 6205 824 6291 880
rect 6347 824 6433 880
rect 6489 824 6575 880
rect 6631 824 6717 880
rect 6773 824 6859 880
rect 6915 824 7001 880
rect 7057 824 7143 880
rect 7199 824 7285 880
rect 7341 824 7351 880
rect -7351 738 7351 824
rect -7351 682 -7341 738
rect -7285 682 -7199 738
rect -7143 682 -7057 738
rect -7001 682 -6915 738
rect -6859 682 -6773 738
rect -6717 682 -6631 738
rect -6575 682 -6489 738
rect -6433 682 -6347 738
rect -6291 682 -6205 738
rect -6149 682 -6063 738
rect -6007 682 -5921 738
rect -5865 682 -5779 738
rect -5723 682 -5637 738
rect -5581 682 -5495 738
rect -5439 682 -5353 738
rect -5297 682 -5211 738
rect -5155 682 -5069 738
rect -5013 682 -4927 738
rect -4871 682 -4785 738
rect -4729 682 -4643 738
rect -4587 682 -4501 738
rect -4445 682 -4359 738
rect -4303 682 -4217 738
rect -4161 682 -4075 738
rect -4019 682 -3933 738
rect -3877 682 -3791 738
rect -3735 682 -3649 738
rect -3593 682 -3507 738
rect -3451 682 -3365 738
rect -3309 682 -3223 738
rect -3167 682 -3081 738
rect -3025 682 -2939 738
rect -2883 682 -2797 738
rect -2741 682 -2655 738
rect -2599 682 -2513 738
rect -2457 682 -2371 738
rect -2315 682 -2229 738
rect -2173 682 -2087 738
rect -2031 682 -1945 738
rect -1889 682 -1803 738
rect -1747 682 -1661 738
rect -1605 682 -1519 738
rect -1463 682 -1377 738
rect -1321 682 -1235 738
rect -1179 682 -1093 738
rect -1037 682 -951 738
rect -895 682 -809 738
rect -753 682 -667 738
rect -611 682 -525 738
rect -469 682 -383 738
rect -327 682 -241 738
rect -185 682 -99 738
rect -43 682 43 738
rect 99 682 185 738
rect 241 682 327 738
rect 383 682 469 738
rect 525 682 611 738
rect 667 682 753 738
rect 809 682 895 738
rect 951 682 1037 738
rect 1093 682 1179 738
rect 1235 682 1321 738
rect 1377 682 1463 738
rect 1519 682 1605 738
rect 1661 682 1747 738
rect 1803 682 1889 738
rect 1945 682 2031 738
rect 2087 682 2173 738
rect 2229 682 2315 738
rect 2371 682 2457 738
rect 2513 682 2599 738
rect 2655 682 2741 738
rect 2797 682 2883 738
rect 2939 682 3025 738
rect 3081 682 3167 738
rect 3223 682 3309 738
rect 3365 682 3451 738
rect 3507 682 3593 738
rect 3649 682 3735 738
rect 3791 682 3877 738
rect 3933 682 4019 738
rect 4075 682 4161 738
rect 4217 682 4303 738
rect 4359 682 4445 738
rect 4501 682 4587 738
rect 4643 682 4729 738
rect 4785 682 4871 738
rect 4927 682 5013 738
rect 5069 682 5155 738
rect 5211 682 5297 738
rect 5353 682 5439 738
rect 5495 682 5581 738
rect 5637 682 5723 738
rect 5779 682 5865 738
rect 5921 682 6007 738
rect 6063 682 6149 738
rect 6205 682 6291 738
rect 6347 682 6433 738
rect 6489 682 6575 738
rect 6631 682 6717 738
rect 6773 682 6859 738
rect 6915 682 7001 738
rect 7057 682 7143 738
rect 7199 682 7285 738
rect 7341 682 7351 738
rect -7351 596 7351 682
rect -7351 540 -7341 596
rect -7285 540 -7199 596
rect -7143 540 -7057 596
rect -7001 540 -6915 596
rect -6859 540 -6773 596
rect -6717 540 -6631 596
rect -6575 540 -6489 596
rect -6433 540 -6347 596
rect -6291 540 -6205 596
rect -6149 540 -6063 596
rect -6007 540 -5921 596
rect -5865 540 -5779 596
rect -5723 540 -5637 596
rect -5581 540 -5495 596
rect -5439 540 -5353 596
rect -5297 540 -5211 596
rect -5155 540 -5069 596
rect -5013 540 -4927 596
rect -4871 540 -4785 596
rect -4729 540 -4643 596
rect -4587 540 -4501 596
rect -4445 540 -4359 596
rect -4303 540 -4217 596
rect -4161 540 -4075 596
rect -4019 540 -3933 596
rect -3877 540 -3791 596
rect -3735 540 -3649 596
rect -3593 540 -3507 596
rect -3451 540 -3365 596
rect -3309 540 -3223 596
rect -3167 540 -3081 596
rect -3025 540 -2939 596
rect -2883 540 -2797 596
rect -2741 540 -2655 596
rect -2599 540 -2513 596
rect -2457 540 -2371 596
rect -2315 540 -2229 596
rect -2173 540 -2087 596
rect -2031 540 -1945 596
rect -1889 540 -1803 596
rect -1747 540 -1661 596
rect -1605 540 -1519 596
rect -1463 540 -1377 596
rect -1321 540 -1235 596
rect -1179 540 -1093 596
rect -1037 540 -951 596
rect -895 540 -809 596
rect -753 540 -667 596
rect -611 540 -525 596
rect -469 540 -383 596
rect -327 540 -241 596
rect -185 540 -99 596
rect -43 540 43 596
rect 99 540 185 596
rect 241 540 327 596
rect 383 540 469 596
rect 525 540 611 596
rect 667 540 753 596
rect 809 540 895 596
rect 951 540 1037 596
rect 1093 540 1179 596
rect 1235 540 1321 596
rect 1377 540 1463 596
rect 1519 540 1605 596
rect 1661 540 1747 596
rect 1803 540 1889 596
rect 1945 540 2031 596
rect 2087 540 2173 596
rect 2229 540 2315 596
rect 2371 540 2457 596
rect 2513 540 2599 596
rect 2655 540 2741 596
rect 2797 540 2883 596
rect 2939 540 3025 596
rect 3081 540 3167 596
rect 3223 540 3309 596
rect 3365 540 3451 596
rect 3507 540 3593 596
rect 3649 540 3735 596
rect 3791 540 3877 596
rect 3933 540 4019 596
rect 4075 540 4161 596
rect 4217 540 4303 596
rect 4359 540 4445 596
rect 4501 540 4587 596
rect 4643 540 4729 596
rect 4785 540 4871 596
rect 4927 540 5013 596
rect 5069 540 5155 596
rect 5211 540 5297 596
rect 5353 540 5439 596
rect 5495 540 5581 596
rect 5637 540 5723 596
rect 5779 540 5865 596
rect 5921 540 6007 596
rect 6063 540 6149 596
rect 6205 540 6291 596
rect 6347 540 6433 596
rect 6489 540 6575 596
rect 6631 540 6717 596
rect 6773 540 6859 596
rect 6915 540 7001 596
rect 7057 540 7143 596
rect 7199 540 7285 596
rect 7341 540 7351 596
rect -7351 454 7351 540
rect -7351 398 -7341 454
rect -7285 398 -7199 454
rect -7143 398 -7057 454
rect -7001 398 -6915 454
rect -6859 398 -6773 454
rect -6717 398 -6631 454
rect -6575 398 -6489 454
rect -6433 398 -6347 454
rect -6291 398 -6205 454
rect -6149 398 -6063 454
rect -6007 398 -5921 454
rect -5865 398 -5779 454
rect -5723 398 -5637 454
rect -5581 398 -5495 454
rect -5439 398 -5353 454
rect -5297 398 -5211 454
rect -5155 398 -5069 454
rect -5013 398 -4927 454
rect -4871 398 -4785 454
rect -4729 398 -4643 454
rect -4587 398 -4501 454
rect -4445 398 -4359 454
rect -4303 398 -4217 454
rect -4161 398 -4075 454
rect -4019 398 -3933 454
rect -3877 398 -3791 454
rect -3735 398 -3649 454
rect -3593 398 -3507 454
rect -3451 398 -3365 454
rect -3309 398 -3223 454
rect -3167 398 -3081 454
rect -3025 398 -2939 454
rect -2883 398 -2797 454
rect -2741 398 -2655 454
rect -2599 398 -2513 454
rect -2457 398 -2371 454
rect -2315 398 -2229 454
rect -2173 398 -2087 454
rect -2031 398 -1945 454
rect -1889 398 -1803 454
rect -1747 398 -1661 454
rect -1605 398 -1519 454
rect -1463 398 -1377 454
rect -1321 398 -1235 454
rect -1179 398 -1093 454
rect -1037 398 -951 454
rect -895 398 -809 454
rect -753 398 -667 454
rect -611 398 -525 454
rect -469 398 -383 454
rect -327 398 -241 454
rect -185 398 -99 454
rect -43 398 43 454
rect 99 398 185 454
rect 241 398 327 454
rect 383 398 469 454
rect 525 398 611 454
rect 667 398 753 454
rect 809 398 895 454
rect 951 398 1037 454
rect 1093 398 1179 454
rect 1235 398 1321 454
rect 1377 398 1463 454
rect 1519 398 1605 454
rect 1661 398 1747 454
rect 1803 398 1889 454
rect 1945 398 2031 454
rect 2087 398 2173 454
rect 2229 398 2315 454
rect 2371 398 2457 454
rect 2513 398 2599 454
rect 2655 398 2741 454
rect 2797 398 2883 454
rect 2939 398 3025 454
rect 3081 398 3167 454
rect 3223 398 3309 454
rect 3365 398 3451 454
rect 3507 398 3593 454
rect 3649 398 3735 454
rect 3791 398 3877 454
rect 3933 398 4019 454
rect 4075 398 4161 454
rect 4217 398 4303 454
rect 4359 398 4445 454
rect 4501 398 4587 454
rect 4643 398 4729 454
rect 4785 398 4871 454
rect 4927 398 5013 454
rect 5069 398 5155 454
rect 5211 398 5297 454
rect 5353 398 5439 454
rect 5495 398 5581 454
rect 5637 398 5723 454
rect 5779 398 5865 454
rect 5921 398 6007 454
rect 6063 398 6149 454
rect 6205 398 6291 454
rect 6347 398 6433 454
rect 6489 398 6575 454
rect 6631 398 6717 454
rect 6773 398 6859 454
rect 6915 398 7001 454
rect 7057 398 7143 454
rect 7199 398 7285 454
rect 7341 398 7351 454
rect -7351 312 7351 398
rect -7351 256 -7341 312
rect -7285 256 -7199 312
rect -7143 256 -7057 312
rect -7001 256 -6915 312
rect -6859 256 -6773 312
rect -6717 256 -6631 312
rect -6575 256 -6489 312
rect -6433 256 -6347 312
rect -6291 256 -6205 312
rect -6149 256 -6063 312
rect -6007 256 -5921 312
rect -5865 256 -5779 312
rect -5723 256 -5637 312
rect -5581 256 -5495 312
rect -5439 256 -5353 312
rect -5297 256 -5211 312
rect -5155 256 -5069 312
rect -5013 256 -4927 312
rect -4871 256 -4785 312
rect -4729 256 -4643 312
rect -4587 256 -4501 312
rect -4445 256 -4359 312
rect -4303 256 -4217 312
rect -4161 256 -4075 312
rect -4019 256 -3933 312
rect -3877 256 -3791 312
rect -3735 256 -3649 312
rect -3593 256 -3507 312
rect -3451 256 -3365 312
rect -3309 256 -3223 312
rect -3167 256 -3081 312
rect -3025 256 -2939 312
rect -2883 256 -2797 312
rect -2741 256 -2655 312
rect -2599 256 -2513 312
rect -2457 256 -2371 312
rect -2315 256 -2229 312
rect -2173 256 -2087 312
rect -2031 256 -1945 312
rect -1889 256 -1803 312
rect -1747 256 -1661 312
rect -1605 256 -1519 312
rect -1463 256 -1377 312
rect -1321 256 -1235 312
rect -1179 256 -1093 312
rect -1037 256 -951 312
rect -895 256 -809 312
rect -753 256 -667 312
rect -611 256 -525 312
rect -469 256 -383 312
rect -327 256 -241 312
rect -185 256 -99 312
rect -43 256 43 312
rect 99 256 185 312
rect 241 256 327 312
rect 383 256 469 312
rect 525 256 611 312
rect 667 256 753 312
rect 809 256 895 312
rect 951 256 1037 312
rect 1093 256 1179 312
rect 1235 256 1321 312
rect 1377 256 1463 312
rect 1519 256 1605 312
rect 1661 256 1747 312
rect 1803 256 1889 312
rect 1945 256 2031 312
rect 2087 256 2173 312
rect 2229 256 2315 312
rect 2371 256 2457 312
rect 2513 256 2599 312
rect 2655 256 2741 312
rect 2797 256 2883 312
rect 2939 256 3025 312
rect 3081 256 3167 312
rect 3223 256 3309 312
rect 3365 256 3451 312
rect 3507 256 3593 312
rect 3649 256 3735 312
rect 3791 256 3877 312
rect 3933 256 4019 312
rect 4075 256 4161 312
rect 4217 256 4303 312
rect 4359 256 4445 312
rect 4501 256 4587 312
rect 4643 256 4729 312
rect 4785 256 4871 312
rect 4927 256 5013 312
rect 5069 256 5155 312
rect 5211 256 5297 312
rect 5353 256 5439 312
rect 5495 256 5581 312
rect 5637 256 5723 312
rect 5779 256 5865 312
rect 5921 256 6007 312
rect 6063 256 6149 312
rect 6205 256 6291 312
rect 6347 256 6433 312
rect 6489 256 6575 312
rect 6631 256 6717 312
rect 6773 256 6859 312
rect 6915 256 7001 312
rect 7057 256 7143 312
rect 7199 256 7285 312
rect 7341 256 7351 312
rect -7351 170 7351 256
rect -7351 114 -7341 170
rect -7285 114 -7199 170
rect -7143 114 -7057 170
rect -7001 114 -6915 170
rect -6859 114 -6773 170
rect -6717 114 -6631 170
rect -6575 114 -6489 170
rect -6433 114 -6347 170
rect -6291 114 -6205 170
rect -6149 114 -6063 170
rect -6007 114 -5921 170
rect -5865 114 -5779 170
rect -5723 114 -5637 170
rect -5581 114 -5495 170
rect -5439 114 -5353 170
rect -5297 114 -5211 170
rect -5155 114 -5069 170
rect -5013 114 -4927 170
rect -4871 114 -4785 170
rect -4729 114 -4643 170
rect -4587 114 -4501 170
rect -4445 114 -4359 170
rect -4303 114 -4217 170
rect -4161 114 -4075 170
rect -4019 114 -3933 170
rect -3877 114 -3791 170
rect -3735 114 -3649 170
rect -3593 114 -3507 170
rect -3451 114 -3365 170
rect -3309 114 -3223 170
rect -3167 114 -3081 170
rect -3025 114 -2939 170
rect -2883 114 -2797 170
rect -2741 114 -2655 170
rect -2599 114 -2513 170
rect -2457 114 -2371 170
rect -2315 114 -2229 170
rect -2173 114 -2087 170
rect -2031 114 -1945 170
rect -1889 114 -1803 170
rect -1747 114 -1661 170
rect -1605 114 -1519 170
rect -1463 114 -1377 170
rect -1321 114 -1235 170
rect -1179 114 -1093 170
rect -1037 114 -951 170
rect -895 114 -809 170
rect -753 114 -667 170
rect -611 114 -525 170
rect -469 114 -383 170
rect -327 114 -241 170
rect -185 114 -99 170
rect -43 114 43 170
rect 99 114 185 170
rect 241 114 327 170
rect 383 114 469 170
rect 525 114 611 170
rect 667 114 753 170
rect 809 114 895 170
rect 951 114 1037 170
rect 1093 114 1179 170
rect 1235 114 1321 170
rect 1377 114 1463 170
rect 1519 114 1605 170
rect 1661 114 1747 170
rect 1803 114 1889 170
rect 1945 114 2031 170
rect 2087 114 2173 170
rect 2229 114 2315 170
rect 2371 114 2457 170
rect 2513 114 2599 170
rect 2655 114 2741 170
rect 2797 114 2883 170
rect 2939 114 3025 170
rect 3081 114 3167 170
rect 3223 114 3309 170
rect 3365 114 3451 170
rect 3507 114 3593 170
rect 3649 114 3735 170
rect 3791 114 3877 170
rect 3933 114 4019 170
rect 4075 114 4161 170
rect 4217 114 4303 170
rect 4359 114 4445 170
rect 4501 114 4587 170
rect 4643 114 4729 170
rect 4785 114 4871 170
rect 4927 114 5013 170
rect 5069 114 5155 170
rect 5211 114 5297 170
rect 5353 114 5439 170
rect 5495 114 5581 170
rect 5637 114 5723 170
rect 5779 114 5865 170
rect 5921 114 6007 170
rect 6063 114 6149 170
rect 6205 114 6291 170
rect 6347 114 6433 170
rect 6489 114 6575 170
rect 6631 114 6717 170
rect 6773 114 6859 170
rect 6915 114 7001 170
rect 7057 114 7143 170
rect 7199 114 7285 170
rect 7341 114 7351 170
rect -7351 28 7351 114
rect -7351 -28 -7341 28
rect -7285 -28 -7199 28
rect -7143 -28 -7057 28
rect -7001 -28 -6915 28
rect -6859 -28 -6773 28
rect -6717 -28 -6631 28
rect -6575 -28 -6489 28
rect -6433 -28 -6347 28
rect -6291 -28 -6205 28
rect -6149 -28 -6063 28
rect -6007 -28 -5921 28
rect -5865 -28 -5779 28
rect -5723 -28 -5637 28
rect -5581 -28 -5495 28
rect -5439 -28 -5353 28
rect -5297 -28 -5211 28
rect -5155 -28 -5069 28
rect -5013 -28 -4927 28
rect -4871 -28 -4785 28
rect -4729 -28 -4643 28
rect -4587 -28 -4501 28
rect -4445 -28 -4359 28
rect -4303 -28 -4217 28
rect -4161 -28 -4075 28
rect -4019 -28 -3933 28
rect -3877 -28 -3791 28
rect -3735 -28 -3649 28
rect -3593 -28 -3507 28
rect -3451 -28 -3365 28
rect -3309 -28 -3223 28
rect -3167 -28 -3081 28
rect -3025 -28 -2939 28
rect -2883 -28 -2797 28
rect -2741 -28 -2655 28
rect -2599 -28 -2513 28
rect -2457 -28 -2371 28
rect -2315 -28 -2229 28
rect -2173 -28 -2087 28
rect -2031 -28 -1945 28
rect -1889 -28 -1803 28
rect -1747 -28 -1661 28
rect -1605 -28 -1519 28
rect -1463 -28 -1377 28
rect -1321 -28 -1235 28
rect -1179 -28 -1093 28
rect -1037 -28 -951 28
rect -895 -28 -809 28
rect -753 -28 -667 28
rect -611 -28 -525 28
rect -469 -28 -383 28
rect -327 -28 -241 28
rect -185 -28 -99 28
rect -43 -28 43 28
rect 99 -28 185 28
rect 241 -28 327 28
rect 383 -28 469 28
rect 525 -28 611 28
rect 667 -28 753 28
rect 809 -28 895 28
rect 951 -28 1037 28
rect 1093 -28 1179 28
rect 1235 -28 1321 28
rect 1377 -28 1463 28
rect 1519 -28 1605 28
rect 1661 -28 1747 28
rect 1803 -28 1889 28
rect 1945 -28 2031 28
rect 2087 -28 2173 28
rect 2229 -28 2315 28
rect 2371 -28 2457 28
rect 2513 -28 2599 28
rect 2655 -28 2741 28
rect 2797 -28 2883 28
rect 2939 -28 3025 28
rect 3081 -28 3167 28
rect 3223 -28 3309 28
rect 3365 -28 3451 28
rect 3507 -28 3593 28
rect 3649 -28 3735 28
rect 3791 -28 3877 28
rect 3933 -28 4019 28
rect 4075 -28 4161 28
rect 4217 -28 4303 28
rect 4359 -28 4445 28
rect 4501 -28 4587 28
rect 4643 -28 4729 28
rect 4785 -28 4871 28
rect 4927 -28 5013 28
rect 5069 -28 5155 28
rect 5211 -28 5297 28
rect 5353 -28 5439 28
rect 5495 -28 5581 28
rect 5637 -28 5723 28
rect 5779 -28 5865 28
rect 5921 -28 6007 28
rect 6063 -28 6149 28
rect 6205 -28 6291 28
rect 6347 -28 6433 28
rect 6489 -28 6575 28
rect 6631 -28 6717 28
rect 6773 -28 6859 28
rect 6915 -28 7001 28
rect 7057 -28 7143 28
rect 7199 -28 7285 28
rect 7341 -28 7351 28
rect -7351 -114 7351 -28
rect -7351 -170 -7341 -114
rect -7285 -170 -7199 -114
rect -7143 -170 -7057 -114
rect -7001 -170 -6915 -114
rect -6859 -170 -6773 -114
rect -6717 -170 -6631 -114
rect -6575 -170 -6489 -114
rect -6433 -170 -6347 -114
rect -6291 -170 -6205 -114
rect -6149 -170 -6063 -114
rect -6007 -170 -5921 -114
rect -5865 -170 -5779 -114
rect -5723 -170 -5637 -114
rect -5581 -170 -5495 -114
rect -5439 -170 -5353 -114
rect -5297 -170 -5211 -114
rect -5155 -170 -5069 -114
rect -5013 -170 -4927 -114
rect -4871 -170 -4785 -114
rect -4729 -170 -4643 -114
rect -4587 -170 -4501 -114
rect -4445 -170 -4359 -114
rect -4303 -170 -4217 -114
rect -4161 -170 -4075 -114
rect -4019 -170 -3933 -114
rect -3877 -170 -3791 -114
rect -3735 -170 -3649 -114
rect -3593 -170 -3507 -114
rect -3451 -170 -3365 -114
rect -3309 -170 -3223 -114
rect -3167 -170 -3081 -114
rect -3025 -170 -2939 -114
rect -2883 -170 -2797 -114
rect -2741 -170 -2655 -114
rect -2599 -170 -2513 -114
rect -2457 -170 -2371 -114
rect -2315 -170 -2229 -114
rect -2173 -170 -2087 -114
rect -2031 -170 -1945 -114
rect -1889 -170 -1803 -114
rect -1747 -170 -1661 -114
rect -1605 -170 -1519 -114
rect -1463 -170 -1377 -114
rect -1321 -170 -1235 -114
rect -1179 -170 -1093 -114
rect -1037 -170 -951 -114
rect -895 -170 -809 -114
rect -753 -170 -667 -114
rect -611 -170 -525 -114
rect -469 -170 -383 -114
rect -327 -170 -241 -114
rect -185 -170 -99 -114
rect -43 -170 43 -114
rect 99 -170 185 -114
rect 241 -170 327 -114
rect 383 -170 469 -114
rect 525 -170 611 -114
rect 667 -170 753 -114
rect 809 -170 895 -114
rect 951 -170 1037 -114
rect 1093 -170 1179 -114
rect 1235 -170 1321 -114
rect 1377 -170 1463 -114
rect 1519 -170 1605 -114
rect 1661 -170 1747 -114
rect 1803 -170 1889 -114
rect 1945 -170 2031 -114
rect 2087 -170 2173 -114
rect 2229 -170 2315 -114
rect 2371 -170 2457 -114
rect 2513 -170 2599 -114
rect 2655 -170 2741 -114
rect 2797 -170 2883 -114
rect 2939 -170 3025 -114
rect 3081 -170 3167 -114
rect 3223 -170 3309 -114
rect 3365 -170 3451 -114
rect 3507 -170 3593 -114
rect 3649 -170 3735 -114
rect 3791 -170 3877 -114
rect 3933 -170 4019 -114
rect 4075 -170 4161 -114
rect 4217 -170 4303 -114
rect 4359 -170 4445 -114
rect 4501 -170 4587 -114
rect 4643 -170 4729 -114
rect 4785 -170 4871 -114
rect 4927 -170 5013 -114
rect 5069 -170 5155 -114
rect 5211 -170 5297 -114
rect 5353 -170 5439 -114
rect 5495 -170 5581 -114
rect 5637 -170 5723 -114
rect 5779 -170 5865 -114
rect 5921 -170 6007 -114
rect 6063 -170 6149 -114
rect 6205 -170 6291 -114
rect 6347 -170 6433 -114
rect 6489 -170 6575 -114
rect 6631 -170 6717 -114
rect 6773 -170 6859 -114
rect 6915 -170 7001 -114
rect 7057 -170 7143 -114
rect 7199 -170 7285 -114
rect 7341 -170 7351 -114
rect -7351 -256 7351 -170
rect -7351 -312 -7341 -256
rect -7285 -312 -7199 -256
rect -7143 -312 -7057 -256
rect -7001 -312 -6915 -256
rect -6859 -312 -6773 -256
rect -6717 -312 -6631 -256
rect -6575 -312 -6489 -256
rect -6433 -312 -6347 -256
rect -6291 -312 -6205 -256
rect -6149 -312 -6063 -256
rect -6007 -312 -5921 -256
rect -5865 -312 -5779 -256
rect -5723 -312 -5637 -256
rect -5581 -312 -5495 -256
rect -5439 -312 -5353 -256
rect -5297 -312 -5211 -256
rect -5155 -312 -5069 -256
rect -5013 -312 -4927 -256
rect -4871 -312 -4785 -256
rect -4729 -312 -4643 -256
rect -4587 -312 -4501 -256
rect -4445 -312 -4359 -256
rect -4303 -312 -4217 -256
rect -4161 -312 -4075 -256
rect -4019 -312 -3933 -256
rect -3877 -312 -3791 -256
rect -3735 -312 -3649 -256
rect -3593 -312 -3507 -256
rect -3451 -312 -3365 -256
rect -3309 -312 -3223 -256
rect -3167 -312 -3081 -256
rect -3025 -312 -2939 -256
rect -2883 -312 -2797 -256
rect -2741 -312 -2655 -256
rect -2599 -312 -2513 -256
rect -2457 -312 -2371 -256
rect -2315 -312 -2229 -256
rect -2173 -312 -2087 -256
rect -2031 -312 -1945 -256
rect -1889 -312 -1803 -256
rect -1747 -312 -1661 -256
rect -1605 -312 -1519 -256
rect -1463 -312 -1377 -256
rect -1321 -312 -1235 -256
rect -1179 -312 -1093 -256
rect -1037 -312 -951 -256
rect -895 -312 -809 -256
rect -753 -312 -667 -256
rect -611 -312 -525 -256
rect -469 -312 -383 -256
rect -327 -312 -241 -256
rect -185 -312 -99 -256
rect -43 -312 43 -256
rect 99 -312 185 -256
rect 241 -312 327 -256
rect 383 -312 469 -256
rect 525 -312 611 -256
rect 667 -312 753 -256
rect 809 -312 895 -256
rect 951 -312 1037 -256
rect 1093 -312 1179 -256
rect 1235 -312 1321 -256
rect 1377 -312 1463 -256
rect 1519 -312 1605 -256
rect 1661 -312 1747 -256
rect 1803 -312 1889 -256
rect 1945 -312 2031 -256
rect 2087 -312 2173 -256
rect 2229 -312 2315 -256
rect 2371 -312 2457 -256
rect 2513 -312 2599 -256
rect 2655 -312 2741 -256
rect 2797 -312 2883 -256
rect 2939 -312 3025 -256
rect 3081 -312 3167 -256
rect 3223 -312 3309 -256
rect 3365 -312 3451 -256
rect 3507 -312 3593 -256
rect 3649 -312 3735 -256
rect 3791 -312 3877 -256
rect 3933 -312 4019 -256
rect 4075 -312 4161 -256
rect 4217 -312 4303 -256
rect 4359 -312 4445 -256
rect 4501 -312 4587 -256
rect 4643 -312 4729 -256
rect 4785 -312 4871 -256
rect 4927 -312 5013 -256
rect 5069 -312 5155 -256
rect 5211 -312 5297 -256
rect 5353 -312 5439 -256
rect 5495 -312 5581 -256
rect 5637 -312 5723 -256
rect 5779 -312 5865 -256
rect 5921 -312 6007 -256
rect 6063 -312 6149 -256
rect 6205 -312 6291 -256
rect 6347 -312 6433 -256
rect 6489 -312 6575 -256
rect 6631 -312 6717 -256
rect 6773 -312 6859 -256
rect 6915 -312 7001 -256
rect 7057 -312 7143 -256
rect 7199 -312 7285 -256
rect 7341 -312 7351 -256
rect -7351 -398 7351 -312
rect -7351 -454 -7341 -398
rect -7285 -454 -7199 -398
rect -7143 -454 -7057 -398
rect -7001 -454 -6915 -398
rect -6859 -454 -6773 -398
rect -6717 -454 -6631 -398
rect -6575 -454 -6489 -398
rect -6433 -454 -6347 -398
rect -6291 -454 -6205 -398
rect -6149 -454 -6063 -398
rect -6007 -454 -5921 -398
rect -5865 -454 -5779 -398
rect -5723 -454 -5637 -398
rect -5581 -454 -5495 -398
rect -5439 -454 -5353 -398
rect -5297 -454 -5211 -398
rect -5155 -454 -5069 -398
rect -5013 -454 -4927 -398
rect -4871 -454 -4785 -398
rect -4729 -454 -4643 -398
rect -4587 -454 -4501 -398
rect -4445 -454 -4359 -398
rect -4303 -454 -4217 -398
rect -4161 -454 -4075 -398
rect -4019 -454 -3933 -398
rect -3877 -454 -3791 -398
rect -3735 -454 -3649 -398
rect -3593 -454 -3507 -398
rect -3451 -454 -3365 -398
rect -3309 -454 -3223 -398
rect -3167 -454 -3081 -398
rect -3025 -454 -2939 -398
rect -2883 -454 -2797 -398
rect -2741 -454 -2655 -398
rect -2599 -454 -2513 -398
rect -2457 -454 -2371 -398
rect -2315 -454 -2229 -398
rect -2173 -454 -2087 -398
rect -2031 -454 -1945 -398
rect -1889 -454 -1803 -398
rect -1747 -454 -1661 -398
rect -1605 -454 -1519 -398
rect -1463 -454 -1377 -398
rect -1321 -454 -1235 -398
rect -1179 -454 -1093 -398
rect -1037 -454 -951 -398
rect -895 -454 -809 -398
rect -753 -454 -667 -398
rect -611 -454 -525 -398
rect -469 -454 -383 -398
rect -327 -454 -241 -398
rect -185 -454 -99 -398
rect -43 -454 43 -398
rect 99 -454 185 -398
rect 241 -454 327 -398
rect 383 -454 469 -398
rect 525 -454 611 -398
rect 667 -454 753 -398
rect 809 -454 895 -398
rect 951 -454 1037 -398
rect 1093 -454 1179 -398
rect 1235 -454 1321 -398
rect 1377 -454 1463 -398
rect 1519 -454 1605 -398
rect 1661 -454 1747 -398
rect 1803 -454 1889 -398
rect 1945 -454 2031 -398
rect 2087 -454 2173 -398
rect 2229 -454 2315 -398
rect 2371 -454 2457 -398
rect 2513 -454 2599 -398
rect 2655 -454 2741 -398
rect 2797 -454 2883 -398
rect 2939 -454 3025 -398
rect 3081 -454 3167 -398
rect 3223 -454 3309 -398
rect 3365 -454 3451 -398
rect 3507 -454 3593 -398
rect 3649 -454 3735 -398
rect 3791 -454 3877 -398
rect 3933 -454 4019 -398
rect 4075 -454 4161 -398
rect 4217 -454 4303 -398
rect 4359 -454 4445 -398
rect 4501 -454 4587 -398
rect 4643 -454 4729 -398
rect 4785 -454 4871 -398
rect 4927 -454 5013 -398
rect 5069 -454 5155 -398
rect 5211 -454 5297 -398
rect 5353 -454 5439 -398
rect 5495 -454 5581 -398
rect 5637 -454 5723 -398
rect 5779 -454 5865 -398
rect 5921 -454 6007 -398
rect 6063 -454 6149 -398
rect 6205 -454 6291 -398
rect 6347 -454 6433 -398
rect 6489 -454 6575 -398
rect 6631 -454 6717 -398
rect 6773 -454 6859 -398
rect 6915 -454 7001 -398
rect 7057 -454 7143 -398
rect 7199 -454 7285 -398
rect 7341 -454 7351 -398
rect -7351 -540 7351 -454
rect -7351 -596 -7341 -540
rect -7285 -596 -7199 -540
rect -7143 -596 -7057 -540
rect -7001 -596 -6915 -540
rect -6859 -596 -6773 -540
rect -6717 -596 -6631 -540
rect -6575 -596 -6489 -540
rect -6433 -596 -6347 -540
rect -6291 -596 -6205 -540
rect -6149 -596 -6063 -540
rect -6007 -596 -5921 -540
rect -5865 -596 -5779 -540
rect -5723 -596 -5637 -540
rect -5581 -596 -5495 -540
rect -5439 -596 -5353 -540
rect -5297 -596 -5211 -540
rect -5155 -596 -5069 -540
rect -5013 -596 -4927 -540
rect -4871 -596 -4785 -540
rect -4729 -596 -4643 -540
rect -4587 -596 -4501 -540
rect -4445 -596 -4359 -540
rect -4303 -596 -4217 -540
rect -4161 -596 -4075 -540
rect -4019 -596 -3933 -540
rect -3877 -596 -3791 -540
rect -3735 -596 -3649 -540
rect -3593 -596 -3507 -540
rect -3451 -596 -3365 -540
rect -3309 -596 -3223 -540
rect -3167 -596 -3081 -540
rect -3025 -596 -2939 -540
rect -2883 -596 -2797 -540
rect -2741 -596 -2655 -540
rect -2599 -596 -2513 -540
rect -2457 -596 -2371 -540
rect -2315 -596 -2229 -540
rect -2173 -596 -2087 -540
rect -2031 -596 -1945 -540
rect -1889 -596 -1803 -540
rect -1747 -596 -1661 -540
rect -1605 -596 -1519 -540
rect -1463 -596 -1377 -540
rect -1321 -596 -1235 -540
rect -1179 -596 -1093 -540
rect -1037 -596 -951 -540
rect -895 -596 -809 -540
rect -753 -596 -667 -540
rect -611 -596 -525 -540
rect -469 -596 -383 -540
rect -327 -596 -241 -540
rect -185 -596 -99 -540
rect -43 -596 43 -540
rect 99 -596 185 -540
rect 241 -596 327 -540
rect 383 -596 469 -540
rect 525 -596 611 -540
rect 667 -596 753 -540
rect 809 -596 895 -540
rect 951 -596 1037 -540
rect 1093 -596 1179 -540
rect 1235 -596 1321 -540
rect 1377 -596 1463 -540
rect 1519 -596 1605 -540
rect 1661 -596 1747 -540
rect 1803 -596 1889 -540
rect 1945 -596 2031 -540
rect 2087 -596 2173 -540
rect 2229 -596 2315 -540
rect 2371 -596 2457 -540
rect 2513 -596 2599 -540
rect 2655 -596 2741 -540
rect 2797 -596 2883 -540
rect 2939 -596 3025 -540
rect 3081 -596 3167 -540
rect 3223 -596 3309 -540
rect 3365 -596 3451 -540
rect 3507 -596 3593 -540
rect 3649 -596 3735 -540
rect 3791 -596 3877 -540
rect 3933 -596 4019 -540
rect 4075 -596 4161 -540
rect 4217 -596 4303 -540
rect 4359 -596 4445 -540
rect 4501 -596 4587 -540
rect 4643 -596 4729 -540
rect 4785 -596 4871 -540
rect 4927 -596 5013 -540
rect 5069 -596 5155 -540
rect 5211 -596 5297 -540
rect 5353 -596 5439 -540
rect 5495 -596 5581 -540
rect 5637 -596 5723 -540
rect 5779 -596 5865 -540
rect 5921 -596 6007 -540
rect 6063 -596 6149 -540
rect 6205 -596 6291 -540
rect 6347 -596 6433 -540
rect 6489 -596 6575 -540
rect 6631 -596 6717 -540
rect 6773 -596 6859 -540
rect 6915 -596 7001 -540
rect 7057 -596 7143 -540
rect 7199 -596 7285 -540
rect 7341 -596 7351 -540
rect -7351 -682 7351 -596
rect -7351 -738 -7341 -682
rect -7285 -738 -7199 -682
rect -7143 -738 -7057 -682
rect -7001 -738 -6915 -682
rect -6859 -738 -6773 -682
rect -6717 -738 -6631 -682
rect -6575 -738 -6489 -682
rect -6433 -738 -6347 -682
rect -6291 -738 -6205 -682
rect -6149 -738 -6063 -682
rect -6007 -738 -5921 -682
rect -5865 -738 -5779 -682
rect -5723 -738 -5637 -682
rect -5581 -738 -5495 -682
rect -5439 -738 -5353 -682
rect -5297 -738 -5211 -682
rect -5155 -738 -5069 -682
rect -5013 -738 -4927 -682
rect -4871 -738 -4785 -682
rect -4729 -738 -4643 -682
rect -4587 -738 -4501 -682
rect -4445 -738 -4359 -682
rect -4303 -738 -4217 -682
rect -4161 -738 -4075 -682
rect -4019 -738 -3933 -682
rect -3877 -738 -3791 -682
rect -3735 -738 -3649 -682
rect -3593 -738 -3507 -682
rect -3451 -738 -3365 -682
rect -3309 -738 -3223 -682
rect -3167 -738 -3081 -682
rect -3025 -738 -2939 -682
rect -2883 -738 -2797 -682
rect -2741 -738 -2655 -682
rect -2599 -738 -2513 -682
rect -2457 -738 -2371 -682
rect -2315 -738 -2229 -682
rect -2173 -738 -2087 -682
rect -2031 -738 -1945 -682
rect -1889 -738 -1803 -682
rect -1747 -738 -1661 -682
rect -1605 -738 -1519 -682
rect -1463 -738 -1377 -682
rect -1321 -738 -1235 -682
rect -1179 -738 -1093 -682
rect -1037 -738 -951 -682
rect -895 -738 -809 -682
rect -753 -738 -667 -682
rect -611 -738 -525 -682
rect -469 -738 -383 -682
rect -327 -738 -241 -682
rect -185 -738 -99 -682
rect -43 -738 43 -682
rect 99 -738 185 -682
rect 241 -738 327 -682
rect 383 -738 469 -682
rect 525 -738 611 -682
rect 667 -738 753 -682
rect 809 -738 895 -682
rect 951 -738 1037 -682
rect 1093 -738 1179 -682
rect 1235 -738 1321 -682
rect 1377 -738 1463 -682
rect 1519 -738 1605 -682
rect 1661 -738 1747 -682
rect 1803 -738 1889 -682
rect 1945 -738 2031 -682
rect 2087 -738 2173 -682
rect 2229 -738 2315 -682
rect 2371 -738 2457 -682
rect 2513 -738 2599 -682
rect 2655 -738 2741 -682
rect 2797 -738 2883 -682
rect 2939 -738 3025 -682
rect 3081 -738 3167 -682
rect 3223 -738 3309 -682
rect 3365 -738 3451 -682
rect 3507 -738 3593 -682
rect 3649 -738 3735 -682
rect 3791 -738 3877 -682
rect 3933 -738 4019 -682
rect 4075 -738 4161 -682
rect 4217 -738 4303 -682
rect 4359 -738 4445 -682
rect 4501 -738 4587 -682
rect 4643 -738 4729 -682
rect 4785 -738 4871 -682
rect 4927 -738 5013 -682
rect 5069 -738 5155 -682
rect 5211 -738 5297 -682
rect 5353 -738 5439 -682
rect 5495 -738 5581 -682
rect 5637 -738 5723 -682
rect 5779 -738 5865 -682
rect 5921 -738 6007 -682
rect 6063 -738 6149 -682
rect 6205 -738 6291 -682
rect 6347 -738 6433 -682
rect 6489 -738 6575 -682
rect 6631 -738 6717 -682
rect 6773 -738 6859 -682
rect 6915 -738 7001 -682
rect 7057 -738 7143 -682
rect 7199 -738 7285 -682
rect 7341 -738 7351 -682
rect -7351 -824 7351 -738
rect -7351 -880 -7341 -824
rect -7285 -880 -7199 -824
rect -7143 -880 -7057 -824
rect -7001 -880 -6915 -824
rect -6859 -880 -6773 -824
rect -6717 -880 -6631 -824
rect -6575 -880 -6489 -824
rect -6433 -880 -6347 -824
rect -6291 -880 -6205 -824
rect -6149 -880 -6063 -824
rect -6007 -880 -5921 -824
rect -5865 -880 -5779 -824
rect -5723 -880 -5637 -824
rect -5581 -880 -5495 -824
rect -5439 -880 -5353 -824
rect -5297 -880 -5211 -824
rect -5155 -880 -5069 -824
rect -5013 -880 -4927 -824
rect -4871 -880 -4785 -824
rect -4729 -880 -4643 -824
rect -4587 -880 -4501 -824
rect -4445 -880 -4359 -824
rect -4303 -880 -4217 -824
rect -4161 -880 -4075 -824
rect -4019 -880 -3933 -824
rect -3877 -880 -3791 -824
rect -3735 -880 -3649 -824
rect -3593 -880 -3507 -824
rect -3451 -880 -3365 -824
rect -3309 -880 -3223 -824
rect -3167 -880 -3081 -824
rect -3025 -880 -2939 -824
rect -2883 -880 -2797 -824
rect -2741 -880 -2655 -824
rect -2599 -880 -2513 -824
rect -2457 -880 -2371 -824
rect -2315 -880 -2229 -824
rect -2173 -880 -2087 -824
rect -2031 -880 -1945 -824
rect -1889 -880 -1803 -824
rect -1747 -880 -1661 -824
rect -1605 -880 -1519 -824
rect -1463 -880 -1377 -824
rect -1321 -880 -1235 -824
rect -1179 -880 -1093 -824
rect -1037 -880 -951 -824
rect -895 -880 -809 -824
rect -753 -880 -667 -824
rect -611 -880 -525 -824
rect -469 -880 -383 -824
rect -327 -880 -241 -824
rect -185 -880 -99 -824
rect -43 -880 43 -824
rect 99 -880 185 -824
rect 241 -880 327 -824
rect 383 -880 469 -824
rect 525 -880 611 -824
rect 667 -880 753 -824
rect 809 -880 895 -824
rect 951 -880 1037 -824
rect 1093 -880 1179 -824
rect 1235 -880 1321 -824
rect 1377 -880 1463 -824
rect 1519 -880 1605 -824
rect 1661 -880 1747 -824
rect 1803 -880 1889 -824
rect 1945 -880 2031 -824
rect 2087 -880 2173 -824
rect 2229 -880 2315 -824
rect 2371 -880 2457 -824
rect 2513 -880 2599 -824
rect 2655 -880 2741 -824
rect 2797 -880 2883 -824
rect 2939 -880 3025 -824
rect 3081 -880 3167 -824
rect 3223 -880 3309 -824
rect 3365 -880 3451 -824
rect 3507 -880 3593 -824
rect 3649 -880 3735 -824
rect 3791 -880 3877 -824
rect 3933 -880 4019 -824
rect 4075 -880 4161 -824
rect 4217 -880 4303 -824
rect 4359 -880 4445 -824
rect 4501 -880 4587 -824
rect 4643 -880 4729 -824
rect 4785 -880 4871 -824
rect 4927 -880 5013 -824
rect 5069 -880 5155 -824
rect 5211 -880 5297 -824
rect 5353 -880 5439 -824
rect 5495 -880 5581 -824
rect 5637 -880 5723 -824
rect 5779 -880 5865 -824
rect 5921 -880 6007 -824
rect 6063 -880 6149 -824
rect 6205 -880 6291 -824
rect 6347 -880 6433 -824
rect 6489 -880 6575 -824
rect 6631 -880 6717 -824
rect 6773 -880 6859 -824
rect 6915 -880 7001 -824
rect 7057 -880 7143 -824
rect 7199 -880 7285 -824
rect 7341 -880 7351 -824
rect -7351 -966 7351 -880
rect -7351 -1022 -7341 -966
rect -7285 -1022 -7199 -966
rect -7143 -1022 -7057 -966
rect -7001 -1022 -6915 -966
rect -6859 -1022 -6773 -966
rect -6717 -1022 -6631 -966
rect -6575 -1022 -6489 -966
rect -6433 -1022 -6347 -966
rect -6291 -1022 -6205 -966
rect -6149 -1022 -6063 -966
rect -6007 -1022 -5921 -966
rect -5865 -1022 -5779 -966
rect -5723 -1022 -5637 -966
rect -5581 -1022 -5495 -966
rect -5439 -1022 -5353 -966
rect -5297 -1022 -5211 -966
rect -5155 -1022 -5069 -966
rect -5013 -1022 -4927 -966
rect -4871 -1022 -4785 -966
rect -4729 -1022 -4643 -966
rect -4587 -1022 -4501 -966
rect -4445 -1022 -4359 -966
rect -4303 -1022 -4217 -966
rect -4161 -1022 -4075 -966
rect -4019 -1022 -3933 -966
rect -3877 -1022 -3791 -966
rect -3735 -1022 -3649 -966
rect -3593 -1022 -3507 -966
rect -3451 -1022 -3365 -966
rect -3309 -1022 -3223 -966
rect -3167 -1022 -3081 -966
rect -3025 -1022 -2939 -966
rect -2883 -1022 -2797 -966
rect -2741 -1022 -2655 -966
rect -2599 -1022 -2513 -966
rect -2457 -1022 -2371 -966
rect -2315 -1022 -2229 -966
rect -2173 -1022 -2087 -966
rect -2031 -1022 -1945 -966
rect -1889 -1022 -1803 -966
rect -1747 -1022 -1661 -966
rect -1605 -1022 -1519 -966
rect -1463 -1022 -1377 -966
rect -1321 -1022 -1235 -966
rect -1179 -1022 -1093 -966
rect -1037 -1022 -951 -966
rect -895 -1022 -809 -966
rect -753 -1022 -667 -966
rect -611 -1022 -525 -966
rect -469 -1022 -383 -966
rect -327 -1022 -241 -966
rect -185 -1022 -99 -966
rect -43 -1022 43 -966
rect 99 -1022 185 -966
rect 241 -1022 327 -966
rect 383 -1022 469 -966
rect 525 -1022 611 -966
rect 667 -1022 753 -966
rect 809 -1022 895 -966
rect 951 -1022 1037 -966
rect 1093 -1022 1179 -966
rect 1235 -1022 1321 -966
rect 1377 -1022 1463 -966
rect 1519 -1022 1605 -966
rect 1661 -1022 1747 -966
rect 1803 -1022 1889 -966
rect 1945 -1022 2031 -966
rect 2087 -1022 2173 -966
rect 2229 -1022 2315 -966
rect 2371 -1022 2457 -966
rect 2513 -1022 2599 -966
rect 2655 -1022 2741 -966
rect 2797 -1022 2883 -966
rect 2939 -1022 3025 -966
rect 3081 -1022 3167 -966
rect 3223 -1022 3309 -966
rect 3365 -1022 3451 -966
rect 3507 -1022 3593 -966
rect 3649 -1022 3735 -966
rect 3791 -1022 3877 -966
rect 3933 -1022 4019 -966
rect 4075 -1022 4161 -966
rect 4217 -1022 4303 -966
rect 4359 -1022 4445 -966
rect 4501 -1022 4587 -966
rect 4643 -1022 4729 -966
rect 4785 -1022 4871 -966
rect 4927 -1022 5013 -966
rect 5069 -1022 5155 -966
rect 5211 -1022 5297 -966
rect 5353 -1022 5439 -966
rect 5495 -1022 5581 -966
rect 5637 -1022 5723 -966
rect 5779 -1022 5865 -966
rect 5921 -1022 6007 -966
rect 6063 -1022 6149 -966
rect 6205 -1022 6291 -966
rect 6347 -1022 6433 -966
rect 6489 -1022 6575 -966
rect 6631 -1022 6717 -966
rect 6773 -1022 6859 -966
rect 6915 -1022 7001 -966
rect 7057 -1022 7143 -966
rect 7199 -1022 7285 -966
rect 7341 -1022 7351 -966
rect -7351 -1108 7351 -1022
rect -7351 -1164 -7341 -1108
rect -7285 -1164 -7199 -1108
rect -7143 -1164 -7057 -1108
rect -7001 -1164 -6915 -1108
rect -6859 -1164 -6773 -1108
rect -6717 -1164 -6631 -1108
rect -6575 -1164 -6489 -1108
rect -6433 -1164 -6347 -1108
rect -6291 -1164 -6205 -1108
rect -6149 -1164 -6063 -1108
rect -6007 -1164 -5921 -1108
rect -5865 -1164 -5779 -1108
rect -5723 -1164 -5637 -1108
rect -5581 -1164 -5495 -1108
rect -5439 -1164 -5353 -1108
rect -5297 -1164 -5211 -1108
rect -5155 -1164 -5069 -1108
rect -5013 -1164 -4927 -1108
rect -4871 -1164 -4785 -1108
rect -4729 -1164 -4643 -1108
rect -4587 -1164 -4501 -1108
rect -4445 -1164 -4359 -1108
rect -4303 -1164 -4217 -1108
rect -4161 -1164 -4075 -1108
rect -4019 -1164 -3933 -1108
rect -3877 -1164 -3791 -1108
rect -3735 -1164 -3649 -1108
rect -3593 -1164 -3507 -1108
rect -3451 -1164 -3365 -1108
rect -3309 -1164 -3223 -1108
rect -3167 -1164 -3081 -1108
rect -3025 -1164 -2939 -1108
rect -2883 -1164 -2797 -1108
rect -2741 -1164 -2655 -1108
rect -2599 -1164 -2513 -1108
rect -2457 -1164 -2371 -1108
rect -2315 -1164 -2229 -1108
rect -2173 -1164 -2087 -1108
rect -2031 -1164 -1945 -1108
rect -1889 -1164 -1803 -1108
rect -1747 -1164 -1661 -1108
rect -1605 -1164 -1519 -1108
rect -1463 -1164 -1377 -1108
rect -1321 -1164 -1235 -1108
rect -1179 -1164 -1093 -1108
rect -1037 -1164 -951 -1108
rect -895 -1164 -809 -1108
rect -753 -1164 -667 -1108
rect -611 -1164 -525 -1108
rect -469 -1164 -383 -1108
rect -327 -1164 -241 -1108
rect -185 -1164 -99 -1108
rect -43 -1164 43 -1108
rect 99 -1164 185 -1108
rect 241 -1164 327 -1108
rect 383 -1164 469 -1108
rect 525 -1164 611 -1108
rect 667 -1164 753 -1108
rect 809 -1164 895 -1108
rect 951 -1164 1037 -1108
rect 1093 -1164 1179 -1108
rect 1235 -1164 1321 -1108
rect 1377 -1164 1463 -1108
rect 1519 -1164 1605 -1108
rect 1661 -1164 1747 -1108
rect 1803 -1164 1889 -1108
rect 1945 -1164 2031 -1108
rect 2087 -1164 2173 -1108
rect 2229 -1164 2315 -1108
rect 2371 -1164 2457 -1108
rect 2513 -1164 2599 -1108
rect 2655 -1164 2741 -1108
rect 2797 -1164 2883 -1108
rect 2939 -1164 3025 -1108
rect 3081 -1164 3167 -1108
rect 3223 -1164 3309 -1108
rect 3365 -1164 3451 -1108
rect 3507 -1164 3593 -1108
rect 3649 -1164 3735 -1108
rect 3791 -1164 3877 -1108
rect 3933 -1164 4019 -1108
rect 4075 -1164 4161 -1108
rect 4217 -1164 4303 -1108
rect 4359 -1164 4445 -1108
rect 4501 -1164 4587 -1108
rect 4643 -1164 4729 -1108
rect 4785 -1164 4871 -1108
rect 4927 -1164 5013 -1108
rect 5069 -1164 5155 -1108
rect 5211 -1164 5297 -1108
rect 5353 -1164 5439 -1108
rect 5495 -1164 5581 -1108
rect 5637 -1164 5723 -1108
rect 5779 -1164 5865 -1108
rect 5921 -1164 6007 -1108
rect 6063 -1164 6149 -1108
rect 6205 -1164 6291 -1108
rect 6347 -1164 6433 -1108
rect 6489 -1164 6575 -1108
rect 6631 -1164 6717 -1108
rect 6773 -1164 6859 -1108
rect 6915 -1164 7001 -1108
rect 7057 -1164 7143 -1108
rect 7199 -1164 7285 -1108
rect 7341 -1164 7351 -1108
rect -7351 -1250 7351 -1164
rect -7351 -1306 -7341 -1250
rect -7285 -1306 -7199 -1250
rect -7143 -1306 -7057 -1250
rect -7001 -1306 -6915 -1250
rect -6859 -1306 -6773 -1250
rect -6717 -1306 -6631 -1250
rect -6575 -1306 -6489 -1250
rect -6433 -1306 -6347 -1250
rect -6291 -1306 -6205 -1250
rect -6149 -1306 -6063 -1250
rect -6007 -1306 -5921 -1250
rect -5865 -1306 -5779 -1250
rect -5723 -1306 -5637 -1250
rect -5581 -1306 -5495 -1250
rect -5439 -1306 -5353 -1250
rect -5297 -1306 -5211 -1250
rect -5155 -1306 -5069 -1250
rect -5013 -1306 -4927 -1250
rect -4871 -1306 -4785 -1250
rect -4729 -1306 -4643 -1250
rect -4587 -1306 -4501 -1250
rect -4445 -1306 -4359 -1250
rect -4303 -1306 -4217 -1250
rect -4161 -1306 -4075 -1250
rect -4019 -1306 -3933 -1250
rect -3877 -1306 -3791 -1250
rect -3735 -1306 -3649 -1250
rect -3593 -1306 -3507 -1250
rect -3451 -1306 -3365 -1250
rect -3309 -1306 -3223 -1250
rect -3167 -1306 -3081 -1250
rect -3025 -1306 -2939 -1250
rect -2883 -1306 -2797 -1250
rect -2741 -1306 -2655 -1250
rect -2599 -1306 -2513 -1250
rect -2457 -1306 -2371 -1250
rect -2315 -1306 -2229 -1250
rect -2173 -1306 -2087 -1250
rect -2031 -1306 -1945 -1250
rect -1889 -1306 -1803 -1250
rect -1747 -1306 -1661 -1250
rect -1605 -1306 -1519 -1250
rect -1463 -1306 -1377 -1250
rect -1321 -1306 -1235 -1250
rect -1179 -1306 -1093 -1250
rect -1037 -1306 -951 -1250
rect -895 -1306 -809 -1250
rect -753 -1306 -667 -1250
rect -611 -1306 -525 -1250
rect -469 -1306 -383 -1250
rect -327 -1306 -241 -1250
rect -185 -1306 -99 -1250
rect -43 -1306 43 -1250
rect 99 -1306 185 -1250
rect 241 -1306 327 -1250
rect 383 -1306 469 -1250
rect 525 -1306 611 -1250
rect 667 -1306 753 -1250
rect 809 -1306 895 -1250
rect 951 -1306 1037 -1250
rect 1093 -1306 1179 -1250
rect 1235 -1306 1321 -1250
rect 1377 -1306 1463 -1250
rect 1519 -1306 1605 -1250
rect 1661 -1306 1747 -1250
rect 1803 -1306 1889 -1250
rect 1945 -1306 2031 -1250
rect 2087 -1306 2173 -1250
rect 2229 -1306 2315 -1250
rect 2371 -1306 2457 -1250
rect 2513 -1306 2599 -1250
rect 2655 -1306 2741 -1250
rect 2797 -1306 2883 -1250
rect 2939 -1306 3025 -1250
rect 3081 -1306 3167 -1250
rect 3223 -1306 3309 -1250
rect 3365 -1306 3451 -1250
rect 3507 -1306 3593 -1250
rect 3649 -1306 3735 -1250
rect 3791 -1306 3877 -1250
rect 3933 -1306 4019 -1250
rect 4075 -1306 4161 -1250
rect 4217 -1306 4303 -1250
rect 4359 -1306 4445 -1250
rect 4501 -1306 4587 -1250
rect 4643 -1306 4729 -1250
rect 4785 -1306 4871 -1250
rect 4927 -1306 5013 -1250
rect 5069 -1306 5155 -1250
rect 5211 -1306 5297 -1250
rect 5353 -1306 5439 -1250
rect 5495 -1306 5581 -1250
rect 5637 -1306 5723 -1250
rect 5779 -1306 5865 -1250
rect 5921 -1306 6007 -1250
rect 6063 -1306 6149 -1250
rect 6205 -1306 6291 -1250
rect 6347 -1306 6433 -1250
rect 6489 -1306 6575 -1250
rect 6631 -1306 6717 -1250
rect 6773 -1306 6859 -1250
rect 6915 -1306 7001 -1250
rect 7057 -1306 7143 -1250
rect 7199 -1306 7285 -1250
rect 7341 -1306 7351 -1250
rect -7351 -1392 7351 -1306
rect -7351 -1448 -7341 -1392
rect -7285 -1448 -7199 -1392
rect -7143 -1448 -7057 -1392
rect -7001 -1448 -6915 -1392
rect -6859 -1448 -6773 -1392
rect -6717 -1448 -6631 -1392
rect -6575 -1448 -6489 -1392
rect -6433 -1448 -6347 -1392
rect -6291 -1448 -6205 -1392
rect -6149 -1448 -6063 -1392
rect -6007 -1448 -5921 -1392
rect -5865 -1448 -5779 -1392
rect -5723 -1448 -5637 -1392
rect -5581 -1448 -5495 -1392
rect -5439 -1448 -5353 -1392
rect -5297 -1448 -5211 -1392
rect -5155 -1448 -5069 -1392
rect -5013 -1448 -4927 -1392
rect -4871 -1448 -4785 -1392
rect -4729 -1448 -4643 -1392
rect -4587 -1448 -4501 -1392
rect -4445 -1448 -4359 -1392
rect -4303 -1448 -4217 -1392
rect -4161 -1448 -4075 -1392
rect -4019 -1448 -3933 -1392
rect -3877 -1448 -3791 -1392
rect -3735 -1448 -3649 -1392
rect -3593 -1448 -3507 -1392
rect -3451 -1448 -3365 -1392
rect -3309 -1448 -3223 -1392
rect -3167 -1448 -3081 -1392
rect -3025 -1448 -2939 -1392
rect -2883 -1448 -2797 -1392
rect -2741 -1448 -2655 -1392
rect -2599 -1448 -2513 -1392
rect -2457 -1448 -2371 -1392
rect -2315 -1448 -2229 -1392
rect -2173 -1448 -2087 -1392
rect -2031 -1448 -1945 -1392
rect -1889 -1448 -1803 -1392
rect -1747 -1448 -1661 -1392
rect -1605 -1448 -1519 -1392
rect -1463 -1448 -1377 -1392
rect -1321 -1448 -1235 -1392
rect -1179 -1448 -1093 -1392
rect -1037 -1448 -951 -1392
rect -895 -1448 -809 -1392
rect -753 -1448 -667 -1392
rect -611 -1448 -525 -1392
rect -469 -1448 -383 -1392
rect -327 -1448 -241 -1392
rect -185 -1448 -99 -1392
rect -43 -1448 43 -1392
rect 99 -1448 185 -1392
rect 241 -1448 327 -1392
rect 383 -1448 469 -1392
rect 525 -1448 611 -1392
rect 667 -1448 753 -1392
rect 809 -1448 895 -1392
rect 951 -1448 1037 -1392
rect 1093 -1448 1179 -1392
rect 1235 -1448 1321 -1392
rect 1377 -1448 1463 -1392
rect 1519 -1448 1605 -1392
rect 1661 -1448 1747 -1392
rect 1803 -1448 1889 -1392
rect 1945 -1448 2031 -1392
rect 2087 -1448 2173 -1392
rect 2229 -1448 2315 -1392
rect 2371 -1448 2457 -1392
rect 2513 -1448 2599 -1392
rect 2655 -1448 2741 -1392
rect 2797 -1448 2883 -1392
rect 2939 -1448 3025 -1392
rect 3081 -1448 3167 -1392
rect 3223 -1448 3309 -1392
rect 3365 -1448 3451 -1392
rect 3507 -1448 3593 -1392
rect 3649 -1448 3735 -1392
rect 3791 -1448 3877 -1392
rect 3933 -1448 4019 -1392
rect 4075 -1448 4161 -1392
rect 4217 -1448 4303 -1392
rect 4359 -1448 4445 -1392
rect 4501 -1448 4587 -1392
rect 4643 -1448 4729 -1392
rect 4785 -1448 4871 -1392
rect 4927 -1448 5013 -1392
rect 5069 -1448 5155 -1392
rect 5211 -1448 5297 -1392
rect 5353 -1448 5439 -1392
rect 5495 -1448 5581 -1392
rect 5637 -1448 5723 -1392
rect 5779 -1448 5865 -1392
rect 5921 -1448 6007 -1392
rect 6063 -1448 6149 -1392
rect 6205 -1448 6291 -1392
rect 6347 -1448 6433 -1392
rect 6489 -1448 6575 -1392
rect 6631 -1448 6717 -1392
rect 6773 -1448 6859 -1392
rect 6915 -1448 7001 -1392
rect 7057 -1448 7143 -1392
rect 7199 -1448 7285 -1392
rect 7341 -1448 7351 -1392
rect -7351 -1458 7351 -1448
<< end >>
