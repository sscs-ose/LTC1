magic
tech gf180mcuC
magscale 1 10
timestamp 1695190274
<< nwell >>
rect -284 -906 284 906
<< nsubdiff >>
rect -260 810 260 882
rect -260 -810 -188 810
rect 188 -810 260 810
rect -260 -882 260 -810
<< polysilicon >>
rect -100 709 100 722
rect -100 663 -87 709
rect 87 663 100 709
rect -100 620 100 663
rect -100 -663 100 -620
rect -100 -709 -87 -663
rect 87 -709 100 -663
rect -100 -722 100 -709
<< polycontact >>
rect -87 663 87 709
rect -87 -709 87 -663
<< ppolyres >>
rect -100 -620 100 620
<< metal1 >>
rect -98 663 -87 709
rect 87 663 98 709
rect -98 -709 -87 -663
rect 87 -709 98 -663
<< properties >>
string FIXED_BBOX -224 -846 224 846
string gencell ppolyf_u
string library gf180mcu
string parameters w 1.0 l 6.2 m 1 nx 1 wmin 0.80 lmin 1.00 rho 315 val 2.1k dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 0 grc 0 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 0
<< end >>
