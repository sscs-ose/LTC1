magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1100 -1019 1100 1019
<< metal1 >>
rect -100 13 100 19
rect -100 -13 -94 13
rect -68 -13 -40 13
rect -14 -13 14 13
rect 40 -13 68 13
rect 94 -13 100 13
rect -100 -19 100 -13
<< via1 >>
rect -94 -13 -68 13
rect -40 -13 -14 13
rect 14 -13 40 13
rect 68 -13 94 13
<< metal2 >>
rect -100 13 100 19
rect -100 -13 -94 13
rect -68 -13 -40 13
rect -14 -13 14 13
rect 40 -13 68 13
rect 94 -13 100 13
rect -100 -19 100 -13
<< end >>
