magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2011 -2000 16989 59600
<< isosubstrate >>
rect 251 53100 14727 57210
rect 2457 47106 12521 53100
rect 601 43110 14377 47106
rect 957 26495 12844 43110
rect 957 1096 14021 26495
<< psubdiff >>
rect 3094 51807 11884 52051
rect 3094 51271 3338 51807
rect 11640 51271 11884 51807
rect 3094 50873 11884 51271
rect 3094 50337 3338 50873
rect 11640 50337 11884 50873
rect 3094 49939 11884 50337
rect 3094 49403 3338 49939
rect 11640 49403 11884 49939
rect 3094 49005 11884 49403
rect 3094 48469 3338 49005
rect 11640 48469 11884 49005
rect 3094 48225 11884 48469
<< metal1 >>
rect 413 57048 499 57116
rect 14479 57048 14565 57116
rect 345 53505 617 56655
rect 14361 53505 14633 56655
rect 345 53194 14633 53505
rect 71 51622 257 52622
rect 2919 52254 3005 52622
rect 11973 52254 12059 52622
rect 3105 51818 11873 52040
rect 71 50422 257 51422
rect 3105 51260 3327 51818
rect 11651 51260 11873 51818
rect 14721 51622 14907 52622
rect 3105 50884 11873 51260
rect 3105 50326 3327 50884
rect 11651 50326 11873 50884
rect 14721 50422 14907 51422
rect 3105 49950 11873 50326
rect 71 48854 257 49854
rect 3105 49392 3327 49950
rect 11651 49392 11873 49950
rect 3105 49016 11873 49392
rect 71 47654 257 48654
rect 3105 48458 3327 49016
rect 11651 48458 11873 49016
rect 14721 48854 14907 49854
rect 3105 48236 11873 48458
rect 2919 47654 3005 48022
rect 11973 47654 12059 48022
rect 14721 47654 14907 48654
rect 71 41658 257 42658
rect 13980 41658 14253 42658
rect 14721 41658 14907 42658
rect 71 40458 257 41458
rect 13980 40458 14253 41458
rect 14721 40458 14907 41458
rect 71 39258 257 40258
rect 13980 39258 14253 40258
rect 14721 39258 14907 40258
rect 71 38058 257 39058
rect 13980 38058 14253 39058
rect 14721 38058 14907 39058
rect 71 36858 257 37858
rect 13980 36858 14253 37858
rect 14721 36858 14907 37858
rect 71 35658 257 36658
rect 13980 35658 14253 36658
rect 14721 35658 14907 36658
rect 71 34458 257 35458
rect 13980 34458 14253 35458
rect 14721 34458 14907 35458
rect 71 33258 257 34258
rect 13980 33258 14253 34258
rect 14721 33258 14907 34258
rect 71 32058 257 33058
rect 13980 32058 14253 33058
rect 14721 32058 14907 33058
rect 71 30858 257 31858
rect 13980 30858 14253 31858
rect 14721 30858 14907 31858
rect 71 29658 257 30658
rect 13980 29658 14253 30658
rect 14721 29658 14907 30658
rect 71 28458 257 29458
rect 13980 28458 14253 29458
rect 14721 28458 14907 29458
rect 71 27258 257 28258
rect 13980 27190 14253 28190
rect 14721 27258 14907 28258
rect 71 26058 257 27058
rect 14721 26058 14907 27058
rect 71 24858 257 25858
rect 14721 24858 14907 25858
rect 71 23658 257 24658
rect 14721 23658 14907 24658
rect 71 22458 257 23458
rect 14721 22458 14907 23458
rect 71 20390 257 21390
rect 14721 20390 14907 21390
rect 71 19190 257 20190
rect 14721 19190 14907 20190
rect 71 17990 257 18990
rect 14721 17990 14907 18990
rect 71 16790 257 17790
rect 14721 16790 14907 17790
rect 71 15590 257 16590
rect 14721 15590 14907 16590
rect 71 14390 257 15390
rect 14721 14390 14907 15390
rect 71 13190 257 14190
rect 14721 13190 14907 14190
rect 71 11990 257 12990
rect 14721 11990 14907 12990
rect 71 10790 257 11790
rect 14721 10790 14907 11790
rect 71 9590 257 10590
rect 14721 9590 14907 10590
rect 71 8390 257 9390
rect 14721 8390 14907 9390
rect 71 7190 257 8190
rect 14721 7190 14907 8190
rect 71 5990 257 6990
rect 14721 5990 14907 6990
rect 71 4790 257 5790
rect 14721 4790 14907 5790
rect 71 3590 257 4590
rect 14721 3590 14907 4590
rect 71 2390 257 3390
rect 14721 2390 14907 3390
rect 71 1190 257 2190
rect 14721 1190 14907 2190
<< metal2 >>
rect -11 56007 10 57271
rect -11 52814 10 54186
rect -11 51200 86 52600
rect -11 48014 10 49386
rect 261 47163 2161 57600
rect -11 44814 10 46186
rect 2292 38400 2368 51000
rect 2481 47163 2681 57278
rect 2741 47163 4791 57600
rect 4851 47163 5051 57278
rect 5111 47163 7161 57600
rect 7221 47163 7757 57278
rect 7817 47163 9867 57600
rect 9927 47163 10127 57278
rect 10187 47163 12237 57600
rect 12297 47163 12497 57278
rect 12817 47163 14717 57600
rect 14968 56007 14989 57271
rect 14968 52814 14989 54186
rect 14892 51200 14989 52600
rect 14968 48014 14989 49386
rect 14968 44814 14989 46186
rect -11 36800 86 38200
rect 14892 36800 14989 38200
rect -11 33604 10 36596
rect 14968 33604 14989 36596
rect -11 27214 10 28586
rect 14968 27214 14989 28586
rect -11 12814 10 14186
rect 14968 12814 14989 14186
rect -11 8004 10 10996
rect 14968 8004 14989 10996
rect -11 4804 10 7796
rect 14968 4804 14989 7796
rect -11 1604 10 4596
rect 14968 1604 14989 4596
rect 261 0 2161 1190
rect 2741 0 4791 1190
rect 5111 0 7161 1190
rect 7817 0 9867 1190
rect 10187 0 12237 1190
rect 12817 0 14717 1190
use comp018green_esd_clamp_v5p0_DVSS  comp018green_esd_clamp_v5p0_DVSS_0
timestamp 1713338890
transform 1 0 1008 0 1 1090
box -747 -51 13709 46134
use M1_NWELL_CDNS_4066195314571  M1_NWELL_CDNS_4066195314571_0
timestamp 1713338890
transform 1 0 12243 0 1 50138
box -278 -2578 278 2578
use M1_NWELL_CDNS_4066195314571  M1_NWELL_CDNS_4066195314571_1
timestamp 1713338890
transform 1 0 2735 0 1 50138
box -278 -2578 278 2578
use M1_NWELL_CDNS_4066195314572  M1_NWELL_CDNS_4066195314572_0
timestamp 1713338890
transform 1 0 7489 0 1 47838
box -4578 -278 4578 278
use M1_NWELL_CDNS_4066195314572  M1_NWELL_CDNS_4066195314572_1
timestamp 1713338890
transform 1 0 7489 0 1 52438
box -4578 -278 4578 278
use M1_PSUB_CDNS_6903358316521  M1_PSUB_CDNS_6903358316521_0
timestamp 1713338890
transform 1 0 7489 0 1 48424
box -4087 -45 4087 45
use M1_PSUB_CDNS_6903358316521  M1_PSUB_CDNS_6903358316521_1
timestamp 1713338890
transform 1 0 7489 0 1 49358
box -4087 -45 4087 45
use M1_PSUB_CDNS_6903358316521  M1_PSUB_CDNS_6903358316521_2
timestamp 1713338890
transform 1 0 7489 0 1 49050
box -4087 -45 4087 45
use M1_PSUB_CDNS_6903358316521  M1_PSUB_CDNS_6903358316521_3
timestamp 1713338890
transform 1 0 7489 0 1 50292
box -4087 -45 4087 45
use M1_PSUB_CDNS_6903358316521  M1_PSUB_CDNS_6903358316521_4
timestamp 1713338890
transform 1 0 7489 0 1 49984
box -4087 -45 4087 45
use M1_PSUB_CDNS_6903358316521  M1_PSUB_CDNS_6903358316521_5
timestamp 1713338890
transform 1 0 7489 0 1 50918
box -4087 -45 4087 45
use M1_PSUB_CDNS_6903358316521  M1_PSUB_CDNS_6903358316521_6
timestamp 1713338890
transform 1 0 7489 0 1 51226
box -4087 -45 4087 45
use M1_PSUB_CDNS_6903358316521  M1_PSUB_CDNS_6903358316521_7
timestamp 1713338890
transform 1 0 7489 0 -1 51852
box -4087 -45 4087 45
use M1_PSUB_CDNS_6903358316522  M1_PSUB_CDNS_6903358316522_0
timestamp 1713338890
transform 1 0 7489 0 1 53228
box -7001 -45 7001 45
use M1_PSUB_CDNS_6903358316522  M1_PSUB_CDNS_6903358316522_1
timestamp 1713338890
transform 1 0 7489 0 1 57082
box -7001 -45 7001 45
use M1_PSUB_CDNS_6903358316545  M1_PSUB_CDNS_6903358316545_0
timestamp 1713338890
transform 1 0 3293 0 1 48737
box -45 -327 45 327
use M1_PSUB_CDNS_6903358316545  M1_PSUB_CDNS_6903358316545_1
timestamp 1713338890
transform 1 0 3293 0 1 49671
box -45 -327 45 327
use M1_PSUB_CDNS_6903358316545  M1_PSUB_CDNS_6903358316545_2
timestamp 1713338890
transform -1 0 11685 0 1 48737
box -45 -327 45 327
use M1_PSUB_CDNS_6903358316545  M1_PSUB_CDNS_6903358316545_3
timestamp 1713338890
transform -1 0 11685 0 1 49671
box -45 -327 45 327
use M1_PSUB_CDNS_6903358316545  M1_PSUB_CDNS_6903358316545_4
timestamp 1713338890
transform -1 0 11685 0 1 50605
box -45 -327 45 327
use M1_PSUB_CDNS_6903358316545  M1_PSUB_CDNS_6903358316545_5
timestamp 1713338890
transform 1 0 3293 0 1 50605
box -45 -327 45 327
use M1_PSUB_CDNS_6903358316545  M1_PSUB_CDNS_6903358316545_6
timestamp 1713338890
transform -1 0 11685 0 1 51539
box -45 -327 45 327
use M1_PSUB_CDNS_6903358316545  M1_PSUB_CDNS_6903358316545_7
timestamp 1713338890
transform 1 0 3293 0 1 51539
box -45 -327 45 327
use M1_PSUB_CDNS_69033583165487  M1_PSUB_CDNS_69033583165487_0
timestamp 1713338890
transform 1 0 491 0 1 21924
box -245 -20745 245 20745
use M1_PSUB_CDNS_69033583165487  M1_PSUB_CDNS_69033583165487_1
timestamp 1713338890
transform -1 0 14487 0 1 21924
box -245 -20745 245 20745
use M1_PSUB_CDNS_69033583165488  M1_PSUB_CDNS_69033583165488_0
timestamp 1713338890
transform -1 0 13496 0 1 34924
box -495 -7745 495 7745
use M1_PSUB_CDNS_69033583165489  M1_PSUB_CDNS_69033583165489_0
timestamp 1713338890
transform 1 0 7489 0 1 48270
box -4369 -45 4369 45
use M1_PSUB_CDNS_69033583165489  M1_PSUB_CDNS_69033583165489_1
timestamp 1713338890
transform 1 0 7489 0 -1 52006
box -4369 -45 4369 45
use M1_PSUB_CDNS_69033583165490  M1_PSUB_CDNS_69033583165490_0
timestamp 1713338890
transform 1 0 7489 0 1 49204
box -4181 -45 4181 45
use M1_PSUB_CDNS_69033583165490  M1_PSUB_CDNS_69033583165490_1
timestamp 1713338890
transform 1 0 7489 0 1 50138
box -4181 -45 4181 45
use M1_PSUB_CDNS_69033583165490  M1_PSUB_CDNS_69033583165490_2
timestamp 1713338890
transform 1 0 7489 0 1 51072
box -4181 -45 4181 45
use M1_PSUB_CDNS_69033583165508  M1_PSUB_CDNS_69033583165508_0
timestamp 1713338890
transform -1 0 11839 0 1 50138
box -45 -1784 45 1784
use M1_PSUB_CDNS_69033583165508  M1_PSUB_CDNS_69033583165508_1
timestamp 1713338890
transform 1 0 3139 0 1 50138
box -45 -1784 45 1784
use M1_PSUB_CDNS_69033583165512  M1_PSUB_CDNS_69033583165512_0
timestamp 1713338890
transform -1 0 13737 0 1 50138
box -995 -2495 995 2495
use M1_PSUB_CDNS_69033583165512  M1_PSUB_CDNS_69033583165512_1
timestamp 1713338890
transform 1 0 1241 0 1 50138
box -995 -2495 995 2495
use M1_PSUB_CDNS_69033583165513  M1_PSUB_CDNS_69033583165513_0
timestamp 1713338890
transform 1 0 379 0 1 55155
box -45 -1972 45 1972
use M1_PSUB_CDNS_69033583165513  M1_PSUB_CDNS_69033583165513_1
timestamp 1713338890
transform 1 0 14599 0 1 55155
box -45 -1972 45 1972
use M2_M1_CDNS_6903358316528  M2_M1_CDNS_6903358316528_0
timestamp 1713338890
transform 1 0 48 0 1 3100
box -38 -1496 38 1496
use M2_M1_CDNS_6903358316528  M2_M1_CDNS_6903358316528_1
timestamp 1713338890
transform 1 0 48 0 1 6300
box -38 -1496 38 1496
use M2_M1_CDNS_6903358316528  M2_M1_CDNS_6903358316528_2
timestamp 1713338890
transform 1 0 48 0 1 9500
box -38 -1496 38 1496
use M2_M1_CDNS_6903358316528  M2_M1_CDNS_6903358316528_3
timestamp 1713338890
transform 1 0 14930 0 1 3100
box -38 -1496 38 1496
use M2_M1_CDNS_6903358316528  M2_M1_CDNS_6903358316528_4
timestamp 1713338890
transform 1 0 14930 0 1 6300
box -38 -1496 38 1496
use M2_M1_CDNS_6903358316528  M2_M1_CDNS_6903358316528_5
timestamp 1713338890
transform 1 0 14930 0 1 9500
box -38 -1496 38 1496
use M2_M1_CDNS_6903358316528  M2_M1_CDNS_6903358316528_6
timestamp 1713338890
transform 1 0 48 0 1 35100
box -38 -1496 38 1496
use M2_M1_CDNS_6903358316528  M2_M1_CDNS_6903358316528_7
timestamp 1713338890
transform 1 0 14930 0 1 35100
box -38 -1496 38 1496
use M2_M1_CDNS_6903358316533  M2_M1_CDNS_6903358316533_0
timestamp 1713338890
transform 1 0 48 0 1 13500
box -38 -686 38 686
use M2_M1_CDNS_6903358316533  M2_M1_CDNS_6903358316533_1
timestamp 1713338890
transform 1 0 48 0 1 27900
box -38 -686 38 686
use M2_M1_CDNS_6903358316533  M2_M1_CDNS_6903358316533_2
timestamp 1713338890
transform 1 0 14930 0 1 13500
box -38 -686 38 686
use M2_M1_CDNS_6903358316533  M2_M1_CDNS_6903358316533_3
timestamp 1713338890
transform 1 0 14930 0 1 27900
box -38 -686 38 686
use M2_M1_CDNS_6903358316533  M2_M1_CDNS_6903358316533_4
timestamp 1713338890
transform 1 0 48 0 1 37500
box -38 -686 38 686
use M2_M1_CDNS_6903358316533  M2_M1_CDNS_6903358316533_5
timestamp 1713338890
transform 1 0 14930 0 1 37500
box -38 -686 38 686
use M2_M1_CDNS_6903358316533  M2_M1_CDNS_6903358316533_6
timestamp 1713338890
transform 1 0 48 0 1 45500
box -38 -686 38 686
use M2_M1_CDNS_6903358316533  M2_M1_CDNS_6903358316533_7
timestamp 1713338890
transform 1 0 14930 0 1 45500
box -38 -686 38 686
use M2_M1_CDNS_6903358316533  M2_M1_CDNS_6903358316533_8
timestamp 1713338890
transform 1 0 48 0 1 48700
box -38 -686 38 686
use M2_M1_CDNS_6903358316533  M2_M1_CDNS_6903358316533_9
timestamp 1713338890
transform 1 0 14930 0 1 48700
box -38 -686 38 686
use M2_M1_CDNS_6903358316533  M2_M1_CDNS_6903358316533_10
timestamp 1713338890
transform 1 0 48 0 1 51900
box -38 -686 38 686
use M2_M1_CDNS_6903358316533  M2_M1_CDNS_6903358316533_11
timestamp 1713338890
transform 1 0 14930 0 1 51900
box -38 -686 38 686
use M2_M1_CDNS_6903358316533  M2_M1_CDNS_6903358316533_12
timestamp 1713338890
transform 1 0 48 0 1 53500
box -38 -686 38 686
use M2_M1_CDNS_6903358316533  M2_M1_CDNS_6903358316533_13
timestamp 1713338890
transform 1 0 14930 0 1 53500
box -38 -686 38 686
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_0
timestamp 1713338890
transform 1 0 7489 0 1 47838
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_1
timestamp 1713338890
transform 1 0 7489 0 1 52438
box -254 -146 254 146
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_0
timestamp 1713338890
transform 1 0 7489 0 1 49671
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_1
timestamp 1713338890
transform 1 0 7489 0 1 48737
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_2
timestamp 1713338890
transform 1 0 7489 0 1 50605
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_3
timestamp 1713338890
transform 1 0 7489 0 1 51539
box -254 -92 254 92
use M2_M1_CDNS_69033583165348  M2_M1_CDNS_69033583165348_0
timestamp 1713338890
transform 1 0 4951 0 1 49671
box -92 -92 92 92
use M2_M1_CDNS_69033583165348  M2_M1_CDNS_69033583165348_1
timestamp 1713338890
transform 1 0 4951 0 1 48737
box -92 -92 92 92
use M2_M1_CDNS_69033583165348  M2_M1_CDNS_69033583165348_2
timestamp 1713338890
transform 1 0 10027 0 1 48737
box -92 -92 92 92
use M2_M1_CDNS_69033583165348  M2_M1_CDNS_69033583165348_3
timestamp 1713338890
transform 1 0 10027 0 1 49671
box -92 -92 92 92
use M2_M1_CDNS_69033583165348  M2_M1_CDNS_69033583165348_4
timestamp 1713338890
transform 1 0 10027 0 1 50605
box -92 -92 92 92
use M2_M1_CDNS_69033583165348  M2_M1_CDNS_69033583165348_5
timestamp 1713338890
transform 1 0 4951 0 1 50605
box -92 -92 92 92
use M2_M1_CDNS_69033583165348  M2_M1_CDNS_69033583165348_6
timestamp 1713338890
transform 1 0 10027 0 1 51539
box -92 -92 92 92
use M2_M1_CDNS_69033583165348  M2_M1_CDNS_69033583165348_7
timestamp 1713338890
transform 1 0 4951 0 1 51539
box -92 -92 92 92
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_0
timestamp 1713338890
transform 1 0 1211 0 1 792
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_1
timestamp 1713338890
transform 1 0 3766 0 1 792
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_2
timestamp 1713338890
transform 1 0 6136 0 1 792
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_3
timestamp 1713338890
transform 1 0 8842 0 1 792
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_4
timestamp 1713338890
transform 1 0 11212 0 1 792
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_5
timestamp 1713338890
transform 1 0 13767 0 1 792
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_6
timestamp 1713338890
transform 1 0 11212 0 1 57473
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_7
timestamp 1713338890
transform 1 0 8842 0 1 57473
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_8
timestamp 1713338890
transform 1 0 13767 0 1 57473
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_9
timestamp 1713338890
transform 1 0 6136 0 1 57473
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_10
timestamp 1713338890
transform 1 0 3766 0 1 57473
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_11
timestamp 1713338890
transform 1 0 1211 0 1 57473
box -902 -38 902 38
use M2_M1_CDNS_69033583165360  M2_M1_CDNS_69033583165360_0
timestamp 1713338890
transform 1 0 3275 0 1 53349
box -524 -146 524 146
use M2_M1_CDNS_69033583165360  M2_M1_CDNS_69033583165360_1
timestamp 1713338890
transform -1 0 11703 0 1 53349
box -524 -146 524 146
use M2_M1_CDNS_69033583165365  M2_M1_CDNS_69033583165365_0
timestamp 1713338890
transform 1 0 3943 0 1 48347
box -794 -92 794 92
use M2_M1_CDNS_69033583165365  M2_M1_CDNS_69033583165365_1
timestamp 1713338890
transform -1 0 11035 0 1 48347
box -794 -92 794 92
use M2_M1_CDNS_69033583165365  M2_M1_CDNS_69033583165365_2
timestamp 1713338890
transform -1 0 11035 0 1 51929
box -794 -92 794 92
use M2_M1_CDNS_69033583165365  M2_M1_CDNS_69033583165365_3
timestamp 1713338890
transform 1 0 3943 0 1 51929
box -794 -92 794 92
use M2_M1_CDNS_69033583165491  M2_M1_CDNS_69033583165491_0
timestamp 1713338890
transform 1 0 581 0 1 54943
box -224 -1712 224 1712
use M2_M1_CDNS_69033583165491  M2_M1_CDNS_69033583165491_1
timestamp 1713338890
transform -1 0 14397 0 1 54943
box -224 -1712 224 1712
use M2_M1_CDNS_69033583165492  M2_M1_CDNS_69033583165492_0
timestamp 1713338890
transform 1 0 4053 0 1 54943
box -162 -1712 162 1712
use M2_M1_CDNS_69033583165492  M2_M1_CDNS_69033583165492_1
timestamp 1713338890
transform -1 0 10925 0 1 54943
box -162 -1712 162 1712
use M2_M1_CDNS_69033583165494  M2_M1_CDNS_69033583165494_0
timestamp 1713338890
transform 1 0 48 0 1 56639
box -38 -632 38 632
use M2_M1_CDNS_69033583165494  M2_M1_CDNS_69033583165494_1
timestamp 1713338890
transform 1 0 14930 0 1 56639
box -38 -632 38 632
use M2_M1_CDNS_69033583165499  M2_M1_CDNS_69033583165499_0
timestamp 1713338890
transform 1 0 12362 0 1 50138
box -38 -2468 38 2468
use M2_M1_CDNS_69033583165499  M2_M1_CDNS_69033583165499_1
timestamp 1713338890
transform 1 0 2616 0 1 50138
box -38 -2468 38 2468
use M2_M1_CDNS_69033583165500  M2_M1_CDNS_69033583165500_0
timestamp 1713338890
transform 1 0 4951 0 1 55155
box -92 -1550 92 1550
use M2_M1_CDNS_69033583165500  M2_M1_CDNS_69033583165500_1
timestamp 1713338890
transform 1 0 10027 0 1 55155
box -92 -1550 92 1550
use M2_M1_CDNS_69033583165501  M2_M1_CDNS_69033583165501_0
timestamp 1713338890
transform 1 0 1489 0 1 53349
box -632 -146 632 146
use M2_M1_CDNS_69033583165501  M2_M1_CDNS_69033583165501_1
timestamp 1713338890
transform -1 0 13489 0 1 53349
box -632 -146 632 146
use M2_M1_CDNS_69033583165502  M2_M1_CDNS_69033583165502_0
timestamp 1713338890
transform -1 0 13767 0 1 57078
box -848 -38 848 38
use M2_M1_CDNS_69033583165502  M2_M1_CDNS_69033583165502_1
timestamp 1713338890
transform 1 0 1211 0 1 57078
box -848 -38 848 38
use M2_M1_CDNS_69033583165503  M2_M1_CDNS_69033583165503_0
timestamp 1713338890
transform 1 0 3943 0 1 49204
box -794 -146 794 146
use M2_M1_CDNS_69033583165503  M2_M1_CDNS_69033583165503_1
timestamp 1713338890
transform -1 0 11035 0 1 49204
box -794 -146 794 146
use M2_M1_CDNS_69033583165503  M2_M1_CDNS_69033583165503_2
timestamp 1713338890
transform -1 0 11035 0 1 50138
box -794 -146 794 146
use M2_M1_CDNS_69033583165503  M2_M1_CDNS_69033583165503_3
timestamp 1713338890
transform 1 0 3943 0 1 50138
box -794 -146 794 146
use M2_M1_CDNS_69033583165503  M2_M1_CDNS_69033583165503_4
timestamp 1713338890
transform -1 0 11035 0 1 51072
box -794 -146 794 146
use M2_M1_CDNS_69033583165503  M2_M1_CDNS_69033583165503_5
timestamp 1713338890
transform 1 0 3943 0 1 51072
box -794 -146 794 146
use M2_M1_CDNS_69033583165506  M2_M1_CDNS_69033583165506_0
timestamp 1713338890
transform 1 0 6136 0 1 48347
box -1010 -92 1010 92
use M2_M1_CDNS_69033583165506  M2_M1_CDNS_69033583165506_1
timestamp 1713338890
transform 1 0 8842 0 1 48347
box -1010 -92 1010 92
use M2_M1_CDNS_69033583165506  M2_M1_CDNS_69033583165506_2
timestamp 1713338890
transform 1 0 8842 0 1 51929
box -1010 -92 1010 92
use M2_M1_CDNS_69033583165506  M2_M1_CDNS_69033583165506_3
timestamp 1713338890
transform 1 0 6136 0 1 51929
box -1010 -92 1010 92
use M2_M1_CDNS_69033583165507  M2_M1_CDNS_69033583165507_0
timestamp 1713338890
transform 1 0 4951 0 1 47838
box -92 -146 92 146
use M2_M1_CDNS_69033583165507  M2_M1_CDNS_69033583165507_1
timestamp 1713338890
transform 1 0 10027 0 1 47838
box -92 -146 92 146
use M2_M1_CDNS_69033583165507  M2_M1_CDNS_69033583165507_2
timestamp 1713338890
transform 1 0 10027 0 1 52438
box -92 -146 92 146
use M2_M1_CDNS_69033583165507  M2_M1_CDNS_69033583165507_3
timestamp 1713338890
transform 1 0 4951 0 1 52438
box -92 -146 92 146
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_0
timestamp 1713338890
transform -1 0 8842 0 1 57078
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_1
timestamp 1713338890
transform -1 0 11212 0 1 57078
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_2
timestamp 1713338890
transform 1 0 3766 0 1 57078
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_3
timestamp 1713338890
transform -1 0 6136 0 1 57078
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165510  M2_M1_CDNS_69033583165510_0
timestamp 1713338890
transform 1 0 6136 0 1 49204
box -1010 -146 1010 146
use M2_M1_CDNS_69033583165510  M2_M1_CDNS_69033583165510_1
timestamp 1713338890
transform 1 0 8842 0 1 49204
box -1010 -146 1010 146
use M2_M1_CDNS_69033583165510  M2_M1_CDNS_69033583165510_2
timestamp 1713338890
transform 1 0 8842 0 1 50138
box -1010 -146 1010 146
use M2_M1_CDNS_69033583165510  M2_M1_CDNS_69033583165510_3
timestamp 1713338890
transform 1 0 6136 0 1 50138
box -1010 -146 1010 146
use M2_M1_CDNS_69033583165510  M2_M1_CDNS_69033583165510_4
timestamp 1713338890
transform 1 0 8842 0 1 51072
box -1010 -146 1010 146
use M2_M1_CDNS_69033583165510  M2_M1_CDNS_69033583165510_5
timestamp 1713338890
transform 1 0 6136 0 1 51072
box -1010 -146 1010 146
use M2_M1_CDNS_69033583165510  M2_M1_CDNS_69033583165510_6
timestamp 1713338890
transform -1 0 6136 0 1 53349
box -1010 -146 1010 146
use M2_M1_CDNS_69033583165510  M2_M1_CDNS_69033583165510_7
timestamp 1713338890
transform -1 0 8842 0 1 53349
box -1010 -146 1010 146
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_0
timestamp 1713338890
transform 1 0 2581 0 1 53595
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_1
timestamp 1713338890
transform 1 0 12397 0 1 53595
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_2
timestamp 1713338890
transform 1 0 12397 0 1 56715
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_3
timestamp 1713338890
transform 1 0 2581 0 1 56715
box -92 -38 92 38
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_0
timestamp 1713338890
transform 1 0 7489 0 1 29500
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_1
timestamp 1713338890
transform 1 0 7489 0 1 11900
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_2
timestamp 1713338890
transform 1 0 7489 0 1 42300
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_3
timestamp 1713338890
transform 1 0 7489 0 1 40700
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_4
timestamp 1713338890
transform 1 0 7489 0 1 43900
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_5
timestamp 1713338890
transform 1 0 7489 0 1 47100
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_6
timestamp 1713338890
transform 1 0 7489 0 1 55100
box -224 -658 224 658
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_0
timestamp 1713338890
transform 1 0 7489 0 1 15900
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_1
timestamp 1713338890
transform 1 0 7489 0 1 19100
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_2
timestamp 1713338890
transform 1 0 7489 0 1 25500
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_3
timestamp 1713338890
transform 1 0 7489 0 1 22300
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_4
timestamp 1713338890
transform 1 0 7489 0 1 31900
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_0
timestamp 1713338890
transform 1 0 2581 0 1 11900
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_1
timestamp 1713338890
transform 1 0 2581 0 1 29500
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_2
timestamp 1713338890
transform 1 0 4951 0 1 11900
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_3
timestamp 1713338890
transform 1 0 4951 0 1 29500
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_4
timestamp 1713338890
transform -1 0 10027 0 1 11900
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_5
timestamp 1713338890
transform -1 0 10027 0 1 29500
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_6
timestamp 1713338890
transform -1 0 12397 0 1 11900
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_7
timestamp 1713338890
transform -1 0 12397 0 1 29500
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_8
timestamp 1713338890
transform 1 0 2581 0 1 42300
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_9
timestamp 1713338890
transform 1 0 2581 0 1 40700
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_10
timestamp 1713338890
transform 1 0 4951 0 1 42300
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_11
timestamp 1713338890
transform 1 0 4951 0 1 40700
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_12
timestamp 1713338890
transform -1 0 10027 0 1 42300
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_13
timestamp 1713338890
transform -1 0 10027 0 1 40700
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_14
timestamp 1713338890
transform -1 0 12397 0 1 42300
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_15
timestamp 1713338890
transform -1 0 12397 0 1 40700
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_16
timestamp 1713338890
transform 1 0 2581 0 1 43900
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_17
timestamp 1713338890
transform 1 0 4951 0 1 43900
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_18
timestamp 1713338890
transform -1 0 10027 0 1 43900
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_19
timestamp 1713338890
transform -1 0 12397 0 1 43900
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_20
timestamp 1713338890
transform 1 0 2581 0 1 47100
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_21
timestamp 1713338890
transform 1 0 4951 0 1 47100
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_22
timestamp 1713338890
transform -1 0 10027 0 1 47100
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_23
timestamp 1713338890
transform -1 0 12397 0 1 47100
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_24
timestamp 1713338890
transform 1 0 2581 0 1 55100
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_25
timestamp 1713338890
transform 1 0 4951 0 1 55100
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_26
timestamp 1713338890
transform -1 0 10027 0 1 55100
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_27
timestamp 1713338890
transform -1 0 12397 0 1 55100
box -100 -658 100 658
use M3_M2_CDNS_6903358316534  M3_M2_CDNS_6903358316534_0
timestamp 1713338890
transform 1 0 48 0 1 13500
box -38 -686 38 686
use M3_M2_CDNS_6903358316534  M3_M2_CDNS_6903358316534_1
timestamp 1713338890
transform 1 0 48 0 1 27900
box -38 -686 38 686
use M3_M2_CDNS_6903358316534  M3_M2_CDNS_6903358316534_2
timestamp 1713338890
transform 1 0 14930 0 1 13500
box -38 -686 38 686
use M3_M2_CDNS_6903358316534  M3_M2_CDNS_6903358316534_3
timestamp 1713338890
transform 1 0 14930 0 1 27900
box -38 -686 38 686
use M3_M2_CDNS_6903358316534  M3_M2_CDNS_6903358316534_4
timestamp 1713338890
transform 1 0 48 0 1 37500
box -38 -686 38 686
use M3_M2_CDNS_6903358316534  M3_M2_CDNS_6903358316534_5
timestamp 1713338890
transform 1 0 14930 0 1 37500
box -38 -686 38 686
use M3_M2_CDNS_6903358316534  M3_M2_CDNS_6903358316534_6
timestamp 1713338890
transform 1 0 48 0 1 45500
box -38 -686 38 686
use M3_M2_CDNS_6903358316534  M3_M2_CDNS_6903358316534_7
timestamp 1713338890
transform 1 0 14930 0 1 45500
box -38 -686 38 686
use M3_M2_CDNS_6903358316534  M3_M2_CDNS_6903358316534_8
timestamp 1713338890
transform 1 0 48 0 1 48700
box -38 -686 38 686
use M3_M2_CDNS_6903358316534  M3_M2_CDNS_6903358316534_9
timestamp 1713338890
transform 1 0 14930 0 1 48700
box -38 -686 38 686
use M3_M2_CDNS_6903358316534  M3_M2_CDNS_6903358316534_10
timestamp 1713338890
transform 1 0 48 0 1 51900
box -38 -686 38 686
use M3_M2_CDNS_6903358316534  M3_M2_CDNS_6903358316534_11
timestamp 1713338890
transform 1 0 14930 0 1 51900
box -38 -686 38 686
use M3_M2_CDNS_6903358316534  M3_M2_CDNS_6903358316534_12
timestamp 1713338890
transform 1 0 48 0 1 53500
box -38 -686 38 686
use M3_M2_CDNS_6903358316534  M3_M2_CDNS_6903358316534_13
timestamp 1713338890
transform 1 0 14930 0 1 53500
box -38 -686 38 686
use M3_M2_CDNS_69033583165372  M3_M2_CDNS_69033583165372_0
timestamp 1713338890
transform 1 0 1211 0 1 3100
box -906 -1464 906 1464
use M3_M2_CDNS_69033583165372  M3_M2_CDNS_69033583165372_1
timestamp 1713338890
transform 1 0 1211 0 1 6300
box -906 -1464 906 1464
use M3_M2_CDNS_69033583165372  M3_M2_CDNS_69033583165372_2
timestamp 1713338890
transform 1 0 1211 0 1 9500
box -906 -1464 906 1464
use M3_M2_CDNS_69033583165372  M3_M2_CDNS_69033583165372_3
timestamp 1713338890
transform -1 0 13767 0 1 3100
box -906 -1464 906 1464
use M3_M2_CDNS_69033583165372  M3_M2_CDNS_69033583165372_4
timestamp 1713338890
transform -1 0 13767 0 1 9500
box -906 -1464 906 1464
use M3_M2_CDNS_69033583165372  M3_M2_CDNS_69033583165372_5
timestamp 1713338890
transform -1 0 13767 0 1 6300
box -906 -1464 906 1464
use M3_M2_CDNS_69033583165372  M3_M2_CDNS_69033583165372_6
timestamp 1713338890
transform 1 0 1211 0 1 35100
box -906 -1464 906 1464
use M3_M2_CDNS_69033583165372  M3_M2_CDNS_69033583165372_7
timestamp 1713338890
transform -1 0 13767 0 1 35100
box -906 -1464 906 1464
use M3_M2_CDNS_69033583165373  M3_M2_CDNS_69033583165373_0
timestamp 1713338890
transform 1 0 1211 0 1 13500
box -906 -658 906 658
use M3_M2_CDNS_69033583165373  M3_M2_CDNS_69033583165373_1
timestamp 1713338890
transform 1 0 1211 0 1 27900
box -906 -658 906 658
use M3_M2_CDNS_69033583165373  M3_M2_CDNS_69033583165373_2
timestamp 1713338890
transform -1 0 13767 0 1 13500
box -906 -658 906 658
use M3_M2_CDNS_69033583165373  M3_M2_CDNS_69033583165373_3
timestamp 1713338890
transform -1 0 13767 0 1 27900
box -906 -658 906 658
use M3_M2_CDNS_69033583165373  M3_M2_CDNS_69033583165373_4
timestamp 1713338890
transform 1 0 1211 0 1 37500
box -906 -658 906 658
use M3_M2_CDNS_69033583165373  M3_M2_CDNS_69033583165373_5
timestamp 1713338890
transform -1 0 13767 0 1 37500
box -906 -658 906 658
use M3_M2_CDNS_69033583165373  M3_M2_CDNS_69033583165373_6
timestamp 1713338890
transform 1 0 1211 0 1 45500
box -906 -658 906 658
use M3_M2_CDNS_69033583165373  M3_M2_CDNS_69033583165373_7
timestamp 1713338890
transform -1 0 13767 0 1 45500
box -906 -658 906 658
use M3_M2_CDNS_69033583165373  M3_M2_CDNS_69033583165373_8
timestamp 1713338890
transform 1 0 1211 0 1 48700
box -906 -658 906 658
use M3_M2_CDNS_69033583165373  M3_M2_CDNS_69033583165373_9
timestamp 1713338890
transform -1 0 13767 0 1 48700
box -906 -658 906 658
use M3_M2_CDNS_69033583165373  M3_M2_CDNS_69033583165373_10
timestamp 1713338890
transform 1 0 1211 0 1 51900
box -906 -658 906 658
use M3_M2_CDNS_69033583165373  M3_M2_CDNS_69033583165373_11
timestamp 1713338890
transform -1 0 13767 0 1 51900
box -906 -658 906 658
use M3_M2_CDNS_69033583165373  M3_M2_CDNS_69033583165373_12
timestamp 1713338890
transform 1 0 1211 0 1 53500
box -906 -658 906 658
use M3_M2_CDNS_69033583165373  M3_M2_CDNS_69033583165373_13
timestamp 1713338890
transform -1 0 13767 0 1 53500
box -906 -658 906 658
use M3_M2_CDNS_69033583165493  M3_M2_CDNS_69033583165493_0
timestamp 1713338890
transform 1 0 3766 0 1 56639
box -968 -596 968 596
use M3_M2_CDNS_69033583165493  M3_M2_CDNS_69033583165493_1
timestamp 1713338890
transform 1 0 6136 0 1 56639
box -968 -596 968 596
use M3_M2_CDNS_69033583165493  M3_M2_CDNS_69033583165493_2
timestamp 1713338890
transform -1 0 8842 0 1 56639
box -968 -596 968 596
use M3_M2_CDNS_69033583165493  M3_M2_CDNS_69033583165493_3
timestamp 1713338890
transform -1 0 11212 0 1 56639
box -968 -596 968 596
use M3_M2_CDNS_69033583165495  M3_M2_CDNS_69033583165495_0
timestamp 1713338890
transform 1 0 48 0 1 56639
box -38 -632 38 632
use M3_M2_CDNS_69033583165495  M3_M2_CDNS_69033583165495_1
timestamp 1713338890
transform 1 0 14930 0 1 56639
box -38 -632 38 632
use M3_M2_CDNS_69033583165496  M3_M2_CDNS_69033583165496_0
timestamp 1713338890
transform 1 0 48 0 1 3100
box -38 -1496 38 1496
use M3_M2_CDNS_69033583165496  M3_M2_CDNS_69033583165496_1
timestamp 1713338890
transform 1 0 48 0 1 6300
box -38 -1496 38 1496
use M3_M2_CDNS_69033583165496  M3_M2_CDNS_69033583165496_2
timestamp 1713338890
transform 1 0 48 0 1 9500
box -38 -1496 38 1496
use M3_M2_CDNS_69033583165496  M3_M2_CDNS_69033583165496_3
timestamp 1713338890
transform 1 0 14930 0 1 3100
box -38 -1496 38 1496
use M3_M2_CDNS_69033583165496  M3_M2_CDNS_69033583165496_4
timestamp 1713338890
transform 1 0 14930 0 1 6300
box -38 -1496 38 1496
use M3_M2_CDNS_69033583165496  M3_M2_CDNS_69033583165496_5
timestamp 1713338890
transform 1 0 14930 0 1 9500
box -38 -1496 38 1496
use M3_M2_CDNS_69033583165496  M3_M2_CDNS_69033583165496_6
timestamp 1713338890
transform 1 0 48 0 1 35100
box -38 -1496 38 1496
use M3_M2_CDNS_69033583165496  M3_M2_CDNS_69033583165496_7
timestamp 1713338890
transform 1 0 14930 0 1 35100
box -38 -1496 38 1496
use M3_M2_CDNS_69033583165497  M3_M2_CDNS_69033583165497_0
timestamp 1713338890
transform 1 0 2581 0 1 15900
box -100 -1464 100 1464
use M3_M2_CDNS_69033583165497  M3_M2_CDNS_69033583165497_1
timestamp 1713338890
transform 1 0 2581 0 1 19100
box -100 -1464 100 1464
use M3_M2_CDNS_69033583165497  M3_M2_CDNS_69033583165497_2
timestamp 1713338890
transform 1 0 2581 0 1 22300
box -100 -1464 100 1464
use M3_M2_CDNS_69033583165497  M3_M2_CDNS_69033583165497_3
timestamp 1713338890
transform 1 0 2581 0 1 25500
box -100 -1464 100 1464
use M3_M2_CDNS_69033583165497  M3_M2_CDNS_69033583165497_4
timestamp 1713338890
transform 1 0 4951 0 1 15900
box -100 -1464 100 1464
use M3_M2_CDNS_69033583165497  M3_M2_CDNS_69033583165497_5
timestamp 1713338890
transform 1 0 4951 0 1 19100
box -100 -1464 100 1464
use M3_M2_CDNS_69033583165497  M3_M2_CDNS_69033583165497_6
timestamp 1713338890
transform 1 0 4951 0 1 22300
box -100 -1464 100 1464
use M3_M2_CDNS_69033583165497  M3_M2_CDNS_69033583165497_7
timestamp 1713338890
transform 1 0 4951 0 1 25500
box -100 -1464 100 1464
use M3_M2_CDNS_69033583165497  M3_M2_CDNS_69033583165497_8
timestamp 1713338890
transform -1 0 10027 0 1 15900
box -100 -1464 100 1464
use M3_M2_CDNS_69033583165497  M3_M2_CDNS_69033583165497_9
timestamp 1713338890
transform -1 0 10027 0 1 19100
box -100 -1464 100 1464
use M3_M2_CDNS_69033583165497  M3_M2_CDNS_69033583165497_10
timestamp 1713338890
transform -1 0 10027 0 1 22300
box -100 -1464 100 1464
use M3_M2_CDNS_69033583165497  M3_M2_CDNS_69033583165497_11
timestamp 1713338890
transform -1 0 10027 0 1 25500
box -100 -1464 100 1464
use M3_M2_CDNS_69033583165497  M3_M2_CDNS_69033583165497_12
timestamp 1713338890
transform -1 0 12397 0 1 15900
box -100 -1464 100 1464
use M3_M2_CDNS_69033583165497  M3_M2_CDNS_69033583165497_13
timestamp 1713338890
transform -1 0 12397 0 1 19100
box -100 -1464 100 1464
use M3_M2_CDNS_69033583165497  M3_M2_CDNS_69033583165497_14
timestamp 1713338890
transform -1 0 12397 0 1 22300
box -100 -1464 100 1464
use M3_M2_CDNS_69033583165497  M3_M2_CDNS_69033583165497_15
timestamp 1713338890
transform -1 0 12397 0 1 25500
box -100 -1464 100 1464
use M3_M2_CDNS_69033583165497  M3_M2_CDNS_69033583165497_16
timestamp 1713338890
transform 1 0 2581 0 1 31900
box -100 -1464 100 1464
use M3_M2_CDNS_69033583165497  M3_M2_CDNS_69033583165497_17
timestamp 1713338890
transform 1 0 4951 0 1 31900
box -100 -1464 100 1464
use M3_M2_CDNS_69033583165497  M3_M2_CDNS_69033583165497_18
timestamp 1713338890
transform -1 0 10027 0 1 31900
box -100 -1464 100 1464
use M3_M2_CDNS_69033583165497  M3_M2_CDNS_69033583165497_19
timestamp 1713338890
transform -1 0 12397 0 1 31900
box -100 -1464 100 1464
use M3_M2_CDNS_69033583165498  M3_M2_CDNS_69033583165498_0
timestamp 1713338890
transform 1 0 1211 0 1 56639
box -906 -596 906 596
use M3_M2_CDNS_69033583165498  M3_M2_CDNS_69033583165498_1
timestamp 1713338890
transform -1 0 13767 0 1 56639
box -906 -596 906 596
use M3_M2_CDNS_69033583165504  M3_M2_CDNS_69033583165504_0
timestamp 1713338890
transform 1 0 3766 0 1 3100
box -968 -1464 968 1464
use M3_M2_CDNS_69033583165504  M3_M2_CDNS_69033583165504_1
timestamp 1713338890
transform 1 0 3766 0 1 6300
box -968 -1464 968 1464
use M3_M2_CDNS_69033583165504  M3_M2_CDNS_69033583165504_2
timestamp 1713338890
transform 1 0 3766 0 1 9500
box -968 -1464 968 1464
use M3_M2_CDNS_69033583165504  M3_M2_CDNS_69033583165504_3
timestamp 1713338890
transform 1 0 6136 0 1 3100
box -968 -1464 968 1464
use M3_M2_CDNS_69033583165504  M3_M2_CDNS_69033583165504_4
timestamp 1713338890
transform 1 0 6136 0 1 6300
box -968 -1464 968 1464
use M3_M2_CDNS_69033583165504  M3_M2_CDNS_69033583165504_5
timestamp 1713338890
transform 1 0 6136 0 1 9500
box -968 -1464 968 1464
use M3_M2_CDNS_69033583165504  M3_M2_CDNS_69033583165504_6
timestamp 1713338890
transform -1 0 8842 0 1 9500
box -968 -1464 968 1464
use M3_M2_CDNS_69033583165504  M3_M2_CDNS_69033583165504_7
timestamp 1713338890
transform -1 0 8842 0 1 3100
box -968 -1464 968 1464
use M3_M2_CDNS_69033583165504  M3_M2_CDNS_69033583165504_8
timestamp 1713338890
transform -1 0 8842 0 1 6300
box -968 -1464 968 1464
use M3_M2_CDNS_69033583165504  M3_M2_CDNS_69033583165504_9
timestamp 1713338890
transform -1 0 11212 0 1 3100
box -968 -1464 968 1464
use M3_M2_CDNS_69033583165504  M3_M2_CDNS_69033583165504_10
timestamp 1713338890
transform -1 0 11212 0 1 6300
box -968 -1464 968 1464
use M3_M2_CDNS_69033583165504  M3_M2_CDNS_69033583165504_11
timestamp 1713338890
transform -1 0 11212 0 1 9500
box -968 -1464 968 1464
use M3_M2_CDNS_69033583165504  M3_M2_CDNS_69033583165504_12
timestamp 1713338890
transform 1 0 3766 0 1 35100
box -968 -1464 968 1464
use M3_M2_CDNS_69033583165504  M3_M2_CDNS_69033583165504_13
timestamp 1713338890
transform 1 0 6136 0 1 35100
box -968 -1464 968 1464
use M3_M2_CDNS_69033583165504  M3_M2_CDNS_69033583165504_14
timestamp 1713338890
transform -1 0 8842 0 1 35100
box -968 -1464 968 1464
use M3_M2_CDNS_69033583165504  M3_M2_CDNS_69033583165504_15
timestamp 1713338890
transform -1 0 11212 0 1 35100
box -968 -1464 968 1464
use M3_M2_CDNS_69033583165505  M3_M2_CDNS_69033583165505_0
timestamp 1713338890
transform 1 0 3766 0 1 13500
box -968 -658 968 658
use M3_M2_CDNS_69033583165505  M3_M2_CDNS_69033583165505_1
timestamp 1713338890
transform 1 0 3766 0 1 27900
box -968 -658 968 658
use M3_M2_CDNS_69033583165505  M3_M2_CDNS_69033583165505_2
timestamp 1713338890
transform 1 0 6136 0 1 13500
box -968 -658 968 658
use M3_M2_CDNS_69033583165505  M3_M2_CDNS_69033583165505_3
timestamp 1713338890
transform 1 0 6136 0 1 27900
box -968 -658 968 658
use M3_M2_CDNS_69033583165505  M3_M2_CDNS_69033583165505_4
timestamp 1713338890
transform -1 0 8842 0 1 13500
box -968 -658 968 658
use M3_M2_CDNS_69033583165505  M3_M2_CDNS_69033583165505_5
timestamp 1713338890
transform -1 0 8842 0 1 27900
box -968 -658 968 658
use M3_M2_CDNS_69033583165505  M3_M2_CDNS_69033583165505_6
timestamp 1713338890
transform -1 0 11212 0 1 13500
box -968 -658 968 658
use M3_M2_CDNS_69033583165505  M3_M2_CDNS_69033583165505_7
timestamp 1713338890
transform -1 0 11212 0 1 27900
box -968 -658 968 658
use M3_M2_CDNS_69033583165505  M3_M2_CDNS_69033583165505_8
timestamp 1713338890
transform 1 0 3766 0 1 37500
box -968 -658 968 658
use M3_M2_CDNS_69033583165505  M3_M2_CDNS_69033583165505_9
timestamp 1713338890
transform 1 0 6136 0 1 37500
box -968 -658 968 658
use M3_M2_CDNS_69033583165505  M3_M2_CDNS_69033583165505_10
timestamp 1713338890
transform -1 0 8842 0 1 37500
box -968 -658 968 658
use M3_M2_CDNS_69033583165505  M3_M2_CDNS_69033583165505_11
timestamp 1713338890
transform -1 0 11212 0 1 37500
box -968 -658 968 658
use M3_M2_CDNS_69033583165505  M3_M2_CDNS_69033583165505_12
timestamp 1713338890
transform 1 0 3766 0 1 45500
box -968 -658 968 658
use M3_M2_CDNS_69033583165505  M3_M2_CDNS_69033583165505_13
timestamp 1713338890
transform 1 0 6136 0 1 45500
box -968 -658 968 658
use M3_M2_CDNS_69033583165505  M3_M2_CDNS_69033583165505_14
timestamp 1713338890
transform -1 0 8842 0 1 45500
box -968 -658 968 658
use M3_M2_CDNS_69033583165505  M3_M2_CDNS_69033583165505_15
timestamp 1713338890
transform -1 0 11212 0 1 45500
box -968 -658 968 658
use M3_M2_CDNS_69033583165505  M3_M2_CDNS_69033583165505_16
timestamp 1713338890
transform 1 0 3766 0 1 48700
box -968 -658 968 658
use M3_M2_CDNS_69033583165505  M3_M2_CDNS_69033583165505_17
timestamp 1713338890
transform 1 0 6136 0 1 48700
box -968 -658 968 658
use M3_M2_CDNS_69033583165505  M3_M2_CDNS_69033583165505_18
timestamp 1713338890
transform -1 0 8842 0 1 48700
box -968 -658 968 658
use M3_M2_CDNS_69033583165505  M3_M2_CDNS_69033583165505_19
timestamp 1713338890
transform -1 0 11212 0 1 48700
box -968 -658 968 658
use M3_M2_CDNS_69033583165505  M3_M2_CDNS_69033583165505_20
timestamp 1713338890
transform 1 0 3766 0 1 51900
box -968 -658 968 658
use M3_M2_CDNS_69033583165505  M3_M2_CDNS_69033583165505_21
timestamp 1713338890
transform 1 0 6136 0 1 51900
box -968 -658 968 658
use M3_M2_CDNS_69033583165505  M3_M2_CDNS_69033583165505_22
timestamp 1713338890
transform -1 0 8842 0 1 51900
box -968 -658 968 658
use M3_M2_CDNS_69033583165505  M3_M2_CDNS_69033583165505_23
timestamp 1713338890
transform -1 0 11212 0 1 51900
box -968 -658 968 658
use M3_M2_CDNS_69033583165505  M3_M2_CDNS_69033583165505_24
timestamp 1713338890
transform 1 0 3766 0 1 53500
box -968 -658 968 658
use M3_M2_CDNS_69033583165505  M3_M2_CDNS_69033583165505_25
timestamp 1713338890
transform 1 0 6136 0 1 53500
box -968 -658 968 658
use M3_M2_CDNS_69033583165505  M3_M2_CDNS_69033583165505_26
timestamp 1713338890
transform -1 0 8842 0 1 53500
box -968 -658 968 658
use M3_M2_CDNS_69033583165505  M3_M2_CDNS_69033583165505_27
timestamp 1713338890
transform -1 0 11212 0 1 53500
box -968 -658 968 658
use M3_M2_CDNS_69033583165514  M3_M2_CDNS_69033583165514_0
timestamp 1713338890
transform 1 0 2330 0 1 39105
box -38 -632 38 632
use M3_M2_CDNS_69033583165514  M3_M2_CDNS_69033583165514_1
timestamp 1713338890
transform 1 0 2330 0 1 50304
box -38 -632 38 632
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_0
timestamp 1713338890
transform 1 0 835 0 1 53655
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_1
timestamp 1713338890
transform 1 0 4271 0 1 53655
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_2
timestamp 1713338890
transform 1 0 7707 0 1 53655
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_3
timestamp 1713338890
transform 1 0 11143 0 1 53655
box -218 -350 3218 3092
use np_6p0_CDNS_406619531451  np_6p0_CDNS_406619531451_0
timestamp 1713338890
transform 1 0 3489 0 1 48637
box 0 0 8000 200
use np_6p0_CDNS_406619531451  np_6p0_CDNS_406619531451_1
timestamp 1713338890
transform 1 0 3489 0 1 49571
box 0 0 8000 200
use np_6p0_CDNS_406619531451  np_6p0_CDNS_406619531451_2
timestamp 1713338890
transform 1 0 3489 0 1 50505
box 0 0 8000 200
use np_6p0_CDNS_406619531451  np_6p0_CDNS_406619531451_3
timestamp 1713338890
transform 1 0 3489 0 1 51439
box 0 0 8000 200
<< labels >>
rlabel metal3 s 774 11795 774 11795 4 DVDD
port 1 nsew
rlabel metal3 s 774 22234 774 22234 4 DVDD
port 1 nsew
rlabel metal3 s 774 19120 774 19120 4 DVDD
port 1 nsew
rlabel metal3 s 774 15905 774 15905 4 DVDD
port 1 nsew
rlabel metal3 s 774 29488 774 29488 4 DVDD
port 1 nsew
rlabel metal3 s 774 25470 774 25470 4 DVDD
port 1 nsew
rlabel metal3 s 774 31879 774 31879 4 DVDD
port 1 nsew
rlabel metal3 s 774 43934 774 43934 4 DVDD
port 1 nsew
rlabel metal3 s 774 42169 774 42169 4 DVDD
port 1 nsew
rlabel metal3 s 774 40734 774 40734 4 DVDD
port 1 nsew
rlabel metal3 s 774 54969 774 54969 4 DVDD
port 1 nsew
rlabel metal3 s 774 47134 774 47134 4 DVDD
port 1 nsew
rlabel metal3 s 705 6432 705 6432 4 DVSS
port 2 nsew
rlabel metal3 s 752 3261 752 3261 4 DVSS
port 2 nsew
rlabel metal3 s 774 9418 774 9418 4 DVSS
port 2 nsew
rlabel metal3 s 774 13611 774 13611 4 DVSS
port 2 nsew
rlabel metal3 s 774 27853 774 27853 4 DVSS
port 2 nsew
rlabel metal3 s 774 35106 774 35106 4 DVSS
port 2 nsew
rlabel metal3 s 774 37534 774 37534 4 DVSS
port 2 nsew
rlabel metal3 s 774 45369 774 45369 4 DVSS
port 2 nsew
rlabel metal3 s 774 51769 774 51769 4 DVSS
port 2 nsew
rlabel metal3 s 774 48569 774 48569 4 DVSS
port 2 nsew
rlabel metal3 s 774 53534 774 53534 4 DVSS
port 2 nsew
rlabel metal3 s 774 56560 774 56560 4 DVSS
port 2 nsew
rlabel metal3 s 774 38969 774 38969 4 VDD
port 3 nsew
rlabel metal3 s 774 50334 774 50334 4 VDD
port 3 nsew
<< end >>
