* NGSPICE file created from CP_LF_mag_flat.ext - technology: gf180mcuC

.subckt CP_mag_flat VSS VCNTL PU PD IPD_ IPD+ VDD
X0 VDD IPD_.t0 IPD_.t1 VDD.t9 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.56u
X1 IPD_ IPD_.t2 VDD.t8 VDD.t7 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.56u
X2 IPD+ IPD+.t2 VSS.t9 VSS.t8 nfet_03v3 ad=92.8f pd=0.92u as=0.158p ps=1.64u w=0.28u l=0.56u
X3 inv_0.OUT PU.t0 VSS.t11 VSS.t10 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X4 a_1365_994# PD.t0 VCNTL.t3 VSS.t12 nfet_03v3 ad=0.158p pd=1.64u as=92.8f ps=0.92u w=0.28u l=0.56u
X5 a_1365_994# IPD+.t5 VSS.t7 VSS.t6 nfet_03v3 ad=92.8f pd=0.92u as=92.8f ps=0.92u w=0.28u l=0.56u
X6 VDD IPD_.t5 a_1358_1409# VDD.t4 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.56u
X7 a_1358_1409# IPD_.t6 VDD.t3 VDD.t2 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.56u
X8 a_1358_1409# inv_0.OUT VCNTL.t1 VDD.t1 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.56u
X9 VCNTL PD.t1 a_1365_994# VSS.t13 nfet_03v3 ad=92.8f pd=0.92u as=0.158p ps=1.64u w=0.28u l=0.56u
X10 inv_0.OUT PU.t1 VDD.t13 VDD.t12 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X11 VCNTL inv_0.OUT a_1358_1409# VDD.t0 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.56u
X12 VSS IPD+.t0 IPD+.t1 VSS.t2 nfet_03v3 ad=92.8f pd=0.92u as=92.8f ps=0.92u w=0.28u l=0.56u
X13 VSS IPD+.t6 a_1365_994# VSS.t0 nfet_03v3 ad=0.158p pd=1.64u as=92.8f ps=0.92u w=0.28u l=0.56u
R0 IPD_.n0 IPD_.t5 16.5741
R1 IPD_.n2 IPD_.t2 11.4186
R2 IPD_.n1 IPD_.n0 10.5125
R3 IPD_.n0 IPD_.t6 6.06211
R4 IPD_.n1 IPD_.t0 6.06211
R5 IPD_.n2 IPD_.n1 5.27348
R6 IPD_.n5 IPD_.n2 4.21062
R7 IPD_.n4 IPD_.t1 3.6405
R8 IPD_.n4 IPD_.n3 3.6405
R9 IPD_.n7 IPD_.n6 2.2572
R10 IPD_.n7 IPD_.n5 1.93868
R11 IPD_.n5 IPD_.n4 1.64004
R12 IPD_ IPD_.n7 0.00720213
R13 VDD.t4 VDD.n5 768.971
R14 VDD.n5 VDD.t0 677.782
R15 VDD.t2 VDD.t4 387.098
R16 VDD.t0 VDD.t1 386.404
R17 VDD.n6 VDD.t2 261.649
R18 VDD.n9 VDD.t7 213.262
R19 VDD.n6 VDD.t9 125.448
R20 VDD.n8 VDD.t8 6.51327
R21 VDD.n4 VDD.n3 6.51327
R22 VDD.n5 VDD.n4 6.39746
R23 VDD.n7 VDD.n6 6.3005
R24 VDD.n10 VDD.n9 6.3005
R25 VDD VDD.n11 6.3005
R26 VDD VDD.t13 5.21168
R27 VDD.n1 VDD.t3 3.6405
R28 VDD.n1 VDD.n0 3.6405
R29 VDD.n11 VDD.t12 3.58471
R30 VDD.n2 VDD.n1 2.87327
R31 VDD.n8 VDD.n7 0.196412
R32 VDD VDD.n10 0.155141
R33 VDD.n4 VDD 0.115362
R34 VDD VDD.n2 0.100445
R35 VDD.n7 VDD.n2 0.0184006
R36 VDD.n10 VDD.n8 0.00596961
R37 IPD+.n2 IPD+.t6 19.4169
R38 IPD+.n3 IPD+.n2 14.623
R39 IPD+.n4 IPD+.t2 11.2885
R40 IPD+.n4 IPD+.n3 6.54523
R41 IPD+.n1 IPD+.n0 5.4005
R42 IPD+.n1 IPD+.t1 5.4005
R43 IPD+.n5 IPD+.n4 4.10363
R44 IPD+.n5 IPD+.n1 2.6255
R45 IPD+.n7 IPD+.n6 2.27277
R46 IPD+.n7 IPD+.n5 1.84106
R47 IPD+.n2 IPD+.t5 1.8255
R48 IPD+.n3 IPD+.t0 1.8255
R49 IPD+ IPD+.n7 0.022768
R50 VSS.t13 VSS.t12 1187.6
R51 VSS.t2 VSS.t6 1185.67
R52 VSS.t6 VSS.t0 1173.2
R53 VSS.n12 VSS.t10 864.362
R54 VSS.n8 VSS.t8 672.231
R55 VSS.n8 VSS.t2 513.437
R56 VSS.t0 VSS.n7 365.825
R57 VSS.n13 VSS.n12 288.122
R58 VSS.n4 VSS.t13 121.942
R59 VSS.n14 VSS.t11 9.47848
R60 VSS.n5 VSS.n3 8.84542
R61 VSS.n10 VSS.t9 8.84542
R62 VSS.n5 VSS.n4 5.47425
R63 VSS.n1 VSS.n0 5.4005
R64 VSS.n1 VSS.t7 5.4005
R65 VSS.n14 VSS.n13 5.2005
R66 VSS.n9 VSS.n8 5.2005
R67 VSS.n7 VSS.n6 5.2005
R68 VSS.n2 VSS.n1 3.44542
R69 VSS.n11 VSS.n10 2.45271
R70 VSS.n6 VSS 0.174875
R71 VSS.n10 VSS.n9 0.1505
R72 VSS.n9 VSS.n2 0.1305
R73 VSS VSS.n2 0.079875
R74 VSS.n6 VSS.n5 0.02675
R75 VSS VSS.n11 0.0167581
R76 VSS VSS.n14 0.000790323
R77 PU.n0 PU.t1 25.4398
R78 PU.n0 PU.t0 17.6975
R79 PU PU.n0 4.24656
R80 PD.n0 PD.t1 18.5164
R81 PD.n2 PD.n0 5.96897
R82 PD.n0 PD.t0 4.95003
R83 PD.n2 PD.n1 2.26661
R84 PD PD.n2 0.0166053
R85 VCNTL.n2 VCNTL.n1 5.4005
R86 VCNTL.n2 VCNTL.t3 5.4005
R87 VCNTL.n5 VCNTL.n2 3.71064
R88 VCNTL.n4 VCNTL.t1 3.6405
R89 VCNTL.n4 VCNTL.n3 3.6405
R90 VCNTL VCNTL.n0 2.2555
R91 VCNTL.n5 VCNTL.n4 1.6852
R92 VCNTL VCNTL.n5 1.33738
C0 a_1365_994# PD 0.144f
C1 PU VDD 0.195f
C2 IPD_ PU 0.0872f
C3 a_1365_994# PU 2.18e-19
C4 IPD+ VCNTL 2.35e-19
C5 a_1358_1409# VDD 0.768f
C6 IPD+ inv_0.OUT 0.127f
C7 IPD_ a_1358_1409# 0.111f
C8 a_1365_994# a_1358_1409# 0.279f
C9 VCNTL inv_0.OUT 0.281f
C10 IPD+ PD 0.49f
C11 IPD_ VDD 1.02f
C12 a_1365_994# VDD 0.00964f
C13 IPD+ PU 0.0527f
C14 VCNTL PD 0.0331f
C15 IPD_ a_1365_994# 0.00945f
C16 PD inv_0.OUT 0.164f
C17 PU inv_0.OUT 0.121f
C18 IPD+ a_1358_1409# 3.09e-19
C19 VCNTL a_1358_1409# 0.215f
C20 PU PD 9.18e-19
C21 IPD+ VDD 0.0131f
C22 a_1358_1409# inv_0.OUT 0.183f
C23 IPD_ IPD+ 0.145f
C24 a_1365_994# IPD+ 0.0463f
C25 VCNTL VDD 0.0486f
C26 PD a_1358_1409# 0.00441f
C27 IPD_ VCNTL 0.00567f
C28 a_1365_994# VCNTL 0.15f
C29 inv_0.OUT VDD 0.559f
C30 IPD_ inv_0.OUT 0.27f
C31 PU a_1358_1409# 1.69e-20
C32 a_1365_994# inv_0.OUT 0.211f
C33 PD VDD 0.00174f
C34 IPD_ PD 9.39e-19
C35 PD VSS 1.69f
C36 IPD+ VSS 1.65f
C37 VCNTL VSS 0.223f
C38 IPD_ VSS 0.747f
C39 a_1365_994# VSS 0.458f
C40 a_1358_1409# VSS 0.104f
C41 inv_0.OUT VSS 0.646f
C42 PU VSS 0.368f
C43 VDD VSS 4.35f
.ends

