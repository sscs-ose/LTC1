magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -3455 -2045 3455 2045
<< psubdiff >>
rect -1455 23 1455 45
rect -1455 -23 -1433 23
rect 1433 -23 1455 23
rect -1455 -45 1455 -23
<< psubdiffcont >>
rect -1433 -23 1433 23
<< metal1 >>
rect -1444 23 1444 34
rect -1444 -23 -1433 23
rect 1433 -23 1444 23
rect -1444 -34 1444 -23
<< end >>
