magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2127 -2235 2772 2615
<< polysilicon >>
rect 25 339 599 615
rect 25 -235 599 41
<< metal1 >>
rect -127 -134 772 514
use M1_POLY2_CDNS_69033583165701  M1_POLY2_CDNS_69033583165701_0
timestamp 1713338890
transform 1 0 557 0 1 474
box -42 -42 42 42
use M1_POLY2_CDNS_69033583165701  M1_POLY2_CDNS_69033583165701_1
timestamp 1713338890
transform 1 0 67 0 1 474
box -42 -42 42 42
use M1_POLY2_CDNS_69033583165701  M1_POLY2_CDNS_69033583165701_2
timestamp 1713338890
transform 1 0 67 0 -1 -100
box -42 -42 42 42
use M1_POLY2_CDNS_69033583165701  M1_POLY2_CDNS_69033583165701_3
timestamp 1713338890
transform 1 0 557 0 -1 -100
box -42 -42 42 42
use M1_PSUB_CDNS_69033583165700  M1_PSUB_CDNS_69033583165700_0
timestamp 1713338890
transform 1 0 308 0 1 190
box -280 -45 280 45
use M1_PSUB_CDNS_69033583165700  M1_PSUB_CDNS_69033583165700_1
timestamp 1713338890
transform 1 0 308 0 -1 190
box -280 -45 280 45
<< end >>
