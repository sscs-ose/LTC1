magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1232 -1090 1232 1090
<< metal2 >>
rect -232 85 232 90
rect -232 57 -227 85
rect -199 57 -156 85
rect -128 57 -85 85
rect -57 57 -14 85
rect 14 57 57 85
rect 85 57 128 85
rect 156 57 199 85
rect 227 57 232 85
rect -232 14 232 57
rect -232 -14 -227 14
rect -199 -14 -156 14
rect -128 -14 -85 14
rect -57 -14 -14 14
rect 14 -14 57 14
rect 85 -14 128 14
rect 156 -14 199 14
rect 227 -14 232 14
rect -232 -57 232 -14
rect -232 -85 -227 -57
rect -199 -85 -156 -57
rect -128 -85 -85 -57
rect -57 -85 -14 -57
rect 14 -85 57 -57
rect 85 -85 128 -57
rect 156 -85 199 -57
rect 227 -85 232 -57
rect -232 -90 232 -85
<< via2 >>
rect -227 57 -199 85
rect -156 57 -128 85
rect -85 57 -57 85
rect -14 57 14 85
rect 57 57 85 85
rect 128 57 156 85
rect 199 57 227 85
rect -227 -14 -199 14
rect -156 -14 -128 14
rect -85 -14 -57 14
rect -14 -14 14 14
rect 57 -14 85 14
rect 128 -14 156 14
rect 199 -14 227 14
rect -227 -85 -199 -57
rect -156 -85 -128 -57
rect -85 -85 -57 -57
rect -14 -85 14 -57
rect 57 -85 85 -57
rect 128 -85 156 -57
rect 199 -85 227 -57
<< metal3 >>
rect -232 85 232 90
rect -232 57 -227 85
rect -199 57 -156 85
rect -128 57 -85 85
rect -57 57 -14 85
rect 14 57 57 85
rect 85 57 128 85
rect 156 57 199 85
rect 227 57 232 85
rect -232 14 232 57
rect -232 -14 -227 14
rect -199 -14 -156 14
rect -128 -14 -85 14
rect -57 -14 -14 14
rect 14 -14 57 14
rect 85 -14 128 14
rect 156 -14 199 14
rect 227 -14 232 14
rect -232 -57 232 -14
rect -232 -85 -227 -57
rect -199 -85 -156 -57
rect -128 -85 -85 -57
rect -57 -85 -14 -57
rect 14 -85 57 -57
rect 85 -85 128 -57
rect 156 -85 199 -57
rect 227 -85 232 -57
rect -232 -90 232 -85
<< end >>
