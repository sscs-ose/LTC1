magic
tech gf180mcuC
magscale 1 10
timestamp 1698660008
<< nwell >>
rect 1677 1096 1832 2749
rect 3436 1096 3644 2749
rect 5251 1096 5512 2748
rect 3438 -4064 3644 -932
rect 5251 -4064 5511 -933
rect 1653 -6660 1892 -6091
rect 1678 -7745 1831 -6660
rect 3438 -7744 3645 -6092
rect 5250 -7747 5512 -6093
<< metal1 >>
rect -2960 2568 -2171 2740
rect -611 2573 178 2745
rect 1675 2575 1840 2749
rect 3435 2575 3664 2749
rect 5249 2575 5528 2748
rect 7116 2574 7118 2748
rect 7503 2731 7676 2748
rect 7503 2675 7507 2731
rect 7563 2675 7617 2731
rect 7673 2675 7676 2731
rect 7503 2621 7676 2675
rect 7503 2565 7507 2621
rect 7563 2565 7617 2621
rect 7673 2565 7676 2621
rect 7503 2511 7676 2565
rect 7503 2455 7507 2511
rect 7563 2455 7617 2511
rect 7673 2455 7676 2511
rect 7503 2443 7676 2455
rect 2995 1319 3070 1331
rect 2995 1265 3002 1319
rect 3056 1265 3070 1319
rect -5214 1204 -5093 1208
rect -5214 1174 -5197 1204
rect -5352 1147 -5197 1174
rect -5140 1147 -5093 1204
rect -3028 1161 -2840 1172
rect -5352 1117 -5093 1147
rect -5214 1094 -5093 1117
rect -3030 1105 -3020 1161
rect -2964 1105 -2909 1161
rect -2853 1105 -2840 1161
rect -3028 1097 -2840 1105
rect -637 1170 -437 1179
rect -637 1169 -505 1170
rect -637 1113 -625 1169
rect -569 1114 -505 1169
rect -449 1114 -437 1170
rect 43 1134 45 1188
rect -569 1113 -437 1114
rect -637 1104 -437 1113
rect 46 1100 125 1214
rect -5214 1037 -5197 1094
rect -5140 1037 -5093 1094
rect -5214 1026 -5093 1037
rect 46 1044 58 1100
rect 114 1044 125 1100
rect 46 1028 125 1044
rect 438 1099 517 1221
rect 1724 1158 1770 1180
rect 438 1045 453 1099
rect 507 1045 517 1099
rect 438 1033 517 1045
rect -5040 969 -4978 977
rect -5111 941 -4887 969
rect -5114 885 -5104 941
rect -5048 885 -4994 941
rect -4938 885 -4887 941
rect -2689 930 -2481 974
rect -5111 853 -4887 885
rect -2691 874 -2681 930
rect -2625 874 -2571 930
rect -2515 874 -2481 930
rect -5197 711 -5101 714
rect -5197 661 -5170 711
rect -5368 654 -5170 661
rect -5113 654 -5101 711
rect -5368 604 -5101 654
rect -5197 601 -5101 604
rect -5197 544 -5170 601
rect -5113 544 -5101 601
rect -5197 540 -5101 544
rect -5040 -615 -4978 853
rect -2689 830 -2481 874
rect -86 896 8 945
rect -86 821 -40 896
rect -102 805 -13 821
rect -102 748 -84 805
rect -27 748 -13 805
rect -102 732 -13 748
rect -2973 161 -2265 162
rect -3054 -10 -2265 161
rect -1019 53 -1009 109
rect -953 53 -943 109
rect -5041 -623 -4935 -615
rect -5041 -679 -5016 -623
rect -4960 -679 -4935 -623
rect -5041 -733 -4935 -679
rect -5041 -789 -5016 -733
rect -4960 -789 -4935 -733
rect -5041 -804 -4935 -789
rect -2601 -624 -2501 -611
rect -2601 -680 -2582 -624
rect -2526 -680 -2501 -624
rect -2601 -734 -2501 -680
rect -2601 -790 -2582 -734
rect -2526 -790 -2501 -734
rect -5194 -914 -5099 -878
rect -5194 -965 -5181 -914
rect -5324 -972 -5181 -965
rect -5123 -972 -5099 -914
rect -5324 -1024 -5099 -972
rect -5324 -1025 -5181 -1024
rect -5194 -1082 -5181 -1025
rect -5123 -1082 -5099 -1024
rect -5194 -1094 -5099 -1082
rect -5189 -1391 -5094 -1381
rect -5189 -1439 -5164 -1391
rect -5254 -1447 -5164 -1439
rect -5108 -1447 -5094 -1391
rect -5254 -1493 -5094 -1447
rect -5189 -1501 -5094 -1493
rect -5189 -1557 -5164 -1501
rect -5108 -1557 -5094 -1501
rect -5189 -1567 -5094 -1557
rect -5209 -3275 -5121 -3268
rect -5209 -3323 -5193 -3275
rect -5288 -3331 -5193 -3323
rect -5137 -3331 -5121 -3275
rect -5288 -3377 -5121 -3331
rect -5209 -3385 -5121 -3377
rect -5209 -3441 -5193 -3385
rect -5137 -3441 -5121 -3385
rect -5209 -3458 -5121 -3441
rect -5189 -3959 -5107 -3947
rect -5336 -3960 -5107 -3959
rect -5336 -4014 -5177 -3960
rect -5189 -4018 -5177 -4014
rect -5119 -4018 -5107 -3960
rect -5189 -4070 -5107 -4018
rect -5189 -4128 -5177 -4070
rect -5119 -4128 -5107 -4070
rect -5189 -4135 -5107 -4128
rect -5040 -4199 -4978 -804
rect -2601 -806 -2501 -790
rect -3049 -958 -2839 -948
rect -630 -950 -436 -942
rect -3049 -1014 -3039 -958
rect -2983 -959 -2839 -958
rect -2983 -1014 -2921 -959
rect -3049 -1015 -2921 -1014
rect -2865 -1015 -2839 -959
rect -631 -1006 -621 -950
rect -565 -1006 -502 -950
rect -446 -1006 -436 -950
rect -3049 -1025 -2839 -1015
rect -630 -1017 -436 -1006
rect -98 -983 -40 732
rect 1708 415 1788 1158
rect 2995 1142 3070 1265
rect 3385 1320 3462 1332
rect 3385 1264 3395 1320
rect 3451 1264 3462 1320
rect 3385 1135 3462 1264
rect 3620 1320 3696 1332
rect 3620 1264 3631 1320
rect 3687 1264 3696 1320
rect 3620 1134 3696 1264
rect 6673 1328 6750 1339
rect 6673 1274 6685 1328
rect 6739 1274 6750 1328
rect 5305 1165 5445 1179
rect 5284 1153 5445 1165
rect 5284 1104 5461 1153
rect 6673 1142 6750 1274
rect 7065 1319 7142 1357
rect 7065 1263 7075 1319
rect 7131 1263 7142 1319
rect 7065 1134 7142 1263
rect 3484 895 3575 945
rect 3484 466 3530 895
rect 1708 360 1721 415
rect 1776 360 1788 415
rect 1708 305 1788 360
rect 1708 250 1721 305
rect 1776 250 1788 305
rect 3470 454 3543 466
rect 3470 400 3480 454
rect 3534 400 3543 454
rect 5284 415 5364 1104
rect 7113 915 7234 944
rect 7113 884 7161 915
rect 7144 858 7161 884
rect 7218 858 7234 915
rect 7144 805 7234 858
rect 7144 748 7161 805
rect 7218 748 7234 805
rect 7144 739 7234 748
rect 7505 791 7676 2443
rect 7505 774 7678 791
rect 7505 718 7509 774
rect 7565 718 7619 774
rect 7675 718 7678 774
rect 7505 664 7678 718
rect 7505 608 7509 664
rect 7565 608 7619 664
rect 7675 608 7678 664
rect 7505 554 7678 608
rect 7505 498 7509 554
rect 7565 498 7619 554
rect 7675 498 7678 554
rect 7505 486 7678 498
rect 3470 344 3543 400
rect 3470 290 3480 344
rect 3534 290 3543 344
rect 3470 277 3543 290
rect 5285 402 5365 415
rect 5285 346 5297 402
rect 5353 346 5365 402
rect 5285 292 5365 346
rect 1708 238 1788 250
rect 5285 236 5297 292
rect 5353 236 5365 292
rect 5285 224 5365 236
rect 70 58 80 114
rect 136 58 146 114
rect 342 -159 352 -103
rect 408 -159 418 -103
rect 467 -161 477 -105
rect 533 -161 543 -105
rect 582 -161 592 -105
rect 648 -161 658 -105
rect 709 -160 719 -104
rect 775 -160 785 -104
rect 839 -158 849 -102
rect 905 -158 915 -102
rect 991 -354 1178 -341
rect 991 -408 1004 -354
rect 1058 -408 1114 -354
rect 1168 -408 1178 -354
rect 991 -420 1178 -408
rect -98 -1029 60 -983
rect 1008 -984 1054 -420
rect 1326 -491 1407 -481
rect 1326 -548 1338 -491
rect 1395 -548 1407 -491
rect 1326 -601 1407 -548
rect 1106 -618 1178 -607
rect 1106 -672 1115 -618
rect 1169 -672 1178 -618
rect 1326 -658 1338 -601
rect 1395 -658 1407 -601
rect 1326 -670 1407 -658
rect 1106 -728 1178 -672
rect 1106 -782 1115 -728
rect 1169 -782 1178 -728
rect 1106 -795 1178 -782
rect -98 -1030 51 -1029
rect 925 -1030 1054 -984
rect -98 -1509 -40 -1030
rect -126 -1519 -31 -1509
rect -126 -1575 -101 -1519
rect -45 -1575 -31 -1519
rect -126 -1629 -31 -1575
rect -126 -1685 -101 -1629
rect -45 -1685 -31 -1629
rect 442 -1634 452 -1578
rect 508 -1634 518 -1578
rect 577 -1633 587 -1577
rect 643 -1633 653 -1577
rect 707 -1632 717 -1576
rect 773 -1632 783 -1576
rect 850 -1633 860 -1577
rect 916 -1633 926 -1577
rect -126 -1695 -31 -1685
rect -340 -2019 -150 -2011
rect -340 -2075 -328 -2019
rect -272 -2075 -218 -2019
rect -162 -2075 -150 -2019
rect -340 -2082 -150 -2075
rect -3010 -2586 -2435 -2419
rect -1090 -2527 -1080 -2471
rect -1024 -2527 -1014 -2471
rect -3050 -3997 -2840 -3988
rect -3050 -4053 -3040 -3997
rect -2984 -4053 -2919 -3997
rect -2863 -4053 -2840 -3997
rect -3050 -4063 -2840 -4053
rect -673 -3989 -437 -3981
rect -673 -3990 -520 -3989
rect -673 -4046 -658 -3990
rect -602 -4045 -520 -3990
rect -464 -4045 -437 -3989
rect -602 -4046 -437 -4045
rect -673 -4057 -437 -4046
rect -5055 -4209 -4960 -4199
rect -5055 -4265 -5030 -4209
rect -4974 -4265 -4960 -4209
rect -5055 -4319 -4960 -4265
rect -5055 -4375 -5030 -4319
rect -4974 -4375 -4960 -4319
rect -5055 -4385 -4960 -4375
rect -2620 -4200 -2525 -4190
rect -2620 -4256 -2595 -4200
rect -2539 -4256 -2525 -4200
rect -2620 -4310 -2525 -4256
rect -2620 -4366 -2595 -4310
rect -2539 -4366 -2525 -4310
rect -2620 -4376 -2525 -4366
rect -340 -4336 -151 -4324
rect -5235 -5518 -5162 -5506
rect -5376 -5575 -5225 -5518
rect -5168 -5575 -5162 -5518
rect -5235 -5628 -5162 -5575
rect -5235 -5685 -5225 -5628
rect -5168 -5685 -5162 -5628
rect -5235 -5697 -5162 -5685
rect -5040 -5768 -4978 -4385
rect -340 -4396 -331 -4336
rect -271 -4396 -218 -4336
rect -158 -4396 -151 -4336
rect -340 -4408 -151 -4396
rect -2969 -5173 -2378 -5000
rect -1199 -5106 -1189 -5050
rect -1133 -5106 -1123 -5050
rect -98 -5642 -40 -1695
rect 7 -2019 92 -2007
rect 7 -2075 24 -2019
rect 80 -2075 92 -2019
rect 7 -2129 92 -2075
rect 7 -2185 24 -2129
rect 80 -2185 92 -2129
rect 7 -2195 92 -2185
rect 746 -2170 935 -2155
rect 17 -2223 76 -2195
rect 746 -2224 756 -2170
rect 810 -2224 866 -2170
rect 920 -2224 935 -2170
rect 746 -2238 935 -2224
rect 385 -3103 395 -3047
rect 451 -3103 461 -3047
rect 503 -3101 513 -3045
rect 569 -3101 579 -3045
rect 627 -3100 637 -3044
rect 693 -3100 703 -3044
rect 736 -3100 746 -3044
rect 802 -3100 812 -3044
rect 856 -3102 866 -3046
rect 922 -3102 932 -3046
rect 749 -3921 941 -3906
rect 23 -4207 69 -3924
rect 75 -3970 83 -3924
rect 749 -3975 765 -3921
rect 819 -3975 875 -3921
rect 929 -3975 941 -3921
rect 749 -3987 941 -3975
rect 7 -4223 86 -4207
rect 7 -4277 19 -4223
rect 73 -4277 86 -4223
rect 7 -4333 86 -4277
rect 7 -4387 19 -4333
rect 73 -4387 86 -4333
rect 7 -4399 86 -4387
rect 1008 -4500 1054 -1030
rect 1118 -2153 1165 -795
rect 1213 -860 1293 -848
rect 1213 -916 1225 -860
rect 1281 -916 1293 -860
rect 1213 -970 1293 -916
rect 1213 -1026 1225 -970
rect 1281 -1026 1293 -970
rect 1213 -1033 1293 -1026
rect 1225 -1898 1272 -1033
rect 1216 -1910 1287 -1898
rect 1216 -1964 1226 -1910
rect 1280 -1964 1287 -1910
rect 1216 -2020 1287 -1964
rect 1216 -2074 1226 -2020
rect 1280 -2074 1287 -2020
rect 1216 -2087 1287 -2074
rect 1104 -2165 1180 -2153
rect 1104 -2219 1115 -2165
rect 1169 -2219 1180 -2165
rect 1104 -2275 1180 -2219
rect 1104 -2329 1115 -2275
rect 1169 -2329 1180 -2275
rect 1104 -2340 1180 -2329
rect 1118 -4072 1165 -2340
rect 1103 -4085 1180 -4072
rect 1103 -4139 1115 -4085
rect 1169 -4139 1180 -4085
rect 1103 -4195 1180 -4139
rect 1103 -4249 1115 -4195
rect 1169 -4249 1180 -4195
rect 1103 -4263 1180 -4249
rect 1226 -4215 1272 -2087
rect 1344 -3796 1391 -670
rect 1469 -1389 1569 79
rect 1673 -5 1841 169
rect 3433 -6 3660 169
rect 5250 -5 5519 168
rect 7118 -6 7412 168
rect 2333 -71 2381 -51
rect 2320 -86 2396 -71
rect 2320 -140 2330 -86
rect 2384 -140 2396 -86
rect 2320 -154 2396 -140
rect 2632 -89 2714 -85
rect 2632 -145 2646 -89
rect 2702 -145 2714 -89
rect 2632 -147 2714 -145
rect 2953 -89 3035 -85
rect 2953 -145 2966 -89
rect 3022 -145 3035 -89
rect 3275 -88 3357 -83
rect 3275 -144 3288 -88
rect 3344 -144 3357 -88
rect 3275 -145 3357 -144
rect 3718 -90 3804 -80
rect 2953 -147 3035 -145
rect 3718 -146 3735 -90
rect 3791 -146 3804 -90
rect 3718 -151 3804 -146
rect 4041 -91 4127 -80
rect 4041 -147 4057 -91
rect 4113 -147 4127 -91
rect 4361 -88 4447 -75
rect 4361 -144 4378 -88
rect 4434 -144 4447 -88
rect 4361 -146 4447 -144
rect 4686 -99 4768 -86
rect 4041 -151 4127 -147
rect 4686 -153 4699 -99
rect 4753 -153 4768 -99
rect 4686 -164 4768 -153
rect 5384 -460 5457 -444
rect 5384 -514 5394 -460
rect 5448 -514 5457 -460
rect 5384 -570 5457 -514
rect 5384 -624 5394 -570
rect 5448 -624 5457 -570
rect 1623 -729 1856 -718
rect 1623 -783 1635 -729
rect 1689 -783 1745 -729
rect 1799 -783 1856 -729
rect 1623 -795 1856 -783
rect 5227 -733 5337 -720
rect 5227 -789 5269 -733
rect 5325 -789 5337 -733
rect 5384 -733 5457 -624
rect 5384 -782 5487 -733
rect 7066 -747 7145 -731
rect 7066 -754 7078 -747
rect 5227 -801 5337 -789
rect 5255 -843 5337 -801
rect 5255 -899 5269 -843
rect 5325 -899 5337 -843
rect 5255 -914 5337 -899
rect 6661 -801 7078 -754
rect 7132 -801 7145 -747
rect 6661 -857 7145 -801
rect 6661 -911 7078 -857
rect 7132 -911 7145 -857
rect 3492 -1065 3604 -941
rect 6661 -950 7145 -911
rect 6661 -967 7146 -950
rect 3492 -1119 3512 -1065
rect 3566 -1119 3604 -1065
rect 3492 -1175 3604 -1119
rect 3492 -1229 3512 -1175
rect 3566 -1229 3604 -1175
rect 3492 -1254 3604 -1229
rect 5461 -1101 5564 -970
rect 5461 -1157 5498 -1101
rect 5554 -1157 5564 -1101
rect 5461 -1254 5564 -1157
rect 5878 -1102 5956 -980
rect 6661 -990 7078 -967
rect 7066 -1021 7078 -990
rect 7132 -1021 7146 -967
rect 7066 -1034 7146 -1021
rect 5878 -1156 5893 -1102
rect 5947 -1156 5956 -1102
rect 5878 -1175 5956 -1156
rect 1458 -1391 1584 -1389
rect 1458 -1447 1492 -1391
rect 1548 -1447 1584 -1391
rect 1458 -1501 1584 -1447
rect 1458 -1557 1492 -1501
rect 1548 -1557 1584 -1501
rect 1458 -1611 1584 -1557
rect 1458 -1667 1492 -1611
rect 1548 -1667 1584 -1611
rect 1458 -1674 1584 -1667
rect 1682 -2550 1935 -2450
rect 1682 -2850 1782 -2550
rect 3416 -2586 3682 -2411
rect 5246 -2585 5515 -2412
rect 1666 -2861 1794 -2850
rect 1666 -2917 1702 -2861
rect 1758 -2917 1794 -2861
rect 1666 -2971 1794 -2917
rect 1666 -3027 1702 -2971
rect 1758 -3027 1794 -2971
rect 1666 -3081 1794 -3027
rect 1666 -3137 1702 -3081
rect 1758 -3137 1794 -3081
rect 1666 -3143 1794 -3137
rect 1323 -3808 1405 -3796
rect 1323 -3865 1333 -3808
rect 1390 -3865 1405 -3808
rect 1323 -3918 1405 -3865
rect 1323 -3975 1333 -3918
rect 1390 -3975 1405 -3918
rect 1323 -3989 1405 -3975
rect 3520 -3823 3602 -3810
rect 3520 -3881 3533 -3823
rect 3591 -3881 3602 -3823
rect 3520 -3933 3602 -3881
rect 3520 -3980 3533 -3933
rect 3390 -3991 3533 -3980
rect 3591 -3980 3602 -3933
rect 5487 -3841 5564 -3822
rect 5487 -3897 5498 -3841
rect 5554 -3897 5564 -3841
rect 3591 -3991 3644 -3980
rect 3390 -4055 3644 -3991
rect 5487 -4027 5564 -3897
rect 5876 -3842 5956 -3836
rect 5876 -3896 5889 -3842
rect 5943 -3896 5956 -3842
rect 5876 -4018 5956 -3896
rect 7084 -3977 7162 -3964
rect 7084 -3995 7096 -3977
rect 6675 -4031 7096 -3995
rect 7150 -4031 7162 -3977
rect 5244 -4099 5322 -4083
rect 5244 -4155 5253 -4099
rect 5309 -4155 5322 -4099
rect 5244 -4202 5322 -4155
rect 6675 -4087 7162 -4031
rect 6675 -4141 7096 -4087
rect 7150 -4141 7162 -4087
rect 6675 -4197 7162 -4141
rect 5244 -4203 5324 -4202
rect 5243 -4209 5324 -4203
rect 1226 -4264 1801 -4215
rect 5243 -4265 5253 -4209
rect 5309 -4265 5324 -4209
rect 5243 -4276 5324 -4265
rect 5421 -4329 5470 -4215
rect 6675 -4231 7096 -4197
rect 7084 -4251 7096 -4231
rect 7150 -4251 7162 -4197
rect 7084 -4268 7162 -4251
rect 5412 -4343 5484 -4329
rect 5412 -4397 5419 -4343
rect 5473 -4397 5484 -4343
rect 5412 -4453 5484 -4397
rect 991 -4512 1180 -4500
rect 991 -4566 1004 -4512
rect 1058 -4566 1114 -4512
rect 1168 -4566 1180 -4512
rect 5412 -4507 5419 -4453
rect 5473 -4507 5484 -4453
rect 5412 -4522 5484 -4507
rect 991 -4579 1180 -4566
rect 311 -5020 405 -4597
rect 2625 -4832 2717 -4822
rect 2327 -4837 2403 -4833
rect 2327 -4891 2337 -4837
rect 2391 -4891 2403 -4837
rect 2327 -4906 2403 -4891
rect 2625 -4888 2645 -4832
rect 2701 -4888 2717 -4832
rect 2625 -4900 2717 -4888
rect 2952 -4845 3037 -4835
rect 2952 -4901 2966 -4845
rect 3022 -4901 3037 -4845
rect 2952 -4910 3037 -4901
rect 3271 -4848 3349 -4837
rect 3271 -4904 3283 -4848
rect 3339 -4904 3349 -4848
rect 3271 -4916 3349 -4904
rect 3732 -4848 3813 -4834
rect 3732 -4904 3745 -4848
rect 3801 -4904 3813 -4848
rect 3732 -4920 3813 -4904
rect 4044 -4846 4125 -4828
rect 4044 -4902 4057 -4846
rect 4113 -4902 4125 -4846
rect 4044 -4914 4125 -4902
rect 4364 -4843 4445 -4830
rect 4364 -4899 4377 -4843
rect 4433 -4899 4445 -4843
rect 4364 -4916 4445 -4899
rect 4683 -4843 4771 -4828
rect 4683 -4897 4699 -4843
rect 4753 -4897 4771 -4843
rect 4683 -4909 4771 -4897
rect 76 -5106 86 -5050
rect 142 -5106 152 -5050
rect 1674 -5165 1837 -4990
rect 3437 -5164 3653 -4991
rect 7245 -4992 7412 -6
rect 5247 -5166 5522 -4992
rect 7114 -5166 7412 -4992
rect 7505 -2281 7676 486
rect 7747 -746 7936 -730
rect 7747 -802 7758 -746
rect 7814 -802 7868 -746
rect 7924 -802 7936 -746
rect 7747 -856 7936 -802
rect 7747 -912 7758 -856
rect 7814 -912 7868 -856
rect 7924 -912 7936 -856
rect 7747 -966 7936 -912
rect 7747 -1022 7758 -966
rect 7814 -1022 7868 -966
rect 7924 -1022 7936 -966
rect 7747 -1034 7936 -1022
rect 7505 -2298 7678 -2281
rect 7505 -2354 7509 -2298
rect 7565 -2354 7619 -2298
rect 7675 -2354 7678 -2298
rect 7505 -2408 7678 -2354
rect 7505 -2464 7509 -2408
rect 7565 -2464 7619 -2408
rect 7675 -2464 7678 -2408
rect 7505 -2518 7678 -2464
rect 7505 -2574 7509 -2518
rect 7565 -2574 7619 -2518
rect 7675 -2574 7678 -2518
rect 7505 -2586 7678 -2574
rect 3470 -5310 3543 -5297
rect 1715 -5337 1795 -5324
rect 1715 -5392 1728 -5337
rect 1783 -5392 1795 -5337
rect 1715 -5447 1795 -5392
rect 1715 -5502 1728 -5447
rect 1783 -5502 1795 -5447
rect 3470 -5364 3480 -5310
rect 3534 -5364 3543 -5310
rect 3470 -5420 3543 -5364
rect 3470 -5474 3480 -5420
rect 3534 -5474 3543 -5420
rect 3470 -5493 3543 -5474
rect 5321 -5342 5408 -5327
rect 5321 -5398 5335 -5342
rect 5391 -5398 5408 -5342
rect 5321 -5452 5408 -5398
rect -97 -5646 -16 -5642
rect -97 -5703 -85 -5646
rect -28 -5703 -16 -5646
rect -97 -5756 -16 -5703
rect -5044 -5778 -4949 -5768
rect -5044 -5834 -5019 -5778
rect -4963 -5834 -4949 -5778
rect -5044 -5888 -4949 -5834
rect -5044 -5944 -5019 -5888
rect -4963 -5944 -4949 -5888
rect -5044 -5954 -4949 -5944
rect -2626 -5782 -2531 -5772
rect -2626 -5838 -2601 -5782
rect -2545 -5838 -2531 -5782
rect -97 -5813 -85 -5756
rect -28 -5813 -16 -5756
rect -97 -5823 -16 -5813
rect -2626 -5892 -2531 -5838
rect -2626 -5948 -2601 -5892
rect -2545 -5948 -2531 -5892
rect -86 -5892 -40 -5823
rect -86 -5941 -6 -5892
rect -5040 -5986 -4978 -5954
rect -2626 -5958 -2531 -5948
rect 47 -6041 124 -6027
rect -5128 -6049 -5051 -6041
rect -5128 -6106 -5119 -6049
rect -5062 -6106 -5051 -6049
rect 47 -6097 57 -6041
rect 113 -6097 124 -6041
rect -5128 -6157 -5051 -6106
rect -3046 -6117 -2840 -6109
rect -641 -6110 -437 -6102
rect -5382 -6159 -5051 -6157
rect -5382 -6216 -5119 -6159
rect -5062 -6216 -5051 -6159
rect -3048 -6173 -3038 -6117
rect -2982 -6173 -2908 -6117
rect -2852 -6173 -2840 -6117
rect -643 -6166 -633 -6110
rect -577 -6166 -508 -6110
rect -452 -6166 -437 -6110
rect -3046 -6184 -2840 -6173
rect -641 -6177 -437 -6166
rect -5128 -6228 -5051 -6216
rect 47 -6220 124 -6097
rect 439 -6040 516 -6028
rect 439 -6096 448 -6040
rect 504 -6096 516 -6040
rect 439 -6154 516 -6096
rect 1715 -6177 1795 -5502
rect 3484 -5892 3530 -5493
rect 5321 -5508 5335 -5452
rect 5391 -5508 5408 -5452
rect 3484 -5941 3579 -5892
rect 2990 -6041 3070 -6034
rect 2990 -6095 3002 -6041
rect 3056 -6095 3070 -6041
rect 2990 -6217 3070 -6095
rect 3620 -6040 3697 -6028
rect 3620 -6096 3631 -6040
rect 3687 -6096 3697 -6040
rect 4012 -6041 4089 -6033
rect 3620 -6219 3697 -6096
rect 4011 -6097 4021 -6041
rect 4077 -6097 4089 -6041
rect 4012 -6217 4089 -6097
rect 5321 -6101 5408 -5508
rect 7085 -5756 7176 -5742
rect 7085 -5810 7108 -5756
rect 7162 -5810 7176 -5756
rect 7085 -5866 7176 -5810
rect 7085 -5920 7108 -5866
rect 7162 -5920 7176 -5866
rect 7085 -5944 7176 -5920
rect 6673 -6042 6750 -6030
rect 6673 -6096 6682 -6042
rect 6736 -6096 6750 -6042
rect 5256 -6176 5539 -6101
rect 6673 -6150 6750 -6096
rect 5285 -6177 5531 -6176
rect 7066 -6261 7143 -6130
rect 7066 -6317 7075 -6261
rect 7131 -6317 7143 -6261
rect 7066 -6334 7143 -6317
rect 7505 -7441 7676 -2586
rect 7753 -3963 7936 -1034
rect 7744 -3976 7936 -3963
rect 7744 -4032 7753 -3976
rect 7809 -4032 7863 -3976
rect 7919 -4032 7936 -3976
rect 7744 -4086 7936 -4032
rect 7744 -4142 7753 -4086
rect 7809 -4142 7863 -4086
rect 7919 -4142 7936 -4086
rect 7744 -4196 7936 -4142
rect 7744 -4252 7753 -4196
rect 7809 -4252 7863 -4196
rect 7919 -4252 7936 -4196
rect 7744 -4267 7936 -4252
rect 7505 -7458 7678 -7441
rect 7505 -7514 7509 -7458
rect 7565 -7514 7619 -7458
rect 7675 -7514 7678 -7458
rect 7505 -7568 7678 -7514
rect 126 -7572 136 -7571
rect -2997 -7752 -2426 -7579
rect -538 -7742 136 -7572
rect 1675 -7745 1838 -7570
rect 3434 -7747 3656 -7571
rect 5247 -7745 5533 -7572
rect 7505 -7624 7509 -7568
rect 7565 -7624 7619 -7568
rect 7675 -7624 7678 -7568
rect 7505 -7678 7678 -7624
rect 7505 -7734 7509 -7678
rect 7565 -7734 7619 -7678
rect 7675 -7734 7678 -7678
rect 7505 -7746 7678 -7734
<< via1 >>
rect 6507 2635 6561 2687
rect 6627 2635 6681 2687
rect 6747 2635 6801 2687
rect 6867 2635 6921 2687
rect 6987 2635 7041 2687
rect 7507 2675 7563 2731
rect 7617 2675 7673 2731
rect 7507 2565 7563 2621
rect 7617 2565 7673 2621
rect 7507 2455 7563 2511
rect 7617 2455 7673 2511
rect 3002 1265 3056 1319
rect -5197 1147 -5140 1204
rect -3020 1105 -2964 1161
rect -2909 1105 -2853 1161
rect -625 1113 -569 1169
rect -505 1114 -449 1170
rect -5197 1037 -5140 1094
rect 58 1044 114 1100
rect 453 1045 507 1099
rect -5104 885 -5048 941
rect -4994 885 -4938 941
rect -2681 874 -2625 930
rect -2571 874 -2515 930
rect -5170 654 -5113 711
rect -5170 544 -5113 601
rect -84 748 -27 805
rect -1009 53 -953 109
rect -899 53 -843 109
rect -789 53 -733 109
rect -679 53 -623 109
rect -5016 -679 -4960 -623
rect -5016 -789 -4960 -733
rect -2582 -680 -2526 -624
rect -2582 -790 -2526 -734
rect -5181 -972 -5123 -914
rect -5181 -1082 -5123 -1024
rect -5164 -1447 -5108 -1391
rect -5164 -1557 -5108 -1501
rect -5193 -3331 -5137 -3275
rect -5193 -3441 -5137 -3385
rect -5177 -4018 -5119 -3960
rect -5177 -4128 -5119 -4070
rect -3039 -1014 -2983 -958
rect -2921 -1015 -2865 -959
rect -621 -1006 -565 -950
rect -502 -1006 -446 -950
rect 3395 1264 3451 1320
rect 3631 1264 3687 1320
rect 6685 1274 6739 1328
rect 7075 1263 7131 1319
rect 1721 360 1776 415
rect 1721 250 1776 305
rect 3480 400 3534 454
rect 7161 858 7218 915
rect 7161 748 7218 805
rect 7509 718 7565 774
rect 7619 718 7675 774
rect 7509 608 7565 664
rect 7619 608 7675 664
rect 7509 498 7565 554
rect 7619 498 7675 554
rect 3480 290 3534 344
rect 5297 346 5353 402
rect 5297 236 5353 292
rect 80 58 136 114
rect 190 58 246 114
rect 300 58 356 114
rect 410 58 466 114
rect 520 58 576 114
rect 352 -159 408 -103
rect 477 -161 533 -105
rect 592 -161 648 -105
rect 719 -160 775 -104
rect 849 -158 905 -102
rect 1004 -408 1058 -354
rect 1114 -408 1168 -354
rect 1338 -548 1395 -491
rect 1115 -672 1169 -618
rect 1338 -658 1395 -601
rect 1115 -782 1169 -728
rect -101 -1575 -45 -1519
rect -101 -1685 -45 -1629
rect 452 -1634 508 -1578
rect 587 -1633 643 -1577
rect 717 -1632 773 -1576
rect 860 -1633 916 -1577
rect -328 -2075 -272 -2019
rect -218 -2075 -162 -2019
rect -1080 -2527 -1024 -2471
rect -970 -2527 -914 -2471
rect -860 -2527 -804 -2471
rect -750 -2527 -694 -2471
rect -640 -2527 -584 -2471
rect -3040 -4053 -2984 -3997
rect -2919 -4053 -2863 -3997
rect -658 -4046 -602 -3990
rect -520 -4045 -464 -3989
rect -5030 -4265 -4974 -4209
rect -5030 -4375 -4974 -4319
rect -2595 -4256 -2539 -4200
rect -2595 -4366 -2539 -4310
rect -5225 -5575 -5168 -5518
rect -5225 -5685 -5168 -5628
rect -331 -4396 -271 -4336
rect -218 -4396 -158 -4336
rect -1189 -5106 -1133 -5050
rect -1079 -5106 -1023 -5050
rect -969 -5106 -913 -5050
rect -859 -5106 -803 -5050
rect -749 -5106 -693 -5050
rect -639 -5106 -583 -5050
rect 24 -2075 80 -2019
rect 24 -2185 80 -2129
rect 756 -2224 810 -2170
rect 866 -2224 920 -2170
rect 395 -3103 451 -3047
rect 513 -3101 569 -3045
rect 637 -3100 693 -3044
rect 746 -3100 802 -3044
rect 866 -3102 922 -3046
rect 765 -3975 819 -3921
rect 875 -3975 929 -3921
rect 19 -4277 73 -4223
rect 19 -4387 73 -4333
rect 1225 -916 1281 -860
rect 1225 -1026 1281 -970
rect 1226 -1964 1280 -1910
rect 1226 -2074 1280 -2020
rect 1115 -2219 1169 -2165
rect 1115 -2329 1169 -2275
rect 1115 -4139 1169 -4085
rect 1115 -4249 1169 -4195
rect 2330 -140 2384 -86
rect 2646 -145 2702 -89
rect 2966 -145 3022 -89
rect 3288 -144 3344 -88
rect 3735 -146 3791 -90
rect 4057 -147 4113 -91
rect 4378 -144 4434 -88
rect 4699 -153 4753 -99
rect 5394 -514 5448 -460
rect 5394 -624 5448 -570
rect 1635 -783 1689 -729
rect 1745 -783 1799 -729
rect 5269 -789 5325 -733
rect 5269 -899 5325 -843
rect 7078 -801 7132 -747
rect 7078 -911 7132 -857
rect 3512 -1119 3566 -1065
rect 3512 -1229 3566 -1175
rect 5498 -1157 5554 -1101
rect 7078 -1021 7132 -967
rect 5893 -1156 5947 -1102
rect 1492 -1447 1548 -1391
rect 1492 -1557 1548 -1501
rect 1492 -1667 1548 -1611
rect 6507 -2525 6561 -2473
rect 6627 -2525 6681 -2473
rect 6747 -2525 6801 -2473
rect 6867 -2525 6921 -2473
rect 6987 -2525 7041 -2473
rect 1702 -2917 1758 -2861
rect 1702 -3027 1758 -2971
rect 1702 -3137 1758 -3081
rect 1333 -3865 1390 -3808
rect 1333 -3975 1390 -3918
rect 3533 -3881 3591 -3823
rect 3533 -3991 3591 -3933
rect 5498 -3897 5554 -3841
rect 5889 -3896 5943 -3842
rect 7096 -4031 7150 -3977
rect 5253 -4155 5309 -4099
rect 7096 -4141 7150 -4087
rect 5253 -4265 5309 -4209
rect 7096 -4251 7150 -4197
rect 5419 -4397 5473 -4343
rect 1004 -4566 1058 -4512
rect 1114 -4566 1168 -4512
rect 5419 -4507 5473 -4453
rect 2337 -4891 2391 -4837
rect 2645 -4888 2701 -4832
rect 2966 -4901 3022 -4845
rect 3283 -4904 3339 -4848
rect 3745 -4904 3801 -4848
rect 4057 -4902 4113 -4846
rect 4377 -4899 4433 -4843
rect 4699 -4897 4753 -4843
rect 86 -5106 142 -5050
rect 196 -5106 252 -5050
rect 306 -5106 362 -5050
rect 416 -5106 472 -5050
rect 526 -5106 582 -5050
rect 636 -5106 692 -5050
rect 746 -5106 802 -5050
rect 7758 -802 7814 -746
rect 7868 -802 7924 -746
rect 7758 -912 7814 -856
rect 7868 -912 7924 -856
rect 7758 -1022 7814 -966
rect 7868 -1022 7924 -966
rect 7509 -2354 7565 -2298
rect 7619 -2354 7675 -2298
rect 7509 -2464 7565 -2408
rect 7619 -2464 7675 -2408
rect 7509 -2574 7565 -2518
rect 7619 -2574 7675 -2518
rect 1728 -5392 1783 -5337
rect 1728 -5502 1783 -5447
rect 3480 -5364 3534 -5310
rect 3480 -5474 3534 -5420
rect 5335 -5398 5391 -5342
rect -85 -5703 -28 -5646
rect -5019 -5834 -4963 -5778
rect -5019 -5944 -4963 -5888
rect -2601 -5838 -2545 -5782
rect -85 -5813 -28 -5756
rect -2601 -5948 -2545 -5892
rect -5119 -6106 -5062 -6049
rect 57 -6097 113 -6041
rect -5119 -6216 -5062 -6159
rect -3038 -6173 -2982 -6117
rect -2908 -6173 -2852 -6117
rect -633 -6166 -577 -6110
rect -508 -6166 -452 -6110
rect 448 -6096 504 -6040
rect 5335 -5508 5391 -5452
rect 3002 -6095 3056 -6041
rect 3631 -6096 3687 -6040
rect 4021 -6097 4077 -6041
rect 7108 -5810 7162 -5756
rect 7108 -5920 7162 -5866
rect 6682 -6096 6736 -6042
rect 7075 -6317 7131 -6261
rect 7753 -4032 7809 -3976
rect 7863 -4032 7919 -3976
rect 7753 -4142 7809 -4086
rect 7863 -4142 7919 -4086
rect 7753 -4252 7809 -4196
rect 7863 -4252 7919 -4196
rect 7509 -7514 7565 -7458
rect 7619 -7514 7675 -7458
rect 7509 -7624 7565 -7568
rect 7619 -7624 7675 -7568
rect 6507 -7685 6561 -7633
rect 6627 -7685 6681 -7633
rect 6747 -7685 6801 -7633
rect 6867 -7685 6921 -7633
rect 6987 -7685 7041 -7633
rect 7509 -7734 7565 -7678
rect 7619 -7734 7675 -7678
<< metal2 >>
rect 6445 2731 7676 2748
rect 6445 2687 7507 2731
rect 6445 2635 6507 2687
rect 6561 2635 6627 2687
rect 6681 2635 6747 2687
rect 6801 2635 6867 2687
rect 6921 2635 6987 2687
rect 7041 2675 7507 2687
rect 7563 2675 7617 2731
rect 7673 2675 7676 2731
rect 7041 2635 7676 2675
rect 6445 2621 7676 2635
rect 6445 2574 7507 2621
rect 7503 2565 7507 2574
rect 7563 2565 7617 2621
rect 7673 2565 7676 2621
rect 7503 2511 7676 2565
rect -3019 2367 7142 2480
rect 7503 2455 7507 2511
rect 7563 2455 7617 2511
rect 7673 2455 7676 2511
rect 7503 2443 7676 2455
rect -5214 1204 -5093 1208
rect -5214 1147 -5197 1204
rect -5140 1202 -5093 1204
rect -5140 1147 -4773 1202
rect -3019 1172 -2906 2367
rect -591 1933 3696 2047
rect -591 1180 -477 1933
rect -174 1655 3070 1684
rect -174 1599 -159 1655
rect -103 1653 3070 1655
rect -103 1599 -40 1653
rect -174 1597 -40 1599
rect 16 1597 67 1653
rect 123 1597 3070 1653
rect -174 1568 3070 1597
rect 2943 1319 3070 1568
rect 3385 1320 3462 1332
rect 3385 1319 3395 1320
rect 2943 1265 3002 1319
rect 3056 1265 3395 1319
rect 2943 1264 3395 1265
rect 3451 1264 3462 1320
rect -59 1221 129 1223
rect -59 1210 517 1221
rect -59 1206 57 1210
rect -591 1179 -449 1180
rect -5214 1094 -4773 1147
rect -3028 1161 -2840 1172
rect -3028 1105 -3020 1161
rect -2964 1105 -2909 1161
rect -2853 1105 -2840 1161
rect -3028 1097 -2840 1105
rect -3020 1095 -2964 1097
rect -5214 1037 -5197 1094
rect -5140 1037 -4773 1094
rect -5214 1026 -4773 1037
rect -5111 958 -4887 969
rect -2689 958 -2481 974
rect -5111 941 -2481 958
rect -5111 885 -5104 941
rect -5048 885 -4994 941
rect -4938 930 -2481 941
rect -4938 885 -2681 930
rect -5111 874 -2681 885
rect -2625 874 -2571 930
rect -2515 874 -2481 930
rect -5111 868 -2481 874
rect -5111 853 -4887 868
rect -2689 830 -2481 868
rect -5197 711 -5101 714
rect -5197 654 -5170 711
rect -5113 699 -5101 711
rect -2219 699 -2062 1177
rect -637 1170 -437 1179
rect -637 1169 -505 1170
rect -637 1113 -625 1169
rect -569 1114 -505 1169
rect -449 1114 -437 1170
rect -569 1113 -437 1114
rect -637 1104 -437 1113
rect -59 1150 -47 1206
rect 9 1154 57 1206
rect 113 1154 517 1210
rect 9 1150 517 1154
rect -625 1103 -569 1104
rect -59 1101 517 1150
rect 2943 1195 3462 1264
rect 2943 1142 3070 1195
rect 3385 1135 3462 1195
rect 3573 1320 3696 1933
rect 3573 1264 3631 1320
rect 3687 1264 3696 1320
rect 3573 1134 3696 1264
rect 6673 1328 6750 1339
rect 6673 1274 6685 1328
rect 6739 1306 6750 1328
rect 7018 1319 7142 2367
rect 7018 1306 7075 1319
rect 6739 1274 7075 1306
rect 6673 1263 7075 1274
rect 7131 1263 7142 1319
rect 6673 1201 7142 1263
rect 6673 1142 6750 1201
rect 7018 1126 7142 1201
rect -59 1045 -47 1101
rect 9 1100 517 1101
rect 9 1045 58 1100
rect -59 1044 58 1045
rect 114 1099 517 1100
rect 114 1053 453 1099
rect 114 1044 129 1053
rect -59 1028 129 1044
rect 438 1045 453 1053
rect 507 1045 517 1099
rect 438 1033 517 1045
rect 7144 915 7234 944
rect 7144 858 7161 915
rect 7218 858 7234 915
rect -102 805 -13 821
rect 7144 805 7234 858
rect -102 748 -84 805
rect -27 748 7161 805
rect 7218 748 7234 805
rect -102 732 -13 748
rect 7144 739 7234 748
rect 7505 774 7678 791
rect -5113 654 -2062 699
rect 7505 718 7509 774
rect 7565 718 7619 774
rect 7675 718 7678 774
rect 7505 682 7678 718
rect -5197 601 -2062 654
rect -5197 544 -5170 601
rect -5113 544 -2062 601
rect -5197 542 -2062 544
rect 824 664 7678 682
rect 824 608 7509 664
rect 7565 608 7619 664
rect 7675 608 7678 664
rect 824 554 7678 608
rect -5197 540 -5101 542
rect 824 540 7509 554
rect -1023 114 645 170
rect -1023 109 80 114
rect -1023 53 -1009 109
rect -953 53 -899 109
rect -843 53 -789 109
rect -733 53 -679 109
rect -623 58 80 109
rect 136 58 190 114
rect 246 58 300 114
rect 356 58 410 114
rect 466 58 520 114
rect 576 58 645 114
rect -623 53 645 58
rect -1023 -6 645 53
rect 824 -74 966 540
rect 7505 498 7509 540
rect 7565 498 7619 554
rect 7675 498 7678 554
rect 7505 486 7678 498
rect 3470 454 3543 466
rect 342 -102 966 -74
rect 342 -103 849 -102
rect 342 -159 352 -103
rect 408 -104 849 -103
rect 408 -105 719 -104
rect 408 -159 477 -105
rect 342 -161 477 -159
rect 533 -161 592 -105
rect 648 -160 719 -105
rect 775 -158 849 -104
rect 905 -158 966 -102
rect 1708 415 1788 430
rect 1708 360 1721 415
rect 1776 360 1788 415
rect 1708 305 1788 360
rect 1708 250 1721 305
rect 1776 250 1788 305
rect 3470 400 3480 454
rect 3534 400 3543 454
rect 3470 344 3543 400
rect 3470 290 3480 344
rect 3534 290 3543 344
rect 3470 277 3543 290
rect 5285 402 5365 415
rect 5285 346 5297 402
rect 5353 346 5365 402
rect 5285 292 5365 346
rect 1708 -71 1788 250
rect 1708 -86 3363 -71
rect 1708 -140 2330 -86
rect 2384 -88 3363 -86
rect 2384 -89 3288 -88
rect 2384 -140 2646 -89
rect 1708 -145 2646 -140
rect 2702 -145 2966 -89
rect 3022 -144 3288 -89
rect 3344 -144 3363 -88
rect 3022 -145 3363 -144
rect 1708 -154 3363 -145
rect 2646 -155 2702 -154
rect 2966 -155 3022 -154
rect 775 -160 966 -158
rect 648 -161 966 -160
rect 342 -174 966 -161
rect 991 -350 1178 -341
rect 3482 -350 3538 277
rect 5285 236 5297 292
rect 5353 236 5365 292
rect 3718 -86 3804 -80
rect 4041 -86 4127 -80
rect 4361 -86 4447 -75
rect 5285 -86 5365 236
rect 3718 -88 5365 -86
rect 3718 -90 4378 -88
rect 3718 -146 3735 -90
rect 3791 -91 4378 -90
rect 3791 -146 4057 -91
rect 3718 -147 4057 -146
rect 4113 -144 4378 -91
rect 4434 -99 5365 -88
rect 4434 -144 4699 -99
rect 4113 -147 4699 -144
rect 3718 -153 4699 -147
rect 4753 -153 5365 -99
rect 3718 -164 5365 -153
rect 991 -354 3538 -350
rect 991 -408 1004 -354
rect 1058 -408 1114 -354
rect 1168 -406 3538 -354
rect 1168 -408 1178 -406
rect 991 -420 1178 -408
rect 5384 -460 5457 -444
rect 1326 -491 1407 -481
rect 1326 -548 1338 -491
rect 1395 -548 1407 -491
rect 1326 -568 1407 -548
rect 5384 -514 5394 -460
rect 5448 -514 5457 -460
rect 5384 -568 5457 -514
rect 1326 -570 5457 -568
rect 1326 -601 5394 -570
rect -5041 -623 -4935 -615
rect -5041 -679 -5016 -623
rect -4960 -659 -4935 -623
rect -2601 -624 -2501 -611
rect -2601 -659 -2582 -624
rect -4960 -679 -2582 -659
rect -5041 -680 -2582 -679
rect -2526 -680 -2501 -624
rect -5041 -733 -2501 -680
rect -5041 -789 -5016 -733
rect -4960 -734 -2501 -733
rect -4960 -770 -2582 -734
rect -4960 -789 -4935 -770
rect -5041 -804 -4935 -789
rect -2601 -790 -2582 -770
rect -2526 -790 -2501 -734
rect -2601 -806 -2501 -790
rect 1106 -618 1178 -607
rect 1106 -672 1115 -618
rect 1169 -672 1178 -618
rect 1326 -658 1338 -601
rect 1395 -624 5394 -601
rect 5448 -624 5457 -570
rect 1395 -625 5457 -624
rect 1395 -658 1407 -625
rect 5384 -635 5457 -625
rect 1326 -670 1407 -658
rect 1106 -726 1178 -672
rect 1623 -726 1856 -718
rect 1106 -728 1856 -726
rect 1106 -782 1115 -728
rect 1169 -729 1856 -728
rect 1169 -782 1635 -729
rect 1106 -795 1178 -782
rect 1623 -783 1635 -782
rect 1689 -783 1745 -729
rect 1799 -783 1856 -729
rect 1623 -795 1856 -783
rect 5255 -733 5337 -720
rect 5255 -789 5269 -733
rect 5325 -789 5337 -733
rect 5255 -843 5337 -789
rect 1213 -858 1293 -848
rect 5255 -858 5269 -843
rect 1213 -860 5269 -858
rect -5194 -914 -4716 -878
rect -5194 -972 -5181 -914
rect -5123 -972 -4716 -914
rect 1213 -916 1225 -860
rect 1281 -899 5269 -860
rect 5325 -899 5337 -843
rect 1281 -914 5337 -899
rect 7066 -747 7145 -731
rect 7066 -801 7078 -747
rect 7132 -801 7145 -747
rect 7066 -808 7145 -801
rect 7747 -746 7936 -730
rect 7747 -802 7758 -746
rect 7814 -802 7868 -746
rect 7924 -802 7936 -746
rect 7747 -808 7936 -802
rect 7066 -856 7936 -808
rect 7066 -857 7758 -856
rect 7066 -911 7078 -857
rect 7132 -911 7758 -857
rect 7066 -912 7758 -911
rect 7814 -912 7868 -856
rect 7924 -912 7936 -856
rect 1281 -916 1293 -914
rect -5194 -1024 -4716 -972
rect -5194 -1082 -5181 -1024
rect -5123 -1054 -4716 -1024
rect -3049 -958 -2839 -948
rect -3049 -1014 -3039 -958
rect -2983 -959 -2839 -958
rect -2983 -1014 -2921 -959
rect -3049 -1015 -2921 -1014
rect -2865 -1015 -2839 -959
rect -3049 -1025 -2839 -1015
rect -5123 -1082 -5099 -1054
rect -5194 -1094 -5099 -1082
rect -5189 -1386 -5094 -1381
rect -2279 -1386 -2122 -932
rect -621 -942 -565 -940
rect -502 -942 -446 -940
rect -630 -950 -436 -942
rect -630 -1006 -621 -950
rect -565 -1006 -502 -950
rect -446 -1006 -436 -950
rect -630 -1017 -436 -1006
rect 1213 -970 1293 -916
rect 7066 -966 7936 -912
rect 7066 -967 7758 -966
rect 1213 -1026 1225 -970
rect 1281 -1026 1293 -970
rect 5442 -980 5564 -970
rect 1213 -1033 1293 -1026
rect 3492 -1065 3604 -1016
rect 3492 -1119 3512 -1065
rect 3566 -1119 3604 -1065
rect 3492 -1142 3604 -1119
rect 5442 -1101 5956 -980
rect 7066 -1021 7078 -967
rect 7132 -1021 7758 -967
rect 7066 -1022 7758 -1021
rect 7814 -1022 7868 -966
rect 7924 -1022 7936 -966
rect 7066 -1034 7146 -1022
rect 7747 -1034 7936 -1022
rect 5442 -1142 5498 -1101
rect 3492 -1157 5498 -1142
rect 5554 -1102 5956 -1101
rect 5554 -1156 5893 -1102
rect 5947 -1156 5956 -1102
rect 5554 -1157 5956 -1156
rect 3492 -1174 5956 -1157
rect 3492 -1175 5564 -1174
rect 5878 -1175 5956 -1174
rect 3492 -1229 3512 -1175
rect 3566 -1229 5564 -1175
rect 3492 -1254 5564 -1229
rect -5189 -1391 -2122 -1386
rect -5189 -1447 -5164 -1391
rect -5108 -1447 -2122 -1391
rect -5189 -1501 -2122 -1447
rect -5189 -1557 -5164 -1501
rect -5108 -1543 -2122 -1501
rect 1458 -1391 1584 -1389
rect 1458 -1447 1492 -1391
rect 1548 -1447 1584 -1391
rect 1458 -1501 1584 -1447
rect -126 -1519 -31 -1509
rect -5108 -1557 -5094 -1543
rect -5189 -1567 -5094 -1557
rect -126 -1575 -101 -1519
rect -45 -1575 -31 -1519
rect 1458 -1557 1492 -1501
rect 1548 -1557 1584 -1501
rect 1458 -1559 1584 -1557
rect -126 -1629 -31 -1575
rect -126 -1635 -101 -1629
rect -5286 -1685 -101 -1635
rect -45 -1685 -31 -1629
rect 441 -1576 1584 -1559
rect 441 -1577 717 -1576
rect 441 -1578 587 -1577
rect 441 -1634 452 -1578
rect 508 -1633 587 -1578
rect 643 -1632 717 -1577
rect 773 -1577 1584 -1576
rect 773 -1632 860 -1577
rect 643 -1633 860 -1632
rect 916 -1611 1584 -1577
rect 916 -1633 1492 -1611
rect 508 -1634 1492 -1633
rect 441 -1667 1492 -1634
rect 1548 -1667 1584 -1611
rect 441 -1674 1584 -1667
rect -5286 -1691 -31 -1685
rect -126 -1695 -31 -1691
rect 1216 -1910 1287 -1898
rect 1216 -1964 1226 -1910
rect 1280 -1964 1287 -1910
rect -340 -2019 -150 -2011
rect 7 -2019 92 -2007
rect 1216 -2019 1287 -1964
rect -5292 -2075 -328 -2019
rect -272 -2075 -218 -2019
rect -162 -2075 24 -2019
rect 80 -2020 1287 -2019
rect 80 -2074 1226 -2020
rect 1280 -2074 1287 -2020
rect 80 -2075 1287 -2074
rect -340 -2082 -150 -2075
rect 7 -2129 92 -2075
rect 1216 -2087 1287 -2075
rect 7 -2185 24 -2129
rect 80 -2185 92 -2129
rect 7 -2195 92 -2185
rect 746 -2166 935 -2155
rect 1104 -2165 1180 -2153
rect 1104 -2166 1115 -2165
rect 746 -2170 1115 -2166
rect 746 -2224 756 -2170
rect 810 -2224 866 -2170
rect 920 -2219 1115 -2170
rect 1169 -2219 1180 -2165
rect 920 -2222 1180 -2219
rect 920 -2224 935 -2222
rect 746 -2238 935 -2224
rect 1104 -2275 1180 -2222
rect 1104 -2329 1115 -2275
rect 1169 -2329 1180 -2275
rect 1104 -2340 1180 -2329
rect 7505 -2298 7678 -2281
rect 7505 -2354 7509 -2298
rect 7565 -2354 7619 -2298
rect 7675 -2354 7678 -2298
rect 7505 -2408 7678 -2354
rect 7505 -2412 7509 -2408
rect -1090 -2428 -518 -2412
rect -1090 -2471 -258 -2428
rect -1090 -2527 -1080 -2471
rect -1024 -2527 -970 -2471
rect -914 -2527 -860 -2471
rect -804 -2527 -750 -2471
rect -694 -2527 -640 -2471
rect -584 -2527 -258 -2471
rect -1090 -2552 -258 -2527
rect -1090 -2585 -518 -2552
rect -382 -3020 -258 -2552
rect 6445 -2464 7509 -2412
rect 7565 -2464 7619 -2408
rect 7675 -2464 7678 -2408
rect 6445 -2473 7678 -2464
rect 6445 -2525 6507 -2473
rect 6561 -2525 6627 -2473
rect 6681 -2525 6747 -2473
rect 6801 -2525 6867 -2473
rect 6921 -2525 6987 -2473
rect 7041 -2518 7678 -2473
rect 7041 -2525 7509 -2518
rect 6445 -2574 7509 -2525
rect 7565 -2574 7619 -2518
rect 7675 -2574 7678 -2518
rect 6445 -2586 7678 -2574
rect 1666 -2861 1794 -2850
rect 1666 -2917 1702 -2861
rect 1758 -2917 1794 -2861
rect 1666 -2971 1794 -2917
rect 373 -3020 922 -3019
rect 1666 -3020 1702 -2971
rect -382 -3027 1702 -3020
rect 1758 -3027 1794 -2971
rect -382 -3044 1794 -3027
rect -382 -3045 637 -3044
rect -382 -3047 513 -3045
rect -382 -3103 395 -3047
rect 451 -3101 513 -3047
rect 569 -3100 637 -3045
rect 693 -3100 746 -3044
rect 802 -3046 1794 -3044
rect 802 -3100 866 -3046
rect 569 -3101 866 -3100
rect 451 -3102 866 -3101
rect 922 -3081 1794 -3046
rect 922 -3102 1702 -3081
rect 451 -3103 1702 -3102
rect -382 -3137 1702 -3103
rect 1758 -3137 1794 -3081
rect -382 -3143 1794 -3137
rect -382 -3144 1702 -3143
rect -5193 -3268 -5137 -3265
rect -5209 -3275 -5121 -3268
rect -5209 -3331 -5193 -3275
rect -5137 -3293 -5121 -3275
rect -5137 -3331 -2150 -3293
rect -5209 -3385 -2150 -3331
rect -5209 -3441 -5193 -3385
rect -5137 -3407 -2150 -3385
rect -5137 -3441 -5121 -3407
rect -5209 -3458 -5121 -3441
rect -5189 -3958 -5107 -3947
rect -5189 -3960 -4706 -3958
rect -5189 -4018 -5177 -3960
rect -5119 -4018 -4706 -3960
rect -3040 -3988 -2984 -3987
rect -2919 -3988 -2863 -3987
rect -5189 -4070 -4706 -4018
rect -3050 -3997 -2840 -3988
rect -3050 -4053 -3040 -3997
rect -2984 -4053 -2919 -3997
rect -2863 -4053 -2840 -3997
rect -3050 -4063 -2840 -4053
rect -5189 -4128 -5177 -4070
rect -5119 -4128 -4706 -4070
rect -2264 -4093 -2150 -3407
rect 1323 -3808 1405 -3796
rect 1323 -3865 1333 -3808
rect 1390 -3865 1405 -3808
rect 749 -3918 941 -3906
rect 1323 -3918 1405 -3865
rect 749 -3921 1333 -3918
rect 749 -3975 765 -3921
rect 819 -3975 875 -3921
rect 929 -3975 1333 -3921
rect 1390 -3975 1405 -3918
rect -658 -3981 -602 -3980
rect -520 -3981 -464 -3979
rect -673 -3989 -437 -3981
rect 749 -3987 941 -3975
rect 1323 -3989 1405 -3975
rect 3520 -3823 5564 -3765
rect 3520 -3881 3533 -3823
rect 3591 -3838 5564 -3823
rect 5876 -3838 5956 -3836
rect 3591 -3841 5956 -3838
rect 3591 -3881 5498 -3841
rect 3520 -3933 3602 -3881
rect -673 -3990 -520 -3989
rect -673 -4046 -658 -3990
rect -602 -4045 -520 -3990
rect -464 -4045 -437 -3989
rect 3520 -3991 3533 -3933
rect 3591 -3991 3602 -3933
rect 3520 -4017 3602 -3991
rect 5487 -3897 5498 -3881
rect 5554 -3842 5956 -3841
rect 5554 -3896 5889 -3842
rect 5943 -3896 5956 -3842
rect 5554 -3897 5956 -3896
rect 5487 -3957 5956 -3897
rect 5487 -4027 5564 -3957
rect 5876 -4018 5956 -3957
rect 7084 -3976 7162 -3964
rect 7744 -3976 7933 -3963
rect 7084 -3977 7753 -3976
rect -602 -4046 -437 -4045
rect -673 -4057 -437 -4046
rect 7084 -4031 7096 -3977
rect 7150 -4031 7753 -3977
rect 7084 -4032 7753 -4031
rect 7809 -4032 7863 -3976
rect 7919 -4032 7933 -3976
rect 1103 -4084 1180 -4072
rect 5244 -4084 5322 -4083
rect 1103 -4085 5322 -4084
rect -5189 -4134 -4706 -4128
rect -5189 -4135 -5107 -4134
rect 1103 -4139 1115 -4085
rect 1169 -4099 5322 -4085
rect 1169 -4139 5253 -4099
rect 1103 -4140 5253 -4139
rect -5055 -4209 -4960 -4199
rect -5055 -4265 -5030 -4209
rect -4974 -4224 -4960 -4209
rect -2620 -4200 -2525 -4190
rect -2620 -4224 -2595 -4200
rect -4974 -4256 -2595 -4224
rect -2539 -4256 -2525 -4200
rect 1103 -4195 1180 -4140
rect -4974 -4265 -2525 -4256
rect -5055 -4310 -2525 -4265
rect -5055 -4319 -2595 -4310
rect -5055 -4375 -5030 -4319
rect -4974 -4344 -2595 -4319
rect -4974 -4375 -4960 -4344
rect -5055 -4385 -4960 -4375
rect -2620 -4366 -2595 -4344
rect -2539 -4366 -2525 -4310
rect 7 -4223 86 -4207
rect 7 -4277 19 -4223
rect 73 -4277 86 -4223
rect 1103 -4249 1115 -4195
rect 1169 -4249 1180 -4195
rect 1103 -4263 1180 -4249
rect 5244 -4155 5253 -4140
rect 5309 -4155 5322 -4099
rect 5244 -4202 5322 -4155
rect 7084 -4086 7933 -4032
rect 7084 -4087 7753 -4086
rect 7084 -4141 7096 -4087
rect 7150 -4141 7753 -4087
rect 7084 -4142 7753 -4141
rect 7809 -4142 7863 -4086
rect 7919 -4142 7933 -4086
rect 7084 -4175 7933 -4142
rect 7084 -4197 7162 -4175
rect 5244 -4209 5324 -4202
rect 5244 -4265 5253 -4209
rect 5309 -4265 5324 -4209
rect 5244 -4276 5324 -4265
rect 7084 -4251 7096 -4197
rect 7150 -4251 7162 -4197
rect 7084 -4268 7162 -4251
rect 7744 -4196 7933 -4175
rect 7744 -4252 7753 -4196
rect 7809 -4252 7863 -4196
rect 7919 -4252 7933 -4196
rect 7744 -4267 7933 -4252
rect -2620 -4376 -2525 -4366
rect -340 -4336 -151 -4324
rect 7 -4333 86 -4277
rect 7 -4336 19 -4333
rect -340 -4396 -331 -4336
rect -271 -4396 -218 -4336
rect -158 -4387 19 -4336
rect 73 -4336 86 -4333
rect 5412 -4336 5484 -4329
rect 73 -4343 5484 -4336
rect 73 -4387 5419 -4343
rect -158 -4396 5419 -4387
rect -340 -4408 -79 -4396
rect 7 -4399 86 -4396
rect 5412 -4397 5419 -4396
rect 5473 -4397 5484 -4343
rect -139 -4513 -79 -4408
rect 5412 -4453 5484 -4397
rect -5306 -4573 -79 -4513
rect 991 -4512 1180 -4500
rect 991 -4566 1004 -4512
rect 1058 -4566 1114 -4512
rect 1168 -4514 1180 -4512
rect 5412 -4507 5419 -4453
rect 5473 -4507 5484 -4453
rect 1168 -4566 3535 -4514
rect 5412 -4522 5484 -4507
rect 991 -4570 3535 -4566
rect 991 -4579 1180 -4570
rect 2625 -4832 2717 -4822
rect 1715 -4837 2403 -4833
rect 2625 -4837 2645 -4832
rect 1715 -4891 2337 -4837
rect 2391 -4888 2645 -4837
rect 2701 -4837 2717 -4832
rect 2952 -4837 3037 -4835
rect 2701 -4845 3349 -4837
rect 2701 -4888 2966 -4845
rect 2391 -4891 2966 -4888
rect 1715 -4901 2966 -4891
rect 3022 -4848 3349 -4845
rect 3022 -4901 3283 -4848
rect 1715 -4904 3283 -4901
rect 3339 -4904 3349 -4848
rect 1715 -4906 3349 -4904
rect -1209 -5050 867 -4988
rect -1209 -5106 -1189 -5050
rect -1133 -5106 -1079 -5050
rect -1023 -5106 -969 -5050
rect -913 -5106 -859 -5050
rect -803 -5106 -749 -5050
rect -693 -5106 -639 -5050
rect -583 -5106 86 -5050
rect 142 -5106 196 -5050
rect 252 -5106 306 -5050
rect 362 -5106 416 -5050
rect 472 -5106 526 -5050
rect 582 -5106 636 -5050
rect 692 -5106 746 -5050
rect 802 -5106 867 -5050
rect -1209 -5165 867 -5106
rect 1715 -5337 1795 -4906
rect 2371 -4916 3349 -4906
rect 2371 -4917 3325 -4916
rect 3479 -5297 3535 -4570
rect 4708 -4828 5408 -4827
rect 3732 -4842 3813 -4834
rect 4044 -4842 4125 -4828
rect 4364 -4842 4445 -4830
rect 4683 -4842 5408 -4828
rect 3732 -4843 5408 -4842
rect 3732 -4846 4377 -4843
rect 3732 -4848 4057 -4846
rect 3732 -4904 3745 -4848
rect 3801 -4898 4057 -4848
rect 3801 -4904 3813 -4898
rect 3732 -4920 3813 -4904
rect 4044 -4902 4057 -4898
rect 4113 -4898 4377 -4846
rect 4113 -4902 4125 -4898
rect 4044 -4914 4125 -4902
rect 4364 -4899 4377 -4898
rect 4433 -4897 4699 -4843
rect 4753 -4897 5408 -4843
rect 4433 -4898 5408 -4897
rect 4433 -4899 4445 -4898
rect 4364 -4916 4445 -4899
rect 4683 -4909 5408 -4898
rect 4708 -4929 5408 -4909
rect 1715 -5392 1728 -5337
rect 1783 -5392 1795 -5337
rect 1715 -5447 1795 -5392
rect 1715 -5502 1728 -5447
rect 1783 -5502 1795 -5447
rect 3470 -5310 3543 -5297
rect 3470 -5364 3480 -5310
rect 3534 -5364 3543 -5310
rect 3470 -5420 3543 -5364
rect 3470 -5474 3480 -5420
rect 3534 -5474 3543 -5420
rect 3470 -5493 3543 -5474
rect 5321 -5342 5408 -4929
rect 5321 -5398 5335 -5342
rect 5391 -5398 5408 -5342
rect 5321 -5452 5408 -5398
rect 1715 -5504 1795 -5502
rect -5235 -5518 -5162 -5506
rect 5321 -5508 5335 -5452
rect 5391 -5508 5408 -5452
rect 5321 -5515 5408 -5508
rect -5235 -5575 -5225 -5518
rect -5168 -5575 -2149 -5518
rect -5235 -5628 -2149 -5575
rect -5235 -5685 -5225 -5628
rect -5168 -5632 -2149 -5628
rect -5168 -5685 -5162 -5632
rect -5235 -5697 -5162 -5685
rect -5044 -5778 -4949 -5768
rect -5044 -5834 -5019 -5778
rect -4963 -5824 -4949 -5778
rect -2626 -5782 -2531 -5772
rect -2626 -5824 -2601 -5782
rect -4963 -5834 -2601 -5824
rect -5044 -5838 -2601 -5834
rect -2545 -5838 -2531 -5782
rect -5044 -5888 -2531 -5838
rect -5044 -5944 -5019 -5888
rect -4963 -5892 -2531 -5888
rect -4963 -5944 -2601 -5892
rect -5044 -5954 -4949 -5944
rect -2626 -5948 -2601 -5944
rect -2545 -5948 -2531 -5892
rect -2626 -5958 -2531 -5948
rect -5128 -6049 -4798 -6038
rect -5128 -6106 -5119 -6049
rect -5062 -6106 -4798 -6049
rect -5128 -6159 -4798 -6106
rect -3038 -6109 -2982 -6107
rect -2908 -6109 -2852 -6107
rect -5128 -6216 -5119 -6159
rect -5062 -6214 -4798 -6159
rect -3046 -6117 -2840 -6109
rect -3046 -6173 -3038 -6117
rect -2982 -6173 -2908 -6117
rect -2852 -6173 -2840 -6117
rect -2263 -6160 -2149 -5632
rect -97 -5646 -16 -5642
rect -97 -5703 -85 -5646
rect -28 -5703 -16 -5646
rect -97 -5704 -16 -5703
rect -97 -5756 7176 -5704
rect -97 -5813 -85 -5756
rect -28 -5810 7108 -5756
rect 7162 -5810 7176 -5756
rect -28 -5813 7176 -5810
rect -97 -5823 -16 -5813
rect 7085 -5866 7176 -5813
rect 7085 -5920 7108 -5866
rect 7162 -5920 7176 -5866
rect 7085 -5944 7176 -5920
rect -80 -6041 124 -6026
rect -80 -6047 57 -6041
rect -633 -6102 -577 -6100
rect -508 -6102 -452 -6100
rect -641 -6110 -437 -6102
rect -3046 -6184 -2840 -6173
rect -641 -6166 -633 -6110
rect -577 -6166 -508 -6110
rect -452 -6166 -437 -6110
rect -641 -6177 -437 -6166
rect -80 -6103 -61 -6047
rect -5 -6097 57 -6047
rect 113 -6071 124 -6041
rect 439 -6040 516 -6028
rect 439 -6071 448 -6040
rect 113 -6096 448 -6071
rect 504 -6096 516 -6040
rect 113 -6097 516 -6096
rect -5 -6103 516 -6097
rect -80 -6150 516 -6103
rect -80 -6157 58 -6150
rect -5062 -6216 -5035 -6214
rect -5128 -6228 -5051 -6216
rect -2981 -7364 -2867 -6184
rect -574 -6986 -460 -6177
rect -80 -6213 -61 -6157
rect -5 -6206 58 -6157
rect 114 -6206 124 -6150
rect 439 -6154 516 -6150
rect 2943 -6041 3070 -6034
rect 2943 -6095 3002 -6041
rect 3056 -6095 3070 -6041
rect 2943 -6150 3070 -6095
rect 3573 -6040 3697 -6028
rect 4021 -6033 4077 -6031
rect 3573 -6096 3631 -6040
rect 3687 -6073 3697 -6040
rect 4012 -6041 4089 -6033
rect 4012 -6073 4021 -6041
rect 3687 -6096 4021 -6073
rect 3573 -6097 4021 -6096
rect 4077 -6097 4089 -6041
rect 3385 -6150 3462 -6131
rect -5 -6213 124 -6206
rect -80 -6220 124 -6213
rect 2943 -6206 3395 -6150
rect 3451 -6206 3462 -6150
rect 2943 -6217 3070 -6206
rect 2943 -6564 3059 -6217
rect 3385 -6219 3462 -6206
rect 3573 -6206 4089 -6097
rect 3573 -6219 3697 -6206
rect 4012 -6217 4089 -6206
rect 6673 -6042 6750 -6030
rect 6673 -6096 6682 -6042
rect 6736 -6096 6750 -6042
rect 6673 -6151 6750 -6096
rect 7066 -6132 7143 -6130
rect 7017 -6151 7143 -6132
rect 6673 -6152 7143 -6151
rect 6673 -6206 6682 -6152
rect 6736 -6206 7143 -6152
rect 6673 -6207 7143 -6206
rect 6673 -6218 6750 -6207
rect -315 -6592 3059 -6564
rect -315 -6648 -300 -6592
rect -244 -6593 3059 -6592
rect -244 -6594 -84 -6593
rect -244 -6648 -189 -6594
rect -315 -6650 -189 -6648
rect -133 -6649 -84 -6594
rect -28 -6649 3059 -6593
rect -133 -6650 3059 -6649
rect -315 -6680 3059 -6650
rect 3573 -6986 3687 -6219
rect -574 -7100 3687 -6986
rect 7017 -6261 7143 -6207
rect 7017 -6317 7075 -6261
rect 7131 -6317 7143 -6261
rect 7017 -6334 7143 -6317
rect 7017 -7364 7142 -6334
rect -2981 -7478 7142 -7364
rect 7505 -7458 7678 -7441
rect 7505 -7514 7509 -7458
rect 7565 -7514 7619 -7458
rect 7675 -7514 7678 -7458
rect 7505 -7568 7678 -7514
rect 7505 -7572 7509 -7568
rect 6445 -7624 7509 -7572
rect 7565 -7624 7619 -7568
rect 7675 -7624 7678 -7568
rect 6445 -7633 7678 -7624
rect 6445 -7685 6507 -7633
rect 6561 -7685 6627 -7633
rect 6681 -7685 6747 -7633
rect 6801 -7685 6867 -7633
rect 6921 -7685 6987 -7633
rect 7041 -7678 7678 -7633
rect 7041 -7685 7509 -7678
rect 6445 -7734 7509 -7685
rect 7565 -7734 7619 -7678
rect 7675 -7734 7678 -7678
rect 6445 -7746 7678 -7734
<< via2 >>
rect -159 1599 -103 1655
rect -40 1597 16 1653
rect 67 1597 123 1653
rect -47 1150 9 1206
rect 57 1154 113 1210
rect -47 1045 9 1101
rect 58 1044 114 1100
rect -3039 -1014 -2983 -958
rect -2921 -1015 -2865 -959
rect -621 -1006 -565 -950
rect -502 -1006 -446 -950
rect -3040 -4053 -2984 -3997
rect -2919 -4053 -2863 -3997
rect -658 -4046 -602 -3990
rect -520 -4045 -464 -3989
rect -61 -6103 -5 -6047
rect 57 -6097 113 -6041
rect -61 -6213 -5 -6157
rect 58 -6206 114 -6150
rect -300 -6648 -244 -6592
rect -189 -6650 -133 -6594
rect -84 -6649 -28 -6593
<< metal3 >>
rect -2973 1655 138 1684
rect -2973 1599 -159 1655
rect -103 1653 138 1655
rect -103 1599 -40 1653
rect -2973 1597 -40 1599
rect 16 1597 67 1653
rect 123 1597 138 1653
rect -2973 1568 138 1597
rect -2973 -948 -2857 1568
rect -59 1210 129 1223
rect -59 1207 57 1210
rect -609 1206 57 1207
rect -609 1150 -47 1206
rect 9 1154 57 1206
rect 113 1154 129 1210
rect 9 1150 129 1154
rect -609 1101 129 1150
rect -609 1063 -47 1101
rect -609 -942 -465 1063
rect -59 1045 -47 1063
rect 9 1100 129 1101
rect 9 1045 58 1100
rect -59 1044 58 1045
rect 114 1044 129 1100
rect -59 1028 129 1044
rect -3049 -958 -2839 -948
rect -630 -950 -436 -942
rect -3049 -1014 -3039 -958
rect -2983 -959 -2839 -958
rect -2983 -1014 -2921 -959
rect -3049 -1015 -2921 -1014
rect -2865 -1015 -2839 -959
rect -631 -1006 -621 -950
rect -565 -1006 -502 -950
rect -446 -1006 -436 -950
rect -3049 -1025 -2839 -1015
rect -630 -1017 -436 -1006
rect -3050 -3997 -2840 -3988
rect -3050 -4053 -3040 -3997
rect -2984 -4053 -2919 -3997
rect -2863 -4053 -2840 -3997
rect -3050 -4063 -2840 -4053
rect -673 -3989 -437 -3981
rect -673 -3990 -520 -3989
rect -673 -4046 -658 -3990
rect -602 -4045 -520 -3990
rect -464 -4045 -437 -3989
rect -602 -4046 -437 -4045
rect -673 -4057 -437 -4046
rect -2998 -6564 -2882 -4063
rect -612 -6038 -454 -4057
rect -80 -6038 124 -6026
rect -612 -6041 124 -6038
rect -612 -6047 57 -6041
rect -612 -6103 -61 -6047
rect -5 -6097 57 -6047
rect 113 -6097 124 -6041
rect -5 -6103 124 -6097
rect -612 -6150 124 -6103
rect -612 -6157 58 -6150
rect -612 -6196 -61 -6157
rect -80 -6213 -61 -6196
rect -5 -6206 58 -6157
rect 114 -6206 124 -6150
rect -5 -6213 124 -6206
rect -80 -6220 124 -6213
rect -2998 -6592 -15 -6564
rect -2998 -6648 -300 -6592
rect -244 -6593 -15 -6592
rect -244 -6594 -84 -6593
rect -244 -6648 -189 -6594
rect -2998 -6650 -189 -6648
rect -133 -6649 -84 -6594
rect -28 -6649 -15 -6593
rect -133 -6650 -15 -6649
rect -2998 -6680 -15 -6650
use INVERTER_MUX  INVERTER_MUX_0
timestamp 1691428809
transform 1 0 61 0 1 -996
box -1 -674 885 935
use INVERTER_MUX  INVERTER_MUX_1
timestamp 1691428809
transform 1 0 61 0 1 -3937
box -1 -674 885 935
use INVERTER_MUX  INVERTER_MUX_2
timestamp 1691428809
transform 1 0 61 0 -1 -2211
box -1 -674 885 935
use TG_GATE_SWITCH_magic  TG_GATE_SWITCH_magic_0
timestamp 1698649173
transform 1 0 -4564 0 -1 -720
box -439 -881 1724 1873
use TG_GATE_SWITCH_magic  TG_GATE_SWITCH_magic_1
timestamp 1698649173
transform 1 0 -4564 0 1 -4292
box -439 -881 1724 1873
use TG_GATE_SWITCH_magic  TG_GATE_SWITCH_magic_2
timestamp 1698649173
transform 1 0 -4564 0 -1 -5880
box -439 -881 1724 1873
use TG_GATE_SWITCH_magic  TG_GATE_SWITCH_magic_3
timestamp 1698649173
transform 1 0 -4564 0 1 868
box -439 -881 1724 1873
use TG_GATE_SWITCH_magic  TG_GATE_SWITCH_magic_4
timestamp 1698649173
transform 1 0 -2161 0 -1 -5873
box -439 -881 1724 1873
use TG_GATE_SWITCH_magic  TG_GATE_SWITCH_magic_5
timestamp 1698649173
transform 1 0 -2161 0 1 -4285
box -439 -881 1724 1873
use TG_GATE_SWITCH_magic  TG_GATE_SWITCH_magic_6
timestamp 1698649173
transform 1 0 -2161 0 -1 -713
box -439 -881 1724 1873
use TG_GATE_SWITCH_magic  TG_GATE_SWITCH_magic_7
timestamp 1698649173
transform 1 0 -2161 0 1 875
box -439 -881 1724 1873
use TG_magic  TG_magic_0
timestamp 1695364382
transform 1 0 1794 0 -1 -712
box -43 -881 1724 1873
use TG_magic  TG_magic_1
timestamp 1695364382
transform -1 0 3475 0 -1 -5872
box -43 -881 1724 1873
use TG_magic  TG_magic_2
timestamp 1695364382
transform 1 0 3607 0 -1 -5872
box -43 -881 1724 1873
use TG_magic  TG_magic_3
timestamp 1695364382
transform -1 0 7155 0 1 875
box -43 -881 1724 1873
use TG_magic  TG_magic_4
timestamp 1695364382
transform 1 0 34 0 -1 -5872
box -43 -881 1724 1873
use TG_magic  TG_magic_5
timestamp 1695364382
transform -1 0 5288 0 -1 -712
box -43 -881 1724 1873
use TG_magic  TG_magic_6
timestamp 1695364382
transform -1 0 3475 0 1 876
box -43 -881 1724 1873
use TG_magic  TG_magic_7
timestamp 1695364382
transform -1 0 5288 0 1 -4284
box -43 -881 1724 1873
use TG_magic  TG_magic_8
timestamp 1695364382
transform 1 0 5474 0 -1 -713
box -43 -881 1724 1873
use TG_magic  TG_magic_9
timestamp 1695364382
transform 1 0 1794 0 1 -4284
box -43 -881 1724 1873
use TG_magic  TG_magic_10
timestamp 1695364382
transform 1 0 34 0 1 876
box -43 -881 1724 1873
use TG_magic  TG_magic_11
timestamp 1695364382
transform 1 0 3607 0 1 876
box -43 -881 1724 1873
use TG_magic  TG_magic_12
timestamp 1695364382
transform 1 0 5474 0 1 -4285
box -43 -881 1724 1873
use TG_magic  TG_magic_13
timestamp 1695364382
transform -1 0 7155 0 -1 -5873
box -43 -881 1724 1873
<< labels >>
flabel metal1 -249 -4375 -249 -4375 0 FreeSans 800 0 0 0 S2
port 33 nsew
flabel via1 -286 -2051 -286 -2051 0 FreeSans 800 0 0 0 S1
port 34 nsew
flabel metal1 -62 -890 -62 -890 0 FreeSans 800 0 0 0 S0
port 3 nsew
flabel metal1 7779 -1906 7779 -1906 0 FreeSans 1120 0 0 0 Vout
port 36 nsew
flabel metal1 5373 2647 5373 2647 0 FreeSans 1600 0 0 0 VDD
port 38 nsew
flabel metal1 7170 -5116 7170 -5116 0 FreeSans 1600 0 0 0 VSS
port 40 nsew
flabel metal1 -5348 -6192 -5348 -6192 0 FreeSans 480 0 0 0 A5
port 29 nsew
flabel metal1 -5362 -5551 -5362 -5551 0 FreeSans 480 0 0 0 A1
port 30 nsew
flabel metal1 -5266 -3998 -5266 -3998 0 FreeSans 480 0 0 0 A3
port 43 nsew
flabel metal1 -5266 1147 -5266 1147 0 FreeSans 480 0 0 0 A6
port 27 nsew
flabel metal1 -5320 626 -5320 626 0 FreeSans 480 0 0 0 A2
port 26 nsew
flabel metal1 -5235 -1468 -5235 -1468 0 FreeSans 480 0 0 0 A4
port 28 nsew
flabel metal1 -5242 -3352 -5242 -3352 0 FreeSans 480 0 0 0 A7
port 45 nsew
flabel metal1 -5245 -994 -5245 -994 0 FreeSans 480 0 0 0 A0
port 6 nsew
flabel metal1 -5011 -24 -5010 -23 0 FreeSans 1600 0 0 0 ENA
port 47 nsew
<< end >>
