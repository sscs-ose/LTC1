magic
tech gf180mcuC
magscale 1 10
timestamp 1691496070
<< nwell >>
rect 540 4324 575 4336
<< metal1 >>
rect -590 8663 -510 8677
rect -590 8662 96 8663
rect -590 8608 -576 8662
rect -522 8608 96 8662
rect -590 8607 96 8608
rect -590 8598 -510 8607
rect 608 8296 694 8306
rect 608 8292 624 8296
rect 593 8246 624 8292
rect 608 8242 624 8246
rect 678 8242 694 8296
rect 76 8110 122 8241
rect 608 8231 694 8242
rect -409 7870 -330 7883
rect -409 7814 -397 7870
rect -341 7814 80 7870
rect -409 7808 -330 7814
rect -591 7687 -511 7699
rect -591 7631 -577 7687
rect -521 7631 98 7687
rect -591 7620 -511 7631
rect 600 7311 680 7323
rect 600 7307 613 7311
rect 49 7263 127 7267
rect 49 7207 61 7263
rect 117 7207 127 7263
rect 593 7261 613 7307
rect 600 7257 613 7261
rect 667 7257 680 7311
rect 600 7252 680 7257
rect 49 7196 127 7207
rect 76 7171 127 7196
rect 76 7125 122 7171
rect -407 6898 -328 6909
rect -407 6842 -397 6898
rect -341 6842 72 6898
rect -407 6834 -328 6842
rect -592 6716 -512 6728
rect -592 6660 -577 6716
rect -521 6660 98 6716
rect -592 6649 -512 6660
rect 873 6335 953 6347
rect 873 6331 886 6335
rect 43 6312 127 6320
rect 43 6256 55 6312
rect 111 6256 127 6312
rect 586 6285 886 6331
rect 873 6281 886 6285
rect 940 6281 953 6335
rect 873 6277 953 6281
rect 43 6243 127 6256
rect 352 6216 440 6228
rect 352 6160 365 6216
rect 421 6160 440 6216
rect 352 6152 440 6160
rect 364 6151 422 6152
rect -408 5911 -329 5920
rect -408 5855 -397 5911
rect -341 5855 70 5911
rect -408 5845 -329 5855
rect -589 5740 -509 5752
rect -589 5684 -577 5740
rect -521 5684 94 5740
rect -589 5673 -509 5684
rect 692 5360 780 5373
rect 692 5356 703 5360
rect 23 5333 103 5344
rect 23 5277 37 5333
rect 93 5277 103 5333
rect 593 5310 703 5356
rect 692 5306 703 5310
rect 757 5306 780 5360
rect 692 5297 780 5306
rect 23 5269 103 5277
rect 351 5244 439 5254
rect 351 5188 362 5244
rect 418 5188 439 5244
rect 351 5176 439 5188
rect -407 4939 -328 4950
rect -407 4883 -397 4939
rect -341 4883 70 4939
rect -407 4875 -328 4883
rect -588 4740 -508 4752
rect -588 4684 -577 4740
rect -521 4684 154 4740
rect -588 4673 -508 4684
rect 574 4386 662 4396
rect 574 4336 588 4386
rect 540 4332 588 4336
rect 642 4332 662 4386
rect 76 4200 122 4327
rect 540 4324 662 4332
rect -408 3970 -329 3981
rect -408 3914 -397 3970
rect -341 3914 70 3970
rect -408 3906 -329 3914
rect -588 3773 -508 3786
rect -588 3717 -577 3773
rect -521 3717 85 3773
rect -588 3707 -508 3717
rect 735 3416 815 3427
rect 735 3412 745 3416
rect 593 3366 745 3412
rect 735 3362 745 3366
rect 799 3362 815 3416
rect 76 3230 122 3355
rect 735 3352 815 3362
rect -408 3000 -329 3008
rect -408 2944 -397 3000
rect -341 2944 69 3000
rect -408 2933 -329 2944
rect -588 2839 -508 2852
rect -588 2783 -577 2839
rect -521 2783 132 2839
rect -588 2773 -508 2783
rect 761 2441 848 2457
rect 761 2437 776 2441
rect -63 2406 16 2417
rect -63 2350 -52 2406
rect 4 2395 16 2406
rect 4 2350 120 2395
rect 591 2391 776 2437
rect 761 2387 776 2391
rect 830 2387 848 2441
rect 761 2381 848 2387
rect -63 2349 120 2350
rect -63 2338 16 2349
rect -237 2281 -156 2292
rect -237 2225 -224 2281
rect -168 2274 -156 2281
rect 76 2274 122 2301
rect -168 2228 122 2274
rect -168 2225 -156 2228
rect -237 2218 -156 2225
rect -411 2013 -332 2022
rect -411 1957 -397 2013
rect -341 1957 67 2013
rect -411 1947 -332 1957
rect -587 1852 -507 1864
rect -587 1796 -577 1852
rect -521 1796 92 1852
rect -587 1785 -507 1796
rect -63 1394 13 1404
rect 76 1394 122 1403
rect -63 1338 -52 1394
rect 4 1338 122 1394
rect -63 1328 13 1338
rect 76 1284 122 1338
rect 587 1212 669 1225
rect 587 1208 600 1212
rect 494 1162 600 1208
rect 587 1158 600 1162
rect 654 1158 669 1212
rect 587 1153 669 1158
rect -411 1041 -332 1051
rect -411 985 -397 1041
rect -341 985 69 1041
rect -411 976 -332 985
rect -587 876 -507 888
rect -587 820 -577 876
rect -521 820 103 876
rect -587 809 -507 820
rect 955 495 1033 504
rect 955 491 966 495
rect 42 464 124 475
rect 42 408 54 464
rect 110 408 124 464
rect 593 445 966 491
rect 955 441 966 445
rect 1020 441 1033 495
rect 955 430 1033 441
rect 42 403 124 408
rect -121 355 -45 357
rect -121 346 122 355
rect -121 290 -110 346
rect -54 309 122 346
rect -54 290 -45 309
rect -121 281 -45 290
rect -408 77 -329 85
rect -408 23 -396 77
rect -342 73 -329 77
rect -342 27 72 73
rect -342 23 -329 27
rect -408 10 -329 23
<< via1 >>
rect -576 8608 -522 8662
rect 624 8242 678 8296
rect -397 7814 -341 7870
rect -577 7631 -521 7687
rect 61 7207 117 7263
rect 613 7257 667 7311
rect -397 6842 -341 6898
rect -577 6660 -521 6716
rect 55 6256 111 6312
rect 886 6281 940 6335
rect 365 6160 421 6216
rect -397 5855 -341 5911
rect -577 5684 -521 5740
rect 37 5277 93 5333
rect 703 5306 757 5360
rect 362 5188 418 5244
rect -397 4883 -341 4939
rect -577 4684 -521 4740
rect 588 4332 642 4386
rect -397 3914 -341 3970
rect -577 3717 -521 3773
rect 745 3362 799 3416
rect -397 2944 -341 3000
rect -577 2783 -521 2839
rect -52 2350 4 2406
rect 776 2387 830 2441
rect -224 2225 -168 2281
rect -397 1957 -341 2013
rect -577 1796 -521 1852
rect -52 1338 4 1394
rect 600 1158 654 1212
rect -397 985 -341 1041
rect -577 820 -521 876
rect 54 408 110 464
rect 966 441 1020 495
rect -110 290 -54 346
rect -396 23 -342 77
<< metal2 >>
rect -590 8662 -510 8677
rect -590 8608 -576 8662
rect -522 8608 -510 8662
rect -590 8598 -510 8608
rect -577 7699 -521 8598
rect 608 8296 694 8306
rect 608 8242 624 8296
rect 678 8242 694 8296
rect 608 8231 694 8242
rect -409 7870 -330 7883
rect -409 7814 -397 7870
rect -341 7814 -330 7870
rect -409 7808 -330 7814
rect -591 7687 -511 7699
rect -591 7631 -577 7687
rect -521 7631 -511 7687
rect -591 7620 -511 7631
rect -577 6728 -521 7620
rect -397 6909 -341 7808
rect 46 7550 132 7564
rect 623 7558 679 8231
rect 46 7494 61 7550
rect 117 7494 132 7550
rect 46 7489 132 7494
rect 610 7550 696 7558
rect 610 7494 623 7550
rect 679 7494 696 7550
rect 61 7267 117 7489
rect 610 7483 696 7494
rect 600 7311 680 7323
rect 49 7263 127 7267
rect 49 7207 61 7263
rect 117 7207 127 7263
rect 600 7257 613 7311
rect 667 7257 680 7311
rect 600 7252 680 7257
rect 49 7196 127 7207
rect -407 6898 -328 6909
rect -407 6842 -397 6898
rect -341 6842 -328 6898
rect -407 6834 -328 6842
rect -592 6716 -512 6728
rect -592 6660 -577 6716
rect -521 6660 -512 6716
rect -592 6649 -512 6660
rect -577 5752 -521 6649
rect -397 5920 -341 6834
rect 44 6568 114 6578
rect 612 6574 668 7252
rect 44 6512 55 6568
rect 111 6512 114 6568
rect 44 6507 114 6512
rect 606 6568 676 6574
rect 606 6512 612 6568
rect 668 6512 676 6568
rect 55 6320 111 6507
rect 606 6503 676 6512
rect 873 6335 953 6347
rect 43 6312 127 6320
rect 43 6256 55 6312
rect 111 6256 127 6312
rect 873 6281 886 6335
rect 940 6281 953 6335
rect 873 6277 953 6281
rect 43 6243 127 6256
rect 352 6216 440 6228
rect 352 6160 365 6216
rect 421 6160 758 6216
rect 352 6152 440 6160
rect -408 5911 -329 5920
rect -408 5855 -397 5911
rect -341 5855 -329 5911
rect -408 5845 -329 5855
rect -589 5740 -509 5752
rect -589 5684 -577 5740
rect -521 5684 -509 5740
rect -589 5673 -509 5684
rect -577 4752 -521 5673
rect -397 4950 -341 5845
rect 702 5373 758 6160
rect 692 5360 780 5373
rect 23 5333 103 5344
rect 23 5277 37 5333
rect 93 5277 103 5333
rect 692 5306 703 5360
rect 757 5306 780 5360
rect 692 5297 780 5306
rect 23 5269 103 5277
rect 37 5055 93 5269
rect 351 5244 439 5253
rect 351 5188 362 5244
rect 418 5188 643 5244
rect 351 5176 439 5188
rect 25 5046 105 5055
rect 25 4990 37 5046
rect 93 4990 105 5046
rect 25 4980 105 4990
rect -407 4939 -328 4950
rect -407 4883 -397 4939
rect -341 4883 -328 4939
rect -407 4875 -328 4883
rect -588 4740 -508 4752
rect -588 4684 -577 4740
rect -521 4684 -508 4740
rect -588 4673 -508 4684
rect -577 3786 -521 4673
rect -397 3981 -341 4875
rect 587 4396 643 5188
rect 738 5046 818 5060
rect 738 4990 744 5046
rect 800 4990 818 5046
rect 738 4985 818 4990
rect 574 4386 662 4396
rect 574 4332 588 4386
rect 642 4332 662 4386
rect 574 4324 662 4332
rect -408 3970 -329 3981
rect -408 3914 -397 3970
rect -341 3914 -329 3970
rect -408 3906 -329 3914
rect -588 3773 -508 3786
rect -588 3717 -577 3773
rect -521 3717 -508 3773
rect -588 3707 -508 3717
rect -577 2852 -521 3707
rect -397 3008 -341 3906
rect 744 3427 800 4985
rect 735 3416 815 3427
rect 735 3362 745 3416
rect 799 3362 815 3416
rect 735 3352 815 3362
rect -408 3000 -329 3008
rect -408 2944 -397 3000
rect -341 2944 -329 3000
rect -408 2933 -329 2944
rect -588 2839 -508 2852
rect -588 2783 -577 2839
rect -521 2783 -508 2839
rect -588 2773 -508 2783
rect -577 1864 -521 2773
rect -397 2022 -341 2933
rect -65 2707 13 2721
rect 885 2711 941 6277
rect -65 2651 -52 2707
rect 4 2651 13 2707
rect -65 2644 13 2651
rect 878 2707 952 2711
rect 878 2651 885 2707
rect 941 2651 952 2707
rect -52 2417 4 2644
rect 878 2641 952 2651
rect 761 2441 848 2457
rect -63 2406 16 2417
rect -63 2350 -52 2406
rect 4 2350 16 2406
rect 761 2387 776 2441
rect 830 2387 848 2441
rect 761 2381 848 2387
rect -63 2338 16 2350
rect -237 2281 -156 2292
rect -237 2225 -224 2281
rect -168 2225 -156 2281
rect -237 2218 -156 2225
rect -411 2013 -332 2022
rect -411 1957 -397 2013
rect -341 1957 -332 2013
rect -411 1947 -332 1957
rect -587 1852 -507 1864
rect -587 1796 -577 1852
rect -521 1796 -507 1852
rect -587 1785 -507 1796
rect -577 888 -521 1785
rect -397 1051 -341 1947
rect -224 1129 -168 2218
rect -52 1404 4 2338
rect -63 1394 13 1404
rect -63 1338 -52 1394
rect 4 1338 13 1394
rect -63 1328 13 1338
rect 587 1212 669 1225
rect 587 1158 600 1212
rect 654 1158 669 1212
rect 587 1153 669 1158
rect -235 1122 -157 1129
rect -235 1066 -224 1122
rect -168 1066 -157 1122
rect -235 1055 -157 1066
rect -411 1041 -332 1051
rect -411 985 -397 1041
rect -341 985 -332 1041
rect -411 976 -332 985
rect -587 876 -507 888
rect -587 820 -577 876
rect -521 820 -507 876
rect -587 809 -507 820
rect -397 85 -341 976
rect -120 944 -44 955
rect -120 888 -110 944
rect -54 888 -44 944
rect -120 879 -44 888
rect -110 357 -54 879
rect 39 746 117 757
rect 599 753 655 1153
rect 775 954 831 2381
rect 953 1122 1031 1132
rect 953 1066 965 1122
rect 1021 1066 1031 1122
rect 953 1058 1031 1066
rect 766 944 842 954
rect 766 888 775 944
rect 831 888 842 944
rect 766 878 842 888
rect 39 690 54 746
rect 110 690 117 746
rect 39 685 117 690
rect 592 746 670 753
rect 592 690 599 746
rect 655 690 670 746
rect 54 475 110 685
rect 592 681 670 690
rect 965 504 1021 1058
rect 955 495 1033 504
rect 42 464 124 475
rect 42 408 54 464
rect 110 408 124 464
rect 955 441 966 495
rect 1020 441 1033 495
rect 955 430 1033 441
rect 42 403 124 408
rect -121 346 -45 357
rect -121 290 -110 346
rect -54 290 -45 346
rect -121 281 -45 290
rect -408 77 -329 85
rect -408 23 -396 77
rect -342 23 -329 77
rect -408 10 -329 23
<< via2 >>
rect 61 7494 117 7550
rect 623 7494 679 7550
rect 55 6512 111 6568
rect 612 6512 668 6568
rect 37 4990 93 5046
rect 744 4990 800 5046
rect -52 2651 4 2707
rect 885 2651 941 2707
rect -224 1066 -168 1122
rect -110 888 -54 944
rect 965 1066 1021 1122
rect 775 888 831 944
rect 54 690 110 746
rect 599 690 655 746
<< metal3 >>
rect 46 7550 132 7564
rect 610 7550 696 7558
rect 46 7494 61 7550
rect 117 7494 623 7550
rect 679 7494 696 7550
rect 46 7489 132 7494
rect 610 7483 696 7494
rect 44 6568 114 6578
rect 606 6568 676 6574
rect 44 6512 55 6568
rect 111 6512 612 6568
rect 668 6512 677 6568
rect 44 6507 114 6512
rect 606 6503 676 6512
rect 25 5046 105 5055
rect 738 5046 818 5060
rect 25 4990 37 5046
rect 93 4990 744 5046
rect 800 4990 818 5046
rect 25 4980 105 4990
rect 738 4985 818 4990
rect -65 2707 13 2721
rect 878 2707 952 2711
rect -65 2651 -52 2707
rect 4 2651 885 2707
rect 941 2651 952 2707
rect -65 2644 13 2651
rect 878 2641 952 2651
rect -235 1122 -157 1129
rect 953 1122 1031 1132
rect -235 1066 -224 1122
rect -168 1066 965 1122
rect 1021 1066 1031 1122
rect -235 1055 -157 1066
rect 953 1058 1031 1066
rect -120 944 -44 955
rect 766 944 842 954
rect -120 888 -110 944
rect -54 888 775 944
rect 831 888 842 944
rect -120 879 -44 888
rect 766 878 842 888
rect 39 746 117 757
rect 592 746 670 753
rect 39 690 54 746
rect 110 690 599 746
rect 655 690 670 746
rect 39 685 117 690
rect 592 681 670 690
use NAND  NAND_0
timestamp 1690283021
transform 1 0 137 0 1 3018
box -86 -97 530 818
use NAND  NAND_1
timestamp 1690283021
transform 1 0 137 0 1 6913
box -86 -97 530 818
use NAND  NAND_2
timestamp 1690283021
transform 1 0 137 0 1 1072
box -86 -97 530 818
use NAND  NAND_3
timestamp 1690283021
transform 1 0 137 0 1 97
box -86 -97 530 818
use NAND  NAND_9
timestamp 1690283021
transform 1 0 137 0 1 2043
box -86 -97 530 818
use NAND  NAND_11
timestamp 1690283021
transform 1 0 137 0 1 3988
box -86 -97 530 818
use NAND  NAND_12
timestamp 1690283021
transform 1 0 137 0 1 4962
box -86 -97 530 818
use NAND  NAND_13
timestamp 1690283021
transform 1 0 137 0 1 5937
box -86 -97 530 818
use NAND  NAND_14
timestamp 1690283021
transform 1 0 137 0 1 7898
box -86 -97 530 818
<< labels >>
flabel via1 990 473 990 473 0 FreeSans 480 0 0 0 QB
port 0 nsew
flabel via1 792 2412 792 2412 0 FreeSans 480 0 0 0 Q
port 1 nsew
flabel metal1 90 8176 90 8176 0 FreeSans 480 0 0 0 Ri-1
port 2 nsew
flabel metal1 93 4257 93 4257 0 FreeSans 480 0 0 0 Ri
port 3 nsew
flabel metal1 93 3298 93 3298 0 FreeSans 480 0 0 0 Ci
port 4 nsew
flabel metal1 80 8650 80 8650 0 FreeSans 480 0 0 0 VDD
port 5 nsew
flabel metal1 0 7850 0 7850 0 FreeSans 480 0 0 0 VSS
port 6 nsew
<< end >>
