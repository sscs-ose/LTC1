magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2410 -2128 2410 2128
<< nwell >>
rect -410 -128 410 128
<< nsubdiff >>
rect -327 23 327 45
rect -327 -23 -305 23
rect 305 -23 327 23
rect -327 -45 327 -23
<< nsubdiffcont >>
rect -305 -23 305 23
<< metal1 >>
rect -316 23 316 34
rect -316 -23 -305 23
rect 305 -23 316 23
rect -316 -34 316 -23
<< end >>
