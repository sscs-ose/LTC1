magic
tech gf180mcuC
magscale 1 10
timestamp 1692387345
<< nwell >>
rect -4898 3321 -845 3789
rect -4898 3243 -3608 3321
rect -1249 3243 -845 3321
rect -4492 3198 -3608 3243
rect -4492 2409 -3608 2532
rect -1249 2409 -845 2487
rect -4492 1611 -845 2409
rect -4492 1488 -3608 1611
rect -1249 1533 -845 1611
rect 22 1534 9082 5906
rect -4492 777 -3608 822
rect -4898 699 -3608 777
rect -1249 699 -845 777
rect -4898 -99 -845 699
rect -4898 -177 -3608 -99
rect -1249 -177 -845 -99
rect -4492 -222 -3608 -177
rect -4492 -1011 -3608 -888
rect -1249 -1011 -845 -933
rect -4492 -1479 -845 -1011
rect -4175 -5794 -551 -3548
rect 22 -5794 9082 -1422
<< pwell >>
rect 84 6010 1484 7168
rect 1492 6010 1772 7168
rect 1896 6010 2176 7168
rect 2184 6010 3584 7168
rect 3708 6010 3988 7168
rect 3996 6010 5396 7168
rect 5520 6010 5800 7168
rect 5808 6010 7208 7168
rect 7332 6010 7612 7168
rect 7620 6010 9020 7168
rect -4836 2933 -4556 3169
rect -4270 2921 -3830 3157
rect -3565 2916 -2885 3110
rect -2779 2916 -2099 3110
rect -1993 2916 -1313 3110
rect -1187 2933 -907 3169
rect -4270 2573 -3830 2809
rect -3565 2620 -2885 2814
rect -2779 2620 -2099 2814
rect -1993 2620 -1313 2814
rect -1187 2561 -907 2797
rect -4270 1211 -3830 1447
rect -3565 1206 -2885 1400
rect -2779 1206 -2099 1400
rect -1993 1206 -1313 1400
rect -1187 1223 -907 1459
rect -4836 851 -4556 1087
rect -4270 863 -3830 1099
rect -3565 910 -2885 1104
rect -2779 910 -2099 1104
rect -1993 910 -1313 1104
rect -1187 851 -907 1087
rect 84 272 364 1430
rect 372 272 1772 1430
rect 1896 272 3296 1430
rect 3304 272 3584 1430
rect 3708 272 3988 1430
rect 3996 272 5396 1430
rect 5520 272 6920 1430
rect 6928 272 7208 1430
rect 7332 272 8732 1430
rect 8740 272 9020 1430
rect -4836 -487 -4556 -251
rect -4270 -499 -3830 -263
rect -3565 -504 -2885 -310
rect -2779 -504 -2099 -310
rect -1993 -504 -1313 -310
rect -1187 -487 -907 -251
rect -4270 -847 -3830 -611
rect -3565 -800 -2885 -606
rect -2779 -800 -2099 -606
rect -1993 -800 -1313 -606
rect -1187 -859 -907 -623
rect 84 -1318 364 -160
rect 372 -1318 1772 -160
rect 1896 -1318 3296 -160
rect 3304 -1318 3584 -160
rect 3708 -1318 3988 -160
rect 3996 -1318 5396 -160
rect 5520 -1318 6920 -160
rect 6928 -1318 7208 -160
rect 7332 -1318 8732 -160
rect 8740 -1318 9020 -160
rect -4113 -7056 -3833 -5898
rect -3825 -7056 -2425 -5898
rect -2301 -7056 -901 -5898
rect -893 -7056 -613 -5898
rect 84 -7056 364 -5898
rect 372 -7056 1772 -5898
rect 1896 -7056 3296 -5898
rect 3304 -7056 3584 -5898
rect 3708 -7056 3988 -5898
rect 3996 -7056 5396 -5898
rect 5520 -7056 6920 -5898
rect 6928 -7056 7208 -5898
rect 7332 -7056 8732 -5898
rect 8740 -7056 9020 -5898
<< nmos >>
rect 196 6850 252 7100
rect 356 6850 412 7100
rect 516 6850 572 7100
rect 676 6850 732 7100
rect 836 6850 892 7100
rect 996 6850 1052 7100
rect 1156 6850 1212 7100
rect 1316 6850 1372 7100
rect 1604 6850 1660 7100
rect 2008 6850 2064 7100
rect 2296 6850 2352 7100
rect 2456 6850 2512 7100
rect 2616 6850 2672 7100
rect 2776 6850 2832 7100
rect 2936 6850 2992 7100
rect 3096 6850 3152 7100
rect 3256 6850 3312 7100
rect 3416 6850 3472 7100
rect 3820 6850 3876 7100
rect 4108 6850 4164 7100
rect 4268 6850 4324 7100
rect 4428 6850 4484 7100
rect 4588 6850 4644 7100
rect 4748 6850 4804 7100
rect 4908 6850 4964 7100
rect 5068 6850 5124 7100
rect 5228 6850 5284 7100
rect 5632 6850 5688 7100
rect 5920 6850 5976 7100
rect 6080 6850 6136 7100
rect 6240 6850 6296 7100
rect 6400 6850 6456 7100
rect 6560 6850 6616 7100
rect 6720 6850 6776 7100
rect 6880 6850 6936 7100
rect 7040 6850 7096 7100
rect 7444 6850 7500 7100
rect 7732 6850 7788 7100
rect 7892 6850 7948 7100
rect 8052 6850 8108 7100
rect 8212 6850 8268 7100
rect 8372 6850 8428 7100
rect 8532 6850 8588 7100
rect 8692 6850 8748 7100
rect 8852 6850 8908 7100
rect 196 6464 252 6714
rect 356 6464 412 6714
rect 516 6464 572 6714
rect 676 6464 732 6714
rect 836 6464 892 6714
rect 996 6464 1052 6714
rect 1156 6464 1212 6714
rect 1316 6464 1372 6714
rect 1604 6464 1660 6714
rect 2008 6464 2064 6714
rect 2296 6464 2352 6714
rect 2456 6464 2512 6714
rect 2616 6464 2672 6714
rect 2776 6464 2832 6714
rect 2936 6464 2992 6714
rect 3096 6464 3152 6714
rect 3256 6464 3312 6714
rect 3416 6464 3472 6714
rect 3820 6464 3876 6714
rect 4108 6464 4164 6714
rect 4268 6464 4324 6714
rect 4428 6464 4484 6714
rect 4588 6464 4644 6714
rect 4748 6464 4804 6714
rect 4908 6464 4964 6714
rect 5068 6464 5124 6714
rect 5228 6464 5284 6714
rect 5632 6464 5688 6714
rect 5920 6464 5976 6714
rect 6080 6464 6136 6714
rect 6240 6464 6296 6714
rect 6400 6464 6456 6714
rect 6560 6464 6616 6714
rect 6720 6464 6776 6714
rect 6880 6464 6936 6714
rect 7040 6464 7096 6714
rect 7444 6464 7500 6714
rect 7732 6464 7788 6714
rect 7892 6464 7948 6714
rect 8052 6464 8108 6714
rect 8212 6464 8268 6714
rect 8372 6464 8428 6714
rect 8532 6464 8588 6714
rect 8692 6464 8748 6714
rect 8852 6464 8908 6714
rect 196 6078 252 6328
rect 356 6078 412 6328
rect 516 6078 572 6328
rect 676 6078 732 6328
rect 836 6078 892 6328
rect 996 6078 1052 6328
rect 1156 6078 1212 6328
rect 1316 6078 1372 6328
rect 1604 6078 1660 6328
rect 2008 6078 2064 6328
rect 2296 6078 2352 6328
rect 2456 6078 2512 6328
rect 2616 6078 2672 6328
rect 2776 6078 2832 6328
rect 2936 6078 2992 6328
rect 3096 6078 3152 6328
rect 3256 6078 3312 6328
rect 3416 6078 3472 6328
rect 3820 6078 3876 6328
rect 4108 6078 4164 6328
rect 4268 6078 4324 6328
rect 4428 6078 4484 6328
rect 4588 6078 4644 6328
rect 4748 6078 4804 6328
rect 4908 6078 4964 6328
rect 5068 6078 5124 6328
rect 5228 6078 5284 6328
rect 5632 6078 5688 6328
rect 5920 6078 5976 6328
rect 6080 6078 6136 6328
rect 6240 6078 6296 6328
rect 6400 6078 6456 6328
rect 6560 6078 6616 6328
rect 6720 6078 6776 6328
rect 6880 6078 6936 6328
rect 7040 6078 7096 6328
rect 7444 6078 7500 6328
rect 7732 6078 7788 6328
rect 7892 6078 7948 6328
rect 8052 6078 8108 6328
rect 8212 6078 8268 6328
rect 8372 6078 8428 6328
rect 8532 6078 8588 6328
rect 8692 6078 8748 6328
rect 8852 6078 8908 6328
rect -4724 3001 -4668 3101
rect -4158 2989 -4102 3089
rect -3998 2989 -3942 3089
rect -3449 2991 -3001 3035
rect -2663 2991 -2215 3035
rect -1877 2991 -1429 3035
rect -1075 3001 -1019 3101
rect -4158 2641 -4102 2741
rect -3998 2641 -3942 2741
rect -3449 2695 -3001 2739
rect -2663 2695 -2215 2739
rect -1877 2695 -1429 2739
rect -1075 2629 -1019 2729
rect -4158 1279 -4102 1379
rect -3998 1279 -3942 1379
rect -3449 1281 -3001 1325
rect -2663 1281 -2215 1325
rect -1877 1281 -1429 1325
rect -1075 1291 -1019 1391
rect 196 1112 252 1362
rect 484 1112 540 1362
rect 644 1112 700 1362
rect 804 1112 860 1362
rect 964 1112 1020 1362
rect 1124 1112 1180 1362
rect 1284 1112 1340 1362
rect 1444 1112 1500 1362
rect 1604 1112 1660 1362
rect 2008 1112 2064 1362
rect 2168 1112 2224 1362
rect 2328 1112 2384 1362
rect 2488 1112 2544 1362
rect 2648 1112 2704 1362
rect 2808 1112 2864 1362
rect 2968 1112 3024 1362
rect 3128 1112 3184 1362
rect 3416 1112 3472 1362
rect 3820 1112 3876 1362
rect 4108 1112 4164 1362
rect 4268 1112 4324 1362
rect 4428 1112 4484 1362
rect 4588 1112 4644 1362
rect 4748 1112 4804 1362
rect 4908 1112 4964 1362
rect 5068 1112 5124 1362
rect 5228 1112 5284 1362
rect 5632 1112 5688 1362
rect 5792 1112 5848 1362
rect 5952 1112 6008 1362
rect 6112 1112 6168 1362
rect 6272 1112 6328 1362
rect 6432 1112 6488 1362
rect 6592 1112 6648 1362
rect 6752 1112 6808 1362
rect 7040 1112 7096 1362
rect 7444 1112 7500 1362
rect 7604 1112 7660 1362
rect 7764 1112 7820 1362
rect 7924 1112 7980 1362
rect 8084 1112 8140 1362
rect 8244 1112 8300 1362
rect 8404 1112 8460 1362
rect 8564 1112 8620 1362
rect 8852 1112 8908 1362
rect -4724 919 -4668 1019
rect -4158 931 -4102 1031
rect -3998 931 -3942 1031
rect -3449 985 -3001 1029
rect -2663 985 -2215 1029
rect -1877 985 -1429 1029
rect -1075 919 -1019 1019
rect 196 726 252 976
rect 484 726 540 976
rect 644 726 700 976
rect 804 726 860 976
rect 964 726 1020 976
rect 1124 726 1180 976
rect 1284 726 1340 976
rect 1444 726 1500 976
rect 1604 726 1660 976
rect 2008 726 2064 976
rect 2168 726 2224 976
rect 2328 726 2384 976
rect 2488 726 2544 976
rect 2648 726 2704 976
rect 2808 726 2864 976
rect 2968 726 3024 976
rect 3128 726 3184 976
rect 3416 726 3472 976
rect 3820 726 3876 976
rect 4108 726 4164 976
rect 4268 726 4324 976
rect 4428 726 4484 976
rect 4588 726 4644 976
rect 4748 726 4804 976
rect 4908 726 4964 976
rect 5068 726 5124 976
rect 5228 726 5284 976
rect 5632 726 5688 976
rect 5792 726 5848 976
rect 5952 726 6008 976
rect 6112 726 6168 976
rect 6272 726 6328 976
rect 6432 726 6488 976
rect 6592 726 6648 976
rect 6752 726 6808 976
rect 7040 726 7096 976
rect 7444 726 7500 976
rect 7604 726 7660 976
rect 7764 726 7820 976
rect 7924 726 7980 976
rect 8084 726 8140 976
rect 8244 726 8300 976
rect 8404 726 8460 976
rect 8564 726 8620 976
rect 8852 726 8908 976
rect 196 340 252 590
rect 484 340 540 590
rect 644 340 700 590
rect 804 340 860 590
rect 964 340 1020 590
rect 1124 340 1180 590
rect 1284 340 1340 590
rect 1444 340 1500 590
rect 1604 340 1660 590
rect 2008 340 2064 590
rect 2168 340 2224 590
rect 2328 340 2384 590
rect 2488 340 2544 590
rect 2648 340 2704 590
rect 2808 340 2864 590
rect 2968 340 3024 590
rect 3128 340 3184 590
rect 3416 340 3472 590
rect 3820 340 3876 590
rect 4108 340 4164 590
rect 4268 340 4324 590
rect 4428 340 4484 590
rect 4588 340 4644 590
rect 4748 340 4804 590
rect 4908 340 4964 590
rect 5068 340 5124 590
rect 5228 340 5284 590
rect 5632 340 5688 590
rect 5792 340 5848 590
rect 5952 340 6008 590
rect 6112 340 6168 590
rect 6272 340 6328 590
rect 6432 340 6488 590
rect 6592 340 6648 590
rect 6752 340 6808 590
rect 7040 340 7096 590
rect 7444 340 7500 590
rect 7604 340 7660 590
rect 7764 340 7820 590
rect 7924 340 7980 590
rect 8084 340 8140 590
rect 8244 340 8300 590
rect 8404 340 8460 590
rect 8564 340 8620 590
rect 8852 340 8908 590
rect -4724 -419 -4668 -319
rect -4158 -431 -4102 -331
rect -3998 -431 -3942 -331
rect -3449 -429 -3001 -385
rect -2663 -429 -2215 -385
rect -1877 -429 -1429 -385
rect -1075 -419 -1019 -319
rect 196 -478 252 -228
rect 484 -478 540 -228
rect 644 -478 700 -228
rect 804 -478 860 -228
rect 964 -478 1020 -228
rect 1124 -478 1180 -228
rect 1284 -478 1340 -228
rect 1444 -478 1500 -228
rect 1604 -478 1660 -228
rect 2008 -478 2064 -228
rect 2168 -478 2224 -228
rect 2328 -478 2384 -228
rect 2488 -478 2544 -228
rect 2648 -478 2704 -228
rect 2808 -478 2864 -228
rect 2968 -478 3024 -228
rect 3128 -478 3184 -228
rect 3416 -478 3472 -228
rect 3820 -478 3876 -228
rect 4108 -478 4164 -228
rect 4268 -478 4324 -228
rect 4428 -478 4484 -228
rect 4588 -478 4644 -228
rect 4748 -478 4804 -228
rect 4908 -478 4964 -228
rect 5068 -478 5124 -228
rect 5228 -478 5284 -228
rect 5632 -478 5688 -228
rect 5792 -478 5848 -228
rect 5952 -478 6008 -228
rect 6112 -478 6168 -228
rect 6272 -478 6328 -228
rect 6432 -478 6488 -228
rect 6592 -478 6648 -228
rect 6752 -478 6808 -228
rect 7040 -478 7096 -228
rect 7444 -478 7500 -228
rect 7604 -478 7660 -228
rect 7764 -478 7820 -228
rect 7924 -478 7980 -228
rect 8084 -478 8140 -228
rect 8244 -478 8300 -228
rect 8404 -478 8460 -228
rect 8564 -478 8620 -228
rect 8852 -478 8908 -228
rect -4158 -779 -4102 -679
rect -3998 -779 -3942 -679
rect -3449 -725 -3001 -681
rect -2663 -725 -2215 -681
rect -1877 -725 -1429 -681
rect -1075 -791 -1019 -691
rect 196 -864 252 -614
rect 484 -864 540 -614
rect 644 -864 700 -614
rect 804 -864 860 -614
rect 964 -864 1020 -614
rect 1124 -864 1180 -614
rect 1284 -864 1340 -614
rect 1444 -864 1500 -614
rect 1604 -864 1660 -614
rect 2008 -864 2064 -614
rect 2168 -864 2224 -614
rect 2328 -864 2384 -614
rect 2488 -864 2544 -614
rect 2648 -864 2704 -614
rect 2808 -864 2864 -614
rect 2968 -864 3024 -614
rect 3128 -864 3184 -614
rect 3416 -864 3472 -614
rect 3820 -864 3876 -614
rect 4108 -864 4164 -614
rect 4268 -864 4324 -614
rect 4428 -864 4484 -614
rect 4588 -864 4644 -614
rect 4748 -864 4804 -614
rect 4908 -864 4964 -614
rect 5068 -864 5124 -614
rect 5228 -864 5284 -614
rect 5632 -864 5688 -614
rect 5792 -864 5848 -614
rect 5952 -864 6008 -614
rect 6112 -864 6168 -614
rect 6272 -864 6328 -614
rect 6432 -864 6488 -614
rect 6592 -864 6648 -614
rect 6752 -864 6808 -614
rect 7040 -864 7096 -614
rect 7444 -864 7500 -614
rect 7604 -864 7660 -614
rect 7764 -864 7820 -614
rect 7924 -864 7980 -614
rect 8084 -864 8140 -614
rect 8244 -864 8300 -614
rect 8404 -864 8460 -614
rect 8564 -864 8620 -614
rect 8852 -864 8908 -614
rect 196 -1250 252 -1000
rect 484 -1250 540 -1000
rect 644 -1250 700 -1000
rect 804 -1250 860 -1000
rect 964 -1250 1020 -1000
rect 1124 -1250 1180 -1000
rect 1284 -1250 1340 -1000
rect 1444 -1250 1500 -1000
rect 1604 -1250 1660 -1000
rect 2008 -1250 2064 -1000
rect 2168 -1250 2224 -1000
rect 2328 -1250 2384 -1000
rect 2488 -1250 2544 -1000
rect 2648 -1250 2704 -1000
rect 2808 -1250 2864 -1000
rect 2968 -1250 3024 -1000
rect 3128 -1250 3184 -1000
rect 3416 -1250 3472 -1000
rect 3820 -1250 3876 -1000
rect 4108 -1250 4164 -1000
rect 4268 -1250 4324 -1000
rect 4428 -1250 4484 -1000
rect 4588 -1250 4644 -1000
rect 4748 -1250 4804 -1000
rect 4908 -1250 4964 -1000
rect 5068 -1250 5124 -1000
rect 5228 -1250 5284 -1000
rect 5632 -1250 5688 -1000
rect 5792 -1250 5848 -1000
rect 5952 -1250 6008 -1000
rect 6112 -1250 6168 -1000
rect 6272 -1250 6328 -1000
rect 6432 -1250 6488 -1000
rect 6592 -1250 6648 -1000
rect 6752 -1250 6808 -1000
rect 7040 -1250 7096 -1000
rect 7444 -1250 7500 -1000
rect 7604 -1250 7660 -1000
rect 7764 -1250 7820 -1000
rect 7924 -1250 7980 -1000
rect 8084 -1250 8140 -1000
rect 8244 -1250 8300 -1000
rect 8404 -1250 8460 -1000
rect 8564 -1250 8620 -1000
rect 8852 -1250 8908 -1000
rect -4001 -6216 -3945 -5966
rect -3713 -6216 -3657 -5966
rect -3553 -6216 -3497 -5966
rect -3393 -6216 -3337 -5966
rect -3233 -6216 -3177 -5966
rect -3073 -6216 -3017 -5966
rect -2913 -6216 -2857 -5966
rect -2753 -6216 -2697 -5966
rect -2593 -6216 -2537 -5966
rect -2189 -6216 -2133 -5966
rect -2029 -6216 -1973 -5966
rect -1869 -6216 -1813 -5966
rect -1709 -6216 -1653 -5966
rect -1549 -6216 -1493 -5966
rect -1389 -6216 -1333 -5966
rect -1229 -6216 -1173 -5966
rect -1069 -6216 -1013 -5966
rect -781 -6216 -725 -5966
rect 196 -6216 252 -5966
rect 484 -6216 540 -5966
rect 644 -6216 700 -5966
rect 804 -6216 860 -5966
rect 964 -6216 1020 -5966
rect 1124 -6216 1180 -5966
rect 1284 -6216 1340 -5966
rect 1444 -6216 1500 -5966
rect 1604 -6216 1660 -5966
rect 2008 -6216 2064 -5966
rect 2168 -6216 2224 -5966
rect 2328 -6216 2384 -5966
rect 2488 -6216 2544 -5966
rect 2648 -6216 2704 -5966
rect 2808 -6216 2864 -5966
rect 2968 -6216 3024 -5966
rect 3128 -6216 3184 -5966
rect 3416 -6216 3472 -5966
rect 3820 -6216 3876 -5966
rect 4108 -6216 4164 -5966
rect 4268 -6216 4324 -5966
rect 4428 -6216 4484 -5966
rect 4588 -6216 4644 -5966
rect 4748 -6216 4804 -5966
rect 4908 -6216 4964 -5966
rect 5068 -6216 5124 -5966
rect 5228 -6216 5284 -5966
rect 5632 -6216 5688 -5966
rect 5792 -6216 5848 -5966
rect 5952 -6216 6008 -5966
rect 6112 -6216 6168 -5966
rect 6272 -6216 6328 -5966
rect 6432 -6216 6488 -5966
rect 6592 -6216 6648 -5966
rect 6752 -6216 6808 -5966
rect 7040 -6216 7096 -5966
rect 7444 -6216 7500 -5966
rect 7604 -6216 7660 -5966
rect 7764 -6216 7820 -5966
rect 7924 -6216 7980 -5966
rect 8084 -6216 8140 -5966
rect 8244 -6216 8300 -5966
rect 8404 -6216 8460 -5966
rect 8564 -6216 8620 -5966
rect 8852 -6216 8908 -5966
rect -4001 -6602 -3945 -6352
rect -3713 -6602 -3657 -6352
rect -3553 -6602 -3497 -6352
rect -3393 -6602 -3337 -6352
rect -3233 -6602 -3177 -6352
rect -3073 -6602 -3017 -6352
rect -2913 -6602 -2857 -6352
rect -2753 -6602 -2697 -6352
rect -2593 -6602 -2537 -6352
rect -2189 -6602 -2133 -6352
rect -2029 -6602 -1973 -6352
rect -1869 -6602 -1813 -6352
rect -1709 -6602 -1653 -6352
rect -1549 -6602 -1493 -6352
rect -1389 -6602 -1333 -6352
rect -1229 -6602 -1173 -6352
rect -1069 -6602 -1013 -6352
rect -781 -6602 -725 -6352
rect 196 -6602 252 -6352
rect 484 -6602 540 -6352
rect 644 -6602 700 -6352
rect 804 -6602 860 -6352
rect 964 -6602 1020 -6352
rect 1124 -6602 1180 -6352
rect 1284 -6602 1340 -6352
rect 1444 -6602 1500 -6352
rect 1604 -6602 1660 -6352
rect 2008 -6602 2064 -6352
rect 2168 -6602 2224 -6352
rect 2328 -6602 2384 -6352
rect 2488 -6602 2544 -6352
rect 2648 -6602 2704 -6352
rect 2808 -6602 2864 -6352
rect 2968 -6602 3024 -6352
rect 3128 -6602 3184 -6352
rect 3416 -6602 3472 -6352
rect 3820 -6602 3876 -6352
rect 4108 -6602 4164 -6352
rect 4268 -6602 4324 -6352
rect 4428 -6602 4484 -6352
rect 4588 -6602 4644 -6352
rect 4748 -6602 4804 -6352
rect 4908 -6602 4964 -6352
rect 5068 -6602 5124 -6352
rect 5228 -6602 5284 -6352
rect 5632 -6602 5688 -6352
rect 5792 -6602 5848 -6352
rect 5952 -6602 6008 -6352
rect 6112 -6602 6168 -6352
rect 6272 -6602 6328 -6352
rect 6432 -6602 6488 -6352
rect 6592 -6602 6648 -6352
rect 6752 -6602 6808 -6352
rect 7040 -6602 7096 -6352
rect 7444 -6602 7500 -6352
rect 7604 -6602 7660 -6352
rect 7764 -6602 7820 -6352
rect 7924 -6602 7980 -6352
rect 8084 -6602 8140 -6352
rect 8244 -6602 8300 -6352
rect 8404 -6602 8460 -6352
rect 8564 -6602 8620 -6352
rect 8852 -6602 8908 -6352
rect -4001 -6988 -3945 -6738
rect -3713 -6988 -3657 -6738
rect -3553 -6988 -3497 -6738
rect -3393 -6988 -3337 -6738
rect -3233 -6988 -3177 -6738
rect -3073 -6988 -3017 -6738
rect -2913 -6988 -2857 -6738
rect -2753 -6988 -2697 -6738
rect -2593 -6988 -2537 -6738
rect -2189 -6988 -2133 -6738
rect -2029 -6988 -1973 -6738
rect -1869 -6988 -1813 -6738
rect -1709 -6988 -1653 -6738
rect -1549 -6988 -1493 -6738
rect -1389 -6988 -1333 -6738
rect -1229 -6988 -1173 -6738
rect -1069 -6988 -1013 -6738
rect -781 -6988 -725 -6738
rect 196 -6988 252 -6738
rect 484 -6988 540 -6738
rect 644 -6988 700 -6738
rect 804 -6988 860 -6738
rect 964 -6988 1020 -6738
rect 1124 -6988 1180 -6738
rect 1284 -6988 1340 -6738
rect 1444 -6988 1500 -6738
rect 1604 -6988 1660 -6738
rect 2008 -6988 2064 -6738
rect 2168 -6988 2224 -6738
rect 2328 -6988 2384 -6738
rect 2488 -6988 2544 -6738
rect 2648 -6988 2704 -6738
rect 2808 -6988 2864 -6738
rect 2968 -6988 3024 -6738
rect 3128 -6988 3184 -6738
rect 3416 -6988 3472 -6738
rect 3820 -6988 3876 -6738
rect 4108 -6988 4164 -6738
rect 4268 -6988 4324 -6738
rect 4428 -6988 4484 -6738
rect 4588 -6988 4644 -6738
rect 4748 -6988 4804 -6738
rect 4908 -6988 4964 -6738
rect 5068 -6988 5124 -6738
rect 5228 -6988 5284 -6738
rect 5632 -6988 5688 -6738
rect 5792 -6988 5848 -6738
rect 5952 -6988 6008 -6738
rect 6112 -6988 6168 -6738
rect 6272 -6988 6328 -6738
rect 6432 -6988 6488 -6738
rect 6592 -6988 6648 -6738
rect 6752 -6988 6808 -6738
rect 7040 -6988 7096 -6738
rect 7444 -6988 7500 -6738
rect 7604 -6988 7660 -6738
rect 7764 -6988 7820 -6738
rect 7924 -6988 7980 -6738
rect 8084 -6988 8140 -6738
rect 8244 -6988 8300 -6738
rect 8404 -6988 8460 -6738
rect 8564 -6988 8620 -6738
rect 8852 -6988 8908 -6738
<< pmos >>
rect 196 5276 252 5776
rect 356 5276 412 5776
rect 516 5276 572 5776
rect 676 5276 732 5776
rect 836 5276 892 5776
rect 996 5276 1052 5776
rect 1156 5276 1212 5776
rect 1316 5276 1372 5776
rect 1604 5276 1660 5776
rect 2008 5276 2064 5776
rect 2296 5276 2352 5776
rect 2456 5276 2512 5776
rect 2616 5276 2672 5776
rect 2776 5276 2832 5776
rect 2936 5276 2992 5776
rect 3096 5276 3152 5776
rect 3256 5276 3312 5776
rect 3416 5276 3472 5776
rect 3820 5276 3876 5776
rect 4108 5276 4164 5776
rect 4268 5276 4324 5776
rect 4428 5276 4484 5776
rect 4588 5276 4644 5776
rect 4748 5276 4804 5776
rect 4908 5276 4964 5776
rect 5068 5276 5124 5776
rect 5228 5276 5284 5776
rect 5632 5276 5688 5776
rect 5920 5276 5976 5776
rect 6080 5276 6136 5776
rect 6240 5276 6296 5776
rect 6400 5276 6456 5776
rect 6560 5276 6616 5776
rect 6720 5276 6776 5776
rect 6880 5276 6936 5776
rect 7040 5276 7096 5776
rect 7444 5276 7500 5776
rect 7732 5276 7788 5776
rect 7892 5276 7948 5776
rect 8052 5276 8108 5776
rect 8212 5276 8268 5776
rect 8372 5276 8428 5776
rect 8532 5276 8588 5776
rect 8692 5276 8748 5776
rect 8852 5276 8908 5776
rect 196 4640 252 5140
rect 356 4640 412 5140
rect 516 4640 572 5140
rect 676 4640 732 5140
rect 836 4640 892 5140
rect 996 4640 1052 5140
rect 1156 4640 1212 5140
rect 1316 4640 1372 5140
rect 1604 4640 1660 5140
rect 2008 4640 2064 5140
rect 2296 4640 2352 5140
rect 2456 4640 2512 5140
rect 2616 4640 2672 5140
rect 2776 4640 2832 5140
rect 2936 4640 2992 5140
rect 3096 4640 3152 5140
rect 3256 4640 3312 5140
rect 3416 4640 3472 5140
rect 3820 4640 3876 5140
rect 4108 4640 4164 5140
rect 4268 4640 4324 5140
rect 4428 4640 4484 5140
rect 4588 4640 4644 5140
rect 4748 4640 4804 5140
rect 4908 4640 4964 5140
rect 5068 4640 5124 5140
rect 5228 4640 5284 5140
rect 5632 4640 5688 5140
rect 5920 4640 5976 5140
rect 6080 4640 6136 5140
rect 6240 4640 6296 5140
rect 6400 4640 6456 5140
rect 6560 4640 6616 5140
rect 6720 4640 6776 5140
rect 6880 4640 6936 5140
rect 7040 4640 7096 5140
rect 7444 4640 7500 5140
rect 7732 4640 7788 5140
rect 7892 4640 7948 5140
rect 8052 4640 8108 5140
rect 8212 4640 8268 5140
rect 8372 4640 8428 5140
rect 8532 4640 8588 5140
rect 8692 4640 8748 5140
rect 8852 4640 8908 5140
rect 196 4004 252 4504
rect 356 4004 412 4504
rect 516 4004 572 4504
rect 676 4004 732 4504
rect 836 4004 892 4504
rect 996 4004 1052 4504
rect 1156 4004 1212 4504
rect 1316 4004 1372 4504
rect 1604 4004 1660 4504
rect 2008 4004 2064 4504
rect 2296 4004 2352 4504
rect 2456 4004 2512 4504
rect 2616 4004 2672 4504
rect 2776 4004 2832 4504
rect 2936 4004 2992 4504
rect 3096 4004 3152 4504
rect 3256 4004 3312 4504
rect 3416 4004 3472 4504
rect 3820 4004 3876 4504
rect 4108 4004 4164 4504
rect 4268 4004 4324 4504
rect 4428 4004 4484 4504
rect 4588 4004 4644 4504
rect 4748 4004 4804 4504
rect 4908 4004 4964 4504
rect 5068 4004 5124 4504
rect 5228 4004 5284 4504
rect 5632 4004 5688 4504
rect 5920 4004 5976 4504
rect 6080 4004 6136 4504
rect 6240 4004 6296 4504
rect 6400 4004 6456 4504
rect 6560 4004 6616 4504
rect 6720 4004 6776 4504
rect 6880 4004 6936 4504
rect 7040 4004 7096 4504
rect 7444 4004 7500 4504
rect 7732 4004 7788 4504
rect 7892 4004 7948 4504
rect 8052 4004 8108 4504
rect 8212 4004 8268 4504
rect 8372 4004 8428 4504
rect 8532 4004 8588 4504
rect 8692 4004 8748 4504
rect 8852 4004 8908 4504
rect -4724 3373 -4668 3573
rect -4318 3328 -4262 3528
rect -4158 3328 -4102 3528
rect -3998 3328 -3942 3528
rect -3838 3328 -3782 3528
rect -3445 3451 -2997 3539
rect -2659 3451 -2211 3539
rect -1873 3451 -1425 3539
rect -1075 3373 -1019 3573
rect 196 2936 252 3436
rect 484 2936 540 3436
rect 644 2936 700 3436
rect 804 2936 860 3436
rect 964 2936 1020 3436
rect 1124 2936 1180 3436
rect 1284 2936 1340 3436
rect 1444 2936 1500 3436
rect 1604 2936 1660 3436
rect 2008 2936 2064 3436
rect 2168 2936 2224 3436
rect 2328 2936 2384 3436
rect 2488 2936 2544 3436
rect 2648 2936 2704 3436
rect 2808 2936 2864 3436
rect 2968 2936 3024 3436
rect 3128 2936 3184 3436
rect 3416 2936 3472 3436
rect 3820 2936 3876 3436
rect 4108 2936 4164 3436
rect 4268 2936 4324 3436
rect 4428 2936 4484 3436
rect 4588 2936 4644 3436
rect 4748 2936 4804 3436
rect 4908 2936 4964 3436
rect 5068 2936 5124 3436
rect 5228 2936 5284 3436
rect 5632 2936 5688 3436
rect 5792 2936 5848 3436
rect 5952 2936 6008 3436
rect 6112 2936 6168 3436
rect 6272 2936 6328 3436
rect 6432 2936 6488 3436
rect 6592 2936 6648 3436
rect 6752 2936 6808 3436
rect 7040 2936 7096 3436
rect 7444 2936 7500 3436
rect 7604 2936 7660 3436
rect 7764 2936 7820 3436
rect 7924 2936 7980 3436
rect 8084 2936 8140 3436
rect 8244 2936 8300 3436
rect 8404 2936 8460 3436
rect 8564 2936 8620 3436
rect 8852 2936 8908 3436
rect -4318 2202 -4262 2402
rect -4158 2202 -4102 2402
rect -3998 2202 -3942 2402
rect -3838 2202 -3782 2402
rect -3445 2191 -2997 2279
rect -2659 2191 -2211 2279
rect -1873 2191 -1425 2279
rect -1075 2157 -1019 2357
rect 196 2300 252 2800
rect 484 2300 540 2800
rect 644 2300 700 2800
rect 804 2300 860 2800
rect 964 2300 1020 2800
rect 1124 2300 1180 2800
rect 1284 2300 1340 2800
rect 1444 2300 1500 2800
rect 1604 2300 1660 2800
rect 2008 2300 2064 2800
rect 2168 2300 2224 2800
rect 2328 2300 2384 2800
rect 2488 2300 2544 2800
rect 2648 2300 2704 2800
rect 2808 2300 2864 2800
rect 2968 2300 3024 2800
rect 3128 2300 3184 2800
rect 3416 2300 3472 2800
rect 3820 2300 3876 2800
rect 4108 2300 4164 2800
rect 4268 2300 4324 2800
rect 4428 2300 4484 2800
rect 4588 2300 4644 2800
rect 4748 2300 4804 2800
rect 4908 2300 4964 2800
rect 5068 2300 5124 2800
rect 5228 2300 5284 2800
rect 5632 2300 5688 2800
rect 5792 2300 5848 2800
rect 5952 2300 6008 2800
rect 6112 2300 6168 2800
rect 6272 2300 6328 2800
rect 6432 2300 6488 2800
rect 6592 2300 6648 2800
rect 6752 2300 6808 2800
rect 7040 2300 7096 2800
rect 7444 2300 7500 2800
rect 7604 2300 7660 2800
rect 7764 2300 7820 2800
rect 7924 2300 7980 2800
rect 8084 2300 8140 2800
rect 8244 2300 8300 2800
rect 8404 2300 8460 2800
rect 8564 2300 8620 2800
rect 8852 2300 8908 2800
rect -4318 1618 -4262 1818
rect -4158 1618 -4102 1818
rect -3998 1618 -3942 1818
rect -3838 1618 -3782 1818
rect -3445 1741 -2997 1829
rect -2659 1741 -2211 1829
rect -1873 1741 -1425 1829
rect -1075 1663 -1019 1863
rect 196 1664 252 2164
rect 484 1664 540 2164
rect 644 1664 700 2164
rect 804 1664 860 2164
rect 964 1664 1020 2164
rect 1124 1664 1180 2164
rect 1284 1664 1340 2164
rect 1444 1664 1500 2164
rect 1604 1664 1660 2164
rect 2008 1664 2064 2164
rect 2168 1664 2224 2164
rect 2328 1664 2384 2164
rect 2488 1664 2544 2164
rect 2648 1664 2704 2164
rect 2808 1664 2864 2164
rect 2968 1664 3024 2164
rect 3128 1664 3184 2164
rect 3416 1664 3472 2164
rect 3820 1664 3876 2164
rect 4108 1664 4164 2164
rect 4268 1664 4324 2164
rect 4428 1664 4484 2164
rect 4588 1664 4644 2164
rect 4748 1664 4804 2164
rect 4908 1664 4964 2164
rect 5068 1664 5124 2164
rect 5228 1664 5284 2164
rect 5632 1664 5688 2164
rect 5792 1664 5848 2164
rect 5952 1664 6008 2164
rect 6112 1664 6168 2164
rect 6272 1664 6328 2164
rect 6432 1664 6488 2164
rect 6592 1664 6648 2164
rect 6752 1664 6808 2164
rect 7040 1664 7096 2164
rect 7444 1664 7500 2164
rect 7604 1664 7660 2164
rect 7764 1664 7820 2164
rect 7924 1664 7980 2164
rect 8084 1664 8140 2164
rect 8244 1664 8300 2164
rect 8404 1664 8460 2164
rect 8564 1664 8620 2164
rect 8852 1664 8908 2164
rect -4724 447 -4668 647
rect -4318 492 -4262 692
rect -4158 492 -4102 692
rect -3998 492 -3942 692
rect -3838 492 -3782 692
rect -3445 481 -2997 569
rect -2659 481 -2211 569
rect -1873 481 -1425 569
rect -1075 447 -1019 647
rect -4724 -47 -4668 153
rect -4318 -92 -4262 108
rect -4158 -92 -4102 108
rect -3998 -92 -3942 108
rect -3838 -92 -3782 108
rect -3445 31 -2997 119
rect -2659 31 -2211 119
rect -1873 31 -1425 119
rect -1075 -47 -1019 153
rect -4318 -1218 -4262 -1018
rect -4158 -1218 -4102 -1018
rect -3998 -1218 -3942 -1018
rect -3838 -1218 -3782 -1018
rect -3445 -1229 -2997 -1141
rect -2659 -1229 -2211 -1141
rect -1873 -1229 -1425 -1141
rect -1075 -1263 -1019 -1063
rect 196 -2052 252 -1552
rect 484 -2052 540 -1552
rect 644 -2052 700 -1552
rect 804 -2052 860 -1552
rect 964 -2052 1020 -1552
rect 1124 -2052 1180 -1552
rect 1284 -2052 1340 -1552
rect 1444 -2052 1500 -1552
rect 1604 -2052 1660 -1552
rect 2008 -2052 2064 -1552
rect 2168 -2052 2224 -1552
rect 2328 -2052 2384 -1552
rect 2488 -2052 2544 -1552
rect 2648 -2052 2704 -1552
rect 2808 -2052 2864 -1552
rect 2968 -2052 3024 -1552
rect 3128 -2052 3184 -1552
rect 3416 -2052 3472 -1552
rect 3820 -2052 3876 -1552
rect 4108 -2052 4164 -1552
rect 4268 -2052 4324 -1552
rect 4428 -2052 4484 -1552
rect 4588 -2052 4644 -1552
rect 4748 -2052 4804 -1552
rect 4908 -2052 4964 -1552
rect 5068 -2052 5124 -1552
rect 5228 -2052 5284 -1552
rect 5632 -2052 5688 -1552
rect 5792 -2052 5848 -1552
rect 5952 -2052 6008 -1552
rect 6112 -2052 6168 -1552
rect 6272 -2052 6328 -1552
rect 6432 -2052 6488 -1552
rect 6592 -2052 6648 -1552
rect 6752 -2052 6808 -1552
rect 7040 -2052 7096 -1552
rect 7444 -2052 7500 -1552
rect 7604 -2052 7660 -1552
rect 7764 -2052 7820 -1552
rect 7924 -2052 7980 -1552
rect 8084 -2052 8140 -1552
rect 8244 -2052 8300 -1552
rect 8404 -2052 8460 -1552
rect 8564 -2052 8620 -1552
rect 8852 -2052 8908 -1552
rect 196 -2688 252 -2188
rect 484 -2688 540 -2188
rect 644 -2688 700 -2188
rect 804 -2688 860 -2188
rect 964 -2688 1020 -2188
rect 1124 -2688 1180 -2188
rect 1284 -2688 1340 -2188
rect 1444 -2688 1500 -2188
rect 1604 -2688 1660 -2188
rect 2008 -2688 2064 -2188
rect 2168 -2688 2224 -2188
rect 2328 -2688 2384 -2188
rect 2488 -2688 2544 -2188
rect 2648 -2688 2704 -2188
rect 2808 -2688 2864 -2188
rect 2968 -2688 3024 -2188
rect 3128 -2688 3184 -2188
rect 3416 -2688 3472 -2188
rect 3820 -2688 3876 -2188
rect 4108 -2688 4164 -2188
rect 4268 -2688 4324 -2188
rect 4428 -2688 4484 -2188
rect 4588 -2688 4644 -2188
rect 4748 -2688 4804 -2188
rect 4908 -2688 4964 -2188
rect 5068 -2688 5124 -2188
rect 5228 -2688 5284 -2188
rect 5632 -2688 5688 -2188
rect 5792 -2688 5848 -2188
rect 5952 -2688 6008 -2188
rect 6112 -2688 6168 -2188
rect 6272 -2688 6328 -2188
rect 6432 -2688 6488 -2188
rect 6592 -2688 6648 -2188
rect 6752 -2688 6808 -2188
rect 7040 -2688 7096 -2188
rect 7444 -2688 7500 -2188
rect 7604 -2688 7660 -2188
rect 7764 -2688 7820 -2188
rect 7924 -2688 7980 -2188
rect 8084 -2688 8140 -2188
rect 8244 -2688 8300 -2188
rect 8404 -2688 8460 -2188
rect 8564 -2688 8620 -2188
rect 8852 -2688 8908 -2188
rect 196 -3324 252 -2824
rect 484 -3324 540 -2824
rect 644 -3324 700 -2824
rect 804 -3324 860 -2824
rect 964 -3324 1020 -2824
rect 1124 -3324 1180 -2824
rect 1284 -3324 1340 -2824
rect 1444 -3324 1500 -2824
rect 1604 -3324 1660 -2824
rect 2008 -3324 2064 -2824
rect 2168 -3324 2224 -2824
rect 2328 -3324 2384 -2824
rect 2488 -3324 2544 -2824
rect 2648 -3324 2704 -2824
rect 2808 -3324 2864 -2824
rect 2968 -3324 3024 -2824
rect 3128 -3324 3184 -2824
rect 3416 -3324 3472 -2824
rect 3820 -3324 3876 -2824
rect 4108 -3324 4164 -2824
rect 4268 -3324 4324 -2824
rect 4428 -3324 4484 -2824
rect 4588 -3324 4644 -2824
rect 4748 -3324 4804 -2824
rect 4908 -3324 4964 -2824
rect 5068 -3324 5124 -2824
rect 5228 -3324 5284 -2824
rect 5632 -3324 5688 -2824
rect 5792 -3324 5848 -2824
rect 5952 -3324 6008 -2824
rect 6112 -3324 6168 -2824
rect 6272 -3324 6328 -2824
rect 6432 -3324 6488 -2824
rect 6592 -3324 6648 -2824
rect 6752 -3324 6808 -2824
rect 7040 -3324 7096 -2824
rect 7444 -3324 7500 -2824
rect 7604 -3324 7660 -2824
rect 7764 -3324 7820 -2824
rect 7924 -3324 7980 -2824
rect 8084 -3324 8140 -2824
rect 8244 -3324 8300 -2824
rect 8404 -3324 8460 -2824
rect 8564 -3324 8620 -2824
rect 8852 -3324 8908 -2824
rect -4001 -4392 -3945 -3892
rect -3713 -4392 -3657 -3892
rect -3553 -4392 -3497 -3892
rect -3393 -4392 -3337 -3892
rect -3233 -4392 -3177 -3892
rect -3073 -4392 -3017 -3892
rect -2913 -4392 -2857 -3892
rect -2753 -4392 -2697 -3892
rect -2593 -4392 -2537 -3892
rect -2189 -4392 -2133 -3892
rect -2029 -4392 -1973 -3892
rect -1869 -4392 -1813 -3892
rect -1709 -4392 -1653 -3892
rect -1549 -4392 -1493 -3892
rect -1389 -4392 -1333 -3892
rect -1229 -4392 -1173 -3892
rect -1069 -4392 -1013 -3892
rect -781 -4392 -725 -3892
rect 196 -4392 252 -3892
rect 484 -4392 540 -3892
rect 644 -4392 700 -3892
rect 804 -4392 860 -3892
rect 964 -4392 1020 -3892
rect 1124 -4392 1180 -3892
rect 1284 -4392 1340 -3892
rect 1444 -4392 1500 -3892
rect 1604 -4392 1660 -3892
rect 2008 -4392 2064 -3892
rect 2168 -4392 2224 -3892
rect 2328 -4392 2384 -3892
rect 2488 -4392 2544 -3892
rect 2648 -4392 2704 -3892
rect 2808 -4392 2864 -3892
rect 2968 -4392 3024 -3892
rect 3128 -4392 3184 -3892
rect 3416 -4392 3472 -3892
rect 3820 -4392 3876 -3892
rect 4108 -4392 4164 -3892
rect 4268 -4392 4324 -3892
rect 4428 -4392 4484 -3892
rect 4588 -4392 4644 -3892
rect 4748 -4392 4804 -3892
rect 4908 -4392 4964 -3892
rect 5068 -4392 5124 -3892
rect 5228 -4392 5284 -3892
rect 5632 -4392 5688 -3892
rect 5792 -4392 5848 -3892
rect 5952 -4392 6008 -3892
rect 6112 -4392 6168 -3892
rect 6272 -4392 6328 -3892
rect 6432 -4392 6488 -3892
rect 6592 -4392 6648 -3892
rect 6752 -4392 6808 -3892
rect 7040 -4392 7096 -3892
rect 7444 -4392 7500 -3892
rect 7604 -4392 7660 -3892
rect 7764 -4392 7820 -3892
rect 7924 -4392 7980 -3892
rect 8084 -4392 8140 -3892
rect 8244 -4392 8300 -3892
rect 8404 -4392 8460 -3892
rect 8564 -4392 8620 -3892
rect 8852 -4392 8908 -3892
rect -4001 -5028 -3945 -4528
rect -3713 -5028 -3657 -4528
rect -3553 -5028 -3497 -4528
rect -3393 -5028 -3337 -4528
rect -3233 -5028 -3177 -4528
rect -3073 -5028 -3017 -4528
rect -2913 -5028 -2857 -4528
rect -2753 -5028 -2697 -4528
rect -2593 -5028 -2537 -4528
rect -2189 -5028 -2133 -4528
rect -2029 -5028 -1973 -4528
rect -1869 -5028 -1813 -4528
rect -1709 -5028 -1653 -4528
rect -1549 -5028 -1493 -4528
rect -1389 -5028 -1333 -4528
rect -1229 -5028 -1173 -4528
rect -1069 -5028 -1013 -4528
rect -781 -5028 -725 -4528
rect 196 -5028 252 -4528
rect 484 -5028 540 -4528
rect 644 -5028 700 -4528
rect 804 -5028 860 -4528
rect 964 -5028 1020 -4528
rect 1124 -5028 1180 -4528
rect 1284 -5028 1340 -4528
rect 1444 -5028 1500 -4528
rect 1604 -5028 1660 -4528
rect 2008 -5028 2064 -4528
rect 2168 -5028 2224 -4528
rect 2328 -5028 2384 -4528
rect 2488 -5028 2544 -4528
rect 2648 -5028 2704 -4528
rect 2808 -5028 2864 -4528
rect 2968 -5028 3024 -4528
rect 3128 -5028 3184 -4528
rect 3416 -5028 3472 -4528
rect 3820 -5028 3876 -4528
rect 4108 -5028 4164 -4528
rect 4268 -5028 4324 -4528
rect 4428 -5028 4484 -4528
rect 4588 -5028 4644 -4528
rect 4748 -5028 4804 -4528
rect 4908 -5028 4964 -4528
rect 5068 -5028 5124 -4528
rect 5228 -5028 5284 -4528
rect 5632 -5028 5688 -4528
rect 5792 -5028 5848 -4528
rect 5952 -5028 6008 -4528
rect 6112 -5028 6168 -4528
rect 6272 -5028 6328 -4528
rect 6432 -5028 6488 -4528
rect 6592 -5028 6648 -4528
rect 6752 -5028 6808 -4528
rect 7040 -5028 7096 -4528
rect 7444 -5028 7500 -4528
rect 7604 -5028 7660 -4528
rect 7764 -5028 7820 -4528
rect 7924 -5028 7980 -4528
rect 8084 -5028 8140 -4528
rect 8244 -5028 8300 -4528
rect 8404 -5028 8460 -4528
rect 8564 -5028 8620 -4528
rect 8852 -5028 8908 -4528
rect -4001 -5664 -3945 -5164
rect -3713 -5664 -3657 -5164
rect -3553 -5664 -3497 -5164
rect -3393 -5664 -3337 -5164
rect -3233 -5664 -3177 -5164
rect -3073 -5664 -3017 -5164
rect -2913 -5664 -2857 -5164
rect -2753 -5664 -2697 -5164
rect -2593 -5664 -2537 -5164
rect -2189 -5664 -2133 -5164
rect -2029 -5664 -1973 -5164
rect -1869 -5664 -1813 -5164
rect -1709 -5664 -1653 -5164
rect -1549 -5664 -1493 -5164
rect -1389 -5664 -1333 -5164
rect -1229 -5664 -1173 -5164
rect -1069 -5664 -1013 -5164
rect -781 -5664 -725 -5164
rect 196 -5664 252 -5164
rect 484 -5664 540 -5164
rect 644 -5664 700 -5164
rect 804 -5664 860 -5164
rect 964 -5664 1020 -5164
rect 1124 -5664 1180 -5164
rect 1284 -5664 1340 -5164
rect 1444 -5664 1500 -5164
rect 1604 -5664 1660 -5164
rect 2008 -5664 2064 -5164
rect 2168 -5664 2224 -5164
rect 2328 -5664 2384 -5164
rect 2488 -5664 2544 -5164
rect 2648 -5664 2704 -5164
rect 2808 -5664 2864 -5164
rect 2968 -5664 3024 -5164
rect 3128 -5664 3184 -5164
rect 3416 -5664 3472 -5164
rect 3820 -5664 3876 -5164
rect 4108 -5664 4164 -5164
rect 4268 -5664 4324 -5164
rect 4428 -5664 4484 -5164
rect 4588 -5664 4644 -5164
rect 4748 -5664 4804 -5164
rect 4908 -5664 4964 -5164
rect 5068 -5664 5124 -5164
rect 5228 -5664 5284 -5164
rect 5632 -5664 5688 -5164
rect 5792 -5664 5848 -5164
rect 5952 -5664 6008 -5164
rect 6112 -5664 6168 -5164
rect 6272 -5664 6328 -5164
rect 6432 -5664 6488 -5164
rect 6592 -5664 6648 -5164
rect 6752 -5664 6808 -5164
rect 7040 -5664 7096 -5164
rect 7444 -5664 7500 -5164
rect 7604 -5664 7660 -5164
rect 7764 -5664 7820 -5164
rect 7924 -5664 7980 -5164
rect 8084 -5664 8140 -5164
rect 8244 -5664 8300 -5164
rect 8404 -5664 8460 -5164
rect 8564 -5664 8620 -5164
rect 8852 -5664 8908 -5164
<< ndiff >>
rect 108 7087 196 7100
rect 108 6863 121 7087
rect 167 6863 196 7087
rect 108 6850 196 6863
rect 252 7087 356 7100
rect 252 6863 281 7087
rect 327 6863 356 7087
rect 252 6850 356 6863
rect 412 7087 516 7100
rect 412 6863 441 7087
rect 487 6863 516 7087
rect 412 6850 516 6863
rect 572 7087 676 7100
rect 572 6863 601 7087
rect 647 6863 676 7087
rect 572 6850 676 6863
rect 732 7087 836 7100
rect 732 6863 761 7087
rect 807 6863 836 7087
rect 732 6850 836 6863
rect 892 7087 996 7100
rect 892 6863 921 7087
rect 967 6863 996 7087
rect 892 6850 996 6863
rect 1052 7087 1156 7100
rect 1052 6863 1081 7087
rect 1127 6863 1156 7087
rect 1052 6850 1156 6863
rect 1212 7087 1316 7100
rect 1212 6863 1241 7087
rect 1287 6863 1316 7087
rect 1212 6850 1316 6863
rect 1372 7087 1460 7100
rect 1372 6863 1401 7087
rect 1447 6863 1460 7087
rect 1372 6850 1460 6863
rect 1516 7087 1604 7100
rect 1516 6863 1529 7087
rect 1575 6863 1604 7087
rect 1516 6850 1604 6863
rect 1660 7087 1748 7100
rect 1660 6863 1689 7087
rect 1735 6863 1748 7087
rect 1660 6850 1748 6863
rect 1920 7087 2008 7100
rect 1920 6863 1933 7087
rect 1979 6863 2008 7087
rect 1920 6850 2008 6863
rect 2064 7087 2152 7100
rect 2064 6863 2093 7087
rect 2139 6863 2152 7087
rect 2064 6850 2152 6863
rect 2208 7087 2296 7100
rect 2208 6863 2221 7087
rect 2267 6863 2296 7087
rect 2208 6850 2296 6863
rect 2352 7087 2456 7100
rect 2352 6863 2381 7087
rect 2427 6863 2456 7087
rect 2352 6850 2456 6863
rect 2512 7087 2616 7100
rect 2512 6863 2541 7087
rect 2587 6863 2616 7087
rect 2512 6850 2616 6863
rect 2672 7087 2776 7100
rect 2672 6863 2701 7087
rect 2747 6863 2776 7087
rect 2672 6850 2776 6863
rect 2832 7087 2936 7100
rect 2832 6863 2861 7087
rect 2907 6863 2936 7087
rect 2832 6850 2936 6863
rect 2992 7087 3096 7100
rect 2992 6863 3021 7087
rect 3067 6863 3096 7087
rect 2992 6850 3096 6863
rect 3152 7087 3256 7100
rect 3152 6863 3181 7087
rect 3227 6863 3256 7087
rect 3152 6850 3256 6863
rect 3312 7087 3416 7100
rect 3312 6863 3341 7087
rect 3387 6863 3416 7087
rect 3312 6850 3416 6863
rect 3472 7087 3560 7100
rect 3472 6863 3501 7087
rect 3547 6863 3560 7087
rect 3472 6850 3560 6863
rect 3732 7087 3820 7100
rect 3732 6863 3745 7087
rect 3791 6863 3820 7087
rect 3732 6850 3820 6863
rect 3876 7087 3964 7100
rect 3876 6863 3905 7087
rect 3951 6863 3964 7087
rect 3876 6850 3964 6863
rect 4020 7087 4108 7100
rect 4020 6863 4033 7087
rect 4079 6863 4108 7087
rect 4020 6850 4108 6863
rect 4164 7087 4268 7100
rect 4164 6863 4193 7087
rect 4239 6863 4268 7087
rect 4164 6850 4268 6863
rect 4324 7087 4428 7100
rect 4324 6863 4353 7087
rect 4399 6863 4428 7087
rect 4324 6850 4428 6863
rect 4484 7087 4588 7100
rect 4484 6863 4513 7087
rect 4559 6863 4588 7087
rect 4484 6850 4588 6863
rect 4644 7087 4748 7100
rect 4644 6863 4673 7087
rect 4719 6863 4748 7087
rect 4644 6850 4748 6863
rect 4804 7087 4908 7100
rect 4804 6863 4833 7087
rect 4879 6863 4908 7087
rect 4804 6850 4908 6863
rect 4964 7087 5068 7100
rect 4964 6863 4993 7087
rect 5039 6863 5068 7087
rect 4964 6850 5068 6863
rect 5124 7087 5228 7100
rect 5124 6863 5153 7087
rect 5199 6863 5228 7087
rect 5124 6850 5228 6863
rect 5284 7087 5372 7100
rect 5284 6863 5313 7087
rect 5359 6863 5372 7087
rect 5284 6850 5372 6863
rect 5544 7087 5632 7100
rect 5544 6863 5557 7087
rect 5603 6863 5632 7087
rect 5544 6850 5632 6863
rect 5688 7087 5776 7100
rect 5688 6863 5717 7087
rect 5763 6863 5776 7087
rect 5688 6850 5776 6863
rect 5832 7087 5920 7100
rect 5832 6863 5845 7087
rect 5891 6863 5920 7087
rect 5832 6850 5920 6863
rect 5976 7087 6080 7100
rect 5976 6863 6005 7087
rect 6051 6863 6080 7087
rect 5976 6850 6080 6863
rect 6136 7087 6240 7100
rect 6136 6863 6165 7087
rect 6211 6863 6240 7087
rect 6136 6850 6240 6863
rect 6296 7087 6400 7100
rect 6296 6863 6325 7087
rect 6371 6863 6400 7087
rect 6296 6850 6400 6863
rect 6456 7087 6560 7100
rect 6456 6863 6485 7087
rect 6531 6863 6560 7087
rect 6456 6850 6560 6863
rect 6616 7087 6720 7100
rect 6616 6863 6645 7087
rect 6691 6863 6720 7087
rect 6616 6850 6720 6863
rect 6776 7087 6880 7100
rect 6776 6863 6805 7087
rect 6851 6863 6880 7087
rect 6776 6850 6880 6863
rect 6936 7087 7040 7100
rect 6936 6863 6965 7087
rect 7011 6863 7040 7087
rect 6936 6850 7040 6863
rect 7096 7087 7184 7100
rect 7096 6863 7125 7087
rect 7171 6863 7184 7087
rect 7096 6850 7184 6863
rect 7356 7087 7444 7100
rect 7356 6863 7369 7087
rect 7415 6863 7444 7087
rect 7356 6850 7444 6863
rect 7500 7087 7588 7100
rect 7500 6863 7529 7087
rect 7575 6863 7588 7087
rect 7500 6850 7588 6863
rect 7644 7087 7732 7100
rect 7644 6863 7657 7087
rect 7703 6863 7732 7087
rect 7644 6850 7732 6863
rect 7788 7087 7892 7100
rect 7788 6863 7817 7087
rect 7863 6863 7892 7087
rect 7788 6850 7892 6863
rect 7948 7087 8052 7100
rect 7948 6863 7977 7087
rect 8023 6863 8052 7087
rect 7948 6850 8052 6863
rect 8108 7087 8212 7100
rect 8108 6863 8137 7087
rect 8183 6863 8212 7087
rect 8108 6850 8212 6863
rect 8268 7087 8372 7100
rect 8268 6863 8297 7087
rect 8343 6863 8372 7087
rect 8268 6850 8372 6863
rect 8428 7087 8532 7100
rect 8428 6863 8457 7087
rect 8503 6863 8532 7087
rect 8428 6850 8532 6863
rect 8588 7087 8692 7100
rect 8588 6863 8617 7087
rect 8663 6863 8692 7087
rect 8588 6850 8692 6863
rect 8748 7087 8852 7100
rect 8748 6863 8777 7087
rect 8823 6863 8852 7087
rect 8748 6850 8852 6863
rect 8908 7087 8996 7100
rect 8908 6863 8937 7087
rect 8983 6863 8996 7087
rect 8908 6850 8996 6863
rect 108 6701 196 6714
rect 108 6477 121 6701
rect 167 6477 196 6701
rect 108 6464 196 6477
rect 252 6701 356 6714
rect 252 6477 281 6701
rect 327 6477 356 6701
rect 252 6464 356 6477
rect 412 6701 516 6714
rect 412 6477 441 6701
rect 487 6477 516 6701
rect 412 6464 516 6477
rect 572 6701 676 6714
rect 572 6477 601 6701
rect 647 6477 676 6701
rect 572 6464 676 6477
rect 732 6701 836 6714
rect 732 6477 761 6701
rect 807 6477 836 6701
rect 732 6464 836 6477
rect 892 6701 996 6714
rect 892 6477 921 6701
rect 967 6477 996 6701
rect 892 6464 996 6477
rect 1052 6701 1156 6714
rect 1052 6477 1081 6701
rect 1127 6477 1156 6701
rect 1052 6464 1156 6477
rect 1212 6701 1316 6714
rect 1212 6477 1241 6701
rect 1287 6477 1316 6701
rect 1212 6464 1316 6477
rect 1372 6701 1460 6714
rect 1372 6477 1401 6701
rect 1447 6477 1460 6701
rect 1372 6464 1460 6477
rect 1516 6701 1604 6714
rect 1516 6477 1529 6701
rect 1575 6477 1604 6701
rect 1516 6464 1604 6477
rect 1660 6701 1748 6714
rect 1660 6477 1689 6701
rect 1735 6477 1748 6701
rect 1660 6464 1748 6477
rect 1920 6701 2008 6714
rect 1920 6477 1933 6701
rect 1979 6477 2008 6701
rect 1920 6464 2008 6477
rect 2064 6701 2152 6714
rect 2064 6477 2093 6701
rect 2139 6477 2152 6701
rect 2064 6464 2152 6477
rect 2208 6701 2296 6714
rect 2208 6477 2221 6701
rect 2267 6477 2296 6701
rect 2208 6464 2296 6477
rect 2352 6701 2456 6714
rect 2352 6477 2381 6701
rect 2427 6477 2456 6701
rect 2352 6464 2456 6477
rect 2512 6701 2616 6714
rect 2512 6477 2541 6701
rect 2587 6477 2616 6701
rect 2512 6464 2616 6477
rect 2672 6701 2776 6714
rect 2672 6477 2701 6701
rect 2747 6477 2776 6701
rect 2672 6464 2776 6477
rect 2832 6701 2936 6714
rect 2832 6477 2861 6701
rect 2907 6477 2936 6701
rect 2832 6464 2936 6477
rect 2992 6701 3096 6714
rect 2992 6477 3021 6701
rect 3067 6477 3096 6701
rect 2992 6464 3096 6477
rect 3152 6701 3256 6714
rect 3152 6477 3181 6701
rect 3227 6477 3256 6701
rect 3152 6464 3256 6477
rect 3312 6701 3416 6714
rect 3312 6477 3341 6701
rect 3387 6477 3416 6701
rect 3312 6464 3416 6477
rect 3472 6701 3560 6714
rect 3472 6477 3501 6701
rect 3547 6477 3560 6701
rect 3472 6464 3560 6477
rect 3732 6701 3820 6714
rect 3732 6477 3745 6701
rect 3791 6477 3820 6701
rect 3732 6464 3820 6477
rect 3876 6701 3964 6714
rect 3876 6477 3905 6701
rect 3951 6477 3964 6701
rect 3876 6464 3964 6477
rect 4020 6701 4108 6714
rect 4020 6477 4033 6701
rect 4079 6477 4108 6701
rect 4020 6464 4108 6477
rect 4164 6701 4268 6714
rect 4164 6477 4193 6701
rect 4239 6477 4268 6701
rect 4164 6464 4268 6477
rect 4324 6701 4428 6714
rect 4324 6477 4353 6701
rect 4399 6477 4428 6701
rect 4324 6464 4428 6477
rect 4484 6701 4588 6714
rect 4484 6477 4513 6701
rect 4559 6477 4588 6701
rect 4484 6464 4588 6477
rect 4644 6701 4748 6714
rect 4644 6477 4673 6701
rect 4719 6477 4748 6701
rect 4644 6464 4748 6477
rect 4804 6701 4908 6714
rect 4804 6477 4833 6701
rect 4879 6477 4908 6701
rect 4804 6464 4908 6477
rect 4964 6701 5068 6714
rect 4964 6477 4993 6701
rect 5039 6477 5068 6701
rect 4964 6464 5068 6477
rect 5124 6701 5228 6714
rect 5124 6477 5153 6701
rect 5199 6477 5228 6701
rect 5124 6464 5228 6477
rect 5284 6701 5372 6714
rect 5284 6477 5313 6701
rect 5359 6477 5372 6701
rect 5284 6464 5372 6477
rect 5544 6701 5632 6714
rect 5544 6477 5557 6701
rect 5603 6477 5632 6701
rect 5544 6464 5632 6477
rect 5688 6701 5776 6714
rect 5688 6477 5717 6701
rect 5763 6477 5776 6701
rect 5688 6464 5776 6477
rect 5832 6701 5920 6714
rect 5832 6477 5845 6701
rect 5891 6477 5920 6701
rect 5832 6464 5920 6477
rect 5976 6701 6080 6714
rect 5976 6477 6005 6701
rect 6051 6477 6080 6701
rect 5976 6464 6080 6477
rect 6136 6701 6240 6714
rect 6136 6477 6165 6701
rect 6211 6477 6240 6701
rect 6136 6464 6240 6477
rect 6296 6701 6400 6714
rect 6296 6477 6325 6701
rect 6371 6477 6400 6701
rect 6296 6464 6400 6477
rect 6456 6701 6560 6714
rect 6456 6477 6485 6701
rect 6531 6477 6560 6701
rect 6456 6464 6560 6477
rect 6616 6701 6720 6714
rect 6616 6477 6645 6701
rect 6691 6477 6720 6701
rect 6616 6464 6720 6477
rect 6776 6701 6880 6714
rect 6776 6477 6805 6701
rect 6851 6477 6880 6701
rect 6776 6464 6880 6477
rect 6936 6701 7040 6714
rect 6936 6477 6965 6701
rect 7011 6477 7040 6701
rect 6936 6464 7040 6477
rect 7096 6701 7184 6714
rect 7096 6477 7125 6701
rect 7171 6477 7184 6701
rect 7096 6464 7184 6477
rect 7356 6701 7444 6714
rect 7356 6477 7369 6701
rect 7415 6477 7444 6701
rect 7356 6464 7444 6477
rect 7500 6701 7588 6714
rect 7500 6477 7529 6701
rect 7575 6477 7588 6701
rect 7500 6464 7588 6477
rect 7644 6701 7732 6714
rect 7644 6477 7657 6701
rect 7703 6477 7732 6701
rect 7644 6464 7732 6477
rect 7788 6701 7892 6714
rect 7788 6477 7817 6701
rect 7863 6477 7892 6701
rect 7788 6464 7892 6477
rect 7948 6701 8052 6714
rect 7948 6477 7977 6701
rect 8023 6477 8052 6701
rect 7948 6464 8052 6477
rect 8108 6701 8212 6714
rect 8108 6477 8137 6701
rect 8183 6477 8212 6701
rect 8108 6464 8212 6477
rect 8268 6701 8372 6714
rect 8268 6477 8297 6701
rect 8343 6477 8372 6701
rect 8268 6464 8372 6477
rect 8428 6701 8532 6714
rect 8428 6477 8457 6701
rect 8503 6477 8532 6701
rect 8428 6464 8532 6477
rect 8588 6701 8692 6714
rect 8588 6477 8617 6701
rect 8663 6477 8692 6701
rect 8588 6464 8692 6477
rect 8748 6701 8852 6714
rect 8748 6477 8777 6701
rect 8823 6477 8852 6701
rect 8748 6464 8852 6477
rect 8908 6701 8996 6714
rect 8908 6477 8937 6701
rect 8983 6477 8996 6701
rect 8908 6464 8996 6477
rect 108 6315 196 6328
rect 108 6091 121 6315
rect 167 6091 196 6315
rect 108 6078 196 6091
rect 252 6315 356 6328
rect 252 6091 281 6315
rect 327 6091 356 6315
rect 252 6078 356 6091
rect 412 6315 516 6328
rect 412 6091 441 6315
rect 487 6091 516 6315
rect 412 6078 516 6091
rect 572 6315 676 6328
rect 572 6091 601 6315
rect 647 6091 676 6315
rect 572 6078 676 6091
rect 732 6315 836 6328
rect 732 6091 761 6315
rect 807 6091 836 6315
rect 732 6078 836 6091
rect 892 6315 996 6328
rect 892 6091 921 6315
rect 967 6091 996 6315
rect 892 6078 996 6091
rect 1052 6315 1156 6328
rect 1052 6091 1081 6315
rect 1127 6091 1156 6315
rect 1052 6078 1156 6091
rect 1212 6315 1316 6328
rect 1212 6091 1241 6315
rect 1287 6091 1316 6315
rect 1212 6078 1316 6091
rect 1372 6315 1460 6328
rect 1372 6091 1401 6315
rect 1447 6091 1460 6315
rect 1372 6078 1460 6091
rect 1516 6315 1604 6328
rect 1516 6091 1529 6315
rect 1575 6091 1604 6315
rect 1516 6078 1604 6091
rect 1660 6315 1748 6328
rect 1660 6091 1689 6315
rect 1735 6091 1748 6315
rect 1660 6078 1748 6091
rect 1920 6315 2008 6328
rect 1920 6091 1933 6315
rect 1979 6091 2008 6315
rect 1920 6078 2008 6091
rect 2064 6315 2152 6328
rect 2064 6091 2093 6315
rect 2139 6091 2152 6315
rect 2064 6078 2152 6091
rect 2208 6315 2296 6328
rect 2208 6091 2221 6315
rect 2267 6091 2296 6315
rect 2208 6078 2296 6091
rect 2352 6315 2456 6328
rect 2352 6091 2381 6315
rect 2427 6091 2456 6315
rect 2352 6078 2456 6091
rect 2512 6315 2616 6328
rect 2512 6091 2541 6315
rect 2587 6091 2616 6315
rect 2512 6078 2616 6091
rect 2672 6315 2776 6328
rect 2672 6091 2701 6315
rect 2747 6091 2776 6315
rect 2672 6078 2776 6091
rect 2832 6315 2936 6328
rect 2832 6091 2861 6315
rect 2907 6091 2936 6315
rect 2832 6078 2936 6091
rect 2992 6315 3096 6328
rect 2992 6091 3021 6315
rect 3067 6091 3096 6315
rect 2992 6078 3096 6091
rect 3152 6315 3256 6328
rect 3152 6091 3181 6315
rect 3227 6091 3256 6315
rect 3152 6078 3256 6091
rect 3312 6315 3416 6328
rect 3312 6091 3341 6315
rect 3387 6091 3416 6315
rect 3312 6078 3416 6091
rect 3472 6315 3560 6328
rect 3472 6091 3501 6315
rect 3547 6091 3560 6315
rect 3472 6078 3560 6091
rect 3732 6315 3820 6328
rect 3732 6091 3745 6315
rect 3791 6091 3820 6315
rect 3732 6078 3820 6091
rect 3876 6315 3964 6328
rect 3876 6091 3905 6315
rect 3951 6091 3964 6315
rect 3876 6078 3964 6091
rect 4020 6315 4108 6328
rect 4020 6091 4033 6315
rect 4079 6091 4108 6315
rect 4020 6078 4108 6091
rect 4164 6315 4268 6328
rect 4164 6091 4193 6315
rect 4239 6091 4268 6315
rect 4164 6078 4268 6091
rect 4324 6315 4428 6328
rect 4324 6091 4353 6315
rect 4399 6091 4428 6315
rect 4324 6078 4428 6091
rect 4484 6315 4588 6328
rect 4484 6091 4513 6315
rect 4559 6091 4588 6315
rect 4484 6078 4588 6091
rect 4644 6315 4748 6328
rect 4644 6091 4673 6315
rect 4719 6091 4748 6315
rect 4644 6078 4748 6091
rect 4804 6315 4908 6328
rect 4804 6091 4833 6315
rect 4879 6091 4908 6315
rect 4804 6078 4908 6091
rect 4964 6315 5068 6328
rect 4964 6091 4993 6315
rect 5039 6091 5068 6315
rect 4964 6078 5068 6091
rect 5124 6315 5228 6328
rect 5124 6091 5153 6315
rect 5199 6091 5228 6315
rect 5124 6078 5228 6091
rect 5284 6315 5372 6328
rect 5284 6091 5313 6315
rect 5359 6091 5372 6315
rect 5284 6078 5372 6091
rect 5544 6315 5632 6328
rect 5544 6091 5557 6315
rect 5603 6091 5632 6315
rect 5544 6078 5632 6091
rect 5688 6315 5776 6328
rect 5688 6091 5717 6315
rect 5763 6091 5776 6315
rect 5688 6078 5776 6091
rect 5832 6315 5920 6328
rect 5832 6091 5845 6315
rect 5891 6091 5920 6315
rect 5832 6078 5920 6091
rect 5976 6315 6080 6328
rect 5976 6091 6005 6315
rect 6051 6091 6080 6315
rect 5976 6078 6080 6091
rect 6136 6315 6240 6328
rect 6136 6091 6165 6315
rect 6211 6091 6240 6315
rect 6136 6078 6240 6091
rect 6296 6315 6400 6328
rect 6296 6091 6325 6315
rect 6371 6091 6400 6315
rect 6296 6078 6400 6091
rect 6456 6315 6560 6328
rect 6456 6091 6485 6315
rect 6531 6091 6560 6315
rect 6456 6078 6560 6091
rect 6616 6315 6720 6328
rect 6616 6091 6645 6315
rect 6691 6091 6720 6315
rect 6616 6078 6720 6091
rect 6776 6315 6880 6328
rect 6776 6091 6805 6315
rect 6851 6091 6880 6315
rect 6776 6078 6880 6091
rect 6936 6315 7040 6328
rect 6936 6091 6965 6315
rect 7011 6091 7040 6315
rect 6936 6078 7040 6091
rect 7096 6315 7184 6328
rect 7096 6091 7125 6315
rect 7171 6091 7184 6315
rect 7096 6078 7184 6091
rect 7356 6315 7444 6328
rect 7356 6091 7369 6315
rect 7415 6091 7444 6315
rect 7356 6078 7444 6091
rect 7500 6315 7588 6328
rect 7500 6091 7529 6315
rect 7575 6091 7588 6315
rect 7500 6078 7588 6091
rect 7644 6315 7732 6328
rect 7644 6091 7657 6315
rect 7703 6091 7732 6315
rect 7644 6078 7732 6091
rect 7788 6315 7892 6328
rect 7788 6091 7817 6315
rect 7863 6091 7892 6315
rect 7788 6078 7892 6091
rect 7948 6315 8052 6328
rect 7948 6091 7977 6315
rect 8023 6091 8052 6315
rect 7948 6078 8052 6091
rect 8108 6315 8212 6328
rect 8108 6091 8137 6315
rect 8183 6091 8212 6315
rect 8108 6078 8212 6091
rect 8268 6315 8372 6328
rect 8268 6091 8297 6315
rect 8343 6091 8372 6315
rect 8268 6078 8372 6091
rect 8428 6315 8532 6328
rect 8428 6091 8457 6315
rect 8503 6091 8532 6315
rect 8428 6078 8532 6091
rect 8588 6315 8692 6328
rect 8588 6091 8617 6315
rect 8663 6091 8692 6315
rect 8588 6078 8692 6091
rect 8748 6315 8852 6328
rect 8748 6091 8777 6315
rect 8823 6091 8852 6315
rect 8748 6078 8852 6091
rect 8908 6315 8996 6328
rect 8908 6091 8937 6315
rect 8983 6091 8996 6315
rect 8908 6078 8996 6091
rect -4812 3088 -4724 3101
rect -4812 3014 -4799 3088
rect -4753 3014 -4724 3088
rect -4812 3001 -4724 3014
rect -4668 3088 -4580 3101
rect -4668 3014 -4639 3088
rect -4593 3014 -4580 3088
rect -4668 3001 -4580 3014
rect -4246 3076 -4158 3089
rect -4246 3002 -4233 3076
rect -4187 3002 -4158 3076
rect -4246 2989 -4158 3002
rect -4102 3076 -3998 3089
rect -4102 3002 -4073 3076
rect -4027 3002 -3998 3076
rect -4102 2989 -3998 3002
rect -3942 3076 -3854 3089
rect -1163 3088 -1075 3101
rect -3942 3002 -3913 3076
rect -3867 3002 -3854 3076
rect -3942 2989 -3854 3002
rect -3541 3036 -3469 3049
rect -3541 2990 -3528 3036
rect -3482 3035 -3469 3036
rect -2981 3036 -2909 3049
rect -2981 3035 -2968 3036
rect -3482 2991 -3449 3035
rect -3001 2991 -2968 3035
rect -3482 2990 -3469 2991
rect -3541 2977 -3469 2990
rect -2981 2990 -2968 2991
rect -2922 2990 -2909 3036
rect -2981 2977 -2909 2990
rect -2755 3036 -2683 3049
rect -2755 2990 -2742 3036
rect -2696 3035 -2683 3036
rect -2195 3036 -2123 3049
rect -2195 3035 -2182 3036
rect -2696 2991 -2663 3035
rect -2215 2991 -2182 3035
rect -2696 2990 -2683 2991
rect -2755 2977 -2683 2990
rect -2195 2990 -2182 2991
rect -2136 2990 -2123 3036
rect -2195 2977 -2123 2990
rect -1969 3036 -1897 3049
rect -1969 2990 -1956 3036
rect -1910 3035 -1897 3036
rect -1409 3036 -1337 3049
rect -1409 3035 -1396 3036
rect -1910 2991 -1877 3035
rect -1429 2991 -1396 3035
rect -1910 2990 -1897 2991
rect -1969 2977 -1897 2990
rect -1409 2990 -1396 2991
rect -1350 2990 -1337 3036
rect -1163 3014 -1150 3088
rect -1104 3014 -1075 3088
rect -1163 3001 -1075 3014
rect -1019 3088 -931 3101
rect -1019 3014 -990 3088
rect -944 3014 -931 3088
rect -1019 3001 -931 3014
rect -1409 2977 -1337 2990
rect -4246 2728 -4158 2741
rect -4246 2654 -4233 2728
rect -4187 2654 -4158 2728
rect -4246 2641 -4158 2654
rect -4102 2728 -3998 2741
rect -4102 2654 -4073 2728
rect -4027 2654 -3998 2728
rect -4102 2641 -3998 2654
rect -3942 2728 -3854 2741
rect -3942 2654 -3913 2728
rect -3867 2654 -3854 2728
rect -3541 2740 -3469 2753
rect -3541 2694 -3528 2740
rect -3482 2739 -3469 2740
rect -2981 2740 -2909 2753
rect -2981 2739 -2968 2740
rect -3482 2695 -3449 2739
rect -3001 2695 -2968 2739
rect -3482 2694 -3469 2695
rect -3541 2681 -3469 2694
rect -3942 2641 -3854 2654
rect -2981 2694 -2968 2695
rect -2922 2694 -2909 2740
rect -2981 2681 -2909 2694
rect -2755 2740 -2683 2753
rect -2755 2694 -2742 2740
rect -2696 2739 -2683 2740
rect -2195 2740 -2123 2753
rect -2195 2739 -2182 2740
rect -2696 2695 -2663 2739
rect -2215 2695 -2182 2739
rect -2696 2694 -2683 2695
rect -2755 2681 -2683 2694
rect -2195 2694 -2182 2695
rect -2136 2694 -2123 2740
rect -2195 2681 -2123 2694
rect -1969 2740 -1897 2753
rect -1969 2694 -1956 2740
rect -1910 2739 -1897 2740
rect -1409 2740 -1337 2753
rect -1409 2739 -1396 2740
rect -1910 2695 -1877 2739
rect -1429 2695 -1396 2739
rect -1910 2694 -1897 2695
rect -1969 2681 -1897 2694
rect -1409 2694 -1396 2695
rect -1350 2694 -1337 2740
rect -1409 2681 -1337 2694
rect -1163 2716 -1075 2729
rect -1163 2642 -1150 2716
rect -1104 2642 -1075 2716
rect -1163 2629 -1075 2642
rect -1019 2716 -931 2729
rect -1019 2642 -990 2716
rect -944 2642 -931 2716
rect -1019 2629 -931 2642
rect -4246 1366 -4158 1379
rect -4246 1292 -4233 1366
rect -4187 1292 -4158 1366
rect -4246 1279 -4158 1292
rect -4102 1366 -3998 1379
rect -4102 1292 -4073 1366
rect -4027 1292 -3998 1366
rect -4102 1279 -3998 1292
rect -3942 1366 -3854 1379
rect -1163 1378 -1075 1391
rect -3942 1292 -3913 1366
rect -3867 1292 -3854 1366
rect -3942 1279 -3854 1292
rect -3541 1326 -3469 1339
rect -3541 1280 -3528 1326
rect -3482 1325 -3469 1326
rect -2981 1326 -2909 1339
rect -2981 1325 -2968 1326
rect -3482 1281 -3449 1325
rect -3001 1281 -2968 1325
rect -3482 1280 -3469 1281
rect -3541 1267 -3469 1280
rect -2981 1280 -2968 1281
rect -2922 1280 -2909 1326
rect -2981 1267 -2909 1280
rect -2755 1326 -2683 1339
rect -2755 1280 -2742 1326
rect -2696 1325 -2683 1326
rect -2195 1326 -2123 1339
rect -2195 1325 -2182 1326
rect -2696 1281 -2663 1325
rect -2215 1281 -2182 1325
rect -2696 1280 -2683 1281
rect -2755 1267 -2683 1280
rect -2195 1280 -2182 1281
rect -2136 1280 -2123 1326
rect -2195 1267 -2123 1280
rect -1969 1326 -1897 1339
rect -1969 1280 -1956 1326
rect -1910 1325 -1897 1326
rect -1409 1326 -1337 1339
rect -1409 1325 -1396 1326
rect -1910 1281 -1877 1325
rect -1429 1281 -1396 1325
rect -1910 1280 -1897 1281
rect -1969 1267 -1897 1280
rect -1409 1280 -1396 1281
rect -1350 1280 -1337 1326
rect -1163 1304 -1150 1378
rect -1104 1304 -1075 1378
rect -1163 1291 -1075 1304
rect -1019 1378 -931 1391
rect -1019 1304 -990 1378
rect -944 1304 -931 1378
rect -1019 1291 -931 1304
rect 108 1349 196 1362
rect -1409 1267 -1337 1280
rect 108 1125 121 1349
rect 167 1125 196 1349
rect 108 1112 196 1125
rect 252 1349 340 1362
rect 252 1125 281 1349
rect 327 1125 340 1349
rect 252 1112 340 1125
rect 396 1349 484 1362
rect 396 1125 409 1349
rect 455 1125 484 1349
rect 396 1112 484 1125
rect 540 1349 644 1362
rect 540 1125 569 1349
rect 615 1125 644 1349
rect 540 1112 644 1125
rect 700 1349 804 1362
rect 700 1125 729 1349
rect 775 1125 804 1349
rect 700 1112 804 1125
rect 860 1349 964 1362
rect 860 1125 889 1349
rect 935 1125 964 1349
rect 860 1112 964 1125
rect 1020 1349 1124 1362
rect 1020 1125 1049 1349
rect 1095 1125 1124 1349
rect 1020 1112 1124 1125
rect 1180 1349 1284 1362
rect 1180 1125 1209 1349
rect 1255 1125 1284 1349
rect 1180 1112 1284 1125
rect 1340 1349 1444 1362
rect 1340 1125 1369 1349
rect 1415 1125 1444 1349
rect 1340 1112 1444 1125
rect 1500 1349 1604 1362
rect 1500 1125 1529 1349
rect 1575 1125 1604 1349
rect 1500 1112 1604 1125
rect 1660 1349 1748 1362
rect 1660 1125 1689 1349
rect 1735 1125 1748 1349
rect 1660 1112 1748 1125
rect 1920 1349 2008 1362
rect 1920 1125 1933 1349
rect 1979 1125 2008 1349
rect 1920 1112 2008 1125
rect 2064 1349 2168 1362
rect 2064 1125 2093 1349
rect 2139 1125 2168 1349
rect 2064 1112 2168 1125
rect 2224 1349 2328 1362
rect 2224 1125 2253 1349
rect 2299 1125 2328 1349
rect 2224 1112 2328 1125
rect 2384 1349 2488 1362
rect 2384 1125 2413 1349
rect 2459 1125 2488 1349
rect 2384 1112 2488 1125
rect 2544 1349 2648 1362
rect 2544 1125 2573 1349
rect 2619 1125 2648 1349
rect 2544 1112 2648 1125
rect 2704 1349 2808 1362
rect 2704 1125 2733 1349
rect 2779 1125 2808 1349
rect 2704 1112 2808 1125
rect 2864 1349 2968 1362
rect 2864 1125 2893 1349
rect 2939 1125 2968 1349
rect 2864 1112 2968 1125
rect 3024 1349 3128 1362
rect 3024 1125 3053 1349
rect 3099 1125 3128 1349
rect 3024 1112 3128 1125
rect 3184 1349 3272 1362
rect 3184 1125 3213 1349
rect 3259 1125 3272 1349
rect 3184 1112 3272 1125
rect 3328 1349 3416 1362
rect 3328 1125 3341 1349
rect 3387 1125 3416 1349
rect 3328 1112 3416 1125
rect 3472 1349 3560 1362
rect 3472 1125 3501 1349
rect 3547 1125 3560 1349
rect 3472 1112 3560 1125
rect 3732 1349 3820 1362
rect 3732 1125 3745 1349
rect 3791 1125 3820 1349
rect 3732 1112 3820 1125
rect 3876 1349 3964 1362
rect 3876 1125 3905 1349
rect 3951 1125 3964 1349
rect 3876 1112 3964 1125
rect 4020 1349 4108 1362
rect 4020 1125 4033 1349
rect 4079 1125 4108 1349
rect 4020 1112 4108 1125
rect 4164 1349 4268 1362
rect 4164 1125 4193 1349
rect 4239 1125 4268 1349
rect 4164 1112 4268 1125
rect 4324 1349 4428 1362
rect 4324 1125 4353 1349
rect 4399 1125 4428 1349
rect 4324 1112 4428 1125
rect 4484 1349 4588 1362
rect 4484 1125 4513 1349
rect 4559 1125 4588 1349
rect 4484 1112 4588 1125
rect 4644 1349 4748 1362
rect 4644 1125 4673 1349
rect 4719 1125 4748 1349
rect 4644 1112 4748 1125
rect 4804 1349 4908 1362
rect 4804 1125 4833 1349
rect 4879 1125 4908 1349
rect 4804 1112 4908 1125
rect 4964 1349 5068 1362
rect 4964 1125 4993 1349
rect 5039 1125 5068 1349
rect 4964 1112 5068 1125
rect 5124 1349 5228 1362
rect 5124 1125 5153 1349
rect 5199 1125 5228 1349
rect 5124 1112 5228 1125
rect 5284 1349 5372 1362
rect 5284 1125 5313 1349
rect 5359 1125 5372 1349
rect 5284 1112 5372 1125
rect 5544 1349 5632 1362
rect 5544 1125 5557 1349
rect 5603 1125 5632 1349
rect 5544 1112 5632 1125
rect 5688 1349 5792 1362
rect 5688 1125 5717 1349
rect 5763 1125 5792 1349
rect 5688 1112 5792 1125
rect 5848 1349 5952 1362
rect 5848 1125 5877 1349
rect 5923 1125 5952 1349
rect 5848 1112 5952 1125
rect 6008 1349 6112 1362
rect 6008 1125 6037 1349
rect 6083 1125 6112 1349
rect 6008 1112 6112 1125
rect 6168 1349 6272 1362
rect 6168 1125 6197 1349
rect 6243 1125 6272 1349
rect 6168 1112 6272 1125
rect 6328 1349 6432 1362
rect 6328 1125 6357 1349
rect 6403 1125 6432 1349
rect 6328 1112 6432 1125
rect 6488 1349 6592 1362
rect 6488 1125 6517 1349
rect 6563 1125 6592 1349
rect 6488 1112 6592 1125
rect 6648 1349 6752 1362
rect 6648 1125 6677 1349
rect 6723 1125 6752 1349
rect 6648 1112 6752 1125
rect 6808 1349 6896 1362
rect 6808 1125 6837 1349
rect 6883 1125 6896 1349
rect 6808 1112 6896 1125
rect 6952 1349 7040 1362
rect 6952 1125 6965 1349
rect 7011 1125 7040 1349
rect 6952 1112 7040 1125
rect 7096 1349 7184 1362
rect 7096 1125 7125 1349
rect 7171 1125 7184 1349
rect 7096 1112 7184 1125
rect 7356 1349 7444 1362
rect 7356 1125 7369 1349
rect 7415 1125 7444 1349
rect 7356 1112 7444 1125
rect 7500 1349 7604 1362
rect 7500 1125 7529 1349
rect 7575 1125 7604 1349
rect 7500 1112 7604 1125
rect 7660 1349 7764 1362
rect 7660 1125 7689 1349
rect 7735 1125 7764 1349
rect 7660 1112 7764 1125
rect 7820 1349 7924 1362
rect 7820 1125 7849 1349
rect 7895 1125 7924 1349
rect 7820 1112 7924 1125
rect 7980 1349 8084 1362
rect 7980 1125 8009 1349
rect 8055 1125 8084 1349
rect 7980 1112 8084 1125
rect 8140 1349 8244 1362
rect 8140 1125 8169 1349
rect 8215 1125 8244 1349
rect 8140 1112 8244 1125
rect 8300 1349 8404 1362
rect 8300 1125 8329 1349
rect 8375 1125 8404 1349
rect 8300 1112 8404 1125
rect 8460 1349 8564 1362
rect 8460 1125 8489 1349
rect 8535 1125 8564 1349
rect 8460 1112 8564 1125
rect 8620 1349 8708 1362
rect 8620 1125 8649 1349
rect 8695 1125 8708 1349
rect 8620 1112 8708 1125
rect 8764 1349 8852 1362
rect 8764 1125 8777 1349
rect 8823 1125 8852 1349
rect 8764 1112 8852 1125
rect 8908 1349 8996 1362
rect 8908 1125 8937 1349
rect 8983 1125 8996 1349
rect 8908 1112 8996 1125
rect -4812 1006 -4724 1019
rect -4812 932 -4799 1006
rect -4753 932 -4724 1006
rect -4812 919 -4724 932
rect -4668 1006 -4580 1019
rect -4668 932 -4639 1006
rect -4593 932 -4580 1006
rect -4668 919 -4580 932
rect -4246 1018 -4158 1031
rect -4246 944 -4233 1018
rect -4187 944 -4158 1018
rect -4246 931 -4158 944
rect -4102 1018 -3998 1031
rect -4102 944 -4073 1018
rect -4027 944 -3998 1018
rect -4102 931 -3998 944
rect -3942 1018 -3854 1031
rect -3942 944 -3913 1018
rect -3867 944 -3854 1018
rect -3541 1030 -3469 1043
rect -3541 984 -3528 1030
rect -3482 1029 -3469 1030
rect -2981 1030 -2909 1043
rect -2981 1029 -2968 1030
rect -3482 985 -3449 1029
rect -3001 985 -2968 1029
rect -3482 984 -3469 985
rect -3541 971 -3469 984
rect -3942 931 -3854 944
rect -2981 984 -2968 985
rect -2922 984 -2909 1030
rect -2981 971 -2909 984
rect -2755 1030 -2683 1043
rect -2755 984 -2742 1030
rect -2696 1029 -2683 1030
rect -2195 1030 -2123 1043
rect -2195 1029 -2182 1030
rect -2696 985 -2663 1029
rect -2215 985 -2182 1029
rect -2696 984 -2683 985
rect -2755 971 -2683 984
rect -2195 984 -2182 985
rect -2136 984 -2123 1030
rect -2195 971 -2123 984
rect -1969 1030 -1897 1043
rect -1969 984 -1956 1030
rect -1910 1029 -1897 1030
rect -1409 1030 -1337 1043
rect -1409 1029 -1396 1030
rect -1910 985 -1877 1029
rect -1429 985 -1396 1029
rect -1910 984 -1897 985
rect -1969 971 -1897 984
rect -1409 984 -1396 985
rect -1350 984 -1337 1030
rect -1409 971 -1337 984
rect -1163 1006 -1075 1019
rect -1163 932 -1150 1006
rect -1104 932 -1075 1006
rect -1163 919 -1075 932
rect -1019 1006 -931 1019
rect -1019 932 -990 1006
rect -944 932 -931 1006
rect -1019 919 -931 932
rect 108 963 196 976
rect 108 739 121 963
rect 167 739 196 963
rect 108 726 196 739
rect 252 963 340 976
rect 252 739 281 963
rect 327 739 340 963
rect 252 726 340 739
rect 396 963 484 976
rect 396 739 409 963
rect 455 739 484 963
rect 396 726 484 739
rect 540 963 644 976
rect 540 739 569 963
rect 615 739 644 963
rect 540 726 644 739
rect 700 963 804 976
rect 700 739 729 963
rect 775 739 804 963
rect 700 726 804 739
rect 860 963 964 976
rect 860 739 889 963
rect 935 739 964 963
rect 860 726 964 739
rect 1020 963 1124 976
rect 1020 739 1049 963
rect 1095 739 1124 963
rect 1020 726 1124 739
rect 1180 963 1284 976
rect 1180 739 1209 963
rect 1255 739 1284 963
rect 1180 726 1284 739
rect 1340 963 1444 976
rect 1340 739 1369 963
rect 1415 739 1444 963
rect 1340 726 1444 739
rect 1500 963 1604 976
rect 1500 739 1529 963
rect 1575 739 1604 963
rect 1500 726 1604 739
rect 1660 963 1748 976
rect 1660 739 1689 963
rect 1735 739 1748 963
rect 1660 726 1748 739
rect 1920 963 2008 976
rect 1920 739 1933 963
rect 1979 739 2008 963
rect 1920 726 2008 739
rect 2064 963 2168 976
rect 2064 739 2093 963
rect 2139 739 2168 963
rect 2064 726 2168 739
rect 2224 963 2328 976
rect 2224 739 2253 963
rect 2299 739 2328 963
rect 2224 726 2328 739
rect 2384 963 2488 976
rect 2384 739 2413 963
rect 2459 739 2488 963
rect 2384 726 2488 739
rect 2544 963 2648 976
rect 2544 739 2573 963
rect 2619 739 2648 963
rect 2544 726 2648 739
rect 2704 963 2808 976
rect 2704 739 2733 963
rect 2779 739 2808 963
rect 2704 726 2808 739
rect 2864 963 2968 976
rect 2864 739 2893 963
rect 2939 739 2968 963
rect 2864 726 2968 739
rect 3024 963 3128 976
rect 3024 739 3053 963
rect 3099 739 3128 963
rect 3024 726 3128 739
rect 3184 963 3272 976
rect 3184 739 3213 963
rect 3259 739 3272 963
rect 3184 726 3272 739
rect 3328 963 3416 976
rect 3328 739 3341 963
rect 3387 739 3416 963
rect 3328 726 3416 739
rect 3472 963 3560 976
rect 3472 739 3501 963
rect 3547 739 3560 963
rect 3472 726 3560 739
rect 3732 963 3820 976
rect 3732 739 3745 963
rect 3791 739 3820 963
rect 3732 726 3820 739
rect 3876 963 3964 976
rect 3876 739 3905 963
rect 3951 739 3964 963
rect 3876 726 3964 739
rect 4020 963 4108 976
rect 4020 739 4033 963
rect 4079 739 4108 963
rect 4020 726 4108 739
rect 4164 963 4268 976
rect 4164 739 4193 963
rect 4239 739 4268 963
rect 4164 726 4268 739
rect 4324 963 4428 976
rect 4324 739 4353 963
rect 4399 739 4428 963
rect 4324 726 4428 739
rect 4484 963 4588 976
rect 4484 739 4513 963
rect 4559 739 4588 963
rect 4484 726 4588 739
rect 4644 963 4748 976
rect 4644 739 4673 963
rect 4719 739 4748 963
rect 4644 726 4748 739
rect 4804 963 4908 976
rect 4804 739 4833 963
rect 4879 739 4908 963
rect 4804 726 4908 739
rect 4964 963 5068 976
rect 4964 739 4993 963
rect 5039 739 5068 963
rect 4964 726 5068 739
rect 5124 963 5228 976
rect 5124 739 5153 963
rect 5199 739 5228 963
rect 5124 726 5228 739
rect 5284 963 5372 976
rect 5284 739 5313 963
rect 5359 739 5372 963
rect 5284 726 5372 739
rect 5544 963 5632 976
rect 5544 739 5557 963
rect 5603 739 5632 963
rect 5544 726 5632 739
rect 5688 963 5792 976
rect 5688 739 5717 963
rect 5763 739 5792 963
rect 5688 726 5792 739
rect 5848 963 5952 976
rect 5848 739 5877 963
rect 5923 739 5952 963
rect 5848 726 5952 739
rect 6008 963 6112 976
rect 6008 739 6037 963
rect 6083 739 6112 963
rect 6008 726 6112 739
rect 6168 963 6272 976
rect 6168 739 6197 963
rect 6243 739 6272 963
rect 6168 726 6272 739
rect 6328 963 6432 976
rect 6328 739 6357 963
rect 6403 739 6432 963
rect 6328 726 6432 739
rect 6488 963 6592 976
rect 6488 739 6517 963
rect 6563 739 6592 963
rect 6488 726 6592 739
rect 6648 963 6752 976
rect 6648 739 6677 963
rect 6723 739 6752 963
rect 6648 726 6752 739
rect 6808 963 6896 976
rect 6808 739 6837 963
rect 6883 739 6896 963
rect 6808 726 6896 739
rect 6952 963 7040 976
rect 6952 739 6965 963
rect 7011 739 7040 963
rect 6952 726 7040 739
rect 7096 963 7184 976
rect 7096 739 7125 963
rect 7171 739 7184 963
rect 7096 726 7184 739
rect 7356 963 7444 976
rect 7356 739 7369 963
rect 7415 739 7444 963
rect 7356 726 7444 739
rect 7500 963 7604 976
rect 7500 739 7529 963
rect 7575 739 7604 963
rect 7500 726 7604 739
rect 7660 963 7764 976
rect 7660 739 7689 963
rect 7735 739 7764 963
rect 7660 726 7764 739
rect 7820 963 7924 976
rect 7820 739 7849 963
rect 7895 739 7924 963
rect 7820 726 7924 739
rect 7980 963 8084 976
rect 7980 739 8009 963
rect 8055 739 8084 963
rect 7980 726 8084 739
rect 8140 963 8244 976
rect 8140 739 8169 963
rect 8215 739 8244 963
rect 8140 726 8244 739
rect 8300 963 8404 976
rect 8300 739 8329 963
rect 8375 739 8404 963
rect 8300 726 8404 739
rect 8460 963 8564 976
rect 8460 739 8489 963
rect 8535 739 8564 963
rect 8460 726 8564 739
rect 8620 963 8708 976
rect 8620 739 8649 963
rect 8695 739 8708 963
rect 8620 726 8708 739
rect 8764 963 8852 976
rect 8764 739 8777 963
rect 8823 739 8852 963
rect 8764 726 8852 739
rect 8908 963 8996 976
rect 8908 739 8937 963
rect 8983 739 8996 963
rect 8908 726 8996 739
rect 108 577 196 590
rect 108 353 121 577
rect 167 353 196 577
rect 108 340 196 353
rect 252 577 340 590
rect 252 353 281 577
rect 327 353 340 577
rect 252 340 340 353
rect 396 577 484 590
rect 396 353 409 577
rect 455 353 484 577
rect 396 340 484 353
rect 540 577 644 590
rect 540 353 569 577
rect 615 353 644 577
rect 540 340 644 353
rect 700 577 804 590
rect 700 353 729 577
rect 775 353 804 577
rect 700 340 804 353
rect 860 577 964 590
rect 860 353 889 577
rect 935 353 964 577
rect 860 340 964 353
rect 1020 577 1124 590
rect 1020 353 1049 577
rect 1095 353 1124 577
rect 1020 340 1124 353
rect 1180 577 1284 590
rect 1180 353 1209 577
rect 1255 353 1284 577
rect 1180 340 1284 353
rect 1340 577 1444 590
rect 1340 353 1369 577
rect 1415 353 1444 577
rect 1340 340 1444 353
rect 1500 577 1604 590
rect 1500 353 1529 577
rect 1575 353 1604 577
rect 1500 340 1604 353
rect 1660 577 1748 590
rect 1660 353 1689 577
rect 1735 353 1748 577
rect 1660 340 1748 353
rect 1920 577 2008 590
rect 1920 353 1933 577
rect 1979 353 2008 577
rect 1920 340 2008 353
rect 2064 577 2168 590
rect 2064 353 2093 577
rect 2139 353 2168 577
rect 2064 340 2168 353
rect 2224 577 2328 590
rect 2224 353 2253 577
rect 2299 353 2328 577
rect 2224 340 2328 353
rect 2384 577 2488 590
rect 2384 353 2413 577
rect 2459 353 2488 577
rect 2384 340 2488 353
rect 2544 577 2648 590
rect 2544 353 2573 577
rect 2619 353 2648 577
rect 2544 340 2648 353
rect 2704 577 2808 590
rect 2704 353 2733 577
rect 2779 353 2808 577
rect 2704 340 2808 353
rect 2864 577 2968 590
rect 2864 353 2893 577
rect 2939 353 2968 577
rect 2864 340 2968 353
rect 3024 577 3128 590
rect 3024 353 3053 577
rect 3099 353 3128 577
rect 3024 340 3128 353
rect 3184 577 3272 590
rect 3184 353 3213 577
rect 3259 353 3272 577
rect 3184 340 3272 353
rect 3328 577 3416 590
rect 3328 353 3341 577
rect 3387 353 3416 577
rect 3328 340 3416 353
rect 3472 577 3560 590
rect 3472 353 3501 577
rect 3547 353 3560 577
rect 3472 340 3560 353
rect 3732 577 3820 590
rect 3732 353 3745 577
rect 3791 353 3820 577
rect 3732 340 3820 353
rect 3876 577 3964 590
rect 3876 353 3905 577
rect 3951 353 3964 577
rect 3876 340 3964 353
rect 4020 577 4108 590
rect 4020 353 4033 577
rect 4079 353 4108 577
rect 4020 340 4108 353
rect 4164 577 4268 590
rect 4164 353 4193 577
rect 4239 353 4268 577
rect 4164 340 4268 353
rect 4324 577 4428 590
rect 4324 353 4353 577
rect 4399 353 4428 577
rect 4324 340 4428 353
rect 4484 577 4588 590
rect 4484 353 4513 577
rect 4559 353 4588 577
rect 4484 340 4588 353
rect 4644 577 4748 590
rect 4644 353 4673 577
rect 4719 353 4748 577
rect 4644 340 4748 353
rect 4804 577 4908 590
rect 4804 353 4833 577
rect 4879 353 4908 577
rect 4804 340 4908 353
rect 4964 577 5068 590
rect 4964 353 4993 577
rect 5039 353 5068 577
rect 4964 340 5068 353
rect 5124 577 5228 590
rect 5124 353 5153 577
rect 5199 353 5228 577
rect 5124 340 5228 353
rect 5284 577 5372 590
rect 5284 353 5313 577
rect 5359 353 5372 577
rect 5284 340 5372 353
rect 5544 577 5632 590
rect 5544 353 5557 577
rect 5603 353 5632 577
rect 5544 340 5632 353
rect 5688 577 5792 590
rect 5688 353 5717 577
rect 5763 353 5792 577
rect 5688 340 5792 353
rect 5848 577 5952 590
rect 5848 353 5877 577
rect 5923 353 5952 577
rect 5848 340 5952 353
rect 6008 577 6112 590
rect 6008 353 6037 577
rect 6083 353 6112 577
rect 6008 340 6112 353
rect 6168 577 6272 590
rect 6168 353 6197 577
rect 6243 353 6272 577
rect 6168 340 6272 353
rect 6328 577 6432 590
rect 6328 353 6357 577
rect 6403 353 6432 577
rect 6328 340 6432 353
rect 6488 577 6592 590
rect 6488 353 6517 577
rect 6563 353 6592 577
rect 6488 340 6592 353
rect 6648 577 6752 590
rect 6648 353 6677 577
rect 6723 353 6752 577
rect 6648 340 6752 353
rect 6808 577 6896 590
rect 6808 353 6837 577
rect 6883 353 6896 577
rect 6808 340 6896 353
rect 6952 577 7040 590
rect 6952 353 6965 577
rect 7011 353 7040 577
rect 6952 340 7040 353
rect 7096 577 7184 590
rect 7096 353 7125 577
rect 7171 353 7184 577
rect 7096 340 7184 353
rect 7356 577 7444 590
rect 7356 353 7369 577
rect 7415 353 7444 577
rect 7356 340 7444 353
rect 7500 577 7604 590
rect 7500 353 7529 577
rect 7575 353 7604 577
rect 7500 340 7604 353
rect 7660 577 7764 590
rect 7660 353 7689 577
rect 7735 353 7764 577
rect 7660 340 7764 353
rect 7820 577 7924 590
rect 7820 353 7849 577
rect 7895 353 7924 577
rect 7820 340 7924 353
rect 7980 577 8084 590
rect 7980 353 8009 577
rect 8055 353 8084 577
rect 7980 340 8084 353
rect 8140 577 8244 590
rect 8140 353 8169 577
rect 8215 353 8244 577
rect 8140 340 8244 353
rect 8300 577 8404 590
rect 8300 353 8329 577
rect 8375 353 8404 577
rect 8300 340 8404 353
rect 8460 577 8564 590
rect 8460 353 8489 577
rect 8535 353 8564 577
rect 8460 340 8564 353
rect 8620 577 8708 590
rect 8620 353 8649 577
rect 8695 353 8708 577
rect 8620 340 8708 353
rect 8764 577 8852 590
rect 8764 353 8777 577
rect 8823 353 8852 577
rect 8764 340 8852 353
rect 8908 577 8996 590
rect 8908 353 8937 577
rect 8983 353 8996 577
rect 8908 340 8996 353
rect -4812 -332 -4724 -319
rect -4812 -406 -4799 -332
rect -4753 -406 -4724 -332
rect -4812 -419 -4724 -406
rect -4668 -332 -4580 -319
rect -4668 -406 -4639 -332
rect -4593 -406 -4580 -332
rect -4668 -419 -4580 -406
rect -4246 -344 -4158 -331
rect -4246 -418 -4233 -344
rect -4187 -418 -4158 -344
rect -4246 -431 -4158 -418
rect -4102 -344 -3998 -331
rect -4102 -418 -4073 -344
rect -4027 -418 -3998 -344
rect -4102 -431 -3998 -418
rect -3942 -344 -3854 -331
rect 108 -241 196 -228
rect -1163 -332 -1075 -319
rect -3942 -418 -3913 -344
rect -3867 -418 -3854 -344
rect -3942 -431 -3854 -418
rect -3541 -384 -3469 -371
rect -3541 -430 -3528 -384
rect -3482 -385 -3469 -384
rect -2981 -384 -2909 -371
rect -2981 -385 -2968 -384
rect -3482 -429 -3449 -385
rect -3001 -429 -2968 -385
rect -3482 -430 -3469 -429
rect -3541 -443 -3469 -430
rect -2981 -430 -2968 -429
rect -2922 -430 -2909 -384
rect -2981 -443 -2909 -430
rect -2755 -384 -2683 -371
rect -2755 -430 -2742 -384
rect -2696 -385 -2683 -384
rect -2195 -384 -2123 -371
rect -2195 -385 -2182 -384
rect -2696 -429 -2663 -385
rect -2215 -429 -2182 -385
rect -2696 -430 -2683 -429
rect -2755 -443 -2683 -430
rect -2195 -430 -2182 -429
rect -2136 -430 -2123 -384
rect -2195 -443 -2123 -430
rect -1969 -384 -1897 -371
rect -1969 -430 -1956 -384
rect -1910 -385 -1897 -384
rect -1409 -384 -1337 -371
rect -1409 -385 -1396 -384
rect -1910 -429 -1877 -385
rect -1429 -429 -1396 -385
rect -1910 -430 -1897 -429
rect -1969 -443 -1897 -430
rect -1409 -430 -1396 -429
rect -1350 -430 -1337 -384
rect -1163 -406 -1150 -332
rect -1104 -406 -1075 -332
rect -1163 -419 -1075 -406
rect -1019 -332 -931 -319
rect -1019 -406 -990 -332
rect -944 -406 -931 -332
rect -1019 -419 -931 -406
rect -1409 -443 -1337 -430
rect 108 -465 121 -241
rect 167 -465 196 -241
rect 108 -478 196 -465
rect 252 -241 340 -228
rect 252 -465 281 -241
rect 327 -465 340 -241
rect 252 -478 340 -465
rect 396 -241 484 -228
rect 396 -465 409 -241
rect 455 -465 484 -241
rect 396 -478 484 -465
rect 540 -241 644 -228
rect 540 -465 569 -241
rect 615 -465 644 -241
rect 540 -478 644 -465
rect 700 -241 804 -228
rect 700 -465 729 -241
rect 775 -465 804 -241
rect 700 -478 804 -465
rect 860 -241 964 -228
rect 860 -465 889 -241
rect 935 -465 964 -241
rect 860 -478 964 -465
rect 1020 -241 1124 -228
rect 1020 -465 1049 -241
rect 1095 -465 1124 -241
rect 1020 -478 1124 -465
rect 1180 -241 1284 -228
rect 1180 -465 1209 -241
rect 1255 -465 1284 -241
rect 1180 -478 1284 -465
rect 1340 -241 1444 -228
rect 1340 -465 1369 -241
rect 1415 -465 1444 -241
rect 1340 -478 1444 -465
rect 1500 -241 1604 -228
rect 1500 -465 1529 -241
rect 1575 -465 1604 -241
rect 1500 -478 1604 -465
rect 1660 -241 1748 -228
rect 1660 -465 1689 -241
rect 1735 -465 1748 -241
rect 1660 -478 1748 -465
rect 1920 -241 2008 -228
rect 1920 -465 1933 -241
rect 1979 -465 2008 -241
rect 1920 -478 2008 -465
rect 2064 -241 2168 -228
rect 2064 -465 2093 -241
rect 2139 -465 2168 -241
rect 2064 -478 2168 -465
rect 2224 -241 2328 -228
rect 2224 -465 2253 -241
rect 2299 -465 2328 -241
rect 2224 -478 2328 -465
rect 2384 -241 2488 -228
rect 2384 -465 2413 -241
rect 2459 -465 2488 -241
rect 2384 -478 2488 -465
rect 2544 -241 2648 -228
rect 2544 -465 2573 -241
rect 2619 -465 2648 -241
rect 2544 -478 2648 -465
rect 2704 -241 2808 -228
rect 2704 -465 2733 -241
rect 2779 -465 2808 -241
rect 2704 -478 2808 -465
rect 2864 -241 2968 -228
rect 2864 -465 2893 -241
rect 2939 -465 2968 -241
rect 2864 -478 2968 -465
rect 3024 -241 3128 -228
rect 3024 -465 3053 -241
rect 3099 -465 3128 -241
rect 3024 -478 3128 -465
rect 3184 -241 3272 -228
rect 3184 -465 3213 -241
rect 3259 -465 3272 -241
rect 3184 -478 3272 -465
rect 3328 -241 3416 -228
rect 3328 -465 3341 -241
rect 3387 -465 3416 -241
rect 3328 -478 3416 -465
rect 3472 -241 3560 -228
rect 3472 -465 3501 -241
rect 3547 -465 3560 -241
rect 3472 -478 3560 -465
rect 3732 -241 3820 -228
rect 3732 -465 3745 -241
rect 3791 -465 3820 -241
rect 3732 -478 3820 -465
rect 3876 -241 3964 -228
rect 3876 -465 3905 -241
rect 3951 -465 3964 -241
rect 3876 -478 3964 -465
rect 4020 -241 4108 -228
rect 4020 -465 4033 -241
rect 4079 -465 4108 -241
rect 4020 -478 4108 -465
rect 4164 -241 4268 -228
rect 4164 -465 4193 -241
rect 4239 -465 4268 -241
rect 4164 -478 4268 -465
rect 4324 -241 4428 -228
rect 4324 -465 4353 -241
rect 4399 -465 4428 -241
rect 4324 -478 4428 -465
rect 4484 -241 4588 -228
rect 4484 -465 4513 -241
rect 4559 -465 4588 -241
rect 4484 -478 4588 -465
rect 4644 -241 4748 -228
rect 4644 -465 4673 -241
rect 4719 -465 4748 -241
rect 4644 -478 4748 -465
rect 4804 -241 4908 -228
rect 4804 -465 4833 -241
rect 4879 -465 4908 -241
rect 4804 -478 4908 -465
rect 4964 -241 5068 -228
rect 4964 -465 4993 -241
rect 5039 -465 5068 -241
rect 4964 -478 5068 -465
rect 5124 -241 5228 -228
rect 5124 -465 5153 -241
rect 5199 -465 5228 -241
rect 5124 -478 5228 -465
rect 5284 -241 5372 -228
rect 5284 -465 5313 -241
rect 5359 -465 5372 -241
rect 5284 -478 5372 -465
rect 5544 -241 5632 -228
rect 5544 -465 5557 -241
rect 5603 -465 5632 -241
rect 5544 -478 5632 -465
rect 5688 -241 5792 -228
rect 5688 -465 5717 -241
rect 5763 -465 5792 -241
rect 5688 -478 5792 -465
rect 5848 -241 5952 -228
rect 5848 -465 5877 -241
rect 5923 -465 5952 -241
rect 5848 -478 5952 -465
rect 6008 -241 6112 -228
rect 6008 -465 6037 -241
rect 6083 -465 6112 -241
rect 6008 -478 6112 -465
rect 6168 -241 6272 -228
rect 6168 -465 6197 -241
rect 6243 -465 6272 -241
rect 6168 -478 6272 -465
rect 6328 -241 6432 -228
rect 6328 -465 6357 -241
rect 6403 -465 6432 -241
rect 6328 -478 6432 -465
rect 6488 -241 6592 -228
rect 6488 -465 6517 -241
rect 6563 -465 6592 -241
rect 6488 -478 6592 -465
rect 6648 -241 6752 -228
rect 6648 -465 6677 -241
rect 6723 -465 6752 -241
rect 6648 -478 6752 -465
rect 6808 -241 6896 -228
rect 6808 -465 6837 -241
rect 6883 -465 6896 -241
rect 6808 -478 6896 -465
rect 6952 -241 7040 -228
rect 6952 -465 6965 -241
rect 7011 -465 7040 -241
rect 6952 -478 7040 -465
rect 7096 -241 7184 -228
rect 7096 -465 7125 -241
rect 7171 -465 7184 -241
rect 7096 -478 7184 -465
rect 7356 -241 7444 -228
rect 7356 -465 7369 -241
rect 7415 -465 7444 -241
rect 7356 -478 7444 -465
rect 7500 -241 7604 -228
rect 7500 -465 7529 -241
rect 7575 -465 7604 -241
rect 7500 -478 7604 -465
rect 7660 -241 7764 -228
rect 7660 -465 7689 -241
rect 7735 -465 7764 -241
rect 7660 -478 7764 -465
rect 7820 -241 7924 -228
rect 7820 -465 7849 -241
rect 7895 -465 7924 -241
rect 7820 -478 7924 -465
rect 7980 -241 8084 -228
rect 7980 -465 8009 -241
rect 8055 -465 8084 -241
rect 7980 -478 8084 -465
rect 8140 -241 8244 -228
rect 8140 -465 8169 -241
rect 8215 -465 8244 -241
rect 8140 -478 8244 -465
rect 8300 -241 8404 -228
rect 8300 -465 8329 -241
rect 8375 -465 8404 -241
rect 8300 -478 8404 -465
rect 8460 -241 8564 -228
rect 8460 -465 8489 -241
rect 8535 -465 8564 -241
rect 8460 -478 8564 -465
rect 8620 -241 8708 -228
rect 8620 -465 8649 -241
rect 8695 -465 8708 -241
rect 8620 -478 8708 -465
rect 8764 -241 8852 -228
rect 8764 -465 8777 -241
rect 8823 -465 8852 -241
rect 8764 -478 8852 -465
rect 8908 -241 8996 -228
rect 8908 -465 8937 -241
rect 8983 -465 8996 -241
rect 8908 -478 8996 -465
rect 108 -627 196 -614
rect -4246 -692 -4158 -679
rect -4246 -766 -4233 -692
rect -4187 -766 -4158 -692
rect -4246 -779 -4158 -766
rect -4102 -692 -3998 -679
rect -4102 -766 -4073 -692
rect -4027 -766 -3998 -692
rect -4102 -779 -3998 -766
rect -3942 -692 -3854 -679
rect -3942 -766 -3913 -692
rect -3867 -766 -3854 -692
rect -3541 -680 -3469 -667
rect -3541 -726 -3528 -680
rect -3482 -681 -3469 -680
rect -2981 -680 -2909 -667
rect -2981 -681 -2968 -680
rect -3482 -725 -3449 -681
rect -3001 -725 -2968 -681
rect -3482 -726 -3469 -725
rect -3541 -739 -3469 -726
rect -3942 -779 -3854 -766
rect -2981 -726 -2968 -725
rect -2922 -726 -2909 -680
rect -2981 -739 -2909 -726
rect -2755 -680 -2683 -667
rect -2755 -726 -2742 -680
rect -2696 -681 -2683 -680
rect -2195 -680 -2123 -667
rect -2195 -681 -2182 -680
rect -2696 -725 -2663 -681
rect -2215 -725 -2182 -681
rect -2696 -726 -2683 -725
rect -2755 -739 -2683 -726
rect -2195 -726 -2182 -725
rect -2136 -726 -2123 -680
rect -2195 -739 -2123 -726
rect -1969 -680 -1897 -667
rect -1969 -726 -1956 -680
rect -1910 -681 -1897 -680
rect -1409 -680 -1337 -667
rect -1409 -681 -1396 -680
rect -1910 -725 -1877 -681
rect -1429 -725 -1396 -681
rect -1910 -726 -1897 -725
rect -1969 -739 -1897 -726
rect -1409 -726 -1396 -725
rect -1350 -726 -1337 -680
rect -1409 -739 -1337 -726
rect -1163 -704 -1075 -691
rect -1163 -778 -1150 -704
rect -1104 -778 -1075 -704
rect -1163 -791 -1075 -778
rect -1019 -704 -931 -691
rect -1019 -778 -990 -704
rect -944 -778 -931 -704
rect -1019 -791 -931 -778
rect 108 -851 121 -627
rect 167 -851 196 -627
rect 108 -864 196 -851
rect 252 -627 340 -614
rect 252 -851 281 -627
rect 327 -851 340 -627
rect 252 -864 340 -851
rect 396 -627 484 -614
rect 396 -851 409 -627
rect 455 -851 484 -627
rect 396 -864 484 -851
rect 540 -627 644 -614
rect 540 -851 569 -627
rect 615 -851 644 -627
rect 540 -864 644 -851
rect 700 -627 804 -614
rect 700 -851 729 -627
rect 775 -851 804 -627
rect 700 -864 804 -851
rect 860 -627 964 -614
rect 860 -851 889 -627
rect 935 -851 964 -627
rect 860 -864 964 -851
rect 1020 -627 1124 -614
rect 1020 -851 1049 -627
rect 1095 -851 1124 -627
rect 1020 -864 1124 -851
rect 1180 -627 1284 -614
rect 1180 -851 1209 -627
rect 1255 -851 1284 -627
rect 1180 -864 1284 -851
rect 1340 -627 1444 -614
rect 1340 -851 1369 -627
rect 1415 -851 1444 -627
rect 1340 -864 1444 -851
rect 1500 -627 1604 -614
rect 1500 -851 1529 -627
rect 1575 -851 1604 -627
rect 1500 -864 1604 -851
rect 1660 -627 1748 -614
rect 1660 -851 1689 -627
rect 1735 -851 1748 -627
rect 1660 -864 1748 -851
rect 1920 -627 2008 -614
rect 1920 -851 1933 -627
rect 1979 -851 2008 -627
rect 1920 -864 2008 -851
rect 2064 -627 2168 -614
rect 2064 -851 2093 -627
rect 2139 -851 2168 -627
rect 2064 -864 2168 -851
rect 2224 -627 2328 -614
rect 2224 -851 2253 -627
rect 2299 -851 2328 -627
rect 2224 -864 2328 -851
rect 2384 -627 2488 -614
rect 2384 -851 2413 -627
rect 2459 -851 2488 -627
rect 2384 -864 2488 -851
rect 2544 -627 2648 -614
rect 2544 -851 2573 -627
rect 2619 -851 2648 -627
rect 2544 -864 2648 -851
rect 2704 -627 2808 -614
rect 2704 -851 2733 -627
rect 2779 -851 2808 -627
rect 2704 -864 2808 -851
rect 2864 -627 2968 -614
rect 2864 -851 2893 -627
rect 2939 -851 2968 -627
rect 2864 -864 2968 -851
rect 3024 -627 3128 -614
rect 3024 -851 3053 -627
rect 3099 -851 3128 -627
rect 3024 -864 3128 -851
rect 3184 -627 3272 -614
rect 3184 -851 3213 -627
rect 3259 -851 3272 -627
rect 3184 -864 3272 -851
rect 3328 -627 3416 -614
rect 3328 -851 3341 -627
rect 3387 -851 3416 -627
rect 3328 -864 3416 -851
rect 3472 -627 3560 -614
rect 3472 -851 3501 -627
rect 3547 -851 3560 -627
rect 3472 -864 3560 -851
rect 3732 -627 3820 -614
rect 3732 -851 3745 -627
rect 3791 -851 3820 -627
rect 3732 -864 3820 -851
rect 3876 -627 3964 -614
rect 3876 -851 3905 -627
rect 3951 -851 3964 -627
rect 3876 -864 3964 -851
rect 4020 -627 4108 -614
rect 4020 -851 4033 -627
rect 4079 -851 4108 -627
rect 4020 -864 4108 -851
rect 4164 -627 4268 -614
rect 4164 -851 4193 -627
rect 4239 -851 4268 -627
rect 4164 -864 4268 -851
rect 4324 -627 4428 -614
rect 4324 -851 4353 -627
rect 4399 -851 4428 -627
rect 4324 -864 4428 -851
rect 4484 -627 4588 -614
rect 4484 -851 4513 -627
rect 4559 -851 4588 -627
rect 4484 -864 4588 -851
rect 4644 -627 4748 -614
rect 4644 -851 4673 -627
rect 4719 -851 4748 -627
rect 4644 -864 4748 -851
rect 4804 -627 4908 -614
rect 4804 -851 4833 -627
rect 4879 -851 4908 -627
rect 4804 -864 4908 -851
rect 4964 -627 5068 -614
rect 4964 -851 4993 -627
rect 5039 -851 5068 -627
rect 4964 -864 5068 -851
rect 5124 -627 5228 -614
rect 5124 -851 5153 -627
rect 5199 -851 5228 -627
rect 5124 -864 5228 -851
rect 5284 -627 5372 -614
rect 5284 -851 5313 -627
rect 5359 -851 5372 -627
rect 5284 -864 5372 -851
rect 5544 -627 5632 -614
rect 5544 -851 5557 -627
rect 5603 -851 5632 -627
rect 5544 -864 5632 -851
rect 5688 -627 5792 -614
rect 5688 -851 5717 -627
rect 5763 -851 5792 -627
rect 5688 -864 5792 -851
rect 5848 -627 5952 -614
rect 5848 -851 5877 -627
rect 5923 -851 5952 -627
rect 5848 -864 5952 -851
rect 6008 -627 6112 -614
rect 6008 -851 6037 -627
rect 6083 -851 6112 -627
rect 6008 -864 6112 -851
rect 6168 -627 6272 -614
rect 6168 -851 6197 -627
rect 6243 -851 6272 -627
rect 6168 -864 6272 -851
rect 6328 -627 6432 -614
rect 6328 -851 6357 -627
rect 6403 -851 6432 -627
rect 6328 -864 6432 -851
rect 6488 -627 6592 -614
rect 6488 -851 6517 -627
rect 6563 -851 6592 -627
rect 6488 -864 6592 -851
rect 6648 -627 6752 -614
rect 6648 -851 6677 -627
rect 6723 -851 6752 -627
rect 6648 -864 6752 -851
rect 6808 -627 6896 -614
rect 6808 -851 6837 -627
rect 6883 -851 6896 -627
rect 6808 -864 6896 -851
rect 6952 -627 7040 -614
rect 6952 -851 6965 -627
rect 7011 -851 7040 -627
rect 6952 -864 7040 -851
rect 7096 -627 7184 -614
rect 7096 -851 7125 -627
rect 7171 -851 7184 -627
rect 7096 -864 7184 -851
rect 7356 -627 7444 -614
rect 7356 -851 7369 -627
rect 7415 -851 7444 -627
rect 7356 -864 7444 -851
rect 7500 -627 7604 -614
rect 7500 -851 7529 -627
rect 7575 -851 7604 -627
rect 7500 -864 7604 -851
rect 7660 -627 7764 -614
rect 7660 -851 7689 -627
rect 7735 -851 7764 -627
rect 7660 -864 7764 -851
rect 7820 -627 7924 -614
rect 7820 -851 7849 -627
rect 7895 -851 7924 -627
rect 7820 -864 7924 -851
rect 7980 -627 8084 -614
rect 7980 -851 8009 -627
rect 8055 -851 8084 -627
rect 7980 -864 8084 -851
rect 8140 -627 8244 -614
rect 8140 -851 8169 -627
rect 8215 -851 8244 -627
rect 8140 -864 8244 -851
rect 8300 -627 8404 -614
rect 8300 -851 8329 -627
rect 8375 -851 8404 -627
rect 8300 -864 8404 -851
rect 8460 -627 8564 -614
rect 8460 -851 8489 -627
rect 8535 -851 8564 -627
rect 8460 -864 8564 -851
rect 8620 -627 8708 -614
rect 8620 -851 8649 -627
rect 8695 -851 8708 -627
rect 8620 -864 8708 -851
rect 8764 -627 8852 -614
rect 8764 -851 8777 -627
rect 8823 -851 8852 -627
rect 8764 -864 8852 -851
rect 8908 -627 8996 -614
rect 8908 -851 8937 -627
rect 8983 -851 8996 -627
rect 8908 -864 8996 -851
rect 108 -1013 196 -1000
rect 108 -1237 121 -1013
rect 167 -1237 196 -1013
rect 108 -1250 196 -1237
rect 252 -1013 340 -1000
rect 252 -1237 281 -1013
rect 327 -1237 340 -1013
rect 252 -1250 340 -1237
rect 396 -1013 484 -1000
rect 396 -1237 409 -1013
rect 455 -1237 484 -1013
rect 396 -1250 484 -1237
rect 540 -1013 644 -1000
rect 540 -1237 569 -1013
rect 615 -1237 644 -1013
rect 540 -1250 644 -1237
rect 700 -1013 804 -1000
rect 700 -1237 729 -1013
rect 775 -1237 804 -1013
rect 700 -1250 804 -1237
rect 860 -1013 964 -1000
rect 860 -1237 889 -1013
rect 935 -1237 964 -1013
rect 860 -1250 964 -1237
rect 1020 -1013 1124 -1000
rect 1020 -1237 1049 -1013
rect 1095 -1237 1124 -1013
rect 1020 -1250 1124 -1237
rect 1180 -1013 1284 -1000
rect 1180 -1237 1209 -1013
rect 1255 -1237 1284 -1013
rect 1180 -1250 1284 -1237
rect 1340 -1013 1444 -1000
rect 1340 -1237 1369 -1013
rect 1415 -1237 1444 -1013
rect 1340 -1250 1444 -1237
rect 1500 -1013 1604 -1000
rect 1500 -1237 1529 -1013
rect 1575 -1237 1604 -1013
rect 1500 -1250 1604 -1237
rect 1660 -1013 1748 -1000
rect 1660 -1237 1689 -1013
rect 1735 -1237 1748 -1013
rect 1660 -1250 1748 -1237
rect 1920 -1013 2008 -1000
rect 1920 -1237 1933 -1013
rect 1979 -1237 2008 -1013
rect 1920 -1250 2008 -1237
rect 2064 -1013 2168 -1000
rect 2064 -1237 2093 -1013
rect 2139 -1237 2168 -1013
rect 2064 -1250 2168 -1237
rect 2224 -1013 2328 -1000
rect 2224 -1237 2253 -1013
rect 2299 -1237 2328 -1013
rect 2224 -1250 2328 -1237
rect 2384 -1013 2488 -1000
rect 2384 -1237 2413 -1013
rect 2459 -1237 2488 -1013
rect 2384 -1250 2488 -1237
rect 2544 -1013 2648 -1000
rect 2544 -1237 2573 -1013
rect 2619 -1237 2648 -1013
rect 2544 -1250 2648 -1237
rect 2704 -1013 2808 -1000
rect 2704 -1237 2733 -1013
rect 2779 -1237 2808 -1013
rect 2704 -1250 2808 -1237
rect 2864 -1013 2968 -1000
rect 2864 -1237 2893 -1013
rect 2939 -1237 2968 -1013
rect 2864 -1250 2968 -1237
rect 3024 -1013 3128 -1000
rect 3024 -1237 3053 -1013
rect 3099 -1237 3128 -1013
rect 3024 -1250 3128 -1237
rect 3184 -1013 3272 -1000
rect 3184 -1237 3213 -1013
rect 3259 -1237 3272 -1013
rect 3184 -1250 3272 -1237
rect 3328 -1013 3416 -1000
rect 3328 -1237 3341 -1013
rect 3387 -1237 3416 -1013
rect 3328 -1250 3416 -1237
rect 3472 -1013 3560 -1000
rect 3472 -1237 3501 -1013
rect 3547 -1237 3560 -1013
rect 3472 -1250 3560 -1237
rect 3732 -1013 3820 -1000
rect 3732 -1237 3745 -1013
rect 3791 -1237 3820 -1013
rect 3732 -1250 3820 -1237
rect 3876 -1013 3964 -1000
rect 3876 -1237 3905 -1013
rect 3951 -1237 3964 -1013
rect 3876 -1250 3964 -1237
rect 4020 -1013 4108 -1000
rect 4020 -1237 4033 -1013
rect 4079 -1237 4108 -1013
rect 4020 -1250 4108 -1237
rect 4164 -1013 4268 -1000
rect 4164 -1237 4193 -1013
rect 4239 -1237 4268 -1013
rect 4164 -1250 4268 -1237
rect 4324 -1013 4428 -1000
rect 4324 -1237 4353 -1013
rect 4399 -1237 4428 -1013
rect 4324 -1250 4428 -1237
rect 4484 -1013 4588 -1000
rect 4484 -1237 4513 -1013
rect 4559 -1237 4588 -1013
rect 4484 -1250 4588 -1237
rect 4644 -1013 4748 -1000
rect 4644 -1237 4673 -1013
rect 4719 -1237 4748 -1013
rect 4644 -1250 4748 -1237
rect 4804 -1013 4908 -1000
rect 4804 -1237 4833 -1013
rect 4879 -1237 4908 -1013
rect 4804 -1250 4908 -1237
rect 4964 -1013 5068 -1000
rect 4964 -1237 4993 -1013
rect 5039 -1237 5068 -1013
rect 4964 -1250 5068 -1237
rect 5124 -1013 5228 -1000
rect 5124 -1237 5153 -1013
rect 5199 -1237 5228 -1013
rect 5124 -1250 5228 -1237
rect 5284 -1013 5372 -1000
rect 5284 -1237 5313 -1013
rect 5359 -1237 5372 -1013
rect 5284 -1250 5372 -1237
rect 5544 -1013 5632 -1000
rect 5544 -1237 5557 -1013
rect 5603 -1237 5632 -1013
rect 5544 -1250 5632 -1237
rect 5688 -1013 5792 -1000
rect 5688 -1237 5717 -1013
rect 5763 -1237 5792 -1013
rect 5688 -1250 5792 -1237
rect 5848 -1013 5952 -1000
rect 5848 -1237 5877 -1013
rect 5923 -1237 5952 -1013
rect 5848 -1250 5952 -1237
rect 6008 -1013 6112 -1000
rect 6008 -1237 6037 -1013
rect 6083 -1237 6112 -1013
rect 6008 -1250 6112 -1237
rect 6168 -1013 6272 -1000
rect 6168 -1237 6197 -1013
rect 6243 -1237 6272 -1013
rect 6168 -1250 6272 -1237
rect 6328 -1013 6432 -1000
rect 6328 -1237 6357 -1013
rect 6403 -1237 6432 -1013
rect 6328 -1250 6432 -1237
rect 6488 -1013 6592 -1000
rect 6488 -1237 6517 -1013
rect 6563 -1237 6592 -1013
rect 6488 -1250 6592 -1237
rect 6648 -1013 6752 -1000
rect 6648 -1237 6677 -1013
rect 6723 -1237 6752 -1013
rect 6648 -1250 6752 -1237
rect 6808 -1013 6896 -1000
rect 6808 -1237 6837 -1013
rect 6883 -1237 6896 -1013
rect 6808 -1250 6896 -1237
rect 6952 -1013 7040 -1000
rect 6952 -1237 6965 -1013
rect 7011 -1237 7040 -1013
rect 6952 -1250 7040 -1237
rect 7096 -1013 7184 -1000
rect 7096 -1237 7125 -1013
rect 7171 -1237 7184 -1013
rect 7096 -1250 7184 -1237
rect 7356 -1013 7444 -1000
rect 7356 -1237 7369 -1013
rect 7415 -1237 7444 -1013
rect 7356 -1250 7444 -1237
rect 7500 -1013 7604 -1000
rect 7500 -1237 7529 -1013
rect 7575 -1237 7604 -1013
rect 7500 -1250 7604 -1237
rect 7660 -1013 7764 -1000
rect 7660 -1237 7689 -1013
rect 7735 -1237 7764 -1013
rect 7660 -1250 7764 -1237
rect 7820 -1013 7924 -1000
rect 7820 -1237 7849 -1013
rect 7895 -1237 7924 -1013
rect 7820 -1250 7924 -1237
rect 7980 -1013 8084 -1000
rect 7980 -1237 8009 -1013
rect 8055 -1237 8084 -1013
rect 7980 -1250 8084 -1237
rect 8140 -1013 8244 -1000
rect 8140 -1237 8169 -1013
rect 8215 -1237 8244 -1013
rect 8140 -1250 8244 -1237
rect 8300 -1013 8404 -1000
rect 8300 -1237 8329 -1013
rect 8375 -1237 8404 -1013
rect 8300 -1250 8404 -1237
rect 8460 -1013 8564 -1000
rect 8460 -1237 8489 -1013
rect 8535 -1237 8564 -1013
rect 8460 -1250 8564 -1237
rect 8620 -1013 8708 -1000
rect 8620 -1237 8649 -1013
rect 8695 -1237 8708 -1013
rect 8620 -1250 8708 -1237
rect 8764 -1013 8852 -1000
rect 8764 -1237 8777 -1013
rect 8823 -1237 8852 -1013
rect 8764 -1250 8852 -1237
rect 8908 -1013 8996 -1000
rect 8908 -1237 8937 -1013
rect 8983 -1237 8996 -1013
rect 8908 -1250 8996 -1237
rect -4089 -5979 -4001 -5966
rect -4089 -6203 -4076 -5979
rect -4030 -6203 -4001 -5979
rect -4089 -6216 -4001 -6203
rect -3945 -5979 -3857 -5966
rect -3945 -6203 -3916 -5979
rect -3870 -6203 -3857 -5979
rect -3945 -6216 -3857 -6203
rect -3801 -5979 -3713 -5966
rect -3801 -6203 -3788 -5979
rect -3742 -6203 -3713 -5979
rect -3801 -6216 -3713 -6203
rect -3657 -5979 -3553 -5966
rect -3657 -6203 -3628 -5979
rect -3582 -6203 -3553 -5979
rect -3657 -6216 -3553 -6203
rect -3497 -5979 -3393 -5966
rect -3497 -6203 -3468 -5979
rect -3422 -6203 -3393 -5979
rect -3497 -6216 -3393 -6203
rect -3337 -5979 -3233 -5966
rect -3337 -6203 -3308 -5979
rect -3262 -6203 -3233 -5979
rect -3337 -6216 -3233 -6203
rect -3177 -5979 -3073 -5966
rect -3177 -6203 -3148 -5979
rect -3102 -6203 -3073 -5979
rect -3177 -6216 -3073 -6203
rect -3017 -5979 -2913 -5966
rect -3017 -6203 -2988 -5979
rect -2942 -6203 -2913 -5979
rect -3017 -6216 -2913 -6203
rect -2857 -5979 -2753 -5966
rect -2857 -6203 -2828 -5979
rect -2782 -6203 -2753 -5979
rect -2857 -6216 -2753 -6203
rect -2697 -5979 -2593 -5966
rect -2697 -6203 -2668 -5979
rect -2622 -6203 -2593 -5979
rect -2697 -6216 -2593 -6203
rect -2537 -5979 -2449 -5966
rect -2537 -6203 -2508 -5979
rect -2462 -6203 -2449 -5979
rect -2537 -6216 -2449 -6203
rect -2277 -5979 -2189 -5966
rect -2277 -6203 -2264 -5979
rect -2218 -6203 -2189 -5979
rect -2277 -6216 -2189 -6203
rect -2133 -5979 -2029 -5966
rect -2133 -6203 -2104 -5979
rect -2058 -6203 -2029 -5979
rect -2133 -6216 -2029 -6203
rect -1973 -5979 -1869 -5966
rect -1973 -6203 -1944 -5979
rect -1898 -6203 -1869 -5979
rect -1973 -6216 -1869 -6203
rect -1813 -5979 -1709 -5966
rect -1813 -6203 -1784 -5979
rect -1738 -6203 -1709 -5979
rect -1813 -6216 -1709 -6203
rect -1653 -5979 -1549 -5966
rect -1653 -6203 -1624 -5979
rect -1578 -6203 -1549 -5979
rect -1653 -6216 -1549 -6203
rect -1493 -5979 -1389 -5966
rect -1493 -6203 -1464 -5979
rect -1418 -6203 -1389 -5979
rect -1493 -6216 -1389 -6203
rect -1333 -5979 -1229 -5966
rect -1333 -6203 -1304 -5979
rect -1258 -6203 -1229 -5979
rect -1333 -6216 -1229 -6203
rect -1173 -5979 -1069 -5966
rect -1173 -6203 -1144 -5979
rect -1098 -6203 -1069 -5979
rect -1173 -6216 -1069 -6203
rect -1013 -5979 -925 -5966
rect -1013 -6203 -984 -5979
rect -938 -6203 -925 -5979
rect -1013 -6216 -925 -6203
rect -869 -5979 -781 -5966
rect -869 -6203 -856 -5979
rect -810 -6203 -781 -5979
rect -869 -6216 -781 -6203
rect -725 -5979 -637 -5966
rect -725 -6203 -696 -5979
rect -650 -6203 -637 -5979
rect -725 -6216 -637 -6203
rect 108 -5979 196 -5966
rect 108 -6203 121 -5979
rect 167 -6203 196 -5979
rect 108 -6216 196 -6203
rect 252 -5979 340 -5966
rect 252 -6203 281 -5979
rect 327 -6203 340 -5979
rect 252 -6216 340 -6203
rect 396 -5979 484 -5966
rect 396 -6203 409 -5979
rect 455 -6203 484 -5979
rect 396 -6216 484 -6203
rect 540 -5979 644 -5966
rect 540 -6203 569 -5979
rect 615 -6203 644 -5979
rect 540 -6216 644 -6203
rect 700 -5979 804 -5966
rect 700 -6203 729 -5979
rect 775 -6203 804 -5979
rect 700 -6216 804 -6203
rect 860 -5979 964 -5966
rect 860 -6203 889 -5979
rect 935 -6203 964 -5979
rect 860 -6216 964 -6203
rect 1020 -5979 1124 -5966
rect 1020 -6203 1049 -5979
rect 1095 -6203 1124 -5979
rect 1020 -6216 1124 -6203
rect 1180 -5979 1284 -5966
rect 1180 -6203 1209 -5979
rect 1255 -6203 1284 -5979
rect 1180 -6216 1284 -6203
rect 1340 -5979 1444 -5966
rect 1340 -6203 1369 -5979
rect 1415 -6203 1444 -5979
rect 1340 -6216 1444 -6203
rect 1500 -5979 1604 -5966
rect 1500 -6203 1529 -5979
rect 1575 -6203 1604 -5979
rect 1500 -6216 1604 -6203
rect 1660 -5979 1748 -5966
rect 1660 -6203 1689 -5979
rect 1735 -6203 1748 -5979
rect 1660 -6216 1748 -6203
rect 1920 -5979 2008 -5966
rect 1920 -6203 1933 -5979
rect 1979 -6203 2008 -5979
rect 1920 -6216 2008 -6203
rect 2064 -5979 2168 -5966
rect 2064 -6203 2093 -5979
rect 2139 -6203 2168 -5979
rect 2064 -6216 2168 -6203
rect 2224 -5979 2328 -5966
rect 2224 -6203 2253 -5979
rect 2299 -6203 2328 -5979
rect 2224 -6216 2328 -6203
rect 2384 -5979 2488 -5966
rect 2384 -6203 2413 -5979
rect 2459 -6203 2488 -5979
rect 2384 -6216 2488 -6203
rect 2544 -5979 2648 -5966
rect 2544 -6203 2573 -5979
rect 2619 -6203 2648 -5979
rect 2544 -6216 2648 -6203
rect 2704 -5979 2808 -5966
rect 2704 -6203 2733 -5979
rect 2779 -6203 2808 -5979
rect 2704 -6216 2808 -6203
rect 2864 -5979 2968 -5966
rect 2864 -6203 2893 -5979
rect 2939 -6203 2968 -5979
rect 2864 -6216 2968 -6203
rect 3024 -5979 3128 -5966
rect 3024 -6203 3053 -5979
rect 3099 -6203 3128 -5979
rect 3024 -6216 3128 -6203
rect 3184 -5979 3272 -5966
rect 3184 -6203 3213 -5979
rect 3259 -6203 3272 -5979
rect 3184 -6216 3272 -6203
rect 3328 -5979 3416 -5966
rect 3328 -6203 3341 -5979
rect 3387 -6203 3416 -5979
rect 3328 -6216 3416 -6203
rect 3472 -5979 3560 -5966
rect 3472 -6203 3501 -5979
rect 3547 -6203 3560 -5979
rect 3472 -6216 3560 -6203
rect 3732 -5979 3820 -5966
rect 3732 -6203 3745 -5979
rect 3791 -6203 3820 -5979
rect 3732 -6216 3820 -6203
rect 3876 -5979 3964 -5966
rect 3876 -6203 3905 -5979
rect 3951 -6203 3964 -5979
rect 3876 -6216 3964 -6203
rect 4020 -5979 4108 -5966
rect 4020 -6203 4033 -5979
rect 4079 -6203 4108 -5979
rect 4020 -6216 4108 -6203
rect 4164 -5979 4268 -5966
rect 4164 -6203 4193 -5979
rect 4239 -6203 4268 -5979
rect 4164 -6216 4268 -6203
rect 4324 -5979 4428 -5966
rect 4324 -6203 4353 -5979
rect 4399 -6203 4428 -5979
rect 4324 -6216 4428 -6203
rect 4484 -5979 4588 -5966
rect 4484 -6203 4513 -5979
rect 4559 -6203 4588 -5979
rect 4484 -6216 4588 -6203
rect 4644 -5979 4748 -5966
rect 4644 -6203 4673 -5979
rect 4719 -6203 4748 -5979
rect 4644 -6216 4748 -6203
rect 4804 -5979 4908 -5966
rect 4804 -6203 4833 -5979
rect 4879 -6203 4908 -5979
rect 4804 -6216 4908 -6203
rect 4964 -5979 5068 -5966
rect 4964 -6203 4993 -5979
rect 5039 -6203 5068 -5979
rect 4964 -6216 5068 -6203
rect 5124 -5979 5228 -5966
rect 5124 -6203 5153 -5979
rect 5199 -6203 5228 -5979
rect 5124 -6216 5228 -6203
rect 5284 -5979 5372 -5966
rect 5284 -6203 5313 -5979
rect 5359 -6203 5372 -5979
rect 5284 -6216 5372 -6203
rect 5544 -5979 5632 -5966
rect 5544 -6203 5557 -5979
rect 5603 -6203 5632 -5979
rect 5544 -6216 5632 -6203
rect 5688 -5979 5792 -5966
rect 5688 -6203 5717 -5979
rect 5763 -6203 5792 -5979
rect 5688 -6216 5792 -6203
rect 5848 -5979 5952 -5966
rect 5848 -6203 5877 -5979
rect 5923 -6203 5952 -5979
rect 5848 -6216 5952 -6203
rect 6008 -5979 6112 -5966
rect 6008 -6203 6037 -5979
rect 6083 -6203 6112 -5979
rect 6008 -6216 6112 -6203
rect 6168 -5979 6272 -5966
rect 6168 -6203 6197 -5979
rect 6243 -6203 6272 -5979
rect 6168 -6216 6272 -6203
rect 6328 -5979 6432 -5966
rect 6328 -6203 6357 -5979
rect 6403 -6203 6432 -5979
rect 6328 -6216 6432 -6203
rect 6488 -5979 6592 -5966
rect 6488 -6203 6517 -5979
rect 6563 -6203 6592 -5979
rect 6488 -6216 6592 -6203
rect 6648 -5979 6752 -5966
rect 6648 -6203 6677 -5979
rect 6723 -6203 6752 -5979
rect 6648 -6216 6752 -6203
rect 6808 -5979 6896 -5966
rect 6808 -6203 6837 -5979
rect 6883 -6203 6896 -5979
rect 6808 -6216 6896 -6203
rect 6952 -5979 7040 -5966
rect 6952 -6203 6965 -5979
rect 7011 -6203 7040 -5979
rect 6952 -6216 7040 -6203
rect 7096 -5979 7184 -5966
rect 7096 -6203 7125 -5979
rect 7171 -6203 7184 -5979
rect 7096 -6216 7184 -6203
rect 7356 -5979 7444 -5966
rect 7356 -6203 7369 -5979
rect 7415 -6203 7444 -5979
rect 7356 -6216 7444 -6203
rect 7500 -5979 7604 -5966
rect 7500 -6203 7529 -5979
rect 7575 -6203 7604 -5979
rect 7500 -6216 7604 -6203
rect 7660 -5979 7764 -5966
rect 7660 -6203 7689 -5979
rect 7735 -6203 7764 -5979
rect 7660 -6216 7764 -6203
rect 7820 -5979 7924 -5966
rect 7820 -6203 7849 -5979
rect 7895 -6203 7924 -5979
rect 7820 -6216 7924 -6203
rect 7980 -5979 8084 -5966
rect 7980 -6203 8009 -5979
rect 8055 -6203 8084 -5979
rect 7980 -6216 8084 -6203
rect 8140 -5979 8244 -5966
rect 8140 -6203 8169 -5979
rect 8215 -6203 8244 -5979
rect 8140 -6216 8244 -6203
rect 8300 -5979 8404 -5966
rect 8300 -6203 8329 -5979
rect 8375 -6203 8404 -5979
rect 8300 -6216 8404 -6203
rect 8460 -5979 8564 -5966
rect 8460 -6203 8489 -5979
rect 8535 -6203 8564 -5979
rect 8460 -6216 8564 -6203
rect 8620 -5979 8708 -5966
rect 8620 -6203 8649 -5979
rect 8695 -6203 8708 -5979
rect 8620 -6216 8708 -6203
rect 8764 -5979 8852 -5966
rect 8764 -6203 8777 -5979
rect 8823 -6203 8852 -5979
rect 8764 -6216 8852 -6203
rect 8908 -5979 8996 -5966
rect 8908 -6203 8937 -5979
rect 8983 -6203 8996 -5979
rect 8908 -6216 8996 -6203
rect -4089 -6365 -4001 -6352
rect -4089 -6589 -4076 -6365
rect -4030 -6589 -4001 -6365
rect -4089 -6602 -4001 -6589
rect -3945 -6365 -3857 -6352
rect -3945 -6589 -3916 -6365
rect -3870 -6589 -3857 -6365
rect -3945 -6602 -3857 -6589
rect -3801 -6365 -3713 -6352
rect -3801 -6589 -3788 -6365
rect -3742 -6589 -3713 -6365
rect -3801 -6602 -3713 -6589
rect -3657 -6365 -3553 -6352
rect -3657 -6589 -3628 -6365
rect -3582 -6589 -3553 -6365
rect -3657 -6602 -3553 -6589
rect -3497 -6365 -3393 -6352
rect -3497 -6589 -3468 -6365
rect -3422 -6589 -3393 -6365
rect -3497 -6602 -3393 -6589
rect -3337 -6365 -3233 -6352
rect -3337 -6589 -3308 -6365
rect -3262 -6589 -3233 -6365
rect -3337 -6602 -3233 -6589
rect -3177 -6365 -3073 -6352
rect -3177 -6589 -3148 -6365
rect -3102 -6589 -3073 -6365
rect -3177 -6602 -3073 -6589
rect -3017 -6365 -2913 -6352
rect -3017 -6589 -2988 -6365
rect -2942 -6589 -2913 -6365
rect -3017 -6602 -2913 -6589
rect -2857 -6365 -2753 -6352
rect -2857 -6589 -2828 -6365
rect -2782 -6589 -2753 -6365
rect -2857 -6602 -2753 -6589
rect -2697 -6365 -2593 -6352
rect -2697 -6589 -2668 -6365
rect -2622 -6589 -2593 -6365
rect -2697 -6602 -2593 -6589
rect -2537 -6365 -2449 -6352
rect -2537 -6589 -2508 -6365
rect -2462 -6589 -2449 -6365
rect -2537 -6602 -2449 -6589
rect -2277 -6365 -2189 -6352
rect -2277 -6589 -2264 -6365
rect -2218 -6589 -2189 -6365
rect -2277 -6602 -2189 -6589
rect -2133 -6365 -2029 -6352
rect -2133 -6589 -2104 -6365
rect -2058 -6589 -2029 -6365
rect -2133 -6602 -2029 -6589
rect -1973 -6365 -1869 -6352
rect -1973 -6589 -1944 -6365
rect -1898 -6589 -1869 -6365
rect -1973 -6602 -1869 -6589
rect -1813 -6365 -1709 -6352
rect -1813 -6589 -1784 -6365
rect -1738 -6589 -1709 -6365
rect -1813 -6602 -1709 -6589
rect -1653 -6365 -1549 -6352
rect -1653 -6589 -1624 -6365
rect -1578 -6589 -1549 -6365
rect -1653 -6602 -1549 -6589
rect -1493 -6365 -1389 -6352
rect -1493 -6589 -1464 -6365
rect -1418 -6589 -1389 -6365
rect -1493 -6602 -1389 -6589
rect -1333 -6365 -1229 -6352
rect -1333 -6589 -1304 -6365
rect -1258 -6589 -1229 -6365
rect -1333 -6602 -1229 -6589
rect -1173 -6365 -1069 -6352
rect -1173 -6589 -1144 -6365
rect -1098 -6589 -1069 -6365
rect -1173 -6602 -1069 -6589
rect -1013 -6365 -925 -6352
rect -1013 -6589 -984 -6365
rect -938 -6589 -925 -6365
rect -1013 -6602 -925 -6589
rect -869 -6365 -781 -6352
rect -869 -6589 -856 -6365
rect -810 -6589 -781 -6365
rect -869 -6602 -781 -6589
rect -725 -6365 -637 -6352
rect -725 -6589 -696 -6365
rect -650 -6589 -637 -6365
rect -725 -6602 -637 -6589
rect 108 -6365 196 -6352
rect 108 -6589 121 -6365
rect 167 -6589 196 -6365
rect 108 -6602 196 -6589
rect 252 -6365 340 -6352
rect 252 -6589 281 -6365
rect 327 -6589 340 -6365
rect 252 -6602 340 -6589
rect 396 -6365 484 -6352
rect 396 -6589 409 -6365
rect 455 -6589 484 -6365
rect 396 -6602 484 -6589
rect 540 -6365 644 -6352
rect 540 -6589 569 -6365
rect 615 -6589 644 -6365
rect 540 -6602 644 -6589
rect 700 -6365 804 -6352
rect 700 -6589 729 -6365
rect 775 -6589 804 -6365
rect 700 -6602 804 -6589
rect 860 -6365 964 -6352
rect 860 -6589 889 -6365
rect 935 -6589 964 -6365
rect 860 -6602 964 -6589
rect 1020 -6365 1124 -6352
rect 1020 -6589 1049 -6365
rect 1095 -6589 1124 -6365
rect 1020 -6602 1124 -6589
rect 1180 -6365 1284 -6352
rect 1180 -6589 1209 -6365
rect 1255 -6589 1284 -6365
rect 1180 -6602 1284 -6589
rect 1340 -6365 1444 -6352
rect 1340 -6589 1369 -6365
rect 1415 -6589 1444 -6365
rect 1340 -6602 1444 -6589
rect 1500 -6365 1604 -6352
rect 1500 -6589 1529 -6365
rect 1575 -6589 1604 -6365
rect 1500 -6602 1604 -6589
rect 1660 -6365 1748 -6352
rect 1660 -6589 1689 -6365
rect 1735 -6589 1748 -6365
rect 1660 -6602 1748 -6589
rect 1920 -6365 2008 -6352
rect 1920 -6589 1933 -6365
rect 1979 -6589 2008 -6365
rect 1920 -6602 2008 -6589
rect 2064 -6365 2168 -6352
rect 2064 -6589 2093 -6365
rect 2139 -6589 2168 -6365
rect 2064 -6602 2168 -6589
rect 2224 -6365 2328 -6352
rect 2224 -6589 2253 -6365
rect 2299 -6589 2328 -6365
rect 2224 -6602 2328 -6589
rect 2384 -6365 2488 -6352
rect 2384 -6589 2413 -6365
rect 2459 -6589 2488 -6365
rect 2384 -6602 2488 -6589
rect 2544 -6365 2648 -6352
rect 2544 -6589 2573 -6365
rect 2619 -6589 2648 -6365
rect 2544 -6602 2648 -6589
rect 2704 -6365 2808 -6352
rect 2704 -6589 2733 -6365
rect 2779 -6589 2808 -6365
rect 2704 -6602 2808 -6589
rect 2864 -6365 2968 -6352
rect 2864 -6589 2893 -6365
rect 2939 -6589 2968 -6365
rect 2864 -6602 2968 -6589
rect 3024 -6365 3128 -6352
rect 3024 -6589 3053 -6365
rect 3099 -6589 3128 -6365
rect 3024 -6602 3128 -6589
rect 3184 -6365 3272 -6352
rect 3184 -6589 3213 -6365
rect 3259 -6589 3272 -6365
rect 3184 -6602 3272 -6589
rect 3328 -6365 3416 -6352
rect 3328 -6589 3341 -6365
rect 3387 -6589 3416 -6365
rect 3328 -6602 3416 -6589
rect 3472 -6365 3560 -6352
rect 3472 -6589 3501 -6365
rect 3547 -6589 3560 -6365
rect 3472 -6602 3560 -6589
rect 3732 -6365 3820 -6352
rect 3732 -6589 3745 -6365
rect 3791 -6589 3820 -6365
rect 3732 -6602 3820 -6589
rect 3876 -6365 3964 -6352
rect 3876 -6589 3905 -6365
rect 3951 -6589 3964 -6365
rect 3876 -6602 3964 -6589
rect 4020 -6365 4108 -6352
rect 4020 -6589 4033 -6365
rect 4079 -6589 4108 -6365
rect 4020 -6602 4108 -6589
rect 4164 -6365 4268 -6352
rect 4164 -6589 4193 -6365
rect 4239 -6589 4268 -6365
rect 4164 -6602 4268 -6589
rect 4324 -6365 4428 -6352
rect 4324 -6589 4353 -6365
rect 4399 -6589 4428 -6365
rect 4324 -6602 4428 -6589
rect 4484 -6365 4588 -6352
rect 4484 -6589 4513 -6365
rect 4559 -6589 4588 -6365
rect 4484 -6602 4588 -6589
rect 4644 -6365 4748 -6352
rect 4644 -6589 4673 -6365
rect 4719 -6589 4748 -6365
rect 4644 -6602 4748 -6589
rect 4804 -6365 4908 -6352
rect 4804 -6589 4833 -6365
rect 4879 -6589 4908 -6365
rect 4804 -6602 4908 -6589
rect 4964 -6365 5068 -6352
rect 4964 -6589 4993 -6365
rect 5039 -6589 5068 -6365
rect 4964 -6602 5068 -6589
rect 5124 -6365 5228 -6352
rect 5124 -6589 5153 -6365
rect 5199 -6589 5228 -6365
rect 5124 -6602 5228 -6589
rect 5284 -6365 5372 -6352
rect 5284 -6589 5313 -6365
rect 5359 -6589 5372 -6365
rect 5284 -6602 5372 -6589
rect 5544 -6365 5632 -6352
rect 5544 -6589 5557 -6365
rect 5603 -6589 5632 -6365
rect 5544 -6602 5632 -6589
rect 5688 -6365 5792 -6352
rect 5688 -6589 5717 -6365
rect 5763 -6589 5792 -6365
rect 5688 -6602 5792 -6589
rect 5848 -6365 5952 -6352
rect 5848 -6589 5877 -6365
rect 5923 -6589 5952 -6365
rect 5848 -6602 5952 -6589
rect 6008 -6365 6112 -6352
rect 6008 -6589 6037 -6365
rect 6083 -6589 6112 -6365
rect 6008 -6602 6112 -6589
rect 6168 -6365 6272 -6352
rect 6168 -6589 6197 -6365
rect 6243 -6589 6272 -6365
rect 6168 -6602 6272 -6589
rect 6328 -6365 6432 -6352
rect 6328 -6589 6357 -6365
rect 6403 -6589 6432 -6365
rect 6328 -6602 6432 -6589
rect 6488 -6365 6592 -6352
rect 6488 -6589 6517 -6365
rect 6563 -6589 6592 -6365
rect 6488 -6602 6592 -6589
rect 6648 -6365 6752 -6352
rect 6648 -6589 6677 -6365
rect 6723 -6589 6752 -6365
rect 6648 -6602 6752 -6589
rect 6808 -6365 6896 -6352
rect 6808 -6589 6837 -6365
rect 6883 -6589 6896 -6365
rect 6808 -6602 6896 -6589
rect 6952 -6365 7040 -6352
rect 6952 -6589 6965 -6365
rect 7011 -6589 7040 -6365
rect 6952 -6602 7040 -6589
rect 7096 -6365 7184 -6352
rect 7096 -6589 7125 -6365
rect 7171 -6589 7184 -6365
rect 7096 -6602 7184 -6589
rect 7356 -6365 7444 -6352
rect 7356 -6589 7369 -6365
rect 7415 -6589 7444 -6365
rect 7356 -6602 7444 -6589
rect 7500 -6365 7604 -6352
rect 7500 -6589 7529 -6365
rect 7575 -6589 7604 -6365
rect 7500 -6602 7604 -6589
rect 7660 -6365 7764 -6352
rect 7660 -6589 7689 -6365
rect 7735 -6589 7764 -6365
rect 7660 -6602 7764 -6589
rect 7820 -6365 7924 -6352
rect 7820 -6589 7849 -6365
rect 7895 -6589 7924 -6365
rect 7820 -6602 7924 -6589
rect 7980 -6365 8084 -6352
rect 7980 -6589 8009 -6365
rect 8055 -6589 8084 -6365
rect 7980 -6602 8084 -6589
rect 8140 -6365 8244 -6352
rect 8140 -6589 8169 -6365
rect 8215 -6589 8244 -6365
rect 8140 -6602 8244 -6589
rect 8300 -6365 8404 -6352
rect 8300 -6589 8329 -6365
rect 8375 -6589 8404 -6365
rect 8300 -6602 8404 -6589
rect 8460 -6365 8564 -6352
rect 8460 -6589 8489 -6365
rect 8535 -6589 8564 -6365
rect 8460 -6602 8564 -6589
rect 8620 -6365 8708 -6352
rect 8620 -6589 8649 -6365
rect 8695 -6589 8708 -6365
rect 8620 -6602 8708 -6589
rect 8764 -6365 8852 -6352
rect 8764 -6589 8777 -6365
rect 8823 -6589 8852 -6365
rect 8764 -6602 8852 -6589
rect 8908 -6365 8996 -6352
rect 8908 -6589 8937 -6365
rect 8983 -6589 8996 -6365
rect 8908 -6602 8996 -6589
rect -4089 -6751 -4001 -6738
rect -4089 -6975 -4076 -6751
rect -4030 -6975 -4001 -6751
rect -4089 -6988 -4001 -6975
rect -3945 -6751 -3857 -6738
rect -3945 -6975 -3916 -6751
rect -3870 -6975 -3857 -6751
rect -3945 -6988 -3857 -6975
rect -3801 -6751 -3713 -6738
rect -3801 -6975 -3788 -6751
rect -3742 -6975 -3713 -6751
rect -3801 -6988 -3713 -6975
rect -3657 -6751 -3553 -6738
rect -3657 -6975 -3628 -6751
rect -3582 -6975 -3553 -6751
rect -3657 -6988 -3553 -6975
rect -3497 -6751 -3393 -6738
rect -3497 -6975 -3468 -6751
rect -3422 -6975 -3393 -6751
rect -3497 -6988 -3393 -6975
rect -3337 -6751 -3233 -6738
rect -3337 -6975 -3308 -6751
rect -3262 -6975 -3233 -6751
rect -3337 -6988 -3233 -6975
rect -3177 -6751 -3073 -6738
rect -3177 -6975 -3148 -6751
rect -3102 -6975 -3073 -6751
rect -3177 -6988 -3073 -6975
rect -3017 -6751 -2913 -6738
rect -3017 -6975 -2988 -6751
rect -2942 -6975 -2913 -6751
rect -3017 -6988 -2913 -6975
rect -2857 -6751 -2753 -6738
rect -2857 -6975 -2828 -6751
rect -2782 -6975 -2753 -6751
rect -2857 -6988 -2753 -6975
rect -2697 -6751 -2593 -6738
rect -2697 -6975 -2668 -6751
rect -2622 -6975 -2593 -6751
rect -2697 -6988 -2593 -6975
rect -2537 -6751 -2449 -6738
rect -2537 -6975 -2508 -6751
rect -2462 -6975 -2449 -6751
rect -2537 -6988 -2449 -6975
rect -2277 -6751 -2189 -6738
rect -2277 -6975 -2264 -6751
rect -2218 -6975 -2189 -6751
rect -2277 -6988 -2189 -6975
rect -2133 -6751 -2029 -6738
rect -2133 -6975 -2104 -6751
rect -2058 -6975 -2029 -6751
rect -2133 -6988 -2029 -6975
rect -1973 -6751 -1869 -6738
rect -1973 -6975 -1944 -6751
rect -1898 -6975 -1869 -6751
rect -1973 -6988 -1869 -6975
rect -1813 -6751 -1709 -6738
rect -1813 -6975 -1784 -6751
rect -1738 -6975 -1709 -6751
rect -1813 -6988 -1709 -6975
rect -1653 -6751 -1549 -6738
rect -1653 -6975 -1624 -6751
rect -1578 -6975 -1549 -6751
rect -1653 -6988 -1549 -6975
rect -1493 -6751 -1389 -6738
rect -1493 -6975 -1464 -6751
rect -1418 -6975 -1389 -6751
rect -1493 -6988 -1389 -6975
rect -1333 -6751 -1229 -6738
rect -1333 -6975 -1304 -6751
rect -1258 -6975 -1229 -6751
rect -1333 -6988 -1229 -6975
rect -1173 -6751 -1069 -6738
rect -1173 -6975 -1144 -6751
rect -1098 -6975 -1069 -6751
rect -1173 -6988 -1069 -6975
rect -1013 -6751 -925 -6738
rect -1013 -6975 -984 -6751
rect -938 -6975 -925 -6751
rect -1013 -6988 -925 -6975
rect -869 -6751 -781 -6738
rect -869 -6975 -856 -6751
rect -810 -6975 -781 -6751
rect -869 -6988 -781 -6975
rect -725 -6751 -637 -6738
rect -725 -6975 -696 -6751
rect -650 -6975 -637 -6751
rect -725 -6988 -637 -6975
rect 108 -6751 196 -6738
rect 108 -6975 121 -6751
rect 167 -6975 196 -6751
rect 108 -6988 196 -6975
rect 252 -6751 340 -6738
rect 252 -6975 281 -6751
rect 327 -6975 340 -6751
rect 252 -6988 340 -6975
rect 396 -6751 484 -6738
rect 396 -6975 409 -6751
rect 455 -6975 484 -6751
rect 396 -6988 484 -6975
rect 540 -6751 644 -6738
rect 540 -6975 569 -6751
rect 615 -6975 644 -6751
rect 540 -6988 644 -6975
rect 700 -6751 804 -6738
rect 700 -6975 729 -6751
rect 775 -6975 804 -6751
rect 700 -6988 804 -6975
rect 860 -6751 964 -6738
rect 860 -6975 889 -6751
rect 935 -6975 964 -6751
rect 860 -6988 964 -6975
rect 1020 -6751 1124 -6738
rect 1020 -6975 1049 -6751
rect 1095 -6975 1124 -6751
rect 1020 -6988 1124 -6975
rect 1180 -6751 1284 -6738
rect 1180 -6975 1209 -6751
rect 1255 -6975 1284 -6751
rect 1180 -6988 1284 -6975
rect 1340 -6751 1444 -6738
rect 1340 -6975 1369 -6751
rect 1415 -6975 1444 -6751
rect 1340 -6988 1444 -6975
rect 1500 -6751 1604 -6738
rect 1500 -6975 1529 -6751
rect 1575 -6975 1604 -6751
rect 1500 -6988 1604 -6975
rect 1660 -6751 1748 -6738
rect 1660 -6975 1689 -6751
rect 1735 -6975 1748 -6751
rect 1660 -6988 1748 -6975
rect 1920 -6751 2008 -6738
rect 1920 -6975 1933 -6751
rect 1979 -6975 2008 -6751
rect 1920 -6988 2008 -6975
rect 2064 -6751 2168 -6738
rect 2064 -6975 2093 -6751
rect 2139 -6975 2168 -6751
rect 2064 -6988 2168 -6975
rect 2224 -6751 2328 -6738
rect 2224 -6975 2253 -6751
rect 2299 -6975 2328 -6751
rect 2224 -6988 2328 -6975
rect 2384 -6751 2488 -6738
rect 2384 -6975 2413 -6751
rect 2459 -6975 2488 -6751
rect 2384 -6988 2488 -6975
rect 2544 -6751 2648 -6738
rect 2544 -6975 2573 -6751
rect 2619 -6975 2648 -6751
rect 2544 -6988 2648 -6975
rect 2704 -6751 2808 -6738
rect 2704 -6975 2733 -6751
rect 2779 -6975 2808 -6751
rect 2704 -6988 2808 -6975
rect 2864 -6751 2968 -6738
rect 2864 -6975 2893 -6751
rect 2939 -6975 2968 -6751
rect 2864 -6988 2968 -6975
rect 3024 -6751 3128 -6738
rect 3024 -6975 3053 -6751
rect 3099 -6975 3128 -6751
rect 3024 -6988 3128 -6975
rect 3184 -6751 3272 -6738
rect 3184 -6975 3213 -6751
rect 3259 -6975 3272 -6751
rect 3184 -6988 3272 -6975
rect 3328 -6751 3416 -6738
rect 3328 -6975 3341 -6751
rect 3387 -6975 3416 -6751
rect 3328 -6988 3416 -6975
rect 3472 -6751 3560 -6738
rect 3472 -6975 3501 -6751
rect 3547 -6975 3560 -6751
rect 3472 -6988 3560 -6975
rect 3732 -6751 3820 -6738
rect 3732 -6975 3745 -6751
rect 3791 -6975 3820 -6751
rect 3732 -6988 3820 -6975
rect 3876 -6751 3964 -6738
rect 3876 -6975 3905 -6751
rect 3951 -6975 3964 -6751
rect 3876 -6988 3964 -6975
rect 4020 -6751 4108 -6738
rect 4020 -6975 4033 -6751
rect 4079 -6975 4108 -6751
rect 4020 -6988 4108 -6975
rect 4164 -6751 4268 -6738
rect 4164 -6975 4193 -6751
rect 4239 -6975 4268 -6751
rect 4164 -6988 4268 -6975
rect 4324 -6751 4428 -6738
rect 4324 -6975 4353 -6751
rect 4399 -6975 4428 -6751
rect 4324 -6988 4428 -6975
rect 4484 -6751 4588 -6738
rect 4484 -6975 4513 -6751
rect 4559 -6975 4588 -6751
rect 4484 -6988 4588 -6975
rect 4644 -6751 4748 -6738
rect 4644 -6975 4673 -6751
rect 4719 -6975 4748 -6751
rect 4644 -6988 4748 -6975
rect 4804 -6751 4908 -6738
rect 4804 -6975 4833 -6751
rect 4879 -6975 4908 -6751
rect 4804 -6988 4908 -6975
rect 4964 -6751 5068 -6738
rect 4964 -6975 4993 -6751
rect 5039 -6975 5068 -6751
rect 4964 -6988 5068 -6975
rect 5124 -6751 5228 -6738
rect 5124 -6975 5153 -6751
rect 5199 -6975 5228 -6751
rect 5124 -6988 5228 -6975
rect 5284 -6751 5372 -6738
rect 5284 -6975 5313 -6751
rect 5359 -6975 5372 -6751
rect 5284 -6988 5372 -6975
rect 5544 -6751 5632 -6738
rect 5544 -6975 5557 -6751
rect 5603 -6975 5632 -6751
rect 5544 -6988 5632 -6975
rect 5688 -6751 5792 -6738
rect 5688 -6975 5717 -6751
rect 5763 -6975 5792 -6751
rect 5688 -6988 5792 -6975
rect 5848 -6751 5952 -6738
rect 5848 -6975 5877 -6751
rect 5923 -6975 5952 -6751
rect 5848 -6988 5952 -6975
rect 6008 -6751 6112 -6738
rect 6008 -6975 6037 -6751
rect 6083 -6975 6112 -6751
rect 6008 -6988 6112 -6975
rect 6168 -6751 6272 -6738
rect 6168 -6975 6197 -6751
rect 6243 -6975 6272 -6751
rect 6168 -6988 6272 -6975
rect 6328 -6751 6432 -6738
rect 6328 -6975 6357 -6751
rect 6403 -6975 6432 -6751
rect 6328 -6988 6432 -6975
rect 6488 -6751 6592 -6738
rect 6488 -6975 6517 -6751
rect 6563 -6975 6592 -6751
rect 6488 -6988 6592 -6975
rect 6648 -6751 6752 -6738
rect 6648 -6975 6677 -6751
rect 6723 -6975 6752 -6751
rect 6648 -6988 6752 -6975
rect 6808 -6751 6896 -6738
rect 6808 -6975 6837 -6751
rect 6883 -6975 6896 -6751
rect 6808 -6988 6896 -6975
rect 6952 -6751 7040 -6738
rect 6952 -6975 6965 -6751
rect 7011 -6975 7040 -6751
rect 6952 -6988 7040 -6975
rect 7096 -6751 7184 -6738
rect 7096 -6975 7125 -6751
rect 7171 -6975 7184 -6751
rect 7096 -6988 7184 -6975
rect 7356 -6751 7444 -6738
rect 7356 -6975 7369 -6751
rect 7415 -6975 7444 -6751
rect 7356 -6988 7444 -6975
rect 7500 -6751 7604 -6738
rect 7500 -6975 7529 -6751
rect 7575 -6975 7604 -6751
rect 7500 -6988 7604 -6975
rect 7660 -6751 7764 -6738
rect 7660 -6975 7689 -6751
rect 7735 -6975 7764 -6751
rect 7660 -6988 7764 -6975
rect 7820 -6751 7924 -6738
rect 7820 -6975 7849 -6751
rect 7895 -6975 7924 -6751
rect 7820 -6988 7924 -6975
rect 7980 -6751 8084 -6738
rect 7980 -6975 8009 -6751
rect 8055 -6975 8084 -6751
rect 7980 -6988 8084 -6975
rect 8140 -6751 8244 -6738
rect 8140 -6975 8169 -6751
rect 8215 -6975 8244 -6751
rect 8140 -6988 8244 -6975
rect 8300 -6751 8404 -6738
rect 8300 -6975 8329 -6751
rect 8375 -6975 8404 -6751
rect 8300 -6988 8404 -6975
rect 8460 -6751 8564 -6738
rect 8460 -6975 8489 -6751
rect 8535 -6975 8564 -6751
rect 8460 -6988 8564 -6975
rect 8620 -6751 8708 -6738
rect 8620 -6975 8649 -6751
rect 8695 -6975 8708 -6751
rect 8620 -6988 8708 -6975
rect 8764 -6751 8852 -6738
rect 8764 -6975 8777 -6751
rect 8823 -6975 8852 -6751
rect 8764 -6988 8852 -6975
rect 8908 -6751 8996 -6738
rect 8908 -6975 8937 -6751
rect 8983 -6975 8996 -6751
rect 8908 -6988 8996 -6975
<< pdiff >>
rect 108 5763 196 5776
rect 108 5289 121 5763
rect 167 5289 196 5763
rect 108 5276 196 5289
rect 252 5763 356 5776
rect 252 5289 281 5763
rect 327 5289 356 5763
rect 252 5276 356 5289
rect 412 5763 516 5776
rect 412 5289 441 5763
rect 487 5289 516 5763
rect 412 5276 516 5289
rect 572 5763 676 5776
rect 572 5289 601 5763
rect 647 5289 676 5763
rect 572 5276 676 5289
rect 732 5763 836 5776
rect 732 5289 761 5763
rect 807 5289 836 5763
rect 732 5276 836 5289
rect 892 5763 996 5776
rect 892 5289 921 5763
rect 967 5289 996 5763
rect 892 5276 996 5289
rect 1052 5763 1156 5776
rect 1052 5289 1081 5763
rect 1127 5289 1156 5763
rect 1052 5276 1156 5289
rect 1212 5763 1316 5776
rect 1212 5289 1241 5763
rect 1287 5289 1316 5763
rect 1212 5276 1316 5289
rect 1372 5763 1460 5776
rect 1372 5289 1401 5763
rect 1447 5289 1460 5763
rect 1372 5276 1460 5289
rect 1516 5763 1604 5776
rect 1516 5289 1529 5763
rect 1575 5289 1604 5763
rect 1516 5276 1604 5289
rect 1660 5763 1748 5776
rect 1660 5289 1689 5763
rect 1735 5289 1748 5763
rect 1660 5276 1748 5289
rect 1920 5763 2008 5776
rect 1920 5289 1933 5763
rect 1979 5289 2008 5763
rect 1920 5276 2008 5289
rect 2064 5763 2152 5776
rect 2064 5289 2093 5763
rect 2139 5289 2152 5763
rect 2064 5276 2152 5289
rect 2208 5763 2296 5776
rect 2208 5289 2221 5763
rect 2267 5289 2296 5763
rect 2208 5276 2296 5289
rect 2352 5763 2456 5776
rect 2352 5289 2381 5763
rect 2427 5289 2456 5763
rect 2352 5276 2456 5289
rect 2512 5763 2616 5776
rect 2512 5289 2541 5763
rect 2587 5289 2616 5763
rect 2512 5276 2616 5289
rect 2672 5763 2776 5776
rect 2672 5289 2701 5763
rect 2747 5289 2776 5763
rect 2672 5276 2776 5289
rect 2832 5763 2936 5776
rect 2832 5289 2861 5763
rect 2907 5289 2936 5763
rect 2832 5276 2936 5289
rect 2992 5763 3096 5776
rect 2992 5289 3021 5763
rect 3067 5289 3096 5763
rect 2992 5276 3096 5289
rect 3152 5763 3256 5776
rect 3152 5289 3181 5763
rect 3227 5289 3256 5763
rect 3152 5276 3256 5289
rect 3312 5763 3416 5776
rect 3312 5289 3341 5763
rect 3387 5289 3416 5763
rect 3312 5276 3416 5289
rect 3472 5763 3560 5776
rect 3472 5289 3501 5763
rect 3547 5289 3560 5763
rect 3472 5276 3560 5289
rect 3732 5763 3820 5776
rect 3732 5289 3745 5763
rect 3791 5289 3820 5763
rect 3732 5276 3820 5289
rect 3876 5763 3964 5776
rect 3876 5289 3905 5763
rect 3951 5289 3964 5763
rect 3876 5276 3964 5289
rect 4020 5763 4108 5776
rect 4020 5289 4033 5763
rect 4079 5289 4108 5763
rect 4020 5276 4108 5289
rect 4164 5763 4268 5776
rect 4164 5289 4193 5763
rect 4239 5289 4268 5763
rect 4164 5276 4268 5289
rect 4324 5763 4428 5776
rect 4324 5289 4353 5763
rect 4399 5289 4428 5763
rect 4324 5276 4428 5289
rect 4484 5763 4588 5776
rect 4484 5289 4513 5763
rect 4559 5289 4588 5763
rect 4484 5276 4588 5289
rect 4644 5763 4748 5776
rect 4644 5289 4673 5763
rect 4719 5289 4748 5763
rect 4644 5276 4748 5289
rect 4804 5763 4908 5776
rect 4804 5289 4833 5763
rect 4879 5289 4908 5763
rect 4804 5276 4908 5289
rect 4964 5763 5068 5776
rect 4964 5289 4993 5763
rect 5039 5289 5068 5763
rect 4964 5276 5068 5289
rect 5124 5763 5228 5776
rect 5124 5289 5153 5763
rect 5199 5289 5228 5763
rect 5124 5276 5228 5289
rect 5284 5763 5372 5776
rect 5284 5289 5313 5763
rect 5359 5289 5372 5763
rect 5284 5276 5372 5289
rect 5544 5763 5632 5776
rect 5544 5289 5557 5763
rect 5603 5289 5632 5763
rect 5544 5276 5632 5289
rect 5688 5763 5776 5776
rect 5688 5289 5717 5763
rect 5763 5289 5776 5763
rect 5688 5276 5776 5289
rect 5832 5763 5920 5776
rect 5832 5289 5845 5763
rect 5891 5289 5920 5763
rect 5832 5276 5920 5289
rect 5976 5763 6080 5776
rect 5976 5289 6005 5763
rect 6051 5289 6080 5763
rect 5976 5276 6080 5289
rect 6136 5763 6240 5776
rect 6136 5289 6165 5763
rect 6211 5289 6240 5763
rect 6136 5276 6240 5289
rect 6296 5763 6400 5776
rect 6296 5289 6325 5763
rect 6371 5289 6400 5763
rect 6296 5276 6400 5289
rect 6456 5763 6560 5776
rect 6456 5289 6485 5763
rect 6531 5289 6560 5763
rect 6456 5276 6560 5289
rect 6616 5763 6720 5776
rect 6616 5289 6645 5763
rect 6691 5289 6720 5763
rect 6616 5276 6720 5289
rect 6776 5763 6880 5776
rect 6776 5289 6805 5763
rect 6851 5289 6880 5763
rect 6776 5276 6880 5289
rect 6936 5763 7040 5776
rect 6936 5289 6965 5763
rect 7011 5289 7040 5763
rect 6936 5276 7040 5289
rect 7096 5763 7184 5776
rect 7096 5289 7125 5763
rect 7171 5289 7184 5763
rect 7096 5276 7184 5289
rect 7356 5763 7444 5776
rect 7356 5289 7369 5763
rect 7415 5289 7444 5763
rect 7356 5276 7444 5289
rect 7500 5763 7588 5776
rect 7500 5289 7529 5763
rect 7575 5289 7588 5763
rect 7500 5276 7588 5289
rect 7644 5763 7732 5776
rect 7644 5289 7657 5763
rect 7703 5289 7732 5763
rect 7644 5276 7732 5289
rect 7788 5763 7892 5776
rect 7788 5289 7817 5763
rect 7863 5289 7892 5763
rect 7788 5276 7892 5289
rect 7948 5763 8052 5776
rect 7948 5289 7977 5763
rect 8023 5289 8052 5763
rect 7948 5276 8052 5289
rect 8108 5763 8212 5776
rect 8108 5289 8137 5763
rect 8183 5289 8212 5763
rect 8108 5276 8212 5289
rect 8268 5763 8372 5776
rect 8268 5289 8297 5763
rect 8343 5289 8372 5763
rect 8268 5276 8372 5289
rect 8428 5763 8532 5776
rect 8428 5289 8457 5763
rect 8503 5289 8532 5763
rect 8428 5276 8532 5289
rect 8588 5763 8692 5776
rect 8588 5289 8617 5763
rect 8663 5289 8692 5763
rect 8588 5276 8692 5289
rect 8748 5763 8852 5776
rect 8748 5289 8777 5763
rect 8823 5289 8852 5763
rect 8748 5276 8852 5289
rect 8908 5763 8996 5776
rect 8908 5289 8937 5763
rect 8983 5289 8996 5763
rect 8908 5276 8996 5289
rect 108 5127 196 5140
rect 108 4653 121 5127
rect 167 4653 196 5127
rect 108 4640 196 4653
rect 252 5127 356 5140
rect 252 4653 281 5127
rect 327 4653 356 5127
rect 252 4640 356 4653
rect 412 5127 516 5140
rect 412 4653 441 5127
rect 487 4653 516 5127
rect 412 4640 516 4653
rect 572 5127 676 5140
rect 572 4653 601 5127
rect 647 4653 676 5127
rect 572 4640 676 4653
rect 732 5127 836 5140
rect 732 4653 761 5127
rect 807 4653 836 5127
rect 732 4640 836 4653
rect 892 5127 996 5140
rect 892 4653 921 5127
rect 967 4653 996 5127
rect 892 4640 996 4653
rect 1052 5127 1156 5140
rect 1052 4653 1081 5127
rect 1127 4653 1156 5127
rect 1052 4640 1156 4653
rect 1212 5127 1316 5140
rect 1212 4653 1241 5127
rect 1287 4653 1316 5127
rect 1212 4640 1316 4653
rect 1372 5127 1460 5140
rect 1372 4653 1401 5127
rect 1447 4653 1460 5127
rect 1372 4640 1460 4653
rect 1516 5127 1604 5140
rect 1516 4653 1529 5127
rect 1575 4653 1604 5127
rect 1516 4640 1604 4653
rect 1660 5127 1748 5140
rect 1660 4653 1689 5127
rect 1735 4653 1748 5127
rect 1660 4640 1748 4653
rect 1920 5127 2008 5140
rect 1920 4653 1933 5127
rect 1979 4653 2008 5127
rect 1920 4640 2008 4653
rect 2064 5127 2152 5140
rect 2064 4653 2093 5127
rect 2139 4653 2152 5127
rect 2064 4640 2152 4653
rect 2208 5127 2296 5140
rect 2208 4653 2221 5127
rect 2267 4653 2296 5127
rect 2208 4640 2296 4653
rect 2352 5127 2456 5140
rect 2352 4653 2381 5127
rect 2427 4653 2456 5127
rect 2352 4640 2456 4653
rect 2512 5127 2616 5140
rect 2512 4653 2541 5127
rect 2587 4653 2616 5127
rect 2512 4640 2616 4653
rect 2672 5127 2776 5140
rect 2672 4653 2701 5127
rect 2747 4653 2776 5127
rect 2672 4640 2776 4653
rect 2832 5127 2936 5140
rect 2832 4653 2861 5127
rect 2907 4653 2936 5127
rect 2832 4640 2936 4653
rect 2992 5127 3096 5140
rect 2992 4653 3021 5127
rect 3067 4653 3096 5127
rect 2992 4640 3096 4653
rect 3152 5127 3256 5140
rect 3152 4653 3181 5127
rect 3227 4653 3256 5127
rect 3152 4640 3256 4653
rect 3312 5127 3416 5140
rect 3312 4653 3341 5127
rect 3387 4653 3416 5127
rect 3312 4640 3416 4653
rect 3472 5127 3560 5140
rect 3472 4653 3501 5127
rect 3547 4653 3560 5127
rect 3472 4640 3560 4653
rect 3732 5127 3820 5140
rect 3732 4653 3745 5127
rect 3791 4653 3820 5127
rect 3732 4640 3820 4653
rect 3876 5127 3964 5140
rect 3876 4653 3905 5127
rect 3951 4653 3964 5127
rect 3876 4640 3964 4653
rect 4020 5127 4108 5140
rect 4020 4653 4033 5127
rect 4079 4653 4108 5127
rect 4020 4640 4108 4653
rect 4164 5127 4268 5140
rect 4164 4653 4193 5127
rect 4239 4653 4268 5127
rect 4164 4640 4268 4653
rect 4324 5127 4428 5140
rect 4324 4653 4353 5127
rect 4399 4653 4428 5127
rect 4324 4640 4428 4653
rect 4484 5127 4588 5140
rect 4484 4653 4513 5127
rect 4559 4653 4588 5127
rect 4484 4640 4588 4653
rect 4644 5127 4748 5140
rect 4644 4653 4673 5127
rect 4719 4653 4748 5127
rect 4644 4640 4748 4653
rect 4804 5127 4908 5140
rect 4804 4653 4833 5127
rect 4879 4653 4908 5127
rect 4804 4640 4908 4653
rect 4964 5127 5068 5140
rect 4964 4653 4993 5127
rect 5039 4653 5068 5127
rect 4964 4640 5068 4653
rect 5124 5127 5228 5140
rect 5124 4653 5153 5127
rect 5199 4653 5228 5127
rect 5124 4640 5228 4653
rect 5284 5127 5372 5140
rect 5284 4653 5313 5127
rect 5359 4653 5372 5127
rect 5284 4640 5372 4653
rect 5544 5127 5632 5140
rect 5544 4653 5557 5127
rect 5603 4653 5632 5127
rect 5544 4640 5632 4653
rect 5688 5127 5776 5140
rect 5688 4653 5717 5127
rect 5763 4653 5776 5127
rect 5688 4640 5776 4653
rect 5832 5127 5920 5140
rect 5832 4653 5845 5127
rect 5891 4653 5920 5127
rect 5832 4640 5920 4653
rect 5976 5127 6080 5140
rect 5976 4653 6005 5127
rect 6051 4653 6080 5127
rect 5976 4640 6080 4653
rect 6136 5127 6240 5140
rect 6136 4653 6165 5127
rect 6211 4653 6240 5127
rect 6136 4640 6240 4653
rect 6296 5127 6400 5140
rect 6296 4653 6325 5127
rect 6371 4653 6400 5127
rect 6296 4640 6400 4653
rect 6456 5127 6560 5140
rect 6456 4653 6485 5127
rect 6531 4653 6560 5127
rect 6456 4640 6560 4653
rect 6616 5127 6720 5140
rect 6616 4653 6645 5127
rect 6691 4653 6720 5127
rect 6616 4640 6720 4653
rect 6776 5127 6880 5140
rect 6776 4653 6805 5127
rect 6851 4653 6880 5127
rect 6776 4640 6880 4653
rect 6936 5127 7040 5140
rect 6936 4653 6965 5127
rect 7011 4653 7040 5127
rect 6936 4640 7040 4653
rect 7096 5127 7184 5140
rect 7096 4653 7125 5127
rect 7171 4653 7184 5127
rect 7096 4640 7184 4653
rect 7356 5127 7444 5140
rect 7356 4653 7369 5127
rect 7415 4653 7444 5127
rect 7356 4640 7444 4653
rect 7500 5127 7588 5140
rect 7500 4653 7529 5127
rect 7575 4653 7588 5127
rect 7500 4640 7588 4653
rect 7644 5127 7732 5140
rect 7644 4653 7657 5127
rect 7703 4653 7732 5127
rect 7644 4640 7732 4653
rect 7788 5127 7892 5140
rect 7788 4653 7817 5127
rect 7863 4653 7892 5127
rect 7788 4640 7892 4653
rect 7948 5127 8052 5140
rect 7948 4653 7977 5127
rect 8023 4653 8052 5127
rect 7948 4640 8052 4653
rect 8108 5127 8212 5140
rect 8108 4653 8137 5127
rect 8183 4653 8212 5127
rect 8108 4640 8212 4653
rect 8268 5127 8372 5140
rect 8268 4653 8297 5127
rect 8343 4653 8372 5127
rect 8268 4640 8372 4653
rect 8428 5127 8532 5140
rect 8428 4653 8457 5127
rect 8503 4653 8532 5127
rect 8428 4640 8532 4653
rect 8588 5127 8692 5140
rect 8588 4653 8617 5127
rect 8663 4653 8692 5127
rect 8588 4640 8692 4653
rect 8748 5127 8852 5140
rect 8748 4653 8777 5127
rect 8823 4653 8852 5127
rect 8748 4640 8852 4653
rect 8908 5127 8996 5140
rect 8908 4653 8937 5127
rect 8983 4653 8996 5127
rect 8908 4640 8996 4653
rect 108 4491 196 4504
rect 108 4017 121 4491
rect 167 4017 196 4491
rect 108 4004 196 4017
rect 252 4491 356 4504
rect 252 4017 281 4491
rect 327 4017 356 4491
rect 252 4004 356 4017
rect 412 4491 516 4504
rect 412 4017 441 4491
rect 487 4017 516 4491
rect 412 4004 516 4017
rect 572 4491 676 4504
rect 572 4017 601 4491
rect 647 4017 676 4491
rect 572 4004 676 4017
rect 732 4491 836 4504
rect 732 4017 761 4491
rect 807 4017 836 4491
rect 732 4004 836 4017
rect 892 4491 996 4504
rect 892 4017 921 4491
rect 967 4017 996 4491
rect 892 4004 996 4017
rect 1052 4491 1156 4504
rect 1052 4017 1081 4491
rect 1127 4017 1156 4491
rect 1052 4004 1156 4017
rect 1212 4491 1316 4504
rect 1212 4017 1241 4491
rect 1287 4017 1316 4491
rect 1212 4004 1316 4017
rect 1372 4491 1460 4504
rect 1372 4017 1401 4491
rect 1447 4017 1460 4491
rect 1372 4004 1460 4017
rect 1516 4491 1604 4504
rect 1516 4017 1529 4491
rect 1575 4017 1604 4491
rect 1516 4004 1604 4017
rect 1660 4491 1748 4504
rect 1660 4017 1689 4491
rect 1735 4017 1748 4491
rect 1660 4004 1748 4017
rect 1920 4491 2008 4504
rect 1920 4017 1933 4491
rect 1979 4017 2008 4491
rect 1920 4004 2008 4017
rect 2064 4491 2152 4504
rect 2064 4017 2093 4491
rect 2139 4017 2152 4491
rect 2064 4004 2152 4017
rect 2208 4491 2296 4504
rect 2208 4017 2221 4491
rect 2267 4017 2296 4491
rect 2208 4004 2296 4017
rect 2352 4491 2456 4504
rect 2352 4017 2381 4491
rect 2427 4017 2456 4491
rect 2352 4004 2456 4017
rect 2512 4491 2616 4504
rect 2512 4017 2541 4491
rect 2587 4017 2616 4491
rect 2512 4004 2616 4017
rect 2672 4491 2776 4504
rect 2672 4017 2701 4491
rect 2747 4017 2776 4491
rect 2672 4004 2776 4017
rect 2832 4491 2936 4504
rect 2832 4017 2861 4491
rect 2907 4017 2936 4491
rect 2832 4004 2936 4017
rect 2992 4491 3096 4504
rect 2992 4017 3021 4491
rect 3067 4017 3096 4491
rect 2992 4004 3096 4017
rect 3152 4491 3256 4504
rect 3152 4017 3181 4491
rect 3227 4017 3256 4491
rect 3152 4004 3256 4017
rect 3312 4491 3416 4504
rect 3312 4017 3341 4491
rect 3387 4017 3416 4491
rect 3312 4004 3416 4017
rect 3472 4491 3560 4504
rect 3472 4017 3501 4491
rect 3547 4017 3560 4491
rect 3472 4004 3560 4017
rect 3732 4491 3820 4504
rect 3732 4017 3745 4491
rect 3791 4017 3820 4491
rect 3732 4004 3820 4017
rect 3876 4491 3964 4504
rect 3876 4017 3905 4491
rect 3951 4017 3964 4491
rect 3876 4004 3964 4017
rect 4020 4491 4108 4504
rect 4020 4017 4033 4491
rect 4079 4017 4108 4491
rect 4020 4004 4108 4017
rect 4164 4491 4268 4504
rect 4164 4017 4193 4491
rect 4239 4017 4268 4491
rect 4164 4004 4268 4017
rect 4324 4491 4428 4504
rect 4324 4017 4353 4491
rect 4399 4017 4428 4491
rect 4324 4004 4428 4017
rect 4484 4491 4588 4504
rect 4484 4017 4513 4491
rect 4559 4017 4588 4491
rect 4484 4004 4588 4017
rect 4644 4491 4748 4504
rect 4644 4017 4673 4491
rect 4719 4017 4748 4491
rect 4644 4004 4748 4017
rect 4804 4491 4908 4504
rect 4804 4017 4833 4491
rect 4879 4017 4908 4491
rect 4804 4004 4908 4017
rect 4964 4491 5068 4504
rect 4964 4017 4993 4491
rect 5039 4017 5068 4491
rect 4964 4004 5068 4017
rect 5124 4491 5228 4504
rect 5124 4017 5153 4491
rect 5199 4017 5228 4491
rect 5124 4004 5228 4017
rect 5284 4491 5372 4504
rect 5284 4017 5313 4491
rect 5359 4017 5372 4491
rect 5284 4004 5372 4017
rect 5544 4491 5632 4504
rect 5544 4017 5557 4491
rect 5603 4017 5632 4491
rect 5544 4004 5632 4017
rect 5688 4491 5776 4504
rect 5688 4017 5717 4491
rect 5763 4017 5776 4491
rect 5688 4004 5776 4017
rect 5832 4491 5920 4504
rect 5832 4017 5845 4491
rect 5891 4017 5920 4491
rect 5832 4004 5920 4017
rect 5976 4491 6080 4504
rect 5976 4017 6005 4491
rect 6051 4017 6080 4491
rect 5976 4004 6080 4017
rect 6136 4491 6240 4504
rect 6136 4017 6165 4491
rect 6211 4017 6240 4491
rect 6136 4004 6240 4017
rect 6296 4491 6400 4504
rect 6296 4017 6325 4491
rect 6371 4017 6400 4491
rect 6296 4004 6400 4017
rect 6456 4491 6560 4504
rect 6456 4017 6485 4491
rect 6531 4017 6560 4491
rect 6456 4004 6560 4017
rect 6616 4491 6720 4504
rect 6616 4017 6645 4491
rect 6691 4017 6720 4491
rect 6616 4004 6720 4017
rect 6776 4491 6880 4504
rect 6776 4017 6805 4491
rect 6851 4017 6880 4491
rect 6776 4004 6880 4017
rect 6936 4491 7040 4504
rect 6936 4017 6965 4491
rect 7011 4017 7040 4491
rect 6936 4004 7040 4017
rect 7096 4491 7184 4504
rect 7096 4017 7125 4491
rect 7171 4017 7184 4491
rect 7096 4004 7184 4017
rect 7356 4491 7444 4504
rect 7356 4017 7369 4491
rect 7415 4017 7444 4491
rect 7356 4004 7444 4017
rect 7500 4491 7588 4504
rect 7500 4017 7529 4491
rect 7575 4017 7588 4491
rect 7500 4004 7588 4017
rect 7644 4491 7732 4504
rect 7644 4017 7657 4491
rect 7703 4017 7732 4491
rect 7644 4004 7732 4017
rect 7788 4491 7892 4504
rect 7788 4017 7817 4491
rect 7863 4017 7892 4491
rect 7788 4004 7892 4017
rect 7948 4491 8052 4504
rect 7948 4017 7977 4491
rect 8023 4017 8052 4491
rect 7948 4004 8052 4017
rect 8108 4491 8212 4504
rect 8108 4017 8137 4491
rect 8183 4017 8212 4491
rect 8108 4004 8212 4017
rect 8268 4491 8372 4504
rect 8268 4017 8297 4491
rect 8343 4017 8372 4491
rect 8268 4004 8372 4017
rect 8428 4491 8532 4504
rect 8428 4017 8457 4491
rect 8503 4017 8532 4491
rect 8428 4004 8532 4017
rect 8588 4491 8692 4504
rect 8588 4017 8617 4491
rect 8663 4017 8692 4491
rect 8588 4004 8692 4017
rect 8748 4491 8852 4504
rect 8748 4017 8777 4491
rect 8823 4017 8852 4491
rect 8748 4004 8852 4017
rect 8908 4491 8996 4504
rect 8908 4017 8937 4491
rect 8983 4017 8996 4491
rect 8908 4004 8996 4017
rect -4812 3560 -4724 3573
rect -4812 3386 -4799 3560
rect -4753 3386 -4724 3560
rect -4812 3373 -4724 3386
rect -4668 3560 -4580 3573
rect -4668 3386 -4639 3560
rect -4593 3386 -4580 3560
rect -1163 3560 -1075 3573
rect -4668 3373 -4580 3386
rect -4406 3515 -4318 3528
rect -4406 3341 -4393 3515
rect -4347 3341 -4318 3515
rect -4406 3328 -4318 3341
rect -4262 3515 -4158 3528
rect -4262 3341 -4233 3515
rect -4187 3341 -4158 3515
rect -4262 3328 -4158 3341
rect -4102 3515 -3998 3528
rect -4102 3341 -4073 3515
rect -4027 3341 -3998 3515
rect -4102 3328 -3998 3341
rect -3942 3515 -3838 3528
rect -3942 3341 -3913 3515
rect -3867 3341 -3838 3515
rect -3942 3328 -3838 3341
rect -3782 3515 -3694 3528
rect -3782 3341 -3753 3515
rect -3707 3341 -3694 3515
rect -3533 3526 -3445 3539
rect -3533 3464 -3520 3526
rect -3474 3464 -3445 3526
rect -3533 3451 -3445 3464
rect -2997 3526 -2909 3539
rect -2997 3464 -2968 3526
rect -2922 3464 -2909 3526
rect -2997 3451 -2909 3464
rect -2747 3526 -2659 3539
rect -2747 3464 -2734 3526
rect -2688 3464 -2659 3526
rect -2747 3451 -2659 3464
rect -2211 3526 -2123 3539
rect -2211 3464 -2182 3526
rect -2136 3464 -2123 3526
rect -2211 3451 -2123 3464
rect -1961 3526 -1873 3539
rect -1961 3464 -1948 3526
rect -1902 3464 -1873 3526
rect -1961 3451 -1873 3464
rect -1425 3526 -1337 3539
rect -1425 3464 -1396 3526
rect -1350 3464 -1337 3526
rect -1425 3451 -1337 3464
rect -3782 3328 -3694 3341
rect -1163 3386 -1150 3560
rect -1104 3386 -1075 3560
rect -1163 3373 -1075 3386
rect -1019 3560 -931 3573
rect -1019 3386 -990 3560
rect -944 3386 -931 3560
rect -1019 3373 -931 3386
rect 108 3423 196 3436
rect 108 2949 121 3423
rect 167 2949 196 3423
rect 108 2936 196 2949
rect 252 3423 340 3436
rect 252 2949 281 3423
rect 327 2949 340 3423
rect 252 2936 340 2949
rect 396 3423 484 3436
rect 396 2949 409 3423
rect 455 2949 484 3423
rect 396 2936 484 2949
rect 540 3423 644 3436
rect 540 2949 569 3423
rect 615 2949 644 3423
rect 540 2936 644 2949
rect 700 3423 804 3436
rect 700 2949 729 3423
rect 775 2949 804 3423
rect 700 2936 804 2949
rect 860 3423 964 3436
rect 860 2949 889 3423
rect 935 2949 964 3423
rect 860 2936 964 2949
rect 1020 3423 1124 3436
rect 1020 2949 1049 3423
rect 1095 2949 1124 3423
rect 1020 2936 1124 2949
rect 1180 3423 1284 3436
rect 1180 2949 1209 3423
rect 1255 2949 1284 3423
rect 1180 2936 1284 2949
rect 1340 3423 1444 3436
rect 1340 2949 1369 3423
rect 1415 2949 1444 3423
rect 1340 2936 1444 2949
rect 1500 3423 1604 3436
rect 1500 2949 1529 3423
rect 1575 2949 1604 3423
rect 1500 2936 1604 2949
rect 1660 3423 1748 3436
rect 1660 2949 1689 3423
rect 1735 2949 1748 3423
rect 1660 2936 1748 2949
rect 1920 3423 2008 3436
rect 1920 2949 1933 3423
rect 1979 2949 2008 3423
rect 1920 2936 2008 2949
rect 2064 3423 2168 3436
rect 2064 2949 2093 3423
rect 2139 2949 2168 3423
rect 2064 2936 2168 2949
rect 2224 3423 2328 3436
rect 2224 2949 2253 3423
rect 2299 2949 2328 3423
rect 2224 2936 2328 2949
rect 2384 3423 2488 3436
rect 2384 2949 2413 3423
rect 2459 2949 2488 3423
rect 2384 2936 2488 2949
rect 2544 3423 2648 3436
rect 2544 2949 2573 3423
rect 2619 2949 2648 3423
rect 2544 2936 2648 2949
rect 2704 3423 2808 3436
rect 2704 2949 2733 3423
rect 2779 2949 2808 3423
rect 2704 2936 2808 2949
rect 2864 3423 2968 3436
rect 2864 2949 2893 3423
rect 2939 2949 2968 3423
rect 2864 2936 2968 2949
rect 3024 3423 3128 3436
rect 3024 2949 3053 3423
rect 3099 2949 3128 3423
rect 3024 2936 3128 2949
rect 3184 3423 3272 3436
rect 3184 2949 3213 3423
rect 3259 2949 3272 3423
rect 3184 2936 3272 2949
rect 3328 3423 3416 3436
rect 3328 2949 3341 3423
rect 3387 2949 3416 3423
rect 3328 2936 3416 2949
rect 3472 3423 3560 3436
rect 3472 2949 3501 3423
rect 3547 2949 3560 3423
rect 3472 2936 3560 2949
rect 3732 3423 3820 3436
rect 3732 2949 3745 3423
rect 3791 2949 3820 3423
rect 3732 2936 3820 2949
rect 3876 3423 3964 3436
rect 3876 2949 3905 3423
rect 3951 2949 3964 3423
rect 3876 2936 3964 2949
rect 4020 3423 4108 3436
rect 4020 2949 4033 3423
rect 4079 2949 4108 3423
rect 4020 2936 4108 2949
rect 4164 3423 4268 3436
rect 4164 2949 4193 3423
rect 4239 2949 4268 3423
rect 4164 2936 4268 2949
rect 4324 3423 4428 3436
rect 4324 2949 4353 3423
rect 4399 2949 4428 3423
rect 4324 2936 4428 2949
rect 4484 3423 4588 3436
rect 4484 2949 4513 3423
rect 4559 2949 4588 3423
rect 4484 2936 4588 2949
rect 4644 3423 4748 3436
rect 4644 2949 4673 3423
rect 4719 2949 4748 3423
rect 4644 2936 4748 2949
rect 4804 3423 4908 3436
rect 4804 2949 4833 3423
rect 4879 2949 4908 3423
rect 4804 2936 4908 2949
rect 4964 3423 5068 3436
rect 4964 2949 4993 3423
rect 5039 2949 5068 3423
rect 4964 2936 5068 2949
rect 5124 3423 5228 3436
rect 5124 2949 5153 3423
rect 5199 2949 5228 3423
rect 5124 2936 5228 2949
rect 5284 3423 5372 3436
rect 5284 2949 5313 3423
rect 5359 2949 5372 3423
rect 5284 2936 5372 2949
rect 5544 3423 5632 3436
rect 5544 2949 5557 3423
rect 5603 2949 5632 3423
rect 5544 2936 5632 2949
rect 5688 3423 5792 3436
rect 5688 2949 5717 3423
rect 5763 2949 5792 3423
rect 5688 2936 5792 2949
rect 5848 3423 5952 3436
rect 5848 2949 5877 3423
rect 5923 2949 5952 3423
rect 5848 2936 5952 2949
rect 6008 3423 6112 3436
rect 6008 2949 6037 3423
rect 6083 2949 6112 3423
rect 6008 2936 6112 2949
rect 6168 3423 6272 3436
rect 6168 2949 6197 3423
rect 6243 2949 6272 3423
rect 6168 2936 6272 2949
rect 6328 3423 6432 3436
rect 6328 2949 6357 3423
rect 6403 2949 6432 3423
rect 6328 2936 6432 2949
rect 6488 3423 6592 3436
rect 6488 2949 6517 3423
rect 6563 2949 6592 3423
rect 6488 2936 6592 2949
rect 6648 3423 6752 3436
rect 6648 2949 6677 3423
rect 6723 2949 6752 3423
rect 6648 2936 6752 2949
rect 6808 3423 6896 3436
rect 6808 2949 6837 3423
rect 6883 2949 6896 3423
rect 6808 2936 6896 2949
rect 6952 3423 7040 3436
rect 6952 2949 6965 3423
rect 7011 2949 7040 3423
rect 6952 2936 7040 2949
rect 7096 3423 7184 3436
rect 7096 2949 7125 3423
rect 7171 2949 7184 3423
rect 7096 2936 7184 2949
rect 7356 3423 7444 3436
rect 7356 2949 7369 3423
rect 7415 2949 7444 3423
rect 7356 2936 7444 2949
rect 7500 3423 7604 3436
rect 7500 2949 7529 3423
rect 7575 2949 7604 3423
rect 7500 2936 7604 2949
rect 7660 3423 7764 3436
rect 7660 2949 7689 3423
rect 7735 2949 7764 3423
rect 7660 2936 7764 2949
rect 7820 3423 7924 3436
rect 7820 2949 7849 3423
rect 7895 2949 7924 3423
rect 7820 2936 7924 2949
rect 7980 3423 8084 3436
rect 7980 2949 8009 3423
rect 8055 2949 8084 3423
rect 7980 2936 8084 2949
rect 8140 3423 8244 3436
rect 8140 2949 8169 3423
rect 8215 2949 8244 3423
rect 8140 2936 8244 2949
rect 8300 3423 8404 3436
rect 8300 2949 8329 3423
rect 8375 2949 8404 3423
rect 8300 2936 8404 2949
rect 8460 3423 8564 3436
rect 8460 2949 8489 3423
rect 8535 2949 8564 3423
rect 8460 2936 8564 2949
rect 8620 3423 8708 3436
rect 8620 2949 8649 3423
rect 8695 2949 8708 3423
rect 8620 2936 8708 2949
rect 8764 3423 8852 3436
rect 8764 2949 8777 3423
rect 8823 2949 8852 3423
rect 8764 2936 8852 2949
rect 8908 3423 8996 3436
rect 8908 2949 8937 3423
rect 8983 2949 8996 3423
rect 8908 2936 8996 2949
rect 108 2787 196 2800
rect -4406 2389 -4318 2402
rect -4406 2215 -4393 2389
rect -4347 2215 -4318 2389
rect -4406 2202 -4318 2215
rect -4262 2389 -4158 2402
rect -4262 2215 -4233 2389
rect -4187 2215 -4158 2389
rect -4262 2202 -4158 2215
rect -4102 2389 -3998 2402
rect -4102 2215 -4073 2389
rect -4027 2215 -3998 2389
rect -4102 2202 -3998 2215
rect -3942 2389 -3838 2402
rect -3942 2215 -3913 2389
rect -3867 2215 -3838 2389
rect -3942 2202 -3838 2215
rect -3782 2389 -3694 2402
rect -3782 2215 -3753 2389
rect -3707 2215 -3694 2389
rect -1163 2344 -1075 2357
rect -3782 2202 -3694 2215
rect -3533 2266 -3445 2279
rect -3533 2204 -3520 2266
rect -3474 2204 -3445 2266
rect -3533 2191 -3445 2204
rect -2997 2266 -2909 2279
rect -2997 2204 -2968 2266
rect -2922 2204 -2909 2266
rect -2997 2191 -2909 2204
rect -2747 2266 -2659 2279
rect -2747 2204 -2734 2266
rect -2688 2204 -2659 2266
rect -2747 2191 -2659 2204
rect -2211 2266 -2123 2279
rect -2211 2204 -2182 2266
rect -2136 2204 -2123 2266
rect -2211 2191 -2123 2204
rect -1961 2266 -1873 2279
rect -1961 2204 -1948 2266
rect -1902 2204 -1873 2266
rect -1961 2191 -1873 2204
rect -1425 2266 -1337 2279
rect -1425 2204 -1396 2266
rect -1350 2204 -1337 2266
rect -1425 2191 -1337 2204
rect -1163 2170 -1150 2344
rect -1104 2170 -1075 2344
rect -1163 2157 -1075 2170
rect -1019 2344 -931 2357
rect -1019 2170 -990 2344
rect -944 2170 -931 2344
rect 108 2313 121 2787
rect 167 2313 196 2787
rect 108 2300 196 2313
rect 252 2787 340 2800
rect 252 2313 281 2787
rect 327 2313 340 2787
rect 252 2300 340 2313
rect 396 2787 484 2800
rect 396 2313 409 2787
rect 455 2313 484 2787
rect 396 2300 484 2313
rect 540 2787 644 2800
rect 540 2313 569 2787
rect 615 2313 644 2787
rect 540 2300 644 2313
rect 700 2787 804 2800
rect 700 2313 729 2787
rect 775 2313 804 2787
rect 700 2300 804 2313
rect 860 2787 964 2800
rect 860 2313 889 2787
rect 935 2313 964 2787
rect 860 2300 964 2313
rect 1020 2787 1124 2800
rect 1020 2313 1049 2787
rect 1095 2313 1124 2787
rect 1020 2300 1124 2313
rect 1180 2787 1284 2800
rect 1180 2313 1209 2787
rect 1255 2313 1284 2787
rect 1180 2300 1284 2313
rect 1340 2787 1444 2800
rect 1340 2313 1369 2787
rect 1415 2313 1444 2787
rect 1340 2300 1444 2313
rect 1500 2787 1604 2800
rect 1500 2313 1529 2787
rect 1575 2313 1604 2787
rect 1500 2300 1604 2313
rect 1660 2787 1748 2800
rect 1660 2313 1689 2787
rect 1735 2313 1748 2787
rect 1660 2300 1748 2313
rect 1920 2787 2008 2800
rect 1920 2313 1933 2787
rect 1979 2313 2008 2787
rect 1920 2300 2008 2313
rect 2064 2787 2168 2800
rect 2064 2313 2093 2787
rect 2139 2313 2168 2787
rect 2064 2300 2168 2313
rect 2224 2787 2328 2800
rect 2224 2313 2253 2787
rect 2299 2313 2328 2787
rect 2224 2300 2328 2313
rect 2384 2787 2488 2800
rect 2384 2313 2413 2787
rect 2459 2313 2488 2787
rect 2384 2300 2488 2313
rect 2544 2787 2648 2800
rect 2544 2313 2573 2787
rect 2619 2313 2648 2787
rect 2544 2300 2648 2313
rect 2704 2787 2808 2800
rect 2704 2313 2733 2787
rect 2779 2313 2808 2787
rect 2704 2300 2808 2313
rect 2864 2787 2968 2800
rect 2864 2313 2893 2787
rect 2939 2313 2968 2787
rect 2864 2300 2968 2313
rect 3024 2787 3128 2800
rect 3024 2313 3053 2787
rect 3099 2313 3128 2787
rect 3024 2300 3128 2313
rect 3184 2787 3272 2800
rect 3184 2313 3213 2787
rect 3259 2313 3272 2787
rect 3184 2300 3272 2313
rect 3328 2787 3416 2800
rect 3328 2313 3341 2787
rect 3387 2313 3416 2787
rect 3328 2300 3416 2313
rect 3472 2787 3560 2800
rect 3472 2313 3501 2787
rect 3547 2313 3560 2787
rect 3472 2300 3560 2313
rect 3732 2787 3820 2800
rect 3732 2313 3745 2787
rect 3791 2313 3820 2787
rect 3732 2300 3820 2313
rect 3876 2787 3964 2800
rect 3876 2313 3905 2787
rect 3951 2313 3964 2787
rect 3876 2300 3964 2313
rect 4020 2787 4108 2800
rect 4020 2313 4033 2787
rect 4079 2313 4108 2787
rect 4020 2300 4108 2313
rect 4164 2787 4268 2800
rect 4164 2313 4193 2787
rect 4239 2313 4268 2787
rect 4164 2300 4268 2313
rect 4324 2787 4428 2800
rect 4324 2313 4353 2787
rect 4399 2313 4428 2787
rect 4324 2300 4428 2313
rect 4484 2787 4588 2800
rect 4484 2313 4513 2787
rect 4559 2313 4588 2787
rect 4484 2300 4588 2313
rect 4644 2787 4748 2800
rect 4644 2313 4673 2787
rect 4719 2313 4748 2787
rect 4644 2300 4748 2313
rect 4804 2787 4908 2800
rect 4804 2313 4833 2787
rect 4879 2313 4908 2787
rect 4804 2300 4908 2313
rect 4964 2787 5068 2800
rect 4964 2313 4993 2787
rect 5039 2313 5068 2787
rect 4964 2300 5068 2313
rect 5124 2787 5228 2800
rect 5124 2313 5153 2787
rect 5199 2313 5228 2787
rect 5124 2300 5228 2313
rect 5284 2787 5372 2800
rect 5284 2313 5313 2787
rect 5359 2313 5372 2787
rect 5284 2300 5372 2313
rect 5544 2787 5632 2800
rect 5544 2313 5557 2787
rect 5603 2313 5632 2787
rect 5544 2300 5632 2313
rect 5688 2787 5792 2800
rect 5688 2313 5717 2787
rect 5763 2313 5792 2787
rect 5688 2300 5792 2313
rect 5848 2787 5952 2800
rect 5848 2313 5877 2787
rect 5923 2313 5952 2787
rect 5848 2300 5952 2313
rect 6008 2787 6112 2800
rect 6008 2313 6037 2787
rect 6083 2313 6112 2787
rect 6008 2300 6112 2313
rect 6168 2787 6272 2800
rect 6168 2313 6197 2787
rect 6243 2313 6272 2787
rect 6168 2300 6272 2313
rect 6328 2787 6432 2800
rect 6328 2313 6357 2787
rect 6403 2313 6432 2787
rect 6328 2300 6432 2313
rect 6488 2787 6592 2800
rect 6488 2313 6517 2787
rect 6563 2313 6592 2787
rect 6488 2300 6592 2313
rect 6648 2787 6752 2800
rect 6648 2313 6677 2787
rect 6723 2313 6752 2787
rect 6648 2300 6752 2313
rect 6808 2787 6896 2800
rect 6808 2313 6837 2787
rect 6883 2313 6896 2787
rect 6808 2300 6896 2313
rect 6952 2787 7040 2800
rect 6952 2313 6965 2787
rect 7011 2313 7040 2787
rect 6952 2300 7040 2313
rect 7096 2787 7184 2800
rect 7096 2313 7125 2787
rect 7171 2313 7184 2787
rect 7096 2300 7184 2313
rect 7356 2787 7444 2800
rect 7356 2313 7369 2787
rect 7415 2313 7444 2787
rect 7356 2300 7444 2313
rect 7500 2787 7604 2800
rect 7500 2313 7529 2787
rect 7575 2313 7604 2787
rect 7500 2300 7604 2313
rect 7660 2787 7764 2800
rect 7660 2313 7689 2787
rect 7735 2313 7764 2787
rect 7660 2300 7764 2313
rect 7820 2787 7924 2800
rect 7820 2313 7849 2787
rect 7895 2313 7924 2787
rect 7820 2300 7924 2313
rect 7980 2787 8084 2800
rect 7980 2313 8009 2787
rect 8055 2313 8084 2787
rect 7980 2300 8084 2313
rect 8140 2787 8244 2800
rect 8140 2313 8169 2787
rect 8215 2313 8244 2787
rect 8140 2300 8244 2313
rect 8300 2787 8404 2800
rect 8300 2313 8329 2787
rect 8375 2313 8404 2787
rect 8300 2300 8404 2313
rect 8460 2787 8564 2800
rect 8460 2313 8489 2787
rect 8535 2313 8564 2787
rect 8460 2300 8564 2313
rect 8620 2787 8708 2800
rect 8620 2313 8649 2787
rect 8695 2313 8708 2787
rect 8620 2300 8708 2313
rect 8764 2787 8852 2800
rect 8764 2313 8777 2787
rect 8823 2313 8852 2787
rect 8764 2300 8852 2313
rect 8908 2787 8996 2800
rect 8908 2313 8937 2787
rect 8983 2313 8996 2787
rect 8908 2300 8996 2313
rect -1019 2157 -931 2170
rect 108 2151 196 2164
rect -1163 1850 -1075 1863
rect -4406 1805 -4318 1818
rect -4406 1631 -4393 1805
rect -4347 1631 -4318 1805
rect -4406 1618 -4318 1631
rect -4262 1805 -4158 1818
rect -4262 1631 -4233 1805
rect -4187 1631 -4158 1805
rect -4262 1618 -4158 1631
rect -4102 1805 -3998 1818
rect -4102 1631 -4073 1805
rect -4027 1631 -3998 1805
rect -4102 1618 -3998 1631
rect -3942 1805 -3838 1818
rect -3942 1631 -3913 1805
rect -3867 1631 -3838 1805
rect -3942 1618 -3838 1631
rect -3782 1805 -3694 1818
rect -3782 1631 -3753 1805
rect -3707 1631 -3694 1805
rect -3533 1816 -3445 1829
rect -3533 1754 -3520 1816
rect -3474 1754 -3445 1816
rect -3533 1741 -3445 1754
rect -2997 1816 -2909 1829
rect -2997 1754 -2968 1816
rect -2922 1754 -2909 1816
rect -2997 1741 -2909 1754
rect -2747 1816 -2659 1829
rect -2747 1754 -2734 1816
rect -2688 1754 -2659 1816
rect -2747 1741 -2659 1754
rect -2211 1816 -2123 1829
rect -2211 1754 -2182 1816
rect -2136 1754 -2123 1816
rect -2211 1741 -2123 1754
rect -1961 1816 -1873 1829
rect -1961 1754 -1948 1816
rect -1902 1754 -1873 1816
rect -1961 1741 -1873 1754
rect -1425 1816 -1337 1829
rect -1425 1754 -1396 1816
rect -1350 1754 -1337 1816
rect -1425 1741 -1337 1754
rect -3782 1618 -3694 1631
rect -1163 1676 -1150 1850
rect -1104 1676 -1075 1850
rect -1163 1663 -1075 1676
rect -1019 1850 -931 1863
rect -1019 1676 -990 1850
rect -944 1676 -931 1850
rect -1019 1663 -931 1676
rect 108 1677 121 2151
rect 167 1677 196 2151
rect 108 1664 196 1677
rect 252 2151 340 2164
rect 252 1677 281 2151
rect 327 1677 340 2151
rect 252 1664 340 1677
rect 396 2151 484 2164
rect 396 1677 409 2151
rect 455 1677 484 2151
rect 396 1664 484 1677
rect 540 2151 644 2164
rect 540 1677 569 2151
rect 615 1677 644 2151
rect 540 1664 644 1677
rect 700 2151 804 2164
rect 700 1677 729 2151
rect 775 1677 804 2151
rect 700 1664 804 1677
rect 860 2151 964 2164
rect 860 1677 889 2151
rect 935 1677 964 2151
rect 860 1664 964 1677
rect 1020 2151 1124 2164
rect 1020 1677 1049 2151
rect 1095 1677 1124 2151
rect 1020 1664 1124 1677
rect 1180 2151 1284 2164
rect 1180 1677 1209 2151
rect 1255 1677 1284 2151
rect 1180 1664 1284 1677
rect 1340 2151 1444 2164
rect 1340 1677 1369 2151
rect 1415 1677 1444 2151
rect 1340 1664 1444 1677
rect 1500 2151 1604 2164
rect 1500 1677 1529 2151
rect 1575 1677 1604 2151
rect 1500 1664 1604 1677
rect 1660 2151 1748 2164
rect 1660 1677 1689 2151
rect 1735 1677 1748 2151
rect 1660 1664 1748 1677
rect 1920 2151 2008 2164
rect 1920 1677 1933 2151
rect 1979 1677 2008 2151
rect 1920 1664 2008 1677
rect 2064 2151 2168 2164
rect 2064 1677 2093 2151
rect 2139 1677 2168 2151
rect 2064 1664 2168 1677
rect 2224 2151 2328 2164
rect 2224 1677 2253 2151
rect 2299 1677 2328 2151
rect 2224 1664 2328 1677
rect 2384 2151 2488 2164
rect 2384 1677 2413 2151
rect 2459 1677 2488 2151
rect 2384 1664 2488 1677
rect 2544 2151 2648 2164
rect 2544 1677 2573 2151
rect 2619 1677 2648 2151
rect 2544 1664 2648 1677
rect 2704 2151 2808 2164
rect 2704 1677 2733 2151
rect 2779 1677 2808 2151
rect 2704 1664 2808 1677
rect 2864 2151 2968 2164
rect 2864 1677 2893 2151
rect 2939 1677 2968 2151
rect 2864 1664 2968 1677
rect 3024 2151 3128 2164
rect 3024 1677 3053 2151
rect 3099 1677 3128 2151
rect 3024 1664 3128 1677
rect 3184 2151 3272 2164
rect 3184 1677 3213 2151
rect 3259 1677 3272 2151
rect 3184 1664 3272 1677
rect 3328 2151 3416 2164
rect 3328 1677 3341 2151
rect 3387 1677 3416 2151
rect 3328 1664 3416 1677
rect 3472 2151 3560 2164
rect 3472 1677 3501 2151
rect 3547 1677 3560 2151
rect 3472 1664 3560 1677
rect 3732 2151 3820 2164
rect 3732 1677 3745 2151
rect 3791 1677 3820 2151
rect 3732 1664 3820 1677
rect 3876 2151 3964 2164
rect 3876 1677 3905 2151
rect 3951 1677 3964 2151
rect 3876 1664 3964 1677
rect 4020 2151 4108 2164
rect 4020 1677 4033 2151
rect 4079 1677 4108 2151
rect 4020 1664 4108 1677
rect 4164 2151 4268 2164
rect 4164 1677 4193 2151
rect 4239 1677 4268 2151
rect 4164 1664 4268 1677
rect 4324 2151 4428 2164
rect 4324 1677 4353 2151
rect 4399 1677 4428 2151
rect 4324 1664 4428 1677
rect 4484 2151 4588 2164
rect 4484 1677 4513 2151
rect 4559 1677 4588 2151
rect 4484 1664 4588 1677
rect 4644 2151 4748 2164
rect 4644 1677 4673 2151
rect 4719 1677 4748 2151
rect 4644 1664 4748 1677
rect 4804 2151 4908 2164
rect 4804 1677 4833 2151
rect 4879 1677 4908 2151
rect 4804 1664 4908 1677
rect 4964 2151 5068 2164
rect 4964 1677 4993 2151
rect 5039 1677 5068 2151
rect 4964 1664 5068 1677
rect 5124 2151 5228 2164
rect 5124 1677 5153 2151
rect 5199 1677 5228 2151
rect 5124 1664 5228 1677
rect 5284 2151 5372 2164
rect 5284 1677 5313 2151
rect 5359 1677 5372 2151
rect 5284 1664 5372 1677
rect 5544 2151 5632 2164
rect 5544 1677 5557 2151
rect 5603 1677 5632 2151
rect 5544 1664 5632 1677
rect 5688 2151 5792 2164
rect 5688 1677 5717 2151
rect 5763 1677 5792 2151
rect 5688 1664 5792 1677
rect 5848 2151 5952 2164
rect 5848 1677 5877 2151
rect 5923 1677 5952 2151
rect 5848 1664 5952 1677
rect 6008 2151 6112 2164
rect 6008 1677 6037 2151
rect 6083 1677 6112 2151
rect 6008 1664 6112 1677
rect 6168 2151 6272 2164
rect 6168 1677 6197 2151
rect 6243 1677 6272 2151
rect 6168 1664 6272 1677
rect 6328 2151 6432 2164
rect 6328 1677 6357 2151
rect 6403 1677 6432 2151
rect 6328 1664 6432 1677
rect 6488 2151 6592 2164
rect 6488 1677 6517 2151
rect 6563 1677 6592 2151
rect 6488 1664 6592 1677
rect 6648 2151 6752 2164
rect 6648 1677 6677 2151
rect 6723 1677 6752 2151
rect 6648 1664 6752 1677
rect 6808 2151 6896 2164
rect 6808 1677 6837 2151
rect 6883 1677 6896 2151
rect 6808 1664 6896 1677
rect 6952 2151 7040 2164
rect 6952 1677 6965 2151
rect 7011 1677 7040 2151
rect 6952 1664 7040 1677
rect 7096 2151 7184 2164
rect 7096 1677 7125 2151
rect 7171 1677 7184 2151
rect 7096 1664 7184 1677
rect 7356 2151 7444 2164
rect 7356 1677 7369 2151
rect 7415 1677 7444 2151
rect 7356 1664 7444 1677
rect 7500 2151 7604 2164
rect 7500 1677 7529 2151
rect 7575 1677 7604 2151
rect 7500 1664 7604 1677
rect 7660 2151 7764 2164
rect 7660 1677 7689 2151
rect 7735 1677 7764 2151
rect 7660 1664 7764 1677
rect 7820 2151 7924 2164
rect 7820 1677 7849 2151
rect 7895 1677 7924 2151
rect 7820 1664 7924 1677
rect 7980 2151 8084 2164
rect 7980 1677 8009 2151
rect 8055 1677 8084 2151
rect 7980 1664 8084 1677
rect 8140 2151 8244 2164
rect 8140 1677 8169 2151
rect 8215 1677 8244 2151
rect 8140 1664 8244 1677
rect 8300 2151 8404 2164
rect 8300 1677 8329 2151
rect 8375 1677 8404 2151
rect 8300 1664 8404 1677
rect 8460 2151 8564 2164
rect 8460 1677 8489 2151
rect 8535 1677 8564 2151
rect 8460 1664 8564 1677
rect 8620 2151 8708 2164
rect 8620 1677 8649 2151
rect 8695 1677 8708 2151
rect 8620 1664 8708 1677
rect 8764 2151 8852 2164
rect 8764 1677 8777 2151
rect 8823 1677 8852 2151
rect 8764 1664 8852 1677
rect 8908 2151 8996 2164
rect 8908 1677 8937 2151
rect 8983 1677 8996 2151
rect 8908 1664 8996 1677
rect -4406 679 -4318 692
rect -4812 634 -4724 647
rect -4812 460 -4799 634
rect -4753 460 -4724 634
rect -4812 447 -4724 460
rect -4668 634 -4580 647
rect -4668 460 -4639 634
rect -4593 460 -4580 634
rect -4406 505 -4393 679
rect -4347 505 -4318 679
rect -4406 492 -4318 505
rect -4262 679 -4158 692
rect -4262 505 -4233 679
rect -4187 505 -4158 679
rect -4262 492 -4158 505
rect -4102 679 -3998 692
rect -4102 505 -4073 679
rect -4027 505 -3998 679
rect -4102 492 -3998 505
rect -3942 679 -3838 692
rect -3942 505 -3913 679
rect -3867 505 -3838 679
rect -3942 492 -3838 505
rect -3782 679 -3694 692
rect -3782 505 -3753 679
rect -3707 505 -3694 679
rect -1163 634 -1075 647
rect -3782 492 -3694 505
rect -3533 556 -3445 569
rect -3533 494 -3520 556
rect -3474 494 -3445 556
rect -4668 447 -4580 460
rect -3533 481 -3445 494
rect -2997 556 -2909 569
rect -2997 494 -2968 556
rect -2922 494 -2909 556
rect -2997 481 -2909 494
rect -2747 556 -2659 569
rect -2747 494 -2734 556
rect -2688 494 -2659 556
rect -2747 481 -2659 494
rect -2211 556 -2123 569
rect -2211 494 -2182 556
rect -2136 494 -2123 556
rect -2211 481 -2123 494
rect -1961 556 -1873 569
rect -1961 494 -1948 556
rect -1902 494 -1873 556
rect -1961 481 -1873 494
rect -1425 556 -1337 569
rect -1425 494 -1396 556
rect -1350 494 -1337 556
rect -1425 481 -1337 494
rect -1163 460 -1150 634
rect -1104 460 -1075 634
rect -1163 447 -1075 460
rect -1019 634 -931 647
rect -1019 460 -990 634
rect -944 460 -931 634
rect -1019 447 -931 460
rect -4812 140 -4724 153
rect -4812 -34 -4799 140
rect -4753 -34 -4724 140
rect -4812 -47 -4724 -34
rect -4668 140 -4580 153
rect -4668 -34 -4639 140
rect -4593 -34 -4580 140
rect -1163 140 -1075 153
rect -4668 -47 -4580 -34
rect -4406 95 -4318 108
rect -4406 -79 -4393 95
rect -4347 -79 -4318 95
rect -4406 -92 -4318 -79
rect -4262 95 -4158 108
rect -4262 -79 -4233 95
rect -4187 -79 -4158 95
rect -4262 -92 -4158 -79
rect -4102 95 -3998 108
rect -4102 -79 -4073 95
rect -4027 -79 -3998 95
rect -4102 -92 -3998 -79
rect -3942 95 -3838 108
rect -3942 -79 -3913 95
rect -3867 -79 -3838 95
rect -3942 -92 -3838 -79
rect -3782 95 -3694 108
rect -3782 -79 -3753 95
rect -3707 -79 -3694 95
rect -3533 106 -3445 119
rect -3533 44 -3520 106
rect -3474 44 -3445 106
rect -3533 31 -3445 44
rect -2997 106 -2909 119
rect -2997 44 -2968 106
rect -2922 44 -2909 106
rect -2997 31 -2909 44
rect -2747 106 -2659 119
rect -2747 44 -2734 106
rect -2688 44 -2659 106
rect -2747 31 -2659 44
rect -2211 106 -2123 119
rect -2211 44 -2182 106
rect -2136 44 -2123 106
rect -2211 31 -2123 44
rect -1961 106 -1873 119
rect -1961 44 -1948 106
rect -1902 44 -1873 106
rect -1961 31 -1873 44
rect -1425 106 -1337 119
rect -1425 44 -1396 106
rect -1350 44 -1337 106
rect -1425 31 -1337 44
rect -3782 -92 -3694 -79
rect -1163 -34 -1150 140
rect -1104 -34 -1075 140
rect -1163 -47 -1075 -34
rect -1019 140 -931 153
rect -1019 -34 -990 140
rect -944 -34 -931 140
rect -1019 -47 -931 -34
rect -4406 -1031 -4318 -1018
rect -4406 -1205 -4393 -1031
rect -4347 -1205 -4318 -1031
rect -4406 -1218 -4318 -1205
rect -4262 -1031 -4158 -1018
rect -4262 -1205 -4233 -1031
rect -4187 -1205 -4158 -1031
rect -4262 -1218 -4158 -1205
rect -4102 -1031 -3998 -1018
rect -4102 -1205 -4073 -1031
rect -4027 -1205 -3998 -1031
rect -4102 -1218 -3998 -1205
rect -3942 -1031 -3838 -1018
rect -3942 -1205 -3913 -1031
rect -3867 -1205 -3838 -1031
rect -3942 -1218 -3838 -1205
rect -3782 -1031 -3694 -1018
rect -3782 -1205 -3753 -1031
rect -3707 -1205 -3694 -1031
rect -1163 -1076 -1075 -1063
rect -3782 -1218 -3694 -1205
rect -3533 -1154 -3445 -1141
rect -3533 -1216 -3520 -1154
rect -3474 -1216 -3445 -1154
rect -3533 -1229 -3445 -1216
rect -2997 -1154 -2909 -1141
rect -2997 -1216 -2968 -1154
rect -2922 -1216 -2909 -1154
rect -2997 -1229 -2909 -1216
rect -2747 -1154 -2659 -1141
rect -2747 -1216 -2734 -1154
rect -2688 -1216 -2659 -1154
rect -2747 -1229 -2659 -1216
rect -2211 -1154 -2123 -1141
rect -2211 -1216 -2182 -1154
rect -2136 -1216 -2123 -1154
rect -2211 -1229 -2123 -1216
rect -1961 -1154 -1873 -1141
rect -1961 -1216 -1948 -1154
rect -1902 -1216 -1873 -1154
rect -1961 -1229 -1873 -1216
rect -1425 -1154 -1337 -1141
rect -1425 -1216 -1396 -1154
rect -1350 -1216 -1337 -1154
rect -1425 -1229 -1337 -1216
rect -1163 -1250 -1150 -1076
rect -1104 -1250 -1075 -1076
rect -1163 -1263 -1075 -1250
rect -1019 -1076 -931 -1063
rect -1019 -1250 -990 -1076
rect -944 -1250 -931 -1076
rect -1019 -1263 -931 -1250
rect 108 -1565 196 -1552
rect 108 -2039 121 -1565
rect 167 -2039 196 -1565
rect 108 -2052 196 -2039
rect 252 -1565 340 -1552
rect 252 -2039 281 -1565
rect 327 -2039 340 -1565
rect 252 -2052 340 -2039
rect 396 -1565 484 -1552
rect 396 -2039 409 -1565
rect 455 -2039 484 -1565
rect 396 -2052 484 -2039
rect 540 -1565 644 -1552
rect 540 -2039 569 -1565
rect 615 -2039 644 -1565
rect 540 -2052 644 -2039
rect 700 -1565 804 -1552
rect 700 -2039 729 -1565
rect 775 -2039 804 -1565
rect 700 -2052 804 -2039
rect 860 -1565 964 -1552
rect 860 -2039 889 -1565
rect 935 -2039 964 -1565
rect 860 -2052 964 -2039
rect 1020 -1565 1124 -1552
rect 1020 -2039 1049 -1565
rect 1095 -2039 1124 -1565
rect 1020 -2052 1124 -2039
rect 1180 -1565 1284 -1552
rect 1180 -2039 1209 -1565
rect 1255 -2039 1284 -1565
rect 1180 -2052 1284 -2039
rect 1340 -1565 1444 -1552
rect 1340 -2039 1369 -1565
rect 1415 -2039 1444 -1565
rect 1340 -2052 1444 -2039
rect 1500 -1565 1604 -1552
rect 1500 -2039 1529 -1565
rect 1575 -2039 1604 -1565
rect 1500 -2052 1604 -2039
rect 1660 -1565 1748 -1552
rect 1660 -2039 1689 -1565
rect 1735 -2039 1748 -1565
rect 1660 -2052 1748 -2039
rect 1920 -1565 2008 -1552
rect 1920 -2039 1933 -1565
rect 1979 -2039 2008 -1565
rect 1920 -2052 2008 -2039
rect 2064 -1565 2168 -1552
rect 2064 -2039 2093 -1565
rect 2139 -2039 2168 -1565
rect 2064 -2052 2168 -2039
rect 2224 -1565 2328 -1552
rect 2224 -2039 2253 -1565
rect 2299 -2039 2328 -1565
rect 2224 -2052 2328 -2039
rect 2384 -1565 2488 -1552
rect 2384 -2039 2413 -1565
rect 2459 -2039 2488 -1565
rect 2384 -2052 2488 -2039
rect 2544 -1565 2648 -1552
rect 2544 -2039 2573 -1565
rect 2619 -2039 2648 -1565
rect 2544 -2052 2648 -2039
rect 2704 -1565 2808 -1552
rect 2704 -2039 2733 -1565
rect 2779 -2039 2808 -1565
rect 2704 -2052 2808 -2039
rect 2864 -1565 2968 -1552
rect 2864 -2039 2893 -1565
rect 2939 -2039 2968 -1565
rect 2864 -2052 2968 -2039
rect 3024 -1565 3128 -1552
rect 3024 -2039 3053 -1565
rect 3099 -2039 3128 -1565
rect 3024 -2052 3128 -2039
rect 3184 -1565 3272 -1552
rect 3184 -2039 3213 -1565
rect 3259 -2039 3272 -1565
rect 3184 -2052 3272 -2039
rect 3328 -1565 3416 -1552
rect 3328 -2039 3341 -1565
rect 3387 -2039 3416 -1565
rect 3328 -2052 3416 -2039
rect 3472 -1565 3560 -1552
rect 3472 -2039 3501 -1565
rect 3547 -2039 3560 -1565
rect 3472 -2052 3560 -2039
rect 3732 -1565 3820 -1552
rect 3732 -2039 3745 -1565
rect 3791 -2039 3820 -1565
rect 3732 -2052 3820 -2039
rect 3876 -1565 3964 -1552
rect 3876 -2039 3905 -1565
rect 3951 -2039 3964 -1565
rect 3876 -2052 3964 -2039
rect 4020 -1565 4108 -1552
rect 4020 -2039 4033 -1565
rect 4079 -2039 4108 -1565
rect 4020 -2052 4108 -2039
rect 4164 -1565 4268 -1552
rect 4164 -2039 4193 -1565
rect 4239 -2039 4268 -1565
rect 4164 -2052 4268 -2039
rect 4324 -1565 4428 -1552
rect 4324 -2039 4353 -1565
rect 4399 -2039 4428 -1565
rect 4324 -2052 4428 -2039
rect 4484 -1565 4588 -1552
rect 4484 -2039 4513 -1565
rect 4559 -2039 4588 -1565
rect 4484 -2052 4588 -2039
rect 4644 -1565 4748 -1552
rect 4644 -2039 4673 -1565
rect 4719 -2039 4748 -1565
rect 4644 -2052 4748 -2039
rect 4804 -1565 4908 -1552
rect 4804 -2039 4833 -1565
rect 4879 -2039 4908 -1565
rect 4804 -2052 4908 -2039
rect 4964 -1565 5068 -1552
rect 4964 -2039 4993 -1565
rect 5039 -2039 5068 -1565
rect 4964 -2052 5068 -2039
rect 5124 -1565 5228 -1552
rect 5124 -2039 5153 -1565
rect 5199 -2039 5228 -1565
rect 5124 -2052 5228 -2039
rect 5284 -1565 5372 -1552
rect 5284 -2039 5313 -1565
rect 5359 -2039 5372 -1565
rect 5284 -2052 5372 -2039
rect 5544 -1565 5632 -1552
rect 5544 -2039 5557 -1565
rect 5603 -2039 5632 -1565
rect 5544 -2052 5632 -2039
rect 5688 -1565 5792 -1552
rect 5688 -2039 5717 -1565
rect 5763 -2039 5792 -1565
rect 5688 -2052 5792 -2039
rect 5848 -1565 5952 -1552
rect 5848 -2039 5877 -1565
rect 5923 -2039 5952 -1565
rect 5848 -2052 5952 -2039
rect 6008 -1565 6112 -1552
rect 6008 -2039 6037 -1565
rect 6083 -2039 6112 -1565
rect 6008 -2052 6112 -2039
rect 6168 -1565 6272 -1552
rect 6168 -2039 6197 -1565
rect 6243 -2039 6272 -1565
rect 6168 -2052 6272 -2039
rect 6328 -1565 6432 -1552
rect 6328 -2039 6357 -1565
rect 6403 -2039 6432 -1565
rect 6328 -2052 6432 -2039
rect 6488 -1565 6592 -1552
rect 6488 -2039 6517 -1565
rect 6563 -2039 6592 -1565
rect 6488 -2052 6592 -2039
rect 6648 -1565 6752 -1552
rect 6648 -2039 6677 -1565
rect 6723 -2039 6752 -1565
rect 6648 -2052 6752 -2039
rect 6808 -1565 6896 -1552
rect 6808 -2039 6837 -1565
rect 6883 -2039 6896 -1565
rect 6808 -2052 6896 -2039
rect 6952 -1565 7040 -1552
rect 6952 -2039 6965 -1565
rect 7011 -2039 7040 -1565
rect 6952 -2052 7040 -2039
rect 7096 -1565 7184 -1552
rect 7096 -2039 7125 -1565
rect 7171 -2039 7184 -1565
rect 7096 -2052 7184 -2039
rect 7356 -1565 7444 -1552
rect 7356 -2039 7369 -1565
rect 7415 -2039 7444 -1565
rect 7356 -2052 7444 -2039
rect 7500 -1565 7604 -1552
rect 7500 -2039 7529 -1565
rect 7575 -2039 7604 -1565
rect 7500 -2052 7604 -2039
rect 7660 -1565 7764 -1552
rect 7660 -2039 7689 -1565
rect 7735 -2039 7764 -1565
rect 7660 -2052 7764 -2039
rect 7820 -1565 7924 -1552
rect 7820 -2039 7849 -1565
rect 7895 -2039 7924 -1565
rect 7820 -2052 7924 -2039
rect 7980 -1565 8084 -1552
rect 7980 -2039 8009 -1565
rect 8055 -2039 8084 -1565
rect 7980 -2052 8084 -2039
rect 8140 -1565 8244 -1552
rect 8140 -2039 8169 -1565
rect 8215 -2039 8244 -1565
rect 8140 -2052 8244 -2039
rect 8300 -1565 8404 -1552
rect 8300 -2039 8329 -1565
rect 8375 -2039 8404 -1565
rect 8300 -2052 8404 -2039
rect 8460 -1565 8564 -1552
rect 8460 -2039 8489 -1565
rect 8535 -2039 8564 -1565
rect 8460 -2052 8564 -2039
rect 8620 -1565 8708 -1552
rect 8620 -2039 8649 -1565
rect 8695 -2039 8708 -1565
rect 8620 -2052 8708 -2039
rect 8764 -1565 8852 -1552
rect 8764 -2039 8777 -1565
rect 8823 -2039 8852 -1565
rect 8764 -2052 8852 -2039
rect 8908 -1565 8996 -1552
rect 8908 -2039 8937 -1565
rect 8983 -2039 8996 -1565
rect 8908 -2052 8996 -2039
rect 108 -2201 196 -2188
rect 108 -2675 121 -2201
rect 167 -2675 196 -2201
rect 108 -2688 196 -2675
rect 252 -2201 340 -2188
rect 252 -2675 281 -2201
rect 327 -2675 340 -2201
rect 252 -2688 340 -2675
rect 396 -2201 484 -2188
rect 396 -2675 409 -2201
rect 455 -2675 484 -2201
rect 396 -2688 484 -2675
rect 540 -2201 644 -2188
rect 540 -2675 569 -2201
rect 615 -2675 644 -2201
rect 540 -2688 644 -2675
rect 700 -2201 804 -2188
rect 700 -2675 729 -2201
rect 775 -2675 804 -2201
rect 700 -2688 804 -2675
rect 860 -2201 964 -2188
rect 860 -2675 889 -2201
rect 935 -2675 964 -2201
rect 860 -2688 964 -2675
rect 1020 -2201 1124 -2188
rect 1020 -2675 1049 -2201
rect 1095 -2675 1124 -2201
rect 1020 -2688 1124 -2675
rect 1180 -2201 1284 -2188
rect 1180 -2675 1209 -2201
rect 1255 -2675 1284 -2201
rect 1180 -2688 1284 -2675
rect 1340 -2201 1444 -2188
rect 1340 -2675 1369 -2201
rect 1415 -2675 1444 -2201
rect 1340 -2688 1444 -2675
rect 1500 -2201 1604 -2188
rect 1500 -2675 1529 -2201
rect 1575 -2675 1604 -2201
rect 1500 -2688 1604 -2675
rect 1660 -2201 1748 -2188
rect 1660 -2675 1689 -2201
rect 1735 -2675 1748 -2201
rect 1660 -2688 1748 -2675
rect 1920 -2201 2008 -2188
rect 1920 -2675 1933 -2201
rect 1979 -2675 2008 -2201
rect 1920 -2688 2008 -2675
rect 2064 -2201 2168 -2188
rect 2064 -2675 2093 -2201
rect 2139 -2675 2168 -2201
rect 2064 -2688 2168 -2675
rect 2224 -2201 2328 -2188
rect 2224 -2675 2253 -2201
rect 2299 -2675 2328 -2201
rect 2224 -2688 2328 -2675
rect 2384 -2201 2488 -2188
rect 2384 -2675 2413 -2201
rect 2459 -2675 2488 -2201
rect 2384 -2688 2488 -2675
rect 2544 -2201 2648 -2188
rect 2544 -2675 2573 -2201
rect 2619 -2675 2648 -2201
rect 2544 -2688 2648 -2675
rect 2704 -2201 2808 -2188
rect 2704 -2675 2733 -2201
rect 2779 -2675 2808 -2201
rect 2704 -2688 2808 -2675
rect 2864 -2201 2968 -2188
rect 2864 -2675 2893 -2201
rect 2939 -2675 2968 -2201
rect 2864 -2688 2968 -2675
rect 3024 -2201 3128 -2188
rect 3024 -2675 3053 -2201
rect 3099 -2675 3128 -2201
rect 3024 -2688 3128 -2675
rect 3184 -2201 3272 -2188
rect 3184 -2675 3213 -2201
rect 3259 -2675 3272 -2201
rect 3184 -2688 3272 -2675
rect 3328 -2201 3416 -2188
rect 3328 -2675 3341 -2201
rect 3387 -2675 3416 -2201
rect 3328 -2688 3416 -2675
rect 3472 -2201 3560 -2188
rect 3472 -2675 3501 -2201
rect 3547 -2675 3560 -2201
rect 3472 -2688 3560 -2675
rect 3732 -2201 3820 -2188
rect 3732 -2675 3745 -2201
rect 3791 -2675 3820 -2201
rect 3732 -2688 3820 -2675
rect 3876 -2201 3964 -2188
rect 3876 -2675 3905 -2201
rect 3951 -2675 3964 -2201
rect 3876 -2688 3964 -2675
rect 4020 -2201 4108 -2188
rect 4020 -2675 4033 -2201
rect 4079 -2675 4108 -2201
rect 4020 -2688 4108 -2675
rect 4164 -2201 4268 -2188
rect 4164 -2675 4193 -2201
rect 4239 -2675 4268 -2201
rect 4164 -2688 4268 -2675
rect 4324 -2201 4428 -2188
rect 4324 -2675 4353 -2201
rect 4399 -2675 4428 -2201
rect 4324 -2688 4428 -2675
rect 4484 -2201 4588 -2188
rect 4484 -2675 4513 -2201
rect 4559 -2675 4588 -2201
rect 4484 -2688 4588 -2675
rect 4644 -2201 4748 -2188
rect 4644 -2675 4673 -2201
rect 4719 -2675 4748 -2201
rect 4644 -2688 4748 -2675
rect 4804 -2201 4908 -2188
rect 4804 -2675 4833 -2201
rect 4879 -2675 4908 -2201
rect 4804 -2688 4908 -2675
rect 4964 -2201 5068 -2188
rect 4964 -2675 4993 -2201
rect 5039 -2675 5068 -2201
rect 4964 -2688 5068 -2675
rect 5124 -2201 5228 -2188
rect 5124 -2675 5153 -2201
rect 5199 -2675 5228 -2201
rect 5124 -2688 5228 -2675
rect 5284 -2201 5372 -2188
rect 5284 -2675 5313 -2201
rect 5359 -2675 5372 -2201
rect 5284 -2688 5372 -2675
rect 5544 -2201 5632 -2188
rect 5544 -2675 5557 -2201
rect 5603 -2675 5632 -2201
rect 5544 -2688 5632 -2675
rect 5688 -2201 5792 -2188
rect 5688 -2675 5717 -2201
rect 5763 -2675 5792 -2201
rect 5688 -2688 5792 -2675
rect 5848 -2201 5952 -2188
rect 5848 -2675 5877 -2201
rect 5923 -2675 5952 -2201
rect 5848 -2688 5952 -2675
rect 6008 -2201 6112 -2188
rect 6008 -2675 6037 -2201
rect 6083 -2675 6112 -2201
rect 6008 -2688 6112 -2675
rect 6168 -2201 6272 -2188
rect 6168 -2675 6197 -2201
rect 6243 -2675 6272 -2201
rect 6168 -2688 6272 -2675
rect 6328 -2201 6432 -2188
rect 6328 -2675 6357 -2201
rect 6403 -2675 6432 -2201
rect 6328 -2688 6432 -2675
rect 6488 -2201 6592 -2188
rect 6488 -2675 6517 -2201
rect 6563 -2675 6592 -2201
rect 6488 -2688 6592 -2675
rect 6648 -2201 6752 -2188
rect 6648 -2675 6677 -2201
rect 6723 -2675 6752 -2201
rect 6648 -2688 6752 -2675
rect 6808 -2201 6896 -2188
rect 6808 -2675 6837 -2201
rect 6883 -2675 6896 -2201
rect 6808 -2688 6896 -2675
rect 6952 -2201 7040 -2188
rect 6952 -2675 6965 -2201
rect 7011 -2675 7040 -2201
rect 6952 -2688 7040 -2675
rect 7096 -2201 7184 -2188
rect 7096 -2675 7125 -2201
rect 7171 -2675 7184 -2201
rect 7096 -2688 7184 -2675
rect 7356 -2201 7444 -2188
rect 7356 -2675 7369 -2201
rect 7415 -2675 7444 -2201
rect 7356 -2688 7444 -2675
rect 7500 -2201 7604 -2188
rect 7500 -2675 7529 -2201
rect 7575 -2675 7604 -2201
rect 7500 -2688 7604 -2675
rect 7660 -2201 7764 -2188
rect 7660 -2675 7689 -2201
rect 7735 -2675 7764 -2201
rect 7660 -2688 7764 -2675
rect 7820 -2201 7924 -2188
rect 7820 -2675 7849 -2201
rect 7895 -2675 7924 -2201
rect 7820 -2688 7924 -2675
rect 7980 -2201 8084 -2188
rect 7980 -2675 8009 -2201
rect 8055 -2675 8084 -2201
rect 7980 -2688 8084 -2675
rect 8140 -2201 8244 -2188
rect 8140 -2675 8169 -2201
rect 8215 -2675 8244 -2201
rect 8140 -2688 8244 -2675
rect 8300 -2201 8404 -2188
rect 8300 -2675 8329 -2201
rect 8375 -2675 8404 -2201
rect 8300 -2688 8404 -2675
rect 8460 -2201 8564 -2188
rect 8460 -2675 8489 -2201
rect 8535 -2675 8564 -2201
rect 8460 -2688 8564 -2675
rect 8620 -2201 8708 -2188
rect 8620 -2675 8649 -2201
rect 8695 -2675 8708 -2201
rect 8620 -2688 8708 -2675
rect 8764 -2201 8852 -2188
rect 8764 -2675 8777 -2201
rect 8823 -2675 8852 -2201
rect 8764 -2688 8852 -2675
rect 8908 -2201 8996 -2188
rect 8908 -2675 8937 -2201
rect 8983 -2675 8996 -2201
rect 8908 -2688 8996 -2675
rect 108 -2837 196 -2824
rect 108 -3311 121 -2837
rect 167 -3311 196 -2837
rect 108 -3324 196 -3311
rect 252 -2837 340 -2824
rect 252 -3311 281 -2837
rect 327 -3311 340 -2837
rect 252 -3324 340 -3311
rect 396 -2837 484 -2824
rect 396 -3311 409 -2837
rect 455 -3311 484 -2837
rect 396 -3324 484 -3311
rect 540 -2837 644 -2824
rect 540 -3311 569 -2837
rect 615 -3311 644 -2837
rect 540 -3324 644 -3311
rect 700 -2837 804 -2824
rect 700 -3311 729 -2837
rect 775 -3311 804 -2837
rect 700 -3324 804 -3311
rect 860 -2837 964 -2824
rect 860 -3311 889 -2837
rect 935 -3311 964 -2837
rect 860 -3324 964 -3311
rect 1020 -2837 1124 -2824
rect 1020 -3311 1049 -2837
rect 1095 -3311 1124 -2837
rect 1020 -3324 1124 -3311
rect 1180 -2837 1284 -2824
rect 1180 -3311 1209 -2837
rect 1255 -3311 1284 -2837
rect 1180 -3324 1284 -3311
rect 1340 -2837 1444 -2824
rect 1340 -3311 1369 -2837
rect 1415 -3311 1444 -2837
rect 1340 -3324 1444 -3311
rect 1500 -2837 1604 -2824
rect 1500 -3311 1529 -2837
rect 1575 -3311 1604 -2837
rect 1500 -3324 1604 -3311
rect 1660 -2837 1748 -2824
rect 1660 -3311 1689 -2837
rect 1735 -3311 1748 -2837
rect 1660 -3324 1748 -3311
rect 1920 -2837 2008 -2824
rect 1920 -3311 1933 -2837
rect 1979 -3311 2008 -2837
rect 1920 -3324 2008 -3311
rect 2064 -2837 2168 -2824
rect 2064 -3311 2093 -2837
rect 2139 -3311 2168 -2837
rect 2064 -3324 2168 -3311
rect 2224 -2837 2328 -2824
rect 2224 -3311 2253 -2837
rect 2299 -3311 2328 -2837
rect 2224 -3324 2328 -3311
rect 2384 -2837 2488 -2824
rect 2384 -3311 2413 -2837
rect 2459 -3311 2488 -2837
rect 2384 -3324 2488 -3311
rect 2544 -2837 2648 -2824
rect 2544 -3311 2573 -2837
rect 2619 -3311 2648 -2837
rect 2544 -3324 2648 -3311
rect 2704 -2837 2808 -2824
rect 2704 -3311 2733 -2837
rect 2779 -3311 2808 -2837
rect 2704 -3324 2808 -3311
rect 2864 -2837 2968 -2824
rect 2864 -3311 2893 -2837
rect 2939 -3311 2968 -2837
rect 2864 -3324 2968 -3311
rect 3024 -2837 3128 -2824
rect 3024 -3311 3053 -2837
rect 3099 -3311 3128 -2837
rect 3024 -3324 3128 -3311
rect 3184 -2837 3272 -2824
rect 3184 -3311 3213 -2837
rect 3259 -3311 3272 -2837
rect 3184 -3324 3272 -3311
rect 3328 -2837 3416 -2824
rect 3328 -3311 3341 -2837
rect 3387 -3311 3416 -2837
rect 3328 -3324 3416 -3311
rect 3472 -2837 3560 -2824
rect 3472 -3311 3501 -2837
rect 3547 -3311 3560 -2837
rect 3472 -3324 3560 -3311
rect 3732 -2837 3820 -2824
rect 3732 -3311 3745 -2837
rect 3791 -3311 3820 -2837
rect 3732 -3324 3820 -3311
rect 3876 -2837 3964 -2824
rect 3876 -3311 3905 -2837
rect 3951 -3311 3964 -2837
rect 3876 -3324 3964 -3311
rect 4020 -2837 4108 -2824
rect 4020 -3311 4033 -2837
rect 4079 -3311 4108 -2837
rect 4020 -3324 4108 -3311
rect 4164 -2837 4268 -2824
rect 4164 -3311 4193 -2837
rect 4239 -3311 4268 -2837
rect 4164 -3324 4268 -3311
rect 4324 -2837 4428 -2824
rect 4324 -3311 4353 -2837
rect 4399 -3311 4428 -2837
rect 4324 -3324 4428 -3311
rect 4484 -2837 4588 -2824
rect 4484 -3311 4513 -2837
rect 4559 -3311 4588 -2837
rect 4484 -3324 4588 -3311
rect 4644 -2837 4748 -2824
rect 4644 -3311 4673 -2837
rect 4719 -3311 4748 -2837
rect 4644 -3324 4748 -3311
rect 4804 -2837 4908 -2824
rect 4804 -3311 4833 -2837
rect 4879 -3311 4908 -2837
rect 4804 -3324 4908 -3311
rect 4964 -2837 5068 -2824
rect 4964 -3311 4993 -2837
rect 5039 -3311 5068 -2837
rect 4964 -3324 5068 -3311
rect 5124 -2837 5228 -2824
rect 5124 -3311 5153 -2837
rect 5199 -3311 5228 -2837
rect 5124 -3324 5228 -3311
rect 5284 -2837 5372 -2824
rect 5284 -3311 5313 -2837
rect 5359 -3311 5372 -2837
rect 5284 -3324 5372 -3311
rect 5544 -2837 5632 -2824
rect 5544 -3311 5557 -2837
rect 5603 -3311 5632 -2837
rect 5544 -3324 5632 -3311
rect 5688 -2837 5792 -2824
rect 5688 -3311 5717 -2837
rect 5763 -3311 5792 -2837
rect 5688 -3324 5792 -3311
rect 5848 -2837 5952 -2824
rect 5848 -3311 5877 -2837
rect 5923 -3311 5952 -2837
rect 5848 -3324 5952 -3311
rect 6008 -2837 6112 -2824
rect 6008 -3311 6037 -2837
rect 6083 -3311 6112 -2837
rect 6008 -3324 6112 -3311
rect 6168 -2837 6272 -2824
rect 6168 -3311 6197 -2837
rect 6243 -3311 6272 -2837
rect 6168 -3324 6272 -3311
rect 6328 -2837 6432 -2824
rect 6328 -3311 6357 -2837
rect 6403 -3311 6432 -2837
rect 6328 -3324 6432 -3311
rect 6488 -2837 6592 -2824
rect 6488 -3311 6517 -2837
rect 6563 -3311 6592 -2837
rect 6488 -3324 6592 -3311
rect 6648 -2837 6752 -2824
rect 6648 -3311 6677 -2837
rect 6723 -3311 6752 -2837
rect 6648 -3324 6752 -3311
rect 6808 -2837 6896 -2824
rect 6808 -3311 6837 -2837
rect 6883 -3311 6896 -2837
rect 6808 -3324 6896 -3311
rect 6952 -2837 7040 -2824
rect 6952 -3311 6965 -2837
rect 7011 -3311 7040 -2837
rect 6952 -3324 7040 -3311
rect 7096 -2837 7184 -2824
rect 7096 -3311 7125 -2837
rect 7171 -3311 7184 -2837
rect 7096 -3324 7184 -3311
rect 7356 -2837 7444 -2824
rect 7356 -3311 7369 -2837
rect 7415 -3311 7444 -2837
rect 7356 -3324 7444 -3311
rect 7500 -2837 7604 -2824
rect 7500 -3311 7529 -2837
rect 7575 -3311 7604 -2837
rect 7500 -3324 7604 -3311
rect 7660 -2837 7764 -2824
rect 7660 -3311 7689 -2837
rect 7735 -3311 7764 -2837
rect 7660 -3324 7764 -3311
rect 7820 -2837 7924 -2824
rect 7820 -3311 7849 -2837
rect 7895 -3311 7924 -2837
rect 7820 -3324 7924 -3311
rect 7980 -2837 8084 -2824
rect 7980 -3311 8009 -2837
rect 8055 -3311 8084 -2837
rect 7980 -3324 8084 -3311
rect 8140 -2837 8244 -2824
rect 8140 -3311 8169 -2837
rect 8215 -3311 8244 -2837
rect 8140 -3324 8244 -3311
rect 8300 -2837 8404 -2824
rect 8300 -3311 8329 -2837
rect 8375 -3311 8404 -2837
rect 8300 -3324 8404 -3311
rect 8460 -2837 8564 -2824
rect 8460 -3311 8489 -2837
rect 8535 -3311 8564 -2837
rect 8460 -3324 8564 -3311
rect 8620 -2837 8708 -2824
rect 8620 -3311 8649 -2837
rect 8695 -3311 8708 -2837
rect 8620 -3324 8708 -3311
rect 8764 -2837 8852 -2824
rect 8764 -3311 8777 -2837
rect 8823 -3311 8852 -2837
rect 8764 -3324 8852 -3311
rect 8908 -2837 8996 -2824
rect 8908 -3311 8937 -2837
rect 8983 -3311 8996 -2837
rect 8908 -3324 8996 -3311
rect -4089 -3905 -4001 -3892
rect -4089 -4379 -4076 -3905
rect -4030 -4379 -4001 -3905
rect -4089 -4392 -4001 -4379
rect -3945 -3905 -3857 -3892
rect -3945 -4379 -3916 -3905
rect -3870 -4379 -3857 -3905
rect -3945 -4392 -3857 -4379
rect -3801 -3905 -3713 -3892
rect -3801 -4379 -3788 -3905
rect -3742 -4379 -3713 -3905
rect -3801 -4392 -3713 -4379
rect -3657 -3905 -3553 -3892
rect -3657 -4379 -3628 -3905
rect -3582 -4379 -3553 -3905
rect -3657 -4392 -3553 -4379
rect -3497 -3905 -3393 -3892
rect -3497 -4379 -3468 -3905
rect -3422 -4379 -3393 -3905
rect -3497 -4392 -3393 -4379
rect -3337 -3905 -3233 -3892
rect -3337 -4379 -3308 -3905
rect -3262 -4379 -3233 -3905
rect -3337 -4392 -3233 -4379
rect -3177 -3905 -3073 -3892
rect -3177 -4379 -3148 -3905
rect -3102 -4379 -3073 -3905
rect -3177 -4392 -3073 -4379
rect -3017 -3905 -2913 -3892
rect -3017 -4379 -2988 -3905
rect -2942 -4379 -2913 -3905
rect -3017 -4392 -2913 -4379
rect -2857 -3905 -2753 -3892
rect -2857 -4379 -2828 -3905
rect -2782 -4379 -2753 -3905
rect -2857 -4392 -2753 -4379
rect -2697 -3905 -2593 -3892
rect -2697 -4379 -2668 -3905
rect -2622 -4379 -2593 -3905
rect -2697 -4392 -2593 -4379
rect -2537 -3905 -2449 -3892
rect -2537 -4379 -2508 -3905
rect -2462 -4379 -2449 -3905
rect -2537 -4392 -2449 -4379
rect -2277 -3905 -2189 -3892
rect -2277 -4379 -2264 -3905
rect -2218 -4379 -2189 -3905
rect -2277 -4392 -2189 -4379
rect -2133 -3905 -2029 -3892
rect -2133 -4379 -2104 -3905
rect -2058 -4379 -2029 -3905
rect -2133 -4392 -2029 -4379
rect -1973 -3905 -1869 -3892
rect -1973 -4379 -1944 -3905
rect -1898 -4379 -1869 -3905
rect -1973 -4392 -1869 -4379
rect -1813 -3905 -1709 -3892
rect -1813 -4379 -1784 -3905
rect -1738 -4379 -1709 -3905
rect -1813 -4392 -1709 -4379
rect -1653 -3905 -1549 -3892
rect -1653 -4379 -1624 -3905
rect -1578 -4379 -1549 -3905
rect -1653 -4392 -1549 -4379
rect -1493 -3905 -1389 -3892
rect -1493 -4379 -1464 -3905
rect -1418 -4379 -1389 -3905
rect -1493 -4392 -1389 -4379
rect -1333 -3905 -1229 -3892
rect -1333 -4379 -1304 -3905
rect -1258 -4379 -1229 -3905
rect -1333 -4392 -1229 -4379
rect -1173 -3905 -1069 -3892
rect -1173 -4379 -1144 -3905
rect -1098 -4379 -1069 -3905
rect -1173 -4392 -1069 -4379
rect -1013 -3905 -925 -3892
rect -1013 -4379 -984 -3905
rect -938 -4379 -925 -3905
rect -1013 -4392 -925 -4379
rect -869 -3905 -781 -3892
rect -869 -4379 -856 -3905
rect -810 -4379 -781 -3905
rect -869 -4392 -781 -4379
rect -725 -3905 -637 -3892
rect -725 -4379 -696 -3905
rect -650 -4379 -637 -3905
rect -725 -4392 -637 -4379
rect 108 -3905 196 -3892
rect 108 -4379 121 -3905
rect 167 -4379 196 -3905
rect 108 -4392 196 -4379
rect 252 -3905 340 -3892
rect 252 -4379 281 -3905
rect 327 -4379 340 -3905
rect 252 -4392 340 -4379
rect 396 -3905 484 -3892
rect 396 -4379 409 -3905
rect 455 -4379 484 -3905
rect 396 -4392 484 -4379
rect 540 -3905 644 -3892
rect 540 -4379 569 -3905
rect 615 -4379 644 -3905
rect 540 -4392 644 -4379
rect 700 -3905 804 -3892
rect 700 -4379 729 -3905
rect 775 -4379 804 -3905
rect 700 -4392 804 -4379
rect 860 -3905 964 -3892
rect 860 -4379 889 -3905
rect 935 -4379 964 -3905
rect 860 -4392 964 -4379
rect 1020 -3905 1124 -3892
rect 1020 -4379 1049 -3905
rect 1095 -4379 1124 -3905
rect 1020 -4392 1124 -4379
rect 1180 -3905 1284 -3892
rect 1180 -4379 1209 -3905
rect 1255 -4379 1284 -3905
rect 1180 -4392 1284 -4379
rect 1340 -3905 1444 -3892
rect 1340 -4379 1369 -3905
rect 1415 -4379 1444 -3905
rect 1340 -4392 1444 -4379
rect 1500 -3905 1604 -3892
rect 1500 -4379 1529 -3905
rect 1575 -4379 1604 -3905
rect 1500 -4392 1604 -4379
rect 1660 -3905 1748 -3892
rect 1660 -4379 1689 -3905
rect 1735 -4379 1748 -3905
rect 1660 -4392 1748 -4379
rect 1920 -3905 2008 -3892
rect 1920 -4379 1933 -3905
rect 1979 -4379 2008 -3905
rect 1920 -4392 2008 -4379
rect 2064 -3905 2168 -3892
rect 2064 -4379 2093 -3905
rect 2139 -4379 2168 -3905
rect 2064 -4392 2168 -4379
rect 2224 -3905 2328 -3892
rect 2224 -4379 2253 -3905
rect 2299 -4379 2328 -3905
rect 2224 -4392 2328 -4379
rect 2384 -3905 2488 -3892
rect 2384 -4379 2413 -3905
rect 2459 -4379 2488 -3905
rect 2384 -4392 2488 -4379
rect 2544 -3905 2648 -3892
rect 2544 -4379 2573 -3905
rect 2619 -4379 2648 -3905
rect 2544 -4392 2648 -4379
rect 2704 -3905 2808 -3892
rect 2704 -4379 2733 -3905
rect 2779 -4379 2808 -3905
rect 2704 -4392 2808 -4379
rect 2864 -3905 2968 -3892
rect 2864 -4379 2893 -3905
rect 2939 -4379 2968 -3905
rect 2864 -4392 2968 -4379
rect 3024 -3905 3128 -3892
rect 3024 -4379 3053 -3905
rect 3099 -4379 3128 -3905
rect 3024 -4392 3128 -4379
rect 3184 -3905 3272 -3892
rect 3184 -4379 3213 -3905
rect 3259 -4379 3272 -3905
rect 3184 -4392 3272 -4379
rect 3328 -3905 3416 -3892
rect 3328 -4379 3341 -3905
rect 3387 -4379 3416 -3905
rect 3328 -4392 3416 -4379
rect 3472 -3905 3560 -3892
rect 3472 -4379 3501 -3905
rect 3547 -4379 3560 -3905
rect 3472 -4392 3560 -4379
rect 3732 -3905 3820 -3892
rect 3732 -4379 3745 -3905
rect 3791 -4379 3820 -3905
rect 3732 -4392 3820 -4379
rect 3876 -3905 3964 -3892
rect 3876 -4379 3905 -3905
rect 3951 -4379 3964 -3905
rect 3876 -4392 3964 -4379
rect 4020 -3905 4108 -3892
rect 4020 -4379 4033 -3905
rect 4079 -4379 4108 -3905
rect 4020 -4392 4108 -4379
rect 4164 -3905 4268 -3892
rect 4164 -4379 4193 -3905
rect 4239 -4379 4268 -3905
rect 4164 -4392 4268 -4379
rect 4324 -3905 4428 -3892
rect 4324 -4379 4353 -3905
rect 4399 -4379 4428 -3905
rect 4324 -4392 4428 -4379
rect 4484 -3905 4588 -3892
rect 4484 -4379 4513 -3905
rect 4559 -4379 4588 -3905
rect 4484 -4392 4588 -4379
rect 4644 -3905 4748 -3892
rect 4644 -4379 4673 -3905
rect 4719 -4379 4748 -3905
rect 4644 -4392 4748 -4379
rect 4804 -3905 4908 -3892
rect 4804 -4379 4833 -3905
rect 4879 -4379 4908 -3905
rect 4804 -4392 4908 -4379
rect 4964 -3905 5068 -3892
rect 4964 -4379 4993 -3905
rect 5039 -4379 5068 -3905
rect 4964 -4392 5068 -4379
rect 5124 -3905 5228 -3892
rect 5124 -4379 5153 -3905
rect 5199 -4379 5228 -3905
rect 5124 -4392 5228 -4379
rect 5284 -3905 5372 -3892
rect 5284 -4379 5313 -3905
rect 5359 -4379 5372 -3905
rect 5284 -4392 5372 -4379
rect 5544 -3905 5632 -3892
rect 5544 -4379 5557 -3905
rect 5603 -4379 5632 -3905
rect 5544 -4392 5632 -4379
rect 5688 -3905 5792 -3892
rect 5688 -4379 5717 -3905
rect 5763 -4379 5792 -3905
rect 5688 -4392 5792 -4379
rect 5848 -3905 5952 -3892
rect 5848 -4379 5877 -3905
rect 5923 -4379 5952 -3905
rect 5848 -4392 5952 -4379
rect 6008 -3905 6112 -3892
rect 6008 -4379 6037 -3905
rect 6083 -4379 6112 -3905
rect 6008 -4392 6112 -4379
rect 6168 -3905 6272 -3892
rect 6168 -4379 6197 -3905
rect 6243 -4379 6272 -3905
rect 6168 -4392 6272 -4379
rect 6328 -3905 6432 -3892
rect 6328 -4379 6357 -3905
rect 6403 -4379 6432 -3905
rect 6328 -4392 6432 -4379
rect 6488 -3905 6592 -3892
rect 6488 -4379 6517 -3905
rect 6563 -4379 6592 -3905
rect 6488 -4392 6592 -4379
rect 6648 -3905 6752 -3892
rect 6648 -4379 6677 -3905
rect 6723 -4379 6752 -3905
rect 6648 -4392 6752 -4379
rect 6808 -3905 6896 -3892
rect 6808 -4379 6837 -3905
rect 6883 -4379 6896 -3905
rect 6808 -4392 6896 -4379
rect 6952 -3905 7040 -3892
rect 6952 -4379 6965 -3905
rect 7011 -4379 7040 -3905
rect 6952 -4392 7040 -4379
rect 7096 -3905 7184 -3892
rect 7096 -4379 7125 -3905
rect 7171 -4379 7184 -3905
rect 7096 -4392 7184 -4379
rect 7356 -3905 7444 -3892
rect 7356 -4379 7369 -3905
rect 7415 -4379 7444 -3905
rect 7356 -4392 7444 -4379
rect 7500 -3905 7604 -3892
rect 7500 -4379 7529 -3905
rect 7575 -4379 7604 -3905
rect 7500 -4392 7604 -4379
rect 7660 -3905 7764 -3892
rect 7660 -4379 7689 -3905
rect 7735 -4379 7764 -3905
rect 7660 -4392 7764 -4379
rect 7820 -3905 7924 -3892
rect 7820 -4379 7849 -3905
rect 7895 -4379 7924 -3905
rect 7820 -4392 7924 -4379
rect 7980 -3905 8084 -3892
rect 7980 -4379 8009 -3905
rect 8055 -4379 8084 -3905
rect 7980 -4392 8084 -4379
rect 8140 -3905 8244 -3892
rect 8140 -4379 8169 -3905
rect 8215 -4379 8244 -3905
rect 8140 -4392 8244 -4379
rect 8300 -3905 8404 -3892
rect 8300 -4379 8329 -3905
rect 8375 -4379 8404 -3905
rect 8300 -4392 8404 -4379
rect 8460 -3905 8564 -3892
rect 8460 -4379 8489 -3905
rect 8535 -4379 8564 -3905
rect 8460 -4392 8564 -4379
rect 8620 -3905 8708 -3892
rect 8620 -4379 8649 -3905
rect 8695 -4379 8708 -3905
rect 8620 -4392 8708 -4379
rect 8764 -3905 8852 -3892
rect 8764 -4379 8777 -3905
rect 8823 -4379 8852 -3905
rect 8764 -4392 8852 -4379
rect 8908 -3905 8996 -3892
rect 8908 -4379 8937 -3905
rect 8983 -4379 8996 -3905
rect 8908 -4392 8996 -4379
rect -4089 -4541 -4001 -4528
rect -4089 -5015 -4076 -4541
rect -4030 -5015 -4001 -4541
rect -4089 -5028 -4001 -5015
rect -3945 -4541 -3857 -4528
rect -3945 -5015 -3916 -4541
rect -3870 -5015 -3857 -4541
rect -3945 -5028 -3857 -5015
rect -3801 -4541 -3713 -4528
rect -3801 -5015 -3788 -4541
rect -3742 -5015 -3713 -4541
rect -3801 -5028 -3713 -5015
rect -3657 -4541 -3553 -4528
rect -3657 -5015 -3628 -4541
rect -3582 -5015 -3553 -4541
rect -3657 -5028 -3553 -5015
rect -3497 -4541 -3393 -4528
rect -3497 -5015 -3468 -4541
rect -3422 -5015 -3393 -4541
rect -3497 -5028 -3393 -5015
rect -3337 -4541 -3233 -4528
rect -3337 -5015 -3308 -4541
rect -3262 -5015 -3233 -4541
rect -3337 -5028 -3233 -5015
rect -3177 -4541 -3073 -4528
rect -3177 -5015 -3148 -4541
rect -3102 -5015 -3073 -4541
rect -3177 -5028 -3073 -5015
rect -3017 -4541 -2913 -4528
rect -3017 -5015 -2988 -4541
rect -2942 -5015 -2913 -4541
rect -3017 -5028 -2913 -5015
rect -2857 -4541 -2753 -4528
rect -2857 -5015 -2828 -4541
rect -2782 -5015 -2753 -4541
rect -2857 -5028 -2753 -5015
rect -2697 -4541 -2593 -4528
rect -2697 -5015 -2668 -4541
rect -2622 -5015 -2593 -4541
rect -2697 -5028 -2593 -5015
rect -2537 -4541 -2449 -4528
rect -2537 -5015 -2508 -4541
rect -2462 -5015 -2449 -4541
rect -2537 -5028 -2449 -5015
rect -2277 -4541 -2189 -4528
rect -2277 -5015 -2264 -4541
rect -2218 -5015 -2189 -4541
rect -2277 -5028 -2189 -5015
rect -2133 -4541 -2029 -4528
rect -2133 -5015 -2104 -4541
rect -2058 -5015 -2029 -4541
rect -2133 -5028 -2029 -5015
rect -1973 -4541 -1869 -4528
rect -1973 -5015 -1944 -4541
rect -1898 -5015 -1869 -4541
rect -1973 -5028 -1869 -5015
rect -1813 -4541 -1709 -4528
rect -1813 -5015 -1784 -4541
rect -1738 -5015 -1709 -4541
rect -1813 -5028 -1709 -5015
rect -1653 -4541 -1549 -4528
rect -1653 -5015 -1624 -4541
rect -1578 -5015 -1549 -4541
rect -1653 -5028 -1549 -5015
rect -1493 -4541 -1389 -4528
rect -1493 -5015 -1464 -4541
rect -1418 -5015 -1389 -4541
rect -1493 -5028 -1389 -5015
rect -1333 -4541 -1229 -4528
rect -1333 -5015 -1304 -4541
rect -1258 -5015 -1229 -4541
rect -1333 -5028 -1229 -5015
rect -1173 -4541 -1069 -4528
rect -1173 -5015 -1144 -4541
rect -1098 -5015 -1069 -4541
rect -1173 -5028 -1069 -5015
rect -1013 -4541 -925 -4528
rect -1013 -5015 -984 -4541
rect -938 -5015 -925 -4541
rect -1013 -5028 -925 -5015
rect -869 -4541 -781 -4528
rect -869 -5015 -856 -4541
rect -810 -5015 -781 -4541
rect -869 -5028 -781 -5015
rect -725 -4541 -637 -4528
rect -725 -5015 -696 -4541
rect -650 -5015 -637 -4541
rect -725 -5028 -637 -5015
rect 108 -4541 196 -4528
rect 108 -5015 121 -4541
rect 167 -5015 196 -4541
rect 108 -5028 196 -5015
rect 252 -4541 340 -4528
rect 252 -5015 281 -4541
rect 327 -5015 340 -4541
rect 252 -5028 340 -5015
rect 396 -4541 484 -4528
rect 396 -5015 409 -4541
rect 455 -5015 484 -4541
rect 396 -5028 484 -5015
rect 540 -4541 644 -4528
rect 540 -5015 569 -4541
rect 615 -5015 644 -4541
rect 540 -5028 644 -5015
rect 700 -4541 804 -4528
rect 700 -5015 729 -4541
rect 775 -5015 804 -4541
rect 700 -5028 804 -5015
rect 860 -4541 964 -4528
rect 860 -5015 889 -4541
rect 935 -5015 964 -4541
rect 860 -5028 964 -5015
rect 1020 -4541 1124 -4528
rect 1020 -5015 1049 -4541
rect 1095 -5015 1124 -4541
rect 1020 -5028 1124 -5015
rect 1180 -4541 1284 -4528
rect 1180 -5015 1209 -4541
rect 1255 -5015 1284 -4541
rect 1180 -5028 1284 -5015
rect 1340 -4541 1444 -4528
rect 1340 -5015 1369 -4541
rect 1415 -5015 1444 -4541
rect 1340 -5028 1444 -5015
rect 1500 -4541 1604 -4528
rect 1500 -5015 1529 -4541
rect 1575 -5015 1604 -4541
rect 1500 -5028 1604 -5015
rect 1660 -4541 1748 -4528
rect 1660 -5015 1689 -4541
rect 1735 -5015 1748 -4541
rect 1660 -5028 1748 -5015
rect 1920 -4541 2008 -4528
rect 1920 -5015 1933 -4541
rect 1979 -5015 2008 -4541
rect 1920 -5028 2008 -5015
rect 2064 -4541 2168 -4528
rect 2064 -5015 2093 -4541
rect 2139 -5015 2168 -4541
rect 2064 -5028 2168 -5015
rect 2224 -4541 2328 -4528
rect 2224 -5015 2253 -4541
rect 2299 -5015 2328 -4541
rect 2224 -5028 2328 -5015
rect 2384 -4541 2488 -4528
rect 2384 -5015 2413 -4541
rect 2459 -5015 2488 -4541
rect 2384 -5028 2488 -5015
rect 2544 -4541 2648 -4528
rect 2544 -5015 2573 -4541
rect 2619 -5015 2648 -4541
rect 2544 -5028 2648 -5015
rect 2704 -4541 2808 -4528
rect 2704 -5015 2733 -4541
rect 2779 -5015 2808 -4541
rect 2704 -5028 2808 -5015
rect 2864 -4541 2968 -4528
rect 2864 -5015 2893 -4541
rect 2939 -5015 2968 -4541
rect 2864 -5028 2968 -5015
rect 3024 -4541 3128 -4528
rect 3024 -5015 3053 -4541
rect 3099 -5015 3128 -4541
rect 3024 -5028 3128 -5015
rect 3184 -4541 3272 -4528
rect 3184 -5015 3213 -4541
rect 3259 -5015 3272 -4541
rect 3184 -5028 3272 -5015
rect 3328 -4541 3416 -4528
rect 3328 -5015 3341 -4541
rect 3387 -5015 3416 -4541
rect 3328 -5028 3416 -5015
rect 3472 -4541 3560 -4528
rect 3472 -5015 3501 -4541
rect 3547 -5015 3560 -4541
rect 3472 -5028 3560 -5015
rect 3732 -4541 3820 -4528
rect 3732 -5015 3745 -4541
rect 3791 -5015 3820 -4541
rect 3732 -5028 3820 -5015
rect 3876 -4541 3964 -4528
rect 3876 -5015 3905 -4541
rect 3951 -5015 3964 -4541
rect 3876 -5028 3964 -5015
rect 4020 -4541 4108 -4528
rect 4020 -5015 4033 -4541
rect 4079 -5015 4108 -4541
rect 4020 -5028 4108 -5015
rect 4164 -4541 4268 -4528
rect 4164 -5015 4193 -4541
rect 4239 -5015 4268 -4541
rect 4164 -5028 4268 -5015
rect 4324 -4541 4428 -4528
rect 4324 -5015 4353 -4541
rect 4399 -5015 4428 -4541
rect 4324 -5028 4428 -5015
rect 4484 -4541 4588 -4528
rect 4484 -5015 4513 -4541
rect 4559 -5015 4588 -4541
rect 4484 -5028 4588 -5015
rect 4644 -4541 4748 -4528
rect 4644 -5015 4673 -4541
rect 4719 -5015 4748 -4541
rect 4644 -5028 4748 -5015
rect 4804 -4541 4908 -4528
rect 4804 -5015 4833 -4541
rect 4879 -5015 4908 -4541
rect 4804 -5028 4908 -5015
rect 4964 -4541 5068 -4528
rect 4964 -5015 4993 -4541
rect 5039 -5015 5068 -4541
rect 4964 -5028 5068 -5015
rect 5124 -4541 5228 -4528
rect 5124 -5015 5153 -4541
rect 5199 -5015 5228 -4541
rect 5124 -5028 5228 -5015
rect 5284 -4541 5372 -4528
rect 5284 -5015 5313 -4541
rect 5359 -5015 5372 -4541
rect 5284 -5028 5372 -5015
rect 5544 -4541 5632 -4528
rect 5544 -5015 5557 -4541
rect 5603 -5015 5632 -4541
rect 5544 -5028 5632 -5015
rect 5688 -4541 5792 -4528
rect 5688 -5015 5717 -4541
rect 5763 -5015 5792 -4541
rect 5688 -5028 5792 -5015
rect 5848 -4541 5952 -4528
rect 5848 -5015 5877 -4541
rect 5923 -5015 5952 -4541
rect 5848 -5028 5952 -5015
rect 6008 -4541 6112 -4528
rect 6008 -5015 6037 -4541
rect 6083 -5015 6112 -4541
rect 6008 -5028 6112 -5015
rect 6168 -4541 6272 -4528
rect 6168 -5015 6197 -4541
rect 6243 -5015 6272 -4541
rect 6168 -5028 6272 -5015
rect 6328 -4541 6432 -4528
rect 6328 -5015 6357 -4541
rect 6403 -5015 6432 -4541
rect 6328 -5028 6432 -5015
rect 6488 -4541 6592 -4528
rect 6488 -5015 6517 -4541
rect 6563 -5015 6592 -4541
rect 6488 -5028 6592 -5015
rect 6648 -4541 6752 -4528
rect 6648 -5015 6677 -4541
rect 6723 -5015 6752 -4541
rect 6648 -5028 6752 -5015
rect 6808 -4541 6896 -4528
rect 6808 -5015 6837 -4541
rect 6883 -5015 6896 -4541
rect 6808 -5028 6896 -5015
rect 6952 -4541 7040 -4528
rect 6952 -5015 6965 -4541
rect 7011 -5015 7040 -4541
rect 6952 -5028 7040 -5015
rect 7096 -4541 7184 -4528
rect 7096 -5015 7125 -4541
rect 7171 -5015 7184 -4541
rect 7096 -5028 7184 -5015
rect 7356 -4541 7444 -4528
rect 7356 -5015 7369 -4541
rect 7415 -5015 7444 -4541
rect 7356 -5028 7444 -5015
rect 7500 -4541 7604 -4528
rect 7500 -5015 7529 -4541
rect 7575 -5015 7604 -4541
rect 7500 -5028 7604 -5015
rect 7660 -4541 7764 -4528
rect 7660 -5015 7689 -4541
rect 7735 -5015 7764 -4541
rect 7660 -5028 7764 -5015
rect 7820 -4541 7924 -4528
rect 7820 -5015 7849 -4541
rect 7895 -5015 7924 -4541
rect 7820 -5028 7924 -5015
rect 7980 -4541 8084 -4528
rect 7980 -5015 8009 -4541
rect 8055 -5015 8084 -4541
rect 7980 -5028 8084 -5015
rect 8140 -4541 8244 -4528
rect 8140 -5015 8169 -4541
rect 8215 -5015 8244 -4541
rect 8140 -5028 8244 -5015
rect 8300 -4541 8404 -4528
rect 8300 -5015 8329 -4541
rect 8375 -5015 8404 -4541
rect 8300 -5028 8404 -5015
rect 8460 -4541 8564 -4528
rect 8460 -5015 8489 -4541
rect 8535 -5015 8564 -4541
rect 8460 -5028 8564 -5015
rect 8620 -4541 8708 -4528
rect 8620 -5015 8649 -4541
rect 8695 -5015 8708 -4541
rect 8620 -5028 8708 -5015
rect 8764 -4541 8852 -4528
rect 8764 -5015 8777 -4541
rect 8823 -5015 8852 -4541
rect 8764 -5028 8852 -5015
rect 8908 -4541 8996 -4528
rect 8908 -5015 8937 -4541
rect 8983 -5015 8996 -4541
rect 8908 -5028 8996 -5015
rect -4089 -5177 -4001 -5164
rect -4089 -5651 -4076 -5177
rect -4030 -5651 -4001 -5177
rect -4089 -5664 -4001 -5651
rect -3945 -5177 -3857 -5164
rect -3945 -5651 -3916 -5177
rect -3870 -5651 -3857 -5177
rect -3945 -5664 -3857 -5651
rect -3801 -5177 -3713 -5164
rect -3801 -5651 -3788 -5177
rect -3742 -5651 -3713 -5177
rect -3801 -5664 -3713 -5651
rect -3657 -5177 -3553 -5164
rect -3657 -5651 -3628 -5177
rect -3582 -5651 -3553 -5177
rect -3657 -5664 -3553 -5651
rect -3497 -5177 -3393 -5164
rect -3497 -5651 -3468 -5177
rect -3422 -5651 -3393 -5177
rect -3497 -5664 -3393 -5651
rect -3337 -5177 -3233 -5164
rect -3337 -5651 -3308 -5177
rect -3262 -5651 -3233 -5177
rect -3337 -5664 -3233 -5651
rect -3177 -5177 -3073 -5164
rect -3177 -5651 -3148 -5177
rect -3102 -5651 -3073 -5177
rect -3177 -5664 -3073 -5651
rect -3017 -5177 -2913 -5164
rect -3017 -5651 -2988 -5177
rect -2942 -5651 -2913 -5177
rect -3017 -5664 -2913 -5651
rect -2857 -5177 -2753 -5164
rect -2857 -5651 -2828 -5177
rect -2782 -5651 -2753 -5177
rect -2857 -5664 -2753 -5651
rect -2697 -5177 -2593 -5164
rect -2697 -5651 -2668 -5177
rect -2622 -5651 -2593 -5177
rect -2697 -5664 -2593 -5651
rect -2537 -5177 -2449 -5164
rect -2537 -5651 -2508 -5177
rect -2462 -5651 -2449 -5177
rect -2537 -5664 -2449 -5651
rect -2277 -5177 -2189 -5164
rect -2277 -5651 -2264 -5177
rect -2218 -5651 -2189 -5177
rect -2277 -5664 -2189 -5651
rect -2133 -5177 -2029 -5164
rect -2133 -5651 -2104 -5177
rect -2058 -5651 -2029 -5177
rect -2133 -5664 -2029 -5651
rect -1973 -5177 -1869 -5164
rect -1973 -5651 -1944 -5177
rect -1898 -5651 -1869 -5177
rect -1973 -5664 -1869 -5651
rect -1813 -5177 -1709 -5164
rect -1813 -5651 -1784 -5177
rect -1738 -5651 -1709 -5177
rect -1813 -5664 -1709 -5651
rect -1653 -5177 -1549 -5164
rect -1653 -5651 -1624 -5177
rect -1578 -5651 -1549 -5177
rect -1653 -5664 -1549 -5651
rect -1493 -5177 -1389 -5164
rect -1493 -5651 -1464 -5177
rect -1418 -5651 -1389 -5177
rect -1493 -5664 -1389 -5651
rect -1333 -5177 -1229 -5164
rect -1333 -5651 -1304 -5177
rect -1258 -5651 -1229 -5177
rect -1333 -5664 -1229 -5651
rect -1173 -5177 -1069 -5164
rect -1173 -5651 -1144 -5177
rect -1098 -5651 -1069 -5177
rect -1173 -5664 -1069 -5651
rect -1013 -5177 -925 -5164
rect -1013 -5651 -984 -5177
rect -938 -5651 -925 -5177
rect -1013 -5664 -925 -5651
rect -869 -5177 -781 -5164
rect -869 -5651 -856 -5177
rect -810 -5651 -781 -5177
rect -869 -5664 -781 -5651
rect -725 -5177 -637 -5164
rect -725 -5651 -696 -5177
rect -650 -5651 -637 -5177
rect -725 -5664 -637 -5651
rect 108 -5177 196 -5164
rect 108 -5651 121 -5177
rect 167 -5651 196 -5177
rect 108 -5664 196 -5651
rect 252 -5177 340 -5164
rect 252 -5651 281 -5177
rect 327 -5651 340 -5177
rect 252 -5664 340 -5651
rect 396 -5177 484 -5164
rect 396 -5651 409 -5177
rect 455 -5651 484 -5177
rect 396 -5664 484 -5651
rect 540 -5177 644 -5164
rect 540 -5651 569 -5177
rect 615 -5651 644 -5177
rect 540 -5664 644 -5651
rect 700 -5177 804 -5164
rect 700 -5651 729 -5177
rect 775 -5651 804 -5177
rect 700 -5664 804 -5651
rect 860 -5177 964 -5164
rect 860 -5651 889 -5177
rect 935 -5651 964 -5177
rect 860 -5664 964 -5651
rect 1020 -5177 1124 -5164
rect 1020 -5651 1049 -5177
rect 1095 -5651 1124 -5177
rect 1020 -5664 1124 -5651
rect 1180 -5177 1284 -5164
rect 1180 -5651 1209 -5177
rect 1255 -5651 1284 -5177
rect 1180 -5664 1284 -5651
rect 1340 -5177 1444 -5164
rect 1340 -5651 1369 -5177
rect 1415 -5651 1444 -5177
rect 1340 -5664 1444 -5651
rect 1500 -5177 1604 -5164
rect 1500 -5651 1529 -5177
rect 1575 -5651 1604 -5177
rect 1500 -5664 1604 -5651
rect 1660 -5177 1748 -5164
rect 1660 -5651 1689 -5177
rect 1735 -5651 1748 -5177
rect 1660 -5664 1748 -5651
rect 1920 -5177 2008 -5164
rect 1920 -5651 1933 -5177
rect 1979 -5651 2008 -5177
rect 1920 -5664 2008 -5651
rect 2064 -5177 2168 -5164
rect 2064 -5651 2093 -5177
rect 2139 -5651 2168 -5177
rect 2064 -5664 2168 -5651
rect 2224 -5177 2328 -5164
rect 2224 -5651 2253 -5177
rect 2299 -5651 2328 -5177
rect 2224 -5664 2328 -5651
rect 2384 -5177 2488 -5164
rect 2384 -5651 2413 -5177
rect 2459 -5651 2488 -5177
rect 2384 -5664 2488 -5651
rect 2544 -5177 2648 -5164
rect 2544 -5651 2573 -5177
rect 2619 -5651 2648 -5177
rect 2544 -5664 2648 -5651
rect 2704 -5177 2808 -5164
rect 2704 -5651 2733 -5177
rect 2779 -5651 2808 -5177
rect 2704 -5664 2808 -5651
rect 2864 -5177 2968 -5164
rect 2864 -5651 2893 -5177
rect 2939 -5651 2968 -5177
rect 2864 -5664 2968 -5651
rect 3024 -5177 3128 -5164
rect 3024 -5651 3053 -5177
rect 3099 -5651 3128 -5177
rect 3024 -5664 3128 -5651
rect 3184 -5177 3272 -5164
rect 3184 -5651 3213 -5177
rect 3259 -5651 3272 -5177
rect 3184 -5664 3272 -5651
rect 3328 -5177 3416 -5164
rect 3328 -5651 3341 -5177
rect 3387 -5651 3416 -5177
rect 3328 -5664 3416 -5651
rect 3472 -5177 3560 -5164
rect 3472 -5651 3501 -5177
rect 3547 -5651 3560 -5177
rect 3472 -5664 3560 -5651
rect 3732 -5177 3820 -5164
rect 3732 -5651 3745 -5177
rect 3791 -5651 3820 -5177
rect 3732 -5664 3820 -5651
rect 3876 -5177 3964 -5164
rect 3876 -5651 3905 -5177
rect 3951 -5651 3964 -5177
rect 3876 -5664 3964 -5651
rect 4020 -5177 4108 -5164
rect 4020 -5651 4033 -5177
rect 4079 -5651 4108 -5177
rect 4020 -5664 4108 -5651
rect 4164 -5177 4268 -5164
rect 4164 -5651 4193 -5177
rect 4239 -5651 4268 -5177
rect 4164 -5664 4268 -5651
rect 4324 -5177 4428 -5164
rect 4324 -5651 4353 -5177
rect 4399 -5651 4428 -5177
rect 4324 -5664 4428 -5651
rect 4484 -5177 4588 -5164
rect 4484 -5651 4513 -5177
rect 4559 -5651 4588 -5177
rect 4484 -5664 4588 -5651
rect 4644 -5177 4748 -5164
rect 4644 -5651 4673 -5177
rect 4719 -5651 4748 -5177
rect 4644 -5664 4748 -5651
rect 4804 -5177 4908 -5164
rect 4804 -5651 4833 -5177
rect 4879 -5651 4908 -5177
rect 4804 -5664 4908 -5651
rect 4964 -5177 5068 -5164
rect 4964 -5651 4993 -5177
rect 5039 -5651 5068 -5177
rect 4964 -5664 5068 -5651
rect 5124 -5177 5228 -5164
rect 5124 -5651 5153 -5177
rect 5199 -5651 5228 -5177
rect 5124 -5664 5228 -5651
rect 5284 -5177 5372 -5164
rect 5284 -5651 5313 -5177
rect 5359 -5651 5372 -5177
rect 5284 -5664 5372 -5651
rect 5544 -5177 5632 -5164
rect 5544 -5651 5557 -5177
rect 5603 -5651 5632 -5177
rect 5544 -5664 5632 -5651
rect 5688 -5177 5792 -5164
rect 5688 -5651 5717 -5177
rect 5763 -5651 5792 -5177
rect 5688 -5664 5792 -5651
rect 5848 -5177 5952 -5164
rect 5848 -5651 5877 -5177
rect 5923 -5651 5952 -5177
rect 5848 -5664 5952 -5651
rect 6008 -5177 6112 -5164
rect 6008 -5651 6037 -5177
rect 6083 -5651 6112 -5177
rect 6008 -5664 6112 -5651
rect 6168 -5177 6272 -5164
rect 6168 -5651 6197 -5177
rect 6243 -5651 6272 -5177
rect 6168 -5664 6272 -5651
rect 6328 -5177 6432 -5164
rect 6328 -5651 6357 -5177
rect 6403 -5651 6432 -5177
rect 6328 -5664 6432 -5651
rect 6488 -5177 6592 -5164
rect 6488 -5651 6517 -5177
rect 6563 -5651 6592 -5177
rect 6488 -5664 6592 -5651
rect 6648 -5177 6752 -5164
rect 6648 -5651 6677 -5177
rect 6723 -5651 6752 -5177
rect 6648 -5664 6752 -5651
rect 6808 -5177 6896 -5164
rect 6808 -5651 6837 -5177
rect 6883 -5651 6896 -5177
rect 6808 -5664 6896 -5651
rect 6952 -5177 7040 -5164
rect 6952 -5651 6965 -5177
rect 7011 -5651 7040 -5177
rect 6952 -5664 7040 -5651
rect 7096 -5177 7184 -5164
rect 7096 -5651 7125 -5177
rect 7171 -5651 7184 -5177
rect 7096 -5664 7184 -5651
rect 7356 -5177 7444 -5164
rect 7356 -5651 7369 -5177
rect 7415 -5651 7444 -5177
rect 7356 -5664 7444 -5651
rect 7500 -5177 7604 -5164
rect 7500 -5651 7529 -5177
rect 7575 -5651 7604 -5177
rect 7500 -5664 7604 -5651
rect 7660 -5177 7764 -5164
rect 7660 -5651 7689 -5177
rect 7735 -5651 7764 -5177
rect 7660 -5664 7764 -5651
rect 7820 -5177 7924 -5164
rect 7820 -5651 7849 -5177
rect 7895 -5651 7924 -5177
rect 7820 -5664 7924 -5651
rect 7980 -5177 8084 -5164
rect 7980 -5651 8009 -5177
rect 8055 -5651 8084 -5177
rect 7980 -5664 8084 -5651
rect 8140 -5177 8244 -5164
rect 8140 -5651 8169 -5177
rect 8215 -5651 8244 -5177
rect 8140 -5664 8244 -5651
rect 8300 -5177 8404 -5164
rect 8300 -5651 8329 -5177
rect 8375 -5651 8404 -5177
rect 8300 -5664 8404 -5651
rect 8460 -5177 8564 -5164
rect 8460 -5651 8489 -5177
rect 8535 -5651 8564 -5177
rect 8460 -5664 8564 -5651
rect 8620 -5177 8708 -5164
rect 8620 -5651 8649 -5177
rect 8695 -5651 8708 -5177
rect 8620 -5664 8708 -5651
rect 8764 -5177 8852 -5164
rect 8764 -5651 8777 -5177
rect 8823 -5651 8852 -5177
rect 8764 -5664 8852 -5651
rect 8908 -5177 8996 -5164
rect 8908 -5651 8937 -5177
rect 8983 -5651 8996 -5177
rect 8908 -5664 8996 -5651
<< ndiffc >>
rect 121 6863 167 7087
rect 281 6863 327 7087
rect 441 6863 487 7087
rect 601 6863 647 7087
rect 761 6863 807 7087
rect 921 6863 967 7087
rect 1081 6863 1127 7087
rect 1241 6863 1287 7087
rect 1401 6863 1447 7087
rect 1529 6863 1575 7087
rect 1689 6863 1735 7087
rect 1933 6863 1979 7087
rect 2093 6863 2139 7087
rect 2221 6863 2267 7087
rect 2381 6863 2427 7087
rect 2541 6863 2587 7087
rect 2701 6863 2747 7087
rect 2861 6863 2907 7087
rect 3021 6863 3067 7087
rect 3181 6863 3227 7087
rect 3341 6863 3387 7087
rect 3501 6863 3547 7087
rect 3745 6863 3791 7087
rect 3905 6863 3951 7087
rect 4033 6863 4079 7087
rect 4193 6863 4239 7087
rect 4353 6863 4399 7087
rect 4513 6863 4559 7087
rect 4673 6863 4719 7087
rect 4833 6863 4879 7087
rect 4993 6863 5039 7087
rect 5153 6863 5199 7087
rect 5313 6863 5359 7087
rect 5557 6863 5603 7087
rect 5717 6863 5763 7087
rect 5845 6863 5891 7087
rect 6005 6863 6051 7087
rect 6165 6863 6211 7087
rect 6325 6863 6371 7087
rect 6485 6863 6531 7087
rect 6645 6863 6691 7087
rect 6805 6863 6851 7087
rect 6965 6863 7011 7087
rect 7125 6863 7171 7087
rect 7369 6863 7415 7087
rect 7529 6863 7575 7087
rect 7657 6863 7703 7087
rect 7817 6863 7863 7087
rect 7977 6863 8023 7087
rect 8137 6863 8183 7087
rect 8297 6863 8343 7087
rect 8457 6863 8503 7087
rect 8617 6863 8663 7087
rect 8777 6863 8823 7087
rect 8937 6863 8983 7087
rect 121 6477 167 6701
rect 281 6477 327 6701
rect 441 6477 487 6701
rect 601 6477 647 6701
rect 761 6477 807 6701
rect 921 6477 967 6701
rect 1081 6477 1127 6701
rect 1241 6477 1287 6701
rect 1401 6477 1447 6701
rect 1529 6477 1575 6701
rect 1689 6477 1735 6701
rect 1933 6477 1979 6701
rect 2093 6477 2139 6701
rect 2221 6477 2267 6701
rect 2381 6477 2427 6701
rect 2541 6477 2587 6701
rect 2701 6477 2747 6701
rect 2861 6477 2907 6701
rect 3021 6477 3067 6701
rect 3181 6477 3227 6701
rect 3341 6477 3387 6701
rect 3501 6477 3547 6701
rect 3745 6477 3791 6701
rect 3905 6477 3951 6701
rect 4033 6477 4079 6701
rect 4193 6477 4239 6701
rect 4353 6477 4399 6701
rect 4513 6477 4559 6701
rect 4673 6477 4719 6701
rect 4833 6477 4879 6701
rect 4993 6477 5039 6701
rect 5153 6477 5199 6701
rect 5313 6477 5359 6701
rect 5557 6477 5603 6701
rect 5717 6477 5763 6701
rect 5845 6477 5891 6701
rect 6005 6477 6051 6701
rect 6165 6477 6211 6701
rect 6325 6477 6371 6701
rect 6485 6477 6531 6701
rect 6645 6477 6691 6701
rect 6805 6477 6851 6701
rect 6965 6477 7011 6701
rect 7125 6477 7171 6701
rect 7369 6477 7415 6701
rect 7529 6477 7575 6701
rect 7657 6477 7703 6701
rect 7817 6477 7863 6701
rect 7977 6477 8023 6701
rect 8137 6477 8183 6701
rect 8297 6477 8343 6701
rect 8457 6477 8503 6701
rect 8617 6477 8663 6701
rect 8777 6477 8823 6701
rect 8937 6477 8983 6701
rect 121 6091 167 6315
rect 281 6091 327 6315
rect 441 6091 487 6315
rect 601 6091 647 6315
rect 761 6091 807 6315
rect 921 6091 967 6315
rect 1081 6091 1127 6315
rect 1241 6091 1287 6315
rect 1401 6091 1447 6315
rect 1529 6091 1575 6315
rect 1689 6091 1735 6315
rect 1933 6091 1979 6315
rect 2093 6091 2139 6315
rect 2221 6091 2267 6315
rect 2381 6091 2427 6315
rect 2541 6091 2587 6315
rect 2701 6091 2747 6315
rect 2861 6091 2907 6315
rect 3021 6091 3067 6315
rect 3181 6091 3227 6315
rect 3341 6091 3387 6315
rect 3501 6091 3547 6315
rect 3745 6091 3791 6315
rect 3905 6091 3951 6315
rect 4033 6091 4079 6315
rect 4193 6091 4239 6315
rect 4353 6091 4399 6315
rect 4513 6091 4559 6315
rect 4673 6091 4719 6315
rect 4833 6091 4879 6315
rect 4993 6091 5039 6315
rect 5153 6091 5199 6315
rect 5313 6091 5359 6315
rect 5557 6091 5603 6315
rect 5717 6091 5763 6315
rect 5845 6091 5891 6315
rect 6005 6091 6051 6315
rect 6165 6091 6211 6315
rect 6325 6091 6371 6315
rect 6485 6091 6531 6315
rect 6645 6091 6691 6315
rect 6805 6091 6851 6315
rect 6965 6091 7011 6315
rect 7125 6091 7171 6315
rect 7369 6091 7415 6315
rect 7529 6091 7575 6315
rect 7657 6091 7703 6315
rect 7817 6091 7863 6315
rect 7977 6091 8023 6315
rect 8137 6091 8183 6315
rect 8297 6091 8343 6315
rect 8457 6091 8503 6315
rect 8617 6091 8663 6315
rect 8777 6091 8823 6315
rect 8937 6091 8983 6315
rect -4799 3014 -4753 3088
rect -4639 3014 -4593 3088
rect -4233 3002 -4187 3076
rect -4073 3002 -4027 3076
rect -3913 3002 -3867 3076
rect -3528 2990 -3482 3036
rect -2968 2990 -2922 3036
rect -2742 2990 -2696 3036
rect -2182 2990 -2136 3036
rect -1956 2990 -1910 3036
rect -1396 2990 -1350 3036
rect -1150 3014 -1104 3088
rect -990 3014 -944 3088
rect -4233 2654 -4187 2728
rect -4073 2654 -4027 2728
rect -3913 2654 -3867 2728
rect -3528 2694 -3482 2740
rect -2968 2694 -2922 2740
rect -2742 2694 -2696 2740
rect -2182 2694 -2136 2740
rect -1956 2694 -1910 2740
rect -1396 2694 -1350 2740
rect -1150 2642 -1104 2716
rect -990 2642 -944 2716
rect -4233 1292 -4187 1366
rect -4073 1292 -4027 1366
rect -3913 1292 -3867 1366
rect -3528 1280 -3482 1326
rect -2968 1280 -2922 1326
rect -2742 1280 -2696 1326
rect -2182 1280 -2136 1326
rect -1956 1280 -1910 1326
rect -1396 1280 -1350 1326
rect -1150 1304 -1104 1378
rect -990 1304 -944 1378
rect 121 1125 167 1349
rect 281 1125 327 1349
rect 409 1125 455 1349
rect 569 1125 615 1349
rect 729 1125 775 1349
rect 889 1125 935 1349
rect 1049 1125 1095 1349
rect 1209 1125 1255 1349
rect 1369 1125 1415 1349
rect 1529 1125 1575 1349
rect 1689 1125 1735 1349
rect 1933 1125 1979 1349
rect 2093 1125 2139 1349
rect 2253 1125 2299 1349
rect 2413 1125 2459 1349
rect 2573 1125 2619 1349
rect 2733 1125 2779 1349
rect 2893 1125 2939 1349
rect 3053 1125 3099 1349
rect 3213 1125 3259 1349
rect 3341 1125 3387 1349
rect 3501 1125 3547 1349
rect 3745 1125 3791 1349
rect 3905 1125 3951 1349
rect 4033 1125 4079 1349
rect 4193 1125 4239 1349
rect 4353 1125 4399 1349
rect 4513 1125 4559 1349
rect 4673 1125 4719 1349
rect 4833 1125 4879 1349
rect 4993 1125 5039 1349
rect 5153 1125 5199 1349
rect 5313 1125 5359 1349
rect 5557 1125 5603 1349
rect 5717 1125 5763 1349
rect 5877 1125 5923 1349
rect 6037 1125 6083 1349
rect 6197 1125 6243 1349
rect 6357 1125 6403 1349
rect 6517 1125 6563 1349
rect 6677 1125 6723 1349
rect 6837 1125 6883 1349
rect 6965 1125 7011 1349
rect 7125 1125 7171 1349
rect 7369 1125 7415 1349
rect 7529 1125 7575 1349
rect 7689 1125 7735 1349
rect 7849 1125 7895 1349
rect 8009 1125 8055 1349
rect 8169 1125 8215 1349
rect 8329 1125 8375 1349
rect 8489 1125 8535 1349
rect 8649 1125 8695 1349
rect 8777 1125 8823 1349
rect 8937 1125 8983 1349
rect -4799 932 -4753 1006
rect -4639 932 -4593 1006
rect -4233 944 -4187 1018
rect -4073 944 -4027 1018
rect -3913 944 -3867 1018
rect -3528 984 -3482 1030
rect -2968 984 -2922 1030
rect -2742 984 -2696 1030
rect -2182 984 -2136 1030
rect -1956 984 -1910 1030
rect -1396 984 -1350 1030
rect -1150 932 -1104 1006
rect -990 932 -944 1006
rect 121 739 167 963
rect 281 739 327 963
rect 409 739 455 963
rect 569 739 615 963
rect 729 739 775 963
rect 889 739 935 963
rect 1049 739 1095 963
rect 1209 739 1255 963
rect 1369 739 1415 963
rect 1529 739 1575 963
rect 1689 739 1735 963
rect 1933 739 1979 963
rect 2093 739 2139 963
rect 2253 739 2299 963
rect 2413 739 2459 963
rect 2573 739 2619 963
rect 2733 739 2779 963
rect 2893 739 2939 963
rect 3053 739 3099 963
rect 3213 739 3259 963
rect 3341 739 3387 963
rect 3501 739 3547 963
rect 3745 739 3791 963
rect 3905 739 3951 963
rect 4033 739 4079 963
rect 4193 739 4239 963
rect 4353 739 4399 963
rect 4513 739 4559 963
rect 4673 739 4719 963
rect 4833 739 4879 963
rect 4993 739 5039 963
rect 5153 739 5199 963
rect 5313 739 5359 963
rect 5557 739 5603 963
rect 5717 739 5763 963
rect 5877 739 5923 963
rect 6037 739 6083 963
rect 6197 739 6243 963
rect 6357 739 6403 963
rect 6517 739 6563 963
rect 6677 739 6723 963
rect 6837 739 6883 963
rect 6965 739 7011 963
rect 7125 739 7171 963
rect 7369 739 7415 963
rect 7529 739 7575 963
rect 7689 739 7735 963
rect 7849 739 7895 963
rect 8009 739 8055 963
rect 8169 739 8215 963
rect 8329 739 8375 963
rect 8489 739 8535 963
rect 8649 739 8695 963
rect 8777 739 8823 963
rect 8937 739 8983 963
rect 121 353 167 577
rect 281 353 327 577
rect 409 353 455 577
rect 569 353 615 577
rect 729 353 775 577
rect 889 353 935 577
rect 1049 353 1095 577
rect 1209 353 1255 577
rect 1369 353 1415 577
rect 1529 353 1575 577
rect 1689 353 1735 577
rect 1933 353 1979 577
rect 2093 353 2139 577
rect 2253 353 2299 577
rect 2413 353 2459 577
rect 2573 353 2619 577
rect 2733 353 2779 577
rect 2893 353 2939 577
rect 3053 353 3099 577
rect 3213 353 3259 577
rect 3341 353 3387 577
rect 3501 353 3547 577
rect 3745 353 3791 577
rect 3905 353 3951 577
rect 4033 353 4079 577
rect 4193 353 4239 577
rect 4353 353 4399 577
rect 4513 353 4559 577
rect 4673 353 4719 577
rect 4833 353 4879 577
rect 4993 353 5039 577
rect 5153 353 5199 577
rect 5313 353 5359 577
rect 5557 353 5603 577
rect 5717 353 5763 577
rect 5877 353 5923 577
rect 6037 353 6083 577
rect 6197 353 6243 577
rect 6357 353 6403 577
rect 6517 353 6563 577
rect 6677 353 6723 577
rect 6837 353 6883 577
rect 6965 353 7011 577
rect 7125 353 7171 577
rect 7369 353 7415 577
rect 7529 353 7575 577
rect 7689 353 7735 577
rect 7849 353 7895 577
rect 8009 353 8055 577
rect 8169 353 8215 577
rect 8329 353 8375 577
rect 8489 353 8535 577
rect 8649 353 8695 577
rect 8777 353 8823 577
rect 8937 353 8983 577
rect -4799 -406 -4753 -332
rect -4639 -406 -4593 -332
rect -4233 -418 -4187 -344
rect -4073 -418 -4027 -344
rect -3913 -418 -3867 -344
rect -3528 -430 -3482 -384
rect -2968 -430 -2922 -384
rect -2742 -430 -2696 -384
rect -2182 -430 -2136 -384
rect -1956 -430 -1910 -384
rect -1396 -430 -1350 -384
rect -1150 -406 -1104 -332
rect -990 -406 -944 -332
rect 121 -465 167 -241
rect 281 -465 327 -241
rect 409 -465 455 -241
rect 569 -465 615 -241
rect 729 -465 775 -241
rect 889 -465 935 -241
rect 1049 -465 1095 -241
rect 1209 -465 1255 -241
rect 1369 -465 1415 -241
rect 1529 -465 1575 -241
rect 1689 -465 1735 -241
rect 1933 -465 1979 -241
rect 2093 -465 2139 -241
rect 2253 -465 2299 -241
rect 2413 -465 2459 -241
rect 2573 -465 2619 -241
rect 2733 -465 2779 -241
rect 2893 -465 2939 -241
rect 3053 -465 3099 -241
rect 3213 -465 3259 -241
rect 3341 -465 3387 -241
rect 3501 -465 3547 -241
rect 3745 -465 3791 -241
rect 3905 -465 3951 -241
rect 4033 -465 4079 -241
rect 4193 -465 4239 -241
rect 4353 -465 4399 -241
rect 4513 -465 4559 -241
rect 4673 -465 4719 -241
rect 4833 -465 4879 -241
rect 4993 -465 5039 -241
rect 5153 -465 5199 -241
rect 5313 -465 5359 -241
rect 5557 -465 5603 -241
rect 5717 -465 5763 -241
rect 5877 -465 5923 -241
rect 6037 -465 6083 -241
rect 6197 -465 6243 -241
rect 6357 -465 6403 -241
rect 6517 -465 6563 -241
rect 6677 -465 6723 -241
rect 6837 -465 6883 -241
rect 6965 -465 7011 -241
rect 7125 -465 7171 -241
rect 7369 -465 7415 -241
rect 7529 -465 7575 -241
rect 7689 -465 7735 -241
rect 7849 -465 7895 -241
rect 8009 -465 8055 -241
rect 8169 -465 8215 -241
rect 8329 -465 8375 -241
rect 8489 -465 8535 -241
rect 8649 -465 8695 -241
rect 8777 -465 8823 -241
rect 8937 -465 8983 -241
rect -4233 -766 -4187 -692
rect -4073 -766 -4027 -692
rect -3913 -766 -3867 -692
rect -3528 -726 -3482 -680
rect -2968 -726 -2922 -680
rect -2742 -726 -2696 -680
rect -2182 -726 -2136 -680
rect -1956 -726 -1910 -680
rect -1396 -726 -1350 -680
rect -1150 -778 -1104 -704
rect -990 -778 -944 -704
rect 121 -851 167 -627
rect 281 -851 327 -627
rect 409 -851 455 -627
rect 569 -851 615 -627
rect 729 -851 775 -627
rect 889 -851 935 -627
rect 1049 -851 1095 -627
rect 1209 -851 1255 -627
rect 1369 -851 1415 -627
rect 1529 -851 1575 -627
rect 1689 -851 1735 -627
rect 1933 -851 1979 -627
rect 2093 -851 2139 -627
rect 2253 -851 2299 -627
rect 2413 -851 2459 -627
rect 2573 -851 2619 -627
rect 2733 -851 2779 -627
rect 2893 -851 2939 -627
rect 3053 -851 3099 -627
rect 3213 -851 3259 -627
rect 3341 -851 3387 -627
rect 3501 -851 3547 -627
rect 3745 -851 3791 -627
rect 3905 -851 3951 -627
rect 4033 -851 4079 -627
rect 4193 -851 4239 -627
rect 4353 -851 4399 -627
rect 4513 -851 4559 -627
rect 4673 -851 4719 -627
rect 4833 -851 4879 -627
rect 4993 -851 5039 -627
rect 5153 -851 5199 -627
rect 5313 -851 5359 -627
rect 5557 -851 5603 -627
rect 5717 -851 5763 -627
rect 5877 -851 5923 -627
rect 6037 -851 6083 -627
rect 6197 -851 6243 -627
rect 6357 -851 6403 -627
rect 6517 -851 6563 -627
rect 6677 -851 6723 -627
rect 6837 -851 6883 -627
rect 6965 -851 7011 -627
rect 7125 -851 7171 -627
rect 7369 -851 7415 -627
rect 7529 -851 7575 -627
rect 7689 -851 7735 -627
rect 7849 -851 7895 -627
rect 8009 -851 8055 -627
rect 8169 -851 8215 -627
rect 8329 -851 8375 -627
rect 8489 -851 8535 -627
rect 8649 -851 8695 -627
rect 8777 -851 8823 -627
rect 8937 -851 8983 -627
rect 121 -1237 167 -1013
rect 281 -1237 327 -1013
rect 409 -1237 455 -1013
rect 569 -1237 615 -1013
rect 729 -1237 775 -1013
rect 889 -1237 935 -1013
rect 1049 -1237 1095 -1013
rect 1209 -1237 1255 -1013
rect 1369 -1237 1415 -1013
rect 1529 -1237 1575 -1013
rect 1689 -1237 1735 -1013
rect 1933 -1237 1979 -1013
rect 2093 -1237 2139 -1013
rect 2253 -1237 2299 -1013
rect 2413 -1237 2459 -1013
rect 2573 -1237 2619 -1013
rect 2733 -1237 2779 -1013
rect 2893 -1237 2939 -1013
rect 3053 -1237 3099 -1013
rect 3213 -1237 3259 -1013
rect 3341 -1237 3387 -1013
rect 3501 -1237 3547 -1013
rect 3745 -1237 3791 -1013
rect 3905 -1237 3951 -1013
rect 4033 -1237 4079 -1013
rect 4193 -1237 4239 -1013
rect 4353 -1237 4399 -1013
rect 4513 -1237 4559 -1013
rect 4673 -1237 4719 -1013
rect 4833 -1237 4879 -1013
rect 4993 -1237 5039 -1013
rect 5153 -1237 5199 -1013
rect 5313 -1237 5359 -1013
rect 5557 -1237 5603 -1013
rect 5717 -1237 5763 -1013
rect 5877 -1237 5923 -1013
rect 6037 -1237 6083 -1013
rect 6197 -1237 6243 -1013
rect 6357 -1237 6403 -1013
rect 6517 -1237 6563 -1013
rect 6677 -1237 6723 -1013
rect 6837 -1237 6883 -1013
rect 6965 -1237 7011 -1013
rect 7125 -1237 7171 -1013
rect 7369 -1237 7415 -1013
rect 7529 -1237 7575 -1013
rect 7689 -1237 7735 -1013
rect 7849 -1237 7895 -1013
rect 8009 -1237 8055 -1013
rect 8169 -1237 8215 -1013
rect 8329 -1237 8375 -1013
rect 8489 -1237 8535 -1013
rect 8649 -1237 8695 -1013
rect 8777 -1237 8823 -1013
rect 8937 -1237 8983 -1013
rect -4076 -6203 -4030 -5979
rect -3916 -6203 -3870 -5979
rect -3788 -6203 -3742 -5979
rect -3628 -6203 -3582 -5979
rect -3468 -6203 -3422 -5979
rect -3308 -6203 -3262 -5979
rect -3148 -6203 -3102 -5979
rect -2988 -6203 -2942 -5979
rect -2828 -6203 -2782 -5979
rect -2668 -6203 -2622 -5979
rect -2508 -6203 -2462 -5979
rect -2264 -6203 -2218 -5979
rect -2104 -6203 -2058 -5979
rect -1944 -6203 -1898 -5979
rect -1784 -6203 -1738 -5979
rect -1624 -6203 -1578 -5979
rect -1464 -6203 -1418 -5979
rect -1304 -6203 -1258 -5979
rect -1144 -6203 -1098 -5979
rect -984 -6203 -938 -5979
rect -856 -6203 -810 -5979
rect -696 -6203 -650 -5979
rect 121 -6203 167 -5979
rect 281 -6203 327 -5979
rect 409 -6203 455 -5979
rect 569 -6203 615 -5979
rect 729 -6203 775 -5979
rect 889 -6203 935 -5979
rect 1049 -6203 1095 -5979
rect 1209 -6203 1255 -5979
rect 1369 -6203 1415 -5979
rect 1529 -6203 1575 -5979
rect 1689 -6203 1735 -5979
rect 1933 -6203 1979 -5979
rect 2093 -6203 2139 -5979
rect 2253 -6203 2299 -5979
rect 2413 -6203 2459 -5979
rect 2573 -6203 2619 -5979
rect 2733 -6203 2779 -5979
rect 2893 -6203 2939 -5979
rect 3053 -6203 3099 -5979
rect 3213 -6203 3259 -5979
rect 3341 -6203 3387 -5979
rect 3501 -6203 3547 -5979
rect 3745 -6203 3791 -5979
rect 3905 -6203 3951 -5979
rect 4033 -6203 4079 -5979
rect 4193 -6203 4239 -5979
rect 4353 -6203 4399 -5979
rect 4513 -6203 4559 -5979
rect 4673 -6203 4719 -5979
rect 4833 -6203 4879 -5979
rect 4993 -6203 5039 -5979
rect 5153 -6203 5199 -5979
rect 5313 -6203 5359 -5979
rect 5557 -6203 5603 -5979
rect 5717 -6203 5763 -5979
rect 5877 -6203 5923 -5979
rect 6037 -6203 6083 -5979
rect 6197 -6203 6243 -5979
rect 6357 -6203 6403 -5979
rect 6517 -6203 6563 -5979
rect 6677 -6203 6723 -5979
rect 6837 -6203 6883 -5979
rect 6965 -6203 7011 -5979
rect 7125 -6203 7171 -5979
rect 7369 -6203 7415 -5979
rect 7529 -6203 7575 -5979
rect 7689 -6203 7735 -5979
rect 7849 -6203 7895 -5979
rect 8009 -6203 8055 -5979
rect 8169 -6203 8215 -5979
rect 8329 -6203 8375 -5979
rect 8489 -6203 8535 -5979
rect 8649 -6203 8695 -5979
rect 8777 -6203 8823 -5979
rect 8937 -6203 8983 -5979
rect -4076 -6589 -4030 -6365
rect -3916 -6589 -3870 -6365
rect -3788 -6589 -3742 -6365
rect -3628 -6589 -3582 -6365
rect -3468 -6589 -3422 -6365
rect -3308 -6589 -3262 -6365
rect -3148 -6589 -3102 -6365
rect -2988 -6589 -2942 -6365
rect -2828 -6589 -2782 -6365
rect -2668 -6589 -2622 -6365
rect -2508 -6589 -2462 -6365
rect -2264 -6589 -2218 -6365
rect -2104 -6589 -2058 -6365
rect -1944 -6589 -1898 -6365
rect -1784 -6589 -1738 -6365
rect -1624 -6589 -1578 -6365
rect -1464 -6589 -1418 -6365
rect -1304 -6589 -1258 -6365
rect -1144 -6589 -1098 -6365
rect -984 -6589 -938 -6365
rect -856 -6589 -810 -6365
rect -696 -6589 -650 -6365
rect 121 -6589 167 -6365
rect 281 -6589 327 -6365
rect 409 -6589 455 -6365
rect 569 -6589 615 -6365
rect 729 -6589 775 -6365
rect 889 -6589 935 -6365
rect 1049 -6589 1095 -6365
rect 1209 -6589 1255 -6365
rect 1369 -6589 1415 -6365
rect 1529 -6589 1575 -6365
rect 1689 -6589 1735 -6365
rect 1933 -6589 1979 -6365
rect 2093 -6589 2139 -6365
rect 2253 -6589 2299 -6365
rect 2413 -6589 2459 -6365
rect 2573 -6589 2619 -6365
rect 2733 -6589 2779 -6365
rect 2893 -6589 2939 -6365
rect 3053 -6589 3099 -6365
rect 3213 -6589 3259 -6365
rect 3341 -6589 3387 -6365
rect 3501 -6589 3547 -6365
rect 3745 -6589 3791 -6365
rect 3905 -6589 3951 -6365
rect 4033 -6589 4079 -6365
rect 4193 -6589 4239 -6365
rect 4353 -6589 4399 -6365
rect 4513 -6589 4559 -6365
rect 4673 -6589 4719 -6365
rect 4833 -6589 4879 -6365
rect 4993 -6589 5039 -6365
rect 5153 -6589 5199 -6365
rect 5313 -6589 5359 -6365
rect 5557 -6589 5603 -6365
rect 5717 -6589 5763 -6365
rect 5877 -6589 5923 -6365
rect 6037 -6589 6083 -6365
rect 6197 -6589 6243 -6365
rect 6357 -6589 6403 -6365
rect 6517 -6589 6563 -6365
rect 6677 -6589 6723 -6365
rect 6837 -6589 6883 -6365
rect 6965 -6589 7011 -6365
rect 7125 -6589 7171 -6365
rect 7369 -6589 7415 -6365
rect 7529 -6589 7575 -6365
rect 7689 -6589 7735 -6365
rect 7849 -6589 7895 -6365
rect 8009 -6589 8055 -6365
rect 8169 -6589 8215 -6365
rect 8329 -6589 8375 -6365
rect 8489 -6589 8535 -6365
rect 8649 -6589 8695 -6365
rect 8777 -6589 8823 -6365
rect 8937 -6589 8983 -6365
rect -4076 -6975 -4030 -6751
rect -3916 -6975 -3870 -6751
rect -3788 -6975 -3742 -6751
rect -3628 -6975 -3582 -6751
rect -3468 -6975 -3422 -6751
rect -3308 -6975 -3262 -6751
rect -3148 -6975 -3102 -6751
rect -2988 -6975 -2942 -6751
rect -2828 -6975 -2782 -6751
rect -2668 -6975 -2622 -6751
rect -2508 -6975 -2462 -6751
rect -2264 -6975 -2218 -6751
rect -2104 -6975 -2058 -6751
rect -1944 -6975 -1898 -6751
rect -1784 -6975 -1738 -6751
rect -1624 -6975 -1578 -6751
rect -1464 -6975 -1418 -6751
rect -1304 -6975 -1258 -6751
rect -1144 -6975 -1098 -6751
rect -984 -6975 -938 -6751
rect -856 -6975 -810 -6751
rect -696 -6975 -650 -6751
rect 121 -6975 167 -6751
rect 281 -6975 327 -6751
rect 409 -6975 455 -6751
rect 569 -6975 615 -6751
rect 729 -6975 775 -6751
rect 889 -6975 935 -6751
rect 1049 -6975 1095 -6751
rect 1209 -6975 1255 -6751
rect 1369 -6975 1415 -6751
rect 1529 -6975 1575 -6751
rect 1689 -6975 1735 -6751
rect 1933 -6975 1979 -6751
rect 2093 -6975 2139 -6751
rect 2253 -6975 2299 -6751
rect 2413 -6975 2459 -6751
rect 2573 -6975 2619 -6751
rect 2733 -6975 2779 -6751
rect 2893 -6975 2939 -6751
rect 3053 -6975 3099 -6751
rect 3213 -6975 3259 -6751
rect 3341 -6975 3387 -6751
rect 3501 -6975 3547 -6751
rect 3745 -6975 3791 -6751
rect 3905 -6975 3951 -6751
rect 4033 -6975 4079 -6751
rect 4193 -6975 4239 -6751
rect 4353 -6975 4399 -6751
rect 4513 -6975 4559 -6751
rect 4673 -6975 4719 -6751
rect 4833 -6975 4879 -6751
rect 4993 -6975 5039 -6751
rect 5153 -6975 5199 -6751
rect 5313 -6975 5359 -6751
rect 5557 -6975 5603 -6751
rect 5717 -6975 5763 -6751
rect 5877 -6975 5923 -6751
rect 6037 -6975 6083 -6751
rect 6197 -6975 6243 -6751
rect 6357 -6975 6403 -6751
rect 6517 -6975 6563 -6751
rect 6677 -6975 6723 -6751
rect 6837 -6975 6883 -6751
rect 6965 -6975 7011 -6751
rect 7125 -6975 7171 -6751
rect 7369 -6975 7415 -6751
rect 7529 -6975 7575 -6751
rect 7689 -6975 7735 -6751
rect 7849 -6975 7895 -6751
rect 8009 -6975 8055 -6751
rect 8169 -6975 8215 -6751
rect 8329 -6975 8375 -6751
rect 8489 -6975 8535 -6751
rect 8649 -6975 8695 -6751
rect 8777 -6975 8823 -6751
rect 8937 -6975 8983 -6751
<< pdiffc >>
rect 121 5289 167 5763
rect 281 5289 327 5763
rect 441 5289 487 5763
rect 601 5289 647 5763
rect 761 5289 807 5763
rect 921 5289 967 5763
rect 1081 5289 1127 5763
rect 1241 5289 1287 5763
rect 1401 5289 1447 5763
rect 1529 5289 1575 5763
rect 1689 5289 1735 5763
rect 1933 5289 1979 5763
rect 2093 5289 2139 5763
rect 2221 5289 2267 5763
rect 2381 5289 2427 5763
rect 2541 5289 2587 5763
rect 2701 5289 2747 5763
rect 2861 5289 2907 5763
rect 3021 5289 3067 5763
rect 3181 5289 3227 5763
rect 3341 5289 3387 5763
rect 3501 5289 3547 5763
rect 3745 5289 3791 5763
rect 3905 5289 3951 5763
rect 4033 5289 4079 5763
rect 4193 5289 4239 5763
rect 4353 5289 4399 5763
rect 4513 5289 4559 5763
rect 4673 5289 4719 5763
rect 4833 5289 4879 5763
rect 4993 5289 5039 5763
rect 5153 5289 5199 5763
rect 5313 5289 5359 5763
rect 5557 5289 5603 5763
rect 5717 5289 5763 5763
rect 5845 5289 5891 5763
rect 6005 5289 6051 5763
rect 6165 5289 6211 5763
rect 6325 5289 6371 5763
rect 6485 5289 6531 5763
rect 6645 5289 6691 5763
rect 6805 5289 6851 5763
rect 6965 5289 7011 5763
rect 7125 5289 7171 5763
rect 7369 5289 7415 5763
rect 7529 5289 7575 5763
rect 7657 5289 7703 5763
rect 7817 5289 7863 5763
rect 7977 5289 8023 5763
rect 8137 5289 8183 5763
rect 8297 5289 8343 5763
rect 8457 5289 8503 5763
rect 8617 5289 8663 5763
rect 8777 5289 8823 5763
rect 8937 5289 8983 5763
rect 121 4653 167 5127
rect 281 4653 327 5127
rect 441 4653 487 5127
rect 601 4653 647 5127
rect 761 4653 807 5127
rect 921 4653 967 5127
rect 1081 4653 1127 5127
rect 1241 4653 1287 5127
rect 1401 4653 1447 5127
rect 1529 4653 1575 5127
rect 1689 4653 1735 5127
rect 1933 4653 1979 5127
rect 2093 4653 2139 5127
rect 2221 4653 2267 5127
rect 2381 4653 2427 5127
rect 2541 4653 2587 5127
rect 2701 4653 2747 5127
rect 2861 4653 2907 5127
rect 3021 4653 3067 5127
rect 3181 4653 3227 5127
rect 3341 4653 3387 5127
rect 3501 4653 3547 5127
rect 3745 4653 3791 5127
rect 3905 4653 3951 5127
rect 4033 4653 4079 5127
rect 4193 4653 4239 5127
rect 4353 4653 4399 5127
rect 4513 4653 4559 5127
rect 4673 4653 4719 5127
rect 4833 4653 4879 5127
rect 4993 4653 5039 5127
rect 5153 4653 5199 5127
rect 5313 4653 5359 5127
rect 5557 4653 5603 5127
rect 5717 4653 5763 5127
rect 5845 4653 5891 5127
rect 6005 4653 6051 5127
rect 6165 4653 6211 5127
rect 6325 4653 6371 5127
rect 6485 4653 6531 5127
rect 6645 4653 6691 5127
rect 6805 4653 6851 5127
rect 6965 4653 7011 5127
rect 7125 4653 7171 5127
rect 7369 4653 7415 5127
rect 7529 4653 7575 5127
rect 7657 4653 7703 5127
rect 7817 4653 7863 5127
rect 7977 4653 8023 5127
rect 8137 4653 8183 5127
rect 8297 4653 8343 5127
rect 8457 4653 8503 5127
rect 8617 4653 8663 5127
rect 8777 4653 8823 5127
rect 8937 4653 8983 5127
rect 121 4017 167 4491
rect 281 4017 327 4491
rect 441 4017 487 4491
rect 601 4017 647 4491
rect 761 4017 807 4491
rect 921 4017 967 4491
rect 1081 4017 1127 4491
rect 1241 4017 1287 4491
rect 1401 4017 1447 4491
rect 1529 4017 1575 4491
rect 1689 4017 1735 4491
rect 1933 4017 1979 4491
rect 2093 4017 2139 4491
rect 2221 4017 2267 4491
rect 2381 4017 2427 4491
rect 2541 4017 2587 4491
rect 2701 4017 2747 4491
rect 2861 4017 2907 4491
rect 3021 4017 3067 4491
rect 3181 4017 3227 4491
rect 3341 4017 3387 4491
rect 3501 4017 3547 4491
rect 3745 4017 3791 4491
rect 3905 4017 3951 4491
rect 4033 4017 4079 4491
rect 4193 4017 4239 4491
rect 4353 4017 4399 4491
rect 4513 4017 4559 4491
rect 4673 4017 4719 4491
rect 4833 4017 4879 4491
rect 4993 4017 5039 4491
rect 5153 4017 5199 4491
rect 5313 4017 5359 4491
rect 5557 4017 5603 4491
rect 5717 4017 5763 4491
rect 5845 4017 5891 4491
rect 6005 4017 6051 4491
rect 6165 4017 6211 4491
rect 6325 4017 6371 4491
rect 6485 4017 6531 4491
rect 6645 4017 6691 4491
rect 6805 4017 6851 4491
rect 6965 4017 7011 4491
rect 7125 4017 7171 4491
rect 7369 4017 7415 4491
rect 7529 4017 7575 4491
rect 7657 4017 7703 4491
rect 7817 4017 7863 4491
rect 7977 4017 8023 4491
rect 8137 4017 8183 4491
rect 8297 4017 8343 4491
rect 8457 4017 8503 4491
rect 8617 4017 8663 4491
rect 8777 4017 8823 4491
rect 8937 4017 8983 4491
rect -4799 3386 -4753 3560
rect -4639 3386 -4593 3560
rect -4393 3341 -4347 3515
rect -4233 3341 -4187 3515
rect -4073 3341 -4027 3515
rect -3913 3341 -3867 3515
rect -3753 3341 -3707 3515
rect -3520 3464 -3474 3526
rect -2968 3464 -2922 3526
rect -2734 3464 -2688 3526
rect -2182 3464 -2136 3526
rect -1948 3464 -1902 3526
rect -1396 3464 -1350 3526
rect -1150 3386 -1104 3560
rect -990 3386 -944 3560
rect 121 2949 167 3423
rect 281 2949 327 3423
rect 409 2949 455 3423
rect 569 2949 615 3423
rect 729 2949 775 3423
rect 889 2949 935 3423
rect 1049 2949 1095 3423
rect 1209 2949 1255 3423
rect 1369 2949 1415 3423
rect 1529 2949 1575 3423
rect 1689 2949 1735 3423
rect 1933 2949 1979 3423
rect 2093 2949 2139 3423
rect 2253 2949 2299 3423
rect 2413 2949 2459 3423
rect 2573 2949 2619 3423
rect 2733 2949 2779 3423
rect 2893 2949 2939 3423
rect 3053 2949 3099 3423
rect 3213 2949 3259 3423
rect 3341 2949 3387 3423
rect 3501 2949 3547 3423
rect 3745 2949 3791 3423
rect 3905 2949 3951 3423
rect 4033 2949 4079 3423
rect 4193 2949 4239 3423
rect 4353 2949 4399 3423
rect 4513 2949 4559 3423
rect 4673 2949 4719 3423
rect 4833 2949 4879 3423
rect 4993 2949 5039 3423
rect 5153 2949 5199 3423
rect 5313 2949 5359 3423
rect 5557 2949 5603 3423
rect 5717 2949 5763 3423
rect 5877 2949 5923 3423
rect 6037 2949 6083 3423
rect 6197 2949 6243 3423
rect 6357 2949 6403 3423
rect 6517 2949 6563 3423
rect 6677 2949 6723 3423
rect 6837 2949 6883 3423
rect 6965 2949 7011 3423
rect 7125 2949 7171 3423
rect 7369 2949 7415 3423
rect 7529 2949 7575 3423
rect 7689 2949 7735 3423
rect 7849 2949 7895 3423
rect 8009 2949 8055 3423
rect 8169 2949 8215 3423
rect 8329 2949 8375 3423
rect 8489 2949 8535 3423
rect 8649 2949 8695 3423
rect 8777 2949 8823 3423
rect 8937 2949 8983 3423
rect -4393 2215 -4347 2389
rect -4233 2215 -4187 2389
rect -4073 2215 -4027 2389
rect -3913 2215 -3867 2389
rect -3753 2215 -3707 2389
rect -3520 2204 -3474 2266
rect -2968 2204 -2922 2266
rect -2734 2204 -2688 2266
rect -2182 2204 -2136 2266
rect -1948 2204 -1902 2266
rect -1396 2204 -1350 2266
rect -1150 2170 -1104 2344
rect -990 2170 -944 2344
rect 121 2313 167 2787
rect 281 2313 327 2787
rect 409 2313 455 2787
rect 569 2313 615 2787
rect 729 2313 775 2787
rect 889 2313 935 2787
rect 1049 2313 1095 2787
rect 1209 2313 1255 2787
rect 1369 2313 1415 2787
rect 1529 2313 1575 2787
rect 1689 2313 1735 2787
rect 1933 2313 1979 2787
rect 2093 2313 2139 2787
rect 2253 2313 2299 2787
rect 2413 2313 2459 2787
rect 2573 2313 2619 2787
rect 2733 2313 2779 2787
rect 2893 2313 2939 2787
rect 3053 2313 3099 2787
rect 3213 2313 3259 2787
rect 3341 2313 3387 2787
rect 3501 2313 3547 2787
rect 3745 2313 3791 2787
rect 3905 2313 3951 2787
rect 4033 2313 4079 2787
rect 4193 2313 4239 2787
rect 4353 2313 4399 2787
rect 4513 2313 4559 2787
rect 4673 2313 4719 2787
rect 4833 2313 4879 2787
rect 4993 2313 5039 2787
rect 5153 2313 5199 2787
rect 5313 2313 5359 2787
rect 5557 2313 5603 2787
rect 5717 2313 5763 2787
rect 5877 2313 5923 2787
rect 6037 2313 6083 2787
rect 6197 2313 6243 2787
rect 6357 2313 6403 2787
rect 6517 2313 6563 2787
rect 6677 2313 6723 2787
rect 6837 2313 6883 2787
rect 6965 2313 7011 2787
rect 7125 2313 7171 2787
rect 7369 2313 7415 2787
rect 7529 2313 7575 2787
rect 7689 2313 7735 2787
rect 7849 2313 7895 2787
rect 8009 2313 8055 2787
rect 8169 2313 8215 2787
rect 8329 2313 8375 2787
rect 8489 2313 8535 2787
rect 8649 2313 8695 2787
rect 8777 2313 8823 2787
rect 8937 2313 8983 2787
rect -4393 1631 -4347 1805
rect -4233 1631 -4187 1805
rect -4073 1631 -4027 1805
rect -3913 1631 -3867 1805
rect -3753 1631 -3707 1805
rect -3520 1754 -3474 1816
rect -2968 1754 -2922 1816
rect -2734 1754 -2688 1816
rect -2182 1754 -2136 1816
rect -1948 1754 -1902 1816
rect -1396 1754 -1350 1816
rect -1150 1676 -1104 1850
rect -990 1676 -944 1850
rect 121 1677 167 2151
rect 281 1677 327 2151
rect 409 1677 455 2151
rect 569 1677 615 2151
rect 729 1677 775 2151
rect 889 1677 935 2151
rect 1049 1677 1095 2151
rect 1209 1677 1255 2151
rect 1369 1677 1415 2151
rect 1529 1677 1575 2151
rect 1689 1677 1735 2151
rect 1933 1677 1979 2151
rect 2093 1677 2139 2151
rect 2253 1677 2299 2151
rect 2413 1677 2459 2151
rect 2573 1677 2619 2151
rect 2733 1677 2779 2151
rect 2893 1677 2939 2151
rect 3053 1677 3099 2151
rect 3213 1677 3259 2151
rect 3341 1677 3387 2151
rect 3501 1677 3547 2151
rect 3745 1677 3791 2151
rect 3905 1677 3951 2151
rect 4033 1677 4079 2151
rect 4193 1677 4239 2151
rect 4353 1677 4399 2151
rect 4513 1677 4559 2151
rect 4673 1677 4719 2151
rect 4833 1677 4879 2151
rect 4993 1677 5039 2151
rect 5153 1677 5199 2151
rect 5313 1677 5359 2151
rect 5557 1677 5603 2151
rect 5717 1677 5763 2151
rect 5877 1677 5923 2151
rect 6037 1677 6083 2151
rect 6197 1677 6243 2151
rect 6357 1677 6403 2151
rect 6517 1677 6563 2151
rect 6677 1677 6723 2151
rect 6837 1677 6883 2151
rect 6965 1677 7011 2151
rect 7125 1677 7171 2151
rect 7369 1677 7415 2151
rect 7529 1677 7575 2151
rect 7689 1677 7735 2151
rect 7849 1677 7895 2151
rect 8009 1677 8055 2151
rect 8169 1677 8215 2151
rect 8329 1677 8375 2151
rect 8489 1677 8535 2151
rect 8649 1677 8695 2151
rect 8777 1677 8823 2151
rect 8937 1677 8983 2151
rect -4799 460 -4753 634
rect -4639 460 -4593 634
rect -4393 505 -4347 679
rect -4233 505 -4187 679
rect -4073 505 -4027 679
rect -3913 505 -3867 679
rect -3753 505 -3707 679
rect -3520 494 -3474 556
rect -2968 494 -2922 556
rect -2734 494 -2688 556
rect -2182 494 -2136 556
rect -1948 494 -1902 556
rect -1396 494 -1350 556
rect -1150 460 -1104 634
rect -990 460 -944 634
rect -4799 -34 -4753 140
rect -4639 -34 -4593 140
rect -4393 -79 -4347 95
rect -4233 -79 -4187 95
rect -4073 -79 -4027 95
rect -3913 -79 -3867 95
rect -3753 -79 -3707 95
rect -3520 44 -3474 106
rect -2968 44 -2922 106
rect -2734 44 -2688 106
rect -2182 44 -2136 106
rect -1948 44 -1902 106
rect -1396 44 -1350 106
rect -1150 -34 -1104 140
rect -990 -34 -944 140
rect -4393 -1205 -4347 -1031
rect -4233 -1205 -4187 -1031
rect -4073 -1205 -4027 -1031
rect -3913 -1205 -3867 -1031
rect -3753 -1205 -3707 -1031
rect -3520 -1216 -3474 -1154
rect -2968 -1216 -2922 -1154
rect -2734 -1216 -2688 -1154
rect -2182 -1216 -2136 -1154
rect -1948 -1216 -1902 -1154
rect -1396 -1216 -1350 -1154
rect -1150 -1250 -1104 -1076
rect -990 -1250 -944 -1076
rect 121 -2039 167 -1565
rect 281 -2039 327 -1565
rect 409 -2039 455 -1565
rect 569 -2039 615 -1565
rect 729 -2039 775 -1565
rect 889 -2039 935 -1565
rect 1049 -2039 1095 -1565
rect 1209 -2039 1255 -1565
rect 1369 -2039 1415 -1565
rect 1529 -2039 1575 -1565
rect 1689 -2039 1735 -1565
rect 1933 -2039 1979 -1565
rect 2093 -2039 2139 -1565
rect 2253 -2039 2299 -1565
rect 2413 -2039 2459 -1565
rect 2573 -2039 2619 -1565
rect 2733 -2039 2779 -1565
rect 2893 -2039 2939 -1565
rect 3053 -2039 3099 -1565
rect 3213 -2039 3259 -1565
rect 3341 -2039 3387 -1565
rect 3501 -2039 3547 -1565
rect 3745 -2039 3791 -1565
rect 3905 -2039 3951 -1565
rect 4033 -2039 4079 -1565
rect 4193 -2039 4239 -1565
rect 4353 -2039 4399 -1565
rect 4513 -2039 4559 -1565
rect 4673 -2039 4719 -1565
rect 4833 -2039 4879 -1565
rect 4993 -2039 5039 -1565
rect 5153 -2039 5199 -1565
rect 5313 -2039 5359 -1565
rect 5557 -2039 5603 -1565
rect 5717 -2039 5763 -1565
rect 5877 -2039 5923 -1565
rect 6037 -2039 6083 -1565
rect 6197 -2039 6243 -1565
rect 6357 -2039 6403 -1565
rect 6517 -2039 6563 -1565
rect 6677 -2039 6723 -1565
rect 6837 -2039 6883 -1565
rect 6965 -2039 7011 -1565
rect 7125 -2039 7171 -1565
rect 7369 -2039 7415 -1565
rect 7529 -2039 7575 -1565
rect 7689 -2039 7735 -1565
rect 7849 -2039 7895 -1565
rect 8009 -2039 8055 -1565
rect 8169 -2039 8215 -1565
rect 8329 -2039 8375 -1565
rect 8489 -2039 8535 -1565
rect 8649 -2039 8695 -1565
rect 8777 -2039 8823 -1565
rect 8937 -2039 8983 -1565
rect 121 -2675 167 -2201
rect 281 -2675 327 -2201
rect 409 -2675 455 -2201
rect 569 -2675 615 -2201
rect 729 -2675 775 -2201
rect 889 -2675 935 -2201
rect 1049 -2675 1095 -2201
rect 1209 -2675 1255 -2201
rect 1369 -2675 1415 -2201
rect 1529 -2675 1575 -2201
rect 1689 -2675 1735 -2201
rect 1933 -2675 1979 -2201
rect 2093 -2675 2139 -2201
rect 2253 -2675 2299 -2201
rect 2413 -2675 2459 -2201
rect 2573 -2675 2619 -2201
rect 2733 -2675 2779 -2201
rect 2893 -2675 2939 -2201
rect 3053 -2675 3099 -2201
rect 3213 -2675 3259 -2201
rect 3341 -2675 3387 -2201
rect 3501 -2675 3547 -2201
rect 3745 -2675 3791 -2201
rect 3905 -2675 3951 -2201
rect 4033 -2675 4079 -2201
rect 4193 -2675 4239 -2201
rect 4353 -2675 4399 -2201
rect 4513 -2675 4559 -2201
rect 4673 -2675 4719 -2201
rect 4833 -2675 4879 -2201
rect 4993 -2675 5039 -2201
rect 5153 -2675 5199 -2201
rect 5313 -2675 5359 -2201
rect 5557 -2675 5603 -2201
rect 5717 -2675 5763 -2201
rect 5877 -2675 5923 -2201
rect 6037 -2675 6083 -2201
rect 6197 -2675 6243 -2201
rect 6357 -2675 6403 -2201
rect 6517 -2675 6563 -2201
rect 6677 -2675 6723 -2201
rect 6837 -2675 6883 -2201
rect 6965 -2675 7011 -2201
rect 7125 -2675 7171 -2201
rect 7369 -2675 7415 -2201
rect 7529 -2675 7575 -2201
rect 7689 -2675 7735 -2201
rect 7849 -2675 7895 -2201
rect 8009 -2675 8055 -2201
rect 8169 -2675 8215 -2201
rect 8329 -2675 8375 -2201
rect 8489 -2675 8535 -2201
rect 8649 -2675 8695 -2201
rect 8777 -2675 8823 -2201
rect 8937 -2675 8983 -2201
rect 121 -3311 167 -2837
rect 281 -3311 327 -2837
rect 409 -3311 455 -2837
rect 569 -3311 615 -2837
rect 729 -3311 775 -2837
rect 889 -3311 935 -2837
rect 1049 -3311 1095 -2837
rect 1209 -3311 1255 -2837
rect 1369 -3311 1415 -2837
rect 1529 -3311 1575 -2837
rect 1689 -3311 1735 -2837
rect 1933 -3311 1979 -2837
rect 2093 -3311 2139 -2837
rect 2253 -3311 2299 -2837
rect 2413 -3311 2459 -2837
rect 2573 -3311 2619 -2837
rect 2733 -3311 2779 -2837
rect 2893 -3311 2939 -2837
rect 3053 -3311 3099 -2837
rect 3213 -3311 3259 -2837
rect 3341 -3311 3387 -2837
rect 3501 -3311 3547 -2837
rect 3745 -3311 3791 -2837
rect 3905 -3311 3951 -2837
rect 4033 -3311 4079 -2837
rect 4193 -3311 4239 -2837
rect 4353 -3311 4399 -2837
rect 4513 -3311 4559 -2837
rect 4673 -3311 4719 -2837
rect 4833 -3311 4879 -2837
rect 4993 -3311 5039 -2837
rect 5153 -3311 5199 -2837
rect 5313 -3311 5359 -2837
rect 5557 -3311 5603 -2837
rect 5717 -3311 5763 -2837
rect 5877 -3311 5923 -2837
rect 6037 -3311 6083 -2837
rect 6197 -3311 6243 -2837
rect 6357 -3311 6403 -2837
rect 6517 -3311 6563 -2837
rect 6677 -3311 6723 -2837
rect 6837 -3311 6883 -2837
rect 6965 -3311 7011 -2837
rect 7125 -3311 7171 -2837
rect 7369 -3311 7415 -2837
rect 7529 -3311 7575 -2837
rect 7689 -3311 7735 -2837
rect 7849 -3311 7895 -2837
rect 8009 -3311 8055 -2837
rect 8169 -3311 8215 -2837
rect 8329 -3311 8375 -2837
rect 8489 -3311 8535 -2837
rect 8649 -3311 8695 -2837
rect 8777 -3311 8823 -2837
rect 8937 -3311 8983 -2837
rect -4076 -4379 -4030 -3905
rect -3916 -4379 -3870 -3905
rect -3788 -4379 -3742 -3905
rect -3628 -4379 -3582 -3905
rect -3468 -4379 -3422 -3905
rect -3308 -4379 -3262 -3905
rect -3148 -4379 -3102 -3905
rect -2988 -4379 -2942 -3905
rect -2828 -4379 -2782 -3905
rect -2668 -4379 -2622 -3905
rect -2508 -4379 -2462 -3905
rect -2264 -4379 -2218 -3905
rect -2104 -4379 -2058 -3905
rect -1944 -4379 -1898 -3905
rect -1784 -4379 -1738 -3905
rect -1624 -4379 -1578 -3905
rect -1464 -4379 -1418 -3905
rect -1304 -4379 -1258 -3905
rect -1144 -4379 -1098 -3905
rect -984 -4379 -938 -3905
rect -856 -4379 -810 -3905
rect -696 -4379 -650 -3905
rect 121 -4379 167 -3905
rect 281 -4379 327 -3905
rect 409 -4379 455 -3905
rect 569 -4379 615 -3905
rect 729 -4379 775 -3905
rect 889 -4379 935 -3905
rect 1049 -4379 1095 -3905
rect 1209 -4379 1255 -3905
rect 1369 -4379 1415 -3905
rect 1529 -4379 1575 -3905
rect 1689 -4379 1735 -3905
rect 1933 -4379 1979 -3905
rect 2093 -4379 2139 -3905
rect 2253 -4379 2299 -3905
rect 2413 -4379 2459 -3905
rect 2573 -4379 2619 -3905
rect 2733 -4379 2779 -3905
rect 2893 -4379 2939 -3905
rect 3053 -4379 3099 -3905
rect 3213 -4379 3259 -3905
rect 3341 -4379 3387 -3905
rect 3501 -4379 3547 -3905
rect 3745 -4379 3791 -3905
rect 3905 -4379 3951 -3905
rect 4033 -4379 4079 -3905
rect 4193 -4379 4239 -3905
rect 4353 -4379 4399 -3905
rect 4513 -4379 4559 -3905
rect 4673 -4379 4719 -3905
rect 4833 -4379 4879 -3905
rect 4993 -4379 5039 -3905
rect 5153 -4379 5199 -3905
rect 5313 -4379 5359 -3905
rect 5557 -4379 5603 -3905
rect 5717 -4379 5763 -3905
rect 5877 -4379 5923 -3905
rect 6037 -4379 6083 -3905
rect 6197 -4379 6243 -3905
rect 6357 -4379 6403 -3905
rect 6517 -4379 6563 -3905
rect 6677 -4379 6723 -3905
rect 6837 -4379 6883 -3905
rect 6965 -4379 7011 -3905
rect 7125 -4379 7171 -3905
rect 7369 -4379 7415 -3905
rect 7529 -4379 7575 -3905
rect 7689 -4379 7735 -3905
rect 7849 -4379 7895 -3905
rect 8009 -4379 8055 -3905
rect 8169 -4379 8215 -3905
rect 8329 -4379 8375 -3905
rect 8489 -4379 8535 -3905
rect 8649 -4379 8695 -3905
rect 8777 -4379 8823 -3905
rect 8937 -4379 8983 -3905
rect -4076 -5015 -4030 -4541
rect -3916 -5015 -3870 -4541
rect -3788 -5015 -3742 -4541
rect -3628 -5015 -3582 -4541
rect -3468 -5015 -3422 -4541
rect -3308 -5015 -3262 -4541
rect -3148 -5015 -3102 -4541
rect -2988 -5015 -2942 -4541
rect -2828 -5015 -2782 -4541
rect -2668 -5015 -2622 -4541
rect -2508 -5015 -2462 -4541
rect -2264 -5015 -2218 -4541
rect -2104 -5015 -2058 -4541
rect -1944 -5015 -1898 -4541
rect -1784 -5015 -1738 -4541
rect -1624 -5015 -1578 -4541
rect -1464 -5015 -1418 -4541
rect -1304 -5015 -1258 -4541
rect -1144 -5015 -1098 -4541
rect -984 -5015 -938 -4541
rect -856 -5015 -810 -4541
rect -696 -5015 -650 -4541
rect 121 -5015 167 -4541
rect 281 -5015 327 -4541
rect 409 -5015 455 -4541
rect 569 -5015 615 -4541
rect 729 -5015 775 -4541
rect 889 -5015 935 -4541
rect 1049 -5015 1095 -4541
rect 1209 -5015 1255 -4541
rect 1369 -5015 1415 -4541
rect 1529 -5015 1575 -4541
rect 1689 -5015 1735 -4541
rect 1933 -5015 1979 -4541
rect 2093 -5015 2139 -4541
rect 2253 -5015 2299 -4541
rect 2413 -5015 2459 -4541
rect 2573 -5015 2619 -4541
rect 2733 -5015 2779 -4541
rect 2893 -5015 2939 -4541
rect 3053 -5015 3099 -4541
rect 3213 -5015 3259 -4541
rect 3341 -5015 3387 -4541
rect 3501 -5015 3547 -4541
rect 3745 -5015 3791 -4541
rect 3905 -5015 3951 -4541
rect 4033 -5015 4079 -4541
rect 4193 -5015 4239 -4541
rect 4353 -5015 4399 -4541
rect 4513 -5015 4559 -4541
rect 4673 -5015 4719 -4541
rect 4833 -5015 4879 -4541
rect 4993 -5015 5039 -4541
rect 5153 -5015 5199 -4541
rect 5313 -5015 5359 -4541
rect 5557 -5015 5603 -4541
rect 5717 -5015 5763 -4541
rect 5877 -5015 5923 -4541
rect 6037 -5015 6083 -4541
rect 6197 -5015 6243 -4541
rect 6357 -5015 6403 -4541
rect 6517 -5015 6563 -4541
rect 6677 -5015 6723 -4541
rect 6837 -5015 6883 -4541
rect 6965 -5015 7011 -4541
rect 7125 -5015 7171 -4541
rect 7369 -5015 7415 -4541
rect 7529 -5015 7575 -4541
rect 7689 -5015 7735 -4541
rect 7849 -5015 7895 -4541
rect 8009 -5015 8055 -4541
rect 8169 -5015 8215 -4541
rect 8329 -5015 8375 -4541
rect 8489 -5015 8535 -4541
rect 8649 -5015 8695 -4541
rect 8777 -5015 8823 -4541
rect 8937 -5015 8983 -4541
rect -4076 -5651 -4030 -5177
rect -3916 -5651 -3870 -5177
rect -3788 -5651 -3742 -5177
rect -3628 -5651 -3582 -5177
rect -3468 -5651 -3422 -5177
rect -3308 -5651 -3262 -5177
rect -3148 -5651 -3102 -5177
rect -2988 -5651 -2942 -5177
rect -2828 -5651 -2782 -5177
rect -2668 -5651 -2622 -5177
rect -2508 -5651 -2462 -5177
rect -2264 -5651 -2218 -5177
rect -2104 -5651 -2058 -5177
rect -1944 -5651 -1898 -5177
rect -1784 -5651 -1738 -5177
rect -1624 -5651 -1578 -5177
rect -1464 -5651 -1418 -5177
rect -1304 -5651 -1258 -5177
rect -1144 -5651 -1098 -5177
rect -984 -5651 -938 -5177
rect -856 -5651 -810 -5177
rect -696 -5651 -650 -5177
rect 121 -5651 167 -5177
rect 281 -5651 327 -5177
rect 409 -5651 455 -5177
rect 569 -5651 615 -5177
rect 729 -5651 775 -5177
rect 889 -5651 935 -5177
rect 1049 -5651 1095 -5177
rect 1209 -5651 1255 -5177
rect 1369 -5651 1415 -5177
rect 1529 -5651 1575 -5177
rect 1689 -5651 1735 -5177
rect 1933 -5651 1979 -5177
rect 2093 -5651 2139 -5177
rect 2253 -5651 2299 -5177
rect 2413 -5651 2459 -5177
rect 2573 -5651 2619 -5177
rect 2733 -5651 2779 -5177
rect 2893 -5651 2939 -5177
rect 3053 -5651 3099 -5177
rect 3213 -5651 3259 -5177
rect 3341 -5651 3387 -5177
rect 3501 -5651 3547 -5177
rect 3745 -5651 3791 -5177
rect 3905 -5651 3951 -5177
rect 4033 -5651 4079 -5177
rect 4193 -5651 4239 -5177
rect 4353 -5651 4399 -5177
rect 4513 -5651 4559 -5177
rect 4673 -5651 4719 -5177
rect 4833 -5651 4879 -5177
rect 4993 -5651 5039 -5177
rect 5153 -5651 5199 -5177
rect 5313 -5651 5359 -5177
rect 5557 -5651 5603 -5177
rect 5717 -5651 5763 -5177
rect 5877 -5651 5923 -5177
rect 6037 -5651 6083 -5177
rect 6197 -5651 6243 -5177
rect 6357 -5651 6403 -5177
rect 6517 -5651 6563 -5177
rect 6677 -5651 6723 -5177
rect 6837 -5651 6883 -5177
rect 6965 -5651 7011 -5177
rect 7125 -5651 7171 -5177
rect 7369 -5651 7415 -5177
rect 7529 -5651 7575 -5177
rect 7689 -5651 7735 -5177
rect 7849 -5651 7895 -5177
rect 8009 -5651 8055 -5177
rect 8169 -5651 8215 -5177
rect 8329 -5651 8375 -5177
rect 8489 -5651 8535 -5177
rect 8649 -5651 8695 -5177
rect 8777 -5651 8823 -5177
rect 8937 -5651 8983 -5177
<< psubdiff >>
rect 93 7407 1763 7420
rect 93 7361 106 7407
rect 152 7361 200 7407
rect 246 7361 294 7407
rect 340 7361 388 7407
rect 434 7361 482 7407
rect 528 7361 576 7407
rect 622 7361 670 7407
rect 716 7361 764 7407
rect 810 7361 858 7407
rect 904 7361 952 7407
rect 998 7361 1046 7407
rect 1092 7361 1140 7407
rect 1186 7361 1234 7407
rect 1280 7361 1328 7407
rect 1374 7361 1422 7407
rect 1468 7361 1516 7407
rect 1562 7361 1610 7407
rect 1656 7361 1704 7407
rect 1750 7361 1763 7407
rect 93 7348 1763 7361
rect 1905 7407 3575 7420
rect 1905 7361 1918 7407
rect 1964 7361 2012 7407
rect 2058 7361 2106 7407
rect 2152 7361 2200 7407
rect 2246 7361 2294 7407
rect 2340 7361 2388 7407
rect 2434 7361 2482 7407
rect 2528 7361 2576 7407
rect 2622 7361 2670 7407
rect 2716 7361 2764 7407
rect 2810 7361 2858 7407
rect 2904 7361 2952 7407
rect 2998 7361 3046 7407
rect 3092 7361 3140 7407
rect 3186 7361 3234 7407
rect 3280 7361 3328 7407
rect 3374 7361 3422 7407
rect 3468 7361 3516 7407
rect 3562 7361 3575 7407
rect 1905 7348 3575 7361
rect 3717 7407 5387 7420
rect 3717 7361 3730 7407
rect 3776 7361 3824 7407
rect 3870 7361 3918 7407
rect 3964 7361 4012 7407
rect 4058 7361 4106 7407
rect 4152 7361 4200 7407
rect 4246 7361 4294 7407
rect 4340 7361 4388 7407
rect 4434 7361 4482 7407
rect 4528 7361 4576 7407
rect 4622 7361 4670 7407
rect 4716 7361 4764 7407
rect 4810 7361 4858 7407
rect 4904 7361 4952 7407
rect 4998 7361 5046 7407
rect 5092 7361 5140 7407
rect 5186 7361 5234 7407
rect 5280 7361 5328 7407
rect 5374 7361 5387 7407
rect 3717 7348 5387 7361
rect 5529 7407 7199 7420
rect 5529 7361 5542 7407
rect 5588 7361 5636 7407
rect 5682 7361 5730 7407
rect 5776 7361 5824 7407
rect 5870 7361 5918 7407
rect 5964 7361 6012 7407
rect 6058 7361 6106 7407
rect 6152 7361 6200 7407
rect 6246 7361 6294 7407
rect 6340 7361 6388 7407
rect 6434 7361 6482 7407
rect 6528 7361 6576 7407
rect 6622 7361 6670 7407
rect 6716 7361 6764 7407
rect 6810 7361 6858 7407
rect 6904 7361 6952 7407
rect 6998 7361 7046 7407
rect 7092 7361 7140 7407
rect 7186 7361 7199 7407
rect 5529 7348 7199 7361
rect 7341 7407 9011 7420
rect 7341 7361 7354 7407
rect 7400 7361 7448 7407
rect 7494 7361 7542 7407
rect 7588 7361 7636 7407
rect 7682 7361 7730 7407
rect 7776 7361 7824 7407
rect 7870 7361 7918 7407
rect 7964 7361 8012 7407
rect 8058 7361 8106 7407
rect 8152 7361 8200 7407
rect 8246 7361 8294 7407
rect 8340 7361 8388 7407
rect 8434 7361 8482 7407
rect 8528 7361 8576 7407
rect 8622 7361 8670 7407
rect 8716 7361 8764 7407
rect 8810 7361 8858 7407
rect 8904 7361 8952 7407
rect 8998 7361 9011 7407
rect 7341 7348 9011 7361
rect -4826 2888 -4566 2901
rect -4826 2842 -4813 2888
rect -4767 2842 -4719 2888
rect -4673 2842 -4625 2888
rect -4579 2842 -4566 2888
rect -4826 2829 -4566 2842
rect -4227 2888 -3873 2901
rect -4227 2842 -4214 2888
rect -4168 2842 -4120 2888
rect -4074 2842 -4026 2888
rect -3980 2842 -3932 2888
rect -3886 2842 -3873 2888
rect -4227 2829 -3873 2842
rect -3545 2888 -2905 2901
rect -3545 2842 -3532 2888
rect -3486 2842 -3438 2888
rect -3392 2842 -3344 2888
rect -3298 2842 -3250 2888
rect -3204 2842 -3156 2888
rect -3110 2842 -3062 2888
rect -3016 2842 -2968 2888
rect -2922 2842 -2905 2888
rect -3545 2829 -2905 2842
rect -2759 2888 -2119 2901
rect -2759 2842 -2746 2888
rect -2700 2842 -2652 2888
rect -2606 2842 -2558 2888
rect -2512 2842 -2464 2888
rect -2418 2842 -2370 2888
rect -2324 2842 -2276 2888
rect -2230 2842 -2182 2888
rect -2136 2842 -2119 2888
rect -2759 2829 -2119 2842
rect -1973 2888 -1333 2901
rect -1973 2842 -1960 2888
rect -1914 2842 -1866 2888
rect -1820 2842 -1772 2888
rect -1726 2842 -1678 2888
rect -1632 2842 -1584 2888
rect -1538 2842 -1490 2888
rect -1444 2842 -1396 2888
rect -1350 2842 -1333 2888
rect -1973 2829 -1333 2842
rect -1177 2888 -917 2901
rect -1177 2842 -1164 2888
rect -1118 2842 -1070 2888
rect -1024 2842 -976 2888
rect -930 2842 -917 2888
rect -1177 2829 -917 2842
rect -4826 1178 -4566 1191
rect -4826 1132 -4813 1178
rect -4767 1132 -4719 1178
rect -4673 1132 -4625 1178
rect -4579 1132 -4566 1178
rect -4826 1119 -4566 1132
rect -4227 1178 -3873 1191
rect -4227 1132 -4214 1178
rect -4168 1132 -4120 1178
rect -4074 1132 -4026 1178
rect -3980 1132 -3932 1178
rect -3886 1132 -3873 1178
rect -4227 1119 -3873 1132
rect -3545 1178 -2905 1191
rect -3545 1132 -3532 1178
rect -3486 1132 -3438 1178
rect -3392 1132 -3344 1178
rect -3298 1132 -3250 1178
rect -3204 1132 -3156 1178
rect -3110 1132 -3062 1178
rect -3016 1132 -2968 1178
rect -2922 1132 -2905 1178
rect -3545 1119 -2905 1132
rect -2759 1178 -2119 1191
rect -2759 1132 -2746 1178
rect -2700 1132 -2652 1178
rect -2606 1132 -2558 1178
rect -2512 1132 -2464 1178
rect -2418 1132 -2370 1178
rect -2324 1132 -2276 1178
rect -2230 1132 -2182 1178
rect -2136 1132 -2119 1178
rect -2759 1119 -2119 1132
rect -1973 1178 -1333 1191
rect -1973 1132 -1960 1178
rect -1914 1132 -1866 1178
rect -1820 1132 -1772 1178
rect -1726 1132 -1678 1178
rect -1632 1132 -1584 1178
rect -1538 1132 -1490 1178
rect -1444 1132 -1396 1178
rect -1350 1132 -1333 1178
rect -1973 1119 -1333 1132
rect -1177 1178 -917 1191
rect -1177 1132 -1164 1178
rect -1118 1132 -1070 1178
rect -1024 1132 -976 1178
rect -930 1132 -917 1178
rect -1177 1119 -917 1132
rect 93 79 1763 92
rect 93 33 106 79
rect 152 33 200 79
rect 246 33 294 79
rect 340 33 388 79
rect 434 33 482 79
rect 528 33 576 79
rect 622 33 670 79
rect 716 33 764 79
rect 810 33 858 79
rect 904 33 952 79
rect 998 33 1046 79
rect 1092 33 1140 79
rect 1186 33 1234 79
rect 1280 33 1328 79
rect 1374 33 1422 79
rect 1468 33 1516 79
rect 1562 33 1610 79
rect 1656 33 1704 79
rect 1750 33 1763 79
rect 93 20 1763 33
rect 1905 79 3575 92
rect 1905 33 1918 79
rect 1964 33 2012 79
rect 2058 33 2106 79
rect 2152 33 2200 79
rect 2246 33 2294 79
rect 2340 33 2388 79
rect 2434 33 2482 79
rect 2528 33 2576 79
rect 2622 33 2670 79
rect 2716 33 2764 79
rect 2810 33 2858 79
rect 2904 33 2952 79
rect 2998 33 3046 79
rect 3092 33 3140 79
rect 3186 33 3234 79
rect 3280 33 3328 79
rect 3374 33 3422 79
rect 3468 33 3516 79
rect 3562 33 3575 79
rect 1905 20 3575 33
rect 3717 79 5387 92
rect 3717 33 3730 79
rect 3776 33 3824 79
rect 3870 33 3918 79
rect 3964 33 4012 79
rect 4058 33 4106 79
rect 4152 33 4200 79
rect 4246 33 4294 79
rect 4340 33 4388 79
rect 4434 33 4482 79
rect 4528 33 4576 79
rect 4622 33 4670 79
rect 4716 33 4764 79
rect 4810 33 4858 79
rect 4904 33 4952 79
rect 4998 33 5046 79
rect 5092 33 5140 79
rect 5186 33 5234 79
rect 5280 33 5328 79
rect 5374 33 5387 79
rect 3717 20 5387 33
rect 5529 79 7199 92
rect 5529 33 5542 79
rect 5588 33 5636 79
rect 5682 33 5730 79
rect 5776 33 5824 79
rect 5870 33 5918 79
rect 5964 33 6012 79
rect 6058 33 6106 79
rect 6152 33 6200 79
rect 6246 33 6294 79
rect 6340 33 6388 79
rect 6434 33 6482 79
rect 6528 33 6576 79
rect 6622 33 6670 79
rect 6716 33 6764 79
rect 6810 33 6858 79
rect 6904 33 6952 79
rect 6998 33 7046 79
rect 7092 33 7140 79
rect 7186 33 7199 79
rect 5529 20 7199 33
rect 7341 79 9011 92
rect 7341 33 7354 79
rect 7400 33 7448 79
rect 7494 33 7542 79
rect 7588 33 7636 79
rect 7682 33 7730 79
rect 7776 33 7824 79
rect 7870 33 7918 79
rect 7964 33 8012 79
rect 8058 33 8106 79
rect 8152 33 8200 79
rect 8246 33 8294 79
rect 8340 33 8388 79
rect 8434 33 8482 79
rect 8528 33 8576 79
rect 8622 33 8670 79
rect 8716 33 8764 79
rect 8810 33 8858 79
rect 8904 33 8952 79
rect 8998 33 9011 79
rect 7341 20 9011 33
rect -4826 -532 -4566 -519
rect -4826 -578 -4813 -532
rect -4767 -578 -4719 -532
rect -4673 -578 -4625 -532
rect -4579 -578 -4566 -532
rect -4826 -591 -4566 -578
rect -4227 -532 -3873 -519
rect -4227 -578 -4214 -532
rect -4168 -578 -4120 -532
rect -4074 -578 -4026 -532
rect -3980 -578 -3932 -532
rect -3886 -578 -3873 -532
rect -4227 -591 -3873 -578
rect -3545 -532 -2905 -519
rect -3545 -578 -3532 -532
rect -3486 -578 -3438 -532
rect -3392 -578 -3344 -532
rect -3298 -578 -3250 -532
rect -3204 -578 -3156 -532
rect -3110 -578 -3062 -532
rect -3016 -578 -2968 -532
rect -2922 -578 -2905 -532
rect -3545 -591 -2905 -578
rect -2759 -532 -2119 -519
rect -2759 -578 -2746 -532
rect -2700 -578 -2652 -532
rect -2606 -578 -2558 -532
rect -2512 -578 -2464 -532
rect -2418 -578 -2370 -532
rect -2324 -578 -2276 -532
rect -2230 -578 -2182 -532
rect -2136 -578 -2119 -532
rect -2759 -591 -2119 -578
rect -1973 -532 -1333 -519
rect -1973 -578 -1960 -532
rect -1914 -578 -1866 -532
rect -1820 -578 -1772 -532
rect -1726 -578 -1678 -532
rect -1632 -578 -1584 -532
rect -1538 -578 -1490 -532
rect -1444 -578 -1396 -532
rect -1350 -578 -1333 -532
rect -1973 -591 -1333 -578
rect -1177 -532 -917 -519
rect -1177 -578 -1164 -532
rect -1118 -578 -1070 -532
rect -1024 -578 -976 -532
rect -930 -578 -917 -532
rect -1177 -591 -917 -578
rect -4104 -7249 -2434 -7236
rect -4104 -7295 -4091 -7249
rect -4045 -7295 -3997 -7249
rect -3951 -7295 -3903 -7249
rect -3857 -7295 -3809 -7249
rect -3763 -7295 -3715 -7249
rect -3669 -7295 -3621 -7249
rect -3575 -7295 -3527 -7249
rect -3481 -7295 -3433 -7249
rect -3387 -7295 -3339 -7249
rect -3293 -7295 -3245 -7249
rect -3199 -7295 -3151 -7249
rect -3105 -7295 -3057 -7249
rect -3011 -7295 -2963 -7249
rect -2917 -7295 -2869 -7249
rect -2823 -7295 -2775 -7249
rect -2729 -7295 -2681 -7249
rect -2635 -7295 -2587 -7249
rect -2541 -7295 -2493 -7249
rect -2447 -7295 -2434 -7249
rect -4104 -7308 -2434 -7295
rect -2292 -7249 -622 -7236
rect -2292 -7295 -2279 -7249
rect -2233 -7295 -2185 -7249
rect -2139 -7295 -2091 -7249
rect -2045 -7295 -1997 -7249
rect -1951 -7295 -1903 -7249
rect -1857 -7295 -1809 -7249
rect -1763 -7295 -1715 -7249
rect -1669 -7295 -1621 -7249
rect -1575 -7295 -1527 -7249
rect -1481 -7295 -1433 -7249
rect -1387 -7295 -1339 -7249
rect -1293 -7295 -1245 -7249
rect -1199 -7295 -1151 -7249
rect -1105 -7295 -1057 -7249
rect -1011 -7295 -963 -7249
rect -917 -7295 -869 -7249
rect -823 -7295 -775 -7249
rect -729 -7295 -681 -7249
rect -635 -7295 -622 -7249
rect -2292 -7308 -622 -7295
rect 93 -7249 1763 -7236
rect 93 -7295 106 -7249
rect 152 -7295 200 -7249
rect 246 -7295 294 -7249
rect 340 -7295 388 -7249
rect 434 -7295 482 -7249
rect 528 -7295 576 -7249
rect 622 -7295 670 -7249
rect 716 -7295 764 -7249
rect 810 -7295 858 -7249
rect 904 -7295 952 -7249
rect 998 -7295 1046 -7249
rect 1092 -7295 1140 -7249
rect 1186 -7295 1234 -7249
rect 1280 -7295 1328 -7249
rect 1374 -7295 1422 -7249
rect 1468 -7295 1516 -7249
rect 1562 -7295 1610 -7249
rect 1656 -7295 1704 -7249
rect 1750 -7295 1763 -7249
rect 93 -7308 1763 -7295
rect 1905 -7249 3575 -7236
rect 1905 -7295 1918 -7249
rect 1964 -7295 2012 -7249
rect 2058 -7295 2106 -7249
rect 2152 -7295 2200 -7249
rect 2246 -7295 2294 -7249
rect 2340 -7295 2388 -7249
rect 2434 -7295 2482 -7249
rect 2528 -7295 2576 -7249
rect 2622 -7295 2670 -7249
rect 2716 -7295 2764 -7249
rect 2810 -7295 2858 -7249
rect 2904 -7295 2952 -7249
rect 2998 -7295 3046 -7249
rect 3092 -7295 3140 -7249
rect 3186 -7295 3234 -7249
rect 3280 -7295 3328 -7249
rect 3374 -7295 3422 -7249
rect 3468 -7295 3516 -7249
rect 3562 -7295 3575 -7249
rect 1905 -7308 3575 -7295
rect 3717 -7249 5387 -7236
rect 3717 -7295 3730 -7249
rect 3776 -7295 3824 -7249
rect 3870 -7295 3918 -7249
rect 3964 -7295 4012 -7249
rect 4058 -7295 4106 -7249
rect 4152 -7295 4200 -7249
rect 4246 -7295 4294 -7249
rect 4340 -7295 4388 -7249
rect 4434 -7295 4482 -7249
rect 4528 -7295 4576 -7249
rect 4622 -7295 4670 -7249
rect 4716 -7295 4764 -7249
rect 4810 -7295 4858 -7249
rect 4904 -7295 4952 -7249
rect 4998 -7295 5046 -7249
rect 5092 -7295 5140 -7249
rect 5186 -7295 5234 -7249
rect 5280 -7295 5328 -7249
rect 5374 -7295 5387 -7249
rect 3717 -7308 5387 -7295
rect 5529 -7249 7199 -7236
rect 5529 -7295 5542 -7249
rect 5588 -7295 5636 -7249
rect 5682 -7295 5730 -7249
rect 5776 -7295 5824 -7249
rect 5870 -7295 5918 -7249
rect 5964 -7295 6012 -7249
rect 6058 -7295 6106 -7249
rect 6152 -7295 6200 -7249
rect 6246 -7295 6294 -7249
rect 6340 -7295 6388 -7249
rect 6434 -7295 6482 -7249
rect 6528 -7295 6576 -7249
rect 6622 -7295 6670 -7249
rect 6716 -7295 6764 -7249
rect 6810 -7295 6858 -7249
rect 6904 -7295 6952 -7249
rect 6998 -7295 7046 -7249
rect 7092 -7295 7140 -7249
rect 7186 -7295 7199 -7249
rect 5529 -7308 7199 -7295
rect 7341 -7249 9011 -7236
rect 7341 -7295 7354 -7249
rect 7400 -7295 7448 -7249
rect 7494 -7295 7542 -7249
rect 7588 -7295 7636 -7249
rect 7682 -7295 7730 -7249
rect 7776 -7295 7824 -7249
rect 7870 -7295 7918 -7249
rect 7964 -7295 8012 -7249
rect 8058 -7295 8106 -7249
rect 8152 -7295 8200 -7249
rect 8246 -7295 8294 -7249
rect 8340 -7295 8388 -7249
rect 8434 -7295 8482 -7249
rect 8528 -7295 8576 -7249
rect 8622 -7295 8670 -7249
rect 8716 -7295 8764 -7249
rect 8810 -7295 8858 -7249
rect 8904 -7295 8952 -7249
rect 8998 -7295 9011 -7249
rect 7341 -7308 9011 -7295
<< nsubdiff >>
rect -4873 3743 -4519 3756
rect -4873 3697 -4860 3743
rect -4814 3697 -4766 3743
rect -4720 3697 -4672 3743
rect -4626 3697 -4578 3743
rect -4532 3697 -4519 3743
rect -4873 3684 -4519 3697
rect -4462 3743 -3638 3756
rect -4462 3697 -4449 3743
rect -4403 3697 -4355 3743
rect -4309 3697 -4261 3743
rect -4215 3697 -4167 3743
rect -4121 3697 -4073 3743
rect -4027 3697 -3979 3743
rect -3933 3697 -3885 3743
rect -3839 3697 -3791 3743
rect -3745 3697 -3697 3743
rect -3651 3697 -3638 3743
rect -4462 3684 -3638 3697
rect -3582 3743 -2852 3756
rect -3582 3697 -3569 3743
rect -3523 3697 -3475 3743
rect -3429 3697 -3381 3743
rect -3335 3697 -3287 3743
rect -3241 3697 -3193 3743
rect -3147 3697 -3099 3743
rect -3053 3697 -3005 3743
rect -2959 3697 -2911 3743
rect -2865 3697 -2852 3743
rect -3582 3684 -2852 3697
rect -2796 3743 -2066 3756
rect -2796 3697 -2783 3743
rect -2737 3697 -2689 3743
rect -2643 3697 -2595 3743
rect -2549 3697 -2501 3743
rect -2455 3697 -2407 3743
rect -2361 3697 -2313 3743
rect -2267 3697 -2219 3743
rect -2173 3697 -2125 3743
rect -2079 3697 -2066 3743
rect -2796 3684 -2066 3697
rect -2010 3743 -1280 3756
rect -2010 3697 -1997 3743
rect -1951 3697 -1903 3743
rect -1857 3697 -1809 3743
rect -1763 3697 -1715 3743
rect -1669 3697 -1621 3743
rect -1575 3697 -1527 3743
rect -1481 3697 -1433 3743
rect -1387 3697 -1339 3743
rect -1293 3697 -1280 3743
rect -2010 3684 -1280 3697
rect -1224 3743 -870 3756
rect -1224 3697 -1211 3743
rect -1165 3697 -1117 3743
rect -1071 3697 -1023 3743
rect -977 3697 -929 3743
rect -883 3697 -870 3743
rect -1224 3684 -870 3697
rect 46 3743 9058 3756
rect 46 3697 59 3743
rect 105 3697 153 3743
rect 199 3697 247 3743
rect 293 3697 341 3743
rect 387 3697 435 3743
rect 481 3697 529 3743
rect 575 3697 623 3743
rect 669 3697 717 3743
rect 763 3697 811 3743
rect 857 3697 905 3743
rect 951 3697 999 3743
rect 1045 3697 1093 3743
rect 1139 3697 1187 3743
rect 1233 3697 1281 3743
rect 1327 3697 1375 3743
rect 1421 3697 1469 3743
rect 1515 3697 1563 3743
rect 1609 3697 1657 3743
rect 1703 3697 1751 3743
rect 1797 3697 1871 3743
rect 1917 3697 1965 3743
rect 2011 3697 2059 3743
rect 2105 3697 2153 3743
rect 2199 3697 2247 3743
rect 2293 3697 2341 3743
rect 2387 3697 2435 3743
rect 2481 3697 2529 3743
rect 2575 3697 2623 3743
rect 2669 3697 2717 3743
rect 2763 3697 2811 3743
rect 2857 3697 2905 3743
rect 2951 3697 2999 3743
rect 3045 3697 3093 3743
rect 3139 3697 3187 3743
rect 3233 3697 3281 3743
rect 3327 3697 3375 3743
rect 3421 3697 3469 3743
rect 3515 3697 3563 3743
rect 3609 3697 3683 3743
rect 3729 3697 3777 3743
rect 3823 3697 3871 3743
rect 3917 3697 3965 3743
rect 4011 3697 4059 3743
rect 4105 3697 4153 3743
rect 4199 3697 4247 3743
rect 4293 3697 4341 3743
rect 4387 3697 4435 3743
rect 4481 3697 4529 3743
rect 4575 3697 4623 3743
rect 4669 3697 4717 3743
rect 4763 3697 4811 3743
rect 4857 3697 4905 3743
rect 4951 3697 4999 3743
rect 5045 3697 5093 3743
rect 5139 3697 5187 3743
rect 5233 3697 5281 3743
rect 5327 3697 5375 3743
rect 5421 3697 5495 3743
rect 5541 3697 5589 3743
rect 5635 3697 5683 3743
rect 5729 3697 5777 3743
rect 5823 3697 5871 3743
rect 5917 3697 5965 3743
rect 6011 3697 6059 3743
rect 6105 3697 6153 3743
rect 6199 3697 6247 3743
rect 6293 3697 6341 3743
rect 6387 3697 6435 3743
rect 6481 3697 6529 3743
rect 6575 3697 6623 3743
rect 6669 3697 6717 3743
rect 6763 3697 6811 3743
rect 6857 3697 6905 3743
rect 6951 3697 6999 3743
rect 7045 3697 7093 3743
rect 7139 3697 7187 3743
rect 7233 3697 7307 3743
rect 7353 3697 7401 3743
rect 7447 3697 7495 3743
rect 7541 3697 7589 3743
rect 7635 3697 7683 3743
rect 7729 3697 7777 3743
rect 7823 3697 7871 3743
rect 7917 3697 7965 3743
rect 8011 3697 8059 3743
rect 8105 3697 8153 3743
rect 8199 3697 8247 3743
rect 8293 3697 8341 3743
rect 8387 3697 8435 3743
rect 8481 3697 8529 3743
rect 8575 3697 8623 3743
rect 8669 3697 8717 3743
rect 8763 3697 8811 3743
rect 8857 3697 8905 3743
rect 8951 3697 8999 3743
rect 9045 3697 9058 3743
rect 46 3684 9058 3697
rect -4462 2033 -3638 2046
rect -4462 1987 -4449 2033
rect -4403 1987 -4355 2033
rect -4309 1987 -4261 2033
rect -4215 1987 -4167 2033
rect -4121 1987 -4073 2033
rect -4027 1987 -3979 2033
rect -3933 1987 -3885 2033
rect -3839 1987 -3791 2033
rect -3745 1987 -3697 2033
rect -3651 1987 -3638 2033
rect -4462 1974 -3638 1987
rect -3582 2033 -2852 2046
rect -3582 1987 -3569 2033
rect -3523 1987 -3475 2033
rect -3429 1987 -3381 2033
rect -3335 1987 -3287 2033
rect -3241 1987 -3193 2033
rect -3147 1987 -3099 2033
rect -3053 1987 -3005 2033
rect -2959 1987 -2911 2033
rect -2865 1987 -2852 2033
rect -3582 1974 -2852 1987
rect -2796 2033 -2066 2046
rect -2796 1987 -2783 2033
rect -2737 1987 -2689 2033
rect -2643 1987 -2595 2033
rect -2549 1987 -2501 2033
rect -2455 1987 -2407 2033
rect -2361 1987 -2313 2033
rect -2267 1987 -2219 2033
rect -2173 1987 -2125 2033
rect -2079 1987 -2066 2033
rect -2796 1974 -2066 1987
rect -2010 2033 -1280 2046
rect -2010 1987 -1997 2033
rect -1951 1987 -1903 2033
rect -1857 1987 -1809 2033
rect -1763 1987 -1715 2033
rect -1669 1987 -1621 2033
rect -1575 1987 -1527 2033
rect -1481 1987 -1433 2033
rect -1387 1987 -1339 2033
rect -1293 1987 -1280 2033
rect -2010 1974 -1280 1987
rect -1224 2033 -870 2046
rect -1224 1987 -1211 2033
rect -1165 1987 -1117 2033
rect -1071 1987 -1023 2033
rect -977 1987 -929 2033
rect -883 1987 -870 2033
rect -1224 1974 -870 1987
rect -4873 323 -4519 336
rect -4873 277 -4860 323
rect -4814 277 -4766 323
rect -4720 277 -4672 323
rect -4626 277 -4578 323
rect -4532 277 -4519 323
rect -4873 264 -4519 277
rect -4462 323 -3638 336
rect -4462 277 -4449 323
rect -4403 277 -4355 323
rect -4309 277 -4261 323
rect -4215 277 -4167 323
rect -4121 277 -4073 323
rect -4027 277 -3979 323
rect -3933 277 -3885 323
rect -3839 277 -3791 323
rect -3745 277 -3697 323
rect -3651 277 -3638 323
rect -4462 264 -3638 277
rect -3582 323 -2852 336
rect -3582 277 -3569 323
rect -3523 277 -3475 323
rect -3429 277 -3381 323
rect -3335 277 -3287 323
rect -3241 277 -3193 323
rect -3147 277 -3099 323
rect -3053 277 -3005 323
rect -2959 277 -2911 323
rect -2865 277 -2852 323
rect -3582 264 -2852 277
rect -2796 323 -2066 336
rect -2796 277 -2783 323
rect -2737 277 -2689 323
rect -2643 277 -2595 323
rect -2549 277 -2501 323
rect -2455 277 -2407 323
rect -2361 277 -2313 323
rect -2267 277 -2219 323
rect -2173 277 -2125 323
rect -2079 277 -2066 323
rect -2796 264 -2066 277
rect -2010 323 -1280 336
rect -2010 277 -1997 323
rect -1951 277 -1903 323
rect -1857 277 -1809 323
rect -1763 277 -1715 323
rect -1669 277 -1621 323
rect -1575 277 -1527 323
rect -1481 277 -1433 323
rect -1387 277 -1339 323
rect -1293 277 -1280 323
rect -2010 264 -1280 277
rect -1224 323 -870 336
rect -1224 277 -1211 323
rect -1165 277 -1117 323
rect -1071 277 -1023 323
rect -977 277 -929 323
rect -883 277 -870 323
rect -1224 264 -870 277
rect -4462 -1387 -3638 -1374
rect -4462 -1433 -4449 -1387
rect -4403 -1433 -4355 -1387
rect -4309 -1433 -4261 -1387
rect -4215 -1433 -4167 -1387
rect -4121 -1433 -4073 -1387
rect -4027 -1433 -3979 -1387
rect -3933 -1433 -3885 -1387
rect -3839 -1433 -3791 -1387
rect -3745 -1433 -3697 -1387
rect -3651 -1433 -3638 -1387
rect -4462 -1446 -3638 -1433
rect -3582 -1387 -2852 -1374
rect -3582 -1433 -3569 -1387
rect -3523 -1433 -3475 -1387
rect -3429 -1433 -3381 -1387
rect -3335 -1433 -3287 -1387
rect -3241 -1433 -3193 -1387
rect -3147 -1433 -3099 -1387
rect -3053 -1433 -3005 -1387
rect -2959 -1433 -2911 -1387
rect -2865 -1433 -2852 -1387
rect -3582 -1446 -2852 -1433
rect -2796 -1387 -2066 -1374
rect -2796 -1433 -2783 -1387
rect -2737 -1433 -2689 -1387
rect -2643 -1433 -2595 -1387
rect -2549 -1433 -2501 -1387
rect -2455 -1433 -2407 -1387
rect -2361 -1433 -2313 -1387
rect -2267 -1433 -2219 -1387
rect -2173 -1433 -2125 -1387
rect -2079 -1433 -2066 -1387
rect -2796 -1446 -2066 -1433
rect -2010 -1387 -1280 -1374
rect -2010 -1433 -1997 -1387
rect -1951 -1433 -1903 -1387
rect -1857 -1433 -1809 -1387
rect -1763 -1433 -1715 -1387
rect -1669 -1433 -1621 -1387
rect -1575 -1433 -1527 -1387
rect -1481 -1433 -1433 -1387
rect -1387 -1433 -1339 -1387
rect -1293 -1433 -1280 -1387
rect -2010 -1446 -1280 -1433
rect -1224 -1387 -870 -1374
rect -1224 -1433 -1211 -1387
rect -1165 -1433 -1117 -1387
rect -1071 -1433 -1023 -1387
rect -977 -1433 -929 -1387
rect -883 -1433 -870 -1387
rect -1224 -1446 -870 -1433
rect -4151 -3585 -575 -3572
rect -4151 -3631 -4138 -3585
rect -4092 -3631 -4044 -3585
rect -3998 -3631 -3950 -3585
rect -3904 -3631 -3856 -3585
rect -3810 -3631 -3762 -3585
rect -3716 -3631 -3668 -3585
rect -3622 -3631 -3574 -3585
rect -3528 -3631 -3480 -3585
rect -3434 -3631 -3386 -3585
rect -3340 -3631 -3292 -3585
rect -3246 -3631 -3198 -3585
rect -3152 -3631 -3104 -3585
rect -3058 -3631 -3010 -3585
rect -2964 -3631 -2916 -3585
rect -2870 -3631 -2822 -3585
rect -2776 -3631 -2728 -3585
rect -2682 -3631 -2634 -3585
rect -2588 -3631 -2540 -3585
rect -2494 -3631 -2446 -3585
rect -2400 -3631 -2326 -3585
rect -2280 -3631 -2232 -3585
rect -2186 -3631 -2138 -3585
rect -2092 -3631 -2044 -3585
rect -1998 -3631 -1950 -3585
rect -1904 -3631 -1856 -3585
rect -1810 -3631 -1762 -3585
rect -1716 -3631 -1668 -3585
rect -1622 -3631 -1574 -3585
rect -1528 -3631 -1480 -3585
rect -1434 -3631 -1386 -3585
rect -1340 -3631 -1292 -3585
rect -1246 -3631 -1198 -3585
rect -1152 -3631 -1104 -3585
rect -1058 -3631 -1010 -3585
rect -964 -3631 -916 -3585
rect -870 -3631 -822 -3585
rect -776 -3631 -728 -3585
rect -682 -3631 -634 -3585
rect -588 -3631 -575 -3585
rect -4151 -3644 -575 -3631
rect 46 -3585 9058 -3572
rect 46 -3631 59 -3585
rect 105 -3631 153 -3585
rect 199 -3631 247 -3585
rect 293 -3631 341 -3585
rect 387 -3631 435 -3585
rect 481 -3631 529 -3585
rect 575 -3631 623 -3585
rect 669 -3631 717 -3585
rect 763 -3631 811 -3585
rect 857 -3631 905 -3585
rect 951 -3631 999 -3585
rect 1045 -3631 1093 -3585
rect 1139 -3631 1187 -3585
rect 1233 -3631 1281 -3585
rect 1327 -3631 1375 -3585
rect 1421 -3631 1469 -3585
rect 1515 -3631 1563 -3585
rect 1609 -3631 1657 -3585
rect 1703 -3631 1751 -3585
rect 1797 -3631 1871 -3585
rect 1917 -3631 1965 -3585
rect 2011 -3631 2059 -3585
rect 2105 -3631 2153 -3585
rect 2199 -3631 2247 -3585
rect 2293 -3631 2341 -3585
rect 2387 -3631 2435 -3585
rect 2481 -3631 2529 -3585
rect 2575 -3631 2623 -3585
rect 2669 -3631 2717 -3585
rect 2763 -3631 2811 -3585
rect 2857 -3631 2905 -3585
rect 2951 -3631 2999 -3585
rect 3045 -3631 3093 -3585
rect 3139 -3631 3187 -3585
rect 3233 -3631 3281 -3585
rect 3327 -3631 3375 -3585
rect 3421 -3631 3469 -3585
rect 3515 -3631 3563 -3585
rect 3609 -3631 3683 -3585
rect 3729 -3631 3777 -3585
rect 3823 -3631 3871 -3585
rect 3917 -3631 3965 -3585
rect 4011 -3631 4059 -3585
rect 4105 -3631 4153 -3585
rect 4199 -3631 4247 -3585
rect 4293 -3631 4341 -3585
rect 4387 -3631 4435 -3585
rect 4481 -3631 4529 -3585
rect 4575 -3631 4623 -3585
rect 4669 -3631 4717 -3585
rect 4763 -3631 4811 -3585
rect 4857 -3631 4905 -3585
rect 4951 -3631 4999 -3585
rect 5045 -3631 5093 -3585
rect 5139 -3631 5187 -3585
rect 5233 -3631 5281 -3585
rect 5327 -3631 5375 -3585
rect 5421 -3631 5495 -3585
rect 5541 -3631 5589 -3585
rect 5635 -3631 5683 -3585
rect 5729 -3631 5777 -3585
rect 5823 -3631 5871 -3585
rect 5917 -3631 5965 -3585
rect 6011 -3631 6059 -3585
rect 6105 -3631 6153 -3585
rect 6199 -3631 6247 -3585
rect 6293 -3631 6341 -3585
rect 6387 -3631 6435 -3585
rect 6481 -3631 6529 -3585
rect 6575 -3631 6623 -3585
rect 6669 -3631 6717 -3585
rect 6763 -3631 6811 -3585
rect 6857 -3631 6905 -3585
rect 6951 -3631 6999 -3585
rect 7045 -3631 7093 -3585
rect 7139 -3631 7187 -3585
rect 7233 -3631 7307 -3585
rect 7353 -3631 7401 -3585
rect 7447 -3631 7495 -3585
rect 7541 -3631 7589 -3585
rect 7635 -3631 7683 -3585
rect 7729 -3631 7777 -3585
rect 7823 -3631 7871 -3585
rect 7917 -3631 7965 -3585
rect 8011 -3631 8059 -3585
rect 8105 -3631 8153 -3585
rect 8199 -3631 8247 -3585
rect 8293 -3631 8341 -3585
rect 8387 -3631 8435 -3585
rect 8481 -3631 8529 -3585
rect 8575 -3631 8623 -3585
rect 8669 -3631 8717 -3585
rect 8763 -3631 8811 -3585
rect 8857 -3631 8905 -3585
rect 8951 -3631 8999 -3585
rect 9045 -3631 9058 -3585
rect 46 -3644 9058 -3631
rect -2387 -3645 -2339 -3644
<< psubdiffcont >>
rect 106 7361 152 7407
rect 200 7361 246 7407
rect 294 7361 340 7407
rect 388 7361 434 7407
rect 482 7361 528 7407
rect 576 7361 622 7407
rect 670 7361 716 7407
rect 764 7361 810 7407
rect 858 7361 904 7407
rect 952 7361 998 7407
rect 1046 7361 1092 7407
rect 1140 7361 1186 7407
rect 1234 7361 1280 7407
rect 1328 7361 1374 7407
rect 1422 7361 1468 7407
rect 1516 7361 1562 7407
rect 1610 7361 1656 7407
rect 1704 7361 1750 7407
rect 1918 7361 1964 7407
rect 2012 7361 2058 7407
rect 2106 7361 2152 7407
rect 2200 7361 2246 7407
rect 2294 7361 2340 7407
rect 2388 7361 2434 7407
rect 2482 7361 2528 7407
rect 2576 7361 2622 7407
rect 2670 7361 2716 7407
rect 2764 7361 2810 7407
rect 2858 7361 2904 7407
rect 2952 7361 2998 7407
rect 3046 7361 3092 7407
rect 3140 7361 3186 7407
rect 3234 7361 3280 7407
rect 3328 7361 3374 7407
rect 3422 7361 3468 7407
rect 3516 7361 3562 7407
rect 3730 7361 3776 7407
rect 3824 7361 3870 7407
rect 3918 7361 3964 7407
rect 4012 7361 4058 7407
rect 4106 7361 4152 7407
rect 4200 7361 4246 7407
rect 4294 7361 4340 7407
rect 4388 7361 4434 7407
rect 4482 7361 4528 7407
rect 4576 7361 4622 7407
rect 4670 7361 4716 7407
rect 4764 7361 4810 7407
rect 4858 7361 4904 7407
rect 4952 7361 4998 7407
rect 5046 7361 5092 7407
rect 5140 7361 5186 7407
rect 5234 7361 5280 7407
rect 5328 7361 5374 7407
rect 5542 7361 5588 7407
rect 5636 7361 5682 7407
rect 5730 7361 5776 7407
rect 5824 7361 5870 7407
rect 5918 7361 5964 7407
rect 6012 7361 6058 7407
rect 6106 7361 6152 7407
rect 6200 7361 6246 7407
rect 6294 7361 6340 7407
rect 6388 7361 6434 7407
rect 6482 7361 6528 7407
rect 6576 7361 6622 7407
rect 6670 7361 6716 7407
rect 6764 7361 6810 7407
rect 6858 7361 6904 7407
rect 6952 7361 6998 7407
rect 7046 7361 7092 7407
rect 7140 7361 7186 7407
rect 7354 7361 7400 7407
rect 7448 7361 7494 7407
rect 7542 7361 7588 7407
rect 7636 7361 7682 7407
rect 7730 7361 7776 7407
rect 7824 7361 7870 7407
rect 7918 7361 7964 7407
rect 8012 7361 8058 7407
rect 8106 7361 8152 7407
rect 8200 7361 8246 7407
rect 8294 7361 8340 7407
rect 8388 7361 8434 7407
rect 8482 7361 8528 7407
rect 8576 7361 8622 7407
rect 8670 7361 8716 7407
rect 8764 7361 8810 7407
rect 8858 7361 8904 7407
rect 8952 7361 8998 7407
rect -4813 2842 -4767 2888
rect -4719 2842 -4673 2888
rect -4625 2842 -4579 2888
rect -4214 2842 -4168 2888
rect -4120 2842 -4074 2888
rect -4026 2842 -3980 2888
rect -3932 2842 -3886 2888
rect -3532 2842 -3486 2888
rect -3438 2842 -3392 2888
rect -3344 2842 -3298 2888
rect -3250 2842 -3204 2888
rect -3156 2842 -3110 2888
rect -3062 2842 -3016 2888
rect -2968 2842 -2922 2888
rect -2746 2842 -2700 2888
rect -2652 2842 -2606 2888
rect -2558 2842 -2512 2888
rect -2464 2842 -2418 2888
rect -2370 2842 -2324 2888
rect -2276 2842 -2230 2888
rect -2182 2842 -2136 2888
rect -1960 2842 -1914 2888
rect -1866 2842 -1820 2888
rect -1772 2842 -1726 2888
rect -1678 2842 -1632 2888
rect -1584 2842 -1538 2888
rect -1490 2842 -1444 2888
rect -1396 2842 -1350 2888
rect -1164 2842 -1118 2888
rect -1070 2842 -1024 2888
rect -976 2842 -930 2888
rect -4813 1132 -4767 1178
rect -4719 1132 -4673 1178
rect -4625 1132 -4579 1178
rect -4214 1132 -4168 1178
rect -4120 1132 -4074 1178
rect -4026 1132 -3980 1178
rect -3932 1132 -3886 1178
rect -3532 1132 -3486 1178
rect -3438 1132 -3392 1178
rect -3344 1132 -3298 1178
rect -3250 1132 -3204 1178
rect -3156 1132 -3110 1178
rect -3062 1132 -3016 1178
rect -2968 1132 -2922 1178
rect -2746 1132 -2700 1178
rect -2652 1132 -2606 1178
rect -2558 1132 -2512 1178
rect -2464 1132 -2418 1178
rect -2370 1132 -2324 1178
rect -2276 1132 -2230 1178
rect -2182 1132 -2136 1178
rect -1960 1132 -1914 1178
rect -1866 1132 -1820 1178
rect -1772 1132 -1726 1178
rect -1678 1132 -1632 1178
rect -1584 1132 -1538 1178
rect -1490 1132 -1444 1178
rect -1396 1132 -1350 1178
rect -1164 1132 -1118 1178
rect -1070 1132 -1024 1178
rect -976 1132 -930 1178
rect 106 33 152 79
rect 200 33 246 79
rect 294 33 340 79
rect 388 33 434 79
rect 482 33 528 79
rect 576 33 622 79
rect 670 33 716 79
rect 764 33 810 79
rect 858 33 904 79
rect 952 33 998 79
rect 1046 33 1092 79
rect 1140 33 1186 79
rect 1234 33 1280 79
rect 1328 33 1374 79
rect 1422 33 1468 79
rect 1516 33 1562 79
rect 1610 33 1656 79
rect 1704 33 1750 79
rect 1918 33 1964 79
rect 2012 33 2058 79
rect 2106 33 2152 79
rect 2200 33 2246 79
rect 2294 33 2340 79
rect 2388 33 2434 79
rect 2482 33 2528 79
rect 2576 33 2622 79
rect 2670 33 2716 79
rect 2764 33 2810 79
rect 2858 33 2904 79
rect 2952 33 2998 79
rect 3046 33 3092 79
rect 3140 33 3186 79
rect 3234 33 3280 79
rect 3328 33 3374 79
rect 3422 33 3468 79
rect 3516 33 3562 79
rect 3730 33 3776 79
rect 3824 33 3870 79
rect 3918 33 3964 79
rect 4012 33 4058 79
rect 4106 33 4152 79
rect 4200 33 4246 79
rect 4294 33 4340 79
rect 4388 33 4434 79
rect 4482 33 4528 79
rect 4576 33 4622 79
rect 4670 33 4716 79
rect 4764 33 4810 79
rect 4858 33 4904 79
rect 4952 33 4998 79
rect 5046 33 5092 79
rect 5140 33 5186 79
rect 5234 33 5280 79
rect 5328 33 5374 79
rect 5542 33 5588 79
rect 5636 33 5682 79
rect 5730 33 5776 79
rect 5824 33 5870 79
rect 5918 33 5964 79
rect 6012 33 6058 79
rect 6106 33 6152 79
rect 6200 33 6246 79
rect 6294 33 6340 79
rect 6388 33 6434 79
rect 6482 33 6528 79
rect 6576 33 6622 79
rect 6670 33 6716 79
rect 6764 33 6810 79
rect 6858 33 6904 79
rect 6952 33 6998 79
rect 7046 33 7092 79
rect 7140 33 7186 79
rect 7354 33 7400 79
rect 7448 33 7494 79
rect 7542 33 7588 79
rect 7636 33 7682 79
rect 7730 33 7776 79
rect 7824 33 7870 79
rect 7918 33 7964 79
rect 8012 33 8058 79
rect 8106 33 8152 79
rect 8200 33 8246 79
rect 8294 33 8340 79
rect 8388 33 8434 79
rect 8482 33 8528 79
rect 8576 33 8622 79
rect 8670 33 8716 79
rect 8764 33 8810 79
rect 8858 33 8904 79
rect 8952 33 8998 79
rect -4813 -578 -4767 -532
rect -4719 -578 -4673 -532
rect -4625 -578 -4579 -532
rect -4214 -578 -4168 -532
rect -4120 -578 -4074 -532
rect -4026 -578 -3980 -532
rect -3932 -578 -3886 -532
rect -3532 -578 -3486 -532
rect -3438 -578 -3392 -532
rect -3344 -578 -3298 -532
rect -3250 -578 -3204 -532
rect -3156 -578 -3110 -532
rect -3062 -578 -3016 -532
rect -2968 -578 -2922 -532
rect -2746 -578 -2700 -532
rect -2652 -578 -2606 -532
rect -2558 -578 -2512 -532
rect -2464 -578 -2418 -532
rect -2370 -578 -2324 -532
rect -2276 -578 -2230 -532
rect -2182 -578 -2136 -532
rect -1960 -578 -1914 -532
rect -1866 -578 -1820 -532
rect -1772 -578 -1726 -532
rect -1678 -578 -1632 -532
rect -1584 -578 -1538 -532
rect -1490 -578 -1444 -532
rect -1396 -578 -1350 -532
rect -1164 -578 -1118 -532
rect -1070 -578 -1024 -532
rect -976 -578 -930 -532
rect -4091 -7295 -4045 -7249
rect -3997 -7295 -3951 -7249
rect -3903 -7295 -3857 -7249
rect -3809 -7295 -3763 -7249
rect -3715 -7295 -3669 -7249
rect -3621 -7295 -3575 -7249
rect -3527 -7295 -3481 -7249
rect -3433 -7295 -3387 -7249
rect -3339 -7295 -3293 -7249
rect -3245 -7295 -3199 -7249
rect -3151 -7295 -3105 -7249
rect -3057 -7295 -3011 -7249
rect -2963 -7295 -2917 -7249
rect -2869 -7295 -2823 -7249
rect -2775 -7295 -2729 -7249
rect -2681 -7295 -2635 -7249
rect -2587 -7295 -2541 -7249
rect -2493 -7295 -2447 -7249
rect -2279 -7295 -2233 -7249
rect -2185 -7295 -2139 -7249
rect -2091 -7295 -2045 -7249
rect -1997 -7295 -1951 -7249
rect -1903 -7295 -1857 -7249
rect -1809 -7295 -1763 -7249
rect -1715 -7295 -1669 -7249
rect -1621 -7295 -1575 -7249
rect -1527 -7295 -1481 -7249
rect -1433 -7295 -1387 -7249
rect -1339 -7295 -1293 -7249
rect -1245 -7295 -1199 -7249
rect -1151 -7295 -1105 -7249
rect -1057 -7295 -1011 -7249
rect -963 -7295 -917 -7249
rect -869 -7295 -823 -7249
rect -775 -7295 -729 -7249
rect -681 -7295 -635 -7249
rect 106 -7295 152 -7249
rect 200 -7295 246 -7249
rect 294 -7295 340 -7249
rect 388 -7295 434 -7249
rect 482 -7295 528 -7249
rect 576 -7295 622 -7249
rect 670 -7295 716 -7249
rect 764 -7295 810 -7249
rect 858 -7295 904 -7249
rect 952 -7295 998 -7249
rect 1046 -7295 1092 -7249
rect 1140 -7295 1186 -7249
rect 1234 -7295 1280 -7249
rect 1328 -7295 1374 -7249
rect 1422 -7295 1468 -7249
rect 1516 -7295 1562 -7249
rect 1610 -7295 1656 -7249
rect 1704 -7295 1750 -7249
rect 1918 -7295 1964 -7249
rect 2012 -7295 2058 -7249
rect 2106 -7295 2152 -7249
rect 2200 -7295 2246 -7249
rect 2294 -7295 2340 -7249
rect 2388 -7295 2434 -7249
rect 2482 -7295 2528 -7249
rect 2576 -7295 2622 -7249
rect 2670 -7295 2716 -7249
rect 2764 -7295 2810 -7249
rect 2858 -7295 2904 -7249
rect 2952 -7295 2998 -7249
rect 3046 -7295 3092 -7249
rect 3140 -7295 3186 -7249
rect 3234 -7295 3280 -7249
rect 3328 -7295 3374 -7249
rect 3422 -7295 3468 -7249
rect 3516 -7295 3562 -7249
rect 3730 -7295 3776 -7249
rect 3824 -7295 3870 -7249
rect 3918 -7295 3964 -7249
rect 4012 -7295 4058 -7249
rect 4106 -7295 4152 -7249
rect 4200 -7295 4246 -7249
rect 4294 -7295 4340 -7249
rect 4388 -7295 4434 -7249
rect 4482 -7295 4528 -7249
rect 4576 -7295 4622 -7249
rect 4670 -7295 4716 -7249
rect 4764 -7295 4810 -7249
rect 4858 -7295 4904 -7249
rect 4952 -7295 4998 -7249
rect 5046 -7295 5092 -7249
rect 5140 -7295 5186 -7249
rect 5234 -7295 5280 -7249
rect 5328 -7295 5374 -7249
rect 5542 -7295 5588 -7249
rect 5636 -7295 5682 -7249
rect 5730 -7295 5776 -7249
rect 5824 -7295 5870 -7249
rect 5918 -7295 5964 -7249
rect 6012 -7295 6058 -7249
rect 6106 -7295 6152 -7249
rect 6200 -7295 6246 -7249
rect 6294 -7295 6340 -7249
rect 6388 -7295 6434 -7249
rect 6482 -7295 6528 -7249
rect 6576 -7295 6622 -7249
rect 6670 -7295 6716 -7249
rect 6764 -7295 6810 -7249
rect 6858 -7295 6904 -7249
rect 6952 -7295 6998 -7249
rect 7046 -7295 7092 -7249
rect 7140 -7295 7186 -7249
rect 7354 -7295 7400 -7249
rect 7448 -7295 7494 -7249
rect 7542 -7295 7588 -7249
rect 7636 -7295 7682 -7249
rect 7730 -7295 7776 -7249
rect 7824 -7295 7870 -7249
rect 7918 -7295 7964 -7249
rect 8012 -7295 8058 -7249
rect 8106 -7295 8152 -7249
rect 8200 -7295 8246 -7249
rect 8294 -7295 8340 -7249
rect 8388 -7295 8434 -7249
rect 8482 -7295 8528 -7249
rect 8576 -7295 8622 -7249
rect 8670 -7295 8716 -7249
rect 8764 -7295 8810 -7249
rect 8858 -7295 8904 -7249
rect 8952 -7295 8998 -7249
<< nsubdiffcont >>
rect -4860 3697 -4814 3743
rect -4766 3697 -4720 3743
rect -4672 3697 -4626 3743
rect -4578 3697 -4532 3743
rect -4449 3697 -4403 3743
rect -4355 3697 -4309 3743
rect -4261 3697 -4215 3743
rect -4167 3697 -4121 3743
rect -4073 3697 -4027 3743
rect -3979 3697 -3933 3743
rect -3885 3697 -3839 3743
rect -3791 3697 -3745 3743
rect -3697 3697 -3651 3743
rect -3569 3697 -3523 3743
rect -3475 3697 -3429 3743
rect -3381 3697 -3335 3743
rect -3287 3697 -3241 3743
rect -3193 3697 -3147 3743
rect -3099 3697 -3053 3743
rect -3005 3697 -2959 3743
rect -2911 3697 -2865 3743
rect -2783 3697 -2737 3743
rect -2689 3697 -2643 3743
rect -2595 3697 -2549 3743
rect -2501 3697 -2455 3743
rect -2407 3697 -2361 3743
rect -2313 3697 -2267 3743
rect -2219 3697 -2173 3743
rect -2125 3697 -2079 3743
rect -1997 3697 -1951 3743
rect -1903 3697 -1857 3743
rect -1809 3697 -1763 3743
rect -1715 3697 -1669 3743
rect -1621 3697 -1575 3743
rect -1527 3697 -1481 3743
rect -1433 3697 -1387 3743
rect -1339 3697 -1293 3743
rect -1211 3697 -1165 3743
rect -1117 3697 -1071 3743
rect -1023 3697 -977 3743
rect -929 3697 -883 3743
rect 59 3697 105 3743
rect 153 3697 199 3743
rect 247 3697 293 3743
rect 341 3697 387 3743
rect 435 3697 481 3743
rect 529 3697 575 3743
rect 623 3697 669 3743
rect 717 3697 763 3743
rect 811 3697 857 3743
rect 905 3697 951 3743
rect 999 3697 1045 3743
rect 1093 3697 1139 3743
rect 1187 3697 1233 3743
rect 1281 3697 1327 3743
rect 1375 3697 1421 3743
rect 1469 3697 1515 3743
rect 1563 3697 1609 3743
rect 1657 3697 1703 3743
rect 1751 3697 1797 3743
rect 1871 3697 1917 3743
rect 1965 3697 2011 3743
rect 2059 3697 2105 3743
rect 2153 3697 2199 3743
rect 2247 3697 2293 3743
rect 2341 3697 2387 3743
rect 2435 3697 2481 3743
rect 2529 3697 2575 3743
rect 2623 3697 2669 3743
rect 2717 3697 2763 3743
rect 2811 3697 2857 3743
rect 2905 3697 2951 3743
rect 2999 3697 3045 3743
rect 3093 3697 3139 3743
rect 3187 3697 3233 3743
rect 3281 3697 3327 3743
rect 3375 3697 3421 3743
rect 3469 3697 3515 3743
rect 3563 3697 3609 3743
rect 3683 3697 3729 3743
rect 3777 3697 3823 3743
rect 3871 3697 3917 3743
rect 3965 3697 4011 3743
rect 4059 3697 4105 3743
rect 4153 3697 4199 3743
rect 4247 3697 4293 3743
rect 4341 3697 4387 3743
rect 4435 3697 4481 3743
rect 4529 3697 4575 3743
rect 4623 3697 4669 3743
rect 4717 3697 4763 3743
rect 4811 3697 4857 3743
rect 4905 3697 4951 3743
rect 4999 3697 5045 3743
rect 5093 3697 5139 3743
rect 5187 3697 5233 3743
rect 5281 3697 5327 3743
rect 5375 3697 5421 3743
rect 5495 3697 5541 3743
rect 5589 3697 5635 3743
rect 5683 3697 5729 3743
rect 5777 3697 5823 3743
rect 5871 3697 5917 3743
rect 5965 3697 6011 3743
rect 6059 3697 6105 3743
rect 6153 3697 6199 3743
rect 6247 3697 6293 3743
rect 6341 3697 6387 3743
rect 6435 3697 6481 3743
rect 6529 3697 6575 3743
rect 6623 3697 6669 3743
rect 6717 3697 6763 3743
rect 6811 3697 6857 3743
rect 6905 3697 6951 3743
rect 6999 3697 7045 3743
rect 7093 3697 7139 3743
rect 7187 3697 7233 3743
rect 7307 3697 7353 3743
rect 7401 3697 7447 3743
rect 7495 3697 7541 3743
rect 7589 3697 7635 3743
rect 7683 3697 7729 3743
rect 7777 3697 7823 3743
rect 7871 3697 7917 3743
rect 7965 3697 8011 3743
rect 8059 3697 8105 3743
rect 8153 3697 8199 3743
rect 8247 3697 8293 3743
rect 8341 3697 8387 3743
rect 8435 3697 8481 3743
rect 8529 3697 8575 3743
rect 8623 3697 8669 3743
rect 8717 3697 8763 3743
rect 8811 3697 8857 3743
rect 8905 3697 8951 3743
rect 8999 3697 9045 3743
rect -4449 1987 -4403 2033
rect -4355 1987 -4309 2033
rect -4261 1987 -4215 2033
rect -4167 1987 -4121 2033
rect -4073 1987 -4027 2033
rect -3979 1987 -3933 2033
rect -3885 1987 -3839 2033
rect -3791 1987 -3745 2033
rect -3697 1987 -3651 2033
rect -3569 1987 -3523 2033
rect -3475 1987 -3429 2033
rect -3381 1987 -3335 2033
rect -3287 1987 -3241 2033
rect -3193 1987 -3147 2033
rect -3099 1987 -3053 2033
rect -3005 1987 -2959 2033
rect -2911 1987 -2865 2033
rect -2783 1987 -2737 2033
rect -2689 1987 -2643 2033
rect -2595 1987 -2549 2033
rect -2501 1987 -2455 2033
rect -2407 1987 -2361 2033
rect -2313 1987 -2267 2033
rect -2219 1987 -2173 2033
rect -2125 1987 -2079 2033
rect -1997 1987 -1951 2033
rect -1903 1987 -1857 2033
rect -1809 1987 -1763 2033
rect -1715 1987 -1669 2033
rect -1621 1987 -1575 2033
rect -1527 1987 -1481 2033
rect -1433 1987 -1387 2033
rect -1339 1987 -1293 2033
rect -1211 1987 -1165 2033
rect -1117 1987 -1071 2033
rect -1023 1987 -977 2033
rect -929 1987 -883 2033
rect -4860 277 -4814 323
rect -4766 277 -4720 323
rect -4672 277 -4626 323
rect -4578 277 -4532 323
rect -4449 277 -4403 323
rect -4355 277 -4309 323
rect -4261 277 -4215 323
rect -4167 277 -4121 323
rect -4073 277 -4027 323
rect -3979 277 -3933 323
rect -3885 277 -3839 323
rect -3791 277 -3745 323
rect -3697 277 -3651 323
rect -3569 277 -3523 323
rect -3475 277 -3429 323
rect -3381 277 -3335 323
rect -3287 277 -3241 323
rect -3193 277 -3147 323
rect -3099 277 -3053 323
rect -3005 277 -2959 323
rect -2911 277 -2865 323
rect -2783 277 -2737 323
rect -2689 277 -2643 323
rect -2595 277 -2549 323
rect -2501 277 -2455 323
rect -2407 277 -2361 323
rect -2313 277 -2267 323
rect -2219 277 -2173 323
rect -2125 277 -2079 323
rect -1997 277 -1951 323
rect -1903 277 -1857 323
rect -1809 277 -1763 323
rect -1715 277 -1669 323
rect -1621 277 -1575 323
rect -1527 277 -1481 323
rect -1433 277 -1387 323
rect -1339 277 -1293 323
rect -1211 277 -1165 323
rect -1117 277 -1071 323
rect -1023 277 -977 323
rect -929 277 -883 323
rect -4449 -1433 -4403 -1387
rect -4355 -1433 -4309 -1387
rect -4261 -1433 -4215 -1387
rect -4167 -1433 -4121 -1387
rect -4073 -1433 -4027 -1387
rect -3979 -1433 -3933 -1387
rect -3885 -1433 -3839 -1387
rect -3791 -1433 -3745 -1387
rect -3697 -1433 -3651 -1387
rect -3569 -1433 -3523 -1387
rect -3475 -1433 -3429 -1387
rect -3381 -1433 -3335 -1387
rect -3287 -1433 -3241 -1387
rect -3193 -1433 -3147 -1387
rect -3099 -1433 -3053 -1387
rect -3005 -1433 -2959 -1387
rect -2911 -1433 -2865 -1387
rect -2783 -1433 -2737 -1387
rect -2689 -1433 -2643 -1387
rect -2595 -1433 -2549 -1387
rect -2501 -1433 -2455 -1387
rect -2407 -1433 -2361 -1387
rect -2313 -1433 -2267 -1387
rect -2219 -1433 -2173 -1387
rect -2125 -1433 -2079 -1387
rect -1997 -1433 -1951 -1387
rect -1903 -1433 -1857 -1387
rect -1809 -1433 -1763 -1387
rect -1715 -1433 -1669 -1387
rect -1621 -1433 -1575 -1387
rect -1527 -1433 -1481 -1387
rect -1433 -1433 -1387 -1387
rect -1339 -1433 -1293 -1387
rect -1211 -1433 -1165 -1387
rect -1117 -1433 -1071 -1387
rect -1023 -1433 -977 -1387
rect -929 -1433 -883 -1387
rect -4138 -3631 -4092 -3585
rect -4044 -3631 -3998 -3585
rect -3950 -3631 -3904 -3585
rect -3856 -3631 -3810 -3585
rect -3762 -3631 -3716 -3585
rect -3668 -3631 -3622 -3585
rect -3574 -3631 -3528 -3585
rect -3480 -3631 -3434 -3585
rect -3386 -3631 -3340 -3585
rect -3292 -3631 -3246 -3585
rect -3198 -3631 -3152 -3585
rect -3104 -3631 -3058 -3585
rect -3010 -3631 -2964 -3585
rect -2916 -3631 -2870 -3585
rect -2822 -3631 -2776 -3585
rect -2728 -3631 -2682 -3585
rect -2634 -3631 -2588 -3585
rect -2540 -3631 -2494 -3585
rect -2446 -3631 -2400 -3585
rect -2326 -3631 -2280 -3585
rect -2232 -3631 -2186 -3585
rect -2138 -3631 -2092 -3585
rect -2044 -3631 -1998 -3585
rect -1950 -3631 -1904 -3585
rect -1856 -3631 -1810 -3585
rect -1762 -3631 -1716 -3585
rect -1668 -3631 -1622 -3585
rect -1574 -3631 -1528 -3585
rect -1480 -3631 -1434 -3585
rect -1386 -3631 -1340 -3585
rect -1292 -3631 -1246 -3585
rect -1198 -3631 -1152 -3585
rect -1104 -3631 -1058 -3585
rect -1010 -3631 -964 -3585
rect -916 -3631 -870 -3585
rect -822 -3631 -776 -3585
rect -728 -3631 -682 -3585
rect -634 -3631 -588 -3585
rect 59 -3631 105 -3585
rect 153 -3631 199 -3585
rect 247 -3631 293 -3585
rect 341 -3631 387 -3585
rect 435 -3631 481 -3585
rect 529 -3631 575 -3585
rect 623 -3631 669 -3585
rect 717 -3631 763 -3585
rect 811 -3631 857 -3585
rect 905 -3631 951 -3585
rect 999 -3631 1045 -3585
rect 1093 -3631 1139 -3585
rect 1187 -3631 1233 -3585
rect 1281 -3631 1327 -3585
rect 1375 -3631 1421 -3585
rect 1469 -3631 1515 -3585
rect 1563 -3631 1609 -3585
rect 1657 -3631 1703 -3585
rect 1751 -3631 1797 -3585
rect 1871 -3631 1917 -3585
rect 1965 -3631 2011 -3585
rect 2059 -3631 2105 -3585
rect 2153 -3631 2199 -3585
rect 2247 -3631 2293 -3585
rect 2341 -3631 2387 -3585
rect 2435 -3631 2481 -3585
rect 2529 -3631 2575 -3585
rect 2623 -3631 2669 -3585
rect 2717 -3631 2763 -3585
rect 2811 -3631 2857 -3585
rect 2905 -3631 2951 -3585
rect 2999 -3631 3045 -3585
rect 3093 -3631 3139 -3585
rect 3187 -3631 3233 -3585
rect 3281 -3631 3327 -3585
rect 3375 -3631 3421 -3585
rect 3469 -3631 3515 -3585
rect 3563 -3631 3609 -3585
rect 3683 -3631 3729 -3585
rect 3777 -3631 3823 -3585
rect 3871 -3631 3917 -3585
rect 3965 -3631 4011 -3585
rect 4059 -3631 4105 -3585
rect 4153 -3631 4199 -3585
rect 4247 -3631 4293 -3585
rect 4341 -3631 4387 -3585
rect 4435 -3631 4481 -3585
rect 4529 -3631 4575 -3585
rect 4623 -3631 4669 -3585
rect 4717 -3631 4763 -3585
rect 4811 -3631 4857 -3585
rect 4905 -3631 4951 -3585
rect 4999 -3631 5045 -3585
rect 5093 -3631 5139 -3585
rect 5187 -3631 5233 -3585
rect 5281 -3631 5327 -3585
rect 5375 -3631 5421 -3585
rect 5495 -3631 5541 -3585
rect 5589 -3631 5635 -3585
rect 5683 -3631 5729 -3585
rect 5777 -3631 5823 -3585
rect 5871 -3631 5917 -3585
rect 5965 -3631 6011 -3585
rect 6059 -3631 6105 -3585
rect 6153 -3631 6199 -3585
rect 6247 -3631 6293 -3585
rect 6341 -3631 6387 -3585
rect 6435 -3631 6481 -3585
rect 6529 -3631 6575 -3585
rect 6623 -3631 6669 -3585
rect 6717 -3631 6763 -3585
rect 6811 -3631 6857 -3585
rect 6905 -3631 6951 -3585
rect 6999 -3631 7045 -3585
rect 7093 -3631 7139 -3585
rect 7187 -3631 7233 -3585
rect 7307 -3631 7353 -3585
rect 7401 -3631 7447 -3585
rect 7495 -3631 7541 -3585
rect 7589 -3631 7635 -3585
rect 7683 -3631 7729 -3585
rect 7777 -3631 7823 -3585
rect 7871 -3631 7917 -3585
rect 7965 -3631 8011 -3585
rect 8059 -3631 8105 -3585
rect 8153 -3631 8199 -3585
rect 8247 -3631 8293 -3585
rect 8341 -3631 8387 -3585
rect 8435 -3631 8481 -3585
rect 8529 -3631 8575 -3585
rect 8623 -3631 8669 -3585
rect 8717 -3631 8763 -3585
rect 8811 -3631 8857 -3585
rect 8905 -3631 8951 -3585
rect 8999 -3631 9045 -3585
<< polysilicon >>
rect 196 7120 1660 7176
rect 196 7100 252 7120
rect 356 7100 412 7120
rect 516 7100 572 7120
rect 676 7100 732 7120
rect 836 7100 892 7120
rect 996 7100 1052 7120
rect 1156 7100 1212 7120
rect 1316 7100 1372 7120
rect 1604 7100 1660 7120
rect 2008 7120 3472 7176
rect 2008 7100 2064 7120
rect 2296 7100 2352 7120
rect 2456 7100 2512 7120
rect 2616 7100 2672 7120
rect 2776 7100 2832 7120
rect 2936 7100 2992 7120
rect 3096 7100 3152 7120
rect 3256 7100 3312 7120
rect 3416 7100 3472 7120
rect 3820 7120 5284 7176
rect 3820 7100 3876 7120
rect 4108 7100 4164 7120
rect 4268 7100 4324 7120
rect 4428 7100 4484 7120
rect 4588 7100 4644 7120
rect 4748 7100 4804 7120
rect 4908 7100 4964 7120
rect 5068 7100 5124 7120
rect 5228 7100 5284 7120
rect 5632 7120 7096 7176
rect 5632 7100 5688 7120
rect 5920 7100 5976 7120
rect 6080 7100 6136 7120
rect 6240 7100 6296 7120
rect 6400 7100 6456 7120
rect 6560 7100 6616 7120
rect 6720 7100 6776 7120
rect 6880 7100 6936 7120
rect 7040 7100 7096 7120
rect 7444 7120 8908 7176
rect 7444 7100 7500 7120
rect 7732 7100 7788 7120
rect 7892 7100 7948 7120
rect 8052 7100 8108 7120
rect 8212 7100 8268 7120
rect 8372 7100 8428 7120
rect 8532 7100 8588 7120
rect 8692 7100 8748 7120
rect 8852 7100 8908 7120
rect 196 6714 252 6850
rect 356 6714 412 6850
rect 516 6714 572 6850
rect 676 6714 732 6850
rect 836 6714 892 6850
rect 996 6714 1052 6850
rect 1156 6714 1212 6850
rect 1316 6714 1372 6850
rect 1604 6714 1660 6850
rect 2008 6714 2064 6850
rect 2296 6714 2352 6850
rect 2456 6714 2512 6850
rect 2616 6714 2672 6850
rect 2776 6714 2832 6850
rect 2936 6714 2992 6850
rect 3096 6714 3152 6850
rect 3256 6714 3312 6850
rect 3416 6714 3472 6850
rect 3820 6714 3876 6850
rect 4108 6714 4164 6850
rect 4268 6714 4324 6850
rect 4428 6714 4484 6850
rect 4588 6714 4644 6850
rect 4748 6714 4804 6850
rect 4908 6714 4964 6850
rect 5068 6714 5124 6850
rect 5228 6714 5284 6850
rect 5632 6714 5688 6850
rect 5920 6714 5976 6850
rect 6080 6714 6136 6850
rect 6240 6714 6296 6850
rect 6400 6714 6456 6850
rect 6560 6714 6616 6850
rect 6720 6714 6776 6850
rect 6880 6714 6936 6850
rect 7040 6714 7096 6850
rect 7444 6714 7500 6850
rect 7732 6714 7788 6850
rect 7892 6714 7948 6850
rect 8052 6714 8108 6850
rect 8212 6714 8268 6850
rect 8372 6714 8428 6850
rect 8532 6714 8588 6850
rect 8692 6714 8748 6850
rect 8852 6714 8908 6850
rect 196 6328 252 6464
rect 356 6328 412 6464
rect 516 6328 572 6464
rect 676 6328 732 6464
rect 836 6328 892 6464
rect 996 6328 1052 6464
rect 1156 6328 1212 6464
rect 1316 6328 1372 6464
rect 1604 6328 1660 6464
rect 2008 6328 2064 6464
rect 2296 6328 2352 6464
rect 2456 6328 2512 6464
rect 2616 6328 2672 6464
rect 2776 6328 2832 6464
rect 2936 6328 2992 6464
rect 3096 6328 3152 6464
rect 3256 6328 3312 6464
rect 3416 6328 3472 6464
rect 3820 6328 3876 6464
rect 4108 6328 4164 6464
rect 4268 6328 4324 6464
rect 4428 6328 4484 6464
rect 4588 6328 4644 6464
rect 4748 6328 4804 6464
rect 4908 6328 4964 6464
rect 5068 6328 5124 6464
rect 5228 6328 5284 6464
rect 5632 6328 5688 6464
rect 5920 6328 5976 6464
rect 6080 6328 6136 6464
rect 6240 6328 6296 6464
rect 6400 6328 6456 6464
rect 6560 6328 6616 6464
rect 6720 6328 6776 6464
rect 6880 6328 6936 6464
rect 7040 6328 7096 6464
rect 7444 6328 7500 6464
rect 7732 6328 7788 6464
rect 7892 6328 7948 6464
rect 8052 6328 8108 6464
rect 8212 6328 8268 6464
rect 8372 6328 8428 6464
rect 8532 6328 8588 6464
rect 8692 6328 8748 6464
rect 8852 6328 8908 6464
rect 196 6034 252 6078
rect 356 6034 412 6078
rect 516 6034 572 6078
rect 676 6034 732 6078
rect 836 6034 892 6078
rect 996 6034 1052 6078
rect 1156 6034 1212 6078
rect 1316 6034 1372 6078
rect 1604 5964 1660 6078
rect 1708 5964 1780 5972
rect 1484 5954 1556 5962
rect 1316 5949 1556 5954
rect 1316 5903 1497 5949
rect 1543 5903 1556 5949
rect 1316 5898 1556 5903
rect 196 5776 252 5820
rect 356 5776 412 5820
rect 516 5776 572 5820
rect 676 5776 732 5820
rect 836 5776 892 5820
rect 996 5776 1052 5820
rect 1156 5776 1212 5820
rect 1316 5776 1372 5898
rect 1484 5890 1556 5898
rect 1604 5959 1780 5964
rect 1604 5913 1721 5959
rect 1767 5913 1780 5959
rect 1604 5908 1780 5913
rect 1604 5776 1660 5908
rect 1708 5900 1780 5908
rect 1888 5964 1960 5972
rect 2008 5964 2064 6078
rect 2296 6034 2352 6078
rect 2456 6034 2512 6078
rect 2616 6034 2672 6078
rect 2776 6034 2832 6078
rect 2936 6034 2992 6078
rect 3096 6034 3152 6078
rect 3256 6034 3312 6078
rect 3416 6034 3472 6078
rect 1888 5959 2064 5964
rect 3700 5964 3772 5972
rect 3820 5964 3876 6078
rect 4108 6034 4164 6078
rect 4268 6034 4324 6078
rect 4428 6034 4484 6078
rect 4588 6034 4644 6078
rect 4748 6034 4804 6078
rect 4908 6034 4964 6078
rect 5068 6034 5124 6078
rect 5228 6034 5284 6078
rect 1888 5913 1901 5959
rect 1947 5913 2064 5959
rect 1888 5908 2064 5913
rect 1888 5900 1960 5908
rect 2008 5776 2064 5908
rect 2112 5954 2184 5962
rect 3700 5959 3876 5964
rect 5512 5964 5584 5972
rect 5632 5964 5688 6078
rect 5920 6034 5976 6078
rect 6080 6034 6136 6078
rect 6240 6034 6296 6078
rect 6400 6034 6456 6078
rect 6560 6034 6616 6078
rect 6720 6034 6776 6078
rect 6880 6034 6936 6078
rect 7040 6034 7096 6078
rect 2112 5949 2352 5954
rect 2112 5903 2125 5949
rect 2171 5903 2352 5949
rect 2112 5898 2352 5903
rect 3700 5913 3713 5959
rect 3759 5913 3876 5959
rect 3700 5908 3876 5913
rect 3700 5900 3772 5908
rect 2112 5890 2184 5898
rect 2296 5776 2352 5898
rect 2456 5776 2512 5820
rect 2616 5776 2672 5820
rect 2776 5776 2832 5820
rect 2936 5776 2992 5820
rect 3096 5776 3152 5820
rect 3256 5776 3312 5820
rect 3416 5776 3472 5820
rect 3820 5776 3876 5908
rect 3924 5954 3996 5962
rect 5512 5959 5688 5964
rect 7324 5964 7396 5972
rect 7444 5964 7500 6078
rect 7732 6034 7788 6078
rect 7892 6034 7948 6078
rect 8052 6034 8108 6078
rect 8212 6034 8268 6078
rect 8372 6034 8428 6078
rect 8532 6034 8588 6078
rect 8692 6034 8748 6078
rect 8852 6034 8908 6078
rect 3924 5949 4164 5954
rect 3924 5903 3937 5949
rect 3983 5903 4164 5949
rect 3924 5898 4164 5903
rect 5512 5913 5525 5959
rect 5571 5913 5688 5959
rect 5512 5908 5688 5913
rect 5512 5900 5584 5908
rect 3924 5890 3996 5898
rect 4108 5776 4164 5898
rect 4268 5776 4324 5820
rect 4428 5776 4484 5820
rect 4588 5776 4644 5820
rect 4748 5776 4804 5820
rect 4908 5776 4964 5820
rect 5068 5776 5124 5820
rect 5228 5776 5284 5820
rect 5632 5776 5688 5908
rect 5736 5954 5808 5962
rect 7324 5959 7500 5964
rect 5736 5949 5976 5954
rect 5736 5903 5749 5949
rect 5795 5903 5976 5949
rect 5736 5898 5976 5903
rect 7324 5913 7337 5959
rect 7383 5913 7500 5959
rect 7324 5908 7500 5913
rect 7324 5900 7396 5908
rect 5736 5890 5808 5898
rect 5920 5776 5976 5898
rect 6080 5776 6136 5820
rect 6240 5776 6296 5820
rect 6400 5776 6456 5820
rect 6560 5776 6616 5820
rect 6720 5776 6776 5820
rect 6880 5776 6936 5820
rect 7040 5776 7096 5820
rect 7444 5776 7500 5908
rect 7548 5954 7620 5962
rect 7548 5949 7788 5954
rect 7548 5903 7561 5949
rect 7607 5903 7788 5949
rect 7548 5898 7788 5903
rect 7548 5890 7620 5898
rect 7732 5776 7788 5898
rect 7892 5776 7948 5820
rect 8052 5776 8108 5820
rect 8212 5776 8268 5820
rect 8372 5776 8428 5820
rect 8532 5776 8588 5820
rect 8692 5776 8748 5820
rect 8852 5776 8908 5820
rect 196 5140 252 5276
rect 356 5140 412 5276
rect 516 5140 572 5276
rect 676 5140 732 5276
rect 836 5140 892 5276
rect 996 5140 1052 5276
rect 1156 5140 1212 5276
rect 1316 5140 1372 5276
rect 1604 5140 1660 5276
rect 2008 5140 2064 5276
rect 2296 5140 2352 5276
rect 2456 5140 2512 5276
rect 2616 5140 2672 5276
rect 2776 5140 2832 5276
rect 2936 5140 2992 5276
rect 3096 5140 3152 5276
rect 3256 5140 3312 5276
rect 3416 5140 3472 5276
rect 3820 5140 3876 5276
rect 4108 5140 4164 5276
rect 4268 5140 4324 5276
rect 4428 5140 4484 5276
rect 4588 5140 4644 5276
rect 4748 5140 4804 5276
rect 4908 5140 4964 5276
rect 5068 5140 5124 5276
rect 5228 5140 5284 5276
rect 5632 5140 5688 5276
rect 5920 5140 5976 5276
rect 6080 5140 6136 5276
rect 6240 5140 6296 5276
rect 6400 5140 6456 5276
rect 6560 5140 6616 5276
rect 6720 5140 6776 5276
rect 6880 5140 6936 5276
rect 7040 5140 7096 5276
rect 7444 5140 7500 5276
rect 7732 5140 7788 5276
rect 7892 5140 7948 5276
rect 8052 5140 8108 5276
rect 8212 5140 8268 5276
rect 8372 5140 8428 5276
rect 8532 5140 8588 5276
rect 8692 5140 8748 5276
rect 8852 5140 8908 5276
rect 196 4504 252 4640
rect 356 4504 412 4640
rect 516 4504 572 4640
rect 676 4504 732 4640
rect 836 4504 892 4640
rect 996 4504 1052 4640
rect 1156 4504 1212 4640
rect 1316 4504 1372 4640
rect 1604 4504 1660 4640
rect 2008 4504 2064 4640
rect 2296 4504 2352 4640
rect 2456 4504 2512 4640
rect 2616 4504 2672 4640
rect 2776 4504 2832 4640
rect 2936 4504 2992 4640
rect 3096 4504 3152 4640
rect 3256 4504 3312 4640
rect 3416 4504 3472 4640
rect 3820 4504 3876 4640
rect 4108 4504 4164 4640
rect 4268 4504 4324 4640
rect 4428 4504 4484 4640
rect 4588 4504 4644 4640
rect 4748 4504 4804 4640
rect 4908 4504 4964 4640
rect 5068 4504 5124 4640
rect 5228 4504 5284 4640
rect 5632 4504 5688 4640
rect 5920 4504 5976 4640
rect 6080 4504 6136 4640
rect 6240 4504 6296 4640
rect 6400 4504 6456 4640
rect 6560 4504 6616 4640
rect 6720 4504 6776 4640
rect 6880 4504 6936 4640
rect 7040 4504 7096 4640
rect 7444 4504 7500 4640
rect 7732 4504 7788 4640
rect 7892 4504 7948 4640
rect 8052 4504 8108 4640
rect 8212 4504 8268 4640
rect 8372 4504 8428 4640
rect 8532 4504 8588 4640
rect 8692 4504 8748 4640
rect 8852 4504 8908 4640
rect 196 3984 252 4004
rect 356 3984 412 4004
rect 516 3984 572 4004
rect 676 3984 732 4004
rect 836 3984 892 4004
rect 996 3984 1052 4004
rect 1156 3984 1212 4004
rect 1316 3984 1372 4004
rect 196 3928 1372 3984
rect 1604 3960 1660 4004
rect 2008 3960 2064 4004
rect 2296 3984 2352 4004
rect 2456 3984 2512 4004
rect 2616 3984 2672 4004
rect 2776 3984 2832 4004
rect 2936 3984 2992 4004
rect 3096 3984 3152 4004
rect 3256 3984 3312 4004
rect 3416 3984 3472 4004
rect 2296 3928 3472 3984
rect 3820 3960 3876 4004
rect 4108 3984 4164 4004
rect 4268 3984 4324 4004
rect 4428 3984 4484 4004
rect 4588 3984 4644 4004
rect 4748 3984 4804 4004
rect 4908 3984 4964 4004
rect 5068 3984 5124 4004
rect 5228 3984 5284 4004
rect 4108 3928 5284 3984
rect 5632 3960 5688 4004
rect 5920 3984 5976 4004
rect 6080 3984 6136 4004
rect 6240 3984 6296 4004
rect 6400 3984 6456 4004
rect 6560 3984 6616 4004
rect 6720 3984 6776 4004
rect 6880 3984 6936 4004
rect 7040 3984 7096 4004
rect 5920 3928 7096 3984
rect 7444 3960 7500 4004
rect 7732 3984 7788 4004
rect 7892 3984 7948 4004
rect 8052 3984 8108 4004
rect 8212 3984 8268 4004
rect 8372 3984 8428 4004
rect 8532 3984 8588 4004
rect 8692 3984 8748 4004
rect 8852 3984 8908 4004
rect 7732 3928 8908 3984
rect -4724 3573 -4668 3617
rect -4318 3528 -4262 3572
rect -4158 3528 -4102 3572
rect -3998 3528 -3942 3572
rect -3838 3528 -3782 3572
rect -3445 3539 -2997 3583
rect -2659 3539 -2211 3583
rect -1873 3539 -1425 3583
rect -1075 3573 -1019 3617
rect -4844 3207 -4772 3215
rect -4724 3207 -4668 3373
rect -3445 3407 -2997 3451
rect -2659 3407 -2211 3451
rect -1873 3407 -1425 3451
rect -4844 3202 -4668 3207
rect -4844 3156 -4831 3202
rect -4785 3156 -4668 3202
rect -4318 3189 -4262 3328
rect -4844 3151 -4668 3156
rect -4844 3143 -4772 3151
rect -4724 3101 -4668 3151
rect -4337 3181 -4262 3189
rect -4158 3181 -4102 3328
rect -4337 3176 -4102 3181
rect -4337 3130 -4324 3176
rect -4278 3130 -4102 3176
rect -4337 3125 -4102 3130
rect -4337 3117 -4265 3125
rect -4158 3089 -4102 3125
rect -3998 3264 -3942 3328
rect -3838 3264 -3782 3328
rect -3378 3289 -3306 3297
rect -3258 3289 -3146 3407
rect -3378 3284 -3146 3289
rect -3998 3208 -3778 3264
rect -3378 3238 -3365 3284
rect -3319 3238 -3146 3284
rect -3378 3233 -3146 3238
rect -3378 3225 -3306 3233
rect -3998 3089 -3942 3208
rect -3834 3151 -3778 3208
rect -3730 3151 -3658 3159
rect -3834 3146 -3658 3151
rect -3834 3099 -3717 3146
rect -3671 3099 -3658 3146
rect -3834 3095 -3658 3099
rect -4724 2957 -4668 3001
rect -3730 3086 -3658 3095
rect -3258 3079 -3146 3233
rect -2592 3289 -2520 3297
rect -2472 3289 -2360 3407
rect -2592 3284 -2360 3289
rect -2592 3238 -2579 3284
rect -2533 3238 -2360 3284
rect -2592 3233 -2360 3238
rect -2592 3225 -2520 3233
rect -2472 3079 -2360 3233
rect -1806 3289 -1734 3297
rect -1686 3289 -1574 3407
rect 196 3436 252 3480
rect 484 3456 1660 3512
rect 484 3436 540 3456
rect 644 3436 700 3456
rect 804 3436 860 3456
rect 964 3436 1020 3456
rect 1124 3436 1180 3456
rect 1284 3436 1340 3456
rect 1444 3436 1500 3456
rect 1604 3436 1660 3456
rect 2008 3456 3184 3512
rect 2008 3436 2064 3456
rect 2168 3436 2224 3456
rect 2328 3436 2384 3456
rect 2488 3436 2544 3456
rect 2648 3436 2704 3456
rect 2808 3436 2864 3456
rect 2968 3436 3024 3456
rect 3128 3436 3184 3456
rect 3416 3436 3472 3480
rect 3820 3436 3876 3480
rect 4108 3456 5284 3512
rect 4108 3436 4164 3456
rect 4268 3436 4324 3456
rect 4428 3436 4484 3456
rect 4588 3436 4644 3456
rect 4748 3436 4804 3456
rect 4908 3436 4964 3456
rect 5068 3436 5124 3456
rect 5228 3436 5284 3456
rect 5632 3456 6808 3512
rect 5632 3436 5688 3456
rect 5792 3436 5848 3456
rect 5952 3436 6008 3456
rect 6112 3436 6168 3456
rect 6272 3436 6328 3456
rect 6432 3436 6488 3456
rect 6592 3436 6648 3456
rect 6752 3436 6808 3456
rect 7040 3436 7096 3480
rect 7444 3456 8620 3512
rect 7444 3436 7500 3456
rect 7604 3436 7660 3456
rect 7764 3436 7820 3456
rect 7924 3436 7980 3456
rect 8084 3436 8140 3456
rect 8244 3436 8300 3456
rect 8404 3436 8460 3456
rect 8564 3436 8620 3456
rect 8852 3436 8908 3480
rect -1806 3284 -1574 3289
rect -1806 3238 -1793 3284
rect -1747 3238 -1574 3284
rect -1806 3233 -1574 3238
rect -1806 3225 -1734 3233
rect -1686 3079 -1574 3233
rect -1195 3207 -1123 3215
rect -1075 3207 -1019 3373
rect -1195 3202 -1019 3207
rect -1195 3156 -1182 3202
rect -1136 3156 -1019 3202
rect -1195 3151 -1019 3156
rect -1195 3143 -1123 3151
rect -1075 3101 -1019 3151
rect -3449 3035 -3001 3079
rect -4158 2945 -4102 2989
rect -3998 2945 -3942 2989
rect -3449 2947 -3001 2991
rect -2663 3035 -2215 3079
rect -2663 2947 -2215 2991
rect -1877 3035 -1429 3079
rect -1877 2947 -1429 2991
rect -1075 2957 -1019 3001
rect 196 2800 252 2936
rect 484 2800 540 2936
rect 644 2800 700 2936
rect 804 2800 860 2936
rect 964 2800 1020 2936
rect 1124 2800 1180 2936
rect 1284 2800 1340 2936
rect 1444 2800 1500 2936
rect 1604 2800 1660 2936
rect 2008 2800 2064 2936
rect 2168 2800 2224 2936
rect 2328 2800 2384 2936
rect 2488 2800 2544 2936
rect 2648 2800 2704 2936
rect 2808 2800 2864 2936
rect 2968 2800 3024 2936
rect 3128 2800 3184 2936
rect 3416 2800 3472 2936
rect 3820 2800 3876 2936
rect 4108 2800 4164 2936
rect 4268 2800 4324 2936
rect 4428 2800 4484 2936
rect 4588 2800 4644 2936
rect 4748 2800 4804 2936
rect 4908 2800 4964 2936
rect 5068 2800 5124 2936
rect 5228 2800 5284 2936
rect 5632 2800 5688 2936
rect 5792 2800 5848 2936
rect 5952 2800 6008 2936
rect 6112 2800 6168 2936
rect 6272 2800 6328 2936
rect 6432 2800 6488 2936
rect 6592 2800 6648 2936
rect 6752 2800 6808 2936
rect 7040 2800 7096 2936
rect 7444 2800 7500 2936
rect 7604 2800 7660 2936
rect 7764 2800 7820 2936
rect 7924 2800 7980 2936
rect 8084 2800 8140 2936
rect 8244 2800 8300 2936
rect 8404 2800 8460 2936
rect 8564 2800 8620 2936
rect 8852 2800 8908 2936
rect -4158 2741 -4102 2785
rect -3998 2741 -3942 2785
rect -3449 2739 -3001 2783
rect -3449 2651 -3001 2695
rect -2663 2739 -2215 2783
rect -2663 2651 -2215 2695
rect -1877 2739 -1429 2783
rect -1877 2651 -1429 2695
rect -1075 2729 -1019 2773
rect -4337 2605 -4265 2613
rect -4158 2605 -4102 2641
rect -4337 2600 -4102 2605
rect -4337 2554 -4324 2600
rect -4278 2554 -4102 2600
rect -4337 2549 -4102 2554
rect -4337 2541 -4262 2549
rect -4318 2402 -4262 2541
rect -4158 2402 -4102 2549
rect -3998 2522 -3942 2641
rect -3730 2635 -3658 2644
rect -3834 2631 -3658 2635
rect -3834 2584 -3717 2631
rect -3671 2584 -3658 2631
rect -3834 2579 -3658 2584
rect -3834 2522 -3778 2579
rect -3730 2571 -3658 2579
rect -3998 2466 -3778 2522
rect -3378 2497 -3306 2505
rect -3258 2497 -3146 2651
rect -3378 2492 -3146 2497
rect -3998 2402 -3942 2466
rect -3838 2402 -3782 2466
rect -3378 2446 -3365 2492
rect -3319 2446 -3146 2492
rect -3378 2441 -3146 2446
rect -3378 2433 -3306 2441
rect -3258 2323 -3146 2441
rect -2592 2497 -2520 2505
rect -2472 2497 -2360 2651
rect -2592 2492 -2360 2497
rect -2592 2446 -2579 2492
rect -2533 2446 -2360 2492
rect -2592 2441 -2360 2446
rect -2592 2433 -2520 2441
rect -2472 2323 -2360 2441
rect -1806 2497 -1734 2505
rect -1686 2497 -1574 2651
rect -1195 2579 -1123 2587
rect -1075 2579 -1019 2629
rect -1195 2574 -1019 2579
rect -1195 2528 -1182 2574
rect -1136 2528 -1019 2574
rect -1195 2523 -1019 2528
rect -1195 2515 -1123 2523
rect -1806 2492 -1574 2497
rect -1806 2446 -1793 2492
rect -1747 2446 -1574 2492
rect -1806 2441 -1574 2446
rect -1806 2433 -1734 2441
rect -1686 2323 -1574 2441
rect -1075 2357 -1019 2523
rect -3445 2279 -2997 2323
rect -2659 2279 -2211 2323
rect -1873 2279 -1425 2323
rect -4318 2158 -4262 2202
rect -4158 2158 -4102 2202
rect -3998 2158 -3942 2202
rect -3838 2158 -3782 2202
rect -3445 2147 -2997 2191
rect -2659 2147 -2211 2191
rect -1873 2147 -1425 2191
rect 196 2164 252 2300
rect 484 2164 540 2300
rect 644 2164 700 2300
rect 804 2164 860 2300
rect 964 2164 1020 2300
rect 1124 2164 1180 2300
rect 1284 2164 1340 2300
rect 1444 2164 1500 2300
rect 1604 2164 1660 2300
rect 2008 2164 2064 2300
rect 2168 2164 2224 2300
rect 2328 2164 2384 2300
rect 2488 2164 2544 2300
rect 2648 2164 2704 2300
rect 2808 2164 2864 2300
rect 2968 2164 3024 2300
rect 3128 2164 3184 2300
rect 3416 2164 3472 2300
rect 3820 2164 3876 2300
rect 4108 2164 4164 2300
rect 4268 2164 4324 2300
rect 4428 2164 4484 2300
rect 4588 2164 4644 2300
rect 4748 2164 4804 2300
rect 4908 2164 4964 2300
rect 5068 2164 5124 2300
rect 5228 2164 5284 2300
rect 5632 2164 5688 2300
rect 5792 2164 5848 2300
rect 5952 2164 6008 2300
rect 6112 2164 6168 2300
rect 6272 2164 6328 2300
rect 6432 2164 6488 2300
rect 6592 2164 6648 2300
rect 6752 2164 6808 2300
rect 7040 2164 7096 2300
rect 7444 2164 7500 2300
rect 7604 2164 7660 2300
rect 7764 2164 7820 2300
rect 7924 2164 7980 2300
rect 8084 2164 8140 2300
rect 8244 2164 8300 2300
rect 8404 2164 8460 2300
rect 8564 2164 8620 2300
rect 8852 2164 8908 2300
rect -1075 2113 -1019 2157
rect -4318 1818 -4262 1862
rect -4158 1818 -4102 1862
rect -3998 1818 -3942 1862
rect -3838 1818 -3782 1862
rect -3445 1829 -2997 1873
rect -2659 1829 -2211 1873
rect -1873 1829 -1425 1873
rect -1075 1863 -1019 1907
rect -3445 1697 -2997 1741
rect -2659 1697 -2211 1741
rect -1873 1697 -1425 1741
rect -4318 1479 -4262 1618
rect -4337 1471 -4262 1479
rect -4158 1471 -4102 1618
rect -4337 1466 -4102 1471
rect -4337 1420 -4324 1466
rect -4278 1420 -4102 1466
rect -4337 1415 -4102 1420
rect -4337 1407 -4265 1415
rect -4158 1379 -4102 1415
rect -3998 1554 -3942 1618
rect -3838 1554 -3782 1618
rect -3378 1579 -3306 1587
rect -3258 1579 -3146 1697
rect -3378 1574 -3146 1579
rect -3998 1498 -3778 1554
rect -3378 1528 -3365 1574
rect -3319 1528 -3146 1574
rect -3378 1523 -3146 1528
rect -3378 1515 -3306 1523
rect -3998 1379 -3942 1498
rect -3834 1441 -3778 1498
rect -3730 1441 -3658 1449
rect -3834 1436 -3658 1441
rect -3834 1389 -3717 1436
rect -3671 1389 -3658 1436
rect -3834 1385 -3658 1389
rect -3730 1376 -3658 1385
rect -3258 1369 -3146 1523
rect -2592 1579 -2520 1587
rect -2472 1579 -2360 1697
rect -2592 1574 -2360 1579
rect -2592 1528 -2579 1574
rect -2533 1528 -2360 1574
rect -2592 1523 -2360 1528
rect -2592 1515 -2520 1523
rect -2472 1369 -2360 1523
rect -1806 1579 -1734 1587
rect -1686 1579 -1574 1697
rect -1806 1574 -1574 1579
rect -1806 1528 -1793 1574
rect -1747 1528 -1574 1574
rect -1806 1523 -1574 1528
rect -1806 1515 -1734 1523
rect -1686 1369 -1574 1523
rect -1195 1497 -1123 1505
rect -1075 1497 -1019 1663
rect -1195 1492 -1019 1497
rect -1195 1446 -1182 1492
rect -1136 1446 -1019 1492
rect 76 1532 148 1540
rect 196 1532 252 1664
rect 76 1527 252 1532
rect 76 1481 89 1527
rect 135 1481 252 1527
rect 76 1476 252 1481
rect 300 1542 372 1550
rect 484 1542 540 1664
rect 644 1620 700 1664
rect 804 1620 860 1664
rect 964 1620 1020 1664
rect 1124 1620 1180 1664
rect 1284 1620 1340 1664
rect 1444 1620 1500 1664
rect 1604 1620 1660 1664
rect 2008 1620 2064 1664
rect 2168 1620 2224 1664
rect 2328 1620 2384 1664
rect 2488 1620 2544 1664
rect 2648 1620 2704 1664
rect 2808 1620 2864 1664
rect 2968 1620 3024 1664
rect 300 1537 540 1542
rect 300 1491 313 1537
rect 359 1491 540 1537
rect 300 1486 540 1491
rect 3128 1542 3184 1664
rect 3296 1542 3368 1550
rect 3128 1537 3368 1542
rect 3128 1491 3309 1537
rect 3355 1491 3368 1537
rect 3128 1486 3368 1491
rect 300 1478 372 1486
rect 3296 1478 3368 1486
rect 3416 1532 3472 1664
rect 3520 1532 3592 1540
rect 3416 1527 3592 1532
rect 3416 1481 3533 1527
rect 3579 1481 3592 1527
rect 76 1468 148 1476
rect -1195 1441 -1019 1446
rect -1195 1433 -1123 1441
rect -1075 1391 -1019 1441
rect -3449 1325 -3001 1369
rect -4158 1235 -4102 1279
rect -3998 1235 -3942 1279
rect -3449 1237 -3001 1281
rect -2663 1325 -2215 1369
rect -2663 1237 -2215 1281
rect -1877 1325 -1429 1369
rect -1877 1237 -1429 1281
rect 196 1362 252 1476
rect 3416 1476 3592 1481
rect 484 1362 540 1406
rect 644 1362 700 1406
rect 804 1362 860 1406
rect 964 1362 1020 1406
rect 1124 1362 1180 1406
rect 1284 1362 1340 1406
rect 1444 1362 1500 1406
rect 1604 1362 1660 1406
rect 2008 1362 2064 1406
rect 2168 1362 2224 1406
rect 2328 1362 2384 1406
rect 2488 1362 2544 1406
rect 2648 1362 2704 1406
rect 2808 1362 2864 1406
rect 2968 1362 3024 1406
rect 3128 1362 3184 1406
rect 3416 1362 3472 1476
rect 3520 1468 3592 1476
rect 3700 1532 3772 1540
rect 3820 1532 3876 1664
rect 3700 1527 3876 1532
rect 3700 1481 3713 1527
rect 3759 1481 3876 1527
rect 3700 1476 3876 1481
rect 3924 1542 3996 1550
rect 4108 1542 4164 1664
rect 4268 1620 4324 1664
rect 4428 1620 4484 1664
rect 4588 1620 4644 1664
rect 4748 1620 4804 1664
rect 4908 1620 4964 1664
rect 5068 1620 5124 1664
rect 5228 1620 5284 1664
rect 5632 1620 5688 1664
rect 5792 1620 5848 1664
rect 5952 1620 6008 1664
rect 6112 1620 6168 1664
rect 6272 1620 6328 1664
rect 6432 1620 6488 1664
rect 6592 1620 6648 1664
rect 3924 1537 4164 1542
rect 3924 1491 3937 1537
rect 3983 1491 4164 1537
rect 3924 1486 4164 1491
rect 6752 1542 6808 1664
rect 6920 1542 6992 1550
rect 6752 1537 6992 1542
rect 6752 1491 6933 1537
rect 6979 1491 6992 1537
rect 6752 1486 6992 1491
rect 3924 1478 3996 1486
rect 6920 1478 6992 1486
rect 7040 1532 7096 1664
rect 7444 1620 7500 1664
rect 7604 1620 7660 1664
rect 7764 1620 7820 1664
rect 7924 1620 7980 1664
rect 8084 1620 8140 1664
rect 8244 1620 8300 1664
rect 8404 1620 8460 1664
rect 8564 1542 8620 1664
rect 8732 1542 8804 1550
rect 7144 1532 7216 1540
rect 7040 1527 7216 1532
rect 7040 1481 7157 1527
rect 7203 1481 7216 1527
rect 8564 1537 8804 1542
rect 8564 1491 8745 1537
rect 8791 1491 8804 1537
rect 8564 1486 8804 1491
rect 3700 1468 3772 1476
rect 3820 1362 3876 1476
rect 7040 1476 7216 1481
rect 8732 1478 8804 1486
rect 8852 1532 8908 1664
rect 8956 1532 9028 1540
rect 8852 1527 9028 1532
rect 8852 1481 8969 1527
rect 9015 1481 9028 1527
rect 4108 1362 4164 1406
rect 4268 1362 4324 1406
rect 4428 1362 4484 1406
rect 4588 1362 4644 1406
rect 4748 1362 4804 1406
rect 4908 1362 4964 1406
rect 5068 1362 5124 1406
rect 5228 1362 5284 1406
rect 5632 1362 5688 1406
rect 5792 1362 5848 1406
rect 5952 1362 6008 1406
rect 6112 1362 6168 1406
rect 6272 1362 6328 1406
rect 6432 1362 6488 1406
rect 6592 1362 6648 1406
rect 6752 1362 6808 1406
rect 7040 1362 7096 1476
rect 7144 1468 7216 1476
rect 8852 1476 9028 1481
rect 7444 1362 7500 1406
rect 7604 1362 7660 1406
rect 7764 1362 7820 1406
rect 7924 1362 7980 1406
rect 8084 1362 8140 1406
rect 8244 1362 8300 1406
rect 8404 1362 8460 1406
rect 8564 1362 8620 1406
rect 8852 1362 8908 1476
rect 8956 1468 9028 1476
rect -1075 1247 -1019 1291
rect -4724 1019 -4668 1063
rect -4158 1031 -4102 1075
rect -3998 1031 -3942 1075
rect -3449 1029 -3001 1073
rect -3449 941 -3001 985
rect -2663 1029 -2215 1073
rect -2663 941 -2215 985
rect -1877 1029 -1429 1073
rect -1877 941 -1429 985
rect -1075 1019 -1019 1063
rect -4844 869 -4772 877
rect -4724 869 -4668 919
rect -4844 864 -4668 869
rect -4844 818 -4831 864
rect -4785 818 -4668 864
rect -4337 895 -4265 903
rect -4158 895 -4102 931
rect -4337 890 -4102 895
rect -4337 844 -4324 890
rect -4278 844 -4102 890
rect -4337 839 -4102 844
rect -4337 831 -4262 839
rect -4844 813 -4668 818
rect -4844 805 -4772 813
rect -4724 647 -4668 813
rect -4318 692 -4262 831
rect -4158 692 -4102 839
rect -3998 812 -3942 931
rect -3730 925 -3658 934
rect -3834 921 -3658 925
rect -3834 874 -3717 921
rect -3671 874 -3658 921
rect -3834 869 -3658 874
rect -3834 812 -3778 869
rect -3730 861 -3658 869
rect -3998 756 -3778 812
rect -3378 787 -3306 795
rect -3258 787 -3146 941
rect -3378 782 -3146 787
rect -3998 692 -3942 756
rect -3838 692 -3782 756
rect -3378 736 -3365 782
rect -3319 736 -3146 782
rect -3378 731 -3146 736
rect -3378 723 -3306 731
rect -3258 613 -3146 731
rect -2592 787 -2520 795
rect -2472 787 -2360 941
rect -2592 782 -2360 787
rect -2592 736 -2579 782
rect -2533 736 -2360 782
rect -2592 731 -2360 736
rect -2592 723 -2520 731
rect -2472 613 -2360 731
rect -1806 787 -1734 795
rect -1686 787 -1574 941
rect 196 976 252 1112
rect 484 976 540 1112
rect 644 976 700 1112
rect 804 976 860 1112
rect 964 976 1020 1112
rect 1124 976 1180 1112
rect 1284 976 1340 1112
rect 1444 976 1500 1112
rect 1604 976 1660 1112
rect 2008 976 2064 1112
rect 2168 976 2224 1112
rect 2328 976 2384 1112
rect 2488 976 2544 1112
rect 2648 976 2704 1112
rect 2808 976 2864 1112
rect 2968 976 3024 1112
rect 3128 976 3184 1112
rect 3416 976 3472 1112
rect 3820 976 3876 1112
rect 4108 976 4164 1112
rect 4268 976 4324 1112
rect 4428 976 4484 1112
rect 4588 976 4644 1112
rect 4748 976 4804 1112
rect 4908 976 4964 1112
rect 5068 976 5124 1112
rect 5228 976 5284 1112
rect 5632 976 5688 1112
rect 5792 976 5848 1112
rect 5952 976 6008 1112
rect 6112 976 6168 1112
rect 6272 976 6328 1112
rect 6432 976 6488 1112
rect 6592 976 6648 1112
rect 6752 976 6808 1112
rect 7040 976 7096 1112
rect 7444 976 7500 1112
rect 7604 976 7660 1112
rect 7764 976 7820 1112
rect 7924 976 7980 1112
rect 8084 976 8140 1112
rect 8244 976 8300 1112
rect 8404 976 8460 1112
rect 8564 976 8620 1112
rect 8852 976 8908 1112
rect -1195 869 -1123 877
rect -1075 869 -1019 919
rect -1195 864 -1019 869
rect -1195 818 -1182 864
rect -1136 818 -1019 864
rect -1195 813 -1019 818
rect -1195 805 -1123 813
rect -1806 782 -1574 787
rect -1806 736 -1793 782
rect -1747 736 -1574 782
rect -1806 731 -1574 736
rect -1806 723 -1734 731
rect -1686 613 -1574 731
rect -1075 647 -1019 813
rect -3445 569 -2997 613
rect -2659 569 -2211 613
rect -1873 569 -1425 613
rect -4318 448 -4262 492
rect -4158 448 -4102 492
rect -3998 448 -3942 492
rect -3838 448 -3782 492
rect -4724 403 -4668 447
rect -3445 437 -2997 481
rect -2659 437 -2211 481
rect -1873 437 -1425 481
rect 196 590 252 726
rect 484 590 540 726
rect 644 590 700 726
rect 804 590 860 726
rect 964 590 1020 726
rect 1124 590 1180 726
rect 1284 590 1340 726
rect 1444 590 1500 726
rect 1604 590 1660 726
rect 2008 590 2064 726
rect 2168 590 2224 726
rect 2328 590 2384 726
rect 2488 590 2544 726
rect 2648 590 2704 726
rect 2808 590 2864 726
rect 2968 590 3024 726
rect 3128 590 3184 726
rect 3416 590 3472 726
rect 3820 590 3876 726
rect 4108 590 4164 726
rect 4268 590 4324 726
rect 4428 590 4484 726
rect 4588 590 4644 726
rect 4748 590 4804 726
rect 4908 590 4964 726
rect 5068 590 5124 726
rect 5228 590 5284 726
rect 5632 590 5688 726
rect 5792 590 5848 726
rect 5952 590 6008 726
rect 6112 590 6168 726
rect 6272 590 6328 726
rect 6432 590 6488 726
rect 6592 590 6648 726
rect 6752 590 6808 726
rect 7040 590 7096 726
rect 7444 590 7500 726
rect 7604 590 7660 726
rect 7764 590 7820 726
rect 7924 590 7980 726
rect 8084 590 8140 726
rect 8244 590 8300 726
rect 8404 590 8460 726
rect 8564 590 8620 726
rect 8852 590 8908 726
rect -1075 403 -1019 447
rect 196 320 252 340
rect 484 320 540 340
rect 644 320 700 340
rect 804 320 860 340
rect 964 320 1020 340
rect 1124 320 1180 340
rect 1284 320 1340 340
rect 1444 320 1500 340
rect 1604 320 1660 340
rect 196 264 1660 320
rect 2008 320 2064 340
rect 2168 320 2224 340
rect 2328 320 2384 340
rect 2488 320 2544 340
rect 2648 320 2704 340
rect 2808 320 2864 340
rect 2968 320 3024 340
rect 3128 320 3184 340
rect 3416 320 3472 340
rect 2008 264 3472 320
rect 3820 320 3876 340
rect 4108 320 4164 340
rect 4268 320 4324 340
rect 4428 320 4484 340
rect 4588 320 4644 340
rect 4748 320 4804 340
rect 4908 320 4964 340
rect 5068 320 5124 340
rect 5228 320 5284 340
rect 3820 264 5284 320
rect 5632 320 5688 340
rect 5792 320 5848 340
rect 5952 320 6008 340
rect 6112 320 6168 340
rect 6272 320 6328 340
rect 6432 320 6488 340
rect 6592 320 6648 340
rect 6752 320 6808 340
rect 7040 320 7096 340
rect 5632 264 7096 320
rect 7444 320 7500 340
rect 7604 320 7660 340
rect 7764 320 7820 340
rect 7924 320 7980 340
rect 8084 320 8140 340
rect 8244 320 8300 340
rect 8404 320 8460 340
rect 8564 320 8620 340
rect 8852 320 8908 340
rect 7444 264 8908 320
rect -4724 153 -4668 197
rect -4318 108 -4262 152
rect -4158 108 -4102 152
rect -3998 108 -3942 152
rect -3838 108 -3782 152
rect -3445 119 -2997 163
rect -2659 119 -2211 163
rect -1873 119 -1425 163
rect -1075 153 -1019 197
rect -4844 -213 -4772 -205
rect -4724 -213 -4668 -47
rect -3445 -13 -2997 31
rect -2659 -13 -2211 31
rect -1873 -13 -1425 31
rect -4844 -218 -4668 -213
rect -4844 -264 -4831 -218
rect -4785 -264 -4668 -218
rect -4318 -231 -4262 -92
rect -4844 -269 -4668 -264
rect -4844 -277 -4772 -269
rect -4724 -319 -4668 -269
rect -4337 -239 -4262 -231
rect -4158 -239 -4102 -92
rect -4337 -244 -4102 -239
rect -4337 -290 -4324 -244
rect -4278 -290 -4102 -244
rect -4337 -295 -4102 -290
rect -4337 -303 -4265 -295
rect -4158 -331 -4102 -295
rect -3998 -156 -3942 -92
rect -3838 -156 -3782 -92
rect -3378 -131 -3306 -123
rect -3258 -131 -3146 -13
rect -3378 -136 -3146 -131
rect -3998 -212 -3778 -156
rect -3378 -182 -3365 -136
rect -3319 -182 -3146 -136
rect -3378 -187 -3146 -182
rect -3378 -195 -3306 -187
rect -3998 -331 -3942 -212
rect -3834 -269 -3778 -212
rect -3730 -269 -3658 -261
rect -3834 -274 -3658 -269
rect -3834 -321 -3717 -274
rect -3671 -321 -3658 -274
rect -3834 -325 -3658 -321
rect -4724 -463 -4668 -419
rect -3730 -334 -3658 -325
rect -3258 -341 -3146 -187
rect -2592 -131 -2520 -123
rect -2472 -131 -2360 -13
rect -2592 -136 -2360 -131
rect -2592 -182 -2579 -136
rect -2533 -182 -2360 -136
rect -2592 -187 -2360 -182
rect -2592 -195 -2520 -187
rect -2472 -341 -2360 -187
rect -1806 -131 -1734 -123
rect -1686 -131 -1574 -13
rect -1806 -136 -1574 -131
rect -1806 -182 -1793 -136
rect -1747 -182 -1574 -136
rect -1806 -187 -1574 -182
rect -1806 -195 -1734 -187
rect -1686 -341 -1574 -187
rect -1195 -213 -1123 -205
rect -1075 -213 -1019 -47
rect -1195 -218 -1019 -213
rect -1195 -264 -1182 -218
rect -1136 -264 -1019 -218
rect 196 -208 1660 -152
rect 196 -228 252 -208
rect 484 -228 540 -208
rect 644 -228 700 -208
rect 804 -228 860 -208
rect 964 -228 1020 -208
rect 1124 -228 1180 -208
rect 1284 -228 1340 -208
rect 1444 -228 1500 -208
rect 1604 -228 1660 -208
rect 2008 -208 3472 -152
rect 2008 -228 2064 -208
rect 2168 -228 2224 -208
rect 2328 -228 2384 -208
rect 2488 -228 2544 -208
rect 2648 -228 2704 -208
rect 2808 -228 2864 -208
rect 2968 -228 3024 -208
rect 3128 -228 3184 -208
rect 3416 -228 3472 -208
rect 3820 -208 5284 -152
rect 3820 -228 3876 -208
rect 4108 -228 4164 -208
rect 4268 -228 4324 -208
rect 4428 -228 4484 -208
rect 4588 -228 4644 -208
rect 4748 -228 4804 -208
rect 4908 -228 4964 -208
rect 5068 -228 5124 -208
rect 5228 -228 5284 -208
rect 5632 -208 7096 -152
rect 5632 -228 5688 -208
rect 5792 -228 5848 -208
rect 5952 -228 6008 -208
rect 6112 -228 6168 -208
rect 6272 -228 6328 -208
rect 6432 -228 6488 -208
rect 6592 -228 6648 -208
rect 6752 -228 6808 -208
rect 7040 -228 7096 -208
rect 7444 -208 8908 -152
rect 7444 -228 7500 -208
rect 7604 -228 7660 -208
rect 7764 -228 7820 -208
rect 7924 -228 7980 -208
rect 8084 -228 8140 -208
rect 8244 -228 8300 -208
rect 8404 -228 8460 -208
rect 8564 -228 8620 -208
rect 8852 -228 8908 -208
rect -1195 -269 -1019 -264
rect -1195 -277 -1123 -269
rect -1075 -319 -1019 -269
rect -3449 -385 -3001 -341
rect -4158 -475 -4102 -431
rect -3998 -475 -3942 -431
rect -3449 -473 -3001 -429
rect -2663 -385 -2215 -341
rect -2663 -473 -2215 -429
rect -1877 -385 -1429 -341
rect -1877 -473 -1429 -429
rect -1075 -463 -1019 -419
rect 196 -614 252 -478
rect 484 -614 540 -478
rect 644 -614 700 -478
rect 804 -614 860 -478
rect 964 -614 1020 -478
rect 1124 -614 1180 -478
rect 1284 -614 1340 -478
rect 1444 -614 1500 -478
rect 1604 -614 1660 -478
rect 2008 -614 2064 -478
rect 2168 -614 2224 -478
rect 2328 -614 2384 -478
rect 2488 -614 2544 -478
rect 2648 -614 2704 -478
rect 2808 -614 2864 -478
rect 2968 -614 3024 -478
rect 3128 -614 3184 -478
rect 3416 -614 3472 -478
rect 3820 -614 3876 -478
rect 4108 -614 4164 -478
rect 4268 -614 4324 -478
rect 4428 -614 4484 -478
rect 4588 -614 4644 -478
rect 4748 -614 4804 -478
rect 4908 -614 4964 -478
rect 5068 -614 5124 -478
rect 5228 -614 5284 -478
rect 5632 -614 5688 -478
rect 5792 -614 5848 -478
rect 5952 -614 6008 -478
rect 6112 -614 6168 -478
rect 6272 -614 6328 -478
rect 6432 -614 6488 -478
rect 6592 -614 6648 -478
rect 6752 -614 6808 -478
rect 7040 -614 7096 -478
rect 7444 -614 7500 -478
rect 7604 -614 7660 -478
rect 7764 -614 7820 -478
rect 7924 -614 7980 -478
rect 8084 -614 8140 -478
rect 8244 -614 8300 -478
rect 8404 -614 8460 -478
rect 8564 -614 8620 -478
rect 8852 -614 8908 -478
rect -4158 -679 -4102 -635
rect -3998 -679 -3942 -635
rect -3449 -681 -3001 -637
rect -3449 -769 -3001 -725
rect -2663 -681 -2215 -637
rect -2663 -769 -2215 -725
rect -1877 -681 -1429 -637
rect -1877 -769 -1429 -725
rect -1075 -691 -1019 -647
rect -4337 -815 -4265 -807
rect -4158 -815 -4102 -779
rect -4337 -820 -4102 -815
rect -4337 -866 -4324 -820
rect -4278 -866 -4102 -820
rect -4337 -871 -4102 -866
rect -4337 -879 -4262 -871
rect -4318 -1018 -4262 -879
rect -4158 -1018 -4102 -871
rect -3998 -898 -3942 -779
rect -3730 -785 -3658 -776
rect -3834 -789 -3658 -785
rect -3834 -836 -3717 -789
rect -3671 -836 -3658 -789
rect -3834 -841 -3658 -836
rect -3834 -898 -3778 -841
rect -3730 -849 -3658 -841
rect -3998 -954 -3778 -898
rect -3378 -923 -3306 -915
rect -3258 -923 -3146 -769
rect -3378 -928 -3146 -923
rect -3998 -1018 -3942 -954
rect -3838 -1018 -3782 -954
rect -3378 -974 -3365 -928
rect -3319 -974 -3146 -928
rect -3378 -979 -3146 -974
rect -3378 -987 -3306 -979
rect -3258 -1097 -3146 -979
rect -2592 -923 -2520 -915
rect -2472 -923 -2360 -769
rect -2592 -928 -2360 -923
rect -2592 -974 -2579 -928
rect -2533 -974 -2360 -928
rect -2592 -979 -2360 -974
rect -2592 -987 -2520 -979
rect -2472 -1097 -2360 -979
rect -1806 -923 -1734 -915
rect -1686 -923 -1574 -769
rect -1195 -841 -1123 -833
rect -1075 -841 -1019 -791
rect -1195 -846 -1019 -841
rect -1195 -892 -1182 -846
rect -1136 -892 -1019 -846
rect -1195 -897 -1019 -892
rect -1195 -905 -1123 -897
rect -1806 -928 -1574 -923
rect -1806 -974 -1793 -928
rect -1747 -974 -1574 -928
rect -1806 -979 -1574 -974
rect -1806 -987 -1734 -979
rect -1686 -1097 -1574 -979
rect -1075 -1063 -1019 -897
rect 196 -1000 252 -864
rect 484 -1000 540 -864
rect 644 -1000 700 -864
rect 804 -1000 860 -864
rect 964 -1000 1020 -864
rect 1124 -1000 1180 -864
rect 1284 -1000 1340 -864
rect 1444 -1000 1500 -864
rect 1604 -1000 1660 -864
rect 2008 -1000 2064 -864
rect 2168 -1000 2224 -864
rect 2328 -1000 2384 -864
rect 2488 -1000 2544 -864
rect 2648 -1000 2704 -864
rect 2808 -1000 2864 -864
rect 2968 -1000 3024 -864
rect 3128 -1000 3184 -864
rect 3416 -1000 3472 -864
rect 3820 -1000 3876 -864
rect 4108 -1000 4164 -864
rect 4268 -1000 4324 -864
rect 4428 -1000 4484 -864
rect 4588 -1000 4644 -864
rect 4748 -1000 4804 -864
rect 4908 -1000 4964 -864
rect 5068 -1000 5124 -864
rect 5228 -1000 5284 -864
rect 5632 -1000 5688 -864
rect 5792 -1000 5848 -864
rect 5952 -1000 6008 -864
rect 6112 -1000 6168 -864
rect 6272 -1000 6328 -864
rect 6432 -1000 6488 -864
rect 6592 -1000 6648 -864
rect 6752 -1000 6808 -864
rect 7040 -1000 7096 -864
rect 7444 -1000 7500 -864
rect 7604 -1000 7660 -864
rect 7764 -1000 7820 -864
rect 7924 -1000 7980 -864
rect 8084 -1000 8140 -864
rect 8244 -1000 8300 -864
rect 8404 -1000 8460 -864
rect 8564 -1000 8620 -864
rect 8852 -1000 8908 -864
rect -3445 -1141 -2997 -1097
rect -2659 -1141 -2211 -1097
rect -1873 -1141 -1425 -1097
rect -4318 -1262 -4262 -1218
rect -4158 -1262 -4102 -1218
rect -3998 -1262 -3942 -1218
rect -3838 -1262 -3782 -1218
rect -3445 -1273 -2997 -1229
rect -2659 -1273 -2211 -1229
rect -1873 -1273 -1425 -1229
rect -1075 -1307 -1019 -1263
rect 76 -1364 148 -1356
rect 196 -1364 252 -1250
rect 484 -1294 540 -1250
rect 644 -1294 700 -1250
rect 804 -1294 860 -1250
rect 964 -1294 1020 -1250
rect 1124 -1294 1180 -1250
rect 1284 -1294 1340 -1250
rect 1444 -1294 1500 -1250
rect 1604 -1294 1660 -1250
rect 2008 -1294 2064 -1250
rect 2168 -1294 2224 -1250
rect 2328 -1294 2384 -1250
rect 2488 -1294 2544 -1250
rect 2648 -1294 2704 -1250
rect 2808 -1294 2864 -1250
rect 2968 -1294 3024 -1250
rect 3128 -1294 3184 -1250
rect 76 -1369 252 -1364
rect 3416 -1364 3472 -1250
rect 3520 -1364 3592 -1356
rect 76 -1415 89 -1369
rect 135 -1415 252 -1369
rect 76 -1420 252 -1415
rect 76 -1428 148 -1420
rect 196 -1552 252 -1420
rect 300 -1374 372 -1366
rect 3296 -1374 3368 -1366
rect 300 -1379 540 -1374
rect 300 -1425 313 -1379
rect 359 -1425 540 -1379
rect 300 -1430 540 -1425
rect 300 -1438 372 -1430
rect 484 -1552 540 -1430
rect 3128 -1379 3368 -1374
rect 3128 -1425 3309 -1379
rect 3355 -1425 3368 -1379
rect 3128 -1430 3368 -1425
rect 644 -1552 700 -1508
rect 804 -1552 860 -1508
rect 964 -1552 1020 -1508
rect 1124 -1552 1180 -1508
rect 1284 -1552 1340 -1508
rect 1444 -1552 1500 -1508
rect 1604 -1552 1660 -1508
rect 2008 -1552 2064 -1508
rect 2168 -1552 2224 -1508
rect 2328 -1552 2384 -1508
rect 2488 -1552 2544 -1508
rect 2648 -1552 2704 -1508
rect 2808 -1552 2864 -1508
rect 2968 -1552 3024 -1508
rect 3128 -1552 3184 -1430
rect 3296 -1438 3368 -1430
rect 3416 -1369 3592 -1364
rect 3416 -1415 3533 -1369
rect 3579 -1415 3592 -1369
rect 3416 -1420 3592 -1415
rect 3416 -1552 3472 -1420
rect 3520 -1428 3592 -1420
rect 3700 -1364 3772 -1356
rect 3820 -1364 3876 -1250
rect 4108 -1294 4164 -1250
rect 4268 -1294 4324 -1250
rect 4428 -1294 4484 -1250
rect 4588 -1294 4644 -1250
rect 4748 -1294 4804 -1250
rect 4908 -1294 4964 -1250
rect 5068 -1294 5124 -1250
rect 5228 -1294 5284 -1250
rect 5632 -1294 5688 -1250
rect 5792 -1294 5848 -1250
rect 5952 -1294 6008 -1250
rect 6112 -1294 6168 -1250
rect 6272 -1294 6328 -1250
rect 6432 -1294 6488 -1250
rect 6592 -1294 6648 -1250
rect 6752 -1294 6808 -1250
rect 3700 -1369 3876 -1364
rect 7040 -1364 7096 -1250
rect 7444 -1294 7500 -1250
rect 7604 -1294 7660 -1250
rect 7764 -1294 7820 -1250
rect 7924 -1294 7980 -1250
rect 8084 -1294 8140 -1250
rect 8244 -1294 8300 -1250
rect 8404 -1294 8460 -1250
rect 8564 -1294 8620 -1250
rect 7144 -1364 7216 -1356
rect 8852 -1364 8908 -1250
rect 8956 -1364 9028 -1356
rect 3700 -1415 3713 -1369
rect 3759 -1415 3876 -1369
rect 3700 -1420 3876 -1415
rect 3700 -1428 3772 -1420
rect 3820 -1552 3876 -1420
rect 3924 -1374 3996 -1366
rect 6920 -1374 6992 -1366
rect 3924 -1379 4164 -1374
rect 3924 -1425 3937 -1379
rect 3983 -1425 4164 -1379
rect 3924 -1430 4164 -1425
rect 3924 -1438 3996 -1430
rect 4108 -1552 4164 -1430
rect 6752 -1379 6992 -1374
rect 6752 -1425 6933 -1379
rect 6979 -1425 6992 -1379
rect 6752 -1430 6992 -1425
rect 4268 -1552 4324 -1508
rect 4428 -1552 4484 -1508
rect 4588 -1552 4644 -1508
rect 4748 -1552 4804 -1508
rect 4908 -1552 4964 -1508
rect 5068 -1552 5124 -1508
rect 5228 -1552 5284 -1508
rect 5632 -1552 5688 -1508
rect 5792 -1552 5848 -1508
rect 5952 -1552 6008 -1508
rect 6112 -1552 6168 -1508
rect 6272 -1552 6328 -1508
rect 6432 -1552 6488 -1508
rect 6592 -1552 6648 -1508
rect 6752 -1552 6808 -1430
rect 6920 -1438 6992 -1430
rect 7040 -1369 7218 -1364
rect 7040 -1415 7157 -1369
rect 7203 -1415 7218 -1369
rect 8732 -1374 8804 -1366
rect 7040 -1420 7218 -1415
rect 8564 -1379 8804 -1374
rect 7040 -1552 7096 -1420
rect 7144 -1428 7216 -1420
rect 8564 -1425 8745 -1379
rect 8791 -1425 8804 -1379
rect 8564 -1430 8804 -1425
rect 7444 -1552 7500 -1508
rect 7604 -1552 7660 -1508
rect 7764 -1552 7820 -1508
rect 7924 -1552 7980 -1508
rect 8084 -1552 8140 -1508
rect 8244 -1552 8300 -1508
rect 8404 -1552 8460 -1508
rect 8564 -1552 8620 -1430
rect 8732 -1438 8804 -1430
rect 8852 -1369 9028 -1364
rect 8852 -1415 8969 -1369
rect 9015 -1415 9028 -1369
rect 8852 -1420 9028 -1415
rect 8852 -1552 8908 -1420
rect 8956 -1428 9028 -1420
rect 196 -2188 252 -2052
rect 484 -2188 540 -2052
rect 644 -2188 700 -2052
rect 804 -2188 860 -2052
rect 964 -2188 1020 -2052
rect 1124 -2188 1180 -2052
rect 1284 -2188 1340 -2052
rect 1444 -2188 1500 -2052
rect 1604 -2188 1660 -2052
rect 2008 -2188 2064 -2052
rect 2168 -2188 2224 -2052
rect 2328 -2188 2384 -2052
rect 2488 -2188 2544 -2052
rect 2648 -2188 2704 -2052
rect 2808 -2188 2864 -2052
rect 2968 -2188 3024 -2052
rect 3128 -2188 3184 -2052
rect 3416 -2188 3472 -2052
rect 3820 -2188 3876 -2052
rect 4108 -2188 4164 -2052
rect 4268 -2188 4324 -2052
rect 4428 -2188 4484 -2052
rect 4588 -2188 4644 -2052
rect 4748 -2188 4804 -2052
rect 4908 -2188 4964 -2052
rect 5068 -2188 5124 -2052
rect 5228 -2188 5284 -2052
rect 5632 -2188 5688 -2052
rect 5792 -2188 5848 -2052
rect 5952 -2188 6008 -2052
rect 6112 -2188 6168 -2052
rect 6272 -2188 6328 -2052
rect 6432 -2188 6488 -2052
rect 6592 -2188 6648 -2052
rect 6752 -2188 6808 -2052
rect 7040 -2188 7096 -2052
rect 7444 -2188 7500 -2052
rect 7604 -2188 7660 -2052
rect 7764 -2188 7820 -2052
rect 7924 -2188 7980 -2052
rect 8084 -2188 8140 -2052
rect 8244 -2188 8300 -2052
rect 8404 -2188 8460 -2052
rect 8564 -2188 8620 -2052
rect 8852 -2188 8908 -2052
rect 196 -2824 252 -2688
rect 484 -2824 540 -2688
rect 644 -2824 700 -2688
rect 804 -2824 860 -2688
rect 964 -2824 1020 -2688
rect 1124 -2824 1180 -2688
rect 1284 -2824 1340 -2688
rect 1444 -2824 1500 -2688
rect 1604 -2824 1660 -2688
rect 2008 -2824 2064 -2688
rect 2168 -2824 2224 -2688
rect 2328 -2824 2384 -2688
rect 2488 -2824 2544 -2688
rect 2648 -2824 2704 -2688
rect 2808 -2824 2864 -2688
rect 2968 -2824 3024 -2688
rect 3128 -2824 3184 -2688
rect 3416 -2824 3472 -2688
rect 3820 -2824 3876 -2688
rect 4108 -2824 4164 -2688
rect 4268 -2824 4324 -2688
rect 4428 -2824 4484 -2688
rect 4588 -2824 4644 -2688
rect 4748 -2824 4804 -2688
rect 4908 -2824 4964 -2688
rect 5068 -2824 5124 -2688
rect 5228 -2824 5284 -2688
rect 5632 -2824 5688 -2688
rect 5792 -2824 5848 -2688
rect 5952 -2824 6008 -2688
rect 6112 -2824 6168 -2688
rect 6272 -2824 6328 -2688
rect 6432 -2824 6488 -2688
rect 6592 -2824 6648 -2688
rect 6752 -2824 6808 -2688
rect 7040 -2824 7096 -2688
rect 7444 -2824 7500 -2688
rect 7604 -2824 7660 -2688
rect 7764 -2824 7820 -2688
rect 7924 -2824 7980 -2688
rect 8084 -2824 8140 -2688
rect 8244 -2824 8300 -2688
rect 8404 -2824 8460 -2688
rect 8564 -2824 8620 -2688
rect 8852 -2824 8908 -2688
rect 196 -3368 252 -3324
rect 484 -3344 540 -3324
rect 644 -3344 700 -3324
rect 804 -3344 860 -3324
rect 964 -3344 1020 -3324
rect 1124 -3344 1180 -3324
rect 1284 -3344 1340 -3324
rect 1444 -3344 1500 -3324
rect 1604 -3344 1660 -3324
rect 484 -3400 1660 -3344
rect 2008 -3344 2064 -3324
rect 2168 -3344 2224 -3324
rect 2328 -3344 2384 -3324
rect 2488 -3344 2544 -3324
rect 2648 -3344 2704 -3324
rect 2808 -3344 2864 -3324
rect 2968 -3344 3024 -3324
rect 3128 -3344 3184 -3324
rect 2008 -3400 3184 -3344
rect 3416 -3368 3472 -3324
rect 3820 -3368 3876 -3324
rect 4108 -3344 4164 -3324
rect 4268 -3344 4324 -3324
rect 4428 -3344 4484 -3324
rect 4588 -3344 4644 -3324
rect 4748 -3344 4804 -3324
rect 4908 -3344 4964 -3324
rect 5068 -3344 5124 -3324
rect 5228 -3344 5284 -3324
rect 4108 -3400 5284 -3344
rect 5632 -3344 5688 -3324
rect 5792 -3344 5848 -3324
rect 5952 -3344 6008 -3324
rect 6112 -3344 6168 -3324
rect 6272 -3344 6328 -3324
rect 6432 -3344 6488 -3324
rect 6592 -3344 6648 -3324
rect 6752 -3344 6808 -3324
rect 5632 -3400 6808 -3344
rect 7040 -3368 7096 -3324
rect 7444 -3344 7500 -3324
rect 7604 -3344 7660 -3324
rect 7764 -3344 7820 -3324
rect 7924 -3344 7980 -3324
rect 8084 -3344 8140 -3324
rect 8244 -3344 8300 -3324
rect 8404 -3344 8460 -3324
rect 8564 -3344 8620 -3324
rect 7444 -3400 8620 -3344
rect 8852 -3368 8908 -3324
rect -4001 -3892 -3945 -3848
rect -3713 -3872 -2537 -3816
rect -3713 -3892 -3657 -3872
rect -3553 -3892 -3497 -3872
rect -3393 -3892 -3337 -3872
rect -3233 -3892 -3177 -3872
rect -3073 -3892 -3017 -3872
rect -2913 -3892 -2857 -3872
rect -2753 -3892 -2697 -3872
rect -2593 -3892 -2537 -3872
rect -2189 -3872 -1013 -3816
rect -2189 -3892 -2133 -3872
rect -2029 -3892 -1973 -3872
rect -1869 -3892 -1813 -3872
rect -1709 -3892 -1653 -3872
rect -1549 -3892 -1493 -3872
rect -1389 -3892 -1333 -3872
rect -1229 -3892 -1173 -3872
rect -1069 -3892 -1013 -3872
rect -781 -3892 -725 -3848
rect 196 -3892 252 -3848
rect 484 -3872 1660 -3816
rect 484 -3892 540 -3872
rect 644 -3892 700 -3872
rect 804 -3892 860 -3872
rect 964 -3892 1020 -3872
rect 1124 -3892 1180 -3872
rect 1284 -3892 1340 -3872
rect 1444 -3892 1500 -3872
rect 1604 -3892 1660 -3872
rect 2008 -3872 3184 -3816
rect 2008 -3892 2064 -3872
rect 2168 -3892 2224 -3872
rect 2328 -3892 2384 -3872
rect 2488 -3892 2544 -3872
rect 2648 -3892 2704 -3872
rect 2808 -3892 2864 -3872
rect 2968 -3892 3024 -3872
rect 3128 -3892 3184 -3872
rect 3416 -3892 3472 -3848
rect 3820 -3892 3876 -3848
rect 4108 -3872 5284 -3816
rect 4108 -3892 4164 -3872
rect 4268 -3892 4324 -3872
rect 4428 -3892 4484 -3872
rect 4588 -3892 4644 -3872
rect 4748 -3892 4804 -3872
rect 4908 -3892 4964 -3872
rect 5068 -3892 5124 -3872
rect 5228 -3892 5284 -3872
rect 5632 -3872 6808 -3816
rect 5632 -3892 5688 -3872
rect 5792 -3892 5848 -3872
rect 5952 -3892 6008 -3872
rect 6112 -3892 6168 -3872
rect 6272 -3892 6328 -3872
rect 6432 -3892 6488 -3872
rect 6592 -3892 6648 -3872
rect 6752 -3892 6808 -3872
rect 7040 -3892 7096 -3848
rect 7444 -3872 8620 -3816
rect 7444 -3892 7500 -3872
rect 7604 -3892 7660 -3872
rect 7764 -3892 7820 -3872
rect 7924 -3892 7980 -3872
rect 8084 -3892 8140 -3872
rect 8244 -3892 8300 -3872
rect 8404 -3892 8460 -3872
rect 8564 -3892 8620 -3872
rect 8852 -3892 8908 -3848
rect -4001 -4528 -3945 -4392
rect -3713 -4528 -3657 -4392
rect -3553 -4528 -3497 -4392
rect -3393 -4528 -3337 -4392
rect -3233 -4528 -3177 -4392
rect -3073 -4528 -3017 -4392
rect -2913 -4528 -2857 -4392
rect -2753 -4528 -2697 -4392
rect -2593 -4528 -2537 -4392
rect -2189 -4528 -2133 -4392
rect -2029 -4528 -1973 -4392
rect -1869 -4528 -1813 -4392
rect -1709 -4528 -1653 -4392
rect -1549 -4528 -1493 -4392
rect -1389 -4528 -1333 -4392
rect -1229 -4528 -1173 -4392
rect -1069 -4528 -1013 -4392
rect -781 -4528 -725 -4392
rect 196 -4528 252 -4392
rect 484 -4528 540 -4392
rect 644 -4528 700 -4392
rect 804 -4528 860 -4392
rect 964 -4528 1020 -4392
rect 1124 -4528 1180 -4392
rect 1284 -4528 1340 -4392
rect 1444 -4528 1500 -4392
rect 1604 -4528 1660 -4392
rect 2008 -4528 2064 -4392
rect 2168 -4528 2224 -4392
rect 2328 -4528 2384 -4392
rect 2488 -4528 2544 -4392
rect 2648 -4528 2704 -4392
rect 2808 -4528 2864 -4392
rect 2968 -4528 3024 -4392
rect 3128 -4528 3184 -4392
rect 3416 -4528 3472 -4392
rect 3820 -4528 3876 -4392
rect 4108 -4528 4164 -4392
rect 4268 -4528 4324 -4392
rect 4428 -4528 4484 -4392
rect 4588 -4528 4644 -4392
rect 4748 -4528 4804 -4392
rect 4908 -4528 4964 -4392
rect 5068 -4528 5124 -4392
rect 5228 -4528 5284 -4392
rect 5632 -4528 5688 -4392
rect 5792 -4528 5848 -4392
rect 5952 -4528 6008 -4392
rect 6112 -4528 6168 -4392
rect 6272 -4528 6328 -4392
rect 6432 -4528 6488 -4392
rect 6592 -4528 6648 -4392
rect 6752 -4528 6808 -4392
rect 7040 -4528 7096 -4392
rect 7444 -4528 7500 -4392
rect 7604 -4528 7660 -4392
rect 7764 -4528 7820 -4392
rect 7924 -4528 7980 -4392
rect 8084 -4528 8140 -4392
rect 8244 -4528 8300 -4392
rect 8404 -4528 8460 -4392
rect 8564 -4528 8620 -4392
rect 8852 -4528 8908 -4392
rect -4001 -5164 -3945 -5028
rect -3713 -5164 -3657 -5028
rect -3553 -5164 -3497 -5028
rect -3393 -5164 -3337 -5028
rect -3233 -5164 -3177 -5028
rect -3073 -5164 -3017 -5028
rect -2913 -5164 -2857 -5028
rect -2753 -5164 -2697 -5028
rect -2593 -5164 -2537 -5028
rect -2189 -5164 -2133 -5028
rect -2029 -5164 -1973 -5028
rect -1869 -5164 -1813 -5028
rect -1709 -5164 -1653 -5028
rect -1549 -5164 -1493 -5028
rect -1389 -5164 -1333 -5028
rect -1229 -5164 -1173 -5028
rect -1069 -5164 -1013 -5028
rect -781 -5164 -725 -5028
rect 196 -5164 252 -5028
rect 484 -5164 540 -5028
rect 644 -5164 700 -5028
rect 804 -5164 860 -5028
rect 964 -5164 1020 -5028
rect 1124 -5164 1180 -5028
rect 1284 -5164 1340 -5028
rect 1444 -5164 1500 -5028
rect 1604 -5164 1660 -5028
rect 2008 -5164 2064 -5028
rect 2168 -5164 2224 -5028
rect 2328 -5164 2384 -5028
rect 2488 -5164 2544 -5028
rect 2648 -5164 2704 -5028
rect 2808 -5164 2864 -5028
rect 2968 -5164 3024 -5028
rect 3128 -5164 3184 -5028
rect 3416 -5164 3472 -5028
rect 3820 -5164 3876 -5028
rect 4108 -5164 4164 -5028
rect 4268 -5164 4324 -5028
rect 4428 -5164 4484 -5028
rect 4588 -5164 4644 -5028
rect 4748 -5164 4804 -5028
rect 4908 -5164 4964 -5028
rect 5068 -5164 5124 -5028
rect 5228 -5164 5284 -5028
rect 5632 -5164 5688 -5028
rect 5792 -5164 5848 -5028
rect 5952 -5164 6008 -5028
rect 6112 -5164 6168 -5028
rect 6272 -5164 6328 -5028
rect 6432 -5164 6488 -5028
rect 6592 -5164 6648 -5028
rect 6752 -5164 6808 -5028
rect 7040 -5164 7096 -5028
rect 7444 -5164 7500 -5028
rect 7604 -5164 7660 -5028
rect 7764 -5164 7820 -5028
rect 7924 -5164 7980 -5028
rect 8084 -5164 8140 -5028
rect 8244 -5164 8300 -5028
rect 8404 -5164 8460 -5028
rect 8564 -5164 8620 -5028
rect 8852 -5164 8908 -5028
rect -4121 -5796 -4049 -5788
rect -4001 -5796 -3945 -5664
rect -4121 -5801 -3945 -5796
rect -4121 -5847 -4108 -5801
rect -4062 -5847 -3945 -5801
rect -4121 -5852 -3945 -5847
rect -3897 -5786 -3825 -5778
rect -3713 -5786 -3657 -5664
rect -3553 -5708 -3497 -5664
rect -3393 -5708 -3337 -5664
rect -3233 -5708 -3177 -5664
rect -3073 -5708 -3017 -5664
rect -2913 -5708 -2857 -5664
rect -2753 -5708 -2697 -5664
rect -2593 -5708 -2537 -5664
rect -2189 -5708 -2133 -5664
rect -2029 -5708 -1973 -5664
rect -1869 -5708 -1813 -5664
rect -1709 -5708 -1653 -5664
rect -1549 -5708 -1493 -5664
rect -1389 -5708 -1333 -5664
rect -1229 -5708 -1173 -5664
rect -3897 -5791 -3657 -5786
rect -3897 -5837 -3884 -5791
rect -3838 -5837 -3657 -5791
rect -3897 -5842 -3657 -5837
rect -1069 -5786 -1013 -5664
rect -901 -5786 -829 -5778
rect -1069 -5791 -829 -5786
rect -1069 -5837 -888 -5791
rect -842 -5837 -829 -5791
rect -1069 -5842 -829 -5837
rect -3897 -5850 -3825 -5842
rect -901 -5850 -829 -5842
rect -781 -5796 -725 -5664
rect -677 -5796 -605 -5788
rect -781 -5801 -605 -5796
rect -781 -5847 -664 -5801
rect -618 -5847 -605 -5801
rect -4121 -5860 -4049 -5852
rect -4001 -5966 -3945 -5852
rect -781 -5852 -605 -5847
rect -3713 -5966 -3657 -5922
rect -3553 -5966 -3497 -5922
rect -3393 -5966 -3337 -5922
rect -3233 -5966 -3177 -5922
rect -3073 -5966 -3017 -5922
rect -2913 -5966 -2857 -5922
rect -2753 -5966 -2697 -5922
rect -2593 -5966 -2537 -5922
rect -2189 -5966 -2133 -5922
rect -2029 -5966 -1973 -5922
rect -1869 -5966 -1813 -5922
rect -1709 -5966 -1653 -5922
rect -1549 -5966 -1493 -5922
rect -1389 -5966 -1333 -5922
rect -1229 -5966 -1173 -5922
rect -1069 -5966 -1013 -5922
rect -781 -5966 -725 -5852
rect -677 -5860 -605 -5852
rect 76 -5796 148 -5788
rect 196 -5796 252 -5664
rect 76 -5801 252 -5796
rect 76 -5847 89 -5801
rect 135 -5847 252 -5801
rect 76 -5852 252 -5847
rect 300 -5786 372 -5778
rect 484 -5786 540 -5664
rect 644 -5708 700 -5664
rect 804 -5708 860 -5664
rect 964 -5708 1020 -5664
rect 1124 -5708 1180 -5664
rect 1284 -5708 1340 -5664
rect 1444 -5708 1500 -5664
rect 1604 -5708 1660 -5664
rect 2008 -5708 2064 -5664
rect 2168 -5708 2224 -5664
rect 2328 -5708 2384 -5664
rect 2488 -5708 2544 -5664
rect 2648 -5708 2704 -5664
rect 2808 -5708 2864 -5664
rect 2968 -5708 3024 -5664
rect 300 -5791 540 -5786
rect 300 -5837 313 -5791
rect 359 -5837 540 -5791
rect 300 -5842 540 -5837
rect 3128 -5786 3184 -5664
rect 3296 -5786 3368 -5778
rect 3128 -5791 3368 -5786
rect 3128 -5837 3309 -5791
rect 3355 -5837 3368 -5791
rect 3128 -5842 3368 -5837
rect 300 -5850 372 -5842
rect 3296 -5850 3368 -5842
rect 3416 -5796 3472 -5664
rect 3520 -5796 3592 -5788
rect 3416 -5801 3592 -5796
rect 3416 -5847 3533 -5801
rect 3579 -5847 3592 -5801
rect 76 -5860 148 -5852
rect 196 -5966 252 -5852
rect 3416 -5852 3592 -5847
rect 484 -5966 540 -5922
rect 644 -5966 700 -5922
rect 804 -5966 860 -5922
rect 964 -5966 1020 -5922
rect 1124 -5966 1180 -5922
rect 1284 -5966 1340 -5922
rect 1444 -5966 1500 -5922
rect 1604 -5966 1660 -5922
rect 2008 -5966 2064 -5922
rect 2168 -5966 2224 -5922
rect 2328 -5966 2384 -5922
rect 2488 -5966 2544 -5922
rect 2648 -5966 2704 -5922
rect 2808 -5966 2864 -5922
rect 2968 -5966 3024 -5922
rect 3128 -5966 3184 -5922
rect 3416 -5966 3472 -5852
rect 3520 -5860 3592 -5852
rect 3700 -5796 3772 -5788
rect 3820 -5796 3876 -5664
rect 3700 -5801 3876 -5796
rect 3700 -5847 3713 -5801
rect 3759 -5847 3876 -5801
rect 3700 -5852 3876 -5847
rect 3924 -5786 3996 -5778
rect 4108 -5786 4164 -5664
rect 4268 -5708 4324 -5664
rect 4428 -5708 4484 -5664
rect 4588 -5708 4644 -5664
rect 4748 -5708 4804 -5664
rect 4908 -5708 4964 -5664
rect 5068 -5708 5124 -5664
rect 5228 -5708 5284 -5664
rect 5632 -5708 5688 -5664
rect 5792 -5708 5848 -5664
rect 5952 -5708 6008 -5664
rect 6112 -5708 6168 -5664
rect 6272 -5708 6328 -5664
rect 6432 -5708 6488 -5664
rect 6592 -5708 6648 -5664
rect 3924 -5791 4164 -5786
rect 3924 -5837 3937 -5791
rect 3983 -5837 4164 -5791
rect 3924 -5842 4164 -5837
rect 6752 -5786 6808 -5664
rect 6920 -5786 6992 -5778
rect 6752 -5791 6992 -5786
rect 6752 -5837 6933 -5791
rect 6979 -5837 6992 -5791
rect 6752 -5842 6992 -5837
rect 3924 -5850 3996 -5842
rect 6920 -5850 6992 -5842
rect 7040 -5796 7096 -5664
rect 7444 -5708 7500 -5664
rect 7604 -5708 7660 -5664
rect 7764 -5708 7820 -5664
rect 7924 -5708 7980 -5664
rect 8084 -5708 8140 -5664
rect 8244 -5708 8300 -5664
rect 8404 -5708 8460 -5664
rect 8564 -5786 8620 -5664
rect 8732 -5786 8804 -5778
rect 7144 -5796 7216 -5788
rect 7040 -5801 7216 -5796
rect 7040 -5847 7157 -5801
rect 7203 -5847 7216 -5801
rect 8564 -5791 8804 -5786
rect 8564 -5837 8745 -5791
rect 8791 -5837 8804 -5791
rect 8564 -5842 8804 -5837
rect 3700 -5860 3772 -5852
rect 3820 -5966 3876 -5852
rect 7040 -5852 7216 -5847
rect 8732 -5850 8804 -5842
rect 8852 -5796 8908 -5664
rect 8956 -5796 9028 -5788
rect 8852 -5801 9028 -5796
rect 8852 -5847 8969 -5801
rect 9015 -5847 9028 -5801
rect 4108 -5966 4164 -5922
rect 4268 -5966 4324 -5922
rect 4428 -5966 4484 -5922
rect 4588 -5966 4644 -5922
rect 4748 -5966 4804 -5922
rect 4908 -5966 4964 -5922
rect 5068 -5966 5124 -5922
rect 5228 -5966 5284 -5922
rect 5632 -5966 5688 -5922
rect 5792 -5966 5848 -5922
rect 5952 -5966 6008 -5922
rect 6112 -5966 6168 -5922
rect 6272 -5966 6328 -5922
rect 6432 -5966 6488 -5922
rect 6592 -5966 6648 -5922
rect 6752 -5966 6808 -5922
rect 7040 -5966 7096 -5852
rect 7144 -5860 7216 -5852
rect 8852 -5852 9028 -5847
rect 7444 -5966 7500 -5922
rect 7604 -5966 7660 -5922
rect 7764 -5966 7820 -5922
rect 7924 -5966 7980 -5922
rect 8084 -5966 8140 -5922
rect 8244 -5966 8300 -5922
rect 8404 -5966 8460 -5922
rect 8564 -5966 8620 -5922
rect 8852 -5966 8908 -5852
rect 8956 -5860 9028 -5852
rect -4001 -6352 -3945 -6216
rect -3713 -6352 -3657 -6216
rect -3553 -6352 -3497 -6216
rect -3393 -6352 -3337 -6216
rect -3233 -6352 -3177 -6216
rect -3073 -6352 -3017 -6216
rect -2913 -6352 -2857 -6216
rect -2753 -6352 -2697 -6216
rect -2593 -6352 -2537 -6216
rect -2189 -6352 -2133 -6216
rect -2029 -6352 -1973 -6216
rect -1869 -6352 -1813 -6216
rect -1709 -6352 -1653 -6216
rect -1549 -6352 -1493 -6216
rect -1389 -6352 -1333 -6216
rect -1229 -6352 -1173 -6216
rect -1069 -6352 -1013 -6216
rect -781 -6352 -725 -6216
rect 196 -6352 252 -6216
rect 484 -6352 540 -6216
rect 644 -6352 700 -6216
rect 804 -6352 860 -6216
rect 964 -6352 1020 -6216
rect 1124 -6352 1180 -6216
rect 1284 -6352 1340 -6216
rect 1444 -6352 1500 -6216
rect 1604 -6352 1660 -6216
rect 2008 -6352 2064 -6216
rect 2168 -6352 2224 -6216
rect 2328 -6352 2384 -6216
rect 2488 -6352 2544 -6216
rect 2648 -6352 2704 -6216
rect 2808 -6352 2864 -6216
rect 2968 -6352 3024 -6216
rect 3128 -6352 3184 -6216
rect 3416 -6352 3472 -6216
rect 3820 -6352 3876 -6216
rect 4108 -6352 4164 -6216
rect 4268 -6352 4324 -6216
rect 4428 -6352 4484 -6216
rect 4588 -6352 4644 -6216
rect 4748 -6352 4804 -6216
rect 4908 -6352 4964 -6216
rect 5068 -6352 5124 -6216
rect 5228 -6352 5284 -6216
rect 5632 -6352 5688 -6216
rect 5792 -6352 5848 -6216
rect 5952 -6352 6008 -6216
rect 6112 -6352 6168 -6216
rect 6272 -6352 6328 -6216
rect 6432 -6352 6488 -6216
rect 6592 -6352 6648 -6216
rect 6752 -6352 6808 -6216
rect 7040 -6352 7096 -6216
rect 7444 -6352 7500 -6216
rect 7604 -6352 7660 -6216
rect 7764 -6352 7820 -6216
rect 7924 -6352 7980 -6216
rect 8084 -6352 8140 -6216
rect 8244 -6352 8300 -6216
rect 8404 -6352 8460 -6216
rect 8564 -6352 8620 -6216
rect 8852 -6352 8908 -6216
rect -4001 -6738 -3945 -6602
rect -3713 -6738 -3657 -6602
rect -3553 -6738 -3497 -6602
rect -3393 -6738 -3337 -6602
rect -3233 -6738 -3177 -6602
rect -3073 -6738 -3017 -6602
rect -2913 -6738 -2857 -6602
rect -2753 -6738 -2697 -6602
rect -2593 -6738 -2537 -6602
rect -2189 -6738 -2133 -6602
rect -2029 -6738 -1973 -6602
rect -1869 -6738 -1813 -6602
rect -1709 -6738 -1653 -6602
rect -1549 -6738 -1493 -6602
rect -1389 -6738 -1333 -6602
rect -1229 -6738 -1173 -6602
rect -1069 -6738 -1013 -6602
rect -781 -6738 -725 -6602
rect 196 -6738 252 -6602
rect 484 -6738 540 -6602
rect 644 -6738 700 -6602
rect 804 -6738 860 -6602
rect 964 -6738 1020 -6602
rect 1124 -6738 1180 -6602
rect 1284 -6738 1340 -6602
rect 1444 -6738 1500 -6602
rect 1604 -6738 1660 -6602
rect 2008 -6738 2064 -6602
rect 2168 -6738 2224 -6602
rect 2328 -6738 2384 -6602
rect 2488 -6738 2544 -6602
rect 2648 -6738 2704 -6602
rect 2808 -6738 2864 -6602
rect 2968 -6738 3024 -6602
rect 3128 -6738 3184 -6602
rect 3416 -6738 3472 -6602
rect 3820 -6738 3876 -6602
rect 4108 -6738 4164 -6602
rect 4268 -6738 4324 -6602
rect 4428 -6738 4484 -6602
rect 4588 -6738 4644 -6602
rect 4748 -6738 4804 -6602
rect 4908 -6738 4964 -6602
rect 5068 -6738 5124 -6602
rect 5228 -6738 5284 -6602
rect 5632 -6738 5688 -6602
rect 5792 -6738 5848 -6602
rect 5952 -6738 6008 -6602
rect 6112 -6738 6168 -6602
rect 6272 -6738 6328 -6602
rect 6432 -6738 6488 -6602
rect 6592 -6738 6648 -6602
rect 6752 -6738 6808 -6602
rect 7040 -6738 7096 -6602
rect 7444 -6738 7500 -6602
rect 7604 -6738 7660 -6602
rect 7764 -6738 7820 -6602
rect 7924 -6738 7980 -6602
rect 8084 -6738 8140 -6602
rect 8244 -6738 8300 -6602
rect 8404 -6738 8460 -6602
rect 8564 -6738 8620 -6602
rect 8852 -6738 8908 -6602
rect -4001 -7008 -3945 -6988
rect -3713 -7008 -3657 -6988
rect -3553 -7008 -3497 -6988
rect -3393 -7008 -3337 -6988
rect -3233 -7008 -3177 -6988
rect -3073 -7008 -3017 -6988
rect -2913 -7008 -2857 -6988
rect -2753 -7008 -2697 -6988
rect -2593 -7008 -2537 -6988
rect -4001 -7064 -2537 -7008
rect -2189 -7008 -2133 -6988
rect -2029 -7008 -1973 -6988
rect -1869 -7008 -1813 -6988
rect -1709 -7008 -1653 -6988
rect -1549 -7008 -1493 -6988
rect -1389 -7008 -1333 -6988
rect -1229 -7008 -1173 -6988
rect -1069 -7008 -1013 -6988
rect -781 -7008 -725 -6988
rect -2189 -7064 -725 -7008
rect 196 -7008 252 -6988
rect 484 -7008 540 -6988
rect 644 -7008 700 -6988
rect 804 -7008 860 -6988
rect 964 -7008 1020 -6988
rect 1124 -7008 1180 -6988
rect 1284 -7008 1340 -6988
rect 1444 -7008 1500 -6988
rect 1604 -7008 1660 -6988
rect 196 -7064 1660 -7008
rect 2008 -7008 2064 -6988
rect 2168 -7008 2224 -6988
rect 2328 -7008 2384 -6988
rect 2488 -7008 2544 -6988
rect 2648 -7008 2704 -6988
rect 2808 -7008 2864 -6988
rect 2968 -7008 3024 -6988
rect 3128 -7008 3184 -6988
rect 3416 -7008 3472 -6988
rect 2008 -7064 3472 -7008
rect 3820 -7008 3876 -6988
rect 4108 -7008 4164 -6988
rect 4268 -7008 4324 -6988
rect 4428 -7008 4484 -6988
rect 4588 -7008 4644 -6988
rect 4748 -7008 4804 -6988
rect 4908 -7008 4964 -6988
rect 5068 -7008 5124 -6988
rect 5228 -7008 5284 -6988
rect 3820 -7064 5284 -7008
rect 5632 -7008 5688 -6988
rect 5792 -7008 5848 -6988
rect 5952 -7008 6008 -6988
rect 6112 -7008 6168 -6988
rect 6272 -7008 6328 -6988
rect 6432 -7008 6488 -6988
rect 6592 -7008 6648 -6988
rect 6752 -7008 6808 -6988
rect 7040 -7008 7096 -6988
rect 5632 -7064 7096 -7008
rect 7444 -7008 7500 -6988
rect 7604 -7008 7660 -6988
rect 7764 -7008 7820 -6988
rect 7924 -7008 7980 -6988
rect 8084 -7008 8140 -6988
rect 8244 -7008 8300 -6988
rect 8404 -7008 8460 -6988
rect 8564 -7008 8620 -6988
rect 8852 -7008 8908 -6988
rect 7444 -7064 8908 -7008
<< polycontact >>
rect 1497 5903 1543 5949
rect 1721 5913 1767 5959
rect 1901 5913 1947 5959
rect 2125 5903 2171 5949
rect 3713 5913 3759 5959
rect 3937 5903 3983 5949
rect 5525 5913 5571 5959
rect 5749 5903 5795 5949
rect 7337 5913 7383 5959
rect 7561 5903 7607 5949
rect -4831 3156 -4785 3202
rect -4324 3130 -4278 3176
rect -3365 3238 -3319 3284
rect -3717 3099 -3671 3146
rect -2579 3238 -2533 3284
rect -1793 3238 -1747 3284
rect -1182 3156 -1136 3202
rect -4324 2554 -4278 2600
rect -3717 2584 -3671 2631
rect -3365 2446 -3319 2492
rect -2579 2446 -2533 2492
rect -1182 2528 -1136 2574
rect -1793 2446 -1747 2492
rect -4324 1420 -4278 1466
rect -3365 1528 -3319 1574
rect -3717 1389 -3671 1436
rect -2579 1528 -2533 1574
rect -1793 1528 -1747 1574
rect -1182 1446 -1136 1492
rect 89 1481 135 1527
rect 313 1491 359 1537
rect 3309 1491 3355 1537
rect 3533 1481 3579 1527
rect 3713 1481 3759 1527
rect 3937 1491 3983 1537
rect 6933 1491 6979 1537
rect 7157 1481 7203 1527
rect 8745 1491 8791 1537
rect 8969 1481 9015 1527
rect -4831 818 -4785 864
rect -4324 844 -4278 890
rect -3717 874 -3671 921
rect -3365 736 -3319 782
rect -2579 736 -2533 782
rect -1182 818 -1136 864
rect -1793 736 -1747 782
rect -4831 -264 -4785 -218
rect -4324 -290 -4278 -244
rect -3365 -182 -3319 -136
rect -3717 -321 -3671 -274
rect -2579 -182 -2533 -136
rect -1793 -182 -1747 -136
rect -1182 -264 -1136 -218
rect -4324 -866 -4278 -820
rect -3717 -836 -3671 -789
rect -3365 -974 -3319 -928
rect -2579 -974 -2533 -928
rect -1182 -892 -1136 -846
rect -1793 -974 -1747 -928
rect 89 -1415 135 -1369
rect 313 -1425 359 -1379
rect 3309 -1425 3355 -1379
rect 3533 -1415 3579 -1369
rect 3713 -1415 3759 -1369
rect 3937 -1425 3983 -1379
rect 6933 -1425 6979 -1379
rect 7157 -1415 7203 -1369
rect 8745 -1425 8791 -1379
rect 8969 -1415 9015 -1369
rect -4108 -5847 -4062 -5801
rect -3884 -5837 -3838 -5791
rect -888 -5837 -842 -5791
rect -664 -5847 -618 -5801
rect 89 -5847 135 -5801
rect 313 -5837 359 -5791
rect 3309 -5837 3355 -5791
rect 3533 -5847 3579 -5801
rect 3713 -5847 3759 -5801
rect 3937 -5837 3983 -5791
rect 6933 -5837 6979 -5791
rect 7157 -5847 7203 -5801
rect 8745 -5837 8791 -5791
rect 8969 -5847 9015 -5801
<< metal1 >>
rect 1226 7875 1302 7887
rect 1226 7823 1238 7875
rect 1290 7872 1302 7875
rect 1290 7826 9391 7872
rect 1290 7823 1302 7826
rect 1226 7811 1302 7823
rect 3006 7767 3082 7779
rect 3006 7715 3018 7767
rect 3070 7763 3082 7767
rect 3070 7717 9385 7763
rect 3070 7715 3082 7717
rect 3006 7703 3082 7715
rect 4818 7658 4894 7670
rect 4818 7606 4830 7658
rect 4882 7655 4894 7658
rect 4882 7609 9382 7655
rect 4882 7606 4894 7609
rect 4818 7594 4894 7606
rect 6630 7551 6706 7563
rect 6630 7499 6642 7551
rect 6694 7548 6706 7551
rect 6694 7502 9376 7548
rect 6694 7499 6706 7502
rect 6630 7487 6706 7499
rect 84 7410 9020 7440
rect 84 7407 855 7410
rect 907 7407 8197 7410
rect 8249 7407 9020 7410
rect 84 7361 106 7407
rect 152 7361 200 7407
rect 246 7361 294 7407
rect 340 7361 388 7407
rect 434 7361 482 7407
rect 528 7361 576 7407
rect 622 7361 670 7407
rect 716 7361 764 7407
rect 810 7361 855 7407
rect 907 7361 952 7407
rect 998 7361 1046 7407
rect 1092 7361 1140 7407
rect 1186 7361 1234 7407
rect 1280 7361 1328 7407
rect 1374 7361 1422 7407
rect 1468 7361 1516 7407
rect 1562 7361 1610 7407
rect 1656 7361 1704 7407
rect 1750 7361 1918 7407
rect 1964 7361 2012 7407
rect 2058 7361 2106 7407
rect 2152 7361 2200 7407
rect 2246 7361 2294 7407
rect 2340 7361 2388 7407
rect 2434 7361 2482 7407
rect 2528 7361 2576 7407
rect 2622 7361 2670 7407
rect 2716 7361 2764 7407
rect 2810 7361 2858 7407
rect 2904 7361 2952 7407
rect 2998 7361 3046 7407
rect 3092 7361 3140 7407
rect 3186 7361 3234 7407
rect 3280 7361 3328 7407
rect 3374 7361 3422 7407
rect 3468 7361 3516 7407
rect 3562 7361 3730 7407
rect 3776 7361 3824 7407
rect 3870 7361 3918 7407
rect 3964 7361 4012 7407
rect 4058 7361 4106 7407
rect 4152 7361 4200 7407
rect 4246 7361 4294 7407
rect 4340 7361 4388 7407
rect 4434 7361 4482 7407
rect 4528 7361 4576 7407
rect 4622 7361 4670 7407
rect 4716 7361 4764 7407
rect 4810 7361 4858 7407
rect 4904 7361 4952 7407
rect 4998 7361 5046 7407
rect 5092 7361 5140 7407
rect 5186 7361 5234 7407
rect 5280 7361 5328 7407
rect 5374 7361 5542 7407
rect 5588 7361 5636 7407
rect 5682 7361 5730 7407
rect 5776 7361 5824 7407
rect 5870 7361 5918 7407
rect 5964 7361 6012 7407
rect 6058 7361 6106 7407
rect 6152 7361 6200 7407
rect 6246 7361 6294 7407
rect 6340 7361 6388 7407
rect 6434 7361 6482 7407
rect 6528 7361 6576 7407
rect 6622 7361 6670 7407
rect 6716 7361 6764 7407
rect 6810 7361 6858 7407
rect 6904 7361 6952 7407
rect 6998 7361 7046 7407
rect 7092 7361 7140 7407
rect 7186 7361 7354 7407
rect 7400 7361 7448 7407
rect 7494 7361 7542 7407
rect 7588 7361 7636 7407
rect 7682 7361 7730 7407
rect 7776 7361 7824 7407
rect 7870 7361 7918 7407
rect 7964 7361 8012 7407
rect 8058 7361 8106 7407
rect 8152 7361 8197 7407
rect 8249 7361 8294 7407
rect 8340 7361 8388 7407
rect 8434 7361 8482 7407
rect 8528 7361 8576 7407
rect 8622 7361 8670 7407
rect 8716 7361 8764 7407
rect 8810 7361 8858 7407
rect 8904 7361 8952 7407
rect 8998 7361 9020 7407
rect 84 7358 855 7361
rect 907 7358 8197 7361
rect 8249 7358 9020 7361
rect 84 7328 9020 7358
rect 441 7236 1447 7282
rect 441 7190 487 7236
rect 121 7144 487 7190
rect 121 7087 167 7144
rect 121 6701 167 6863
rect 121 6315 167 6477
rect 121 6080 167 6091
rect 281 7087 327 7098
rect 281 6701 327 6863
rect 281 6315 327 6477
rect 281 5984 327 6091
rect 441 7087 487 7144
rect 441 6701 487 6863
rect 441 6315 487 6477
rect 441 6080 487 6091
rect 601 7178 1302 7190
rect 601 7144 1238 7178
rect 601 7087 647 7144
rect 601 6701 647 6863
rect 601 6315 647 6477
rect 601 5984 647 6091
rect 178 5938 647 5984
rect 13 5763 167 5789
rect 13 5743 121 5763
rect 121 5127 167 5289
rect 121 4491 167 4653
rect 121 3960 167 4017
rect 281 5763 327 5938
rect 281 5127 327 5289
rect 281 4491 327 4653
rect 281 4006 327 4017
rect 441 5763 487 5774
rect 441 5127 487 5289
rect 441 4491 487 4653
rect 441 3960 487 4017
rect 121 3914 487 3960
rect 601 5763 647 5938
rect 601 5127 647 5289
rect 601 4491 647 4653
rect 601 3960 647 4017
rect 761 7087 807 7098
rect 761 6701 807 6863
rect 761 6315 807 6477
rect 761 6034 807 6091
rect 921 7087 967 7144
rect 1226 7126 1238 7144
rect 1290 7126 1302 7178
rect 1226 7114 1302 7126
rect 921 6701 967 6863
rect 921 6315 967 6477
rect 921 6080 967 6091
rect 1081 7087 1127 7098
rect 1081 6701 1127 6863
rect 1081 6315 1127 6477
rect 1081 6034 1127 6091
rect 1241 7087 1287 7114
rect 1241 6701 1287 6863
rect 1241 6315 1287 6477
rect 1241 6080 1287 6091
rect 1401 7087 1447 7236
rect 1401 6701 1447 6863
rect 1401 6315 1447 6477
rect 1401 6034 1447 6091
rect 761 5988 1447 6034
rect 1529 7087 1575 7098
rect 1529 6701 1575 6863
rect 1529 6315 1575 6477
rect 761 5866 807 5988
rect 1529 5960 1575 6091
rect 1689 7087 1735 7328
rect 1689 6701 1735 6863
rect 1689 6315 1735 6477
rect 1689 6080 1735 6091
rect 1933 7087 1979 7328
rect 2221 7236 3227 7282
rect 1933 6701 1979 6863
rect 1933 6315 1979 6477
rect 1933 6080 1979 6091
rect 2093 7087 2139 7098
rect 2093 6701 2139 6863
rect 2093 6315 2139 6477
rect 1486 5949 1575 5960
rect 1486 5903 1497 5949
rect 1543 5903 1575 5949
rect 1486 5892 1575 5903
rect 1710 5959 1778 5970
rect 1886 5962 1962 5974
rect 1886 5959 1898 5962
rect 1710 5913 1721 5959
rect 1767 5913 1898 5959
rect 1710 5902 1778 5913
rect 1886 5910 1898 5913
rect 1950 5910 1962 5962
rect 1886 5898 1962 5910
rect 2093 5960 2139 6091
rect 2221 7087 2267 7236
rect 3181 7190 3227 7236
rect 2221 6701 2267 6863
rect 2221 6315 2267 6477
rect 2221 6034 2267 6091
rect 2381 7178 3082 7190
rect 2381 7144 3018 7178
rect 2381 7087 2427 7144
rect 2381 6701 2427 6863
rect 2381 6315 2427 6477
rect 2381 6080 2427 6091
rect 2541 7087 2587 7098
rect 2541 6701 2587 6863
rect 2541 6315 2587 6477
rect 2541 6034 2587 6091
rect 2701 7087 2747 7144
rect 3006 7126 3018 7144
rect 3070 7126 3082 7178
rect 3006 7114 3082 7126
rect 3181 7144 3547 7190
rect 2701 6701 2747 6863
rect 2701 6315 2747 6477
rect 2701 6080 2747 6091
rect 2861 7087 2907 7098
rect 2861 6701 2907 6863
rect 2861 6315 2907 6477
rect 2861 6034 2907 6091
rect 2221 5988 2907 6034
rect 2093 5949 2182 5960
rect 2093 5903 2125 5949
rect 2171 5903 2182 5949
rect 761 5820 1447 5866
rect 761 5763 807 5820
rect 761 5127 807 5289
rect 761 4491 807 4653
rect 761 4006 807 4017
rect 921 5763 967 5774
rect 921 5127 967 5289
rect 921 4491 967 4653
rect 921 3960 967 4017
rect 1081 5763 1127 5820
rect 1081 5127 1127 5289
rect 1081 4491 1127 4653
rect 1081 4006 1127 4017
rect 1241 5763 1287 5774
rect 1241 5127 1287 5289
rect 1241 4491 1287 4653
rect 1241 3960 1287 4017
rect 601 3914 1287 3960
rect 1401 5763 1447 5820
rect 1401 5127 1447 5289
rect 1401 4491 1447 4653
rect 441 3868 487 3914
rect 1401 3898 1447 4017
rect 1529 5763 1575 5892
rect 2093 5892 2182 5903
rect 1529 5127 1575 5289
rect 1529 4491 1575 4653
rect 1529 4006 1575 4017
rect 1689 5763 1735 5774
rect 1689 5127 1735 5289
rect 1689 4491 1735 4653
rect 1381 3886 1457 3898
rect 1381 3868 1393 3886
rect 441 3834 1393 3868
rect 1445 3834 1457 3886
rect 441 3822 1457 3834
rect 1689 3776 1735 4017
rect 1933 5763 1979 5774
rect 1933 5127 1979 5289
rect 1933 4491 1979 4653
rect 1933 3776 1979 4017
rect 2093 5763 2139 5892
rect 2861 5866 2907 5988
rect 2093 5127 2139 5289
rect 2093 4491 2139 4653
rect 2093 4006 2139 4017
rect 2221 5820 2907 5866
rect 2221 5763 2267 5820
rect 2221 5127 2267 5289
rect 2221 4491 2267 4653
rect 2221 3898 2267 4017
rect 2381 5763 2427 5774
rect 2381 5127 2427 5289
rect 2381 4491 2427 4653
rect 2381 3960 2427 4017
rect 2541 5763 2587 5820
rect 2541 5127 2587 5289
rect 2541 4491 2587 4653
rect 2541 4006 2587 4017
rect 2701 5763 2747 5774
rect 2701 5127 2747 5289
rect 2701 4491 2747 4653
rect 2701 3960 2747 4017
rect 2861 5763 2907 5820
rect 2861 5127 2907 5289
rect 2861 4491 2907 4653
rect 2861 4006 2907 4017
rect 3021 7087 3067 7114
rect 3021 6701 3067 6863
rect 3021 6315 3067 6477
rect 3021 5984 3067 6091
rect 3181 7087 3227 7144
rect 3181 6701 3227 6863
rect 3181 6315 3227 6477
rect 3181 6080 3227 6091
rect 3341 7087 3387 7098
rect 3341 6701 3387 6863
rect 3341 6315 3387 6477
rect 3341 5984 3387 6091
rect 3501 7087 3547 7144
rect 3501 6701 3547 6863
rect 3501 6315 3547 6477
rect 3501 6080 3547 6091
rect 3745 7087 3791 7328
rect 4033 7236 5039 7282
rect 3745 6701 3791 6863
rect 3745 6315 3791 6477
rect 3745 6080 3791 6091
rect 3905 7087 3951 7098
rect 3905 6701 3951 6863
rect 3905 6315 3951 6477
rect 3021 5938 3490 5984
rect 3698 5962 3774 5974
rect 3698 5959 3710 5962
rect 3021 5763 3067 5938
rect 3021 5127 3067 5289
rect 3021 4491 3067 4653
rect 3021 3960 3067 4017
rect 2381 3914 3067 3960
rect 3181 5763 3227 5774
rect 3181 5127 3227 5289
rect 3181 4491 3227 4653
rect 3181 3960 3227 4017
rect 3341 5763 3387 5938
rect 3657 5913 3710 5959
rect 3698 5910 3710 5913
rect 3762 5910 3774 5962
rect 3698 5898 3774 5910
rect 3905 5960 3951 6091
rect 4033 7087 4079 7236
rect 4993 7190 5039 7236
rect 4033 6701 4079 6863
rect 4033 6315 4079 6477
rect 4033 6034 4079 6091
rect 4193 7178 4894 7190
rect 4193 7144 4830 7178
rect 4193 7087 4239 7144
rect 4193 6701 4239 6863
rect 4193 6315 4239 6477
rect 4193 6080 4239 6091
rect 4353 7087 4399 7098
rect 4353 6701 4399 6863
rect 4353 6315 4399 6477
rect 4353 6034 4399 6091
rect 4513 7087 4559 7144
rect 4818 7126 4830 7144
rect 4882 7126 4894 7178
rect 4818 7114 4894 7126
rect 4993 7144 5359 7190
rect 4513 6701 4559 6863
rect 4513 6315 4559 6477
rect 4513 6080 4559 6091
rect 4673 7087 4719 7098
rect 4673 6701 4719 6863
rect 4673 6315 4719 6477
rect 4673 6034 4719 6091
rect 4033 5988 4719 6034
rect 3905 5949 3994 5960
rect 3905 5903 3937 5949
rect 3983 5903 3994 5949
rect 3905 5892 3994 5903
rect 3341 5127 3387 5289
rect 3341 4491 3387 4653
rect 3341 4006 3387 4017
rect 3501 5763 3655 5789
rect 3547 5743 3655 5763
rect 3745 5763 3791 5774
rect 3501 5127 3547 5289
rect 3501 4491 3547 4653
rect 3501 3960 3547 4017
rect 3181 3914 3547 3960
rect 3745 5127 3791 5289
rect 3745 4491 3791 4653
rect 2211 3886 2287 3898
rect 2211 3834 2223 3886
rect 2275 3868 2287 3886
rect 3181 3868 3227 3914
rect 2275 3834 3227 3868
rect 2211 3822 3227 3834
rect 3745 3776 3791 4017
rect 3905 5763 3951 5892
rect 4673 5866 4719 5988
rect 3905 5127 3951 5289
rect 3905 4491 3951 4653
rect 3905 4006 3951 4017
rect 4033 5820 4719 5866
rect 4033 5763 4079 5820
rect 4033 5127 4079 5289
rect 4033 4491 4079 4653
rect 4033 3898 4079 4017
rect 4193 5763 4239 5774
rect 4193 5127 4239 5289
rect 4193 4491 4239 4653
rect 4193 3960 4239 4017
rect 4353 5763 4399 5820
rect 4353 5127 4399 5289
rect 4353 4491 4399 4653
rect 4353 4006 4399 4017
rect 4513 5763 4559 5774
rect 4513 5127 4559 5289
rect 4513 4491 4559 4653
rect 4513 3960 4559 4017
rect 4673 5763 4719 5820
rect 4673 5127 4719 5289
rect 4673 4491 4719 4653
rect 4673 4006 4719 4017
rect 4833 7087 4879 7114
rect 4833 6701 4879 6863
rect 4833 6315 4879 6477
rect 4833 5984 4879 6091
rect 4993 7087 5039 7144
rect 4993 6701 5039 6863
rect 4993 6315 5039 6477
rect 4993 6080 5039 6091
rect 5153 7087 5199 7098
rect 5153 6701 5199 6863
rect 5153 6315 5199 6477
rect 5153 5984 5199 6091
rect 5313 7087 5359 7144
rect 5313 6701 5359 6863
rect 5313 6315 5359 6477
rect 5313 6080 5359 6091
rect 5557 7087 5603 7328
rect 5845 7236 6851 7282
rect 5557 6701 5603 6863
rect 5557 6315 5603 6477
rect 5557 6080 5603 6091
rect 5717 7087 5763 7098
rect 5717 6701 5763 6863
rect 5717 6315 5763 6477
rect 4833 5938 5302 5984
rect 5510 5962 5586 5974
rect 5510 5959 5522 5962
rect 4833 5763 4879 5938
rect 4833 5127 4879 5289
rect 4833 4491 4879 4653
rect 4833 3960 4879 4017
rect 4193 3914 4879 3960
rect 4993 5763 5039 5774
rect 4993 5127 5039 5289
rect 4993 4491 5039 4653
rect 4993 3960 5039 4017
rect 5153 5763 5199 5938
rect 5469 5913 5522 5959
rect 5510 5910 5522 5913
rect 5574 5910 5586 5962
rect 5510 5898 5586 5910
rect 5717 5960 5763 6091
rect 5845 7087 5891 7236
rect 6805 7190 6851 7236
rect 5845 6701 5891 6863
rect 5845 6315 5891 6477
rect 5845 6034 5891 6091
rect 6005 7178 6706 7190
rect 6005 7144 6642 7178
rect 6005 7087 6051 7144
rect 6005 6701 6051 6863
rect 6005 6315 6051 6477
rect 6005 6080 6051 6091
rect 6165 7087 6211 7098
rect 6165 6701 6211 6863
rect 6165 6315 6211 6477
rect 6165 6034 6211 6091
rect 6325 7087 6371 7144
rect 6630 7126 6642 7144
rect 6694 7126 6706 7178
rect 6630 7114 6706 7126
rect 6805 7144 7171 7190
rect 6325 6701 6371 6863
rect 6325 6315 6371 6477
rect 6325 6080 6371 6091
rect 6485 7087 6531 7098
rect 6485 6701 6531 6863
rect 6485 6315 6531 6477
rect 6485 6034 6531 6091
rect 5845 5988 6531 6034
rect 5717 5949 5806 5960
rect 5717 5903 5749 5949
rect 5795 5903 5806 5949
rect 5717 5892 5806 5903
rect 5153 5127 5199 5289
rect 5153 4491 5199 4653
rect 5153 4006 5199 4017
rect 5313 5763 5467 5789
rect 5359 5743 5467 5763
rect 5557 5763 5603 5774
rect 5313 5127 5359 5289
rect 5313 4491 5359 4653
rect 5313 3960 5359 4017
rect 4993 3914 5359 3960
rect 5557 5127 5603 5289
rect 5557 4491 5603 4653
rect 4023 3886 4099 3898
rect 4023 3834 4035 3886
rect 4087 3868 4099 3886
rect 4993 3868 5039 3914
rect 4087 3834 5039 3868
rect 4023 3822 5039 3834
rect 5557 3776 5603 4017
rect 5717 5763 5763 5892
rect 6485 5866 6531 5988
rect 5717 5127 5763 5289
rect 5717 4491 5763 4653
rect 5717 4006 5763 4017
rect 5845 5820 6531 5866
rect 5845 5763 5891 5820
rect 5845 5127 5891 5289
rect 5845 4491 5891 4653
rect 5845 3898 5891 4017
rect 6005 5763 6051 5774
rect 6005 5127 6051 5289
rect 6005 4491 6051 4653
rect 6005 3960 6051 4017
rect 6165 5763 6211 5820
rect 6165 5127 6211 5289
rect 6165 4491 6211 4653
rect 6165 4006 6211 4017
rect 6325 5763 6371 5774
rect 6325 5127 6371 5289
rect 6325 4491 6371 4653
rect 6325 3960 6371 4017
rect 6485 5763 6531 5820
rect 6485 5127 6531 5289
rect 6485 4491 6531 4653
rect 6485 4006 6531 4017
rect 6645 7087 6691 7114
rect 6645 6701 6691 6863
rect 6645 6315 6691 6477
rect 6645 5984 6691 6091
rect 6805 7087 6851 7144
rect 6805 6701 6851 6863
rect 6805 6315 6851 6477
rect 6805 6080 6851 6091
rect 6965 7087 7011 7098
rect 6965 6701 7011 6863
rect 6965 6315 7011 6477
rect 6965 5984 7011 6091
rect 7125 7087 7171 7144
rect 7125 6701 7171 6863
rect 7125 6315 7171 6477
rect 7125 6080 7171 6091
rect 7369 7087 7415 7328
rect 7657 7236 8663 7282
rect 7369 6701 7415 6863
rect 7369 6315 7415 6477
rect 7369 6080 7415 6091
rect 7529 7087 7575 7098
rect 7529 6701 7575 6863
rect 7529 6315 7575 6477
rect 6645 5938 7114 5984
rect 7322 5963 7398 5975
rect 7322 5959 7334 5963
rect 6645 5763 6691 5938
rect 6645 5127 6691 5289
rect 6645 4491 6691 4653
rect 6645 3960 6691 4017
rect 6005 3914 6691 3960
rect 6805 5763 6851 5774
rect 6805 5127 6851 5289
rect 6805 4491 6851 4653
rect 6805 3960 6851 4017
rect 6965 5763 7011 5938
rect 7281 5913 7334 5959
rect 7322 5911 7334 5913
rect 7386 5911 7398 5963
rect 7322 5899 7398 5911
rect 7529 5960 7575 6091
rect 7657 7087 7703 7236
rect 8617 7190 8663 7236
rect 8922 7193 8998 7205
rect 8922 7190 8934 7193
rect 7657 6701 7703 6863
rect 7657 6315 7703 6477
rect 7657 6034 7703 6091
rect 7817 7144 8503 7190
rect 7817 7087 7863 7144
rect 7817 6701 7863 6863
rect 7817 6315 7863 6477
rect 7817 6080 7863 6091
rect 7977 7087 8023 7098
rect 7977 6701 8023 6863
rect 7977 6315 8023 6477
rect 7977 6034 8023 6091
rect 8137 7087 8183 7144
rect 8137 6701 8183 6863
rect 8137 6315 8183 6477
rect 8137 6080 8183 6091
rect 8297 7087 8343 7098
rect 8297 6701 8343 6863
rect 8297 6315 8343 6477
rect 8297 6034 8343 6091
rect 7657 5988 8343 6034
rect 7529 5949 7618 5960
rect 7529 5903 7561 5949
rect 7607 5903 7618 5949
rect 7529 5892 7618 5903
rect 6965 5127 7011 5289
rect 6965 4491 7011 4653
rect 6965 4006 7011 4017
rect 7125 5763 7279 5789
rect 7171 5743 7279 5763
rect 7369 5763 7415 5774
rect 7125 5127 7171 5289
rect 7125 4491 7171 4653
rect 7125 3960 7171 4017
rect 6805 3914 7171 3960
rect 7369 5127 7415 5289
rect 7369 4491 7415 4653
rect 5835 3886 5911 3898
rect 5835 3834 5847 3886
rect 5899 3868 5911 3886
rect 6805 3868 6851 3914
rect 5899 3834 6851 3868
rect 5835 3822 6851 3834
rect 7369 3776 7415 4017
rect 7529 5763 7575 5892
rect 8297 5866 8343 5988
rect 7529 5127 7575 5289
rect 7529 4491 7575 4653
rect 7529 4006 7575 4017
rect 7657 5820 8343 5866
rect 7657 5763 7703 5820
rect 7657 5127 7703 5289
rect 7657 4491 7703 4653
rect 7657 3868 7703 4017
rect 7817 5763 7863 5774
rect 7817 5127 7863 5289
rect 7817 4491 7863 4653
rect 7817 3960 7863 4017
rect 7977 5763 8023 5820
rect 7977 5127 8023 5289
rect 7977 4491 8023 4653
rect 7977 4006 8023 4017
rect 8137 5763 8183 5774
rect 8137 5127 8183 5289
rect 8137 4491 8183 4653
rect 8137 3960 8183 4017
rect 8297 5763 8343 5820
rect 8297 5127 8343 5289
rect 8297 4491 8343 4653
rect 8297 4006 8343 4017
rect 8457 7087 8503 7144
rect 8457 6701 8503 6863
rect 8457 6315 8503 6477
rect 8457 5984 8503 6091
rect 8617 7144 8934 7190
rect 8617 7087 8663 7144
rect 8922 7141 8934 7144
rect 8986 7141 8998 7193
rect 8922 7129 8998 7141
rect 8617 6701 8663 6863
rect 8617 6315 8663 6477
rect 8617 6080 8663 6091
rect 8777 7087 8823 7098
rect 8777 6701 8823 6863
rect 8777 6315 8823 6477
rect 8777 5984 8823 6091
rect 8937 7087 8983 7129
rect 8937 6701 8983 6863
rect 8937 6315 8983 6477
rect 8937 6080 8983 6091
rect 8457 5938 8926 5984
rect 9086 5963 9162 5975
rect 8457 5763 8503 5938
rect 8457 5127 8503 5289
rect 8457 4491 8503 4653
rect 8457 3990 8503 4017
rect 8617 5763 8663 5774
rect 8617 5127 8663 5289
rect 8617 4491 8663 4653
rect 8442 3978 8518 3990
rect 8442 3960 8454 3978
rect 7817 3926 8454 3960
rect 8506 3926 8518 3978
rect 7817 3914 8518 3926
rect 8617 3960 8663 4017
rect 8777 5763 8823 5938
rect 9086 5911 9098 5963
rect 9150 5959 9162 5963
rect 9150 5913 9252 5959
rect 9150 5911 9162 5913
rect 9086 5899 9162 5911
rect 8777 5127 8823 5289
rect 8777 4491 8823 4653
rect 8777 4006 8823 4017
rect 8937 5763 9091 5789
rect 8983 5743 9091 5763
rect 8937 5127 8983 5289
rect 8937 4491 8983 4653
rect 8937 3960 8983 4017
rect 8617 3914 8983 3960
rect 9118 3978 9194 3990
rect 9118 3926 9130 3978
rect 9182 3975 9194 3978
rect 9182 3929 9282 3975
rect 9182 3926 9194 3929
rect 9118 3914 9194 3926
rect 8617 3868 8663 3914
rect 7657 3822 8663 3868
rect -4898 3746 9082 3776
rect -4898 3743 -4452 3746
rect -4400 3743 9082 3746
rect -4898 3697 -4860 3743
rect -4814 3697 -4766 3743
rect -4720 3697 -4672 3743
rect -4626 3697 -4578 3743
rect -4532 3697 -4452 3743
rect -4400 3697 -4355 3743
rect -4309 3697 -4261 3743
rect -4215 3697 -4167 3743
rect -4121 3697 -4073 3743
rect -4027 3697 -3979 3743
rect -3933 3697 -3885 3743
rect -3839 3697 -3791 3743
rect -3745 3697 -3697 3743
rect -3651 3697 -3569 3743
rect -3523 3697 -3475 3743
rect -3429 3697 -3381 3743
rect -3335 3697 -3287 3743
rect -3241 3697 -3193 3743
rect -3147 3697 -3099 3743
rect -3053 3697 -3005 3743
rect -2959 3697 -2911 3743
rect -2865 3697 -2783 3743
rect -2737 3697 -2689 3743
rect -2643 3697 -2595 3743
rect -2549 3697 -2501 3743
rect -2455 3697 -2407 3743
rect -2361 3697 -2313 3743
rect -2267 3697 -2219 3743
rect -2173 3697 -2125 3743
rect -2079 3697 -1997 3743
rect -1951 3697 -1903 3743
rect -1857 3697 -1809 3743
rect -1763 3697 -1715 3743
rect -1669 3697 -1621 3743
rect -1575 3697 -1527 3743
rect -1481 3697 -1433 3743
rect -1387 3697 -1339 3743
rect -1293 3697 -1211 3743
rect -1165 3697 -1117 3743
rect -1071 3697 -1023 3743
rect -977 3697 -929 3743
rect -883 3697 59 3743
rect 105 3697 153 3743
rect 199 3697 247 3743
rect 293 3697 341 3743
rect 387 3697 435 3743
rect 481 3697 529 3743
rect 575 3697 623 3743
rect 669 3697 717 3743
rect 763 3697 811 3743
rect 857 3697 905 3743
rect 951 3697 999 3743
rect 1045 3697 1093 3743
rect 1139 3697 1187 3743
rect 1233 3697 1281 3743
rect 1327 3697 1375 3743
rect 1421 3697 1469 3743
rect 1515 3697 1563 3743
rect 1609 3697 1657 3743
rect 1703 3697 1751 3743
rect 1797 3697 1871 3743
rect 1917 3697 1965 3743
rect 2011 3697 2059 3743
rect 2105 3697 2153 3743
rect 2199 3697 2247 3743
rect 2293 3697 2341 3743
rect 2387 3697 2435 3743
rect 2481 3697 2529 3743
rect 2575 3697 2623 3743
rect 2669 3697 2717 3743
rect 2763 3697 2811 3743
rect 2857 3697 2905 3743
rect 2951 3697 2999 3743
rect 3045 3697 3093 3743
rect 3139 3697 3187 3743
rect 3233 3697 3281 3743
rect 3327 3697 3375 3743
rect 3421 3697 3469 3743
rect 3515 3697 3563 3743
rect 3609 3697 3683 3743
rect 3729 3697 3777 3743
rect 3823 3697 3871 3743
rect 3917 3697 3965 3743
rect 4011 3697 4059 3743
rect 4105 3697 4153 3743
rect 4199 3697 4247 3743
rect 4293 3697 4341 3743
rect 4387 3697 4435 3743
rect 4481 3697 4529 3743
rect 4575 3697 4623 3743
rect 4669 3697 4717 3743
rect 4763 3697 4811 3743
rect 4857 3697 4905 3743
rect 4951 3697 4999 3743
rect 5045 3697 5093 3743
rect 5139 3697 5187 3743
rect 5233 3697 5281 3743
rect 5327 3697 5375 3743
rect 5421 3697 5495 3743
rect 5541 3697 5589 3743
rect 5635 3697 5683 3743
rect 5729 3697 5777 3743
rect 5823 3697 5871 3743
rect 5917 3697 5965 3743
rect 6011 3697 6059 3743
rect 6105 3697 6153 3743
rect 6199 3697 6247 3743
rect 6293 3697 6341 3743
rect 6387 3697 6435 3743
rect 6481 3697 6529 3743
rect 6575 3697 6623 3743
rect 6669 3697 6717 3743
rect 6763 3697 6811 3743
rect 6857 3697 6905 3743
rect 6951 3697 6999 3743
rect 7045 3697 7093 3743
rect 7139 3697 7187 3743
rect 7233 3697 7307 3743
rect 7353 3697 7401 3743
rect 7447 3697 7495 3743
rect 7541 3697 7589 3743
rect 7635 3697 7683 3743
rect 7729 3697 7777 3743
rect 7823 3697 7871 3743
rect 7917 3697 7965 3743
rect 8011 3697 8059 3743
rect 8105 3697 8153 3743
rect 8199 3697 8247 3743
rect 8293 3697 8341 3743
rect 8387 3697 8435 3743
rect 8481 3697 8529 3743
rect 8575 3697 8623 3743
rect 8669 3697 8717 3743
rect 8763 3697 8811 3743
rect 8857 3697 8905 3743
rect 8951 3697 8999 3743
rect 9045 3697 9082 3743
rect -4898 3694 -4452 3697
rect -4400 3694 9082 3697
rect -4898 3664 9082 3694
rect -4799 3560 -4753 3664
rect -4799 3375 -4753 3386
rect -4639 3560 -4593 3571
rect -4639 3329 -4593 3386
rect -4393 3515 -4347 3526
rect -4531 3329 -4485 3330
rect -4639 3283 -4485 3329
rect -4842 3202 -4774 3213
rect -5127 3156 -4831 3202
rect -4785 3156 -4774 3202
rect -4938 2600 -4892 3156
rect -4842 3145 -4774 3156
rect -4799 3088 -4753 3099
rect -4799 2921 -4753 3014
rect -4639 3088 -4593 3283
rect -4531 3176 -4485 3283
rect -4393 3284 -4347 3341
rect -4233 3515 -4187 3664
rect -4233 3330 -4187 3341
rect -4073 3572 -3707 3618
rect -4073 3515 -4027 3572
rect -4073 3284 -4027 3341
rect -4393 3238 -4027 3284
rect -3913 3515 -3867 3526
rect -3913 3284 -3867 3341
rect -3753 3515 -3707 3572
rect -3520 3526 -3474 3664
rect -3520 3453 -3474 3464
rect -2968 3526 -2922 3537
rect -3753 3330 -3707 3341
rect -3378 3284 -3308 3295
rect -3913 3238 -3365 3284
rect -3319 3238 -3308 3284
rect -4335 3176 -4267 3187
rect -3913 3179 -3867 3238
rect -3378 3231 -3308 3238
rect -3376 3227 -3308 3231
rect -2968 3284 -2922 3464
rect -2734 3526 -2688 3664
rect -2734 3453 -2688 3464
rect -2182 3526 -2136 3537
rect -2592 3284 -2522 3295
rect -2968 3238 -2579 3284
rect -2533 3238 -2522 3284
rect -4531 3130 -4324 3176
rect -4278 3130 -4267 3176
rect -4335 3119 -4267 3130
rect -4073 3133 -3867 3179
rect -3728 3148 -3660 3157
rect -4639 3003 -4593 3014
rect -4233 3076 -4187 3087
rect -4233 2921 -4187 3002
rect -4073 3076 -4027 3133
rect -3728 3096 -3720 3148
rect -3668 3146 -3660 3148
rect -3668 3099 -3590 3146
rect -3668 3096 -3660 3099
rect -3728 3088 -3660 3096
rect -4073 2991 -4027 3002
rect -3913 3076 -3867 3087
rect -2968 3036 -2922 3238
rect -2592 3231 -2522 3238
rect -2590 3227 -2522 3231
rect -2182 3284 -2136 3464
rect -1948 3526 -1902 3664
rect -1150 3560 -1104 3664
rect -1948 3453 -1902 3464
rect -1396 3526 -1350 3537
rect -1806 3284 -1736 3295
rect -2182 3238 -1793 3284
rect -1747 3238 -1736 3284
rect -2182 3036 -2136 3238
rect -1806 3231 -1736 3238
rect -1804 3227 -1736 3231
rect -1396 3284 -1350 3464
rect -1150 3375 -1104 3386
rect -990 3560 -944 3571
rect -990 3329 -944 3386
rect 121 3423 167 3664
rect 409 3572 1415 3618
rect -1396 3238 -1258 3284
rect -1396 3036 -1350 3238
rect -1304 3202 -1258 3238
rect -990 3283 -457 3329
rect -1193 3202 -1125 3213
rect -1304 3156 -1182 3202
rect -1136 3156 -1125 3202
rect -1193 3145 -1125 3156
rect -1150 3088 -1104 3099
rect -3913 2921 -3867 3002
rect -3539 2990 -3528 3036
rect -3482 2990 -3471 3036
rect -2979 2990 -2968 3036
rect -2922 2990 -2911 3036
rect -2753 2990 -2742 3036
rect -2696 2990 -2685 3036
rect -2193 2990 -2182 3036
rect -2136 2990 -2125 3036
rect -1967 2990 -1956 3036
rect -1910 2990 -1899 3036
rect -1407 2990 -1396 3036
rect -1350 2990 -1339 3036
rect -3528 2921 -3482 2990
rect -2742 2921 -2696 2990
rect -1956 2921 -1910 2990
rect -1150 2921 -1104 3014
rect -990 3088 -944 3283
rect -801 3148 -725 3160
rect -801 3096 -789 3148
rect -737 3096 -725 3148
rect -801 3084 -725 3096
rect -990 3003 -944 3014
rect -4846 2891 -897 2921
rect -4846 2888 -2749 2891
rect -2697 2888 -2185 2891
rect -2133 2888 -1682 2891
rect -1630 2888 -897 2891
rect -4846 2842 -4813 2888
rect -4767 2842 -4719 2888
rect -4673 2842 -4625 2888
rect -4579 2842 -4214 2888
rect -4168 2842 -4120 2888
rect -4074 2842 -4026 2888
rect -3980 2842 -3932 2888
rect -3886 2842 -3532 2888
rect -3486 2842 -3438 2888
rect -3392 2842 -3344 2888
rect -3298 2842 -3250 2888
rect -3204 2842 -3156 2888
rect -3110 2842 -3062 2888
rect -3016 2842 -2968 2888
rect -2922 2842 -2749 2888
rect -2697 2842 -2652 2888
rect -2606 2842 -2558 2888
rect -2512 2842 -2464 2888
rect -2418 2842 -2370 2888
rect -2324 2842 -2276 2888
rect -2230 2842 -2185 2888
rect -2133 2842 -1960 2888
rect -1914 2842 -1866 2888
rect -1820 2842 -1772 2888
rect -1726 2842 -1682 2888
rect -1630 2842 -1584 2888
rect -1538 2842 -1490 2888
rect -1444 2842 -1396 2888
rect -1350 2842 -1164 2888
rect -1118 2842 -1070 2888
rect -1024 2842 -976 2888
rect -930 2842 -897 2888
rect -4846 2839 -2749 2842
rect -2697 2839 -2185 2842
rect -2133 2839 -1682 2842
rect -1630 2839 -897 2842
rect -4846 2809 -897 2839
rect -4233 2728 -4187 2809
rect -4233 2643 -4187 2654
rect -4073 2728 -4027 2739
rect -4335 2600 -4267 2611
rect -4938 2554 -4324 2600
rect -4278 2554 -4267 2600
rect -4335 2543 -4267 2554
rect -4073 2597 -4027 2654
rect -3913 2728 -3867 2809
rect -3528 2740 -3482 2809
rect -2742 2740 -2696 2809
rect -1956 2740 -1910 2809
rect -3539 2694 -3528 2740
rect -3482 2694 -3471 2740
rect -2979 2694 -2968 2740
rect -2922 2694 -2911 2740
rect -2753 2694 -2742 2740
rect -2696 2694 -2685 2740
rect -2193 2694 -2182 2740
rect -2136 2694 -2125 2740
rect -1967 2694 -1956 2740
rect -1910 2694 -1899 2740
rect -1407 2694 -1396 2740
rect -1350 2694 -1339 2740
rect -1150 2716 -1104 2809
rect -3913 2643 -3867 2654
rect -3728 2633 -3660 2642
rect -4073 2551 -3867 2597
rect -3728 2581 -3720 2633
rect -3668 2631 -3660 2633
rect -3668 2584 -3590 2631
rect -3668 2581 -3660 2584
rect -3728 2573 -3660 2581
rect -3913 2492 -3867 2551
rect -3376 2499 -3308 2503
rect -3378 2492 -3308 2499
rect -4393 2446 -4027 2492
rect -4393 2389 -4347 2446
rect -4393 2204 -4347 2215
rect -4233 2389 -4187 2400
rect -4233 2066 -4187 2215
rect -4073 2389 -4027 2446
rect -4073 2158 -4027 2215
rect -3913 2446 -3365 2492
rect -3319 2446 -3308 2492
rect -3913 2389 -3867 2446
rect -3378 2435 -3308 2446
rect -2968 2492 -2922 2694
rect -2590 2499 -2522 2503
rect -2592 2492 -2522 2499
rect -2968 2446 -2579 2492
rect -2533 2446 -2522 2492
rect -3913 2204 -3867 2215
rect -3753 2389 -3707 2400
rect -3753 2158 -3707 2215
rect -4073 2112 -3707 2158
rect -3520 2266 -3474 2277
rect -3520 2066 -3474 2204
rect -2968 2266 -2922 2446
rect -2592 2435 -2522 2446
rect -2182 2492 -2136 2694
rect -1804 2499 -1736 2503
rect -1806 2492 -1736 2499
rect -2182 2446 -1793 2492
rect -1747 2446 -1736 2492
rect -2968 2193 -2922 2204
rect -2734 2266 -2688 2277
rect -2734 2066 -2688 2204
rect -2182 2266 -2136 2446
rect -1806 2435 -1736 2446
rect -1396 2492 -1350 2694
rect -1150 2631 -1104 2642
rect -990 2716 -944 2727
rect -1193 2574 -1125 2585
rect -1304 2528 -1182 2574
rect -1136 2528 -1125 2574
rect -1304 2492 -1258 2528
rect -1193 2517 -1125 2528
rect -1396 2446 -1258 2492
rect -990 2447 -944 2642
rect -786 2447 -740 3084
rect -679 2645 -633 3283
rect 121 2787 167 2949
rect -690 2633 -614 2645
rect -690 2581 -678 2633
rect -626 2630 -614 2633
rect -59 2633 17 2645
rect -59 2630 -47 2633
rect -626 2584 -47 2630
rect -626 2581 -614 2584
rect -690 2569 -614 2581
rect -59 2581 -47 2584
rect 5 2581 17 2633
rect -59 2569 17 2581
rect -181 2450 -105 2462
rect -181 2447 -169 2450
rect -2182 2193 -2136 2204
rect -1948 2266 -1902 2277
rect -1948 2066 -1902 2204
rect -1396 2266 -1350 2446
rect -990 2401 -169 2447
rect -1396 2193 -1350 2204
rect -1150 2344 -1104 2355
rect -1150 2066 -1104 2170
rect -990 2344 -944 2401
rect -181 2398 -169 2401
rect -117 2398 -105 2450
rect -181 2386 -105 2398
rect -990 2159 -944 2170
rect 121 2151 167 2313
rect -4492 2036 -845 2066
rect -4492 1984 -4452 2036
rect -4400 2033 -845 2036
rect -4400 1987 -4355 2033
rect -4309 1987 -4261 2033
rect -4215 1987 -4167 2033
rect -4121 1987 -4073 2033
rect -4027 1987 -3979 2033
rect -3933 1987 -3885 2033
rect -3839 1987 -3791 2033
rect -3745 1987 -3697 2033
rect -3651 1987 -3569 2033
rect -3523 1987 -3475 2033
rect -3429 1987 -3381 2033
rect -3335 1987 -3287 2033
rect -3241 1987 -3193 2033
rect -3147 1987 -3099 2033
rect -3053 1987 -3005 2033
rect -2959 1987 -2911 2033
rect -2865 1987 -2783 2033
rect -2737 1987 -2689 2033
rect -2643 1987 -2595 2033
rect -2549 1987 -2501 2033
rect -2455 1987 -2407 2033
rect -2361 1987 -2313 2033
rect -2267 1987 -2219 2033
rect -2173 1987 -2125 2033
rect -2079 1987 -1997 2033
rect -1951 1987 -1903 2033
rect -1857 1987 -1809 2033
rect -1763 1987 -1715 2033
rect -1669 1987 -1621 2033
rect -1575 1987 -1527 2033
rect -1481 1987 -1433 2033
rect -1387 1987 -1339 2033
rect -1293 1987 -1211 2033
rect -1165 1987 -1117 2033
rect -1071 1987 -1023 2033
rect -977 1987 -929 2033
rect -883 1987 -845 2033
rect -4400 1984 -845 1987
rect -4492 1954 -845 1984
rect -4393 1805 -4347 1816
rect -4393 1574 -4347 1631
rect -4233 1805 -4187 1954
rect -4233 1620 -4187 1631
rect -4073 1862 -3707 1908
rect -4073 1805 -4027 1862
rect -4073 1574 -4027 1631
rect -4393 1528 -4027 1574
rect -3913 1805 -3867 1816
rect -3913 1574 -3867 1631
rect -3753 1805 -3707 1862
rect -3520 1816 -3474 1954
rect -3520 1743 -3474 1754
rect -2968 1816 -2922 1827
rect -3753 1620 -3707 1631
rect -3378 1574 -3308 1585
rect -3913 1528 -3365 1574
rect -3319 1528 -3308 1574
rect -4335 1466 -4267 1477
rect -3913 1469 -3867 1528
rect -3378 1521 -3308 1528
rect -3376 1517 -3308 1521
rect -2968 1574 -2922 1754
rect -2734 1816 -2688 1954
rect -2734 1743 -2688 1754
rect -2182 1816 -2136 1827
rect -2592 1574 -2522 1585
rect -2968 1528 -2579 1574
rect -2533 1528 -2522 1574
rect -4938 1420 -4324 1466
rect -4278 1420 -4267 1466
rect -4938 864 -4892 1420
rect -4335 1409 -4267 1420
rect -4073 1423 -3867 1469
rect -3728 1439 -3660 1447
rect -4233 1366 -4187 1377
rect -4233 1211 -4187 1292
rect -4073 1366 -4027 1423
rect -3728 1387 -3720 1439
rect -3668 1436 -3660 1439
rect -3668 1389 -3590 1436
rect -3668 1387 -3660 1389
rect -3728 1378 -3660 1387
rect -4073 1281 -4027 1292
rect -3913 1366 -3867 1377
rect -2968 1326 -2922 1528
rect -2592 1521 -2522 1528
rect -2590 1517 -2522 1521
rect -2182 1574 -2136 1754
rect -1948 1816 -1902 1954
rect -1150 1850 -1104 1954
rect -1948 1743 -1902 1754
rect -1396 1816 -1350 1827
rect -1806 1574 -1736 1585
rect -2182 1528 -1793 1574
rect -1747 1528 -1736 1574
rect -2182 1326 -2136 1528
rect -1806 1521 -1736 1528
rect -1804 1517 -1736 1521
rect -1396 1574 -1350 1754
rect -1150 1665 -1104 1676
rect -990 1850 -944 1861
rect -990 1619 -944 1676
rect 121 1666 167 1677
rect 281 3423 327 3434
rect 281 2787 327 2949
rect 281 2151 327 2313
rect -303 1622 -227 1634
rect -303 1619 -291 1622
rect -1396 1528 -1258 1574
rect -1396 1326 -1350 1528
rect -1304 1492 -1258 1528
rect -990 1573 -291 1619
rect -1193 1492 -1125 1503
rect -1304 1446 -1182 1492
rect -1136 1446 -1125 1492
rect -1193 1435 -1125 1446
rect -1150 1378 -1104 1389
rect -3913 1211 -3867 1292
rect -3539 1280 -3528 1326
rect -3482 1280 -3471 1326
rect -2979 1280 -2968 1326
rect -2922 1280 -2911 1326
rect -2753 1280 -2742 1326
rect -2696 1280 -2685 1326
rect -2193 1280 -2182 1326
rect -2136 1280 -2125 1326
rect -1967 1280 -1956 1326
rect -1910 1280 -1899 1326
rect -1407 1280 -1396 1326
rect -1350 1280 -1339 1326
rect -3528 1211 -3482 1280
rect -2742 1211 -2696 1280
rect -1956 1211 -1910 1280
rect -1150 1211 -1104 1304
rect -990 1378 -944 1573
rect -990 1293 -944 1304
rect -4846 1181 -897 1211
rect -4846 1178 -2748 1181
rect -2696 1178 -2184 1181
rect -2132 1178 -1681 1181
rect -1629 1178 -897 1181
rect -4846 1132 -4813 1178
rect -4767 1132 -4719 1178
rect -4673 1132 -4625 1178
rect -4579 1132 -4214 1178
rect -4168 1132 -4120 1178
rect -4074 1132 -4026 1178
rect -3980 1132 -3932 1178
rect -3886 1132 -3532 1178
rect -3486 1132 -3438 1178
rect -3392 1132 -3344 1178
rect -3298 1132 -3250 1178
rect -3204 1132 -3156 1178
rect -3110 1132 -3062 1178
rect -3016 1132 -2968 1178
rect -2922 1132 -2748 1178
rect -2696 1132 -2652 1178
rect -2606 1132 -2558 1178
rect -2512 1132 -2464 1178
rect -2418 1132 -2370 1178
rect -2324 1132 -2276 1178
rect -2230 1132 -2184 1178
rect -2132 1132 -1960 1178
rect -1914 1132 -1866 1178
rect -1820 1132 -1772 1178
rect -1726 1132 -1681 1178
rect -1629 1132 -1584 1178
rect -1538 1132 -1490 1178
rect -1444 1132 -1396 1178
rect -1350 1132 -1164 1178
rect -1118 1132 -1070 1178
rect -1024 1132 -976 1178
rect -930 1132 -897 1178
rect -4846 1129 -2748 1132
rect -2696 1129 -2184 1132
rect -2132 1129 -1681 1132
rect -1629 1129 -897 1132
rect -4846 1099 -897 1129
rect -4799 1006 -4753 1099
rect -4233 1018 -4187 1099
rect -4799 921 -4753 932
rect -4639 1006 -4593 1017
rect -4233 933 -4187 944
rect -4073 1018 -4027 1029
rect -4842 864 -4774 875
rect -5127 818 -4831 864
rect -4785 818 -4774 864
rect -4842 807 -4774 818
rect -4639 737 -4593 932
rect -4335 890 -4267 901
rect -4531 844 -4324 890
rect -4278 844 -4267 890
rect -4531 737 -4485 844
rect -4335 833 -4267 844
rect -4073 887 -4027 944
rect -3913 1018 -3867 1099
rect -3528 1030 -3482 1099
rect -2742 1030 -2696 1099
rect -1956 1030 -1910 1099
rect -3539 984 -3528 1030
rect -3482 984 -3471 1030
rect -2979 984 -2968 1030
rect -2922 984 -2911 1030
rect -2753 984 -2742 1030
rect -2696 984 -2685 1030
rect -2193 984 -2182 1030
rect -2136 984 -2125 1030
rect -1967 984 -1956 1030
rect -1910 984 -1899 1030
rect -1407 984 -1396 1030
rect -1350 984 -1339 1030
rect -1150 1006 -1104 1099
rect -3913 933 -3867 944
rect -3728 924 -3660 932
rect -4073 841 -3867 887
rect -3728 872 -3720 924
rect -3668 921 -3660 924
rect -3668 874 -3590 921
rect -3668 872 -3660 874
rect -3728 863 -3660 872
rect -3913 782 -3867 841
rect -3376 789 -3308 793
rect -3378 782 -3308 789
rect -4639 691 -4485 737
rect -4799 634 -4753 645
rect -4799 356 -4753 460
rect -4639 634 -4593 691
rect -4531 690 -4485 691
rect -4393 736 -4027 782
rect -4393 679 -4347 736
rect -4393 494 -4347 505
rect -4233 679 -4187 690
rect -4639 449 -4593 460
rect -4233 356 -4187 505
rect -4073 679 -4027 736
rect -4073 448 -4027 505
rect -3913 736 -3365 782
rect -3319 736 -3308 782
rect -3913 679 -3867 736
rect -3378 725 -3308 736
rect -2968 782 -2922 984
rect -2590 789 -2522 793
rect -2592 782 -2522 789
rect -2968 736 -2579 782
rect -2533 736 -2522 782
rect -3913 494 -3867 505
rect -3753 679 -3707 690
rect -3753 448 -3707 505
rect -4073 402 -3707 448
rect -3520 556 -3474 567
rect -3520 356 -3474 494
rect -2968 556 -2922 736
rect -2592 725 -2522 736
rect -2182 782 -2136 984
rect -1804 789 -1736 793
rect -1806 782 -1736 789
rect -2182 736 -1793 782
rect -1747 736 -1736 782
rect -2968 483 -2922 494
rect -2734 556 -2688 567
rect -2734 356 -2688 494
rect -2182 556 -2136 736
rect -1806 725 -1736 736
rect -1396 782 -1350 984
rect -1150 921 -1104 932
rect -990 1006 -944 1017
rect -786 936 -740 1573
rect -303 1570 -291 1573
rect -239 1570 -227 1622
rect -303 1558 -227 1570
rect 281 1548 327 1677
rect 409 3423 455 3572
rect 1369 3526 1415 3572
rect 2253 3572 3259 3618
rect 2253 3526 2299 3572
rect 409 2787 455 2949
rect 409 2151 455 2313
rect 409 1620 455 1677
rect 569 3514 1270 3526
rect 569 3480 1206 3514
rect 569 3423 615 3480
rect 569 2787 615 2949
rect 569 2151 615 2313
rect 569 1666 615 1677
rect 729 3423 775 3434
rect 729 2787 775 2949
rect 729 2151 775 2313
rect 729 1620 775 1677
rect 889 3423 935 3480
rect 1194 3462 1206 3480
rect 1258 3462 1270 3514
rect 1194 3450 1270 3462
rect 1369 3480 1735 3526
rect 889 2787 935 2949
rect 889 2151 935 2313
rect 889 1666 935 1677
rect 1049 3423 1095 3434
rect 1049 2787 1095 2949
rect 1049 2151 1095 2313
rect 1049 1620 1095 1677
rect 409 1574 1095 1620
rect -59 1530 17 1542
rect -59 1478 -47 1530
rect 5 1527 17 1530
rect 78 1530 146 1538
rect 78 1527 86 1530
rect 5 1481 86 1527
rect 5 1478 17 1481
rect -59 1466 17 1478
rect 78 1478 86 1481
rect 138 1478 146 1530
rect 78 1470 146 1478
rect 281 1537 370 1548
rect 281 1491 313 1537
rect 359 1491 370 1537
rect 281 1480 370 1491
rect -690 1439 -614 1451
rect -690 1387 -678 1439
rect -626 1387 -614 1439
rect -690 1375 -614 1387
rect -1193 864 -1125 875
rect -1304 818 -1182 864
rect -1136 818 -1125 864
rect -1304 782 -1258 818
rect -1193 807 -1125 818
rect -1396 736 -1258 782
rect -990 737 -944 932
rect -801 924 -725 936
rect -801 872 -789 924
rect -737 872 -725 924
rect -801 860 -725 872
rect -679 737 -633 1375
rect 121 1349 167 1360
rect 121 963 167 1125
rect -425 740 -349 752
rect -425 737 -413 740
rect -2182 483 -2136 494
rect -1948 556 -1902 567
rect -1948 356 -1902 494
rect -1396 556 -1350 736
rect -990 691 -413 737
rect -1396 483 -1350 494
rect -1150 634 -1104 645
rect -1150 356 -1104 460
rect -990 634 -944 691
rect -425 688 -413 691
rect -361 688 -349 740
rect -425 676 -349 688
rect -990 449 -944 460
rect 121 577 167 739
rect -4898 326 -845 356
rect -4898 323 -4452 326
rect -4400 323 -845 326
rect -4898 277 -4860 323
rect -4814 277 -4766 323
rect -4720 277 -4672 323
rect -4626 277 -4578 323
rect -4532 277 -4452 323
rect -4400 277 -4355 323
rect -4309 277 -4261 323
rect -4215 277 -4167 323
rect -4121 277 -4073 323
rect -4027 277 -3979 323
rect -3933 277 -3885 323
rect -3839 277 -3791 323
rect -3745 277 -3697 323
rect -3651 277 -3569 323
rect -3523 277 -3475 323
rect -3429 277 -3381 323
rect -3335 277 -3287 323
rect -3241 277 -3193 323
rect -3147 277 -3099 323
rect -3053 277 -3005 323
rect -2959 277 -2911 323
rect -2865 277 -2783 323
rect -2737 277 -2689 323
rect -2643 277 -2595 323
rect -2549 277 -2501 323
rect -2455 277 -2407 323
rect -2361 277 -2313 323
rect -2267 277 -2219 323
rect -2173 277 -2125 323
rect -2079 277 -1997 323
rect -1951 277 -1903 323
rect -1857 277 -1809 323
rect -1763 277 -1715 323
rect -1669 277 -1621 323
rect -1575 277 -1527 323
rect -1481 277 -1433 323
rect -1387 277 -1339 323
rect -1293 277 -1211 323
rect -1165 277 -1117 323
rect -1071 277 -1023 323
rect -977 277 -929 323
rect -883 277 -845 323
rect -4898 274 -4452 277
rect -4400 274 -845 277
rect -4898 244 -845 274
rect -4799 140 -4753 244
rect -4799 -45 -4753 -34
rect -4639 140 -4593 151
rect -4639 -91 -4593 -34
rect -4393 95 -4347 106
rect -4531 -91 -4485 -90
rect -4639 -137 -4485 -91
rect -4842 -218 -4774 -207
rect -5126 -264 -4831 -218
rect -4785 -264 -4774 -218
rect -4938 -820 -4892 -264
rect -4842 -275 -4774 -264
rect -4799 -332 -4753 -321
rect -4799 -499 -4753 -406
rect -4639 -332 -4593 -137
rect -4531 -244 -4485 -137
rect -4393 -136 -4347 -79
rect -4233 95 -4187 244
rect -4233 -90 -4187 -79
rect -4073 152 -3707 198
rect -4073 95 -4027 152
rect -4073 -136 -4027 -79
rect -4393 -182 -4027 -136
rect -3913 95 -3867 106
rect -3913 -136 -3867 -79
rect -3753 95 -3707 152
rect -3520 106 -3474 244
rect -3520 33 -3474 44
rect -2968 106 -2922 117
rect -3753 -90 -3707 -79
rect -3378 -136 -3308 -125
rect -3913 -182 -3365 -136
rect -3319 -182 -3308 -136
rect -4335 -244 -4267 -233
rect -3913 -241 -3867 -182
rect -3378 -189 -3308 -182
rect -3376 -193 -3308 -189
rect -2968 -136 -2922 44
rect -2734 106 -2688 244
rect -2734 33 -2688 44
rect -2182 106 -2136 117
rect -2592 -136 -2522 -125
rect -2968 -182 -2579 -136
rect -2533 -182 -2522 -136
rect -4531 -290 -4324 -244
rect -4278 -290 -4267 -244
rect -4335 -301 -4267 -290
rect -4073 -287 -3867 -241
rect -3728 -272 -3660 -263
rect -4639 -417 -4593 -406
rect -4233 -344 -4187 -333
rect -4233 -499 -4187 -418
rect -4073 -344 -4027 -287
rect -3728 -324 -3720 -272
rect -3668 -274 -3660 -272
rect -3668 -321 -3590 -274
rect -3668 -324 -3660 -321
rect -3728 -332 -3660 -324
rect -4073 -429 -4027 -418
rect -3913 -344 -3867 -333
rect -2968 -384 -2922 -182
rect -2592 -189 -2522 -182
rect -2590 -193 -2522 -189
rect -2182 -136 -2136 44
rect -1948 106 -1902 244
rect -1150 140 -1104 244
rect -1948 33 -1902 44
rect -1396 106 -1350 117
rect -1806 -136 -1736 -125
rect -2182 -182 -1793 -136
rect -1747 -182 -1736 -136
rect -2182 -384 -2136 -182
rect -1806 -189 -1736 -182
rect -1804 -193 -1736 -189
rect -1396 -136 -1350 44
rect -1150 -45 -1104 -34
rect -990 140 -944 151
rect 121 112 167 353
rect 281 1349 327 1480
rect 1049 1452 1095 1574
rect 281 963 327 1125
rect 281 577 327 739
rect 281 342 327 353
rect 409 1406 1095 1452
rect 409 1349 455 1406
rect 409 963 455 1125
rect 409 577 455 739
rect 409 204 455 353
rect 569 1349 615 1360
rect 569 963 615 1125
rect 569 577 615 739
rect 569 296 615 353
rect 729 1349 775 1406
rect 729 963 775 1125
rect 729 577 775 739
rect 729 342 775 353
rect 889 1349 935 1360
rect 889 963 935 1125
rect 889 577 935 739
rect 889 296 935 353
rect 1049 1349 1095 1406
rect 1049 963 1095 1125
rect 1049 577 1095 739
rect 1049 342 1095 353
rect 1209 3423 1255 3450
rect 1209 2787 1255 2949
rect 1209 2151 1255 2313
rect 1209 1502 1255 1677
rect 1369 3423 1415 3480
rect 1369 2787 1415 2949
rect 1369 2151 1415 2313
rect 1369 1666 1415 1677
rect 1529 3423 1575 3434
rect 1529 2787 1575 2949
rect 1529 2151 1575 2313
rect 1529 1502 1575 1677
rect 1689 3423 1735 3480
rect 1689 2787 1735 2949
rect 1689 2151 1735 2313
rect 1933 3480 2299 3526
rect 1933 3423 1979 3480
rect 1933 2787 1979 2949
rect 1933 2151 1979 2313
rect 1735 1677 1933 1697
rect 1689 1671 1979 1677
rect 1674 1659 1979 1671
rect 1674 1607 1686 1659
rect 1738 1651 1979 1659
rect 2093 3423 2139 3434
rect 2093 2787 2139 2949
rect 2093 2151 2139 2313
rect 1738 1607 1750 1651
rect 1674 1595 1750 1607
rect 2093 1502 2139 1677
rect 2253 3423 2299 3480
rect 2398 3514 3099 3526
rect 2398 3462 2410 3514
rect 2462 3480 3099 3514
rect 2462 3462 2474 3480
rect 2398 3450 2474 3462
rect 2253 2787 2299 2949
rect 2253 2151 2299 2313
rect 2253 1666 2299 1677
rect 2413 3423 2459 3450
rect 2413 2787 2459 2949
rect 2413 2151 2459 2313
rect 2413 1502 2459 1677
rect 1209 1456 1678 1502
rect 1990 1456 2459 1502
rect 1209 1349 1255 1456
rect 1209 963 1255 1125
rect 1209 577 1255 739
rect 1209 296 1255 353
rect 569 250 1255 296
rect 1369 1349 1415 1360
rect 1369 963 1415 1125
rect 1369 577 1415 739
rect 1369 296 1415 353
rect 1529 1349 1575 1456
rect 1529 963 1575 1125
rect 1529 577 1575 739
rect 1529 342 1575 353
rect 1689 1349 1735 1360
rect 1689 963 1735 1125
rect 1689 577 1735 739
rect 1689 296 1735 353
rect 1369 250 1735 296
rect 1933 1349 1979 1360
rect 1933 963 1979 1125
rect 1933 577 1979 739
rect 1933 296 1979 353
rect 2093 1349 2139 1456
rect 2093 963 2139 1125
rect 2093 577 2139 739
rect 2093 342 2139 353
rect 2253 1349 2299 1360
rect 2253 963 2299 1125
rect 2253 577 2299 739
rect 2253 296 2299 353
rect 1933 250 2299 296
rect 2413 1349 2459 1456
rect 2413 963 2459 1125
rect 2413 577 2459 739
rect 2413 296 2459 353
rect 2573 3423 2619 3434
rect 2573 2787 2619 2949
rect 2573 2151 2619 2313
rect 2573 1620 2619 1677
rect 2733 3423 2779 3480
rect 2733 2787 2779 2949
rect 2733 2151 2779 2313
rect 2733 1666 2779 1677
rect 2893 3423 2939 3434
rect 2893 2787 2939 2949
rect 2893 2151 2939 2313
rect 2893 1620 2939 1677
rect 3053 3423 3099 3480
rect 3053 2787 3099 2949
rect 3053 2151 3099 2313
rect 3053 1666 3099 1677
rect 3213 3423 3259 3572
rect 3213 2787 3259 2949
rect 3213 2151 3259 2313
rect 3213 1620 3259 1677
rect 2573 1574 3259 1620
rect 3341 3423 3387 3434
rect 3341 2787 3387 2949
rect 3341 2151 3387 2313
rect 2573 1452 2619 1574
rect 3341 1548 3387 1677
rect 3501 3423 3547 3664
rect 3501 2787 3547 2949
rect 3501 2151 3547 2313
rect 3501 1666 3547 1677
rect 3745 3423 3791 3664
rect 4033 3572 5039 3618
rect 3745 2787 3791 2949
rect 3745 2151 3791 2313
rect 3745 1666 3791 1677
rect 3905 3423 3951 3434
rect 3905 2787 3951 2949
rect 3905 2151 3951 2313
rect 3298 1537 3387 1548
rect 3905 1548 3951 1677
rect 4033 3423 4079 3572
rect 4993 3526 5039 3572
rect 5877 3572 6883 3618
rect 5877 3526 5923 3572
rect 4178 3514 4879 3526
rect 4178 3462 4190 3514
rect 4242 3480 4879 3514
rect 4242 3462 4254 3480
rect 4178 3450 4254 3462
rect 4033 2787 4079 2949
rect 4033 2151 4079 2313
rect 4033 1620 4079 1677
rect 4193 3423 4239 3450
rect 4193 2787 4239 2949
rect 4193 2151 4239 2313
rect 4193 1666 4239 1677
rect 4353 3423 4399 3434
rect 4353 2787 4399 2949
rect 4353 2151 4399 2313
rect 4353 1620 4399 1677
rect 4513 3423 4559 3480
rect 4513 2787 4559 2949
rect 4513 2151 4559 2313
rect 4513 1666 4559 1677
rect 4673 3423 4719 3434
rect 4673 2787 4719 2949
rect 4673 2151 4719 2313
rect 4673 1620 4719 1677
rect 4033 1574 4719 1620
rect 3298 1491 3309 1537
rect 3355 1491 3387 1537
rect 3298 1480 3387 1491
rect 2573 1406 3259 1452
rect 2573 1349 2619 1406
rect 2573 963 2619 1125
rect 2573 577 2619 739
rect 2573 342 2619 353
rect 2733 1349 2779 1360
rect 2733 963 2779 1125
rect 2733 577 2779 739
rect 2733 296 2779 353
rect 2893 1349 2939 1406
rect 2893 963 2939 1125
rect 2893 577 2939 739
rect 2893 342 2939 353
rect 3053 1349 3099 1360
rect 3053 963 3099 1125
rect 3053 577 3099 739
rect 3053 296 3099 353
rect 2413 250 3099 296
rect 3213 1349 3259 1406
rect 3213 963 3259 1125
rect 3213 577 3259 739
rect 1369 204 1415 250
rect 409 158 1415 204
rect 2253 204 2299 250
rect 3213 204 3259 353
rect 3341 1349 3387 1480
rect 3522 1530 3590 1538
rect 3522 1478 3530 1530
rect 3582 1527 3590 1530
rect 3702 1527 3770 1538
rect 3582 1481 3713 1527
rect 3759 1481 3770 1527
rect 3582 1478 3590 1481
rect 3522 1470 3590 1478
rect 3702 1470 3770 1481
rect 3905 1537 3994 1548
rect 3905 1491 3937 1537
rect 3983 1491 3994 1537
rect 3905 1480 3994 1491
rect 3341 963 3387 1125
rect 3341 577 3387 739
rect 3341 342 3387 353
rect 3501 1349 3547 1360
rect 3501 963 3547 1125
rect 3501 577 3547 739
rect 2253 158 3259 204
rect 3501 112 3547 353
rect 3745 1349 3791 1360
rect 3745 963 3791 1125
rect 3745 577 3791 739
rect 3745 112 3791 353
rect 3905 1349 3951 1480
rect 4673 1452 4719 1574
rect 3905 963 3951 1125
rect 3905 577 3951 739
rect 3905 342 3951 353
rect 4033 1406 4719 1452
rect 4033 1349 4079 1406
rect 4033 963 4079 1125
rect 4033 577 4079 739
rect 4033 204 4079 353
rect 4193 1349 4239 1360
rect 4193 963 4239 1125
rect 4193 577 4239 739
rect 4193 296 4239 353
rect 4353 1349 4399 1406
rect 4353 963 4399 1125
rect 4353 577 4399 739
rect 4353 342 4399 353
rect 4513 1349 4559 1360
rect 4513 963 4559 1125
rect 4513 577 4559 739
rect 4513 296 4559 353
rect 4673 1349 4719 1406
rect 4673 963 4719 1125
rect 4673 577 4719 739
rect 4673 342 4719 353
rect 4833 3423 4879 3480
rect 4833 2787 4879 2949
rect 4833 2151 4879 2313
rect 4833 1502 4879 1677
rect 4993 3480 5359 3526
rect 4993 3423 5039 3480
rect 4993 2787 5039 2949
rect 4993 2151 5039 2313
rect 4993 1666 5039 1677
rect 5153 3423 5199 3434
rect 5153 2787 5199 2949
rect 5153 2151 5199 2313
rect 5153 1502 5199 1677
rect 5313 3423 5359 3480
rect 5313 2787 5359 2949
rect 5313 2151 5359 2313
rect 5557 3480 5923 3526
rect 5557 3423 5603 3480
rect 5557 2787 5603 2949
rect 5557 2151 5603 2313
rect 5359 1677 5557 1697
rect 5313 1651 5603 1677
rect 5717 3423 5763 3434
rect 5717 2787 5763 2949
rect 5717 2151 5763 2313
rect 5717 1502 5763 1677
rect 5877 3423 5923 3480
rect 6022 3514 6723 3526
rect 6022 3462 6034 3514
rect 6086 3480 6723 3514
rect 6086 3462 6098 3480
rect 6022 3450 6098 3462
rect 5877 2787 5923 2949
rect 5877 2151 5923 2313
rect 5877 1666 5923 1677
rect 6037 3423 6083 3450
rect 6037 2787 6083 2949
rect 6037 2151 6083 2313
rect 6037 1502 6083 1677
rect 4833 1456 5302 1502
rect 5614 1456 6083 1502
rect 4833 1349 4879 1456
rect 4833 963 4879 1125
rect 4833 577 4879 739
rect 4833 296 4879 353
rect 4193 250 4879 296
rect 4993 1349 5039 1360
rect 4993 963 5039 1125
rect 4993 577 5039 739
rect 4993 296 5039 353
rect 5153 1349 5199 1456
rect 5153 963 5199 1125
rect 5153 577 5199 739
rect 5153 342 5199 353
rect 5313 1349 5359 1360
rect 5313 963 5359 1125
rect 5313 577 5359 739
rect 5313 311 5359 353
rect 5557 1349 5603 1360
rect 5557 963 5603 1125
rect 5557 577 5603 739
rect 5298 299 5374 311
rect 5298 296 5310 299
rect 4993 250 5310 296
rect 4993 204 5039 250
rect 5298 247 5310 250
rect 5362 247 5374 299
rect 5557 296 5603 353
rect 5717 1349 5763 1456
rect 5717 963 5763 1125
rect 5717 577 5763 739
rect 5717 342 5763 353
rect 5877 1349 5923 1360
rect 5877 963 5923 1125
rect 5877 577 5923 739
rect 5877 296 5923 353
rect 5557 250 5923 296
rect 6037 1349 6083 1456
rect 6037 963 6083 1125
rect 6037 577 6083 739
rect 6037 296 6083 353
rect 6197 3423 6243 3434
rect 6197 2787 6243 2949
rect 6197 2151 6243 2313
rect 6197 1620 6243 1677
rect 6357 3423 6403 3480
rect 6357 2787 6403 2949
rect 6357 2151 6403 2313
rect 6357 1666 6403 1677
rect 6517 3423 6563 3434
rect 6517 2787 6563 2949
rect 6517 2151 6563 2313
rect 6517 1620 6563 1677
rect 6677 3423 6723 3480
rect 6677 2787 6723 2949
rect 6677 2151 6723 2313
rect 6677 1666 6723 1677
rect 6837 3423 6883 3572
rect 6837 2787 6883 2949
rect 6837 2151 6883 2313
rect 6837 1620 6883 1677
rect 6197 1574 6883 1620
rect 6965 3423 7011 3434
rect 6965 2787 7011 2949
rect 6965 2151 7011 2313
rect 6197 1452 6243 1574
rect 6965 1548 7011 1677
rect 7125 3423 7171 3664
rect 7689 3572 8695 3618
rect 7689 3526 7735 3572
rect 7349 3514 7735 3526
rect 7349 3462 7361 3514
rect 7413 3480 7735 3514
rect 7413 3462 7425 3480
rect 7349 3450 7425 3462
rect 7125 2787 7171 2949
rect 7125 2151 7171 2313
rect 7369 3423 7415 3450
rect 7369 2787 7415 2949
rect 7369 2151 7415 2313
rect 7125 1666 7171 1677
rect 7261 1677 7369 1697
rect 7261 1651 7415 1677
rect 7529 3423 7575 3434
rect 7529 2787 7575 2949
rect 7529 2151 7575 2313
rect 6922 1537 7011 1548
rect 6922 1491 6933 1537
rect 6979 1491 7011 1537
rect 6922 1480 7011 1491
rect 6197 1406 6883 1452
rect 6197 1349 6243 1406
rect 6197 963 6243 1125
rect 6197 577 6243 739
rect 6197 342 6243 353
rect 6357 1349 6403 1360
rect 6357 963 6403 1125
rect 6357 577 6403 739
rect 6357 296 6403 353
rect 6517 1349 6563 1406
rect 6517 963 6563 1125
rect 6517 577 6563 739
rect 6517 342 6563 353
rect 6677 1349 6723 1360
rect 6677 963 6723 1125
rect 6677 577 6723 739
rect 6677 296 6723 353
rect 6037 250 6723 296
rect 6837 1349 6883 1406
rect 6837 963 6883 1125
rect 6837 577 6883 739
rect 5298 235 5374 247
rect 4033 158 5039 204
rect 5877 204 5923 250
rect 6837 204 6883 353
rect 6965 1349 7011 1480
rect 7146 1530 7214 1538
rect 7146 1478 7154 1530
rect 7206 1527 7214 1530
rect 7206 1481 7259 1527
rect 7529 1502 7575 1677
rect 7689 3423 7735 3480
rect 7689 2787 7735 2949
rect 7689 2151 7735 2313
rect 7689 1666 7735 1677
rect 7849 3480 8535 3526
rect 7849 3423 7895 3480
rect 7849 2787 7895 2949
rect 7849 2151 7895 2313
rect 7849 1517 7895 1677
rect 8009 3423 8055 3434
rect 8009 2787 8055 2949
rect 8009 2151 8055 2313
rect 8009 1620 8055 1677
rect 8169 3423 8215 3480
rect 8169 2787 8215 2949
rect 8169 2151 8215 2313
rect 8169 1666 8215 1677
rect 8329 3423 8375 3434
rect 8329 2787 8375 2949
rect 8329 2151 8375 2313
rect 8329 1620 8375 1677
rect 8489 3423 8535 3480
rect 8489 2787 8535 2949
rect 8489 2151 8535 2313
rect 8489 1666 8535 1677
rect 8649 3423 8695 3572
rect 8649 2787 8695 2949
rect 8649 2151 8695 2313
rect 8649 1620 8695 1677
rect 8009 1574 8695 1620
rect 8777 3423 8823 3434
rect 8777 2787 8823 2949
rect 8777 2151 8823 2313
rect 7834 1505 7910 1517
rect 7834 1502 7846 1505
rect 7206 1478 7214 1481
rect 7146 1470 7214 1478
rect 7426 1456 7846 1502
rect 6965 963 7011 1125
rect 6965 577 7011 739
rect 6965 342 7011 353
rect 7125 1349 7171 1360
rect 7125 963 7171 1125
rect 7125 577 7171 739
rect 5877 158 6883 204
rect 7125 112 7171 353
rect 7369 1349 7415 1360
rect 7369 963 7415 1125
rect 7369 577 7415 739
rect 7369 296 7415 353
rect 7529 1349 7575 1456
rect 7834 1453 7846 1456
rect 7898 1453 7910 1505
rect 7834 1441 7910 1453
rect 8009 1452 8055 1574
rect 8777 1548 8823 1677
rect 8937 3423 8983 3664
rect 8937 2787 8983 2949
rect 8937 2151 8983 2313
rect 8937 1666 8983 1677
rect 8734 1537 8823 1548
rect 8734 1491 8745 1537
rect 8791 1491 8823 1537
rect 8734 1480 8823 1491
rect 7529 963 7575 1125
rect 7529 577 7575 739
rect 7529 342 7575 353
rect 7689 1349 7735 1360
rect 7689 963 7735 1125
rect 7689 577 7735 739
rect 7689 296 7735 353
rect 7369 250 7735 296
rect 7849 1349 7895 1441
rect 7849 963 7895 1125
rect 7849 577 7895 739
rect 7849 296 7895 353
rect 8009 1406 8695 1452
rect 8009 1349 8055 1406
rect 8009 963 8055 1125
rect 8009 577 8055 739
rect 8009 342 8055 353
rect 8169 1349 8215 1360
rect 8169 963 8215 1125
rect 8169 577 8215 739
rect 8169 296 8215 353
rect 8329 1349 8375 1406
rect 8329 963 8375 1125
rect 8329 577 8375 739
rect 8329 342 8375 353
rect 8489 1349 8535 1360
rect 8489 963 8535 1125
rect 8489 577 8535 739
rect 8489 296 8535 353
rect 7849 250 8535 296
rect 8649 1349 8695 1406
rect 8649 963 8695 1125
rect 8649 577 8695 739
rect 7689 204 7735 250
rect 8649 204 8695 353
rect 8777 1349 8823 1480
rect 8958 1530 9026 1538
rect 8958 1478 8966 1530
rect 9018 1527 9026 1530
rect 9018 1481 9071 1527
rect 9118 1505 9194 1517
rect 9018 1478 9026 1481
rect 8958 1470 9026 1478
rect 9118 1453 9130 1505
rect 9182 1502 9194 1505
rect 9182 1456 9282 1502
rect 9182 1453 9194 1456
rect 9118 1441 9194 1453
rect 8777 963 8823 1125
rect 8777 577 8823 739
rect 8777 342 8823 353
rect 8937 1349 8983 1360
rect 8937 963 8983 1125
rect 8937 577 8983 739
rect 7689 158 8695 204
rect 8937 112 8983 353
rect 84 82 9020 112
rect 84 79 855 82
rect 907 79 8197 82
rect 8249 79 9020 82
rect 84 33 106 79
rect 152 33 200 79
rect 246 33 294 79
rect 340 33 388 79
rect 434 33 482 79
rect 528 33 576 79
rect 622 33 670 79
rect 716 33 764 79
rect 810 33 855 79
rect 907 33 952 79
rect 998 33 1046 79
rect 1092 33 1140 79
rect 1186 33 1234 79
rect 1280 33 1328 79
rect 1374 33 1422 79
rect 1468 33 1516 79
rect 1562 33 1610 79
rect 1656 33 1704 79
rect 1750 33 1918 79
rect 1964 33 2012 79
rect 2058 33 2106 79
rect 2152 33 2200 79
rect 2246 33 2294 79
rect 2340 33 2388 79
rect 2434 33 2482 79
rect 2528 33 2576 79
rect 2622 33 2670 79
rect 2716 33 2764 79
rect 2810 33 2858 79
rect 2904 33 2952 79
rect 2998 33 3046 79
rect 3092 33 3140 79
rect 3186 33 3234 79
rect 3280 33 3328 79
rect 3374 33 3422 79
rect 3468 33 3516 79
rect 3562 33 3730 79
rect 3776 33 3824 79
rect 3870 33 3918 79
rect 3964 33 4012 79
rect 4058 33 4106 79
rect 4152 33 4200 79
rect 4246 33 4294 79
rect 4340 33 4388 79
rect 4434 33 4482 79
rect 4528 33 4576 79
rect 4622 33 4670 79
rect 4716 33 4764 79
rect 4810 33 4858 79
rect 4904 33 4952 79
rect 4998 33 5046 79
rect 5092 33 5140 79
rect 5186 33 5234 79
rect 5280 33 5328 79
rect 5374 33 5542 79
rect 5588 33 5636 79
rect 5682 33 5730 79
rect 5776 33 5824 79
rect 5870 33 5918 79
rect 5964 33 6012 79
rect 6058 33 6106 79
rect 6152 33 6200 79
rect 6246 33 6294 79
rect 6340 33 6388 79
rect 6434 33 6482 79
rect 6528 33 6576 79
rect 6622 33 6670 79
rect 6716 33 6764 79
rect 6810 33 6858 79
rect 6904 33 6952 79
rect 6998 33 7046 79
rect 7092 33 7140 79
rect 7186 33 7354 79
rect 7400 33 7448 79
rect 7494 33 7542 79
rect 7588 33 7636 79
rect 7682 33 7730 79
rect 7776 33 7824 79
rect 7870 33 7918 79
rect 7964 33 8012 79
rect 8058 33 8106 79
rect 8152 33 8197 79
rect 8249 33 8294 79
rect 8340 33 8388 79
rect 8434 33 8482 79
rect 8528 33 8576 79
rect 8622 33 8670 79
rect 8716 33 8764 79
rect 8810 33 8858 79
rect 8904 33 8952 79
rect 8998 33 9020 79
rect 84 30 855 33
rect 907 30 8197 33
rect 8249 30 9020 33
rect 84 0 9020 30
rect -990 -91 -944 -34
rect -1396 -182 -1258 -136
rect -1396 -384 -1350 -182
rect -1304 -218 -1258 -182
rect -990 -137 -457 -91
rect -1193 -218 -1125 -207
rect -1304 -264 -1182 -218
rect -1136 -264 -1125 -218
rect -1193 -275 -1125 -264
rect -1150 -332 -1104 -321
rect -3913 -499 -3867 -418
rect -3539 -430 -3528 -384
rect -3482 -430 -3471 -384
rect -2979 -430 -2968 -384
rect -2922 -430 -2911 -384
rect -2753 -430 -2742 -384
rect -2696 -430 -2685 -384
rect -2193 -430 -2182 -384
rect -2136 -430 -2125 -384
rect -1967 -430 -1956 -384
rect -1910 -430 -1899 -384
rect -1407 -430 -1396 -384
rect -1350 -430 -1339 -384
rect -3528 -499 -3482 -430
rect -2742 -499 -2696 -430
rect -1956 -499 -1910 -430
rect -1150 -499 -1104 -406
rect -990 -332 -944 -137
rect -801 -272 -725 -260
rect -801 -324 -789 -272
rect -737 -324 -725 -272
rect -801 -336 -725 -324
rect -990 -417 -944 -406
rect -4846 -529 -897 -499
rect -4846 -532 -2748 -529
rect -2696 -532 -2184 -529
rect -2132 -532 -1681 -529
rect -1629 -532 -897 -529
rect -4846 -578 -4813 -532
rect -4767 -578 -4719 -532
rect -4673 -578 -4625 -532
rect -4579 -578 -4214 -532
rect -4168 -578 -4120 -532
rect -4074 -578 -4026 -532
rect -3980 -578 -3932 -532
rect -3886 -578 -3532 -532
rect -3486 -578 -3438 -532
rect -3392 -578 -3344 -532
rect -3298 -578 -3250 -532
rect -3204 -578 -3156 -532
rect -3110 -578 -3062 -532
rect -3016 -578 -2968 -532
rect -2922 -578 -2748 -532
rect -2696 -578 -2652 -532
rect -2606 -578 -2558 -532
rect -2512 -578 -2464 -532
rect -2418 -578 -2370 -532
rect -2324 -578 -2276 -532
rect -2230 -578 -2184 -532
rect -2132 -578 -1960 -532
rect -1914 -578 -1866 -532
rect -1820 -578 -1772 -532
rect -1726 -578 -1681 -532
rect -1629 -578 -1584 -532
rect -1538 -578 -1490 -532
rect -1444 -578 -1396 -532
rect -1350 -578 -1164 -532
rect -1118 -578 -1070 -532
rect -1024 -578 -976 -532
rect -930 -578 -897 -532
rect -4846 -581 -2748 -578
rect -2696 -581 -2184 -578
rect -2132 -581 -1681 -578
rect -1629 -581 -897 -578
rect -4846 -611 -897 -581
rect -4233 -692 -4187 -611
rect -4233 -777 -4187 -766
rect -4073 -692 -4027 -681
rect -4335 -820 -4267 -809
rect -4938 -866 -4324 -820
rect -4278 -866 -4267 -820
rect -4335 -877 -4267 -866
rect -4073 -823 -4027 -766
rect -3913 -692 -3867 -611
rect -3528 -680 -3482 -611
rect -2742 -680 -2696 -611
rect -1956 -680 -1910 -611
rect -3539 -726 -3528 -680
rect -3482 -726 -3471 -680
rect -2979 -726 -2968 -680
rect -2922 -726 -2911 -680
rect -2753 -726 -2742 -680
rect -2696 -726 -2685 -680
rect -2193 -726 -2182 -680
rect -2136 -726 -2125 -680
rect -1967 -726 -1956 -680
rect -1910 -726 -1899 -680
rect -1407 -726 -1396 -680
rect -1350 -726 -1339 -680
rect -1150 -704 -1104 -611
rect -3913 -777 -3867 -766
rect -3728 -787 -3660 -778
rect -4073 -869 -3867 -823
rect -3728 -839 -3720 -787
rect -3668 -789 -3660 -787
rect -3668 -836 -3590 -789
rect -3668 -839 -3660 -836
rect -3728 -847 -3660 -839
rect -3913 -928 -3867 -869
rect -3376 -921 -3308 -917
rect -3378 -928 -3308 -921
rect -4393 -974 -4027 -928
rect -4393 -1031 -4347 -974
rect -4393 -1216 -4347 -1205
rect -4233 -1031 -4187 -1020
rect -4233 -1354 -4187 -1205
rect -4073 -1031 -4027 -974
rect -4073 -1262 -4027 -1205
rect -3913 -974 -3365 -928
rect -3319 -974 -3308 -928
rect -3913 -1031 -3867 -974
rect -3378 -985 -3308 -974
rect -2968 -928 -2922 -726
rect -2590 -921 -2522 -917
rect -2592 -928 -2522 -921
rect -2968 -974 -2579 -928
rect -2533 -974 -2522 -928
rect -3913 -1216 -3867 -1205
rect -3753 -1031 -3707 -1020
rect -3753 -1262 -3707 -1205
rect -4073 -1308 -3707 -1262
rect -3520 -1154 -3474 -1143
rect -3520 -1354 -3474 -1216
rect -2968 -1154 -2922 -974
rect -2592 -985 -2522 -974
rect -2182 -928 -2136 -726
rect -1804 -921 -1736 -917
rect -1806 -928 -1736 -921
rect -2182 -974 -1793 -928
rect -1747 -974 -1736 -928
rect -2968 -1227 -2922 -1216
rect -2734 -1154 -2688 -1143
rect -2734 -1354 -2688 -1216
rect -2182 -1154 -2136 -974
rect -1806 -985 -1736 -974
rect -1396 -928 -1350 -726
rect -1150 -789 -1104 -778
rect -990 -704 -944 -693
rect -1193 -846 -1125 -835
rect -1304 -892 -1182 -846
rect -1136 -892 -1125 -846
rect -1304 -928 -1258 -892
rect -1193 -903 -1125 -892
rect -1396 -974 -1258 -928
rect -990 -973 -944 -778
rect -786 -973 -740 -336
rect -679 -775 -633 -137
rect 121 -241 167 0
rect 409 -92 1415 -46
rect 121 -627 167 -465
rect -690 -787 -614 -775
rect -690 -839 -678 -787
rect -626 -839 -614 -787
rect -690 -851 -614 -839
rect -547 -970 -471 -958
rect -547 -973 -535 -970
rect -2182 -1227 -2136 -1216
rect -1948 -1154 -1902 -1143
rect -1948 -1354 -1902 -1216
rect -1396 -1154 -1350 -974
rect -990 -1019 -535 -973
rect -1396 -1227 -1350 -1216
rect -1150 -1076 -1104 -1065
rect -1150 -1354 -1104 -1250
rect -990 -1076 -944 -1019
rect -547 -1022 -535 -1019
rect -483 -1022 -471 -970
rect -547 -1034 -471 -1022
rect 121 -1013 167 -851
rect 121 -1248 167 -1237
rect 281 -241 327 -230
rect 281 -627 327 -465
rect 281 -1013 327 -851
rect -990 -1261 -944 -1250
rect -4492 -1384 -845 -1354
rect 78 -1366 146 -1358
rect 78 -1369 86 -1366
rect -4492 -1436 -4452 -1384
rect -4400 -1387 -3953 -1384
rect -3901 -1387 -3653 -1384
rect -3601 -1387 -3353 -1384
rect -3301 -1387 -3053 -1384
rect -3001 -1387 -2753 -1384
rect -2701 -1387 -845 -1384
rect -4400 -1433 -4355 -1387
rect -4309 -1433 -4261 -1387
rect -4215 -1433 -4167 -1387
rect -4121 -1433 -4073 -1387
rect -4027 -1433 -3979 -1387
rect -3901 -1433 -3885 -1387
rect -3839 -1433 -3791 -1387
rect -3745 -1433 -3697 -1387
rect -3601 -1433 -3569 -1387
rect -3523 -1433 -3475 -1387
rect -3429 -1433 -3381 -1387
rect -3301 -1433 -3287 -1387
rect -3241 -1433 -3193 -1387
rect -3147 -1433 -3099 -1387
rect -2959 -1433 -2911 -1387
rect -2865 -1433 -2783 -1387
rect -2701 -1433 -2689 -1387
rect -2643 -1433 -2595 -1387
rect -2549 -1433 -2501 -1387
rect -2455 -1433 -2407 -1387
rect -2361 -1433 -2313 -1387
rect -2267 -1433 -2219 -1387
rect -2173 -1433 -2125 -1387
rect -2079 -1433 -1997 -1387
rect -1951 -1433 -1903 -1387
rect -1857 -1433 -1809 -1387
rect -1763 -1433 -1715 -1387
rect -1669 -1433 -1621 -1387
rect -1575 -1433 -1527 -1387
rect -1481 -1433 -1433 -1387
rect -1387 -1433 -1339 -1387
rect -1293 -1433 -1211 -1387
rect -1165 -1433 -1117 -1387
rect -1071 -1433 -1023 -1387
rect -977 -1433 -929 -1387
rect -883 -1433 -845 -1387
rect 33 -1415 86 -1369
rect 78 -1418 86 -1415
rect 138 -1418 146 -1366
rect 78 -1426 146 -1418
rect 281 -1368 327 -1237
rect 409 -241 455 -92
rect 1369 -138 1415 -92
rect 2253 -92 3259 -46
rect 2253 -138 2299 -92
rect 554 -150 1255 -138
rect 554 -202 566 -150
rect 618 -184 1255 -150
rect 618 -202 630 -184
rect 554 -214 630 -202
rect 409 -627 455 -465
rect 409 -1013 455 -851
rect 409 -1294 455 -1237
rect 569 -241 615 -214
rect 569 -627 615 -465
rect 569 -1013 615 -851
rect 569 -1248 615 -1237
rect 729 -241 775 -230
rect 729 -627 775 -465
rect 729 -1013 775 -851
rect 729 -1294 775 -1237
rect 889 -241 935 -184
rect 889 -627 935 -465
rect 889 -1013 935 -851
rect 889 -1248 935 -1237
rect 1049 -241 1095 -230
rect 1049 -627 1095 -465
rect 1049 -1013 1095 -851
rect 1049 -1294 1095 -1237
rect 409 -1340 1095 -1294
rect 281 -1379 370 -1368
rect 281 -1425 313 -1379
rect 359 -1425 370 -1379
rect -4400 -1436 -3953 -1433
rect -3901 -1436 -3653 -1433
rect -3601 -1436 -3353 -1433
rect -3301 -1436 -3053 -1433
rect -3001 -1436 -2753 -1433
rect -2701 -1436 -845 -1433
rect -4492 -1466 -845 -1436
rect 281 -1436 370 -1425
rect 121 -1565 167 -1554
rect 121 -2201 167 -2039
rect 121 -2837 167 -2675
rect 121 -3552 167 -3311
rect 281 -1565 327 -1436
rect 1049 -1462 1095 -1340
rect 281 -2201 327 -2039
rect 281 -2837 327 -2675
rect 281 -3322 327 -3311
rect 409 -1508 1095 -1462
rect 409 -1565 455 -1508
rect 409 -2201 455 -2039
rect 409 -2837 455 -2675
rect 409 -3460 455 -3311
rect 569 -1565 615 -1554
rect 569 -2201 615 -2039
rect 569 -2837 615 -2675
rect 569 -3368 615 -3311
rect 729 -1565 775 -1508
rect 729 -2201 775 -2039
rect 729 -2837 775 -2675
rect 729 -3322 775 -3311
rect 889 -1565 935 -1554
rect 889 -2201 935 -2039
rect 889 -2837 935 -2675
rect 889 -3368 935 -3311
rect 1049 -1565 1095 -1508
rect 1049 -2201 1095 -2039
rect 1049 -2837 1095 -2675
rect 1049 -3322 1095 -3311
rect 1209 -241 1255 -184
rect 1209 -627 1255 -465
rect 1209 -1013 1255 -851
rect 1209 -1344 1255 -1237
rect 1369 -184 1735 -138
rect 1369 -241 1415 -184
rect 1369 -627 1415 -465
rect 1369 -1013 1415 -851
rect 1369 -1248 1415 -1237
rect 1529 -241 1575 -230
rect 1529 -627 1575 -465
rect 1529 -1013 1575 -851
rect 1529 -1344 1575 -1237
rect 1689 -241 1735 -184
rect 1689 -627 1735 -465
rect 1689 -1013 1735 -851
rect 1689 -1248 1735 -1237
rect 1933 -184 2299 -138
rect 1933 -241 1979 -184
rect 1933 -627 1979 -465
rect 1933 -1013 1979 -851
rect 1933 -1248 1979 -1237
rect 2093 -241 2139 -230
rect 2093 -627 2139 -465
rect 2093 -1013 2139 -851
rect 2093 -1344 2139 -1237
rect 2253 -241 2299 -184
rect 2253 -627 2299 -465
rect 2253 -1013 2299 -851
rect 2253 -1248 2299 -1237
rect 2413 -150 3114 -138
rect 2413 -184 3050 -150
rect 2413 -241 2459 -184
rect 2413 -627 2459 -465
rect 2413 -1013 2459 -851
rect 2413 -1344 2459 -1237
rect 1209 -1390 1678 -1344
rect 1990 -1390 2459 -1344
rect 1209 -1565 1255 -1390
rect 1209 -2201 1255 -2039
rect 1209 -2837 1255 -2675
rect 1209 -3368 1255 -3311
rect 569 -3414 1255 -3368
rect 1369 -1565 1415 -1554
rect 1369 -2201 1415 -2039
rect 1369 -2837 1415 -2675
rect 1369 -3368 1415 -3311
rect 1529 -1565 1575 -1390
rect 1529 -2201 1575 -2039
rect 1529 -2837 1575 -2675
rect 1529 -3322 1575 -3311
rect 1689 -1565 1979 -1539
rect 1735 -1585 1933 -1565
rect 1689 -2201 1735 -2039
rect 1689 -2837 1735 -2675
rect 1689 -3368 1735 -3311
rect 1933 -2201 1979 -2039
rect 1933 -2837 1979 -2675
rect 1933 -3353 1979 -3311
rect 2093 -1565 2139 -1390
rect 2093 -2201 2139 -2039
rect 2093 -2837 2139 -2675
rect 2093 -3322 2139 -3311
rect 2253 -1565 2299 -1554
rect 2253 -2201 2299 -2039
rect 2253 -2837 2299 -2675
rect 1369 -3414 1735 -3368
rect 1918 -3365 1994 -3353
rect 1369 -3460 1415 -3414
rect 1918 -3417 1930 -3365
rect 1982 -3368 1994 -3365
rect 2253 -3368 2299 -3311
rect 1982 -3414 2299 -3368
rect 2413 -1565 2459 -1390
rect 2413 -2201 2459 -2039
rect 2413 -2837 2459 -2675
rect 2413 -3368 2459 -3311
rect 2573 -241 2619 -230
rect 2573 -627 2619 -465
rect 2573 -1013 2619 -851
rect 2573 -1294 2619 -1237
rect 2733 -241 2779 -184
rect 3038 -202 3050 -184
rect 3102 -202 3114 -150
rect 3038 -214 3114 -202
rect 2733 -627 2779 -465
rect 2733 -1013 2779 -851
rect 2733 -1248 2779 -1237
rect 2893 -241 2939 -230
rect 2893 -627 2939 -465
rect 2893 -1013 2939 -851
rect 2893 -1294 2939 -1237
rect 3053 -241 3099 -214
rect 3053 -627 3099 -465
rect 3053 -1013 3099 -851
rect 3053 -1248 3099 -1237
rect 3213 -241 3259 -92
rect 3213 -627 3259 -465
rect 3213 -1013 3259 -851
rect 3213 -1294 3259 -1237
rect 2573 -1340 3259 -1294
rect 3341 -241 3387 -230
rect 3341 -627 3387 -465
rect 3341 -1013 3387 -851
rect 2573 -1462 2619 -1340
rect 3341 -1368 3387 -1237
rect 3501 -241 3547 0
rect 3501 -627 3547 -465
rect 3501 -1013 3547 -851
rect 3501 -1248 3547 -1237
rect 3745 -241 3791 0
rect 4033 -92 5039 -46
rect 3745 -627 3791 -465
rect 3745 -1013 3791 -851
rect 3745 -1248 3791 -1237
rect 3905 -241 3951 -230
rect 3905 -627 3951 -465
rect 3905 -1013 3951 -851
rect 3298 -1379 3387 -1368
rect 3298 -1425 3309 -1379
rect 3355 -1425 3387 -1379
rect 3298 -1436 3387 -1425
rect 3522 -1366 3590 -1358
rect 3522 -1418 3530 -1366
rect 3582 -1369 3590 -1366
rect 3702 -1369 3770 -1358
rect 3582 -1415 3713 -1369
rect 3759 -1415 3770 -1369
rect 3582 -1418 3590 -1415
rect 3522 -1426 3590 -1418
rect 3702 -1426 3770 -1415
rect 3905 -1368 3951 -1237
rect 4033 -241 4079 -92
rect 4993 -138 5039 -92
rect 5877 -92 6883 -46
rect 5877 -138 5923 -92
rect 4033 -627 4079 -465
rect 4033 -1013 4079 -851
rect 4033 -1294 4079 -1237
rect 4193 -150 4894 -138
rect 4193 -184 4830 -150
rect 4193 -241 4239 -184
rect 4193 -627 4239 -465
rect 4193 -1013 4239 -851
rect 4193 -1248 4239 -1237
rect 4353 -241 4399 -230
rect 4353 -627 4399 -465
rect 4353 -1013 4399 -851
rect 4353 -1294 4399 -1237
rect 4513 -241 4559 -184
rect 4818 -202 4830 -184
rect 4882 -202 4894 -150
rect 4818 -214 4894 -202
rect 4993 -184 5359 -138
rect 4513 -627 4559 -465
rect 4513 -1013 4559 -851
rect 4513 -1248 4559 -1237
rect 4673 -241 4719 -230
rect 4673 -627 4719 -465
rect 4673 -1013 4719 -851
rect 4673 -1294 4719 -1237
rect 4033 -1340 4719 -1294
rect 3905 -1379 3994 -1368
rect 3905 -1425 3937 -1379
rect 3983 -1425 3994 -1379
rect 2573 -1508 3259 -1462
rect 2573 -1565 2619 -1508
rect 2573 -2201 2619 -2039
rect 2573 -2837 2619 -2675
rect 2573 -3322 2619 -3311
rect 2733 -1565 2779 -1554
rect 2733 -2201 2779 -2039
rect 2733 -2837 2779 -2675
rect 2733 -3368 2779 -3311
rect 2893 -1565 2939 -1508
rect 2893 -2201 2939 -2039
rect 2893 -2837 2939 -2675
rect 2893 -3322 2939 -3311
rect 3053 -1565 3099 -1554
rect 3053 -2201 3099 -2039
rect 3053 -2837 3099 -2675
rect 3053 -3368 3099 -3311
rect 2413 -3414 3099 -3368
rect 3213 -1565 3259 -1508
rect 3213 -2201 3259 -2039
rect 3213 -2837 3259 -2675
rect 1982 -3417 1994 -3414
rect 1918 -3429 1994 -3417
rect 409 -3506 1415 -3460
rect 2253 -3460 2299 -3414
rect 3213 -3460 3259 -3311
rect 3341 -1565 3387 -1436
rect 3905 -1436 3994 -1425
rect 3341 -2201 3387 -2039
rect 3341 -2837 3387 -2675
rect 3341 -3322 3387 -3311
rect 3501 -1565 3547 -1554
rect 3501 -2201 3547 -2039
rect 3501 -2837 3547 -2675
rect 2253 -3506 3259 -3460
rect 3501 -3552 3547 -3311
rect 3745 -1565 3791 -1554
rect 3745 -2201 3791 -2039
rect 3745 -2837 3791 -2675
rect 3745 -3552 3791 -3311
rect 3905 -1565 3951 -1436
rect 4673 -1462 4719 -1340
rect 3905 -2201 3951 -2039
rect 3905 -2837 3951 -2675
rect 3905 -3322 3951 -3311
rect 4033 -1508 4719 -1462
rect 4033 -1565 4079 -1508
rect 4033 -2201 4079 -2039
rect 4033 -2837 4079 -2675
rect 4033 -3460 4079 -3311
rect 4193 -1565 4239 -1554
rect 4193 -2201 4239 -2039
rect 4193 -2837 4239 -2675
rect 4193 -3368 4239 -3311
rect 4353 -1565 4399 -1508
rect 4353 -2201 4399 -2039
rect 4353 -2837 4399 -2675
rect 4353 -3322 4399 -3311
rect 4513 -1565 4559 -1554
rect 4513 -2201 4559 -2039
rect 4513 -2837 4559 -2675
rect 4513 -3368 4559 -3311
rect 4673 -1565 4719 -1508
rect 4673 -2201 4719 -2039
rect 4673 -2837 4719 -2675
rect 4673 -3322 4719 -3311
rect 4833 -241 4879 -214
rect 4833 -627 4879 -465
rect 4833 -1013 4879 -851
rect 4833 -1344 4879 -1237
rect 4993 -241 5039 -184
rect 4993 -627 5039 -465
rect 4993 -1013 5039 -851
rect 4993 -1248 5039 -1237
rect 5153 -241 5199 -230
rect 5153 -627 5199 -465
rect 5153 -1013 5199 -851
rect 5153 -1344 5199 -1237
rect 5313 -241 5359 -184
rect 5313 -627 5359 -465
rect 5313 -1013 5359 -851
rect 5313 -1248 5359 -1237
rect 5557 -184 5923 -138
rect 5557 -241 5603 -184
rect 5557 -627 5603 -465
rect 5557 -1013 5603 -851
rect 5557 -1248 5603 -1237
rect 5717 -241 5763 -230
rect 5717 -627 5763 -465
rect 5717 -1013 5763 -851
rect 5717 -1344 5763 -1237
rect 5877 -241 5923 -184
rect 5877 -627 5923 -465
rect 5877 -1013 5923 -851
rect 5877 -1248 5923 -1237
rect 6037 -150 6738 -138
rect 6037 -184 6674 -150
rect 6037 -241 6083 -184
rect 6037 -627 6083 -465
rect 6037 -1013 6083 -851
rect 6037 -1344 6083 -1237
rect 4833 -1390 5302 -1344
rect 5614 -1390 6083 -1344
rect 4833 -1565 4879 -1390
rect 4833 -2201 4879 -2039
rect 4833 -2837 4879 -2675
rect 4833 -3368 4879 -3311
rect 4193 -3414 4879 -3368
rect 4993 -1565 5039 -1554
rect 4993 -2201 5039 -2039
rect 4993 -2837 5039 -2675
rect 4993 -3368 5039 -3311
rect 5153 -1565 5199 -1390
rect 5153 -2201 5199 -2039
rect 5153 -2837 5199 -2675
rect 5153 -3322 5199 -3311
rect 5313 -1565 5603 -1539
rect 5359 -1585 5557 -1565
rect 5313 -2201 5359 -2039
rect 5313 -2837 5359 -2675
rect 5313 -3368 5359 -3311
rect 5557 -2201 5603 -2039
rect 5557 -2837 5603 -2675
rect 5557 -3353 5603 -3311
rect 5717 -1565 5763 -1390
rect 5717 -2201 5763 -2039
rect 5717 -2837 5763 -2675
rect 5717 -3322 5763 -3311
rect 5877 -1565 5923 -1554
rect 5877 -2201 5923 -2039
rect 5877 -2837 5923 -2675
rect 4993 -3414 5359 -3368
rect 5542 -3365 5618 -3353
rect 4993 -3460 5039 -3414
rect 5542 -3417 5554 -3365
rect 5606 -3368 5618 -3365
rect 5877 -3368 5923 -3311
rect 5606 -3414 5923 -3368
rect 6037 -1565 6083 -1390
rect 6037 -2201 6083 -2039
rect 6037 -2837 6083 -2675
rect 6037 -3368 6083 -3311
rect 6197 -241 6243 -230
rect 6197 -627 6243 -465
rect 6197 -1013 6243 -851
rect 6197 -1294 6243 -1237
rect 6357 -241 6403 -184
rect 6662 -202 6674 -184
rect 6726 -202 6738 -150
rect 6662 -214 6738 -202
rect 6357 -627 6403 -465
rect 6357 -1013 6403 -851
rect 6357 -1248 6403 -1237
rect 6517 -241 6563 -230
rect 6517 -627 6563 -465
rect 6517 -1013 6563 -851
rect 6517 -1294 6563 -1237
rect 6677 -241 6723 -214
rect 6677 -627 6723 -465
rect 6677 -1013 6723 -851
rect 6677 -1248 6723 -1237
rect 6837 -241 6883 -92
rect 6837 -627 6883 -465
rect 6837 -1013 6883 -851
rect 6837 -1294 6883 -1237
rect 6197 -1340 6883 -1294
rect 6965 -241 7011 -230
rect 6965 -627 7011 -465
rect 6965 -1013 7011 -851
rect 6197 -1462 6243 -1340
rect 6965 -1368 7011 -1237
rect 7125 -241 7171 0
rect 7689 -92 8695 -46
rect 7689 -138 7735 -92
rect 7349 -150 7735 -138
rect 7349 -202 7361 -150
rect 7413 -184 7735 -150
rect 7413 -202 7425 -184
rect 7349 -214 7425 -202
rect 7125 -627 7171 -465
rect 7125 -1013 7171 -851
rect 7125 -1248 7171 -1237
rect 7369 -241 7415 -214
rect 7369 -627 7415 -465
rect 7369 -1013 7415 -851
rect 7369 -1248 7415 -1237
rect 7529 -241 7575 -230
rect 7529 -627 7575 -465
rect 7529 -1013 7575 -851
rect 7529 -1344 7575 -1237
rect 7689 -241 7735 -184
rect 7689 -627 7735 -465
rect 7689 -1013 7735 -851
rect 7689 -1248 7735 -1237
rect 7849 -184 8535 -138
rect 7849 -241 7895 -184
rect 7849 -627 7895 -465
rect 7849 -1013 7895 -851
rect 7849 -1329 7895 -1237
rect 8009 -241 8055 -230
rect 8009 -627 8055 -465
rect 8009 -1013 8055 -851
rect 8009 -1294 8055 -1237
rect 8169 -241 8215 -184
rect 8169 -627 8215 -465
rect 8169 -1013 8215 -851
rect 8169 -1248 8215 -1237
rect 8329 -241 8375 -230
rect 8329 -627 8375 -465
rect 8329 -1013 8375 -851
rect 8329 -1294 8375 -1237
rect 8489 -241 8535 -184
rect 8489 -627 8535 -465
rect 8489 -1013 8535 -851
rect 8489 -1248 8535 -1237
rect 8649 -241 8695 -92
rect 8649 -627 8695 -465
rect 8649 -1013 8695 -851
rect 8649 -1294 8695 -1237
rect 7834 -1341 7910 -1329
rect 7834 -1344 7846 -1341
rect 6922 -1379 7011 -1368
rect 7146 -1366 7214 -1358
rect 7146 -1369 7154 -1366
rect 7206 -1369 7214 -1366
rect 6922 -1425 6933 -1379
rect 6979 -1425 7011 -1379
rect 7142 -1415 7154 -1369
rect 7206 -1415 7259 -1369
rect 7426 -1390 7846 -1344
rect 6922 -1436 7011 -1425
rect 7146 -1418 7154 -1415
rect 7206 -1418 7214 -1415
rect 7146 -1426 7214 -1418
rect 6197 -1508 6883 -1462
rect 6197 -1565 6243 -1508
rect 6197 -2201 6243 -2039
rect 6197 -2837 6243 -2675
rect 6197 -3322 6243 -3311
rect 6357 -1565 6403 -1554
rect 6357 -2201 6403 -2039
rect 6357 -2837 6403 -2675
rect 6357 -3368 6403 -3311
rect 6517 -1565 6563 -1508
rect 6517 -2201 6563 -2039
rect 6517 -2837 6563 -2675
rect 6517 -3322 6563 -3311
rect 6677 -1565 6723 -1554
rect 6677 -2201 6723 -2039
rect 6677 -2837 6723 -2675
rect 6677 -3368 6723 -3311
rect 6037 -3414 6723 -3368
rect 6837 -1565 6883 -1508
rect 6837 -2201 6883 -2039
rect 6837 -2837 6883 -2675
rect 5606 -3417 5618 -3414
rect 5542 -3429 5618 -3417
rect 4033 -3506 5039 -3460
rect 5877 -3460 5923 -3414
rect 6837 -3460 6883 -3311
rect 6965 -1565 7011 -1436
rect 6965 -2201 7011 -2039
rect 6965 -2837 7011 -2675
rect 6965 -3322 7011 -3311
rect 7125 -1565 7171 -1554
rect 7261 -1565 7415 -1539
rect 7261 -1585 7369 -1565
rect 7125 -2201 7171 -2039
rect 7125 -2837 7171 -2675
rect 5877 -3506 6883 -3460
rect 7125 -3552 7171 -3311
rect 7369 -2201 7415 -2039
rect 7369 -2837 7415 -2675
rect 7369 -3368 7415 -3311
rect 7529 -1565 7575 -1390
rect 7834 -1393 7846 -1390
rect 7898 -1393 7910 -1341
rect 7834 -1405 7910 -1393
rect 8009 -1340 8695 -1294
rect 8777 -241 8823 -230
rect 8777 -627 8823 -465
rect 8777 -1013 8823 -851
rect 7529 -2201 7575 -2039
rect 7529 -2837 7575 -2675
rect 7529 -3322 7575 -3311
rect 7689 -1565 7735 -1554
rect 7689 -2201 7735 -2039
rect 7689 -2837 7735 -2675
rect 7689 -3368 7735 -3311
rect 7369 -3414 7735 -3368
rect 7849 -1565 7895 -1405
rect 7849 -2201 7895 -2039
rect 7849 -2837 7895 -2675
rect 7849 -3368 7895 -3311
rect 8009 -1462 8055 -1340
rect 8777 -1368 8823 -1237
rect 8937 -241 8983 0
rect 8937 -627 8983 -465
rect 8937 -1013 8983 -851
rect 8937 -1248 8983 -1237
rect 9118 -1341 9194 -1329
rect 8734 -1379 8823 -1368
rect 8734 -1425 8745 -1379
rect 8791 -1425 8823 -1379
rect 8734 -1436 8823 -1425
rect 8958 -1366 9026 -1358
rect 8958 -1418 8966 -1366
rect 9018 -1369 9026 -1366
rect 9018 -1415 9071 -1369
rect 9118 -1393 9130 -1341
rect 9182 -1344 9194 -1341
rect 9182 -1390 9282 -1344
rect 9182 -1393 9194 -1390
rect 9118 -1405 9194 -1393
rect 9018 -1418 9026 -1415
rect 8958 -1426 9026 -1418
rect 8009 -1508 8695 -1462
rect 8009 -1565 8055 -1508
rect 8009 -2201 8055 -2039
rect 8009 -2837 8055 -2675
rect 8009 -3322 8055 -3311
rect 8169 -1565 8215 -1554
rect 8169 -2201 8215 -2039
rect 8169 -2837 8215 -2675
rect 8169 -3368 8215 -3311
rect 8329 -1565 8375 -1508
rect 8329 -2201 8375 -2039
rect 8329 -2837 8375 -2675
rect 8329 -3322 8375 -3311
rect 8489 -1565 8535 -1554
rect 8489 -2201 8535 -2039
rect 8489 -2837 8535 -2675
rect 8489 -3368 8535 -3311
rect 7849 -3414 8535 -3368
rect 8649 -1565 8695 -1508
rect 8649 -2201 8695 -2039
rect 8649 -2837 8695 -2675
rect 7689 -3460 7735 -3414
rect 8649 -3460 8695 -3311
rect 8777 -1565 8823 -1436
rect 8777 -2201 8823 -2039
rect 8777 -2837 8823 -2675
rect 8777 -3322 8823 -3311
rect 8937 -1565 8983 -1554
rect 8937 -2201 8983 -2039
rect 8937 -2837 8983 -2675
rect 7689 -3506 8695 -3460
rect 8937 -3552 8983 -3311
rect -4175 -3582 9082 -3552
rect -4175 -3585 -3953 -3582
rect -3901 -3585 -3653 -3582
rect -3601 -3585 -3353 -3582
rect -3301 -3585 -3053 -3582
rect -3001 -3585 -2753 -3582
rect -2701 -3585 9082 -3582
rect -4175 -3631 -4138 -3585
rect -4092 -3631 -4044 -3585
rect -3998 -3631 -3953 -3585
rect -3901 -3631 -3856 -3585
rect -3810 -3631 -3762 -3585
rect -3716 -3631 -3668 -3585
rect -3601 -3631 -3574 -3585
rect -3528 -3631 -3480 -3585
rect -3434 -3631 -3386 -3585
rect -3301 -3631 -3292 -3585
rect -3246 -3631 -3198 -3585
rect -3152 -3631 -3104 -3585
rect -3058 -3631 -3053 -3585
rect -2964 -3631 -2916 -3585
rect -2870 -3631 -2822 -3585
rect -2776 -3631 -2753 -3585
rect -2682 -3631 -2634 -3585
rect -2588 -3631 -2540 -3585
rect -2494 -3631 -2446 -3585
rect -2400 -3631 -2326 -3585
rect -2280 -3631 -2232 -3585
rect -2186 -3631 -2138 -3585
rect -2092 -3631 -2044 -3585
rect -1998 -3631 -1950 -3585
rect -1904 -3631 -1856 -3585
rect -1810 -3631 -1762 -3585
rect -1716 -3631 -1668 -3585
rect -1622 -3631 -1574 -3585
rect -1528 -3631 -1480 -3585
rect -1434 -3631 -1386 -3585
rect -1340 -3631 -1292 -3585
rect -1246 -3631 -1198 -3585
rect -1152 -3631 -1104 -3585
rect -1058 -3631 -1010 -3585
rect -964 -3631 -916 -3585
rect -870 -3631 -822 -3585
rect -776 -3631 -728 -3585
rect -682 -3631 -634 -3585
rect -588 -3631 59 -3585
rect 105 -3631 153 -3585
rect 199 -3631 247 -3585
rect 293 -3631 341 -3585
rect 387 -3631 435 -3585
rect 481 -3631 529 -3585
rect 575 -3631 623 -3585
rect 669 -3631 717 -3585
rect 763 -3631 811 -3585
rect 857 -3631 905 -3585
rect 951 -3631 999 -3585
rect 1045 -3631 1093 -3585
rect 1139 -3631 1187 -3585
rect 1233 -3631 1281 -3585
rect 1327 -3631 1375 -3585
rect 1421 -3631 1469 -3585
rect 1515 -3631 1563 -3585
rect 1609 -3631 1657 -3585
rect 1703 -3631 1751 -3585
rect 1797 -3631 1871 -3585
rect 1917 -3631 1965 -3585
rect 2011 -3631 2059 -3585
rect 2105 -3631 2153 -3585
rect 2199 -3631 2247 -3585
rect 2293 -3631 2341 -3585
rect 2387 -3631 2435 -3585
rect 2481 -3631 2529 -3585
rect 2575 -3631 2623 -3585
rect 2669 -3631 2717 -3585
rect 2763 -3631 2811 -3585
rect 2857 -3631 2905 -3585
rect 2951 -3631 2999 -3585
rect 3045 -3631 3093 -3585
rect 3139 -3631 3187 -3585
rect 3233 -3631 3281 -3585
rect 3327 -3631 3375 -3585
rect 3421 -3631 3469 -3585
rect 3515 -3631 3563 -3585
rect 3609 -3631 3683 -3585
rect 3729 -3631 3777 -3585
rect 3823 -3631 3871 -3585
rect 3917 -3631 3965 -3585
rect 4011 -3631 4059 -3585
rect 4105 -3631 4153 -3585
rect 4199 -3631 4247 -3585
rect 4293 -3631 4341 -3585
rect 4387 -3631 4435 -3585
rect 4481 -3631 4529 -3585
rect 4575 -3631 4623 -3585
rect 4669 -3631 4717 -3585
rect 4763 -3631 4811 -3585
rect 4857 -3631 4905 -3585
rect 4951 -3631 4999 -3585
rect 5045 -3631 5093 -3585
rect 5139 -3631 5187 -3585
rect 5233 -3631 5281 -3585
rect 5327 -3631 5375 -3585
rect 5421 -3631 5495 -3585
rect 5541 -3631 5589 -3585
rect 5635 -3631 5683 -3585
rect 5729 -3631 5777 -3585
rect 5823 -3631 5871 -3585
rect 5917 -3631 5965 -3585
rect 6011 -3631 6059 -3585
rect 6105 -3631 6153 -3585
rect 6199 -3631 6247 -3585
rect 6293 -3631 6341 -3585
rect 6387 -3631 6435 -3585
rect 6481 -3631 6529 -3585
rect 6575 -3631 6623 -3585
rect 6669 -3631 6717 -3585
rect 6763 -3631 6811 -3585
rect 6857 -3631 6905 -3585
rect 6951 -3631 6999 -3585
rect 7045 -3631 7093 -3585
rect 7139 -3631 7187 -3585
rect 7233 -3631 7307 -3585
rect 7353 -3631 7401 -3585
rect 7447 -3631 7495 -3585
rect 7541 -3631 7589 -3585
rect 7635 -3631 7683 -3585
rect 7729 -3631 7777 -3585
rect 7823 -3631 7871 -3585
rect 7917 -3631 7965 -3585
rect 8011 -3631 8059 -3585
rect 8105 -3631 8153 -3585
rect 8199 -3631 8247 -3585
rect 8293 -3631 8341 -3585
rect 8387 -3631 8435 -3585
rect 8481 -3631 8529 -3585
rect 8575 -3631 8623 -3585
rect 8669 -3631 8717 -3585
rect 8763 -3631 8811 -3585
rect 8857 -3631 8905 -3585
rect 8951 -3631 8999 -3585
rect 9045 -3631 9082 -3585
rect -4175 -3634 -3953 -3631
rect -3901 -3634 -3653 -3631
rect -3601 -3634 -3353 -3631
rect -3301 -3634 -3053 -3631
rect -3001 -3634 -2753 -3631
rect -2701 -3634 9082 -3631
rect -4175 -3664 9082 -3634
rect -4285 -3799 -4209 -3787
rect -4285 -3802 -4273 -3799
rect -4398 -3848 -4273 -3802
rect -4285 -3851 -4273 -3848
rect -4221 -3851 -4209 -3799
rect -4285 -3863 -4209 -3851
rect -4076 -3905 -4030 -3664
rect -3788 -3756 -2782 -3710
rect -4076 -4541 -4030 -4379
rect -4076 -5177 -4030 -5015
rect -4076 -5662 -4030 -5651
rect -3916 -3905 -3870 -3894
rect -3916 -4541 -3870 -4379
rect -3916 -5177 -3870 -5015
rect -3916 -5780 -3870 -5651
rect -3788 -3905 -3742 -3756
rect -2828 -3802 -2782 -3756
rect -1944 -3756 -938 -3710
rect -2523 -3799 -2447 -3787
rect -2523 -3802 -2511 -3799
rect -3788 -4541 -3742 -4379
rect -3788 -5177 -3742 -5015
rect -3788 -5708 -3742 -5651
rect -3628 -3848 -2942 -3802
rect -3628 -3905 -3582 -3848
rect -3628 -4541 -3582 -4379
rect -3628 -5177 -3582 -5015
rect -3628 -5662 -3582 -5651
rect -3468 -3905 -3422 -3894
rect -3468 -4541 -3422 -4379
rect -3468 -5177 -3422 -5015
rect -3468 -5708 -3422 -5651
rect -3308 -3905 -3262 -3848
rect -3308 -4541 -3262 -4379
rect -3308 -5177 -3262 -5015
rect -3308 -5662 -3262 -5651
rect -3148 -3905 -3102 -3894
rect -3148 -4541 -3102 -4379
rect -3148 -5177 -3102 -5015
rect -3148 -5708 -3102 -5651
rect -3788 -5754 -3102 -5708
rect -4119 -5798 -4051 -5790
rect -4119 -5801 -4111 -5798
rect -4164 -5847 -4111 -5801
rect -4119 -5850 -4111 -5847
rect -4059 -5850 -4051 -5798
rect -4119 -5858 -4051 -5850
rect -3916 -5791 -3827 -5780
rect -3916 -5837 -3884 -5791
rect -3838 -5837 -3827 -5791
rect -3916 -5848 -3827 -5837
rect -4076 -5979 -4030 -5968
rect -4076 -6365 -4030 -6203
rect -4076 -6751 -4030 -6589
rect -4076 -7216 -4030 -6975
rect -3916 -5979 -3870 -5848
rect -3148 -5876 -3102 -5754
rect -3916 -6365 -3870 -6203
rect -3916 -6751 -3870 -6589
rect -3916 -6986 -3870 -6975
rect -3788 -5922 -3102 -5876
rect -3788 -5979 -3742 -5922
rect -3788 -6365 -3742 -6203
rect -3788 -6751 -3742 -6589
rect -3788 -7124 -3742 -6975
rect -3628 -5979 -3582 -5968
rect -3628 -6365 -3582 -6203
rect -3628 -6751 -3582 -6589
rect -3628 -7032 -3582 -6975
rect -3468 -5979 -3422 -5922
rect -3468 -6365 -3422 -6203
rect -3468 -6751 -3422 -6589
rect -3468 -6986 -3422 -6975
rect -3308 -5979 -3262 -5968
rect -3308 -6365 -3262 -6203
rect -3308 -6751 -3262 -6589
rect -3308 -7032 -3262 -6975
rect -3148 -5979 -3102 -5922
rect -3148 -6365 -3102 -6203
rect -3148 -6751 -3102 -6589
rect -3148 -6986 -3102 -6975
rect -2988 -3905 -2942 -3848
rect -2988 -4541 -2942 -4379
rect -2988 -5177 -2942 -5015
rect -2988 -5826 -2942 -5651
rect -2828 -3848 -2511 -3802
rect -2828 -3905 -2782 -3848
rect -2523 -3851 -2511 -3848
rect -2459 -3851 -2447 -3799
rect -1944 -3802 -1898 -3756
rect -2523 -3863 -2447 -3851
rect -2264 -3848 -1898 -3802
rect -2828 -4541 -2782 -4379
rect -2828 -5177 -2782 -5015
rect -2828 -5662 -2782 -5651
rect -2668 -3905 -2622 -3894
rect -2668 -4541 -2622 -4379
rect -2668 -5177 -2622 -5015
rect -2668 -5826 -2622 -5651
rect -2508 -3905 -2462 -3863
rect -2508 -4541 -2462 -4379
rect -2508 -5177 -2462 -5015
rect -2264 -3905 -2218 -3848
rect -2264 -4541 -2218 -4379
rect -2264 -5177 -2218 -5015
rect -2462 -5651 -2264 -5631
rect -2508 -5677 -2218 -5651
rect -2104 -3905 -2058 -3894
rect -2104 -4541 -2058 -4379
rect -2104 -5177 -2058 -5015
rect -2104 -5826 -2058 -5651
rect -1944 -3905 -1898 -3848
rect -1944 -4541 -1898 -4379
rect -1944 -5177 -1898 -5015
rect -1944 -5662 -1898 -5651
rect -1784 -3814 -1083 -3802
rect -1784 -3848 -1147 -3814
rect -1784 -3905 -1738 -3848
rect -1784 -4541 -1738 -4379
rect -1784 -5177 -1738 -5015
rect -1784 -5826 -1738 -5651
rect -2988 -5872 -2519 -5826
rect -2207 -5872 -1738 -5826
rect -2988 -5979 -2942 -5872
rect -2988 -6365 -2942 -6203
rect -2988 -6751 -2942 -6589
rect -2988 -7002 -2942 -6975
rect -2828 -5979 -2782 -5968
rect -2828 -6365 -2782 -6203
rect -2828 -6751 -2782 -6589
rect -3003 -7014 -2927 -7002
rect -3003 -7032 -2991 -7014
rect -3628 -7066 -2991 -7032
rect -2939 -7066 -2927 -7014
rect -3628 -7078 -2927 -7066
rect -2828 -7032 -2782 -6975
rect -2668 -5979 -2622 -5872
rect -2668 -6365 -2622 -6203
rect -2668 -6751 -2622 -6589
rect -2668 -6986 -2622 -6975
rect -2508 -5979 -2462 -5968
rect -2508 -6365 -2462 -6203
rect -2508 -6751 -2462 -6589
rect -2508 -7032 -2462 -6975
rect -2828 -7078 -2462 -7032
rect -2264 -5979 -2218 -5968
rect -2264 -6365 -2218 -6203
rect -2264 -6751 -2218 -6589
rect -2264 -7032 -2218 -6975
rect -2104 -5979 -2058 -5872
rect -2104 -6365 -2058 -6203
rect -2104 -6751 -2058 -6589
rect -2104 -6986 -2058 -6975
rect -1944 -5979 -1898 -5968
rect -1944 -6365 -1898 -6203
rect -1944 -6751 -1898 -6589
rect -1944 -7032 -1898 -6975
rect -2264 -7078 -1898 -7032
rect -1784 -5979 -1738 -5872
rect -1784 -6365 -1738 -6203
rect -1784 -6751 -1738 -6589
rect -1784 -7032 -1738 -6975
rect -1624 -3905 -1578 -3894
rect -1624 -4541 -1578 -4379
rect -1624 -5177 -1578 -5015
rect -1624 -5708 -1578 -5651
rect -1464 -3905 -1418 -3848
rect -1159 -3866 -1147 -3848
rect -1095 -3866 -1083 -3814
rect -1159 -3878 -1083 -3866
rect -1464 -4541 -1418 -4379
rect -1464 -5177 -1418 -5015
rect -1464 -5662 -1418 -5651
rect -1304 -3905 -1258 -3894
rect -1304 -4541 -1258 -4379
rect -1304 -5177 -1258 -5015
rect -1304 -5708 -1258 -5651
rect -1144 -3905 -1098 -3878
rect -1144 -4541 -1098 -4379
rect -1144 -5177 -1098 -5015
rect -1144 -5662 -1098 -5651
rect -984 -3905 -938 -3756
rect -984 -4541 -938 -4379
rect -984 -5177 -938 -5015
rect -984 -5708 -938 -5651
rect -1624 -5754 -938 -5708
rect -856 -3905 -810 -3894
rect -856 -4541 -810 -4379
rect -856 -5177 -810 -5015
rect -1624 -5876 -1578 -5754
rect -856 -5780 -810 -5651
rect -696 -3905 -650 -3664
rect -696 -4541 -650 -4379
rect -696 -5177 -650 -5015
rect -696 -5662 -650 -5651
rect 121 -3905 167 -3664
rect 409 -3756 1415 -3710
rect 121 -4541 167 -4379
rect 121 -5177 167 -5015
rect 121 -5662 167 -5651
rect 281 -3905 327 -3894
rect 281 -4541 327 -4379
rect 281 -5177 327 -5015
rect -899 -5791 -810 -5780
rect 281 -5780 327 -5651
rect 409 -3905 455 -3756
rect 1369 -3802 1415 -3756
rect 2253 -3756 3259 -3710
rect 2253 -3802 2299 -3756
rect 409 -4541 455 -4379
rect 409 -5177 455 -5015
rect 409 -5708 455 -5651
rect 569 -3848 1255 -3802
rect 569 -3905 615 -3848
rect 569 -4541 615 -4379
rect 569 -5177 615 -5015
rect 569 -5662 615 -5651
rect 729 -3905 775 -3894
rect 729 -4541 775 -4379
rect 729 -5177 775 -5015
rect 729 -5708 775 -5651
rect 889 -3905 935 -3848
rect 889 -4541 935 -4379
rect 889 -5177 935 -5015
rect 889 -5662 935 -5651
rect 1049 -3905 1095 -3894
rect 1049 -4541 1095 -4379
rect 1049 -5177 1095 -5015
rect 1049 -5708 1095 -5651
rect 409 -5754 1095 -5708
rect -899 -5837 -888 -5791
rect -842 -5837 -810 -5791
rect -899 -5848 -810 -5837
rect -1624 -5922 -938 -5876
rect -1624 -5979 -1578 -5922
rect -1624 -6365 -1578 -6203
rect -1624 -6751 -1578 -6589
rect -1624 -6986 -1578 -6975
rect -1464 -5979 -1418 -5968
rect -1464 -6365 -1418 -6203
rect -1464 -6751 -1418 -6589
rect -1464 -7032 -1418 -6975
rect -1304 -5979 -1258 -5922
rect -1304 -6365 -1258 -6203
rect -1304 -6751 -1258 -6589
rect -1304 -6986 -1258 -6975
rect -1144 -5979 -1098 -5968
rect -1144 -6365 -1098 -6203
rect -1144 -6751 -1098 -6589
rect -1144 -7032 -1098 -6975
rect -1784 -7078 -1098 -7032
rect -984 -5979 -938 -5922
rect -984 -6365 -938 -6203
rect -984 -6751 -938 -6589
rect -2828 -7124 -2782 -7078
rect -3788 -7170 -2782 -7124
rect -1944 -7124 -1898 -7078
rect -984 -7124 -938 -6975
rect -856 -5979 -810 -5848
rect -679 -5798 -603 -5786
rect -679 -5850 -667 -5798
rect -615 -5801 -603 -5798
rect -303 -5798 -227 -5786
rect -615 -5847 -562 -5801
rect -615 -5850 -603 -5847
rect -679 -5862 -603 -5850
rect -303 -5850 -291 -5798
rect -239 -5801 -227 -5798
rect 78 -5798 146 -5790
rect 78 -5801 86 -5798
rect -239 -5847 86 -5801
rect -239 -5850 -227 -5847
rect -303 -5862 -227 -5850
rect 78 -5850 86 -5847
rect 138 -5850 146 -5798
rect 78 -5858 146 -5850
rect 281 -5791 370 -5780
rect 281 -5837 313 -5791
rect 359 -5837 370 -5791
rect 281 -5848 370 -5837
rect -856 -6365 -810 -6203
rect -856 -6751 -810 -6589
rect -856 -6986 -810 -6975
rect -696 -5979 -650 -5968
rect -696 -6365 -650 -6203
rect -696 -6751 -650 -6589
rect -1944 -7170 -938 -7124
rect -696 -7216 -650 -6975
rect 121 -5979 167 -5968
rect 121 -6365 167 -6203
rect 121 -6751 167 -6589
rect 121 -7216 167 -6975
rect 281 -5979 327 -5848
rect 1049 -5876 1095 -5754
rect 281 -6365 327 -6203
rect 281 -6751 327 -6589
rect 281 -6986 327 -6975
rect 409 -5922 1095 -5876
rect 409 -5979 455 -5922
rect 409 -6365 455 -6203
rect 409 -6751 455 -6589
rect 409 -7002 455 -6975
rect 569 -5979 615 -5968
rect 569 -6365 615 -6203
rect 569 -6751 615 -6589
rect 389 -7014 465 -7002
rect 389 -7066 401 -7014
rect 453 -7066 465 -7014
rect 389 -7078 465 -7066
rect 569 -7032 615 -6975
rect 729 -5979 775 -5922
rect 729 -6365 775 -6203
rect 729 -6751 775 -6589
rect 729 -6986 775 -6975
rect 889 -5979 935 -5968
rect 889 -6365 935 -6203
rect 889 -6751 935 -6589
rect 889 -7032 935 -6975
rect 1049 -5979 1095 -5922
rect 1049 -6365 1095 -6203
rect 1049 -6751 1095 -6589
rect 1049 -6986 1095 -6975
rect 1209 -3905 1255 -3848
rect 1209 -4541 1255 -4379
rect 1209 -5177 1255 -5015
rect 1209 -5826 1255 -5651
rect 1369 -3848 1735 -3802
rect 1369 -3905 1415 -3848
rect 1369 -4541 1415 -4379
rect 1369 -5177 1415 -5015
rect 1369 -5662 1415 -5651
rect 1529 -3905 1575 -3894
rect 1529 -4541 1575 -4379
rect 1529 -5177 1575 -5015
rect 1529 -5826 1575 -5651
rect 1689 -3905 1735 -3848
rect 1689 -4541 1735 -4379
rect 1689 -5177 1735 -5015
rect 1933 -3848 2299 -3802
rect 1933 -3905 1979 -3848
rect 1933 -4541 1979 -4379
rect 1933 -5177 1979 -5015
rect 1735 -5651 1933 -5631
rect 1689 -5677 1979 -5651
rect 2093 -3905 2139 -3894
rect 2093 -4541 2139 -4379
rect 2093 -5177 2139 -5015
rect 1674 -5823 1750 -5811
rect 1674 -5826 1686 -5823
rect 1209 -5872 1686 -5826
rect 1209 -5979 1255 -5872
rect 1209 -6365 1255 -6203
rect 1209 -6751 1255 -6589
rect 1209 -7032 1255 -6975
rect 569 -7078 1255 -7032
rect 1369 -5979 1415 -5968
rect 1369 -6365 1415 -6203
rect 1369 -6751 1415 -6589
rect 1369 -7032 1415 -6975
rect 1529 -5979 1575 -5872
rect 1674 -5875 1686 -5872
rect 1738 -5875 1750 -5823
rect 1674 -5887 1750 -5875
rect 1918 -5823 1994 -5811
rect 1918 -5875 1930 -5823
rect 1982 -5826 1994 -5823
rect 2093 -5826 2139 -5651
rect 2253 -3905 2299 -3848
rect 2253 -4541 2299 -4379
rect 2253 -5177 2299 -5015
rect 2253 -5662 2299 -5651
rect 2413 -3848 3099 -3802
rect 2413 -3905 2459 -3848
rect 2413 -4541 2459 -4379
rect 2413 -5177 2459 -5015
rect 2413 -5826 2459 -5651
rect 1982 -5872 2459 -5826
rect 1982 -5875 1994 -5872
rect 1918 -5887 1994 -5875
rect 1529 -6365 1575 -6203
rect 1529 -6751 1575 -6589
rect 1529 -6986 1575 -6975
rect 1689 -5979 1735 -5968
rect 1689 -6365 1735 -6203
rect 1689 -6751 1735 -6589
rect 1689 -7032 1735 -6975
rect 1369 -7078 1735 -7032
rect 1933 -5979 1979 -5968
rect 1933 -6365 1979 -6203
rect 1933 -6751 1979 -6589
rect 1933 -7032 1979 -6975
rect 2093 -5979 2139 -5872
rect 2093 -6365 2139 -6203
rect 2093 -6751 2139 -6589
rect 2093 -6986 2139 -6975
rect 2253 -5979 2299 -5968
rect 2253 -6365 2299 -6203
rect 2253 -6751 2299 -6589
rect 2253 -7032 2299 -6975
rect 1933 -7078 2299 -7032
rect 2413 -5979 2459 -5872
rect 2413 -6365 2459 -6203
rect 2413 -6751 2459 -6589
rect 2413 -7032 2459 -6975
rect 2573 -3905 2619 -3894
rect 2573 -4541 2619 -4379
rect 2573 -5177 2619 -5015
rect 2573 -5708 2619 -5651
rect 2733 -3905 2779 -3848
rect 2733 -4541 2779 -4379
rect 2733 -5177 2779 -5015
rect 2733 -5662 2779 -5651
rect 2893 -3905 2939 -3894
rect 2893 -4541 2939 -4379
rect 2893 -5177 2939 -5015
rect 2893 -5708 2939 -5651
rect 3053 -3905 3099 -3848
rect 3053 -4541 3099 -4379
rect 3053 -5177 3099 -5015
rect 3053 -5662 3099 -5651
rect 3213 -3905 3259 -3756
rect 3213 -4541 3259 -4379
rect 3213 -5177 3259 -5015
rect 3213 -5708 3259 -5651
rect 2573 -5754 3259 -5708
rect 3341 -3905 3387 -3894
rect 3341 -4541 3387 -4379
rect 3341 -5177 3387 -5015
rect 2573 -5876 2619 -5754
rect 3341 -5780 3387 -5651
rect 3501 -3905 3547 -3664
rect 3501 -4541 3547 -4379
rect 3501 -5177 3547 -5015
rect 3501 -5662 3547 -5651
rect 3745 -3905 3791 -3664
rect 4033 -3756 5039 -3710
rect 4033 -3802 4079 -3756
rect 4993 -3802 5039 -3756
rect 5877 -3756 6883 -3710
rect 5877 -3802 5923 -3756
rect 4013 -3814 4089 -3802
rect 4013 -3866 4025 -3814
rect 4077 -3866 4089 -3814
rect 4013 -3878 4089 -3866
rect 4193 -3848 4879 -3802
rect 3745 -4541 3791 -4379
rect 3745 -5177 3791 -5015
rect 3745 -5662 3791 -5651
rect 3905 -3905 3951 -3894
rect 3905 -4541 3951 -4379
rect 3905 -5177 3951 -5015
rect 3298 -5791 3387 -5780
rect 3905 -5780 3951 -5651
rect 4033 -3905 4079 -3878
rect 4033 -4541 4079 -4379
rect 4033 -5177 4079 -5015
rect 4033 -5708 4079 -5651
rect 4193 -3905 4239 -3848
rect 4193 -4541 4239 -4379
rect 4193 -5177 4239 -5015
rect 4193 -5662 4239 -5651
rect 4353 -3905 4399 -3894
rect 4353 -4541 4399 -4379
rect 4353 -5177 4399 -5015
rect 4353 -5708 4399 -5651
rect 4513 -3905 4559 -3848
rect 4513 -4541 4559 -4379
rect 4513 -5177 4559 -5015
rect 4513 -5662 4559 -5651
rect 4673 -3905 4719 -3894
rect 4673 -4541 4719 -4379
rect 4673 -5177 4719 -5015
rect 4673 -5708 4719 -5651
rect 4033 -5754 4719 -5708
rect 3298 -5837 3309 -5791
rect 3355 -5837 3387 -5791
rect 3298 -5848 3387 -5837
rect 2573 -5922 3259 -5876
rect 2573 -5979 2619 -5922
rect 2573 -6365 2619 -6203
rect 2573 -6751 2619 -6589
rect 2573 -6986 2619 -6975
rect 2733 -5979 2779 -5968
rect 2733 -6365 2779 -6203
rect 2733 -6751 2779 -6589
rect 2733 -7032 2779 -6975
rect 2893 -5979 2939 -5922
rect 2893 -6365 2939 -6203
rect 2893 -6751 2939 -6589
rect 2893 -6986 2939 -6975
rect 3053 -5979 3099 -5968
rect 3053 -6365 3099 -6203
rect 3053 -6751 3099 -6589
rect 3053 -7032 3099 -6975
rect 2413 -7078 3099 -7032
rect 3213 -5979 3259 -5922
rect 3213 -6365 3259 -6203
rect 3213 -6751 3259 -6589
rect 409 -7124 455 -7078
rect 1369 -7124 1415 -7078
rect 409 -7170 1415 -7124
rect 2253 -7124 2299 -7078
rect 3213 -7124 3259 -6975
rect 3341 -5979 3387 -5848
rect 3518 -5798 3594 -5786
rect 3518 -5850 3530 -5798
rect 3582 -5801 3594 -5798
rect 3702 -5801 3770 -5790
rect 3582 -5847 3713 -5801
rect 3759 -5847 3770 -5801
rect 3582 -5850 3594 -5847
rect 3518 -5862 3594 -5850
rect 3702 -5858 3770 -5847
rect 3905 -5791 3994 -5780
rect 3905 -5837 3937 -5791
rect 3983 -5837 3994 -5791
rect 3905 -5848 3994 -5837
rect 3341 -6365 3387 -6203
rect 3341 -6751 3387 -6589
rect 3341 -6986 3387 -6975
rect 3501 -5979 3547 -5968
rect 3501 -6365 3547 -6203
rect 3501 -6751 3547 -6589
rect 2253 -7170 3259 -7124
rect 3501 -7216 3547 -6975
rect 3745 -5979 3791 -5968
rect 3745 -6365 3791 -6203
rect 3745 -6751 3791 -6589
rect 3745 -7216 3791 -6975
rect 3905 -5979 3951 -5848
rect 4673 -5876 4719 -5754
rect 3905 -6365 3951 -6203
rect 3905 -6751 3951 -6589
rect 3905 -6986 3951 -6975
rect 4033 -5922 4719 -5876
rect 4033 -5979 4079 -5922
rect 4033 -6365 4079 -6203
rect 4033 -6751 4079 -6589
rect 4033 -7124 4079 -6975
rect 4193 -5979 4239 -5968
rect 4193 -6365 4239 -6203
rect 4193 -6751 4239 -6589
rect 4193 -7032 4239 -6975
rect 4353 -5979 4399 -5922
rect 4353 -6365 4399 -6203
rect 4353 -6751 4399 -6589
rect 4353 -6986 4399 -6975
rect 4513 -5979 4559 -5968
rect 4513 -6365 4559 -6203
rect 4513 -6751 4559 -6589
rect 4513 -7032 4559 -6975
rect 4673 -5979 4719 -5922
rect 4673 -6365 4719 -6203
rect 4673 -6751 4719 -6589
rect 4673 -6986 4719 -6975
rect 4833 -3905 4879 -3848
rect 4833 -4541 4879 -4379
rect 4833 -5177 4879 -5015
rect 4833 -5826 4879 -5651
rect 4993 -3848 5359 -3802
rect 4993 -3905 5039 -3848
rect 4993 -4541 5039 -4379
rect 4993 -5177 5039 -5015
rect 4993 -5662 5039 -5651
rect 5153 -3905 5199 -3894
rect 5153 -4541 5199 -4379
rect 5153 -5177 5199 -5015
rect 5153 -5826 5199 -5651
rect 5313 -3905 5359 -3848
rect 5313 -4541 5359 -4379
rect 5313 -5177 5359 -5015
rect 5557 -3848 5923 -3802
rect 5557 -3905 5603 -3848
rect 5557 -4541 5603 -4379
rect 5557 -5177 5603 -5015
rect 5359 -5651 5557 -5631
rect 5313 -5677 5603 -5651
rect 5717 -3905 5763 -3894
rect 5717 -4541 5763 -4379
rect 5717 -5177 5763 -5015
rect 5298 -5823 5374 -5811
rect 5298 -5826 5310 -5823
rect 4833 -5872 5310 -5826
rect 4833 -5979 4879 -5872
rect 4833 -6365 4879 -6203
rect 4833 -6751 4879 -6589
rect 4833 -7032 4879 -6975
rect 4193 -7078 4879 -7032
rect 4993 -5979 5039 -5968
rect 4993 -6365 5039 -6203
rect 4993 -6751 5039 -6589
rect 4993 -7032 5039 -6975
rect 5153 -5979 5199 -5872
rect 5298 -5875 5310 -5872
rect 5362 -5875 5374 -5823
rect 5298 -5887 5374 -5875
rect 5542 -5823 5618 -5811
rect 5542 -5875 5554 -5823
rect 5606 -5826 5618 -5823
rect 5717 -5826 5763 -5651
rect 5877 -3905 5923 -3848
rect 5877 -4541 5923 -4379
rect 5877 -5177 5923 -5015
rect 5877 -5662 5923 -5651
rect 6037 -3848 6723 -3802
rect 6037 -3905 6083 -3848
rect 6037 -4541 6083 -4379
rect 6037 -5177 6083 -5015
rect 6037 -5826 6083 -5651
rect 5606 -5872 6083 -5826
rect 5606 -5875 5618 -5872
rect 5542 -5887 5618 -5875
rect 5153 -6365 5199 -6203
rect 5153 -6751 5199 -6589
rect 5153 -6986 5199 -6975
rect 5313 -5979 5359 -5968
rect 5313 -6365 5359 -6203
rect 5313 -6751 5359 -6589
rect 5313 -7032 5359 -6975
rect 4993 -7078 5359 -7032
rect 5557 -5979 5603 -5968
rect 5557 -6365 5603 -6203
rect 5557 -6751 5603 -6589
rect 5557 -7032 5603 -6975
rect 5717 -5979 5763 -5872
rect 5717 -6365 5763 -6203
rect 5717 -6751 5763 -6589
rect 5717 -6986 5763 -6975
rect 5877 -5979 5923 -5968
rect 5877 -6365 5923 -6203
rect 5877 -6751 5923 -6589
rect 5877 -7032 5923 -6975
rect 5557 -7078 5923 -7032
rect 6037 -5979 6083 -5872
rect 6037 -6365 6083 -6203
rect 6037 -6751 6083 -6589
rect 6037 -7032 6083 -6975
rect 6197 -3905 6243 -3894
rect 6197 -4541 6243 -4379
rect 6197 -5177 6243 -5015
rect 6197 -5708 6243 -5651
rect 6357 -3905 6403 -3848
rect 6357 -4541 6403 -4379
rect 6357 -5177 6403 -5015
rect 6357 -5662 6403 -5651
rect 6517 -3905 6563 -3894
rect 6517 -4541 6563 -4379
rect 6517 -5177 6563 -5015
rect 6517 -5708 6563 -5651
rect 6677 -3905 6723 -3848
rect 6677 -4541 6723 -4379
rect 6677 -5177 6723 -5015
rect 6677 -5662 6723 -5651
rect 6837 -3905 6883 -3756
rect 6837 -4541 6883 -4379
rect 6837 -5177 6883 -5015
rect 6837 -5708 6883 -5651
rect 6197 -5754 6883 -5708
rect 6965 -3905 7011 -3894
rect 6965 -4541 7011 -4379
rect 6965 -5177 7011 -5015
rect 6197 -5876 6243 -5754
rect 6965 -5780 7011 -5651
rect 7125 -3905 7171 -3664
rect 7689 -3756 8695 -3710
rect 7689 -3802 7735 -3756
rect 7125 -4541 7171 -4379
rect 7125 -5177 7171 -5015
rect 7369 -3848 7735 -3802
rect 7369 -3905 7415 -3848
rect 7369 -4541 7415 -4379
rect 7369 -5177 7415 -5015
rect 7125 -5662 7171 -5651
rect 7261 -5651 7369 -5631
rect 7261 -5677 7415 -5651
rect 7529 -3905 7575 -3894
rect 7529 -4541 7575 -4379
rect 7529 -5177 7575 -5015
rect 6922 -5791 7011 -5780
rect 6922 -5837 6933 -5791
rect 6979 -5837 7011 -5791
rect 6922 -5848 7011 -5837
rect 6197 -5922 6883 -5876
rect 6197 -5979 6243 -5922
rect 6197 -6365 6243 -6203
rect 6197 -6751 6243 -6589
rect 6197 -6986 6243 -6975
rect 6357 -5979 6403 -5968
rect 6357 -6365 6403 -6203
rect 6357 -6751 6403 -6589
rect 6357 -7032 6403 -6975
rect 6517 -5979 6563 -5922
rect 6517 -6365 6563 -6203
rect 6517 -6751 6563 -6589
rect 6517 -6986 6563 -6975
rect 6677 -5979 6723 -5968
rect 6677 -6365 6723 -6203
rect 6677 -6751 6723 -6589
rect 6677 -7032 6723 -6975
rect 6037 -7078 6723 -7032
rect 6837 -5979 6883 -5922
rect 6837 -6365 6883 -6203
rect 6837 -6751 6883 -6589
rect 4993 -7124 5039 -7078
rect 4033 -7170 5039 -7124
rect 5877 -7124 5923 -7078
rect 6837 -7124 6883 -6975
rect 6965 -5979 7011 -5848
rect 7146 -5798 7214 -5790
rect 7146 -5850 7154 -5798
rect 7206 -5801 7214 -5798
rect 7206 -5847 7259 -5801
rect 7529 -5826 7575 -5651
rect 7689 -3905 7735 -3848
rect 7689 -4541 7735 -4379
rect 7689 -5177 7735 -5015
rect 7689 -5662 7735 -5651
rect 7849 -3848 8535 -3802
rect 7849 -3905 7895 -3848
rect 7849 -4541 7895 -4379
rect 7849 -5177 7895 -5015
rect 7849 -5811 7895 -5651
rect 8009 -3905 8055 -3894
rect 8009 -4541 8055 -4379
rect 8009 -5177 8055 -5015
rect 8009 -5708 8055 -5651
rect 8169 -3905 8215 -3848
rect 8169 -4541 8215 -4379
rect 8169 -5177 8215 -5015
rect 8169 -5662 8215 -5651
rect 8329 -3905 8375 -3894
rect 8329 -4541 8375 -4379
rect 8329 -5177 8375 -5015
rect 8329 -5708 8375 -5651
rect 8489 -3905 8535 -3848
rect 8489 -4541 8535 -4379
rect 8489 -5177 8535 -5015
rect 8489 -5662 8535 -5651
rect 8649 -3905 8695 -3756
rect 8649 -4541 8695 -4379
rect 8649 -5177 8695 -5015
rect 8649 -5708 8695 -5651
rect 8009 -5754 8695 -5708
rect 8777 -3905 8823 -3894
rect 8777 -4541 8823 -4379
rect 8777 -5177 8823 -5015
rect 7834 -5823 7910 -5811
rect 7834 -5826 7846 -5823
rect 7206 -5850 7214 -5847
rect 7146 -5858 7214 -5850
rect 7426 -5872 7846 -5826
rect 6965 -6365 7011 -6203
rect 6965 -6751 7011 -6589
rect 6965 -6986 7011 -6975
rect 7125 -5979 7171 -5968
rect 7125 -6365 7171 -6203
rect 7125 -6751 7171 -6589
rect 5877 -7170 6883 -7124
rect 7125 -7216 7171 -6975
rect 7369 -5979 7415 -5968
rect 7369 -6365 7415 -6203
rect 7369 -6751 7415 -6589
rect 7369 -7016 7415 -6975
rect 7529 -5979 7575 -5872
rect 7834 -5875 7846 -5872
rect 7898 -5875 7910 -5823
rect 7834 -5887 7910 -5875
rect 8009 -5876 8055 -5754
rect 8777 -5780 8823 -5651
rect 8937 -3905 8983 -3664
rect 8937 -4541 8983 -4379
rect 8937 -5177 8983 -5015
rect 8937 -5662 8983 -5651
rect 8734 -5791 8823 -5780
rect 8734 -5837 8745 -5791
rect 8791 -5837 8823 -5791
rect 8734 -5848 8823 -5837
rect 7529 -6365 7575 -6203
rect 7529 -6751 7575 -6589
rect 7529 -6986 7575 -6975
rect 7689 -5979 7735 -5968
rect 7689 -6365 7735 -6203
rect 7689 -6751 7735 -6589
rect 7354 -7028 7430 -7016
rect 7354 -7080 7366 -7028
rect 7418 -7032 7430 -7028
rect 7689 -7032 7735 -6975
rect 7418 -7078 7735 -7032
rect 7849 -5979 7895 -5887
rect 7849 -6365 7895 -6203
rect 7849 -6751 7895 -6589
rect 7849 -7032 7895 -6975
rect 8009 -5922 8695 -5876
rect 8009 -5979 8055 -5922
rect 8009 -6365 8055 -6203
rect 8009 -6751 8055 -6589
rect 8009 -6986 8055 -6975
rect 8169 -5979 8215 -5968
rect 8169 -6365 8215 -6203
rect 8169 -6751 8215 -6589
rect 8169 -7032 8215 -6975
rect 8329 -5979 8375 -5922
rect 8329 -6365 8375 -6203
rect 8329 -6751 8375 -6589
rect 8329 -6986 8375 -6975
rect 8489 -5979 8535 -5968
rect 8489 -6365 8535 -6203
rect 8489 -6751 8535 -6589
rect 8489 -7032 8535 -6975
rect 7849 -7078 8535 -7032
rect 8649 -5979 8695 -5922
rect 8649 -6365 8695 -6203
rect 8649 -6751 8695 -6589
rect 7418 -7080 7430 -7078
rect 7354 -7092 7430 -7080
rect 7689 -7124 7735 -7078
rect 8649 -7124 8695 -6975
rect 8777 -5979 8823 -5848
rect 8954 -5798 9030 -5786
rect 8954 -5850 8966 -5798
rect 9018 -5801 9030 -5798
rect 9018 -5847 9071 -5801
rect 9118 -5823 9194 -5811
rect 9018 -5850 9030 -5847
rect 8954 -5862 9030 -5850
rect 9118 -5875 9130 -5823
rect 9182 -5826 9194 -5823
rect 9182 -5872 9282 -5826
rect 9182 -5875 9194 -5872
rect 9118 -5887 9194 -5875
rect 8777 -6365 8823 -6203
rect 8777 -6751 8823 -6589
rect 8777 -6986 8823 -6975
rect 8937 -5979 8983 -5968
rect 8937 -6365 8983 -6203
rect 8937 -6751 8983 -6589
rect 7689 -7170 8695 -7124
rect 8937 -7216 8983 -6975
rect -4113 -7246 9020 -7216
rect -4113 -7249 -2188 -7246
rect -2136 -7249 -1682 -7246
rect -1630 -7249 855 -7246
rect 907 -7249 8197 -7246
rect 8249 -7249 9020 -7246
rect -4113 -7295 -4091 -7249
rect -4045 -7295 -3997 -7249
rect -3951 -7295 -3903 -7249
rect -3857 -7295 -3809 -7249
rect -3763 -7295 -3715 -7249
rect -3669 -7295 -3621 -7249
rect -3575 -7295 -3527 -7249
rect -3481 -7295 -3433 -7249
rect -3387 -7295 -3339 -7249
rect -3293 -7295 -3245 -7249
rect -3199 -7295 -3151 -7249
rect -3105 -7295 -3057 -7249
rect -3011 -7295 -2963 -7249
rect -2917 -7295 -2869 -7249
rect -2823 -7295 -2775 -7249
rect -2729 -7295 -2681 -7249
rect -2635 -7295 -2587 -7249
rect -2541 -7295 -2493 -7249
rect -2447 -7295 -2279 -7249
rect -2233 -7295 -2188 -7249
rect -2136 -7295 -2091 -7249
rect -2045 -7295 -1997 -7249
rect -1951 -7295 -1903 -7249
rect -1857 -7295 -1809 -7249
rect -1763 -7295 -1715 -7249
rect -1630 -7295 -1621 -7249
rect -1575 -7295 -1527 -7249
rect -1481 -7295 -1433 -7249
rect -1387 -7295 -1339 -7249
rect -1293 -7295 -1245 -7249
rect -1199 -7295 -1151 -7249
rect -1105 -7295 -1057 -7249
rect -1011 -7295 -963 -7249
rect -917 -7295 -869 -7249
rect -823 -7295 -775 -7249
rect -729 -7295 -681 -7249
rect -635 -7295 106 -7249
rect 152 -7295 200 -7249
rect 246 -7295 294 -7249
rect 340 -7295 388 -7249
rect 434 -7295 482 -7249
rect 528 -7295 576 -7249
rect 622 -7295 670 -7249
rect 716 -7295 764 -7249
rect 810 -7295 855 -7249
rect 907 -7295 952 -7249
rect 998 -7295 1046 -7249
rect 1092 -7295 1140 -7249
rect 1186 -7295 1234 -7249
rect 1280 -7295 1328 -7249
rect 1374 -7295 1422 -7249
rect 1468 -7295 1516 -7249
rect 1562 -7295 1610 -7249
rect 1656 -7295 1704 -7249
rect 1750 -7295 1918 -7249
rect 1964 -7295 2012 -7249
rect 2058 -7295 2106 -7249
rect 2152 -7295 2200 -7249
rect 2246 -7295 2294 -7249
rect 2340 -7295 2388 -7249
rect 2434 -7295 2482 -7249
rect 2528 -7295 2576 -7249
rect 2622 -7295 2670 -7249
rect 2716 -7295 2764 -7249
rect 2810 -7295 2858 -7249
rect 2904 -7295 2952 -7249
rect 2998 -7295 3046 -7249
rect 3092 -7295 3140 -7249
rect 3186 -7295 3234 -7249
rect 3280 -7295 3328 -7249
rect 3374 -7295 3422 -7249
rect 3468 -7295 3516 -7249
rect 3562 -7295 3730 -7249
rect 3776 -7295 3824 -7249
rect 3870 -7295 3918 -7249
rect 3964 -7295 4012 -7249
rect 4058 -7295 4106 -7249
rect 4152 -7295 4200 -7249
rect 4246 -7295 4294 -7249
rect 4340 -7295 4388 -7249
rect 4434 -7295 4482 -7249
rect 4528 -7295 4576 -7249
rect 4622 -7295 4670 -7249
rect 4716 -7295 4764 -7249
rect 4810 -7295 4858 -7249
rect 4904 -7295 4952 -7249
rect 4998 -7295 5046 -7249
rect 5092 -7295 5140 -7249
rect 5186 -7295 5234 -7249
rect 5280 -7295 5328 -7249
rect 5374 -7295 5542 -7249
rect 5588 -7295 5636 -7249
rect 5682 -7295 5730 -7249
rect 5776 -7295 5824 -7249
rect 5870 -7295 5918 -7249
rect 5964 -7295 6012 -7249
rect 6058 -7295 6106 -7249
rect 6152 -7295 6200 -7249
rect 6246 -7295 6294 -7249
rect 6340 -7295 6388 -7249
rect 6434 -7295 6482 -7249
rect 6528 -7295 6576 -7249
rect 6622 -7295 6670 -7249
rect 6716 -7295 6764 -7249
rect 6810 -7295 6858 -7249
rect 6904 -7295 6952 -7249
rect 6998 -7295 7046 -7249
rect 7092 -7295 7140 -7249
rect 7186 -7295 7354 -7249
rect 7400 -7295 7448 -7249
rect 7494 -7295 7542 -7249
rect 7588 -7295 7636 -7249
rect 7682 -7295 7730 -7249
rect 7776 -7295 7824 -7249
rect 7870 -7295 7918 -7249
rect 7964 -7295 8012 -7249
rect 8058 -7295 8106 -7249
rect 8152 -7295 8197 -7249
rect 8249 -7295 8294 -7249
rect 8340 -7295 8388 -7249
rect 8434 -7295 8482 -7249
rect 8528 -7295 8576 -7249
rect 8622 -7295 8670 -7249
rect 8716 -7295 8764 -7249
rect 8810 -7295 8858 -7249
rect 8904 -7295 8952 -7249
rect 8998 -7295 9020 -7249
rect -4113 -7298 -2188 -7295
rect -2136 -7298 -1682 -7295
rect -1630 -7298 855 -7295
rect 907 -7298 8197 -7295
rect 8249 -7298 9020 -7295
rect -4113 -7328 9020 -7298
<< via1 >>
rect 1238 7823 1290 7875
rect 3018 7715 3070 7767
rect 4830 7606 4882 7658
rect 6642 7499 6694 7551
rect 855 7407 907 7410
rect 8197 7407 8249 7410
rect 855 7361 858 7407
rect 858 7361 904 7407
rect 904 7361 907 7407
rect 8197 7361 8200 7407
rect 8200 7361 8246 7407
rect 8246 7361 8249 7407
rect 855 7358 907 7361
rect 8197 7358 8249 7361
rect 1238 7126 1290 7178
rect 1898 5959 1950 5962
rect 1898 5913 1901 5959
rect 1901 5913 1947 5959
rect 1947 5913 1950 5959
rect 1898 5910 1950 5913
rect 3018 7126 3070 7178
rect 1393 3834 1445 3886
rect 3710 5959 3762 5962
rect 3710 5913 3713 5959
rect 3713 5913 3759 5959
rect 3759 5913 3762 5959
rect 3710 5910 3762 5913
rect 4830 7126 4882 7178
rect 2223 3834 2275 3886
rect 5522 5959 5574 5962
rect 5522 5913 5525 5959
rect 5525 5913 5571 5959
rect 5571 5913 5574 5959
rect 5522 5910 5574 5913
rect 6642 7126 6694 7178
rect 4035 3834 4087 3886
rect 7334 5959 7386 5963
rect 7334 5913 7337 5959
rect 7337 5913 7383 5959
rect 7383 5913 7386 5959
rect 7334 5911 7386 5913
rect 5847 3834 5899 3886
rect 8934 7141 8986 7193
rect 8454 3926 8506 3978
rect 9098 5911 9150 5963
rect 9130 3926 9182 3978
rect -4452 3743 -4400 3746
rect -4452 3697 -4449 3743
rect -4449 3697 -4403 3743
rect -4403 3697 -4400 3743
rect -4452 3694 -4400 3697
rect -3720 3146 -3668 3148
rect -3720 3099 -3717 3146
rect -3717 3099 -3671 3146
rect -3671 3099 -3668 3146
rect -3720 3096 -3668 3099
rect -789 3096 -737 3148
rect -2749 2888 -2697 2891
rect -2185 2888 -2133 2891
rect -1682 2888 -1630 2891
rect -2749 2842 -2746 2888
rect -2746 2842 -2700 2888
rect -2700 2842 -2697 2888
rect -2185 2842 -2182 2888
rect -2182 2842 -2136 2888
rect -2136 2842 -2133 2888
rect -1682 2842 -1678 2888
rect -1678 2842 -1632 2888
rect -1632 2842 -1630 2888
rect -2749 2839 -2697 2842
rect -2185 2839 -2133 2842
rect -1682 2839 -1630 2842
rect -3720 2631 -3668 2633
rect -3720 2584 -3717 2631
rect -3717 2584 -3671 2631
rect -3671 2584 -3668 2631
rect -3720 2581 -3668 2584
rect -678 2581 -626 2633
rect -47 2581 5 2633
rect -169 2398 -117 2450
rect -4452 2033 -4400 2036
rect -4452 1987 -4449 2033
rect -4449 1987 -4403 2033
rect -4403 1987 -4400 2033
rect -4452 1984 -4400 1987
rect -3720 1436 -3668 1439
rect -3720 1389 -3717 1436
rect -3717 1389 -3671 1436
rect -3671 1389 -3668 1436
rect -3720 1387 -3668 1389
rect -2748 1178 -2696 1181
rect -2184 1178 -2132 1181
rect -1681 1178 -1629 1181
rect -2748 1132 -2746 1178
rect -2746 1132 -2700 1178
rect -2700 1132 -2696 1178
rect -2184 1132 -2182 1178
rect -2182 1132 -2136 1178
rect -2136 1132 -2132 1178
rect -1681 1132 -1678 1178
rect -1678 1132 -1632 1178
rect -1632 1132 -1629 1178
rect -2748 1129 -2696 1132
rect -2184 1129 -2132 1132
rect -1681 1129 -1629 1132
rect -3720 921 -3668 924
rect -3720 874 -3717 921
rect -3717 874 -3671 921
rect -3671 874 -3668 921
rect -3720 872 -3668 874
rect -291 1570 -239 1622
rect 1206 3462 1258 3514
rect -47 1478 5 1530
rect 86 1527 138 1530
rect 86 1481 89 1527
rect 89 1481 135 1527
rect 135 1481 138 1527
rect 86 1478 138 1481
rect -678 1387 -626 1439
rect -789 872 -737 924
rect -413 688 -361 740
rect -4452 323 -4400 326
rect -4452 277 -4449 323
rect -4449 277 -4403 323
rect -4403 277 -4400 323
rect -4452 274 -4400 277
rect -3720 -274 -3668 -272
rect -3720 -321 -3717 -274
rect -3717 -321 -3671 -274
rect -3671 -321 -3668 -274
rect -3720 -324 -3668 -321
rect 1686 1607 1738 1659
rect 2410 3462 2462 3514
rect 4190 3462 4242 3514
rect 3530 1527 3582 1530
rect 3530 1481 3533 1527
rect 3533 1481 3579 1527
rect 3579 1481 3582 1527
rect 3530 1478 3582 1481
rect 6034 3462 6086 3514
rect 5310 247 5362 299
rect 7361 3462 7413 3514
rect 7154 1527 7206 1530
rect 7154 1481 7157 1527
rect 7157 1481 7203 1527
rect 7203 1481 7206 1527
rect 7154 1478 7206 1481
rect 7846 1453 7898 1505
rect 8966 1527 9018 1530
rect 8966 1481 8969 1527
rect 8969 1481 9015 1527
rect 9015 1481 9018 1527
rect 8966 1478 9018 1481
rect 9130 1453 9182 1505
rect 855 79 907 82
rect 8197 79 8249 82
rect 855 33 858 79
rect 858 33 904 79
rect 904 33 907 79
rect 8197 33 8200 79
rect 8200 33 8246 79
rect 8246 33 8249 79
rect 855 30 907 33
rect 8197 30 8249 33
rect -789 -324 -737 -272
rect -2748 -532 -2696 -529
rect -2184 -532 -2132 -529
rect -1681 -532 -1629 -529
rect -2748 -578 -2746 -532
rect -2746 -578 -2700 -532
rect -2700 -578 -2696 -532
rect -2184 -578 -2182 -532
rect -2182 -578 -2136 -532
rect -2136 -578 -2132 -532
rect -1681 -578 -1678 -532
rect -1678 -578 -1632 -532
rect -1632 -578 -1629 -532
rect -2748 -581 -2696 -578
rect -2184 -581 -2132 -578
rect -1681 -581 -1629 -578
rect -3720 -789 -3668 -787
rect -3720 -836 -3717 -789
rect -3717 -836 -3671 -789
rect -3671 -836 -3668 -789
rect -3720 -839 -3668 -836
rect -678 -839 -626 -787
rect -535 -1022 -483 -970
rect 86 -1369 138 -1366
rect -4452 -1387 -4400 -1384
rect -3953 -1387 -3901 -1384
rect -3653 -1387 -3601 -1384
rect -3353 -1387 -3301 -1384
rect -3053 -1387 -3001 -1384
rect -2753 -1387 -2701 -1384
rect -4452 -1433 -4449 -1387
rect -4449 -1433 -4403 -1387
rect -4403 -1433 -4400 -1387
rect -3953 -1433 -3933 -1387
rect -3933 -1433 -3901 -1387
rect -3653 -1433 -3651 -1387
rect -3651 -1433 -3601 -1387
rect -3353 -1433 -3335 -1387
rect -3335 -1433 -3301 -1387
rect -3053 -1433 -3005 -1387
rect -3005 -1433 -3001 -1387
rect -2753 -1433 -2737 -1387
rect -2737 -1433 -2701 -1387
rect 86 -1415 89 -1369
rect 89 -1415 135 -1369
rect 135 -1415 138 -1369
rect 86 -1418 138 -1415
rect 566 -202 618 -150
rect -4452 -1436 -4400 -1433
rect -3953 -1436 -3901 -1433
rect -3653 -1436 -3601 -1433
rect -3353 -1436 -3301 -1433
rect -3053 -1436 -3001 -1433
rect -2753 -1436 -2701 -1433
rect 1930 -3417 1982 -3365
rect 3050 -202 3102 -150
rect 3530 -1369 3582 -1366
rect 3530 -1415 3533 -1369
rect 3533 -1415 3579 -1369
rect 3579 -1415 3582 -1369
rect 3530 -1418 3582 -1415
rect 4830 -202 4882 -150
rect 5554 -3417 5606 -3365
rect 6674 -202 6726 -150
rect 7361 -202 7413 -150
rect 7154 -1369 7206 -1366
rect 7154 -1415 7157 -1369
rect 7157 -1415 7203 -1369
rect 7203 -1415 7206 -1369
rect 7154 -1418 7206 -1415
rect 7846 -1393 7898 -1341
rect 8966 -1369 9018 -1366
rect 8966 -1415 8969 -1369
rect 8969 -1415 9015 -1369
rect 9015 -1415 9018 -1369
rect 9130 -1393 9182 -1341
rect 8966 -1418 9018 -1415
rect -3953 -3585 -3901 -3582
rect -3653 -3585 -3601 -3582
rect -3353 -3585 -3301 -3582
rect -3053 -3585 -3001 -3582
rect -2753 -3585 -2701 -3582
rect -3953 -3631 -3950 -3585
rect -3950 -3631 -3904 -3585
rect -3904 -3631 -3901 -3585
rect -3653 -3631 -3622 -3585
rect -3622 -3631 -3601 -3585
rect -3353 -3631 -3340 -3585
rect -3340 -3631 -3301 -3585
rect -3053 -3631 -3010 -3585
rect -3010 -3631 -3001 -3585
rect -2753 -3631 -2728 -3585
rect -2728 -3631 -2701 -3585
rect -3953 -3634 -3901 -3631
rect -3653 -3634 -3601 -3631
rect -3353 -3634 -3301 -3631
rect -3053 -3634 -3001 -3631
rect -2753 -3634 -2701 -3631
rect -4273 -3851 -4221 -3799
rect -4111 -5801 -4059 -5798
rect -4111 -5847 -4108 -5801
rect -4108 -5847 -4062 -5801
rect -4062 -5847 -4059 -5801
rect -4111 -5850 -4059 -5847
rect -2511 -3851 -2459 -3799
rect -2991 -7066 -2939 -7014
rect -1147 -3866 -1095 -3814
rect -667 -5801 -615 -5798
rect -667 -5847 -664 -5801
rect -664 -5847 -618 -5801
rect -618 -5847 -615 -5801
rect -667 -5850 -615 -5847
rect -291 -5850 -239 -5798
rect 86 -5801 138 -5798
rect 86 -5847 89 -5801
rect 89 -5847 135 -5801
rect 135 -5847 138 -5801
rect 86 -5850 138 -5847
rect 401 -7066 453 -7014
rect 1686 -5875 1738 -5823
rect 1930 -5875 1982 -5823
rect 4025 -3866 4077 -3814
rect 3530 -5801 3582 -5798
rect 3530 -5847 3533 -5801
rect 3533 -5847 3579 -5801
rect 3579 -5847 3582 -5801
rect 3530 -5850 3582 -5847
rect 5310 -5875 5362 -5823
rect 5554 -5875 5606 -5823
rect 7154 -5801 7206 -5798
rect 7154 -5847 7157 -5801
rect 7157 -5847 7203 -5801
rect 7203 -5847 7206 -5801
rect 7154 -5850 7206 -5847
rect 7846 -5875 7898 -5823
rect 7366 -7080 7418 -7028
rect 8966 -5801 9018 -5798
rect 8966 -5847 8969 -5801
rect 8969 -5847 9015 -5801
rect 9015 -5847 9018 -5801
rect 8966 -5850 9018 -5847
rect 9130 -5875 9182 -5823
rect -2188 -7249 -2136 -7246
rect -1682 -7249 -1630 -7246
rect 855 -7249 907 -7246
rect 8197 -7249 8249 -7246
rect -2188 -7295 -2185 -7249
rect -2185 -7295 -2139 -7249
rect -2139 -7295 -2136 -7249
rect -1682 -7295 -1669 -7249
rect -1669 -7295 -1630 -7249
rect 855 -7295 858 -7249
rect 858 -7295 904 -7249
rect 904 -7295 907 -7249
rect 8197 -7295 8200 -7249
rect 8200 -7295 8246 -7249
rect 8246 -7295 8249 -7249
rect -2188 -7298 -2136 -7295
rect -1682 -7298 -1630 -7295
rect 855 -7298 907 -7295
rect 8197 -7298 8249 -7295
<< metal2 >>
rect 1226 7875 1302 7887
rect 1226 7823 1238 7875
rect 1290 7823 1302 7875
rect 1226 7811 1302 7823
rect 825 7410 937 7440
rect 825 7358 855 7410
rect 907 7358 937 7410
rect 554 7195 630 7205
rect 554 7139 564 7195
rect 620 7139 630 7195
rect 554 7129 630 7139
rect -4464 3746 -4388 3758
rect -4464 3694 -4452 3746
rect -4400 3694 -4388 3746
rect -4464 3682 -4388 3694
rect -4454 2048 -4398 3682
rect -3732 3150 -3656 3160
rect -801 3150 -725 3160
rect -3732 3148 -725 3150
rect -3732 3096 -3720 3148
rect -3668 3096 -789 3148
rect -737 3096 -725 3148
rect -3732 3094 -725 3096
rect -3732 3084 -3656 3094
rect -801 3084 -725 3094
rect -2761 2893 -2685 2903
rect -2761 2837 -2751 2893
rect -2695 2837 -2685 2893
rect -2761 2827 -2685 2837
rect -2197 2893 -2121 2903
rect -2197 2837 -2187 2893
rect -2131 2837 -2121 2893
rect -2197 2827 -2121 2837
rect -1694 2893 -1618 2903
rect -1694 2837 -1684 2893
rect -1628 2837 -1618 2893
rect -1694 2827 -1618 2837
rect -3732 2635 -3656 2645
rect -690 2635 -614 2645
rect -3732 2633 -614 2635
rect -3732 2581 -3720 2633
rect -3668 2581 -678 2633
rect -626 2581 -614 2633
rect -3732 2579 -614 2581
rect -3732 2569 -3656 2579
rect -690 2569 -614 2579
rect -59 2633 17 2645
rect -59 2581 -47 2633
rect 5 2581 17 2633
rect -59 2569 17 2581
rect -181 2450 -105 2462
rect -181 2398 -169 2450
rect -117 2398 -105 2450
rect -181 2386 -105 2398
rect -4464 2036 -4388 2048
rect -4464 1984 -4452 2036
rect -4400 1984 -4388 2036
rect -4464 1972 -4388 1984
rect -4454 338 -4398 1972
rect -303 1622 -227 1634
rect -303 1570 -291 1622
rect -239 1570 -227 1622
rect -303 1558 -227 1570
rect -3732 1441 -3656 1451
rect -690 1441 -614 1451
rect -3732 1439 -614 1441
rect -3732 1387 -3720 1439
rect -3668 1387 -678 1439
rect -626 1387 -614 1439
rect -3732 1385 -614 1387
rect -3732 1375 -3656 1385
rect -690 1375 -614 1385
rect -2760 1183 -2684 1193
rect -2760 1127 -2750 1183
rect -2694 1127 -2684 1183
rect -2760 1117 -2684 1127
rect -2196 1183 -2120 1193
rect -2196 1127 -2186 1183
rect -2130 1127 -2120 1183
rect -2196 1117 -2120 1127
rect -1693 1183 -1617 1193
rect -1693 1127 -1683 1183
rect -1627 1127 -1617 1183
rect -1693 1117 -1617 1127
rect -3732 926 -3656 936
rect -801 926 -725 936
rect -3732 924 -725 926
rect -3732 872 -3720 924
rect -3668 872 -789 924
rect -737 872 -725 924
rect -3732 870 -725 872
rect -3732 860 -3656 870
rect -801 860 -725 870
rect -425 740 -349 752
rect -425 688 -413 740
rect -361 688 -349 740
rect -425 676 -349 688
rect -4464 326 -4388 338
rect -4464 274 -4452 326
rect -4400 274 -4388 326
rect -4464 262 -4388 274
rect -4454 -1372 -4398 262
rect -3732 -270 -3656 -260
rect -801 -270 -725 -260
rect -3732 -272 -725 -270
rect -3732 -324 -3720 -272
rect -3668 -324 -789 -272
rect -737 -324 -725 -272
rect -3732 -326 -725 -324
rect -3732 -336 -3656 -326
rect -801 -336 -725 -326
rect -2760 -527 -2684 -517
rect -2760 -583 -2750 -527
rect -2694 -583 -2684 -527
rect -2760 -593 -2684 -583
rect -2196 -527 -2120 -517
rect -2196 -583 -2186 -527
rect -2130 -583 -2120 -527
rect -2196 -593 -2120 -583
rect -1693 -527 -1617 -517
rect -1693 -583 -1683 -527
rect -1627 -583 -1617 -527
rect -1693 -593 -1617 -583
rect -3732 -785 -3656 -775
rect -690 -776 -614 -775
rect -690 -785 -613 -776
rect -3732 -787 -613 -785
rect -3732 -839 -3720 -787
rect -3668 -839 -678 -787
rect -626 -839 -613 -787
rect -3732 -841 -613 -839
rect -3732 -851 -3656 -841
rect -690 -851 -613 -841
rect -4464 -1384 -4388 -1372
rect -4464 -1436 -4452 -1384
rect -4400 -1436 -4388 -1384
rect -4464 -1448 -4388 -1436
rect -3983 -1384 -3871 -1374
rect -3983 -1436 -3953 -1384
rect -3901 -1436 -3871 -1384
rect -3983 -3582 -3871 -1436
rect -3983 -3634 -3953 -3582
rect -3901 -3634 -3871 -3582
rect -3983 -3646 -3871 -3634
rect -3683 -1384 -3571 -1374
rect -3683 -1436 -3653 -1384
rect -3601 -1436 -3571 -1384
rect -3683 -3582 -3571 -1436
rect -3683 -3634 -3653 -3582
rect -3601 -3634 -3571 -3582
rect -3683 -3646 -3571 -3634
rect -3383 -1384 -3271 -1374
rect -3383 -1436 -3353 -1384
rect -3301 -1436 -3271 -1384
rect -3383 -3582 -3271 -1436
rect -3383 -3634 -3353 -3582
rect -3301 -3634 -3271 -3582
rect -3383 -3646 -3271 -3634
rect -3083 -1384 -2971 -1374
rect -3083 -1436 -3053 -1384
rect -3001 -1436 -2971 -1384
rect -3083 -3582 -2971 -1436
rect -3083 -3634 -3053 -3582
rect -3001 -3634 -2971 -3582
rect -3083 -3646 -2971 -3634
rect -2783 -1384 -2671 -1374
rect -2783 -1436 -2753 -1384
rect -2701 -1436 -2671 -1384
rect -2783 -3582 -2671 -1436
rect -2783 -3634 -2753 -3582
rect -2701 -3634 -2671 -3582
rect -2783 -3646 -2671 -3634
rect -2215 -2849 -2103 -2841
rect -2215 -2905 -2187 -2849
rect -2131 -2905 -2103 -2849
rect -2215 -2953 -2103 -2905
rect -2215 -3009 -2187 -2953
rect -2131 -3009 -2103 -2953
rect -4285 -3797 -4209 -3787
rect -4285 -3853 -4275 -3797
rect -4219 -3853 -4209 -3797
rect -4285 -3863 -4209 -3853
rect -2523 -3797 -2447 -3787
rect -2523 -3853 -2513 -3797
rect -2457 -3853 -2447 -3797
rect -2523 -3863 -2447 -3853
rect -4123 -5796 -4047 -5786
rect -4123 -5852 -4113 -5796
rect -4057 -5852 -4047 -5796
rect -4123 -5862 -4047 -5852
rect -3003 -7012 -2927 -7002
rect -3003 -7068 -2993 -7012
rect -2937 -7068 -2927 -7012
rect -3003 -7078 -2927 -7068
rect -2215 -7246 -2103 -3009
rect -2215 -7298 -2188 -7246
rect -2136 -7298 -2103 -7246
rect -2215 -7328 -2103 -7298
rect -1712 -2849 -1600 -2840
rect -1712 -2905 -1684 -2849
rect -1628 -2905 -1600 -2849
rect -1712 -2953 -1600 -2905
rect -1712 -3009 -1684 -2953
rect -1628 -3009 -1600 -2953
rect -1712 -7246 -1600 -3009
rect -1159 -3812 -1083 -3802
rect -1159 -3868 -1149 -3812
rect -1093 -3868 -1083 -3812
rect -1159 -3878 -1083 -3868
rect -669 -5786 -613 -851
rect -547 -970 -471 -958
rect -547 -1022 -535 -970
rect -483 -1022 -471 -970
rect -547 -1034 -471 -1022
rect -537 -5786 -481 -1034
rect -415 -3245 -359 676
rect -425 -3255 -349 -3245
rect -425 -3311 -415 -3255
rect -359 -3311 -349 -3255
rect -425 -3321 -349 -3311
rect -293 -5786 -237 1558
rect -171 -1354 -115 2386
rect -49 1542 7 2569
rect -59 1530 17 1542
rect -59 1478 -47 1530
rect 5 1478 17 1530
rect -59 1466 17 1478
rect 74 1532 150 1542
rect 74 1476 84 1532
rect 140 1476 150 1532
rect 74 1466 150 1476
rect 84 -1354 140 1466
rect 564 -138 620 7129
rect 825 82 937 7358
rect 1236 7190 1292 7811
rect 3006 7767 3082 7779
rect 3006 7715 3018 7767
rect 3070 7715 3082 7767
rect 3006 7703 3082 7715
rect 3016 7190 3072 7703
rect 4818 7658 4894 7670
rect 4818 7606 4830 7658
rect 4882 7606 4894 7658
rect 4818 7594 4894 7606
rect 4828 7190 4884 7594
rect 6630 7551 6706 7563
rect 6630 7499 6642 7551
rect 6694 7499 6706 7551
rect 6630 7487 6706 7499
rect 6640 7190 6696 7487
rect 8167 7410 8279 7440
rect 8167 7358 8197 7410
rect 8249 7358 8279 7410
rect 1226 7178 1302 7190
rect 1226 7126 1238 7178
rect 1290 7126 1302 7178
rect 1226 7114 1302 7126
rect 3006 7178 3082 7190
rect 3006 7126 3018 7178
rect 3070 7126 3082 7178
rect 3006 7114 3082 7126
rect 4818 7178 4894 7190
rect 4818 7126 4830 7178
rect 4882 7126 4894 7178
rect 4818 7114 4894 7126
rect 6630 7178 6706 7190
rect 6630 7126 6642 7178
rect 6694 7126 6706 7178
rect 6630 7114 6706 7126
rect 1886 5964 1962 5974
rect 1886 5908 1896 5964
rect 1952 5908 1962 5964
rect 1886 5898 1962 5908
rect 3698 5964 3774 5974
rect 3698 5908 3708 5964
rect 3764 5908 3774 5964
rect 3698 5898 3774 5908
rect 5510 5964 5586 5974
rect 5510 5908 5520 5964
rect 5576 5908 5586 5964
rect 5510 5898 5586 5908
rect 7322 5965 7398 5975
rect 7322 5909 7332 5965
rect 7388 5909 7398 5965
rect 7322 5899 7398 5909
rect 1381 3888 1457 3898
rect 1204 3886 1457 3888
rect 1204 3834 1393 3886
rect 1445 3834 1457 3886
rect 1204 3832 1457 3834
rect 1204 3526 1260 3832
rect 1381 3822 1457 3832
rect 2211 3888 2287 3898
rect 4023 3888 4099 3898
rect 4818 3888 4894 3898
rect 2211 3886 2464 3888
rect 2211 3834 2223 3886
rect 2275 3834 2464 3886
rect 2211 3832 2464 3834
rect 2211 3822 2287 3832
rect 2408 3526 2464 3832
rect 4023 3886 4244 3888
rect 4023 3834 4035 3886
rect 4087 3834 4244 3886
rect 4023 3832 4244 3834
rect 4023 3822 4099 3832
rect 4188 3526 4244 3832
rect 4818 3832 4828 3888
rect 4884 3832 4894 3888
rect 4818 3822 4894 3832
rect 5835 3888 5911 3898
rect 5835 3832 5845 3888
rect 5901 3832 5911 3888
rect 5835 3822 5911 3832
rect 1194 3514 1270 3526
rect 1194 3462 1206 3514
rect 1258 3462 1270 3514
rect 1194 3450 1270 3462
rect 2398 3514 2474 3526
rect 2398 3462 2410 3514
rect 2462 3462 2474 3514
rect 2398 3450 2474 3462
rect 4178 3514 4254 3526
rect 4178 3462 4190 3514
rect 4242 3462 4254 3514
rect 4178 3450 4254 3462
rect 1674 1659 1750 1671
rect 1674 1607 1686 1659
rect 1738 1607 1750 1659
rect 1674 1595 1750 1607
rect 825 30 855 82
rect 907 30 937 82
rect 554 -150 630 -138
rect 554 -202 566 -150
rect 618 -202 630 -150
rect 554 -214 630 -202
rect -181 -1364 -105 -1354
rect -181 -1420 -171 -1364
rect -115 -1420 -105 -1364
rect -181 -1430 -105 -1420
rect 74 -1366 150 -1354
rect 74 -1418 86 -1366
rect 138 -1418 150 -1366
rect 74 -1430 150 -1418
rect -679 -5798 -603 -5786
rect -679 -5850 -667 -5798
rect -615 -5850 -603 -5798
rect -679 -5862 -603 -5850
rect -547 -5796 -471 -5786
rect -547 -5852 -537 -5796
rect -481 -5852 -471 -5796
rect -547 -5862 -471 -5852
rect -303 -5798 -227 -5786
rect -303 -5850 -291 -5798
rect -239 -5850 -227 -5798
rect -303 -5862 -227 -5850
rect 74 -5796 150 -5786
rect 74 -5852 84 -5796
rect 140 -5852 150 -5796
rect 74 -5862 150 -5852
rect 389 -7012 465 -7002
rect 389 -7068 399 -7012
rect 455 -7068 465 -7012
rect 389 -7078 465 -7068
rect -1712 -7298 -1682 -7246
rect -1630 -7298 -1600 -7246
rect -1712 -7328 -1600 -7298
rect 825 -7246 937 30
rect 1684 -5811 1740 1595
rect 3518 1530 3594 1542
rect 3518 1478 3530 1530
rect 3582 1478 3594 1530
rect 3518 1466 3594 1478
rect 3038 -150 3114 -138
rect 3038 -202 3050 -150
rect 3102 -202 3114 -150
rect 3038 -214 3114 -202
rect 1918 -3365 1994 -3353
rect 1918 -3417 1930 -3365
rect 1982 -3417 1994 -3365
rect 1918 -3429 1994 -3417
rect 1928 -5811 1984 -3429
rect 1674 -5823 1750 -5811
rect 1674 -5875 1686 -5823
rect 1738 -5875 1750 -5823
rect 1674 -5887 1750 -5875
rect 1918 -5823 1994 -5811
rect 1918 -5875 1930 -5823
rect 1982 -5875 1994 -5823
rect 1918 -5887 1994 -5875
rect 3048 -7016 3104 -214
rect 3528 -1354 3584 1466
rect 4828 -138 4884 3822
rect 6022 3516 6098 3526
rect 6022 3460 6032 3516
rect 6088 3460 6098 3516
rect 6022 3450 6098 3460
rect 7349 3516 7425 3526
rect 7349 3460 7359 3516
rect 7415 3460 7425 3516
rect 7349 3450 7425 3460
rect 7142 1532 7218 1542
rect 7142 1476 7152 1532
rect 7208 1476 7218 1532
rect 7142 1466 7218 1476
rect 7834 1507 7910 1517
rect 5298 299 5374 311
rect 5298 247 5310 299
rect 5362 247 5374 299
rect 5298 235 5374 247
rect 4818 -150 4894 -138
rect 4818 -202 4830 -150
rect 4882 -202 4894 -150
rect 4818 -214 4894 -202
rect 3518 -1364 3594 -1354
rect 3518 -1420 3528 -1364
rect 3584 -1420 3594 -1364
rect 3518 -1430 3594 -1420
rect 3518 -3255 3594 -3245
rect 3518 -3311 3528 -3255
rect 3584 -3311 3594 -3255
rect 3518 -3321 3594 -3311
rect 3528 -5786 3584 -3321
rect 4013 -3812 4089 -3802
rect 4013 -3868 4023 -3812
rect 4079 -3868 4089 -3812
rect 4013 -3878 4089 -3868
rect 3518 -5798 3594 -5786
rect 3518 -5850 3530 -5798
rect 3582 -5850 3594 -5798
rect 5308 -5811 5364 235
rect 6662 -148 6738 -138
rect 6662 -204 6672 -148
rect 6728 -204 6738 -148
rect 6662 -214 6738 -204
rect 7152 -1354 7208 1466
rect 7834 1451 7844 1507
rect 7900 1451 7910 1507
rect 7834 1441 7910 1451
rect 8167 82 8279 7358
rect 8922 7195 8998 7205
rect 8922 7139 8932 7195
rect 8988 7139 8998 7195
rect 8922 7129 8998 7139
rect 8954 5965 9030 5975
rect 8954 5909 8964 5965
rect 9020 5909 9030 5965
rect 8954 5899 9030 5909
rect 9086 5965 9162 5975
rect 9086 5909 9096 5965
rect 9152 5909 9162 5965
rect 9086 5899 9162 5909
rect 8442 3980 8518 3990
rect 8442 3924 8452 3980
rect 8508 3924 8518 3980
rect 8442 3914 8518 3924
rect 8964 1542 9020 5899
rect 9118 3980 9194 3990
rect 9118 3924 9128 3980
rect 9184 3924 9194 3980
rect 9118 3914 9194 3924
rect 8954 1530 9030 1542
rect 8954 1478 8966 1530
rect 9018 1478 9030 1530
rect 8954 1466 9030 1478
rect 9118 1507 9194 1517
rect 8167 30 8197 82
rect 8249 30 8279 82
rect 7349 -148 7425 -138
rect 7349 -204 7359 -148
rect 7415 -204 7425 -148
rect 7349 -214 7425 -204
rect 7834 -1339 7910 -1329
rect 7142 -1366 7218 -1354
rect 7142 -1418 7154 -1366
rect 7206 -1418 7218 -1366
rect 7834 -1395 7844 -1339
rect 7900 -1395 7910 -1339
rect 7834 -1405 7910 -1395
rect 7142 -1430 7218 -1418
rect 5542 -3365 5618 -3353
rect 5542 -3417 5554 -3365
rect 5606 -3417 5618 -3365
rect 5542 -3429 5618 -3417
rect 5552 -5811 5608 -3429
rect 7142 -5796 7218 -5786
rect 3518 -5862 3594 -5850
rect 5298 -5823 5374 -5811
rect 5298 -5875 5310 -5823
rect 5362 -5875 5374 -5823
rect 5298 -5887 5374 -5875
rect 5542 -5823 5618 -5811
rect 5542 -5875 5554 -5823
rect 5606 -5875 5618 -5823
rect 7142 -5852 7152 -5796
rect 7208 -5852 7218 -5796
rect 7142 -5862 7218 -5852
rect 7834 -5821 7910 -5811
rect 5542 -5887 5618 -5875
rect 7834 -5877 7844 -5821
rect 7900 -5877 7910 -5821
rect 7834 -5887 7910 -5877
rect 3038 -7026 3114 -7016
rect 3038 -7082 3048 -7026
rect 3104 -7082 3114 -7026
rect 3038 -7092 3114 -7082
rect 7354 -7026 7430 -7016
rect 7354 -7082 7364 -7026
rect 7420 -7082 7430 -7026
rect 7354 -7092 7430 -7082
rect 825 -7298 855 -7246
rect 907 -7298 937 -7246
rect 825 -7328 937 -7298
rect 8167 -7246 8279 30
rect 8964 -1354 9020 1466
rect 9118 1451 9128 1507
rect 9184 1451 9194 1507
rect 9118 1441 9194 1451
rect 9118 -1339 9194 -1329
rect 8954 -1366 9030 -1354
rect 8954 -1418 8966 -1366
rect 9018 -1418 9030 -1366
rect 9118 -1395 9128 -1339
rect 9184 -1395 9194 -1339
rect 9118 -1405 9194 -1395
rect 8954 -1430 9030 -1418
rect 8964 -5786 9020 -1430
rect 8954 -5798 9030 -5786
rect 8954 -5850 8966 -5798
rect 9018 -5850 9030 -5798
rect 8954 -5862 9030 -5850
rect 9118 -5821 9194 -5811
rect 9118 -5877 9128 -5821
rect 9184 -5877 9194 -5821
rect 9118 -5887 9194 -5877
rect 8167 -7298 8197 -7246
rect 8249 -7298 8279 -7246
rect 8167 -7328 8279 -7298
<< via2 >>
rect 564 7139 620 7195
rect -2751 2891 -2695 2893
rect -2751 2839 -2749 2891
rect -2749 2839 -2697 2891
rect -2697 2839 -2695 2891
rect -2751 2837 -2695 2839
rect -2187 2891 -2131 2893
rect -2187 2839 -2185 2891
rect -2185 2839 -2133 2891
rect -2133 2839 -2131 2891
rect -2187 2837 -2131 2839
rect -1684 2891 -1628 2893
rect -1684 2839 -1682 2891
rect -1682 2839 -1630 2891
rect -1630 2839 -1628 2891
rect -1684 2837 -1628 2839
rect -2750 1181 -2694 1183
rect -2750 1129 -2748 1181
rect -2748 1129 -2696 1181
rect -2696 1129 -2694 1181
rect -2750 1127 -2694 1129
rect -2186 1181 -2130 1183
rect -2186 1129 -2184 1181
rect -2184 1129 -2132 1181
rect -2132 1129 -2130 1181
rect -2186 1127 -2130 1129
rect -1683 1181 -1627 1183
rect -1683 1129 -1681 1181
rect -1681 1129 -1629 1181
rect -1629 1129 -1627 1181
rect -1683 1127 -1627 1129
rect -2750 -529 -2694 -527
rect -2750 -581 -2748 -529
rect -2748 -581 -2696 -529
rect -2696 -581 -2694 -529
rect -2750 -583 -2694 -581
rect -2186 -529 -2130 -527
rect -2186 -581 -2184 -529
rect -2184 -581 -2132 -529
rect -2132 -581 -2130 -529
rect -2186 -583 -2130 -581
rect -1683 -529 -1627 -527
rect -1683 -581 -1681 -529
rect -1681 -581 -1629 -529
rect -1629 -581 -1627 -529
rect -1683 -583 -1627 -581
rect -2187 -2905 -2131 -2849
rect -2187 -3009 -2131 -2953
rect -4275 -3799 -4219 -3797
rect -4275 -3851 -4273 -3799
rect -4273 -3851 -4221 -3799
rect -4221 -3851 -4219 -3799
rect -4275 -3853 -4219 -3851
rect -2513 -3799 -2457 -3797
rect -2513 -3851 -2511 -3799
rect -2511 -3851 -2459 -3799
rect -2459 -3851 -2457 -3799
rect -2513 -3853 -2457 -3851
rect -4113 -5798 -4057 -5796
rect -4113 -5850 -4111 -5798
rect -4111 -5850 -4059 -5798
rect -4059 -5850 -4057 -5798
rect -4113 -5852 -4057 -5850
rect -2993 -7014 -2937 -7012
rect -2993 -7066 -2991 -7014
rect -2991 -7066 -2939 -7014
rect -2939 -7066 -2937 -7014
rect -2993 -7068 -2937 -7066
rect -1684 -2905 -1628 -2849
rect -1684 -3009 -1628 -2953
rect -1149 -3814 -1093 -3812
rect -1149 -3866 -1147 -3814
rect -1147 -3866 -1095 -3814
rect -1095 -3866 -1093 -3814
rect -1149 -3868 -1093 -3866
rect -415 -3311 -359 -3255
rect 84 1530 140 1532
rect 84 1478 86 1530
rect 86 1478 138 1530
rect 138 1478 140 1530
rect 84 1476 140 1478
rect 1896 5962 1952 5964
rect 1896 5910 1898 5962
rect 1898 5910 1950 5962
rect 1950 5910 1952 5962
rect 1896 5908 1952 5910
rect 3708 5962 3764 5964
rect 3708 5910 3710 5962
rect 3710 5910 3762 5962
rect 3762 5910 3764 5962
rect 3708 5908 3764 5910
rect 5520 5962 5576 5964
rect 5520 5910 5522 5962
rect 5522 5910 5574 5962
rect 5574 5910 5576 5962
rect 5520 5908 5576 5910
rect 7332 5963 7388 5965
rect 7332 5911 7334 5963
rect 7334 5911 7386 5963
rect 7386 5911 7388 5963
rect 7332 5909 7388 5911
rect 4828 3832 4884 3888
rect 5845 3886 5901 3888
rect 5845 3834 5847 3886
rect 5847 3834 5899 3886
rect 5899 3834 5901 3886
rect 5845 3832 5901 3834
rect -171 -1420 -115 -1364
rect -537 -5852 -481 -5796
rect 84 -5798 140 -5796
rect 84 -5850 86 -5798
rect 86 -5850 138 -5798
rect 138 -5850 140 -5798
rect 84 -5852 140 -5850
rect 399 -7014 455 -7012
rect 399 -7066 401 -7014
rect 401 -7066 453 -7014
rect 453 -7066 455 -7014
rect 399 -7068 455 -7066
rect 6032 3514 6088 3516
rect 6032 3462 6034 3514
rect 6034 3462 6086 3514
rect 6086 3462 6088 3514
rect 6032 3460 6088 3462
rect 7359 3514 7415 3516
rect 7359 3462 7361 3514
rect 7361 3462 7413 3514
rect 7413 3462 7415 3514
rect 7359 3460 7415 3462
rect 7152 1530 7208 1532
rect 7152 1478 7154 1530
rect 7154 1478 7206 1530
rect 7206 1478 7208 1530
rect 7152 1476 7208 1478
rect 3528 -1366 3584 -1364
rect 3528 -1418 3530 -1366
rect 3530 -1418 3582 -1366
rect 3582 -1418 3584 -1366
rect 3528 -1420 3584 -1418
rect 3528 -3311 3584 -3255
rect 4023 -3814 4079 -3812
rect 4023 -3866 4025 -3814
rect 4025 -3866 4077 -3814
rect 4077 -3866 4079 -3814
rect 4023 -3868 4079 -3866
rect 6672 -150 6728 -148
rect 6672 -202 6674 -150
rect 6674 -202 6726 -150
rect 6726 -202 6728 -150
rect 6672 -204 6728 -202
rect 7844 1505 7900 1507
rect 7844 1453 7846 1505
rect 7846 1453 7898 1505
rect 7898 1453 7900 1505
rect 7844 1451 7900 1453
rect 8932 7193 8988 7195
rect 8932 7141 8934 7193
rect 8934 7141 8986 7193
rect 8986 7141 8988 7193
rect 8932 7139 8988 7141
rect 8964 5909 9020 5965
rect 9096 5963 9152 5965
rect 9096 5911 9098 5963
rect 9098 5911 9150 5963
rect 9150 5911 9152 5963
rect 9096 5909 9152 5911
rect 8452 3978 8508 3980
rect 8452 3926 8454 3978
rect 8454 3926 8506 3978
rect 8506 3926 8508 3978
rect 8452 3924 8508 3926
rect 9128 3978 9184 3980
rect 9128 3926 9130 3978
rect 9130 3926 9182 3978
rect 9182 3926 9184 3978
rect 9128 3924 9184 3926
rect 7359 -150 7415 -148
rect 7359 -202 7361 -150
rect 7361 -202 7413 -150
rect 7413 -202 7415 -150
rect 7359 -204 7415 -202
rect 7844 -1341 7900 -1339
rect 7844 -1393 7846 -1341
rect 7846 -1393 7898 -1341
rect 7898 -1393 7900 -1341
rect 7844 -1395 7900 -1393
rect 7152 -5798 7208 -5796
rect 7152 -5850 7154 -5798
rect 7154 -5850 7206 -5798
rect 7206 -5850 7208 -5798
rect 7152 -5852 7208 -5850
rect 7844 -5823 7900 -5821
rect 7844 -5875 7846 -5823
rect 7846 -5875 7898 -5823
rect 7898 -5875 7900 -5823
rect 7844 -5877 7900 -5875
rect 3048 -7082 3104 -7026
rect 7364 -7028 7420 -7026
rect 7364 -7080 7366 -7028
rect 7366 -7080 7418 -7028
rect 7418 -7080 7420 -7028
rect 7364 -7082 7420 -7080
rect 9128 1505 9184 1507
rect 9128 1453 9130 1505
rect 9130 1453 9182 1505
rect 9182 1453 9184 1505
rect 9128 1451 9184 1453
rect 9128 -1341 9184 -1339
rect 9128 -1393 9130 -1341
rect 9130 -1393 9182 -1341
rect 9182 -1393 9184 -1341
rect 9128 -1395 9184 -1393
rect 9128 -5823 9184 -5821
rect 9128 -5875 9130 -5823
rect 9130 -5875 9182 -5823
rect 9182 -5875 9184 -5823
rect 9128 -5877 9184 -5875
<< metal3 >>
rect 554 7195 630 7205
rect 8922 7195 8998 7205
rect 554 7139 564 7195
rect 620 7139 8932 7195
rect 8988 7139 8998 7195
rect 554 7129 630 7139
rect 8922 7129 8998 7139
rect 1886 5964 1962 5974
rect 3698 5964 3774 5974
rect 5510 5964 5586 5974
rect 7322 5965 7398 5975
rect 8954 5965 9030 5975
rect 9086 5965 9162 5975
rect 7322 5964 7332 5965
rect 1886 5908 1896 5964
rect 1952 5908 3708 5964
rect 3764 5908 5520 5964
rect 5576 5909 7332 5964
rect 7388 5909 8964 5965
rect 9020 5909 9096 5965
rect 9152 5909 9162 5965
rect 5576 5908 7398 5909
rect 1886 5898 1962 5908
rect 3698 5898 3774 5908
rect 5510 5898 5586 5908
rect 7322 5899 7398 5908
rect 8954 5899 9030 5909
rect 9086 5899 9162 5909
rect 8442 3980 8518 3990
rect 9118 3980 9194 3990
rect 8442 3924 8452 3980
rect 8508 3924 9128 3980
rect 9184 3924 9194 3980
rect 8442 3914 8518 3924
rect 9118 3914 9194 3924
rect 4818 3888 4894 3898
rect 5835 3888 5911 3898
rect 4818 3832 4828 3888
rect 4884 3832 5845 3888
rect 5901 3832 5911 3888
rect 4818 3822 4894 3832
rect 5835 3822 5911 3832
rect 6022 3516 6098 3526
rect 7349 3516 7425 3526
rect 6022 3460 6032 3516
rect 6088 3460 7359 3516
rect 7415 3460 7425 3516
rect 6022 3450 6098 3460
rect 7349 3450 7425 3460
rect -2779 2893 -2667 2921
rect -2779 2837 -2751 2893
rect -2695 2837 -2667 2893
rect -2779 1183 -2667 2837
rect -2779 1127 -2750 1183
rect -2694 1127 -2667 1183
rect -2779 -527 -2667 1127
rect -2779 -583 -2750 -527
rect -2694 -583 -2667 -527
rect -2779 -611 -2667 -583
rect -2215 2893 -2103 2921
rect -2215 2837 -2187 2893
rect -2131 2837 -2103 2893
rect -2215 1183 -2103 2837
rect -2215 1127 -2186 1183
rect -2130 1127 -2103 1183
rect -2215 -527 -2103 1127
rect -2215 -583 -2186 -527
rect -2130 -583 -2103 -527
rect -2215 -2849 -2103 -583
rect -2215 -2905 -2187 -2849
rect -2131 -2905 -2103 -2849
rect -2215 -2953 -2103 -2905
rect -2215 -3009 -2187 -2953
rect -2131 -3009 -2103 -2953
rect -2215 -3037 -2103 -3009
rect -1712 2893 -1600 2921
rect -1712 2837 -1684 2893
rect -1628 2837 -1600 2893
rect -1712 1183 -1600 2837
rect 74 1532 150 1542
rect 7142 1532 7218 1542
rect 74 1476 84 1532
rect 140 1476 7152 1532
rect 7208 1476 7218 1532
rect 74 1466 150 1476
rect 7142 1466 7218 1476
rect 7834 1507 7910 1517
rect 9118 1507 9194 1517
rect 7834 1451 7844 1507
rect 7900 1451 9128 1507
rect 9184 1451 9194 1507
rect 7834 1441 7910 1451
rect 9118 1441 9194 1451
rect -1712 1127 -1683 1183
rect -1627 1127 -1600 1183
rect -1712 -527 -1600 1127
rect 6662 -148 6738 -138
rect 7349 -148 7425 -138
rect 6662 -204 6672 -148
rect 6728 -204 7359 -148
rect 7415 -204 7425 -148
rect 6662 -214 6738 -204
rect 7349 -214 7425 -204
rect -1712 -583 -1683 -527
rect -1627 -583 -1600 -527
rect -1712 -2849 -1600 -583
rect 7834 -1339 7910 -1329
rect 9118 -1339 9194 -1329
rect -181 -1364 -105 -1354
rect 3518 -1364 3594 -1354
rect -181 -1420 -171 -1364
rect -115 -1420 3528 -1364
rect 3584 -1420 3594 -1364
rect 7834 -1395 7844 -1339
rect 7900 -1395 9128 -1339
rect 9184 -1395 9194 -1339
rect 7834 -1405 7910 -1395
rect 9118 -1405 9194 -1395
rect -181 -1430 -105 -1420
rect 3518 -1430 3594 -1420
rect -1712 -2905 -1684 -2849
rect -1628 -2905 -1600 -2849
rect -1712 -2953 -1600 -2905
rect -1712 -3009 -1684 -2953
rect -1628 -3009 -1600 -2953
rect -1712 -3037 -1600 -3009
rect -425 -3255 -349 -3245
rect 3518 -3255 3594 -3245
rect -425 -3311 -415 -3255
rect -359 -3311 3528 -3255
rect 3584 -3311 3594 -3255
rect -425 -3321 -349 -3311
rect 3518 -3321 3594 -3311
rect -4285 -3797 -4209 -3787
rect -2523 -3797 -2447 -3787
rect -4285 -3853 -4275 -3797
rect -4219 -3853 -2513 -3797
rect -2457 -3853 -2447 -3797
rect -4285 -3863 -4209 -3853
rect -2523 -3863 -2447 -3853
rect -1159 -3812 -1083 -3802
rect 4013 -3812 4089 -3802
rect -1159 -3868 -1149 -3812
rect -1093 -3868 4023 -3812
rect 4079 -3868 4089 -3812
rect -1159 -3878 -1083 -3868
rect 4013 -3878 4089 -3868
rect -4123 -5796 -4047 -5786
rect -547 -5796 -471 -5786
rect -4123 -5852 -4113 -5796
rect -4057 -5852 -537 -5796
rect -481 -5852 -471 -5796
rect -4123 -5862 -4047 -5852
rect -547 -5862 -471 -5852
rect 74 -5796 150 -5786
rect 7142 -5796 7218 -5786
rect 74 -5852 84 -5796
rect 140 -5852 7152 -5796
rect 7208 -5852 7218 -5796
rect 74 -5862 150 -5852
rect 7142 -5862 7218 -5852
rect 7834 -5821 7910 -5811
rect 9118 -5821 9194 -5811
rect 7834 -5877 7844 -5821
rect 7900 -5877 9128 -5821
rect 9184 -5877 9194 -5821
rect 7834 -5887 7910 -5877
rect 9118 -5887 9194 -5877
rect -3003 -7012 -2927 -7002
rect 389 -7012 465 -7002
rect -3003 -7068 -2993 -7012
rect -2937 -7068 399 -7012
rect 455 -7068 465 -7012
rect -3003 -7078 -2927 -7068
rect 389 -7078 465 -7068
rect 3038 -7026 3114 -7016
rect 7354 -7026 7430 -7016
rect 3038 -7082 3048 -7026
rect 3104 -7082 7364 -7026
rect 7420 -7082 7430 -7026
rect 3038 -7092 3114 -7082
rect 7354 -7092 7430 -7082
<< labels >>
flabel metal1 9297 7848 9297 7848 0 FreeSans 320 0 0 0 IN2
port 4 nsew
flabel metal1 9320 7742 9320 7742 0 FreeSans 320 0 0 0 IN1
port 5 nsew
flabel metal1 9217 5937 9217 5937 0 FreeSans 320 0 0 0 EN
port 14 nsew
flabel metal1 -5082 3176 -5082 3176 0 FreeSans 320 0 0 0 A1
port 15 nsew
flabel metal1 -5088 841 -5088 841 0 FreeSans 320 0 0 0 B1
port 16 nsew
flabel metal1 -5079 -243 -5079 -243 0 FreeSans 320 0 0 0 C1
port 18 nsew
flabel metal1 3634 7382 3634 7382 0 FreeSans 320 0 0 0 VSS
port 19 nsew
flabel metal1 1831 -3615 1831 -3615 0 FreeSans 320 0 0 0 VDD
port 20 nsew
flabel metal1 9233 3946 9233 3946 0 FreeSans 320 0 0 0 IN4
port 21 nsew
flabel metal1 9226 -5845 9226 -5845 0 FreeSans 320 0 0 0 IN3
port 22 nsew
flabel metal1 -4346 -3826 -4346 -3826 0 FreeSans 320 0 0 0 OUT
port 33 nsew
flabel metal1 9281 7634 9281 7634 0 FreeSans 320 0 0 0 IN7
port 34 nsew
flabel metal1 9301 7522 9301 7522 0 FreeSans 320 0 0 0 IN5
port 35 nsew
flabel metal1 9237 1477 9237 1477 0 FreeSans 320 0 0 0 IN8
port 36 nsew
flabel metal1 9240 -1365 9240 -1365 0 FreeSans 320 0 0 0 IN6
port 37 nsew
flabel metal1 -1462 -7272 -1462 -7272 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_12.VSS
flabel nsubdiffcont -1363 -3608 -1363 -3608 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_12.VDD
flabel polycontact -641 -5824 -641 -5824 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_12.CLK
flabel metal1 -2151 -5848 -2151 -5848 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_12.VIN
flabel metal1 -2298 -5652 -2298 -5652 0 FreeSans 320 180 0 0 Transmission_Gate_Layout_12.VOUT
flabel metal1 -3264 -7272 -3264 -7272 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_13.VSS
flabel nsubdiffcont -3363 -3608 -3363 -3608 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_13.VDD
flabel polycontact -4085 -5824 -4085 -5824 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_13.CLK
flabel metal1 -2575 -5848 -2575 -5848 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_13.VIN
flabel metal1 -2428 -5652 -2428 -5652 0 FreeSans 320 180 0 0 Transmission_Gate_Layout_13.VOUT
flabel metal1 4557 -7272 4557 -7272 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_1.VSS
flabel nsubdiffcont 4458 -3608 4458 -3608 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_1.VDD
flabel polycontact 3736 -5824 3736 -5824 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_1.CLK
flabel metal1 5246 -5848 5246 -5848 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_1.VIN
flabel metal1 5393 -5652 5393 -5652 0 FreeSans 320 180 0 0 Transmission_Gate_Layout_1.VOUT
flabel metal1 2735 -7272 2735 -7272 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_2.VSS
flabel nsubdiffcont 2834 -3608 2834 -3608 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_2.VDD
flabel polycontact 3556 -5824 3556 -5824 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_2.CLK
flabel metal1 2046 -5848 2046 -5848 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_2.VIN
flabel metal1 1899 -5652 1899 -5652 0 FreeSans 320 180 0 0 Transmission_Gate_Layout_2.VOUT
flabel metal1 933 -7272 933 -7272 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_3.VSS
flabel nsubdiffcont 834 -3608 834 -3608 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_3.VDD
flabel polycontact 112 -5824 112 -5824 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_3.CLK
flabel metal1 1622 -5848 1622 -5848 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_3.VIN
flabel metal1 1769 -5652 1769 -5652 0 FreeSans 320 180 0 0 Transmission_Gate_Layout_3.VOUT
flabel metal1 4557 56 4557 56 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_9.VSS
flabel nsubdiffcont 4458 -3608 4458 -3608 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_9.VDD
flabel polycontact 3736 -1392 3736 -1392 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_9.CLK
flabel metal1 5246 -1368 5246 -1368 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_9.VIN
flabel metal1 5393 -1564 5393 -1564 0 FreeSans 320 180 0 0 Transmission_Gate_Layout_9.VOUT
flabel metal1 2735 56 2735 56 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_10.VSS
flabel nsubdiffcont 2834 -3608 2834 -3608 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_10.VDD
flabel polycontact 3556 -1392 3556 -1392 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_10.CLK
flabel metal1 2046 -1368 2046 -1368 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_10.VIN
flabel metal1 1899 -1564 1899 -1564 0 FreeSans 320 180 0 0 Transmission_Gate_Layout_10.VOUT
flabel metal1 933 56 933 56 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_11.VSS
flabel nsubdiffcont 834 -3608 834 -3608 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_11.VDD
flabel polycontact 112 -1392 112 -1392 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_11.CLK
flabel metal1 1622 -1368 1622 -1368 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_11.VIN
flabel metal1 1769 -1564 1769 -1564 0 FreeSans 320 180 0 0 Transmission_Gate_Layout_11.VOUT
flabel metal1 6359 -7272 6359 -7272 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_0.VSS
flabel nsubdiffcont 6458 -3608 6458 -3608 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_0.VDD
flabel polycontact 7180 -5824 7180 -5824 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_0.CLK
flabel metal1 5670 -5848 5670 -5848 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_0.VIN
flabel metal1 5523 -5652 5523 -5652 0 FreeSans 320 180 0 0 Transmission_Gate_Layout_0.VOUT
flabel metal1 6359 56 6359 56 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_8.VSS
flabel nsubdiffcont 6458 -3608 6458 -3608 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_8.VDD
flabel polycontact 7180 -1392 7180 -1392 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_8.CLK
flabel metal1 5670 -1368 5670 -1368 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_8.VIN
flabel metal1 5523 -1564 5523 -1564 0 FreeSans 320 180 0 0 Transmission_Gate_Layout_8.VOUT
flabel metal1 8171 -7272 8171 -7272 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_14.VSS
flabel nsubdiffcont 8270 -3608 8270 -3608 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_14.VDD
flabel polycontact 8992 -5824 8992 -5824 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_14.CLK
flabel metal1 7482 -5848 7482 -5848 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_14.VIN
flabel metal1 7335 -5652 7335 -5652 0 FreeSans 320 180 0 0 Transmission_Gate_Layout_14.VOUT
flabel metal1 8171 56 8171 56 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_21.VSS
flabel nsubdiffcont 8270 -3608 8270 -3608 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_21.VDD
flabel polycontact 8992 -1392 8992 -1392 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_21.CLK
flabel metal1 7482 -1368 7482 -1368 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_21.VIN
flabel metal1 7335 -1564 7335 -1564 0 FreeSans 320 180 0 0 Transmission_Gate_Layout_21.VOUT
flabel metal1 -5067 -234 -5067 -234 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.VIN
flabel metal1 -657 -995 -657 -995 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.PH2
flabel metal1 -3227 -553 -3227 -553 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.VSS
flabel metal1 -3264 301 -3264 301 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.VDD
flabel metal1 -529 -114 -529 -114 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.PH1
flabel psubdiffcont -4696 -555 -4696 -555 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_2.VSS
flabel metal1 -4696 303 -4696 303 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_2.VDD
flabel metal1 -4876 -241 -4876 -241 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_2.IN
flabel metal1 -4557 -114 -4557 -114 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_2.OUT
flabel metal1 -4055 -555 -4055 -555 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.VSS
flabel nsubdiffcont -4050 -1410 -4050 -1410 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.VDD
flabel metal1 -4369 -843 -4369 -843 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.A
flabel metal1 -3604 -813 -3604 -813 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.B
flabel metal1 -3811 -951 -3811 -951 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.OUT
flabel metal1 -4055 -555 -4055 -555 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.VSS
flabel nsubdiffcont -4050 300 -4050 300 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.VDD
flabel metal1 -4369 -267 -4369 -267 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.A
flabel metal1 -3604 -297 -3604 -297 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.B
flabel metal1 -3811 -159 -3811 -159 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT
flabel psubdiffcont -3227 -555 -3227 -555 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_1.VSS
flabel nsubdiffcont -3264 -1410 -3264 -1410 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_1.VDD
flabel metal1 -3418 -951 -3418 -951 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_1.IN
flabel metal1 -2910 -951 -2910 -951 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_1.OUT
flabel psubdiffcont -3227 -555 -3227 -555 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_5.VSS
flabel nsubdiffcont -3264 300 -3264 300 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_5.VDD
flabel metal1 -3418 -159 -3418 -159 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_5.IN
flabel metal1 -2910 -159 -2910 -159 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_5.OUT
flabel psubdiffcont -2441 -555 -2441 -555 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_2.VSS
flabel nsubdiffcont -2478 -1410 -2478 -1410 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_2.VDD
flabel metal1 -2632 -951 -2632 -951 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_2.IN
flabel metal1 -2124 -951 -2124 -951 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_2.OUT
flabel psubdiffcont -2441 -555 -2441 -555 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_4.VSS
flabel nsubdiffcont -2478 300 -2478 300 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_4.VDD
flabel metal1 -2632 -159 -2632 -159 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_4.IN
flabel metal1 -2124 -159 -2124 -159 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_4.OUT
flabel psubdiffcont -1655 -555 -1655 -555 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_0.VSS
flabel nsubdiffcont -1692 -1410 -1692 -1410 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_0.VDD
flabel metal1 -1846 -951 -1846 -951 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_0.IN
flabel metal1 -1338 -951 -1338 -951 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_0.OUT
flabel psubdiffcont -1655 -555 -1655 -555 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_3.VSS
flabel nsubdiffcont -1692 300 -1692 300 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_3.VDD
flabel metal1 -1846 -159 -1846 -159 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_3.IN
flabel metal1 -1338 -159 -1338 -159 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_3.OUT
flabel psubdiffcont -1047 -555 -1047 -555 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_0.VSS
flabel metal1 -1047 -1413 -1047 -1413 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_0.VDD
flabel metal1 -1227 -869 -1227 -869 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_0.IN
flabel metal1 -908 -996 -908 -996 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_0.OUT
flabel psubdiffcont -1047 -555 -1047 -555 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_1.VSS
flabel metal1 -1047 303 -1047 303 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_1.VDD
flabel metal1 -1227 -241 -1227 -241 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_1.IN
flabel metal1 -908 -114 -908 -114 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_1.OUT
flabel metal1 -5067 834 -5067 834 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.VIN
flabel metal1 -657 1595 -657 1595 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.PH2
flabel metal1 -3227 1153 -3227 1153 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.VSS
flabel metal1 -3264 299 -3264 299 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.VDD
flabel metal1 -529 714 -529 714 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.PH1
flabel psubdiffcont -4696 1155 -4696 1155 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_2.VSS
flabel metal1 -4696 297 -4696 297 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_2.VDD
flabel metal1 -4876 841 -4876 841 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_2.IN
flabel metal1 -4557 714 -4557 714 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_2.OUT
flabel metal1 -4055 1155 -4055 1155 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.VSS
flabel nsubdiffcont -4050 2010 -4050 2010 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.VDD
flabel metal1 -4369 1443 -4369 1443 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.A
flabel metal1 -3604 1413 -3604 1413 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.B
flabel metal1 -3811 1551 -3811 1551 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.OUT
flabel metal1 -4055 1155 -4055 1155 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.VSS
flabel nsubdiffcont -4050 300 -4050 300 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.VDD
flabel metal1 -4369 867 -4369 867 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.A
flabel metal1 -3604 897 -3604 897 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.B
flabel metal1 -3811 759 -3811 759 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT
flabel psubdiffcont -3227 1155 -3227 1155 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_1.VSS
flabel nsubdiffcont -3264 2010 -3264 2010 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_1.VDD
flabel metal1 -3418 1551 -3418 1551 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_1.IN
flabel metal1 -2910 1551 -2910 1551 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_1.OUT
flabel psubdiffcont -3227 1155 -3227 1155 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_5.VSS
flabel nsubdiffcont -3264 300 -3264 300 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_5.VDD
flabel metal1 -3418 759 -3418 759 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_5.IN
flabel metal1 -2910 759 -2910 759 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_5.OUT
flabel psubdiffcont -2441 1155 -2441 1155 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_2.VSS
flabel nsubdiffcont -2478 2010 -2478 2010 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_2.VDD
flabel metal1 -2632 1551 -2632 1551 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_2.IN
flabel metal1 -2124 1551 -2124 1551 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_2.OUT
flabel psubdiffcont -2441 1155 -2441 1155 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_4.VSS
flabel nsubdiffcont -2478 300 -2478 300 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_4.VDD
flabel metal1 -2632 759 -2632 759 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_4.IN
flabel metal1 -2124 759 -2124 759 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_4.OUT
flabel psubdiffcont -1655 1155 -1655 1155 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_0.VSS
flabel nsubdiffcont -1692 2010 -1692 2010 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_0.VDD
flabel metal1 -1846 1551 -1846 1551 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_0.IN
flabel metal1 -1338 1551 -1338 1551 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_0.OUT
flabel psubdiffcont -1655 1155 -1655 1155 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_3.VSS
flabel nsubdiffcont -1692 300 -1692 300 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_3.VDD
flabel metal1 -1846 759 -1846 759 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_3.IN
flabel metal1 -1338 759 -1338 759 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_3.OUT
flabel psubdiffcont -1047 1155 -1047 1155 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_0.VSS
flabel metal1 -1047 2013 -1047 2013 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_0.VDD
flabel metal1 -1227 1469 -1227 1469 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_0.IN
flabel metal1 -908 1596 -908 1596 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_0.OUT
flabel psubdiffcont -1047 1155 -1047 1155 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_1.VSS
flabel metal1 -1047 297 -1047 297 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_1.VDD
flabel metal1 -1227 841 -1227 841 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_1.IN
flabel metal1 -908 714 -908 714 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_1.OUT
flabel metal1 4557 56 4557 56 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_4.VSS
flabel nsubdiffcont 4458 3720 4458 3720 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_4.VDD
flabel polycontact 3736 1504 3736 1504 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_4.CLK
flabel metal1 5246 1480 5246 1480 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_4.VIN
flabel metal1 5393 1676 5393 1676 0 FreeSans 320 180 0 0 Transmission_Gate_Layout_4.VOUT
flabel metal1 2735 56 2735 56 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_6.VSS
flabel nsubdiffcont 2834 3720 2834 3720 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_6.VDD
flabel polycontact 3556 1504 3556 1504 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_6.CLK
flabel metal1 2046 1480 2046 1480 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_6.VIN
flabel metal1 1899 1676 1899 1676 0 FreeSans 320 180 0 0 Transmission_Gate_Layout_6.VOUT
flabel metal1 933 56 933 56 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_7.VSS
flabel nsubdiffcont 834 3720 834 3720 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_7.VDD
flabel polycontact 112 1504 112 1504 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_7.CLK
flabel metal1 1622 1480 1622 1480 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_7.VIN
flabel metal1 1769 1676 1769 1676 0 FreeSans 320 180 0 0 Transmission_Gate_Layout_7.VOUT
flabel metal1 6359 56 6359 56 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_5.VSS
flabel nsubdiffcont 6458 3720 6458 3720 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_5.VDD
flabel polycontact 7180 1504 7180 1504 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_5.CLK
flabel metal1 5670 1480 5670 1480 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_5.VIN
flabel metal1 5523 1676 5523 1676 0 FreeSans 320 180 0 0 Transmission_Gate_Layout_5.VOUT
flabel metal1 8171 56 8171 56 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_20.VSS
flabel nsubdiffcont 8270 3720 8270 3720 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_20.VDD
flabel polycontact 8992 1504 8992 1504 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_20.CLK
flabel metal1 7482 1480 7482 1480 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_20.VIN
flabel metal1 7335 1676 7335 1676 0 FreeSans 320 180 0 0 Transmission_Gate_Layout_20.VOUT
flabel metal1 -5067 3186 -5067 3186 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.VIN
flabel metal1 -657 2425 -657 2425 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.PH2
flabel metal1 -3227 2867 -3227 2867 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.VSS
flabel metal1 -3264 3721 -3264 3721 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.VDD
flabel metal1 -529 3306 -529 3306 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.PH1
flabel psubdiffcont -4696 2865 -4696 2865 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_2.VSS
flabel metal1 -4696 3723 -4696 3723 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_2.VDD
flabel metal1 -4876 3179 -4876 3179 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_2.IN
flabel metal1 -4557 3306 -4557 3306 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_2.OUT
flabel metal1 -4055 2865 -4055 2865 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.VSS
flabel nsubdiffcont -4050 2010 -4050 2010 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.VDD
flabel metal1 -4369 2577 -4369 2577 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.A
flabel metal1 -3604 2607 -3604 2607 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.B
flabel metal1 -3811 2469 -3811 2469 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.OUT
flabel metal1 -4055 2865 -4055 2865 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.VSS
flabel nsubdiffcont -4050 3720 -4050 3720 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.VDD
flabel metal1 -4369 3153 -4369 3153 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.A
flabel metal1 -3604 3123 -3604 3123 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.B
flabel metal1 -3811 3261 -3811 3261 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.OUT
flabel psubdiffcont -3227 2865 -3227 2865 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_1.VSS
flabel nsubdiffcont -3264 2010 -3264 2010 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_1.VDD
flabel metal1 -3418 2469 -3418 2469 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_1.IN
flabel metal1 -2910 2469 -2910 2469 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_1.OUT
flabel psubdiffcont -3227 2865 -3227 2865 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_5.VSS
flabel nsubdiffcont -3264 3720 -3264 3720 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_5.VDD
flabel metal1 -3418 3261 -3418 3261 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_5.IN
flabel metal1 -2910 3261 -2910 3261 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_5.OUT
flabel psubdiffcont -2441 2865 -2441 2865 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_2.VSS
flabel nsubdiffcont -2478 2010 -2478 2010 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_2.VDD
flabel metal1 -2632 2469 -2632 2469 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_2.IN
flabel metal1 -2124 2469 -2124 2469 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_2.OUT
flabel psubdiffcont -2441 2865 -2441 2865 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_4.VSS
flabel nsubdiffcont -2478 3720 -2478 3720 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_4.VDD
flabel metal1 -2632 3261 -2632 3261 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_4.IN
flabel metal1 -2124 3261 -2124 3261 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_4.OUT
flabel psubdiffcont -1655 2865 -1655 2865 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_0.VSS
flabel nsubdiffcont -1692 2010 -1692 2010 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_0.VDD
flabel metal1 -1846 2469 -1846 2469 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_0.IN
flabel metal1 -1338 2469 -1338 2469 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_0.OUT
flabel psubdiffcont -1655 2865 -1655 2865 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_3.VSS
flabel nsubdiffcont -1692 3720 -1692 3720 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_3.VDD
flabel metal1 -1846 3261 -1846 3261 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_3.IN
flabel metal1 -1338 3261 -1338 3261 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_3.OUT
flabel psubdiffcont -1047 2865 -1047 2865 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_0.VSS
flabel metal1 -1047 2007 -1047 2007 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_0.VDD
flabel metal1 -1227 2551 -1227 2551 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_0.IN
flabel metal1 -908 2424 -908 2424 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_0.OUT
flabel psubdiffcont -1047 2865 -1047 2865 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_1.VSS
flabel metal1 -1047 3723 -1047 3723 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_1.VDD
flabel metal1 -1227 3179 -1227 3179 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_1.IN
flabel metal1 -908 3306 -908 3306 0 FreeSans 320 0 0 0 Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_1.OUT
flabel metal1 2745 7384 2745 7384 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_16.VSS
flabel nsubdiffcont 2646 3720 2646 3720 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_16.VDD
flabel polycontact 1924 5936 1924 5936 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_16.CLK
flabel metal1 3434 5960 3434 5960 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_16.VIN
flabel metal1 3581 5764 3581 5764 0 FreeSans 320 180 0 0 Transmission_Gate_Layout_16.VOUT
flabel metal1 4557 7384 4557 7384 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_17.VSS
flabel nsubdiffcont 4458 3720 4458 3720 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_17.VDD
flabel polycontact 3736 5936 3736 5936 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_17.CLK
flabel metal1 5246 5960 5246 5960 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_17.VIN
flabel metal1 5393 5764 5393 5764 0 FreeSans 320 180 0 0 Transmission_Gate_Layout_17.VOUT
flabel metal1 923 7384 923 7384 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_18.VSS
flabel nsubdiffcont 1022 3720 1022 3720 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_18.VDD
flabel polycontact 1744 5936 1744 5936 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_18.CLK
flabel metal1 234 5960 234 5960 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_18.VIN
flabel metal1 87 5764 87 5764 0 FreeSans 320 180 0 0 Transmission_Gate_Layout_18.VOUT
flabel metal1 6369 7384 6369 7384 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_15.VSS
flabel nsubdiffcont 6270 3720 6270 3720 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_15.VDD
flabel polycontact 5548 5936 5548 5936 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_15.CLK
flabel metal1 7058 5960 7058 5960 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_15.VIN
flabel metal1 7205 5764 7205 5764 0 FreeSans 320 180 0 0 Transmission_Gate_Layout_15.VOUT
flabel metal1 8181 7384 8181 7384 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_19.VSS
flabel nsubdiffcont 8082 3720 8082 3720 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_19.VDD
flabel polycontact 7360 5936 7360 5936 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_19.CLK
flabel metal1 8870 5960 8870 5960 0 FreeSans 320 0 0 0 Transmission_Gate_Layout_19.VIN
flabel metal1 9017 5764 9017 5764 0 FreeSans 320 180 0 0 Transmission_Gate_Layout_19.VOUT
<< end >>
