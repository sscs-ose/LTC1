magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -4057 -1143 4057 1143
<< metal3 >>
rect -3057 138 3057 143
rect -3057 110 -3052 138
rect -3024 110 -2990 138
rect -2962 110 -2928 138
rect -2900 110 -2866 138
rect -2838 110 -2804 138
rect -2776 110 -2742 138
rect -2714 110 -2680 138
rect -2652 110 -2618 138
rect -2590 110 -2556 138
rect -2528 110 -2494 138
rect -2466 110 -2432 138
rect -2404 110 -2370 138
rect -2342 110 -2308 138
rect -2280 110 -2246 138
rect -2218 110 -2184 138
rect -2156 110 -2122 138
rect -2094 110 -2060 138
rect -2032 110 -1998 138
rect -1970 110 -1936 138
rect -1908 110 -1874 138
rect -1846 110 -1812 138
rect -1784 110 -1750 138
rect -1722 110 -1688 138
rect -1660 110 -1626 138
rect -1598 110 -1564 138
rect -1536 110 -1502 138
rect -1474 110 -1440 138
rect -1412 110 -1378 138
rect -1350 110 -1316 138
rect -1288 110 -1254 138
rect -1226 110 -1192 138
rect -1164 110 -1130 138
rect -1102 110 -1068 138
rect -1040 110 -1006 138
rect -978 110 -944 138
rect -916 110 -882 138
rect -854 110 -820 138
rect -792 110 -758 138
rect -730 110 -696 138
rect -668 110 -634 138
rect -606 110 -572 138
rect -544 110 -510 138
rect -482 110 -448 138
rect -420 110 -386 138
rect -358 110 -324 138
rect -296 110 -262 138
rect -234 110 -200 138
rect -172 110 -138 138
rect -110 110 -76 138
rect -48 110 -14 138
rect 14 110 48 138
rect 76 110 110 138
rect 138 110 172 138
rect 200 110 234 138
rect 262 110 296 138
rect 324 110 358 138
rect 386 110 420 138
rect 448 110 482 138
rect 510 110 544 138
rect 572 110 606 138
rect 634 110 668 138
rect 696 110 730 138
rect 758 110 792 138
rect 820 110 854 138
rect 882 110 916 138
rect 944 110 978 138
rect 1006 110 1040 138
rect 1068 110 1102 138
rect 1130 110 1164 138
rect 1192 110 1226 138
rect 1254 110 1288 138
rect 1316 110 1350 138
rect 1378 110 1412 138
rect 1440 110 1474 138
rect 1502 110 1536 138
rect 1564 110 1598 138
rect 1626 110 1660 138
rect 1688 110 1722 138
rect 1750 110 1784 138
rect 1812 110 1846 138
rect 1874 110 1908 138
rect 1936 110 1970 138
rect 1998 110 2032 138
rect 2060 110 2094 138
rect 2122 110 2156 138
rect 2184 110 2218 138
rect 2246 110 2280 138
rect 2308 110 2342 138
rect 2370 110 2404 138
rect 2432 110 2466 138
rect 2494 110 2528 138
rect 2556 110 2590 138
rect 2618 110 2652 138
rect 2680 110 2714 138
rect 2742 110 2776 138
rect 2804 110 2838 138
rect 2866 110 2900 138
rect 2928 110 2962 138
rect 2990 110 3024 138
rect 3052 110 3057 138
rect -3057 76 3057 110
rect -3057 48 -3052 76
rect -3024 48 -2990 76
rect -2962 48 -2928 76
rect -2900 48 -2866 76
rect -2838 48 -2804 76
rect -2776 48 -2742 76
rect -2714 48 -2680 76
rect -2652 48 -2618 76
rect -2590 48 -2556 76
rect -2528 48 -2494 76
rect -2466 48 -2432 76
rect -2404 48 -2370 76
rect -2342 48 -2308 76
rect -2280 48 -2246 76
rect -2218 48 -2184 76
rect -2156 48 -2122 76
rect -2094 48 -2060 76
rect -2032 48 -1998 76
rect -1970 48 -1936 76
rect -1908 48 -1874 76
rect -1846 48 -1812 76
rect -1784 48 -1750 76
rect -1722 48 -1688 76
rect -1660 48 -1626 76
rect -1598 48 -1564 76
rect -1536 48 -1502 76
rect -1474 48 -1440 76
rect -1412 48 -1378 76
rect -1350 48 -1316 76
rect -1288 48 -1254 76
rect -1226 48 -1192 76
rect -1164 48 -1130 76
rect -1102 48 -1068 76
rect -1040 48 -1006 76
rect -978 48 -944 76
rect -916 48 -882 76
rect -854 48 -820 76
rect -792 48 -758 76
rect -730 48 -696 76
rect -668 48 -634 76
rect -606 48 -572 76
rect -544 48 -510 76
rect -482 48 -448 76
rect -420 48 -386 76
rect -358 48 -324 76
rect -296 48 -262 76
rect -234 48 -200 76
rect -172 48 -138 76
rect -110 48 -76 76
rect -48 48 -14 76
rect 14 48 48 76
rect 76 48 110 76
rect 138 48 172 76
rect 200 48 234 76
rect 262 48 296 76
rect 324 48 358 76
rect 386 48 420 76
rect 448 48 482 76
rect 510 48 544 76
rect 572 48 606 76
rect 634 48 668 76
rect 696 48 730 76
rect 758 48 792 76
rect 820 48 854 76
rect 882 48 916 76
rect 944 48 978 76
rect 1006 48 1040 76
rect 1068 48 1102 76
rect 1130 48 1164 76
rect 1192 48 1226 76
rect 1254 48 1288 76
rect 1316 48 1350 76
rect 1378 48 1412 76
rect 1440 48 1474 76
rect 1502 48 1536 76
rect 1564 48 1598 76
rect 1626 48 1660 76
rect 1688 48 1722 76
rect 1750 48 1784 76
rect 1812 48 1846 76
rect 1874 48 1908 76
rect 1936 48 1970 76
rect 1998 48 2032 76
rect 2060 48 2094 76
rect 2122 48 2156 76
rect 2184 48 2218 76
rect 2246 48 2280 76
rect 2308 48 2342 76
rect 2370 48 2404 76
rect 2432 48 2466 76
rect 2494 48 2528 76
rect 2556 48 2590 76
rect 2618 48 2652 76
rect 2680 48 2714 76
rect 2742 48 2776 76
rect 2804 48 2838 76
rect 2866 48 2900 76
rect 2928 48 2962 76
rect 2990 48 3024 76
rect 3052 48 3057 76
rect -3057 14 3057 48
rect -3057 -14 -3052 14
rect -3024 -14 -2990 14
rect -2962 -14 -2928 14
rect -2900 -14 -2866 14
rect -2838 -14 -2804 14
rect -2776 -14 -2742 14
rect -2714 -14 -2680 14
rect -2652 -14 -2618 14
rect -2590 -14 -2556 14
rect -2528 -14 -2494 14
rect -2466 -14 -2432 14
rect -2404 -14 -2370 14
rect -2342 -14 -2308 14
rect -2280 -14 -2246 14
rect -2218 -14 -2184 14
rect -2156 -14 -2122 14
rect -2094 -14 -2060 14
rect -2032 -14 -1998 14
rect -1970 -14 -1936 14
rect -1908 -14 -1874 14
rect -1846 -14 -1812 14
rect -1784 -14 -1750 14
rect -1722 -14 -1688 14
rect -1660 -14 -1626 14
rect -1598 -14 -1564 14
rect -1536 -14 -1502 14
rect -1474 -14 -1440 14
rect -1412 -14 -1378 14
rect -1350 -14 -1316 14
rect -1288 -14 -1254 14
rect -1226 -14 -1192 14
rect -1164 -14 -1130 14
rect -1102 -14 -1068 14
rect -1040 -14 -1006 14
rect -978 -14 -944 14
rect -916 -14 -882 14
rect -854 -14 -820 14
rect -792 -14 -758 14
rect -730 -14 -696 14
rect -668 -14 -634 14
rect -606 -14 -572 14
rect -544 -14 -510 14
rect -482 -14 -448 14
rect -420 -14 -386 14
rect -358 -14 -324 14
rect -296 -14 -262 14
rect -234 -14 -200 14
rect -172 -14 -138 14
rect -110 -14 -76 14
rect -48 -14 -14 14
rect 14 -14 48 14
rect 76 -14 110 14
rect 138 -14 172 14
rect 200 -14 234 14
rect 262 -14 296 14
rect 324 -14 358 14
rect 386 -14 420 14
rect 448 -14 482 14
rect 510 -14 544 14
rect 572 -14 606 14
rect 634 -14 668 14
rect 696 -14 730 14
rect 758 -14 792 14
rect 820 -14 854 14
rect 882 -14 916 14
rect 944 -14 978 14
rect 1006 -14 1040 14
rect 1068 -14 1102 14
rect 1130 -14 1164 14
rect 1192 -14 1226 14
rect 1254 -14 1288 14
rect 1316 -14 1350 14
rect 1378 -14 1412 14
rect 1440 -14 1474 14
rect 1502 -14 1536 14
rect 1564 -14 1598 14
rect 1626 -14 1660 14
rect 1688 -14 1722 14
rect 1750 -14 1784 14
rect 1812 -14 1846 14
rect 1874 -14 1908 14
rect 1936 -14 1970 14
rect 1998 -14 2032 14
rect 2060 -14 2094 14
rect 2122 -14 2156 14
rect 2184 -14 2218 14
rect 2246 -14 2280 14
rect 2308 -14 2342 14
rect 2370 -14 2404 14
rect 2432 -14 2466 14
rect 2494 -14 2528 14
rect 2556 -14 2590 14
rect 2618 -14 2652 14
rect 2680 -14 2714 14
rect 2742 -14 2776 14
rect 2804 -14 2838 14
rect 2866 -14 2900 14
rect 2928 -14 2962 14
rect 2990 -14 3024 14
rect 3052 -14 3057 14
rect -3057 -48 3057 -14
rect -3057 -76 -3052 -48
rect -3024 -76 -2990 -48
rect -2962 -76 -2928 -48
rect -2900 -76 -2866 -48
rect -2838 -76 -2804 -48
rect -2776 -76 -2742 -48
rect -2714 -76 -2680 -48
rect -2652 -76 -2618 -48
rect -2590 -76 -2556 -48
rect -2528 -76 -2494 -48
rect -2466 -76 -2432 -48
rect -2404 -76 -2370 -48
rect -2342 -76 -2308 -48
rect -2280 -76 -2246 -48
rect -2218 -76 -2184 -48
rect -2156 -76 -2122 -48
rect -2094 -76 -2060 -48
rect -2032 -76 -1998 -48
rect -1970 -76 -1936 -48
rect -1908 -76 -1874 -48
rect -1846 -76 -1812 -48
rect -1784 -76 -1750 -48
rect -1722 -76 -1688 -48
rect -1660 -76 -1626 -48
rect -1598 -76 -1564 -48
rect -1536 -76 -1502 -48
rect -1474 -76 -1440 -48
rect -1412 -76 -1378 -48
rect -1350 -76 -1316 -48
rect -1288 -76 -1254 -48
rect -1226 -76 -1192 -48
rect -1164 -76 -1130 -48
rect -1102 -76 -1068 -48
rect -1040 -76 -1006 -48
rect -978 -76 -944 -48
rect -916 -76 -882 -48
rect -854 -76 -820 -48
rect -792 -76 -758 -48
rect -730 -76 -696 -48
rect -668 -76 -634 -48
rect -606 -76 -572 -48
rect -544 -76 -510 -48
rect -482 -76 -448 -48
rect -420 -76 -386 -48
rect -358 -76 -324 -48
rect -296 -76 -262 -48
rect -234 -76 -200 -48
rect -172 -76 -138 -48
rect -110 -76 -76 -48
rect -48 -76 -14 -48
rect 14 -76 48 -48
rect 76 -76 110 -48
rect 138 -76 172 -48
rect 200 -76 234 -48
rect 262 -76 296 -48
rect 324 -76 358 -48
rect 386 -76 420 -48
rect 448 -76 482 -48
rect 510 -76 544 -48
rect 572 -76 606 -48
rect 634 -76 668 -48
rect 696 -76 730 -48
rect 758 -76 792 -48
rect 820 -76 854 -48
rect 882 -76 916 -48
rect 944 -76 978 -48
rect 1006 -76 1040 -48
rect 1068 -76 1102 -48
rect 1130 -76 1164 -48
rect 1192 -76 1226 -48
rect 1254 -76 1288 -48
rect 1316 -76 1350 -48
rect 1378 -76 1412 -48
rect 1440 -76 1474 -48
rect 1502 -76 1536 -48
rect 1564 -76 1598 -48
rect 1626 -76 1660 -48
rect 1688 -76 1722 -48
rect 1750 -76 1784 -48
rect 1812 -76 1846 -48
rect 1874 -76 1908 -48
rect 1936 -76 1970 -48
rect 1998 -76 2032 -48
rect 2060 -76 2094 -48
rect 2122 -76 2156 -48
rect 2184 -76 2218 -48
rect 2246 -76 2280 -48
rect 2308 -76 2342 -48
rect 2370 -76 2404 -48
rect 2432 -76 2466 -48
rect 2494 -76 2528 -48
rect 2556 -76 2590 -48
rect 2618 -76 2652 -48
rect 2680 -76 2714 -48
rect 2742 -76 2776 -48
rect 2804 -76 2838 -48
rect 2866 -76 2900 -48
rect 2928 -76 2962 -48
rect 2990 -76 3024 -48
rect 3052 -76 3057 -48
rect -3057 -110 3057 -76
rect -3057 -138 -3052 -110
rect -3024 -138 -2990 -110
rect -2962 -138 -2928 -110
rect -2900 -138 -2866 -110
rect -2838 -138 -2804 -110
rect -2776 -138 -2742 -110
rect -2714 -138 -2680 -110
rect -2652 -138 -2618 -110
rect -2590 -138 -2556 -110
rect -2528 -138 -2494 -110
rect -2466 -138 -2432 -110
rect -2404 -138 -2370 -110
rect -2342 -138 -2308 -110
rect -2280 -138 -2246 -110
rect -2218 -138 -2184 -110
rect -2156 -138 -2122 -110
rect -2094 -138 -2060 -110
rect -2032 -138 -1998 -110
rect -1970 -138 -1936 -110
rect -1908 -138 -1874 -110
rect -1846 -138 -1812 -110
rect -1784 -138 -1750 -110
rect -1722 -138 -1688 -110
rect -1660 -138 -1626 -110
rect -1598 -138 -1564 -110
rect -1536 -138 -1502 -110
rect -1474 -138 -1440 -110
rect -1412 -138 -1378 -110
rect -1350 -138 -1316 -110
rect -1288 -138 -1254 -110
rect -1226 -138 -1192 -110
rect -1164 -138 -1130 -110
rect -1102 -138 -1068 -110
rect -1040 -138 -1006 -110
rect -978 -138 -944 -110
rect -916 -138 -882 -110
rect -854 -138 -820 -110
rect -792 -138 -758 -110
rect -730 -138 -696 -110
rect -668 -138 -634 -110
rect -606 -138 -572 -110
rect -544 -138 -510 -110
rect -482 -138 -448 -110
rect -420 -138 -386 -110
rect -358 -138 -324 -110
rect -296 -138 -262 -110
rect -234 -138 -200 -110
rect -172 -138 -138 -110
rect -110 -138 -76 -110
rect -48 -138 -14 -110
rect 14 -138 48 -110
rect 76 -138 110 -110
rect 138 -138 172 -110
rect 200 -138 234 -110
rect 262 -138 296 -110
rect 324 -138 358 -110
rect 386 -138 420 -110
rect 448 -138 482 -110
rect 510 -138 544 -110
rect 572 -138 606 -110
rect 634 -138 668 -110
rect 696 -138 730 -110
rect 758 -138 792 -110
rect 820 -138 854 -110
rect 882 -138 916 -110
rect 944 -138 978 -110
rect 1006 -138 1040 -110
rect 1068 -138 1102 -110
rect 1130 -138 1164 -110
rect 1192 -138 1226 -110
rect 1254 -138 1288 -110
rect 1316 -138 1350 -110
rect 1378 -138 1412 -110
rect 1440 -138 1474 -110
rect 1502 -138 1536 -110
rect 1564 -138 1598 -110
rect 1626 -138 1660 -110
rect 1688 -138 1722 -110
rect 1750 -138 1784 -110
rect 1812 -138 1846 -110
rect 1874 -138 1908 -110
rect 1936 -138 1970 -110
rect 1998 -138 2032 -110
rect 2060 -138 2094 -110
rect 2122 -138 2156 -110
rect 2184 -138 2218 -110
rect 2246 -138 2280 -110
rect 2308 -138 2342 -110
rect 2370 -138 2404 -110
rect 2432 -138 2466 -110
rect 2494 -138 2528 -110
rect 2556 -138 2590 -110
rect 2618 -138 2652 -110
rect 2680 -138 2714 -110
rect 2742 -138 2776 -110
rect 2804 -138 2838 -110
rect 2866 -138 2900 -110
rect 2928 -138 2962 -110
rect 2990 -138 3024 -110
rect 3052 -138 3057 -110
rect -3057 -143 3057 -138
<< via3 >>
rect -3052 110 -3024 138
rect -2990 110 -2962 138
rect -2928 110 -2900 138
rect -2866 110 -2838 138
rect -2804 110 -2776 138
rect -2742 110 -2714 138
rect -2680 110 -2652 138
rect -2618 110 -2590 138
rect -2556 110 -2528 138
rect -2494 110 -2466 138
rect -2432 110 -2404 138
rect -2370 110 -2342 138
rect -2308 110 -2280 138
rect -2246 110 -2218 138
rect -2184 110 -2156 138
rect -2122 110 -2094 138
rect -2060 110 -2032 138
rect -1998 110 -1970 138
rect -1936 110 -1908 138
rect -1874 110 -1846 138
rect -1812 110 -1784 138
rect -1750 110 -1722 138
rect -1688 110 -1660 138
rect -1626 110 -1598 138
rect -1564 110 -1536 138
rect -1502 110 -1474 138
rect -1440 110 -1412 138
rect -1378 110 -1350 138
rect -1316 110 -1288 138
rect -1254 110 -1226 138
rect -1192 110 -1164 138
rect -1130 110 -1102 138
rect -1068 110 -1040 138
rect -1006 110 -978 138
rect -944 110 -916 138
rect -882 110 -854 138
rect -820 110 -792 138
rect -758 110 -730 138
rect -696 110 -668 138
rect -634 110 -606 138
rect -572 110 -544 138
rect -510 110 -482 138
rect -448 110 -420 138
rect -386 110 -358 138
rect -324 110 -296 138
rect -262 110 -234 138
rect -200 110 -172 138
rect -138 110 -110 138
rect -76 110 -48 138
rect -14 110 14 138
rect 48 110 76 138
rect 110 110 138 138
rect 172 110 200 138
rect 234 110 262 138
rect 296 110 324 138
rect 358 110 386 138
rect 420 110 448 138
rect 482 110 510 138
rect 544 110 572 138
rect 606 110 634 138
rect 668 110 696 138
rect 730 110 758 138
rect 792 110 820 138
rect 854 110 882 138
rect 916 110 944 138
rect 978 110 1006 138
rect 1040 110 1068 138
rect 1102 110 1130 138
rect 1164 110 1192 138
rect 1226 110 1254 138
rect 1288 110 1316 138
rect 1350 110 1378 138
rect 1412 110 1440 138
rect 1474 110 1502 138
rect 1536 110 1564 138
rect 1598 110 1626 138
rect 1660 110 1688 138
rect 1722 110 1750 138
rect 1784 110 1812 138
rect 1846 110 1874 138
rect 1908 110 1936 138
rect 1970 110 1998 138
rect 2032 110 2060 138
rect 2094 110 2122 138
rect 2156 110 2184 138
rect 2218 110 2246 138
rect 2280 110 2308 138
rect 2342 110 2370 138
rect 2404 110 2432 138
rect 2466 110 2494 138
rect 2528 110 2556 138
rect 2590 110 2618 138
rect 2652 110 2680 138
rect 2714 110 2742 138
rect 2776 110 2804 138
rect 2838 110 2866 138
rect 2900 110 2928 138
rect 2962 110 2990 138
rect 3024 110 3052 138
rect -3052 48 -3024 76
rect -2990 48 -2962 76
rect -2928 48 -2900 76
rect -2866 48 -2838 76
rect -2804 48 -2776 76
rect -2742 48 -2714 76
rect -2680 48 -2652 76
rect -2618 48 -2590 76
rect -2556 48 -2528 76
rect -2494 48 -2466 76
rect -2432 48 -2404 76
rect -2370 48 -2342 76
rect -2308 48 -2280 76
rect -2246 48 -2218 76
rect -2184 48 -2156 76
rect -2122 48 -2094 76
rect -2060 48 -2032 76
rect -1998 48 -1970 76
rect -1936 48 -1908 76
rect -1874 48 -1846 76
rect -1812 48 -1784 76
rect -1750 48 -1722 76
rect -1688 48 -1660 76
rect -1626 48 -1598 76
rect -1564 48 -1536 76
rect -1502 48 -1474 76
rect -1440 48 -1412 76
rect -1378 48 -1350 76
rect -1316 48 -1288 76
rect -1254 48 -1226 76
rect -1192 48 -1164 76
rect -1130 48 -1102 76
rect -1068 48 -1040 76
rect -1006 48 -978 76
rect -944 48 -916 76
rect -882 48 -854 76
rect -820 48 -792 76
rect -758 48 -730 76
rect -696 48 -668 76
rect -634 48 -606 76
rect -572 48 -544 76
rect -510 48 -482 76
rect -448 48 -420 76
rect -386 48 -358 76
rect -324 48 -296 76
rect -262 48 -234 76
rect -200 48 -172 76
rect -138 48 -110 76
rect -76 48 -48 76
rect -14 48 14 76
rect 48 48 76 76
rect 110 48 138 76
rect 172 48 200 76
rect 234 48 262 76
rect 296 48 324 76
rect 358 48 386 76
rect 420 48 448 76
rect 482 48 510 76
rect 544 48 572 76
rect 606 48 634 76
rect 668 48 696 76
rect 730 48 758 76
rect 792 48 820 76
rect 854 48 882 76
rect 916 48 944 76
rect 978 48 1006 76
rect 1040 48 1068 76
rect 1102 48 1130 76
rect 1164 48 1192 76
rect 1226 48 1254 76
rect 1288 48 1316 76
rect 1350 48 1378 76
rect 1412 48 1440 76
rect 1474 48 1502 76
rect 1536 48 1564 76
rect 1598 48 1626 76
rect 1660 48 1688 76
rect 1722 48 1750 76
rect 1784 48 1812 76
rect 1846 48 1874 76
rect 1908 48 1936 76
rect 1970 48 1998 76
rect 2032 48 2060 76
rect 2094 48 2122 76
rect 2156 48 2184 76
rect 2218 48 2246 76
rect 2280 48 2308 76
rect 2342 48 2370 76
rect 2404 48 2432 76
rect 2466 48 2494 76
rect 2528 48 2556 76
rect 2590 48 2618 76
rect 2652 48 2680 76
rect 2714 48 2742 76
rect 2776 48 2804 76
rect 2838 48 2866 76
rect 2900 48 2928 76
rect 2962 48 2990 76
rect 3024 48 3052 76
rect -3052 -14 -3024 14
rect -2990 -14 -2962 14
rect -2928 -14 -2900 14
rect -2866 -14 -2838 14
rect -2804 -14 -2776 14
rect -2742 -14 -2714 14
rect -2680 -14 -2652 14
rect -2618 -14 -2590 14
rect -2556 -14 -2528 14
rect -2494 -14 -2466 14
rect -2432 -14 -2404 14
rect -2370 -14 -2342 14
rect -2308 -14 -2280 14
rect -2246 -14 -2218 14
rect -2184 -14 -2156 14
rect -2122 -14 -2094 14
rect -2060 -14 -2032 14
rect -1998 -14 -1970 14
rect -1936 -14 -1908 14
rect -1874 -14 -1846 14
rect -1812 -14 -1784 14
rect -1750 -14 -1722 14
rect -1688 -14 -1660 14
rect -1626 -14 -1598 14
rect -1564 -14 -1536 14
rect -1502 -14 -1474 14
rect -1440 -14 -1412 14
rect -1378 -14 -1350 14
rect -1316 -14 -1288 14
rect -1254 -14 -1226 14
rect -1192 -14 -1164 14
rect -1130 -14 -1102 14
rect -1068 -14 -1040 14
rect -1006 -14 -978 14
rect -944 -14 -916 14
rect -882 -14 -854 14
rect -820 -14 -792 14
rect -758 -14 -730 14
rect -696 -14 -668 14
rect -634 -14 -606 14
rect -572 -14 -544 14
rect -510 -14 -482 14
rect -448 -14 -420 14
rect -386 -14 -358 14
rect -324 -14 -296 14
rect -262 -14 -234 14
rect -200 -14 -172 14
rect -138 -14 -110 14
rect -76 -14 -48 14
rect -14 -14 14 14
rect 48 -14 76 14
rect 110 -14 138 14
rect 172 -14 200 14
rect 234 -14 262 14
rect 296 -14 324 14
rect 358 -14 386 14
rect 420 -14 448 14
rect 482 -14 510 14
rect 544 -14 572 14
rect 606 -14 634 14
rect 668 -14 696 14
rect 730 -14 758 14
rect 792 -14 820 14
rect 854 -14 882 14
rect 916 -14 944 14
rect 978 -14 1006 14
rect 1040 -14 1068 14
rect 1102 -14 1130 14
rect 1164 -14 1192 14
rect 1226 -14 1254 14
rect 1288 -14 1316 14
rect 1350 -14 1378 14
rect 1412 -14 1440 14
rect 1474 -14 1502 14
rect 1536 -14 1564 14
rect 1598 -14 1626 14
rect 1660 -14 1688 14
rect 1722 -14 1750 14
rect 1784 -14 1812 14
rect 1846 -14 1874 14
rect 1908 -14 1936 14
rect 1970 -14 1998 14
rect 2032 -14 2060 14
rect 2094 -14 2122 14
rect 2156 -14 2184 14
rect 2218 -14 2246 14
rect 2280 -14 2308 14
rect 2342 -14 2370 14
rect 2404 -14 2432 14
rect 2466 -14 2494 14
rect 2528 -14 2556 14
rect 2590 -14 2618 14
rect 2652 -14 2680 14
rect 2714 -14 2742 14
rect 2776 -14 2804 14
rect 2838 -14 2866 14
rect 2900 -14 2928 14
rect 2962 -14 2990 14
rect 3024 -14 3052 14
rect -3052 -76 -3024 -48
rect -2990 -76 -2962 -48
rect -2928 -76 -2900 -48
rect -2866 -76 -2838 -48
rect -2804 -76 -2776 -48
rect -2742 -76 -2714 -48
rect -2680 -76 -2652 -48
rect -2618 -76 -2590 -48
rect -2556 -76 -2528 -48
rect -2494 -76 -2466 -48
rect -2432 -76 -2404 -48
rect -2370 -76 -2342 -48
rect -2308 -76 -2280 -48
rect -2246 -76 -2218 -48
rect -2184 -76 -2156 -48
rect -2122 -76 -2094 -48
rect -2060 -76 -2032 -48
rect -1998 -76 -1970 -48
rect -1936 -76 -1908 -48
rect -1874 -76 -1846 -48
rect -1812 -76 -1784 -48
rect -1750 -76 -1722 -48
rect -1688 -76 -1660 -48
rect -1626 -76 -1598 -48
rect -1564 -76 -1536 -48
rect -1502 -76 -1474 -48
rect -1440 -76 -1412 -48
rect -1378 -76 -1350 -48
rect -1316 -76 -1288 -48
rect -1254 -76 -1226 -48
rect -1192 -76 -1164 -48
rect -1130 -76 -1102 -48
rect -1068 -76 -1040 -48
rect -1006 -76 -978 -48
rect -944 -76 -916 -48
rect -882 -76 -854 -48
rect -820 -76 -792 -48
rect -758 -76 -730 -48
rect -696 -76 -668 -48
rect -634 -76 -606 -48
rect -572 -76 -544 -48
rect -510 -76 -482 -48
rect -448 -76 -420 -48
rect -386 -76 -358 -48
rect -324 -76 -296 -48
rect -262 -76 -234 -48
rect -200 -76 -172 -48
rect -138 -76 -110 -48
rect -76 -76 -48 -48
rect -14 -76 14 -48
rect 48 -76 76 -48
rect 110 -76 138 -48
rect 172 -76 200 -48
rect 234 -76 262 -48
rect 296 -76 324 -48
rect 358 -76 386 -48
rect 420 -76 448 -48
rect 482 -76 510 -48
rect 544 -76 572 -48
rect 606 -76 634 -48
rect 668 -76 696 -48
rect 730 -76 758 -48
rect 792 -76 820 -48
rect 854 -76 882 -48
rect 916 -76 944 -48
rect 978 -76 1006 -48
rect 1040 -76 1068 -48
rect 1102 -76 1130 -48
rect 1164 -76 1192 -48
rect 1226 -76 1254 -48
rect 1288 -76 1316 -48
rect 1350 -76 1378 -48
rect 1412 -76 1440 -48
rect 1474 -76 1502 -48
rect 1536 -76 1564 -48
rect 1598 -76 1626 -48
rect 1660 -76 1688 -48
rect 1722 -76 1750 -48
rect 1784 -76 1812 -48
rect 1846 -76 1874 -48
rect 1908 -76 1936 -48
rect 1970 -76 1998 -48
rect 2032 -76 2060 -48
rect 2094 -76 2122 -48
rect 2156 -76 2184 -48
rect 2218 -76 2246 -48
rect 2280 -76 2308 -48
rect 2342 -76 2370 -48
rect 2404 -76 2432 -48
rect 2466 -76 2494 -48
rect 2528 -76 2556 -48
rect 2590 -76 2618 -48
rect 2652 -76 2680 -48
rect 2714 -76 2742 -48
rect 2776 -76 2804 -48
rect 2838 -76 2866 -48
rect 2900 -76 2928 -48
rect 2962 -76 2990 -48
rect 3024 -76 3052 -48
rect -3052 -138 -3024 -110
rect -2990 -138 -2962 -110
rect -2928 -138 -2900 -110
rect -2866 -138 -2838 -110
rect -2804 -138 -2776 -110
rect -2742 -138 -2714 -110
rect -2680 -138 -2652 -110
rect -2618 -138 -2590 -110
rect -2556 -138 -2528 -110
rect -2494 -138 -2466 -110
rect -2432 -138 -2404 -110
rect -2370 -138 -2342 -110
rect -2308 -138 -2280 -110
rect -2246 -138 -2218 -110
rect -2184 -138 -2156 -110
rect -2122 -138 -2094 -110
rect -2060 -138 -2032 -110
rect -1998 -138 -1970 -110
rect -1936 -138 -1908 -110
rect -1874 -138 -1846 -110
rect -1812 -138 -1784 -110
rect -1750 -138 -1722 -110
rect -1688 -138 -1660 -110
rect -1626 -138 -1598 -110
rect -1564 -138 -1536 -110
rect -1502 -138 -1474 -110
rect -1440 -138 -1412 -110
rect -1378 -138 -1350 -110
rect -1316 -138 -1288 -110
rect -1254 -138 -1226 -110
rect -1192 -138 -1164 -110
rect -1130 -138 -1102 -110
rect -1068 -138 -1040 -110
rect -1006 -138 -978 -110
rect -944 -138 -916 -110
rect -882 -138 -854 -110
rect -820 -138 -792 -110
rect -758 -138 -730 -110
rect -696 -138 -668 -110
rect -634 -138 -606 -110
rect -572 -138 -544 -110
rect -510 -138 -482 -110
rect -448 -138 -420 -110
rect -386 -138 -358 -110
rect -324 -138 -296 -110
rect -262 -138 -234 -110
rect -200 -138 -172 -110
rect -138 -138 -110 -110
rect -76 -138 -48 -110
rect -14 -138 14 -110
rect 48 -138 76 -110
rect 110 -138 138 -110
rect 172 -138 200 -110
rect 234 -138 262 -110
rect 296 -138 324 -110
rect 358 -138 386 -110
rect 420 -138 448 -110
rect 482 -138 510 -110
rect 544 -138 572 -110
rect 606 -138 634 -110
rect 668 -138 696 -110
rect 730 -138 758 -110
rect 792 -138 820 -110
rect 854 -138 882 -110
rect 916 -138 944 -110
rect 978 -138 1006 -110
rect 1040 -138 1068 -110
rect 1102 -138 1130 -110
rect 1164 -138 1192 -110
rect 1226 -138 1254 -110
rect 1288 -138 1316 -110
rect 1350 -138 1378 -110
rect 1412 -138 1440 -110
rect 1474 -138 1502 -110
rect 1536 -138 1564 -110
rect 1598 -138 1626 -110
rect 1660 -138 1688 -110
rect 1722 -138 1750 -110
rect 1784 -138 1812 -110
rect 1846 -138 1874 -110
rect 1908 -138 1936 -110
rect 1970 -138 1998 -110
rect 2032 -138 2060 -110
rect 2094 -138 2122 -110
rect 2156 -138 2184 -110
rect 2218 -138 2246 -110
rect 2280 -138 2308 -110
rect 2342 -138 2370 -110
rect 2404 -138 2432 -110
rect 2466 -138 2494 -110
rect 2528 -138 2556 -110
rect 2590 -138 2618 -110
rect 2652 -138 2680 -110
rect 2714 -138 2742 -110
rect 2776 -138 2804 -110
rect 2838 -138 2866 -110
rect 2900 -138 2928 -110
rect 2962 -138 2990 -110
rect 3024 -138 3052 -110
<< metal4 >>
rect -3057 138 3057 143
rect -3057 110 -3052 138
rect -3024 110 -2990 138
rect -2962 110 -2928 138
rect -2900 110 -2866 138
rect -2838 110 -2804 138
rect -2776 110 -2742 138
rect -2714 110 -2680 138
rect -2652 110 -2618 138
rect -2590 110 -2556 138
rect -2528 110 -2494 138
rect -2466 110 -2432 138
rect -2404 110 -2370 138
rect -2342 110 -2308 138
rect -2280 110 -2246 138
rect -2218 110 -2184 138
rect -2156 110 -2122 138
rect -2094 110 -2060 138
rect -2032 110 -1998 138
rect -1970 110 -1936 138
rect -1908 110 -1874 138
rect -1846 110 -1812 138
rect -1784 110 -1750 138
rect -1722 110 -1688 138
rect -1660 110 -1626 138
rect -1598 110 -1564 138
rect -1536 110 -1502 138
rect -1474 110 -1440 138
rect -1412 110 -1378 138
rect -1350 110 -1316 138
rect -1288 110 -1254 138
rect -1226 110 -1192 138
rect -1164 110 -1130 138
rect -1102 110 -1068 138
rect -1040 110 -1006 138
rect -978 110 -944 138
rect -916 110 -882 138
rect -854 110 -820 138
rect -792 110 -758 138
rect -730 110 -696 138
rect -668 110 -634 138
rect -606 110 -572 138
rect -544 110 -510 138
rect -482 110 -448 138
rect -420 110 -386 138
rect -358 110 -324 138
rect -296 110 -262 138
rect -234 110 -200 138
rect -172 110 -138 138
rect -110 110 -76 138
rect -48 110 -14 138
rect 14 110 48 138
rect 76 110 110 138
rect 138 110 172 138
rect 200 110 234 138
rect 262 110 296 138
rect 324 110 358 138
rect 386 110 420 138
rect 448 110 482 138
rect 510 110 544 138
rect 572 110 606 138
rect 634 110 668 138
rect 696 110 730 138
rect 758 110 792 138
rect 820 110 854 138
rect 882 110 916 138
rect 944 110 978 138
rect 1006 110 1040 138
rect 1068 110 1102 138
rect 1130 110 1164 138
rect 1192 110 1226 138
rect 1254 110 1288 138
rect 1316 110 1350 138
rect 1378 110 1412 138
rect 1440 110 1474 138
rect 1502 110 1536 138
rect 1564 110 1598 138
rect 1626 110 1660 138
rect 1688 110 1722 138
rect 1750 110 1784 138
rect 1812 110 1846 138
rect 1874 110 1908 138
rect 1936 110 1970 138
rect 1998 110 2032 138
rect 2060 110 2094 138
rect 2122 110 2156 138
rect 2184 110 2218 138
rect 2246 110 2280 138
rect 2308 110 2342 138
rect 2370 110 2404 138
rect 2432 110 2466 138
rect 2494 110 2528 138
rect 2556 110 2590 138
rect 2618 110 2652 138
rect 2680 110 2714 138
rect 2742 110 2776 138
rect 2804 110 2838 138
rect 2866 110 2900 138
rect 2928 110 2962 138
rect 2990 110 3024 138
rect 3052 110 3057 138
rect -3057 76 3057 110
rect -3057 48 -3052 76
rect -3024 48 -2990 76
rect -2962 48 -2928 76
rect -2900 48 -2866 76
rect -2838 48 -2804 76
rect -2776 48 -2742 76
rect -2714 48 -2680 76
rect -2652 48 -2618 76
rect -2590 48 -2556 76
rect -2528 48 -2494 76
rect -2466 48 -2432 76
rect -2404 48 -2370 76
rect -2342 48 -2308 76
rect -2280 48 -2246 76
rect -2218 48 -2184 76
rect -2156 48 -2122 76
rect -2094 48 -2060 76
rect -2032 48 -1998 76
rect -1970 48 -1936 76
rect -1908 48 -1874 76
rect -1846 48 -1812 76
rect -1784 48 -1750 76
rect -1722 48 -1688 76
rect -1660 48 -1626 76
rect -1598 48 -1564 76
rect -1536 48 -1502 76
rect -1474 48 -1440 76
rect -1412 48 -1378 76
rect -1350 48 -1316 76
rect -1288 48 -1254 76
rect -1226 48 -1192 76
rect -1164 48 -1130 76
rect -1102 48 -1068 76
rect -1040 48 -1006 76
rect -978 48 -944 76
rect -916 48 -882 76
rect -854 48 -820 76
rect -792 48 -758 76
rect -730 48 -696 76
rect -668 48 -634 76
rect -606 48 -572 76
rect -544 48 -510 76
rect -482 48 -448 76
rect -420 48 -386 76
rect -358 48 -324 76
rect -296 48 -262 76
rect -234 48 -200 76
rect -172 48 -138 76
rect -110 48 -76 76
rect -48 48 -14 76
rect 14 48 48 76
rect 76 48 110 76
rect 138 48 172 76
rect 200 48 234 76
rect 262 48 296 76
rect 324 48 358 76
rect 386 48 420 76
rect 448 48 482 76
rect 510 48 544 76
rect 572 48 606 76
rect 634 48 668 76
rect 696 48 730 76
rect 758 48 792 76
rect 820 48 854 76
rect 882 48 916 76
rect 944 48 978 76
rect 1006 48 1040 76
rect 1068 48 1102 76
rect 1130 48 1164 76
rect 1192 48 1226 76
rect 1254 48 1288 76
rect 1316 48 1350 76
rect 1378 48 1412 76
rect 1440 48 1474 76
rect 1502 48 1536 76
rect 1564 48 1598 76
rect 1626 48 1660 76
rect 1688 48 1722 76
rect 1750 48 1784 76
rect 1812 48 1846 76
rect 1874 48 1908 76
rect 1936 48 1970 76
rect 1998 48 2032 76
rect 2060 48 2094 76
rect 2122 48 2156 76
rect 2184 48 2218 76
rect 2246 48 2280 76
rect 2308 48 2342 76
rect 2370 48 2404 76
rect 2432 48 2466 76
rect 2494 48 2528 76
rect 2556 48 2590 76
rect 2618 48 2652 76
rect 2680 48 2714 76
rect 2742 48 2776 76
rect 2804 48 2838 76
rect 2866 48 2900 76
rect 2928 48 2962 76
rect 2990 48 3024 76
rect 3052 48 3057 76
rect -3057 14 3057 48
rect -3057 -14 -3052 14
rect -3024 -14 -2990 14
rect -2962 -14 -2928 14
rect -2900 -14 -2866 14
rect -2838 -14 -2804 14
rect -2776 -14 -2742 14
rect -2714 -14 -2680 14
rect -2652 -14 -2618 14
rect -2590 -14 -2556 14
rect -2528 -14 -2494 14
rect -2466 -14 -2432 14
rect -2404 -14 -2370 14
rect -2342 -14 -2308 14
rect -2280 -14 -2246 14
rect -2218 -14 -2184 14
rect -2156 -14 -2122 14
rect -2094 -14 -2060 14
rect -2032 -14 -1998 14
rect -1970 -14 -1936 14
rect -1908 -14 -1874 14
rect -1846 -14 -1812 14
rect -1784 -14 -1750 14
rect -1722 -14 -1688 14
rect -1660 -14 -1626 14
rect -1598 -14 -1564 14
rect -1536 -14 -1502 14
rect -1474 -14 -1440 14
rect -1412 -14 -1378 14
rect -1350 -14 -1316 14
rect -1288 -14 -1254 14
rect -1226 -14 -1192 14
rect -1164 -14 -1130 14
rect -1102 -14 -1068 14
rect -1040 -14 -1006 14
rect -978 -14 -944 14
rect -916 -14 -882 14
rect -854 -14 -820 14
rect -792 -14 -758 14
rect -730 -14 -696 14
rect -668 -14 -634 14
rect -606 -14 -572 14
rect -544 -14 -510 14
rect -482 -14 -448 14
rect -420 -14 -386 14
rect -358 -14 -324 14
rect -296 -14 -262 14
rect -234 -14 -200 14
rect -172 -14 -138 14
rect -110 -14 -76 14
rect -48 -14 -14 14
rect 14 -14 48 14
rect 76 -14 110 14
rect 138 -14 172 14
rect 200 -14 234 14
rect 262 -14 296 14
rect 324 -14 358 14
rect 386 -14 420 14
rect 448 -14 482 14
rect 510 -14 544 14
rect 572 -14 606 14
rect 634 -14 668 14
rect 696 -14 730 14
rect 758 -14 792 14
rect 820 -14 854 14
rect 882 -14 916 14
rect 944 -14 978 14
rect 1006 -14 1040 14
rect 1068 -14 1102 14
rect 1130 -14 1164 14
rect 1192 -14 1226 14
rect 1254 -14 1288 14
rect 1316 -14 1350 14
rect 1378 -14 1412 14
rect 1440 -14 1474 14
rect 1502 -14 1536 14
rect 1564 -14 1598 14
rect 1626 -14 1660 14
rect 1688 -14 1722 14
rect 1750 -14 1784 14
rect 1812 -14 1846 14
rect 1874 -14 1908 14
rect 1936 -14 1970 14
rect 1998 -14 2032 14
rect 2060 -14 2094 14
rect 2122 -14 2156 14
rect 2184 -14 2218 14
rect 2246 -14 2280 14
rect 2308 -14 2342 14
rect 2370 -14 2404 14
rect 2432 -14 2466 14
rect 2494 -14 2528 14
rect 2556 -14 2590 14
rect 2618 -14 2652 14
rect 2680 -14 2714 14
rect 2742 -14 2776 14
rect 2804 -14 2838 14
rect 2866 -14 2900 14
rect 2928 -14 2962 14
rect 2990 -14 3024 14
rect 3052 -14 3057 14
rect -3057 -48 3057 -14
rect -3057 -76 -3052 -48
rect -3024 -76 -2990 -48
rect -2962 -76 -2928 -48
rect -2900 -76 -2866 -48
rect -2838 -76 -2804 -48
rect -2776 -76 -2742 -48
rect -2714 -76 -2680 -48
rect -2652 -76 -2618 -48
rect -2590 -76 -2556 -48
rect -2528 -76 -2494 -48
rect -2466 -76 -2432 -48
rect -2404 -76 -2370 -48
rect -2342 -76 -2308 -48
rect -2280 -76 -2246 -48
rect -2218 -76 -2184 -48
rect -2156 -76 -2122 -48
rect -2094 -76 -2060 -48
rect -2032 -76 -1998 -48
rect -1970 -76 -1936 -48
rect -1908 -76 -1874 -48
rect -1846 -76 -1812 -48
rect -1784 -76 -1750 -48
rect -1722 -76 -1688 -48
rect -1660 -76 -1626 -48
rect -1598 -76 -1564 -48
rect -1536 -76 -1502 -48
rect -1474 -76 -1440 -48
rect -1412 -76 -1378 -48
rect -1350 -76 -1316 -48
rect -1288 -76 -1254 -48
rect -1226 -76 -1192 -48
rect -1164 -76 -1130 -48
rect -1102 -76 -1068 -48
rect -1040 -76 -1006 -48
rect -978 -76 -944 -48
rect -916 -76 -882 -48
rect -854 -76 -820 -48
rect -792 -76 -758 -48
rect -730 -76 -696 -48
rect -668 -76 -634 -48
rect -606 -76 -572 -48
rect -544 -76 -510 -48
rect -482 -76 -448 -48
rect -420 -76 -386 -48
rect -358 -76 -324 -48
rect -296 -76 -262 -48
rect -234 -76 -200 -48
rect -172 -76 -138 -48
rect -110 -76 -76 -48
rect -48 -76 -14 -48
rect 14 -76 48 -48
rect 76 -76 110 -48
rect 138 -76 172 -48
rect 200 -76 234 -48
rect 262 -76 296 -48
rect 324 -76 358 -48
rect 386 -76 420 -48
rect 448 -76 482 -48
rect 510 -76 544 -48
rect 572 -76 606 -48
rect 634 -76 668 -48
rect 696 -76 730 -48
rect 758 -76 792 -48
rect 820 -76 854 -48
rect 882 -76 916 -48
rect 944 -76 978 -48
rect 1006 -76 1040 -48
rect 1068 -76 1102 -48
rect 1130 -76 1164 -48
rect 1192 -76 1226 -48
rect 1254 -76 1288 -48
rect 1316 -76 1350 -48
rect 1378 -76 1412 -48
rect 1440 -76 1474 -48
rect 1502 -76 1536 -48
rect 1564 -76 1598 -48
rect 1626 -76 1660 -48
rect 1688 -76 1722 -48
rect 1750 -76 1784 -48
rect 1812 -76 1846 -48
rect 1874 -76 1908 -48
rect 1936 -76 1970 -48
rect 1998 -76 2032 -48
rect 2060 -76 2094 -48
rect 2122 -76 2156 -48
rect 2184 -76 2218 -48
rect 2246 -76 2280 -48
rect 2308 -76 2342 -48
rect 2370 -76 2404 -48
rect 2432 -76 2466 -48
rect 2494 -76 2528 -48
rect 2556 -76 2590 -48
rect 2618 -76 2652 -48
rect 2680 -76 2714 -48
rect 2742 -76 2776 -48
rect 2804 -76 2838 -48
rect 2866 -76 2900 -48
rect 2928 -76 2962 -48
rect 2990 -76 3024 -48
rect 3052 -76 3057 -48
rect -3057 -110 3057 -76
rect -3057 -138 -3052 -110
rect -3024 -138 -2990 -110
rect -2962 -138 -2928 -110
rect -2900 -138 -2866 -110
rect -2838 -138 -2804 -110
rect -2776 -138 -2742 -110
rect -2714 -138 -2680 -110
rect -2652 -138 -2618 -110
rect -2590 -138 -2556 -110
rect -2528 -138 -2494 -110
rect -2466 -138 -2432 -110
rect -2404 -138 -2370 -110
rect -2342 -138 -2308 -110
rect -2280 -138 -2246 -110
rect -2218 -138 -2184 -110
rect -2156 -138 -2122 -110
rect -2094 -138 -2060 -110
rect -2032 -138 -1998 -110
rect -1970 -138 -1936 -110
rect -1908 -138 -1874 -110
rect -1846 -138 -1812 -110
rect -1784 -138 -1750 -110
rect -1722 -138 -1688 -110
rect -1660 -138 -1626 -110
rect -1598 -138 -1564 -110
rect -1536 -138 -1502 -110
rect -1474 -138 -1440 -110
rect -1412 -138 -1378 -110
rect -1350 -138 -1316 -110
rect -1288 -138 -1254 -110
rect -1226 -138 -1192 -110
rect -1164 -138 -1130 -110
rect -1102 -138 -1068 -110
rect -1040 -138 -1006 -110
rect -978 -138 -944 -110
rect -916 -138 -882 -110
rect -854 -138 -820 -110
rect -792 -138 -758 -110
rect -730 -138 -696 -110
rect -668 -138 -634 -110
rect -606 -138 -572 -110
rect -544 -138 -510 -110
rect -482 -138 -448 -110
rect -420 -138 -386 -110
rect -358 -138 -324 -110
rect -296 -138 -262 -110
rect -234 -138 -200 -110
rect -172 -138 -138 -110
rect -110 -138 -76 -110
rect -48 -138 -14 -110
rect 14 -138 48 -110
rect 76 -138 110 -110
rect 138 -138 172 -110
rect 200 -138 234 -110
rect 262 -138 296 -110
rect 324 -138 358 -110
rect 386 -138 420 -110
rect 448 -138 482 -110
rect 510 -138 544 -110
rect 572 -138 606 -110
rect 634 -138 668 -110
rect 696 -138 730 -110
rect 758 -138 792 -110
rect 820 -138 854 -110
rect 882 -138 916 -110
rect 944 -138 978 -110
rect 1006 -138 1040 -110
rect 1068 -138 1102 -110
rect 1130 -138 1164 -110
rect 1192 -138 1226 -110
rect 1254 -138 1288 -110
rect 1316 -138 1350 -110
rect 1378 -138 1412 -110
rect 1440 -138 1474 -110
rect 1502 -138 1536 -110
rect 1564 -138 1598 -110
rect 1626 -138 1660 -110
rect 1688 -138 1722 -110
rect 1750 -138 1784 -110
rect 1812 -138 1846 -110
rect 1874 -138 1908 -110
rect 1936 -138 1970 -110
rect 1998 -138 2032 -110
rect 2060 -138 2094 -110
rect 2122 -138 2156 -110
rect 2184 -138 2218 -110
rect 2246 -138 2280 -110
rect 2308 -138 2342 -110
rect 2370 -138 2404 -110
rect 2432 -138 2466 -110
rect 2494 -138 2528 -110
rect 2556 -138 2590 -110
rect 2618 -138 2652 -110
rect 2680 -138 2714 -110
rect 2742 -138 2776 -110
rect 2804 -138 2838 -110
rect 2866 -138 2900 -110
rect 2928 -138 2962 -110
rect 2990 -138 3024 -110
rect 3052 -138 3057 -110
rect -3057 -143 3057 -138
<< end >>
