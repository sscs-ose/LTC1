magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1046 -1019 1046 1019
<< metal1 >>
rect -46 13 46 19
rect -46 -13 -40 13
rect -14 -13 14 13
rect 40 -13 46 13
rect -46 -19 46 -13
<< via1 >>
rect -40 -13 -14 13
rect 14 -13 40 13
<< metal2 >>
rect -46 13 46 19
rect -46 -13 -40 13
rect -14 -13 14 13
rect 40 -13 46 13
rect -46 -19 46 -13
<< end >>
