* NGSPICE file created from AND_3_In_Layout_flat.ext - technology: gf180mcuC

.subckt AND_3_In_Layout_flat A B C OUT VDD VSS
X0 OUT a_24_68# VDD.t1 VDD.t0 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_24_68# A.t0 a_168_68# VSS.t11 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X2 a_648_68# B.t0 a_168_68# VSS.t12 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X3 a_168_68# A.t1 a_24_68# VSS.t10 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X4 OUT a_24_68# VSS.t1 VSS.t0 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X5 a_24_68# B.t1 VDD.t3 VDD.t2 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X6 a_168_68# B.t2 a_648_68# VSS.t4 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X7 VSS C.t0 a_648_68# VSS.t6 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X8 a_648_68# B.t3 a_168_68# VSS.t5 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X9 a_648_68# C.t1 VSS.t3 VSS.t2 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X10 VDD C.t2 a_24_68# VDD.t4 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X11 a_168_68# A.t2 a_24_68# VSS.t9 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X12 VSS C.t3 a_648_68# VSS.t13 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X13 VDD A.t3 a_24_68# VDD.t7 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
R0 VDD.n9 VDD.t4 154.44
R1 VDD.n4 VDD.t0 85.6379
R2 VDD.n15 VDD.t7 85.6365
R3 VDD.t4 VDD.n8 27.0275
R4 VDD.n17 VDD.t2 27.0275
R5 VDD.n10 VDD.n7 8.2255
R6 VDD.n18 VDD.n10 8.2255
R7 VDD VDD.n10 6.3005
R8 VDD VDD.n10 6.3005
R9 VDD.n3 VDD.n2 3.1505
R10 VDD.n7 VDD.n6 3.1505
R11 VDD.n8 VDD.n7 3.1505
R12 VDD.n10 VDD.n9 3.1505
R13 VDD.n19 VDD.n18 3.1505
R14 VDD.n18 VDD.n17 3.1505
R15 VDD.n14 VDD.n13 3.1505
R16 VDD.n5 VDD.n1 2.91941
R17 VDD.n16 VDD.n12 2.91705
R18 VDD.n4 VDD.n3 1.87098
R19 VDD.n15 VDD.n14 1.8708
R20 VDD.n12 VDD.t3 1.8205
R21 VDD.n12 VDD.n11 1.8205
R22 VDD.n1 VDD.t1 1.8205
R23 VDD.n1 VDD.n0 1.8205
R24 VDD.n5 VDD.n4 0.58998
R25 VDD.n16 VDD.n15 0.588573
R26 VDD VDD.n6 0.0760357
R27 VDD VDD.n19 0.0760357
R28 VDD.n19 VDD.n16 0.0551429
R29 VDD.n6 VDD.n5 0.0535357
R30 OUT.n2 OUT.n0 7.06041
R31 OUT.n2 OUT.n1 5.46137
R32 OUT OUT.n2 0.196152
R33 A.n1 A.t3 39.6291
R34 A.n0 A.t1 29.9826
R35 A.t2 A.n0 29.9826
R36 A.n1 A.t2 28.9398
R37 A A.n1 21.7803
R38 A.n0 A.t0 9.1255
R39 VSS.n13 VSS.t6 231.768
R40 VSS.n36 VSS.t11 221.232
R41 VSS.n0 VSS.t12 179.093
R42 VSS.n52 VSS.t4 168.559
R43 VSS.n39 VSS.t9 126.418
R44 VSS.n16 VSS.t2 115.883
R45 VSS.n6 VSS.t0 84.2793
R46 VSS.n30 VSS.t10 73.7444
R47 VSS.n23 VSS.t13 31.605
R48 VSS.n45 VSS.t5 21.0702
R49 VSS VSS.n1 4.66717
R50 VSS VSS.n53 4.47272
R51 VSS.n9 VSS.n5 3.76289
R52 VSS.n22 VSS.n3 3.76289
R53 VSS.n5 VSS.t1 3.2765
R54 VSS.n5 VSS.n4 3.2765
R55 VSS.n3 VSS.t3 3.2765
R56 VSS.n3 VSS.n2 3.2765
R57 VSS.n7 VSS.n6 2.6005
R58 VSS.n12 VSS.n11 2.6005
R59 VSS.n11 VSS.n10 2.6005
R60 VSS.n15 VSS.n14 2.6005
R61 VSS.n14 VSS.n13 2.6005
R62 VSS.n18 VSS.n17 2.6005
R63 VSS.n17 VSS.n16 2.6005
R64 VSS.n21 VSS.n20 2.6005
R65 VSS.n20 VSS.n19 2.6005
R66 VSS.n25 VSS.n24 2.6005
R67 VSS.n24 VSS.n23 2.6005
R68 VSS.n28 VSS.n27 2.6005
R69 VSS.n27 VSS.n26 2.6005
R70 VSS.n1 VSS.n0 2.6005
R71 VSS.n53 VSS.n51 2.6005
R72 VSS.n53 VSS.n52 2.6005
R73 VSS.n50 VSS.n49 2.6005
R74 VSS.n49 VSS.n48 2.6005
R75 VSS.n47 VSS.n46 2.6005
R76 VSS.n46 VSS.n45 2.6005
R77 VSS.n44 VSS.n43 2.6005
R78 VSS.n43 VSS.n42 2.6005
R79 VSS.n41 VSS.n40 2.6005
R80 VSS.n40 VSS.n39 2.6005
R81 VSS.n38 VSS.n37 2.6005
R82 VSS.n37 VSS.n36 2.6005
R83 VSS.n35 VSS.n34 2.6005
R84 VSS.n34 VSS.n33 2.6005
R85 VSS.n31 VSS.n30 2.6005
R86 VSS.n8 VSS.n7 1.64943
R87 VSS.n32 VSS.n31 1.64943
R88 VSS.n35 VSS.n32 0.559135
R89 VSS.n9 VSS.n8 0.535028
R90 VSS.n15 VSS.n12 0.0760357
R91 VSS.n18 VSS.n15 0.0760357
R92 VSS.n21 VSS.n18 0.0760357
R93 VSS.n28 VSS.n25 0.0760357
R94 VSS.n29 VSS.n28 0.0760357
R95 VSS.n51 VSS.n29 0.0760357
R96 VSS.n51 VSS.n50 0.0760357
R97 VSS.n50 VSS.n47 0.0760357
R98 VSS.n47 VSS.n44 0.0760357
R99 VSS.n44 VSS.n41 0.0760357
R100 VSS.n41 VSS.n38 0.0760357
R101 VSS.n38 VSS.n35 0.0760357
R102 VSS.n25 VSS.n22 0.0696071
R103 VSS.n12 VSS.n9 0.0246071
R104 VSS.n22 VSS.n21 0.00692857
R105 B.t2 B.t1 55.0112
R106 B.n0 B.t0 29.9826
R107 B B.n1 27.1952
R108 B.n1 B.t3 22.5523
R109 B.n0 B.t2 9.1255
R110 B.n1 B.n0 7.43086
R111 C.t3 C.t2 68.5684
R112 C C.n1 37.2709
R113 C.n0 C.t3 29.9826
R114 C.n1 C.n0 20.8576
R115 C.n1 C.t0 9.1255
R116 C.n0 C.t1 9.1255
C0 a_168_68# a_648_68# 0.248f
C1 a_24_68# B 0.0309f
C2 OUT B 1.47e-19
C3 a_168_68# A 0.0498f
C4 B a_648_68# 0.0405f
C5 a_168_68# C 0.002f
C6 B A 0.0428f
C7 B C 0.061f
C8 VDD a_24_68# 0.687f
C9 VDD OUT 0.147f
C10 VDD a_648_68# 0.00487f
C11 a_168_68# B 0.193f
C12 OUT a_24_68# 0.259f
C13 VDD A 0.17f
C14 VDD C 0.136f
C15 a_24_68# a_648_68# 0.429f
C16 OUT a_648_68# 0.0155f
C17 a_24_68# A 0.201f
C18 a_24_68# C 0.107f
C19 OUT C 0.0364f
C20 A a_648_68# 0.00131f
C21 VDD a_168_68# 6.85e-19
C22 C a_648_68# 0.0543f
C23 VDD B 0.109f
C24 a_24_68# a_168_68# 0.343f
.ends

