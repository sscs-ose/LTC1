magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1045 -1123 1045 1123
<< metal1 >>
rect -45 117 45 123
rect -45 -117 -39 117
rect 39 -117 45 117
rect -45 -123 45 -117
<< via1 >>
rect -39 -117 39 117
<< metal2 >>
rect -45 117 45 123
rect -45 -117 -39 117
rect 39 -117 45 117
rect -45 -123 45 -117
<< end >>
