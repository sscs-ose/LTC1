** sch_path: /home/shahid/GF180Projects/dff_inv_nand/Xschem/inv_my_pex_tb.sym
**.subckt inv_my_pex_tb
C1 OUT VSS 50f m=1
V1 IN VSS pulse (0 3.3 0 100p 100p 100n 200n)
.save i(v1)
V2 VSS GND 0
.save i(v2)
V3 VDD VSS 3.3
.save i(v3)
x1 VSS IN OUT VDD inv_my_pex
**** begin user architecture code

.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical



.include pex_inv.spice
.control
save all
dc v1 0 3.3 0.1
plot v(IN) v(OUT)

tran 10p 1u
plot v(IN) v(OUT)
*write test_nfet_03v3.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
