magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -20335 -2665 20335 2665
<< psubdiff >>
rect -18335 643 18335 665
rect -18335 597 -18313 643
rect -18267 597 -18189 643
rect -18143 597 -18065 643
rect -18019 597 -17941 643
rect -17895 597 -17817 643
rect -17771 597 -17693 643
rect -17647 597 -17569 643
rect -17523 597 -17445 643
rect -17399 597 -17321 643
rect -17275 597 -17197 643
rect -17151 597 -17073 643
rect -17027 597 -16949 643
rect -16903 597 -16825 643
rect -16779 597 -16701 643
rect -16655 597 -16577 643
rect -16531 597 -16453 643
rect -16407 597 -16329 643
rect -16283 597 -16205 643
rect -16159 597 -16081 643
rect -16035 597 -15957 643
rect -15911 597 -15833 643
rect -15787 597 -15709 643
rect -15663 597 -15585 643
rect -15539 597 -15461 643
rect -15415 597 -15337 643
rect -15291 597 -15213 643
rect -15167 597 -15089 643
rect -15043 597 -14965 643
rect -14919 597 -14841 643
rect -14795 597 -14717 643
rect -14671 597 -14593 643
rect -14547 597 -14469 643
rect -14423 597 -14345 643
rect -14299 597 -14221 643
rect -14175 597 -14097 643
rect -14051 597 -13973 643
rect -13927 597 -13849 643
rect -13803 597 -13725 643
rect -13679 597 -13601 643
rect -13555 597 -13477 643
rect -13431 597 -13353 643
rect -13307 597 -13229 643
rect -13183 597 -13105 643
rect -13059 597 -12981 643
rect -12935 597 -12857 643
rect -12811 597 -12733 643
rect -12687 597 -12609 643
rect -12563 597 -12485 643
rect -12439 597 -12361 643
rect -12315 597 -12237 643
rect -12191 597 -12113 643
rect -12067 597 -11989 643
rect -11943 597 -11865 643
rect -11819 597 -11741 643
rect -11695 597 -11617 643
rect -11571 597 -11493 643
rect -11447 597 -11369 643
rect -11323 597 -11245 643
rect -11199 597 -11121 643
rect -11075 597 -10997 643
rect -10951 597 -10873 643
rect -10827 597 -10749 643
rect -10703 597 -10625 643
rect -10579 597 -10501 643
rect -10455 597 -10377 643
rect -10331 597 -10253 643
rect -10207 597 -10129 643
rect -10083 597 -10005 643
rect -9959 597 -9881 643
rect -9835 597 -9757 643
rect -9711 597 -9633 643
rect -9587 597 -9509 643
rect -9463 597 -9385 643
rect -9339 597 -9261 643
rect -9215 597 -9137 643
rect -9091 597 -9013 643
rect -8967 597 -8889 643
rect -8843 597 -8765 643
rect -8719 597 -8641 643
rect -8595 597 -8517 643
rect -8471 597 -8393 643
rect -8347 597 -8269 643
rect -8223 597 -8145 643
rect -8099 597 -8021 643
rect -7975 597 -7897 643
rect -7851 597 -7773 643
rect -7727 597 -7649 643
rect -7603 597 -7525 643
rect -7479 597 -7401 643
rect -7355 597 -7277 643
rect -7231 597 -7153 643
rect -7107 597 -7029 643
rect -6983 597 -6905 643
rect -6859 597 -6781 643
rect -6735 597 -6657 643
rect -6611 597 -6533 643
rect -6487 597 -6409 643
rect -6363 597 -6285 643
rect -6239 597 -6161 643
rect -6115 597 -6037 643
rect -5991 597 -5913 643
rect -5867 597 -5789 643
rect -5743 597 -5665 643
rect -5619 597 -5541 643
rect -5495 597 -5417 643
rect -5371 597 -5293 643
rect -5247 597 -5169 643
rect -5123 597 -5045 643
rect -4999 597 -4921 643
rect -4875 597 -4797 643
rect -4751 597 -4673 643
rect -4627 597 -4549 643
rect -4503 597 -4425 643
rect -4379 597 -4301 643
rect -4255 597 -4177 643
rect -4131 597 -4053 643
rect -4007 597 -3929 643
rect -3883 597 -3805 643
rect -3759 597 -3681 643
rect -3635 597 -3557 643
rect -3511 597 -3433 643
rect -3387 597 -3309 643
rect -3263 597 -3185 643
rect -3139 597 -3061 643
rect -3015 597 -2937 643
rect -2891 597 -2813 643
rect -2767 597 -2689 643
rect -2643 597 -2565 643
rect -2519 597 -2441 643
rect -2395 597 -2317 643
rect -2271 597 -2193 643
rect -2147 597 -2069 643
rect -2023 597 -1945 643
rect -1899 597 -1821 643
rect -1775 597 -1697 643
rect -1651 597 -1573 643
rect -1527 597 -1449 643
rect -1403 597 -1325 643
rect -1279 597 -1201 643
rect -1155 597 -1077 643
rect -1031 597 -953 643
rect -907 597 -829 643
rect -783 597 -705 643
rect -659 597 -581 643
rect -535 597 -457 643
rect -411 597 -333 643
rect -287 597 -209 643
rect -163 597 -85 643
rect -39 597 39 643
rect 85 597 163 643
rect 209 597 287 643
rect 333 597 411 643
rect 457 597 535 643
rect 581 597 659 643
rect 705 597 783 643
rect 829 597 907 643
rect 953 597 1031 643
rect 1077 597 1155 643
rect 1201 597 1279 643
rect 1325 597 1403 643
rect 1449 597 1527 643
rect 1573 597 1651 643
rect 1697 597 1775 643
rect 1821 597 1899 643
rect 1945 597 2023 643
rect 2069 597 2147 643
rect 2193 597 2271 643
rect 2317 597 2395 643
rect 2441 597 2519 643
rect 2565 597 2643 643
rect 2689 597 2767 643
rect 2813 597 2891 643
rect 2937 597 3015 643
rect 3061 597 3139 643
rect 3185 597 3263 643
rect 3309 597 3387 643
rect 3433 597 3511 643
rect 3557 597 3635 643
rect 3681 597 3759 643
rect 3805 597 3883 643
rect 3929 597 4007 643
rect 4053 597 4131 643
rect 4177 597 4255 643
rect 4301 597 4379 643
rect 4425 597 4503 643
rect 4549 597 4627 643
rect 4673 597 4751 643
rect 4797 597 4875 643
rect 4921 597 4999 643
rect 5045 597 5123 643
rect 5169 597 5247 643
rect 5293 597 5371 643
rect 5417 597 5495 643
rect 5541 597 5619 643
rect 5665 597 5743 643
rect 5789 597 5867 643
rect 5913 597 5991 643
rect 6037 597 6115 643
rect 6161 597 6239 643
rect 6285 597 6363 643
rect 6409 597 6487 643
rect 6533 597 6611 643
rect 6657 597 6735 643
rect 6781 597 6859 643
rect 6905 597 6983 643
rect 7029 597 7107 643
rect 7153 597 7231 643
rect 7277 597 7355 643
rect 7401 597 7479 643
rect 7525 597 7603 643
rect 7649 597 7727 643
rect 7773 597 7851 643
rect 7897 597 7975 643
rect 8021 597 8099 643
rect 8145 597 8223 643
rect 8269 597 8347 643
rect 8393 597 8471 643
rect 8517 597 8595 643
rect 8641 597 8719 643
rect 8765 597 8843 643
rect 8889 597 8967 643
rect 9013 597 9091 643
rect 9137 597 9215 643
rect 9261 597 9339 643
rect 9385 597 9463 643
rect 9509 597 9587 643
rect 9633 597 9711 643
rect 9757 597 9835 643
rect 9881 597 9959 643
rect 10005 597 10083 643
rect 10129 597 10207 643
rect 10253 597 10331 643
rect 10377 597 10455 643
rect 10501 597 10579 643
rect 10625 597 10703 643
rect 10749 597 10827 643
rect 10873 597 10951 643
rect 10997 597 11075 643
rect 11121 597 11199 643
rect 11245 597 11323 643
rect 11369 597 11447 643
rect 11493 597 11571 643
rect 11617 597 11695 643
rect 11741 597 11819 643
rect 11865 597 11943 643
rect 11989 597 12067 643
rect 12113 597 12191 643
rect 12237 597 12315 643
rect 12361 597 12439 643
rect 12485 597 12563 643
rect 12609 597 12687 643
rect 12733 597 12811 643
rect 12857 597 12935 643
rect 12981 597 13059 643
rect 13105 597 13183 643
rect 13229 597 13307 643
rect 13353 597 13431 643
rect 13477 597 13555 643
rect 13601 597 13679 643
rect 13725 597 13803 643
rect 13849 597 13927 643
rect 13973 597 14051 643
rect 14097 597 14175 643
rect 14221 597 14299 643
rect 14345 597 14423 643
rect 14469 597 14547 643
rect 14593 597 14671 643
rect 14717 597 14795 643
rect 14841 597 14919 643
rect 14965 597 15043 643
rect 15089 597 15167 643
rect 15213 597 15291 643
rect 15337 597 15415 643
rect 15461 597 15539 643
rect 15585 597 15663 643
rect 15709 597 15787 643
rect 15833 597 15911 643
rect 15957 597 16035 643
rect 16081 597 16159 643
rect 16205 597 16283 643
rect 16329 597 16407 643
rect 16453 597 16531 643
rect 16577 597 16655 643
rect 16701 597 16779 643
rect 16825 597 16903 643
rect 16949 597 17027 643
rect 17073 597 17151 643
rect 17197 597 17275 643
rect 17321 597 17399 643
rect 17445 597 17523 643
rect 17569 597 17647 643
rect 17693 597 17771 643
rect 17817 597 17895 643
rect 17941 597 18019 643
rect 18065 597 18143 643
rect 18189 597 18267 643
rect 18313 597 18335 643
rect -18335 519 18335 597
rect -18335 473 -18313 519
rect -18267 473 -18189 519
rect -18143 473 -18065 519
rect -18019 473 -17941 519
rect -17895 473 -17817 519
rect -17771 473 -17693 519
rect -17647 473 -17569 519
rect -17523 473 -17445 519
rect -17399 473 -17321 519
rect -17275 473 -17197 519
rect -17151 473 -17073 519
rect -17027 473 -16949 519
rect -16903 473 -16825 519
rect -16779 473 -16701 519
rect -16655 473 -16577 519
rect -16531 473 -16453 519
rect -16407 473 -16329 519
rect -16283 473 -16205 519
rect -16159 473 -16081 519
rect -16035 473 -15957 519
rect -15911 473 -15833 519
rect -15787 473 -15709 519
rect -15663 473 -15585 519
rect -15539 473 -15461 519
rect -15415 473 -15337 519
rect -15291 473 -15213 519
rect -15167 473 -15089 519
rect -15043 473 -14965 519
rect -14919 473 -14841 519
rect -14795 473 -14717 519
rect -14671 473 -14593 519
rect -14547 473 -14469 519
rect -14423 473 -14345 519
rect -14299 473 -14221 519
rect -14175 473 -14097 519
rect -14051 473 -13973 519
rect -13927 473 -13849 519
rect -13803 473 -13725 519
rect -13679 473 -13601 519
rect -13555 473 -13477 519
rect -13431 473 -13353 519
rect -13307 473 -13229 519
rect -13183 473 -13105 519
rect -13059 473 -12981 519
rect -12935 473 -12857 519
rect -12811 473 -12733 519
rect -12687 473 -12609 519
rect -12563 473 -12485 519
rect -12439 473 -12361 519
rect -12315 473 -12237 519
rect -12191 473 -12113 519
rect -12067 473 -11989 519
rect -11943 473 -11865 519
rect -11819 473 -11741 519
rect -11695 473 -11617 519
rect -11571 473 -11493 519
rect -11447 473 -11369 519
rect -11323 473 -11245 519
rect -11199 473 -11121 519
rect -11075 473 -10997 519
rect -10951 473 -10873 519
rect -10827 473 -10749 519
rect -10703 473 -10625 519
rect -10579 473 -10501 519
rect -10455 473 -10377 519
rect -10331 473 -10253 519
rect -10207 473 -10129 519
rect -10083 473 -10005 519
rect -9959 473 -9881 519
rect -9835 473 -9757 519
rect -9711 473 -9633 519
rect -9587 473 -9509 519
rect -9463 473 -9385 519
rect -9339 473 -9261 519
rect -9215 473 -9137 519
rect -9091 473 -9013 519
rect -8967 473 -8889 519
rect -8843 473 -8765 519
rect -8719 473 -8641 519
rect -8595 473 -8517 519
rect -8471 473 -8393 519
rect -8347 473 -8269 519
rect -8223 473 -8145 519
rect -8099 473 -8021 519
rect -7975 473 -7897 519
rect -7851 473 -7773 519
rect -7727 473 -7649 519
rect -7603 473 -7525 519
rect -7479 473 -7401 519
rect -7355 473 -7277 519
rect -7231 473 -7153 519
rect -7107 473 -7029 519
rect -6983 473 -6905 519
rect -6859 473 -6781 519
rect -6735 473 -6657 519
rect -6611 473 -6533 519
rect -6487 473 -6409 519
rect -6363 473 -6285 519
rect -6239 473 -6161 519
rect -6115 473 -6037 519
rect -5991 473 -5913 519
rect -5867 473 -5789 519
rect -5743 473 -5665 519
rect -5619 473 -5541 519
rect -5495 473 -5417 519
rect -5371 473 -5293 519
rect -5247 473 -5169 519
rect -5123 473 -5045 519
rect -4999 473 -4921 519
rect -4875 473 -4797 519
rect -4751 473 -4673 519
rect -4627 473 -4549 519
rect -4503 473 -4425 519
rect -4379 473 -4301 519
rect -4255 473 -4177 519
rect -4131 473 -4053 519
rect -4007 473 -3929 519
rect -3883 473 -3805 519
rect -3759 473 -3681 519
rect -3635 473 -3557 519
rect -3511 473 -3433 519
rect -3387 473 -3309 519
rect -3263 473 -3185 519
rect -3139 473 -3061 519
rect -3015 473 -2937 519
rect -2891 473 -2813 519
rect -2767 473 -2689 519
rect -2643 473 -2565 519
rect -2519 473 -2441 519
rect -2395 473 -2317 519
rect -2271 473 -2193 519
rect -2147 473 -2069 519
rect -2023 473 -1945 519
rect -1899 473 -1821 519
rect -1775 473 -1697 519
rect -1651 473 -1573 519
rect -1527 473 -1449 519
rect -1403 473 -1325 519
rect -1279 473 -1201 519
rect -1155 473 -1077 519
rect -1031 473 -953 519
rect -907 473 -829 519
rect -783 473 -705 519
rect -659 473 -581 519
rect -535 473 -457 519
rect -411 473 -333 519
rect -287 473 -209 519
rect -163 473 -85 519
rect -39 473 39 519
rect 85 473 163 519
rect 209 473 287 519
rect 333 473 411 519
rect 457 473 535 519
rect 581 473 659 519
rect 705 473 783 519
rect 829 473 907 519
rect 953 473 1031 519
rect 1077 473 1155 519
rect 1201 473 1279 519
rect 1325 473 1403 519
rect 1449 473 1527 519
rect 1573 473 1651 519
rect 1697 473 1775 519
rect 1821 473 1899 519
rect 1945 473 2023 519
rect 2069 473 2147 519
rect 2193 473 2271 519
rect 2317 473 2395 519
rect 2441 473 2519 519
rect 2565 473 2643 519
rect 2689 473 2767 519
rect 2813 473 2891 519
rect 2937 473 3015 519
rect 3061 473 3139 519
rect 3185 473 3263 519
rect 3309 473 3387 519
rect 3433 473 3511 519
rect 3557 473 3635 519
rect 3681 473 3759 519
rect 3805 473 3883 519
rect 3929 473 4007 519
rect 4053 473 4131 519
rect 4177 473 4255 519
rect 4301 473 4379 519
rect 4425 473 4503 519
rect 4549 473 4627 519
rect 4673 473 4751 519
rect 4797 473 4875 519
rect 4921 473 4999 519
rect 5045 473 5123 519
rect 5169 473 5247 519
rect 5293 473 5371 519
rect 5417 473 5495 519
rect 5541 473 5619 519
rect 5665 473 5743 519
rect 5789 473 5867 519
rect 5913 473 5991 519
rect 6037 473 6115 519
rect 6161 473 6239 519
rect 6285 473 6363 519
rect 6409 473 6487 519
rect 6533 473 6611 519
rect 6657 473 6735 519
rect 6781 473 6859 519
rect 6905 473 6983 519
rect 7029 473 7107 519
rect 7153 473 7231 519
rect 7277 473 7355 519
rect 7401 473 7479 519
rect 7525 473 7603 519
rect 7649 473 7727 519
rect 7773 473 7851 519
rect 7897 473 7975 519
rect 8021 473 8099 519
rect 8145 473 8223 519
rect 8269 473 8347 519
rect 8393 473 8471 519
rect 8517 473 8595 519
rect 8641 473 8719 519
rect 8765 473 8843 519
rect 8889 473 8967 519
rect 9013 473 9091 519
rect 9137 473 9215 519
rect 9261 473 9339 519
rect 9385 473 9463 519
rect 9509 473 9587 519
rect 9633 473 9711 519
rect 9757 473 9835 519
rect 9881 473 9959 519
rect 10005 473 10083 519
rect 10129 473 10207 519
rect 10253 473 10331 519
rect 10377 473 10455 519
rect 10501 473 10579 519
rect 10625 473 10703 519
rect 10749 473 10827 519
rect 10873 473 10951 519
rect 10997 473 11075 519
rect 11121 473 11199 519
rect 11245 473 11323 519
rect 11369 473 11447 519
rect 11493 473 11571 519
rect 11617 473 11695 519
rect 11741 473 11819 519
rect 11865 473 11943 519
rect 11989 473 12067 519
rect 12113 473 12191 519
rect 12237 473 12315 519
rect 12361 473 12439 519
rect 12485 473 12563 519
rect 12609 473 12687 519
rect 12733 473 12811 519
rect 12857 473 12935 519
rect 12981 473 13059 519
rect 13105 473 13183 519
rect 13229 473 13307 519
rect 13353 473 13431 519
rect 13477 473 13555 519
rect 13601 473 13679 519
rect 13725 473 13803 519
rect 13849 473 13927 519
rect 13973 473 14051 519
rect 14097 473 14175 519
rect 14221 473 14299 519
rect 14345 473 14423 519
rect 14469 473 14547 519
rect 14593 473 14671 519
rect 14717 473 14795 519
rect 14841 473 14919 519
rect 14965 473 15043 519
rect 15089 473 15167 519
rect 15213 473 15291 519
rect 15337 473 15415 519
rect 15461 473 15539 519
rect 15585 473 15663 519
rect 15709 473 15787 519
rect 15833 473 15911 519
rect 15957 473 16035 519
rect 16081 473 16159 519
rect 16205 473 16283 519
rect 16329 473 16407 519
rect 16453 473 16531 519
rect 16577 473 16655 519
rect 16701 473 16779 519
rect 16825 473 16903 519
rect 16949 473 17027 519
rect 17073 473 17151 519
rect 17197 473 17275 519
rect 17321 473 17399 519
rect 17445 473 17523 519
rect 17569 473 17647 519
rect 17693 473 17771 519
rect 17817 473 17895 519
rect 17941 473 18019 519
rect 18065 473 18143 519
rect 18189 473 18267 519
rect 18313 473 18335 519
rect -18335 395 18335 473
rect -18335 349 -18313 395
rect -18267 349 -18189 395
rect -18143 349 -18065 395
rect -18019 349 -17941 395
rect -17895 349 -17817 395
rect -17771 349 -17693 395
rect -17647 349 -17569 395
rect -17523 349 -17445 395
rect -17399 349 -17321 395
rect -17275 349 -17197 395
rect -17151 349 -17073 395
rect -17027 349 -16949 395
rect -16903 349 -16825 395
rect -16779 349 -16701 395
rect -16655 349 -16577 395
rect -16531 349 -16453 395
rect -16407 349 -16329 395
rect -16283 349 -16205 395
rect -16159 349 -16081 395
rect -16035 349 -15957 395
rect -15911 349 -15833 395
rect -15787 349 -15709 395
rect -15663 349 -15585 395
rect -15539 349 -15461 395
rect -15415 349 -15337 395
rect -15291 349 -15213 395
rect -15167 349 -15089 395
rect -15043 349 -14965 395
rect -14919 349 -14841 395
rect -14795 349 -14717 395
rect -14671 349 -14593 395
rect -14547 349 -14469 395
rect -14423 349 -14345 395
rect -14299 349 -14221 395
rect -14175 349 -14097 395
rect -14051 349 -13973 395
rect -13927 349 -13849 395
rect -13803 349 -13725 395
rect -13679 349 -13601 395
rect -13555 349 -13477 395
rect -13431 349 -13353 395
rect -13307 349 -13229 395
rect -13183 349 -13105 395
rect -13059 349 -12981 395
rect -12935 349 -12857 395
rect -12811 349 -12733 395
rect -12687 349 -12609 395
rect -12563 349 -12485 395
rect -12439 349 -12361 395
rect -12315 349 -12237 395
rect -12191 349 -12113 395
rect -12067 349 -11989 395
rect -11943 349 -11865 395
rect -11819 349 -11741 395
rect -11695 349 -11617 395
rect -11571 349 -11493 395
rect -11447 349 -11369 395
rect -11323 349 -11245 395
rect -11199 349 -11121 395
rect -11075 349 -10997 395
rect -10951 349 -10873 395
rect -10827 349 -10749 395
rect -10703 349 -10625 395
rect -10579 349 -10501 395
rect -10455 349 -10377 395
rect -10331 349 -10253 395
rect -10207 349 -10129 395
rect -10083 349 -10005 395
rect -9959 349 -9881 395
rect -9835 349 -9757 395
rect -9711 349 -9633 395
rect -9587 349 -9509 395
rect -9463 349 -9385 395
rect -9339 349 -9261 395
rect -9215 349 -9137 395
rect -9091 349 -9013 395
rect -8967 349 -8889 395
rect -8843 349 -8765 395
rect -8719 349 -8641 395
rect -8595 349 -8517 395
rect -8471 349 -8393 395
rect -8347 349 -8269 395
rect -8223 349 -8145 395
rect -8099 349 -8021 395
rect -7975 349 -7897 395
rect -7851 349 -7773 395
rect -7727 349 -7649 395
rect -7603 349 -7525 395
rect -7479 349 -7401 395
rect -7355 349 -7277 395
rect -7231 349 -7153 395
rect -7107 349 -7029 395
rect -6983 349 -6905 395
rect -6859 349 -6781 395
rect -6735 349 -6657 395
rect -6611 349 -6533 395
rect -6487 349 -6409 395
rect -6363 349 -6285 395
rect -6239 349 -6161 395
rect -6115 349 -6037 395
rect -5991 349 -5913 395
rect -5867 349 -5789 395
rect -5743 349 -5665 395
rect -5619 349 -5541 395
rect -5495 349 -5417 395
rect -5371 349 -5293 395
rect -5247 349 -5169 395
rect -5123 349 -5045 395
rect -4999 349 -4921 395
rect -4875 349 -4797 395
rect -4751 349 -4673 395
rect -4627 349 -4549 395
rect -4503 349 -4425 395
rect -4379 349 -4301 395
rect -4255 349 -4177 395
rect -4131 349 -4053 395
rect -4007 349 -3929 395
rect -3883 349 -3805 395
rect -3759 349 -3681 395
rect -3635 349 -3557 395
rect -3511 349 -3433 395
rect -3387 349 -3309 395
rect -3263 349 -3185 395
rect -3139 349 -3061 395
rect -3015 349 -2937 395
rect -2891 349 -2813 395
rect -2767 349 -2689 395
rect -2643 349 -2565 395
rect -2519 349 -2441 395
rect -2395 349 -2317 395
rect -2271 349 -2193 395
rect -2147 349 -2069 395
rect -2023 349 -1945 395
rect -1899 349 -1821 395
rect -1775 349 -1697 395
rect -1651 349 -1573 395
rect -1527 349 -1449 395
rect -1403 349 -1325 395
rect -1279 349 -1201 395
rect -1155 349 -1077 395
rect -1031 349 -953 395
rect -907 349 -829 395
rect -783 349 -705 395
rect -659 349 -581 395
rect -535 349 -457 395
rect -411 349 -333 395
rect -287 349 -209 395
rect -163 349 -85 395
rect -39 349 39 395
rect 85 349 163 395
rect 209 349 287 395
rect 333 349 411 395
rect 457 349 535 395
rect 581 349 659 395
rect 705 349 783 395
rect 829 349 907 395
rect 953 349 1031 395
rect 1077 349 1155 395
rect 1201 349 1279 395
rect 1325 349 1403 395
rect 1449 349 1527 395
rect 1573 349 1651 395
rect 1697 349 1775 395
rect 1821 349 1899 395
rect 1945 349 2023 395
rect 2069 349 2147 395
rect 2193 349 2271 395
rect 2317 349 2395 395
rect 2441 349 2519 395
rect 2565 349 2643 395
rect 2689 349 2767 395
rect 2813 349 2891 395
rect 2937 349 3015 395
rect 3061 349 3139 395
rect 3185 349 3263 395
rect 3309 349 3387 395
rect 3433 349 3511 395
rect 3557 349 3635 395
rect 3681 349 3759 395
rect 3805 349 3883 395
rect 3929 349 4007 395
rect 4053 349 4131 395
rect 4177 349 4255 395
rect 4301 349 4379 395
rect 4425 349 4503 395
rect 4549 349 4627 395
rect 4673 349 4751 395
rect 4797 349 4875 395
rect 4921 349 4999 395
rect 5045 349 5123 395
rect 5169 349 5247 395
rect 5293 349 5371 395
rect 5417 349 5495 395
rect 5541 349 5619 395
rect 5665 349 5743 395
rect 5789 349 5867 395
rect 5913 349 5991 395
rect 6037 349 6115 395
rect 6161 349 6239 395
rect 6285 349 6363 395
rect 6409 349 6487 395
rect 6533 349 6611 395
rect 6657 349 6735 395
rect 6781 349 6859 395
rect 6905 349 6983 395
rect 7029 349 7107 395
rect 7153 349 7231 395
rect 7277 349 7355 395
rect 7401 349 7479 395
rect 7525 349 7603 395
rect 7649 349 7727 395
rect 7773 349 7851 395
rect 7897 349 7975 395
rect 8021 349 8099 395
rect 8145 349 8223 395
rect 8269 349 8347 395
rect 8393 349 8471 395
rect 8517 349 8595 395
rect 8641 349 8719 395
rect 8765 349 8843 395
rect 8889 349 8967 395
rect 9013 349 9091 395
rect 9137 349 9215 395
rect 9261 349 9339 395
rect 9385 349 9463 395
rect 9509 349 9587 395
rect 9633 349 9711 395
rect 9757 349 9835 395
rect 9881 349 9959 395
rect 10005 349 10083 395
rect 10129 349 10207 395
rect 10253 349 10331 395
rect 10377 349 10455 395
rect 10501 349 10579 395
rect 10625 349 10703 395
rect 10749 349 10827 395
rect 10873 349 10951 395
rect 10997 349 11075 395
rect 11121 349 11199 395
rect 11245 349 11323 395
rect 11369 349 11447 395
rect 11493 349 11571 395
rect 11617 349 11695 395
rect 11741 349 11819 395
rect 11865 349 11943 395
rect 11989 349 12067 395
rect 12113 349 12191 395
rect 12237 349 12315 395
rect 12361 349 12439 395
rect 12485 349 12563 395
rect 12609 349 12687 395
rect 12733 349 12811 395
rect 12857 349 12935 395
rect 12981 349 13059 395
rect 13105 349 13183 395
rect 13229 349 13307 395
rect 13353 349 13431 395
rect 13477 349 13555 395
rect 13601 349 13679 395
rect 13725 349 13803 395
rect 13849 349 13927 395
rect 13973 349 14051 395
rect 14097 349 14175 395
rect 14221 349 14299 395
rect 14345 349 14423 395
rect 14469 349 14547 395
rect 14593 349 14671 395
rect 14717 349 14795 395
rect 14841 349 14919 395
rect 14965 349 15043 395
rect 15089 349 15167 395
rect 15213 349 15291 395
rect 15337 349 15415 395
rect 15461 349 15539 395
rect 15585 349 15663 395
rect 15709 349 15787 395
rect 15833 349 15911 395
rect 15957 349 16035 395
rect 16081 349 16159 395
rect 16205 349 16283 395
rect 16329 349 16407 395
rect 16453 349 16531 395
rect 16577 349 16655 395
rect 16701 349 16779 395
rect 16825 349 16903 395
rect 16949 349 17027 395
rect 17073 349 17151 395
rect 17197 349 17275 395
rect 17321 349 17399 395
rect 17445 349 17523 395
rect 17569 349 17647 395
rect 17693 349 17771 395
rect 17817 349 17895 395
rect 17941 349 18019 395
rect 18065 349 18143 395
rect 18189 349 18267 395
rect 18313 349 18335 395
rect -18335 271 18335 349
rect -18335 225 -18313 271
rect -18267 225 -18189 271
rect -18143 225 -18065 271
rect -18019 225 -17941 271
rect -17895 225 -17817 271
rect -17771 225 -17693 271
rect -17647 225 -17569 271
rect -17523 225 -17445 271
rect -17399 225 -17321 271
rect -17275 225 -17197 271
rect -17151 225 -17073 271
rect -17027 225 -16949 271
rect -16903 225 -16825 271
rect -16779 225 -16701 271
rect -16655 225 -16577 271
rect -16531 225 -16453 271
rect -16407 225 -16329 271
rect -16283 225 -16205 271
rect -16159 225 -16081 271
rect -16035 225 -15957 271
rect -15911 225 -15833 271
rect -15787 225 -15709 271
rect -15663 225 -15585 271
rect -15539 225 -15461 271
rect -15415 225 -15337 271
rect -15291 225 -15213 271
rect -15167 225 -15089 271
rect -15043 225 -14965 271
rect -14919 225 -14841 271
rect -14795 225 -14717 271
rect -14671 225 -14593 271
rect -14547 225 -14469 271
rect -14423 225 -14345 271
rect -14299 225 -14221 271
rect -14175 225 -14097 271
rect -14051 225 -13973 271
rect -13927 225 -13849 271
rect -13803 225 -13725 271
rect -13679 225 -13601 271
rect -13555 225 -13477 271
rect -13431 225 -13353 271
rect -13307 225 -13229 271
rect -13183 225 -13105 271
rect -13059 225 -12981 271
rect -12935 225 -12857 271
rect -12811 225 -12733 271
rect -12687 225 -12609 271
rect -12563 225 -12485 271
rect -12439 225 -12361 271
rect -12315 225 -12237 271
rect -12191 225 -12113 271
rect -12067 225 -11989 271
rect -11943 225 -11865 271
rect -11819 225 -11741 271
rect -11695 225 -11617 271
rect -11571 225 -11493 271
rect -11447 225 -11369 271
rect -11323 225 -11245 271
rect -11199 225 -11121 271
rect -11075 225 -10997 271
rect -10951 225 -10873 271
rect -10827 225 -10749 271
rect -10703 225 -10625 271
rect -10579 225 -10501 271
rect -10455 225 -10377 271
rect -10331 225 -10253 271
rect -10207 225 -10129 271
rect -10083 225 -10005 271
rect -9959 225 -9881 271
rect -9835 225 -9757 271
rect -9711 225 -9633 271
rect -9587 225 -9509 271
rect -9463 225 -9385 271
rect -9339 225 -9261 271
rect -9215 225 -9137 271
rect -9091 225 -9013 271
rect -8967 225 -8889 271
rect -8843 225 -8765 271
rect -8719 225 -8641 271
rect -8595 225 -8517 271
rect -8471 225 -8393 271
rect -8347 225 -8269 271
rect -8223 225 -8145 271
rect -8099 225 -8021 271
rect -7975 225 -7897 271
rect -7851 225 -7773 271
rect -7727 225 -7649 271
rect -7603 225 -7525 271
rect -7479 225 -7401 271
rect -7355 225 -7277 271
rect -7231 225 -7153 271
rect -7107 225 -7029 271
rect -6983 225 -6905 271
rect -6859 225 -6781 271
rect -6735 225 -6657 271
rect -6611 225 -6533 271
rect -6487 225 -6409 271
rect -6363 225 -6285 271
rect -6239 225 -6161 271
rect -6115 225 -6037 271
rect -5991 225 -5913 271
rect -5867 225 -5789 271
rect -5743 225 -5665 271
rect -5619 225 -5541 271
rect -5495 225 -5417 271
rect -5371 225 -5293 271
rect -5247 225 -5169 271
rect -5123 225 -5045 271
rect -4999 225 -4921 271
rect -4875 225 -4797 271
rect -4751 225 -4673 271
rect -4627 225 -4549 271
rect -4503 225 -4425 271
rect -4379 225 -4301 271
rect -4255 225 -4177 271
rect -4131 225 -4053 271
rect -4007 225 -3929 271
rect -3883 225 -3805 271
rect -3759 225 -3681 271
rect -3635 225 -3557 271
rect -3511 225 -3433 271
rect -3387 225 -3309 271
rect -3263 225 -3185 271
rect -3139 225 -3061 271
rect -3015 225 -2937 271
rect -2891 225 -2813 271
rect -2767 225 -2689 271
rect -2643 225 -2565 271
rect -2519 225 -2441 271
rect -2395 225 -2317 271
rect -2271 225 -2193 271
rect -2147 225 -2069 271
rect -2023 225 -1945 271
rect -1899 225 -1821 271
rect -1775 225 -1697 271
rect -1651 225 -1573 271
rect -1527 225 -1449 271
rect -1403 225 -1325 271
rect -1279 225 -1201 271
rect -1155 225 -1077 271
rect -1031 225 -953 271
rect -907 225 -829 271
rect -783 225 -705 271
rect -659 225 -581 271
rect -535 225 -457 271
rect -411 225 -333 271
rect -287 225 -209 271
rect -163 225 -85 271
rect -39 225 39 271
rect 85 225 163 271
rect 209 225 287 271
rect 333 225 411 271
rect 457 225 535 271
rect 581 225 659 271
rect 705 225 783 271
rect 829 225 907 271
rect 953 225 1031 271
rect 1077 225 1155 271
rect 1201 225 1279 271
rect 1325 225 1403 271
rect 1449 225 1527 271
rect 1573 225 1651 271
rect 1697 225 1775 271
rect 1821 225 1899 271
rect 1945 225 2023 271
rect 2069 225 2147 271
rect 2193 225 2271 271
rect 2317 225 2395 271
rect 2441 225 2519 271
rect 2565 225 2643 271
rect 2689 225 2767 271
rect 2813 225 2891 271
rect 2937 225 3015 271
rect 3061 225 3139 271
rect 3185 225 3263 271
rect 3309 225 3387 271
rect 3433 225 3511 271
rect 3557 225 3635 271
rect 3681 225 3759 271
rect 3805 225 3883 271
rect 3929 225 4007 271
rect 4053 225 4131 271
rect 4177 225 4255 271
rect 4301 225 4379 271
rect 4425 225 4503 271
rect 4549 225 4627 271
rect 4673 225 4751 271
rect 4797 225 4875 271
rect 4921 225 4999 271
rect 5045 225 5123 271
rect 5169 225 5247 271
rect 5293 225 5371 271
rect 5417 225 5495 271
rect 5541 225 5619 271
rect 5665 225 5743 271
rect 5789 225 5867 271
rect 5913 225 5991 271
rect 6037 225 6115 271
rect 6161 225 6239 271
rect 6285 225 6363 271
rect 6409 225 6487 271
rect 6533 225 6611 271
rect 6657 225 6735 271
rect 6781 225 6859 271
rect 6905 225 6983 271
rect 7029 225 7107 271
rect 7153 225 7231 271
rect 7277 225 7355 271
rect 7401 225 7479 271
rect 7525 225 7603 271
rect 7649 225 7727 271
rect 7773 225 7851 271
rect 7897 225 7975 271
rect 8021 225 8099 271
rect 8145 225 8223 271
rect 8269 225 8347 271
rect 8393 225 8471 271
rect 8517 225 8595 271
rect 8641 225 8719 271
rect 8765 225 8843 271
rect 8889 225 8967 271
rect 9013 225 9091 271
rect 9137 225 9215 271
rect 9261 225 9339 271
rect 9385 225 9463 271
rect 9509 225 9587 271
rect 9633 225 9711 271
rect 9757 225 9835 271
rect 9881 225 9959 271
rect 10005 225 10083 271
rect 10129 225 10207 271
rect 10253 225 10331 271
rect 10377 225 10455 271
rect 10501 225 10579 271
rect 10625 225 10703 271
rect 10749 225 10827 271
rect 10873 225 10951 271
rect 10997 225 11075 271
rect 11121 225 11199 271
rect 11245 225 11323 271
rect 11369 225 11447 271
rect 11493 225 11571 271
rect 11617 225 11695 271
rect 11741 225 11819 271
rect 11865 225 11943 271
rect 11989 225 12067 271
rect 12113 225 12191 271
rect 12237 225 12315 271
rect 12361 225 12439 271
rect 12485 225 12563 271
rect 12609 225 12687 271
rect 12733 225 12811 271
rect 12857 225 12935 271
rect 12981 225 13059 271
rect 13105 225 13183 271
rect 13229 225 13307 271
rect 13353 225 13431 271
rect 13477 225 13555 271
rect 13601 225 13679 271
rect 13725 225 13803 271
rect 13849 225 13927 271
rect 13973 225 14051 271
rect 14097 225 14175 271
rect 14221 225 14299 271
rect 14345 225 14423 271
rect 14469 225 14547 271
rect 14593 225 14671 271
rect 14717 225 14795 271
rect 14841 225 14919 271
rect 14965 225 15043 271
rect 15089 225 15167 271
rect 15213 225 15291 271
rect 15337 225 15415 271
rect 15461 225 15539 271
rect 15585 225 15663 271
rect 15709 225 15787 271
rect 15833 225 15911 271
rect 15957 225 16035 271
rect 16081 225 16159 271
rect 16205 225 16283 271
rect 16329 225 16407 271
rect 16453 225 16531 271
rect 16577 225 16655 271
rect 16701 225 16779 271
rect 16825 225 16903 271
rect 16949 225 17027 271
rect 17073 225 17151 271
rect 17197 225 17275 271
rect 17321 225 17399 271
rect 17445 225 17523 271
rect 17569 225 17647 271
rect 17693 225 17771 271
rect 17817 225 17895 271
rect 17941 225 18019 271
rect 18065 225 18143 271
rect 18189 225 18267 271
rect 18313 225 18335 271
rect -18335 147 18335 225
rect -18335 101 -18313 147
rect -18267 101 -18189 147
rect -18143 101 -18065 147
rect -18019 101 -17941 147
rect -17895 101 -17817 147
rect -17771 101 -17693 147
rect -17647 101 -17569 147
rect -17523 101 -17445 147
rect -17399 101 -17321 147
rect -17275 101 -17197 147
rect -17151 101 -17073 147
rect -17027 101 -16949 147
rect -16903 101 -16825 147
rect -16779 101 -16701 147
rect -16655 101 -16577 147
rect -16531 101 -16453 147
rect -16407 101 -16329 147
rect -16283 101 -16205 147
rect -16159 101 -16081 147
rect -16035 101 -15957 147
rect -15911 101 -15833 147
rect -15787 101 -15709 147
rect -15663 101 -15585 147
rect -15539 101 -15461 147
rect -15415 101 -15337 147
rect -15291 101 -15213 147
rect -15167 101 -15089 147
rect -15043 101 -14965 147
rect -14919 101 -14841 147
rect -14795 101 -14717 147
rect -14671 101 -14593 147
rect -14547 101 -14469 147
rect -14423 101 -14345 147
rect -14299 101 -14221 147
rect -14175 101 -14097 147
rect -14051 101 -13973 147
rect -13927 101 -13849 147
rect -13803 101 -13725 147
rect -13679 101 -13601 147
rect -13555 101 -13477 147
rect -13431 101 -13353 147
rect -13307 101 -13229 147
rect -13183 101 -13105 147
rect -13059 101 -12981 147
rect -12935 101 -12857 147
rect -12811 101 -12733 147
rect -12687 101 -12609 147
rect -12563 101 -12485 147
rect -12439 101 -12361 147
rect -12315 101 -12237 147
rect -12191 101 -12113 147
rect -12067 101 -11989 147
rect -11943 101 -11865 147
rect -11819 101 -11741 147
rect -11695 101 -11617 147
rect -11571 101 -11493 147
rect -11447 101 -11369 147
rect -11323 101 -11245 147
rect -11199 101 -11121 147
rect -11075 101 -10997 147
rect -10951 101 -10873 147
rect -10827 101 -10749 147
rect -10703 101 -10625 147
rect -10579 101 -10501 147
rect -10455 101 -10377 147
rect -10331 101 -10253 147
rect -10207 101 -10129 147
rect -10083 101 -10005 147
rect -9959 101 -9881 147
rect -9835 101 -9757 147
rect -9711 101 -9633 147
rect -9587 101 -9509 147
rect -9463 101 -9385 147
rect -9339 101 -9261 147
rect -9215 101 -9137 147
rect -9091 101 -9013 147
rect -8967 101 -8889 147
rect -8843 101 -8765 147
rect -8719 101 -8641 147
rect -8595 101 -8517 147
rect -8471 101 -8393 147
rect -8347 101 -8269 147
rect -8223 101 -8145 147
rect -8099 101 -8021 147
rect -7975 101 -7897 147
rect -7851 101 -7773 147
rect -7727 101 -7649 147
rect -7603 101 -7525 147
rect -7479 101 -7401 147
rect -7355 101 -7277 147
rect -7231 101 -7153 147
rect -7107 101 -7029 147
rect -6983 101 -6905 147
rect -6859 101 -6781 147
rect -6735 101 -6657 147
rect -6611 101 -6533 147
rect -6487 101 -6409 147
rect -6363 101 -6285 147
rect -6239 101 -6161 147
rect -6115 101 -6037 147
rect -5991 101 -5913 147
rect -5867 101 -5789 147
rect -5743 101 -5665 147
rect -5619 101 -5541 147
rect -5495 101 -5417 147
rect -5371 101 -5293 147
rect -5247 101 -5169 147
rect -5123 101 -5045 147
rect -4999 101 -4921 147
rect -4875 101 -4797 147
rect -4751 101 -4673 147
rect -4627 101 -4549 147
rect -4503 101 -4425 147
rect -4379 101 -4301 147
rect -4255 101 -4177 147
rect -4131 101 -4053 147
rect -4007 101 -3929 147
rect -3883 101 -3805 147
rect -3759 101 -3681 147
rect -3635 101 -3557 147
rect -3511 101 -3433 147
rect -3387 101 -3309 147
rect -3263 101 -3185 147
rect -3139 101 -3061 147
rect -3015 101 -2937 147
rect -2891 101 -2813 147
rect -2767 101 -2689 147
rect -2643 101 -2565 147
rect -2519 101 -2441 147
rect -2395 101 -2317 147
rect -2271 101 -2193 147
rect -2147 101 -2069 147
rect -2023 101 -1945 147
rect -1899 101 -1821 147
rect -1775 101 -1697 147
rect -1651 101 -1573 147
rect -1527 101 -1449 147
rect -1403 101 -1325 147
rect -1279 101 -1201 147
rect -1155 101 -1077 147
rect -1031 101 -953 147
rect -907 101 -829 147
rect -783 101 -705 147
rect -659 101 -581 147
rect -535 101 -457 147
rect -411 101 -333 147
rect -287 101 -209 147
rect -163 101 -85 147
rect -39 101 39 147
rect 85 101 163 147
rect 209 101 287 147
rect 333 101 411 147
rect 457 101 535 147
rect 581 101 659 147
rect 705 101 783 147
rect 829 101 907 147
rect 953 101 1031 147
rect 1077 101 1155 147
rect 1201 101 1279 147
rect 1325 101 1403 147
rect 1449 101 1527 147
rect 1573 101 1651 147
rect 1697 101 1775 147
rect 1821 101 1899 147
rect 1945 101 2023 147
rect 2069 101 2147 147
rect 2193 101 2271 147
rect 2317 101 2395 147
rect 2441 101 2519 147
rect 2565 101 2643 147
rect 2689 101 2767 147
rect 2813 101 2891 147
rect 2937 101 3015 147
rect 3061 101 3139 147
rect 3185 101 3263 147
rect 3309 101 3387 147
rect 3433 101 3511 147
rect 3557 101 3635 147
rect 3681 101 3759 147
rect 3805 101 3883 147
rect 3929 101 4007 147
rect 4053 101 4131 147
rect 4177 101 4255 147
rect 4301 101 4379 147
rect 4425 101 4503 147
rect 4549 101 4627 147
rect 4673 101 4751 147
rect 4797 101 4875 147
rect 4921 101 4999 147
rect 5045 101 5123 147
rect 5169 101 5247 147
rect 5293 101 5371 147
rect 5417 101 5495 147
rect 5541 101 5619 147
rect 5665 101 5743 147
rect 5789 101 5867 147
rect 5913 101 5991 147
rect 6037 101 6115 147
rect 6161 101 6239 147
rect 6285 101 6363 147
rect 6409 101 6487 147
rect 6533 101 6611 147
rect 6657 101 6735 147
rect 6781 101 6859 147
rect 6905 101 6983 147
rect 7029 101 7107 147
rect 7153 101 7231 147
rect 7277 101 7355 147
rect 7401 101 7479 147
rect 7525 101 7603 147
rect 7649 101 7727 147
rect 7773 101 7851 147
rect 7897 101 7975 147
rect 8021 101 8099 147
rect 8145 101 8223 147
rect 8269 101 8347 147
rect 8393 101 8471 147
rect 8517 101 8595 147
rect 8641 101 8719 147
rect 8765 101 8843 147
rect 8889 101 8967 147
rect 9013 101 9091 147
rect 9137 101 9215 147
rect 9261 101 9339 147
rect 9385 101 9463 147
rect 9509 101 9587 147
rect 9633 101 9711 147
rect 9757 101 9835 147
rect 9881 101 9959 147
rect 10005 101 10083 147
rect 10129 101 10207 147
rect 10253 101 10331 147
rect 10377 101 10455 147
rect 10501 101 10579 147
rect 10625 101 10703 147
rect 10749 101 10827 147
rect 10873 101 10951 147
rect 10997 101 11075 147
rect 11121 101 11199 147
rect 11245 101 11323 147
rect 11369 101 11447 147
rect 11493 101 11571 147
rect 11617 101 11695 147
rect 11741 101 11819 147
rect 11865 101 11943 147
rect 11989 101 12067 147
rect 12113 101 12191 147
rect 12237 101 12315 147
rect 12361 101 12439 147
rect 12485 101 12563 147
rect 12609 101 12687 147
rect 12733 101 12811 147
rect 12857 101 12935 147
rect 12981 101 13059 147
rect 13105 101 13183 147
rect 13229 101 13307 147
rect 13353 101 13431 147
rect 13477 101 13555 147
rect 13601 101 13679 147
rect 13725 101 13803 147
rect 13849 101 13927 147
rect 13973 101 14051 147
rect 14097 101 14175 147
rect 14221 101 14299 147
rect 14345 101 14423 147
rect 14469 101 14547 147
rect 14593 101 14671 147
rect 14717 101 14795 147
rect 14841 101 14919 147
rect 14965 101 15043 147
rect 15089 101 15167 147
rect 15213 101 15291 147
rect 15337 101 15415 147
rect 15461 101 15539 147
rect 15585 101 15663 147
rect 15709 101 15787 147
rect 15833 101 15911 147
rect 15957 101 16035 147
rect 16081 101 16159 147
rect 16205 101 16283 147
rect 16329 101 16407 147
rect 16453 101 16531 147
rect 16577 101 16655 147
rect 16701 101 16779 147
rect 16825 101 16903 147
rect 16949 101 17027 147
rect 17073 101 17151 147
rect 17197 101 17275 147
rect 17321 101 17399 147
rect 17445 101 17523 147
rect 17569 101 17647 147
rect 17693 101 17771 147
rect 17817 101 17895 147
rect 17941 101 18019 147
rect 18065 101 18143 147
rect 18189 101 18267 147
rect 18313 101 18335 147
rect -18335 23 18335 101
rect -18335 -23 -18313 23
rect -18267 -23 -18189 23
rect -18143 -23 -18065 23
rect -18019 -23 -17941 23
rect -17895 -23 -17817 23
rect -17771 -23 -17693 23
rect -17647 -23 -17569 23
rect -17523 -23 -17445 23
rect -17399 -23 -17321 23
rect -17275 -23 -17197 23
rect -17151 -23 -17073 23
rect -17027 -23 -16949 23
rect -16903 -23 -16825 23
rect -16779 -23 -16701 23
rect -16655 -23 -16577 23
rect -16531 -23 -16453 23
rect -16407 -23 -16329 23
rect -16283 -23 -16205 23
rect -16159 -23 -16081 23
rect -16035 -23 -15957 23
rect -15911 -23 -15833 23
rect -15787 -23 -15709 23
rect -15663 -23 -15585 23
rect -15539 -23 -15461 23
rect -15415 -23 -15337 23
rect -15291 -23 -15213 23
rect -15167 -23 -15089 23
rect -15043 -23 -14965 23
rect -14919 -23 -14841 23
rect -14795 -23 -14717 23
rect -14671 -23 -14593 23
rect -14547 -23 -14469 23
rect -14423 -23 -14345 23
rect -14299 -23 -14221 23
rect -14175 -23 -14097 23
rect -14051 -23 -13973 23
rect -13927 -23 -13849 23
rect -13803 -23 -13725 23
rect -13679 -23 -13601 23
rect -13555 -23 -13477 23
rect -13431 -23 -13353 23
rect -13307 -23 -13229 23
rect -13183 -23 -13105 23
rect -13059 -23 -12981 23
rect -12935 -23 -12857 23
rect -12811 -23 -12733 23
rect -12687 -23 -12609 23
rect -12563 -23 -12485 23
rect -12439 -23 -12361 23
rect -12315 -23 -12237 23
rect -12191 -23 -12113 23
rect -12067 -23 -11989 23
rect -11943 -23 -11865 23
rect -11819 -23 -11741 23
rect -11695 -23 -11617 23
rect -11571 -23 -11493 23
rect -11447 -23 -11369 23
rect -11323 -23 -11245 23
rect -11199 -23 -11121 23
rect -11075 -23 -10997 23
rect -10951 -23 -10873 23
rect -10827 -23 -10749 23
rect -10703 -23 -10625 23
rect -10579 -23 -10501 23
rect -10455 -23 -10377 23
rect -10331 -23 -10253 23
rect -10207 -23 -10129 23
rect -10083 -23 -10005 23
rect -9959 -23 -9881 23
rect -9835 -23 -9757 23
rect -9711 -23 -9633 23
rect -9587 -23 -9509 23
rect -9463 -23 -9385 23
rect -9339 -23 -9261 23
rect -9215 -23 -9137 23
rect -9091 -23 -9013 23
rect -8967 -23 -8889 23
rect -8843 -23 -8765 23
rect -8719 -23 -8641 23
rect -8595 -23 -8517 23
rect -8471 -23 -8393 23
rect -8347 -23 -8269 23
rect -8223 -23 -8145 23
rect -8099 -23 -8021 23
rect -7975 -23 -7897 23
rect -7851 -23 -7773 23
rect -7727 -23 -7649 23
rect -7603 -23 -7525 23
rect -7479 -23 -7401 23
rect -7355 -23 -7277 23
rect -7231 -23 -7153 23
rect -7107 -23 -7029 23
rect -6983 -23 -6905 23
rect -6859 -23 -6781 23
rect -6735 -23 -6657 23
rect -6611 -23 -6533 23
rect -6487 -23 -6409 23
rect -6363 -23 -6285 23
rect -6239 -23 -6161 23
rect -6115 -23 -6037 23
rect -5991 -23 -5913 23
rect -5867 -23 -5789 23
rect -5743 -23 -5665 23
rect -5619 -23 -5541 23
rect -5495 -23 -5417 23
rect -5371 -23 -5293 23
rect -5247 -23 -5169 23
rect -5123 -23 -5045 23
rect -4999 -23 -4921 23
rect -4875 -23 -4797 23
rect -4751 -23 -4673 23
rect -4627 -23 -4549 23
rect -4503 -23 -4425 23
rect -4379 -23 -4301 23
rect -4255 -23 -4177 23
rect -4131 -23 -4053 23
rect -4007 -23 -3929 23
rect -3883 -23 -3805 23
rect -3759 -23 -3681 23
rect -3635 -23 -3557 23
rect -3511 -23 -3433 23
rect -3387 -23 -3309 23
rect -3263 -23 -3185 23
rect -3139 -23 -3061 23
rect -3015 -23 -2937 23
rect -2891 -23 -2813 23
rect -2767 -23 -2689 23
rect -2643 -23 -2565 23
rect -2519 -23 -2441 23
rect -2395 -23 -2317 23
rect -2271 -23 -2193 23
rect -2147 -23 -2069 23
rect -2023 -23 -1945 23
rect -1899 -23 -1821 23
rect -1775 -23 -1697 23
rect -1651 -23 -1573 23
rect -1527 -23 -1449 23
rect -1403 -23 -1325 23
rect -1279 -23 -1201 23
rect -1155 -23 -1077 23
rect -1031 -23 -953 23
rect -907 -23 -829 23
rect -783 -23 -705 23
rect -659 -23 -581 23
rect -535 -23 -457 23
rect -411 -23 -333 23
rect -287 -23 -209 23
rect -163 -23 -85 23
rect -39 -23 39 23
rect 85 -23 163 23
rect 209 -23 287 23
rect 333 -23 411 23
rect 457 -23 535 23
rect 581 -23 659 23
rect 705 -23 783 23
rect 829 -23 907 23
rect 953 -23 1031 23
rect 1077 -23 1155 23
rect 1201 -23 1279 23
rect 1325 -23 1403 23
rect 1449 -23 1527 23
rect 1573 -23 1651 23
rect 1697 -23 1775 23
rect 1821 -23 1899 23
rect 1945 -23 2023 23
rect 2069 -23 2147 23
rect 2193 -23 2271 23
rect 2317 -23 2395 23
rect 2441 -23 2519 23
rect 2565 -23 2643 23
rect 2689 -23 2767 23
rect 2813 -23 2891 23
rect 2937 -23 3015 23
rect 3061 -23 3139 23
rect 3185 -23 3263 23
rect 3309 -23 3387 23
rect 3433 -23 3511 23
rect 3557 -23 3635 23
rect 3681 -23 3759 23
rect 3805 -23 3883 23
rect 3929 -23 4007 23
rect 4053 -23 4131 23
rect 4177 -23 4255 23
rect 4301 -23 4379 23
rect 4425 -23 4503 23
rect 4549 -23 4627 23
rect 4673 -23 4751 23
rect 4797 -23 4875 23
rect 4921 -23 4999 23
rect 5045 -23 5123 23
rect 5169 -23 5247 23
rect 5293 -23 5371 23
rect 5417 -23 5495 23
rect 5541 -23 5619 23
rect 5665 -23 5743 23
rect 5789 -23 5867 23
rect 5913 -23 5991 23
rect 6037 -23 6115 23
rect 6161 -23 6239 23
rect 6285 -23 6363 23
rect 6409 -23 6487 23
rect 6533 -23 6611 23
rect 6657 -23 6735 23
rect 6781 -23 6859 23
rect 6905 -23 6983 23
rect 7029 -23 7107 23
rect 7153 -23 7231 23
rect 7277 -23 7355 23
rect 7401 -23 7479 23
rect 7525 -23 7603 23
rect 7649 -23 7727 23
rect 7773 -23 7851 23
rect 7897 -23 7975 23
rect 8021 -23 8099 23
rect 8145 -23 8223 23
rect 8269 -23 8347 23
rect 8393 -23 8471 23
rect 8517 -23 8595 23
rect 8641 -23 8719 23
rect 8765 -23 8843 23
rect 8889 -23 8967 23
rect 9013 -23 9091 23
rect 9137 -23 9215 23
rect 9261 -23 9339 23
rect 9385 -23 9463 23
rect 9509 -23 9587 23
rect 9633 -23 9711 23
rect 9757 -23 9835 23
rect 9881 -23 9959 23
rect 10005 -23 10083 23
rect 10129 -23 10207 23
rect 10253 -23 10331 23
rect 10377 -23 10455 23
rect 10501 -23 10579 23
rect 10625 -23 10703 23
rect 10749 -23 10827 23
rect 10873 -23 10951 23
rect 10997 -23 11075 23
rect 11121 -23 11199 23
rect 11245 -23 11323 23
rect 11369 -23 11447 23
rect 11493 -23 11571 23
rect 11617 -23 11695 23
rect 11741 -23 11819 23
rect 11865 -23 11943 23
rect 11989 -23 12067 23
rect 12113 -23 12191 23
rect 12237 -23 12315 23
rect 12361 -23 12439 23
rect 12485 -23 12563 23
rect 12609 -23 12687 23
rect 12733 -23 12811 23
rect 12857 -23 12935 23
rect 12981 -23 13059 23
rect 13105 -23 13183 23
rect 13229 -23 13307 23
rect 13353 -23 13431 23
rect 13477 -23 13555 23
rect 13601 -23 13679 23
rect 13725 -23 13803 23
rect 13849 -23 13927 23
rect 13973 -23 14051 23
rect 14097 -23 14175 23
rect 14221 -23 14299 23
rect 14345 -23 14423 23
rect 14469 -23 14547 23
rect 14593 -23 14671 23
rect 14717 -23 14795 23
rect 14841 -23 14919 23
rect 14965 -23 15043 23
rect 15089 -23 15167 23
rect 15213 -23 15291 23
rect 15337 -23 15415 23
rect 15461 -23 15539 23
rect 15585 -23 15663 23
rect 15709 -23 15787 23
rect 15833 -23 15911 23
rect 15957 -23 16035 23
rect 16081 -23 16159 23
rect 16205 -23 16283 23
rect 16329 -23 16407 23
rect 16453 -23 16531 23
rect 16577 -23 16655 23
rect 16701 -23 16779 23
rect 16825 -23 16903 23
rect 16949 -23 17027 23
rect 17073 -23 17151 23
rect 17197 -23 17275 23
rect 17321 -23 17399 23
rect 17445 -23 17523 23
rect 17569 -23 17647 23
rect 17693 -23 17771 23
rect 17817 -23 17895 23
rect 17941 -23 18019 23
rect 18065 -23 18143 23
rect 18189 -23 18267 23
rect 18313 -23 18335 23
rect -18335 -101 18335 -23
rect -18335 -147 -18313 -101
rect -18267 -147 -18189 -101
rect -18143 -147 -18065 -101
rect -18019 -147 -17941 -101
rect -17895 -147 -17817 -101
rect -17771 -147 -17693 -101
rect -17647 -147 -17569 -101
rect -17523 -147 -17445 -101
rect -17399 -147 -17321 -101
rect -17275 -147 -17197 -101
rect -17151 -147 -17073 -101
rect -17027 -147 -16949 -101
rect -16903 -147 -16825 -101
rect -16779 -147 -16701 -101
rect -16655 -147 -16577 -101
rect -16531 -147 -16453 -101
rect -16407 -147 -16329 -101
rect -16283 -147 -16205 -101
rect -16159 -147 -16081 -101
rect -16035 -147 -15957 -101
rect -15911 -147 -15833 -101
rect -15787 -147 -15709 -101
rect -15663 -147 -15585 -101
rect -15539 -147 -15461 -101
rect -15415 -147 -15337 -101
rect -15291 -147 -15213 -101
rect -15167 -147 -15089 -101
rect -15043 -147 -14965 -101
rect -14919 -147 -14841 -101
rect -14795 -147 -14717 -101
rect -14671 -147 -14593 -101
rect -14547 -147 -14469 -101
rect -14423 -147 -14345 -101
rect -14299 -147 -14221 -101
rect -14175 -147 -14097 -101
rect -14051 -147 -13973 -101
rect -13927 -147 -13849 -101
rect -13803 -147 -13725 -101
rect -13679 -147 -13601 -101
rect -13555 -147 -13477 -101
rect -13431 -147 -13353 -101
rect -13307 -147 -13229 -101
rect -13183 -147 -13105 -101
rect -13059 -147 -12981 -101
rect -12935 -147 -12857 -101
rect -12811 -147 -12733 -101
rect -12687 -147 -12609 -101
rect -12563 -147 -12485 -101
rect -12439 -147 -12361 -101
rect -12315 -147 -12237 -101
rect -12191 -147 -12113 -101
rect -12067 -147 -11989 -101
rect -11943 -147 -11865 -101
rect -11819 -147 -11741 -101
rect -11695 -147 -11617 -101
rect -11571 -147 -11493 -101
rect -11447 -147 -11369 -101
rect -11323 -147 -11245 -101
rect -11199 -147 -11121 -101
rect -11075 -147 -10997 -101
rect -10951 -147 -10873 -101
rect -10827 -147 -10749 -101
rect -10703 -147 -10625 -101
rect -10579 -147 -10501 -101
rect -10455 -147 -10377 -101
rect -10331 -147 -10253 -101
rect -10207 -147 -10129 -101
rect -10083 -147 -10005 -101
rect -9959 -147 -9881 -101
rect -9835 -147 -9757 -101
rect -9711 -147 -9633 -101
rect -9587 -147 -9509 -101
rect -9463 -147 -9385 -101
rect -9339 -147 -9261 -101
rect -9215 -147 -9137 -101
rect -9091 -147 -9013 -101
rect -8967 -147 -8889 -101
rect -8843 -147 -8765 -101
rect -8719 -147 -8641 -101
rect -8595 -147 -8517 -101
rect -8471 -147 -8393 -101
rect -8347 -147 -8269 -101
rect -8223 -147 -8145 -101
rect -8099 -147 -8021 -101
rect -7975 -147 -7897 -101
rect -7851 -147 -7773 -101
rect -7727 -147 -7649 -101
rect -7603 -147 -7525 -101
rect -7479 -147 -7401 -101
rect -7355 -147 -7277 -101
rect -7231 -147 -7153 -101
rect -7107 -147 -7029 -101
rect -6983 -147 -6905 -101
rect -6859 -147 -6781 -101
rect -6735 -147 -6657 -101
rect -6611 -147 -6533 -101
rect -6487 -147 -6409 -101
rect -6363 -147 -6285 -101
rect -6239 -147 -6161 -101
rect -6115 -147 -6037 -101
rect -5991 -147 -5913 -101
rect -5867 -147 -5789 -101
rect -5743 -147 -5665 -101
rect -5619 -147 -5541 -101
rect -5495 -147 -5417 -101
rect -5371 -147 -5293 -101
rect -5247 -147 -5169 -101
rect -5123 -147 -5045 -101
rect -4999 -147 -4921 -101
rect -4875 -147 -4797 -101
rect -4751 -147 -4673 -101
rect -4627 -147 -4549 -101
rect -4503 -147 -4425 -101
rect -4379 -147 -4301 -101
rect -4255 -147 -4177 -101
rect -4131 -147 -4053 -101
rect -4007 -147 -3929 -101
rect -3883 -147 -3805 -101
rect -3759 -147 -3681 -101
rect -3635 -147 -3557 -101
rect -3511 -147 -3433 -101
rect -3387 -147 -3309 -101
rect -3263 -147 -3185 -101
rect -3139 -147 -3061 -101
rect -3015 -147 -2937 -101
rect -2891 -147 -2813 -101
rect -2767 -147 -2689 -101
rect -2643 -147 -2565 -101
rect -2519 -147 -2441 -101
rect -2395 -147 -2317 -101
rect -2271 -147 -2193 -101
rect -2147 -147 -2069 -101
rect -2023 -147 -1945 -101
rect -1899 -147 -1821 -101
rect -1775 -147 -1697 -101
rect -1651 -147 -1573 -101
rect -1527 -147 -1449 -101
rect -1403 -147 -1325 -101
rect -1279 -147 -1201 -101
rect -1155 -147 -1077 -101
rect -1031 -147 -953 -101
rect -907 -147 -829 -101
rect -783 -147 -705 -101
rect -659 -147 -581 -101
rect -535 -147 -457 -101
rect -411 -147 -333 -101
rect -287 -147 -209 -101
rect -163 -147 -85 -101
rect -39 -147 39 -101
rect 85 -147 163 -101
rect 209 -147 287 -101
rect 333 -147 411 -101
rect 457 -147 535 -101
rect 581 -147 659 -101
rect 705 -147 783 -101
rect 829 -147 907 -101
rect 953 -147 1031 -101
rect 1077 -147 1155 -101
rect 1201 -147 1279 -101
rect 1325 -147 1403 -101
rect 1449 -147 1527 -101
rect 1573 -147 1651 -101
rect 1697 -147 1775 -101
rect 1821 -147 1899 -101
rect 1945 -147 2023 -101
rect 2069 -147 2147 -101
rect 2193 -147 2271 -101
rect 2317 -147 2395 -101
rect 2441 -147 2519 -101
rect 2565 -147 2643 -101
rect 2689 -147 2767 -101
rect 2813 -147 2891 -101
rect 2937 -147 3015 -101
rect 3061 -147 3139 -101
rect 3185 -147 3263 -101
rect 3309 -147 3387 -101
rect 3433 -147 3511 -101
rect 3557 -147 3635 -101
rect 3681 -147 3759 -101
rect 3805 -147 3883 -101
rect 3929 -147 4007 -101
rect 4053 -147 4131 -101
rect 4177 -147 4255 -101
rect 4301 -147 4379 -101
rect 4425 -147 4503 -101
rect 4549 -147 4627 -101
rect 4673 -147 4751 -101
rect 4797 -147 4875 -101
rect 4921 -147 4999 -101
rect 5045 -147 5123 -101
rect 5169 -147 5247 -101
rect 5293 -147 5371 -101
rect 5417 -147 5495 -101
rect 5541 -147 5619 -101
rect 5665 -147 5743 -101
rect 5789 -147 5867 -101
rect 5913 -147 5991 -101
rect 6037 -147 6115 -101
rect 6161 -147 6239 -101
rect 6285 -147 6363 -101
rect 6409 -147 6487 -101
rect 6533 -147 6611 -101
rect 6657 -147 6735 -101
rect 6781 -147 6859 -101
rect 6905 -147 6983 -101
rect 7029 -147 7107 -101
rect 7153 -147 7231 -101
rect 7277 -147 7355 -101
rect 7401 -147 7479 -101
rect 7525 -147 7603 -101
rect 7649 -147 7727 -101
rect 7773 -147 7851 -101
rect 7897 -147 7975 -101
rect 8021 -147 8099 -101
rect 8145 -147 8223 -101
rect 8269 -147 8347 -101
rect 8393 -147 8471 -101
rect 8517 -147 8595 -101
rect 8641 -147 8719 -101
rect 8765 -147 8843 -101
rect 8889 -147 8967 -101
rect 9013 -147 9091 -101
rect 9137 -147 9215 -101
rect 9261 -147 9339 -101
rect 9385 -147 9463 -101
rect 9509 -147 9587 -101
rect 9633 -147 9711 -101
rect 9757 -147 9835 -101
rect 9881 -147 9959 -101
rect 10005 -147 10083 -101
rect 10129 -147 10207 -101
rect 10253 -147 10331 -101
rect 10377 -147 10455 -101
rect 10501 -147 10579 -101
rect 10625 -147 10703 -101
rect 10749 -147 10827 -101
rect 10873 -147 10951 -101
rect 10997 -147 11075 -101
rect 11121 -147 11199 -101
rect 11245 -147 11323 -101
rect 11369 -147 11447 -101
rect 11493 -147 11571 -101
rect 11617 -147 11695 -101
rect 11741 -147 11819 -101
rect 11865 -147 11943 -101
rect 11989 -147 12067 -101
rect 12113 -147 12191 -101
rect 12237 -147 12315 -101
rect 12361 -147 12439 -101
rect 12485 -147 12563 -101
rect 12609 -147 12687 -101
rect 12733 -147 12811 -101
rect 12857 -147 12935 -101
rect 12981 -147 13059 -101
rect 13105 -147 13183 -101
rect 13229 -147 13307 -101
rect 13353 -147 13431 -101
rect 13477 -147 13555 -101
rect 13601 -147 13679 -101
rect 13725 -147 13803 -101
rect 13849 -147 13927 -101
rect 13973 -147 14051 -101
rect 14097 -147 14175 -101
rect 14221 -147 14299 -101
rect 14345 -147 14423 -101
rect 14469 -147 14547 -101
rect 14593 -147 14671 -101
rect 14717 -147 14795 -101
rect 14841 -147 14919 -101
rect 14965 -147 15043 -101
rect 15089 -147 15167 -101
rect 15213 -147 15291 -101
rect 15337 -147 15415 -101
rect 15461 -147 15539 -101
rect 15585 -147 15663 -101
rect 15709 -147 15787 -101
rect 15833 -147 15911 -101
rect 15957 -147 16035 -101
rect 16081 -147 16159 -101
rect 16205 -147 16283 -101
rect 16329 -147 16407 -101
rect 16453 -147 16531 -101
rect 16577 -147 16655 -101
rect 16701 -147 16779 -101
rect 16825 -147 16903 -101
rect 16949 -147 17027 -101
rect 17073 -147 17151 -101
rect 17197 -147 17275 -101
rect 17321 -147 17399 -101
rect 17445 -147 17523 -101
rect 17569 -147 17647 -101
rect 17693 -147 17771 -101
rect 17817 -147 17895 -101
rect 17941 -147 18019 -101
rect 18065 -147 18143 -101
rect 18189 -147 18267 -101
rect 18313 -147 18335 -101
rect -18335 -225 18335 -147
rect -18335 -271 -18313 -225
rect -18267 -271 -18189 -225
rect -18143 -271 -18065 -225
rect -18019 -271 -17941 -225
rect -17895 -271 -17817 -225
rect -17771 -271 -17693 -225
rect -17647 -271 -17569 -225
rect -17523 -271 -17445 -225
rect -17399 -271 -17321 -225
rect -17275 -271 -17197 -225
rect -17151 -271 -17073 -225
rect -17027 -271 -16949 -225
rect -16903 -271 -16825 -225
rect -16779 -271 -16701 -225
rect -16655 -271 -16577 -225
rect -16531 -271 -16453 -225
rect -16407 -271 -16329 -225
rect -16283 -271 -16205 -225
rect -16159 -271 -16081 -225
rect -16035 -271 -15957 -225
rect -15911 -271 -15833 -225
rect -15787 -271 -15709 -225
rect -15663 -271 -15585 -225
rect -15539 -271 -15461 -225
rect -15415 -271 -15337 -225
rect -15291 -271 -15213 -225
rect -15167 -271 -15089 -225
rect -15043 -271 -14965 -225
rect -14919 -271 -14841 -225
rect -14795 -271 -14717 -225
rect -14671 -271 -14593 -225
rect -14547 -271 -14469 -225
rect -14423 -271 -14345 -225
rect -14299 -271 -14221 -225
rect -14175 -271 -14097 -225
rect -14051 -271 -13973 -225
rect -13927 -271 -13849 -225
rect -13803 -271 -13725 -225
rect -13679 -271 -13601 -225
rect -13555 -271 -13477 -225
rect -13431 -271 -13353 -225
rect -13307 -271 -13229 -225
rect -13183 -271 -13105 -225
rect -13059 -271 -12981 -225
rect -12935 -271 -12857 -225
rect -12811 -271 -12733 -225
rect -12687 -271 -12609 -225
rect -12563 -271 -12485 -225
rect -12439 -271 -12361 -225
rect -12315 -271 -12237 -225
rect -12191 -271 -12113 -225
rect -12067 -271 -11989 -225
rect -11943 -271 -11865 -225
rect -11819 -271 -11741 -225
rect -11695 -271 -11617 -225
rect -11571 -271 -11493 -225
rect -11447 -271 -11369 -225
rect -11323 -271 -11245 -225
rect -11199 -271 -11121 -225
rect -11075 -271 -10997 -225
rect -10951 -271 -10873 -225
rect -10827 -271 -10749 -225
rect -10703 -271 -10625 -225
rect -10579 -271 -10501 -225
rect -10455 -271 -10377 -225
rect -10331 -271 -10253 -225
rect -10207 -271 -10129 -225
rect -10083 -271 -10005 -225
rect -9959 -271 -9881 -225
rect -9835 -271 -9757 -225
rect -9711 -271 -9633 -225
rect -9587 -271 -9509 -225
rect -9463 -271 -9385 -225
rect -9339 -271 -9261 -225
rect -9215 -271 -9137 -225
rect -9091 -271 -9013 -225
rect -8967 -271 -8889 -225
rect -8843 -271 -8765 -225
rect -8719 -271 -8641 -225
rect -8595 -271 -8517 -225
rect -8471 -271 -8393 -225
rect -8347 -271 -8269 -225
rect -8223 -271 -8145 -225
rect -8099 -271 -8021 -225
rect -7975 -271 -7897 -225
rect -7851 -271 -7773 -225
rect -7727 -271 -7649 -225
rect -7603 -271 -7525 -225
rect -7479 -271 -7401 -225
rect -7355 -271 -7277 -225
rect -7231 -271 -7153 -225
rect -7107 -271 -7029 -225
rect -6983 -271 -6905 -225
rect -6859 -271 -6781 -225
rect -6735 -271 -6657 -225
rect -6611 -271 -6533 -225
rect -6487 -271 -6409 -225
rect -6363 -271 -6285 -225
rect -6239 -271 -6161 -225
rect -6115 -271 -6037 -225
rect -5991 -271 -5913 -225
rect -5867 -271 -5789 -225
rect -5743 -271 -5665 -225
rect -5619 -271 -5541 -225
rect -5495 -271 -5417 -225
rect -5371 -271 -5293 -225
rect -5247 -271 -5169 -225
rect -5123 -271 -5045 -225
rect -4999 -271 -4921 -225
rect -4875 -271 -4797 -225
rect -4751 -271 -4673 -225
rect -4627 -271 -4549 -225
rect -4503 -271 -4425 -225
rect -4379 -271 -4301 -225
rect -4255 -271 -4177 -225
rect -4131 -271 -4053 -225
rect -4007 -271 -3929 -225
rect -3883 -271 -3805 -225
rect -3759 -271 -3681 -225
rect -3635 -271 -3557 -225
rect -3511 -271 -3433 -225
rect -3387 -271 -3309 -225
rect -3263 -271 -3185 -225
rect -3139 -271 -3061 -225
rect -3015 -271 -2937 -225
rect -2891 -271 -2813 -225
rect -2767 -271 -2689 -225
rect -2643 -271 -2565 -225
rect -2519 -271 -2441 -225
rect -2395 -271 -2317 -225
rect -2271 -271 -2193 -225
rect -2147 -271 -2069 -225
rect -2023 -271 -1945 -225
rect -1899 -271 -1821 -225
rect -1775 -271 -1697 -225
rect -1651 -271 -1573 -225
rect -1527 -271 -1449 -225
rect -1403 -271 -1325 -225
rect -1279 -271 -1201 -225
rect -1155 -271 -1077 -225
rect -1031 -271 -953 -225
rect -907 -271 -829 -225
rect -783 -271 -705 -225
rect -659 -271 -581 -225
rect -535 -271 -457 -225
rect -411 -271 -333 -225
rect -287 -271 -209 -225
rect -163 -271 -85 -225
rect -39 -271 39 -225
rect 85 -271 163 -225
rect 209 -271 287 -225
rect 333 -271 411 -225
rect 457 -271 535 -225
rect 581 -271 659 -225
rect 705 -271 783 -225
rect 829 -271 907 -225
rect 953 -271 1031 -225
rect 1077 -271 1155 -225
rect 1201 -271 1279 -225
rect 1325 -271 1403 -225
rect 1449 -271 1527 -225
rect 1573 -271 1651 -225
rect 1697 -271 1775 -225
rect 1821 -271 1899 -225
rect 1945 -271 2023 -225
rect 2069 -271 2147 -225
rect 2193 -271 2271 -225
rect 2317 -271 2395 -225
rect 2441 -271 2519 -225
rect 2565 -271 2643 -225
rect 2689 -271 2767 -225
rect 2813 -271 2891 -225
rect 2937 -271 3015 -225
rect 3061 -271 3139 -225
rect 3185 -271 3263 -225
rect 3309 -271 3387 -225
rect 3433 -271 3511 -225
rect 3557 -271 3635 -225
rect 3681 -271 3759 -225
rect 3805 -271 3883 -225
rect 3929 -271 4007 -225
rect 4053 -271 4131 -225
rect 4177 -271 4255 -225
rect 4301 -271 4379 -225
rect 4425 -271 4503 -225
rect 4549 -271 4627 -225
rect 4673 -271 4751 -225
rect 4797 -271 4875 -225
rect 4921 -271 4999 -225
rect 5045 -271 5123 -225
rect 5169 -271 5247 -225
rect 5293 -271 5371 -225
rect 5417 -271 5495 -225
rect 5541 -271 5619 -225
rect 5665 -271 5743 -225
rect 5789 -271 5867 -225
rect 5913 -271 5991 -225
rect 6037 -271 6115 -225
rect 6161 -271 6239 -225
rect 6285 -271 6363 -225
rect 6409 -271 6487 -225
rect 6533 -271 6611 -225
rect 6657 -271 6735 -225
rect 6781 -271 6859 -225
rect 6905 -271 6983 -225
rect 7029 -271 7107 -225
rect 7153 -271 7231 -225
rect 7277 -271 7355 -225
rect 7401 -271 7479 -225
rect 7525 -271 7603 -225
rect 7649 -271 7727 -225
rect 7773 -271 7851 -225
rect 7897 -271 7975 -225
rect 8021 -271 8099 -225
rect 8145 -271 8223 -225
rect 8269 -271 8347 -225
rect 8393 -271 8471 -225
rect 8517 -271 8595 -225
rect 8641 -271 8719 -225
rect 8765 -271 8843 -225
rect 8889 -271 8967 -225
rect 9013 -271 9091 -225
rect 9137 -271 9215 -225
rect 9261 -271 9339 -225
rect 9385 -271 9463 -225
rect 9509 -271 9587 -225
rect 9633 -271 9711 -225
rect 9757 -271 9835 -225
rect 9881 -271 9959 -225
rect 10005 -271 10083 -225
rect 10129 -271 10207 -225
rect 10253 -271 10331 -225
rect 10377 -271 10455 -225
rect 10501 -271 10579 -225
rect 10625 -271 10703 -225
rect 10749 -271 10827 -225
rect 10873 -271 10951 -225
rect 10997 -271 11075 -225
rect 11121 -271 11199 -225
rect 11245 -271 11323 -225
rect 11369 -271 11447 -225
rect 11493 -271 11571 -225
rect 11617 -271 11695 -225
rect 11741 -271 11819 -225
rect 11865 -271 11943 -225
rect 11989 -271 12067 -225
rect 12113 -271 12191 -225
rect 12237 -271 12315 -225
rect 12361 -271 12439 -225
rect 12485 -271 12563 -225
rect 12609 -271 12687 -225
rect 12733 -271 12811 -225
rect 12857 -271 12935 -225
rect 12981 -271 13059 -225
rect 13105 -271 13183 -225
rect 13229 -271 13307 -225
rect 13353 -271 13431 -225
rect 13477 -271 13555 -225
rect 13601 -271 13679 -225
rect 13725 -271 13803 -225
rect 13849 -271 13927 -225
rect 13973 -271 14051 -225
rect 14097 -271 14175 -225
rect 14221 -271 14299 -225
rect 14345 -271 14423 -225
rect 14469 -271 14547 -225
rect 14593 -271 14671 -225
rect 14717 -271 14795 -225
rect 14841 -271 14919 -225
rect 14965 -271 15043 -225
rect 15089 -271 15167 -225
rect 15213 -271 15291 -225
rect 15337 -271 15415 -225
rect 15461 -271 15539 -225
rect 15585 -271 15663 -225
rect 15709 -271 15787 -225
rect 15833 -271 15911 -225
rect 15957 -271 16035 -225
rect 16081 -271 16159 -225
rect 16205 -271 16283 -225
rect 16329 -271 16407 -225
rect 16453 -271 16531 -225
rect 16577 -271 16655 -225
rect 16701 -271 16779 -225
rect 16825 -271 16903 -225
rect 16949 -271 17027 -225
rect 17073 -271 17151 -225
rect 17197 -271 17275 -225
rect 17321 -271 17399 -225
rect 17445 -271 17523 -225
rect 17569 -271 17647 -225
rect 17693 -271 17771 -225
rect 17817 -271 17895 -225
rect 17941 -271 18019 -225
rect 18065 -271 18143 -225
rect 18189 -271 18267 -225
rect 18313 -271 18335 -225
rect -18335 -349 18335 -271
rect -18335 -395 -18313 -349
rect -18267 -395 -18189 -349
rect -18143 -395 -18065 -349
rect -18019 -395 -17941 -349
rect -17895 -395 -17817 -349
rect -17771 -395 -17693 -349
rect -17647 -395 -17569 -349
rect -17523 -395 -17445 -349
rect -17399 -395 -17321 -349
rect -17275 -395 -17197 -349
rect -17151 -395 -17073 -349
rect -17027 -395 -16949 -349
rect -16903 -395 -16825 -349
rect -16779 -395 -16701 -349
rect -16655 -395 -16577 -349
rect -16531 -395 -16453 -349
rect -16407 -395 -16329 -349
rect -16283 -395 -16205 -349
rect -16159 -395 -16081 -349
rect -16035 -395 -15957 -349
rect -15911 -395 -15833 -349
rect -15787 -395 -15709 -349
rect -15663 -395 -15585 -349
rect -15539 -395 -15461 -349
rect -15415 -395 -15337 -349
rect -15291 -395 -15213 -349
rect -15167 -395 -15089 -349
rect -15043 -395 -14965 -349
rect -14919 -395 -14841 -349
rect -14795 -395 -14717 -349
rect -14671 -395 -14593 -349
rect -14547 -395 -14469 -349
rect -14423 -395 -14345 -349
rect -14299 -395 -14221 -349
rect -14175 -395 -14097 -349
rect -14051 -395 -13973 -349
rect -13927 -395 -13849 -349
rect -13803 -395 -13725 -349
rect -13679 -395 -13601 -349
rect -13555 -395 -13477 -349
rect -13431 -395 -13353 -349
rect -13307 -395 -13229 -349
rect -13183 -395 -13105 -349
rect -13059 -395 -12981 -349
rect -12935 -395 -12857 -349
rect -12811 -395 -12733 -349
rect -12687 -395 -12609 -349
rect -12563 -395 -12485 -349
rect -12439 -395 -12361 -349
rect -12315 -395 -12237 -349
rect -12191 -395 -12113 -349
rect -12067 -395 -11989 -349
rect -11943 -395 -11865 -349
rect -11819 -395 -11741 -349
rect -11695 -395 -11617 -349
rect -11571 -395 -11493 -349
rect -11447 -395 -11369 -349
rect -11323 -395 -11245 -349
rect -11199 -395 -11121 -349
rect -11075 -395 -10997 -349
rect -10951 -395 -10873 -349
rect -10827 -395 -10749 -349
rect -10703 -395 -10625 -349
rect -10579 -395 -10501 -349
rect -10455 -395 -10377 -349
rect -10331 -395 -10253 -349
rect -10207 -395 -10129 -349
rect -10083 -395 -10005 -349
rect -9959 -395 -9881 -349
rect -9835 -395 -9757 -349
rect -9711 -395 -9633 -349
rect -9587 -395 -9509 -349
rect -9463 -395 -9385 -349
rect -9339 -395 -9261 -349
rect -9215 -395 -9137 -349
rect -9091 -395 -9013 -349
rect -8967 -395 -8889 -349
rect -8843 -395 -8765 -349
rect -8719 -395 -8641 -349
rect -8595 -395 -8517 -349
rect -8471 -395 -8393 -349
rect -8347 -395 -8269 -349
rect -8223 -395 -8145 -349
rect -8099 -395 -8021 -349
rect -7975 -395 -7897 -349
rect -7851 -395 -7773 -349
rect -7727 -395 -7649 -349
rect -7603 -395 -7525 -349
rect -7479 -395 -7401 -349
rect -7355 -395 -7277 -349
rect -7231 -395 -7153 -349
rect -7107 -395 -7029 -349
rect -6983 -395 -6905 -349
rect -6859 -395 -6781 -349
rect -6735 -395 -6657 -349
rect -6611 -395 -6533 -349
rect -6487 -395 -6409 -349
rect -6363 -395 -6285 -349
rect -6239 -395 -6161 -349
rect -6115 -395 -6037 -349
rect -5991 -395 -5913 -349
rect -5867 -395 -5789 -349
rect -5743 -395 -5665 -349
rect -5619 -395 -5541 -349
rect -5495 -395 -5417 -349
rect -5371 -395 -5293 -349
rect -5247 -395 -5169 -349
rect -5123 -395 -5045 -349
rect -4999 -395 -4921 -349
rect -4875 -395 -4797 -349
rect -4751 -395 -4673 -349
rect -4627 -395 -4549 -349
rect -4503 -395 -4425 -349
rect -4379 -395 -4301 -349
rect -4255 -395 -4177 -349
rect -4131 -395 -4053 -349
rect -4007 -395 -3929 -349
rect -3883 -395 -3805 -349
rect -3759 -395 -3681 -349
rect -3635 -395 -3557 -349
rect -3511 -395 -3433 -349
rect -3387 -395 -3309 -349
rect -3263 -395 -3185 -349
rect -3139 -395 -3061 -349
rect -3015 -395 -2937 -349
rect -2891 -395 -2813 -349
rect -2767 -395 -2689 -349
rect -2643 -395 -2565 -349
rect -2519 -395 -2441 -349
rect -2395 -395 -2317 -349
rect -2271 -395 -2193 -349
rect -2147 -395 -2069 -349
rect -2023 -395 -1945 -349
rect -1899 -395 -1821 -349
rect -1775 -395 -1697 -349
rect -1651 -395 -1573 -349
rect -1527 -395 -1449 -349
rect -1403 -395 -1325 -349
rect -1279 -395 -1201 -349
rect -1155 -395 -1077 -349
rect -1031 -395 -953 -349
rect -907 -395 -829 -349
rect -783 -395 -705 -349
rect -659 -395 -581 -349
rect -535 -395 -457 -349
rect -411 -395 -333 -349
rect -287 -395 -209 -349
rect -163 -395 -85 -349
rect -39 -395 39 -349
rect 85 -395 163 -349
rect 209 -395 287 -349
rect 333 -395 411 -349
rect 457 -395 535 -349
rect 581 -395 659 -349
rect 705 -395 783 -349
rect 829 -395 907 -349
rect 953 -395 1031 -349
rect 1077 -395 1155 -349
rect 1201 -395 1279 -349
rect 1325 -395 1403 -349
rect 1449 -395 1527 -349
rect 1573 -395 1651 -349
rect 1697 -395 1775 -349
rect 1821 -395 1899 -349
rect 1945 -395 2023 -349
rect 2069 -395 2147 -349
rect 2193 -395 2271 -349
rect 2317 -395 2395 -349
rect 2441 -395 2519 -349
rect 2565 -395 2643 -349
rect 2689 -395 2767 -349
rect 2813 -395 2891 -349
rect 2937 -395 3015 -349
rect 3061 -395 3139 -349
rect 3185 -395 3263 -349
rect 3309 -395 3387 -349
rect 3433 -395 3511 -349
rect 3557 -395 3635 -349
rect 3681 -395 3759 -349
rect 3805 -395 3883 -349
rect 3929 -395 4007 -349
rect 4053 -395 4131 -349
rect 4177 -395 4255 -349
rect 4301 -395 4379 -349
rect 4425 -395 4503 -349
rect 4549 -395 4627 -349
rect 4673 -395 4751 -349
rect 4797 -395 4875 -349
rect 4921 -395 4999 -349
rect 5045 -395 5123 -349
rect 5169 -395 5247 -349
rect 5293 -395 5371 -349
rect 5417 -395 5495 -349
rect 5541 -395 5619 -349
rect 5665 -395 5743 -349
rect 5789 -395 5867 -349
rect 5913 -395 5991 -349
rect 6037 -395 6115 -349
rect 6161 -395 6239 -349
rect 6285 -395 6363 -349
rect 6409 -395 6487 -349
rect 6533 -395 6611 -349
rect 6657 -395 6735 -349
rect 6781 -395 6859 -349
rect 6905 -395 6983 -349
rect 7029 -395 7107 -349
rect 7153 -395 7231 -349
rect 7277 -395 7355 -349
rect 7401 -395 7479 -349
rect 7525 -395 7603 -349
rect 7649 -395 7727 -349
rect 7773 -395 7851 -349
rect 7897 -395 7975 -349
rect 8021 -395 8099 -349
rect 8145 -395 8223 -349
rect 8269 -395 8347 -349
rect 8393 -395 8471 -349
rect 8517 -395 8595 -349
rect 8641 -395 8719 -349
rect 8765 -395 8843 -349
rect 8889 -395 8967 -349
rect 9013 -395 9091 -349
rect 9137 -395 9215 -349
rect 9261 -395 9339 -349
rect 9385 -395 9463 -349
rect 9509 -395 9587 -349
rect 9633 -395 9711 -349
rect 9757 -395 9835 -349
rect 9881 -395 9959 -349
rect 10005 -395 10083 -349
rect 10129 -395 10207 -349
rect 10253 -395 10331 -349
rect 10377 -395 10455 -349
rect 10501 -395 10579 -349
rect 10625 -395 10703 -349
rect 10749 -395 10827 -349
rect 10873 -395 10951 -349
rect 10997 -395 11075 -349
rect 11121 -395 11199 -349
rect 11245 -395 11323 -349
rect 11369 -395 11447 -349
rect 11493 -395 11571 -349
rect 11617 -395 11695 -349
rect 11741 -395 11819 -349
rect 11865 -395 11943 -349
rect 11989 -395 12067 -349
rect 12113 -395 12191 -349
rect 12237 -395 12315 -349
rect 12361 -395 12439 -349
rect 12485 -395 12563 -349
rect 12609 -395 12687 -349
rect 12733 -395 12811 -349
rect 12857 -395 12935 -349
rect 12981 -395 13059 -349
rect 13105 -395 13183 -349
rect 13229 -395 13307 -349
rect 13353 -395 13431 -349
rect 13477 -395 13555 -349
rect 13601 -395 13679 -349
rect 13725 -395 13803 -349
rect 13849 -395 13927 -349
rect 13973 -395 14051 -349
rect 14097 -395 14175 -349
rect 14221 -395 14299 -349
rect 14345 -395 14423 -349
rect 14469 -395 14547 -349
rect 14593 -395 14671 -349
rect 14717 -395 14795 -349
rect 14841 -395 14919 -349
rect 14965 -395 15043 -349
rect 15089 -395 15167 -349
rect 15213 -395 15291 -349
rect 15337 -395 15415 -349
rect 15461 -395 15539 -349
rect 15585 -395 15663 -349
rect 15709 -395 15787 -349
rect 15833 -395 15911 -349
rect 15957 -395 16035 -349
rect 16081 -395 16159 -349
rect 16205 -395 16283 -349
rect 16329 -395 16407 -349
rect 16453 -395 16531 -349
rect 16577 -395 16655 -349
rect 16701 -395 16779 -349
rect 16825 -395 16903 -349
rect 16949 -395 17027 -349
rect 17073 -395 17151 -349
rect 17197 -395 17275 -349
rect 17321 -395 17399 -349
rect 17445 -395 17523 -349
rect 17569 -395 17647 -349
rect 17693 -395 17771 -349
rect 17817 -395 17895 -349
rect 17941 -395 18019 -349
rect 18065 -395 18143 -349
rect 18189 -395 18267 -349
rect 18313 -395 18335 -349
rect -18335 -473 18335 -395
rect -18335 -519 -18313 -473
rect -18267 -519 -18189 -473
rect -18143 -519 -18065 -473
rect -18019 -519 -17941 -473
rect -17895 -519 -17817 -473
rect -17771 -519 -17693 -473
rect -17647 -519 -17569 -473
rect -17523 -519 -17445 -473
rect -17399 -519 -17321 -473
rect -17275 -519 -17197 -473
rect -17151 -519 -17073 -473
rect -17027 -519 -16949 -473
rect -16903 -519 -16825 -473
rect -16779 -519 -16701 -473
rect -16655 -519 -16577 -473
rect -16531 -519 -16453 -473
rect -16407 -519 -16329 -473
rect -16283 -519 -16205 -473
rect -16159 -519 -16081 -473
rect -16035 -519 -15957 -473
rect -15911 -519 -15833 -473
rect -15787 -519 -15709 -473
rect -15663 -519 -15585 -473
rect -15539 -519 -15461 -473
rect -15415 -519 -15337 -473
rect -15291 -519 -15213 -473
rect -15167 -519 -15089 -473
rect -15043 -519 -14965 -473
rect -14919 -519 -14841 -473
rect -14795 -519 -14717 -473
rect -14671 -519 -14593 -473
rect -14547 -519 -14469 -473
rect -14423 -519 -14345 -473
rect -14299 -519 -14221 -473
rect -14175 -519 -14097 -473
rect -14051 -519 -13973 -473
rect -13927 -519 -13849 -473
rect -13803 -519 -13725 -473
rect -13679 -519 -13601 -473
rect -13555 -519 -13477 -473
rect -13431 -519 -13353 -473
rect -13307 -519 -13229 -473
rect -13183 -519 -13105 -473
rect -13059 -519 -12981 -473
rect -12935 -519 -12857 -473
rect -12811 -519 -12733 -473
rect -12687 -519 -12609 -473
rect -12563 -519 -12485 -473
rect -12439 -519 -12361 -473
rect -12315 -519 -12237 -473
rect -12191 -519 -12113 -473
rect -12067 -519 -11989 -473
rect -11943 -519 -11865 -473
rect -11819 -519 -11741 -473
rect -11695 -519 -11617 -473
rect -11571 -519 -11493 -473
rect -11447 -519 -11369 -473
rect -11323 -519 -11245 -473
rect -11199 -519 -11121 -473
rect -11075 -519 -10997 -473
rect -10951 -519 -10873 -473
rect -10827 -519 -10749 -473
rect -10703 -519 -10625 -473
rect -10579 -519 -10501 -473
rect -10455 -519 -10377 -473
rect -10331 -519 -10253 -473
rect -10207 -519 -10129 -473
rect -10083 -519 -10005 -473
rect -9959 -519 -9881 -473
rect -9835 -519 -9757 -473
rect -9711 -519 -9633 -473
rect -9587 -519 -9509 -473
rect -9463 -519 -9385 -473
rect -9339 -519 -9261 -473
rect -9215 -519 -9137 -473
rect -9091 -519 -9013 -473
rect -8967 -519 -8889 -473
rect -8843 -519 -8765 -473
rect -8719 -519 -8641 -473
rect -8595 -519 -8517 -473
rect -8471 -519 -8393 -473
rect -8347 -519 -8269 -473
rect -8223 -519 -8145 -473
rect -8099 -519 -8021 -473
rect -7975 -519 -7897 -473
rect -7851 -519 -7773 -473
rect -7727 -519 -7649 -473
rect -7603 -519 -7525 -473
rect -7479 -519 -7401 -473
rect -7355 -519 -7277 -473
rect -7231 -519 -7153 -473
rect -7107 -519 -7029 -473
rect -6983 -519 -6905 -473
rect -6859 -519 -6781 -473
rect -6735 -519 -6657 -473
rect -6611 -519 -6533 -473
rect -6487 -519 -6409 -473
rect -6363 -519 -6285 -473
rect -6239 -519 -6161 -473
rect -6115 -519 -6037 -473
rect -5991 -519 -5913 -473
rect -5867 -519 -5789 -473
rect -5743 -519 -5665 -473
rect -5619 -519 -5541 -473
rect -5495 -519 -5417 -473
rect -5371 -519 -5293 -473
rect -5247 -519 -5169 -473
rect -5123 -519 -5045 -473
rect -4999 -519 -4921 -473
rect -4875 -519 -4797 -473
rect -4751 -519 -4673 -473
rect -4627 -519 -4549 -473
rect -4503 -519 -4425 -473
rect -4379 -519 -4301 -473
rect -4255 -519 -4177 -473
rect -4131 -519 -4053 -473
rect -4007 -519 -3929 -473
rect -3883 -519 -3805 -473
rect -3759 -519 -3681 -473
rect -3635 -519 -3557 -473
rect -3511 -519 -3433 -473
rect -3387 -519 -3309 -473
rect -3263 -519 -3185 -473
rect -3139 -519 -3061 -473
rect -3015 -519 -2937 -473
rect -2891 -519 -2813 -473
rect -2767 -519 -2689 -473
rect -2643 -519 -2565 -473
rect -2519 -519 -2441 -473
rect -2395 -519 -2317 -473
rect -2271 -519 -2193 -473
rect -2147 -519 -2069 -473
rect -2023 -519 -1945 -473
rect -1899 -519 -1821 -473
rect -1775 -519 -1697 -473
rect -1651 -519 -1573 -473
rect -1527 -519 -1449 -473
rect -1403 -519 -1325 -473
rect -1279 -519 -1201 -473
rect -1155 -519 -1077 -473
rect -1031 -519 -953 -473
rect -907 -519 -829 -473
rect -783 -519 -705 -473
rect -659 -519 -581 -473
rect -535 -519 -457 -473
rect -411 -519 -333 -473
rect -287 -519 -209 -473
rect -163 -519 -85 -473
rect -39 -519 39 -473
rect 85 -519 163 -473
rect 209 -519 287 -473
rect 333 -519 411 -473
rect 457 -519 535 -473
rect 581 -519 659 -473
rect 705 -519 783 -473
rect 829 -519 907 -473
rect 953 -519 1031 -473
rect 1077 -519 1155 -473
rect 1201 -519 1279 -473
rect 1325 -519 1403 -473
rect 1449 -519 1527 -473
rect 1573 -519 1651 -473
rect 1697 -519 1775 -473
rect 1821 -519 1899 -473
rect 1945 -519 2023 -473
rect 2069 -519 2147 -473
rect 2193 -519 2271 -473
rect 2317 -519 2395 -473
rect 2441 -519 2519 -473
rect 2565 -519 2643 -473
rect 2689 -519 2767 -473
rect 2813 -519 2891 -473
rect 2937 -519 3015 -473
rect 3061 -519 3139 -473
rect 3185 -519 3263 -473
rect 3309 -519 3387 -473
rect 3433 -519 3511 -473
rect 3557 -519 3635 -473
rect 3681 -519 3759 -473
rect 3805 -519 3883 -473
rect 3929 -519 4007 -473
rect 4053 -519 4131 -473
rect 4177 -519 4255 -473
rect 4301 -519 4379 -473
rect 4425 -519 4503 -473
rect 4549 -519 4627 -473
rect 4673 -519 4751 -473
rect 4797 -519 4875 -473
rect 4921 -519 4999 -473
rect 5045 -519 5123 -473
rect 5169 -519 5247 -473
rect 5293 -519 5371 -473
rect 5417 -519 5495 -473
rect 5541 -519 5619 -473
rect 5665 -519 5743 -473
rect 5789 -519 5867 -473
rect 5913 -519 5991 -473
rect 6037 -519 6115 -473
rect 6161 -519 6239 -473
rect 6285 -519 6363 -473
rect 6409 -519 6487 -473
rect 6533 -519 6611 -473
rect 6657 -519 6735 -473
rect 6781 -519 6859 -473
rect 6905 -519 6983 -473
rect 7029 -519 7107 -473
rect 7153 -519 7231 -473
rect 7277 -519 7355 -473
rect 7401 -519 7479 -473
rect 7525 -519 7603 -473
rect 7649 -519 7727 -473
rect 7773 -519 7851 -473
rect 7897 -519 7975 -473
rect 8021 -519 8099 -473
rect 8145 -519 8223 -473
rect 8269 -519 8347 -473
rect 8393 -519 8471 -473
rect 8517 -519 8595 -473
rect 8641 -519 8719 -473
rect 8765 -519 8843 -473
rect 8889 -519 8967 -473
rect 9013 -519 9091 -473
rect 9137 -519 9215 -473
rect 9261 -519 9339 -473
rect 9385 -519 9463 -473
rect 9509 -519 9587 -473
rect 9633 -519 9711 -473
rect 9757 -519 9835 -473
rect 9881 -519 9959 -473
rect 10005 -519 10083 -473
rect 10129 -519 10207 -473
rect 10253 -519 10331 -473
rect 10377 -519 10455 -473
rect 10501 -519 10579 -473
rect 10625 -519 10703 -473
rect 10749 -519 10827 -473
rect 10873 -519 10951 -473
rect 10997 -519 11075 -473
rect 11121 -519 11199 -473
rect 11245 -519 11323 -473
rect 11369 -519 11447 -473
rect 11493 -519 11571 -473
rect 11617 -519 11695 -473
rect 11741 -519 11819 -473
rect 11865 -519 11943 -473
rect 11989 -519 12067 -473
rect 12113 -519 12191 -473
rect 12237 -519 12315 -473
rect 12361 -519 12439 -473
rect 12485 -519 12563 -473
rect 12609 -519 12687 -473
rect 12733 -519 12811 -473
rect 12857 -519 12935 -473
rect 12981 -519 13059 -473
rect 13105 -519 13183 -473
rect 13229 -519 13307 -473
rect 13353 -519 13431 -473
rect 13477 -519 13555 -473
rect 13601 -519 13679 -473
rect 13725 -519 13803 -473
rect 13849 -519 13927 -473
rect 13973 -519 14051 -473
rect 14097 -519 14175 -473
rect 14221 -519 14299 -473
rect 14345 -519 14423 -473
rect 14469 -519 14547 -473
rect 14593 -519 14671 -473
rect 14717 -519 14795 -473
rect 14841 -519 14919 -473
rect 14965 -519 15043 -473
rect 15089 -519 15167 -473
rect 15213 -519 15291 -473
rect 15337 -519 15415 -473
rect 15461 -519 15539 -473
rect 15585 -519 15663 -473
rect 15709 -519 15787 -473
rect 15833 -519 15911 -473
rect 15957 -519 16035 -473
rect 16081 -519 16159 -473
rect 16205 -519 16283 -473
rect 16329 -519 16407 -473
rect 16453 -519 16531 -473
rect 16577 -519 16655 -473
rect 16701 -519 16779 -473
rect 16825 -519 16903 -473
rect 16949 -519 17027 -473
rect 17073 -519 17151 -473
rect 17197 -519 17275 -473
rect 17321 -519 17399 -473
rect 17445 -519 17523 -473
rect 17569 -519 17647 -473
rect 17693 -519 17771 -473
rect 17817 -519 17895 -473
rect 17941 -519 18019 -473
rect 18065 -519 18143 -473
rect 18189 -519 18267 -473
rect 18313 -519 18335 -473
rect -18335 -597 18335 -519
rect -18335 -643 -18313 -597
rect -18267 -643 -18189 -597
rect -18143 -643 -18065 -597
rect -18019 -643 -17941 -597
rect -17895 -643 -17817 -597
rect -17771 -643 -17693 -597
rect -17647 -643 -17569 -597
rect -17523 -643 -17445 -597
rect -17399 -643 -17321 -597
rect -17275 -643 -17197 -597
rect -17151 -643 -17073 -597
rect -17027 -643 -16949 -597
rect -16903 -643 -16825 -597
rect -16779 -643 -16701 -597
rect -16655 -643 -16577 -597
rect -16531 -643 -16453 -597
rect -16407 -643 -16329 -597
rect -16283 -643 -16205 -597
rect -16159 -643 -16081 -597
rect -16035 -643 -15957 -597
rect -15911 -643 -15833 -597
rect -15787 -643 -15709 -597
rect -15663 -643 -15585 -597
rect -15539 -643 -15461 -597
rect -15415 -643 -15337 -597
rect -15291 -643 -15213 -597
rect -15167 -643 -15089 -597
rect -15043 -643 -14965 -597
rect -14919 -643 -14841 -597
rect -14795 -643 -14717 -597
rect -14671 -643 -14593 -597
rect -14547 -643 -14469 -597
rect -14423 -643 -14345 -597
rect -14299 -643 -14221 -597
rect -14175 -643 -14097 -597
rect -14051 -643 -13973 -597
rect -13927 -643 -13849 -597
rect -13803 -643 -13725 -597
rect -13679 -643 -13601 -597
rect -13555 -643 -13477 -597
rect -13431 -643 -13353 -597
rect -13307 -643 -13229 -597
rect -13183 -643 -13105 -597
rect -13059 -643 -12981 -597
rect -12935 -643 -12857 -597
rect -12811 -643 -12733 -597
rect -12687 -643 -12609 -597
rect -12563 -643 -12485 -597
rect -12439 -643 -12361 -597
rect -12315 -643 -12237 -597
rect -12191 -643 -12113 -597
rect -12067 -643 -11989 -597
rect -11943 -643 -11865 -597
rect -11819 -643 -11741 -597
rect -11695 -643 -11617 -597
rect -11571 -643 -11493 -597
rect -11447 -643 -11369 -597
rect -11323 -643 -11245 -597
rect -11199 -643 -11121 -597
rect -11075 -643 -10997 -597
rect -10951 -643 -10873 -597
rect -10827 -643 -10749 -597
rect -10703 -643 -10625 -597
rect -10579 -643 -10501 -597
rect -10455 -643 -10377 -597
rect -10331 -643 -10253 -597
rect -10207 -643 -10129 -597
rect -10083 -643 -10005 -597
rect -9959 -643 -9881 -597
rect -9835 -643 -9757 -597
rect -9711 -643 -9633 -597
rect -9587 -643 -9509 -597
rect -9463 -643 -9385 -597
rect -9339 -643 -9261 -597
rect -9215 -643 -9137 -597
rect -9091 -643 -9013 -597
rect -8967 -643 -8889 -597
rect -8843 -643 -8765 -597
rect -8719 -643 -8641 -597
rect -8595 -643 -8517 -597
rect -8471 -643 -8393 -597
rect -8347 -643 -8269 -597
rect -8223 -643 -8145 -597
rect -8099 -643 -8021 -597
rect -7975 -643 -7897 -597
rect -7851 -643 -7773 -597
rect -7727 -643 -7649 -597
rect -7603 -643 -7525 -597
rect -7479 -643 -7401 -597
rect -7355 -643 -7277 -597
rect -7231 -643 -7153 -597
rect -7107 -643 -7029 -597
rect -6983 -643 -6905 -597
rect -6859 -643 -6781 -597
rect -6735 -643 -6657 -597
rect -6611 -643 -6533 -597
rect -6487 -643 -6409 -597
rect -6363 -643 -6285 -597
rect -6239 -643 -6161 -597
rect -6115 -643 -6037 -597
rect -5991 -643 -5913 -597
rect -5867 -643 -5789 -597
rect -5743 -643 -5665 -597
rect -5619 -643 -5541 -597
rect -5495 -643 -5417 -597
rect -5371 -643 -5293 -597
rect -5247 -643 -5169 -597
rect -5123 -643 -5045 -597
rect -4999 -643 -4921 -597
rect -4875 -643 -4797 -597
rect -4751 -643 -4673 -597
rect -4627 -643 -4549 -597
rect -4503 -643 -4425 -597
rect -4379 -643 -4301 -597
rect -4255 -643 -4177 -597
rect -4131 -643 -4053 -597
rect -4007 -643 -3929 -597
rect -3883 -643 -3805 -597
rect -3759 -643 -3681 -597
rect -3635 -643 -3557 -597
rect -3511 -643 -3433 -597
rect -3387 -643 -3309 -597
rect -3263 -643 -3185 -597
rect -3139 -643 -3061 -597
rect -3015 -643 -2937 -597
rect -2891 -643 -2813 -597
rect -2767 -643 -2689 -597
rect -2643 -643 -2565 -597
rect -2519 -643 -2441 -597
rect -2395 -643 -2317 -597
rect -2271 -643 -2193 -597
rect -2147 -643 -2069 -597
rect -2023 -643 -1945 -597
rect -1899 -643 -1821 -597
rect -1775 -643 -1697 -597
rect -1651 -643 -1573 -597
rect -1527 -643 -1449 -597
rect -1403 -643 -1325 -597
rect -1279 -643 -1201 -597
rect -1155 -643 -1077 -597
rect -1031 -643 -953 -597
rect -907 -643 -829 -597
rect -783 -643 -705 -597
rect -659 -643 -581 -597
rect -535 -643 -457 -597
rect -411 -643 -333 -597
rect -287 -643 -209 -597
rect -163 -643 -85 -597
rect -39 -643 39 -597
rect 85 -643 163 -597
rect 209 -643 287 -597
rect 333 -643 411 -597
rect 457 -643 535 -597
rect 581 -643 659 -597
rect 705 -643 783 -597
rect 829 -643 907 -597
rect 953 -643 1031 -597
rect 1077 -643 1155 -597
rect 1201 -643 1279 -597
rect 1325 -643 1403 -597
rect 1449 -643 1527 -597
rect 1573 -643 1651 -597
rect 1697 -643 1775 -597
rect 1821 -643 1899 -597
rect 1945 -643 2023 -597
rect 2069 -643 2147 -597
rect 2193 -643 2271 -597
rect 2317 -643 2395 -597
rect 2441 -643 2519 -597
rect 2565 -643 2643 -597
rect 2689 -643 2767 -597
rect 2813 -643 2891 -597
rect 2937 -643 3015 -597
rect 3061 -643 3139 -597
rect 3185 -643 3263 -597
rect 3309 -643 3387 -597
rect 3433 -643 3511 -597
rect 3557 -643 3635 -597
rect 3681 -643 3759 -597
rect 3805 -643 3883 -597
rect 3929 -643 4007 -597
rect 4053 -643 4131 -597
rect 4177 -643 4255 -597
rect 4301 -643 4379 -597
rect 4425 -643 4503 -597
rect 4549 -643 4627 -597
rect 4673 -643 4751 -597
rect 4797 -643 4875 -597
rect 4921 -643 4999 -597
rect 5045 -643 5123 -597
rect 5169 -643 5247 -597
rect 5293 -643 5371 -597
rect 5417 -643 5495 -597
rect 5541 -643 5619 -597
rect 5665 -643 5743 -597
rect 5789 -643 5867 -597
rect 5913 -643 5991 -597
rect 6037 -643 6115 -597
rect 6161 -643 6239 -597
rect 6285 -643 6363 -597
rect 6409 -643 6487 -597
rect 6533 -643 6611 -597
rect 6657 -643 6735 -597
rect 6781 -643 6859 -597
rect 6905 -643 6983 -597
rect 7029 -643 7107 -597
rect 7153 -643 7231 -597
rect 7277 -643 7355 -597
rect 7401 -643 7479 -597
rect 7525 -643 7603 -597
rect 7649 -643 7727 -597
rect 7773 -643 7851 -597
rect 7897 -643 7975 -597
rect 8021 -643 8099 -597
rect 8145 -643 8223 -597
rect 8269 -643 8347 -597
rect 8393 -643 8471 -597
rect 8517 -643 8595 -597
rect 8641 -643 8719 -597
rect 8765 -643 8843 -597
rect 8889 -643 8967 -597
rect 9013 -643 9091 -597
rect 9137 -643 9215 -597
rect 9261 -643 9339 -597
rect 9385 -643 9463 -597
rect 9509 -643 9587 -597
rect 9633 -643 9711 -597
rect 9757 -643 9835 -597
rect 9881 -643 9959 -597
rect 10005 -643 10083 -597
rect 10129 -643 10207 -597
rect 10253 -643 10331 -597
rect 10377 -643 10455 -597
rect 10501 -643 10579 -597
rect 10625 -643 10703 -597
rect 10749 -643 10827 -597
rect 10873 -643 10951 -597
rect 10997 -643 11075 -597
rect 11121 -643 11199 -597
rect 11245 -643 11323 -597
rect 11369 -643 11447 -597
rect 11493 -643 11571 -597
rect 11617 -643 11695 -597
rect 11741 -643 11819 -597
rect 11865 -643 11943 -597
rect 11989 -643 12067 -597
rect 12113 -643 12191 -597
rect 12237 -643 12315 -597
rect 12361 -643 12439 -597
rect 12485 -643 12563 -597
rect 12609 -643 12687 -597
rect 12733 -643 12811 -597
rect 12857 -643 12935 -597
rect 12981 -643 13059 -597
rect 13105 -643 13183 -597
rect 13229 -643 13307 -597
rect 13353 -643 13431 -597
rect 13477 -643 13555 -597
rect 13601 -643 13679 -597
rect 13725 -643 13803 -597
rect 13849 -643 13927 -597
rect 13973 -643 14051 -597
rect 14097 -643 14175 -597
rect 14221 -643 14299 -597
rect 14345 -643 14423 -597
rect 14469 -643 14547 -597
rect 14593 -643 14671 -597
rect 14717 -643 14795 -597
rect 14841 -643 14919 -597
rect 14965 -643 15043 -597
rect 15089 -643 15167 -597
rect 15213 -643 15291 -597
rect 15337 -643 15415 -597
rect 15461 -643 15539 -597
rect 15585 -643 15663 -597
rect 15709 -643 15787 -597
rect 15833 -643 15911 -597
rect 15957 -643 16035 -597
rect 16081 -643 16159 -597
rect 16205 -643 16283 -597
rect 16329 -643 16407 -597
rect 16453 -643 16531 -597
rect 16577 -643 16655 -597
rect 16701 -643 16779 -597
rect 16825 -643 16903 -597
rect 16949 -643 17027 -597
rect 17073 -643 17151 -597
rect 17197 -643 17275 -597
rect 17321 -643 17399 -597
rect 17445 -643 17523 -597
rect 17569 -643 17647 -597
rect 17693 -643 17771 -597
rect 17817 -643 17895 -597
rect 17941 -643 18019 -597
rect 18065 -643 18143 -597
rect 18189 -643 18267 -597
rect 18313 -643 18335 -597
rect -18335 -665 18335 -643
<< psubdiffcont >>
rect -18313 597 -18267 643
rect -18189 597 -18143 643
rect -18065 597 -18019 643
rect -17941 597 -17895 643
rect -17817 597 -17771 643
rect -17693 597 -17647 643
rect -17569 597 -17523 643
rect -17445 597 -17399 643
rect -17321 597 -17275 643
rect -17197 597 -17151 643
rect -17073 597 -17027 643
rect -16949 597 -16903 643
rect -16825 597 -16779 643
rect -16701 597 -16655 643
rect -16577 597 -16531 643
rect -16453 597 -16407 643
rect -16329 597 -16283 643
rect -16205 597 -16159 643
rect -16081 597 -16035 643
rect -15957 597 -15911 643
rect -15833 597 -15787 643
rect -15709 597 -15663 643
rect -15585 597 -15539 643
rect -15461 597 -15415 643
rect -15337 597 -15291 643
rect -15213 597 -15167 643
rect -15089 597 -15043 643
rect -14965 597 -14919 643
rect -14841 597 -14795 643
rect -14717 597 -14671 643
rect -14593 597 -14547 643
rect -14469 597 -14423 643
rect -14345 597 -14299 643
rect -14221 597 -14175 643
rect -14097 597 -14051 643
rect -13973 597 -13927 643
rect -13849 597 -13803 643
rect -13725 597 -13679 643
rect -13601 597 -13555 643
rect -13477 597 -13431 643
rect -13353 597 -13307 643
rect -13229 597 -13183 643
rect -13105 597 -13059 643
rect -12981 597 -12935 643
rect -12857 597 -12811 643
rect -12733 597 -12687 643
rect -12609 597 -12563 643
rect -12485 597 -12439 643
rect -12361 597 -12315 643
rect -12237 597 -12191 643
rect -12113 597 -12067 643
rect -11989 597 -11943 643
rect -11865 597 -11819 643
rect -11741 597 -11695 643
rect -11617 597 -11571 643
rect -11493 597 -11447 643
rect -11369 597 -11323 643
rect -11245 597 -11199 643
rect -11121 597 -11075 643
rect -10997 597 -10951 643
rect -10873 597 -10827 643
rect -10749 597 -10703 643
rect -10625 597 -10579 643
rect -10501 597 -10455 643
rect -10377 597 -10331 643
rect -10253 597 -10207 643
rect -10129 597 -10083 643
rect -10005 597 -9959 643
rect -9881 597 -9835 643
rect -9757 597 -9711 643
rect -9633 597 -9587 643
rect -9509 597 -9463 643
rect -9385 597 -9339 643
rect -9261 597 -9215 643
rect -9137 597 -9091 643
rect -9013 597 -8967 643
rect -8889 597 -8843 643
rect -8765 597 -8719 643
rect -8641 597 -8595 643
rect -8517 597 -8471 643
rect -8393 597 -8347 643
rect -8269 597 -8223 643
rect -8145 597 -8099 643
rect -8021 597 -7975 643
rect -7897 597 -7851 643
rect -7773 597 -7727 643
rect -7649 597 -7603 643
rect -7525 597 -7479 643
rect -7401 597 -7355 643
rect -7277 597 -7231 643
rect -7153 597 -7107 643
rect -7029 597 -6983 643
rect -6905 597 -6859 643
rect -6781 597 -6735 643
rect -6657 597 -6611 643
rect -6533 597 -6487 643
rect -6409 597 -6363 643
rect -6285 597 -6239 643
rect -6161 597 -6115 643
rect -6037 597 -5991 643
rect -5913 597 -5867 643
rect -5789 597 -5743 643
rect -5665 597 -5619 643
rect -5541 597 -5495 643
rect -5417 597 -5371 643
rect -5293 597 -5247 643
rect -5169 597 -5123 643
rect -5045 597 -4999 643
rect -4921 597 -4875 643
rect -4797 597 -4751 643
rect -4673 597 -4627 643
rect -4549 597 -4503 643
rect -4425 597 -4379 643
rect -4301 597 -4255 643
rect -4177 597 -4131 643
rect -4053 597 -4007 643
rect -3929 597 -3883 643
rect -3805 597 -3759 643
rect -3681 597 -3635 643
rect -3557 597 -3511 643
rect -3433 597 -3387 643
rect -3309 597 -3263 643
rect -3185 597 -3139 643
rect -3061 597 -3015 643
rect -2937 597 -2891 643
rect -2813 597 -2767 643
rect -2689 597 -2643 643
rect -2565 597 -2519 643
rect -2441 597 -2395 643
rect -2317 597 -2271 643
rect -2193 597 -2147 643
rect -2069 597 -2023 643
rect -1945 597 -1899 643
rect -1821 597 -1775 643
rect -1697 597 -1651 643
rect -1573 597 -1527 643
rect -1449 597 -1403 643
rect -1325 597 -1279 643
rect -1201 597 -1155 643
rect -1077 597 -1031 643
rect -953 597 -907 643
rect -829 597 -783 643
rect -705 597 -659 643
rect -581 597 -535 643
rect -457 597 -411 643
rect -333 597 -287 643
rect -209 597 -163 643
rect -85 597 -39 643
rect 39 597 85 643
rect 163 597 209 643
rect 287 597 333 643
rect 411 597 457 643
rect 535 597 581 643
rect 659 597 705 643
rect 783 597 829 643
rect 907 597 953 643
rect 1031 597 1077 643
rect 1155 597 1201 643
rect 1279 597 1325 643
rect 1403 597 1449 643
rect 1527 597 1573 643
rect 1651 597 1697 643
rect 1775 597 1821 643
rect 1899 597 1945 643
rect 2023 597 2069 643
rect 2147 597 2193 643
rect 2271 597 2317 643
rect 2395 597 2441 643
rect 2519 597 2565 643
rect 2643 597 2689 643
rect 2767 597 2813 643
rect 2891 597 2937 643
rect 3015 597 3061 643
rect 3139 597 3185 643
rect 3263 597 3309 643
rect 3387 597 3433 643
rect 3511 597 3557 643
rect 3635 597 3681 643
rect 3759 597 3805 643
rect 3883 597 3929 643
rect 4007 597 4053 643
rect 4131 597 4177 643
rect 4255 597 4301 643
rect 4379 597 4425 643
rect 4503 597 4549 643
rect 4627 597 4673 643
rect 4751 597 4797 643
rect 4875 597 4921 643
rect 4999 597 5045 643
rect 5123 597 5169 643
rect 5247 597 5293 643
rect 5371 597 5417 643
rect 5495 597 5541 643
rect 5619 597 5665 643
rect 5743 597 5789 643
rect 5867 597 5913 643
rect 5991 597 6037 643
rect 6115 597 6161 643
rect 6239 597 6285 643
rect 6363 597 6409 643
rect 6487 597 6533 643
rect 6611 597 6657 643
rect 6735 597 6781 643
rect 6859 597 6905 643
rect 6983 597 7029 643
rect 7107 597 7153 643
rect 7231 597 7277 643
rect 7355 597 7401 643
rect 7479 597 7525 643
rect 7603 597 7649 643
rect 7727 597 7773 643
rect 7851 597 7897 643
rect 7975 597 8021 643
rect 8099 597 8145 643
rect 8223 597 8269 643
rect 8347 597 8393 643
rect 8471 597 8517 643
rect 8595 597 8641 643
rect 8719 597 8765 643
rect 8843 597 8889 643
rect 8967 597 9013 643
rect 9091 597 9137 643
rect 9215 597 9261 643
rect 9339 597 9385 643
rect 9463 597 9509 643
rect 9587 597 9633 643
rect 9711 597 9757 643
rect 9835 597 9881 643
rect 9959 597 10005 643
rect 10083 597 10129 643
rect 10207 597 10253 643
rect 10331 597 10377 643
rect 10455 597 10501 643
rect 10579 597 10625 643
rect 10703 597 10749 643
rect 10827 597 10873 643
rect 10951 597 10997 643
rect 11075 597 11121 643
rect 11199 597 11245 643
rect 11323 597 11369 643
rect 11447 597 11493 643
rect 11571 597 11617 643
rect 11695 597 11741 643
rect 11819 597 11865 643
rect 11943 597 11989 643
rect 12067 597 12113 643
rect 12191 597 12237 643
rect 12315 597 12361 643
rect 12439 597 12485 643
rect 12563 597 12609 643
rect 12687 597 12733 643
rect 12811 597 12857 643
rect 12935 597 12981 643
rect 13059 597 13105 643
rect 13183 597 13229 643
rect 13307 597 13353 643
rect 13431 597 13477 643
rect 13555 597 13601 643
rect 13679 597 13725 643
rect 13803 597 13849 643
rect 13927 597 13973 643
rect 14051 597 14097 643
rect 14175 597 14221 643
rect 14299 597 14345 643
rect 14423 597 14469 643
rect 14547 597 14593 643
rect 14671 597 14717 643
rect 14795 597 14841 643
rect 14919 597 14965 643
rect 15043 597 15089 643
rect 15167 597 15213 643
rect 15291 597 15337 643
rect 15415 597 15461 643
rect 15539 597 15585 643
rect 15663 597 15709 643
rect 15787 597 15833 643
rect 15911 597 15957 643
rect 16035 597 16081 643
rect 16159 597 16205 643
rect 16283 597 16329 643
rect 16407 597 16453 643
rect 16531 597 16577 643
rect 16655 597 16701 643
rect 16779 597 16825 643
rect 16903 597 16949 643
rect 17027 597 17073 643
rect 17151 597 17197 643
rect 17275 597 17321 643
rect 17399 597 17445 643
rect 17523 597 17569 643
rect 17647 597 17693 643
rect 17771 597 17817 643
rect 17895 597 17941 643
rect 18019 597 18065 643
rect 18143 597 18189 643
rect 18267 597 18313 643
rect -18313 473 -18267 519
rect -18189 473 -18143 519
rect -18065 473 -18019 519
rect -17941 473 -17895 519
rect -17817 473 -17771 519
rect -17693 473 -17647 519
rect -17569 473 -17523 519
rect -17445 473 -17399 519
rect -17321 473 -17275 519
rect -17197 473 -17151 519
rect -17073 473 -17027 519
rect -16949 473 -16903 519
rect -16825 473 -16779 519
rect -16701 473 -16655 519
rect -16577 473 -16531 519
rect -16453 473 -16407 519
rect -16329 473 -16283 519
rect -16205 473 -16159 519
rect -16081 473 -16035 519
rect -15957 473 -15911 519
rect -15833 473 -15787 519
rect -15709 473 -15663 519
rect -15585 473 -15539 519
rect -15461 473 -15415 519
rect -15337 473 -15291 519
rect -15213 473 -15167 519
rect -15089 473 -15043 519
rect -14965 473 -14919 519
rect -14841 473 -14795 519
rect -14717 473 -14671 519
rect -14593 473 -14547 519
rect -14469 473 -14423 519
rect -14345 473 -14299 519
rect -14221 473 -14175 519
rect -14097 473 -14051 519
rect -13973 473 -13927 519
rect -13849 473 -13803 519
rect -13725 473 -13679 519
rect -13601 473 -13555 519
rect -13477 473 -13431 519
rect -13353 473 -13307 519
rect -13229 473 -13183 519
rect -13105 473 -13059 519
rect -12981 473 -12935 519
rect -12857 473 -12811 519
rect -12733 473 -12687 519
rect -12609 473 -12563 519
rect -12485 473 -12439 519
rect -12361 473 -12315 519
rect -12237 473 -12191 519
rect -12113 473 -12067 519
rect -11989 473 -11943 519
rect -11865 473 -11819 519
rect -11741 473 -11695 519
rect -11617 473 -11571 519
rect -11493 473 -11447 519
rect -11369 473 -11323 519
rect -11245 473 -11199 519
rect -11121 473 -11075 519
rect -10997 473 -10951 519
rect -10873 473 -10827 519
rect -10749 473 -10703 519
rect -10625 473 -10579 519
rect -10501 473 -10455 519
rect -10377 473 -10331 519
rect -10253 473 -10207 519
rect -10129 473 -10083 519
rect -10005 473 -9959 519
rect -9881 473 -9835 519
rect -9757 473 -9711 519
rect -9633 473 -9587 519
rect -9509 473 -9463 519
rect -9385 473 -9339 519
rect -9261 473 -9215 519
rect -9137 473 -9091 519
rect -9013 473 -8967 519
rect -8889 473 -8843 519
rect -8765 473 -8719 519
rect -8641 473 -8595 519
rect -8517 473 -8471 519
rect -8393 473 -8347 519
rect -8269 473 -8223 519
rect -8145 473 -8099 519
rect -8021 473 -7975 519
rect -7897 473 -7851 519
rect -7773 473 -7727 519
rect -7649 473 -7603 519
rect -7525 473 -7479 519
rect -7401 473 -7355 519
rect -7277 473 -7231 519
rect -7153 473 -7107 519
rect -7029 473 -6983 519
rect -6905 473 -6859 519
rect -6781 473 -6735 519
rect -6657 473 -6611 519
rect -6533 473 -6487 519
rect -6409 473 -6363 519
rect -6285 473 -6239 519
rect -6161 473 -6115 519
rect -6037 473 -5991 519
rect -5913 473 -5867 519
rect -5789 473 -5743 519
rect -5665 473 -5619 519
rect -5541 473 -5495 519
rect -5417 473 -5371 519
rect -5293 473 -5247 519
rect -5169 473 -5123 519
rect -5045 473 -4999 519
rect -4921 473 -4875 519
rect -4797 473 -4751 519
rect -4673 473 -4627 519
rect -4549 473 -4503 519
rect -4425 473 -4379 519
rect -4301 473 -4255 519
rect -4177 473 -4131 519
rect -4053 473 -4007 519
rect -3929 473 -3883 519
rect -3805 473 -3759 519
rect -3681 473 -3635 519
rect -3557 473 -3511 519
rect -3433 473 -3387 519
rect -3309 473 -3263 519
rect -3185 473 -3139 519
rect -3061 473 -3015 519
rect -2937 473 -2891 519
rect -2813 473 -2767 519
rect -2689 473 -2643 519
rect -2565 473 -2519 519
rect -2441 473 -2395 519
rect -2317 473 -2271 519
rect -2193 473 -2147 519
rect -2069 473 -2023 519
rect -1945 473 -1899 519
rect -1821 473 -1775 519
rect -1697 473 -1651 519
rect -1573 473 -1527 519
rect -1449 473 -1403 519
rect -1325 473 -1279 519
rect -1201 473 -1155 519
rect -1077 473 -1031 519
rect -953 473 -907 519
rect -829 473 -783 519
rect -705 473 -659 519
rect -581 473 -535 519
rect -457 473 -411 519
rect -333 473 -287 519
rect -209 473 -163 519
rect -85 473 -39 519
rect 39 473 85 519
rect 163 473 209 519
rect 287 473 333 519
rect 411 473 457 519
rect 535 473 581 519
rect 659 473 705 519
rect 783 473 829 519
rect 907 473 953 519
rect 1031 473 1077 519
rect 1155 473 1201 519
rect 1279 473 1325 519
rect 1403 473 1449 519
rect 1527 473 1573 519
rect 1651 473 1697 519
rect 1775 473 1821 519
rect 1899 473 1945 519
rect 2023 473 2069 519
rect 2147 473 2193 519
rect 2271 473 2317 519
rect 2395 473 2441 519
rect 2519 473 2565 519
rect 2643 473 2689 519
rect 2767 473 2813 519
rect 2891 473 2937 519
rect 3015 473 3061 519
rect 3139 473 3185 519
rect 3263 473 3309 519
rect 3387 473 3433 519
rect 3511 473 3557 519
rect 3635 473 3681 519
rect 3759 473 3805 519
rect 3883 473 3929 519
rect 4007 473 4053 519
rect 4131 473 4177 519
rect 4255 473 4301 519
rect 4379 473 4425 519
rect 4503 473 4549 519
rect 4627 473 4673 519
rect 4751 473 4797 519
rect 4875 473 4921 519
rect 4999 473 5045 519
rect 5123 473 5169 519
rect 5247 473 5293 519
rect 5371 473 5417 519
rect 5495 473 5541 519
rect 5619 473 5665 519
rect 5743 473 5789 519
rect 5867 473 5913 519
rect 5991 473 6037 519
rect 6115 473 6161 519
rect 6239 473 6285 519
rect 6363 473 6409 519
rect 6487 473 6533 519
rect 6611 473 6657 519
rect 6735 473 6781 519
rect 6859 473 6905 519
rect 6983 473 7029 519
rect 7107 473 7153 519
rect 7231 473 7277 519
rect 7355 473 7401 519
rect 7479 473 7525 519
rect 7603 473 7649 519
rect 7727 473 7773 519
rect 7851 473 7897 519
rect 7975 473 8021 519
rect 8099 473 8145 519
rect 8223 473 8269 519
rect 8347 473 8393 519
rect 8471 473 8517 519
rect 8595 473 8641 519
rect 8719 473 8765 519
rect 8843 473 8889 519
rect 8967 473 9013 519
rect 9091 473 9137 519
rect 9215 473 9261 519
rect 9339 473 9385 519
rect 9463 473 9509 519
rect 9587 473 9633 519
rect 9711 473 9757 519
rect 9835 473 9881 519
rect 9959 473 10005 519
rect 10083 473 10129 519
rect 10207 473 10253 519
rect 10331 473 10377 519
rect 10455 473 10501 519
rect 10579 473 10625 519
rect 10703 473 10749 519
rect 10827 473 10873 519
rect 10951 473 10997 519
rect 11075 473 11121 519
rect 11199 473 11245 519
rect 11323 473 11369 519
rect 11447 473 11493 519
rect 11571 473 11617 519
rect 11695 473 11741 519
rect 11819 473 11865 519
rect 11943 473 11989 519
rect 12067 473 12113 519
rect 12191 473 12237 519
rect 12315 473 12361 519
rect 12439 473 12485 519
rect 12563 473 12609 519
rect 12687 473 12733 519
rect 12811 473 12857 519
rect 12935 473 12981 519
rect 13059 473 13105 519
rect 13183 473 13229 519
rect 13307 473 13353 519
rect 13431 473 13477 519
rect 13555 473 13601 519
rect 13679 473 13725 519
rect 13803 473 13849 519
rect 13927 473 13973 519
rect 14051 473 14097 519
rect 14175 473 14221 519
rect 14299 473 14345 519
rect 14423 473 14469 519
rect 14547 473 14593 519
rect 14671 473 14717 519
rect 14795 473 14841 519
rect 14919 473 14965 519
rect 15043 473 15089 519
rect 15167 473 15213 519
rect 15291 473 15337 519
rect 15415 473 15461 519
rect 15539 473 15585 519
rect 15663 473 15709 519
rect 15787 473 15833 519
rect 15911 473 15957 519
rect 16035 473 16081 519
rect 16159 473 16205 519
rect 16283 473 16329 519
rect 16407 473 16453 519
rect 16531 473 16577 519
rect 16655 473 16701 519
rect 16779 473 16825 519
rect 16903 473 16949 519
rect 17027 473 17073 519
rect 17151 473 17197 519
rect 17275 473 17321 519
rect 17399 473 17445 519
rect 17523 473 17569 519
rect 17647 473 17693 519
rect 17771 473 17817 519
rect 17895 473 17941 519
rect 18019 473 18065 519
rect 18143 473 18189 519
rect 18267 473 18313 519
rect -18313 349 -18267 395
rect -18189 349 -18143 395
rect -18065 349 -18019 395
rect -17941 349 -17895 395
rect -17817 349 -17771 395
rect -17693 349 -17647 395
rect -17569 349 -17523 395
rect -17445 349 -17399 395
rect -17321 349 -17275 395
rect -17197 349 -17151 395
rect -17073 349 -17027 395
rect -16949 349 -16903 395
rect -16825 349 -16779 395
rect -16701 349 -16655 395
rect -16577 349 -16531 395
rect -16453 349 -16407 395
rect -16329 349 -16283 395
rect -16205 349 -16159 395
rect -16081 349 -16035 395
rect -15957 349 -15911 395
rect -15833 349 -15787 395
rect -15709 349 -15663 395
rect -15585 349 -15539 395
rect -15461 349 -15415 395
rect -15337 349 -15291 395
rect -15213 349 -15167 395
rect -15089 349 -15043 395
rect -14965 349 -14919 395
rect -14841 349 -14795 395
rect -14717 349 -14671 395
rect -14593 349 -14547 395
rect -14469 349 -14423 395
rect -14345 349 -14299 395
rect -14221 349 -14175 395
rect -14097 349 -14051 395
rect -13973 349 -13927 395
rect -13849 349 -13803 395
rect -13725 349 -13679 395
rect -13601 349 -13555 395
rect -13477 349 -13431 395
rect -13353 349 -13307 395
rect -13229 349 -13183 395
rect -13105 349 -13059 395
rect -12981 349 -12935 395
rect -12857 349 -12811 395
rect -12733 349 -12687 395
rect -12609 349 -12563 395
rect -12485 349 -12439 395
rect -12361 349 -12315 395
rect -12237 349 -12191 395
rect -12113 349 -12067 395
rect -11989 349 -11943 395
rect -11865 349 -11819 395
rect -11741 349 -11695 395
rect -11617 349 -11571 395
rect -11493 349 -11447 395
rect -11369 349 -11323 395
rect -11245 349 -11199 395
rect -11121 349 -11075 395
rect -10997 349 -10951 395
rect -10873 349 -10827 395
rect -10749 349 -10703 395
rect -10625 349 -10579 395
rect -10501 349 -10455 395
rect -10377 349 -10331 395
rect -10253 349 -10207 395
rect -10129 349 -10083 395
rect -10005 349 -9959 395
rect -9881 349 -9835 395
rect -9757 349 -9711 395
rect -9633 349 -9587 395
rect -9509 349 -9463 395
rect -9385 349 -9339 395
rect -9261 349 -9215 395
rect -9137 349 -9091 395
rect -9013 349 -8967 395
rect -8889 349 -8843 395
rect -8765 349 -8719 395
rect -8641 349 -8595 395
rect -8517 349 -8471 395
rect -8393 349 -8347 395
rect -8269 349 -8223 395
rect -8145 349 -8099 395
rect -8021 349 -7975 395
rect -7897 349 -7851 395
rect -7773 349 -7727 395
rect -7649 349 -7603 395
rect -7525 349 -7479 395
rect -7401 349 -7355 395
rect -7277 349 -7231 395
rect -7153 349 -7107 395
rect -7029 349 -6983 395
rect -6905 349 -6859 395
rect -6781 349 -6735 395
rect -6657 349 -6611 395
rect -6533 349 -6487 395
rect -6409 349 -6363 395
rect -6285 349 -6239 395
rect -6161 349 -6115 395
rect -6037 349 -5991 395
rect -5913 349 -5867 395
rect -5789 349 -5743 395
rect -5665 349 -5619 395
rect -5541 349 -5495 395
rect -5417 349 -5371 395
rect -5293 349 -5247 395
rect -5169 349 -5123 395
rect -5045 349 -4999 395
rect -4921 349 -4875 395
rect -4797 349 -4751 395
rect -4673 349 -4627 395
rect -4549 349 -4503 395
rect -4425 349 -4379 395
rect -4301 349 -4255 395
rect -4177 349 -4131 395
rect -4053 349 -4007 395
rect -3929 349 -3883 395
rect -3805 349 -3759 395
rect -3681 349 -3635 395
rect -3557 349 -3511 395
rect -3433 349 -3387 395
rect -3309 349 -3263 395
rect -3185 349 -3139 395
rect -3061 349 -3015 395
rect -2937 349 -2891 395
rect -2813 349 -2767 395
rect -2689 349 -2643 395
rect -2565 349 -2519 395
rect -2441 349 -2395 395
rect -2317 349 -2271 395
rect -2193 349 -2147 395
rect -2069 349 -2023 395
rect -1945 349 -1899 395
rect -1821 349 -1775 395
rect -1697 349 -1651 395
rect -1573 349 -1527 395
rect -1449 349 -1403 395
rect -1325 349 -1279 395
rect -1201 349 -1155 395
rect -1077 349 -1031 395
rect -953 349 -907 395
rect -829 349 -783 395
rect -705 349 -659 395
rect -581 349 -535 395
rect -457 349 -411 395
rect -333 349 -287 395
rect -209 349 -163 395
rect -85 349 -39 395
rect 39 349 85 395
rect 163 349 209 395
rect 287 349 333 395
rect 411 349 457 395
rect 535 349 581 395
rect 659 349 705 395
rect 783 349 829 395
rect 907 349 953 395
rect 1031 349 1077 395
rect 1155 349 1201 395
rect 1279 349 1325 395
rect 1403 349 1449 395
rect 1527 349 1573 395
rect 1651 349 1697 395
rect 1775 349 1821 395
rect 1899 349 1945 395
rect 2023 349 2069 395
rect 2147 349 2193 395
rect 2271 349 2317 395
rect 2395 349 2441 395
rect 2519 349 2565 395
rect 2643 349 2689 395
rect 2767 349 2813 395
rect 2891 349 2937 395
rect 3015 349 3061 395
rect 3139 349 3185 395
rect 3263 349 3309 395
rect 3387 349 3433 395
rect 3511 349 3557 395
rect 3635 349 3681 395
rect 3759 349 3805 395
rect 3883 349 3929 395
rect 4007 349 4053 395
rect 4131 349 4177 395
rect 4255 349 4301 395
rect 4379 349 4425 395
rect 4503 349 4549 395
rect 4627 349 4673 395
rect 4751 349 4797 395
rect 4875 349 4921 395
rect 4999 349 5045 395
rect 5123 349 5169 395
rect 5247 349 5293 395
rect 5371 349 5417 395
rect 5495 349 5541 395
rect 5619 349 5665 395
rect 5743 349 5789 395
rect 5867 349 5913 395
rect 5991 349 6037 395
rect 6115 349 6161 395
rect 6239 349 6285 395
rect 6363 349 6409 395
rect 6487 349 6533 395
rect 6611 349 6657 395
rect 6735 349 6781 395
rect 6859 349 6905 395
rect 6983 349 7029 395
rect 7107 349 7153 395
rect 7231 349 7277 395
rect 7355 349 7401 395
rect 7479 349 7525 395
rect 7603 349 7649 395
rect 7727 349 7773 395
rect 7851 349 7897 395
rect 7975 349 8021 395
rect 8099 349 8145 395
rect 8223 349 8269 395
rect 8347 349 8393 395
rect 8471 349 8517 395
rect 8595 349 8641 395
rect 8719 349 8765 395
rect 8843 349 8889 395
rect 8967 349 9013 395
rect 9091 349 9137 395
rect 9215 349 9261 395
rect 9339 349 9385 395
rect 9463 349 9509 395
rect 9587 349 9633 395
rect 9711 349 9757 395
rect 9835 349 9881 395
rect 9959 349 10005 395
rect 10083 349 10129 395
rect 10207 349 10253 395
rect 10331 349 10377 395
rect 10455 349 10501 395
rect 10579 349 10625 395
rect 10703 349 10749 395
rect 10827 349 10873 395
rect 10951 349 10997 395
rect 11075 349 11121 395
rect 11199 349 11245 395
rect 11323 349 11369 395
rect 11447 349 11493 395
rect 11571 349 11617 395
rect 11695 349 11741 395
rect 11819 349 11865 395
rect 11943 349 11989 395
rect 12067 349 12113 395
rect 12191 349 12237 395
rect 12315 349 12361 395
rect 12439 349 12485 395
rect 12563 349 12609 395
rect 12687 349 12733 395
rect 12811 349 12857 395
rect 12935 349 12981 395
rect 13059 349 13105 395
rect 13183 349 13229 395
rect 13307 349 13353 395
rect 13431 349 13477 395
rect 13555 349 13601 395
rect 13679 349 13725 395
rect 13803 349 13849 395
rect 13927 349 13973 395
rect 14051 349 14097 395
rect 14175 349 14221 395
rect 14299 349 14345 395
rect 14423 349 14469 395
rect 14547 349 14593 395
rect 14671 349 14717 395
rect 14795 349 14841 395
rect 14919 349 14965 395
rect 15043 349 15089 395
rect 15167 349 15213 395
rect 15291 349 15337 395
rect 15415 349 15461 395
rect 15539 349 15585 395
rect 15663 349 15709 395
rect 15787 349 15833 395
rect 15911 349 15957 395
rect 16035 349 16081 395
rect 16159 349 16205 395
rect 16283 349 16329 395
rect 16407 349 16453 395
rect 16531 349 16577 395
rect 16655 349 16701 395
rect 16779 349 16825 395
rect 16903 349 16949 395
rect 17027 349 17073 395
rect 17151 349 17197 395
rect 17275 349 17321 395
rect 17399 349 17445 395
rect 17523 349 17569 395
rect 17647 349 17693 395
rect 17771 349 17817 395
rect 17895 349 17941 395
rect 18019 349 18065 395
rect 18143 349 18189 395
rect 18267 349 18313 395
rect -18313 225 -18267 271
rect -18189 225 -18143 271
rect -18065 225 -18019 271
rect -17941 225 -17895 271
rect -17817 225 -17771 271
rect -17693 225 -17647 271
rect -17569 225 -17523 271
rect -17445 225 -17399 271
rect -17321 225 -17275 271
rect -17197 225 -17151 271
rect -17073 225 -17027 271
rect -16949 225 -16903 271
rect -16825 225 -16779 271
rect -16701 225 -16655 271
rect -16577 225 -16531 271
rect -16453 225 -16407 271
rect -16329 225 -16283 271
rect -16205 225 -16159 271
rect -16081 225 -16035 271
rect -15957 225 -15911 271
rect -15833 225 -15787 271
rect -15709 225 -15663 271
rect -15585 225 -15539 271
rect -15461 225 -15415 271
rect -15337 225 -15291 271
rect -15213 225 -15167 271
rect -15089 225 -15043 271
rect -14965 225 -14919 271
rect -14841 225 -14795 271
rect -14717 225 -14671 271
rect -14593 225 -14547 271
rect -14469 225 -14423 271
rect -14345 225 -14299 271
rect -14221 225 -14175 271
rect -14097 225 -14051 271
rect -13973 225 -13927 271
rect -13849 225 -13803 271
rect -13725 225 -13679 271
rect -13601 225 -13555 271
rect -13477 225 -13431 271
rect -13353 225 -13307 271
rect -13229 225 -13183 271
rect -13105 225 -13059 271
rect -12981 225 -12935 271
rect -12857 225 -12811 271
rect -12733 225 -12687 271
rect -12609 225 -12563 271
rect -12485 225 -12439 271
rect -12361 225 -12315 271
rect -12237 225 -12191 271
rect -12113 225 -12067 271
rect -11989 225 -11943 271
rect -11865 225 -11819 271
rect -11741 225 -11695 271
rect -11617 225 -11571 271
rect -11493 225 -11447 271
rect -11369 225 -11323 271
rect -11245 225 -11199 271
rect -11121 225 -11075 271
rect -10997 225 -10951 271
rect -10873 225 -10827 271
rect -10749 225 -10703 271
rect -10625 225 -10579 271
rect -10501 225 -10455 271
rect -10377 225 -10331 271
rect -10253 225 -10207 271
rect -10129 225 -10083 271
rect -10005 225 -9959 271
rect -9881 225 -9835 271
rect -9757 225 -9711 271
rect -9633 225 -9587 271
rect -9509 225 -9463 271
rect -9385 225 -9339 271
rect -9261 225 -9215 271
rect -9137 225 -9091 271
rect -9013 225 -8967 271
rect -8889 225 -8843 271
rect -8765 225 -8719 271
rect -8641 225 -8595 271
rect -8517 225 -8471 271
rect -8393 225 -8347 271
rect -8269 225 -8223 271
rect -8145 225 -8099 271
rect -8021 225 -7975 271
rect -7897 225 -7851 271
rect -7773 225 -7727 271
rect -7649 225 -7603 271
rect -7525 225 -7479 271
rect -7401 225 -7355 271
rect -7277 225 -7231 271
rect -7153 225 -7107 271
rect -7029 225 -6983 271
rect -6905 225 -6859 271
rect -6781 225 -6735 271
rect -6657 225 -6611 271
rect -6533 225 -6487 271
rect -6409 225 -6363 271
rect -6285 225 -6239 271
rect -6161 225 -6115 271
rect -6037 225 -5991 271
rect -5913 225 -5867 271
rect -5789 225 -5743 271
rect -5665 225 -5619 271
rect -5541 225 -5495 271
rect -5417 225 -5371 271
rect -5293 225 -5247 271
rect -5169 225 -5123 271
rect -5045 225 -4999 271
rect -4921 225 -4875 271
rect -4797 225 -4751 271
rect -4673 225 -4627 271
rect -4549 225 -4503 271
rect -4425 225 -4379 271
rect -4301 225 -4255 271
rect -4177 225 -4131 271
rect -4053 225 -4007 271
rect -3929 225 -3883 271
rect -3805 225 -3759 271
rect -3681 225 -3635 271
rect -3557 225 -3511 271
rect -3433 225 -3387 271
rect -3309 225 -3263 271
rect -3185 225 -3139 271
rect -3061 225 -3015 271
rect -2937 225 -2891 271
rect -2813 225 -2767 271
rect -2689 225 -2643 271
rect -2565 225 -2519 271
rect -2441 225 -2395 271
rect -2317 225 -2271 271
rect -2193 225 -2147 271
rect -2069 225 -2023 271
rect -1945 225 -1899 271
rect -1821 225 -1775 271
rect -1697 225 -1651 271
rect -1573 225 -1527 271
rect -1449 225 -1403 271
rect -1325 225 -1279 271
rect -1201 225 -1155 271
rect -1077 225 -1031 271
rect -953 225 -907 271
rect -829 225 -783 271
rect -705 225 -659 271
rect -581 225 -535 271
rect -457 225 -411 271
rect -333 225 -287 271
rect -209 225 -163 271
rect -85 225 -39 271
rect 39 225 85 271
rect 163 225 209 271
rect 287 225 333 271
rect 411 225 457 271
rect 535 225 581 271
rect 659 225 705 271
rect 783 225 829 271
rect 907 225 953 271
rect 1031 225 1077 271
rect 1155 225 1201 271
rect 1279 225 1325 271
rect 1403 225 1449 271
rect 1527 225 1573 271
rect 1651 225 1697 271
rect 1775 225 1821 271
rect 1899 225 1945 271
rect 2023 225 2069 271
rect 2147 225 2193 271
rect 2271 225 2317 271
rect 2395 225 2441 271
rect 2519 225 2565 271
rect 2643 225 2689 271
rect 2767 225 2813 271
rect 2891 225 2937 271
rect 3015 225 3061 271
rect 3139 225 3185 271
rect 3263 225 3309 271
rect 3387 225 3433 271
rect 3511 225 3557 271
rect 3635 225 3681 271
rect 3759 225 3805 271
rect 3883 225 3929 271
rect 4007 225 4053 271
rect 4131 225 4177 271
rect 4255 225 4301 271
rect 4379 225 4425 271
rect 4503 225 4549 271
rect 4627 225 4673 271
rect 4751 225 4797 271
rect 4875 225 4921 271
rect 4999 225 5045 271
rect 5123 225 5169 271
rect 5247 225 5293 271
rect 5371 225 5417 271
rect 5495 225 5541 271
rect 5619 225 5665 271
rect 5743 225 5789 271
rect 5867 225 5913 271
rect 5991 225 6037 271
rect 6115 225 6161 271
rect 6239 225 6285 271
rect 6363 225 6409 271
rect 6487 225 6533 271
rect 6611 225 6657 271
rect 6735 225 6781 271
rect 6859 225 6905 271
rect 6983 225 7029 271
rect 7107 225 7153 271
rect 7231 225 7277 271
rect 7355 225 7401 271
rect 7479 225 7525 271
rect 7603 225 7649 271
rect 7727 225 7773 271
rect 7851 225 7897 271
rect 7975 225 8021 271
rect 8099 225 8145 271
rect 8223 225 8269 271
rect 8347 225 8393 271
rect 8471 225 8517 271
rect 8595 225 8641 271
rect 8719 225 8765 271
rect 8843 225 8889 271
rect 8967 225 9013 271
rect 9091 225 9137 271
rect 9215 225 9261 271
rect 9339 225 9385 271
rect 9463 225 9509 271
rect 9587 225 9633 271
rect 9711 225 9757 271
rect 9835 225 9881 271
rect 9959 225 10005 271
rect 10083 225 10129 271
rect 10207 225 10253 271
rect 10331 225 10377 271
rect 10455 225 10501 271
rect 10579 225 10625 271
rect 10703 225 10749 271
rect 10827 225 10873 271
rect 10951 225 10997 271
rect 11075 225 11121 271
rect 11199 225 11245 271
rect 11323 225 11369 271
rect 11447 225 11493 271
rect 11571 225 11617 271
rect 11695 225 11741 271
rect 11819 225 11865 271
rect 11943 225 11989 271
rect 12067 225 12113 271
rect 12191 225 12237 271
rect 12315 225 12361 271
rect 12439 225 12485 271
rect 12563 225 12609 271
rect 12687 225 12733 271
rect 12811 225 12857 271
rect 12935 225 12981 271
rect 13059 225 13105 271
rect 13183 225 13229 271
rect 13307 225 13353 271
rect 13431 225 13477 271
rect 13555 225 13601 271
rect 13679 225 13725 271
rect 13803 225 13849 271
rect 13927 225 13973 271
rect 14051 225 14097 271
rect 14175 225 14221 271
rect 14299 225 14345 271
rect 14423 225 14469 271
rect 14547 225 14593 271
rect 14671 225 14717 271
rect 14795 225 14841 271
rect 14919 225 14965 271
rect 15043 225 15089 271
rect 15167 225 15213 271
rect 15291 225 15337 271
rect 15415 225 15461 271
rect 15539 225 15585 271
rect 15663 225 15709 271
rect 15787 225 15833 271
rect 15911 225 15957 271
rect 16035 225 16081 271
rect 16159 225 16205 271
rect 16283 225 16329 271
rect 16407 225 16453 271
rect 16531 225 16577 271
rect 16655 225 16701 271
rect 16779 225 16825 271
rect 16903 225 16949 271
rect 17027 225 17073 271
rect 17151 225 17197 271
rect 17275 225 17321 271
rect 17399 225 17445 271
rect 17523 225 17569 271
rect 17647 225 17693 271
rect 17771 225 17817 271
rect 17895 225 17941 271
rect 18019 225 18065 271
rect 18143 225 18189 271
rect 18267 225 18313 271
rect -18313 101 -18267 147
rect -18189 101 -18143 147
rect -18065 101 -18019 147
rect -17941 101 -17895 147
rect -17817 101 -17771 147
rect -17693 101 -17647 147
rect -17569 101 -17523 147
rect -17445 101 -17399 147
rect -17321 101 -17275 147
rect -17197 101 -17151 147
rect -17073 101 -17027 147
rect -16949 101 -16903 147
rect -16825 101 -16779 147
rect -16701 101 -16655 147
rect -16577 101 -16531 147
rect -16453 101 -16407 147
rect -16329 101 -16283 147
rect -16205 101 -16159 147
rect -16081 101 -16035 147
rect -15957 101 -15911 147
rect -15833 101 -15787 147
rect -15709 101 -15663 147
rect -15585 101 -15539 147
rect -15461 101 -15415 147
rect -15337 101 -15291 147
rect -15213 101 -15167 147
rect -15089 101 -15043 147
rect -14965 101 -14919 147
rect -14841 101 -14795 147
rect -14717 101 -14671 147
rect -14593 101 -14547 147
rect -14469 101 -14423 147
rect -14345 101 -14299 147
rect -14221 101 -14175 147
rect -14097 101 -14051 147
rect -13973 101 -13927 147
rect -13849 101 -13803 147
rect -13725 101 -13679 147
rect -13601 101 -13555 147
rect -13477 101 -13431 147
rect -13353 101 -13307 147
rect -13229 101 -13183 147
rect -13105 101 -13059 147
rect -12981 101 -12935 147
rect -12857 101 -12811 147
rect -12733 101 -12687 147
rect -12609 101 -12563 147
rect -12485 101 -12439 147
rect -12361 101 -12315 147
rect -12237 101 -12191 147
rect -12113 101 -12067 147
rect -11989 101 -11943 147
rect -11865 101 -11819 147
rect -11741 101 -11695 147
rect -11617 101 -11571 147
rect -11493 101 -11447 147
rect -11369 101 -11323 147
rect -11245 101 -11199 147
rect -11121 101 -11075 147
rect -10997 101 -10951 147
rect -10873 101 -10827 147
rect -10749 101 -10703 147
rect -10625 101 -10579 147
rect -10501 101 -10455 147
rect -10377 101 -10331 147
rect -10253 101 -10207 147
rect -10129 101 -10083 147
rect -10005 101 -9959 147
rect -9881 101 -9835 147
rect -9757 101 -9711 147
rect -9633 101 -9587 147
rect -9509 101 -9463 147
rect -9385 101 -9339 147
rect -9261 101 -9215 147
rect -9137 101 -9091 147
rect -9013 101 -8967 147
rect -8889 101 -8843 147
rect -8765 101 -8719 147
rect -8641 101 -8595 147
rect -8517 101 -8471 147
rect -8393 101 -8347 147
rect -8269 101 -8223 147
rect -8145 101 -8099 147
rect -8021 101 -7975 147
rect -7897 101 -7851 147
rect -7773 101 -7727 147
rect -7649 101 -7603 147
rect -7525 101 -7479 147
rect -7401 101 -7355 147
rect -7277 101 -7231 147
rect -7153 101 -7107 147
rect -7029 101 -6983 147
rect -6905 101 -6859 147
rect -6781 101 -6735 147
rect -6657 101 -6611 147
rect -6533 101 -6487 147
rect -6409 101 -6363 147
rect -6285 101 -6239 147
rect -6161 101 -6115 147
rect -6037 101 -5991 147
rect -5913 101 -5867 147
rect -5789 101 -5743 147
rect -5665 101 -5619 147
rect -5541 101 -5495 147
rect -5417 101 -5371 147
rect -5293 101 -5247 147
rect -5169 101 -5123 147
rect -5045 101 -4999 147
rect -4921 101 -4875 147
rect -4797 101 -4751 147
rect -4673 101 -4627 147
rect -4549 101 -4503 147
rect -4425 101 -4379 147
rect -4301 101 -4255 147
rect -4177 101 -4131 147
rect -4053 101 -4007 147
rect -3929 101 -3883 147
rect -3805 101 -3759 147
rect -3681 101 -3635 147
rect -3557 101 -3511 147
rect -3433 101 -3387 147
rect -3309 101 -3263 147
rect -3185 101 -3139 147
rect -3061 101 -3015 147
rect -2937 101 -2891 147
rect -2813 101 -2767 147
rect -2689 101 -2643 147
rect -2565 101 -2519 147
rect -2441 101 -2395 147
rect -2317 101 -2271 147
rect -2193 101 -2147 147
rect -2069 101 -2023 147
rect -1945 101 -1899 147
rect -1821 101 -1775 147
rect -1697 101 -1651 147
rect -1573 101 -1527 147
rect -1449 101 -1403 147
rect -1325 101 -1279 147
rect -1201 101 -1155 147
rect -1077 101 -1031 147
rect -953 101 -907 147
rect -829 101 -783 147
rect -705 101 -659 147
rect -581 101 -535 147
rect -457 101 -411 147
rect -333 101 -287 147
rect -209 101 -163 147
rect -85 101 -39 147
rect 39 101 85 147
rect 163 101 209 147
rect 287 101 333 147
rect 411 101 457 147
rect 535 101 581 147
rect 659 101 705 147
rect 783 101 829 147
rect 907 101 953 147
rect 1031 101 1077 147
rect 1155 101 1201 147
rect 1279 101 1325 147
rect 1403 101 1449 147
rect 1527 101 1573 147
rect 1651 101 1697 147
rect 1775 101 1821 147
rect 1899 101 1945 147
rect 2023 101 2069 147
rect 2147 101 2193 147
rect 2271 101 2317 147
rect 2395 101 2441 147
rect 2519 101 2565 147
rect 2643 101 2689 147
rect 2767 101 2813 147
rect 2891 101 2937 147
rect 3015 101 3061 147
rect 3139 101 3185 147
rect 3263 101 3309 147
rect 3387 101 3433 147
rect 3511 101 3557 147
rect 3635 101 3681 147
rect 3759 101 3805 147
rect 3883 101 3929 147
rect 4007 101 4053 147
rect 4131 101 4177 147
rect 4255 101 4301 147
rect 4379 101 4425 147
rect 4503 101 4549 147
rect 4627 101 4673 147
rect 4751 101 4797 147
rect 4875 101 4921 147
rect 4999 101 5045 147
rect 5123 101 5169 147
rect 5247 101 5293 147
rect 5371 101 5417 147
rect 5495 101 5541 147
rect 5619 101 5665 147
rect 5743 101 5789 147
rect 5867 101 5913 147
rect 5991 101 6037 147
rect 6115 101 6161 147
rect 6239 101 6285 147
rect 6363 101 6409 147
rect 6487 101 6533 147
rect 6611 101 6657 147
rect 6735 101 6781 147
rect 6859 101 6905 147
rect 6983 101 7029 147
rect 7107 101 7153 147
rect 7231 101 7277 147
rect 7355 101 7401 147
rect 7479 101 7525 147
rect 7603 101 7649 147
rect 7727 101 7773 147
rect 7851 101 7897 147
rect 7975 101 8021 147
rect 8099 101 8145 147
rect 8223 101 8269 147
rect 8347 101 8393 147
rect 8471 101 8517 147
rect 8595 101 8641 147
rect 8719 101 8765 147
rect 8843 101 8889 147
rect 8967 101 9013 147
rect 9091 101 9137 147
rect 9215 101 9261 147
rect 9339 101 9385 147
rect 9463 101 9509 147
rect 9587 101 9633 147
rect 9711 101 9757 147
rect 9835 101 9881 147
rect 9959 101 10005 147
rect 10083 101 10129 147
rect 10207 101 10253 147
rect 10331 101 10377 147
rect 10455 101 10501 147
rect 10579 101 10625 147
rect 10703 101 10749 147
rect 10827 101 10873 147
rect 10951 101 10997 147
rect 11075 101 11121 147
rect 11199 101 11245 147
rect 11323 101 11369 147
rect 11447 101 11493 147
rect 11571 101 11617 147
rect 11695 101 11741 147
rect 11819 101 11865 147
rect 11943 101 11989 147
rect 12067 101 12113 147
rect 12191 101 12237 147
rect 12315 101 12361 147
rect 12439 101 12485 147
rect 12563 101 12609 147
rect 12687 101 12733 147
rect 12811 101 12857 147
rect 12935 101 12981 147
rect 13059 101 13105 147
rect 13183 101 13229 147
rect 13307 101 13353 147
rect 13431 101 13477 147
rect 13555 101 13601 147
rect 13679 101 13725 147
rect 13803 101 13849 147
rect 13927 101 13973 147
rect 14051 101 14097 147
rect 14175 101 14221 147
rect 14299 101 14345 147
rect 14423 101 14469 147
rect 14547 101 14593 147
rect 14671 101 14717 147
rect 14795 101 14841 147
rect 14919 101 14965 147
rect 15043 101 15089 147
rect 15167 101 15213 147
rect 15291 101 15337 147
rect 15415 101 15461 147
rect 15539 101 15585 147
rect 15663 101 15709 147
rect 15787 101 15833 147
rect 15911 101 15957 147
rect 16035 101 16081 147
rect 16159 101 16205 147
rect 16283 101 16329 147
rect 16407 101 16453 147
rect 16531 101 16577 147
rect 16655 101 16701 147
rect 16779 101 16825 147
rect 16903 101 16949 147
rect 17027 101 17073 147
rect 17151 101 17197 147
rect 17275 101 17321 147
rect 17399 101 17445 147
rect 17523 101 17569 147
rect 17647 101 17693 147
rect 17771 101 17817 147
rect 17895 101 17941 147
rect 18019 101 18065 147
rect 18143 101 18189 147
rect 18267 101 18313 147
rect -18313 -23 -18267 23
rect -18189 -23 -18143 23
rect -18065 -23 -18019 23
rect -17941 -23 -17895 23
rect -17817 -23 -17771 23
rect -17693 -23 -17647 23
rect -17569 -23 -17523 23
rect -17445 -23 -17399 23
rect -17321 -23 -17275 23
rect -17197 -23 -17151 23
rect -17073 -23 -17027 23
rect -16949 -23 -16903 23
rect -16825 -23 -16779 23
rect -16701 -23 -16655 23
rect -16577 -23 -16531 23
rect -16453 -23 -16407 23
rect -16329 -23 -16283 23
rect -16205 -23 -16159 23
rect -16081 -23 -16035 23
rect -15957 -23 -15911 23
rect -15833 -23 -15787 23
rect -15709 -23 -15663 23
rect -15585 -23 -15539 23
rect -15461 -23 -15415 23
rect -15337 -23 -15291 23
rect -15213 -23 -15167 23
rect -15089 -23 -15043 23
rect -14965 -23 -14919 23
rect -14841 -23 -14795 23
rect -14717 -23 -14671 23
rect -14593 -23 -14547 23
rect -14469 -23 -14423 23
rect -14345 -23 -14299 23
rect -14221 -23 -14175 23
rect -14097 -23 -14051 23
rect -13973 -23 -13927 23
rect -13849 -23 -13803 23
rect -13725 -23 -13679 23
rect -13601 -23 -13555 23
rect -13477 -23 -13431 23
rect -13353 -23 -13307 23
rect -13229 -23 -13183 23
rect -13105 -23 -13059 23
rect -12981 -23 -12935 23
rect -12857 -23 -12811 23
rect -12733 -23 -12687 23
rect -12609 -23 -12563 23
rect -12485 -23 -12439 23
rect -12361 -23 -12315 23
rect -12237 -23 -12191 23
rect -12113 -23 -12067 23
rect -11989 -23 -11943 23
rect -11865 -23 -11819 23
rect -11741 -23 -11695 23
rect -11617 -23 -11571 23
rect -11493 -23 -11447 23
rect -11369 -23 -11323 23
rect -11245 -23 -11199 23
rect -11121 -23 -11075 23
rect -10997 -23 -10951 23
rect -10873 -23 -10827 23
rect -10749 -23 -10703 23
rect -10625 -23 -10579 23
rect -10501 -23 -10455 23
rect -10377 -23 -10331 23
rect -10253 -23 -10207 23
rect -10129 -23 -10083 23
rect -10005 -23 -9959 23
rect -9881 -23 -9835 23
rect -9757 -23 -9711 23
rect -9633 -23 -9587 23
rect -9509 -23 -9463 23
rect -9385 -23 -9339 23
rect -9261 -23 -9215 23
rect -9137 -23 -9091 23
rect -9013 -23 -8967 23
rect -8889 -23 -8843 23
rect -8765 -23 -8719 23
rect -8641 -23 -8595 23
rect -8517 -23 -8471 23
rect -8393 -23 -8347 23
rect -8269 -23 -8223 23
rect -8145 -23 -8099 23
rect -8021 -23 -7975 23
rect -7897 -23 -7851 23
rect -7773 -23 -7727 23
rect -7649 -23 -7603 23
rect -7525 -23 -7479 23
rect -7401 -23 -7355 23
rect -7277 -23 -7231 23
rect -7153 -23 -7107 23
rect -7029 -23 -6983 23
rect -6905 -23 -6859 23
rect -6781 -23 -6735 23
rect -6657 -23 -6611 23
rect -6533 -23 -6487 23
rect -6409 -23 -6363 23
rect -6285 -23 -6239 23
rect -6161 -23 -6115 23
rect -6037 -23 -5991 23
rect -5913 -23 -5867 23
rect -5789 -23 -5743 23
rect -5665 -23 -5619 23
rect -5541 -23 -5495 23
rect -5417 -23 -5371 23
rect -5293 -23 -5247 23
rect -5169 -23 -5123 23
rect -5045 -23 -4999 23
rect -4921 -23 -4875 23
rect -4797 -23 -4751 23
rect -4673 -23 -4627 23
rect -4549 -23 -4503 23
rect -4425 -23 -4379 23
rect -4301 -23 -4255 23
rect -4177 -23 -4131 23
rect -4053 -23 -4007 23
rect -3929 -23 -3883 23
rect -3805 -23 -3759 23
rect -3681 -23 -3635 23
rect -3557 -23 -3511 23
rect -3433 -23 -3387 23
rect -3309 -23 -3263 23
rect -3185 -23 -3139 23
rect -3061 -23 -3015 23
rect -2937 -23 -2891 23
rect -2813 -23 -2767 23
rect -2689 -23 -2643 23
rect -2565 -23 -2519 23
rect -2441 -23 -2395 23
rect -2317 -23 -2271 23
rect -2193 -23 -2147 23
rect -2069 -23 -2023 23
rect -1945 -23 -1899 23
rect -1821 -23 -1775 23
rect -1697 -23 -1651 23
rect -1573 -23 -1527 23
rect -1449 -23 -1403 23
rect -1325 -23 -1279 23
rect -1201 -23 -1155 23
rect -1077 -23 -1031 23
rect -953 -23 -907 23
rect -829 -23 -783 23
rect -705 -23 -659 23
rect -581 -23 -535 23
rect -457 -23 -411 23
rect -333 -23 -287 23
rect -209 -23 -163 23
rect -85 -23 -39 23
rect 39 -23 85 23
rect 163 -23 209 23
rect 287 -23 333 23
rect 411 -23 457 23
rect 535 -23 581 23
rect 659 -23 705 23
rect 783 -23 829 23
rect 907 -23 953 23
rect 1031 -23 1077 23
rect 1155 -23 1201 23
rect 1279 -23 1325 23
rect 1403 -23 1449 23
rect 1527 -23 1573 23
rect 1651 -23 1697 23
rect 1775 -23 1821 23
rect 1899 -23 1945 23
rect 2023 -23 2069 23
rect 2147 -23 2193 23
rect 2271 -23 2317 23
rect 2395 -23 2441 23
rect 2519 -23 2565 23
rect 2643 -23 2689 23
rect 2767 -23 2813 23
rect 2891 -23 2937 23
rect 3015 -23 3061 23
rect 3139 -23 3185 23
rect 3263 -23 3309 23
rect 3387 -23 3433 23
rect 3511 -23 3557 23
rect 3635 -23 3681 23
rect 3759 -23 3805 23
rect 3883 -23 3929 23
rect 4007 -23 4053 23
rect 4131 -23 4177 23
rect 4255 -23 4301 23
rect 4379 -23 4425 23
rect 4503 -23 4549 23
rect 4627 -23 4673 23
rect 4751 -23 4797 23
rect 4875 -23 4921 23
rect 4999 -23 5045 23
rect 5123 -23 5169 23
rect 5247 -23 5293 23
rect 5371 -23 5417 23
rect 5495 -23 5541 23
rect 5619 -23 5665 23
rect 5743 -23 5789 23
rect 5867 -23 5913 23
rect 5991 -23 6037 23
rect 6115 -23 6161 23
rect 6239 -23 6285 23
rect 6363 -23 6409 23
rect 6487 -23 6533 23
rect 6611 -23 6657 23
rect 6735 -23 6781 23
rect 6859 -23 6905 23
rect 6983 -23 7029 23
rect 7107 -23 7153 23
rect 7231 -23 7277 23
rect 7355 -23 7401 23
rect 7479 -23 7525 23
rect 7603 -23 7649 23
rect 7727 -23 7773 23
rect 7851 -23 7897 23
rect 7975 -23 8021 23
rect 8099 -23 8145 23
rect 8223 -23 8269 23
rect 8347 -23 8393 23
rect 8471 -23 8517 23
rect 8595 -23 8641 23
rect 8719 -23 8765 23
rect 8843 -23 8889 23
rect 8967 -23 9013 23
rect 9091 -23 9137 23
rect 9215 -23 9261 23
rect 9339 -23 9385 23
rect 9463 -23 9509 23
rect 9587 -23 9633 23
rect 9711 -23 9757 23
rect 9835 -23 9881 23
rect 9959 -23 10005 23
rect 10083 -23 10129 23
rect 10207 -23 10253 23
rect 10331 -23 10377 23
rect 10455 -23 10501 23
rect 10579 -23 10625 23
rect 10703 -23 10749 23
rect 10827 -23 10873 23
rect 10951 -23 10997 23
rect 11075 -23 11121 23
rect 11199 -23 11245 23
rect 11323 -23 11369 23
rect 11447 -23 11493 23
rect 11571 -23 11617 23
rect 11695 -23 11741 23
rect 11819 -23 11865 23
rect 11943 -23 11989 23
rect 12067 -23 12113 23
rect 12191 -23 12237 23
rect 12315 -23 12361 23
rect 12439 -23 12485 23
rect 12563 -23 12609 23
rect 12687 -23 12733 23
rect 12811 -23 12857 23
rect 12935 -23 12981 23
rect 13059 -23 13105 23
rect 13183 -23 13229 23
rect 13307 -23 13353 23
rect 13431 -23 13477 23
rect 13555 -23 13601 23
rect 13679 -23 13725 23
rect 13803 -23 13849 23
rect 13927 -23 13973 23
rect 14051 -23 14097 23
rect 14175 -23 14221 23
rect 14299 -23 14345 23
rect 14423 -23 14469 23
rect 14547 -23 14593 23
rect 14671 -23 14717 23
rect 14795 -23 14841 23
rect 14919 -23 14965 23
rect 15043 -23 15089 23
rect 15167 -23 15213 23
rect 15291 -23 15337 23
rect 15415 -23 15461 23
rect 15539 -23 15585 23
rect 15663 -23 15709 23
rect 15787 -23 15833 23
rect 15911 -23 15957 23
rect 16035 -23 16081 23
rect 16159 -23 16205 23
rect 16283 -23 16329 23
rect 16407 -23 16453 23
rect 16531 -23 16577 23
rect 16655 -23 16701 23
rect 16779 -23 16825 23
rect 16903 -23 16949 23
rect 17027 -23 17073 23
rect 17151 -23 17197 23
rect 17275 -23 17321 23
rect 17399 -23 17445 23
rect 17523 -23 17569 23
rect 17647 -23 17693 23
rect 17771 -23 17817 23
rect 17895 -23 17941 23
rect 18019 -23 18065 23
rect 18143 -23 18189 23
rect 18267 -23 18313 23
rect -18313 -147 -18267 -101
rect -18189 -147 -18143 -101
rect -18065 -147 -18019 -101
rect -17941 -147 -17895 -101
rect -17817 -147 -17771 -101
rect -17693 -147 -17647 -101
rect -17569 -147 -17523 -101
rect -17445 -147 -17399 -101
rect -17321 -147 -17275 -101
rect -17197 -147 -17151 -101
rect -17073 -147 -17027 -101
rect -16949 -147 -16903 -101
rect -16825 -147 -16779 -101
rect -16701 -147 -16655 -101
rect -16577 -147 -16531 -101
rect -16453 -147 -16407 -101
rect -16329 -147 -16283 -101
rect -16205 -147 -16159 -101
rect -16081 -147 -16035 -101
rect -15957 -147 -15911 -101
rect -15833 -147 -15787 -101
rect -15709 -147 -15663 -101
rect -15585 -147 -15539 -101
rect -15461 -147 -15415 -101
rect -15337 -147 -15291 -101
rect -15213 -147 -15167 -101
rect -15089 -147 -15043 -101
rect -14965 -147 -14919 -101
rect -14841 -147 -14795 -101
rect -14717 -147 -14671 -101
rect -14593 -147 -14547 -101
rect -14469 -147 -14423 -101
rect -14345 -147 -14299 -101
rect -14221 -147 -14175 -101
rect -14097 -147 -14051 -101
rect -13973 -147 -13927 -101
rect -13849 -147 -13803 -101
rect -13725 -147 -13679 -101
rect -13601 -147 -13555 -101
rect -13477 -147 -13431 -101
rect -13353 -147 -13307 -101
rect -13229 -147 -13183 -101
rect -13105 -147 -13059 -101
rect -12981 -147 -12935 -101
rect -12857 -147 -12811 -101
rect -12733 -147 -12687 -101
rect -12609 -147 -12563 -101
rect -12485 -147 -12439 -101
rect -12361 -147 -12315 -101
rect -12237 -147 -12191 -101
rect -12113 -147 -12067 -101
rect -11989 -147 -11943 -101
rect -11865 -147 -11819 -101
rect -11741 -147 -11695 -101
rect -11617 -147 -11571 -101
rect -11493 -147 -11447 -101
rect -11369 -147 -11323 -101
rect -11245 -147 -11199 -101
rect -11121 -147 -11075 -101
rect -10997 -147 -10951 -101
rect -10873 -147 -10827 -101
rect -10749 -147 -10703 -101
rect -10625 -147 -10579 -101
rect -10501 -147 -10455 -101
rect -10377 -147 -10331 -101
rect -10253 -147 -10207 -101
rect -10129 -147 -10083 -101
rect -10005 -147 -9959 -101
rect -9881 -147 -9835 -101
rect -9757 -147 -9711 -101
rect -9633 -147 -9587 -101
rect -9509 -147 -9463 -101
rect -9385 -147 -9339 -101
rect -9261 -147 -9215 -101
rect -9137 -147 -9091 -101
rect -9013 -147 -8967 -101
rect -8889 -147 -8843 -101
rect -8765 -147 -8719 -101
rect -8641 -147 -8595 -101
rect -8517 -147 -8471 -101
rect -8393 -147 -8347 -101
rect -8269 -147 -8223 -101
rect -8145 -147 -8099 -101
rect -8021 -147 -7975 -101
rect -7897 -147 -7851 -101
rect -7773 -147 -7727 -101
rect -7649 -147 -7603 -101
rect -7525 -147 -7479 -101
rect -7401 -147 -7355 -101
rect -7277 -147 -7231 -101
rect -7153 -147 -7107 -101
rect -7029 -147 -6983 -101
rect -6905 -147 -6859 -101
rect -6781 -147 -6735 -101
rect -6657 -147 -6611 -101
rect -6533 -147 -6487 -101
rect -6409 -147 -6363 -101
rect -6285 -147 -6239 -101
rect -6161 -147 -6115 -101
rect -6037 -147 -5991 -101
rect -5913 -147 -5867 -101
rect -5789 -147 -5743 -101
rect -5665 -147 -5619 -101
rect -5541 -147 -5495 -101
rect -5417 -147 -5371 -101
rect -5293 -147 -5247 -101
rect -5169 -147 -5123 -101
rect -5045 -147 -4999 -101
rect -4921 -147 -4875 -101
rect -4797 -147 -4751 -101
rect -4673 -147 -4627 -101
rect -4549 -147 -4503 -101
rect -4425 -147 -4379 -101
rect -4301 -147 -4255 -101
rect -4177 -147 -4131 -101
rect -4053 -147 -4007 -101
rect -3929 -147 -3883 -101
rect -3805 -147 -3759 -101
rect -3681 -147 -3635 -101
rect -3557 -147 -3511 -101
rect -3433 -147 -3387 -101
rect -3309 -147 -3263 -101
rect -3185 -147 -3139 -101
rect -3061 -147 -3015 -101
rect -2937 -147 -2891 -101
rect -2813 -147 -2767 -101
rect -2689 -147 -2643 -101
rect -2565 -147 -2519 -101
rect -2441 -147 -2395 -101
rect -2317 -147 -2271 -101
rect -2193 -147 -2147 -101
rect -2069 -147 -2023 -101
rect -1945 -147 -1899 -101
rect -1821 -147 -1775 -101
rect -1697 -147 -1651 -101
rect -1573 -147 -1527 -101
rect -1449 -147 -1403 -101
rect -1325 -147 -1279 -101
rect -1201 -147 -1155 -101
rect -1077 -147 -1031 -101
rect -953 -147 -907 -101
rect -829 -147 -783 -101
rect -705 -147 -659 -101
rect -581 -147 -535 -101
rect -457 -147 -411 -101
rect -333 -147 -287 -101
rect -209 -147 -163 -101
rect -85 -147 -39 -101
rect 39 -147 85 -101
rect 163 -147 209 -101
rect 287 -147 333 -101
rect 411 -147 457 -101
rect 535 -147 581 -101
rect 659 -147 705 -101
rect 783 -147 829 -101
rect 907 -147 953 -101
rect 1031 -147 1077 -101
rect 1155 -147 1201 -101
rect 1279 -147 1325 -101
rect 1403 -147 1449 -101
rect 1527 -147 1573 -101
rect 1651 -147 1697 -101
rect 1775 -147 1821 -101
rect 1899 -147 1945 -101
rect 2023 -147 2069 -101
rect 2147 -147 2193 -101
rect 2271 -147 2317 -101
rect 2395 -147 2441 -101
rect 2519 -147 2565 -101
rect 2643 -147 2689 -101
rect 2767 -147 2813 -101
rect 2891 -147 2937 -101
rect 3015 -147 3061 -101
rect 3139 -147 3185 -101
rect 3263 -147 3309 -101
rect 3387 -147 3433 -101
rect 3511 -147 3557 -101
rect 3635 -147 3681 -101
rect 3759 -147 3805 -101
rect 3883 -147 3929 -101
rect 4007 -147 4053 -101
rect 4131 -147 4177 -101
rect 4255 -147 4301 -101
rect 4379 -147 4425 -101
rect 4503 -147 4549 -101
rect 4627 -147 4673 -101
rect 4751 -147 4797 -101
rect 4875 -147 4921 -101
rect 4999 -147 5045 -101
rect 5123 -147 5169 -101
rect 5247 -147 5293 -101
rect 5371 -147 5417 -101
rect 5495 -147 5541 -101
rect 5619 -147 5665 -101
rect 5743 -147 5789 -101
rect 5867 -147 5913 -101
rect 5991 -147 6037 -101
rect 6115 -147 6161 -101
rect 6239 -147 6285 -101
rect 6363 -147 6409 -101
rect 6487 -147 6533 -101
rect 6611 -147 6657 -101
rect 6735 -147 6781 -101
rect 6859 -147 6905 -101
rect 6983 -147 7029 -101
rect 7107 -147 7153 -101
rect 7231 -147 7277 -101
rect 7355 -147 7401 -101
rect 7479 -147 7525 -101
rect 7603 -147 7649 -101
rect 7727 -147 7773 -101
rect 7851 -147 7897 -101
rect 7975 -147 8021 -101
rect 8099 -147 8145 -101
rect 8223 -147 8269 -101
rect 8347 -147 8393 -101
rect 8471 -147 8517 -101
rect 8595 -147 8641 -101
rect 8719 -147 8765 -101
rect 8843 -147 8889 -101
rect 8967 -147 9013 -101
rect 9091 -147 9137 -101
rect 9215 -147 9261 -101
rect 9339 -147 9385 -101
rect 9463 -147 9509 -101
rect 9587 -147 9633 -101
rect 9711 -147 9757 -101
rect 9835 -147 9881 -101
rect 9959 -147 10005 -101
rect 10083 -147 10129 -101
rect 10207 -147 10253 -101
rect 10331 -147 10377 -101
rect 10455 -147 10501 -101
rect 10579 -147 10625 -101
rect 10703 -147 10749 -101
rect 10827 -147 10873 -101
rect 10951 -147 10997 -101
rect 11075 -147 11121 -101
rect 11199 -147 11245 -101
rect 11323 -147 11369 -101
rect 11447 -147 11493 -101
rect 11571 -147 11617 -101
rect 11695 -147 11741 -101
rect 11819 -147 11865 -101
rect 11943 -147 11989 -101
rect 12067 -147 12113 -101
rect 12191 -147 12237 -101
rect 12315 -147 12361 -101
rect 12439 -147 12485 -101
rect 12563 -147 12609 -101
rect 12687 -147 12733 -101
rect 12811 -147 12857 -101
rect 12935 -147 12981 -101
rect 13059 -147 13105 -101
rect 13183 -147 13229 -101
rect 13307 -147 13353 -101
rect 13431 -147 13477 -101
rect 13555 -147 13601 -101
rect 13679 -147 13725 -101
rect 13803 -147 13849 -101
rect 13927 -147 13973 -101
rect 14051 -147 14097 -101
rect 14175 -147 14221 -101
rect 14299 -147 14345 -101
rect 14423 -147 14469 -101
rect 14547 -147 14593 -101
rect 14671 -147 14717 -101
rect 14795 -147 14841 -101
rect 14919 -147 14965 -101
rect 15043 -147 15089 -101
rect 15167 -147 15213 -101
rect 15291 -147 15337 -101
rect 15415 -147 15461 -101
rect 15539 -147 15585 -101
rect 15663 -147 15709 -101
rect 15787 -147 15833 -101
rect 15911 -147 15957 -101
rect 16035 -147 16081 -101
rect 16159 -147 16205 -101
rect 16283 -147 16329 -101
rect 16407 -147 16453 -101
rect 16531 -147 16577 -101
rect 16655 -147 16701 -101
rect 16779 -147 16825 -101
rect 16903 -147 16949 -101
rect 17027 -147 17073 -101
rect 17151 -147 17197 -101
rect 17275 -147 17321 -101
rect 17399 -147 17445 -101
rect 17523 -147 17569 -101
rect 17647 -147 17693 -101
rect 17771 -147 17817 -101
rect 17895 -147 17941 -101
rect 18019 -147 18065 -101
rect 18143 -147 18189 -101
rect 18267 -147 18313 -101
rect -18313 -271 -18267 -225
rect -18189 -271 -18143 -225
rect -18065 -271 -18019 -225
rect -17941 -271 -17895 -225
rect -17817 -271 -17771 -225
rect -17693 -271 -17647 -225
rect -17569 -271 -17523 -225
rect -17445 -271 -17399 -225
rect -17321 -271 -17275 -225
rect -17197 -271 -17151 -225
rect -17073 -271 -17027 -225
rect -16949 -271 -16903 -225
rect -16825 -271 -16779 -225
rect -16701 -271 -16655 -225
rect -16577 -271 -16531 -225
rect -16453 -271 -16407 -225
rect -16329 -271 -16283 -225
rect -16205 -271 -16159 -225
rect -16081 -271 -16035 -225
rect -15957 -271 -15911 -225
rect -15833 -271 -15787 -225
rect -15709 -271 -15663 -225
rect -15585 -271 -15539 -225
rect -15461 -271 -15415 -225
rect -15337 -271 -15291 -225
rect -15213 -271 -15167 -225
rect -15089 -271 -15043 -225
rect -14965 -271 -14919 -225
rect -14841 -271 -14795 -225
rect -14717 -271 -14671 -225
rect -14593 -271 -14547 -225
rect -14469 -271 -14423 -225
rect -14345 -271 -14299 -225
rect -14221 -271 -14175 -225
rect -14097 -271 -14051 -225
rect -13973 -271 -13927 -225
rect -13849 -271 -13803 -225
rect -13725 -271 -13679 -225
rect -13601 -271 -13555 -225
rect -13477 -271 -13431 -225
rect -13353 -271 -13307 -225
rect -13229 -271 -13183 -225
rect -13105 -271 -13059 -225
rect -12981 -271 -12935 -225
rect -12857 -271 -12811 -225
rect -12733 -271 -12687 -225
rect -12609 -271 -12563 -225
rect -12485 -271 -12439 -225
rect -12361 -271 -12315 -225
rect -12237 -271 -12191 -225
rect -12113 -271 -12067 -225
rect -11989 -271 -11943 -225
rect -11865 -271 -11819 -225
rect -11741 -271 -11695 -225
rect -11617 -271 -11571 -225
rect -11493 -271 -11447 -225
rect -11369 -271 -11323 -225
rect -11245 -271 -11199 -225
rect -11121 -271 -11075 -225
rect -10997 -271 -10951 -225
rect -10873 -271 -10827 -225
rect -10749 -271 -10703 -225
rect -10625 -271 -10579 -225
rect -10501 -271 -10455 -225
rect -10377 -271 -10331 -225
rect -10253 -271 -10207 -225
rect -10129 -271 -10083 -225
rect -10005 -271 -9959 -225
rect -9881 -271 -9835 -225
rect -9757 -271 -9711 -225
rect -9633 -271 -9587 -225
rect -9509 -271 -9463 -225
rect -9385 -271 -9339 -225
rect -9261 -271 -9215 -225
rect -9137 -271 -9091 -225
rect -9013 -271 -8967 -225
rect -8889 -271 -8843 -225
rect -8765 -271 -8719 -225
rect -8641 -271 -8595 -225
rect -8517 -271 -8471 -225
rect -8393 -271 -8347 -225
rect -8269 -271 -8223 -225
rect -8145 -271 -8099 -225
rect -8021 -271 -7975 -225
rect -7897 -271 -7851 -225
rect -7773 -271 -7727 -225
rect -7649 -271 -7603 -225
rect -7525 -271 -7479 -225
rect -7401 -271 -7355 -225
rect -7277 -271 -7231 -225
rect -7153 -271 -7107 -225
rect -7029 -271 -6983 -225
rect -6905 -271 -6859 -225
rect -6781 -271 -6735 -225
rect -6657 -271 -6611 -225
rect -6533 -271 -6487 -225
rect -6409 -271 -6363 -225
rect -6285 -271 -6239 -225
rect -6161 -271 -6115 -225
rect -6037 -271 -5991 -225
rect -5913 -271 -5867 -225
rect -5789 -271 -5743 -225
rect -5665 -271 -5619 -225
rect -5541 -271 -5495 -225
rect -5417 -271 -5371 -225
rect -5293 -271 -5247 -225
rect -5169 -271 -5123 -225
rect -5045 -271 -4999 -225
rect -4921 -271 -4875 -225
rect -4797 -271 -4751 -225
rect -4673 -271 -4627 -225
rect -4549 -271 -4503 -225
rect -4425 -271 -4379 -225
rect -4301 -271 -4255 -225
rect -4177 -271 -4131 -225
rect -4053 -271 -4007 -225
rect -3929 -271 -3883 -225
rect -3805 -271 -3759 -225
rect -3681 -271 -3635 -225
rect -3557 -271 -3511 -225
rect -3433 -271 -3387 -225
rect -3309 -271 -3263 -225
rect -3185 -271 -3139 -225
rect -3061 -271 -3015 -225
rect -2937 -271 -2891 -225
rect -2813 -271 -2767 -225
rect -2689 -271 -2643 -225
rect -2565 -271 -2519 -225
rect -2441 -271 -2395 -225
rect -2317 -271 -2271 -225
rect -2193 -271 -2147 -225
rect -2069 -271 -2023 -225
rect -1945 -271 -1899 -225
rect -1821 -271 -1775 -225
rect -1697 -271 -1651 -225
rect -1573 -271 -1527 -225
rect -1449 -271 -1403 -225
rect -1325 -271 -1279 -225
rect -1201 -271 -1155 -225
rect -1077 -271 -1031 -225
rect -953 -271 -907 -225
rect -829 -271 -783 -225
rect -705 -271 -659 -225
rect -581 -271 -535 -225
rect -457 -271 -411 -225
rect -333 -271 -287 -225
rect -209 -271 -163 -225
rect -85 -271 -39 -225
rect 39 -271 85 -225
rect 163 -271 209 -225
rect 287 -271 333 -225
rect 411 -271 457 -225
rect 535 -271 581 -225
rect 659 -271 705 -225
rect 783 -271 829 -225
rect 907 -271 953 -225
rect 1031 -271 1077 -225
rect 1155 -271 1201 -225
rect 1279 -271 1325 -225
rect 1403 -271 1449 -225
rect 1527 -271 1573 -225
rect 1651 -271 1697 -225
rect 1775 -271 1821 -225
rect 1899 -271 1945 -225
rect 2023 -271 2069 -225
rect 2147 -271 2193 -225
rect 2271 -271 2317 -225
rect 2395 -271 2441 -225
rect 2519 -271 2565 -225
rect 2643 -271 2689 -225
rect 2767 -271 2813 -225
rect 2891 -271 2937 -225
rect 3015 -271 3061 -225
rect 3139 -271 3185 -225
rect 3263 -271 3309 -225
rect 3387 -271 3433 -225
rect 3511 -271 3557 -225
rect 3635 -271 3681 -225
rect 3759 -271 3805 -225
rect 3883 -271 3929 -225
rect 4007 -271 4053 -225
rect 4131 -271 4177 -225
rect 4255 -271 4301 -225
rect 4379 -271 4425 -225
rect 4503 -271 4549 -225
rect 4627 -271 4673 -225
rect 4751 -271 4797 -225
rect 4875 -271 4921 -225
rect 4999 -271 5045 -225
rect 5123 -271 5169 -225
rect 5247 -271 5293 -225
rect 5371 -271 5417 -225
rect 5495 -271 5541 -225
rect 5619 -271 5665 -225
rect 5743 -271 5789 -225
rect 5867 -271 5913 -225
rect 5991 -271 6037 -225
rect 6115 -271 6161 -225
rect 6239 -271 6285 -225
rect 6363 -271 6409 -225
rect 6487 -271 6533 -225
rect 6611 -271 6657 -225
rect 6735 -271 6781 -225
rect 6859 -271 6905 -225
rect 6983 -271 7029 -225
rect 7107 -271 7153 -225
rect 7231 -271 7277 -225
rect 7355 -271 7401 -225
rect 7479 -271 7525 -225
rect 7603 -271 7649 -225
rect 7727 -271 7773 -225
rect 7851 -271 7897 -225
rect 7975 -271 8021 -225
rect 8099 -271 8145 -225
rect 8223 -271 8269 -225
rect 8347 -271 8393 -225
rect 8471 -271 8517 -225
rect 8595 -271 8641 -225
rect 8719 -271 8765 -225
rect 8843 -271 8889 -225
rect 8967 -271 9013 -225
rect 9091 -271 9137 -225
rect 9215 -271 9261 -225
rect 9339 -271 9385 -225
rect 9463 -271 9509 -225
rect 9587 -271 9633 -225
rect 9711 -271 9757 -225
rect 9835 -271 9881 -225
rect 9959 -271 10005 -225
rect 10083 -271 10129 -225
rect 10207 -271 10253 -225
rect 10331 -271 10377 -225
rect 10455 -271 10501 -225
rect 10579 -271 10625 -225
rect 10703 -271 10749 -225
rect 10827 -271 10873 -225
rect 10951 -271 10997 -225
rect 11075 -271 11121 -225
rect 11199 -271 11245 -225
rect 11323 -271 11369 -225
rect 11447 -271 11493 -225
rect 11571 -271 11617 -225
rect 11695 -271 11741 -225
rect 11819 -271 11865 -225
rect 11943 -271 11989 -225
rect 12067 -271 12113 -225
rect 12191 -271 12237 -225
rect 12315 -271 12361 -225
rect 12439 -271 12485 -225
rect 12563 -271 12609 -225
rect 12687 -271 12733 -225
rect 12811 -271 12857 -225
rect 12935 -271 12981 -225
rect 13059 -271 13105 -225
rect 13183 -271 13229 -225
rect 13307 -271 13353 -225
rect 13431 -271 13477 -225
rect 13555 -271 13601 -225
rect 13679 -271 13725 -225
rect 13803 -271 13849 -225
rect 13927 -271 13973 -225
rect 14051 -271 14097 -225
rect 14175 -271 14221 -225
rect 14299 -271 14345 -225
rect 14423 -271 14469 -225
rect 14547 -271 14593 -225
rect 14671 -271 14717 -225
rect 14795 -271 14841 -225
rect 14919 -271 14965 -225
rect 15043 -271 15089 -225
rect 15167 -271 15213 -225
rect 15291 -271 15337 -225
rect 15415 -271 15461 -225
rect 15539 -271 15585 -225
rect 15663 -271 15709 -225
rect 15787 -271 15833 -225
rect 15911 -271 15957 -225
rect 16035 -271 16081 -225
rect 16159 -271 16205 -225
rect 16283 -271 16329 -225
rect 16407 -271 16453 -225
rect 16531 -271 16577 -225
rect 16655 -271 16701 -225
rect 16779 -271 16825 -225
rect 16903 -271 16949 -225
rect 17027 -271 17073 -225
rect 17151 -271 17197 -225
rect 17275 -271 17321 -225
rect 17399 -271 17445 -225
rect 17523 -271 17569 -225
rect 17647 -271 17693 -225
rect 17771 -271 17817 -225
rect 17895 -271 17941 -225
rect 18019 -271 18065 -225
rect 18143 -271 18189 -225
rect 18267 -271 18313 -225
rect -18313 -395 -18267 -349
rect -18189 -395 -18143 -349
rect -18065 -395 -18019 -349
rect -17941 -395 -17895 -349
rect -17817 -395 -17771 -349
rect -17693 -395 -17647 -349
rect -17569 -395 -17523 -349
rect -17445 -395 -17399 -349
rect -17321 -395 -17275 -349
rect -17197 -395 -17151 -349
rect -17073 -395 -17027 -349
rect -16949 -395 -16903 -349
rect -16825 -395 -16779 -349
rect -16701 -395 -16655 -349
rect -16577 -395 -16531 -349
rect -16453 -395 -16407 -349
rect -16329 -395 -16283 -349
rect -16205 -395 -16159 -349
rect -16081 -395 -16035 -349
rect -15957 -395 -15911 -349
rect -15833 -395 -15787 -349
rect -15709 -395 -15663 -349
rect -15585 -395 -15539 -349
rect -15461 -395 -15415 -349
rect -15337 -395 -15291 -349
rect -15213 -395 -15167 -349
rect -15089 -395 -15043 -349
rect -14965 -395 -14919 -349
rect -14841 -395 -14795 -349
rect -14717 -395 -14671 -349
rect -14593 -395 -14547 -349
rect -14469 -395 -14423 -349
rect -14345 -395 -14299 -349
rect -14221 -395 -14175 -349
rect -14097 -395 -14051 -349
rect -13973 -395 -13927 -349
rect -13849 -395 -13803 -349
rect -13725 -395 -13679 -349
rect -13601 -395 -13555 -349
rect -13477 -395 -13431 -349
rect -13353 -395 -13307 -349
rect -13229 -395 -13183 -349
rect -13105 -395 -13059 -349
rect -12981 -395 -12935 -349
rect -12857 -395 -12811 -349
rect -12733 -395 -12687 -349
rect -12609 -395 -12563 -349
rect -12485 -395 -12439 -349
rect -12361 -395 -12315 -349
rect -12237 -395 -12191 -349
rect -12113 -395 -12067 -349
rect -11989 -395 -11943 -349
rect -11865 -395 -11819 -349
rect -11741 -395 -11695 -349
rect -11617 -395 -11571 -349
rect -11493 -395 -11447 -349
rect -11369 -395 -11323 -349
rect -11245 -395 -11199 -349
rect -11121 -395 -11075 -349
rect -10997 -395 -10951 -349
rect -10873 -395 -10827 -349
rect -10749 -395 -10703 -349
rect -10625 -395 -10579 -349
rect -10501 -395 -10455 -349
rect -10377 -395 -10331 -349
rect -10253 -395 -10207 -349
rect -10129 -395 -10083 -349
rect -10005 -395 -9959 -349
rect -9881 -395 -9835 -349
rect -9757 -395 -9711 -349
rect -9633 -395 -9587 -349
rect -9509 -395 -9463 -349
rect -9385 -395 -9339 -349
rect -9261 -395 -9215 -349
rect -9137 -395 -9091 -349
rect -9013 -395 -8967 -349
rect -8889 -395 -8843 -349
rect -8765 -395 -8719 -349
rect -8641 -395 -8595 -349
rect -8517 -395 -8471 -349
rect -8393 -395 -8347 -349
rect -8269 -395 -8223 -349
rect -8145 -395 -8099 -349
rect -8021 -395 -7975 -349
rect -7897 -395 -7851 -349
rect -7773 -395 -7727 -349
rect -7649 -395 -7603 -349
rect -7525 -395 -7479 -349
rect -7401 -395 -7355 -349
rect -7277 -395 -7231 -349
rect -7153 -395 -7107 -349
rect -7029 -395 -6983 -349
rect -6905 -395 -6859 -349
rect -6781 -395 -6735 -349
rect -6657 -395 -6611 -349
rect -6533 -395 -6487 -349
rect -6409 -395 -6363 -349
rect -6285 -395 -6239 -349
rect -6161 -395 -6115 -349
rect -6037 -395 -5991 -349
rect -5913 -395 -5867 -349
rect -5789 -395 -5743 -349
rect -5665 -395 -5619 -349
rect -5541 -395 -5495 -349
rect -5417 -395 -5371 -349
rect -5293 -395 -5247 -349
rect -5169 -395 -5123 -349
rect -5045 -395 -4999 -349
rect -4921 -395 -4875 -349
rect -4797 -395 -4751 -349
rect -4673 -395 -4627 -349
rect -4549 -395 -4503 -349
rect -4425 -395 -4379 -349
rect -4301 -395 -4255 -349
rect -4177 -395 -4131 -349
rect -4053 -395 -4007 -349
rect -3929 -395 -3883 -349
rect -3805 -395 -3759 -349
rect -3681 -395 -3635 -349
rect -3557 -395 -3511 -349
rect -3433 -395 -3387 -349
rect -3309 -395 -3263 -349
rect -3185 -395 -3139 -349
rect -3061 -395 -3015 -349
rect -2937 -395 -2891 -349
rect -2813 -395 -2767 -349
rect -2689 -395 -2643 -349
rect -2565 -395 -2519 -349
rect -2441 -395 -2395 -349
rect -2317 -395 -2271 -349
rect -2193 -395 -2147 -349
rect -2069 -395 -2023 -349
rect -1945 -395 -1899 -349
rect -1821 -395 -1775 -349
rect -1697 -395 -1651 -349
rect -1573 -395 -1527 -349
rect -1449 -395 -1403 -349
rect -1325 -395 -1279 -349
rect -1201 -395 -1155 -349
rect -1077 -395 -1031 -349
rect -953 -395 -907 -349
rect -829 -395 -783 -349
rect -705 -395 -659 -349
rect -581 -395 -535 -349
rect -457 -395 -411 -349
rect -333 -395 -287 -349
rect -209 -395 -163 -349
rect -85 -395 -39 -349
rect 39 -395 85 -349
rect 163 -395 209 -349
rect 287 -395 333 -349
rect 411 -395 457 -349
rect 535 -395 581 -349
rect 659 -395 705 -349
rect 783 -395 829 -349
rect 907 -395 953 -349
rect 1031 -395 1077 -349
rect 1155 -395 1201 -349
rect 1279 -395 1325 -349
rect 1403 -395 1449 -349
rect 1527 -395 1573 -349
rect 1651 -395 1697 -349
rect 1775 -395 1821 -349
rect 1899 -395 1945 -349
rect 2023 -395 2069 -349
rect 2147 -395 2193 -349
rect 2271 -395 2317 -349
rect 2395 -395 2441 -349
rect 2519 -395 2565 -349
rect 2643 -395 2689 -349
rect 2767 -395 2813 -349
rect 2891 -395 2937 -349
rect 3015 -395 3061 -349
rect 3139 -395 3185 -349
rect 3263 -395 3309 -349
rect 3387 -395 3433 -349
rect 3511 -395 3557 -349
rect 3635 -395 3681 -349
rect 3759 -395 3805 -349
rect 3883 -395 3929 -349
rect 4007 -395 4053 -349
rect 4131 -395 4177 -349
rect 4255 -395 4301 -349
rect 4379 -395 4425 -349
rect 4503 -395 4549 -349
rect 4627 -395 4673 -349
rect 4751 -395 4797 -349
rect 4875 -395 4921 -349
rect 4999 -395 5045 -349
rect 5123 -395 5169 -349
rect 5247 -395 5293 -349
rect 5371 -395 5417 -349
rect 5495 -395 5541 -349
rect 5619 -395 5665 -349
rect 5743 -395 5789 -349
rect 5867 -395 5913 -349
rect 5991 -395 6037 -349
rect 6115 -395 6161 -349
rect 6239 -395 6285 -349
rect 6363 -395 6409 -349
rect 6487 -395 6533 -349
rect 6611 -395 6657 -349
rect 6735 -395 6781 -349
rect 6859 -395 6905 -349
rect 6983 -395 7029 -349
rect 7107 -395 7153 -349
rect 7231 -395 7277 -349
rect 7355 -395 7401 -349
rect 7479 -395 7525 -349
rect 7603 -395 7649 -349
rect 7727 -395 7773 -349
rect 7851 -395 7897 -349
rect 7975 -395 8021 -349
rect 8099 -395 8145 -349
rect 8223 -395 8269 -349
rect 8347 -395 8393 -349
rect 8471 -395 8517 -349
rect 8595 -395 8641 -349
rect 8719 -395 8765 -349
rect 8843 -395 8889 -349
rect 8967 -395 9013 -349
rect 9091 -395 9137 -349
rect 9215 -395 9261 -349
rect 9339 -395 9385 -349
rect 9463 -395 9509 -349
rect 9587 -395 9633 -349
rect 9711 -395 9757 -349
rect 9835 -395 9881 -349
rect 9959 -395 10005 -349
rect 10083 -395 10129 -349
rect 10207 -395 10253 -349
rect 10331 -395 10377 -349
rect 10455 -395 10501 -349
rect 10579 -395 10625 -349
rect 10703 -395 10749 -349
rect 10827 -395 10873 -349
rect 10951 -395 10997 -349
rect 11075 -395 11121 -349
rect 11199 -395 11245 -349
rect 11323 -395 11369 -349
rect 11447 -395 11493 -349
rect 11571 -395 11617 -349
rect 11695 -395 11741 -349
rect 11819 -395 11865 -349
rect 11943 -395 11989 -349
rect 12067 -395 12113 -349
rect 12191 -395 12237 -349
rect 12315 -395 12361 -349
rect 12439 -395 12485 -349
rect 12563 -395 12609 -349
rect 12687 -395 12733 -349
rect 12811 -395 12857 -349
rect 12935 -395 12981 -349
rect 13059 -395 13105 -349
rect 13183 -395 13229 -349
rect 13307 -395 13353 -349
rect 13431 -395 13477 -349
rect 13555 -395 13601 -349
rect 13679 -395 13725 -349
rect 13803 -395 13849 -349
rect 13927 -395 13973 -349
rect 14051 -395 14097 -349
rect 14175 -395 14221 -349
rect 14299 -395 14345 -349
rect 14423 -395 14469 -349
rect 14547 -395 14593 -349
rect 14671 -395 14717 -349
rect 14795 -395 14841 -349
rect 14919 -395 14965 -349
rect 15043 -395 15089 -349
rect 15167 -395 15213 -349
rect 15291 -395 15337 -349
rect 15415 -395 15461 -349
rect 15539 -395 15585 -349
rect 15663 -395 15709 -349
rect 15787 -395 15833 -349
rect 15911 -395 15957 -349
rect 16035 -395 16081 -349
rect 16159 -395 16205 -349
rect 16283 -395 16329 -349
rect 16407 -395 16453 -349
rect 16531 -395 16577 -349
rect 16655 -395 16701 -349
rect 16779 -395 16825 -349
rect 16903 -395 16949 -349
rect 17027 -395 17073 -349
rect 17151 -395 17197 -349
rect 17275 -395 17321 -349
rect 17399 -395 17445 -349
rect 17523 -395 17569 -349
rect 17647 -395 17693 -349
rect 17771 -395 17817 -349
rect 17895 -395 17941 -349
rect 18019 -395 18065 -349
rect 18143 -395 18189 -349
rect 18267 -395 18313 -349
rect -18313 -519 -18267 -473
rect -18189 -519 -18143 -473
rect -18065 -519 -18019 -473
rect -17941 -519 -17895 -473
rect -17817 -519 -17771 -473
rect -17693 -519 -17647 -473
rect -17569 -519 -17523 -473
rect -17445 -519 -17399 -473
rect -17321 -519 -17275 -473
rect -17197 -519 -17151 -473
rect -17073 -519 -17027 -473
rect -16949 -519 -16903 -473
rect -16825 -519 -16779 -473
rect -16701 -519 -16655 -473
rect -16577 -519 -16531 -473
rect -16453 -519 -16407 -473
rect -16329 -519 -16283 -473
rect -16205 -519 -16159 -473
rect -16081 -519 -16035 -473
rect -15957 -519 -15911 -473
rect -15833 -519 -15787 -473
rect -15709 -519 -15663 -473
rect -15585 -519 -15539 -473
rect -15461 -519 -15415 -473
rect -15337 -519 -15291 -473
rect -15213 -519 -15167 -473
rect -15089 -519 -15043 -473
rect -14965 -519 -14919 -473
rect -14841 -519 -14795 -473
rect -14717 -519 -14671 -473
rect -14593 -519 -14547 -473
rect -14469 -519 -14423 -473
rect -14345 -519 -14299 -473
rect -14221 -519 -14175 -473
rect -14097 -519 -14051 -473
rect -13973 -519 -13927 -473
rect -13849 -519 -13803 -473
rect -13725 -519 -13679 -473
rect -13601 -519 -13555 -473
rect -13477 -519 -13431 -473
rect -13353 -519 -13307 -473
rect -13229 -519 -13183 -473
rect -13105 -519 -13059 -473
rect -12981 -519 -12935 -473
rect -12857 -519 -12811 -473
rect -12733 -519 -12687 -473
rect -12609 -519 -12563 -473
rect -12485 -519 -12439 -473
rect -12361 -519 -12315 -473
rect -12237 -519 -12191 -473
rect -12113 -519 -12067 -473
rect -11989 -519 -11943 -473
rect -11865 -519 -11819 -473
rect -11741 -519 -11695 -473
rect -11617 -519 -11571 -473
rect -11493 -519 -11447 -473
rect -11369 -519 -11323 -473
rect -11245 -519 -11199 -473
rect -11121 -519 -11075 -473
rect -10997 -519 -10951 -473
rect -10873 -519 -10827 -473
rect -10749 -519 -10703 -473
rect -10625 -519 -10579 -473
rect -10501 -519 -10455 -473
rect -10377 -519 -10331 -473
rect -10253 -519 -10207 -473
rect -10129 -519 -10083 -473
rect -10005 -519 -9959 -473
rect -9881 -519 -9835 -473
rect -9757 -519 -9711 -473
rect -9633 -519 -9587 -473
rect -9509 -519 -9463 -473
rect -9385 -519 -9339 -473
rect -9261 -519 -9215 -473
rect -9137 -519 -9091 -473
rect -9013 -519 -8967 -473
rect -8889 -519 -8843 -473
rect -8765 -519 -8719 -473
rect -8641 -519 -8595 -473
rect -8517 -519 -8471 -473
rect -8393 -519 -8347 -473
rect -8269 -519 -8223 -473
rect -8145 -519 -8099 -473
rect -8021 -519 -7975 -473
rect -7897 -519 -7851 -473
rect -7773 -519 -7727 -473
rect -7649 -519 -7603 -473
rect -7525 -519 -7479 -473
rect -7401 -519 -7355 -473
rect -7277 -519 -7231 -473
rect -7153 -519 -7107 -473
rect -7029 -519 -6983 -473
rect -6905 -519 -6859 -473
rect -6781 -519 -6735 -473
rect -6657 -519 -6611 -473
rect -6533 -519 -6487 -473
rect -6409 -519 -6363 -473
rect -6285 -519 -6239 -473
rect -6161 -519 -6115 -473
rect -6037 -519 -5991 -473
rect -5913 -519 -5867 -473
rect -5789 -519 -5743 -473
rect -5665 -519 -5619 -473
rect -5541 -519 -5495 -473
rect -5417 -519 -5371 -473
rect -5293 -519 -5247 -473
rect -5169 -519 -5123 -473
rect -5045 -519 -4999 -473
rect -4921 -519 -4875 -473
rect -4797 -519 -4751 -473
rect -4673 -519 -4627 -473
rect -4549 -519 -4503 -473
rect -4425 -519 -4379 -473
rect -4301 -519 -4255 -473
rect -4177 -519 -4131 -473
rect -4053 -519 -4007 -473
rect -3929 -519 -3883 -473
rect -3805 -519 -3759 -473
rect -3681 -519 -3635 -473
rect -3557 -519 -3511 -473
rect -3433 -519 -3387 -473
rect -3309 -519 -3263 -473
rect -3185 -519 -3139 -473
rect -3061 -519 -3015 -473
rect -2937 -519 -2891 -473
rect -2813 -519 -2767 -473
rect -2689 -519 -2643 -473
rect -2565 -519 -2519 -473
rect -2441 -519 -2395 -473
rect -2317 -519 -2271 -473
rect -2193 -519 -2147 -473
rect -2069 -519 -2023 -473
rect -1945 -519 -1899 -473
rect -1821 -519 -1775 -473
rect -1697 -519 -1651 -473
rect -1573 -519 -1527 -473
rect -1449 -519 -1403 -473
rect -1325 -519 -1279 -473
rect -1201 -519 -1155 -473
rect -1077 -519 -1031 -473
rect -953 -519 -907 -473
rect -829 -519 -783 -473
rect -705 -519 -659 -473
rect -581 -519 -535 -473
rect -457 -519 -411 -473
rect -333 -519 -287 -473
rect -209 -519 -163 -473
rect -85 -519 -39 -473
rect 39 -519 85 -473
rect 163 -519 209 -473
rect 287 -519 333 -473
rect 411 -519 457 -473
rect 535 -519 581 -473
rect 659 -519 705 -473
rect 783 -519 829 -473
rect 907 -519 953 -473
rect 1031 -519 1077 -473
rect 1155 -519 1201 -473
rect 1279 -519 1325 -473
rect 1403 -519 1449 -473
rect 1527 -519 1573 -473
rect 1651 -519 1697 -473
rect 1775 -519 1821 -473
rect 1899 -519 1945 -473
rect 2023 -519 2069 -473
rect 2147 -519 2193 -473
rect 2271 -519 2317 -473
rect 2395 -519 2441 -473
rect 2519 -519 2565 -473
rect 2643 -519 2689 -473
rect 2767 -519 2813 -473
rect 2891 -519 2937 -473
rect 3015 -519 3061 -473
rect 3139 -519 3185 -473
rect 3263 -519 3309 -473
rect 3387 -519 3433 -473
rect 3511 -519 3557 -473
rect 3635 -519 3681 -473
rect 3759 -519 3805 -473
rect 3883 -519 3929 -473
rect 4007 -519 4053 -473
rect 4131 -519 4177 -473
rect 4255 -519 4301 -473
rect 4379 -519 4425 -473
rect 4503 -519 4549 -473
rect 4627 -519 4673 -473
rect 4751 -519 4797 -473
rect 4875 -519 4921 -473
rect 4999 -519 5045 -473
rect 5123 -519 5169 -473
rect 5247 -519 5293 -473
rect 5371 -519 5417 -473
rect 5495 -519 5541 -473
rect 5619 -519 5665 -473
rect 5743 -519 5789 -473
rect 5867 -519 5913 -473
rect 5991 -519 6037 -473
rect 6115 -519 6161 -473
rect 6239 -519 6285 -473
rect 6363 -519 6409 -473
rect 6487 -519 6533 -473
rect 6611 -519 6657 -473
rect 6735 -519 6781 -473
rect 6859 -519 6905 -473
rect 6983 -519 7029 -473
rect 7107 -519 7153 -473
rect 7231 -519 7277 -473
rect 7355 -519 7401 -473
rect 7479 -519 7525 -473
rect 7603 -519 7649 -473
rect 7727 -519 7773 -473
rect 7851 -519 7897 -473
rect 7975 -519 8021 -473
rect 8099 -519 8145 -473
rect 8223 -519 8269 -473
rect 8347 -519 8393 -473
rect 8471 -519 8517 -473
rect 8595 -519 8641 -473
rect 8719 -519 8765 -473
rect 8843 -519 8889 -473
rect 8967 -519 9013 -473
rect 9091 -519 9137 -473
rect 9215 -519 9261 -473
rect 9339 -519 9385 -473
rect 9463 -519 9509 -473
rect 9587 -519 9633 -473
rect 9711 -519 9757 -473
rect 9835 -519 9881 -473
rect 9959 -519 10005 -473
rect 10083 -519 10129 -473
rect 10207 -519 10253 -473
rect 10331 -519 10377 -473
rect 10455 -519 10501 -473
rect 10579 -519 10625 -473
rect 10703 -519 10749 -473
rect 10827 -519 10873 -473
rect 10951 -519 10997 -473
rect 11075 -519 11121 -473
rect 11199 -519 11245 -473
rect 11323 -519 11369 -473
rect 11447 -519 11493 -473
rect 11571 -519 11617 -473
rect 11695 -519 11741 -473
rect 11819 -519 11865 -473
rect 11943 -519 11989 -473
rect 12067 -519 12113 -473
rect 12191 -519 12237 -473
rect 12315 -519 12361 -473
rect 12439 -519 12485 -473
rect 12563 -519 12609 -473
rect 12687 -519 12733 -473
rect 12811 -519 12857 -473
rect 12935 -519 12981 -473
rect 13059 -519 13105 -473
rect 13183 -519 13229 -473
rect 13307 -519 13353 -473
rect 13431 -519 13477 -473
rect 13555 -519 13601 -473
rect 13679 -519 13725 -473
rect 13803 -519 13849 -473
rect 13927 -519 13973 -473
rect 14051 -519 14097 -473
rect 14175 -519 14221 -473
rect 14299 -519 14345 -473
rect 14423 -519 14469 -473
rect 14547 -519 14593 -473
rect 14671 -519 14717 -473
rect 14795 -519 14841 -473
rect 14919 -519 14965 -473
rect 15043 -519 15089 -473
rect 15167 -519 15213 -473
rect 15291 -519 15337 -473
rect 15415 -519 15461 -473
rect 15539 -519 15585 -473
rect 15663 -519 15709 -473
rect 15787 -519 15833 -473
rect 15911 -519 15957 -473
rect 16035 -519 16081 -473
rect 16159 -519 16205 -473
rect 16283 -519 16329 -473
rect 16407 -519 16453 -473
rect 16531 -519 16577 -473
rect 16655 -519 16701 -473
rect 16779 -519 16825 -473
rect 16903 -519 16949 -473
rect 17027 -519 17073 -473
rect 17151 -519 17197 -473
rect 17275 -519 17321 -473
rect 17399 -519 17445 -473
rect 17523 -519 17569 -473
rect 17647 -519 17693 -473
rect 17771 -519 17817 -473
rect 17895 -519 17941 -473
rect 18019 -519 18065 -473
rect 18143 -519 18189 -473
rect 18267 -519 18313 -473
rect -18313 -643 -18267 -597
rect -18189 -643 -18143 -597
rect -18065 -643 -18019 -597
rect -17941 -643 -17895 -597
rect -17817 -643 -17771 -597
rect -17693 -643 -17647 -597
rect -17569 -643 -17523 -597
rect -17445 -643 -17399 -597
rect -17321 -643 -17275 -597
rect -17197 -643 -17151 -597
rect -17073 -643 -17027 -597
rect -16949 -643 -16903 -597
rect -16825 -643 -16779 -597
rect -16701 -643 -16655 -597
rect -16577 -643 -16531 -597
rect -16453 -643 -16407 -597
rect -16329 -643 -16283 -597
rect -16205 -643 -16159 -597
rect -16081 -643 -16035 -597
rect -15957 -643 -15911 -597
rect -15833 -643 -15787 -597
rect -15709 -643 -15663 -597
rect -15585 -643 -15539 -597
rect -15461 -643 -15415 -597
rect -15337 -643 -15291 -597
rect -15213 -643 -15167 -597
rect -15089 -643 -15043 -597
rect -14965 -643 -14919 -597
rect -14841 -643 -14795 -597
rect -14717 -643 -14671 -597
rect -14593 -643 -14547 -597
rect -14469 -643 -14423 -597
rect -14345 -643 -14299 -597
rect -14221 -643 -14175 -597
rect -14097 -643 -14051 -597
rect -13973 -643 -13927 -597
rect -13849 -643 -13803 -597
rect -13725 -643 -13679 -597
rect -13601 -643 -13555 -597
rect -13477 -643 -13431 -597
rect -13353 -643 -13307 -597
rect -13229 -643 -13183 -597
rect -13105 -643 -13059 -597
rect -12981 -643 -12935 -597
rect -12857 -643 -12811 -597
rect -12733 -643 -12687 -597
rect -12609 -643 -12563 -597
rect -12485 -643 -12439 -597
rect -12361 -643 -12315 -597
rect -12237 -643 -12191 -597
rect -12113 -643 -12067 -597
rect -11989 -643 -11943 -597
rect -11865 -643 -11819 -597
rect -11741 -643 -11695 -597
rect -11617 -643 -11571 -597
rect -11493 -643 -11447 -597
rect -11369 -643 -11323 -597
rect -11245 -643 -11199 -597
rect -11121 -643 -11075 -597
rect -10997 -643 -10951 -597
rect -10873 -643 -10827 -597
rect -10749 -643 -10703 -597
rect -10625 -643 -10579 -597
rect -10501 -643 -10455 -597
rect -10377 -643 -10331 -597
rect -10253 -643 -10207 -597
rect -10129 -643 -10083 -597
rect -10005 -643 -9959 -597
rect -9881 -643 -9835 -597
rect -9757 -643 -9711 -597
rect -9633 -643 -9587 -597
rect -9509 -643 -9463 -597
rect -9385 -643 -9339 -597
rect -9261 -643 -9215 -597
rect -9137 -643 -9091 -597
rect -9013 -643 -8967 -597
rect -8889 -643 -8843 -597
rect -8765 -643 -8719 -597
rect -8641 -643 -8595 -597
rect -8517 -643 -8471 -597
rect -8393 -643 -8347 -597
rect -8269 -643 -8223 -597
rect -8145 -643 -8099 -597
rect -8021 -643 -7975 -597
rect -7897 -643 -7851 -597
rect -7773 -643 -7727 -597
rect -7649 -643 -7603 -597
rect -7525 -643 -7479 -597
rect -7401 -643 -7355 -597
rect -7277 -643 -7231 -597
rect -7153 -643 -7107 -597
rect -7029 -643 -6983 -597
rect -6905 -643 -6859 -597
rect -6781 -643 -6735 -597
rect -6657 -643 -6611 -597
rect -6533 -643 -6487 -597
rect -6409 -643 -6363 -597
rect -6285 -643 -6239 -597
rect -6161 -643 -6115 -597
rect -6037 -643 -5991 -597
rect -5913 -643 -5867 -597
rect -5789 -643 -5743 -597
rect -5665 -643 -5619 -597
rect -5541 -643 -5495 -597
rect -5417 -643 -5371 -597
rect -5293 -643 -5247 -597
rect -5169 -643 -5123 -597
rect -5045 -643 -4999 -597
rect -4921 -643 -4875 -597
rect -4797 -643 -4751 -597
rect -4673 -643 -4627 -597
rect -4549 -643 -4503 -597
rect -4425 -643 -4379 -597
rect -4301 -643 -4255 -597
rect -4177 -643 -4131 -597
rect -4053 -643 -4007 -597
rect -3929 -643 -3883 -597
rect -3805 -643 -3759 -597
rect -3681 -643 -3635 -597
rect -3557 -643 -3511 -597
rect -3433 -643 -3387 -597
rect -3309 -643 -3263 -597
rect -3185 -643 -3139 -597
rect -3061 -643 -3015 -597
rect -2937 -643 -2891 -597
rect -2813 -643 -2767 -597
rect -2689 -643 -2643 -597
rect -2565 -643 -2519 -597
rect -2441 -643 -2395 -597
rect -2317 -643 -2271 -597
rect -2193 -643 -2147 -597
rect -2069 -643 -2023 -597
rect -1945 -643 -1899 -597
rect -1821 -643 -1775 -597
rect -1697 -643 -1651 -597
rect -1573 -643 -1527 -597
rect -1449 -643 -1403 -597
rect -1325 -643 -1279 -597
rect -1201 -643 -1155 -597
rect -1077 -643 -1031 -597
rect -953 -643 -907 -597
rect -829 -643 -783 -597
rect -705 -643 -659 -597
rect -581 -643 -535 -597
rect -457 -643 -411 -597
rect -333 -643 -287 -597
rect -209 -643 -163 -597
rect -85 -643 -39 -597
rect 39 -643 85 -597
rect 163 -643 209 -597
rect 287 -643 333 -597
rect 411 -643 457 -597
rect 535 -643 581 -597
rect 659 -643 705 -597
rect 783 -643 829 -597
rect 907 -643 953 -597
rect 1031 -643 1077 -597
rect 1155 -643 1201 -597
rect 1279 -643 1325 -597
rect 1403 -643 1449 -597
rect 1527 -643 1573 -597
rect 1651 -643 1697 -597
rect 1775 -643 1821 -597
rect 1899 -643 1945 -597
rect 2023 -643 2069 -597
rect 2147 -643 2193 -597
rect 2271 -643 2317 -597
rect 2395 -643 2441 -597
rect 2519 -643 2565 -597
rect 2643 -643 2689 -597
rect 2767 -643 2813 -597
rect 2891 -643 2937 -597
rect 3015 -643 3061 -597
rect 3139 -643 3185 -597
rect 3263 -643 3309 -597
rect 3387 -643 3433 -597
rect 3511 -643 3557 -597
rect 3635 -643 3681 -597
rect 3759 -643 3805 -597
rect 3883 -643 3929 -597
rect 4007 -643 4053 -597
rect 4131 -643 4177 -597
rect 4255 -643 4301 -597
rect 4379 -643 4425 -597
rect 4503 -643 4549 -597
rect 4627 -643 4673 -597
rect 4751 -643 4797 -597
rect 4875 -643 4921 -597
rect 4999 -643 5045 -597
rect 5123 -643 5169 -597
rect 5247 -643 5293 -597
rect 5371 -643 5417 -597
rect 5495 -643 5541 -597
rect 5619 -643 5665 -597
rect 5743 -643 5789 -597
rect 5867 -643 5913 -597
rect 5991 -643 6037 -597
rect 6115 -643 6161 -597
rect 6239 -643 6285 -597
rect 6363 -643 6409 -597
rect 6487 -643 6533 -597
rect 6611 -643 6657 -597
rect 6735 -643 6781 -597
rect 6859 -643 6905 -597
rect 6983 -643 7029 -597
rect 7107 -643 7153 -597
rect 7231 -643 7277 -597
rect 7355 -643 7401 -597
rect 7479 -643 7525 -597
rect 7603 -643 7649 -597
rect 7727 -643 7773 -597
rect 7851 -643 7897 -597
rect 7975 -643 8021 -597
rect 8099 -643 8145 -597
rect 8223 -643 8269 -597
rect 8347 -643 8393 -597
rect 8471 -643 8517 -597
rect 8595 -643 8641 -597
rect 8719 -643 8765 -597
rect 8843 -643 8889 -597
rect 8967 -643 9013 -597
rect 9091 -643 9137 -597
rect 9215 -643 9261 -597
rect 9339 -643 9385 -597
rect 9463 -643 9509 -597
rect 9587 -643 9633 -597
rect 9711 -643 9757 -597
rect 9835 -643 9881 -597
rect 9959 -643 10005 -597
rect 10083 -643 10129 -597
rect 10207 -643 10253 -597
rect 10331 -643 10377 -597
rect 10455 -643 10501 -597
rect 10579 -643 10625 -597
rect 10703 -643 10749 -597
rect 10827 -643 10873 -597
rect 10951 -643 10997 -597
rect 11075 -643 11121 -597
rect 11199 -643 11245 -597
rect 11323 -643 11369 -597
rect 11447 -643 11493 -597
rect 11571 -643 11617 -597
rect 11695 -643 11741 -597
rect 11819 -643 11865 -597
rect 11943 -643 11989 -597
rect 12067 -643 12113 -597
rect 12191 -643 12237 -597
rect 12315 -643 12361 -597
rect 12439 -643 12485 -597
rect 12563 -643 12609 -597
rect 12687 -643 12733 -597
rect 12811 -643 12857 -597
rect 12935 -643 12981 -597
rect 13059 -643 13105 -597
rect 13183 -643 13229 -597
rect 13307 -643 13353 -597
rect 13431 -643 13477 -597
rect 13555 -643 13601 -597
rect 13679 -643 13725 -597
rect 13803 -643 13849 -597
rect 13927 -643 13973 -597
rect 14051 -643 14097 -597
rect 14175 -643 14221 -597
rect 14299 -643 14345 -597
rect 14423 -643 14469 -597
rect 14547 -643 14593 -597
rect 14671 -643 14717 -597
rect 14795 -643 14841 -597
rect 14919 -643 14965 -597
rect 15043 -643 15089 -597
rect 15167 -643 15213 -597
rect 15291 -643 15337 -597
rect 15415 -643 15461 -597
rect 15539 -643 15585 -597
rect 15663 -643 15709 -597
rect 15787 -643 15833 -597
rect 15911 -643 15957 -597
rect 16035 -643 16081 -597
rect 16159 -643 16205 -597
rect 16283 -643 16329 -597
rect 16407 -643 16453 -597
rect 16531 -643 16577 -597
rect 16655 -643 16701 -597
rect 16779 -643 16825 -597
rect 16903 -643 16949 -597
rect 17027 -643 17073 -597
rect 17151 -643 17197 -597
rect 17275 -643 17321 -597
rect 17399 -643 17445 -597
rect 17523 -643 17569 -597
rect 17647 -643 17693 -597
rect 17771 -643 17817 -597
rect 17895 -643 17941 -597
rect 18019 -643 18065 -597
rect 18143 -643 18189 -597
rect 18267 -643 18313 -597
<< metal1 >>
rect -18324 643 18324 654
rect -18324 597 -18313 643
rect -18267 597 -18189 643
rect -18143 597 -18065 643
rect -18019 597 -17941 643
rect -17895 597 -17817 643
rect -17771 597 -17693 643
rect -17647 597 -17569 643
rect -17523 597 -17445 643
rect -17399 597 -17321 643
rect -17275 597 -17197 643
rect -17151 597 -17073 643
rect -17027 597 -16949 643
rect -16903 597 -16825 643
rect -16779 597 -16701 643
rect -16655 597 -16577 643
rect -16531 597 -16453 643
rect -16407 597 -16329 643
rect -16283 597 -16205 643
rect -16159 597 -16081 643
rect -16035 597 -15957 643
rect -15911 597 -15833 643
rect -15787 597 -15709 643
rect -15663 597 -15585 643
rect -15539 597 -15461 643
rect -15415 597 -15337 643
rect -15291 597 -15213 643
rect -15167 597 -15089 643
rect -15043 597 -14965 643
rect -14919 597 -14841 643
rect -14795 597 -14717 643
rect -14671 597 -14593 643
rect -14547 597 -14469 643
rect -14423 597 -14345 643
rect -14299 597 -14221 643
rect -14175 597 -14097 643
rect -14051 597 -13973 643
rect -13927 597 -13849 643
rect -13803 597 -13725 643
rect -13679 597 -13601 643
rect -13555 597 -13477 643
rect -13431 597 -13353 643
rect -13307 597 -13229 643
rect -13183 597 -13105 643
rect -13059 597 -12981 643
rect -12935 597 -12857 643
rect -12811 597 -12733 643
rect -12687 597 -12609 643
rect -12563 597 -12485 643
rect -12439 597 -12361 643
rect -12315 597 -12237 643
rect -12191 597 -12113 643
rect -12067 597 -11989 643
rect -11943 597 -11865 643
rect -11819 597 -11741 643
rect -11695 597 -11617 643
rect -11571 597 -11493 643
rect -11447 597 -11369 643
rect -11323 597 -11245 643
rect -11199 597 -11121 643
rect -11075 597 -10997 643
rect -10951 597 -10873 643
rect -10827 597 -10749 643
rect -10703 597 -10625 643
rect -10579 597 -10501 643
rect -10455 597 -10377 643
rect -10331 597 -10253 643
rect -10207 597 -10129 643
rect -10083 597 -10005 643
rect -9959 597 -9881 643
rect -9835 597 -9757 643
rect -9711 597 -9633 643
rect -9587 597 -9509 643
rect -9463 597 -9385 643
rect -9339 597 -9261 643
rect -9215 597 -9137 643
rect -9091 597 -9013 643
rect -8967 597 -8889 643
rect -8843 597 -8765 643
rect -8719 597 -8641 643
rect -8595 597 -8517 643
rect -8471 597 -8393 643
rect -8347 597 -8269 643
rect -8223 597 -8145 643
rect -8099 597 -8021 643
rect -7975 597 -7897 643
rect -7851 597 -7773 643
rect -7727 597 -7649 643
rect -7603 597 -7525 643
rect -7479 597 -7401 643
rect -7355 597 -7277 643
rect -7231 597 -7153 643
rect -7107 597 -7029 643
rect -6983 597 -6905 643
rect -6859 597 -6781 643
rect -6735 597 -6657 643
rect -6611 597 -6533 643
rect -6487 597 -6409 643
rect -6363 597 -6285 643
rect -6239 597 -6161 643
rect -6115 597 -6037 643
rect -5991 597 -5913 643
rect -5867 597 -5789 643
rect -5743 597 -5665 643
rect -5619 597 -5541 643
rect -5495 597 -5417 643
rect -5371 597 -5293 643
rect -5247 597 -5169 643
rect -5123 597 -5045 643
rect -4999 597 -4921 643
rect -4875 597 -4797 643
rect -4751 597 -4673 643
rect -4627 597 -4549 643
rect -4503 597 -4425 643
rect -4379 597 -4301 643
rect -4255 597 -4177 643
rect -4131 597 -4053 643
rect -4007 597 -3929 643
rect -3883 597 -3805 643
rect -3759 597 -3681 643
rect -3635 597 -3557 643
rect -3511 597 -3433 643
rect -3387 597 -3309 643
rect -3263 597 -3185 643
rect -3139 597 -3061 643
rect -3015 597 -2937 643
rect -2891 597 -2813 643
rect -2767 597 -2689 643
rect -2643 597 -2565 643
rect -2519 597 -2441 643
rect -2395 597 -2317 643
rect -2271 597 -2193 643
rect -2147 597 -2069 643
rect -2023 597 -1945 643
rect -1899 597 -1821 643
rect -1775 597 -1697 643
rect -1651 597 -1573 643
rect -1527 597 -1449 643
rect -1403 597 -1325 643
rect -1279 597 -1201 643
rect -1155 597 -1077 643
rect -1031 597 -953 643
rect -907 597 -829 643
rect -783 597 -705 643
rect -659 597 -581 643
rect -535 597 -457 643
rect -411 597 -333 643
rect -287 597 -209 643
rect -163 597 -85 643
rect -39 597 39 643
rect 85 597 163 643
rect 209 597 287 643
rect 333 597 411 643
rect 457 597 535 643
rect 581 597 659 643
rect 705 597 783 643
rect 829 597 907 643
rect 953 597 1031 643
rect 1077 597 1155 643
rect 1201 597 1279 643
rect 1325 597 1403 643
rect 1449 597 1527 643
rect 1573 597 1651 643
rect 1697 597 1775 643
rect 1821 597 1899 643
rect 1945 597 2023 643
rect 2069 597 2147 643
rect 2193 597 2271 643
rect 2317 597 2395 643
rect 2441 597 2519 643
rect 2565 597 2643 643
rect 2689 597 2767 643
rect 2813 597 2891 643
rect 2937 597 3015 643
rect 3061 597 3139 643
rect 3185 597 3263 643
rect 3309 597 3387 643
rect 3433 597 3511 643
rect 3557 597 3635 643
rect 3681 597 3759 643
rect 3805 597 3883 643
rect 3929 597 4007 643
rect 4053 597 4131 643
rect 4177 597 4255 643
rect 4301 597 4379 643
rect 4425 597 4503 643
rect 4549 597 4627 643
rect 4673 597 4751 643
rect 4797 597 4875 643
rect 4921 597 4999 643
rect 5045 597 5123 643
rect 5169 597 5247 643
rect 5293 597 5371 643
rect 5417 597 5495 643
rect 5541 597 5619 643
rect 5665 597 5743 643
rect 5789 597 5867 643
rect 5913 597 5991 643
rect 6037 597 6115 643
rect 6161 597 6239 643
rect 6285 597 6363 643
rect 6409 597 6487 643
rect 6533 597 6611 643
rect 6657 597 6735 643
rect 6781 597 6859 643
rect 6905 597 6983 643
rect 7029 597 7107 643
rect 7153 597 7231 643
rect 7277 597 7355 643
rect 7401 597 7479 643
rect 7525 597 7603 643
rect 7649 597 7727 643
rect 7773 597 7851 643
rect 7897 597 7975 643
rect 8021 597 8099 643
rect 8145 597 8223 643
rect 8269 597 8347 643
rect 8393 597 8471 643
rect 8517 597 8595 643
rect 8641 597 8719 643
rect 8765 597 8843 643
rect 8889 597 8967 643
rect 9013 597 9091 643
rect 9137 597 9215 643
rect 9261 597 9339 643
rect 9385 597 9463 643
rect 9509 597 9587 643
rect 9633 597 9711 643
rect 9757 597 9835 643
rect 9881 597 9959 643
rect 10005 597 10083 643
rect 10129 597 10207 643
rect 10253 597 10331 643
rect 10377 597 10455 643
rect 10501 597 10579 643
rect 10625 597 10703 643
rect 10749 597 10827 643
rect 10873 597 10951 643
rect 10997 597 11075 643
rect 11121 597 11199 643
rect 11245 597 11323 643
rect 11369 597 11447 643
rect 11493 597 11571 643
rect 11617 597 11695 643
rect 11741 597 11819 643
rect 11865 597 11943 643
rect 11989 597 12067 643
rect 12113 597 12191 643
rect 12237 597 12315 643
rect 12361 597 12439 643
rect 12485 597 12563 643
rect 12609 597 12687 643
rect 12733 597 12811 643
rect 12857 597 12935 643
rect 12981 597 13059 643
rect 13105 597 13183 643
rect 13229 597 13307 643
rect 13353 597 13431 643
rect 13477 597 13555 643
rect 13601 597 13679 643
rect 13725 597 13803 643
rect 13849 597 13927 643
rect 13973 597 14051 643
rect 14097 597 14175 643
rect 14221 597 14299 643
rect 14345 597 14423 643
rect 14469 597 14547 643
rect 14593 597 14671 643
rect 14717 597 14795 643
rect 14841 597 14919 643
rect 14965 597 15043 643
rect 15089 597 15167 643
rect 15213 597 15291 643
rect 15337 597 15415 643
rect 15461 597 15539 643
rect 15585 597 15663 643
rect 15709 597 15787 643
rect 15833 597 15911 643
rect 15957 597 16035 643
rect 16081 597 16159 643
rect 16205 597 16283 643
rect 16329 597 16407 643
rect 16453 597 16531 643
rect 16577 597 16655 643
rect 16701 597 16779 643
rect 16825 597 16903 643
rect 16949 597 17027 643
rect 17073 597 17151 643
rect 17197 597 17275 643
rect 17321 597 17399 643
rect 17445 597 17523 643
rect 17569 597 17647 643
rect 17693 597 17771 643
rect 17817 597 17895 643
rect 17941 597 18019 643
rect 18065 597 18143 643
rect 18189 597 18267 643
rect 18313 597 18324 643
rect -18324 519 18324 597
rect -18324 473 -18313 519
rect -18267 473 -18189 519
rect -18143 473 -18065 519
rect -18019 473 -17941 519
rect -17895 473 -17817 519
rect -17771 473 -17693 519
rect -17647 473 -17569 519
rect -17523 473 -17445 519
rect -17399 473 -17321 519
rect -17275 473 -17197 519
rect -17151 473 -17073 519
rect -17027 473 -16949 519
rect -16903 473 -16825 519
rect -16779 473 -16701 519
rect -16655 473 -16577 519
rect -16531 473 -16453 519
rect -16407 473 -16329 519
rect -16283 473 -16205 519
rect -16159 473 -16081 519
rect -16035 473 -15957 519
rect -15911 473 -15833 519
rect -15787 473 -15709 519
rect -15663 473 -15585 519
rect -15539 473 -15461 519
rect -15415 473 -15337 519
rect -15291 473 -15213 519
rect -15167 473 -15089 519
rect -15043 473 -14965 519
rect -14919 473 -14841 519
rect -14795 473 -14717 519
rect -14671 473 -14593 519
rect -14547 473 -14469 519
rect -14423 473 -14345 519
rect -14299 473 -14221 519
rect -14175 473 -14097 519
rect -14051 473 -13973 519
rect -13927 473 -13849 519
rect -13803 473 -13725 519
rect -13679 473 -13601 519
rect -13555 473 -13477 519
rect -13431 473 -13353 519
rect -13307 473 -13229 519
rect -13183 473 -13105 519
rect -13059 473 -12981 519
rect -12935 473 -12857 519
rect -12811 473 -12733 519
rect -12687 473 -12609 519
rect -12563 473 -12485 519
rect -12439 473 -12361 519
rect -12315 473 -12237 519
rect -12191 473 -12113 519
rect -12067 473 -11989 519
rect -11943 473 -11865 519
rect -11819 473 -11741 519
rect -11695 473 -11617 519
rect -11571 473 -11493 519
rect -11447 473 -11369 519
rect -11323 473 -11245 519
rect -11199 473 -11121 519
rect -11075 473 -10997 519
rect -10951 473 -10873 519
rect -10827 473 -10749 519
rect -10703 473 -10625 519
rect -10579 473 -10501 519
rect -10455 473 -10377 519
rect -10331 473 -10253 519
rect -10207 473 -10129 519
rect -10083 473 -10005 519
rect -9959 473 -9881 519
rect -9835 473 -9757 519
rect -9711 473 -9633 519
rect -9587 473 -9509 519
rect -9463 473 -9385 519
rect -9339 473 -9261 519
rect -9215 473 -9137 519
rect -9091 473 -9013 519
rect -8967 473 -8889 519
rect -8843 473 -8765 519
rect -8719 473 -8641 519
rect -8595 473 -8517 519
rect -8471 473 -8393 519
rect -8347 473 -8269 519
rect -8223 473 -8145 519
rect -8099 473 -8021 519
rect -7975 473 -7897 519
rect -7851 473 -7773 519
rect -7727 473 -7649 519
rect -7603 473 -7525 519
rect -7479 473 -7401 519
rect -7355 473 -7277 519
rect -7231 473 -7153 519
rect -7107 473 -7029 519
rect -6983 473 -6905 519
rect -6859 473 -6781 519
rect -6735 473 -6657 519
rect -6611 473 -6533 519
rect -6487 473 -6409 519
rect -6363 473 -6285 519
rect -6239 473 -6161 519
rect -6115 473 -6037 519
rect -5991 473 -5913 519
rect -5867 473 -5789 519
rect -5743 473 -5665 519
rect -5619 473 -5541 519
rect -5495 473 -5417 519
rect -5371 473 -5293 519
rect -5247 473 -5169 519
rect -5123 473 -5045 519
rect -4999 473 -4921 519
rect -4875 473 -4797 519
rect -4751 473 -4673 519
rect -4627 473 -4549 519
rect -4503 473 -4425 519
rect -4379 473 -4301 519
rect -4255 473 -4177 519
rect -4131 473 -4053 519
rect -4007 473 -3929 519
rect -3883 473 -3805 519
rect -3759 473 -3681 519
rect -3635 473 -3557 519
rect -3511 473 -3433 519
rect -3387 473 -3309 519
rect -3263 473 -3185 519
rect -3139 473 -3061 519
rect -3015 473 -2937 519
rect -2891 473 -2813 519
rect -2767 473 -2689 519
rect -2643 473 -2565 519
rect -2519 473 -2441 519
rect -2395 473 -2317 519
rect -2271 473 -2193 519
rect -2147 473 -2069 519
rect -2023 473 -1945 519
rect -1899 473 -1821 519
rect -1775 473 -1697 519
rect -1651 473 -1573 519
rect -1527 473 -1449 519
rect -1403 473 -1325 519
rect -1279 473 -1201 519
rect -1155 473 -1077 519
rect -1031 473 -953 519
rect -907 473 -829 519
rect -783 473 -705 519
rect -659 473 -581 519
rect -535 473 -457 519
rect -411 473 -333 519
rect -287 473 -209 519
rect -163 473 -85 519
rect -39 473 39 519
rect 85 473 163 519
rect 209 473 287 519
rect 333 473 411 519
rect 457 473 535 519
rect 581 473 659 519
rect 705 473 783 519
rect 829 473 907 519
rect 953 473 1031 519
rect 1077 473 1155 519
rect 1201 473 1279 519
rect 1325 473 1403 519
rect 1449 473 1527 519
rect 1573 473 1651 519
rect 1697 473 1775 519
rect 1821 473 1899 519
rect 1945 473 2023 519
rect 2069 473 2147 519
rect 2193 473 2271 519
rect 2317 473 2395 519
rect 2441 473 2519 519
rect 2565 473 2643 519
rect 2689 473 2767 519
rect 2813 473 2891 519
rect 2937 473 3015 519
rect 3061 473 3139 519
rect 3185 473 3263 519
rect 3309 473 3387 519
rect 3433 473 3511 519
rect 3557 473 3635 519
rect 3681 473 3759 519
rect 3805 473 3883 519
rect 3929 473 4007 519
rect 4053 473 4131 519
rect 4177 473 4255 519
rect 4301 473 4379 519
rect 4425 473 4503 519
rect 4549 473 4627 519
rect 4673 473 4751 519
rect 4797 473 4875 519
rect 4921 473 4999 519
rect 5045 473 5123 519
rect 5169 473 5247 519
rect 5293 473 5371 519
rect 5417 473 5495 519
rect 5541 473 5619 519
rect 5665 473 5743 519
rect 5789 473 5867 519
rect 5913 473 5991 519
rect 6037 473 6115 519
rect 6161 473 6239 519
rect 6285 473 6363 519
rect 6409 473 6487 519
rect 6533 473 6611 519
rect 6657 473 6735 519
rect 6781 473 6859 519
rect 6905 473 6983 519
rect 7029 473 7107 519
rect 7153 473 7231 519
rect 7277 473 7355 519
rect 7401 473 7479 519
rect 7525 473 7603 519
rect 7649 473 7727 519
rect 7773 473 7851 519
rect 7897 473 7975 519
rect 8021 473 8099 519
rect 8145 473 8223 519
rect 8269 473 8347 519
rect 8393 473 8471 519
rect 8517 473 8595 519
rect 8641 473 8719 519
rect 8765 473 8843 519
rect 8889 473 8967 519
rect 9013 473 9091 519
rect 9137 473 9215 519
rect 9261 473 9339 519
rect 9385 473 9463 519
rect 9509 473 9587 519
rect 9633 473 9711 519
rect 9757 473 9835 519
rect 9881 473 9959 519
rect 10005 473 10083 519
rect 10129 473 10207 519
rect 10253 473 10331 519
rect 10377 473 10455 519
rect 10501 473 10579 519
rect 10625 473 10703 519
rect 10749 473 10827 519
rect 10873 473 10951 519
rect 10997 473 11075 519
rect 11121 473 11199 519
rect 11245 473 11323 519
rect 11369 473 11447 519
rect 11493 473 11571 519
rect 11617 473 11695 519
rect 11741 473 11819 519
rect 11865 473 11943 519
rect 11989 473 12067 519
rect 12113 473 12191 519
rect 12237 473 12315 519
rect 12361 473 12439 519
rect 12485 473 12563 519
rect 12609 473 12687 519
rect 12733 473 12811 519
rect 12857 473 12935 519
rect 12981 473 13059 519
rect 13105 473 13183 519
rect 13229 473 13307 519
rect 13353 473 13431 519
rect 13477 473 13555 519
rect 13601 473 13679 519
rect 13725 473 13803 519
rect 13849 473 13927 519
rect 13973 473 14051 519
rect 14097 473 14175 519
rect 14221 473 14299 519
rect 14345 473 14423 519
rect 14469 473 14547 519
rect 14593 473 14671 519
rect 14717 473 14795 519
rect 14841 473 14919 519
rect 14965 473 15043 519
rect 15089 473 15167 519
rect 15213 473 15291 519
rect 15337 473 15415 519
rect 15461 473 15539 519
rect 15585 473 15663 519
rect 15709 473 15787 519
rect 15833 473 15911 519
rect 15957 473 16035 519
rect 16081 473 16159 519
rect 16205 473 16283 519
rect 16329 473 16407 519
rect 16453 473 16531 519
rect 16577 473 16655 519
rect 16701 473 16779 519
rect 16825 473 16903 519
rect 16949 473 17027 519
rect 17073 473 17151 519
rect 17197 473 17275 519
rect 17321 473 17399 519
rect 17445 473 17523 519
rect 17569 473 17647 519
rect 17693 473 17771 519
rect 17817 473 17895 519
rect 17941 473 18019 519
rect 18065 473 18143 519
rect 18189 473 18267 519
rect 18313 473 18324 519
rect -18324 395 18324 473
rect -18324 349 -18313 395
rect -18267 349 -18189 395
rect -18143 349 -18065 395
rect -18019 349 -17941 395
rect -17895 349 -17817 395
rect -17771 349 -17693 395
rect -17647 349 -17569 395
rect -17523 349 -17445 395
rect -17399 349 -17321 395
rect -17275 349 -17197 395
rect -17151 349 -17073 395
rect -17027 349 -16949 395
rect -16903 349 -16825 395
rect -16779 349 -16701 395
rect -16655 349 -16577 395
rect -16531 349 -16453 395
rect -16407 349 -16329 395
rect -16283 349 -16205 395
rect -16159 349 -16081 395
rect -16035 349 -15957 395
rect -15911 349 -15833 395
rect -15787 349 -15709 395
rect -15663 349 -15585 395
rect -15539 349 -15461 395
rect -15415 349 -15337 395
rect -15291 349 -15213 395
rect -15167 349 -15089 395
rect -15043 349 -14965 395
rect -14919 349 -14841 395
rect -14795 349 -14717 395
rect -14671 349 -14593 395
rect -14547 349 -14469 395
rect -14423 349 -14345 395
rect -14299 349 -14221 395
rect -14175 349 -14097 395
rect -14051 349 -13973 395
rect -13927 349 -13849 395
rect -13803 349 -13725 395
rect -13679 349 -13601 395
rect -13555 349 -13477 395
rect -13431 349 -13353 395
rect -13307 349 -13229 395
rect -13183 349 -13105 395
rect -13059 349 -12981 395
rect -12935 349 -12857 395
rect -12811 349 -12733 395
rect -12687 349 -12609 395
rect -12563 349 -12485 395
rect -12439 349 -12361 395
rect -12315 349 -12237 395
rect -12191 349 -12113 395
rect -12067 349 -11989 395
rect -11943 349 -11865 395
rect -11819 349 -11741 395
rect -11695 349 -11617 395
rect -11571 349 -11493 395
rect -11447 349 -11369 395
rect -11323 349 -11245 395
rect -11199 349 -11121 395
rect -11075 349 -10997 395
rect -10951 349 -10873 395
rect -10827 349 -10749 395
rect -10703 349 -10625 395
rect -10579 349 -10501 395
rect -10455 349 -10377 395
rect -10331 349 -10253 395
rect -10207 349 -10129 395
rect -10083 349 -10005 395
rect -9959 349 -9881 395
rect -9835 349 -9757 395
rect -9711 349 -9633 395
rect -9587 349 -9509 395
rect -9463 349 -9385 395
rect -9339 349 -9261 395
rect -9215 349 -9137 395
rect -9091 349 -9013 395
rect -8967 349 -8889 395
rect -8843 349 -8765 395
rect -8719 349 -8641 395
rect -8595 349 -8517 395
rect -8471 349 -8393 395
rect -8347 349 -8269 395
rect -8223 349 -8145 395
rect -8099 349 -8021 395
rect -7975 349 -7897 395
rect -7851 349 -7773 395
rect -7727 349 -7649 395
rect -7603 349 -7525 395
rect -7479 349 -7401 395
rect -7355 349 -7277 395
rect -7231 349 -7153 395
rect -7107 349 -7029 395
rect -6983 349 -6905 395
rect -6859 349 -6781 395
rect -6735 349 -6657 395
rect -6611 349 -6533 395
rect -6487 349 -6409 395
rect -6363 349 -6285 395
rect -6239 349 -6161 395
rect -6115 349 -6037 395
rect -5991 349 -5913 395
rect -5867 349 -5789 395
rect -5743 349 -5665 395
rect -5619 349 -5541 395
rect -5495 349 -5417 395
rect -5371 349 -5293 395
rect -5247 349 -5169 395
rect -5123 349 -5045 395
rect -4999 349 -4921 395
rect -4875 349 -4797 395
rect -4751 349 -4673 395
rect -4627 349 -4549 395
rect -4503 349 -4425 395
rect -4379 349 -4301 395
rect -4255 349 -4177 395
rect -4131 349 -4053 395
rect -4007 349 -3929 395
rect -3883 349 -3805 395
rect -3759 349 -3681 395
rect -3635 349 -3557 395
rect -3511 349 -3433 395
rect -3387 349 -3309 395
rect -3263 349 -3185 395
rect -3139 349 -3061 395
rect -3015 349 -2937 395
rect -2891 349 -2813 395
rect -2767 349 -2689 395
rect -2643 349 -2565 395
rect -2519 349 -2441 395
rect -2395 349 -2317 395
rect -2271 349 -2193 395
rect -2147 349 -2069 395
rect -2023 349 -1945 395
rect -1899 349 -1821 395
rect -1775 349 -1697 395
rect -1651 349 -1573 395
rect -1527 349 -1449 395
rect -1403 349 -1325 395
rect -1279 349 -1201 395
rect -1155 349 -1077 395
rect -1031 349 -953 395
rect -907 349 -829 395
rect -783 349 -705 395
rect -659 349 -581 395
rect -535 349 -457 395
rect -411 349 -333 395
rect -287 349 -209 395
rect -163 349 -85 395
rect -39 349 39 395
rect 85 349 163 395
rect 209 349 287 395
rect 333 349 411 395
rect 457 349 535 395
rect 581 349 659 395
rect 705 349 783 395
rect 829 349 907 395
rect 953 349 1031 395
rect 1077 349 1155 395
rect 1201 349 1279 395
rect 1325 349 1403 395
rect 1449 349 1527 395
rect 1573 349 1651 395
rect 1697 349 1775 395
rect 1821 349 1899 395
rect 1945 349 2023 395
rect 2069 349 2147 395
rect 2193 349 2271 395
rect 2317 349 2395 395
rect 2441 349 2519 395
rect 2565 349 2643 395
rect 2689 349 2767 395
rect 2813 349 2891 395
rect 2937 349 3015 395
rect 3061 349 3139 395
rect 3185 349 3263 395
rect 3309 349 3387 395
rect 3433 349 3511 395
rect 3557 349 3635 395
rect 3681 349 3759 395
rect 3805 349 3883 395
rect 3929 349 4007 395
rect 4053 349 4131 395
rect 4177 349 4255 395
rect 4301 349 4379 395
rect 4425 349 4503 395
rect 4549 349 4627 395
rect 4673 349 4751 395
rect 4797 349 4875 395
rect 4921 349 4999 395
rect 5045 349 5123 395
rect 5169 349 5247 395
rect 5293 349 5371 395
rect 5417 349 5495 395
rect 5541 349 5619 395
rect 5665 349 5743 395
rect 5789 349 5867 395
rect 5913 349 5991 395
rect 6037 349 6115 395
rect 6161 349 6239 395
rect 6285 349 6363 395
rect 6409 349 6487 395
rect 6533 349 6611 395
rect 6657 349 6735 395
rect 6781 349 6859 395
rect 6905 349 6983 395
rect 7029 349 7107 395
rect 7153 349 7231 395
rect 7277 349 7355 395
rect 7401 349 7479 395
rect 7525 349 7603 395
rect 7649 349 7727 395
rect 7773 349 7851 395
rect 7897 349 7975 395
rect 8021 349 8099 395
rect 8145 349 8223 395
rect 8269 349 8347 395
rect 8393 349 8471 395
rect 8517 349 8595 395
rect 8641 349 8719 395
rect 8765 349 8843 395
rect 8889 349 8967 395
rect 9013 349 9091 395
rect 9137 349 9215 395
rect 9261 349 9339 395
rect 9385 349 9463 395
rect 9509 349 9587 395
rect 9633 349 9711 395
rect 9757 349 9835 395
rect 9881 349 9959 395
rect 10005 349 10083 395
rect 10129 349 10207 395
rect 10253 349 10331 395
rect 10377 349 10455 395
rect 10501 349 10579 395
rect 10625 349 10703 395
rect 10749 349 10827 395
rect 10873 349 10951 395
rect 10997 349 11075 395
rect 11121 349 11199 395
rect 11245 349 11323 395
rect 11369 349 11447 395
rect 11493 349 11571 395
rect 11617 349 11695 395
rect 11741 349 11819 395
rect 11865 349 11943 395
rect 11989 349 12067 395
rect 12113 349 12191 395
rect 12237 349 12315 395
rect 12361 349 12439 395
rect 12485 349 12563 395
rect 12609 349 12687 395
rect 12733 349 12811 395
rect 12857 349 12935 395
rect 12981 349 13059 395
rect 13105 349 13183 395
rect 13229 349 13307 395
rect 13353 349 13431 395
rect 13477 349 13555 395
rect 13601 349 13679 395
rect 13725 349 13803 395
rect 13849 349 13927 395
rect 13973 349 14051 395
rect 14097 349 14175 395
rect 14221 349 14299 395
rect 14345 349 14423 395
rect 14469 349 14547 395
rect 14593 349 14671 395
rect 14717 349 14795 395
rect 14841 349 14919 395
rect 14965 349 15043 395
rect 15089 349 15167 395
rect 15213 349 15291 395
rect 15337 349 15415 395
rect 15461 349 15539 395
rect 15585 349 15663 395
rect 15709 349 15787 395
rect 15833 349 15911 395
rect 15957 349 16035 395
rect 16081 349 16159 395
rect 16205 349 16283 395
rect 16329 349 16407 395
rect 16453 349 16531 395
rect 16577 349 16655 395
rect 16701 349 16779 395
rect 16825 349 16903 395
rect 16949 349 17027 395
rect 17073 349 17151 395
rect 17197 349 17275 395
rect 17321 349 17399 395
rect 17445 349 17523 395
rect 17569 349 17647 395
rect 17693 349 17771 395
rect 17817 349 17895 395
rect 17941 349 18019 395
rect 18065 349 18143 395
rect 18189 349 18267 395
rect 18313 349 18324 395
rect -18324 271 18324 349
rect -18324 225 -18313 271
rect -18267 225 -18189 271
rect -18143 225 -18065 271
rect -18019 225 -17941 271
rect -17895 225 -17817 271
rect -17771 225 -17693 271
rect -17647 225 -17569 271
rect -17523 225 -17445 271
rect -17399 225 -17321 271
rect -17275 225 -17197 271
rect -17151 225 -17073 271
rect -17027 225 -16949 271
rect -16903 225 -16825 271
rect -16779 225 -16701 271
rect -16655 225 -16577 271
rect -16531 225 -16453 271
rect -16407 225 -16329 271
rect -16283 225 -16205 271
rect -16159 225 -16081 271
rect -16035 225 -15957 271
rect -15911 225 -15833 271
rect -15787 225 -15709 271
rect -15663 225 -15585 271
rect -15539 225 -15461 271
rect -15415 225 -15337 271
rect -15291 225 -15213 271
rect -15167 225 -15089 271
rect -15043 225 -14965 271
rect -14919 225 -14841 271
rect -14795 225 -14717 271
rect -14671 225 -14593 271
rect -14547 225 -14469 271
rect -14423 225 -14345 271
rect -14299 225 -14221 271
rect -14175 225 -14097 271
rect -14051 225 -13973 271
rect -13927 225 -13849 271
rect -13803 225 -13725 271
rect -13679 225 -13601 271
rect -13555 225 -13477 271
rect -13431 225 -13353 271
rect -13307 225 -13229 271
rect -13183 225 -13105 271
rect -13059 225 -12981 271
rect -12935 225 -12857 271
rect -12811 225 -12733 271
rect -12687 225 -12609 271
rect -12563 225 -12485 271
rect -12439 225 -12361 271
rect -12315 225 -12237 271
rect -12191 225 -12113 271
rect -12067 225 -11989 271
rect -11943 225 -11865 271
rect -11819 225 -11741 271
rect -11695 225 -11617 271
rect -11571 225 -11493 271
rect -11447 225 -11369 271
rect -11323 225 -11245 271
rect -11199 225 -11121 271
rect -11075 225 -10997 271
rect -10951 225 -10873 271
rect -10827 225 -10749 271
rect -10703 225 -10625 271
rect -10579 225 -10501 271
rect -10455 225 -10377 271
rect -10331 225 -10253 271
rect -10207 225 -10129 271
rect -10083 225 -10005 271
rect -9959 225 -9881 271
rect -9835 225 -9757 271
rect -9711 225 -9633 271
rect -9587 225 -9509 271
rect -9463 225 -9385 271
rect -9339 225 -9261 271
rect -9215 225 -9137 271
rect -9091 225 -9013 271
rect -8967 225 -8889 271
rect -8843 225 -8765 271
rect -8719 225 -8641 271
rect -8595 225 -8517 271
rect -8471 225 -8393 271
rect -8347 225 -8269 271
rect -8223 225 -8145 271
rect -8099 225 -8021 271
rect -7975 225 -7897 271
rect -7851 225 -7773 271
rect -7727 225 -7649 271
rect -7603 225 -7525 271
rect -7479 225 -7401 271
rect -7355 225 -7277 271
rect -7231 225 -7153 271
rect -7107 225 -7029 271
rect -6983 225 -6905 271
rect -6859 225 -6781 271
rect -6735 225 -6657 271
rect -6611 225 -6533 271
rect -6487 225 -6409 271
rect -6363 225 -6285 271
rect -6239 225 -6161 271
rect -6115 225 -6037 271
rect -5991 225 -5913 271
rect -5867 225 -5789 271
rect -5743 225 -5665 271
rect -5619 225 -5541 271
rect -5495 225 -5417 271
rect -5371 225 -5293 271
rect -5247 225 -5169 271
rect -5123 225 -5045 271
rect -4999 225 -4921 271
rect -4875 225 -4797 271
rect -4751 225 -4673 271
rect -4627 225 -4549 271
rect -4503 225 -4425 271
rect -4379 225 -4301 271
rect -4255 225 -4177 271
rect -4131 225 -4053 271
rect -4007 225 -3929 271
rect -3883 225 -3805 271
rect -3759 225 -3681 271
rect -3635 225 -3557 271
rect -3511 225 -3433 271
rect -3387 225 -3309 271
rect -3263 225 -3185 271
rect -3139 225 -3061 271
rect -3015 225 -2937 271
rect -2891 225 -2813 271
rect -2767 225 -2689 271
rect -2643 225 -2565 271
rect -2519 225 -2441 271
rect -2395 225 -2317 271
rect -2271 225 -2193 271
rect -2147 225 -2069 271
rect -2023 225 -1945 271
rect -1899 225 -1821 271
rect -1775 225 -1697 271
rect -1651 225 -1573 271
rect -1527 225 -1449 271
rect -1403 225 -1325 271
rect -1279 225 -1201 271
rect -1155 225 -1077 271
rect -1031 225 -953 271
rect -907 225 -829 271
rect -783 225 -705 271
rect -659 225 -581 271
rect -535 225 -457 271
rect -411 225 -333 271
rect -287 225 -209 271
rect -163 225 -85 271
rect -39 225 39 271
rect 85 225 163 271
rect 209 225 287 271
rect 333 225 411 271
rect 457 225 535 271
rect 581 225 659 271
rect 705 225 783 271
rect 829 225 907 271
rect 953 225 1031 271
rect 1077 225 1155 271
rect 1201 225 1279 271
rect 1325 225 1403 271
rect 1449 225 1527 271
rect 1573 225 1651 271
rect 1697 225 1775 271
rect 1821 225 1899 271
rect 1945 225 2023 271
rect 2069 225 2147 271
rect 2193 225 2271 271
rect 2317 225 2395 271
rect 2441 225 2519 271
rect 2565 225 2643 271
rect 2689 225 2767 271
rect 2813 225 2891 271
rect 2937 225 3015 271
rect 3061 225 3139 271
rect 3185 225 3263 271
rect 3309 225 3387 271
rect 3433 225 3511 271
rect 3557 225 3635 271
rect 3681 225 3759 271
rect 3805 225 3883 271
rect 3929 225 4007 271
rect 4053 225 4131 271
rect 4177 225 4255 271
rect 4301 225 4379 271
rect 4425 225 4503 271
rect 4549 225 4627 271
rect 4673 225 4751 271
rect 4797 225 4875 271
rect 4921 225 4999 271
rect 5045 225 5123 271
rect 5169 225 5247 271
rect 5293 225 5371 271
rect 5417 225 5495 271
rect 5541 225 5619 271
rect 5665 225 5743 271
rect 5789 225 5867 271
rect 5913 225 5991 271
rect 6037 225 6115 271
rect 6161 225 6239 271
rect 6285 225 6363 271
rect 6409 225 6487 271
rect 6533 225 6611 271
rect 6657 225 6735 271
rect 6781 225 6859 271
rect 6905 225 6983 271
rect 7029 225 7107 271
rect 7153 225 7231 271
rect 7277 225 7355 271
rect 7401 225 7479 271
rect 7525 225 7603 271
rect 7649 225 7727 271
rect 7773 225 7851 271
rect 7897 225 7975 271
rect 8021 225 8099 271
rect 8145 225 8223 271
rect 8269 225 8347 271
rect 8393 225 8471 271
rect 8517 225 8595 271
rect 8641 225 8719 271
rect 8765 225 8843 271
rect 8889 225 8967 271
rect 9013 225 9091 271
rect 9137 225 9215 271
rect 9261 225 9339 271
rect 9385 225 9463 271
rect 9509 225 9587 271
rect 9633 225 9711 271
rect 9757 225 9835 271
rect 9881 225 9959 271
rect 10005 225 10083 271
rect 10129 225 10207 271
rect 10253 225 10331 271
rect 10377 225 10455 271
rect 10501 225 10579 271
rect 10625 225 10703 271
rect 10749 225 10827 271
rect 10873 225 10951 271
rect 10997 225 11075 271
rect 11121 225 11199 271
rect 11245 225 11323 271
rect 11369 225 11447 271
rect 11493 225 11571 271
rect 11617 225 11695 271
rect 11741 225 11819 271
rect 11865 225 11943 271
rect 11989 225 12067 271
rect 12113 225 12191 271
rect 12237 225 12315 271
rect 12361 225 12439 271
rect 12485 225 12563 271
rect 12609 225 12687 271
rect 12733 225 12811 271
rect 12857 225 12935 271
rect 12981 225 13059 271
rect 13105 225 13183 271
rect 13229 225 13307 271
rect 13353 225 13431 271
rect 13477 225 13555 271
rect 13601 225 13679 271
rect 13725 225 13803 271
rect 13849 225 13927 271
rect 13973 225 14051 271
rect 14097 225 14175 271
rect 14221 225 14299 271
rect 14345 225 14423 271
rect 14469 225 14547 271
rect 14593 225 14671 271
rect 14717 225 14795 271
rect 14841 225 14919 271
rect 14965 225 15043 271
rect 15089 225 15167 271
rect 15213 225 15291 271
rect 15337 225 15415 271
rect 15461 225 15539 271
rect 15585 225 15663 271
rect 15709 225 15787 271
rect 15833 225 15911 271
rect 15957 225 16035 271
rect 16081 225 16159 271
rect 16205 225 16283 271
rect 16329 225 16407 271
rect 16453 225 16531 271
rect 16577 225 16655 271
rect 16701 225 16779 271
rect 16825 225 16903 271
rect 16949 225 17027 271
rect 17073 225 17151 271
rect 17197 225 17275 271
rect 17321 225 17399 271
rect 17445 225 17523 271
rect 17569 225 17647 271
rect 17693 225 17771 271
rect 17817 225 17895 271
rect 17941 225 18019 271
rect 18065 225 18143 271
rect 18189 225 18267 271
rect 18313 225 18324 271
rect -18324 147 18324 225
rect -18324 101 -18313 147
rect -18267 101 -18189 147
rect -18143 101 -18065 147
rect -18019 101 -17941 147
rect -17895 101 -17817 147
rect -17771 101 -17693 147
rect -17647 101 -17569 147
rect -17523 101 -17445 147
rect -17399 101 -17321 147
rect -17275 101 -17197 147
rect -17151 101 -17073 147
rect -17027 101 -16949 147
rect -16903 101 -16825 147
rect -16779 101 -16701 147
rect -16655 101 -16577 147
rect -16531 101 -16453 147
rect -16407 101 -16329 147
rect -16283 101 -16205 147
rect -16159 101 -16081 147
rect -16035 101 -15957 147
rect -15911 101 -15833 147
rect -15787 101 -15709 147
rect -15663 101 -15585 147
rect -15539 101 -15461 147
rect -15415 101 -15337 147
rect -15291 101 -15213 147
rect -15167 101 -15089 147
rect -15043 101 -14965 147
rect -14919 101 -14841 147
rect -14795 101 -14717 147
rect -14671 101 -14593 147
rect -14547 101 -14469 147
rect -14423 101 -14345 147
rect -14299 101 -14221 147
rect -14175 101 -14097 147
rect -14051 101 -13973 147
rect -13927 101 -13849 147
rect -13803 101 -13725 147
rect -13679 101 -13601 147
rect -13555 101 -13477 147
rect -13431 101 -13353 147
rect -13307 101 -13229 147
rect -13183 101 -13105 147
rect -13059 101 -12981 147
rect -12935 101 -12857 147
rect -12811 101 -12733 147
rect -12687 101 -12609 147
rect -12563 101 -12485 147
rect -12439 101 -12361 147
rect -12315 101 -12237 147
rect -12191 101 -12113 147
rect -12067 101 -11989 147
rect -11943 101 -11865 147
rect -11819 101 -11741 147
rect -11695 101 -11617 147
rect -11571 101 -11493 147
rect -11447 101 -11369 147
rect -11323 101 -11245 147
rect -11199 101 -11121 147
rect -11075 101 -10997 147
rect -10951 101 -10873 147
rect -10827 101 -10749 147
rect -10703 101 -10625 147
rect -10579 101 -10501 147
rect -10455 101 -10377 147
rect -10331 101 -10253 147
rect -10207 101 -10129 147
rect -10083 101 -10005 147
rect -9959 101 -9881 147
rect -9835 101 -9757 147
rect -9711 101 -9633 147
rect -9587 101 -9509 147
rect -9463 101 -9385 147
rect -9339 101 -9261 147
rect -9215 101 -9137 147
rect -9091 101 -9013 147
rect -8967 101 -8889 147
rect -8843 101 -8765 147
rect -8719 101 -8641 147
rect -8595 101 -8517 147
rect -8471 101 -8393 147
rect -8347 101 -8269 147
rect -8223 101 -8145 147
rect -8099 101 -8021 147
rect -7975 101 -7897 147
rect -7851 101 -7773 147
rect -7727 101 -7649 147
rect -7603 101 -7525 147
rect -7479 101 -7401 147
rect -7355 101 -7277 147
rect -7231 101 -7153 147
rect -7107 101 -7029 147
rect -6983 101 -6905 147
rect -6859 101 -6781 147
rect -6735 101 -6657 147
rect -6611 101 -6533 147
rect -6487 101 -6409 147
rect -6363 101 -6285 147
rect -6239 101 -6161 147
rect -6115 101 -6037 147
rect -5991 101 -5913 147
rect -5867 101 -5789 147
rect -5743 101 -5665 147
rect -5619 101 -5541 147
rect -5495 101 -5417 147
rect -5371 101 -5293 147
rect -5247 101 -5169 147
rect -5123 101 -5045 147
rect -4999 101 -4921 147
rect -4875 101 -4797 147
rect -4751 101 -4673 147
rect -4627 101 -4549 147
rect -4503 101 -4425 147
rect -4379 101 -4301 147
rect -4255 101 -4177 147
rect -4131 101 -4053 147
rect -4007 101 -3929 147
rect -3883 101 -3805 147
rect -3759 101 -3681 147
rect -3635 101 -3557 147
rect -3511 101 -3433 147
rect -3387 101 -3309 147
rect -3263 101 -3185 147
rect -3139 101 -3061 147
rect -3015 101 -2937 147
rect -2891 101 -2813 147
rect -2767 101 -2689 147
rect -2643 101 -2565 147
rect -2519 101 -2441 147
rect -2395 101 -2317 147
rect -2271 101 -2193 147
rect -2147 101 -2069 147
rect -2023 101 -1945 147
rect -1899 101 -1821 147
rect -1775 101 -1697 147
rect -1651 101 -1573 147
rect -1527 101 -1449 147
rect -1403 101 -1325 147
rect -1279 101 -1201 147
rect -1155 101 -1077 147
rect -1031 101 -953 147
rect -907 101 -829 147
rect -783 101 -705 147
rect -659 101 -581 147
rect -535 101 -457 147
rect -411 101 -333 147
rect -287 101 -209 147
rect -163 101 -85 147
rect -39 101 39 147
rect 85 101 163 147
rect 209 101 287 147
rect 333 101 411 147
rect 457 101 535 147
rect 581 101 659 147
rect 705 101 783 147
rect 829 101 907 147
rect 953 101 1031 147
rect 1077 101 1155 147
rect 1201 101 1279 147
rect 1325 101 1403 147
rect 1449 101 1527 147
rect 1573 101 1651 147
rect 1697 101 1775 147
rect 1821 101 1899 147
rect 1945 101 2023 147
rect 2069 101 2147 147
rect 2193 101 2271 147
rect 2317 101 2395 147
rect 2441 101 2519 147
rect 2565 101 2643 147
rect 2689 101 2767 147
rect 2813 101 2891 147
rect 2937 101 3015 147
rect 3061 101 3139 147
rect 3185 101 3263 147
rect 3309 101 3387 147
rect 3433 101 3511 147
rect 3557 101 3635 147
rect 3681 101 3759 147
rect 3805 101 3883 147
rect 3929 101 4007 147
rect 4053 101 4131 147
rect 4177 101 4255 147
rect 4301 101 4379 147
rect 4425 101 4503 147
rect 4549 101 4627 147
rect 4673 101 4751 147
rect 4797 101 4875 147
rect 4921 101 4999 147
rect 5045 101 5123 147
rect 5169 101 5247 147
rect 5293 101 5371 147
rect 5417 101 5495 147
rect 5541 101 5619 147
rect 5665 101 5743 147
rect 5789 101 5867 147
rect 5913 101 5991 147
rect 6037 101 6115 147
rect 6161 101 6239 147
rect 6285 101 6363 147
rect 6409 101 6487 147
rect 6533 101 6611 147
rect 6657 101 6735 147
rect 6781 101 6859 147
rect 6905 101 6983 147
rect 7029 101 7107 147
rect 7153 101 7231 147
rect 7277 101 7355 147
rect 7401 101 7479 147
rect 7525 101 7603 147
rect 7649 101 7727 147
rect 7773 101 7851 147
rect 7897 101 7975 147
rect 8021 101 8099 147
rect 8145 101 8223 147
rect 8269 101 8347 147
rect 8393 101 8471 147
rect 8517 101 8595 147
rect 8641 101 8719 147
rect 8765 101 8843 147
rect 8889 101 8967 147
rect 9013 101 9091 147
rect 9137 101 9215 147
rect 9261 101 9339 147
rect 9385 101 9463 147
rect 9509 101 9587 147
rect 9633 101 9711 147
rect 9757 101 9835 147
rect 9881 101 9959 147
rect 10005 101 10083 147
rect 10129 101 10207 147
rect 10253 101 10331 147
rect 10377 101 10455 147
rect 10501 101 10579 147
rect 10625 101 10703 147
rect 10749 101 10827 147
rect 10873 101 10951 147
rect 10997 101 11075 147
rect 11121 101 11199 147
rect 11245 101 11323 147
rect 11369 101 11447 147
rect 11493 101 11571 147
rect 11617 101 11695 147
rect 11741 101 11819 147
rect 11865 101 11943 147
rect 11989 101 12067 147
rect 12113 101 12191 147
rect 12237 101 12315 147
rect 12361 101 12439 147
rect 12485 101 12563 147
rect 12609 101 12687 147
rect 12733 101 12811 147
rect 12857 101 12935 147
rect 12981 101 13059 147
rect 13105 101 13183 147
rect 13229 101 13307 147
rect 13353 101 13431 147
rect 13477 101 13555 147
rect 13601 101 13679 147
rect 13725 101 13803 147
rect 13849 101 13927 147
rect 13973 101 14051 147
rect 14097 101 14175 147
rect 14221 101 14299 147
rect 14345 101 14423 147
rect 14469 101 14547 147
rect 14593 101 14671 147
rect 14717 101 14795 147
rect 14841 101 14919 147
rect 14965 101 15043 147
rect 15089 101 15167 147
rect 15213 101 15291 147
rect 15337 101 15415 147
rect 15461 101 15539 147
rect 15585 101 15663 147
rect 15709 101 15787 147
rect 15833 101 15911 147
rect 15957 101 16035 147
rect 16081 101 16159 147
rect 16205 101 16283 147
rect 16329 101 16407 147
rect 16453 101 16531 147
rect 16577 101 16655 147
rect 16701 101 16779 147
rect 16825 101 16903 147
rect 16949 101 17027 147
rect 17073 101 17151 147
rect 17197 101 17275 147
rect 17321 101 17399 147
rect 17445 101 17523 147
rect 17569 101 17647 147
rect 17693 101 17771 147
rect 17817 101 17895 147
rect 17941 101 18019 147
rect 18065 101 18143 147
rect 18189 101 18267 147
rect 18313 101 18324 147
rect -18324 23 18324 101
rect -18324 -23 -18313 23
rect -18267 -23 -18189 23
rect -18143 -23 -18065 23
rect -18019 -23 -17941 23
rect -17895 -23 -17817 23
rect -17771 -23 -17693 23
rect -17647 -23 -17569 23
rect -17523 -23 -17445 23
rect -17399 -23 -17321 23
rect -17275 -23 -17197 23
rect -17151 -23 -17073 23
rect -17027 -23 -16949 23
rect -16903 -23 -16825 23
rect -16779 -23 -16701 23
rect -16655 -23 -16577 23
rect -16531 -23 -16453 23
rect -16407 -23 -16329 23
rect -16283 -23 -16205 23
rect -16159 -23 -16081 23
rect -16035 -23 -15957 23
rect -15911 -23 -15833 23
rect -15787 -23 -15709 23
rect -15663 -23 -15585 23
rect -15539 -23 -15461 23
rect -15415 -23 -15337 23
rect -15291 -23 -15213 23
rect -15167 -23 -15089 23
rect -15043 -23 -14965 23
rect -14919 -23 -14841 23
rect -14795 -23 -14717 23
rect -14671 -23 -14593 23
rect -14547 -23 -14469 23
rect -14423 -23 -14345 23
rect -14299 -23 -14221 23
rect -14175 -23 -14097 23
rect -14051 -23 -13973 23
rect -13927 -23 -13849 23
rect -13803 -23 -13725 23
rect -13679 -23 -13601 23
rect -13555 -23 -13477 23
rect -13431 -23 -13353 23
rect -13307 -23 -13229 23
rect -13183 -23 -13105 23
rect -13059 -23 -12981 23
rect -12935 -23 -12857 23
rect -12811 -23 -12733 23
rect -12687 -23 -12609 23
rect -12563 -23 -12485 23
rect -12439 -23 -12361 23
rect -12315 -23 -12237 23
rect -12191 -23 -12113 23
rect -12067 -23 -11989 23
rect -11943 -23 -11865 23
rect -11819 -23 -11741 23
rect -11695 -23 -11617 23
rect -11571 -23 -11493 23
rect -11447 -23 -11369 23
rect -11323 -23 -11245 23
rect -11199 -23 -11121 23
rect -11075 -23 -10997 23
rect -10951 -23 -10873 23
rect -10827 -23 -10749 23
rect -10703 -23 -10625 23
rect -10579 -23 -10501 23
rect -10455 -23 -10377 23
rect -10331 -23 -10253 23
rect -10207 -23 -10129 23
rect -10083 -23 -10005 23
rect -9959 -23 -9881 23
rect -9835 -23 -9757 23
rect -9711 -23 -9633 23
rect -9587 -23 -9509 23
rect -9463 -23 -9385 23
rect -9339 -23 -9261 23
rect -9215 -23 -9137 23
rect -9091 -23 -9013 23
rect -8967 -23 -8889 23
rect -8843 -23 -8765 23
rect -8719 -23 -8641 23
rect -8595 -23 -8517 23
rect -8471 -23 -8393 23
rect -8347 -23 -8269 23
rect -8223 -23 -8145 23
rect -8099 -23 -8021 23
rect -7975 -23 -7897 23
rect -7851 -23 -7773 23
rect -7727 -23 -7649 23
rect -7603 -23 -7525 23
rect -7479 -23 -7401 23
rect -7355 -23 -7277 23
rect -7231 -23 -7153 23
rect -7107 -23 -7029 23
rect -6983 -23 -6905 23
rect -6859 -23 -6781 23
rect -6735 -23 -6657 23
rect -6611 -23 -6533 23
rect -6487 -23 -6409 23
rect -6363 -23 -6285 23
rect -6239 -23 -6161 23
rect -6115 -23 -6037 23
rect -5991 -23 -5913 23
rect -5867 -23 -5789 23
rect -5743 -23 -5665 23
rect -5619 -23 -5541 23
rect -5495 -23 -5417 23
rect -5371 -23 -5293 23
rect -5247 -23 -5169 23
rect -5123 -23 -5045 23
rect -4999 -23 -4921 23
rect -4875 -23 -4797 23
rect -4751 -23 -4673 23
rect -4627 -23 -4549 23
rect -4503 -23 -4425 23
rect -4379 -23 -4301 23
rect -4255 -23 -4177 23
rect -4131 -23 -4053 23
rect -4007 -23 -3929 23
rect -3883 -23 -3805 23
rect -3759 -23 -3681 23
rect -3635 -23 -3557 23
rect -3511 -23 -3433 23
rect -3387 -23 -3309 23
rect -3263 -23 -3185 23
rect -3139 -23 -3061 23
rect -3015 -23 -2937 23
rect -2891 -23 -2813 23
rect -2767 -23 -2689 23
rect -2643 -23 -2565 23
rect -2519 -23 -2441 23
rect -2395 -23 -2317 23
rect -2271 -23 -2193 23
rect -2147 -23 -2069 23
rect -2023 -23 -1945 23
rect -1899 -23 -1821 23
rect -1775 -23 -1697 23
rect -1651 -23 -1573 23
rect -1527 -23 -1449 23
rect -1403 -23 -1325 23
rect -1279 -23 -1201 23
rect -1155 -23 -1077 23
rect -1031 -23 -953 23
rect -907 -23 -829 23
rect -783 -23 -705 23
rect -659 -23 -581 23
rect -535 -23 -457 23
rect -411 -23 -333 23
rect -287 -23 -209 23
rect -163 -23 -85 23
rect -39 -23 39 23
rect 85 -23 163 23
rect 209 -23 287 23
rect 333 -23 411 23
rect 457 -23 535 23
rect 581 -23 659 23
rect 705 -23 783 23
rect 829 -23 907 23
rect 953 -23 1031 23
rect 1077 -23 1155 23
rect 1201 -23 1279 23
rect 1325 -23 1403 23
rect 1449 -23 1527 23
rect 1573 -23 1651 23
rect 1697 -23 1775 23
rect 1821 -23 1899 23
rect 1945 -23 2023 23
rect 2069 -23 2147 23
rect 2193 -23 2271 23
rect 2317 -23 2395 23
rect 2441 -23 2519 23
rect 2565 -23 2643 23
rect 2689 -23 2767 23
rect 2813 -23 2891 23
rect 2937 -23 3015 23
rect 3061 -23 3139 23
rect 3185 -23 3263 23
rect 3309 -23 3387 23
rect 3433 -23 3511 23
rect 3557 -23 3635 23
rect 3681 -23 3759 23
rect 3805 -23 3883 23
rect 3929 -23 4007 23
rect 4053 -23 4131 23
rect 4177 -23 4255 23
rect 4301 -23 4379 23
rect 4425 -23 4503 23
rect 4549 -23 4627 23
rect 4673 -23 4751 23
rect 4797 -23 4875 23
rect 4921 -23 4999 23
rect 5045 -23 5123 23
rect 5169 -23 5247 23
rect 5293 -23 5371 23
rect 5417 -23 5495 23
rect 5541 -23 5619 23
rect 5665 -23 5743 23
rect 5789 -23 5867 23
rect 5913 -23 5991 23
rect 6037 -23 6115 23
rect 6161 -23 6239 23
rect 6285 -23 6363 23
rect 6409 -23 6487 23
rect 6533 -23 6611 23
rect 6657 -23 6735 23
rect 6781 -23 6859 23
rect 6905 -23 6983 23
rect 7029 -23 7107 23
rect 7153 -23 7231 23
rect 7277 -23 7355 23
rect 7401 -23 7479 23
rect 7525 -23 7603 23
rect 7649 -23 7727 23
rect 7773 -23 7851 23
rect 7897 -23 7975 23
rect 8021 -23 8099 23
rect 8145 -23 8223 23
rect 8269 -23 8347 23
rect 8393 -23 8471 23
rect 8517 -23 8595 23
rect 8641 -23 8719 23
rect 8765 -23 8843 23
rect 8889 -23 8967 23
rect 9013 -23 9091 23
rect 9137 -23 9215 23
rect 9261 -23 9339 23
rect 9385 -23 9463 23
rect 9509 -23 9587 23
rect 9633 -23 9711 23
rect 9757 -23 9835 23
rect 9881 -23 9959 23
rect 10005 -23 10083 23
rect 10129 -23 10207 23
rect 10253 -23 10331 23
rect 10377 -23 10455 23
rect 10501 -23 10579 23
rect 10625 -23 10703 23
rect 10749 -23 10827 23
rect 10873 -23 10951 23
rect 10997 -23 11075 23
rect 11121 -23 11199 23
rect 11245 -23 11323 23
rect 11369 -23 11447 23
rect 11493 -23 11571 23
rect 11617 -23 11695 23
rect 11741 -23 11819 23
rect 11865 -23 11943 23
rect 11989 -23 12067 23
rect 12113 -23 12191 23
rect 12237 -23 12315 23
rect 12361 -23 12439 23
rect 12485 -23 12563 23
rect 12609 -23 12687 23
rect 12733 -23 12811 23
rect 12857 -23 12935 23
rect 12981 -23 13059 23
rect 13105 -23 13183 23
rect 13229 -23 13307 23
rect 13353 -23 13431 23
rect 13477 -23 13555 23
rect 13601 -23 13679 23
rect 13725 -23 13803 23
rect 13849 -23 13927 23
rect 13973 -23 14051 23
rect 14097 -23 14175 23
rect 14221 -23 14299 23
rect 14345 -23 14423 23
rect 14469 -23 14547 23
rect 14593 -23 14671 23
rect 14717 -23 14795 23
rect 14841 -23 14919 23
rect 14965 -23 15043 23
rect 15089 -23 15167 23
rect 15213 -23 15291 23
rect 15337 -23 15415 23
rect 15461 -23 15539 23
rect 15585 -23 15663 23
rect 15709 -23 15787 23
rect 15833 -23 15911 23
rect 15957 -23 16035 23
rect 16081 -23 16159 23
rect 16205 -23 16283 23
rect 16329 -23 16407 23
rect 16453 -23 16531 23
rect 16577 -23 16655 23
rect 16701 -23 16779 23
rect 16825 -23 16903 23
rect 16949 -23 17027 23
rect 17073 -23 17151 23
rect 17197 -23 17275 23
rect 17321 -23 17399 23
rect 17445 -23 17523 23
rect 17569 -23 17647 23
rect 17693 -23 17771 23
rect 17817 -23 17895 23
rect 17941 -23 18019 23
rect 18065 -23 18143 23
rect 18189 -23 18267 23
rect 18313 -23 18324 23
rect -18324 -101 18324 -23
rect -18324 -147 -18313 -101
rect -18267 -147 -18189 -101
rect -18143 -147 -18065 -101
rect -18019 -147 -17941 -101
rect -17895 -147 -17817 -101
rect -17771 -147 -17693 -101
rect -17647 -147 -17569 -101
rect -17523 -147 -17445 -101
rect -17399 -147 -17321 -101
rect -17275 -147 -17197 -101
rect -17151 -147 -17073 -101
rect -17027 -147 -16949 -101
rect -16903 -147 -16825 -101
rect -16779 -147 -16701 -101
rect -16655 -147 -16577 -101
rect -16531 -147 -16453 -101
rect -16407 -147 -16329 -101
rect -16283 -147 -16205 -101
rect -16159 -147 -16081 -101
rect -16035 -147 -15957 -101
rect -15911 -147 -15833 -101
rect -15787 -147 -15709 -101
rect -15663 -147 -15585 -101
rect -15539 -147 -15461 -101
rect -15415 -147 -15337 -101
rect -15291 -147 -15213 -101
rect -15167 -147 -15089 -101
rect -15043 -147 -14965 -101
rect -14919 -147 -14841 -101
rect -14795 -147 -14717 -101
rect -14671 -147 -14593 -101
rect -14547 -147 -14469 -101
rect -14423 -147 -14345 -101
rect -14299 -147 -14221 -101
rect -14175 -147 -14097 -101
rect -14051 -147 -13973 -101
rect -13927 -147 -13849 -101
rect -13803 -147 -13725 -101
rect -13679 -147 -13601 -101
rect -13555 -147 -13477 -101
rect -13431 -147 -13353 -101
rect -13307 -147 -13229 -101
rect -13183 -147 -13105 -101
rect -13059 -147 -12981 -101
rect -12935 -147 -12857 -101
rect -12811 -147 -12733 -101
rect -12687 -147 -12609 -101
rect -12563 -147 -12485 -101
rect -12439 -147 -12361 -101
rect -12315 -147 -12237 -101
rect -12191 -147 -12113 -101
rect -12067 -147 -11989 -101
rect -11943 -147 -11865 -101
rect -11819 -147 -11741 -101
rect -11695 -147 -11617 -101
rect -11571 -147 -11493 -101
rect -11447 -147 -11369 -101
rect -11323 -147 -11245 -101
rect -11199 -147 -11121 -101
rect -11075 -147 -10997 -101
rect -10951 -147 -10873 -101
rect -10827 -147 -10749 -101
rect -10703 -147 -10625 -101
rect -10579 -147 -10501 -101
rect -10455 -147 -10377 -101
rect -10331 -147 -10253 -101
rect -10207 -147 -10129 -101
rect -10083 -147 -10005 -101
rect -9959 -147 -9881 -101
rect -9835 -147 -9757 -101
rect -9711 -147 -9633 -101
rect -9587 -147 -9509 -101
rect -9463 -147 -9385 -101
rect -9339 -147 -9261 -101
rect -9215 -147 -9137 -101
rect -9091 -147 -9013 -101
rect -8967 -147 -8889 -101
rect -8843 -147 -8765 -101
rect -8719 -147 -8641 -101
rect -8595 -147 -8517 -101
rect -8471 -147 -8393 -101
rect -8347 -147 -8269 -101
rect -8223 -147 -8145 -101
rect -8099 -147 -8021 -101
rect -7975 -147 -7897 -101
rect -7851 -147 -7773 -101
rect -7727 -147 -7649 -101
rect -7603 -147 -7525 -101
rect -7479 -147 -7401 -101
rect -7355 -147 -7277 -101
rect -7231 -147 -7153 -101
rect -7107 -147 -7029 -101
rect -6983 -147 -6905 -101
rect -6859 -147 -6781 -101
rect -6735 -147 -6657 -101
rect -6611 -147 -6533 -101
rect -6487 -147 -6409 -101
rect -6363 -147 -6285 -101
rect -6239 -147 -6161 -101
rect -6115 -147 -6037 -101
rect -5991 -147 -5913 -101
rect -5867 -147 -5789 -101
rect -5743 -147 -5665 -101
rect -5619 -147 -5541 -101
rect -5495 -147 -5417 -101
rect -5371 -147 -5293 -101
rect -5247 -147 -5169 -101
rect -5123 -147 -5045 -101
rect -4999 -147 -4921 -101
rect -4875 -147 -4797 -101
rect -4751 -147 -4673 -101
rect -4627 -147 -4549 -101
rect -4503 -147 -4425 -101
rect -4379 -147 -4301 -101
rect -4255 -147 -4177 -101
rect -4131 -147 -4053 -101
rect -4007 -147 -3929 -101
rect -3883 -147 -3805 -101
rect -3759 -147 -3681 -101
rect -3635 -147 -3557 -101
rect -3511 -147 -3433 -101
rect -3387 -147 -3309 -101
rect -3263 -147 -3185 -101
rect -3139 -147 -3061 -101
rect -3015 -147 -2937 -101
rect -2891 -147 -2813 -101
rect -2767 -147 -2689 -101
rect -2643 -147 -2565 -101
rect -2519 -147 -2441 -101
rect -2395 -147 -2317 -101
rect -2271 -147 -2193 -101
rect -2147 -147 -2069 -101
rect -2023 -147 -1945 -101
rect -1899 -147 -1821 -101
rect -1775 -147 -1697 -101
rect -1651 -147 -1573 -101
rect -1527 -147 -1449 -101
rect -1403 -147 -1325 -101
rect -1279 -147 -1201 -101
rect -1155 -147 -1077 -101
rect -1031 -147 -953 -101
rect -907 -147 -829 -101
rect -783 -147 -705 -101
rect -659 -147 -581 -101
rect -535 -147 -457 -101
rect -411 -147 -333 -101
rect -287 -147 -209 -101
rect -163 -147 -85 -101
rect -39 -147 39 -101
rect 85 -147 163 -101
rect 209 -147 287 -101
rect 333 -147 411 -101
rect 457 -147 535 -101
rect 581 -147 659 -101
rect 705 -147 783 -101
rect 829 -147 907 -101
rect 953 -147 1031 -101
rect 1077 -147 1155 -101
rect 1201 -147 1279 -101
rect 1325 -147 1403 -101
rect 1449 -147 1527 -101
rect 1573 -147 1651 -101
rect 1697 -147 1775 -101
rect 1821 -147 1899 -101
rect 1945 -147 2023 -101
rect 2069 -147 2147 -101
rect 2193 -147 2271 -101
rect 2317 -147 2395 -101
rect 2441 -147 2519 -101
rect 2565 -147 2643 -101
rect 2689 -147 2767 -101
rect 2813 -147 2891 -101
rect 2937 -147 3015 -101
rect 3061 -147 3139 -101
rect 3185 -147 3263 -101
rect 3309 -147 3387 -101
rect 3433 -147 3511 -101
rect 3557 -147 3635 -101
rect 3681 -147 3759 -101
rect 3805 -147 3883 -101
rect 3929 -147 4007 -101
rect 4053 -147 4131 -101
rect 4177 -147 4255 -101
rect 4301 -147 4379 -101
rect 4425 -147 4503 -101
rect 4549 -147 4627 -101
rect 4673 -147 4751 -101
rect 4797 -147 4875 -101
rect 4921 -147 4999 -101
rect 5045 -147 5123 -101
rect 5169 -147 5247 -101
rect 5293 -147 5371 -101
rect 5417 -147 5495 -101
rect 5541 -147 5619 -101
rect 5665 -147 5743 -101
rect 5789 -147 5867 -101
rect 5913 -147 5991 -101
rect 6037 -147 6115 -101
rect 6161 -147 6239 -101
rect 6285 -147 6363 -101
rect 6409 -147 6487 -101
rect 6533 -147 6611 -101
rect 6657 -147 6735 -101
rect 6781 -147 6859 -101
rect 6905 -147 6983 -101
rect 7029 -147 7107 -101
rect 7153 -147 7231 -101
rect 7277 -147 7355 -101
rect 7401 -147 7479 -101
rect 7525 -147 7603 -101
rect 7649 -147 7727 -101
rect 7773 -147 7851 -101
rect 7897 -147 7975 -101
rect 8021 -147 8099 -101
rect 8145 -147 8223 -101
rect 8269 -147 8347 -101
rect 8393 -147 8471 -101
rect 8517 -147 8595 -101
rect 8641 -147 8719 -101
rect 8765 -147 8843 -101
rect 8889 -147 8967 -101
rect 9013 -147 9091 -101
rect 9137 -147 9215 -101
rect 9261 -147 9339 -101
rect 9385 -147 9463 -101
rect 9509 -147 9587 -101
rect 9633 -147 9711 -101
rect 9757 -147 9835 -101
rect 9881 -147 9959 -101
rect 10005 -147 10083 -101
rect 10129 -147 10207 -101
rect 10253 -147 10331 -101
rect 10377 -147 10455 -101
rect 10501 -147 10579 -101
rect 10625 -147 10703 -101
rect 10749 -147 10827 -101
rect 10873 -147 10951 -101
rect 10997 -147 11075 -101
rect 11121 -147 11199 -101
rect 11245 -147 11323 -101
rect 11369 -147 11447 -101
rect 11493 -147 11571 -101
rect 11617 -147 11695 -101
rect 11741 -147 11819 -101
rect 11865 -147 11943 -101
rect 11989 -147 12067 -101
rect 12113 -147 12191 -101
rect 12237 -147 12315 -101
rect 12361 -147 12439 -101
rect 12485 -147 12563 -101
rect 12609 -147 12687 -101
rect 12733 -147 12811 -101
rect 12857 -147 12935 -101
rect 12981 -147 13059 -101
rect 13105 -147 13183 -101
rect 13229 -147 13307 -101
rect 13353 -147 13431 -101
rect 13477 -147 13555 -101
rect 13601 -147 13679 -101
rect 13725 -147 13803 -101
rect 13849 -147 13927 -101
rect 13973 -147 14051 -101
rect 14097 -147 14175 -101
rect 14221 -147 14299 -101
rect 14345 -147 14423 -101
rect 14469 -147 14547 -101
rect 14593 -147 14671 -101
rect 14717 -147 14795 -101
rect 14841 -147 14919 -101
rect 14965 -147 15043 -101
rect 15089 -147 15167 -101
rect 15213 -147 15291 -101
rect 15337 -147 15415 -101
rect 15461 -147 15539 -101
rect 15585 -147 15663 -101
rect 15709 -147 15787 -101
rect 15833 -147 15911 -101
rect 15957 -147 16035 -101
rect 16081 -147 16159 -101
rect 16205 -147 16283 -101
rect 16329 -147 16407 -101
rect 16453 -147 16531 -101
rect 16577 -147 16655 -101
rect 16701 -147 16779 -101
rect 16825 -147 16903 -101
rect 16949 -147 17027 -101
rect 17073 -147 17151 -101
rect 17197 -147 17275 -101
rect 17321 -147 17399 -101
rect 17445 -147 17523 -101
rect 17569 -147 17647 -101
rect 17693 -147 17771 -101
rect 17817 -147 17895 -101
rect 17941 -147 18019 -101
rect 18065 -147 18143 -101
rect 18189 -147 18267 -101
rect 18313 -147 18324 -101
rect -18324 -225 18324 -147
rect -18324 -271 -18313 -225
rect -18267 -271 -18189 -225
rect -18143 -271 -18065 -225
rect -18019 -271 -17941 -225
rect -17895 -271 -17817 -225
rect -17771 -271 -17693 -225
rect -17647 -271 -17569 -225
rect -17523 -271 -17445 -225
rect -17399 -271 -17321 -225
rect -17275 -271 -17197 -225
rect -17151 -271 -17073 -225
rect -17027 -271 -16949 -225
rect -16903 -271 -16825 -225
rect -16779 -271 -16701 -225
rect -16655 -271 -16577 -225
rect -16531 -271 -16453 -225
rect -16407 -271 -16329 -225
rect -16283 -271 -16205 -225
rect -16159 -271 -16081 -225
rect -16035 -271 -15957 -225
rect -15911 -271 -15833 -225
rect -15787 -271 -15709 -225
rect -15663 -271 -15585 -225
rect -15539 -271 -15461 -225
rect -15415 -271 -15337 -225
rect -15291 -271 -15213 -225
rect -15167 -271 -15089 -225
rect -15043 -271 -14965 -225
rect -14919 -271 -14841 -225
rect -14795 -271 -14717 -225
rect -14671 -271 -14593 -225
rect -14547 -271 -14469 -225
rect -14423 -271 -14345 -225
rect -14299 -271 -14221 -225
rect -14175 -271 -14097 -225
rect -14051 -271 -13973 -225
rect -13927 -271 -13849 -225
rect -13803 -271 -13725 -225
rect -13679 -271 -13601 -225
rect -13555 -271 -13477 -225
rect -13431 -271 -13353 -225
rect -13307 -271 -13229 -225
rect -13183 -271 -13105 -225
rect -13059 -271 -12981 -225
rect -12935 -271 -12857 -225
rect -12811 -271 -12733 -225
rect -12687 -271 -12609 -225
rect -12563 -271 -12485 -225
rect -12439 -271 -12361 -225
rect -12315 -271 -12237 -225
rect -12191 -271 -12113 -225
rect -12067 -271 -11989 -225
rect -11943 -271 -11865 -225
rect -11819 -271 -11741 -225
rect -11695 -271 -11617 -225
rect -11571 -271 -11493 -225
rect -11447 -271 -11369 -225
rect -11323 -271 -11245 -225
rect -11199 -271 -11121 -225
rect -11075 -271 -10997 -225
rect -10951 -271 -10873 -225
rect -10827 -271 -10749 -225
rect -10703 -271 -10625 -225
rect -10579 -271 -10501 -225
rect -10455 -271 -10377 -225
rect -10331 -271 -10253 -225
rect -10207 -271 -10129 -225
rect -10083 -271 -10005 -225
rect -9959 -271 -9881 -225
rect -9835 -271 -9757 -225
rect -9711 -271 -9633 -225
rect -9587 -271 -9509 -225
rect -9463 -271 -9385 -225
rect -9339 -271 -9261 -225
rect -9215 -271 -9137 -225
rect -9091 -271 -9013 -225
rect -8967 -271 -8889 -225
rect -8843 -271 -8765 -225
rect -8719 -271 -8641 -225
rect -8595 -271 -8517 -225
rect -8471 -271 -8393 -225
rect -8347 -271 -8269 -225
rect -8223 -271 -8145 -225
rect -8099 -271 -8021 -225
rect -7975 -271 -7897 -225
rect -7851 -271 -7773 -225
rect -7727 -271 -7649 -225
rect -7603 -271 -7525 -225
rect -7479 -271 -7401 -225
rect -7355 -271 -7277 -225
rect -7231 -271 -7153 -225
rect -7107 -271 -7029 -225
rect -6983 -271 -6905 -225
rect -6859 -271 -6781 -225
rect -6735 -271 -6657 -225
rect -6611 -271 -6533 -225
rect -6487 -271 -6409 -225
rect -6363 -271 -6285 -225
rect -6239 -271 -6161 -225
rect -6115 -271 -6037 -225
rect -5991 -271 -5913 -225
rect -5867 -271 -5789 -225
rect -5743 -271 -5665 -225
rect -5619 -271 -5541 -225
rect -5495 -271 -5417 -225
rect -5371 -271 -5293 -225
rect -5247 -271 -5169 -225
rect -5123 -271 -5045 -225
rect -4999 -271 -4921 -225
rect -4875 -271 -4797 -225
rect -4751 -271 -4673 -225
rect -4627 -271 -4549 -225
rect -4503 -271 -4425 -225
rect -4379 -271 -4301 -225
rect -4255 -271 -4177 -225
rect -4131 -271 -4053 -225
rect -4007 -271 -3929 -225
rect -3883 -271 -3805 -225
rect -3759 -271 -3681 -225
rect -3635 -271 -3557 -225
rect -3511 -271 -3433 -225
rect -3387 -271 -3309 -225
rect -3263 -271 -3185 -225
rect -3139 -271 -3061 -225
rect -3015 -271 -2937 -225
rect -2891 -271 -2813 -225
rect -2767 -271 -2689 -225
rect -2643 -271 -2565 -225
rect -2519 -271 -2441 -225
rect -2395 -271 -2317 -225
rect -2271 -271 -2193 -225
rect -2147 -271 -2069 -225
rect -2023 -271 -1945 -225
rect -1899 -271 -1821 -225
rect -1775 -271 -1697 -225
rect -1651 -271 -1573 -225
rect -1527 -271 -1449 -225
rect -1403 -271 -1325 -225
rect -1279 -271 -1201 -225
rect -1155 -271 -1077 -225
rect -1031 -271 -953 -225
rect -907 -271 -829 -225
rect -783 -271 -705 -225
rect -659 -271 -581 -225
rect -535 -271 -457 -225
rect -411 -271 -333 -225
rect -287 -271 -209 -225
rect -163 -271 -85 -225
rect -39 -271 39 -225
rect 85 -271 163 -225
rect 209 -271 287 -225
rect 333 -271 411 -225
rect 457 -271 535 -225
rect 581 -271 659 -225
rect 705 -271 783 -225
rect 829 -271 907 -225
rect 953 -271 1031 -225
rect 1077 -271 1155 -225
rect 1201 -271 1279 -225
rect 1325 -271 1403 -225
rect 1449 -271 1527 -225
rect 1573 -271 1651 -225
rect 1697 -271 1775 -225
rect 1821 -271 1899 -225
rect 1945 -271 2023 -225
rect 2069 -271 2147 -225
rect 2193 -271 2271 -225
rect 2317 -271 2395 -225
rect 2441 -271 2519 -225
rect 2565 -271 2643 -225
rect 2689 -271 2767 -225
rect 2813 -271 2891 -225
rect 2937 -271 3015 -225
rect 3061 -271 3139 -225
rect 3185 -271 3263 -225
rect 3309 -271 3387 -225
rect 3433 -271 3511 -225
rect 3557 -271 3635 -225
rect 3681 -271 3759 -225
rect 3805 -271 3883 -225
rect 3929 -271 4007 -225
rect 4053 -271 4131 -225
rect 4177 -271 4255 -225
rect 4301 -271 4379 -225
rect 4425 -271 4503 -225
rect 4549 -271 4627 -225
rect 4673 -271 4751 -225
rect 4797 -271 4875 -225
rect 4921 -271 4999 -225
rect 5045 -271 5123 -225
rect 5169 -271 5247 -225
rect 5293 -271 5371 -225
rect 5417 -271 5495 -225
rect 5541 -271 5619 -225
rect 5665 -271 5743 -225
rect 5789 -271 5867 -225
rect 5913 -271 5991 -225
rect 6037 -271 6115 -225
rect 6161 -271 6239 -225
rect 6285 -271 6363 -225
rect 6409 -271 6487 -225
rect 6533 -271 6611 -225
rect 6657 -271 6735 -225
rect 6781 -271 6859 -225
rect 6905 -271 6983 -225
rect 7029 -271 7107 -225
rect 7153 -271 7231 -225
rect 7277 -271 7355 -225
rect 7401 -271 7479 -225
rect 7525 -271 7603 -225
rect 7649 -271 7727 -225
rect 7773 -271 7851 -225
rect 7897 -271 7975 -225
rect 8021 -271 8099 -225
rect 8145 -271 8223 -225
rect 8269 -271 8347 -225
rect 8393 -271 8471 -225
rect 8517 -271 8595 -225
rect 8641 -271 8719 -225
rect 8765 -271 8843 -225
rect 8889 -271 8967 -225
rect 9013 -271 9091 -225
rect 9137 -271 9215 -225
rect 9261 -271 9339 -225
rect 9385 -271 9463 -225
rect 9509 -271 9587 -225
rect 9633 -271 9711 -225
rect 9757 -271 9835 -225
rect 9881 -271 9959 -225
rect 10005 -271 10083 -225
rect 10129 -271 10207 -225
rect 10253 -271 10331 -225
rect 10377 -271 10455 -225
rect 10501 -271 10579 -225
rect 10625 -271 10703 -225
rect 10749 -271 10827 -225
rect 10873 -271 10951 -225
rect 10997 -271 11075 -225
rect 11121 -271 11199 -225
rect 11245 -271 11323 -225
rect 11369 -271 11447 -225
rect 11493 -271 11571 -225
rect 11617 -271 11695 -225
rect 11741 -271 11819 -225
rect 11865 -271 11943 -225
rect 11989 -271 12067 -225
rect 12113 -271 12191 -225
rect 12237 -271 12315 -225
rect 12361 -271 12439 -225
rect 12485 -271 12563 -225
rect 12609 -271 12687 -225
rect 12733 -271 12811 -225
rect 12857 -271 12935 -225
rect 12981 -271 13059 -225
rect 13105 -271 13183 -225
rect 13229 -271 13307 -225
rect 13353 -271 13431 -225
rect 13477 -271 13555 -225
rect 13601 -271 13679 -225
rect 13725 -271 13803 -225
rect 13849 -271 13927 -225
rect 13973 -271 14051 -225
rect 14097 -271 14175 -225
rect 14221 -271 14299 -225
rect 14345 -271 14423 -225
rect 14469 -271 14547 -225
rect 14593 -271 14671 -225
rect 14717 -271 14795 -225
rect 14841 -271 14919 -225
rect 14965 -271 15043 -225
rect 15089 -271 15167 -225
rect 15213 -271 15291 -225
rect 15337 -271 15415 -225
rect 15461 -271 15539 -225
rect 15585 -271 15663 -225
rect 15709 -271 15787 -225
rect 15833 -271 15911 -225
rect 15957 -271 16035 -225
rect 16081 -271 16159 -225
rect 16205 -271 16283 -225
rect 16329 -271 16407 -225
rect 16453 -271 16531 -225
rect 16577 -271 16655 -225
rect 16701 -271 16779 -225
rect 16825 -271 16903 -225
rect 16949 -271 17027 -225
rect 17073 -271 17151 -225
rect 17197 -271 17275 -225
rect 17321 -271 17399 -225
rect 17445 -271 17523 -225
rect 17569 -271 17647 -225
rect 17693 -271 17771 -225
rect 17817 -271 17895 -225
rect 17941 -271 18019 -225
rect 18065 -271 18143 -225
rect 18189 -271 18267 -225
rect 18313 -271 18324 -225
rect -18324 -349 18324 -271
rect -18324 -395 -18313 -349
rect -18267 -395 -18189 -349
rect -18143 -395 -18065 -349
rect -18019 -395 -17941 -349
rect -17895 -395 -17817 -349
rect -17771 -395 -17693 -349
rect -17647 -395 -17569 -349
rect -17523 -395 -17445 -349
rect -17399 -395 -17321 -349
rect -17275 -395 -17197 -349
rect -17151 -395 -17073 -349
rect -17027 -395 -16949 -349
rect -16903 -395 -16825 -349
rect -16779 -395 -16701 -349
rect -16655 -395 -16577 -349
rect -16531 -395 -16453 -349
rect -16407 -395 -16329 -349
rect -16283 -395 -16205 -349
rect -16159 -395 -16081 -349
rect -16035 -395 -15957 -349
rect -15911 -395 -15833 -349
rect -15787 -395 -15709 -349
rect -15663 -395 -15585 -349
rect -15539 -395 -15461 -349
rect -15415 -395 -15337 -349
rect -15291 -395 -15213 -349
rect -15167 -395 -15089 -349
rect -15043 -395 -14965 -349
rect -14919 -395 -14841 -349
rect -14795 -395 -14717 -349
rect -14671 -395 -14593 -349
rect -14547 -395 -14469 -349
rect -14423 -395 -14345 -349
rect -14299 -395 -14221 -349
rect -14175 -395 -14097 -349
rect -14051 -395 -13973 -349
rect -13927 -395 -13849 -349
rect -13803 -395 -13725 -349
rect -13679 -395 -13601 -349
rect -13555 -395 -13477 -349
rect -13431 -395 -13353 -349
rect -13307 -395 -13229 -349
rect -13183 -395 -13105 -349
rect -13059 -395 -12981 -349
rect -12935 -395 -12857 -349
rect -12811 -395 -12733 -349
rect -12687 -395 -12609 -349
rect -12563 -395 -12485 -349
rect -12439 -395 -12361 -349
rect -12315 -395 -12237 -349
rect -12191 -395 -12113 -349
rect -12067 -395 -11989 -349
rect -11943 -395 -11865 -349
rect -11819 -395 -11741 -349
rect -11695 -395 -11617 -349
rect -11571 -395 -11493 -349
rect -11447 -395 -11369 -349
rect -11323 -395 -11245 -349
rect -11199 -395 -11121 -349
rect -11075 -395 -10997 -349
rect -10951 -395 -10873 -349
rect -10827 -395 -10749 -349
rect -10703 -395 -10625 -349
rect -10579 -395 -10501 -349
rect -10455 -395 -10377 -349
rect -10331 -395 -10253 -349
rect -10207 -395 -10129 -349
rect -10083 -395 -10005 -349
rect -9959 -395 -9881 -349
rect -9835 -395 -9757 -349
rect -9711 -395 -9633 -349
rect -9587 -395 -9509 -349
rect -9463 -395 -9385 -349
rect -9339 -395 -9261 -349
rect -9215 -395 -9137 -349
rect -9091 -395 -9013 -349
rect -8967 -395 -8889 -349
rect -8843 -395 -8765 -349
rect -8719 -395 -8641 -349
rect -8595 -395 -8517 -349
rect -8471 -395 -8393 -349
rect -8347 -395 -8269 -349
rect -8223 -395 -8145 -349
rect -8099 -395 -8021 -349
rect -7975 -395 -7897 -349
rect -7851 -395 -7773 -349
rect -7727 -395 -7649 -349
rect -7603 -395 -7525 -349
rect -7479 -395 -7401 -349
rect -7355 -395 -7277 -349
rect -7231 -395 -7153 -349
rect -7107 -395 -7029 -349
rect -6983 -395 -6905 -349
rect -6859 -395 -6781 -349
rect -6735 -395 -6657 -349
rect -6611 -395 -6533 -349
rect -6487 -395 -6409 -349
rect -6363 -395 -6285 -349
rect -6239 -395 -6161 -349
rect -6115 -395 -6037 -349
rect -5991 -395 -5913 -349
rect -5867 -395 -5789 -349
rect -5743 -395 -5665 -349
rect -5619 -395 -5541 -349
rect -5495 -395 -5417 -349
rect -5371 -395 -5293 -349
rect -5247 -395 -5169 -349
rect -5123 -395 -5045 -349
rect -4999 -395 -4921 -349
rect -4875 -395 -4797 -349
rect -4751 -395 -4673 -349
rect -4627 -395 -4549 -349
rect -4503 -395 -4425 -349
rect -4379 -395 -4301 -349
rect -4255 -395 -4177 -349
rect -4131 -395 -4053 -349
rect -4007 -395 -3929 -349
rect -3883 -395 -3805 -349
rect -3759 -395 -3681 -349
rect -3635 -395 -3557 -349
rect -3511 -395 -3433 -349
rect -3387 -395 -3309 -349
rect -3263 -395 -3185 -349
rect -3139 -395 -3061 -349
rect -3015 -395 -2937 -349
rect -2891 -395 -2813 -349
rect -2767 -395 -2689 -349
rect -2643 -395 -2565 -349
rect -2519 -395 -2441 -349
rect -2395 -395 -2317 -349
rect -2271 -395 -2193 -349
rect -2147 -395 -2069 -349
rect -2023 -395 -1945 -349
rect -1899 -395 -1821 -349
rect -1775 -395 -1697 -349
rect -1651 -395 -1573 -349
rect -1527 -395 -1449 -349
rect -1403 -395 -1325 -349
rect -1279 -395 -1201 -349
rect -1155 -395 -1077 -349
rect -1031 -395 -953 -349
rect -907 -395 -829 -349
rect -783 -395 -705 -349
rect -659 -395 -581 -349
rect -535 -395 -457 -349
rect -411 -395 -333 -349
rect -287 -395 -209 -349
rect -163 -395 -85 -349
rect -39 -395 39 -349
rect 85 -395 163 -349
rect 209 -395 287 -349
rect 333 -395 411 -349
rect 457 -395 535 -349
rect 581 -395 659 -349
rect 705 -395 783 -349
rect 829 -395 907 -349
rect 953 -395 1031 -349
rect 1077 -395 1155 -349
rect 1201 -395 1279 -349
rect 1325 -395 1403 -349
rect 1449 -395 1527 -349
rect 1573 -395 1651 -349
rect 1697 -395 1775 -349
rect 1821 -395 1899 -349
rect 1945 -395 2023 -349
rect 2069 -395 2147 -349
rect 2193 -395 2271 -349
rect 2317 -395 2395 -349
rect 2441 -395 2519 -349
rect 2565 -395 2643 -349
rect 2689 -395 2767 -349
rect 2813 -395 2891 -349
rect 2937 -395 3015 -349
rect 3061 -395 3139 -349
rect 3185 -395 3263 -349
rect 3309 -395 3387 -349
rect 3433 -395 3511 -349
rect 3557 -395 3635 -349
rect 3681 -395 3759 -349
rect 3805 -395 3883 -349
rect 3929 -395 4007 -349
rect 4053 -395 4131 -349
rect 4177 -395 4255 -349
rect 4301 -395 4379 -349
rect 4425 -395 4503 -349
rect 4549 -395 4627 -349
rect 4673 -395 4751 -349
rect 4797 -395 4875 -349
rect 4921 -395 4999 -349
rect 5045 -395 5123 -349
rect 5169 -395 5247 -349
rect 5293 -395 5371 -349
rect 5417 -395 5495 -349
rect 5541 -395 5619 -349
rect 5665 -395 5743 -349
rect 5789 -395 5867 -349
rect 5913 -395 5991 -349
rect 6037 -395 6115 -349
rect 6161 -395 6239 -349
rect 6285 -395 6363 -349
rect 6409 -395 6487 -349
rect 6533 -395 6611 -349
rect 6657 -395 6735 -349
rect 6781 -395 6859 -349
rect 6905 -395 6983 -349
rect 7029 -395 7107 -349
rect 7153 -395 7231 -349
rect 7277 -395 7355 -349
rect 7401 -395 7479 -349
rect 7525 -395 7603 -349
rect 7649 -395 7727 -349
rect 7773 -395 7851 -349
rect 7897 -395 7975 -349
rect 8021 -395 8099 -349
rect 8145 -395 8223 -349
rect 8269 -395 8347 -349
rect 8393 -395 8471 -349
rect 8517 -395 8595 -349
rect 8641 -395 8719 -349
rect 8765 -395 8843 -349
rect 8889 -395 8967 -349
rect 9013 -395 9091 -349
rect 9137 -395 9215 -349
rect 9261 -395 9339 -349
rect 9385 -395 9463 -349
rect 9509 -395 9587 -349
rect 9633 -395 9711 -349
rect 9757 -395 9835 -349
rect 9881 -395 9959 -349
rect 10005 -395 10083 -349
rect 10129 -395 10207 -349
rect 10253 -395 10331 -349
rect 10377 -395 10455 -349
rect 10501 -395 10579 -349
rect 10625 -395 10703 -349
rect 10749 -395 10827 -349
rect 10873 -395 10951 -349
rect 10997 -395 11075 -349
rect 11121 -395 11199 -349
rect 11245 -395 11323 -349
rect 11369 -395 11447 -349
rect 11493 -395 11571 -349
rect 11617 -395 11695 -349
rect 11741 -395 11819 -349
rect 11865 -395 11943 -349
rect 11989 -395 12067 -349
rect 12113 -395 12191 -349
rect 12237 -395 12315 -349
rect 12361 -395 12439 -349
rect 12485 -395 12563 -349
rect 12609 -395 12687 -349
rect 12733 -395 12811 -349
rect 12857 -395 12935 -349
rect 12981 -395 13059 -349
rect 13105 -395 13183 -349
rect 13229 -395 13307 -349
rect 13353 -395 13431 -349
rect 13477 -395 13555 -349
rect 13601 -395 13679 -349
rect 13725 -395 13803 -349
rect 13849 -395 13927 -349
rect 13973 -395 14051 -349
rect 14097 -395 14175 -349
rect 14221 -395 14299 -349
rect 14345 -395 14423 -349
rect 14469 -395 14547 -349
rect 14593 -395 14671 -349
rect 14717 -395 14795 -349
rect 14841 -395 14919 -349
rect 14965 -395 15043 -349
rect 15089 -395 15167 -349
rect 15213 -395 15291 -349
rect 15337 -395 15415 -349
rect 15461 -395 15539 -349
rect 15585 -395 15663 -349
rect 15709 -395 15787 -349
rect 15833 -395 15911 -349
rect 15957 -395 16035 -349
rect 16081 -395 16159 -349
rect 16205 -395 16283 -349
rect 16329 -395 16407 -349
rect 16453 -395 16531 -349
rect 16577 -395 16655 -349
rect 16701 -395 16779 -349
rect 16825 -395 16903 -349
rect 16949 -395 17027 -349
rect 17073 -395 17151 -349
rect 17197 -395 17275 -349
rect 17321 -395 17399 -349
rect 17445 -395 17523 -349
rect 17569 -395 17647 -349
rect 17693 -395 17771 -349
rect 17817 -395 17895 -349
rect 17941 -395 18019 -349
rect 18065 -395 18143 -349
rect 18189 -395 18267 -349
rect 18313 -395 18324 -349
rect -18324 -473 18324 -395
rect -18324 -519 -18313 -473
rect -18267 -519 -18189 -473
rect -18143 -519 -18065 -473
rect -18019 -519 -17941 -473
rect -17895 -519 -17817 -473
rect -17771 -519 -17693 -473
rect -17647 -519 -17569 -473
rect -17523 -519 -17445 -473
rect -17399 -519 -17321 -473
rect -17275 -519 -17197 -473
rect -17151 -519 -17073 -473
rect -17027 -519 -16949 -473
rect -16903 -519 -16825 -473
rect -16779 -519 -16701 -473
rect -16655 -519 -16577 -473
rect -16531 -519 -16453 -473
rect -16407 -519 -16329 -473
rect -16283 -519 -16205 -473
rect -16159 -519 -16081 -473
rect -16035 -519 -15957 -473
rect -15911 -519 -15833 -473
rect -15787 -519 -15709 -473
rect -15663 -519 -15585 -473
rect -15539 -519 -15461 -473
rect -15415 -519 -15337 -473
rect -15291 -519 -15213 -473
rect -15167 -519 -15089 -473
rect -15043 -519 -14965 -473
rect -14919 -519 -14841 -473
rect -14795 -519 -14717 -473
rect -14671 -519 -14593 -473
rect -14547 -519 -14469 -473
rect -14423 -519 -14345 -473
rect -14299 -519 -14221 -473
rect -14175 -519 -14097 -473
rect -14051 -519 -13973 -473
rect -13927 -519 -13849 -473
rect -13803 -519 -13725 -473
rect -13679 -519 -13601 -473
rect -13555 -519 -13477 -473
rect -13431 -519 -13353 -473
rect -13307 -519 -13229 -473
rect -13183 -519 -13105 -473
rect -13059 -519 -12981 -473
rect -12935 -519 -12857 -473
rect -12811 -519 -12733 -473
rect -12687 -519 -12609 -473
rect -12563 -519 -12485 -473
rect -12439 -519 -12361 -473
rect -12315 -519 -12237 -473
rect -12191 -519 -12113 -473
rect -12067 -519 -11989 -473
rect -11943 -519 -11865 -473
rect -11819 -519 -11741 -473
rect -11695 -519 -11617 -473
rect -11571 -519 -11493 -473
rect -11447 -519 -11369 -473
rect -11323 -519 -11245 -473
rect -11199 -519 -11121 -473
rect -11075 -519 -10997 -473
rect -10951 -519 -10873 -473
rect -10827 -519 -10749 -473
rect -10703 -519 -10625 -473
rect -10579 -519 -10501 -473
rect -10455 -519 -10377 -473
rect -10331 -519 -10253 -473
rect -10207 -519 -10129 -473
rect -10083 -519 -10005 -473
rect -9959 -519 -9881 -473
rect -9835 -519 -9757 -473
rect -9711 -519 -9633 -473
rect -9587 -519 -9509 -473
rect -9463 -519 -9385 -473
rect -9339 -519 -9261 -473
rect -9215 -519 -9137 -473
rect -9091 -519 -9013 -473
rect -8967 -519 -8889 -473
rect -8843 -519 -8765 -473
rect -8719 -519 -8641 -473
rect -8595 -519 -8517 -473
rect -8471 -519 -8393 -473
rect -8347 -519 -8269 -473
rect -8223 -519 -8145 -473
rect -8099 -519 -8021 -473
rect -7975 -519 -7897 -473
rect -7851 -519 -7773 -473
rect -7727 -519 -7649 -473
rect -7603 -519 -7525 -473
rect -7479 -519 -7401 -473
rect -7355 -519 -7277 -473
rect -7231 -519 -7153 -473
rect -7107 -519 -7029 -473
rect -6983 -519 -6905 -473
rect -6859 -519 -6781 -473
rect -6735 -519 -6657 -473
rect -6611 -519 -6533 -473
rect -6487 -519 -6409 -473
rect -6363 -519 -6285 -473
rect -6239 -519 -6161 -473
rect -6115 -519 -6037 -473
rect -5991 -519 -5913 -473
rect -5867 -519 -5789 -473
rect -5743 -519 -5665 -473
rect -5619 -519 -5541 -473
rect -5495 -519 -5417 -473
rect -5371 -519 -5293 -473
rect -5247 -519 -5169 -473
rect -5123 -519 -5045 -473
rect -4999 -519 -4921 -473
rect -4875 -519 -4797 -473
rect -4751 -519 -4673 -473
rect -4627 -519 -4549 -473
rect -4503 -519 -4425 -473
rect -4379 -519 -4301 -473
rect -4255 -519 -4177 -473
rect -4131 -519 -4053 -473
rect -4007 -519 -3929 -473
rect -3883 -519 -3805 -473
rect -3759 -519 -3681 -473
rect -3635 -519 -3557 -473
rect -3511 -519 -3433 -473
rect -3387 -519 -3309 -473
rect -3263 -519 -3185 -473
rect -3139 -519 -3061 -473
rect -3015 -519 -2937 -473
rect -2891 -519 -2813 -473
rect -2767 -519 -2689 -473
rect -2643 -519 -2565 -473
rect -2519 -519 -2441 -473
rect -2395 -519 -2317 -473
rect -2271 -519 -2193 -473
rect -2147 -519 -2069 -473
rect -2023 -519 -1945 -473
rect -1899 -519 -1821 -473
rect -1775 -519 -1697 -473
rect -1651 -519 -1573 -473
rect -1527 -519 -1449 -473
rect -1403 -519 -1325 -473
rect -1279 -519 -1201 -473
rect -1155 -519 -1077 -473
rect -1031 -519 -953 -473
rect -907 -519 -829 -473
rect -783 -519 -705 -473
rect -659 -519 -581 -473
rect -535 -519 -457 -473
rect -411 -519 -333 -473
rect -287 -519 -209 -473
rect -163 -519 -85 -473
rect -39 -519 39 -473
rect 85 -519 163 -473
rect 209 -519 287 -473
rect 333 -519 411 -473
rect 457 -519 535 -473
rect 581 -519 659 -473
rect 705 -519 783 -473
rect 829 -519 907 -473
rect 953 -519 1031 -473
rect 1077 -519 1155 -473
rect 1201 -519 1279 -473
rect 1325 -519 1403 -473
rect 1449 -519 1527 -473
rect 1573 -519 1651 -473
rect 1697 -519 1775 -473
rect 1821 -519 1899 -473
rect 1945 -519 2023 -473
rect 2069 -519 2147 -473
rect 2193 -519 2271 -473
rect 2317 -519 2395 -473
rect 2441 -519 2519 -473
rect 2565 -519 2643 -473
rect 2689 -519 2767 -473
rect 2813 -519 2891 -473
rect 2937 -519 3015 -473
rect 3061 -519 3139 -473
rect 3185 -519 3263 -473
rect 3309 -519 3387 -473
rect 3433 -519 3511 -473
rect 3557 -519 3635 -473
rect 3681 -519 3759 -473
rect 3805 -519 3883 -473
rect 3929 -519 4007 -473
rect 4053 -519 4131 -473
rect 4177 -519 4255 -473
rect 4301 -519 4379 -473
rect 4425 -519 4503 -473
rect 4549 -519 4627 -473
rect 4673 -519 4751 -473
rect 4797 -519 4875 -473
rect 4921 -519 4999 -473
rect 5045 -519 5123 -473
rect 5169 -519 5247 -473
rect 5293 -519 5371 -473
rect 5417 -519 5495 -473
rect 5541 -519 5619 -473
rect 5665 -519 5743 -473
rect 5789 -519 5867 -473
rect 5913 -519 5991 -473
rect 6037 -519 6115 -473
rect 6161 -519 6239 -473
rect 6285 -519 6363 -473
rect 6409 -519 6487 -473
rect 6533 -519 6611 -473
rect 6657 -519 6735 -473
rect 6781 -519 6859 -473
rect 6905 -519 6983 -473
rect 7029 -519 7107 -473
rect 7153 -519 7231 -473
rect 7277 -519 7355 -473
rect 7401 -519 7479 -473
rect 7525 -519 7603 -473
rect 7649 -519 7727 -473
rect 7773 -519 7851 -473
rect 7897 -519 7975 -473
rect 8021 -519 8099 -473
rect 8145 -519 8223 -473
rect 8269 -519 8347 -473
rect 8393 -519 8471 -473
rect 8517 -519 8595 -473
rect 8641 -519 8719 -473
rect 8765 -519 8843 -473
rect 8889 -519 8967 -473
rect 9013 -519 9091 -473
rect 9137 -519 9215 -473
rect 9261 -519 9339 -473
rect 9385 -519 9463 -473
rect 9509 -519 9587 -473
rect 9633 -519 9711 -473
rect 9757 -519 9835 -473
rect 9881 -519 9959 -473
rect 10005 -519 10083 -473
rect 10129 -519 10207 -473
rect 10253 -519 10331 -473
rect 10377 -519 10455 -473
rect 10501 -519 10579 -473
rect 10625 -519 10703 -473
rect 10749 -519 10827 -473
rect 10873 -519 10951 -473
rect 10997 -519 11075 -473
rect 11121 -519 11199 -473
rect 11245 -519 11323 -473
rect 11369 -519 11447 -473
rect 11493 -519 11571 -473
rect 11617 -519 11695 -473
rect 11741 -519 11819 -473
rect 11865 -519 11943 -473
rect 11989 -519 12067 -473
rect 12113 -519 12191 -473
rect 12237 -519 12315 -473
rect 12361 -519 12439 -473
rect 12485 -519 12563 -473
rect 12609 -519 12687 -473
rect 12733 -519 12811 -473
rect 12857 -519 12935 -473
rect 12981 -519 13059 -473
rect 13105 -519 13183 -473
rect 13229 -519 13307 -473
rect 13353 -519 13431 -473
rect 13477 -519 13555 -473
rect 13601 -519 13679 -473
rect 13725 -519 13803 -473
rect 13849 -519 13927 -473
rect 13973 -519 14051 -473
rect 14097 -519 14175 -473
rect 14221 -519 14299 -473
rect 14345 -519 14423 -473
rect 14469 -519 14547 -473
rect 14593 -519 14671 -473
rect 14717 -519 14795 -473
rect 14841 -519 14919 -473
rect 14965 -519 15043 -473
rect 15089 -519 15167 -473
rect 15213 -519 15291 -473
rect 15337 -519 15415 -473
rect 15461 -519 15539 -473
rect 15585 -519 15663 -473
rect 15709 -519 15787 -473
rect 15833 -519 15911 -473
rect 15957 -519 16035 -473
rect 16081 -519 16159 -473
rect 16205 -519 16283 -473
rect 16329 -519 16407 -473
rect 16453 -519 16531 -473
rect 16577 -519 16655 -473
rect 16701 -519 16779 -473
rect 16825 -519 16903 -473
rect 16949 -519 17027 -473
rect 17073 -519 17151 -473
rect 17197 -519 17275 -473
rect 17321 -519 17399 -473
rect 17445 -519 17523 -473
rect 17569 -519 17647 -473
rect 17693 -519 17771 -473
rect 17817 -519 17895 -473
rect 17941 -519 18019 -473
rect 18065 -519 18143 -473
rect 18189 -519 18267 -473
rect 18313 -519 18324 -473
rect -18324 -597 18324 -519
rect -18324 -643 -18313 -597
rect -18267 -643 -18189 -597
rect -18143 -643 -18065 -597
rect -18019 -643 -17941 -597
rect -17895 -643 -17817 -597
rect -17771 -643 -17693 -597
rect -17647 -643 -17569 -597
rect -17523 -643 -17445 -597
rect -17399 -643 -17321 -597
rect -17275 -643 -17197 -597
rect -17151 -643 -17073 -597
rect -17027 -643 -16949 -597
rect -16903 -643 -16825 -597
rect -16779 -643 -16701 -597
rect -16655 -643 -16577 -597
rect -16531 -643 -16453 -597
rect -16407 -643 -16329 -597
rect -16283 -643 -16205 -597
rect -16159 -643 -16081 -597
rect -16035 -643 -15957 -597
rect -15911 -643 -15833 -597
rect -15787 -643 -15709 -597
rect -15663 -643 -15585 -597
rect -15539 -643 -15461 -597
rect -15415 -643 -15337 -597
rect -15291 -643 -15213 -597
rect -15167 -643 -15089 -597
rect -15043 -643 -14965 -597
rect -14919 -643 -14841 -597
rect -14795 -643 -14717 -597
rect -14671 -643 -14593 -597
rect -14547 -643 -14469 -597
rect -14423 -643 -14345 -597
rect -14299 -643 -14221 -597
rect -14175 -643 -14097 -597
rect -14051 -643 -13973 -597
rect -13927 -643 -13849 -597
rect -13803 -643 -13725 -597
rect -13679 -643 -13601 -597
rect -13555 -643 -13477 -597
rect -13431 -643 -13353 -597
rect -13307 -643 -13229 -597
rect -13183 -643 -13105 -597
rect -13059 -643 -12981 -597
rect -12935 -643 -12857 -597
rect -12811 -643 -12733 -597
rect -12687 -643 -12609 -597
rect -12563 -643 -12485 -597
rect -12439 -643 -12361 -597
rect -12315 -643 -12237 -597
rect -12191 -643 -12113 -597
rect -12067 -643 -11989 -597
rect -11943 -643 -11865 -597
rect -11819 -643 -11741 -597
rect -11695 -643 -11617 -597
rect -11571 -643 -11493 -597
rect -11447 -643 -11369 -597
rect -11323 -643 -11245 -597
rect -11199 -643 -11121 -597
rect -11075 -643 -10997 -597
rect -10951 -643 -10873 -597
rect -10827 -643 -10749 -597
rect -10703 -643 -10625 -597
rect -10579 -643 -10501 -597
rect -10455 -643 -10377 -597
rect -10331 -643 -10253 -597
rect -10207 -643 -10129 -597
rect -10083 -643 -10005 -597
rect -9959 -643 -9881 -597
rect -9835 -643 -9757 -597
rect -9711 -643 -9633 -597
rect -9587 -643 -9509 -597
rect -9463 -643 -9385 -597
rect -9339 -643 -9261 -597
rect -9215 -643 -9137 -597
rect -9091 -643 -9013 -597
rect -8967 -643 -8889 -597
rect -8843 -643 -8765 -597
rect -8719 -643 -8641 -597
rect -8595 -643 -8517 -597
rect -8471 -643 -8393 -597
rect -8347 -643 -8269 -597
rect -8223 -643 -8145 -597
rect -8099 -643 -8021 -597
rect -7975 -643 -7897 -597
rect -7851 -643 -7773 -597
rect -7727 -643 -7649 -597
rect -7603 -643 -7525 -597
rect -7479 -643 -7401 -597
rect -7355 -643 -7277 -597
rect -7231 -643 -7153 -597
rect -7107 -643 -7029 -597
rect -6983 -643 -6905 -597
rect -6859 -643 -6781 -597
rect -6735 -643 -6657 -597
rect -6611 -643 -6533 -597
rect -6487 -643 -6409 -597
rect -6363 -643 -6285 -597
rect -6239 -643 -6161 -597
rect -6115 -643 -6037 -597
rect -5991 -643 -5913 -597
rect -5867 -643 -5789 -597
rect -5743 -643 -5665 -597
rect -5619 -643 -5541 -597
rect -5495 -643 -5417 -597
rect -5371 -643 -5293 -597
rect -5247 -643 -5169 -597
rect -5123 -643 -5045 -597
rect -4999 -643 -4921 -597
rect -4875 -643 -4797 -597
rect -4751 -643 -4673 -597
rect -4627 -643 -4549 -597
rect -4503 -643 -4425 -597
rect -4379 -643 -4301 -597
rect -4255 -643 -4177 -597
rect -4131 -643 -4053 -597
rect -4007 -643 -3929 -597
rect -3883 -643 -3805 -597
rect -3759 -643 -3681 -597
rect -3635 -643 -3557 -597
rect -3511 -643 -3433 -597
rect -3387 -643 -3309 -597
rect -3263 -643 -3185 -597
rect -3139 -643 -3061 -597
rect -3015 -643 -2937 -597
rect -2891 -643 -2813 -597
rect -2767 -643 -2689 -597
rect -2643 -643 -2565 -597
rect -2519 -643 -2441 -597
rect -2395 -643 -2317 -597
rect -2271 -643 -2193 -597
rect -2147 -643 -2069 -597
rect -2023 -643 -1945 -597
rect -1899 -643 -1821 -597
rect -1775 -643 -1697 -597
rect -1651 -643 -1573 -597
rect -1527 -643 -1449 -597
rect -1403 -643 -1325 -597
rect -1279 -643 -1201 -597
rect -1155 -643 -1077 -597
rect -1031 -643 -953 -597
rect -907 -643 -829 -597
rect -783 -643 -705 -597
rect -659 -643 -581 -597
rect -535 -643 -457 -597
rect -411 -643 -333 -597
rect -287 -643 -209 -597
rect -163 -643 -85 -597
rect -39 -643 39 -597
rect 85 -643 163 -597
rect 209 -643 287 -597
rect 333 -643 411 -597
rect 457 -643 535 -597
rect 581 -643 659 -597
rect 705 -643 783 -597
rect 829 -643 907 -597
rect 953 -643 1031 -597
rect 1077 -643 1155 -597
rect 1201 -643 1279 -597
rect 1325 -643 1403 -597
rect 1449 -643 1527 -597
rect 1573 -643 1651 -597
rect 1697 -643 1775 -597
rect 1821 -643 1899 -597
rect 1945 -643 2023 -597
rect 2069 -643 2147 -597
rect 2193 -643 2271 -597
rect 2317 -643 2395 -597
rect 2441 -643 2519 -597
rect 2565 -643 2643 -597
rect 2689 -643 2767 -597
rect 2813 -643 2891 -597
rect 2937 -643 3015 -597
rect 3061 -643 3139 -597
rect 3185 -643 3263 -597
rect 3309 -643 3387 -597
rect 3433 -643 3511 -597
rect 3557 -643 3635 -597
rect 3681 -643 3759 -597
rect 3805 -643 3883 -597
rect 3929 -643 4007 -597
rect 4053 -643 4131 -597
rect 4177 -643 4255 -597
rect 4301 -643 4379 -597
rect 4425 -643 4503 -597
rect 4549 -643 4627 -597
rect 4673 -643 4751 -597
rect 4797 -643 4875 -597
rect 4921 -643 4999 -597
rect 5045 -643 5123 -597
rect 5169 -643 5247 -597
rect 5293 -643 5371 -597
rect 5417 -643 5495 -597
rect 5541 -643 5619 -597
rect 5665 -643 5743 -597
rect 5789 -643 5867 -597
rect 5913 -643 5991 -597
rect 6037 -643 6115 -597
rect 6161 -643 6239 -597
rect 6285 -643 6363 -597
rect 6409 -643 6487 -597
rect 6533 -643 6611 -597
rect 6657 -643 6735 -597
rect 6781 -643 6859 -597
rect 6905 -643 6983 -597
rect 7029 -643 7107 -597
rect 7153 -643 7231 -597
rect 7277 -643 7355 -597
rect 7401 -643 7479 -597
rect 7525 -643 7603 -597
rect 7649 -643 7727 -597
rect 7773 -643 7851 -597
rect 7897 -643 7975 -597
rect 8021 -643 8099 -597
rect 8145 -643 8223 -597
rect 8269 -643 8347 -597
rect 8393 -643 8471 -597
rect 8517 -643 8595 -597
rect 8641 -643 8719 -597
rect 8765 -643 8843 -597
rect 8889 -643 8967 -597
rect 9013 -643 9091 -597
rect 9137 -643 9215 -597
rect 9261 -643 9339 -597
rect 9385 -643 9463 -597
rect 9509 -643 9587 -597
rect 9633 -643 9711 -597
rect 9757 -643 9835 -597
rect 9881 -643 9959 -597
rect 10005 -643 10083 -597
rect 10129 -643 10207 -597
rect 10253 -643 10331 -597
rect 10377 -643 10455 -597
rect 10501 -643 10579 -597
rect 10625 -643 10703 -597
rect 10749 -643 10827 -597
rect 10873 -643 10951 -597
rect 10997 -643 11075 -597
rect 11121 -643 11199 -597
rect 11245 -643 11323 -597
rect 11369 -643 11447 -597
rect 11493 -643 11571 -597
rect 11617 -643 11695 -597
rect 11741 -643 11819 -597
rect 11865 -643 11943 -597
rect 11989 -643 12067 -597
rect 12113 -643 12191 -597
rect 12237 -643 12315 -597
rect 12361 -643 12439 -597
rect 12485 -643 12563 -597
rect 12609 -643 12687 -597
rect 12733 -643 12811 -597
rect 12857 -643 12935 -597
rect 12981 -643 13059 -597
rect 13105 -643 13183 -597
rect 13229 -643 13307 -597
rect 13353 -643 13431 -597
rect 13477 -643 13555 -597
rect 13601 -643 13679 -597
rect 13725 -643 13803 -597
rect 13849 -643 13927 -597
rect 13973 -643 14051 -597
rect 14097 -643 14175 -597
rect 14221 -643 14299 -597
rect 14345 -643 14423 -597
rect 14469 -643 14547 -597
rect 14593 -643 14671 -597
rect 14717 -643 14795 -597
rect 14841 -643 14919 -597
rect 14965 -643 15043 -597
rect 15089 -643 15167 -597
rect 15213 -643 15291 -597
rect 15337 -643 15415 -597
rect 15461 -643 15539 -597
rect 15585 -643 15663 -597
rect 15709 -643 15787 -597
rect 15833 -643 15911 -597
rect 15957 -643 16035 -597
rect 16081 -643 16159 -597
rect 16205 -643 16283 -597
rect 16329 -643 16407 -597
rect 16453 -643 16531 -597
rect 16577 -643 16655 -597
rect 16701 -643 16779 -597
rect 16825 -643 16903 -597
rect 16949 -643 17027 -597
rect 17073 -643 17151 -597
rect 17197 -643 17275 -597
rect 17321 -643 17399 -597
rect 17445 -643 17523 -597
rect 17569 -643 17647 -597
rect 17693 -643 17771 -597
rect 17817 -643 17895 -597
rect 17941 -643 18019 -597
rect 18065 -643 18143 -597
rect 18189 -643 18267 -597
rect 18313 -643 18324 -597
rect -18324 -654 18324 -643
<< end >>
