magic
tech gf180mcuC
magscale 1 10
timestamp 1693222705
<< pwell >>
rect -162 -3908 162 3908
<< nmos >>
rect -50 -3840 50 3840
<< ndiff >>
rect -138 3827 -50 3840
rect -138 -3827 -125 3827
rect -79 -3827 -50 3827
rect -138 -3840 -50 -3827
rect 50 3827 138 3840
rect 50 -3827 79 3827
rect 125 -3827 138 3827
rect 50 -3840 138 -3827
<< ndiffc >>
rect -125 -3827 -79 3827
rect 79 -3827 125 3827
<< polysilicon >>
rect -50 3840 50 3884
rect -50 -3884 50 -3840
<< metal1 >>
rect -125 3827 -79 3838
rect -125 -3838 -79 -3827
rect 79 3827 125 3838
rect 79 -3838 125 -3827
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 38.4 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
