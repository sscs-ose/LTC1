magic
tech gf180mcuC
magscale 1 10
timestamp 1714140926
<< nwell >>
rect -1376 -1318 1376 1318
<< nsubdiff >>
rect -1352 1222 1352 1294
rect -1352 1178 -1280 1222
rect -1352 -1178 -1339 1178
rect -1293 -1178 -1280 1178
rect 1280 1178 1352 1222
rect -1352 -1222 -1280 -1178
rect 1280 -1178 1293 1178
rect 1339 -1178 1352 1178
rect 1280 -1222 1352 -1178
rect -1352 -1294 1352 -1222
<< nsubdiffcont >>
rect -1339 -1178 -1293 1178
rect 1293 -1178 1339 1178
<< polysilicon >>
rect -1160 1089 -1000 1102
rect -1160 1043 -1147 1089
rect -1013 1043 -1000 1089
rect -1160 1000 -1000 1043
rect -1160 -1043 -1000 -1000
rect -1160 -1089 -1147 -1043
rect -1013 -1089 -1000 -1043
rect -1160 -1102 -1000 -1089
rect -920 1089 -760 1102
rect -920 1043 -907 1089
rect -773 1043 -760 1089
rect -920 1000 -760 1043
rect -920 -1043 -760 -1000
rect -920 -1089 -907 -1043
rect -773 -1089 -760 -1043
rect -920 -1102 -760 -1089
rect -680 1089 -520 1102
rect -680 1043 -667 1089
rect -533 1043 -520 1089
rect -680 1000 -520 1043
rect -680 -1043 -520 -1000
rect -680 -1089 -667 -1043
rect -533 -1089 -520 -1043
rect -680 -1102 -520 -1089
rect -440 1089 -280 1102
rect -440 1043 -427 1089
rect -293 1043 -280 1089
rect -440 1000 -280 1043
rect -440 -1043 -280 -1000
rect -440 -1089 -427 -1043
rect -293 -1089 -280 -1043
rect -440 -1102 -280 -1089
rect -200 1089 -40 1102
rect -200 1043 -187 1089
rect -53 1043 -40 1089
rect -200 1000 -40 1043
rect -200 -1043 -40 -1000
rect -200 -1089 -187 -1043
rect -53 -1089 -40 -1043
rect -200 -1102 -40 -1089
rect 40 1089 200 1102
rect 40 1043 53 1089
rect 187 1043 200 1089
rect 40 1000 200 1043
rect 40 -1043 200 -1000
rect 40 -1089 53 -1043
rect 187 -1089 200 -1043
rect 40 -1102 200 -1089
rect 280 1089 440 1102
rect 280 1043 293 1089
rect 427 1043 440 1089
rect 280 1000 440 1043
rect 280 -1043 440 -1000
rect 280 -1089 293 -1043
rect 427 -1089 440 -1043
rect 280 -1102 440 -1089
rect 520 1089 680 1102
rect 520 1043 533 1089
rect 667 1043 680 1089
rect 520 1000 680 1043
rect 520 -1043 680 -1000
rect 520 -1089 533 -1043
rect 667 -1089 680 -1043
rect 520 -1102 680 -1089
rect 760 1089 920 1102
rect 760 1043 773 1089
rect 907 1043 920 1089
rect 760 1000 920 1043
rect 760 -1043 920 -1000
rect 760 -1089 773 -1043
rect 907 -1089 920 -1043
rect 760 -1102 920 -1089
rect 1000 1089 1160 1102
rect 1000 1043 1013 1089
rect 1147 1043 1160 1089
rect 1000 1000 1160 1043
rect 1000 -1043 1160 -1000
rect 1000 -1089 1013 -1043
rect 1147 -1089 1160 -1043
rect 1000 -1102 1160 -1089
<< polycontact >>
rect -1147 1043 -1013 1089
rect -1147 -1089 -1013 -1043
rect -907 1043 -773 1089
rect -907 -1089 -773 -1043
rect -667 1043 -533 1089
rect -667 -1089 -533 -1043
rect -427 1043 -293 1089
rect -427 -1089 -293 -1043
rect -187 1043 -53 1089
rect -187 -1089 -53 -1043
rect 53 1043 187 1089
rect 53 -1089 187 -1043
rect 293 1043 427 1089
rect 293 -1089 427 -1043
rect 533 1043 667 1089
rect 533 -1089 667 -1043
rect 773 1043 907 1089
rect 773 -1089 907 -1043
rect 1013 1043 1147 1089
rect 1013 -1089 1147 -1043
<< ppolyres >>
rect -1160 -1000 -1000 1000
rect -920 -1000 -760 1000
rect -680 -1000 -520 1000
rect -440 -1000 -280 1000
rect -200 -1000 -40 1000
rect 40 -1000 200 1000
rect 280 -1000 440 1000
rect 520 -1000 680 1000
rect 760 -1000 920 1000
rect 1000 -1000 1160 1000
<< metal1 >>
rect -1339 1235 1339 1281
rect -1339 1178 -1293 1235
rect 1293 1178 1339 1235
rect -1158 1043 -1147 1089
rect -1013 1043 -1002 1089
rect -918 1043 -907 1089
rect -773 1043 -762 1089
rect -678 1043 -667 1089
rect -533 1043 -522 1089
rect -438 1043 -427 1089
rect -293 1043 -282 1089
rect -198 1043 -187 1089
rect -53 1043 -42 1089
rect 42 1043 53 1089
rect 187 1043 198 1089
rect 282 1043 293 1089
rect 427 1043 438 1089
rect 522 1043 533 1089
rect 667 1043 678 1089
rect 762 1043 773 1089
rect 907 1043 918 1089
rect 1002 1043 1013 1089
rect 1147 1043 1158 1089
rect -1158 -1089 -1147 -1043
rect -1013 -1089 -1002 -1043
rect -918 -1089 -907 -1043
rect -773 -1089 -762 -1043
rect -678 -1089 -667 -1043
rect -533 -1089 -522 -1043
rect -438 -1089 -427 -1043
rect -293 -1089 -282 -1043
rect -198 -1089 -187 -1043
rect -53 -1089 -42 -1043
rect 42 -1089 53 -1043
rect 187 -1089 198 -1043
rect 282 -1089 293 -1043
rect 427 -1089 438 -1043
rect 522 -1089 533 -1043
rect 667 -1089 678 -1043
rect 762 -1089 773 -1043
rect 907 -1089 918 -1043
rect 1002 -1089 1013 -1043
rect 1147 -1089 1158 -1043
rect -1339 -1235 -1293 -1178
rect 1293 -1235 1339 -1178
rect -1339 -1281 1339 -1235
<< properties >>
string FIXED_BBOX -1316 -1258 1316 1258
string gencell ppolyf_u
string library gf180mcu
string parameters w 0.80 l 10 m 1 nx 10 wmin 0.80 lmin 1.00 rho 315 val 4.315k dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 1 grc 1 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 1
<< end >>
