* NGSPICE file created from Buffer_delayed_mag_flat.ext - technology: gf180mcuC

.subckt pex_Buffer_delayed_mag VSS IN OUT VDD
X0 OUT Inverter_delayed_mag_0.IN VDD.t1 VDD.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X1 Inverter_delayed_mag_0.IN IN.t0 VDD.t3 VDD.t2 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X2 Inverter_delayed_mag_0.IN IN.t1 VSS.t3 VSS.t2 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X3 OUT Inverter_delayed_mag_0.IN VSS.t1 VSS.t0 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
R0 VDD.n2 VDD.t0 1105.93
R1 VDD.t0 VDD 61.3852
R2 VDD.n2 VDD.t2 55.0852
R3 VDD VDD.t3 5.24355
R4 VDD.n0 VDD.t1 5.09693
R5 VDD.n4 VDD.n3 3.1505
R6 VDD.n3 VDD.n2 3.1505
R7 VDD.n4 VDD.n0 0.317357
R8 VDD VDD.n0 0.147133
R9 VDD.n3 VDD.n1 0.0785186
R10 VDD VDD.n4 0.00219811
R11 OUT OUT.n1 9.33985
R12 OUT OUT.n0 5.17407
R13 IN.n0 IN.t0 7.483
R14 IN.n0 IN.t1 4.636
R15 IN IN.n0 4.17425
R16 VSS.n0 VSS.t0 219.273
R17 VSS.n3 VSS.t2 214.072
R18 VSS.n5 VSS.t3 9.45851
R19 VSS.n1 VSS.t1 9.30518
R20 VSS.n5 VSS.n4 2.6005
R21 VSS.n4 VSS.n3 2.6005
R22 VSS VSS.n1 0.310668
R23 VSS.n4 VSS.n2 0.177715
R24 VSS.n1 VSS.n0 0.152211
R25 VSS.n0 VSS 0.00219811
R26 VSS VSS.n5 0.00219811
C0 IN VDD 0.311f
C1 OUT VDD 0.103f
C2 VDD Inverter_delayed_mag_0.IN 0.495f
C3 IN Inverter_delayed_mag_0.IN 0.0985f
C4 OUT Inverter_delayed_mag_0.IN 0.0995f
C5 IN VSS 0.562f
C6 OUT VSS 0.147f
C7 Inverter_delayed_mag_0.IN VSS 0.702f
C8 VDD VSS 1.75f
.ends

