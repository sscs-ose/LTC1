magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2000 -2000 2764 2500
<< polysilicon >>
rect 0 487 102 500
rect 0 441 13 487
rect 59 441 102 487
rect 0 380 102 441
rect 0 334 13 380
rect 59 334 102 380
rect 0 273 102 334
rect 0 227 13 273
rect 59 227 102 273
rect 0 166 102 227
rect 0 120 13 166
rect 59 120 102 166
rect 0 59 102 120
rect 0 13 13 59
rect 59 13 102 59
rect 0 0 102 13
rect 662 487 764 500
rect 662 441 705 487
rect 751 441 764 487
rect 662 380 764 441
rect 662 334 705 380
rect 751 334 764 380
rect 662 273 764 334
rect 662 227 705 273
rect 751 227 764 273
rect 662 166 764 227
rect 662 120 705 166
rect 751 120 764 166
rect 662 59 764 120
rect 662 13 705 59
rect 751 13 764 59
rect 662 0 764 13
<< polycontact >>
rect 13 441 59 487
rect 13 334 59 380
rect 13 227 59 273
rect 13 120 59 166
rect 13 13 59 59
rect 705 441 751 487
rect 705 334 751 380
rect 705 227 751 273
rect 705 120 751 166
rect 705 13 751 59
<< ppolyres >>
rect 102 0 662 500
<< metal1 >>
rect 2 487 70 498
rect 2 441 13 487
rect 59 441 70 487
rect 2 380 70 441
rect 2 334 13 380
rect 59 334 70 380
rect 2 273 70 334
rect 2 227 13 273
rect 59 227 70 273
rect 2 166 70 227
rect 2 120 13 166
rect 59 120 70 166
rect 2 59 70 120
rect 2 13 13 59
rect 59 13 70 59
rect 2 2 70 13
rect 694 487 762 498
rect 694 441 705 487
rect 751 441 762 487
rect 694 380 762 441
rect 694 334 705 380
rect 751 334 762 380
rect 694 273 762 334
rect 694 227 705 273
rect 751 227 762 273
rect 694 166 762 227
rect 694 120 705 166
rect 751 120 762 166
rect 694 59 762 120
rect 694 13 705 59
rect 751 13 762 59
rect 694 2 762 13
<< labels >>
rlabel polycontact 728 250 728 250 4 MINUS
rlabel polycontact 36 250 36 250 4 PLUS
<< end >>
