magic
tech gf180mcuC
magscale 1 10
timestamp 1692518709
<< nwell >>
rect 0 0 1924 531
<< pwell >>
rect 62 -270 1862 -72
<< nmos >>
rect 178 -196 234 -146
rect 346 -196 402 -146
rect 514 -196 570 -146
rect 682 -196 738 -146
rect 850 -196 906 -146
rect 1018 -196 1074 -146
rect 1186 -196 1242 -146
rect 1354 -196 1410 -146
rect 1522 -196 1578 -146
rect 1690 -196 1746 -146
<< pmos >>
rect 178 136 234 186
rect 346 136 402 186
rect 514 136 570 186
rect 682 136 738 186
rect 850 136 906 186
rect 1018 136 1074 186
rect 1186 136 1242 186
rect 1354 136 1410 186
rect 1522 136 1578 186
rect 1690 136 1746 186
<< ndiff >>
rect 86 -146 158 -135
rect 254 -146 326 -135
rect 422 -146 494 -135
rect 590 -146 662 -135
rect 758 -146 830 -135
rect 926 -146 998 -135
rect 1094 -146 1166 -135
rect 1262 -146 1334 -135
rect 1430 -146 1502 -135
rect 1598 -146 1670 -135
rect 1766 -146 1838 -135
rect 86 -148 178 -146
rect 86 -194 99 -148
rect 145 -194 178 -148
rect 86 -196 178 -194
rect 234 -148 346 -146
rect 234 -194 267 -148
rect 313 -194 346 -148
rect 234 -196 346 -194
rect 402 -148 514 -146
rect 402 -194 435 -148
rect 481 -194 514 -148
rect 402 -196 514 -194
rect 570 -148 682 -146
rect 570 -194 603 -148
rect 649 -194 682 -148
rect 570 -196 682 -194
rect 738 -148 850 -146
rect 738 -194 771 -148
rect 817 -194 850 -148
rect 738 -196 850 -194
rect 906 -148 1018 -146
rect 906 -194 939 -148
rect 985 -194 1018 -148
rect 906 -196 1018 -194
rect 1074 -148 1186 -146
rect 1074 -194 1107 -148
rect 1153 -194 1186 -148
rect 1074 -196 1186 -194
rect 1242 -148 1354 -146
rect 1242 -194 1275 -148
rect 1321 -194 1354 -148
rect 1242 -196 1354 -194
rect 1410 -148 1522 -146
rect 1410 -194 1443 -148
rect 1489 -194 1522 -148
rect 1410 -196 1522 -194
rect 1578 -148 1690 -146
rect 1578 -194 1611 -148
rect 1657 -194 1690 -148
rect 1578 -196 1690 -194
rect 1746 -148 1838 -146
rect 1746 -194 1779 -148
rect 1825 -194 1838 -148
rect 1746 -196 1838 -194
rect 86 -207 158 -196
rect 254 -207 326 -196
rect 422 -207 494 -196
rect 590 -207 662 -196
rect 758 -207 830 -196
rect 926 -207 998 -196
rect 1094 -207 1166 -196
rect 1262 -207 1334 -196
rect 1430 -207 1502 -196
rect 1598 -207 1670 -196
rect 1766 -207 1838 -196
<< pdiff >>
rect 86 186 158 197
rect 254 186 326 197
rect 422 186 494 197
rect 590 186 662 197
rect 758 186 830 197
rect 926 186 998 197
rect 1094 186 1166 197
rect 1262 186 1334 197
rect 1430 186 1502 197
rect 1598 186 1670 197
rect 1766 186 1838 197
rect 86 184 178 186
rect 86 138 99 184
rect 145 138 178 184
rect 86 136 178 138
rect 234 184 346 186
rect 234 138 267 184
rect 313 138 346 184
rect 234 136 346 138
rect 402 184 514 186
rect 402 138 435 184
rect 481 138 514 184
rect 402 136 514 138
rect 570 184 682 186
rect 570 138 603 184
rect 649 138 682 184
rect 570 136 682 138
rect 738 184 850 186
rect 738 138 771 184
rect 817 138 850 184
rect 738 136 850 138
rect 906 184 1018 186
rect 906 138 939 184
rect 985 138 1018 184
rect 906 136 1018 138
rect 1074 184 1186 186
rect 1074 138 1107 184
rect 1153 138 1186 184
rect 1074 136 1186 138
rect 1242 184 1354 186
rect 1242 138 1275 184
rect 1321 138 1354 184
rect 1242 136 1354 138
rect 1410 184 1522 186
rect 1410 138 1443 184
rect 1489 138 1522 184
rect 1410 136 1522 138
rect 1578 184 1690 186
rect 1578 138 1611 184
rect 1657 138 1690 184
rect 1578 136 1690 138
rect 1746 184 1838 186
rect 1746 138 1779 184
rect 1825 138 1838 184
rect 1746 136 1838 138
rect 86 125 158 136
rect 254 125 326 136
rect 422 125 494 136
rect 590 125 662 136
rect 758 125 830 136
rect 926 125 998 136
rect 1094 125 1166 136
rect 1262 125 1334 136
rect 1430 125 1502 136
rect 1598 125 1670 136
rect 1766 125 1838 136
<< ndiffc >>
rect 99 -194 145 -148
rect 267 -194 313 -148
rect 435 -194 481 -148
rect 603 -194 649 -148
rect 771 -194 817 -148
rect 939 -194 985 -148
rect 1107 -194 1153 -148
rect 1275 -194 1321 -148
rect 1443 -194 1489 -148
rect 1611 -194 1657 -148
rect 1779 -194 1825 -148
<< pdiffc >>
rect 99 138 145 184
rect 267 138 313 184
rect 435 138 481 184
rect 603 138 649 184
rect 771 138 817 184
rect 939 138 985 184
rect 1107 138 1153 184
rect 1275 138 1321 184
rect 1443 138 1489 184
rect 1611 138 1657 184
rect 1779 138 1825 184
<< psubdiff >>
rect 31 -478 1884 -464
rect 31 -525 44 -478
rect 96 -525 154 -478
rect 206 -525 264 -478
rect 316 -525 374 -478
rect 426 -525 484 -478
rect 536 -525 594 -478
rect 646 -525 704 -478
rect 756 -525 814 -478
rect 866 -525 924 -478
rect 976 -525 1034 -478
rect 1086 -525 1144 -478
rect 1196 -525 1254 -478
rect 1306 -525 1364 -478
rect 1416 -525 1474 -478
rect 1526 -525 1584 -478
rect 1636 -525 1694 -478
rect 1746 -525 1804 -478
rect 1856 -525 1884 -478
rect 31 -538 1884 -525
<< nsubdiff >>
rect 30 481 1887 494
rect 30 430 44 481
rect 95 430 154 481
rect 205 430 264 481
rect 315 430 374 481
rect 425 430 484 481
rect 535 430 594 481
rect 645 430 704 481
rect 755 430 814 481
rect 865 430 924 481
rect 975 430 1034 481
rect 1085 430 1144 481
rect 1195 430 1254 481
rect 1305 430 1364 481
rect 1415 430 1474 481
rect 1525 430 1584 481
rect 1635 430 1694 481
rect 1745 430 1804 481
rect 1855 430 1887 481
rect 30 416 1887 430
<< psubdiffcont >>
rect 44 -525 96 -478
rect 154 -525 206 -478
rect 264 -525 316 -478
rect 374 -525 426 -478
rect 484 -525 536 -478
rect 594 -525 646 -478
rect 704 -525 756 -478
rect 814 -525 866 -478
rect 924 -525 976 -478
rect 1034 -525 1086 -478
rect 1144 -525 1196 -478
rect 1254 -525 1306 -478
rect 1364 -525 1416 -478
rect 1474 -525 1526 -478
rect 1584 -525 1636 -478
rect 1694 -525 1746 -478
rect 1804 -525 1856 -478
<< nsubdiffcont >>
rect 44 430 95 481
rect 154 430 205 481
rect 264 430 315 481
rect 374 430 425 481
rect 484 430 535 481
rect 594 430 645 481
rect 704 430 755 481
rect 814 430 865 481
rect 924 430 975 481
rect 1034 430 1085 481
rect 1144 430 1195 481
rect 1254 430 1305 481
rect 1364 430 1415 481
rect 1474 430 1525 481
rect 1584 430 1635 481
rect 1694 430 1745 481
rect 1804 430 1855 481
<< polysilicon >>
rect -32 338 40 346
rect -32 333 570 338
rect -32 287 -19 333
rect 27 287 570 333
rect -32 282 570 287
rect -32 274 40 282
rect 178 186 234 230
rect 346 186 402 230
rect 514 186 570 282
rect 842 303 914 316
rect 842 257 855 303
rect 901 257 914 303
rect 1346 303 1418 316
rect 842 244 914 257
rect 682 186 738 230
rect 850 186 906 244
rect 1018 230 1242 266
rect 1346 257 1359 303
rect 1405 257 1418 303
rect 1346 244 1418 257
rect 1018 186 1074 230
rect 1186 186 1242 230
rect 1354 186 1410 244
rect 1522 186 1578 230
rect 1690 186 1746 230
rect 178 92 234 136
rect 346 92 402 136
rect 178 78 402 92
rect 120 65 402 78
rect 120 19 133 65
rect 179 55 402 65
rect 514 92 570 136
rect 682 92 738 136
rect 850 92 906 136
rect 1018 92 1074 136
rect 514 56 738 92
rect 179 19 234 55
rect 120 6 234 19
rect 178 -69 234 6
rect 178 -105 570 -69
rect 178 -146 234 -105
rect 346 -146 402 -105
rect 514 -146 570 -105
rect 682 -79 738 56
rect 682 -115 1074 -79
rect 682 -146 738 -115
rect 850 -146 906 -115
rect 1018 -146 1074 -115
rect 1186 -146 1242 136
rect 1354 92 1410 136
rect 1522 92 1578 136
rect 1690 92 1746 136
rect 1522 62 1746 92
rect 1469 56 1746 62
rect 1469 49 1578 56
rect 1469 3 1482 49
rect 1528 3 1578 49
rect 1469 -10 1578 3
rect 1354 -146 1410 -102
rect 1522 -146 1578 -102
rect 1690 -146 1746 56
rect 178 -240 234 -196
rect 346 -240 402 -196
rect 514 -240 570 -196
rect 682 -240 738 -196
rect 850 -240 906 -196
rect 1018 -240 1074 -196
rect 1186 -230 1242 -196
rect 1354 -230 1410 -196
rect 1522 -230 1578 -196
rect 1186 -266 1578 -230
rect 1690 -240 1746 -196
rect 1186 -332 1242 -266
rect 1170 -345 1242 -332
rect 1170 -391 1183 -345
rect 1229 -391 1242 -345
rect 1170 -404 1242 -391
<< polycontact >>
rect -19 287 27 333
rect 855 257 901 303
rect 1359 257 1405 303
rect 133 19 179 65
rect 1482 3 1528 49
rect 1183 -391 1229 -345
<< metal1 >>
rect 18 481 1899 506
rect 18 430 44 481
rect 95 430 154 481
rect 205 430 264 481
rect 315 430 374 481
rect 425 430 484 481
rect 535 430 594 481
rect 645 430 704 481
rect 755 430 814 481
rect 865 430 924 481
rect 975 430 1034 481
rect 1085 430 1144 481
rect 1195 430 1254 481
rect 1305 430 1364 481
rect 1415 430 1474 481
rect 1525 430 1584 481
rect 1635 430 1694 481
rect 1745 430 1804 481
rect 1855 430 1899 481
rect 18 404 1899 430
rect -32 333 40 346
rect -111 287 -19 333
rect 27 287 40 333
rect -32 274 40 287
rect 99 184 145 404
rect 435 184 481 404
rect 855 316 901 404
rect 1359 316 1405 404
rect 842 303 914 316
rect 1346 303 1418 316
rect 771 257 855 303
rect 901 257 985 303
rect 771 244 985 257
rect 771 184 817 244
rect 939 184 985 244
rect 1275 257 1359 303
rect 1405 257 1489 303
rect 1275 244 1489 257
rect 1275 184 1321 244
rect 1443 184 1489 244
rect 1779 184 1825 404
rect 88 138 99 184
rect 145 138 156 184
rect 256 138 267 184
rect 313 138 324 184
rect 424 138 435 184
rect 481 138 492 184
rect 592 138 603 184
rect 649 138 660 184
rect 760 138 771 184
rect 817 138 828 184
rect 928 138 939 184
rect 985 138 996 184
rect 1096 138 1107 184
rect 1153 138 1164 184
rect 1264 138 1275 184
rect 1321 138 1332 184
rect 1432 138 1443 184
rect 1489 138 1500 184
rect 1600 138 1611 184
rect 1657 138 1668 184
rect 1768 138 1779 184
rect 1825 138 1836 184
rect 267 92 313 138
rect 603 92 649 138
rect 1107 92 1153 138
rect 120 65 192 78
rect -111 19 133 65
rect 179 19 192 65
rect 267 49 1313 92
rect 1611 90 1657 138
rect 1469 49 1539 62
rect 267 46 1482 49
rect 120 6 192 19
rect 395 -56 441 46
rect 1267 3 1482 46
rect 1528 3 1539 49
rect 1611 44 1825 90
rect 1469 -10 1539 3
rect 1779 -43 1825 44
rect 99 -102 481 -56
rect 99 -148 145 -102
rect 435 -148 481 -102
rect 603 -102 985 -56
rect 603 -148 649 -102
rect 939 -148 985 -102
rect 1107 -102 1489 -56
rect 1107 -148 1153 -102
rect 1443 -148 1489 -102
rect 1779 -89 1925 -43
rect 1779 -148 1825 -89
rect 88 -194 99 -148
rect 145 -194 156 -148
rect 256 -194 267 -148
rect 313 -194 324 -148
rect 424 -194 435 -148
rect 481 -194 492 -148
rect 592 -194 603 -148
rect 649 -194 660 -148
rect 760 -194 771 -148
rect 817 -194 828 -148
rect 928 -194 939 -148
rect 985 -194 996 -148
rect 1096 -194 1107 -148
rect 1153 -194 1164 -148
rect 1264 -194 1275 -148
rect 1321 -194 1332 -148
rect 1432 -194 1443 -148
rect 1489 -194 1500 -148
rect 1600 -194 1611 -148
rect 1657 -194 1668 -148
rect 1768 -194 1779 -148
rect 1825 -194 1836 -148
rect 267 -240 313 -194
rect 603 -240 649 -194
rect 267 -286 649 -240
rect 771 -240 817 -194
rect 1107 -240 1153 -194
rect 771 -286 1153 -240
rect 1275 -240 1321 -194
rect 1611 -240 1657 -194
rect 1779 -196 1825 -194
rect 1275 -286 1657 -240
rect -111 -345 1242 -332
rect -111 -378 1183 -345
rect 1170 -391 1183 -378
rect 1229 -391 1242 -345
rect 1170 -404 1242 -391
rect 1611 -450 1657 -286
rect 17 -478 1898 -450
rect 17 -525 44 -478
rect 96 -525 154 -478
rect 206 -525 264 -478
rect 316 -525 374 -478
rect 426 -525 484 -478
rect 536 -525 594 -478
rect 646 -525 704 -478
rect 756 -525 814 -478
rect 866 -525 924 -478
rect 976 -525 1034 -478
rect 1086 -525 1144 -478
rect 1196 -525 1254 -478
rect 1306 -525 1364 -478
rect 1416 -525 1474 -478
rect 1526 -525 1584 -478
rect 1636 -525 1694 -478
rect 1746 -525 1804 -478
rect 1856 -525 1898 -478
rect 17 -552 1898 -525
<< labels >>
flabel metal1 -94 311 -94 311 0 FreeSans 480 0 0 0 B
port 0 nsew
flabel metal1 1841 -70 1841 -70 0 FreeSans 480 0 0 0 OUT
port 6 nsew
flabel nsubdiffcont 951 457 951 457 0 FreeSans 480 0 0 0 VDD
port 7 nsew
flabel metal1 -92 -356 -92 -356 0 FreeSans 480 0 0 0 C
port 4 nsew
flabel psubdiffcont 949 -498 949 -498 0 FreeSans 480 0 0 0 VSS
port 9 nsew
flabel metal1 -91 45 -91 45 0 FreeSans 480 0 0 0 A
port 10 nsew
<< end >>
