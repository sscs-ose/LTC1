magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect 1261 -2000 58836 2069
<< labels >>
rlabel metal3 s 45743 69 45743 69 4 DVSS
port 1 nsew
rlabel metal3 s 48934 69 48934 69 4 DVSS
port 1 nsew
rlabel metal3 s 6432 0 6432 0 4 DVSS
port 1 nsew
rlabel metal3 s 3261 47 3261 47 4 DVSS
port 1 nsew
rlabel metal3 s 9418 69 9418 69 4 DVSS
port 1 nsew
rlabel metal3 s 13611 69 13611 69 4 DVSS
port 1 nsew
rlabel metal3 s 28150 69 28150 69 4 DVSS
port 1 nsew
rlabel metal3 s 35334 69 35334 69 4 DVSS
port 1 nsew
rlabel metal3 s 53701 69 53701 69 4 DVSS
port 1 nsew
rlabel metal3 s 56836 69 56836 69 4 DVSS
port 1 nsew
rlabel metal3 s 44136 69 44136 69 4 DVDD
port 2 nsew
rlabel metal3 s 47320 69 47320 69 4 DVDD
port 2 nsew
rlabel metal3 s 42501 69 42501 69 4 DVDD
port 2 nsew
rlabel metal3 s 11795 69 11795 69 4 DVDD
port 2 nsew
rlabel metal3 s 22234 69 22234 69 4 DVDD
port 2 nsew
rlabel metal3 s 19120 69 19120 69 4 DVDD
port 2 nsew
rlabel metal3 s 15905 69 15905 69 4 DVDD
port 2 nsew
rlabel metal3 s 29692 69 29692 69 4 DVDD
port 2 nsew
rlabel metal3 s 25470 69 25470 69 4 DVDD
port 2 nsew
rlabel metal3 s 32104 69 32104 69 4 DVDD
port 2 nsew
rlabel metal3 s 55292 69 55292 69 4 DVDD
port 2 nsew
rlabel metal3 s 40880 69 40880 69 4 DVDD
port 2 nsew
rlabel metal3 s 37660 69 37660 69 4 VSS
port 3 nsew
rlabel metal3 s 52136 69 52136 69 4 VSS
port 3 nsew
rlabel metal3 s 50526 69 50526 69 4 VDD
port 4 nsew
rlabel metal3 s 39308 69 39308 69 4 VDD
port 4 nsew
<< end >>
