magic
tech gf180mcuC
magscale 1 10
timestamp 1691428906
<< nwell >>
rect 0 0 884 935
<< pwell >>
rect 62 -523 822 -51
<< nmos >>
rect 174 -219 230 -119
rect 334 -219 390 -119
rect 494 -219 550 -119
rect 654 -219 710 -119
rect 174 -455 230 -355
rect 334 -455 390 -355
rect 494 -455 550 -355
rect 654 -455 710 -355
<< pmos >>
rect 174 466 230 666
rect 334 466 390 666
rect 494 466 550 666
rect 654 466 710 666
rect 174 130 230 330
rect 334 130 390 330
rect 494 130 550 330
rect 654 130 710 330
<< ndiff >>
rect 86 -132 174 -119
rect 86 -206 99 -132
rect 145 -206 174 -132
rect 86 -219 174 -206
rect 230 -132 334 -119
rect 230 -206 259 -132
rect 305 -206 334 -132
rect 230 -219 334 -206
rect 390 -132 494 -119
rect 390 -206 419 -132
rect 465 -206 494 -132
rect 390 -219 494 -206
rect 550 -132 654 -119
rect 550 -206 579 -132
rect 625 -206 654 -132
rect 550 -219 654 -206
rect 710 -132 798 -119
rect 710 -206 739 -132
rect 785 -206 798 -132
rect 710 -219 798 -206
rect 86 -368 174 -355
rect 86 -442 99 -368
rect 145 -442 174 -368
rect 86 -455 174 -442
rect 230 -368 334 -355
rect 230 -442 259 -368
rect 305 -442 334 -368
rect 230 -455 334 -442
rect 390 -368 494 -355
rect 390 -442 419 -368
rect 465 -442 494 -368
rect 390 -455 494 -442
rect 550 -368 654 -355
rect 550 -442 579 -368
rect 625 -442 654 -368
rect 550 -455 654 -442
rect 710 -368 798 -355
rect 710 -442 739 -368
rect 785 -442 798 -368
rect 710 -455 798 -442
<< pdiff >>
rect 86 653 174 666
rect 86 479 99 653
rect 145 479 174 653
rect 86 466 174 479
rect 230 653 334 666
rect 230 479 259 653
rect 305 479 334 653
rect 230 466 334 479
rect 390 653 494 666
rect 390 479 419 653
rect 465 479 494 653
rect 390 466 494 479
rect 550 653 654 666
rect 550 479 579 653
rect 625 479 654 653
rect 550 466 654 479
rect 710 653 798 666
rect 710 479 739 653
rect 785 479 798 653
rect 710 466 798 479
rect 86 317 174 330
rect 86 143 99 317
rect 145 143 174 317
rect 86 130 174 143
rect 230 317 334 330
rect 230 143 259 317
rect 305 143 334 317
rect 230 130 334 143
rect 390 317 494 330
rect 390 143 419 317
rect 465 143 494 317
rect 390 130 494 143
rect 550 317 654 330
rect 550 143 579 317
rect 625 143 654 317
rect 550 130 654 143
rect 710 317 798 330
rect 710 143 739 317
rect 785 143 798 317
rect 710 130 798 143
<< ndiffc >>
rect 99 -206 145 -132
rect 259 -206 305 -132
rect 419 -206 465 -132
rect 579 -206 625 -132
rect 739 -206 785 -132
rect 99 -442 145 -368
rect 259 -442 305 -368
rect 419 -442 465 -368
rect 579 -442 625 -368
rect 739 -442 785 -368
<< pdiffc >>
rect 99 479 145 653
rect 259 479 305 653
rect 419 479 465 653
rect 579 479 625 653
rect 739 479 785 653
rect 99 143 145 317
rect 259 143 305 317
rect 419 143 465 317
rect 579 143 625 317
rect 739 143 785 317
<< psubdiff >>
rect 32 -580 847 -562
rect 32 -635 54 -580
rect 818 -635 847 -580
rect 32 -653 847 -635
<< nsubdiff >>
rect 34 893 849 910
rect 34 833 63 893
rect 810 833 849 893
rect 34 820 849 833
<< psubdiffcont >>
rect 54 -635 818 -580
<< nsubdiffcont >>
rect 63 833 810 893
<< polysilicon >>
rect 174 666 230 710
rect 334 666 390 710
rect 494 666 550 710
rect 654 666 710 710
rect 174 330 230 466
rect 334 330 390 466
rect 494 330 550 466
rect 654 330 710 466
rect 174 86 230 130
rect 334 86 390 130
rect 494 86 550 130
rect 654 86 710 130
rect 174 42 710 86
rect 174 23 230 42
rect 128 10 230 23
rect 128 -39 144 10
rect 191 -39 230 10
rect 128 -54 230 -39
rect 174 -119 230 -54
rect 334 -119 390 42
rect 494 -119 550 42
rect 654 -119 710 42
rect 174 -355 230 -219
rect 334 -355 390 -219
rect 494 -355 550 -219
rect 654 -355 710 -219
rect 174 -499 230 -455
rect 334 -499 390 -455
rect 494 -499 550 -455
rect 654 -499 710 -455
<< polycontact >>
rect 144 -39 191 10
<< metal1 >>
rect 0 893 884 935
rect 0 833 63 893
rect 810 833 884 893
rect 0 796 884 833
rect 99 653 145 796
rect 99 317 145 479
rect 99 132 145 143
rect 259 653 305 664
rect 259 317 305 479
rect 128 13 205 23
rect -1 10 205 13
rect -1 -33 144 10
rect 128 -39 144 -33
rect 191 -39 205 10
rect 128 -54 205 -39
rect 259 12 305 143
rect 419 653 465 796
rect 419 317 465 479
rect 419 132 465 143
rect 579 653 625 664
rect 579 317 625 479
rect 579 12 625 143
rect 739 653 785 796
rect 739 317 785 479
rect 739 132 785 143
rect 259 -34 885 12
rect 99 -132 145 -121
rect 99 -368 145 -206
rect 99 -535 145 -442
rect 259 -132 305 -34
rect 259 -368 305 -206
rect 259 -453 305 -442
rect 419 -132 465 -121
rect 419 -368 465 -206
rect 419 -535 465 -442
rect 579 -132 625 -34
rect 579 -368 625 -206
rect 579 -453 625 -442
rect 739 -132 785 -121
rect 739 -368 785 -206
rect 739 -535 785 -442
rect 0 -580 884 -535
rect 0 -635 54 -580
rect 818 -635 884 -580
rect 0 -674 884 -635
<< labels >>
flabel nsubdiffcont 434 863 434 863 0 FreeSans 800 0 0 0 VDD
port 0 nsew
flabel psubdiffcont 425 -618 428 -615 0 FreeSans 800 0 0 0 VSS
port 1 nsew
flabel metal1 27 -17 27 -17 0 FreeSans 800 0 0 0 IN
port 3 nsew
flabel metal1 851 -11 851 -11 0 FreeSans 800 0 0 0 OUT
port 5 nsew
<< end >>
