magic
tech gf180mcuC
magscale 1 10
timestamp 1692168538
<< nwell >>
rect 0 1710 442 1828
rect 404 1328 442 1710
rect 1250 423 1362 891
<< metal1 >>
rect 0 1710 442 1828
rect 1481 1706 1956 1828
rect -132 1542 -52 1553
rect -132 1486 -120 1542
rect -64 1486 -52 1542
rect -132 1473 -52 1486
rect 415 1501 489 1502
rect 415 1445 424 1501
rect 480 1445 489 1501
rect 415 1444 489 1445
rect -119 1375 129 1390
rect -119 1319 52 1375
rect 108 1319 129 1375
rect 1640 1372 1713 1385
rect 322 1355 404 1359
rect -119 1309 129 1319
rect 1640 1316 1647 1372
rect 1703 1316 1713 1372
rect 1640 1302 1713 1316
rect 404 1024 443 1050
rect 404 1023 488 1024
rect 404 959 415 1023
rect 479 959 488 1023
rect 404 958 488 959
rect 404 937 443 958
rect 1197 792 1352 891
rect 1834 867 1956 1706
rect 1848 834 1896 867
rect -146 511 68 564
rect 1264 543 1343 548
rect 1264 489 1276 543
rect 1330 539 1343 543
rect 1330 489 1378 539
rect 1264 477 1378 489
rect 1332 459 1378 477
rect 41 426 119 434
rect 41 372 53 426
rect 107 422 119 426
rect 107 376 182 422
rect 107 372 119 376
rect 41 361 119 372
rect 1234 373 1281 418
rect 1234 326 1360 373
rect 2846 350 2920 397
rect 415 81 479 90
rect 415 43 416 81
rect 38 19 416 43
rect 478 43 479 81
rect 1244 50 1391 92
rect 1200 43 1391 50
rect 478 19 1391 43
rect 38 -21 1391 19
<< via1 >>
rect -120 1486 -64 1542
rect 424 1445 480 1501
rect 52 1319 108 1375
rect 1647 1316 1703 1372
rect 415 959 479 1023
rect 1276 489 1330 543
rect 53 372 107 426
rect 416 19 478 81
<< metal2 >>
rect -132 1542 -52 1553
rect -132 1486 -120 1542
rect -64 1512 480 1542
rect -64 1501 491 1512
rect -64 1486 424 1501
rect -132 1473 -52 1486
rect 412 1445 424 1486
rect 480 1445 491 1501
rect 412 1437 491 1445
rect 424 1436 480 1437
rect 44 1375 114 1391
rect 44 1319 52 1375
rect 108 1319 114 1375
rect 1640 1372 1713 1385
rect 44 1309 114 1319
rect 1275 1316 1647 1372
rect 1703 1316 1713 1372
rect 52 434 108 1309
rect 403 1023 492 1039
rect 403 959 415 1023
rect 479 959 492 1023
rect 403 944 492 959
rect 41 426 119 434
rect 41 372 53 426
rect 107 372 119 426
rect 41 361 119 372
rect 415 94 479 944
rect 1275 548 1331 1316
rect 1640 1302 1713 1316
rect 1264 543 1343 548
rect 1264 489 1276 543
rect 1330 489 1343 543
rect 1264 477 1343 489
rect 396 81 499 94
rect 396 19 416 81
rect 478 19 499 81
rect 396 7 499 19
use AND  AND_0
timestamp 1692166961
transform 1 0 422 0 1 1074
box -18 -137 1331 754
use AND  AND_1
timestamp 1692166961
transform 1 0 18 0 1 137
box -18 -137 1331 754
use Inverter  Inverter_0
timestamp 1692166831
transform 1 0 118 0 1 1151
box -118 -214 286 599
use OR  OR_0 ~/GF180Projects/GF_INV/Magic
timestamp 1692166961
transform 1 0 1327 0 1 129
box 0 -150 1631 762
<< labels >>
flabel metal1 -113 548 -113 548 0 FreeSans 480 0 0 0 A
port 0 nsew
flabel via1 -89 1523 -89 1523 0 FreeSans 480 0 0 0 B
port 1 nsew
flabel metal1 274 1774 274 1774 0 FreeSans 480 0 0 0 VDD
port 2 nsew
flabel metal1 804 8 804 8 0 FreeSans 480 0 0 0 VSS
port 3 nsew
flabel metal1 -97 1358 -97 1358 0 FreeSans 480 0 0 0 SEL
port 4 nsew
flabel metal1 2907 383 2907 383 0 FreeSans 480 0 0 0 OUT
port 5 nsew
<< end >>
