magic
tech gf180mcuC
magscale 1 10
timestamp 1697518002
<< pwell >>
rect -2916 -348 2916 348
<< nmos >>
rect -2804 -280 -2704 280
rect -2600 -280 -2500 280
rect -2396 -280 -2296 280
rect -2192 -280 -2092 280
rect -1988 -280 -1888 280
rect -1784 -280 -1684 280
rect -1580 -280 -1480 280
rect -1376 -280 -1276 280
rect -1172 -280 -1072 280
rect -968 -280 -868 280
rect -764 -280 -664 280
rect -560 -280 -460 280
rect -356 -280 -256 280
rect -152 -280 -52 280
rect 52 -280 152 280
rect 256 -280 356 280
rect 460 -280 560 280
rect 664 -280 764 280
rect 868 -280 968 280
rect 1072 -280 1172 280
rect 1276 -280 1376 280
rect 1480 -280 1580 280
rect 1684 -280 1784 280
rect 1888 -280 1988 280
rect 2092 -280 2192 280
rect 2296 -280 2396 280
rect 2500 -280 2600 280
rect 2704 -280 2804 280
<< ndiff >>
rect -2892 267 -2804 280
rect -2892 -267 -2879 267
rect -2833 -267 -2804 267
rect -2892 -280 -2804 -267
rect -2704 267 -2600 280
rect -2704 -267 -2675 267
rect -2629 -267 -2600 267
rect -2704 -280 -2600 -267
rect -2500 267 -2396 280
rect -2500 -267 -2471 267
rect -2425 -267 -2396 267
rect -2500 -280 -2396 -267
rect -2296 267 -2192 280
rect -2296 -267 -2267 267
rect -2221 -267 -2192 267
rect -2296 -280 -2192 -267
rect -2092 267 -1988 280
rect -2092 -267 -2063 267
rect -2017 -267 -1988 267
rect -2092 -280 -1988 -267
rect -1888 267 -1784 280
rect -1888 -267 -1859 267
rect -1813 -267 -1784 267
rect -1888 -280 -1784 -267
rect -1684 267 -1580 280
rect -1684 -267 -1655 267
rect -1609 -267 -1580 267
rect -1684 -280 -1580 -267
rect -1480 267 -1376 280
rect -1480 -267 -1451 267
rect -1405 -267 -1376 267
rect -1480 -280 -1376 -267
rect -1276 267 -1172 280
rect -1276 -267 -1247 267
rect -1201 -267 -1172 267
rect -1276 -280 -1172 -267
rect -1072 267 -968 280
rect -1072 -267 -1043 267
rect -997 -267 -968 267
rect -1072 -280 -968 -267
rect -868 267 -764 280
rect -868 -267 -839 267
rect -793 -267 -764 267
rect -868 -280 -764 -267
rect -664 267 -560 280
rect -664 -267 -635 267
rect -589 -267 -560 267
rect -664 -280 -560 -267
rect -460 267 -356 280
rect -460 -267 -431 267
rect -385 -267 -356 267
rect -460 -280 -356 -267
rect -256 267 -152 280
rect -256 -267 -227 267
rect -181 -267 -152 267
rect -256 -280 -152 -267
rect -52 267 52 280
rect -52 -267 -23 267
rect 23 -267 52 267
rect -52 -280 52 -267
rect 152 267 256 280
rect 152 -267 181 267
rect 227 -267 256 267
rect 152 -280 256 -267
rect 356 267 460 280
rect 356 -267 385 267
rect 431 -267 460 267
rect 356 -280 460 -267
rect 560 267 664 280
rect 560 -267 589 267
rect 635 -267 664 267
rect 560 -280 664 -267
rect 764 267 868 280
rect 764 -267 793 267
rect 839 -267 868 267
rect 764 -280 868 -267
rect 968 267 1072 280
rect 968 -267 997 267
rect 1043 -267 1072 267
rect 968 -280 1072 -267
rect 1172 267 1276 280
rect 1172 -267 1201 267
rect 1247 -267 1276 267
rect 1172 -280 1276 -267
rect 1376 267 1480 280
rect 1376 -267 1405 267
rect 1451 -267 1480 267
rect 1376 -280 1480 -267
rect 1580 267 1684 280
rect 1580 -267 1609 267
rect 1655 -267 1684 267
rect 1580 -280 1684 -267
rect 1784 267 1888 280
rect 1784 -267 1813 267
rect 1859 -267 1888 267
rect 1784 -280 1888 -267
rect 1988 267 2092 280
rect 1988 -267 2017 267
rect 2063 -267 2092 267
rect 1988 -280 2092 -267
rect 2192 267 2296 280
rect 2192 -267 2221 267
rect 2267 -267 2296 267
rect 2192 -280 2296 -267
rect 2396 267 2500 280
rect 2396 -267 2425 267
rect 2471 -267 2500 267
rect 2396 -280 2500 -267
rect 2600 267 2704 280
rect 2600 -267 2629 267
rect 2675 -267 2704 267
rect 2600 -280 2704 -267
rect 2804 267 2892 280
rect 2804 -267 2833 267
rect 2879 -267 2892 267
rect 2804 -280 2892 -267
<< ndiffc >>
rect -2879 -267 -2833 267
rect -2675 -267 -2629 267
rect -2471 -267 -2425 267
rect -2267 -267 -2221 267
rect -2063 -267 -2017 267
rect -1859 -267 -1813 267
rect -1655 -267 -1609 267
rect -1451 -267 -1405 267
rect -1247 -267 -1201 267
rect -1043 -267 -997 267
rect -839 -267 -793 267
rect -635 -267 -589 267
rect -431 -267 -385 267
rect -227 -267 -181 267
rect -23 -267 23 267
rect 181 -267 227 267
rect 385 -267 431 267
rect 589 -267 635 267
rect 793 -267 839 267
rect 997 -267 1043 267
rect 1201 -267 1247 267
rect 1405 -267 1451 267
rect 1609 -267 1655 267
rect 1813 -267 1859 267
rect 2017 -267 2063 267
rect 2221 -267 2267 267
rect 2425 -267 2471 267
rect 2629 -267 2675 267
rect 2833 -267 2879 267
<< polysilicon >>
rect -2804 280 -2704 324
rect -2600 280 -2500 324
rect -2396 280 -2296 324
rect -2192 280 -2092 324
rect -1988 280 -1888 324
rect -1784 280 -1684 324
rect -1580 280 -1480 324
rect -1376 280 -1276 324
rect -1172 280 -1072 324
rect -968 280 -868 324
rect -764 280 -664 324
rect -560 280 -460 324
rect -356 280 -256 324
rect -152 280 -52 324
rect 52 280 152 324
rect 256 280 356 324
rect 460 280 560 324
rect 664 280 764 324
rect 868 280 968 324
rect 1072 280 1172 324
rect 1276 280 1376 324
rect 1480 280 1580 324
rect 1684 280 1784 324
rect 1888 280 1988 324
rect 2092 280 2192 324
rect 2296 280 2396 324
rect 2500 280 2600 324
rect 2704 280 2804 324
rect -2804 -324 -2704 -280
rect -2600 -324 -2500 -280
rect -2396 -324 -2296 -280
rect -2192 -324 -2092 -280
rect -1988 -324 -1888 -280
rect -1784 -324 -1684 -280
rect -1580 -324 -1480 -280
rect -1376 -324 -1276 -280
rect -1172 -324 -1072 -280
rect -968 -324 -868 -280
rect -764 -324 -664 -280
rect -560 -324 -460 -280
rect -356 -324 -256 -280
rect -152 -324 -52 -280
rect 52 -324 152 -280
rect 256 -324 356 -280
rect 460 -324 560 -280
rect 664 -324 764 -280
rect 868 -324 968 -280
rect 1072 -324 1172 -280
rect 1276 -324 1376 -280
rect 1480 -324 1580 -280
rect 1684 -324 1784 -280
rect 1888 -324 1988 -280
rect 2092 -324 2192 -280
rect 2296 -324 2396 -280
rect 2500 -324 2600 -280
rect 2704 -324 2804 -280
<< metal1 >>
rect -2879 267 -2833 278
rect -2879 -278 -2833 -267
rect -2675 267 -2629 278
rect -2675 -278 -2629 -267
rect -2471 267 -2425 278
rect -2471 -278 -2425 -267
rect -2267 267 -2221 278
rect -2267 -278 -2221 -267
rect -2063 267 -2017 278
rect -2063 -278 -2017 -267
rect -1859 267 -1813 278
rect -1859 -278 -1813 -267
rect -1655 267 -1609 278
rect -1655 -278 -1609 -267
rect -1451 267 -1405 278
rect -1451 -278 -1405 -267
rect -1247 267 -1201 278
rect -1247 -278 -1201 -267
rect -1043 267 -997 278
rect -1043 -278 -997 -267
rect -839 267 -793 278
rect -839 -278 -793 -267
rect -635 267 -589 278
rect -635 -278 -589 -267
rect -431 267 -385 278
rect -431 -278 -385 -267
rect -227 267 -181 278
rect -227 -278 -181 -267
rect -23 267 23 278
rect -23 -278 23 -267
rect 181 267 227 278
rect 181 -278 227 -267
rect 385 267 431 278
rect 385 -278 431 -267
rect 589 267 635 278
rect 589 -278 635 -267
rect 793 267 839 278
rect 793 -278 839 -267
rect 997 267 1043 278
rect 997 -278 1043 -267
rect 1201 267 1247 278
rect 1201 -278 1247 -267
rect 1405 267 1451 278
rect 1405 -278 1451 -267
rect 1609 267 1655 278
rect 1609 -278 1655 -267
rect 1813 267 1859 278
rect 1813 -278 1859 -267
rect 2017 267 2063 278
rect 2017 -278 2063 -267
rect 2221 267 2267 278
rect 2221 -278 2267 -267
rect 2425 267 2471 278
rect 2425 -278 2471 -267
rect 2629 267 2675 278
rect 2629 -278 2675 -267
rect 2833 267 2879 278
rect 2833 -278 2879 -267
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 2.8 l 0.5 m 1 nf 28 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
