magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2245 -5495 2245 5495
<< psubdiff >>
rect -245 3473 245 3495
rect -245 -3473 -223 3473
rect 223 -3473 245 3473
rect -245 -3495 245 -3473
<< psubdiffcont >>
rect -223 -3473 223 3473
<< metal1 >>
rect -234 3473 234 3484
rect -234 -3473 -223 3473
rect 223 -3473 234 3473
rect -234 -3484 234 -3473
<< end >>
