* NGSPICE file created from DAC_12_Bit.ext - technology: gf180mcuC

.subckt nmos_3p3_AGPLV7 a_n138_n60# a_50_n60# a_n50_n104# VSUBS
X0 a_50_n60# a_n50_n104# a_n138_n60# VSUBS nfet_03v3 ad=0.264p pd=2.08u as=0.264p ps=2.08u w=0.6u l=0.5u
.ends

.subckt nmos_3p3_AQEADK a_n138_n60# a_50_n60# a_n50_n104# VSUBS
X0 a_50_n60# a_n50_n104# a_n138_n60# VSUBS nfet_03v3 ad=0.264p pd=2.08u as=0.264p ps=2.08u w=0.6u l=0.5u
.ends

.subckt MSB_Unit_Cell_p2 m1_34_n336# a_316_n480# a_51_258# a_316_26# m1_23_6# a_3095_69#
+ VSUBS
Xnmos_3p3_AGPLV7_5 m1_34_n336# a_3095_69# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_6 a_3095_69# m1_23_6# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_7 m1_23_6# a_3095_69# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_8 a_3095_69# m1_34_n336# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_9 m1_34_n336# a_3095_69# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AQEADK_0 a_3095_69# m1_34_n336# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_1 m1_23_6# a_3095_69# a_51_258# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_2 a_3095_69# m1_34_n336# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_4 a_3095_69# m1_23_6# a_51_258# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_3 m1_34_n336# a_3095_69# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_5 m1_23_6# a_3095_69# a_51_258# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_10 a_3095_69# m1_23_6# a_51_258# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_6 a_3095_69# m1_34_n336# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_11 m1_34_n336# a_3095_69# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_7 m1_34_n336# a_3095_69# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_12 a_3095_69# m1_23_6# a_51_258# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_8 a_3095_69# m1_23_6# a_51_258# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_13 m1_23_6# a_3095_69# a_51_258# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_9 m1_23_6# a_3095_69# a_51_258# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_15 m1_34_n336# a_3095_69# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_14 a_3095_69# m1_34_n336# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AGPLV7_10 a_3095_69# m1_23_6# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_12 a_3095_69# m1_23_6# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_11 m1_23_6# a_3095_69# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_13 m1_34_n336# a_3095_69# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_14 m1_23_6# a_3095_69# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_15 a_3095_69# m1_34_n336# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_0 a_3095_69# m1_34_n336# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_1 m1_34_n336# a_3095_69# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_2 a_3095_69# m1_23_6# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_3 m1_23_6# a_3095_69# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_4 a_3095_69# m1_34_n336# a_316_26# VSUBS nmos_3p3_AGPLV7
.ends

.subckt pmos_3p3_M8RWPS a_n28_n94# w_n202_n180# a_n116_n50# a_28_n50#
X0 a_28_n50# a_n28_n94# a_n116_n50# w_n202_n180# pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
.ends

.subckt nmos_3p3_HZS5UA a_n28_n94# a_n116_n50# a_28_n50# VSUBS
X0 a_28_n50# a_n28_n94# a_n116_n50# VSUBS nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
.ends

.subckt NAND VDD VSS B A OUT SD
Xpmos_3p3_M8RWPS_0 A VDD VDD OUT pmos_3p3_M8RWPS
Xpmos_3p3_M8RWPS_1 B VDD VDD OUT pmos_3p3_M8RWPS
Xnmos_3p3_HZS5UA_0 A SD OUT VSS nmos_3p3_HZS5UA
Xnmos_3p3_HZS5UA_1 B VSS SD VSS nmos_3p3_HZS5UA
.ends

.subckt Local_Enc Q QB Ci Ri Ri-1 VDD VSS
XNAND_0 VDD VSS Ri-1 Ri-1 NAND_1/B NAND_0/SD NAND
XNAND_1 VDD VSS NAND_1/B NAND_1/B NAND_5/B NAND_1/SD NAND
XNAND_2 VDD VSS Ci Ci NAND_6/B NAND_2/SD NAND
XNAND_3 VDD VSS Ri Ri NAND_6/A NAND_3/SD NAND
XNAND_4 VDD VSS NAND_4/B Q QB NAND_4/SD NAND
XNAND_5 VDD VSS NAND_5/B NAND_5/A NAND_8/A NAND_5/SD NAND
XNAND_6 VDD VSS NAND_6/B NAND_6/A NAND_5/A NAND_6/SD NAND
XNAND_7 VDD VSS NAND_8/A NAND_8/A NAND_4/B NAND_7/SD NAND
XNAND_8 VDD VSS QB NAND_8/A Q NAND_8/SD NAND
.ends

.subckt nmos_3p3_LNPLVM a_2192_n120# a_3112_n164# a_n2296_n120# a_2092_n164# a_n968_n164#
+ a_1172_n120# a_n256_n120# a_n1988_n164# a_n1276_n120# a_1072_n164# a_1988_n120#
+ a_2908_n164# a_1888_n164# a_n460_n120# a_n2500_n120# a_n1480_n120# a_764_n120# a_664_n164#
+ a_n2092_n120# a_n3112_n120# a_n764_n164# a_n2804_n164# a_n1784_n164# a_n52_n120#
+ a_n1072_n120# a_2804_n120# a_1784_n120# a_356_n120# a_n868_n120# a_n2908_n120# a_2704_n164#
+ a_1684_n164# a_n1888_n120# a_256_n164# a_n2396_n164# a_n356_n164# a_560_n120# a_n1376_n164#
+ a_2396_n120# a_460_n164# a_2296_n164# a_1376_n120# a_n560_n164# a_1276_n164# a_n1580_n164#
+ a_n2600_n164# a_n3008_n164# a_2600_n120# a_1580_n120# a_3008_n120# a_152_n120# a_n664_n120#
+ a_n2704_n120# a_2500_n164# a_1480_n164# a_n1684_n120# a_968_n120# a_52_n164# a_n2192_n164#
+ a_n3212_n164# a_868_n164# a_n152_n164# a_3212_n120# a_n3300_n120# a_n1172_n164#
+ VSUBS
X0 a_n460_n120# a_n560_n164# a_n664_n120# VSUBS nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X1 a_n52_n120# a_n152_n164# a_n256_n120# VSUBS nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X2 a_n1480_n120# a_n1580_n164# a_n1684_n120# VSUBS nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X3 a_n1072_n120# a_n1172_n164# a_n1276_n120# VSUBS nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X4 a_1172_n120# a_1072_n164# a_968_n120# VSUBS nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X5 a_n868_n120# a_n968_n164# a_n1072_n120# VSUBS nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X6 a_n1888_n120# a_n1988_n164# a_n2092_n120# VSUBS nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X7 a_1988_n120# a_1888_n164# a_1784_n120# VSUBS nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X8 a_1580_n120# a_1480_n164# a_1376_n120# VSUBS nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X9 a_968_n120# a_868_n164# a_764_n120# VSUBS nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X10 a_3008_n120# a_2908_n164# a_2804_n120# VSUBS nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X11 a_n2500_n120# a_n2600_n164# a_n2704_n120# VSUBS nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X12 a_n2092_n120# a_n2192_n164# a_n2296_n120# VSUBS nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X13 a_560_n120# a_460_n164# a_356_n120# VSUBS nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X14 a_2192_n120# a_2092_n164# a_1988_n120# VSUBS nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X15 a_2600_n120# a_2500_n164# a_2396_n120# VSUBS nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X16 a_n3112_n120# a_n3212_n164# a_n3300_n120# VSUBS nfet_03v3 ad=0.312p pd=1.72u as=0.528p ps=3.28u w=1.2u l=0.5u
X17 a_3212_n120# a_3112_n164# a_3008_n120# VSUBS nfet_03v3 ad=0.528p pd=3.28u as=0.312p ps=1.72u w=1.2u l=0.5u
X18 a_n256_n120# a_n356_n164# a_n460_n120# VSUBS nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X19 a_n1276_n120# a_n1376_n164# a_n1480_n120# VSUBS nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X20 a_1376_n120# a_1276_n164# a_1172_n120# VSUBS nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X21 a_356_n120# a_256_n164# a_152_n120# VSUBS nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X22 a_n2908_n120# a_n3008_n164# a_n3112_n120# VSUBS nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X23 a_n664_n120# a_n764_n164# a_n868_n120# VSUBS nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X24 a_152_n120# a_52_n164# a_n52_n120# VSUBS nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X25 a_n1684_n120# a_n1784_n164# a_n1888_n120# VSUBS nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X26 a_1784_n120# a_1684_n164# a_1580_n120# VSUBS nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X27 a_764_n120# a_664_n164# a_560_n120# VSUBS nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X28 a_2804_n120# a_2704_n164# a_2600_n120# VSUBS nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X29 a_n2704_n120# a_n2804_n164# a_n2908_n120# VSUBS nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X30 a_n2296_n120# a_n2396_n164# a_n2500_n120# VSUBS nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X31 a_2396_n120# a_2296_n164# a_2192_n120# VSUBS nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
.ends

.subckt CM_MSB_V2 IM_T VSS OUT IM SD
Xnmos_3p3_LNPLVM_0 SD IM_T SD IM IM_T VSS SD IM VSS IM VSS IM IM VSS OUT SD OUT IM_T
+ VSS SD IM_T IM IM_T OUT SD VSS SD VSS OUT VSS IM IM_T SD IM IM_T IM SD IM OUT IM
+ IM_T SD IM IM IM_T IM_T IM SD OUT SD SD SD SD IM_T IM_T OUT SD IM_T IM IM_T IM_T
+ IM_T OUT OUT IM VSS nmos_3p3_LNPLVM
Xnmos_3p3_LNPLVM_1 SD IM SD IM_T IM OUT SD IM_T OUT IM_T OUT IM_T IM_T OUT VSS SD
+ VSS IM OUT SD IM IM_T IM VSS SD OUT SD OUT VSS OUT IM_T IM SD IM_T IM IM_T SD IM_T
+ VSS IM_T IM SD IM_T IM_T IM IM IM_T SD VSS SD SD SD SD IM IM VSS SD IM IM_T IM IM
+ IM VSS VSS IM_T VSS nmos_3p3_LNPLVM
.ends

.subckt MSB_Unit_Cell IM Ri Ci VDD QB Q OUT OUT+ OUT- SD Ri-1 IM_T VSS
XMSB_Unit_Cell_p2_3 OUT- Q Q QB OUT+ OUT VSS MSB_Unit_Cell_p2
XLocal_Enc_0 Q QB Ci Ri Ri-1 VDD VSS Local_Enc
XCM_MSB_V2_0 IM_T VSS OUT IM SD CM_MSB_V2
XMSB_Unit_Cell_p2_0 OUT- Q Q QB OUT+ OUT VSS MSB_Unit_Cell_p2
XMSB_Unit_Cell_p2_1 OUT- Q Q QB OUT+ OUT VSS MSB_Unit_Cell_p2
XMSB_Unit_Cell_p2_2 OUT- Q Q QB OUT+ OUT VSS MSB_Unit_Cell_p2
.ends

.subckt nmos_3p3_H9QVWA a_n120_n36# a_28_n25# a_n28_n69# VSUBS
X0 a_28_n25# a_n28_n69# a_n120_n36# VSUBS nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
.ends

.subckt Inverter VDD VSS IN OUT
Xnmos_3p3_H9QVWA_0 VSS OUT IN VSS nmos_3p3_H9QVWA
Xpmos_3p3_M8RWPS_0 IN VDD VDD OUT pmos_3p3_M8RWPS
.ends

.subckt INV_BUFF IN SD1 OUT VDD VSS
XInverter_0 VDD VSS SD1 OUT Inverter
XInverter_1 VDD VSS IN SD1 Inverter
.ends

.subckt nmos_3p3_9NPLV7 a_3008_n60# a_764_n60# a_n664_n60# a_2192_n60# a_n2092_n60#
+ a_664_n104# a_2804_n60# a_n2704_n60# a_560_n60# a_n460_n60# a_n764_n104# a_n2804_n104#
+ a_1988_n60# a_n1888_n60# a_n1784_n104# a_2600_n60# a_n2500_n60# a_2704_n104# a_1684_n104#
+ a_256_n104# a_1784_n60# a_n256_n60# a_n1684_n60# a_356_n60# a_n2396_n104# a_n356_n104#
+ a_460_n104# a_n1376_n104# a_1580_n60# a_n1480_n60# a_2296_n104# a_152_n60# a_1276_n104#
+ a_n560_n104# a_n2600_n104# a_n1580_n104# a_n3008_n104# a_n52_n60# a_2500_n104# a_1376_n60#
+ a_n1276_n60# a_1480_n104# a_n3212_n104# a_52_n104# a_n2192_n104# a_868_n104# a_n152_n104#
+ a_1172_n60# a_n1072_n60# a_n1172_n104# a_3112_n104# a_2092_n104# a_n968_n104# a_n1988_n104#
+ a_3212_n60# a_n3112_n60# a_n3300_n60# a_1072_n104# a_968_n60# a_n868_n60# a_2908_n104#
+ a_2396_n60# a_n2296_n60# a_1888_n104# a_n2908_n60# VSUBS
X0 a_n2908_n60# a_n3008_n104# a_n3112_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X1 a_n256_n60# a_n356_n104# a_n460_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X2 a_1376_n60# a_1276_n104# a_1172_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X3 a_n3112_n60# a_n3212_n104# a_n3300_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X4 a_1580_n60# a_1480_n104# a_1376_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X5 a_n2704_n60# a_n2804_n104# a_n2908_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X6 a_n460_n60# a_n560_n104# a_n664_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X7 a_2192_n60# a_2092_n104# a_1988_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X8 a_n664_n60# a_n764_n104# a_n868_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X9 a_1784_n60# a_1684_n104# a_1580_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X10 a_2396_n60# a_2296_n104# a_2192_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X11 a_n1072_n60# a_n1172_n104# a_n1276_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X12 a_n868_n60# a_n968_n104# a_n1072_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X13 a_1988_n60# a_1888_n104# a_1784_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X14 a_356_n60# a_256_n104# a_152_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X15 a_n1276_n60# a_n1376_n104# a_n1480_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X16 a_560_n60# a_460_n104# a_356_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X17 a_n1480_n60# a_n1580_n104# a_n1684_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X18 a_n2092_n60# a_n2192_n104# a_n2296_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X19 a_2600_n60# a_2500_n104# a_2396_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X20 a_764_n60# a_664_n104# a_560_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X21 a_n1684_n60# a_n1784_n104# a_n1888_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X22 a_3212_n60# a_3112_n104# a_3008_n60# VSUBS nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X23 a_152_n60# a_52_n104# a_n52_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X24 a_n2296_n60# a_n2396_n104# a_n2500_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X25 a_2804_n60# a_2704_n104# a_2600_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X26 a_n1888_n60# a_n1988_n104# a_n2092_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X27 a_968_n60# a_868_n104# a_764_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X28 a_n2500_n60# a_n2600_n104# a_n2704_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X29 a_3008_n60# a_2908_n104# a_2804_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X30 a_n52_n60# a_n152_n104# a_n256_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X31 a_1172_n60# a_1072_n104# a_968_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
.ends

.subckt pmos_3p3_DVR9E7 a_3008_n60# a_764_n60# a_n664_n60# a_2192_n60# a_n2092_n60#
+ a_664_n104# w_n3386_n190# a_2804_n60# a_n2704_n60# a_560_n60# a_n460_n60# a_n764_n104#
+ a_n2804_n104# a_1988_n60# a_n1888_n60# a_n1784_n104# a_2600_n60# a_n2500_n60# a_2704_n104#
+ a_1684_n104# a_256_n104# a_1784_n60# a_n256_n60# a_n1684_n60# a_356_n60# a_n2396_n104#
+ a_n356_n104# a_460_n104# a_n1376_n104# a_1580_n60# a_n1480_n60# a_2296_n104# a_152_n60#
+ a_1276_n104# a_n560_n104# a_n2600_n104# a_n1580_n104# a_n3008_n104# a_n52_n60# a_2500_n104#
+ a_1376_n60# a_n1276_n60# a_1480_n104# a_n3212_n104# a_52_n104# a_n2192_n104# a_868_n104#
+ a_n152_n104# a_1172_n60# a_n1072_n60# a_n1172_n104# a_3112_n104# a_2092_n104# a_n968_n104#
+ a_n1988_n104# a_3212_n60# a_n3112_n60# a_n3300_n60# a_1072_n104# a_968_n60# a_n868_n60#
+ a_2908_n104# a_2396_n60# a_n2296_n60# a_1888_n104# a_n2908_n60#
X0 a_n2908_n60# a_n3008_n104# a_n3112_n60# w_n3386_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X1 a_n256_n60# a_n356_n104# a_n460_n60# w_n3386_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X2 a_1376_n60# a_1276_n104# a_1172_n60# w_n3386_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X3 a_n3112_n60# a_n3212_n104# a_n3300_n60# w_n3386_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X4 a_1580_n60# a_1480_n104# a_1376_n60# w_n3386_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X5 a_n2704_n60# a_n2804_n104# a_n2908_n60# w_n3386_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X6 a_n460_n60# a_n560_n104# a_n664_n60# w_n3386_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X7 a_2192_n60# a_2092_n104# a_1988_n60# w_n3386_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X8 a_n664_n60# a_n764_n104# a_n868_n60# w_n3386_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X9 a_1784_n60# a_1684_n104# a_1580_n60# w_n3386_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X10 a_2396_n60# a_2296_n104# a_2192_n60# w_n3386_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X11 a_n1072_n60# a_n1172_n104# a_n1276_n60# w_n3386_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X12 a_n868_n60# a_n968_n104# a_n1072_n60# w_n3386_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X13 a_1988_n60# a_1888_n104# a_1784_n60# w_n3386_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X14 a_356_n60# a_256_n104# a_152_n60# w_n3386_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X15 a_n1276_n60# a_n1376_n104# a_n1480_n60# w_n3386_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X16 a_560_n60# a_460_n104# a_356_n60# w_n3386_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X17 a_n1480_n60# a_n1580_n104# a_n1684_n60# w_n3386_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X18 a_n2092_n60# a_n2192_n104# a_n2296_n60# w_n3386_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X19 a_2600_n60# a_2500_n104# a_2396_n60# w_n3386_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X20 a_764_n60# a_664_n104# a_560_n60# w_n3386_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X21 a_n1684_n60# a_n1784_n104# a_n1888_n60# w_n3386_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X22 a_3212_n60# a_3112_n104# a_3008_n60# w_n3386_n190# pfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X23 a_n2296_n60# a_n2396_n104# a_n2500_n60# w_n3386_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X24 a_152_n60# a_52_n104# a_n52_n60# w_n3386_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X25 a_2804_n60# a_2704_n104# a_2600_n60# w_n3386_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X26 a_n1888_n60# a_n1988_n104# a_n2092_n60# w_n3386_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X27 a_968_n60# a_868_n104# a_764_n60# w_n3386_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X28 a_n2500_n60# a_n2600_n104# a_n2704_n60# w_n3386_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X29 a_3008_n60# a_2908_n104# a_2804_n60# w_n3386_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X30 a_n52_n60# a_n152_n104# a_n256_n60# w_n3386_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X31 a_1172_n60# a_1072_n104# a_968_n60# w_n3386_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
.ends

.subckt CM_32_C SD0_1 G1_2 G1_1 SD2_0 G0_1 G0_2 VSS VDD G3_1 G3_2
Xnmos_3p3_9NPLV7_0 G3_1 G3_2 G3_1 G3_1 VSS G3_2 VSS G3_1 G3_1 VSS G3_2 G3_1 VSS G3_1
+ G3_2 G3_1 G3_2 G3_1 G3_2 G3_1 G3_1 G3_1 G3_2 VSS G3_2 G3_1 G3_1 G3_1 G3_2 G3_1 G3_2
+ G3_1 G3_1 G3_1 G3_2 G3_2 G3_1 G3_2 G3_2 G3_1 VSS G3_2 G3_2 G3_2 G3_1 G3_2 G3_2 VSS
+ G3_1 G3_1 G3_2 G3_1 G3_2 G3_1 G3_2 G3_1 G3_2 G3_1 G3_1 G3_2 G3_1 G3_2 G3_1 G3_1
+ VSS VSS nmos_3p3_9NPLV7
Xnmos_3p3_9NPLV7_1 SD0_1 VSS SD0_1 SD0_1 G1_1 G0_1 G1_1 SD0_1 SD0_1 G1_1 G0_1 G0_2
+ G1_1 SD0_1 G0_1 SD0_1 VSS G0_2 G0_1 G0_2 SD0_1 SD0_1 VSS G1_1 G0_1 G0_2 G0_2 G0_2
+ VSS SD0_1 G0_1 SD0_1 G0_2 G0_2 G0_1 G0_1 G0_2 VSS G0_1 SD0_1 G1_1 G0_1 G0_1 G0_1
+ G0_2 G0_1 G0_1 G1_1 SD0_1 G0_2 G0_1 G0_2 G0_1 G0_2 VSS SD0_1 VSS G0_2 SD0_1 VSS
+ G0_2 VSS SD0_1 G0_2 G1_1 VSS nmos_3p3_9NPLV7
Xnmos_3p3_9NPLV7_2 SD0_1 G1_1 SD0_1 SD0_1 VSS G0_2 VSS SD0_1 SD0_1 VSS G0_2 G0_1 VSS
+ SD0_1 G0_2 SD0_1 G1_1 G0_1 G0_2 G0_1 SD0_1 SD0_1 G1_1 VSS G0_2 G0_1 G0_1 G0_1 G1_1
+ SD0_1 G0_2 SD0_1 G0_1 G0_1 G0_2 G0_2 G0_1 G1_1 G0_2 SD0_1 VSS G0_2 G0_2 G0_2 G0_1
+ G0_2 G0_2 VSS SD0_1 G0_1 G0_2 G0_1 G0_2 G0_1 G1_1 SD0_1 G1_1 G0_1 SD0_1 G1_1 G0_1
+ G1_1 SD0_1 G0_1 VSS VSS nmos_3p3_9NPLV7
Xnmos_3p3_9NPLV7_3 G3_1 VSS G3_1 G3_1 G3_2 G3_1 G3_2 G3_1 G3_1 G3_2 G3_1 G3_2 G3_2
+ G3_1 G3_1 G3_1 VSS G3_2 G3_1 G3_2 G3_1 G3_1 VSS G3_2 G3_1 G3_2 G3_2 G3_2 VSS G3_1
+ G3_1 G3_1 G3_2 G3_2 G3_1 G3_1 G3_2 VSS G3_1 G3_1 G3_2 G3_1 G3_1 G3_1 G3_2 G3_1 G3_1
+ G3_2 G3_1 G3_2 G3_1 G3_2 G3_1 G3_2 VSS G3_1 VSS G3_2 G3_1 VSS G3_2 VSS G3_1 G3_2
+ G3_2 VSS nmos_3p3_9NPLV7
Xpmos_3p3_DVR9E7_0 G1_2 VDD G1_2 G1_2 G1_1 G1_2 VDD G1_1 G1_2 G1_2 G1_1 G1_2 G1_1
+ G1_1 G1_2 G1_2 G1_2 VDD G1_1 G1_2 G1_1 G1_2 G1_2 VDD G1_1 G1_2 G1_1 G1_1 G1_1 VDD
+ G1_2 G1_2 G1_2 G1_1 G1_1 G1_2 G1_2 G1_1 VDD G1_2 G1_2 G1_1 G1_2 G1_2 G1_2 G1_1 G1_2
+ G1_2 G1_1 G1_2 G1_1 G1_2 G1_1 G1_2 G1_1 VDD G1_2 VDD G1_1 G1_2 VDD G1_1 VDD G1_2
+ G1_1 G1_1 pmos_3p3_DVR9E7
Xpmos_3p3_DVR9E7_1 SD2_0 VDD SD2_0 SD2_0 G3_2 G1_2 VDD G3_2 SD2_0 SD2_0 G3_2 G1_2
+ G1_1 G3_2 SD2_0 G1_2 SD2_0 VDD G1_1 G1_2 G1_1 SD2_0 SD2_0 VDD G3_2 G1_2 G1_1 G1_1
+ G1_1 VDD SD2_0 G1_2 SD2_0 G1_1 G1_1 G1_2 G1_2 G1_1 VDD G1_2 SD2_0 G3_2 G1_2 G1_2
+ G1_2 G1_1 G1_2 G1_2 G3_2 SD2_0 G1_1 G1_2 G1_1 G1_2 G1_1 VDD SD2_0 VDD G1_1 SD2_0
+ VDD G1_1 VDD SD2_0 G1_1 G3_2 pmos_3p3_DVR9E7
Xpmos_3p3_DVR9E7_2 G1_2 G1_1 G1_2 G1_2 VDD G1_1 VDD VDD G1_2 G1_2 VDD G1_1 G1_2 VDD
+ G1_2 G1_1 G1_2 G1_1 G1_2 G1_1 G1_2 G1_2 G1_2 G1_1 VDD G1_1 G1_2 G1_2 G1_2 G1_1 G1_2
+ G1_1 G1_2 G1_2 G1_2 G1_1 G1_1 G1_2 G1_1 G1_1 G1_2 VDD G1_1 G1_1 G1_1 G1_2 G1_1 G1_1
+ VDD G1_2 G1_2 G1_1 G1_2 G1_1 G1_2 G1_1 G1_2 G1_1 G1_2 G1_2 G1_1 G1_2 G1_1 G1_2 G1_2
+ VDD pmos_3p3_DVR9E7
Xpmos_3p3_DVR9E7_3 SD2_0 G3_2 SD2_0 SD2_0 VDD G1_1 VDD VDD SD2_0 SD2_0 VDD G1_1 G1_2
+ VDD SD2_0 G1_1 SD2_0 G3_2 G1_2 G1_1 G1_2 SD2_0 SD2_0 G3_2 VDD G1_1 G1_2 G1_2 G1_2
+ G3_2 SD2_0 G1_1 SD2_0 G1_2 G1_2 G1_1 G1_1 G1_2 G3_2 G1_1 SD2_0 VDD G1_1 G1_1 G1_1
+ G1_2 G1_1 G1_1 VDD SD2_0 G1_2 G1_1 G1_2 G1_1 G1_2 G3_2 SD2_0 G3_2 G1_2 SD2_0 G3_2
+ G1_2 G3_2 SD2_0 G1_2 VDD pmos_3p3_DVR9E7
.ends

.subckt pmos_3p3_MGRWPS a_n52_n50# a_n196_n50# a_52_n94# a_108_n50# a_n108_n94# w_n282_n180#
X0 a_108_n50# a_52_n94# a_n52_n50# w_n282_n180# pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X1 a_n52_n50# a_n108_n94# a_n196_n50# w_n282_n180# pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
.ends

.subckt OR A B VSS VDD OUT SD1 SD2
Xnmos_3p3_H9QVWA_0 VSS SD2 A VSS nmos_3p3_H9QVWA
Xpmos_3p3_MGRWPS_0 SD2 SD1 A SD1 A VDD pmos_3p3_MGRWPS
Xnmos_3p3_H9QVWA_1 VSS SD2 B VSS nmos_3p3_H9QVWA
Xpmos_3p3_MGRWPS_1 SD1 VDD B VDD B VDD pmos_3p3_MGRWPS
XInverter_0 VDD VSS SD2 OUT Inverter
.ends

.subckt AND VDD VSS OUT A B SD1 SD2
XInverter_0 VDD VSS SD2 OUT Inverter
Xpmos_3p3_M8RWPS_0 B VDD SD2 VDD pmos_3p3_M8RWPS
Xpmos_3p3_M8RWPS_1 A VDD VDD SD2 pmos_3p3_M8RWPS
Xnmos_3p3_HZS5UA_0 A VSS SD1 VSS nmos_3p3_HZS5UA
Xnmos_3p3_HZS5UA_1 B SD1 SD2 VSS nmos_3p3_HZS5UA
.ends

.subckt therm_Dec B1 VDD D1 D2 D4 D3 D5 D6 D7 B3 B2 VSS
XOR_4 B1 B2 VSS VDD OR_3/B OR_4/SD1 OR_4/SD2 OR
XINV_BUFF_0 AND_0/OUT INV_BUFF_0/SD1 D1 VDD VSS INV_BUFF
XINV_BUFF_1 AND_2/OUT INV_BUFF_1/SD1 D2 VDD VSS INV_BUFF
XINV_BUFF_2 AND_3/OUT INV_BUFF_2/SD1 D3 VDD VSS INV_BUFF
XINV_BUFF_3 B1 INV_BUFF_3/SD1 D4 VDD VSS INV_BUFF
XINV_BUFF_4 OR_1/OUT INV_BUFF_4/SD1 D5 VDD VSS INV_BUFF
XAND_0 VDD VSS AND_0/OUT B3 AND_0/B AND_0/SD1 AND_0/SD2 AND
XINV_BUFF_5 OR_2/OUT INV_BUFF_5/SD1 D6 VDD VSS INV_BUFF
XAND_1 VDD VSS AND_0/B B1 B2 AND_1/SD1 AND_1/SD2 AND
XINV_BUFF_6 OR_3/OUT INV_BUFF_6/SD1 D7 VDD VSS INV_BUFF
XAND_2 VDD VSS AND_2/OUT B1 B2 AND_2/SD1 AND_2/SD2 AND
XAND_3 VDD VSS AND_3/OUT B1 AND_3/B AND_3/SD1 AND_3/SD2 AND
XAND_4 VDD VSS OR_1/B B2 B3 AND_4/SD1 AND_4/SD2 AND
XOR_0 B2 B3 VSS VDD AND_3/B OR_0/SD1 OR_0/SD2 OR
XOR_1 B1 OR_1/B VSS VDD OR_1/OUT OR_1/SD1 OR_1/SD2 OR
XOR_2 B1 B2 VSS VDD OR_2/OUT OR_2/SD1 OR_2/SD2 OR
XOR_3 B3 OR_3/B VSS VDD OR_3/OUT OR_3/SD1 OR_3/SD2 OR
.ends

.subckt nmos_3p3_MGEA3B a_n138_n60# a_50_n60# a_n50_n104# VSUBS
X0 a_50_n60# a_n50_n104# a_n138_n60# VSUBS nfet_03v3 ad=0.264p pd=2.08u as=0.264p ps=2.08u w=0.6u l=0.5u
.ends

.subckt nmos_3p3_MGEAJ7 a_50_n30# a_n50_n74# a_n142_n36# VSUBS
X0 a_50_n30# a_n50_n74# a_n142_n36# VSUBS nfet_03v3 ad=0.16p pd=1.64u as=0.16p ps=1.64u w=0.3u l=0.5u
.ends

.subckt pmos_3p3_M8LTNG a_n120_n36# a_28_n22# a_n28_n66# w_n206_n159#
X0 a_28_n22# a_n28_n66# a_n120_n36# w_n206_n159# pfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
.ends

.subckt nmos_3p3_DDNVWA a_n120_n36# a_28_n22# a_n28_n66# VSUBS
X0 a_28_n22# a_n28_n66# a_n120_n36# VSUBS nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
.ends

.subckt Balance_Inverter VDD VSS OUT OUT_B VIN
Xpmos_3p3_M8LTNG_0 OUT VDD OUT_B VDD pmos_3p3_M8LTNG
Xpmos_3p3_M8LTNG_1 VDD OUT_B OUT VDD pmos_3p3_M8LTNG
XInverter_0 VDD VSS VIN Inverter_0/OUT Inverter
Xnmos_3p3_DDNVWA_0 OUT VSS Inverter_0/OUT VSS nmos_3p3_DDNVWA
Xnmos_3p3_DDNVWA_1 VSS OUT_B VIN VSS nmos_3p3_DDNVWA
.ends

.subckt CM_32 VSS G0_2 G0_1 VDD G1_2 G1_1 SD2_0 G3_2 G3_1 SD0_1
Xnmos_3p3_9NPLV7_0 G3_1 G3_2 G3_1 G3_1 VSS G3_2 VSS G3_1 G3_1 VSS G3_2 G3_1 VSS G3_1
+ G3_2 G3_1 G3_2 G3_1 G3_2 G3_1 G3_1 G3_1 G3_2 VSS G3_2 G3_1 G3_1 G3_1 G3_2 G3_1 G3_2
+ G3_1 G3_1 G3_1 G3_2 G3_2 G3_1 G3_2 G3_2 G3_1 VSS G3_2 G3_2 G3_2 G3_1 G3_2 G3_2 VSS
+ G3_1 G3_1 G3_2 G3_1 G3_2 G3_1 G3_2 G3_1 G3_2 G3_1 G3_1 G3_2 G3_1 G3_2 G3_1 G3_1
+ VSS VSS nmos_3p3_9NPLV7
Xnmos_3p3_9NPLV7_1 SD0_1 VSS SD0_1 SD0_1 G1_1 G0_1 G1_1 SD0_1 SD0_1 G1_1 G0_1 G0_2
+ G1_1 SD0_1 G0_1 SD0_1 VSS G0_2 G0_1 G0_2 SD0_1 SD0_1 VSS G1_1 G0_1 G0_2 G0_2 G0_2
+ VSS SD0_1 G0_1 SD0_1 G0_2 G0_2 G0_1 G0_1 G0_2 VSS G0_1 SD0_1 G1_1 G0_1 G0_1 G0_1
+ G0_2 G0_1 G0_1 G1_1 SD0_1 G0_2 G0_1 G0_2 G0_1 G0_2 VSS SD0_1 VSS G0_2 SD0_1 VSS
+ G0_2 VSS SD0_1 G0_2 G1_1 VSS nmos_3p3_9NPLV7
Xnmos_3p3_9NPLV7_2 SD0_1 G1_1 SD0_1 SD0_1 VSS G0_2 VSS SD0_1 SD0_1 VSS G0_2 G0_1 VSS
+ SD0_1 G0_2 SD0_1 G1_1 G0_1 G0_2 G0_1 SD0_1 SD0_1 G1_1 VSS G0_2 G0_1 G0_1 G0_1 G1_1
+ SD0_1 G0_2 SD0_1 G0_1 G0_1 G0_2 G0_2 G0_1 G1_1 G0_2 SD0_1 VSS G0_2 G0_2 G0_2 G0_1
+ G0_2 G0_2 VSS SD0_1 G0_1 G0_2 G0_1 G0_2 G0_1 G1_1 SD0_1 G1_1 G0_1 SD0_1 G1_1 G0_1
+ G1_1 SD0_1 G0_1 VSS VSS nmos_3p3_9NPLV7
Xnmos_3p3_9NPLV7_3 G3_1 VSS G3_1 G3_1 G3_2 G3_1 G3_2 G3_1 G3_1 G3_2 G3_1 G3_2 G3_2
+ G3_1 G3_1 G3_1 VSS G3_2 G3_1 G3_2 G3_1 G3_1 VSS G3_2 G3_1 G3_2 G3_2 G3_2 VSS G3_1
+ G3_1 G3_1 G3_2 G3_2 G3_1 G3_1 G3_2 VSS G3_1 G3_1 G3_2 G3_1 G3_1 G3_1 G3_2 G3_1 G3_1
+ G3_2 G3_1 G3_2 G3_1 G3_2 G3_1 G3_2 VSS G3_1 VSS G3_2 G3_1 VSS G3_2 VSS G3_1 G3_2
+ G3_2 VSS nmos_3p3_9NPLV7
Xpmos_3p3_DVR9E7_0 G1_2 VDD G1_2 G1_2 G1_1 G1_2 VDD G1_1 G1_2 G1_2 G1_1 G1_2 G1_1
+ G1_1 G1_2 G1_2 G1_2 VDD G1_1 G1_2 G1_1 G1_2 G1_2 VDD G1_1 G1_2 G1_1 G1_1 G1_1 VDD
+ G1_2 G1_2 G1_2 G1_1 G1_1 G1_2 G1_2 G1_1 VDD G1_2 G1_2 G1_1 G1_2 G1_2 G1_2 G1_1 G1_2
+ G1_2 G1_1 G1_2 G1_1 G1_2 G1_1 G1_2 G1_1 VDD G1_2 VDD G1_1 G1_2 VDD G1_1 VDD G1_2
+ G1_1 G1_1 pmos_3p3_DVR9E7
Xpmos_3p3_DVR9E7_1 SD2_0 VDD SD2_0 SD2_0 G3_2 G1_2 VDD G3_2 SD2_0 SD2_0 G3_2 G1_2
+ G1_1 G3_2 SD2_0 G1_2 SD2_0 VDD G1_1 G1_2 G1_1 SD2_0 SD2_0 VDD G3_2 G1_2 G1_1 G1_1
+ G1_1 VDD SD2_0 G1_2 SD2_0 G1_1 G1_1 G1_2 G1_2 G1_1 VDD G1_2 SD2_0 G3_2 G1_2 G1_2
+ G1_2 G1_1 G1_2 G1_2 G3_2 SD2_0 G1_1 G1_2 G1_1 G1_2 G1_1 VDD SD2_0 VDD G1_1 SD2_0
+ VDD G1_1 VDD SD2_0 G1_1 G3_2 pmos_3p3_DVR9E7
Xpmos_3p3_DVR9E7_2 G1_2 G1_1 G1_2 G1_2 VDD G1_1 VDD VDD G1_2 G1_2 VDD G1_1 G1_2 VDD
+ G1_2 G1_1 G1_2 G1_1 G1_2 G1_1 G1_2 G1_2 G1_2 G1_1 VDD G1_1 G1_2 G1_2 G1_2 G1_1 G1_2
+ G1_1 G1_2 G1_2 G1_2 G1_1 G1_1 G1_2 G1_1 G1_1 G1_2 VDD G1_1 G1_1 G1_1 G1_2 G1_1 G1_1
+ VDD G1_2 G1_2 G1_1 G1_2 G1_1 G1_2 G1_1 G1_2 G1_1 G1_2 G1_2 G1_1 G1_2 G1_1 G1_2 G1_2
+ VDD pmos_3p3_DVR9E7
Xpmos_3p3_DVR9E7_3 SD2_0 G3_2 SD2_0 SD2_0 VDD G1_1 VDD VDD SD2_0 SD2_0 VDD G1_1 G1_2
+ VDD SD2_0 G1_1 SD2_0 G3_2 G1_2 G1_1 G1_2 SD2_0 SD2_0 G3_2 VDD G1_1 G1_2 G1_2 G1_2
+ G3_2 SD2_0 G1_1 SD2_0 G1_2 G1_2 G1_1 G1_1 G1_2 G3_2 G1_1 SD2_0 VDD G1_1 G1_1 G1_1
+ G1_2 G1_1 G1_1 VDD SD2_0 G1_2 G1_1 G1_2 G1_1 G1_2 G3_2 SD2_0 G3_2 G1_2 SD2_0 G3_2
+ G1_2 G3_2 SD2_0 G1_2 VDD pmos_3p3_DVR9E7
.ends

.subckt nmos_3p3_ECASTA a_n52_n200# a_n212_n200# a_108_n200# a_52_n244# a_n108_n244#
+ a_212_n244# a_268_n200# a_n268_n244# a_n356_n200# VSUBS
X0 a_108_n200# a_52_n244# a_n52_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_268_n200# a_212_n244# a_108_n200# VSUBS nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_n212_n200# a_n268_n244# a_n356_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.28u
X3 a_n52_n200# a_n108_n244# a_n212_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt nmos_3p3_AEBEG7 a_2988_n200# a_1228_n200# a_n52_n200# a_n852_n200# a_n428_n244#
+ a_n1012_n200# a_532_n244# a_n2772_n200# a_n1388_n244# a_588_n200# a_n1812_n200#
+ a_2292_n244# a_1332_n244# a_n2348_n244# a_2348_n200# a_1388_n200# a_n212_n200# a_n588_n244#
+ a_n1172_n200# a_n3092_n200# a_692_n244# a_n2132_n200# a_n1972_n200# a_n2932_n200#
+ a_1492_n244# a_n1548_n244# a_748_n200# a_2452_n244# a_n2508_n244# a_n372_n200# a_2508_n200#
+ a_1548_n200# a_n748_n244# a_n2292_n200# a_108_n200# a_n1332_n200# a_852_n244# a_52_n244#
+ a_n2668_n244# a_908_n200# a_2612_n244# a_1652_n244# a_n1708_n244# a_2668_n200# a_1708_n200#
+ a_n532_n200# a_n108_n244# a_212_n244# a_268_n200# a_n1492_n200# a_n2452_n200# a_n908_n244#
+ a_n1068_n244# a_n2028_n244# a_1012_n244# a_n1868_n244# a_1068_n200# a_2772_n244#
+ a_n2828_n244# a_2028_n200# a_1812_n244# a_2828_n200# a_1868_n200# a_n692_n200# a_n268_n244#
+ a_372_n244# a_n2188_n244# a_n1652_n200# a_n2612_n200# a_3092_n244# a_1172_n244#
+ a_n1228_n244# a_n3148_n244# a_428_n200# a_2132_n244# a_n2988_n244# a_3148_n200#
+ a_2188_n200# a_n3236_n200# a_2932_n244# a_1972_n244# VSUBS
X0 a_1548_n200# a_1492_n244# a_1388_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_n2612_n200# a_n2668_n244# a_n2772_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_588_n200# a_532_n244# a_428_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X3 a_1388_n200# a_1332_n244# a_1228_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X4 a_n2452_n200# a_n2508_n244# a_n2612_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X5 a_2508_n200# a_2452_n244# a_2348_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X6 a_n532_n200# a_n588_n244# a_n692_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X7 a_n372_n200# a_n428_n244# a_n532_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X8 a_n1332_n200# a_n1388_n244# a_n1492_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X9 a_n1172_n200# a_n1228_n244# a_n1332_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X10 a_108_n200# a_52_n244# a_n52_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X11 a_428_n200# a_372_n244# a_268_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X12 a_268_n200# a_212_n244# a_108_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X13 a_1228_n200# a_1172_n244# a_1068_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X14 a_n2292_n200# a_n2348_n244# a_n2452_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X15 a_1068_n200# a_1012_n244# a_908_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X16 a_2028_n200# a_1972_n244# a_1868_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X17 a_2348_n200# a_2292_n244# a_2188_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X18 a_1868_n200# a_1812_n244# a_1708_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X19 a_2188_n200# a_2132_n244# a_2028_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X20 a_n212_n200# a_n268_n244# a_n372_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X21 a_2988_n200# a_2932_n244# a_2828_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X22 a_n52_n200# a_n108_n244# a_n212_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X23 a_n852_n200# a_n908_n244# a_n1012_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X24 a_n1012_n200# a_n1068_n244# a_n1172_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X25 a_n2132_n200# a_n2188_n244# a_n2292_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X26 a_n1812_n200# a_n1868_n244# a_n1972_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X27 a_n1972_n200# a_n2028_n244# a_n2132_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X28 a_n1652_n200# a_n1708_n244# a_n1812_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X29 a_908_n200# a_852_n244# a_748_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X30 a_n2932_n200# a_n2988_n244# a_n3092_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X31 a_1708_n200# a_1652_n244# a_1548_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X32 a_n3092_n200# a_n3148_n244# a_n3236_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.28u
X33 a_n2772_n200# a_n2828_n244# a_n2932_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X34 a_2828_n200# a_2772_n244# a_2668_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X35 a_2668_n200# a_2612_n244# a_2508_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X36 a_3148_n200# a_3092_n244# a_2988_n200# VSUBS nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.28u
X37 a_n692_n200# a_n748_n244# a_n852_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X38 a_n1492_n200# a_n1548_n244# a_n1652_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X39 a_748_n200# a_692_n244# a_588_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt pmos_3p3_MLZUAR a_n52_n200# a_n428_n244# a_532_n244# a_588_n200# a_n212_n200#
+ a_n588_n244# a_n676_n200# a_n372_n200# a_108_n200# a_52_n244# a_n532_n200# a_n108_n244#
+ a_212_n244# a_268_n200# a_n268_n244# a_372_n244# w_n762_n330# a_428_n200#
X0 a_588_n200# a_532_n244# a_428_n200# w_n762_n330# pfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_n532_n200# a_n588_n244# a_n676_n200# w_n762_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.28u
X2 a_n372_n200# a_n428_n244# a_n532_n200# w_n762_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X3 a_108_n200# a_52_n244# a_n52_n200# w_n762_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X4 a_428_n200# a_372_n244# a_268_n200# w_n762_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X5 a_268_n200# a_212_n244# a_108_n200# w_n762_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X6 a_n212_n200# a_n268_n244# a_n372_n200# w_n762_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X7 a_n52_n200# a_n108_n244# a_n212_n200# w_n762_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt pmos_3p3_Q3Y3KU a_2988_n200# a_1228_n200# a_n52_n200# a_n852_n200# a_n428_n244#
+ a_n1012_n200# a_532_n244# w_n3322_n330# a_n2772_n200# a_n1388_n244# a_588_n200#
+ a_n1812_n200# a_2292_n244# a_1332_n244# a_n2348_n244# a_2348_n200# a_1388_n200#
+ a_n212_n200# a_n588_n244# a_n1172_n200# a_n3092_n200# a_692_n244# a_n2132_n200#
+ a_n1972_n200# a_n2932_n200# a_1492_n244# a_n1548_n244# a_748_n200# a_2452_n244#
+ a_n2508_n244# a_n372_n200# a_2508_n200# a_1548_n200# a_n748_n244# a_n2292_n200#
+ a_108_n200# a_n1332_n200# a_852_n244# a_52_n244# a_n2668_n244# a_908_n200# a_2612_n244#
+ a_1652_n244# a_n1708_n244# a_2668_n200# a_1708_n200# a_n532_n200# a_n108_n244# a_212_n244#
+ a_268_n200# a_n1492_n200# a_n2452_n200# a_n908_n244# a_n1068_n244# a_n2028_n244#
+ a_1012_n244# a_n1868_n244# a_1068_n200# a_2772_n244# a_n2828_n244# a_2028_n200#
+ a_1812_n244# a_2828_n200# a_1868_n200# a_n692_n200# a_n268_n244# a_372_n244# a_n2188_n244#
+ a_n1652_n200# a_n2612_n200# a_3092_n244# a_1172_n244# a_n1228_n244# a_n3148_n244#
+ a_428_n200# a_2132_n244# a_n2988_n244# a_3148_n200# a_2188_n200# a_n3236_n200# a_2932_n244#
+ a_1972_n244#
X0 a_n1492_n200# a_n1548_n244# a_n1652_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_748_n200# a_692_n244# a_588_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_1548_n200# a_1492_n244# a_1388_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X3 a_n2612_n200# a_n2668_n244# a_n2772_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X4 a_588_n200# a_532_n244# a_428_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X5 a_1388_n200# a_1332_n244# a_1228_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X6 a_n2452_n200# a_n2508_n244# a_n2612_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X7 a_2508_n200# a_2452_n244# a_2348_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X8 a_n532_n200# a_n588_n244# a_n692_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X9 a_n372_n200# a_n428_n244# a_n532_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X10 a_n1332_n200# a_n1388_n244# a_n1492_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X11 a_108_n200# a_52_n244# a_n52_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X12 a_n1172_n200# a_n1228_n244# a_n1332_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X13 a_428_n200# a_372_n244# a_268_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X14 a_268_n200# a_212_n244# a_108_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X15 a_1228_n200# a_1172_n244# a_1068_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X16 a_n2292_n200# a_n2348_n244# a_n2452_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X17 a_1068_n200# a_1012_n244# a_908_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X18 a_2028_n200# a_1972_n244# a_1868_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X19 a_2348_n200# a_2292_n244# a_2188_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X20 a_1868_n200# a_1812_n244# a_1708_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X21 a_2188_n200# a_2132_n244# a_2028_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X22 a_n212_n200# a_n268_n244# a_n372_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X23 a_n52_n200# a_n108_n244# a_n212_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X24 a_2988_n200# a_2932_n244# a_2828_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X25 a_n852_n200# a_n908_n244# a_n1012_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X26 a_n1012_n200# a_n1068_n244# a_n1172_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X27 a_n2132_n200# a_n2188_n244# a_n2292_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X28 a_n1812_n200# a_n1868_n244# a_n1972_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X29 a_n1972_n200# a_n2028_n244# a_n2132_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X30 a_n1652_n200# a_n1708_n244# a_n1812_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X31 a_908_n200# a_852_n244# a_748_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X32 a_n2932_n200# a_n2988_n244# a_n3092_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X33 a_1708_n200# a_1652_n244# a_1548_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X34 a_n3092_n200# a_n3148_n244# a_n3236_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.28u
X35 a_n2772_n200# a_n2828_n244# a_n2932_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X36 a_2828_n200# a_2772_n244# a_2668_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X37 a_3148_n200# a_3092_n244# a_2988_n200# w_n3322_n330# pfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.28u
X38 a_2668_n200# a_2612_n244# a_2508_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X39 a_n692_n200# a_n748_n244# a_n852_n200# w_n3322_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt TG VDD VSS SEL IN OUT
Xnmos_3p3_ECASTA_0 VSS a_n941_n129# a_n941_n129# SEL SEL SEL VSS SEL VSS VSS nmos_3p3_ECASTA
Xnmos_3p3_AEBEG7_0 OUT IN IN OUT SEL IN SEL OUT SEL IN OUT SEL SEL SEL OUT OUT OUT
+ SEL OUT OUT SEL OUT IN IN SEL SEL OUT SEL SEL IN IN IN SEL IN OUT IN SEL SEL SEL
+ IN SEL SEL SEL OUT OUT OUT SEL SEL IN OUT OUT SEL SEL SEL SEL SEL OUT SEL SEL OUT
+ SEL IN IN IN SEL SEL SEL IN IN SEL SEL SEL SEL OUT SEL SEL IN IN IN SEL SEL VSS
+ nmos_3p3_AEBEG7
Xpmos_3p3_MLZUAR_0 VDD SEL SEL VDD a_n941_n129# SEL VDD VDD a_n941_n129# SEL a_n941_n129#
+ SEL SEL VDD SEL SEL VDD a_n941_n129# pmos_3p3_MLZUAR
Xpmos_3p3_Q3Y3KU_0 OUT IN IN OUT a_n941_n129# IN a_n941_n129# VDD OUT a_n941_n129#
+ IN OUT a_n941_n129# a_n941_n129# a_n941_n129# OUT OUT OUT a_n941_n129# OUT OUT a_n941_n129#
+ OUT IN IN a_n941_n129# a_n941_n129# OUT a_n941_n129# a_n941_n129# IN IN IN a_n941_n129#
+ IN OUT IN a_n941_n129# a_n941_n129# a_n941_n129# IN a_n941_n129# a_n941_n129# a_n941_n129#
+ OUT OUT OUT a_n941_n129# a_n941_n129# IN OUT OUT a_n941_n129# a_n941_n129# a_n941_n129#
+ a_n941_n129# a_n941_n129# OUT a_n941_n129# a_n941_n129# OUT a_n941_n129# IN IN IN
+ a_n941_n129# a_n941_n129# a_n941_n129# IN IN a_n941_n129# a_n941_n129# a_n941_n129#
+ a_n941_n129# OUT a_n941_n129# a_n941_n129# IN IN IN a_n941_n129# a_n941_n129# pmos_3p3_Q3Y3KU
.ends

.subckt pmos_3p3_DVJ9E7 a_764_n60# a_n664_n60# a_664_n104# a_560_n60# a_n460_n60#
+ a_n764_n104# a_256_n104# a_n256_n60# a_356_n60# a_n356_n104# a_460_n104# a_n1376_n104#
+ a_1580_n60# a_n1480_n60# a_152_n60# a_n1668_n60# a_1276_n104# a_n560_n104# a_n1580_n104#
+ a_n52_n60# a_1376_n60# a_n1276_n60# a_1480_n104# a_52_n104# a_868_n104# a_n152_n104#
+ a_1172_n60# a_n1072_n60# a_n1172_n104# a_n968_n104# a_1072_n104# a_968_n60# a_n868_n60#
+ w_n1754_n190#
X0 a_n256_n60# a_n356_n104# a_n460_n60# w_n1754_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X1 a_1376_n60# a_1276_n104# a_1172_n60# w_n1754_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X2 a_1580_n60# a_1480_n104# a_1376_n60# w_n1754_n190# pfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X3 a_n460_n60# a_n560_n104# a_n664_n60# w_n1754_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X4 a_n664_n60# a_n764_n104# a_n868_n60# w_n1754_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X5 a_n1072_n60# a_n1172_n104# a_n1276_n60# w_n1754_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X6 a_n868_n60# a_n968_n104# a_n1072_n60# w_n1754_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X7 a_356_n60# a_256_n104# a_152_n60# w_n1754_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X8 a_n1276_n60# a_n1376_n104# a_n1480_n60# w_n1754_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X9 a_560_n60# a_460_n104# a_356_n60# w_n1754_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X10 a_n1480_n60# a_n1580_n104# a_n1668_n60# w_n1754_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X11 a_764_n60# a_664_n104# a_560_n60# w_n1754_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X12 a_152_n60# a_52_n104# a_n52_n60# w_n1754_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X13 a_968_n60# a_868_n104# a_764_n60# w_n1754_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X14 a_n52_n60# a_n152_n104# a_n256_n60# w_n1754_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X15 a_1172_n60# a_1072_n104# a_968_n60# w_n1754_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
.ends

.subckt pmos_3p3_KYXSLM a_764_n60# a_n664_n60# a_n852_n60# a_664_n104# w_n938_n190#
+ a_560_n60# a_n460_n60# a_n764_n104# a_256_n104# a_n256_n60# a_356_n60# a_n356_n104#
+ a_460_n104# a_152_n60# a_n560_n104# a_n52_n60# a_52_n104# a_n152_n104#
X0 a_n256_n60# a_n356_n104# a_n460_n60# w_n938_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X1 a_n460_n60# a_n560_n104# a_n664_n60# w_n938_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X2 a_n664_n60# a_n764_n104# a_n852_n60# w_n938_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X3 a_356_n60# a_256_n104# a_152_n60# w_n938_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X4 a_560_n60# a_460_n104# a_356_n60# w_n938_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X5 a_764_n60# a_664_n104# a_560_n60# w_n938_n190# pfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X6 a_152_n60# a_52_n104# a_n52_n60# w_n938_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X7 a_n52_n60# a_n152_n104# a_n256_n60# w_n938_n190# pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
.ends

.subckt nmos_3p3_AJEA3B a_764_n60# a_n664_n60# a_n852_n60# a_664_n104# a_560_n60#
+ a_n460_n60# a_n764_n104# a_256_n104# a_n256_n60# a_356_n60# a_n356_n104# a_460_n104#
+ a_152_n60# a_n560_n104# a_n52_n60# a_52_n104# a_n152_n104# VSUBS
X0 a_n256_n60# a_n356_n104# a_n460_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X1 a_n460_n60# a_n560_n104# a_n664_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X2 a_n664_n60# a_n764_n104# a_n852_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X3 a_356_n60# a_256_n104# a_152_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X4 a_560_n60# a_460_n104# a_356_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X5 a_764_n60# a_664_n104# a_560_n60# VSUBS nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X6 a_152_n60# a_52_n104# a_n52_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X7 a_n52_n60# a_n152_n104# a_n256_n60# VSUBS nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
.ends

.subckt CM_LSB_mod ITAIL_1 SD0_1 VDD G1_1 G1_2 SD1_1 SD2_1 ITAIL G2_1 OUT_2 OUT_1
+ SD2_3 SD2_4 OUT_3 OUT_4 SD2_5 SD0_2 OUT_5 SD3_1 OUT_6 VSS SD2_2
Xnmos_3p3_MGEA3B_19 OUT_4 SD2_5 ITAIL VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_4 VSS SD2_4 G2_1 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_5 SD2_3 OUT_2 ITAIL VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_6 VSS SD2_3 G2_1 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_7 SD2_3 VSS G2_1 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_8 OUT_2 SD2_3 ITAIL VSS nmos_3p3_MGEA3B
Xpmos_3p3_DVJ9E7_0 VDD G1_1 G1_1 G1_1 G1_2 G1_1 G1_2 G1_1 G1_2 G1_2 G1_2 G1_2 VDD
+ G1_1 G1_1 VDD G1_2 G1_2 G1_1 VDD G1_1 G1_2 G1_1 G1_1 G1_1 G1_1 G1_2 G1_1 G1_2 G1_1
+ G1_2 G1_1 VDD VDD pmos_3p3_DVJ9E7
Xnmos_3p3_MGEA3B_9 VSS SD2_4 G2_1 VSS nmos_3p3_MGEA3B
Xnmos_3p3_9NPLV7_0 SD3_1 OUT_6 SD3_1 SD3_1 VSS ITAIL_1 VSS SD3_1 SD3_1 VSS ITAIL_1
+ SD0_2 VSS SD3_1 ITAIL_1 SD3_1 OUT_6 SD0_2 ITAIL_1 SD0_2 SD3_1 SD3_1 OUT_6 VSS ITAIL_1
+ SD0_2 SD0_2 SD0_2 OUT_6 SD3_1 ITAIL_1 SD3_1 SD0_2 SD0_2 ITAIL_1 ITAIL_1 SD0_2 OUT_6
+ ITAIL_1 SD3_1 VSS ITAIL_1 ITAIL_1 ITAIL_1 SD0_2 ITAIL_1 ITAIL_1 VSS SD3_1 SD0_2
+ ITAIL_1 SD0_2 ITAIL_1 SD0_2 OUT_6 SD3_1 OUT_6 SD0_2 SD3_1 OUT_6 SD0_2 OUT_6 SD3_1
+ SD0_2 VSS VSS nmos_3p3_9NPLV7
Xnmos_3p3_9NPLV7_1 SD3_1 VSS SD3_1 SD3_1 OUT_6 SD0_2 OUT_6 SD3_1 SD3_1 OUT_6 SD0_2
+ ITAIL_1 OUT_6 SD3_1 SD0_2 SD3_1 VSS ITAIL_1 SD0_2 ITAIL_1 SD3_1 SD3_1 VSS OUT_6
+ SD0_2 ITAIL_1 ITAIL_1 ITAIL_1 VSS SD3_1 SD0_2 SD3_1 ITAIL_1 ITAIL_1 SD0_2 SD0_2
+ ITAIL_1 VSS SD0_2 SD3_1 OUT_6 SD0_2 SD0_2 SD0_2 ITAIL_1 SD0_2 SD0_2 OUT_6 SD3_1
+ ITAIL_1 SD0_2 ITAIL_1 SD0_2 ITAIL_1 VSS SD3_1 VSS ITAIL_1 SD3_1 VSS ITAIL_1 VSS
+ SD3_1 ITAIL_1 OUT_6 VSS nmos_3p3_9NPLV7
Xpmos_3p3_KYXSLM_0 VDD SD1_1 VDD G1_1 VDD SD1_1 ITAIL_1 G1_1 G1_2 SD1_1 ITAIL_1 G1_2
+ G1_2 SD1_1 G1_2 VDD G1_1 G1_1 pmos_3p3_KYXSLM
Xpmos_3p3_KYXSLM_1 VDD SD1_1 VDD G1_1 VDD SD1_1 ITAIL_1 G1_1 G1_2 SD1_1 ITAIL_1 G1_2
+ G1_2 SD1_1 G1_2 VDD G1_1 G1_1 pmos_3p3_KYXSLM
Xnmos_3p3_AJEA3B_0 OUT_5 SD0_1 OUT_5 ITAIL_1 SD0_1 VSS ITAIL_1 SD0_2 SD0_1 VSS SD0_2
+ SD0_2 SD0_1 SD0_2 OUT_5 ITAIL_1 ITAIL_1 VSS nmos_3p3_AJEA3B
Xnmos_3p3_MGEA3B_40 VSS SD2_1 G2_1 VSS nmos_3p3_MGEA3B
Xnmos_3p3_AJEA3B_1 VSS SD0_1 VSS SD0_2 SD0_1 OUT_5 SD0_2 ITAIL_1 SD0_1 OUT_5 ITAIL_1
+ ITAIL_1 SD0_1 ITAIL_1 VSS SD0_2 SD0_2 VSS nmos_3p3_AJEA3B
Xnmos_3p3_MGEA3B_30 SD2_5 OUT_4 ITAIL VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_41 SD2_1 VSS G2_1 VSS nmos_3p3_MGEA3B
Xnmos_3p3_AJEA3B_2 OUT_5 SD0_1 OUT_5 ITAIL_1 SD0_1 VSS ITAIL_1 SD0_2 SD0_1 VSS SD0_2
+ SD0_2 SD0_1 SD0_2 OUT_5 ITAIL_1 ITAIL_1 VSS nmos_3p3_AJEA3B
Xnmos_3p3_MGEA3B_31 OUT_4 SD2_5 ITAIL VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_20 SD2_5 OUT_4 ITAIL VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_42 VSS SD2_1 G2_1 VSS nmos_3p3_MGEA3B
Xnmos_3p3_AJEA3B_4 ITAIL_1 SD0_2 ITAIL_1 ITAIL_1 SD0_2 VSS ITAIL_1 SD0_2 SD0_2 VSS
+ SD0_2 SD0_2 SD0_2 SD0_2 ITAIL_1 ITAIL_1 ITAIL_1 VSS nmos_3p3_AJEA3B
Xnmos_3p3_AJEA3B_3 VSS SD0_1 VSS SD0_2 SD0_1 OUT_5 SD0_2 ITAIL_1 SD0_1 OUT_5 ITAIL_1
+ ITAIL_1 SD0_1 ITAIL_1 VSS SD0_2 SD0_2 VSS nmos_3p3_AJEA3B
Xnmos_3p3_MGEA3B_32 SD2_5 VSS G2_1 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_10 SD2_4 OUT_3 ITAIL VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_21 VSS SD2_5 G2_1 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_43 SD2_1 VSS G2_1 VSS nmos_3p3_MGEA3B
Xnmos_3p3_AJEA3B_5 VSS SD0_2 VSS SD0_2 SD0_2 ITAIL_1 SD0_2 ITAIL_1 SD0_2 ITAIL_1 ITAIL_1
+ ITAIL_1 SD0_2 ITAIL_1 VSS SD0_2 SD0_2 VSS nmos_3p3_AJEA3B
Xnmos_3p3_MGEA3B_44 SD2_1 G1_2 ITAIL VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_33 VSS SD2_5 G2_1 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_11 SD2_4 OUT_3 ITAIL VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_22 SD2_5 VSS G2_1 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_46 SD2_1 G1_2 ITAIL VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_45 VSS SD2_1 G2_1 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_23 G1_2 SD2_1 ITAIL VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_12 SD2_5 OUT_4 ITAIL VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_34 SD2_5 OUT_4 ITAIL VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_13 SD2_4 VSS G2_1 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_24 OUT_4 SD2_5 ITAIL VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_35 SD2_1 G1_2 ITAIL VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_47 VSS SD2_1 G2_1 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_36 SD2_1 VSS G2_1 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_14 SD2_4 VSS G2_1 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_25 SD2_1 G1_2 ITAIL VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_26 G1_2 SD2_1 ITAIL VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_37 SD2_1 VSS G2_1 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_15 OUT_3 SD2_4 ITAIL VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_0 G2_1 VSS G2_1 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_16 OUT_3 SD2_4 ITAIL VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_27 OUT_4 SD2_5 ITAIL VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_38 G1_2 SD2_1 ITAIL VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_17 VSS SD2_5 G2_1 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_1 OUT_1 SD2_2 ITAIL VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_28 SD2_5 VSS G2_1 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_39 G1_2 SD2_1 ITAIL VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_18 SD2_5 VSS G2_1 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_2 SD2_2 VSS G2_1 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_3 ITAIL G2_1 ITAIL VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_29 VSS SD2_5 G2_1 VSS nmos_3p3_MGEA3B
.ends

.subckt LSBs_magic_TG B2 b1 b1b b2 b2b b3 b3b b4 b4b b5 b5b b6 b6b OUT1 OUT2 OUT3
+ OUT4 OUT5 OUT6 G2 SD2_2 SD2_3 SD2_5 SD2_1 SD2_4 G1_2 SD1_1 G1_1 SD3_1 SDn_1 SDn_2
+ IT B1 B3 B4 B5 B6 OUT- OUT+ VSS VDD ITAIL C32_D SEL_L SDc_1 Gc_1 Gc_2 SDc_2 C32_U
Xnmos_3p3_MGEA3B_169 OUT4 TG_0/IN b4 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_158 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_147 OUT2 TG_1/IN b2b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEAJ7_12 TG_0/IN b3b TG_0/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEAJ7_23 TG_0/IN b4b TG_0/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEAJ7_34 TG_0/IN b4b TG_0/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEA3B_159 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_148 TG_1/IN OUT2 b2b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_307 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_318 OUT5 TG_1/IN b5b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_329 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEAJ7_13 TG_1/IN b3 TG_1/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEAJ7_35 TG_1/IN b4 TG_1/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEAJ7_24 TG_0/IN b4b TG_0/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEA3B_308 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_319 TG_1/IN OUT5 b5b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_149 OUT2 TG_0/IN b2 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEAJ7_14 TG_1/IN b1 TG_1/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEAJ7_36 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEAJ7_25 TG_1/IN b4 TG_1/IN VSS nmos_3p3_MGEAJ7
XBalance_Inverter_0 VDD VSS b4 b4b B4 Balance_Inverter
Xnmos_3p3_MGEA3B_309 OUT5 TG_1/IN b5b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEAJ7_15 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEAJ7_37 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEAJ7_26 TG_1/IN b4 TG_1/IN VSS nmos_3p3_MGEAJ7
XBalance_Inverter_1 VDD VSS b3 b3b B3 Balance_Inverter
Xnmos_3p3_MGEA3B_290 TG_1/IN TG_1/IN b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEAJ7_16 TG_1/IN b3 TG_1/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEAJ7_38 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEAJ7_27 TG_0/IN b4b TG_0/IN VSS nmos_3p3_MGEAJ7
XBalance_Inverter_2 VDD VSS b2 b2b B2 Balance_Inverter
Xnmos_3p3_MGEA3B_291 TG_1/IN TG_1/IN b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_280 TG_1/IN TG_1/IN b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEAJ7_17 TG_1/IN b3 TG_1/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEAJ7_39 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEAJ7_28 TG_1/IN b4 TG_1/IN VSS nmos_3p3_MGEAJ7
XBalance_Inverter_3 VDD VSS b1 b1b B1 Balance_Inverter
Xnmos_3p3_MGEA3B_292 TG_0/IN TG_0/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_281 TG_1/IN TG_1/IN b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_270 TG_0/IN TG_0/IN b5b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEAJ7_18 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEAJ7_29 TG_0/IN b4b TG_0/IN VSS nmos_3p3_MGEAJ7
XBalance_Inverter_4 VDD VSS b5 b5b B5 Balance_Inverter
Xnmos_3p3_MGEA3B_293 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_282 TG_1/IN TG_1/IN b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_271 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_260 TG_0/IN TG_0/IN b5b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEAJ7_19 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEAJ7
XBalance_Inverter_5 VDD VSS b6 b6b B6 Balance_Inverter
Xnmos_3p3_MGEA3B_294 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_283 TG_0/IN TG_0/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_261 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_272 TG_1/IN TG_1/IN b5 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_250 TG_0/IN OUT6 b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_284 TG_0/IN TG_0/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_273 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_262 TG_0/IN TG_0/IN b5b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_295 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_251 OUT6 TG_1/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_240 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_285 TG_0/IN TG_0/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_274 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_263 TG_1/IN TG_1/IN b5 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_296 TG_1/IN OUT6 b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_241 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_252 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_230 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_286 TG_1/IN TG_1/IN b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_275 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_264 TG_1/IN TG_1/IN b5 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_297 OUT6 TG_0/IN b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_242 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_253 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_220 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_287 TG_1/IN TG_1/IN b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_276 TG_0/IN TG_0/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_265 TG_1/IN TG_1/IN b5 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_298 OUT6 TG_1/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_243 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_232 TG_0/IN OUT6 b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_254 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_210 TG_1/IN OUT5 b5b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_221 OUT6 TG_0/IN b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_288 TG_0/IN TG_0/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_200 TG_1/IN TG_1/IN b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_277 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_266 TG_0/IN TG_0/IN b5b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_255 TG_1/IN TG_1/IN b5 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_299 TG_1/IN OUT6 b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_244 TG_1/IN OUT6 b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_233 OUT6 TG_1/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_211 OUT5 TG_1/IN b5b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_222 TG_0/IN OUT6 b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_201 TG_0/IN TG_0/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_289 TG_0/IN TG_0/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_278 TG_1/IN TG_1/IN b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_267 TG_1/IN TG_1/IN b5 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_256 TG_1/IN TG_1/IN b5 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_245 OUT6 TG_0/IN b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_234 TG_1/IN OUT6 b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_212 TG_1/IN OUT5 b5b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_223 TG_1/IN OUT6 b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_279 TG_0/IN TG_0/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_202 TG_1/IN TG_1/IN b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_268 TG_0/IN TG_0/IN b5b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_257 TG_0/IN TG_0/IN b5b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_246 TG_0/IN OUT6 b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_235 OUT6 TG_0/IN b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_213 OUT5 TG_0/IN b5 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_224 OUT6 TG_1/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_203 TG_1/IN TG_1/IN b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_269 TG_0/IN TG_0/IN b5b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_258 TG_1/IN TG_1/IN b5 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_247 OUT6 TG_1/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_236 TG_0/IN OUT6 b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_214 TG_0/IN OUT5 b5 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_225 TG_1/IN OUT6 b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_204 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_259 TG_0/IN TG_0/IN b5b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_248 TG_1/IN OUT6 b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_237 OUT6 TG_1/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_215 OUT5 TG_1/IN b5b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_226 OUT6 TG_0/IN b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_205 TG_1/IN TG_1/IN b6 VSS nmos_3p3_MGEA3B
XCM_32_0 VSS IT SDn_2 VDD Gc_2 Gc_1 SDc_2 C32_U C32_D SDc_1 CM_32
Xnmos_3p3_MGEA3B_238 TG_1/IN OUT6 b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_249 OUT6 TG_0/IN b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_216 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_227 TG_0/IN OUT6 b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_206 TG_0/IN TG_0/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_239 OUT6 TG_0/IN b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_217 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_228 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_207 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_218 OUT6 TG_1/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_229 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
XTG_0 VDD VSS SEL_L TG_0/IN OUT+ TG
Xnmos_3p3_MGEA3B_390 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_208 TG_0/IN TG_0/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_219 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_380 OUT6 TG_1/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_391 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
XTG_1 VDD VSS SEL_L TG_1/IN OUT- TG
Xnmos_3p3_MGEA3B_209 OUT5 TG_0/IN b5 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_381 OUT6 TG_0/IN b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_370 TG_1/IN OUT6 b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_382 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_371 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_360 TG_0/IN OUT6 b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_190 TG_1/IN TG_1/IN b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_383 TG_0/IN OUT6 b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_372 OUT6 TG_0/IN b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_361 OUT6 TG_1/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_350 TG_0/IN OUT6 b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_180 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_191 TG_1/IN TG_1/IN b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEAJ7_0 TG_1/IN b2 TG_1/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEA3B_170 OUT4 TG_1/IN b4b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_181 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_192 TG_0/IN TG_0/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_384 OUT6 TG_0/IN b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_373 OUT6 TG_0/IN b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_340 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_362 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_351 TG_1/IN OUT6 b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEAJ7_1 TG_0/IN b1b TG_0/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEA3B_385 OUT6 TG_1/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_374 TG_0/IN OUT6 b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_341 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_330 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_363 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_352 OUT6 TG_1/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_160 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_182 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_171 TG_0/IN OUT4 b4 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_193 TG_0/IN TG_0/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEAJ7_2 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEA3B_161 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_150 TG_0/IN OUT3 b3 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_183 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_172 OUT4 TG_1/IN b4b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_194 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_386 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_375 OUT6 TG_1/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_342 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_331 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_364 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_320 OUT5 TG_0/IN b5 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_353 TG_0/IN OUT6 b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEAJ7_3 TG_0/IN b4b TG_0/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEA3B_387 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_376 TG_1/IN OUT6 b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_321 TG_0/IN OUT5 b5 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_332 OUT5 TG_0/IN b5 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_310 TG_0/IN OUT5 b5 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_354 TG_1/IN OUT6 b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_365 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_343 TG_0/IN OUT6 b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_162 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_151 OUT3 TG_1/IN b3b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_140 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_173 TG_1/IN OUT4 b4b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_184 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_195 TG_1/IN TG_1/IN b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEAJ7_4 TG_0/IN b3b TG_0/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEA3B_141 OUT3 TG_1/IN b3b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_152 TG_1/IN OUT3 b3b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_163 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_185 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_174 OUT4 TG_0/IN b4 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_196 TG_0/IN TG_0/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_388 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_377 TG_1/IN OUT6 b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_333 TG_0/IN OUT5 b5 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_322 OUT5 TG_1/IN b5b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_355 TG_1/IN OUT6 b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_300 TG_0/IN OUT6 b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_311 TG_1/IN OUT5 b5b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_366 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_344 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEAJ7_5 TG_0/IN b3b TG_0/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEA3B_389 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_378 TG_0/IN OUT6 b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_367 TG_0/IN OUT6 b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_334 OUT5 TG_1/IN b5b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_323 TG_1/IN OUT5 b5b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_356 OUT6 TG_0/IN b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_301 TG_0/IN OUT6 b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_312 OUT5 TG_0/IN b5 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_345 OUT6 TG_1/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_142 OUT1 TG_1/IN b1b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_153 OUT3 TG_0/IN b3 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_186 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_175 TG_0/IN OUT4 b4 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_164 OUT4 TG_1/IN b4b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_197 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEAJ7_6 TG_1/IN b2 TG_1/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEA3B_154 TG_0/IN OUT1 b1 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_143 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_176 OUT4 TG_1/IN b4b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_165 TG_1/IN OUT4 b4b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_379 TG_1/IN OUT6 b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_368 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_324 OUT5 TG_0/IN b5 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_335 TG_1/IN OUT5 b5b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_313 OUT5 TG_1/IN b5b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_357 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_302 OUT6 TG_1/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_187 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_346 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_198 TG_0/IN TG_0/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEAJ7_7 TG_0/IN b2b TG_0/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEAJ7_30 TG_0/IN b4b TG_0/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEA3B_369 OUT6 TG_1/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_336 OUT5 TG_1/IN b5b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_314 TG_0/IN OUT5 b5 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_358 OUT6 TG_1/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_303 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_325 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_347 TG_1/IN OUT6 b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_144 TG_1/IN OUT3 b3b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_155 TG_0/IN OUT2 b2 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_177 TG_1/IN OUT4 b4b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_166 OUT4 TG_0/IN b4 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_199 TG_0/IN TG_0/IN b6b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_188 TG_1/IN TG_1/IN b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEAJ7_8 TG_0/IN b2b TG_0/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEAJ7_20 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEAJ7_31 TG_1/IN b4 TG_1/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEA3B_337 TG_1/IN OUT5 b5b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_315 TG_1/IN OUT5 b5b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_304 OUT6 TG_0/IN b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_326 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_348 OUT6 TG_0/IN b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_359 OUT6 TG_0/IN b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_145 OUT3 TG_0/IN b3 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_156 TG_0/IN OUT3 b3 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_167 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_178 OUT4 TG_0/IN b4 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_189 TG_0/IN OUT5 b5 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEAJ7_9 TG_1/IN b3 TG_1/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEAJ7_10 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEAJ7_21 TG_1/IN b4 TG_1/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEAJ7_32 TG_1/IN b4 TG_1/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEA3B_327 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_338 OUT5 TG_0/IN b5 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_316 OUT5 TG_0/IN b5 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_305 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_349 OUT6 TG_0/IN b6 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_157 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_179 TG_1/IN OUT4 b4b VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_168 TG_0/IN OUT4 b4 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_146 TG_0/IN OUT4 b4 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEAJ7_11 TG_0/IN b3b TG_0/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEAJ7_22 TG_1/IN b4 TG_1/IN VSS nmos_3p3_MGEAJ7
Xnmos_3p3_MGEAJ7_33 TG_0/IN b4b TG_0/IN VSS nmos_3p3_MGEAJ7
XCM_LSB_mod_0 IT SDn_1 VDD G1_1 G1_2 SD1_1 SD2_1 ITAIL G2 OUT2 OUT1 SD2_3 SD2_4 OUT3
+ OUT4 SD2_5 SDn_2 OUT5 SD3_1 OUT6 VSS SD2_2 CM_LSB_mod
Xnmos_3p3_MGEA3B_328 TG_0/IN TG_0/IN TG_0/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_339 TG_0/IN OUT5 b5 VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_306 TG_1/IN TG_1/IN TG_1/IN VSS nmos_3p3_MGEA3B
Xnmos_3p3_MGEA3B_317 TG_0/IN OUT5 b5 VSS nmos_3p3_MGEA3B
.ends

.subckt DAC_12_Bit R6 R5 R3 R4 R2 R1 R0 C6 C5 C3 C4 C2 C1 C0 VDD VSS OUT+ OUT- B12
+ B11 B10 B12D B11D B10D B9 B8 B7 B9D B8D B7D SEL_L SEL B1 B2 B3 B4 B5 B6 B1D B2D
+ B3D B4D B5D B6D ITAIL B10M B11M B12M B1M B2M B3M B5M B6M B9M B8M B7M cur_1_d cur_1_u
+ cur_2_u cur_2_d cur_3_u cur_3_d cur_6_u cur_6_d cur_7_d cur_7_u cur_8_d cur_8_u
+ cur_9_u cur_9_d cur_10_d cur_10_u cur_11_u cur_11_d cur_12_d cur_12_u cur_13_u cur_13_d
+ cur_14_u cur_14_d cur_15_d cur_15_u cur_16_d cur_16_u cur_17_d cur_17_u cur_18_d
+ cur_18_u cur_19_u cur_19_d cur_20_u cur_20_d cur_21_d cur_21_u SEL_M cur_4_d cur_4_u
+ cur_5_u cur_5_d B4M
XMSB_Unit_Cell_49 cur_7_d R3 VSS VDD MSB_Unit_Cell_49/QB MSB_Unit_Cell_49/Q MSB_Unit_Cell_49/OUT
+ OUT+ OUT- MSB_Unit_Cell_49/SD R2 cur_7_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_38 cur_21_d R4 C6 VDD MSB_Unit_Cell_38/QB MSB_Unit_Cell_38/Q MSB_Unit_Cell_38/OUT
+ OUT+ OUT- MSB_Unit_Cell_38/SD R3 cur_21_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_27 cur_14_d R6 C1 VDD MSB_Unit_Cell_27/QB MSB_Unit_Cell_27/Q MSB_Unit_Cell_27/OUT
+ OUT+ OUT- MSB_Unit_Cell_27/SD R5 cur_14_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_16 cur_16_d R6 C3 VDD MSB_Unit_Cell_16/QB MSB_Unit_Cell_16/Q MSB_Unit_Cell_16/OUT
+ OUT+ OUT- MSB_Unit_Cell_16/SD R5 cur_16_u VSS MSB_Unit_Cell
XINV_BUFF_16 B11M INV_BUFF_16/SD1 B11D VDD VSS INV_BUFF
XCM_32_C_17 CM_32_C_17/SD0_1 CM_32_C_17/G1_2 CM_32_C_17/G1_1 CM_32_C_17/SD2_0 cur_6_d
+ cur_6_u VSS VDD cur_7_d cur_7_u CM_32_C
XMSB_Unit_Cell_39 cur_7_d R0 VSS VDD MSB_Unit_Cell_39/QB MSB_Unit_Cell_39/Q MSB_Unit_Cell_39/OUT
+ OUT+ OUT- MSB_Unit_Cell_39/SD VDD cur_7_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_28 cur_4_d R4 C3 VDD MSB_Unit_Cell_28/QB MSB_Unit_Cell_28/Q MSB_Unit_Cell_28/OUT
+ OUT+ OUT- MSB_Unit_Cell_28/SD R3 cur_4_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_17 cur_16_d R6 C2 VDD MSB_Unit_Cell_17/QB MSB_Unit_Cell_17/Q MSB_Unit_Cell_17/OUT
+ OUT+ OUT- MSB_Unit_Cell_17/SD R5 cur_16_u VSS MSB_Unit_Cell
XINV_BUFF_17 B8M INV_BUFF_17/SD1 B8D VDD VSS INV_BUFF
XCM_32_C_18 CM_32_C_18/SD0_1 CM_32_C_18/G1_2 CM_32_C_18/G1_1 CM_32_C_18/SD2_0 cur_9_d
+ cur_9_u VSS VDD cur_8_d cur_8_u CM_32_C
XMSB_Unit_Cell_29 cur_14_d R4 C1 VDD MSB_Unit_Cell_29/QB MSB_Unit_Cell_29/Q MSB_Unit_Cell_29/OUT
+ OUT+ OUT- MSB_Unit_Cell_29/SD R3 cur_14_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_18 cur_4_d R5 C0 VDD MSB_Unit_Cell_18/QB MSB_Unit_Cell_18/Q MSB_Unit_Cell_18/OUT
+ OUT+ OUT- MSB_Unit_Cell_18/SD R4 cur_4_u VSS MSB_Unit_Cell
XINV_BUFF_18 B12 INV_BUFF_18/SD1 B12M VDD VSS INV_BUFF
XCM_32_C_19 CM_32_C_19/SD0_1 CM_32_C_19/G1_2 CM_32_C_19/G1_1 CM_32_C_19/SD2_0 cur_14_d
+ cur_14_u VSS VDD cur_15_d cur_15_u CM_32_C
XINV_BUFF_0 B6M INV_BUFF_0/SD1 B6D VDD VSS INV_BUFF
XMSB_Unit_Cell_19 cur_14_d R4 C2 VDD MSB_Unit_Cell_19/QB MSB_Unit_Cell_19/Q MSB_Unit_Cell_19/OUT
+ OUT+ OUT- MSB_Unit_Cell_19/SD R3 cur_14_u VSS MSB_Unit_Cell
XINV_BUFF_19 B11 INV_BUFF_19/SD1 B11M VDD VSS INV_BUFF
XINV_BUFF_1 B6 INV_BUFF_1/SD1 B6M VDD VSS INV_BUFF
XMSB_Unit_Cell_0 cur_3_d R3 C3 VDD MSB_Unit_Cell_0/QB MSB_Unit_Cell_0/Q MSB_Unit_Cell_0/OUT
+ OUT+ OUT- MSB_Unit_Cell_0/SD R2 cur_3_u VSS MSB_Unit_Cell
XINV_BUFF_2 B1M INV_BUFF_2/SD1 B1D VDD VSS INV_BUFF
XMSB_Unit_Cell_1 cur_10_d R2 C2 VDD MSB_Unit_Cell_1/QB MSB_Unit_Cell_1/Q MSB_Unit_Cell_1/OUT
+ OUT+ OUT- MSB_Unit_Cell_1/SD R1 cur_10_u VSS MSB_Unit_Cell
XINV_BUFF_3 B5 INV_BUFF_3/SD1 B5M VDD VSS INV_BUFF
XMSB_Unit_Cell_2 cur_2_d R3 C4 VDD MSB_Unit_Cell_2/QB MSB_Unit_Cell_2/Q MSB_Unit_Cell_2/OUT
+ OUT+ OUT- MSB_Unit_Cell_2/SD R2 cur_2_u VSS MSB_Unit_Cell
XINV_BUFF_4 B4 INV_BUFF_4/SD1 B4M VDD VSS INV_BUFF
XMSB_Unit_Cell_3 cur_13_d R2 C3 VDD MSB_Unit_Cell_3/QB MSB_Unit_Cell_3/Q MSB_Unit_Cell_3/OUT
+ OUT+ OUT- MSB_Unit_Cell_3/SD R1 cur_13_u VSS MSB_Unit_Cell
XINV_BUFF_5 B3 INV_BUFF_5/SD1 B3M VDD VSS INV_BUFF
XMSB_Unit_Cell_4 cur_5_d R4 C4 VDD MSB_Unit_Cell_4/QB MSB_Unit_Cell_4/Q MSB_Unit_Cell_4/OUT
+ OUT+ OUT- MSB_Unit_Cell_4/SD R3 cur_5_u VSS MSB_Unit_Cell
Xtherm_Dec_0 B12D VDD R6 R5 R3 R4 R2 R1 R0 B10D B11D VSS therm_Dec
XINV_BUFF_6 B2 INV_BUFF_6/SD1 B2M VDD VSS INV_BUFF
XMSB_Unit_Cell_5 cur_18_d R6 C4 VDD MSB_Unit_Cell_5/QB MSB_Unit_Cell_5/Q MSB_Unit_Cell_5/OUT
+ OUT+ OUT- MSB_Unit_Cell_5/SD R5 cur_18_u VSS MSB_Unit_Cell
XINV_BUFF_7 SEL_L INV_BUFF_7/SD1 SEL_M VDD VSS INV_BUFF
Xtherm_Dec_1 B9D VDD C6 C5 C3 C4 C2 C1 C0 B7D B8D VSS therm_Dec
XMSB_Unit_Cell_6 cur_18_d R6 C5 VDD MSB_Unit_Cell_6/QB MSB_Unit_Cell_6/Q MSB_Unit_Cell_6/OUT
+ OUT+ OUT- MSB_Unit_Cell_6/SD R5 cur_18_u VSS MSB_Unit_Cell
XINV_BUFF_8 B1 INV_BUFF_8/SD1 B1M VDD VSS INV_BUFF
XMSB_Unit_Cell_7 cur_20_d R6 C6 VDD MSB_Unit_Cell_7/QB MSB_Unit_Cell_7/Q MSB_Unit_Cell_7/OUT
+ OUT+ OUT- MSB_Unit_Cell_7/SD R5 cur_20_u VSS MSB_Unit_Cell
XINV_BUFF_9 B5M INV_BUFF_9/SD1 B5D VDD VSS INV_BUFF
XMSB_Unit_Cell_8 cur_20_d R5 C2 VDD MSB_Unit_Cell_8/QB MSB_Unit_Cell_8/Q MSB_Unit_Cell_8/OUT
+ OUT+ OUT- MSB_Unit_Cell_8/SD R4 cur_20_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_9 cur_20_d R4 C5 VDD MSB_Unit_Cell_9/QB MSB_Unit_Cell_9/Q MSB_Unit_Cell_9/OUT
+ OUT+ OUT- MSB_Unit_Cell_9/SD R3 cur_20_u VSS MSB_Unit_Cell
XCM_32_C_0 CM_32_C_0/SD0_1 CM_32_C_0/G1_2 CM_32_C_0/G1_1 CM_32_C_0/SD2_0 cur_1_d cur_1_u
+ VSS VDD cur_3_d cur_3_u CM_32_C
XCM_32_C_1 CM_32_C_1/SD0_1 CM_32_C_1/G1_2 CM_32_C_1/G1_1 CM_32_C_1/SD2_0 cur_1_d cur_1_u
+ VSS VDD cur_4_d cur_4_u CM_32_C
XCM_32_C_2 CM_32_C_2/SD0_1 CM_32_C_2/G1_2 CM_32_C_2/G1_1 CM_32_C_2/SD2_0 cur_1_d cur_1_u
+ VSS VDD cur_5_d cur_5_u CM_32_C
XMSB_Unit_Cell_60 cur_11_d R0 C2 VDD MSB_Unit_Cell_60/QB MSB_Unit_Cell_60/Q MSB_Unit_Cell_60/OUT
+ OUT+ OUT- MSB_Unit_Cell_60/SD VDD cur_11_u VSS MSB_Unit_Cell
XCM_32_C_3 CM_32_C_3/SD0_1 CM_32_C_3/G1_2 CM_32_C_3/G1_1 CM_32_C_3/SD2_0 cur_1_d cur_1_u
+ VSS VDD cur_2_d cur_2_u CM_32_C
XMSB_Unit_Cell_61 cur_8_d R0 C3 VDD MSB_Unit_Cell_61/QB MSB_Unit_Cell_61/Q MSB_Unit_Cell_61/OUT
+ OUT+ OUT- MSB_Unit_Cell_61/SD VDD cur_8_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_50 cur_7_d R1 VSS VDD MSB_Unit_Cell_50/QB MSB_Unit_Cell_50/Q MSB_Unit_Cell_50/OUT
+ OUT+ OUT- MSB_Unit_Cell_50/SD R0 cur_7_u VSS MSB_Unit_Cell
XCM_32_C_4 CM_32_C_4/SD0_1 CM_32_C_4/G1_2 CM_32_C_4/G1_1 CM_32_C_4/SD2_0 cur_4_d cur_4_u
+ VSS VDD cur_16_d cur_16_u CM_32_C
XMSB_Unit_Cell_40 cur_17_d VSS C0 VDD MSB_Unit_Cell_40/QB MSB_Unit_Cell_40/Q MSB_Unit_Cell_40/OUT
+ OUT+ OUT- MSB_Unit_Cell_40/SD R6 cur_17_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_51 cur_12_d R1 C0 VDD MSB_Unit_Cell_51/QB MSB_Unit_Cell_51/Q MSB_Unit_Cell_51/OUT
+ OUT+ OUT- MSB_Unit_Cell_51/SD R0 cur_12_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_62 cur_8_d R0 C6 VDD MSB_Unit_Cell_62/QB MSB_Unit_Cell_62/Q MSB_Unit_Cell_62/OUT
+ OUT+ OUT- MSB_Unit_Cell_62/SD VDD cur_8_u VSS MSB_Unit_Cell
XCM_32_C_5 CM_32_C_5/SD0_1 CM_32_C_5/G1_2 CM_32_C_5/G1_1 CM_32_C_5/SD2_0 cur_13_d
+ cur_13_u VSS VDD cur_12_d cur_12_u CM_32_C
XMSB_Unit_Cell_41 cur_17_d VSS C3 VDD MSB_Unit_Cell_41/QB MSB_Unit_Cell_41/Q MSB_Unit_Cell_41/OUT
+ OUT+ OUT- MSB_Unit_Cell_41/SD R6 cur_17_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_30 cur_13_d R3 C1 VDD MSB_Unit_Cell_30/QB MSB_Unit_Cell_30/Q MSB_Unit_Cell_30/OUT
+ OUT+ OUT- MSB_Unit_Cell_30/SD R2 cur_13_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_52 cur_15_d R6 C0 VDD MSB_Unit_Cell_52/QB MSB_Unit_Cell_52/Q MSB_Unit_Cell_52/OUT
+ OUT+ OUT- MSB_Unit_Cell_52/SD R5 cur_15_u VSS MSB_Unit_Cell
XCM_32_C_6 CM_32_C_6/SD0_1 CM_32_C_6/G1_2 CM_32_C_6/G1_1 CM_32_C_6/SD2_0 cur_5_d cur_5_u
+ VSS VDD cur_18_d cur_18_u CM_32_C
XMSB_Unit_Cell_31 cur_12_d R1 C1 VDD MSB_Unit_Cell_31/QB MSB_Unit_Cell_31/Q MSB_Unit_Cell_31/OUT
+ OUT+ OUT- MSB_Unit_Cell_31/SD R0 cur_12_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_20 cur_13_d R3 C2 VDD MSB_Unit_Cell_20/QB MSB_Unit_Cell_20/Q MSB_Unit_Cell_20/OUT
+ OUT+ OUT- MSB_Unit_Cell_20/SD R2 cur_13_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_42 cur_3_d R2 C6 VDD MSB_Unit_Cell_42/QB MSB_Unit_Cell_42/Q MSB_Unit_Cell_42/OUT
+ OUT+ OUT- MSB_Unit_Cell_42/SD R1 cur_3_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_53 cur_15_d R4 C0 VDD MSB_Unit_Cell_53/QB MSB_Unit_Cell_53/Q MSB_Unit_Cell_53/OUT
+ OUT+ OUT- MSB_Unit_Cell_53/SD R3 cur_15_u VSS MSB_Unit_Cell
XCM_32_C_7 CM_32_C_7/SD0_1 CM_32_C_7/G1_2 CM_32_C_7/G1_1 CM_32_C_7/SD2_0 cur_5_d cur_5_u
+ VSS VDD cur_20_d cur_20_u CM_32_C
XINV_BUFF_20 B10 INV_BUFF_20/SD1 B10M VDD VSS INV_BUFF
XCM_32_C_10 CM_32_C_10/SD0_1 CM_32_C_10/G1_2 CM_32_C_10/G1_1 CM_32_C_10/SD2_0 cur_3_d
+ cur_3_u VSS VDD cur_10_d cur_10_u CM_32_C
XMSB_Unit_Cell_43 cur_17_d VSS C5 VDD MSB_Unit_Cell_43/QB MSB_Unit_Cell_43/Q MSB_Unit_Cell_43/OUT
+ OUT+ OUT- MSB_Unit_Cell_43/SD R6 cur_17_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_21 cur_9_d R1 C3 VDD MSB_Unit_Cell_21/QB MSB_Unit_Cell_21/Q MSB_Unit_Cell_21/OUT
+ OUT+ OUT- MSB_Unit_Cell_21/SD R0 cur_9_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_54 cur_15_d R3 C0 VDD MSB_Unit_Cell_54/QB MSB_Unit_Cell_54/Q MSB_Unit_Cell_54/OUT
+ OUT+ OUT- MSB_Unit_Cell_54/SD R2 cur_15_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_10 cur_6_d R3 C5 VDD MSB_Unit_Cell_10/QB MSB_Unit_Cell_10/Q MSB_Unit_Cell_10/OUT
+ OUT+ OUT- MSB_Unit_Cell_10/SD R2 cur_6_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_32 cur_19_d R5 C6 VDD MSB_Unit_Cell_32/QB MSB_Unit_Cell_32/Q MSB_Unit_Cell_32/OUT
+ OUT+ OUT- MSB_Unit_Cell_32/SD R4 cur_19_u VSS MSB_Unit_Cell
XINV_BUFF_21 B9M INV_BUFF_21/SD1 B9D VDD VSS INV_BUFF
XCM_32_C_8 CM_32_C_8/SD0_1 CM_32_C_8/G1_2 CM_32_C_8/G1_1 CM_32_C_8/SD2_0 cur_2_d cur_2_u
+ VSS VDD cur_6_d cur_6_u CM_32_C
XINV_BUFF_10 B4M INV_BUFF_10/SD1 B4D VDD VSS INV_BUFF
XCM_32_C_11 CM_32_C_11/SD0_1 CM_32_C_11/G1_2 CM_32_C_11/G1_1 CM_32_C_11/SD2_0 cur_3_d
+ cur_3_u VSS VDD cur_13_d cur_13_u CM_32_C
XMSB_Unit_Cell_44 cur_19_d VSS C6 VDD MSB_Unit_Cell_44/QB MSB_Unit_Cell_44/Q MSB_Unit_Cell_44/OUT
+ OUT+ OUT- MSB_Unit_Cell_44/SD R6 cur_19_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_22 cur_11_d R1 C2 VDD MSB_Unit_Cell_22/QB MSB_Unit_Cell_22/Q MSB_Unit_Cell_22/OUT
+ OUT+ OUT- MSB_Unit_Cell_22/SD R0 cur_11_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_33 cur_6_d R1 C6 VDD MSB_Unit_Cell_33/QB MSB_Unit_Cell_33/Q MSB_Unit_Cell_33/OUT
+ OUT+ OUT- MSB_Unit_Cell_33/SD R0 cur_6_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_55 cur_12_d R2 C1 VDD MSB_Unit_Cell_55/QB MSB_Unit_Cell_55/Q MSB_Unit_Cell_55/OUT
+ OUT+ OUT- MSB_Unit_Cell_55/SD R1 cur_12_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_11 cur_2_d R2 VSS VDD MSB_Unit_Cell_11/QB MSB_Unit_Cell_11/Q MSB_Unit_Cell_11/OUT
+ OUT+ OUT- MSB_Unit_Cell_11/SD R1 cur_2_u VSS MSB_Unit_Cell
XCM_32_C_9 CM_32_C_9/SD0_1 CM_32_C_9/G1_2 CM_32_C_9/G1_1 CM_32_C_9/SD2_0 cur_2_d cur_2_u
+ VSS VDD cur_9_d cur_9_u CM_32_C
XLSBs_magic_TG_0 B2D LSBs_magic_TG_0/b1 LSBs_magic_TG_0/b1b LSBs_magic_TG_0/b2 LSBs_magic_TG_0/b2b
+ LSBs_magic_TG_0/b3 LSBs_magic_TG_0/b3b LSBs_magic_TG_0/b4 LSBs_magic_TG_0/b4b LSBs_magic_TG_0/b5
+ LSBs_magic_TG_0/b5b LSBs_magic_TG_0/b6 LSBs_magic_TG_0/b6b LSBs_magic_TG_0/OUT1
+ LSBs_magic_TG_0/OUT2 LSBs_magic_TG_0/OUT3 LSBs_magic_TG_0/OUT4 LSBs_magic_TG_0/OUT5
+ LSBs_magic_TG_0/OUT6 LSBs_magic_TG_0/G2 LSBs_magic_TG_0/SD2_2 LSBs_magic_TG_0/SD2_3
+ LSBs_magic_TG_0/SD2_5 LSBs_magic_TG_0/SD2_1 LSBs_magic_TG_0/SD2_4 LSBs_magic_TG_0/G1_2
+ LSBs_magic_TG_0/SD1_1 LSBs_magic_TG_0/G1_1 LSBs_magic_TG_0/SD3_1 LSBs_magic_TG_0/SDn_1
+ LSBs_magic_TG_0/SDn_2 LSBs_magic_TG_0/IT B1D B3D B4D B5D B6D OUT- OUT+ VSS VDD ITAIL
+ cur_1_d SEL LSBs_magic_TG_0/SDc_1 LSBs_magic_TG_0/Gc_1 LSBs_magic_TG_0/Gc_2 LSBs_magic_TG_0/SDc_2
+ cur_1_u LSBs_magic_TG
XINV_BUFF_22 B9 INV_BUFF_22/SD1 B9M VDD VSS INV_BUFF
XCM_32_C_12 CM_32_C_12/SD0_1 CM_32_C_12/G1_2 CM_32_C_12/G1_1 CM_32_C_12/SD2_0 cur_4_d
+ cur_4_u VSS VDD cur_14_d cur_14_u CM_32_C
XINV_BUFF_11 B3M INV_BUFF_11/SD1 B3D VDD VSS INV_BUFF
XMSB_Unit_Cell_45 cur_19_d R5 VSS VDD MSB_Unit_Cell_45/QB MSB_Unit_Cell_45/Q MSB_Unit_Cell_45/OUT
+ OUT+ OUT- MSB_Unit_Cell_45/SD R4 cur_19_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_56 cur_12_d R2 C0 VDD MSB_Unit_Cell_56/QB MSB_Unit_Cell_56/Q MSB_Unit_Cell_56/OUT
+ OUT+ OUT- MSB_Unit_Cell_56/SD R1 cur_12_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_34 cur_8_d R0 C4 VDD MSB_Unit_Cell_34/QB MSB_Unit_Cell_34/Q MSB_Unit_Cell_34/OUT
+ OUT+ OUT- MSB_Unit_Cell_34/SD VDD cur_8_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_12 cur_9_d R1 C5 VDD MSB_Unit_Cell_12/QB MSB_Unit_Cell_12/Q MSB_Unit_Cell_12/OUT
+ OUT+ OUT- MSB_Unit_Cell_12/SD R0 cur_9_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_23 cur_18_d VSS C4 VDD MSB_Unit_Cell_23/QB MSB_Unit_Cell_23/Q MSB_Unit_Cell_23/OUT
+ OUT+ OUT- MSB_Unit_Cell_23/SD R6 cur_18_u VSS MSB_Unit_Cell
XINV_BUFF_23 B7M INV_BUFF_23/SD1 B7D VDD VSS INV_BUFF
XINV_BUFF_12 B2M INV_BUFF_12/SD1 B2D VDD VSS INV_BUFF
XCM_32_C_13 CM_32_C_13/SD0_1 CM_32_C_13/G1_2 CM_32_C_13/G1_1 CM_32_C_13/SD2_0 cur_16_d
+ cur_16_u VSS VDD cur_17_d cur_17_u CM_32_C
XMSB_Unit_Cell_46 cur_21_d R5 C5 VDD MSB_Unit_Cell_46/QB MSB_Unit_Cell_46/Q MSB_Unit_Cell_46/OUT
+ OUT+ OUT- MSB_Unit_Cell_46/SD R4 cur_21_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_57 cur_11_d R0 C1 VDD MSB_Unit_Cell_57/QB MSB_Unit_Cell_57/Q MSB_Unit_Cell_57/OUT
+ OUT+ OUT- MSB_Unit_Cell_57/SD VDD cur_11_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_13 cur_9_d R1 C4 VDD MSB_Unit_Cell_13/QB MSB_Unit_Cell_13/Q MSB_Unit_Cell_13/OUT
+ OUT+ OUT- MSB_Unit_Cell_13/SD R0 cur_9_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_35 cur_8_d R0 C5 VDD MSB_Unit_Cell_35/QB MSB_Unit_Cell_35/Q MSB_Unit_Cell_35/OUT
+ OUT+ OUT- MSB_Unit_Cell_35/SD VDD cur_8_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_24 cur_19_d R6 VSS VDD MSB_Unit_Cell_24/QB MSB_Unit_Cell_24/Q MSB_Unit_Cell_24/OUT
+ OUT+ OUT- MSB_Unit_Cell_24/SD R5 cur_19_u VSS MSB_Unit_Cell
XINV_BUFF_24 B7 INV_BUFF_24/SD1 B7M VDD VSS INV_BUFF
XCM_32_C_14 CM_32_C_14/SD0_1 CM_32_C_14/G1_2 CM_32_C_14/G1_1 CM_32_C_14/SD2_0 cur_10_d
+ cur_10_u VSS VDD cur_11_d cur_11_u CM_32_C
XINV_BUFF_13 SEL_M INV_BUFF_13/SD1 SEL VDD VSS INV_BUFF
XMSB_Unit_Cell_47 cur_21_d R5 C4 VDD MSB_Unit_Cell_47/QB MSB_Unit_Cell_47/Q MSB_Unit_Cell_47/OUT
+ OUT+ OUT- MSB_Unit_Cell_47/SD R4 cur_21_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_14 cur_10_d R2 C5 VDD MSB_Unit_Cell_14/QB MSB_Unit_Cell_14/Q MSB_Unit_Cell_14/OUT
+ OUT+ OUT- MSB_Unit_Cell_14/SD R1 cur_10_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_36 cur_6_d R3 C6 VDD MSB_Unit_Cell_36/QB MSB_Unit_Cell_36/Q MSB_Unit_Cell_36/OUT
+ OUT+ OUT- MSB_Unit_Cell_36/SD R2 cur_6_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_58 cur_5_d R5 C1 VDD MSB_Unit_Cell_58/QB MSB_Unit_Cell_58/Q MSB_Unit_Cell_58/OUT
+ OUT+ OUT- MSB_Unit_Cell_58/SD R4 cur_5_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_25 cur_16_d VSS C2 VDD MSB_Unit_Cell_25/QB MSB_Unit_Cell_25/Q MSB_Unit_Cell_25/OUT
+ OUT+ OUT- MSB_Unit_Cell_25/SD R6 cur_16_u VSS MSB_Unit_Cell
XINV_BUFF_14 B10M INV_BUFF_14/SD1 B10D VDD VSS INV_BUFF
XINV_BUFF_25 B8 INV_BUFF_25/SD1 B8M VDD VSS INV_BUFF
XCM_32_C_15 CM_32_C_15/SD0_1 CM_32_C_15/G1_2 CM_32_C_15/G1_1 CM_32_C_15/SD2_0 cur_18_d
+ cur_18_u VSS VDD cur_19_d cur_19_u CM_32_C
XMSB_Unit_Cell_59 cur_11_d R0 C0 VDD MSB_Unit_Cell_59/QB MSB_Unit_Cell_59/Q MSB_Unit_Cell_59/OUT
+ OUT+ OUT- MSB_Unit_Cell_59/SD VDD cur_11_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_15 cur_10_d R2 C4 VDD MSB_Unit_Cell_15/QB MSB_Unit_Cell_15/Q MSB_Unit_Cell_15/OUT
+ OUT+ OUT- MSB_Unit_Cell_15/SD R1 cur_10_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_48 cur_7_d R4 VSS VDD MSB_Unit_Cell_48/QB MSB_Unit_Cell_48/Q MSB_Unit_Cell_48/OUT
+ OUT+ OUT- MSB_Unit_Cell_48/SD R3 cur_7_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_26 cur_15_d VSS C1 VDD MSB_Unit_Cell_26/QB MSB_Unit_Cell_26/Q MSB_Unit_Cell_26/OUT
+ OUT+ OUT- MSB_Unit_Cell_26/SD R6 cur_15_u VSS MSB_Unit_Cell
XMSB_Unit_Cell_37 cur_21_d R5 C3 VDD MSB_Unit_Cell_37/QB MSB_Unit_Cell_37/Q MSB_Unit_Cell_37/OUT
+ OUT+ OUT- MSB_Unit_Cell_37/SD R4 cur_21_u VSS MSB_Unit_Cell
XINV_BUFF_15 B12M INV_BUFF_15/SD1 B12D VDD VSS INV_BUFF
XCM_32_C_16 CM_32_C_16/SD0_1 CM_32_C_16/G1_2 CM_32_C_16/G1_1 CM_32_C_16/SD2_0 cur_20_d
+ cur_20_u VSS VDD cur_21_d cur_21_u CM_32_C
.ends

