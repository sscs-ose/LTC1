magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1453 -1298 1453 1298
<< metal3 >>
rect -453 293 453 298
rect -453 265 -448 293
rect -420 265 -386 293
rect -358 265 -324 293
rect -296 265 -262 293
rect -234 265 -200 293
rect -172 265 -138 293
rect -110 265 -76 293
rect -48 265 -14 293
rect 14 265 48 293
rect 76 265 110 293
rect 138 265 172 293
rect 200 265 234 293
rect 262 265 296 293
rect 324 265 358 293
rect 386 265 420 293
rect 448 265 453 293
rect -453 231 453 265
rect -453 203 -448 231
rect -420 203 -386 231
rect -358 203 -324 231
rect -296 203 -262 231
rect -234 203 -200 231
rect -172 203 -138 231
rect -110 203 -76 231
rect -48 203 -14 231
rect 14 203 48 231
rect 76 203 110 231
rect 138 203 172 231
rect 200 203 234 231
rect 262 203 296 231
rect 324 203 358 231
rect 386 203 420 231
rect 448 203 453 231
rect -453 169 453 203
rect -453 141 -448 169
rect -420 141 -386 169
rect -358 141 -324 169
rect -296 141 -262 169
rect -234 141 -200 169
rect -172 141 -138 169
rect -110 141 -76 169
rect -48 141 -14 169
rect 14 141 48 169
rect 76 141 110 169
rect 138 141 172 169
rect 200 141 234 169
rect 262 141 296 169
rect 324 141 358 169
rect 386 141 420 169
rect 448 141 453 169
rect -453 107 453 141
rect -453 79 -448 107
rect -420 79 -386 107
rect -358 79 -324 107
rect -296 79 -262 107
rect -234 79 -200 107
rect -172 79 -138 107
rect -110 79 -76 107
rect -48 79 -14 107
rect 14 79 48 107
rect 76 79 110 107
rect 138 79 172 107
rect 200 79 234 107
rect 262 79 296 107
rect 324 79 358 107
rect 386 79 420 107
rect 448 79 453 107
rect -453 45 453 79
rect -453 17 -448 45
rect -420 17 -386 45
rect -358 17 -324 45
rect -296 17 -262 45
rect -234 17 -200 45
rect -172 17 -138 45
rect -110 17 -76 45
rect -48 17 -14 45
rect 14 17 48 45
rect 76 17 110 45
rect 138 17 172 45
rect 200 17 234 45
rect 262 17 296 45
rect 324 17 358 45
rect 386 17 420 45
rect 448 17 453 45
rect -453 -17 453 17
rect -453 -45 -448 -17
rect -420 -45 -386 -17
rect -358 -45 -324 -17
rect -296 -45 -262 -17
rect -234 -45 -200 -17
rect -172 -45 -138 -17
rect -110 -45 -76 -17
rect -48 -45 -14 -17
rect 14 -45 48 -17
rect 76 -45 110 -17
rect 138 -45 172 -17
rect 200 -45 234 -17
rect 262 -45 296 -17
rect 324 -45 358 -17
rect 386 -45 420 -17
rect 448 -45 453 -17
rect -453 -79 453 -45
rect -453 -107 -448 -79
rect -420 -107 -386 -79
rect -358 -107 -324 -79
rect -296 -107 -262 -79
rect -234 -107 -200 -79
rect -172 -107 -138 -79
rect -110 -107 -76 -79
rect -48 -107 -14 -79
rect 14 -107 48 -79
rect 76 -107 110 -79
rect 138 -107 172 -79
rect 200 -107 234 -79
rect 262 -107 296 -79
rect 324 -107 358 -79
rect 386 -107 420 -79
rect 448 -107 453 -79
rect -453 -141 453 -107
rect -453 -169 -448 -141
rect -420 -169 -386 -141
rect -358 -169 -324 -141
rect -296 -169 -262 -141
rect -234 -169 -200 -141
rect -172 -169 -138 -141
rect -110 -169 -76 -141
rect -48 -169 -14 -141
rect 14 -169 48 -141
rect 76 -169 110 -141
rect 138 -169 172 -141
rect 200 -169 234 -141
rect 262 -169 296 -141
rect 324 -169 358 -141
rect 386 -169 420 -141
rect 448 -169 453 -141
rect -453 -203 453 -169
rect -453 -231 -448 -203
rect -420 -231 -386 -203
rect -358 -231 -324 -203
rect -296 -231 -262 -203
rect -234 -231 -200 -203
rect -172 -231 -138 -203
rect -110 -231 -76 -203
rect -48 -231 -14 -203
rect 14 -231 48 -203
rect 76 -231 110 -203
rect 138 -231 172 -203
rect 200 -231 234 -203
rect 262 -231 296 -203
rect 324 -231 358 -203
rect 386 -231 420 -203
rect 448 -231 453 -203
rect -453 -265 453 -231
rect -453 -293 -448 -265
rect -420 -293 -386 -265
rect -358 -293 -324 -265
rect -296 -293 -262 -265
rect -234 -293 -200 -265
rect -172 -293 -138 -265
rect -110 -293 -76 -265
rect -48 -293 -14 -265
rect 14 -293 48 -265
rect 76 -293 110 -265
rect 138 -293 172 -265
rect 200 -293 234 -265
rect 262 -293 296 -265
rect 324 -293 358 -265
rect 386 -293 420 -265
rect 448 -293 453 -265
rect -453 -298 453 -293
<< via3 >>
rect -448 265 -420 293
rect -386 265 -358 293
rect -324 265 -296 293
rect -262 265 -234 293
rect -200 265 -172 293
rect -138 265 -110 293
rect -76 265 -48 293
rect -14 265 14 293
rect 48 265 76 293
rect 110 265 138 293
rect 172 265 200 293
rect 234 265 262 293
rect 296 265 324 293
rect 358 265 386 293
rect 420 265 448 293
rect -448 203 -420 231
rect -386 203 -358 231
rect -324 203 -296 231
rect -262 203 -234 231
rect -200 203 -172 231
rect -138 203 -110 231
rect -76 203 -48 231
rect -14 203 14 231
rect 48 203 76 231
rect 110 203 138 231
rect 172 203 200 231
rect 234 203 262 231
rect 296 203 324 231
rect 358 203 386 231
rect 420 203 448 231
rect -448 141 -420 169
rect -386 141 -358 169
rect -324 141 -296 169
rect -262 141 -234 169
rect -200 141 -172 169
rect -138 141 -110 169
rect -76 141 -48 169
rect -14 141 14 169
rect 48 141 76 169
rect 110 141 138 169
rect 172 141 200 169
rect 234 141 262 169
rect 296 141 324 169
rect 358 141 386 169
rect 420 141 448 169
rect -448 79 -420 107
rect -386 79 -358 107
rect -324 79 -296 107
rect -262 79 -234 107
rect -200 79 -172 107
rect -138 79 -110 107
rect -76 79 -48 107
rect -14 79 14 107
rect 48 79 76 107
rect 110 79 138 107
rect 172 79 200 107
rect 234 79 262 107
rect 296 79 324 107
rect 358 79 386 107
rect 420 79 448 107
rect -448 17 -420 45
rect -386 17 -358 45
rect -324 17 -296 45
rect -262 17 -234 45
rect -200 17 -172 45
rect -138 17 -110 45
rect -76 17 -48 45
rect -14 17 14 45
rect 48 17 76 45
rect 110 17 138 45
rect 172 17 200 45
rect 234 17 262 45
rect 296 17 324 45
rect 358 17 386 45
rect 420 17 448 45
rect -448 -45 -420 -17
rect -386 -45 -358 -17
rect -324 -45 -296 -17
rect -262 -45 -234 -17
rect -200 -45 -172 -17
rect -138 -45 -110 -17
rect -76 -45 -48 -17
rect -14 -45 14 -17
rect 48 -45 76 -17
rect 110 -45 138 -17
rect 172 -45 200 -17
rect 234 -45 262 -17
rect 296 -45 324 -17
rect 358 -45 386 -17
rect 420 -45 448 -17
rect -448 -107 -420 -79
rect -386 -107 -358 -79
rect -324 -107 -296 -79
rect -262 -107 -234 -79
rect -200 -107 -172 -79
rect -138 -107 -110 -79
rect -76 -107 -48 -79
rect -14 -107 14 -79
rect 48 -107 76 -79
rect 110 -107 138 -79
rect 172 -107 200 -79
rect 234 -107 262 -79
rect 296 -107 324 -79
rect 358 -107 386 -79
rect 420 -107 448 -79
rect -448 -169 -420 -141
rect -386 -169 -358 -141
rect -324 -169 -296 -141
rect -262 -169 -234 -141
rect -200 -169 -172 -141
rect -138 -169 -110 -141
rect -76 -169 -48 -141
rect -14 -169 14 -141
rect 48 -169 76 -141
rect 110 -169 138 -141
rect 172 -169 200 -141
rect 234 -169 262 -141
rect 296 -169 324 -141
rect 358 -169 386 -141
rect 420 -169 448 -141
rect -448 -231 -420 -203
rect -386 -231 -358 -203
rect -324 -231 -296 -203
rect -262 -231 -234 -203
rect -200 -231 -172 -203
rect -138 -231 -110 -203
rect -76 -231 -48 -203
rect -14 -231 14 -203
rect 48 -231 76 -203
rect 110 -231 138 -203
rect 172 -231 200 -203
rect 234 -231 262 -203
rect 296 -231 324 -203
rect 358 -231 386 -203
rect 420 -231 448 -203
rect -448 -293 -420 -265
rect -386 -293 -358 -265
rect -324 -293 -296 -265
rect -262 -293 -234 -265
rect -200 -293 -172 -265
rect -138 -293 -110 -265
rect -76 -293 -48 -265
rect -14 -293 14 -265
rect 48 -293 76 -265
rect 110 -293 138 -265
rect 172 -293 200 -265
rect 234 -293 262 -265
rect 296 -293 324 -265
rect 358 -293 386 -265
rect 420 -293 448 -265
<< metal4 >>
rect -453 293 453 298
rect -453 265 -448 293
rect -420 265 -386 293
rect -358 265 -324 293
rect -296 265 -262 293
rect -234 265 -200 293
rect -172 265 -138 293
rect -110 265 -76 293
rect -48 265 -14 293
rect 14 265 48 293
rect 76 265 110 293
rect 138 265 172 293
rect 200 265 234 293
rect 262 265 296 293
rect 324 265 358 293
rect 386 265 420 293
rect 448 265 453 293
rect -453 231 453 265
rect -453 203 -448 231
rect -420 203 -386 231
rect -358 203 -324 231
rect -296 203 -262 231
rect -234 203 -200 231
rect -172 203 -138 231
rect -110 203 -76 231
rect -48 203 -14 231
rect 14 203 48 231
rect 76 203 110 231
rect 138 203 172 231
rect 200 203 234 231
rect 262 203 296 231
rect 324 203 358 231
rect 386 203 420 231
rect 448 203 453 231
rect -453 169 453 203
rect -453 141 -448 169
rect -420 141 -386 169
rect -358 141 -324 169
rect -296 141 -262 169
rect -234 141 -200 169
rect -172 141 -138 169
rect -110 141 -76 169
rect -48 141 -14 169
rect 14 141 48 169
rect 76 141 110 169
rect 138 141 172 169
rect 200 141 234 169
rect 262 141 296 169
rect 324 141 358 169
rect 386 141 420 169
rect 448 141 453 169
rect -453 107 453 141
rect -453 79 -448 107
rect -420 79 -386 107
rect -358 79 -324 107
rect -296 79 -262 107
rect -234 79 -200 107
rect -172 79 -138 107
rect -110 79 -76 107
rect -48 79 -14 107
rect 14 79 48 107
rect 76 79 110 107
rect 138 79 172 107
rect 200 79 234 107
rect 262 79 296 107
rect 324 79 358 107
rect 386 79 420 107
rect 448 79 453 107
rect -453 45 453 79
rect -453 17 -448 45
rect -420 17 -386 45
rect -358 17 -324 45
rect -296 17 -262 45
rect -234 17 -200 45
rect -172 17 -138 45
rect -110 17 -76 45
rect -48 17 -14 45
rect 14 17 48 45
rect 76 17 110 45
rect 138 17 172 45
rect 200 17 234 45
rect 262 17 296 45
rect 324 17 358 45
rect 386 17 420 45
rect 448 17 453 45
rect -453 -17 453 17
rect -453 -45 -448 -17
rect -420 -45 -386 -17
rect -358 -45 -324 -17
rect -296 -45 -262 -17
rect -234 -45 -200 -17
rect -172 -45 -138 -17
rect -110 -45 -76 -17
rect -48 -45 -14 -17
rect 14 -45 48 -17
rect 76 -45 110 -17
rect 138 -45 172 -17
rect 200 -45 234 -17
rect 262 -45 296 -17
rect 324 -45 358 -17
rect 386 -45 420 -17
rect 448 -45 453 -17
rect -453 -79 453 -45
rect -453 -107 -448 -79
rect -420 -107 -386 -79
rect -358 -107 -324 -79
rect -296 -107 -262 -79
rect -234 -107 -200 -79
rect -172 -107 -138 -79
rect -110 -107 -76 -79
rect -48 -107 -14 -79
rect 14 -107 48 -79
rect 76 -107 110 -79
rect 138 -107 172 -79
rect 200 -107 234 -79
rect 262 -107 296 -79
rect 324 -107 358 -79
rect 386 -107 420 -79
rect 448 -107 453 -79
rect -453 -141 453 -107
rect -453 -169 -448 -141
rect -420 -169 -386 -141
rect -358 -169 -324 -141
rect -296 -169 -262 -141
rect -234 -169 -200 -141
rect -172 -169 -138 -141
rect -110 -169 -76 -141
rect -48 -169 -14 -141
rect 14 -169 48 -141
rect 76 -169 110 -141
rect 138 -169 172 -141
rect 200 -169 234 -141
rect 262 -169 296 -141
rect 324 -169 358 -141
rect 386 -169 420 -141
rect 448 -169 453 -141
rect -453 -203 453 -169
rect -453 -231 -448 -203
rect -420 -231 -386 -203
rect -358 -231 -324 -203
rect -296 -231 -262 -203
rect -234 -231 -200 -203
rect -172 -231 -138 -203
rect -110 -231 -76 -203
rect -48 -231 -14 -203
rect 14 -231 48 -203
rect 76 -231 110 -203
rect 138 -231 172 -203
rect 200 -231 234 -203
rect 262 -231 296 -203
rect 324 -231 358 -203
rect 386 -231 420 -203
rect 448 -231 453 -203
rect -453 -265 453 -231
rect -453 -293 -448 -265
rect -420 -293 -386 -265
rect -358 -293 -324 -265
rect -296 -293 -262 -265
rect -234 -293 -200 -265
rect -172 -293 -138 -265
rect -110 -293 -76 -265
rect -48 -293 -14 -265
rect 14 -293 48 -265
rect 76 -293 110 -265
rect 138 -293 172 -265
rect 200 -293 234 -265
rect 262 -293 296 -265
rect 324 -293 358 -265
rect 386 -293 420 -265
rect 448 -293 453 -265
rect -453 -298 453 -293
<< end >>
