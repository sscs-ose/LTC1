* NGSPICE file created from Folded_Diff_Op_Amp_Layout_flat.ext - technology: gf180mcuC

.subckt Folded_Diff_Op_Amp_Layout_flat VDD BD IND IPD VSS VB4 VB2 VB3 VB1 VND VPD
+ IBIAS1 VBIASN VOUT VBM VCD IBIAS4 IBIAS3 IBS OUT_P OUT_N IBIAS2 IBIAS VCM IVS IB4
+ IB2 IB3 IB5 IN_P IN_N OUT1 OUT2
X0 VSS VB4.t32 IND.t42 VSS.t221 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X1 VDD.t1396 VDD.t1395 VDD.t1396 VDD.t1228 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X2 VDD IBIAS2.t122 OUT_N.t243 VDD.t43 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X3 VSS.t598 VSS.t597 VSS.t598 VSS.t493 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.28u
X4 VDD IBIAS2.t123 OUT_N.t242 VDD.t311 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X5 VDD IBIAS2.t124 OUT_P.t230 VDD.t314 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X6 VCD VCM.t0 VBM.t25 VSS.t599 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X7 IND IN_N.t0 BD.t58 VDD.t519 pfet_03v3 ad=1.65p pd=8.38u as=0.975p ps=4.27u w=3.75u l=0.28u
X8 VDD IBIAS2.t125 OUT_P.t229 VDD.t317 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X9 VDD IBIAS2.t126 OUT_P.t228 VDD.t91 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X10 IVS IBIAS3.t21 VDD.t807 VDD.t306 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X11 VDD VB1.t34 VPD.t16 VDD.t209 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X12 VDD.t1394 VDD.t1393 VDD.t1394 VDD.t1182 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X13 VB4 VB4.t12 VSS.t295 VSS.t294 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X14 VDD.t1392 VDD.t1391 VDD.t1392 VDD.t1209 pfet_03v3 ad=1.65p pd=8.38u as=0 ps=0 w=3.75u l=0.28u
X15 OUT_N OUT1.t36 VSS.t664 VSS.t313 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X16 OUT_N IBIAS2.t127 VDD.t276 VDD.t275 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X17 OUT_P IBIAS2.t128 VDD.t277 VDD.t50 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X18 OUT_N IBIAS2.t129 VDD.t18 VDD.t17 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X19 OUT_N IBIAS2.t130 VDD.t20 VDD.t19 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X20 a_29248_n7510.t3 OUT_N.t253 cap_mim_2f0fF c_width=21u c_length=21u
X21 OUT_N OUT1.t37 VSS.t665 VSS.t112 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X22 VSS OUT1.t38 OUT_N.t263 VSS.t7 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X23 OUT_P IBIAS2.t131 VDD.t22 VDD.t21 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X24 OUT_N IBIAS2.t132 VDD.t1088 VDD.t461 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X25 BD IBIAS.t12 VDD.t326 VDD.t114 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X26 OUT_P IBIAS2.t133 VDD.t1089 VDD.t263 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X27 BD IBIAS.t13 VDD.t521 VDD.t520 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X28 OUT_N IBIAS2.t134 VDD.t1090 VDD.t551 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X29 VCD VOUT.t2 VB1.t12 VSS.t6 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X30 VPD VB1.t35 VDD.t404 VDD.t290 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X31 VSS OUT2.t36 OUT_P.t16 VSS.t33 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X32 VDD IBIAS2.t135 OUT_N.t236 VDD.t355 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X33 OUT_P IBIAS2.t136 VDD.t659 VDD.t587 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X34 VDD IBIAS2.t137 OUT_N.t235 VDD.t28 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X35 IBIAS IBS.t9 VSS.t390 VSS.t389 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=1u
X36 VSS VB4.t34 IPD.t32 VSS.t221 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X37 VPD VB2.t33 OUT2.t25 VDD.t104 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X38 VSS.t596 VSS.t595 VSS.t596 VSS.t407 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X39 VDD IBIAS2.t138 OUT_P.t223 VDD.t98 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X40 IB5 IBIAS1.t2 VDD.t791 VDD.t790 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X41 VSS OUT1.t39 OUT_N.t264 VSS.t33 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X42 OUT1 VB2.t34 VND.t15 VDD.t102 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X43 VSS OUT2.t37 OUT_P.t17 VSS.t114 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X44 OUT_P IBIAS2.t139 VDD.t1055 VDD.t161 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X45 VDD IBIAS2.t140 OUT_P.t221 VDD.t577 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X46 VDD IBIAS4.t5 IB4.t17 VDD.t1013 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X47 VSS.t594 VSS.t593 VSS.t594 VSS.t413 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X48 VSS.t592 VSS.t591 VSS.t592 VSS.t456 nfet_03v3 ad=0.88p pd=4.88u as=0 ps=0 w=2u l=1u
X49 VSS VB4.t35 IND.t41 VSS.t192 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X50 VPD VB1.t36 VDD.t1133 VDD.t770 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X51 VDD IBIAS3.t22 IVS.t54 VDD.t406 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X52 OUT_P OUT2.t38 VSS.t134 VSS.t71 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X53 BD IBIAS.t14 VDD.t523 VDD.t522 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X54 VSS OUT2.t39 OUT_P.t4 VSS.t40 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X55 BD IN_P.t0 IPD.t51 VDD.t293 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X56 VSS.t590 VSS.t589 VSS.t590 VSS.t425 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X57 VDD IBIAS2.t141 OUT_N.t234 VDD.t176 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X58 VDD IBIAS3.t23 IVS.t53 VDD.t401 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X59 VB3 VB3.t10 IB3.t6 VSS.t331 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X60 VDD IBIAS2.t142 OUT_P.t220 VDD.t179 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X61 OUT_N IBIAS2.t143 VDD.t182 VDD.t86 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X62 VDD.t1390 VDD.t1389 VDD.t1390 VDD.t1174 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.56u
X63 IPD VB3.t17 OUT2.t17 VSS.t388 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X64 OUT1 VB3.t18 IND.t58 VSS.t392 nfet_03v3 ad=1.27p pd=6.64u as=1.27p ps=6.64u w=2.88u l=0.28u
X65 VDD IBIAS2.t144 OUT_N.t232 VDD.t241 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X66 VDD.t1388 VDD.t1387 VDD.t1388 VDD.t1191 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X67 VDD IBIAS3.t24 IVS.t52 VDD.t412 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X68 VB1 VOUT.t3 VCD.t11 VSS.t353 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X69 OUT_N OUT1.t40 VSS.t113 VSS.t112 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X70 VDD IBIAS2.t145 OUT_P.t219 VDD.t317 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X71 VDD IBIAS2.t110 IBIAS2.t111 VDD.t7 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X72 VDD.t1386 VDD.t1385 VDD.t1386 VDD.t1250 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X73 VBM VCM.t1 VCD.t41 VSS.t3 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X74 VSS VB4.t36 IPD.t31 VSS.t221 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X75 OUT_N IBIAS2.t146 VDD.t561 VDD.t433 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X76 VSS VBIASN.t5 VCD.t53 VSS.t659 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X77 VCD VCM.t2 VBM.t24 VSS.t5 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X78 OUT_N IBIAS2.t147 VDD.t260 VDD.t252 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X79 IPD IN_P.t1 BD.t26 VDD.t108 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X80 IND VB4.t37 VSS.t287 VSS.t164 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X81 VDD IBIAS2.t108 IBIAS2.t109 VDD.t1107 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X82 OUT_P IBIAS2.t148 VDD.t262 VDD.t261 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X83 OUT_P IBIAS2.t149 VDD.t264 VDD.t263 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X84 VDD IBIAS2.t150 OUT_N.t229 VDD.t457 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X85 VCD VBIASN.t6 VSS.t663 VSS.t662 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X86 VDD IBIAS.t15 BD.t4 VDD.t111 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X87 OUT_P IBIAS2.t151 VDD.t682 VDD.t163 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X88 VDD IBIAS2.t152 OUT_N.t228 VDD.t46 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X89 VSS VBIASN.t7 IBIAS4.t0 VSS.t46 nfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=1u
X90 VSS IVS.t74 IVS.t75 VSS.t620 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X91 VSS.t588 VSS.t587 VSS.t588 VSS.t404 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X92 VSS VB4.t38 IND.t40 VSS.t192 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X93 IPD VB4.t39 VSS.t284 VSS.t209 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X94 VDD.t1384 VDD.t1383 VDD.t1384 VDD.t1284 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X95 VDD IBIAS2.t153 OUT_N.t227 VDD.t577 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X96 a_25078_n6312# a_24798_n7414# VDD.t580 ppolyf_u r_width=1u r_length=5u
X97 IND IN_N.t1 BD.t57 VDD.t353 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X98 VND VB2.t35 OUT1.t26 VDD.t309 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X99 VSS OUT1.t41 OUT_N.t31 VSS.t114 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X100 VCD VOUT.t4 VB1.t24 VSS.t141 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X101 OUT_N IBIAS2.t154 VDD.t1025 VDD.t86 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X102 VDD IBIAS2.t155 OUT_N.t225 VDD.t88 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X103 OUT_N OUT1.t42 VSS.t117 VSS.t89 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X104 VSS OUT1.t43 OUT_N.t33 VSS.t93 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X105 VDD IBIAS2.t156 OUT_N.t224 VDD.t127 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X106 IVS IBIAS3.t25 VDD.t170 VDD.t109 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X107 IND VB4.t40 VSS.t283 VSS.t197 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X108 VDD.t1382 VDD.t1381 VDD.t1382 VDD.t1228 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X109 VDD.t1380 VDD.t1379 VDD.t1380 VDD.t1182 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X110 VDD VB1.t37 VPD.t13 VDD.t282 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X111 VSS OUT1.t44 OUT_N.t34 VSS.t7 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X112 VDD IBIAS.t16 BD.t5 VDD.t267 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X113 VSS.t586 VSS.t585 VSS.t586 VSS.t433 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X114 VDD IBIAS2.t106 IBIAS2.t107 VDD.t199 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X115 a_29248_n5498.t1 OUT_P.t270 cap_mim_2f0fF c_width=21u c_length=21u
X116 OUT_N IBIAS2.t157 VDD.t962 VDD.t465 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X117 VCD VOUT.t5 VB1.t30 VSS.t599 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X118 VSS.t584 VSS.t583 VSS.t584 VSS.t430 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X119 VDD.t1378 VDD.t1376 VDD.t1378 VDD.t1377 pfet_03v3 ad=1.76p pd=8.88u as=0 ps=0 w=4u l=0.28u
X120 VB4 VB4.t10 VSS.t282 VSS.t281 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X121 VB1 VOUT.t6 VCD.t7 VSS.t142 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X122 VDD.t1375 VDD.t1374 VDD.t1375 VDD.t1194 pfet_03v3 ad=1.65p pd=8.38u as=0 ps=0 w=3.75u l=0.28u
X123 VDD IBIAS2.t158 OUT_P.t215 VDD.t675 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X124 IPD VB4.t42 VSS.t280 VSS.t209 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X125 VSS OUT2.t40 OUT_P.t5 VSS.t24 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X126 VDD.t1373 VDD.t1372 VDD.t1373 VDD.t1291 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X127 VDD.t1371 VDD.t1370 VDD.t1371 VDD.t1169 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X128 VDD IBIAS2.t159 OUT_N.t222 VDD.t0 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X129 OUT_P IBIAS2.t160 VDD.t1412 VDD.t52 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X130 VDD IBIAS2.t161 OUT_N.t221 VDD.t457 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X131 OUT_N IBIAS2.t162 VDD.t733 VDD.t465 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X132 VDD IBIAS2.t163 OUT_N.t219 VDD.t67 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X133 VDD.t1369 VDD.t1368 VDD.t1369 VDD.t1279 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X134 VB3 VB3.t12 IB3.t5 VSS.t332 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X135 VSS.t582 VSS.t581 VSS.t582 VSS.t407 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X136 OUT_N IBIAS2.t164 VDD.t736 VDD.t227 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X137 VDD IBIAS4.t6 IB4.t16 VDD.t1013 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X138 VSS OUT1.t45 OUT_N.t35 VSS.t13 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X139 VDD IBIAS2.t165 OUT_N.t217 VDD.t43 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X140 BD IBIAS.t17 VDD.t1102 VDD.t520 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X141 IND VB4.t43 VSS.t279 VSS.t162 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X142 OUT_P IBIAS2.t166 VDD.t967 VDD.t19 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X143 VBM VCM.t3 VCD.t39 VSS.t3 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X144 VB1 VOUT.t7 VCD.t55 VSS.t140 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X145 IND VB4.t44 VSS.t278 VSS.t197 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X146 OUT_P IBIAS2.t167 VDD.t968 VDD.t81 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X147 VDD IBIAS4.t7 IB4.t15 VDD.t1013 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X148 IVS IVS.t72 VSS.t637 VSS.t636 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X149 VDD IBIAS2.t168 OUT_P.t211 VDD.t28 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X150 VSS IVS.t77 IBIAS2.t112 VSS.t346 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X151 BD IN_P.t2 IPD.t39 VDD.t107 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X152 OUT_N OUT1.t46 VSS.t92 VSS.t91 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X153 OUT_P IBIAS2.t169 VDD.t31 VDD.t17 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X154 VDD IBIAS2.t170 OUT_P.t209 VDD.t32 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X155 VND VB2.t36 OUT1.t30 VDD.t104 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X156 OUT_N IBIAS2.t171 VDD.t566 VDD.t437 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X157 VDD IBIAS3.t26 IVS.t50 VDD.t401 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X158 OUT_N IBIAS2.t172 VDD.t568 VDD.t567 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X159 VSS.t580 VSS.t579 VSS.t580 VSS.t477 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.28u
X160 BD IN_P.t3 IPD.t40 VDD.t530 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X161 OUT_N IBIAS2.t173 VDD.t569 VDD.t148 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X162 VDD IBIAS2.t174 OUT_P.t208 VDD.t295 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X163 OUT_N IBIAS2.t175 VDD.t455 VDD.t454 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X164 OUT2.t24 a_29248_n5498.t1 VDD.t697 ppolyf_u r_width=1u r_length=6.2u
X165 IBIAS3 IBIAS3.t19 VDD.t575 VDD.t574 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X166 VSS.t578 VSS.t576 VSS.t578 VSS.t577 nfet_03v3 ad=0.26p pd=1.52u as=0 ps=0 w=1u l=0.28u
X167 OUT_N IBIAS2.t176 VDD.t456 VDD.t435 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X168 OUT2 VB2.t37 VPD.t31 VDD.t102 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X169 VDD IBIAS3.t28 IVS.t49 VDD.t401 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X170 OUT_P IBIAS2.t177 VDD.t482 VDD.t433 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X171 VND VB1.t38 VDD.t1406 VDD.t770 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X172 VDD IBIAS2.t104 IBIAS2.t105 VDD.t199 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X173 IBIAS2 IBIAS2.t102 VDD.t518 VDD.t336 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X174 VDD IBIAS2.t179 OUT_N.t211 VDD.t483 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X175 VSS.t575 VSS.t574 VSS.t575 VSS.t416 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X176 VSS.t573 VSS.t572 VSS.t573 VSS.t493 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.28u
X177 IND VB4.t45 VSS.t277 VSS.t164 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X178 OUT_N IBIAS2.t180 VDD.t486 VDD.t275 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X179 VSS.t571 VSS.t570 VSS.t571 VSS.t413 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X180 OUT_P OUT2.t41 VSS.t80 VSS.t79 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X181 VSS OUT1.t47 OUT_N.t19 VSS.t93 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X182 OUT_P IBIAS2.t181 VDD.t118 VDD.t117 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X183 IVS IBIAS3.t29 VDD.t1091 VDD.t364 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X184 IB3 VB3.t4 VB3.t5 VSS.t399 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X185 OUT_N OUT1.t48 VSS.t96 VSS.t79 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X186 VDD IBIAS2.t182 OUT_P.t205 VDD.t119 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X187 VSS.t569 VSS.t568 VSS.t569 VSS.t410 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X188 VSS VB4.t46 IPD.t28 VSS.t192 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X189 VB1 VB1.t4 VDD.t789 VDD.t788 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X190 IPD VB3.t20 OUT2.t18 VSS.t1 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X191 OUT2 VB3.t21 IPD.t48 VSS.t392 nfet_03v3 ad=1.27p pd=6.64u as=1.27p ps=6.64u w=2.88u l=0.28u
X192 VDD IBIAS2.t183 OUT_N.t209 VDD.t122 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X193 VCD VOUT.t8 VB1.t17 VSS.t599 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X194 IND VB3.t22 OUT1.t15 VSS.t1 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X195 VDD IBIAS2.t184 OUT_P.t204 VDD.t60 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X196 VCD VOUT.t9 VB1.t6 VSS.t5 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X197 OUT1 VB2.t38 VND.t12 VDD.t103 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X198 OUT_P IBIAS2.t185 VDD.t64 VDD.t63 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X199 VB4 VB4.t8 VSS.t274 VSS.t273 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X200 VDD.t1367 VDD.t1366 VDD.t1367 VDD.t1179 pfet_03v3 ad=1.65p pd=8.38u as=0 ps=0 w=3.75u l=0.28u
X201 VSS.t567 VSS.t566 VSS.t567 VSS.t404 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X202 VSS OUT2.t42 OUT_P.t7 VSS.t10 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X203 VDD IBIAS2.t100 IBIAS2.t101 VDD.t515 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X204 VSS.t565 VSS.t564 VSS.t565 VSS.t413 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X205 VSS VB4.t48 IPD.t27 VSS.t159 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X206 IND VB3.t23 OUT1.t16 VSS.t385 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X207 IVS IBIAS3.t30 VDD.t360 VDD.t109 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X208 a_24798_n4340# a_23622_n5442# VDD.t766 ppolyf_u r_width=1u r_length=5u
X209 BD IBIAS.t18 VDD.t1103 VDD.t522 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X210 VSS OUT2.t43 OUT_P.t31 VSS.t24 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X211 OUT_P IBIAS2.t186 VDD.t65 VDD.t5 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X212 VDD.t1365 VDD.t1364 VDD.t1365 VDD.t1174 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.56u
X213 VDD IBIAS2.t187 OUT_P.t201 VDD.t88 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X214 IBIAS2 IVS.t78 VSS.t642 VSS.t342 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X215 VSS.t563 VSS.t562 VSS.t563 VSS.t416 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X216 OUT_N OUT1.t49 VSS.t97 VSS.t38 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X217 OUT_P IBIAS2.t188 VDD.t612 VDD.t117 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X218 IVS IBIAS3.t31 VDD.t110 VDD.t109 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X219 VDD IBIAS2.t189 OUT_P.t199 VDD.t469 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X220 VSS.t561 VSS.t560 VSS.t561 VSS.t419 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X221 VPD VB2.t39 OUT2.t6 VDD.t309 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X222 VSS OUT1.t50 OUT_N.t22 VSS.t98 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X223 VSS OUT2.t44 OUT_P.t32 VSS.t28 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X224 VSS VB4.t49 IPD.t26 VSS.t221 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X225 OUT_P IBIAS2.t190 VDD.t741 VDD.t72 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X226 VDD IBIAS1.t3 VBIASN.t0 VDD.t746 pfet_03v3 ad=1.04p pd=4.52u as=1.76p ps=8.88u w=4u l=0.56u
X227 VSS OUT2.t45 OUT_P.t33 VSS.t98 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X228 VDD.t1363 VDD.t1362 VDD.t1363 VDD.t1145 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X229 VDD.t1361 VDD.t1360 VDD.t1361 VDD.t1279 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X230 IB2 VB2.t30 VB2.t31 VDD.t792 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X231 VSS OUT2.t46 OUT_P.t34 VSS.t16 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X232 VDD IBIAS2.t191 OUT_P.t197 VDD.t38 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X233 VSS.t559 VSS.t558 VSS.t559 VSS.t404 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X234 VSS VB4.t50 IND.t39 VSS.t192 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X235 VDD.t1359 VDD.t1358 VDD.t1359 VDD.t1279 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X236 VSS VB4.t26 VB4.t27 VSS.t264 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X237 VDD IBIAS2.t98 IBIAS2.t99 VDD.t173 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X238 VDD.t1357 VDD.t1356 VDD.t1357 VDD.t1270 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X239 VDD IBIAS2.t192 OUT_N.t208 VDD.t179 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X240 VPD VB2.t40 OUT2.t7 VDD.t354 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X241 VDD IBIAS2.t193 OUT_P.t196 VDD.t376 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X242 OUT_P OUT2.t47 VSS.t333 VSS.t91 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X243 OUT_N IBIAS2.t194 VDD.t631 VDD.t461 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X244 VDD.t1355 VDD.t1354 VDD.t1355 VDD.t1206 pfet_03v3 ad=0.13p pd=1.02u as=0 ps=0 w=0.5u l=0.28u
X245 VDD IBIAS2.t195 OUT_N.t206 VDD.t60 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X246 OUT1.t20 a_29248_n7510.t1 VDD.t697 ppolyf_u r_width=1u r_length=6.2u
X247 IPD IN_P.t4 BD.t20 VDD.t294 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X248 VDD IBIAS2.t196 OUT_P.t195 VDD.t0 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X249 OUT_P IBIAS2.t197 VDD.t822 VDD.t780 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X250 VSS VB4.t51 IND.t38 VSS.t159 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X251 IBIAS3 IBIAS3.t17 VDD.t831 VDD.t574 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X252 VDD IBIAS3.t33 IVS.t45 VDD.t186 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X253 OUT2 VB3.t24 IPD.t42 VSS.t391 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X254 VDD IBIAS2.t198 OUT_P.t193 VDD.t221 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X255 VSS.t557 VSS.t556 VSS.t557 VSS.t419 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X256 VCD VOUT.t10 VB1.t9 VSS.t5 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X257 IBS IBIAS1.t4 VDD.t696 VDD.t695 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X258 IBIAS3 IBIAS3.t15 VDD.t1132 VDD.t574 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X259 VDD.t1353 VDD.t1352 VDD.t1353 VDD.t1145 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X260 VDD IBIAS2.t199 OUT_N.t205 VDD.t57 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X261 VDD IBIAS2.t200 OUT_N.t204 VDD.t469 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X262 VB4 IB5.t10 IB5.t11 VSS.t616 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X263 IND IN_N.t2 BD.t56 VDD.t37 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X264 VDD IBIAS2.t201 OUT_P.t192 VDD.t224 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X265 VDD IBIAS2.t202 OUT_N.t203 VDD.t54 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X266 VDD IBIAS2.t203 OUT_P.t191 VDD.t28 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X267 IVS IBIAS3.t35 VDD.t365 VDD.t364 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X268 VSS IVS.t70 IVS.t71 VSS.t624 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X269 VDD IBIAS.t19 BD.t7 VDD.t137 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X270 IPD VB4.t52 VSS.t261 VSS.t209 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X271 IND VB4.t53 VSS.t260 VSS.t209 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X272 OUT_P OUT2.t48 VSS.t334 VSS.t103 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X273 OUT_N OUT1.t51 VSS.t102 VSS.t101 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X274 VDD IBIAS2.t204 OUT_N.t202 VDD.t67 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X275 VB2 VB2.t14 IB2.t14 VDD.t783 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X276 OUT_P IBIAS2.t205 VDD.t491 VDD.t41 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X277 IVS IBIAS3.t36 VDD.t1078 VDD.t364 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X278 IBIAS2 IVS.t79 VSS.t643 VSS.t344 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X279 OUT2 VB2.t42 VPD.t22 VDD.t103 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X280 OUT2 VB3.t25 IPD.t43 VSS.t0 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X281 OUT_N OUT1.t52 VSS.t104 VSS.t103 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X282 VDD.t1351 VDD.t1350 VDD.t1351 VDD.t1247 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X283 VPD VB2.t43 OUT2.t31 VDD.t354 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X284 OUT_N IBIAS2.t206 VDD.t493 VDD.t492 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X285 IBIAS2 IBIAS2.t96 VDD.t196 VDD.t195 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X286 VSS OUT2.t49 OUT_P.t238 VSS.t40 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X287 VSS OUT2.t50 OUT_P.t239 VSS.t10 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X288 IBIAS2 IBIAS2.t94 VDD.t143 VDD.t142 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X289 IND VB4.t54 VSS.t259 VSS.t197 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X290 IPD VB4.t55 VSS.t258 VSS.t164 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X291 VDD IBIAS2.t209 OUT_N.t200 VDD.t494 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X292 OUT_N IBIAS2.t210 VDD.t487 VDD.t385 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X293 VSS.t555 VSS.t554 VSS.t555 VSS.t425 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X294 OUT_P IBIAS2.t211 VDD.t488 VDD.t94 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X295 IBIAS2 IBIAS2.t92 VDD.t141 VDD.t140 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X296 IVS IBIAS3.t37 VDD.t946 VDD.t184 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X297 OUT_P OUT2.t51 VSS.t84 VSS.t83 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X298 VDD.t1349 VDD.t1348 VDD.t1349 VDD.t1212 pfet_03v3 ad=1.76p pd=8.88u as=0 ps=0 w=4u l=0.28u
X299 VDD IBIAS2.t213 OUT_N.t198 VDD.t83 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X300 VBM VCM.t4 VCD.t38 VSS.t142 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X301 OUT_P IBIAS2.t214 VDD.t53 VDD.t52 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X302 VDD.t399 VDD.t400 VDD.t396 ppolyf_u r_width=1u r_length=5u
X303 VCD VBIASN.t8 VSS.t50 VSS.t49 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X304 VSS VB4.t24 VB4.t25 VSS.t255 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X305 BD IN_N.t3 IND.t44 VDD.t361 pfet_03v3 ad=0.975p pd=4.27u as=1.65p ps=8.38u w=3.75u l=0.28u
X306 VDD.t1347 VDD.t1346 VDD.t1347 VDD.t1261 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X307 VDD IBIAS2.t215 OUT_P.t187 VDD.t54 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X308 VDD IBIAS2.t216 OUT_P.t186 VDD.t57 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X309 VDD.t1345 VDD.t1344 VDD.t1345 VDD.t1242 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X310 VSS.t553 VSS.t552 VSS.t553 VSS.t442 nfet_03v3 ad=0.52p pd=2.52u as=0 ps=0 w=2u l=1u
X311 VDD.t1343 VDD.t1342 VDD.t1343 VDD.t1188 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X312 OUT1 VB3.t26 IND.t55 VSS.t384 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X313 VDD IBIAS2.t217 OUT_P.t185 VDD.t38 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X314 BD IN_P.t5 IPD.t65 VDD.t537 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X315 OUT_P IBIAS2.t218 VDD.t42 VDD.t41 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X316 VDD IBIAS2.t219 OUT_P.t183 VDD.t43 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X317 VB1 VOUT.t11 VCD.t0 VSS.t3 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X318 VSS VB4.t56 IND.t37 VSS.t221 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X319 VSS OUT2.t52 OUT_P.t9 VSS.t33 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X320 VSS OUT2.t53 OUT_P.t10 VSS.t10 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X321 VDD.t1341 VDD.t1340 VDD.t1341 VDD.t1284 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X322 VSS.t551 VSS.t550 VSS.t551 VSS.t477 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.28u
X323 VDD IBIAS2.t220 OUT_N.t197 VDD.t46 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X324 VDD.t1339 VDD.t1338 VDD.t1339 VDD.t1270 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X325 VSS.t549 VSS.t548 VSS.t549 VSS.t540 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.28u
X326 OUT_P OUT2.t54 VSS.t90 VSS.t89 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X327 OUT_P IBIAS2.t221 VDD.t49 VDD.t17 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X328 OUT_N IBIAS2.t222 VDD.t51 VDD.t50 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X329 OUT_P IBIAS2.t223 VDD.t463 VDD.t461 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X330 VDD.t1337 VDD.t1336 VDD.t1337 VDD.t1284 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X331 OUT_P IBIAS2.t224 VDD.t464 VDD.t70 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X332 OUT_P IBIAS2.t225 VDD.t466 VDD.t465 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X333 a_24798_n4340# a_25078_n5442# VDD.t580 ppolyf_u r_width=1u r_length=5u
X334 VDD.t1335 VDD.t1334 VDD.t1335 VDD.t1270 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X335 VSS VB4.t57 IPD.t23 VSS.t192 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X336 VDD IBIAS2.t226 OUT_N.t195 VDD.t91 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X337 VSS.t547 VSS.t546 VSS.t547 VSS.t416 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X338 BD IBIAS.t20 VDD.t330 VDD.t329 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X339 OUT_P OUT2.t55 VSS.t368 VSS.t89 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X340 VSS.t545 VSS.t544 VSS.t545 VSS.t430 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X341 VDD.t1333 VDD.t1332 VDD.t1333 VDD.t1182 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X342 IVS IBIAS3.t38 VDD.t539 VDD.t531 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X343 VSS.t543 VSS.t542 VSS.t543 VSS.t493 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.28u
X344 OUT_P IBIAS2.t227 VDD.t95 VDD.t94 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X345 IVS IBIAS3.t39 VDD.t208 VDD.t207 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X346 OUT_P IBIAS2.t228 VDD.t97 VDD.t96 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X347 VDD.t1331 VDD.t1330 VDD.t1331 VDD.t1142 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X348 IBIAS1 IBIAS1.t0 VDD.t784 VDD.t581 pfet_03v3 ad=1.76p pd=8.88u as=1.04p ps=4.52u w=4u l=0.56u
X349 OUT_P IBIAS2.t229 VDD.t73 VDD.t72 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X350 IVS IBIAS3.t40 VDD.t213 VDD.t130 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X351 VCD VCM.t5 VBM.t23 VSS.t599 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X352 IND VB3.t27 OUT1.t34 VSS.t385 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X353 VDD IBIAS2.t230 OUT_P.t175 VDD.t74 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X354 VDD IBIAS.t21 BD.t65 VDD.t111 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X355 VDD IBIAS2.t231 OUT_N.t194 VDD.t77 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X356 IND VB4.t58 VSS.t250 VSS.t209 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X357 VDD IBIAS2.t90 IBIAS2.t91 VDD.t199 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X358 OUT_N IBIAS2.t232 VDD.t815 VDD.t72 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X359 VDD IBIAS2.t233 OUT_N.t192 VDD.t311 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X360 VSS OUT2.t56 OUT_P.t245 VSS.t114 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X361 VDD IBIAS2.t234 OUT_P.t174 VDD.t666 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X362 OUT1 VB2.t44 VND.t11 VDD.t305 pfet_03v3 ad=1.38p pd=7.14u as=1.38p ps=7.14u w=3.13u l=0.28u
X363 VDD IBIAS2.t235 OUT_P.t173 VDD.t241 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X364 VDD IBIAS2.t88 IBIAS2.t89 VDD.t7 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X365 VDD.t1329 VDD.t1328 VDD.t1329 VDD.t1169 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X366 VDD IBIAS2.t236 OUT_N.t191 VDD.t317 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X367 VDD.t1327 VDD.t1326 VDD.t1327 VDD.t1250 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X368 OUT_P IBIAS2.t237 VDD.t930 VDD.t430 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X369 VPD VB2.t45 OUT2.t32 VDD.t310 pfet_03v3 ad=1.38p pd=7.14u as=1.38p ps=7.14u w=3.13u l=0.28u
X370 VDD IBIAS3.t13 IBIAS3.t14 VDD.t320 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X371 VSS.t541 VSS.t539 VSS.t541 VSS.t540 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.28u
X372 VDD IBIAS2.t238 OUT_N.t190 VDD.t669 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X373 IPD VB4.t59 VSS.t249 VSS.t197 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X374 VDD IBIAS2.t239 OUT_P.t171 VDD.t119 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X375 OUT_N IBIAS2.t240 VDD.t925 VDD.t261 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X376 VND VB2.t46 OUT1.t8 VDD.t354 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X377 VSS OUT1.t53 OUT_N.t25 VSS.t16 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X378 IND IN_N.t4 BD.t54 VDD.t519 pfet_03v3 ad=1.65p pd=8.38u as=0.975p ps=4.27u w=3.75u l=0.28u
X379 VDD IBIAS3.t41 IVS.t38 VDD.t204 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X380 VDD IBIAS2.t241 OUT_N.t188 VDD.t83 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X381 BD IN_N.t5 IND.t51 VDD.t537 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X382 VSS.t538 VSS.t537 VSS.t538 VSS.t413 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X383 VSS OUT1.t54 OUT_N.t26 VSS.t93 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X384 IVS IVS.t68 VSS.t623 VSS.t62 nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=1u
X385 IB4 IB4.t8 VSS.t671 VSS.t618 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X386 VDD.t1325 VDD.t1324 VDD.t1325 VDD.t1185 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X387 OUT_P IBIAS2.t242 VDD.t87 VDD.t86 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X388 VB1 VOUT.t12 VCD.t59 VSS.t142 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X389 VDD IBIAS2.t243 OUT_P.t169 VDD.t88 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X390 VSS IB4.t19 IBIAS3.t0 VSS.t339 nfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=1u
X391 VSS IVS.t81 IBIAS2.t115 VSS.t349 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X392 IBIAS IBIAS.t10 VDD.t325 VDD.t324 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X393 IBIAS2 IBIAS2.t86 VDD.t203 VDD.t202 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X394 VSS OUT2.t57 OUT_P.t246 VSS.t10 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X395 BD IN_P.t6 IPD.t66 VDD.t292 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X396 VDD IBIAS2.t245 OUT_P.t168 VDD.t355 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X397 OUT_N IBIAS2.t246 VDD.t863 VDD.t63 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X398 OUT_P OUT2.t58 VSS.t373 VSS.t22 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X399 OUT1 VB3.t28 IND.t70 VSS.t391 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X400 VSS.t536 VSS.t535 VSS.t536 VSS.t416 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X401 VDD IBIAS2.t84 IBIAS2.t85 VDD.t199 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X402 OUT_N IBIAS2.t247 VDD.t864 VDD.t492 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X403 IPD VB3.t29 OUT2.t35 VSS.t385 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X404 OUT1 VB3.t30 IND.t67 VSS.t0 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X405 VDD.t1323 VDD.t1322 VDD.t1323 VDD.t1291 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X406 OUT_P OUT2.t59 VSS.t135 VSS.t91 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X407 VCD VCM.t6 VBM.t22 VSS.t5 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X408 VDD IBIAS2.t248 OUT_N.t185 VDD.t675 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X409 VDD IBIAS2.t249 OUT_P.t167 VDD.t675 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X410 OUT2 VB2.t47 VPD.t23 VDD.t102 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X411 OUT_N OUT1.t55 VSS.t109 VSS.t22 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X412 VSS.t534 VSS.t533 VSS.t534 VSS.t404 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X413 OUT_P OUT2.t60 VSS.t136 VSS.t68 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X414 OUT_N OUT1.t56 VSS.t110 VSS.t89 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X415 OUT_P IBIAS2.t250 VDD.t689 VDD.t433 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X416 VDD.t1321 VDD.t1320 VDD.t1321 VDD.t1247 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X417 VDD.t1319 VDD.t1318 VDD.t1319 VDD.t1291 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X418 VDD IBIAS2.t251 OUT_N.t184 VDD.t179 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X419 VDD IBIAS2.t252 OUT_P.t165 VDD.t483 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X420 IVS IBIAS3.t42 VDD.t1085 VDD.t207 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X421 IND IN_N.t6 BD.t52 VDD.t108 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X422 OUT_P IBIAS2.t253 VDD.t501 VDD.t227 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X423 VSS.t532 VSS.t531 VSS.t532 VSS.t433 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X424 VSS.t530 VSS.t528 VSS.t530 VSS.t529 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.28u
X425 VB2 VB2.t12 IB2.t13 VDD.t36 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X426 BD IN_P.t7 IPD.t67 VDD.t293 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X427 OUT1 VB3.t31 IND.t68 VSS.t392 nfet_03v3 ad=1.27p pd=6.64u as=1.27p ps=6.64u w=2.88u l=0.28u
X428 OUT_P IBIAS2.t254 VDD.t506 VDD.t275 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X429 IVS IBIAS3.t43 VDD.t1106 VDD.t207 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X430 VDD VB1.t40 VND.t30 VDD.t209 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X431 VB4 VB4.t6 VSS.t248 VSS.t247 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X432 OUT_N IBIAS2.t255 VDD.t507 VDD.t358 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X433 IBIAS2 IBIAS2.t82 VDD.t527 VDD.t526 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X434 VSS.t527 VSS.t526 VSS.t527 VSS.t493 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.28u
X435 OUT_P OUT2.t61 VSS.t137 VSS.t79 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X436 IPD IN_P.t8 BD.t59 VDD.t353 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X437 VDD IBIAS2.t257 OUT_P.t162 VDD.t508 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X438 OUT_P IBIAS2.t258 VDD.t502 VDD.t379 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X439 VDD IBIAS2.t259 OUT_N.t182 VDD.t32 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X440 VSS VB4.t61 IND.t36 VSS.t221 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X441 OUT_P IBIAS2.t260 VDD.t505 VDD.t437 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X442 IB5 IBIAS1.t6 VDD.t1398 VDD.t1397 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X443 OUT_P IBIAS2.t261 VDD.t431 VDD.t430 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X444 OUT_N IBIAS2.t262 VDD.t432 VDD.t5 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X445 IBIAS2 IBIAS2.t80 VDD.t525 VDD.t171 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X446 VDD.t1071 VDD.t1072 VDD.t934 ppolyf_u r_width=1u r_length=6.2u
X447 VDD.t15 VDD.t16 VDD.t14 ppolyf_u r_width=1u r_length=5u
X448 VDD.t1317 VDD.t1316 VDD.t1317 VDD.t1201 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X449 VB1 VOUT.t13 VCD.t48 VSS.t142 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X450 VDD.t1315 VDD.t1314 VDD.t1315 VDD.t1153 pfet_03v3 ad=0.814p pd=3.65u as=0 ps=0 w=3.13u l=0.56u
X451 IPD VB4.t62 VSS.t241 VSS.t162 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X452 OUT_N IBIAS2.t264 VDD.t434 VDD.t433 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X453 BD IN_N.t7 IND.t5 VDD.t166 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X454 VSS VB4.t63 IPD.t20 VSS.t192 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X455 IBIAS2 IBIAS2.t78 VDD.t524 VDD.t336 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X456 VDD.t1313 VDD.t1312 VDD.t1313 VDD.t1188 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X457 VDD IBIAS2.t266 OUT_N.t179 VDD.t669 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X458 VDD.t1311 VDD.t1310 VDD.t1311 VDD.t1237 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X459 VDD IBIAS3.t44 IVS.t35 VDD.t204 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X460 VPD VB1.t41 VDD.t1140 VDD.t759 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X461 VDD IBIAS2.t267 OUT_N.t178 VDD.t119 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X462 OUT_N IBIAS2.t268 VDD.t674 VDD.t117 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X463 VDD IBIAS2.t269 OUT_P.t158 VDD.t494 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X464 OUT_P IBIAS2.t270 VDD.t1047 VDD.t454 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X465 VSS VB4.t64 IND.t35 VSS.t175 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X466 VSS.t525 VSS.t524 VSS.t525 VSS.t419 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X467 VSS.t523 VSS.t521 VSS.t523 VSS.t522 nfet_03v3 ad=0.26p pd=1.52u as=0 ps=0 w=1u l=0.28u
X468 IB2 VB2.t28 VB2.t29 VDD.t1095 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X469 VDD.t1309 VDD.t1308 VDD.t1309 VDD.t1261 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X470 OUT_N OUT1.t57 VSS.t111 VSS.t101 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X471 VDD IBIAS3.t45 IVS.t34 VDD.t204 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X472 VBM VCM.t7 VCD.t35 VSS.t352 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X473 VSS OUT2.t62 OUT_P.t22 VSS.t98 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X474 OUT1 VB2.t49 VND.t9 VDD.t103 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X475 OUT2 VB2.t50 VPD.t27 VDD.t305 pfet_03v3 ad=1.38p pd=7.14u as=1.38p ps=7.14u w=3.13u l=0.28u
X476 VSS.t520 VSS.t519 VSS.t520 VSS.t477 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.28u
X477 VSS VB4.t65 IND.t34 VSS.t221 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X478 VPD VB1.t42 VDD.t782 VDD.t759 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X479 VDD IBIAS2.t271 OUT_N.t176 VDD.t60 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X480 OUT_P IBIAS2.t272 VDD.t601 VDD.t389 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X481 VDD IBIAS.t8 IBIAS.t9 VDD.t1066 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X482 VSS OUT2.t63 OUT_P.t265 VSS.t19 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X483 VDD.t1307 VDD.t1306 VDD.t1307 VDD.t1237 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X484 VDD IBIAS2.t273 OUT_N.t175 VDD.t32 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X485 VND VB1.t43 VDD.t538 VDD.t105 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X486 OUT_P IBIAS2.t274 VDD.t604 VDD.t163 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X487 VDD IBIAS2.t76 IBIAS2.t77 VDD.t515 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X488 VSS IBS.t2 IBS.t3 VSS.t607 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=1u
X489 OUT_P OUT2.t64 VSS.t652 VSS.t103 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X490 OUT_N IBIAS2.t275 VDD.t698 VDD.t301 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X491 VSS.t518 VSS.t517 VSS.t518 VSS.t46 nfet_03v3 ad=0.88p pd=4.88u as=0 ps=0 w=2u l=1u
X492 IB3 VB3.t2 VB3.t3 VSS.t398 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X493 VDD.t1305 VDD.t1304 VDD.t1305 VDD.t1194 pfet_03v3 ad=1.65p pd=8.38u as=0 ps=0 w=3.75u l=0.28u
X494 IPD IN_P.t9 BD.t60 VDD.t620 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X495 VDD IBIAS2.t276 OUT_N.t173 VDD.t77 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X496 VSS OUT1.t58 OUT_N.t12 VSS.t16 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X497 VDD IBIAS2.t74 IBIAS2.t75 VDD.t7 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X498 VDD IBIAS2.t277 OUT_P.t154 VDD.t127 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X499 VBIASN VBIASN.t3 VSS.t658 VSS.t657 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X500 BD IN_N.t8 IND.t49 VDD.t107 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X501 IND VB4.t66 VSS.t237 VSS.t209 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X502 OUT1 VB2.t51 VND.t8 VDD.t304 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X503 VB2 VB2.t10 IB2.t11 VDD.t1101 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X504 VDD IBIAS2.t278 OUT_N.t172 VDD.t241 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X505 VDD IBIAS2.t279 OUT_P.t153 VDD.t244 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X506 VDD IBIAS2.t280 OUT_N.t171 VDD.t236 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X507 VB4 VB4.t4 VSS.t236 VSS.t235 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X508 VSS.t516 VSS.t515 VSS.t516 VSS.t493 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.28u
X509 VSS VB4.t68 IND.t33 VSS.t175 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X510 VDD.t1303 VDD.t1301 VDD.t1303 VDD.t1302 pfet_03v3 ad=1.04p pd=4.52u as=0 ps=0 w=4u l=0.28u
X511 OUT2 VB2.t53 VPD.t28 VDD.t304 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X512 OUT_N IBIAS2.t281 VDD.t1041 VDD.t72 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X513 OUT_N IBIAS2.t282 VDD.t1042 VDD.t50 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X514 VSS IVS.t66 IVS.t67 VSS.t620 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X515 VSS OUT1.t59 OUT_N.t13 VSS.t28 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X516 VDD IBIAS2.t283 OUT_P.t152 VDD.t216 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X517 OUT_N IBIAS2.t284 VDD.t543 VDD.t435 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X518 IND IN_N.t9 BD.t49 VDD.t411 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X519 IPD VB4.t69 VSS.t232 VSS.t197 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X520 VSS.t514 VSS.t513 VSS.t514 VSS.t401 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X521 OUT_P IBIAS2.t285 VDD.t544 VDD.t150 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X522 VCD VOUT.t14 VB1.t32 VSS.t4 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X523 OUT_N OUT1.t60 VSS.t69 VSS.t68 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X524 VDD IBIAS2.t286 OUT_N.t167 VDD.t38 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X525 VDD.t397 VDD.t398 VDD.t396 ppolyf_u r_width=1u r_length=5u
X526 VSS OUT2.t65 OUT_P.t267 VSS.t33 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X527 VSS OUT2.t66 OUT_P.t268 VSS.t28 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X528 VDD IBIAS2.t287 OUT_P.t150 VDD.t224 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X529 OUT1 VB2.t54 VND.t7 VDD.t102 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X530 VDD IBIAS1.t7 VB3.t15 VDD.t192 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X531 OUT_P OUT2.t67 VSS.t325 VSS.t313 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X532 VDD IBIAS2.t288 OUT_N.t166 VDD.t0 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X533 VDD.t1300 VDD.t1299 VDD.t1300 VDD.t1242 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X534 VDD.t935 VDD.t936 VDD.t934 ppolyf_u r_width=1u r_length=6.2u
X535 VDD IBIAS2.t289 OUT_P.t149 VDD.t216 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X536 VSS.t512 VSS.t511 VSS.t512 VSS.t433 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X537 OUT_N IBIAS2.t290 VDD.t725 VDD.t256 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X538 IB2 VB2.t26 VB2.t27 VDD.t652 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X539 VDD IBIAS.t23 BD.t66 VDD.t134 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X540 VDD IBIAS2.t291 OUT_N.t164 VDD.t74 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X541 VDD IBIAS2.t292 OUT_P.t148 VDD.t176 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X542 VDD IBIAS4.t8 IB4.t14 VDD.t1013 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X543 IPD VB3.t32 OUT2.t34 VSS.t388 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X544 VDD VB1.t44 VPD.t10 VDD.t209 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X545 VSS VB4.t22 VB4.t23 VSS.t229 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X546 VDD IBIAS2.t293 OUT_P.t147 VDD.t54 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X547 VDD IBIAS2.t294 OUT_P.t146 VDD.t236 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X548 VDD IBIAS2.t295 OUT_P.t145 VDD.t43 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X549 VDD IBIAS.t24 BD.t2 VDD.t134 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X550 VSS.t510 VSS.t509 VSS.t510 VSS.t407 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X551 OUT_N OUT1.t61 VSS.t70 VSS.t38 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X552 VDD IBIAS2.t296 OUT_N.t163 VDD.t158 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X553 VDD IBIAS2.t297 OUT_P.t144 VDD.t624 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X554 VDD IBIAS2.t298 OUT_P.t143 VDD.t577 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X555 OUT_P IBIAS2.t299 VDD.t596 VDD.t214 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X556 OUT_P IBIAS2.t300 VDD.t598 VDD.t597 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X557 VSS.t508 VSS.t507 VSS.t508 VSS.t456 nfet_03v3 ad=0.88p pd=4.88u as=0 ps=0 w=2u l=1u
X558 VDD VB1.t45 VND.t28 VDD.t285 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X559 VDD IBIAS2.t301 OUT_N.t162 VDD.t317 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X560 VDD IBIAS2.t302 OUT_P.t140 VDD.t67 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X561 OUT_N IBIAS2.t303 VDD.t859 VDD.t117 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X562 OUT_N IBIAS2.t304 VDD.t860 VDD.t41 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X563 VDD IBIAS3.t46 IVS.t33 VDD.t401 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X564 VDD IBIAS3.t47 IVS.t32 VDD.t167 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X565 IBIAS2 IBIAS2.t72 VDD.t1400 VDD.t195 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X566 VSS IVS.t82 IBIAS2.t116 VSS.t346 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X567 OUT_N IBIAS2.t306 VDD.t951 VDD.t94 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X568 a_25526_n6312# a_24350_n7414# VDD.t183 ppolyf_u r_width=1u r_length=5u
X569 VDD.t1298 VDD.t1297 VDD.t1298 VDD.t1247 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X570 IBIAS2 IBIAS2.t70 VDD.t1399 VDD.t195 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X571 IB3 VB3.t33 VSS.t387 VSS.t386 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X572 OUT_N OUT1.t62 VSS.t72 VSS.t71 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X573 OUT_P IBIAS2.t308 VDD.t952 VDD.t645 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X574 IBIAS2 IBIAS2.t68 VDD.t1405 VDD.t140 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X575 VDD.t1296 VDD.t1295 VDD.t1296 VDD.t1185 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X576 VND VB1.t46 VDD.t771 VDD.t770 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X577 VSS OUT2.t68 OUT_P.t233 VSS.t114 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X578 OUT_P IBIAS2.t310 VDD.t953 VDD.t150 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X579 VND VB1.t47 VDD.t969 VDD.t759 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X580 VSS.t506 VSS.t505 VSS.t506 VSS.t477 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.28u
X581 VSS OUT1.t63 OUT_N.t17 VSS.t28 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X582 VDD.t1294 VDD.t1293 VDD.t1294 VDD.t1261 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X583 OUT2 VB2.t55 VPD.t0 VDD.t103 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X584 OUT_N OUT1.t64 VSS.t360 VSS.t103 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X585 OUT_P OUT2.t69 VSS.t328 VSS.t112 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X586 VDD.t1292 VDD.t1290 VDD.t1292 VDD.t1291 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X587 VSS OUT1.t65 OUT_N.t248 VSS.t19 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X588 VDD IBIAS2.t311 OUT_P.t137 VDD.t494 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X589 OUT_P IBIAS2.t312 VDD.t710 VDD.t435 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X590 VSS.t504 VSS.t503 VSS.t504 VSS.t401 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X591 OUT_N IBIAS2.t313 VDD.t711 VDD.t125 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X592 VPD VB1.t48 VDD.t133 VDD.t105 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X593 VDD.t1289 VDD.t1288 VDD.t1289 VDD.t1188 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X594 OUT_P IBIAS2.t314 VDD.t637 VDD.t374 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X595 VDD.t1287 VDD.t1286 VDD.t1287 VDD.t1166 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X596 VDD IBIAS.t25 BD.t3 VDD.t137 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X597 IVS IBIAS3.t48 VDD.t534 VDD.t109 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X598 OUT_P OUT2.t70 VSS.t329 VSS.t83 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X599 OUT_N OUT1.t66 VSS.t363 VSS.t38 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X600 VND VB2.t56 OUT1.t2 VDD.t104 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X601 VDD IBIAS2.t315 OUT_N.t157 VDD.t508 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X602 VDD.t1285 VDD.t1283 VDD.t1285 VDD.t1284 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X603 VDD IBIAS2.t316 OUT_P.t134 VDD.t46 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X604 VSS VB4.t20 VB4.t21 VSS.t226 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X605 VDD IBIAS.t26 BD.t11 VDD.t134 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X606 VDD IBIAS2.t317 OUT_N.t156 VDD.t666 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X607 VDD IBIAS2.t66 IBIAS2.t67 VDD.t1107 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X608 VDD IBIAS2.t318 OUT_N.t155 VDD.t483 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X609 BD IN_N.t10 IND.t50 VDD.t530 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X610 OUT_P OUT2.t71 VSS.t601 VSS.t71 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X611 OUT_P IBIAS2.t319 VDD.t707 VDD.t63 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X612 IND IN_N.t11 BD.t47 VDD.t230 pfet_03v3 ad=1.65p pd=8.38u as=0.975p ps=4.27u w=3.75u l=0.28u
X613 VSS OUT2.t72 OUT_P.t261 VSS.t7 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X614 VDD.t1282 VDD.t1281 VDD.t1282 VDD.t1156 pfet_03v3 ad=1.65p pd=8.38u as=0 ps=0 w=3.75u l=0.28u
X615 VDD.t1280 VDD.t1278 VDD.t1280 VDD.t1279 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X616 VBM VCM.t8 VCD.t34 VSS.t142 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X617 VDD IBIAS2.t320 OUT_N.t154 VDD.t314 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X618 IBIAS2 IBIAS2.t64 VDD.t1409 VDD.t526 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X619 BD IBIAS.t27 VDD.t395 VDD.t329 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X620 OUT2 VB3.t34 IPD.t38 VSS.t384 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X621 OUT_P OUT2.t73 VSS.t604 VSS.t91 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X622 VDD IBIAS2.t62 IBIAS2.t63 VDD.t1107 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X623 VDD.t419 VDD.t420 VDD.t10 ppolyf_u r_width=1u r_length=6.2u
X624 OUT_N OUT1.t67 VSS.t364 VSS.t101 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X625 OUT_N IBIAS2.t322 VDD.t1038 VDD.t645 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X626 VDD.t1277 VDD.t1276 VDD.t1277 VDD.t1250 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X627 VDD IBIAS2.t323 OUT_P.t132 VDD.t60 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X628 VB1 VOUT.t15 VCD.t61 VSS.t352 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X629 OUT_N IBIAS2.t324 VDD.t1009 VDD.t645 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X630 VSS OUT1.t68 OUT_N.t251 VSS.t24 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X631 IB4 IB4.t6 VSS.t670 VSS.t636 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X632 VSS VB4.t70 IND.t32 VSS.t175 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X633 VSS VB4.t71 IPD.t18 VSS.t221 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X634 OUT_N IBIAS2.t325 VDD.t1010 VDD.t161 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X635 a_24070_n6312# OUT_N.t244 VDD.t415 ppolyf_u r_width=1u r_length=5u
X636 a_29248_n7510.t4 OUT_N.t254 cap_mim_2f0fF c_width=21u c_length=21u
X637 VDD IBIAS3.t49 IVS.t30 VDD.t167 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X638 VSS.t502 VSS.t501 VSS.t502 VSS.t477 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.28u
X639 VDD IBIAS.t28 BD.t69 VDD.t137 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X640 VSS.t500 VSS.t499 VSS.t500 VSS.t413 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X641 VDD IBIAS.t29 BD.t70 VDD.t137 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X642 VND VB1.t49 VDD.t106 VDD.t105 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X643 VSS OUT2.t74 OUT_P.t263 VSS.t13 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X644 IBIAS3 IBIAS3.t11 VDD.t593 VDD.t574 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X645 OUT2 VB2.t57 VPD.t17 VDD.t304 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X646 VDD IBIAS2.t326 OUT_N.t150 VDD.t152 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X647 BD IBIAS.t30 VDD.t655 VDD.t522 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X648 OUT_P OUT2.t75 VSS.t143 VSS.t79 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X649 VDD IBIAS2.t327 OUT_P.t131 VDD.t469 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X650 VDD IBIAS3.t51 IVS.t29 VDD.t167 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X651 VSS VB4.t72 IND.t31 VSS.t192 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X652 OUT_N OUT1.t69 VSS.t367 VSS.t83 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X653 OUT_N IBIAS2.t328 VDD.t997 VDD.t21 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X654 VDD IBIAS2.t329 OUT_P.t130 VDD.t77 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X655 OUT_N IBIAS2.t330 VDD.t836 VDD.t430 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X656 VDD IBIAS2.t331 OUT_N.t147 VDD.t666 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X657 VDD IBIAS2.t332 OUT_P.t129 VDD.t311 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X658 VDD IBIAS1.t8 IBS.t6 VDD.t753 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X659 VDD IBIAS2.t333 OUT_N.t146 VDD.t624 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X660 OUT2.t26 a_29248_n5498.t2 VDD.t116 ppolyf_u r_width=1u r_length=6.2u
X661 BD IBIAS.t31 VDD.t656 VDD.t114 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X662 VDD IBIAS2.t334 OUT_N.t145 VDD.t216 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X663 IVS IBIAS3.t52 VDD.t514 VDD.t364 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X664 VDD IBIAS2.t335 OUT_N.t144 VDD.t812 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X665 VDD IBIAS2.t60 IBIAS2.t61 VDD.t145 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X666 IND IN_N.t12 BD.t46 VDD.t620 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X667 VND VB1.t50 VDD.t760 VDD.t759 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X668 OUT_N IBIAS2.t336 VDD.t634 VDD.t430 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X669 VSS.t498 VSS.t497 VSS.t498 VSS.t425 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X670 VSS.t496 VSS.t495 VSS.t496 VSS.t401 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X671 VSS.t494 VSS.t492 VSS.t494 VSS.t493 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.28u
X672 VCD VCM.t9 VBM.t21 VSS.t4 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X673 VSS OUT1.t70 OUT_N.t36 VSS.t7 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X674 IBIAS2 IBIAS2.t58 VDD.t797 VDD.t202 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X675 VB2 VB2.t8 IB2.t9 VDD.t740 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X676 VDD.t367 VDD.t368 VDD.t14 ppolyf_u r_width=1u r_length=5u
X677 VCD VOUT.t16 VB1.t20 VSS.t6 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X678 IND VB3.t35 OUT1.t13 VSS.t388 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X679 OUT_N IBIAS2.t338 VDD.t635 VDD.t256 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X680 VDD IBIAS.t6 IBIAS.t7 VDD.t189 pfet_03v3 ad=1.04p pd=4.52u as=1.76p ps=8.88u w=4u l=0.56u
X681 VSS.t491 VSS.t490 VSS.t491 VSS.t410 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X682 VSS VB4.t73 IND.t30 VSS.t159 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X683 VSS.t489 VSS.t488 VSS.t489 VSS.t419 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X684 VDD.t1275 VDD.t1274 VDD.t1275 VDD.t1209 pfet_03v3 ad=1.65p pd=8.38u as=0 ps=0 w=3.75u l=0.28u
X685 VDD VB1.t51 VPD.t8 VDD.t761 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X686 VSS OUT2.t76 OUT_P.t24 VSS.t98 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X687 OUT_P OUT2.t77 VSS.t146 VSS.t89 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X688 VDD IBIAS2.t56 IBIAS2.t57 VDD.t145 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X689 BD IN_N.t13 IND.t66 VDD.t418 pfet_03v3 ad=0.975p pd=4.27u as=1.65p ps=8.38u w=3.75u l=0.28u
X690 IPD VB4.t74 VSS.t216 VSS.t209 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X691 OUT_N IBIAS2.t339 VDD.t636 VDD.t254 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X692 VSS.t487 VSS.t486 VSS.t487 VSS.t442 nfet_03v3 ad=0.52p pd=2.52u as=0 ps=0 w=2u l=1u
X693 VDD IBIAS2.t340 OUT_P.t128 VDD.t46 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X694 OUT_P IBIAS2.t341 VDD.t1123 VDD.t492 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X695 IBIAS3 IB4.t21 VSS.t343 VSS.t342 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X696 IBIAS2 IBIAS2.t54 VDD.t144 VDD.t142 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X697 VSS OUT2.t78 OUT_P.t26 VSS.t40 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X698 VDD IBIAS3.t53 IVS.t27 VDD.t331 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X699 VCD VBIASN.t10 VSS.t52 VSS.t51 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X700 BD IN_P.t10 IPD.t64 VDD.t292 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X701 OUT_N IBIAS2.t343 VDD.t1124 VDD.t379 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X702 IBIAS2 IBIAS2.t52 VDD.t427 VDD.t140 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X703 VSS OUT1.t71 OUT_N.t37 VSS.t16 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X704 OUT_P IBIAS2.t345 VDD.t642 VDD.t492 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X705 VB3 IBIAS1.t9 VDD.t971 VDD.t970 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X706 IPD VB4.t75 VSS.t215 VSS.t197 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X707 IND VB4.t76 VSS.t214 VSS.t197 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X708 OUT_N OUT1.t72 VSS.t153 VSS.t83 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X709 VDD.t11 VDD.t12 VDD.t10 ppolyf_u r_width=1u r_length=6.2u
X710 OUT_P OUT2.t79 VSS.t39 VSS.t38 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X711 OUT_N IBIAS2.t346 VDD.t643 VDD.t17 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X712 VSS VB4.t18 VB4.t19 VSS.t211 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X713 IND IN_N.t14 BD.t44 VDD.t294 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X714 IPD VB3.t36 OUT2.t22 VSS.t2 nfet_03v3 ad=1.27p pd=6.64u as=1.27p ps=6.64u w=2.88u l=0.28u
X715 OUT_P IBIAS2.t347 VDD.t644 VDD.t50 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X716 VDD IBIAS2.t348 OUT_P.t124 VDD.t179 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X717 OUT_N IBIAS2.t349 VDD.t607 VDD.t263 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X718 VDD.t1273 VDD.t1272 VDD.t1273 VDD.t1242 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X719 VDD IBIAS2.t350 OUT_N.t137 VDD.t176 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X720 VSS.t485 VSS.t484 VSS.t485 VSS.t430 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X721 VDD.t1271 VDD.t1269 VDD.t1271 VDD.t1270 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X722 a_25078_n6312# a_26254_n7414# VDD.t13 ppolyf_u r_width=1u r_length=5u
X723 VB1 VOUT.t17 VCD.t43 VSS.t353 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X724 VDD.t1268 VDD.t1267 VDD.t1268 VDD.t1156 pfet_03v3 ad=1.65p pd=8.38u as=0 ps=0 w=3.75u l=0.28u
X725 VDD.t1266 VDD.t1265 VDD.t1266 VDD.t1166 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X726 OUT_P IBIAS2.t351 VDD.t954 VDD.t70 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X727 BD IBIAS.t32 VDD.t972 VDD.t114 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X728 IND VB4.t77 VSS.t210 VSS.t209 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X729 VSS OUT2.t80 OUT_P.t1 VSS.t40 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X730 OUT_P OUT2.t81 VSS.t43 VSS.t22 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X731 OUT_N IBIAS2.t352 VDD.t955 VDD.t301 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X732 OUT_P IBIAS2.t353 VDD.t956 VDD.t358 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X733 VSS IBS.t10 IBIAS.t1 VSS.t610 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=1u
X734 VDD IBIAS1.t10 IB5.t1 VDD.t1134 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X735 VSS VB4.t78 IPD.t15 VSS.t175 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X736 VDD IBIAS2.t354 OUT_P.t121 VDD.t0 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X737 OUT_N IBIAS2.t355 VDD.t4 VDD.t3 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X738 OUT1.t4 a_29248_n7510.t0 VDD.t116 ppolyf_u r_width=1u r_length=6.2u
X739 VDD.t1264 VDD.t1263 VDD.t1264 VDD.t1228 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X740 OUT_P IBIAS2.t356 VDD.t6 VDD.t5 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X741 VB2 VB2.t6 IB2.t8 VDD.t212 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X742 IBIAS2 IBIAS2.t50 VDD.t426 VDD.t171 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X743 VSS.t483 VSS.t481 VSS.t483 VSS.t482 nfet_03v3 ad=0.26p pd=1.52u as=0 ps=0 w=1u l=0.28u
X744 VCD VOUT.t18 VB1.t14 VSS.t141 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X745 VB4 VB4.t2 VSS.t206 VSS.t205 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X746 OUT2 VB3.t37 IPD.t69 VSS.t391 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X747 VDD IBIAS.t33 BD.t68 VDD.t267 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X748 VDD VB1.t52 VND.t23 VDD.t282 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X749 VDD IBIAS2.t358 OUT_P.t119 VDD.t669 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X750 VSS IB4.t4 IB4.t5 VSS.t624 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X751 OUT1 VB2.t60 VND.t5 VDD.t304 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X752 VDD IBIAS2.t359 OUT_N.t134 VDD.t119 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X753 IBIAS2 IBIAS2.t48 VDD.t425 VDD.t195 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X754 a_23622_n6312# OUT_P.t231 VDD.t405 ppolyf_u r_width=1u r_length=5u
X755 IBIAS3 IB4.t22 VSS.t345 VSS.t344 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X756 VSS OUT1.t73 OUT_N.t39 VSS.t13 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X757 OUT_N IBIAS2.t361 VDD.t724 VDD.t567 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X758 BD IN_N.t15 IND.t47 VDD.t418 pfet_03v3 ad=0.975p pd=4.27u as=1.65p ps=8.38u w=3.75u l=0.28u
X759 VDD IBIAS2.t362 OUT_N.t132 VDD.t91 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X760 VDD IBIAS2.t46 IBIAS2.t47 VDD.t145 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X761 IBIAS IBIAS.t4 VDD.t1070 VDD.t1069 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X762 OUT2 VB2.t61 VPD.t18 VDD.t305 pfet_03v3 ad=1.38p pd=7.14u as=1.38p ps=7.14u w=3.13u l=0.28u
X763 VDD.t1262 VDD.t1260 VDD.t1262 VDD.t1261 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X764 VDD.t1259 VDD.t1258 VDD.t1259 VDD.t1201 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X765 OUT_N IBIAS2.t363 VDD.t718 VDD.t3 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X766 OUT_P IBIAS2.t364 VDD.t719 VDD.t81 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X767 IB4 IBIAS4.t9 VDD.t1016 VDD.t895 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X768 VDD.t1257 VDD.t1256 VDD.t1257 VDD.t1237 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X769 VDD IBIAS2.t365 OUT_N.t130 VDD.t127 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X770 OUT_P IBIAS2.t366 VDD.t375 VDD.t374 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X771 OUT1 VB3.t38 IND.t63 VSS.t384 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X772 VDD IBIAS2.t367 OUT_N.t129 VDD.t376 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X773 OUT_P IBIAS2.t368 VDD.t441 VDD.t301 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X774 VDD IBIAS3.t54 IVS.t26 VDD.t331 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X775 VSS VBIASN.t11 VCD.t4 VSS.t53 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X776 VDD.t1255 VDD.t1254 VDD.t1255 VDD.t1179 pfet_03v3 ad=1.65p pd=8.38u as=0 ps=0 w=3.75u l=0.28u
X777 OUT_N OUT1.t74 VSS.t156 VSS.t112 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X778 IVS IVS.t64 VSS.t619 VSS.t618 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X779 VSS OUT1.t75 OUT_N.t41 VSS.t40 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X780 IB2 VB2.t24 VB2.t25 VDD.t623 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X781 VSS.t480 VSS.t479 VSS.t480 VSS.t425 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X782 VDD IBIAS2.t44 IBIAS2.t45 VDD.t173 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X783 VDD IBIAS2.t369 OUT_P.t115 VDD.t442 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X784 VB1 VOUT.t19 VCD.t60 VSS.t140 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X785 IND VB3.t39 OUT1.t21 VSS.t388 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X786 VDD IBIAS2.t370 OUT_N.t128 VDD.t445 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X787 VDD IBIAS2.t371 OUT_P.t114 VDD.t624 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X788 a_24350_n4340# a_25526_n5442# VDD.t183 ppolyf_u r_width=1u r_length=5u
X789 VDD IBIAS3.t55 IVS.t25 VDD.t331 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X790 VSS IVS.t84 IBIAS2.t117 VSS.t339 nfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=1u
X791 OUT2 VB3.t40 IPD.t57 VSS.t392 nfet_03v3 ad=1.27p pd=6.64u as=1.27p ps=6.64u w=2.88u l=0.28u
X792 VSS OUT1.t76 OUT_N.t265 VSS.t28 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X793 VDD.t1253 VDD.t1252 VDD.t1253 VDD.t843 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X794 IND IN_N.t16 BD.t42 VDD.t108 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X795 VDD IBIAS2.t372 OUT_N.t127 VDD.t244 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X796 VDD IBIAS2.t373 OUT_P.t113 VDD.t236 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X797 VDD.t1251 VDD.t1249 VDD.t1251 VDD.t1250 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X798 VBM VCM.t10 VCD.t32 VSS.t352 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X799 VDD IBIAS2.t374 OUT_P.t112 VDD.t314 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X800 VSS OUT2.t82 OUT_P.t3 VSS.t19 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X801 OUT_N IBIAS2.t375 VDD.t714 VDD.t358 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X802 IBIAS2 IBIAS2.t42 VDD.t1116 VDD.t202 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X803 OUT_N IBIAS2.t377 VDD.t715 VDD.t96 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X804 IVS IVS.t62 VSS.t617 VSS.t62 nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=1u
X805 BD IN_P.t11 IPD.t33 VDD.t166 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X806 IND IN_N.t17 BD.t41 VDD.t294 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X807 OUT_P IBIAS2.t378 VDD.t436 VDD.t435 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X808 a_29248_n5498.t1 OUT_P.t269 cap_mim_2f0fF c_width=21u c_length=21u
X809 IPD IN_P.t12 BD.t16 VDD.t353 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X810 OUT_N IBIAS2.t379 VDD.t438 VDD.t437 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X811 VSS IVS.t86 IBIAS2.t118 VSS.t349 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X812 VB2 VB2.t4 IB2.t6 VDD.t591 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X813 VSS.t478 VSS.t476 VSS.t478 VSS.t477 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.28u
X814 VDD IBIAS2.t380 OUT_N.t123 VDD.t57 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X815 VDD IBIAS2.t381 OUT_P.t110 VDD.t221 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X816 VB4 VB4.t0 VSS.t204 VSS.t203 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X817 VSS OUT2.t83 OUT_P.t248 VSS.t98 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X818 VPD VB2.t63 OUT2.t5 VDD.t309 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X819 VSS OUT2.t84 OUT_P.t249 VSS.t114 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X820 VDD IBIAS2.t382 OUT_N.t122 VDD.t224 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X821 VDD.t1248 VDD.t1246 VDD.t1248 VDD.t1247 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X822 VDD.t1245 VDD.t1244 VDD.t1245 VDD.t1191 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X823 VDD.t1243 VDD.t1241 VDD.t1243 VDD.t1242 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X824 OUT_P IBIAS2.t383 VDD.t228 VDD.t227 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X825 VSS.t475 VSS.t474 VSS.t475 VSS.t419 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X826 OUT_P IBIAS2.t384 VDD.t215 VDD.t214 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X827 VSS.t473 VSS.t472 VSS.t473 VSS.t401 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X828 VDD IBIAS2.t385 OUT_N.t121 VDD.t216 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X829 VDD IBIAS2.t386 OUT_P.t107 VDD.t158 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X830 IVS IBIAS3.t56 VDD.t334 VDD.t207 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X831 VDD.t1240 VDD.t1239 VDD.t1240 VDD.t1142 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X832 OUT_P IBIAS2.t387 VDD.t257 VDD.t256 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X833 IVS IBIAS3.t57 VDD.t943 VDD.t306 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X834 OUT_N OUT1.t77 VSS.t674 VSS.t68 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X835 VDD IBIAS2.t388 OUT_P.t105 VDD.t74 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X836 BD IBIAS.t35 VDD.t1137 VDD.t329 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X837 VCD VCM.t11 VBM.t20 VSS.t6 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X838 VCD VOUT.t20 VB1.t19 VSS.t4 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X839 OUT_P IBIAS2.t389 VDD.t253 VDD.t252 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X840 VSS.t471 VSS.t470 VSS.t471 VSS.t430 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X841 OUT_N IBIAS2.t390 VDD.t255 VDD.t254 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X842 VDD.t1238 VDD.t1236 VDD.t1238 VDD.t1237 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X843 a_25526_n6312# a_25806_n7414# VDD.t366 ppolyf_u r_width=1u r_length=5u
X844 VDD.t1235 VDD.t1234 VDD.t1235 VDD.t1212 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.28u
X845 VDD.t1233 VDD.t1232 VDD.t1233 VDD.t1191 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X846 VDD.t1231 VDD.t1230 VDD.t1231 VDD.t1153 pfet_03v3 ad=0.814p pd=3.65u as=0 ps=0 w=3.13u l=0.56u
X847 VDD VB1.t53 VND.t22 VDD.t282 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X848 VDD IBIAS2.t391 OUT_P.t103 VDD.t158 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X849 OUT_N IBIAS2.t392 VDD.t251 VDD.t227 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X850 IND VB4.t81 VSS.t202 VSS.t162 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X851 VDD.t1229 VDD.t1227 VDD.t1229 VDD.t1228 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X852 OUT_N IBIAS2.t393 VDD.t871 VDD.t597 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X853 OUT_P OUT2.t85 VSS.t378 VSS.t313 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X854 IB4 IBIAS4.t10 VDD.t1017 VDD.t895 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X855 IB2 VB2.t22 VB2.t23 VDD.t749 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X856 OUT_P OUT2.t86 VSS.t379 VSS.t103 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X857 IPD IN_P.t13 BD.t17 VDD.t411 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X858 OUT_N IBIAS2.t394 VDD.t872 VDD.t81 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X859 OUT1 VB2.t64 VND.t4 VDD.t305 pfet_03v3 ad=1.38p pd=7.14u as=1.38p ps=7.14u w=3.13u l=0.28u
X860 BD IN_N.t18 IND.t3 VDD.t107 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X861 VDD VB1.t54 VPD.t7 VDD.t285 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X862 VDD IBIAS2.t395 OUT_P.t102 VDD.t122 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X863 IB4 IBIAS4.t11 VDD.t896 VDD.t895 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X864 VDD IBIAS1.t11 IBS.t8 VDD.t772 pfet_03v3 ad=1.04p pd=4.52u as=1.76p ps=8.88u w=4u l=0.56u
X865 OUT_N OUT1.t78 VSS.t675 VSS.t313 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X866 OUT_P IBIAS2.t396 VDD.t233 VDD.t21 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X867 VDD IBIAS2.t40 IBIAS2.t41 VDD.t7 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X868 OUT_N IBIAS2.t397 VDD.t883 VDD.t551 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X869 VDD IBIAS2.t38 IBIAS2.t39 VDD.t23 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X870 OUT_P IBIAS2.t398 VDD.t884 VDD.t256 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X871 VDD.t1226 VDD.t1225 VDD.t1226 VDD.t1185 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X872 VOUT.t1 a_24070_n5442# VDD.t415 ppolyf_u r_width=1u r_length=5u
X873 OUT_N OUT1.t79 VSS.t676 VSS.t83 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X874 VSS.t469 VSS.t468 VSS.t469 VSS.t407 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X875 OUT_N IBIAS2.t399 VDD.t868 VDD.t150 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X876 VND VB2.t65 OUT1.t7 VDD.t310 pfet_03v3 ad=1.38p pd=7.14u as=1.38p ps=7.14u w=3.13u l=0.28u
X877 VDD IBIAS2.t400 OUT_P.t99 VDD.t445 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X878 OUT_P IBIAS2.t401 VDD.t913 VDD.t587 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X879 VDD IBIAS3.t58 IVS.t22 VDD.t204 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X880 VSS VB4.t82 IPD.t14 VSS.t175 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X881 IPD VB3.t41 OUT2.t21 VSS.t2 nfet_03v3 ad=1.27p pd=6.64u as=1.27p ps=6.64u w=2.88u l=0.28u
X882 VDD IBIAS3.t59 IVS.t21 VDD.t406 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X883 VDD.t1224 VDD.t1223 VDD.t1224 VDD.t843 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X884 OUT_P IBIAS2.t402 VDD.t914 VDD.t389 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X885 VBM VCM.t12 VCD.t30 VSS.t353 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X886 IND VB4.t83 VSS.t199 VSS.t162 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X887 VDD IBIAS2.t403 OUT_N.t114 VDD.t494 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X888 OUT_N IBIAS2.t404 VDD.t867 VDD.t161 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X889 VDD IBIAS.t36 BD.t79 VDD.t267 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X890 OUT_P IBIAS2.t405 VDD.t983 VDD.t125 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X891 VDD.t1222 VDD.t1221 VDD.t1222 VDD.t1166 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X892 VSS OUT2.t87 OUT_P.t240 VSS.t33 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X893 OUT_N OUT1.t80 VSS.t677 VSS.t71 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X894 VDD IBIAS4.t3 IBIAS4.t4 VDD.t843 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X895 VDD IBIAS2.t36 IBIAS2.t37 VDD.t23 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X896 BD IN_P.t14 IPD.t45 VDD.t361 pfet_03v3 ad=0.975p pd=4.27u as=1.65p ps=8.38u w=3.75u l=0.28u
X897 OUT_P OUT2.t88 VSS.t356 VSS.t71 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X898 VDD IBIAS3.t60 IVS.t20 VDD.t412 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X899 VB3 VB3.t6 IB3.t2 VSS.t683 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X900 VDD.t1220 VDD.t1219 VDD.t1220 VDD.t1148 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X901 IPD VB4.t84 VSS.t198 VSS.t197 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X902 VSS OUT2.t89 OUT_P.t242 VSS.t93 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X903 VSS.t467 VSS.t466 VSS.t467 VSS.t453 nfet_03v3 ad=0.26p pd=1.52u as=0 ps=0 w=1u l=0.28u
X904 VDD VBM.t2 VBM.t3 VDD.t1092 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X905 VSS VB4.t85 IPD.t12 VSS.t159 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X906 VDD IBIAS2.t406 OUT_P.t95 VDD.t508 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X907 VDD.t1218 VDD.t1217 VDD.t1218 VDD.t1201 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X908 IND VB3.t43 OUT1.t18 VSS.t1 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X909 VB1 VOUT.t21 VCD.t51 VSS.t352 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X910 OUT_P OUT2.t90 VSS.t359 VSS.t89 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X911 OUT_P OUT2.t91 VSS.t124 VSS.t112 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X912 VDD IBIAS2.t407 OUT_P.t94 VDD.t457 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X913 OUT_N IBIAS2.t408 VDD.t982 VDD.t214 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X914 VSS.t465 VSS.t464 VSS.t465 VSS.t46 nfet_03v3 ad=0.88p pd=4.88u as=0 ps=0 w=2u l=1u
X915 VDD.t1216 VDD.t1214 VDD.t1216 VDD.t1215 pfet_03v3 ad=1.04p pd=4.52u as=0 ps=0 w=4u l=0.28u
X916 OUT_P IBIAS2.t409 VDD.t149 VDD.t148 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X917 OUT_N IBIAS2.t410 VDD.t151 VDD.t150 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X918 VCD VCM.t13 VBM.t19 VSS.t141 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X919 OUT_N IBIAS2.t411 VDD.t562 VDD.t261 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X920 VSS VBIASN.t12 VB2.t32 VSS.t56 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X921 VSS OUT1.t81 OUT_N.t270 VSS.t10 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X922 OUT_N IBIAS2.t412 VDD.t563 VDD.t63 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X923 VDD IBIAS2.t413 OUT_N.t108 VDD.t244 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X924 VDD IBIAS2.t34 IBIAS2.t35 VDD.t23 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X925 OUT_P IBIAS2.t414 VDD.t586 VDD.t437 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X926 VDD IBIAS2.t415 OUT_N.t107 VDD.t508 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X927 IVS IBIAS3.t61 VDD.t307 VDD.t306 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X928 a_24070_n6312# a_24350_n7414# VDD.t35 ppolyf_u r_width=1u r_length=5u
X929 VSS.t463 VSS.t462 VSS.t463 VSS.t404 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X930 VDD VB1.t55 VPD.t6 VDD.t285 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X931 VSS.t461 VSS.t460 VSS.t461 VSS.t416 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X932 VDD IBIAS2.t32 IBIAS2.t33 VDD.t1107 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X933 IBIAS2 IBIAS2.t30 VDD.t758 VDD.t526 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X934 VDD IBIAS.t37 BD.t9 VDD.t111 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X935 VSS VB4.t86 IPD.t11 VSS.t192 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X936 OUT_P IBIAS2.t417 VDD.t646 VDD.t645 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X937 IVS IBIAS3.t62 VDD.t308 VDD.t306 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X938 VDD IBIAS2.t418 OUT_P.t90 VDD.t376 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X939 VDD.t1213 VDD.t1211 VDD.t1213 VDD.t1212 pfet_03v3 ad=1.76p pd=8.88u as=0 ps=0 w=4u l=0.28u
X940 OUT_P IBIAS2.t419 VDD.t649 VDD.t261 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X941 VSS VB4.t87 IPD.t10 VSS.t159 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X942 OUT_P IBIAS2.t420 VDD.t162 VDD.t161 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X943 OUT_N IBIAS2.t421 VDD.t164 VDD.t163 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X944 VND VB1.t56 VDD.t291 VDD.t290 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X945 BD IN_N.t19 IND.t54 VDD.t537 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X946 VDD.t1210 VDD.t1208 VDD.t1210 VDD.t1209 pfet_03v3 ad=1.65p pd=8.38u as=0 ps=0 w=3.75u l=0.28u
X947 VSS OUT2.t92 OUT_P.t13 VSS.t7 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X948 OUT2.t2 a_29248_n5498.t0 VDD.t165 ppolyf_u r_width=1u r_length=6.2u
X949 IBIAS2 IBIAS2.t28 VDD.t757 VDD.t142 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X950 VCD VCM.t14 VBM.t18 VSS.t4 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X951 VDD IBIAS2.t423 OUT_P.t87 VDD.t152 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X952 VSS.t459 VSS.t458 VSS.t459 VSS.t430 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X953 VSS.t457 VSS.t455 VSS.t457 VSS.t456 nfet_03v3 ad=0.88p pd=4.88u as=0 ps=0 w=2u l=1u
X954 VBM VCM.t15 VCD.t27 VSS.t140 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X955 IBS IBIAS1.t12 VDD.t622 VDD.t621 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X956 a_26254_n4340# a_25078_n5442# VDD.t13 ppolyf_u r_width=1u r_length=5u
X957 VSS OUT1.t82 OUT_N.t6 VSS.t24 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X958 VDD IBIAS2.t424 OUT_N.t105 VDD.t155 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X959 VDD IBIAS2.t425 OUT_N.t104 VDD.t158 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X960 IB2 VB2.t20 VB2.t21 VDD.t885 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X961 VDD VB1.t57 VPD.t5 VDD.t282 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X962 OUT_N IBIAS2.t426 VDD.t977 VDD.t125 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X963 VDD IBIAS2.t427 OUT_N.t102 VDD.t445 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X964 VSS.t454 VSS.t452 VSS.t454 VSS.t453 nfet_03v3 ad=0.26p pd=1.52u as=0 ps=0 w=1u l=0.28u
X965 VB1 VOUT.t22 VCD.t46 VSS.t3 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X966 BD IBIAS.t38 VDD.t346 VDD.t329 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X967 VDD IBIAS3.t63 IVS.t17 VDD.t406 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X968 VPD VB1.t58 VDD.t802 VDD.t770 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X969 VDD IBIAS2.t428 OUT_P.t86 VDD.t812 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X970 OUT1 VB3.t44 IND.t60 VSS.t391 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X971 VSS OUT2.t93 OUT_P.t14 VSS.t13 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X972 VB1 VOUT.t23 VCD.t57 VSS.t352 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X973 VDD IBIAS2.t429 OUT_N.t101 VDD.t442 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X974 VDD IBIAS3.t64 IVS.t16 VDD.t406 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X975 OUT_P OUT2.t94 VSS.t129 VSS.t79 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X976 VDD IBIAS2.t430 OUT_P.t85 VDD.t355 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X977 OUT_P IBIAS2.t431 VDD.t359 VDD.t358 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X978 OUT_P IBIAS2.t432 VDD.t911 VDD.t254 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X979 IB5 IB5.t8 VB4.t29 VSS.t615 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X980 OUT_P IBIAS2.t433 VDD.t912 VDD.t780 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X981 VDD VB1.t59 VND.t20 VDD.t285 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X982 IBIAS2 IBIAS2.t26 VDD.t756 VDD.t202 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X983 IPD IN_P.t15 BD.t23 VDD.t37 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X984 OUT_N IBIAS2.t435 VDD.t873 VDD.t587 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X985 VDD IBIAS3.t65 IVS.t15 VDD.t412 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X986 IPD IN_P.t16 BD.t24 VDD.t519 pfet_03v3 ad=1.65p pd=8.38u as=0.975p ps=4.27u w=3.75u l=0.28u
X987 VDD IBIAS2.t436 OUT_P.t81 VDD.t311 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X988 OUT_P IBIAS2.t437 VDD.t876 VDD.t252 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X989 OUT_N IBIAS2.t438 VDD.t383 VDD.t96 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X990 OUT_P OUT2.t95 VSS.t380 VSS.t101 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X991 VDD IBIAS2.t24 IBIAS2.t25 VDD.t145 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X992 VDD IBIAS3.t66 IVS.t14 VDD.t412 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X993 VDD.t1207 VDD.t1205 VDD.t1207 VDD.t1206 pfet_03v3 ad=1.76p pd=8.88u as=0 ps=0 w=4u l=0.28u
X994 IPD VB4.t88 VSS.t189 VSS.t164 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X995 VDD VB1.t60 VPD.t3 VDD.t761 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X996 OUT_P IBIAS2.t439 VDD.t384 VDD.t254 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X997 VOUT.t0 a_23622_n5442# VDD.t405 ppolyf_u r_width=1u r_length=5u
X998 VDD IBIAS1.t13 IB5.t0 VDD.t581 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X999 OUT_N OUT1.t83 VSS.t27 VSS.t22 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X1000 OUT_P IBIAS2.t440 VDD.t380 VDD.t379 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1001 VDD VB2.t66 IB2.t16 VDD.t540 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=1u
X1002 VSS.t451 VSS.t450 VSS.t451 VSS.t410 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X1003 VCD VCM.t16 VBM.t17 VSS.t599 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1004 OUT2 VB3.t45 IPD.t56 VSS.t0 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X1005 VSS VB4.t89 IPD.t8 VSS.t175 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X1006 a_26534_n6312# a_26254_n7414# VDD.t229 ppolyf_u r_width=1u r_length=5u
X1007 VDD IBIAS2.t441 OUT_P.t77 VDD.t83 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1008 VDD IBIAS2.t442 OUT_N.t98 VDD.t295 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1009 VSS IB4.t2 IB4.t3 VSS.t620 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X1010 VSS OUT1.t84 OUT_N.t8 VSS.t28 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1011 VCD VCM.t17 VBM.t16 VSS.t4 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1012 OUT_P IBIAS2.t443 VDD.t1052 VDD.t148 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1013 OUT_N IBIAS2.t444 VDD.t386 VDD.t385 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X1014 VCD VOUT.t24 VB1.t1 VSS.t6 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1015 VDD IBIAS2.t445 OUT_N.t96 VDD.t122 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1016 VB4 IB5.t6 IB5.t7 VSS.t695 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1017 VSS VB4.t90 IPD.t7 VSS.t175 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X1018 VSS OUT1.t85 OUT_N.t9 VSS.t13 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X1019 IND VB4.t91 VSS.t184 VSS.t162 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X1020 OUT_P IBIAS2.t446 VDD.t552 VDD.t551 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1021 OUT1.t24 a_29248_n7510.t2 VDD.t165 ppolyf_u r_width=1u r_length=6.2u
X1022 IPD VB4.t92 VSS.t183 VSS.t164 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X1023 OUT_N IBIAS2.t447 VDD.t553 VDD.t70 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1024 IB2 VB2.t18 VB2.t19 VDD.t592 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X1025 OUT2 VB3.t46 IPD.t36 VSS.t384 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X1026 VDD IBIAS2.t448 OUT_P.t74 VDD.t442 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1027 a_26534_n5442# a_25806_n7414# VDD.t573 ppolyf_u r_width=1u r_length=5u
X1028 VSS VB4.t16 VB4.t17 VSS.t180 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1029 BD IN_N.t20 IND.t8 VDD.t293 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X1030 OUT_P OUT2.t96 VSS.t381 VSS.t38 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X1031 VDD IBIAS2.t449 OUT_N.t94 VDD.t88 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1032 VDD IBIAS2.t450 OUT_N.t93 VDD.t236 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1033 VDD IBIAS2.t451 OUT_N.t92 VDD.t314 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1034 VSS OUT1.t86 OUT_N.t10 VSS.t33 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1035 OUT_N IBIAS2.t452 VDD.t890 VDD.t597 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1036 VDD IBIAS2.t453 OUT_P.t73 VDD.t152 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1037 IVS IVS.t60 VSS.t649 VSS.t636 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X1038 OUT_P IBIAS2.t454 VDD.t270 VDD.t3 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1039 VDD IBIAS2.t455 OUT_P.t71 VDD.t244 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1040 VDD IBIAS2.t456 OUT_N.t90 VDD.t38 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X1041 OUT_N IBIAS2.t457 VDD.t371 VDD.t263 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1042 BD IN_P.t17 IPD.t59 VDD.t418 pfet_03v3 ad=0.975p pd=4.27u as=1.65p ps=8.38u w=3.75u l=0.28u
X1043 VPD VB1.t61 VDD.t937 VDD.t290 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X1044 OUT_P IBIAS2.t458 VDD.t957 VDD.t385 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X1045 VB1 VOUT.t25 VCD.t63 VSS.t353 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X1046 VND VB2.t67 OUT1.t10 VDD.t354 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X1047 VDD IBIAS3.t67 IVS.t13 VDD.t167 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1048 VDD.t1204 VDD.t1203 VDD.t1204 VDD.t1174 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.56u
X1049 VDD IBIAS2.t459 OUT_N.t88 VDD.t98 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1050 OUT_N IBIAS2.t460 VDD.t588 VDD.t587 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1051 VDD IBIAS2.t461 OUT_P.t69 VDD.t91 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1052 OUT_P IBIAS2.t462 VDD.t576 VDD.t567 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1053 VDD IBIAS3.t68 IVS.t12 VDD.t186 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1054 VSS IB4.t23 IBIAS3.t3 VSS.t346 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X1055 VDD IBIAS2.t463 OUT_N.t86 VDD.t577 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1056 VB2 VB2.t2 IB2.t2 VDD.t886 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X1057 VDD.t1202 VDD.t1200 VDD.t1202 VDD.t1201 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1058 VCD VCM.t18 VBM.t15 VSS.t5 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1059 VDD VB1.t2 VB1.t3 VDD.t730 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X1060 OUT_P OUT2.t97 VSS.t382 VSS.t103 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1061 VSS OUT1.t87 OUT_N.t11 VSS.t19 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1062 VSS VB4.t93 IPD.t5 VSS.t159 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X1063 VSS VB4.t94 IND.t29 VSS.t175 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X1064 VDD.t1199 VDD.t1198 VDD.t1199 VDD.t1169 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X1065 a_25806_n4340# a_25526_n5442# VDD.t366 ppolyf_u r_width=1u r_length=5u
X1066 BD IBIAS.t39 VDD.t1098 VDD.t520 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X1067 IPD VB3.t47 OUT2.t12 VSS.t385 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X1068 OUT_P IBIAS2.t464 VDD.t126 VDD.t125 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1069 VDD IBIAS2.t465 OUT_P.t66 VDD.t127 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1070 OUT_P IBIAS2.t466 VDD.t855 VDD.t86 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1071 VDD.t1197 VDD.t1196 VDD.t1197 VDD.t1148 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X1072 OUT_N IBIAS2.t467 VDD.t856 VDD.t374 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X1073 VDD IBIAS2.t468 OUT_P.t64 VDD.t98 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1074 OUT_P IBIAS2.t469 VDD.t101 VDD.t19 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1075 VCD VOUT.t26 VB1.t22 VSS.t141 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X1076 VDD IBIAS2.t470 OUT_P.t62 VDD.t176 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1077 BD IN_P.t18 IPD.t60 VDD.t530 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X1078 IBIAS2 IBIAS2.t22 VDD.t1125 VDD.t336 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1079 OUT_N IBIAS2.t472 VDD.t66 VDD.t52 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1080 VDD IBIAS2.t473 OUT_P.t61 VDD.t67 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1081 OUT_N OUT1.t88 VSS.t305 VSS.t83 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1082 VSS OUT1.t89 OUT_N.t43 VSS.t19 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1083 OUT_N IBIAS2.t474 VDD.t71 VDD.t70 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1084 VDD.t1195 VDD.t1193 VDD.t1195 VDD.t1194 pfet_03v3 ad=1.65p pd=8.38u as=0 ps=0 w=3.75u l=0.28u
X1085 VDD IBIAS2.t475 OUT_N.t82 VDD.t624 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1086 VDD IBIAS2.t476 OUT_N.t81 VDD.t442 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1087 VDD.t1192 VDD.t1190 VDD.t1192 VDD.t1191 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1088 VDD IBIAS.t40 BD.t75 VDD.t267 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X1089 VSS OUT1.t90 OUT_N.t44 VSS.t114 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1090 IBIAS2 IVS.t88 VSS.t691 VSS.t342 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X1091 VDD IBIAS.t2 IBIAS.t3 VDD.t750 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X1092 VDD.t1189 VDD.t1187 VDD.t1189 VDD.t1188 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1093 VSS.t449 VSS.t448 VSS.t449 VSS.t413 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X1094 VDD VB1.t62 VND.t19 VDD.t761 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X1095 OUT_N IBIAS2.t477 VDD.t474 VDD.t379 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1096 OUT_P IBIAS2.t478 VDD.t475 VDD.t96 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1097 VSS.t447 VSS.t446 VSS.t447 VSS.t401 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1098 IBS IBS.t0 VSS.t614 VSS.t613 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=1u
X1099 IVS IBIAS3.t69 VDD.t185 VDD.t184 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1100 OUT_P OUT2.t98 VSS.t383 VSS.t68 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1101 OUT_N OUT1.t91 VSS.t310 VSS.t101 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X1102 VDD.t1186 VDD.t1184 VDD.t1186 VDD.t1185 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1103 BD IBIAS.t41 VDD.t1073 VDD.t522 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X1104 VSS OUT1.t92 OUT_N.t46 VSS.t40 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1105 OUT_N IBIAS2.t479 VDD.t692 VDD.t163 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1106 VSS.t445 VSS.t444 VSS.t445 VSS.t425 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1107 VSS.t443 VSS.t441 VSS.t443 VSS.t442 nfet_03v3 ad=0.52p pd=2.52u as=0 ps=0 w=2u l=1u
X1108 VDD IBIAS2.t480 OUT_N.t78 VDD.t221 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1109 VDD IBIAS2.t481 OUT_P.t59 VDD.t57 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1110 VCD VCM.t19 VBM.t14 VSS.t6 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1111 VPD VB1.t63 VDD.t940 VDD.t105 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X1112 BD IBIAS.t42 VDD.t1074 VDD.t520 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X1113 VDD IBIAS2.t20 IBIAS2.t21 VDD.t515 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1114 VBM VCM.t20 VCD.t22 VSS.t3 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1115 VB1 VOUT.t27 VCD.t65 VSS.t140 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1116 IPD VB4.t95 VSS.t174 VSS.t162 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X1117 OUT_N OUT1.t93 VSS.t314 VSS.t313 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1118 VSS OUT2.t99 OUT_P.t256 VSS.t24 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1119 IND VB3.t48 OUT1.t12 VSS.t2 nfet_03v3 ad=1.27p pd=6.64u as=1.27p ps=6.64u w=2.88u l=0.28u
X1120 VDD.t1183 VDD.t1181 VDD.t1183 VDD.t1182 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1121 VDD IBIAS2.t482 OUT_P.t58 VDD.t812 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1122 OUT_P IBIAS2.t483 VDD.t893 VDD.t567 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1123 OUT_N IBIAS2.t484 VDD.t894 VDD.t214 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X1124 VDD.t1180 VDD.t1178 VDD.t1180 VDD.t1179 pfet_03v3 ad=1.65p pd=8.38u as=0 ps=0 w=3.75u l=0.28u
X1125 VSS.t440 VSS.t439 VSS.t440 VSS.t413 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X1126 VDD.t1177 VDD.t1176 VDD.t1177 VDD.t1142 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1127 OUT_P IBIAS2.t485 VDD.t650 VDD.t597 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1128 OUT_P IBIAS2.t486 VDD.t651 VDD.t465 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1129 VSS.t438 VSS.t437 VSS.t438 VSS.t404 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X1130 IPD IN_P.t19 BD.t34 VDD.t230 pfet_03v3 ad=1.65p pd=8.38u as=0.975p ps=4.27u w=3.75u l=0.28u
X1131 VDD VB1.t64 VND.t18 VDD.t761 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X1132 VBM VCM.t21 VCD.t21 VSS.t352 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1133 VSS.t436 VSS.t435 VSS.t436 VSS.t407 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1134 OUT_N OUT1.t94 VSS.t627 VSS.t91 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1135 OUT_P OUT2.t100 VSS.t395 VSS.t91 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1136 IBIAS2 IBIAS2.t18 VDD.t785 VDD.t171 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1137 OUT_P OUT2.t101 VSS.t396 VSS.t68 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1138 VDD IBIAS2.t488 OUT_P.t54 VDD.t457 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1139 OUT_N IBIAS2.t489 VDD.t460 VDD.t52 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1140 VDD IBIAS3.t70 IVS.t10 VDD.t186 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1141 VDD.t1175 VDD.t1173 VDD.t1175 VDD.t1174 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.56u
X1142 OUT_P IBIAS2.t490 VDD.t462 VDD.t461 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1143 VDD IBIAS2.t491 OUT_N.t75 VDD.t675 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1144 a_24350_n4340# a_24070_n5442# VDD.t35 ppolyf_u r_width=1u r_length=5u
X1145 VDD.t1172 VDD.t1171 VDD.t1172 VDD.t1148 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X1146 VDD IBIAS2.t492 OUT_N.t74 VDD.t98 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1147 IVS IBIAS3.t71 VDD.t794 VDD.t531 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1148 VSS IVS.t58 IVS.t59 VSS.t624 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X1149 VSS.t434 VSS.t432 VSS.t434 VSS.t433 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X1150 OUT_N IBIAS2.t493 VDD.t80 VDD.t19 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1151 VDD IBIAS3.t72 IVS.t8 VDD.t186 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1152 VBM VCM.t22 VCD.t20 VSS.t353 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X1153 OUT_N IBIAS2.t494 VDD.t82 VDD.t81 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1154 VCD VOUT.t28 VB1.t26 VSS.t599 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1155 IPD IN_P.t20 BD.t29 VDD.t37 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X1156 IPD VB4.t96 VSS.t173 VSS.t164 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X1157 OUT_P OUT2.t102 VSS.t397 VSS.t71 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1158 VDD IBIAS2.t495 OUT_N.t71 VDD.t28 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1159 IBIAS2 IVS.t89 VSS.t692 VSS.t344 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X1160 VDD IBIAS.t43 BD.t0 VDD.t111 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X1161 OUT_P IBIAS2.t496 VDD.t572 VDD.t551 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1162 VDD IBIAS2.t497 OUT_P.t51 VDD.t32 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1163 VSS.t431 VSS.t429 VSS.t431 VSS.t430 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1164 OUT_N IBIAS2.t498 VDD.t739 VDD.t21 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1165 OUT_N OUT1.t95 VSS.t628 VSS.t79 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1166 IB3 VB3.t0 VB3.t1 VSS.t600 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1167 VSS.t428 VSS.t427 VSS.t428 VSS.t404 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X1168 OUT_P IBIAS2.t499 VDD.t1000 VDD.t454 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1169 IVS IBIAS3.t73 VDD.t362 VDD.t130 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1170 VSS VB4.t97 IND.t28 VSS.t159 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X1171 VBM VBM.t0 VDD.t352 VDD.t351 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X1172 VSS.t426 VSS.t424 VSS.t426 VSS.t425 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1173 OUT_N OUT1.t96 VSS.t629 VSS.t112 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1174 VSS.t423 VSS.t421 VSS.t423 VSS.t422 nfet_03v3 ad=0.26p pd=1.52u as=0 ps=0 w=1u l=0.28u
X1175 BD IN_P.t21 IPD.t54 VDD.t166 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X1176 VSS OUT1.t97 OUT_N.t258 VSS.t93 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X1177 VDD IBIAS2.t500 OUT_N.t69 VDD.t74 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1178 OUT_N IBIAS2.t501 VDD.t931 VDD.t389 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1179 VCD VCM.t23 VBM.t13 VSS.t6 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1180 VCD VOUT.t29 VB1.t8 VSS.t4 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1181 IPD VB3.t49 OUT2.t1 VSS.t1 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X1182 VND VB2.t69 OUT1.t11 VDD.t310 pfet_03v3 ad=1.38p pd=7.14u as=1.38p ps=7.14u w=3.13u l=0.28u
X1183 VCD VCM.t24 VBM.t12 VSS.t141 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X1184 VDD.t1170 VDD.t1168 VDD.t1170 VDD.t1169 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X1185 VDD IBIAS2.t502 OUT_P.t49 VDD.t155 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1186 VDD IBIAS2.t503 OUT_P.t48 VDD.t669 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1187 VDD IBIAS2.t504 OUT_P.t47 VDD.t483 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X1188 VDD.t1167 VDD.t1165 VDD.t1167 VDD.t1166 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1189 BD IN_N.t21 IND.t7 VDD.t292 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X1190 VDD IBIAS2.t505 OUT_N.t67 VDD.t54 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1191 OUT_P IBIAS2.t506 VDD.t1020 VDD.t275 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X1192 OUT_N IBIAS2.t507 VDD.t390 VDD.t389 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1193 VDD IBIAS2.t16 IBIAS2.t17 VDD.t23 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1194 IVS IBIAS3.t74 VDD.t363 VDD.t184 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1195 VSS VBIASN.t1 VBIASN.t2 VSS.t680 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X1196 VDD IBIAS2.t508 OUT_N.t65 VDD.t224 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1197 IBIAS2 IBIAS2.t14 VDD.t1075 VDD.t526 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1198 VDD IBIAS3.t75 IVS.t5 VDD.t331 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1199 VDD IBIAS3.t9 IBIAS3.t10 VDD.t320 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1200 VDD IBIAS2.t510 OUT_N.t64 VDD.t295 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1201 VDD IBIAS2.t511 OUT_P.t45 VDD.t122 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1202 IVS IBIAS3.t76 VDD.t920 VDD.t184 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1203 VPD VB2.t70 OUT2.t27 VDD.t104 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X1204 VSS.t420 VSS.t418 VSS.t420 VSS.t419 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1205 VSS OUT1.t98 OUT_N.t259 VSS.t98 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1206 IVS IVS.t56 VSS.t646 VSS.t618 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X1207 VDD.t1164 VDD.t1163 VDD.t1164 VDD.t1153 pfet_03v3 ad=0.814p pd=3.65u as=0 ps=0 w=3.13u l=0.56u
X1208 OUT_N IBIAS2.t512 VDD.t300 VDD.t148 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1209 VDD.t1162 VDD.t1161 VDD.t1162 VDD.t1145 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1210 VDD IBIAS2.t12 IBIAS2.t13 VDD.t515 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1211 OUT_N OUT1.t99 VSS.t634 VSS.t22 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X1212 VSS OUT1.t100 OUT_N.t0 VSS.t7 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X1213 VB3 VB3.t8 IB3.t0 VSS.t684 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1214 VSS IVS.t91 IBIAS2.t121 VSS.t339 nfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=1u
X1215 IND VB4.t98 VSS.t170 VSS.t164 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X1216 BD IBIAS.t44 VDD.t115 VDD.t114 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X1217 VSS OUT2.t103 OUT_P.t27 VSS.t16 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1218 VSS OUT2.t104 OUT_P.t28 VSS.t93 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X1219 VBM VCM.t25 VCD.t17 VSS.t353 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X1220 VDD IBIAS2.t513 OUT_N.t62 VDD.t469 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1221 OUT2.t10 a_29248_n5498.t1 VDD.t511 ppolyf_u r_width=1u r_length=6.2u
X1222 VBM VCM.t26 VCD.t16 VSS.t140 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1223 OUT_N IBIAS2.t514 VDD.t781 VDD.t780 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1224 VDD IBIAS.t45 BD.t73 VDD.t134 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X1225 VND VB2.t71 OUT1.t27 VDD.t309 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X1226 VSS OUT2.t105 OUT_P.t29 VSS.t24 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1227 VSS VB4.t14 VB4.t15 VSS.t167 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1228 VCD VOUT.t30 VB1.t15 VSS.t5 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1229 VDD.t1160 VDD.t1158 VDD.t1160 VDD.t1159 pfet_03v3 ad=1.04p pd=4.52u as=0 ps=0 w=4u l=0.28u
X1230 IPD IN_P.t22 BD.t31 VDD.t411 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X1231 VDD IBIAS2.t515 OUT_P.t44 VDD.t241 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1232 a_26254_n4340# a_26534_n5442# VDD.t229 ppolyf_u r_width=1u r_length=5u
X1233 VB2 VB2.t0 IB2.t1 VDD.t793 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X1234 VSS OUT1.t101 OUT_N.t1 VSS.t10 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1235 VSS OUT1.t102 OUT_N.t2 VSS.t13 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X1236 IBIAS2 IBIAS2.t10 VDD.t915 VDD.t142 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1237 IVS IBIAS3.t77 VDD.t532 VDD.t531 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1238 BD IN_N.t22 IND.t71 VDD.t361 pfet_03v3 ad=0.975p pd=4.27u as=1.65p ps=8.38u w=3.75u l=0.28u
X1239 OUT1 VB3.t51 IND.t0 VSS.t0 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X1240 VDD VB1.t65 VND.t17 VDD.t209 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X1241 VSS.t417 VSS.t415 VSS.t417 VSS.t416 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1242 VDD.t1157 VDD.t1155 VDD.t1157 VDD.t1156 pfet_03v3 ad=1.65p pd=8.38u as=0 ps=0 w=3.75u l=0.28u
X1243 VCD VCM.t27 VBM.t11 VSS.t141 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X1244 VDD.t1154 VDD.t1152 VDD.t1154 VDD.t1153 pfet_03v3 ad=0.814p pd=3.65u as=0 ps=0 w=3.13u l=0.56u
X1245 VDD IBIAS2.t517 OUT_N.t60 VDD.t376 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1246 VDD IBIAS2.t8 IBIAS2.t9 VDD.t173 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1247 OUT_N IBIAS2.t518 VDD.t775 VDD.t454 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1248 IVS IBIAS3.t78 VDD.t533 VDD.t531 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1249 IPD IN_P.t23 BD.t21 VDD.t620 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X1250 IBIAS2 IBIAS2.t6 VDD.t172 VDD.t171 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1251 VDD IBIAS2.t520 OUT_N.t58 VDD.t221 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1252 VDD.t1151 VDD.t1150 VDD.t1151 VDD.t1101 pfet_03v3 ad=1.76p pd=8.88u as=0 ps=0 w=4u l=0.28u
X1253 VDD IBIAS2.t521 OUT_P.t43 VDD.t155 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1254 VDD IBIAS2.t522 OUT_P.t42 VDD.t445 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1255 OUT_P IBIAS2.t523 VDD.t854 VDD.t3 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1256 IVS IBIAS3.t79 VDD.t131 VDD.t130 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1257 IPD VB4.t99 VSS.t166 VSS.t162 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X1258 OUT_P IBIAS2.t524 VDD.t302 VDD.t301 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1259 OUT_N IBIAS2.t525 VDD.t303 VDD.t5 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1260 a_25806_n4340# a_26534_n6312# VDD.t573 ppolyf_u r_width=1u r_length=5u
X1261 OUT_N IBIAS2.t526 VDD.t887 VDD.t780 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1262 IND VB4.t100 VSS.t165 VSS.t164 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X1263 VDD.t1149 VDD.t1147 VDD.t1149 VDD.t1148 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X1264 IBIAS2 IBIAS2.t4 VDD.t337 VDD.t336 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1265 IVS IBIAS3.t80 VDD.t132 VDD.t130 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1266 IB4 IBIAS4.t12 VDD.t897 VDD.t895 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1267 VSS.t414 VSS.t412 VSS.t414 VSS.t413 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X1268 VSS OUT1.t103 OUT_N.t3 VSS.t16 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1269 VDD IBIAS2.t528 OUT_N.t55 VDD.t355 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1270 VDD IBIAS2.t529 OUT_N.t54 VDD.t155 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1271 VDD.t1146 VDD.t1144 VDD.t1146 VDD.t1145 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1272 VDD IBIAS1.t14 IBS.t7 VDD.t767 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X1273 VDD.t1143 VDD.t1141 VDD.t1143 VDD.t1142 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1274 IB2 VB2.t16 VB2.t17 VDD.t323 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X1275 a_23622_n6312# a_24798_n7414# VDD.t766 ppolyf_u r_width=1u r_length=5u
X1276 VBM VCM.t28 VCD.t14 VSS.t142 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1277 VSS.t411 VSS.t409 VSS.t411 VSS.t410 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X1278 OUT_N IBIAS2.t530 VDD.t904 VDD.t252 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X1279 VDD IBIAS3.t7 IBIAS3.t8 VDD.t320 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1280 IPD VB4.t101 VSS.t163 VSS.t162 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X1281 VDD IBIAS2.t531 OUT_N.t52 VDD.t812 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1282 VND VB1.t66 VDD.t994 VDD.t290 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X1283 VSS OUT1.t104 OUT_N.t4 VSS.t19 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1284 VBM VCM.t29 VCD.t13 VSS.t140 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1285 VB1 VOUT.t31 VCD.t10 VSS.t3 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1286 OUT_N OUT1.t105 VSS.t23 VSS.t22 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X1287 OUT_N IBIAS2.t532 VDD.t554 VDD.t41 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1288 VDD IBIAS2.t533 OUT_P.t39 VDD.t77 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1289 VDD IBIAS3.t5 IBIAS3.t6 VDD.t320 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1290 VDD IBIAS4.t1 IBIAS4.t2 VDD.t843 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X1291 VPD VB2.t73 OUT2.t28 VDD.t310 pfet_03v3 ad=1.38p pd=7.14u as=1.38p ps=7.14u w=3.13u l=0.28u
X1292 IB5 IB5.t4 VB4.t28 VSS.t330 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1293 IND IN_N.t23 BD.t35 VDD.t230 pfet_03v3 ad=1.65p pd=8.38u as=0.975p ps=4.27u w=3.75u l=0.28u
X1294 OUT_N IBIAS2.t534 VDD.t564 VDD.t374 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X1295 OUT_P IBIAS2.t535 VDD.t565 VDD.t385 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X1296 IBIAS2 IBIAS2.t2 VDD.t335 VDD.t140 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1297 VDD IBIAS2.t0 IBIAS2.t1 VDD.t173 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1298 OUT_N OUT1.t106 VSS.t323 VSS.t38 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X1299 OUT_N IBIAS2.t537 VDD.t615 VDD.t94 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1300 OUT1.t22 a_29248_n7510.t1 VDD.t511 ppolyf_u r_width=1u r_length=6.2u
X1301 VSS.t408 VSS.t406 VSS.t408 VSS.t407 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1302 VDD IBIAS2.t538 OUT_P.t37 VDD.t295 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1303 IB4 IB4.t0 VSS.t63 VSS.t62 nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=1u
X1304 VSS.t405 VSS.t403 VSS.t405 VSS.t404 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X1305 IND VB3.t52 OUT1.t3 VSS.t2 nfet_03v3 ad=1.27p pd=6.64u as=1.27p ps=6.64u w=2.88u l=0.28u
X1306 OUT_P OUT2.t106 VSS.t304 VSS.t101 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X1307 VDD IBIAS2.t539 OUT_P.t36 VDD.t83 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1308 VSS VB4.t102 IND.t27 VSS.t159 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X1309 OUT_N OUT1.t107 VSS.t324 VSS.t313 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1310 VSS IB4.t25 IBIAS3.t4 VSS.t349 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X1311 VSS.t402 VSS.t400 VSS.t402 VSS.t401 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1312 VDD IBIAS2.t540 OUT_N.t48 VDD.t152 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1313 VSS VBIASN.t13 VCD.t5 VSS.t59 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X1314 OUT_P OUT2.t107 VSS.t635 VSS.t68 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1315 VDD IBIAS2.t541 OUT_P.t35 VDD.t666 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
R0 VB4.n130 VB4.t72 52.1434
R1 VB4.n129 VB4.t76 52.1434
R2 VB4.n128 VB4.t71 52.1434
R3 VB4.n127 VB4.t74 52.1434
R4 VB4.n126 VB4.t94 52.1434
R5 VB4.n125 VB4.t43 52.1434
R6 VB4.n124 VB4.t48 52.1434
R7 VB4.t37 VB4.n86 51.2309
R8 VB4.t61 VB4.n94 51.2309
R9 VB4.t82 VB4.n102 51.2309
R10 VB4.t96 VB4.n89 50.188
R11 VB4.t49 VB4.n96 50.188
R12 VB4.t70 VB4.n105 50.188
R13 VB4.t55 VB4.n123 49.6666
R14 VB4.t45 VB4.n91 48.8844
R15 VB4.t86 VB4.n111 48.8844
R16 VB4.t51 VB4.n115 48.8844
R17 VB4.t62 VB4.n114 48.8844
R18 VB4.t88 VB4.n90 48.6237
R19 VB4.t35 VB4.n92 48.6237
R20 VB4.t40 VB4.n99 48.6237
R21 VB4.t64 VB4.n106 48.6237
R22 VB4.t81 VB4.n113 48.6237
R23 VB4.n90 VB4.t96 48.1023
R24 VB4.n92 VB4.t50 48.1023
R25 VB4.n99 VB4.t54 48.1023
R26 VB4.n98 VB4.t49 48.1023
R27 VB4.n97 VB4.t52 48.1023
R28 VB4.n106 VB4.t70 48.1023
R29 VB4.n112 VB4.t93 48.1023
R30 VB4.n113 VB4.t91 48.1023
R31 VB4.n91 VB4.t88 47.8416
R32 VB4.n111 VB4.t35 47.8416
R33 VB4.n110 VB4.t40 47.8416
R34 VB4.n109 VB4.t34 47.8416
R35 VB4.n108 VB4.t39 47.8416
R36 VB4.n107 VB4.t64 47.8416
R37 VB4.n114 VB4.t81 47.8416
R38 VB4.n115 VB4.t85 47.8416
R39 VB4.n133 VB4.t55 47.3393
R40 VB4.n123 VB4.t45 47.0594
R41 VB4.n122 VB4.t86 47.0594
R42 VB4.n121 VB4.t75 47.0594
R43 VB4.n120 VB4.t65 47.0594
R44 VB4.n119 VB4.t53 47.0594
R45 VB4.n118 VB4.t90 47.0594
R46 VB4.n116 VB4.t51 47.0594
R47 VB4.n117 VB4.t62 47.0594
R48 VB4.n89 VB4.t37 46.538
R49 VB4.n88 VB4.t63 46.538
R50 VB4.n87 VB4.t69 46.538
R51 VB4.n96 VB4.t61 46.538
R52 VB4.n95 VB4.t66 46.538
R53 VB4.n105 VB4.t82 46.538
R54 VB4.n104 VB4.t99 46.538
R55 VB4.n103 VB4.t102 46.538
R56 VB4.t92 VB4.n83 45.8862
R57 VB4.n86 VB4.t92 45.4951
R58 VB4.n85 VB4.t38 45.4951
R59 VB4.n84 VB4.t44 45.4951
R60 VB4.n94 VB4.t36 45.4951
R61 VB4.n93 VB4.t42 45.4951
R62 VB4.n102 VB4.t68 45.4951
R63 VB4.n100 VB4.t87 45.4951
R64 VB4.n101 VB4.t83 45.4951
R65 VB4.n77 VB4.t95 45.2344
R66 VB4.n83 VB4.t100 45.2344
R67 VB4.n82 VB4.t57 45.2344
R68 VB4.n81 VB4.t59 45.2344
R69 VB4.n80 VB4.t56 45.2344
R70 VB4.n79 VB4.t58 45.2344
R71 VB4.n78 VB4.t78 45.2344
R72 VB4.n76 VB4.t97 45.2344
R73 VB4.n130 VB4.t46 44.5826
R74 VB4.n129 VB4.t84 44.5826
R75 VB4.n128 VB4.t32 44.5826
R76 VB4.n127 VB4.t77 44.5826
R77 VB4.n126 VB4.t89 44.5826
R78 VB4.n125 VB4.t101 44.5826
R79 VB4.n124 VB4.t73 44.5826
R80 VB4.n131 VB4.t98 44.5826
R81 VB4.n61 VB4.t20 17.0773
R82 VB4.n43 VB4.t8 17.0773
R83 VB4.n40 VB4.t14 17.0773
R84 VB4.n38 VB4.t4 17.0773
R85 VB4.n35 VB4.t26 17.0773
R86 VB4.n33 VB4.t0 17.0773
R87 VB4.n30 VB4.t22 17.0773
R88 VB4.n28 VB4.t10 17.0773
R89 VB4.n25 VB4.t18 17.0773
R90 VB4.n23 VB4.t6 17.0773
R91 VB4.n20 VB4.t16 17.0773
R92 VB4.n18 VB4.t2 17.0773
R93 VB4.n56 VB4.t12 17.0773
R94 VB4.n54 VB4.t24 17.0773
R95 VB4.n78 VB4.n77 9.73383
R96 VB4.n77 VB4.n76 9.73383
R97 VB4.n86 VB4.n85 9.73383
R98 VB4.n85 VB4.n84 9.73383
R99 VB4.n94 VB4.n93 9.73383
R100 VB4.n102 VB4.n101 9.73383
R101 VB4.n101 VB4.n100 9.73383
R102 VB4.n89 VB4.n88 9.73383
R103 VB4.n88 VB4.n87 9.73383
R104 VB4.n96 VB4.n95 9.73383
R105 VB4.n105 VB4.n104 9.73383
R106 VB4.n104 VB4.n103 9.73383
R107 VB4.n99 VB4.n98 9.73383
R108 VB4.n98 VB4.n97 9.73383
R109 VB4.n113 VB4.n112 9.73383
R110 VB4.n111 VB4.n110 9.73383
R111 VB4.n110 VB4.n109 9.73383
R112 VB4.n109 VB4.n108 9.73383
R113 VB4.n108 VB4.n107 9.73383
R114 VB4.n123 VB4.n122 9.73383
R115 VB4.n122 VB4.n121 9.73383
R116 VB4.n121 VB4.n120 9.73383
R117 VB4.n120 VB4.n119 9.73383
R118 VB4.n119 VB4.n118 9.73383
R119 VB4.n118 VB4.n117 9.73383
R120 VB4.n117 VB4.n116 9.73383
R121 VB4.n131 VB4.n130 9.73383
R122 VB4.n130 VB4.n129 9.73383
R123 VB4.n129 VB4.n128 9.73383
R124 VB4.n128 VB4.n127 9.73383
R125 VB4.n127 VB4.n126 9.73383
R126 VB4.n126 VB4.n125 9.73383
R127 VB4.n125 VB4.n124 9.73383
R128 VB4.n79 VB4.n78 9.28449
R129 VB4.n83 VB4.n82 7.16614
R130 VB4.n82 VB4.n81 7.16614
R131 VB4.n81 VB4.n80 7.16614
R132 VB4.n80 VB4.n79 7.16614
R133 VB4.n136 VB4.n135 6.78515
R134 VB4.n52 VB4.t29 5.69633
R135 VB4.n19 VB4.n17 5.22676
R136 VB4.n64 VB4.n63 4.5005
R137 VB4.n55 VB4.n54 4.0005
R138 VB4.n57 VB4.n56 4.0005
R139 VB4.n19 VB4.n18 4.0005
R140 VB4.n21 VB4.n20 4.0005
R141 VB4.n24 VB4.n23 4.0005
R142 VB4.n26 VB4.n25 4.0005
R143 VB4.n29 VB4.n28 4.0005
R144 VB4.n31 VB4.n30 4.0005
R145 VB4.n34 VB4.n33 4.0005
R146 VB4.n36 VB4.n35 4.0005
R147 VB4.n39 VB4.n38 4.0005
R148 VB4.n41 VB4.n40 4.0005
R149 VB4.n44 VB4.n43 4.0005
R150 VB4.n62 VB4.n61 4.0005
R151 VB4.n58 VB4.n47 3.43224
R152 VB4.n52 VB4.n51 3.43224
R153 VB4.n42 VB4.n8 3.43224
R154 VB4.n37 VB4.n10 3.43224
R155 VB4.n32 VB4.n12 3.43224
R156 VB4.n27 VB4.n14 3.43224
R157 VB4.n22 VB4.n16 3.43224
R158 VB4.n53 VB4.n49 3.1505
R159 VB4.n70 VB4.n69 3.0736
R160 VB4.n139 VB4.n134 2.8805
R161 VB4.n133 VB4.n132 2.82317
R162 VB4.n150 VB4.n149 1.81328
R163 VB4.n47 VB4.t21 1.6385
R164 VB4.n47 VB4.n46 1.6385
R165 VB4.n49 VB4.t25 1.6385
R166 VB4.n49 VB4.n48 1.6385
R167 VB4.n51 VB4.t28 1.6385
R168 VB4.n51 VB4.n50 1.6385
R169 VB4.n8 VB4.t15 1.6385
R170 VB4.n8 VB4.n7 1.6385
R171 VB4.n10 VB4.t27 1.6385
R172 VB4.n10 VB4.n9 1.6385
R173 VB4.n12 VB4.t23 1.6385
R174 VB4.n12 VB4.n11 1.6385
R175 VB4.n14 VB4.t19 1.6385
R176 VB4.n14 VB4.n13 1.6385
R177 VB4.n16 VB4.t17 1.6385
R178 VB4.n16 VB4.n15 1.6385
R179 VB4.n147 VB4.n146 1.50393
R180 VB4.n73 VB4.n72 1.49812
R181 VB4.n61 VB4.n60 1.31856
R182 VB4.n134 VB4.n133 1.18887
R183 VB4.n154 VB4.n153 1.12675
R184 VB4.n154 VB4.n74 1.126
R185 VB4.n68 VB4.n65 1.11382
R186 VB4.n53 VB4.n52 0.908326
R187 VB4.n146 VB4.n139 0.901294
R188 VB4.n132 VB4.n131 0.548
R189 VB4.n55 VB4.n53 0.438761
R190 VB4.n57 VB4.n55 0.313543
R191 VB4.n21 VB4.n19 0.313543
R192 VB4.n26 VB4.n24 0.313543
R193 VB4.n31 VB4.n29 0.313543
R194 VB4.n36 VB4.n34 0.313543
R195 VB4.n41 VB4.n39 0.313543
R196 VB4.n45 VB4.n44 0.202326
R197 VB4.n22 VB4.n21 0.157022
R198 VB4.n24 VB4.n22 0.157022
R199 VB4.n27 VB4.n26 0.157022
R200 VB4.n29 VB4.n27 0.157022
R201 VB4.n32 VB4.n31 0.157022
R202 VB4.n34 VB4.n32 0.157022
R203 VB4.n37 VB4.n36 0.157022
R204 VB4.n39 VB4.n37 0.157022
R205 VB4.n42 VB4.n41 0.157022
R206 VB4.n44 VB4.n42 0.157022
R207 VB4 VB4.n154 0.111701
R208 VB4.n58 VB4.n57 0.104587
R209 VB4.n138 VB4.n137 0.0656316
R210 VB4.n59 VB4.n58 0.034
R211 VB4.n143 VB4.n142 0.0339644
R212 VB4.n144 VB4.n143 0.0327802
R213 VB4.n139 VB4.n138 0.0301053
R214 VB4.n145 VB4.n144 0.0301053
R215 VB4.n68 VB4.n67 0.0298454
R216 VB4.n137 VB4.n136 0.0289211
R217 VB4.n142 VB4.n141 0.0289211
R218 VB4.n69 VB4.n68 0.0256315
R219 VB4.n6 VB4.n5 0.0207053
R220 VB4.n1 VB4.n0 0.0207053
R221 VB4.n4 VB4.n3 0.014
R222 VB4.n5 VB4.n4 0.0134654
R223 VB4.n149 VB4.n148 0.00858096
R224 VB4.n148 VB4.n147 0.00858096
R225 VB4.n147 VB4.n75 0.00858096
R226 VB4.n153 VB4.n151 0.00773989
R227 VB4.n71 VB4.n70 0.00773989
R228 VB4.n151 VB4.n150 0.00773989
R229 VB4.n72 VB4.n71 0.00773989
R230 VB4.n3 VB4.n2 0.00773989
R231 VB4.n153 VB4.n152 0.00773989
R232 VB4.n72 VB4.n6 0.00773989
R233 VB4.n74 VB4.n1 0.00773989
R234 VB4.n65 VB4.n64 0.0075
R235 VB4.n62 VB4.n59 0.007
R236 VB4.n141 VB4.n140 0.00685938
R237 VB4.n65 VB4.n45 0.0065
R238 VB4.n74 VB4.n73 0.00582347
R239 VB4.n64 VB4.n62 0.0055
R240 VB4.n67 VB4.n66 0.0045
R241 VB4.n146 VB4.n145 0.0030309
R242 IND.n318 IND.t66 4.62366
R243 IND.n344 IND.n343 4.62366
R244 IND.n56 IND.n55 4.37688
R245 IND.n110 IND.n109 4.34373
R246 IND.n96 IND.n95 4.34373
R247 IND.n62 IND.n61 4.34007
R248 IND.n330 IND.n329 4.13833
R249 IND.n313 IND.n312 2.31142
R250 IND.n436 IND.n435 1.66567
R251 IND.n460 IND.t28 1.66567
R252 IND.n365 IND.n363 1.6654
R253 IND.n390 IND.t27 1.6654
R254 IND.n200 IND.n198 1.66411
R255 IND.n225 IND.t30 1.66411
R256 IND.n473 IND.n472 1.49812
R257 IND.n91 IND.n90 1.49201
R258 IND.n80 IND.t38 1.49201
R259 IND.n298 IND.n297 1.49175
R260 IND.n287 IND.t58 1.49175
R261 IND.n177 IND.n176 1.49048
R262 IND.n166 IND.t68 1.49048
R263 IND.n106 IND.n105 1.47245
R264 IND.n101 IND.n100 1.47245
R265 IND.n52 IND.n51 1.46565
R266 IND.n2 IND.n1 1.31982
R267 IND.n13 IND.t44 1.31982
R268 IND.n142 IND.t47 1.31982
R269 IND.n138 IND.n137 1.31982
R270 IND.n259 IND.n258 1.23423
R271 IND.n403 IND.n402 1.19479
R272 IND.n294 IND.n293 1.19462
R273 IND.n92 IND.n91 1.19459
R274 IND.n81 IND.n80 1.19459
R275 IND.n173 IND.n172 1.19439
R276 IND.n9 IND.n8 1.19395
R277 IND.n154 IND.n153 1.19395
R278 IND.n143 IND.n142 1.19393
R279 IND.n87 IND.n86 1.17958
R280 IND.n44 IND.n43 1.17929
R281 IND.n276 IND.n275 1.17929
R282 IND.n299 IND.n298 1.17924
R283 IND.n288 IND.n287 1.17924
R284 IND.n178 IND.n177 1.17917
R285 IND.n167 IND.n166 1.17917
R286 IND.n409 IND.n408 1.17907
R287 IND.n33 IND.n32 1.17902
R288 IND.n265 IND.n264 1.17902
R289 IND.n3 IND.n2 1.1787
R290 IND.n14 IND.n13 1.1787
R291 IND.n139 IND.n138 1.1787
R292 IND.n474 IND.n425 1.1775
R293 IND.n216 IND.n215 1.16728
R294 IND.n381 IND.n380 1.16675
R295 IND.n242 IND.n241 1.16675
R296 IND.n254 IND.n253 1.16675
R297 IND.n68 IND.n67 1.16667
R298 IND.n201 IND.n200 1.16641
R299 IND.n226 IND.n225 1.16641
R300 IND.n450 IND.n449 1.16617
R301 IND.n366 IND.n365 1.16588
R302 IND.n391 IND.n390 1.16588
R303 IND.n317 IND.n316 1.1658
R304 IND.n336 IND.n335 1.1658
R305 IND.n350 IND.n349 1.1658
R306 IND.n437 IND.n436 1.1656
R307 IND.n461 IND.n460 1.1656
R308 IND.n422 IND.n28 1.1515
R309 IND.n358 IND.n78 1.1515
R310 IND.n285 IND.n135 1.1515
R311 IND.n107 IND.n106 1.14066
R312 IND.n102 IND.n101 1.14066
R313 IND.n53 IND.n52 1.14059
R314 IND.n15 IND.n14 1.12717
R315 IND.n382 IND.n381 1.1257
R316 IND.n243 IND.n242 1.1257
R317 IND.n217 IND.n216 1.1257
R318 IND.n320 IND.n319 1.1255
R319 IND.n332 IND.n331 1.1255
R320 IND.n346 IND.n345 1.1255
R321 IND.n58 IND.n57 1.1255
R322 IND.n64 IND.n63 1.1255
R323 IND.n112 IND.n111 1.1255
R324 IND.n98 IND.n97 1.1255
R325 IND.n284 IND.n283 1.1255
R326 IND.n357 IND.n356 1.1255
R327 IND.n421 IND.n420 1.1255
R328 IND.n474 IND.n473 1.1255
R329 IND.n452 IND.n451 1.10737
R330 IND.n368 IND.n367 1.1073
R331 IND.n393 IND.n392 1.1073
R332 IND.n256 IND.n255 1.1073
R333 IND.n203 IND.n202 1.1073
R334 IND.n228 IND.n227 1.1073
R335 IND.n449 IND.n448 1.09663
R336 IND.n380 IND.n378 1.09644
R337 IND.n241 IND.n239 1.09644
R338 IND.n253 IND.n252 1.09644
R339 IND.n215 IND.n213 1.09514
R340 IND.n67 IND.n66 1.08656
R341 IND.n396 IND.n395 1.05423
R342 IND.n397 IND.n49 1.05265
R343 IND.n259 IND.n231 1.0087
R344 IND.n316 IND.n315 1.00677
R345 IND.n335 IND.n334 1.00677
R346 IND.n349 IND.n348 1.00677
R347 IND.n293 IND.n292 0.922998
R348 IND.n86 IND.n85 0.922926
R349 IND.n172 IND.n171 0.92139
R350 IND.n408 IND.n407 0.920264
R351 IND.n402 IND.n401 0.920264
R352 IND.n439 IND.n438 0.88565
R353 IND.n463 IND.n462 0.88565
R354 IND.n43 IND.n42 0.834379
R355 IND.n275 IND.n274 0.834379
R356 IND.n32 IND.n31 0.834365
R357 IND.n264 IND.n263 0.834365
R358 IND.n8 IND.n7 0.834193
R359 IND.n153 IND.n152 0.834193
R360 IND.n122 IND.n121 0.759312
R361 IND.n47 IND.n46 0.727916
R362 IND.n338 IND.n337 0.727916
R363 IND.n352 IND.n351 0.727916
R364 IND.n279 IND.n278 0.727916
R365 IND.n157 IND.n156 0.727916
R366 IND.n25 IND.n4 0.727104
R367 IND.n416 IND.n404 0.727104
R368 IND.n71 IND.n69 0.727104
R369 IND.n306 IND.n295 0.727104
R370 IND.n119 IND.n103 0.727104
R371 IND.n128 IND.n88 0.727104
R372 IND.n162 IND.n140 0.727104
R373 IND.n181 IND.n179 0.727104
R374 IND.n190 IND.n168 0.727104
R375 IND.n313 IND.n285 0.656743
R376 IND.n419 IND.n418 0.650188
R377 IND.n78 IND.n77 0.650188
R378 IND.n20 IND.n10 0.616779
R379 IND.n412 IND.n410 0.616779
R380 IND.n36 IND.n34 0.616779
R381 IND.n323 IND.n321 0.616779
R382 IND.n76 IND.n59 0.616779
R383 IND.n302 IND.n300 0.616779
R384 IND.n311 IND.n289 0.616779
R385 IND.n268 IND.n266 0.616779
R386 IND.n115 IND.n113 0.616779
R387 IND.n124 IND.n93 0.616779
R388 IND.n133 IND.n82 0.616779
R389 IND.n146 IND.n144 0.616779
R390 IND.n186 IND.n174 0.616779
R391 IND.n407 IND.t40 0.56925
R392 IND.n407 IND.n406 0.56925
R393 IND.n401 IND.t33 0.56925
R394 IND.n401 IND.n400 0.56925
R395 IND.n378 IND.t36 0.56925
R396 IND.n378 IND.n377 0.56925
R397 IND.n66 IND.t39 0.56925
R398 IND.n66 IND.n65 0.56925
R399 IND.n61 IND.t41 0.56925
R400 IND.n61 IND.n60 0.56925
R401 IND.n51 IND.t32 0.56925
R402 IND.n51 IND.n50 0.56925
R403 IND.n55 IND.t35 0.56925
R404 IND.n55 IND.n54 0.56925
R405 IND.n292 IND.t55 0.56925
R406 IND.n292 IND.n291 0.56925
R407 IND.n105 IND.t0 0.56925
R408 IND.n105 IND.n104 0.56925
R409 IND.n109 IND.t67 0.56925
R410 IND.n109 IND.n108 0.56925
R411 IND.n100 IND.t70 0.56925
R412 IND.n100 IND.n99 0.56925
R413 IND.n95 IND.t60 0.56925
R414 IND.n95 IND.n94 0.56925
R415 IND.n85 IND.t34 0.56925
R416 IND.n85 IND.n84 0.56925
R417 IND.n239 IND.t31 0.56925
R418 IND.n239 IND.n238 0.56925
R419 IND.n252 IND.t29 0.56925
R420 IND.n252 IND.n251 0.56925
R421 IND.n171 IND.t63 0.56925
R422 IND.n171 IND.n170 0.56925
R423 IND.n213 IND.t42 0.56925
R424 IND.n213 IND.n212 0.56925
R425 IND.n448 IND.t37 0.56925
R426 IND.n448 IND.n447 0.56925
R427 IND.n231 IND.n230 0.516159
R428 IND.n193 IND.n192 0.507313
R429 IND.n7 IND.t3 0.485833
R430 IND.n7 IND.n6 0.485833
R431 IND.n31 IND.t5 0.485833
R432 IND.n31 IND.n30 0.485833
R433 IND.n42 IND.t8 0.485833
R434 IND.n42 IND.n41 0.485833
R435 IND.n315 IND.t71 0.485833
R436 IND.n334 IND.t49 0.485833
R437 IND.n334 IND.n333 0.485833
R438 IND.n329 IND.t54 0.485833
R439 IND.n329 IND.n328 0.485833
R440 IND.n348 IND.n347 0.485833
R441 IND.n263 IND.t50 0.485833
R442 IND.n263 IND.n262 0.485833
R443 IND.n274 IND.t7 0.485833
R444 IND.n274 IND.n273 0.485833
R445 IND.n152 IND.t51 0.485833
R446 IND.n152 IND.n151 0.485833
R447 IND.n465 IND.n464 0.475688
R448 IND.n304 IND.n303 0.474125
R449 IND.n309 IND.n308 0.474125
R450 IND.n117 IND.n116 0.474125
R451 IND.n184 IND.n183 0.474125
R452 IND.n188 IND.n187 0.474125
R453 IND.n282 IND.n281 0.470187
R454 IND.n135 IND.n134 0.470187
R455 IND.n396 IND.n358 0.419368
R456 IND.n260 IND.n259 0.395709
R457 IND.n397 IND.n396 0.390055
R458 IND.n423 IND.n422 0.368687
R459 IND.n231 IND.n164 0.336564
R460 IND.n39 IND.n38 0.330687
R461 IND.n271 IND.n270 0.330687
R462 IND.n23 IND.n22 0.330125
R463 IND.n19 IND.n18 0.330125
R464 IND.n414 IND.n413 0.330125
R465 IND.n371 IND.n370 0.330125
R466 IND.n384 IND.n383 0.330125
R467 IND.n341 IND.n340 0.330125
R468 IND.n326 IND.n325 0.330125
R469 IND.n74 IND.n73 0.330125
R470 IND.n126 IND.n125 0.330125
R471 IND.n131 IND.n130 0.330125
R472 IND.n245 IND.n244 0.330125
R473 IND.n160 IND.n159 0.330125
R474 IND.n149 IND.n148 0.330125
R475 IND.n206 IND.n205 0.330125
R476 IND.n219 IND.n218 0.330125
R477 IND.n441 IND.n440 0.330125
R478 IND.n455 IND.n454 0.330125
R479 IND.n28 IND.n27 0.29075
R480 IND.n355 IND.n354 0.29075
R481 IND.n398 IND.n397 0.262189
R482 IND.n314 IND.n313 0.203334
R483 IND.n462 IND.n458 0.0936537
R484 IND.n438 IND.n433 0.0936537
R485 IND.n202 IND.n197 0.0910426
R486 IND.n227 IND.n223 0.0910426
R487 IND.n367 IND.n362 0.0886741
R488 IND.n392 IND.n388 0.0886741
R489 IND.n255 IND.n249 0.0886741
R490 IND.n451 IND.n445 0.0880141
R491 IND.n14 IND.n12 0.0832399
R492 IND.n46 IND.n45 0.0826464
R493 IND.n337 IND.n336 0.0826464
R494 IND.n351 IND.n350 0.0826464
R495 IND.n278 IND.n277 0.0826464
R496 IND.n156 IND.n155 0.0826464
R497 IND.n4 IND.n0 0.0823987
R498 IND.n404 IND.n399 0.0823987
R499 IND.n69 IND.n64 0.0823987
R500 IND.n295 IND.n290 0.0823987
R501 IND.n103 IND.n98 0.0823987
R502 IND.n88 IND.n83 0.0823987
R503 IND.n140 IND.n136 0.0823987
R504 IND.n179 IND.n175 0.0823987
R505 IND.n168 IND.n165 0.0823987
R506 IND.n215 IND.n214 0.0801656
R507 IND.n200 IND.n199 0.0800575
R508 IND.n225 IND.n224 0.0800575
R509 IND.n380 IND.n379 0.0784141
R510 IND.n241 IND.n240 0.0784141
R511 IND.n253 IND.n250 0.0784141
R512 IND.n365 IND.n364 0.0783056
R513 IND.n390 IND.n389 0.0783056
R514 IND.n449 IND.n446 0.0778549
R515 IND.n436 IND.n434 0.0774429
R516 IND.n460 IND.n459 0.0774429
R517 IND.n10 IND.n5 0.0712285
R518 IND.n410 IND.n405 0.0712285
R519 IND.n34 IND.n29 0.0712285
R520 IND.n321 IND.n317 0.0712285
R521 IND.n59 IND.n53 0.0712285
R522 IND.n289 IND.n286 0.0712285
R523 IND.n300 IND.n296 0.0712285
R524 IND.n266 IND.n261 0.0712285
R525 IND.n82 IND.n79 0.0712285
R526 IND.n93 IND.n89 0.0712285
R527 IND.n113 IND.n107 0.0712285
R528 IND.n144 IND.n141 0.0712285
R529 IND.n174 IND.n169 0.0712285
R530 IND.n63 IND.n62 0.0631087
R531 IND.n381 IND.n376 0.0623855
R532 IND.n242 IND.n237 0.0623855
R533 IND.n216 IND.n211 0.0623855
R534 IND.n211 IND.n210 0.060017
R535 IND IND.n474 0.058875
R536 IND.n376 IND.n375 0.0576486
R537 IND.n237 IND.n236 0.0576486
R538 IND.n319 IND.n318 0.0572391
R539 IND.n331 IND.n330 0.0572391
R540 IND.n345 IND.n344 0.0572391
R541 IND.n10 IND.n9 0.0534597
R542 IND.n410 IND.n409 0.0534597
R543 IND.n34 IND.n33 0.0534597
R544 IND.n321 IND.n320 0.0534597
R545 IND.n59 IND.n58 0.0534597
R546 IND.n300 IND.n299 0.0534597
R547 IND.n289 IND.n288 0.0534597
R548 IND.n266 IND.n265 0.0534597
R549 IND.n113 IND.n112 0.0534597
R550 IND.n93 IND.n92 0.0534597
R551 IND.n82 IND.n81 0.0534597
R552 IND.n144 IND.n143 0.0534597
R553 IND.n174 IND.n173 0.0534597
R554 IND.n285 IND.n284 0.0525
R555 IND.n284 IND.n260 0.0525
R556 IND.n358 IND.n357 0.0525
R557 IND.n357 IND.n314 0.0525
R558 IND.n422 IND.n421 0.0525
R559 IND.n421 IND.n398 0.0525
R560 IND.n46 IND.n44 0.0423164
R561 IND.n337 IND.n332 0.0423164
R562 IND.n351 IND.n346 0.0423164
R563 IND.n278 IND.n276 0.0423164
R564 IND.n156 IND.n154 0.0423164
R565 IND.n12 IND.n11 0.0419676
R566 IND.n4 IND.n3 0.0415773
R567 IND.n404 IND.n403 0.0415773
R568 IND.n69 IND.n68 0.0415773
R569 IND.n295 IND.n294 0.0415773
R570 IND.n88 IND.n87 0.0415773
R571 IND.n103 IND.n102 0.0415773
R572 IND.n140 IND.n139 0.0415773
R573 IND.n168 IND.n167 0.0415773
R574 IND.n179 IND.n178 0.0415773
R575 IND.n392 IND.n391 0.032498
R576 IND.n367 IND.n366 0.032498
R577 IND.n255 IND.n254 0.032498
R578 IND.n227 IND.n226 0.032498
R579 IND.n202 IND.n201 0.032498
R580 IND.n451 IND.n450 0.0319869
R581 IND.n57 IND.n56 0.0269366
R582 IND.n420 IND.n419 0.0265
R583 IND.n356 IND.n355 0.0265
R584 IND.n283 IND.n282 0.0265
R585 IND.n462 IND.n461 0.0261793
R586 IND.n438 IND.n437 0.0261793
R587 IND.n472 IND.n471 0.0236139
R588 IND.n428 IND.n427 0.0207053
R589 IND.n471 IND.n470 0.0207053
R590 IND.n111 IND.n110 0.0191828
R591 IND.n97 IND.n96 0.0191828
R592 IND.n20 IND.n19 0.0156875
R593 IND.n413 IND.n412 0.0156875
R594 IND.n36 IND.n35 0.0156875
R595 IND.n372 IND.n371 0.0156875
R596 IND.n323 IND.n322 0.0156875
R597 IND.n77 IND.n76 0.0156875
R598 IND.n303 IND.n302 0.0156875
R599 IND.n312 IND.n311 0.0156875
R600 IND.n268 IND.n267 0.0156875
R601 IND.n116 IND.n115 0.0156875
R602 IND.n125 IND.n124 0.0156875
R603 IND.n134 IND.n133 0.0156875
R604 IND.n233 IND.n232 0.0156875
R605 IND.n146 IND.n145 0.0156875
R606 IND.n187 IND.n186 0.0156875
R607 IND.n207 IND.n206 0.0156875
R608 IND.n439 IND.n430 0.0156875
R609 IND.n440 IND.n439 0.0156875
R610 IND.n463 IND.n455 0.0156875
R611 IND.n464 IND.n463 0.0156875
R612 IND.n222 IND.n221 0.0151213
R613 IND.n196 IND.n195 0.0151213
R614 IND.n473 IND.n429 0.014
R615 IND.n387 IND.n386 0.0139513
R616 IND.n361 IND.n360 0.0139513
R617 IND.n248 IND.n247 0.0139513
R618 IND.n429 IND.n428 0.0134654
R619 IND.n444 IND.n443 0.0133659
R620 IND.n383 IND.n382 0.0123533
R621 IND.n244 IND.n243 0.0123533
R622 IND.n218 IND.n217 0.0123533
R623 IND.n370 IND.n369 0.0111023
R624 IND.n395 IND.n394 0.0111023
R625 IND.n258 IND.n257 0.0111023
R626 IND.n205 IND.n204 0.0111023
R627 IND.n230 IND.n229 0.0111023
R628 IND.n454 IND.n453 0.0111023
R629 IND.n25 IND.n24 0.00860784
R630 IND.n21 IND.n20 0.00860784
R631 IND.n17 IND.n16 0.00860784
R632 IND.n412 IND.n411 0.00860784
R633 IND.n417 IND.n416 0.00860784
R634 IND.n37 IND.n36 0.00860784
R635 IND.n368 IND.n359 0.00860784
R636 IND.n393 IND.n385 0.00860784
R637 IND.n324 IND.n323 0.00860784
R638 IND.n72 IND.n71 0.00860784
R639 IND.n76 IND.n75 0.00860784
R640 IND.n302 IND.n301 0.00860784
R641 IND.n307 IND.n306 0.00860784
R642 IND.n311 IND.n310 0.00860784
R643 IND.n269 IND.n268 0.00860784
R644 IND.n115 IND.n114 0.00860784
R645 IND.n120 IND.n119 0.00860784
R646 IND.n124 IND.n123 0.00860784
R647 IND.n129 IND.n128 0.00860784
R648 IND.n133 IND.n132 0.00860784
R649 IND.n256 IND.n246 0.00860784
R650 IND.n147 IND.n146 0.00860784
R651 IND.n162 IND.n161 0.00860784
R652 IND.n182 IND.n181 0.00860784
R653 IND.n186 IND.n185 0.00860784
R654 IND.n191 IND.n190 0.00860784
R655 IND.n203 IND.n194 0.00860784
R656 IND.n228 IND.n220 0.00860784
R657 IND.n452 IND.n442 0.00860784
R658 IND.n27 IND.n26 0.00858096
R659 IND.n26 IND.n25 0.00858096
R660 IND.n415 IND.n414 0.00858096
R661 IND.n416 IND.n415 0.00858096
R662 IND.n48 IND.n47 0.00858096
R663 IND.n40 IND.n39 0.00858096
R664 IND.n49 IND.n48 0.00858096
R665 IND.n47 IND.n40 0.00858096
R666 IND.n353 IND.n352 0.00858096
R667 IND.n342 IND.n341 0.00858096
R668 IND.n339 IND.n338 0.00858096
R669 IND.n327 IND.n326 0.00858096
R670 IND.n354 IND.n353 0.00858096
R671 IND.n352 IND.n342 0.00858096
R672 IND.n340 IND.n339 0.00858096
R673 IND.n338 IND.n327 0.00858096
R674 IND.n71 IND.n70 0.00858096
R675 IND.n305 IND.n304 0.00858096
R676 IND.n306 IND.n305 0.00858096
R677 IND.n280 IND.n279 0.00858096
R678 IND.n272 IND.n271 0.00858096
R679 IND.n281 IND.n280 0.00858096
R680 IND.n279 IND.n272 0.00858096
R681 IND.n118 IND.n117 0.00858096
R682 IND.n127 IND.n126 0.00858096
R683 IND.n128 IND.n127 0.00858096
R684 IND.n119 IND.n118 0.00858096
R685 IND.n164 IND.n163 0.00858096
R686 IND.n158 IND.n157 0.00858096
R687 IND.n150 IND.n149 0.00858096
R688 IND.n163 IND.n162 0.00858096
R689 IND.n159 IND.n158 0.00858096
R690 IND.n157 IND.n150 0.00858096
R691 IND.n189 IND.n188 0.00858096
R692 IND.n190 IND.n189 0.00858096
R693 IND.n181 IND.n180 0.00858096
R694 IND.n24 IND.n23 0.00855417
R695 IND.n22 IND.n21 0.00855417
R696 IND.n18 IND.n17 0.00855417
R697 IND.n418 IND.n417 0.00855417
R698 IND.n38 IND.n37 0.00855417
R699 IND.n385 IND.n384 0.00855417
R700 IND.n325 IND.n324 0.00855417
R701 IND.n73 IND.n72 0.00855417
R702 IND.n75 IND.n74 0.00855417
R703 IND.n308 IND.n307 0.00855417
R704 IND.n310 IND.n309 0.00855417
R705 IND.n270 IND.n269 0.00855417
R706 IND.n121 IND.n120 0.00855417
R707 IND.n123 IND.n122 0.00855417
R708 IND.n130 IND.n129 0.00855417
R709 IND.n132 IND.n131 0.00855417
R710 IND.n246 IND.n245 0.00855417
R711 IND.n161 IND.n160 0.00855417
R712 IND.n148 IND.n147 0.00855417
R713 IND.n183 IND.n182 0.00855417
R714 IND.n185 IND.n184 0.00855417
R715 IND.n192 IND.n191 0.00855417
R716 IND.n194 IND.n193 0.00855417
R717 IND.n220 IND.n219 0.00855417
R718 IND.n442 IND.n441 0.00855417
R719 IND.n473 IND.n426 0.00773989
R720 IND.n424 IND.n423 0.00773989
R721 IND.n466 IND.n465 0.00773989
R722 IND.n467 IND.n466 0.00773989
R723 IND.n469 IND.n468 0.00773989
R724 IND.n425 IND.n424 0.00773989
R725 IND.n470 IND.n469 0.00773989
R726 IND.n433 IND.n432 0.00642105
R727 IND.n445 IND.n444 0.00642105
R728 IND.n458 IND.n457 0.00642105
R729 IND.n209 IND.n208 0.006097
R730 IND.n394 IND.n393 0.00605114
R731 IND.n369 IND.n368 0.00605114
R732 IND.n257 IND.n256 0.00605114
R733 IND.n229 IND.n228 0.00605114
R734 IND.n204 IND.n203 0.00605114
R735 IND.n453 IND.n452 0.00605114
R736 IND.n472 IND.n467 0.00582347
R737 IND.n374 IND.n373 0.00570918
R738 IND.n235 IND.n234 0.00570918
R739 IND.n457 IND.n456 0.00551512
R740 IND.n432 IND.n431 0.00551512
R741 IND.n362 IND.n361 0.00523684
R742 IND.n375 IND.n374 0.00523684
R743 IND.n388 IND.n387 0.00523684
R744 IND.n236 IND.n235 0.00523684
R745 IND.n249 IND.n248 0.00523684
R746 IND.n382 IND.n372 0.00479588
R747 IND.n243 IND.n233 0.00479588
R748 IND.n217 IND.n207 0.00479588
R749 IND.n16 IND.n15 0.00364318
R750 IND.n197 IND.n196 0.00286842
R751 IND.n210 IND.n209 0.00286842
R752 IND.n223 IND.n222 0.00286842
R753 VSS.t460 VSS.t535 122.014
R754 VSS.t415 VSS.t546 122.014
R755 VSS.t472 VSS.t495 122.014
R756 VSS.t513 VSS.t400 122.014
R757 VSS.t560 VSS.t474 122.014
R758 VSS.t418 VSS.t488 122.014
R759 VSS.t444 VSS.t424 122.014
R760 VSS.t479 VSS.t554 122.014
R761 VSS.t429 VSS.t458 122.014
R762 VSS.t470 VSS.t544 122.014
R763 VSS.t468 VSS.t406 122.014
R764 VSS.t509 VSS.t595 122.014
R765 VSS.t427 VSS.t587 112.368
R766 VSS.t558 VSS.t427 112.368
R767 VSS.t403 VSS.t558 112.368
R768 VSS.t437 VSS.t403 112.368
R769 VSS.t566 VSS.t437 112.368
R770 VSS.t533 VSS.t566 112.368
R771 VSS.t439 VSS.t593 112.368
R772 VSS.t564 VSS.t439 112.368
R773 VSS.t412 VSS.t564 112.368
R774 VSS.t448 VSS.t412 112.368
R775 VSS.t570 VSS.t448 112.368
R776 VSS.t537 VSS.t570 112.368
R777 VSS.t568 VSS.t409 112.368
R778 VSS.t490 VSS.t568 112.368
R779 VSS.t511 VSS.t531 112.368
R780 VSS.t432 VSS.t511 112.368
R781 VSS.t519 VSS.t505 69.8719
R782 VSS.t550 VSS.t519 69.8719
R783 VSS.t476 VSS.t550 69.8719
R784 VSS.t501 VSS.t579 69.8719
R785 VSS.t542 VSS.t526 69.8719
R786 VSS.t572 VSS.t542 69.8719
R787 VSS.t492 VSS.t572 69.8719
R788 VSS.t515 VSS.t597 69.8719
R789 VSS.n690 VSS.t562 59.9648
R790 VSS.n690 VSS.t460 59.9648
R791 VSS.n1651 VSS.t415 59.9648
R792 VSS.n1651 VSS.t574 59.9648
R793 VSS.n680 VSS.t446 59.9648
R794 VSS.n1557 VSS.t503 59.9648
R795 VSS.n1557 VSS.t472 59.9648
R796 VSS.n680 VSS.t513 59.9648
R797 VSS.n423 VSS.t524 59.9648
R798 VSS.n1521 VSS.t556 59.9648
R799 VSS.n1521 VSS.t560 59.9648
R800 VSS.n423 VSS.t418 59.9648
R801 VSS.n413 VSS.t589 59.9648
R802 VSS.n1425 VSS.t497 59.9648
R803 VSS.n1425 VSS.t444 59.9648
R804 VSS.n413 VSS.t479 59.9648
R805 VSS.n156 VSS.t583 59.9648
R806 VSS.n1389 VSS.t484 59.9648
R807 VSS.n1389 VSS.t429 59.9648
R808 VSS.n156 VSS.t470 59.9648
R809 VSS.n146 VSS.t435 59.9648
R810 VSS.n1293 VSS.t581 59.9648
R811 VSS.n1293 VSS.t468 59.9648
R812 VSS.n146 VSS.t509 59.9648
R813 VSS.n3786 VSS.t533 55.1416
R814 VSS.n3786 VSS.t462 55.1416
R815 VSS.n3426 VSS.t537 55.1416
R816 VSS.n3426 VSS.t499 55.1416
R817 VSS.n2245 VSS.t490 55.1416
R818 VSS.n2245 VSS.t450 55.1416
R819 VSS.n2375 VSS.t432 55.1416
R820 VSS.n2375 VSS.t585 55.1416
R821 VSS.n3543 VSS.t539 40.5416
R822 VSS.n2418 VSS.t452 40.5416
R823 VSS.n3543 VSS.t548 40.4112
R824 VSS.n2413 VSS.t528 36.5005
R825 VSS.n3480 VSS.t476 33.8934
R826 VSS.n3480 VSS.t501 33.8934
R827 VSS.n3269 VSS.t492 33.8434
R828 VSS.n3269 VSS.t515 33.8434
R829 VSS.n2044 VSS.n2023 27.2315
R830 VSS.n3113 VSS.t62 21.0957
R831 VSS.n2485 VSS.t453 21.0957
R832 VSS.n3306 VSS.t205 21.0957
R833 VSS.n3652 VSS.t540 21.0957
R834 VSS.n2417 VSS.n2416 20.8576
R835 VSS.n2416 VSS.n2415 20.8576
R836 VSS.n2415 VSS.n2414 20.8576
R837 VSS.n2414 VSS.n2413 20.8576
R838 VSS.t464 VSS.t517 19.5645
R839 VSS.t486 VSS.t441 19.5645
R840 VSS.t455 VSS.t591 19.5645
R841 VSS.n3288 VSS.t332 19.3003
R842 VSS.n3282 VSS.t386 19.3003
R843 VSS.n3761 VSS.t59 19.3003
R844 VSS.n3297 VSS.t599 18.8515
R845 VSS.n3076 VSS.t349 18.4027
R846 VSS.n3151 VSS.t636 18.4027
R847 VSS.n3376 VSS.n3375 18.022
R848 VSS.n3037 VSS.n3036 17.9538
R849 VSS.t529 VSS.t610 17.9538
R850 VSS.n3502 VSS.t264 17.505
R851 VSS.n2418 VSS.n2417 17.4684
R852 VSS.n2501 VSS.t482 16.6073
R853 VSS.n4032 VSS.t197 16.1048
R854 VSS.n4012 VSS.t175 16.1048
R855 VSS.n3537 VSS.t255 15.7097
R856 VSS.n2417 VSS.t466 15.6434
R857 VSS.n2413 VSS.t576 15.6434
R858 VSS.n2414 VSS.t481 15.6434
R859 VSS.n2415 VSS.t521 15.6434
R860 VSS.n2416 VSS.t421 15.6434
R861 VSS.n2401 VSS.t388 14.9545
R862 VSS.n3347 VSS.t391 14.9545
R863 VSS.n3306 VSS.t684 14.812
R864 VSS.n3303 VSS.t399 14.812
R865 VSS.t229 VSS.t4 14.812
R866 VSS.t235 VSS.t352 14.812
R867 VSS.n3511 VSS.t53 14.812
R868 VSS.n3520 VSS.t662 14.812
R869 VSS.n3282 VSS.t3 14.3632
R870 VSS.n3088 VSS.t344 13.9143
R871 VSS.n3165 VSS.t46 13.9143
R872 VSS.n3316 VSS.t389 13.9143
R873 VSS.n3540 VSS.t695 13.9143
R874 VSS.n890 VSS.t91 13.78
R875 VSS.n908 VSS.t24 13.78
R876 VSS.n1051 VSS.t89 13.78
R877 VSS.n1069 VSS.t10 13.78
R878 VSS.n1212 VSS.t79 13.78
R879 VSS.n1230 VSS.t98 13.78
R880 VSS.n2571 VSS.t486 13.542
R881 VSS.n2573 VSS.t552 13.542
R882 VSS.n2551 VSS.t455 13.542
R883 VSS.n2553 VSS.t507 13.542
R884 VSS.n2504 VSS.t577 13.0167
R885 VSS.n3285 VSS.t281 13.0167
R886 VSS.n3164 VSS.t464 12.7007
R887 VSS.n3335 VSS.t384 12.6539
R888 VSS.n3338 VSS.t385 12.6539
R889 VSS.t56 VSS.t615 12.5678
R890 VSS.n3047 VSS.t442 11.2213
R891 VSS.n3123 VSS.t624 11.2213
R892 VSS.n3179 VSS.t456 11.2213
R893 VSS.n3665 VSS.t616 11.2213
R894 VSS.n3294 VSS.t142 10.7725
R895 VSS.n3320 VSS.t331 10.3237
R896 VSS.n3291 VSS.t600 10.3237
R897 VSS.n3499 VSS.t680 10.3237
R898 VSS.n3534 VSS.t51 10.3237
R899 VSS.n3505 VSS.t5 9.87483
R900 VSS.n3524 VSS.t226 9.42599
R901 VSS.n4035 VSS.t192 9.20295
R902 VSS.n4009 VSS.t162 9.20295
R903 VSS.n3425 VSS.n3424 9.13939
R904 VSS.n4066 VSS.n3425 9.13939
R905 VSS.n2370 VSS.t433 8.81952
R906 VSS.n3372 VSS.t410 8.81952
R907 VSS.n3066 VSS.t342 8.52833
R908 VSS.n3142 VSS.t620 8.52833
R909 VSS.n2489 VSS.t422 8.52833
R910 VSS.n2501 VSS.t613 8.52833
R911 VSS.n3300 VSS.t180 8.52833
R912 VSS.n887 VSS.t114 7.87452
R913 VSS.n911 VSS.t71 7.87452
R914 VSS.n1048 VSS.t33 7.87452
R915 VSS.n1072 VSS.t68 7.87452
R916 VSS.n1209 VSS.t40 7.87452
R917 VSS.n1233 VSS.t103 7.87452
R918 VSS.n3514 VSS.t167 7.63066
R919 VSS.n3514 VSS.t141 7.18183
R920 VSS.t398 VSS.t493 6.733
R921 VSS.n3668 VSS.t49 6.733
R922 VSS.n2386 VSS.t2 6.5189
R923 VSS.n3362 VSS.t392 6.5189
R924 VSS.n3303 VSS.t353 6.28416
R925 VSS.n3479 VSS.t580 5.8372
R926 VSS.n3268 VSS.t598 5.8372
R927 VSS.n3662 VSS.t56 5.83533
R928 VSS.t662 VSS.t273 5.3865
R929 VSS.n4025 VSS.t221 5.3686
R930 VSS.n4019 VSS.t209 5.3686
R931 VSS VSS.n3425 5.2005
R932 VSS VSS.n3425 5.2005
R933 VSS.n2443 VSS.t390 5.07024
R934 VSS.n2902 VSS.t518 5.0182
R935 VSS.n3508 VSS.t235 4.93766
R936 VSS.n3546 VSS.t541 4.7885
R937 VSS.n3592 VSS.t549 4.7885
R938 VSS.n2743 VSS.t467 4.7885
R939 VSS.n3479 VSS.t502 4.7885
R940 VSS.n3483 VSS.t478 4.7885
R941 VSS.n3484 VSS.t551 4.7885
R942 VSS.n3485 VSS.t520 4.7885
R943 VSS.n3486 VSS.t506 4.7885
R944 VSS.n3275 VSS.t527 4.7885
R945 VSS.n3274 VSS.t543 4.7885
R946 VSS.n3273 VSS.t573 4.7885
R947 VSS.n3272 VSS.t494 4.7885
R948 VSS.n3268 VSS.t516 4.7885
R949 VSS.n2907 VSS.n2906 4.78615
R950 VSS.n896 VSS.t28 4.59368
R951 VSS.n902 VSS.t112 4.59368
R952 VSS.n1057 VSS.t19 4.59368
R953 VSS.n1063 VSS.t313 4.59368
R954 VSS.n1218 VSS.t16 4.59368
R955 VSS.n1224 VSS.t83 4.59368
R956 VSS.n2640 VSS.n2570 4.45746
R957 VSS.n2655 VSS.n2568 4.45746
R958 VSS.n1576 VSS.n1575 4.44992
R959 VSS.n1596 VSS.n1595 4.44992
R960 VSS.n1444 VSS.n1443 4.44992
R961 VSS.n1464 VSS.n1463 4.44992
R962 VSS.n1312 VSS.n1311 4.44992
R963 VSS.n1332 VSS.n1331 4.44992
R964 VSS.n2395 VSS.t0 4.21829
R965 VSS.n3353 VSS.t1 4.21829
R966 VSS.n2925 VSS.n2924 4.1992
R967 VSS.n2930 VSS.n2929 4.1992
R968 VSS.n2437 VSS.n2436 4.05833
R969 VSS.n3098 VSS.t339 4.04
R970 VSS.n2495 VSS.t522 4.04
R971 VSS.n3294 VSS.t247 4.04
R972 VSS.n2246 VSS.n2245 4.0005
R973 VSS.n681 VSS.n680 4.0005
R974 VSS.n1558 VSS.n1557 4.0005
R975 VSS.n424 VSS.n423 4.0005
R976 VSS.n1522 VSS.n1521 4.0005
R977 VSS.n414 VSS.n413 4.0005
R978 VSS.n1426 VSS.n1425 4.0005
R979 VSS.n157 VSS.n156 4.0005
R980 VSS.n1390 VSS.n1389 4.0005
R981 VSS.n147 VSS.n146 4.0005
R982 VSS.n1294 VSS.n1293 4.0005
R983 VSS.n1652 VSS.n1651 4.0005
R984 VSS.n691 VSS.n690 4.0005
R985 VSS.n2419 VSS.n2418 4.0005
R986 VSS.n3544 VSS.n3543 4.0005
R987 VSS.n3481 VSS.n3480 4.0005
R988 VSS.n3270 VSS.n3269 4.0005
R989 VSS.n2376 VSS.n2375 4.0005
R990 VSS.n3427 VSS.n3426 4.0005
R991 VSS.n3787 VSS.n3786 4.0005
R992 VSS.n2902 VSS.t465 3.9695
R993 VSS.n2558 VSS.t508 3.9695
R994 VSS.n2898 VSS.t457 3.9695
R995 VSS.n2899 VSS.t592 3.9695
R996 VSS.n2820 VSS.n2746 3.75898
R997 VSS.n2817 VSS.n2747 3.75898
R998 VSS.n2812 VSS.n2748 3.75898
R999 VSS.n2807 VSS.n2749 3.75898
R1000 VSS.n2771 VSS.n2751 3.75898
R1001 VSS.n2760 VSS.n2753 3.75898
R1002 VSS.n3558 VSS.n3555 3.75898
R1003 VSS.n3569 VSS.n3553 3.75898
R1004 VSS.n3578 VSS.n3551 3.75898
R1005 VSS.n3789 VSS.t463 3.71925
R1006 VSS.n3785 VSS.t534 3.71925
R1007 VSS.n3784 VSS.t567 3.71925
R1008 VSS.n3783 VSS.t438 3.71925
R1009 VSS.n3782 VSS.t405 3.71925
R1010 VSS.n68 VSS.t559 3.71925
R1011 VSS.n69 VSS.t428 3.71925
R1012 VSS.n70 VSS.t588 3.71925
R1013 VSS.n3431 VSS.t538 3.71925
R1014 VSS.n3430 VSS.t571 3.71925
R1015 VSS.n3429 VSS.t449 3.71925
R1016 VSS.n3428 VSS.t414 3.71925
R1017 VSS.n5 VSS.t565 3.71925
R1018 VSS.n6 VSS.t440 3.71925
R1019 VSS.n7 VSS.t594 3.71925
R1020 VSS.n3433 VSS.t500 3.71925
R1021 VSS.n2248 VSS.t451 3.71925
R1022 VSS.n2244 VSS.t491 3.71925
R1023 VSS.n2243 VSS.t569 3.71925
R1024 VSS.n2089 VSS.t411 3.71925
R1025 VSS.n2378 VSS.t586 3.71925
R1026 VSS.n2374 VSS.t434 3.71925
R1027 VSS.n2373 VSS.t512 3.71925
R1028 VSS.n2091 VSS.t532 3.71925
R1029 VSS.n689 VSS.t461 3.6965
R1030 VSS.n688 VSS.t536 3.6965
R1031 VSS.n1653 VSS.t547 3.6965
R1032 VSS.n1654 VSS.t417 3.6965
R1033 VSS.n1656 VSS.t575 3.6965
R1034 VSS.n1560 VSS.t504 3.6965
R1035 VSS.n679 VSS.t514 3.6965
R1036 VSS.n678 VSS.t402 3.6965
R1037 VSS.n1555 VSS.t496 3.6965
R1038 VSS.n1556 VSS.t473 3.6965
R1039 VSS.n683 VSS.t447 3.6965
R1040 VSS.n1524 VSS.t557 3.6965
R1041 VSS.n422 VSS.t420 3.6965
R1042 VSS.n421 VSS.t489 3.6965
R1043 VSS.n1519 VSS.t475 3.6965
R1044 VSS.n1520 VSS.t561 3.6965
R1045 VSS.n426 VSS.t525 3.6965
R1046 VSS.n1428 VSS.t498 3.6965
R1047 VSS.n412 VSS.t480 3.6965
R1048 VSS.n411 VSS.t555 3.6965
R1049 VSS.n1423 VSS.t426 3.6965
R1050 VSS.n1424 VSS.t445 3.6965
R1051 VSS.n416 VSS.t590 3.6965
R1052 VSS.n1392 VSS.t485 3.6965
R1053 VSS.n155 VSS.t471 3.6965
R1054 VSS.n154 VSS.t545 3.6965
R1055 VSS.n1387 VSS.t459 3.6965
R1056 VSS.n1388 VSS.t431 3.6965
R1057 VSS.n159 VSS.t584 3.6965
R1058 VSS.n1296 VSS.t582 3.6965
R1059 VSS.n145 VSS.t510 3.6965
R1060 VSS.n144 VSS.t596 3.6965
R1061 VSS.n1291 VSS.t408 3.6965
R1062 VSS.n1292 VSS.t469 3.6965
R1063 VSS.n149 VSS.t436 3.6965
R1064 VSS.n693 VSS.t563 3.6965
R1065 VSS.n2444 VSS.n2422 3.43224
R1066 VSS.n2442 VSS.n2424 3.43224
R1067 VSS.n2441 VSS.n2426 3.43224
R1068 VSS.n2440 VSS.n2428 3.43224
R1069 VSS.n2439 VSS.n2430 3.43224
R1070 VSS.n2438 VSS.n2432 3.43224
R1071 VSS.n2437 VSS.n2434 3.43224
R1072 VSS.n2732 VSS.n2730 3.31707
R1073 VSS.n2046 VSS.n2022 3.3165
R1074 VSS.n2046 VSS.n2045 3.3165
R1075 VSS.n2471 VSS.n2470 3.3165
R1076 VSS.n2547 VSS.n2544 3.3164
R1077 VSS.n2868 VSS.n2866 3.3164
R1078 VSS.n2865 VSS.n2864 3.3164
R1079 VSS.n2547 VSS.n2546 3.31583
R1080 VSS.n2868 VSS.n2867 3.31583
R1081 VSS.n19 VSS.n12 3.1505
R1082 VSS.n18 VSS.n14 3.1505
R1083 VSS.n17 VSS.n16 3.1505
R1084 VSS.n3436 VSS.n3435 3.1505
R1085 VSS.n3439 VSS.n3438 3.1505
R1086 VSS.n3442 VSS.n3441 3.1505
R1087 VSS.n3445 VSS.n3444 3.1505
R1088 VSS.n3448 VSS.n3447 3.1505
R1089 VSS.n28 VSS.n21 3.1505
R1090 VSS.n27 VSS.n23 3.1505
R1091 VSS.n26 VSS.n25 3.1505
R1092 VSS.n3451 VSS.n3450 3.1505
R1093 VSS.n3454 VSS.n3453 3.1505
R1094 VSS.n3457 VSS.n3456 3.1505
R1095 VSS.n3460 VSS.n3459 3.1505
R1096 VSS.n3463 VSS.n3462 3.1505
R1097 VSS.n37 VSS.n30 3.1505
R1098 VSS.n36 VSS.n32 3.1505
R1099 VSS.n35 VSS.n34 3.1505
R1100 VSS.n3466 VSS.n3465 3.1505
R1101 VSS.n3469 VSS.n3468 3.1505
R1102 VSS.n3472 VSS.n3471 3.1505
R1103 VSS.n3475 VSS.n3474 3.1505
R1104 VSS.n3478 VSS.n3477 3.1505
R1105 VSS.n2907 VSS.n2904 3.1505
R1106 VSS.n2908 VSS.n2903 3.1505
R1107 VSS.n2925 VSS.n2922 3.1505
R1108 VSS.n2930 VSS.n2927 3.1505
R1109 VSS.n1629 VSS.n1628 3.1505
R1110 VSS.n1630 VSS.n1624 3.1505
R1111 VSS.n1497 VSS.n1496 3.1505
R1112 VSS.n1498 VSS.n1492 3.1505
R1113 VSS.n1365 VSS.n1364 3.1505
R1114 VSS.n1366 VSS.n1360 3.1505
R1115 VSS.n2936 VSS.n2932 3.1505
R1116 VSS.n2935 VSS.n2934 3.1505
R1117 VSS.n2580 VSS.n2579 3.1505
R1118 VSS.n2920 VSS.n2916 3.1505
R1119 VSS.n2919 VSS.n2918 3.1505
R1120 VSS.n2566 VSS.n2565 3.1505
R1121 VSS.n2914 VSS.n2910 3.1505
R1122 VSS.n2913 VSS.n2912 3.1505
R1123 VSS.n2563 VSS.n2562 3.1505
R1124 VSS.n2446 VSS.n2412 3.1505
R1125 VSS.n2745 VSS.n2744 3.1505
R1126 VSS.n46 VSS.n39 3.1505
R1127 VSS.n45 VSS.n41 3.1505
R1128 VSS.n44 VSS.n43 3.1505
R1129 VSS.n3769 VSS.n3768 3.1505
R1130 VSS.n3772 VSS.n3771 3.1505
R1131 VSS.n3775 VSS.n3774 3.1505
R1132 VSS.n3778 VSS.n3777 3.1505
R1133 VSS.n3781 VSS.n3780 3.1505
R1134 VSS.n3531 VSS.t294 3.14233
R1135 VSS.n3216 VSS.n3214 3.06136
R1136 VSS.n1170 VSS.n1169 3.01258
R1137 VSS.n1009 VSS.n1008 3.01258
R1138 VSS.n848 VSS.n847 3.01258
R1139 VSS.n2732 VSS.n2731 3.01202
R1140 VSS.n2742 VSS.n2741 3.01202
R1141 VSS.n2471 VSS.n2469 3.0115
R1142 VSS.n1569 VSS.n1566 2.91104
R1143 VSS.n1589 VSS.n1586 2.91104
R1144 VSS.n1437 VSS.n1434 2.91104
R1145 VSS.n1457 VSS.n1454 2.91104
R1146 VSS.n1305 VSS.n1302 2.91104
R1147 VSS.n1325 VSS.n1322 2.91104
R1148 VSS.n1581 VSS.n1578 2.86846
R1149 VSS.n1601 VSS.n1598 2.86846
R1150 VSS.n1449 VSS.n1446 2.86846
R1151 VSS.n1469 VSS.n1466 2.86846
R1152 VSS.n1317 VSS.n1314 2.86846
R1153 VSS.n1337 VSS.n1334 2.86846
R1154 VSS.n1634 VSS.n1633 2.80979
R1155 VSS.n1502 VSS.n1501 2.80979
R1156 VSS.n1370 VSS.n1369 2.80979
R1157 VSS.n976 VSS.n975 2.80714
R1158 VSS.n1137 VSS.n1136 2.80714
R1159 VSS.n1272 VSS.n1271 2.80714
R1160 VSS.n2522 VSS.n2521 2.80714
R1161 VSS.n2522 VSS.n2520 2.80651
R1162 VSS.n3018 VSS.n3017 2.74966
R1163 VSS.n3499 VSS.t140 2.6935
R1164 VSS.n2575 VSS.n2573 2.65431
R1165 VSS.n2555 VSS.n2553 2.65431
R1166 VSS.n3602 VSS.n3601 2.6005
R1167 VSS.n3637 VSS.n3636 2.6005
R1168 VSS.n3635 VSS.n3634 2.6005
R1169 VSS.n3632 VSS.n3631 2.6005
R1170 VSS.n3630 VSS.n3629 2.6005
R1171 VSS.n3627 VSS.n3626 2.6005
R1172 VSS.n3625 VSS.n3624 2.6005
R1173 VSS.n3622 VSS.n3621 2.6005
R1174 VSS.n3620 VSS.n3619 2.6005
R1175 VSS.n3617 VSS.n3616 2.6005
R1176 VSS.n3615 VSS.n3614 2.6005
R1177 VSS.n3612 VSS.n3611 2.6005
R1178 VSS.n3610 VSS.n3609 2.6005
R1179 VSS.n3607 VSS.n3606 2.6005
R1180 VSS.n3605 VSS.n3604 2.6005
R1181 VSS.n2465 VSS.n2464 2.6005
R1182 VSS.n2897 VSS.n2896 2.6005
R1183 VSS.n2881 VSS.n2880 2.6005
R1184 VSS.n2883 VSS.n2882 2.6005
R1185 VSS.n2886 VSS.n2885 2.6005
R1186 VSS.n2889 VSS.n2888 2.6005
R1187 VSS.n2892 VSS.n2891 2.6005
R1188 VSS.n2895 VSS.n2894 2.6005
R1189 VSS.n2463 VSS.n2462 2.6005
R1190 VSS.n2460 VSS.n2459 2.6005
R1191 VSS.n2458 VSS.n2457 2.6005
R1192 VSS.n2455 VSS.n2454 2.6005
R1193 VSS.n2453 VSS.n2452 2.6005
R1194 VSS.n2450 VSS.n2449 2.6005
R1195 VSS.n2448 VSS.n2447 2.6005
R1196 VSS.n2734 VSS.n2733 2.6005
R1197 VSS.n2736 VSS.n2735 2.6005
R1198 VSS.n2739 VSS.n2738 2.6005
R1199 VSS.n2260 VSS.n2259 2.6005
R1200 VSS.n3807 VSS.n3806 2.6005
R1201 VSS.n3809 VSS.n3808 2.6005
R1202 VSS.n3811 VSS.n3810 2.6005
R1203 VSS.n3813 VSS.n3812 2.6005
R1204 VSS.n3815 VSS.n3814 2.6005
R1205 VSS.n3817 VSS.n3816 2.6005
R1206 VSS.n3819 VSS.n3818 2.6005
R1207 VSS.n3821 VSS.n3820 2.6005
R1208 VSS.n3823 VSS.n3822 2.6005
R1209 VSS.n3825 VSS.n3824 2.6005
R1210 VSS.n3827 VSS.n3826 2.6005
R1211 VSS.n3829 VSS.n3828 2.6005
R1212 VSS.n3831 VSS.n3830 2.6005
R1213 VSS.n3833 VSS.n3832 2.6005
R1214 VSS.n3835 VSS.n3834 2.6005
R1215 VSS.n3837 VSS.n3836 2.6005
R1216 VSS.n3839 VSS.n3838 2.6005
R1217 VSS.n3841 VSS.n3840 2.6005
R1218 VSS.n3843 VSS.n3842 2.6005
R1219 VSS.n3845 VSS.n3844 2.6005
R1220 VSS.n3847 VSS.n3846 2.6005
R1221 VSS.n3849 VSS.n3848 2.6005
R1222 VSS.n3851 VSS.n3850 2.6005
R1223 VSS.n3853 VSS.n3852 2.6005
R1224 VSS.n3855 VSS.n3854 2.6005
R1225 VSS.n3857 VSS.n3856 2.6005
R1226 VSS.n3859 VSS.n3858 2.6005
R1227 VSS.n3861 VSS.n3860 2.6005
R1228 VSS.n3863 VSS.n3862 2.6005
R1229 VSS.n3865 VSS.n3864 2.6005
R1230 VSS.n3867 VSS.n3866 2.6005
R1231 VSS.n3869 VSS.n3868 2.6005
R1232 VSS.n3871 VSS.n3870 2.6005
R1233 VSS.n3873 VSS.n3872 2.6005
R1234 VSS.n3875 VSS.n3874 2.6005
R1235 VSS.n3877 VSS.n3876 2.6005
R1236 VSS.n3879 VSS.n3878 2.6005
R1237 VSS.n3881 VSS.n3880 2.6005
R1238 VSS.n3883 VSS.n3882 2.6005
R1239 VSS.n3885 VSS.n3884 2.6005
R1240 VSS.n3887 VSS.n3886 2.6005
R1241 VSS.n3889 VSS.n3888 2.6005
R1242 VSS.n3891 VSS.n3890 2.6005
R1243 VSS.n3893 VSS.n3892 2.6005
R1244 VSS.n3896 VSS.n3895 2.6005
R1245 VSS.n3898 VSS.n3897 2.6005
R1246 VSS.n3901 VSS.n3900 2.6005
R1247 VSS.n3903 VSS.n3902 2.6005
R1248 VSS.n3906 VSS.n3905 2.6005
R1249 VSS.n3908 VSS.n3907 2.6005
R1250 VSS.n3911 VSS.n3910 2.6005
R1251 VSS.n3913 VSS.n3912 2.6005
R1252 VSS.n3916 VSS.n3915 2.6005
R1253 VSS.n3918 VSS.n3917 2.6005
R1254 VSS.n3921 VSS.n3920 2.6005
R1255 VSS.n3923 VSS.n3922 2.6005
R1256 VSS.n3980 VSS.n3979 2.6005
R1257 VSS.n2262 VSS.n2261 2.6005
R1258 VSS.n2264 VSS.n2263 2.6005
R1259 VSS.n2266 VSS.n2265 2.6005
R1260 VSS.n2268 VSS.n2267 2.6005
R1261 VSS.n2270 VSS.n2269 2.6005
R1262 VSS.n2272 VSS.n2271 2.6005
R1263 VSS.n2274 VSS.n2273 2.6005
R1264 VSS.n2276 VSS.n2275 2.6005
R1265 VSS.n2278 VSS.n2277 2.6005
R1266 VSS.n2280 VSS.n2279 2.6005
R1267 VSS.n2282 VSS.n2281 2.6005
R1268 VSS.n2284 VSS.n2283 2.6005
R1269 VSS.n2286 VSS.n2285 2.6005
R1270 VSS.n2288 VSS.n2287 2.6005
R1271 VSS.n2290 VSS.n2289 2.6005
R1272 VSS.n2292 VSS.n2291 2.6005
R1273 VSS.n2294 VSS.n2293 2.6005
R1274 VSS.n2296 VSS.n2295 2.6005
R1275 VSS.n2298 VSS.n2297 2.6005
R1276 VSS.n2300 VSS.n2299 2.6005
R1277 VSS.n2302 VSS.n2301 2.6005
R1278 VSS.n2304 VSS.n2303 2.6005
R1279 VSS.n2306 VSS.n2305 2.6005
R1280 VSS.n2308 VSS.n2307 2.6005
R1281 VSS.n2310 VSS.n2309 2.6005
R1282 VSS.n2312 VSS.n2311 2.6005
R1283 VSS.n2314 VSS.n2313 2.6005
R1284 VSS.n2316 VSS.n2315 2.6005
R1285 VSS.n2318 VSS.n2317 2.6005
R1286 VSS.n2321 VSS.n2320 2.6005
R1287 VSS.n2323 VSS.n2322 2.6005
R1288 VSS.n2326 VSS.n2325 2.6005
R1289 VSS.n2328 VSS.n2327 2.6005
R1290 VSS.n2331 VSS.n2330 2.6005
R1291 VSS.n2333 VSS.n2332 2.6005
R1292 VSS.n2336 VSS.n2335 2.6005
R1293 VSS.n2338 VSS.n2337 2.6005
R1294 VSS.n2341 VSS.n2340 2.6005
R1295 VSS.n2343 VSS.n2342 2.6005
R1296 VSS.n126 VSS.n125 2.6005
R1297 VSS.n143 VSS.n142 2.6005
R1298 VSS.n137 VSS.n136 2.6005
R1299 VSS.n139 VSS.n138 2.6005
R1300 VSS.n141 VSS.n140 2.6005
R1301 VSS.n135 VSS.n134 2.6005
R1302 VSS.n2088 VSS.n2087 2.6005
R1303 VSS.n2060 VSS.n2059 2.6005
R1304 VSS.n2062 VSS.n2061 2.6005
R1305 VSS.n2064 VSS.n2063 2.6005
R1306 VSS.n2066 VSS.n2065 2.6005
R1307 VSS.n2068 VSS.n2067 2.6005
R1308 VSS.n2070 VSS.n2069 2.6005
R1309 VSS.n2072 VSS.n2071 2.6005
R1310 VSS.n2074 VSS.n2073 2.6005
R1311 VSS.n2076 VSS.n2075 2.6005
R1312 VSS.n2078 VSS.n2077 2.6005
R1313 VSS.n2080 VSS.n2079 2.6005
R1314 VSS.n2082 VSS.n2081 2.6005
R1315 VSS.n2084 VSS.n2083 2.6005
R1316 VSS.n2086 VSS.n2085 2.6005
R1317 VSS.n2058 VSS.n2057 2.6005
R1318 VSS.n2055 VSS.n2052 2.6005
R1319 VSS.n2055 VSS.n2054 2.6005
R1320 VSS.n132 VSS.n131 2.6005
R1321 VSS.n1900 VSS.n1899 2.6005
R1322 VSS.n1900 VSS.n1897 2.6005
R1323 VSS.n1901 VSS.n1290 2.6005
R1324 VSS.n1282 VSS.n1281 2.6005
R1325 VSS.n1284 VSS.n1283 2.6005
R1326 VSS.n1287 VSS.n1286 2.6005
R1327 VSS.n1289 VSS.n1288 2.6005
R1328 VSS.n2048 VSS.n2047 2.6005
R1329 VSS.n2020 VSS.n2019 2.6005
R1330 VSS.n2017 VSS.n2016 2.6005
R1331 VSS.n2015 VSS.n2014 2.6005
R1332 VSS.n2012 VSS.n2011 2.6005
R1333 VSS.n2010 VSS.n2009 2.6005
R1334 VSS.n2007 VSS.n2006 2.6005
R1335 VSS.n2005 VSS.n2004 2.6005
R1336 VSS.n2002 VSS.n2001 2.6005
R1337 VSS.n2000 VSS.n1999 2.6005
R1338 VSS.n1997 VSS.n1996 2.6005
R1339 VSS.n1995 VSS.n1994 2.6005
R1340 VSS.n1992 VSS.n1991 2.6005
R1341 VSS.n1990 VSS.n1989 2.6005
R1342 VSS.n1987 VSS.n1986 2.6005
R1343 VSS.n1985 VSS.n1984 2.6005
R1344 VSS.n1982 VSS.n1981 2.6005
R1345 VSS.n1980 VSS.n1979 2.6005
R1346 VSS.n1977 VSS.n1976 2.6005
R1347 VSS.n1975 VSS.n1974 2.6005
R1348 VSS.n1973 VSS.n1972 2.6005
R1349 VSS.n1971 VSS.n1970 2.6005
R1350 VSS.n1969 VSS.n1968 2.6005
R1351 VSS.n1967 VSS.n1966 2.6005
R1352 VSS.n1965 VSS.n1964 2.6005
R1353 VSS.n1963 VSS.n1962 2.6005
R1354 VSS.n1961 VSS.n1960 2.6005
R1355 VSS.n1959 VSS.n1958 2.6005
R1356 VSS.n1957 VSS.n1956 2.6005
R1357 VSS.n1955 VSS.n1954 2.6005
R1358 VSS.n1953 VSS.n1952 2.6005
R1359 VSS.n1951 VSS.n1950 2.6005
R1360 VSS.n1949 VSS.n1948 2.6005
R1361 VSS.n1947 VSS.n1946 2.6005
R1362 VSS.n1945 VSS.n1944 2.6005
R1363 VSS.n1943 VSS.n1942 2.6005
R1364 VSS.n1941 VSS.n1940 2.6005
R1365 VSS.n1939 VSS.n1938 2.6005
R1366 VSS.n1937 VSS.n1936 2.6005
R1367 VSS.n1935 VSS.n1934 2.6005
R1368 VSS.n1933 VSS.n1932 2.6005
R1369 VSS.n1931 VSS.n1930 2.6005
R1370 VSS.n1929 VSS.n1928 2.6005
R1371 VSS.n1927 VSS.n1926 2.6005
R1372 VSS.n1925 VSS.n1924 2.6005
R1373 VSS.n1923 VSS.n1922 2.6005
R1374 VSS.n1921 VSS.n1920 2.6005
R1375 VSS.n1919 VSS.n1918 2.6005
R1376 VSS.n1917 VSS.n1916 2.6005
R1377 VSS.n1915 VSS.n1914 2.6005
R1378 VSS.n1913 VSS.n1912 2.6005
R1379 VSS.n1911 VSS.n1910 2.6005
R1380 VSS.n1909 VSS.n1908 2.6005
R1381 VSS.n1907 VSS.n1906 2.6005
R1382 VSS.n1905 VSS.n1904 2.6005
R1383 VSS.n1903 VSS.n1902 2.6005
R1384 VSS.n1279 VSS.n1278 2.6005
R1385 VSS.n1176 VSS.n1175 2.6005
R1386 VSS.n1175 VSS.n1174 2.6005
R1387 VSS.n1179 VSS.n1178 2.6005
R1388 VSS.n1178 VSS.n1177 2.6005
R1389 VSS.n1182 VSS.n1181 2.6005
R1390 VSS.n1181 VSS.n1180 2.6005
R1391 VSS.n1185 VSS.n1184 2.6005
R1392 VSS.n1184 VSS.n1183 2.6005
R1393 VSS.n1188 VSS.n1187 2.6005
R1394 VSS.n1187 VSS.n1186 2.6005
R1395 VSS.n1191 VSS.n1190 2.6005
R1396 VSS.n1190 VSS.n1189 2.6005
R1397 VSS.n1195 VSS.n1194 2.6005
R1398 VSS.n1194 VSS.n1193 2.6005
R1399 VSS.n1199 VSS.n1198 2.6005
R1400 VSS.n1198 VSS.n1197 2.6005
R1401 VSS.n1202 VSS.n1201 2.6005
R1402 VSS.n1201 VSS.n1200 2.6005
R1403 VSS.n1205 VSS.n1204 2.6005
R1404 VSS.n1204 VSS.n1203 2.6005
R1405 VSS.n1208 VSS.n1207 2.6005
R1406 VSS.n1207 VSS.n1206 2.6005
R1407 VSS.n1211 VSS.n1210 2.6005
R1408 VSS.n1210 VSS.n1209 2.6005
R1409 VSS.n1214 VSS.n1213 2.6005
R1410 VSS.n1213 VSS.n1212 2.6005
R1411 VSS.n1217 VSS.n1216 2.6005
R1412 VSS.n1216 VSS.n1215 2.6005
R1413 VSS.n1220 VSS.n1219 2.6005
R1414 VSS.n1219 VSS.n1218 2.6005
R1415 VSS.n1223 VSS.n1222 2.6005
R1416 VSS.n1222 VSS.n1221 2.6005
R1417 VSS.n1226 VSS.n1225 2.6005
R1418 VSS.n1225 VSS.n1224 2.6005
R1419 VSS.n1229 VSS.n1228 2.6005
R1420 VSS.n1228 VSS.n1227 2.6005
R1421 VSS.n1232 VSS.n1231 2.6005
R1422 VSS.n1231 VSS.n1230 2.6005
R1423 VSS.n1235 VSS.n1234 2.6005
R1424 VSS.n1234 VSS.n1233 2.6005
R1425 VSS.n1238 VSS.n1237 2.6005
R1426 VSS.n1237 VSS.n1236 2.6005
R1427 VSS.n1241 VSS.n1240 2.6005
R1428 VSS.n1240 VSS.n1239 2.6005
R1429 VSS.n1244 VSS.n1243 2.6005
R1430 VSS.n1243 VSS.n1242 2.6005
R1431 VSS.n1247 VSS.n1246 2.6005
R1432 VSS.n1246 VSS.n1245 2.6005
R1433 VSS.n1251 VSS.n1250 2.6005
R1434 VSS.n1250 VSS.n1249 2.6005
R1435 VSS.n1255 VSS.n1254 2.6005
R1436 VSS.n1254 VSS.n1253 2.6005
R1437 VSS.n1258 VSS.n1257 2.6005
R1438 VSS.n1257 VSS.n1256 2.6005
R1439 VSS.n1261 VSS.n1260 2.6005
R1440 VSS.n1260 VSS.n1259 2.6005
R1441 VSS.n1264 VSS.n1263 2.6005
R1442 VSS.n1263 VSS.n1262 2.6005
R1443 VSS.n1267 VSS.n1266 2.6005
R1444 VSS.n1266 VSS.n1265 2.6005
R1445 VSS.n1270 VSS.n1269 2.6005
R1446 VSS.n1269 VSS.n1268 2.6005
R1447 VSS.n1172 VSS.n1171 2.6005
R1448 VSS.n1406 VSS.n1405 2.6005
R1449 VSS.n1404 VSS.n1403 2.6005
R1450 VSS.n1402 VSS.n1401 2.6005
R1451 VSS.n1400 VSS.n1399 2.6005
R1452 VSS.n1398 VSS.n1397 2.6005
R1453 VSS.n165 VSS.n164 2.6005
R1454 VSS.n167 VSS.n166 2.6005
R1455 VSS.n169 VSS.n168 2.6005
R1456 VSS.n171 VSS.n170 2.6005
R1457 VSS.n173 VSS.n172 2.6005
R1458 VSS.n175 VSS.n174 2.6005
R1459 VSS.n177 VSS.n176 2.6005
R1460 VSS.n179 VSS.n178 2.6005
R1461 VSS.n181 VSS.n180 2.6005
R1462 VSS.n183 VSS.n182 2.6005
R1463 VSS.n185 VSS.n184 2.6005
R1464 VSS.n187 VSS.n186 2.6005
R1465 VSS.n189 VSS.n188 2.6005
R1466 VSS.n191 VSS.n190 2.6005
R1467 VSS.n193 VSS.n192 2.6005
R1468 VSS.n195 VSS.n194 2.6005
R1469 VSS.n197 VSS.n196 2.6005
R1470 VSS.n199 VSS.n198 2.6005
R1471 VSS.n201 VSS.n200 2.6005
R1472 VSS.n203 VSS.n202 2.6005
R1473 VSS.n205 VSS.n204 2.6005
R1474 VSS.n207 VSS.n206 2.6005
R1475 VSS.n209 VSS.n208 2.6005
R1476 VSS.n211 VSS.n210 2.6005
R1477 VSS.n213 VSS.n212 2.6005
R1478 VSS.n215 VSS.n214 2.6005
R1479 VSS.n217 VSS.n216 2.6005
R1480 VSS.n219 VSS.n218 2.6005
R1481 VSS.n221 VSS.n220 2.6005
R1482 VSS.n223 VSS.n222 2.6005
R1483 VSS.n225 VSS.n224 2.6005
R1484 VSS.n227 VSS.n226 2.6005
R1485 VSS.n229 VSS.n228 2.6005
R1486 VSS.n231 VSS.n230 2.6005
R1487 VSS.n233 VSS.n232 2.6005
R1488 VSS.n235 VSS.n234 2.6005
R1489 VSS.n237 VSS.n236 2.6005
R1490 VSS.n239 VSS.n238 2.6005
R1491 VSS.n241 VSS.n240 2.6005
R1492 VSS.n243 VSS.n242 2.6005
R1493 VSS.n245 VSS.n244 2.6005
R1494 VSS.n247 VSS.n246 2.6005
R1495 VSS.n249 VSS.n248 2.6005
R1496 VSS.n251 VSS.n250 2.6005
R1497 VSS.n253 VSS.n252 2.6005
R1498 VSS.n255 VSS.n254 2.6005
R1499 VSS.n258 VSS.n257 2.6005
R1500 VSS.n260 VSS.n259 2.6005
R1501 VSS.n263 VSS.n262 2.6005
R1502 VSS.n265 VSS.n264 2.6005
R1503 VSS.n268 VSS.n267 2.6005
R1504 VSS.n270 VSS.n269 2.6005
R1505 VSS.n273 VSS.n272 2.6005
R1506 VSS.n275 VSS.n274 2.6005
R1507 VSS.n278 VSS.n277 2.6005
R1508 VSS.n280 VSS.n279 2.6005
R1509 VSS.n283 VSS.n282 2.6005
R1510 VSS.n1408 VSS.n1407 2.6005
R1511 VSS.n1829 VSS.n1409 2.6005
R1512 VSS.n1828 VSS.n1826 2.6005
R1513 VSS.n1831 VSS.n1830 2.6005
R1514 VSS.n1833 VSS.n1832 2.6005
R1515 VSS.n1835 VSS.n1834 2.6005
R1516 VSS.n1837 VSS.n1836 2.6005
R1517 VSS.n1839 VSS.n1838 2.6005
R1518 VSS.n1841 VSS.n1840 2.6005
R1519 VSS.n1844 VSS.n1843 2.6005
R1520 VSS.n1847 VSS.n1846 2.6005
R1521 VSS.n1849 VSS.n1848 2.6005
R1522 VSS.n1851 VSS.n1850 2.6005
R1523 VSS.n1854 VSS.n1853 2.6005
R1524 VSS.n1856 VSS.n1855 2.6005
R1525 VSS.n1858 VSS.n1857 2.6005
R1526 VSS.n1860 VSS.n1859 2.6005
R1527 VSS.n1862 VSS.n1861 2.6005
R1528 VSS.n1864 VSS.n1863 2.6005
R1529 VSS.n1866 VSS.n1865 2.6005
R1530 VSS.n1868 VSS.n1867 2.6005
R1531 VSS.n1870 VSS.n1869 2.6005
R1532 VSS.n1872 VSS.n1871 2.6005
R1533 VSS.n1874 VSS.n1873 2.6005
R1534 VSS.n1876 VSS.n1875 2.6005
R1535 VSS.n1878 VSS.n1877 2.6005
R1536 VSS.n1880 VSS.n1879 2.6005
R1537 VSS.n1883 VSS.n1882 2.6005
R1538 VSS.n1886 VSS.n1885 2.6005
R1539 VSS.n1888 VSS.n1887 2.6005
R1540 VSS.n1890 VSS.n1889 2.6005
R1541 VSS.n1892 VSS.n1891 2.6005
R1542 VSS.n1894 VSS.n1893 2.6005
R1543 VSS.n1896 VSS.n1895 2.6005
R1544 VSS.n1828 VSS.n1827 2.6005
R1545 VSS.n1825 VSS.n1824 2.6005
R1546 VSS.n1825 VSS.n1822 2.6005
R1547 VSS.n1821 VSS.n1422 2.6005
R1548 VSS.n408 VSS.n407 2.6005
R1549 VSS.n405 VSS.n404 2.6005
R1550 VSS.n402 VSS.n401 2.6005
R1551 VSS.n400 VSS.n399 2.6005
R1552 VSS.n397 VSS.n396 2.6005
R1553 VSS.n395 VSS.n394 2.6005
R1554 VSS.n392 VSS.n391 2.6005
R1555 VSS.n390 VSS.n389 2.6005
R1556 VSS.n387 VSS.n386 2.6005
R1557 VSS.n385 VSS.n384 2.6005
R1558 VSS.n382 VSS.n381 2.6005
R1559 VSS.n380 VSS.n379 2.6005
R1560 VSS.n377 VSS.n376 2.6005
R1561 VSS.n375 VSS.n374 2.6005
R1562 VSS.n372 VSS.n371 2.6005
R1563 VSS.n370 VSS.n369 2.6005
R1564 VSS.n367 VSS.n366 2.6005
R1565 VSS.n365 VSS.n364 2.6005
R1566 VSS.n362 VSS.n361 2.6005
R1567 VSS.n360 VSS.n359 2.6005
R1568 VSS.n357 VSS.n356 2.6005
R1569 VSS.n355 VSS.n354 2.6005
R1570 VSS.n352 VSS.n351 2.6005
R1571 VSS.n350 VSS.n349 2.6005
R1572 VSS.n348 VSS.n347 2.6005
R1573 VSS.n346 VSS.n345 2.6005
R1574 VSS.n344 VSS.n343 2.6005
R1575 VSS.n342 VSS.n341 2.6005
R1576 VSS.n340 VSS.n339 2.6005
R1577 VSS.n338 VSS.n337 2.6005
R1578 VSS.n336 VSS.n335 2.6005
R1579 VSS.n334 VSS.n333 2.6005
R1580 VSS.n332 VSS.n331 2.6005
R1581 VSS.n330 VSS.n329 2.6005
R1582 VSS.n328 VSS.n327 2.6005
R1583 VSS.n326 VSS.n325 2.6005
R1584 VSS.n324 VSS.n323 2.6005
R1585 VSS.n322 VSS.n321 2.6005
R1586 VSS.n320 VSS.n319 2.6005
R1587 VSS.n318 VSS.n317 2.6005
R1588 VSS.n316 VSS.n315 2.6005
R1589 VSS.n314 VSS.n313 2.6005
R1590 VSS.n312 VSS.n311 2.6005
R1591 VSS.n310 VSS.n309 2.6005
R1592 VSS.n308 VSS.n307 2.6005
R1593 VSS.n306 VSS.n305 2.6005
R1594 VSS.n304 VSS.n303 2.6005
R1595 VSS.n302 VSS.n301 2.6005
R1596 VSS.n300 VSS.n299 2.6005
R1597 VSS.n298 VSS.n297 2.6005
R1598 VSS.n296 VSS.n295 2.6005
R1599 VSS.n294 VSS.n293 2.6005
R1600 VSS.n292 VSS.n291 2.6005
R1601 VSS.n290 VSS.n289 2.6005
R1602 VSS.n288 VSS.n287 2.6005
R1603 VSS.n286 VSS.n285 2.6005
R1604 VSS.n1411 VSS.n1410 2.6005
R1605 VSS.n1413 VSS.n1412 2.6005
R1606 VSS.n1415 VSS.n1414 2.6005
R1607 VSS.n1417 VSS.n1416 2.6005
R1608 VSS.n1419 VSS.n1418 2.6005
R1609 VSS.n1421 VSS.n1420 2.6005
R1610 VSS.n410 VSS.n409 2.6005
R1611 VSS.n1015 VSS.n1014 2.6005
R1612 VSS.n1014 VSS.n1013 2.6005
R1613 VSS.n1018 VSS.n1017 2.6005
R1614 VSS.n1017 VSS.n1016 2.6005
R1615 VSS.n1021 VSS.n1020 2.6005
R1616 VSS.n1020 VSS.n1019 2.6005
R1617 VSS.n1024 VSS.n1023 2.6005
R1618 VSS.n1023 VSS.n1022 2.6005
R1619 VSS.n1027 VSS.n1026 2.6005
R1620 VSS.n1026 VSS.n1025 2.6005
R1621 VSS.n1030 VSS.n1029 2.6005
R1622 VSS.n1029 VSS.n1028 2.6005
R1623 VSS.n1034 VSS.n1033 2.6005
R1624 VSS.n1033 VSS.n1032 2.6005
R1625 VSS.n1038 VSS.n1037 2.6005
R1626 VSS.n1037 VSS.n1036 2.6005
R1627 VSS.n1041 VSS.n1040 2.6005
R1628 VSS.n1040 VSS.n1039 2.6005
R1629 VSS.n1044 VSS.n1043 2.6005
R1630 VSS.n1043 VSS.n1042 2.6005
R1631 VSS.n1047 VSS.n1046 2.6005
R1632 VSS.n1046 VSS.n1045 2.6005
R1633 VSS.n1050 VSS.n1049 2.6005
R1634 VSS.n1049 VSS.n1048 2.6005
R1635 VSS.n1053 VSS.n1052 2.6005
R1636 VSS.n1052 VSS.n1051 2.6005
R1637 VSS.n1056 VSS.n1055 2.6005
R1638 VSS.n1055 VSS.n1054 2.6005
R1639 VSS.n1059 VSS.n1058 2.6005
R1640 VSS.n1058 VSS.n1057 2.6005
R1641 VSS.n1062 VSS.n1061 2.6005
R1642 VSS.n1061 VSS.n1060 2.6005
R1643 VSS.n1065 VSS.n1064 2.6005
R1644 VSS.n1064 VSS.n1063 2.6005
R1645 VSS.n1068 VSS.n1067 2.6005
R1646 VSS.n1067 VSS.n1066 2.6005
R1647 VSS.n1071 VSS.n1070 2.6005
R1648 VSS.n1070 VSS.n1069 2.6005
R1649 VSS.n1074 VSS.n1073 2.6005
R1650 VSS.n1073 VSS.n1072 2.6005
R1651 VSS.n1077 VSS.n1076 2.6005
R1652 VSS.n1076 VSS.n1075 2.6005
R1653 VSS.n1080 VSS.n1079 2.6005
R1654 VSS.n1079 VSS.n1078 2.6005
R1655 VSS.n1083 VSS.n1082 2.6005
R1656 VSS.n1082 VSS.n1081 2.6005
R1657 VSS.n1086 VSS.n1085 2.6005
R1658 VSS.n1085 VSS.n1084 2.6005
R1659 VSS.n1090 VSS.n1089 2.6005
R1660 VSS.n1089 VSS.n1088 2.6005
R1661 VSS.n1094 VSS.n1093 2.6005
R1662 VSS.n1093 VSS.n1092 2.6005
R1663 VSS.n1097 VSS.n1096 2.6005
R1664 VSS.n1096 VSS.n1095 2.6005
R1665 VSS.n1100 VSS.n1099 2.6005
R1666 VSS.n1099 VSS.n1098 2.6005
R1667 VSS.n1103 VSS.n1102 2.6005
R1668 VSS.n1102 VSS.n1101 2.6005
R1669 VSS.n1106 VSS.n1105 2.6005
R1670 VSS.n1105 VSS.n1104 2.6005
R1671 VSS.n1109 VSS.n1108 2.6005
R1672 VSS.n1108 VSS.n1107 2.6005
R1673 VSS.n1011 VSS.n1010 2.6005
R1674 VSS.n1538 VSS.n1537 2.6005
R1675 VSS.n1536 VSS.n1535 2.6005
R1676 VSS.n1534 VSS.n1533 2.6005
R1677 VSS.n1532 VSS.n1531 2.6005
R1678 VSS.n1530 VSS.n1529 2.6005
R1679 VSS.n432 VSS.n431 2.6005
R1680 VSS.n434 VSS.n433 2.6005
R1681 VSS.n436 VSS.n435 2.6005
R1682 VSS.n438 VSS.n437 2.6005
R1683 VSS.n440 VSS.n439 2.6005
R1684 VSS.n442 VSS.n441 2.6005
R1685 VSS.n444 VSS.n443 2.6005
R1686 VSS.n446 VSS.n445 2.6005
R1687 VSS.n448 VSS.n447 2.6005
R1688 VSS.n450 VSS.n449 2.6005
R1689 VSS.n452 VSS.n451 2.6005
R1690 VSS.n454 VSS.n453 2.6005
R1691 VSS.n456 VSS.n455 2.6005
R1692 VSS.n458 VSS.n457 2.6005
R1693 VSS.n460 VSS.n459 2.6005
R1694 VSS.n462 VSS.n461 2.6005
R1695 VSS.n464 VSS.n463 2.6005
R1696 VSS.n466 VSS.n465 2.6005
R1697 VSS.n468 VSS.n467 2.6005
R1698 VSS.n470 VSS.n469 2.6005
R1699 VSS.n472 VSS.n471 2.6005
R1700 VSS.n474 VSS.n473 2.6005
R1701 VSS.n476 VSS.n475 2.6005
R1702 VSS.n478 VSS.n477 2.6005
R1703 VSS.n480 VSS.n479 2.6005
R1704 VSS.n482 VSS.n481 2.6005
R1705 VSS.n484 VSS.n483 2.6005
R1706 VSS.n486 VSS.n485 2.6005
R1707 VSS.n488 VSS.n487 2.6005
R1708 VSS.n490 VSS.n489 2.6005
R1709 VSS.n492 VSS.n491 2.6005
R1710 VSS.n494 VSS.n493 2.6005
R1711 VSS.n496 VSS.n495 2.6005
R1712 VSS.n498 VSS.n497 2.6005
R1713 VSS.n500 VSS.n499 2.6005
R1714 VSS.n502 VSS.n501 2.6005
R1715 VSS.n504 VSS.n503 2.6005
R1716 VSS.n506 VSS.n505 2.6005
R1717 VSS.n508 VSS.n507 2.6005
R1718 VSS.n510 VSS.n509 2.6005
R1719 VSS.n512 VSS.n511 2.6005
R1720 VSS.n514 VSS.n513 2.6005
R1721 VSS.n516 VSS.n515 2.6005
R1722 VSS.n518 VSS.n517 2.6005
R1723 VSS.n520 VSS.n519 2.6005
R1724 VSS.n522 VSS.n521 2.6005
R1725 VSS.n525 VSS.n524 2.6005
R1726 VSS.n527 VSS.n526 2.6005
R1727 VSS.n530 VSS.n529 2.6005
R1728 VSS.n532 VSS.n531 2.6005
R1729 VSS.n535 VSS.n534 2.6005
R1730 VSS.n537 VSS.n536 2.6005
R1731 VSS.n540 VSS.n539 2.6005
R1732 VSS.n542 VSS.n541 2.6005
R1733 VSS.n545 VSS.n544 2.6005
R1734 VSS.n547 VSS.n546 2.6005
R1735 VSS.n550 VSS.n549 2.6005
R1736 VSS.n1540 VSS.n1539 2.6005
R1737 VSS.n1753 VSS.n1541 2.6005
R1738 VSS.n1752 VSS.n1750 2.6005
R1739 VSS.n1755 VSS.n1754 2.6005
R1740 VSS.n1757 VSS.n1756 2.6005
R1741 VSS.n1759 VSS.n1758 2.6005
R1742 VSS.n1761 VSS.n1760 2.6005
R1743 VSS.n1763 VSS.n1762 2.6005
R1744 VSS.n1765 VSS.n1764 2.6005
R1745 VSS.n1768 VSS.n1767 2.6005
R1746 VSS.n1771 VSS.n1770 2.6005
R1747 VSS.n1773 VSS.n1772 2.6005
R1748 VSS.n1775 VSS.n1774 2.6005
R1749 VSS.n1777 VSS.n1776 2.6005
R1750 VSS.n1779 VSS.n1778 2.6005
R1751 VSS.n1781 VSS.n1780 2.6005
R1752 VSS.n1783 VSS.n1782 2.6005
R1753 VSS.n1785 VSS.n1784 2.6005
R1754 VSS.n1787 VSS.n1786 2.6005
R1755 VSS.n1789 VSS.n1788 2.6005
R1756 VSS.n1791 VSS.n1790 2.6005
R1757 VSS.n1793 VSS.n1792 2.6005
R1758 VSS.n1795 VSS.n1794 2.6005
R1759 VSS.n1797 VSS.n1796 2.6005
R1760 VSS.n1800 VSS.n1799 2.6005
R1761 VSS.n1802 VSS.n1801 2.6005
R1762 VSS.n1804 VSS.n1803 2.6005
R1763 VSS.n1807 VSS.n1806 2.6005
R1764 VSS.n1810 VSS.n1809 2.6005
R1765 VSS.n1812 VSS.n1811 2.6005
R1766 VSS.n1814 VSS.n1813 2.6005
R1767 VSS.n1816 VSS.n1815 2.6005
R1768 VSS.n1818 VSS.n1817 2.6005
R1769 VSS.n1820 VSS.n1819 2.6005
R1770 VSS.n1752 VSS.n1751 2.6005
R1771 VSS.n1749 VSS.n1748 2.6005
R1772 VSS.n1749 VSS.n1746 2.6005
R1773 VSS.n1745 VSS.n1554 2.6005
R1774 VSS.n675 VSS.n674 2.6005
R1775 VSS.n672 VSS.n671 2.6005
R1776 VSS.n669 VSS.n668 2.6005
R1777 VSS.n667 VSS.n666 2.6005
R1778 VSS.n664 VSS.n663 2.6005
R1779 VSS.n662 VSS.n661 2.6005
R1780 VSS.n659 VSS.n658 2.6005
R1781 VSS.n657 VSS.n656 2.6005
R1782 VSS.n654 VSS.n653 2.6005
R1783 VSS.n652 VSS.n651 2.6005
R1784 VSS.n649 VSS.n648 2.6005
R1785 VSS.n647 VSS.n646 2.6005
R1786 VSS.n644 VSS.n643 2.6005
R1787 VSS.n642 VSS.n641 2.6005
R1788 VSS.n639 VSS.n638 2.6005
R1789 VSS.n637 VSS.n636 2.6005
R1790 VSS.n634 VSS.n633 2.6005
R1791 VSS.n632 VSS.n631 2.6005
R1792 VSS.n629 VSS.n628 2.6005
R1793 VSS.n627 VSS.n626 2.6005
R1794 VSS.n624 VSS.n623 2.6005
R1795 VSS.n622 VSS.n621 2.6005
R1796 VSS.n619 VSS.n618 2.6005
R1797 VSS.n617 VSS.n616 2.6005
R1798 VSS.n615 VSS.n614 2.6005
R1799 VSS.n613 VSS.n612 2.6005
R1800 VSS.n611 VSS.n610 2.6005
R1801 VSS.n609 VSS.n608 2.6005
R1802 VSS.n607 VSS.n606 2.6005
R1803 VSS.n605 VSS.n604 2.6005
R1804 VSS.n603 VSS.n602 2.6005
R1805 VSS.n601 VSS.n600 2.6005
R1806 VSS.n599 VSS.n598 2.6005
R1807 VSS.n597 VSS.n596 2.6005
R1808 VSS.n595 VSS.n594 2.6005
R1809 VSS.n593 VSS.n592 2.6005
R1810 VSS.n591 VSS.n590 2.6005
R1811 VSS.n589 VSS.n588 2.6005
R1812 VSS.n587 VSS.n586 2.6005
R1813 VSS.n585 VSS.n584 2.6005
R1814 VSS.n583 VSS.n582 2.6005
R1815 VSS.n581 VSS.n580 2.6005
R1816 VSS.n579 VSS.n578 2.6005
R1817 VSS.n577 VSS.n576 2.6005
R1818 VSS.n575 VSS.n574 2.6005
R1819 VSS.n573 VSS.n572 2.6005
R1820 VSS.n571 VSS.n570 2.6005
R1821 VSS.n569 VSS.n568 2.6005
R1822 VSS.n567 VSS.n566 2.6005
R1823 VSS.n565 VSS.n564 2.6005
R1824 VSS.n563 VSS.n562 2.6005
R1825 VSS.n561 VSS.n560 2.6005
R1826 VSS.n559 VSS.n558 2.6005
R1827 VSS.n557 VSS.n556 2.6005
R1828 VSS.n555 VSS.n554 2.6005
R1829 VSS.n553 VSS.n552 2.6005
R1830 VSS.n1543 VSS.n1542 2.6005
R1831 VSS.n1545 VSS.n1544 2.6005
R1832 VSS.n1547 VSS.n1546 2.6005
R1833 VSS.n1549 VSS.n1548 2.6005
R1834 VSS.n1551 VSS.n1550 2.6005
R1835 VSS.n1553 VSS.n1552 2.6005
R1836 VSS.n677 VSS.n676 2.6005
R1837 VSS.n854 VSS.n853 2.6005
R1838 VSS.n853 VSS.n852 2.6005
R1839 VSS.n857 VSS.n856 2.6005
R1840 VSS.n856 VSS.n855 2.6005
R1841 VSS.n860 VSS.n859 2.6005
R1842 VSS.n859 VSS.n858 2.6005
R1843 VSS.n863 VSS.n862 2.6005
R1844 VSS.n862 VSS.n861 2.6005
R1845 VSS.n866 VSS.n865 2.6005
R1846 VSS.n865 VSS.n864 2.6005
R1847 VSS.n869 VSS.n868 2.6005
R1848 VSS.n868 VSS.n867 2.6005
R1849 VSS.n873 VSS.n872 2.6005
R1850 VSS.n872 VSS.n871 2.6005
R1851 VSS.n877 VSS.n876 2.6005
R1852 VSS.n876 VSS.n875 2.6005
R1853 VSS.n880 VSS.n879 2.6005
R1854 VSS.n879 VSS.n878 2.6005
R1855 VSS.n883 VSS.n882 2.6005
R1856 VSS.n882 VSS.n881 2.6005
R1857 VSS.n886 VSS.n885 2.6005
R1858 VSS.n885 VSS.n884 2.6005
R1859 VSS.n889 VSS.n888 2.6005
R1860 VSS.n888 VSS.n887 2.6005
R1861 VSS.n892 VSS.n891 2.6005
R1862 VSS.n891 VSS.n890 2.6005
R1863 VSS.n895 VSS.n894 2.6005
R1864 VSS.n894 VSS.n893 2.6005
R1865 VSS.n898 VSS.n897 2.6005
R1866 VSS.n897 VSS.n896 2.6005
R1867 VSS.n901 VSS.n900 2.6005
R1868 VSS.n900 VSS.n899 2.6005
R1869 VSS.n904 VSS.n903 2.6005
R1870 VSS.n903 VSS.n902 2.6005
R1871 VSS.n907 VSS.n906 2.6005
R1872 VSS.n906 VSS.n905 2.6005
R1873 VSS.n910 VSS.n909 2.6005
R1874 VSS.n909 VSS.n908 2.6005
R1875 VSS.n913 VSS.n912 2.6005
R1876 VSS.n912 VSS.n911 2.6005
R1877 VSS.n916 VSS.n915 2.6005
R1878 VSS.n915 VSS.n914 2.6005
R1879 VSS.n919 VSS.n918 2.6005
R1880 VSS.n918 VSS.n917 2.6005
R1881 VSS.n922 VSS.n921 2.6005
R1882 VSS.n921 VSS.n920 2.6005
R1883 VSS.n925 VSS.n924 2.6005
R1884 VSS.n924 VSS.n923 2.6005
R1885 VSS.n929 VSS.n928 2.6005
R1886 VSS.n928 VSS.n927 2.6005
R1887 VSS.n933 VSS.n932 2.6005
R1888 VSS.n932 VSS.n931 2.6005
R1889 VSS.n936 VSS.n935 2.6005
R1890 VSS.n935 VSS.n934 2.6005
R1891 VSS.n939 VSS.n938 2.6005
R1892 VSS.n938 VSS.n937 2.6005
R1893 VSS.n942 VSS.n941 2.6005
R1894 VSS.n941 VSS.n940 2.6005
R1895 VSS.n945 VSS.n944 2.6005
R1896 VSS.n944 VSS.n943 2.6005
R1897 VSS.n948 VSS.n947 2.6005
R1898 VSS.n947 VSS.n946 2.6005
R1899 VSS.n850 VSS.n849 2.6005
R1900 VSS.n817 VSS.n816 2.6005
R1901 VSS.n814 VSS.n813 2.6005
R1902 VSS.n812 VSS.n811 2.6005
R1903 VSS.n809 VSS.n808 2.6005
R1904 VSS.n807 VSS.n806 2.6005
R1905 VSS.n804 VSS.n803 2.6005
R1906 VSS.n802 VSS.n801 2.6005
R1907 VSS.n799 VSS.n798 2.6005
R1908 VSS.n797 VSS.n796 2.6005
R1909 VSS.n794 VSS.n793 2.6005
R1910 VSS.n792 VSS.n791 2.6005
R1911 VSS.n789 VSS.n788 2.6005
R1912 VSS.n787 VSS.n786 2.6005
R1913 VSS.n785 VSS.n784 2.6005
R1914 VSS.n783 VSS.n782 2.6005
R1915 VSS.n781 VSS.n780 2.6005
R1916 VSS.n779 VSS.n778 2.6005
R1917 VSS.n777 VSS.n776 2.6005
R1918 VSS.n775 VSS.n774 2.6005
R1919 VSS.n773 VSS.n772 2.6005
R1920 VSS.n771 VSS.n770 2.6005
R1921 VSS.n769 VSS.n768 2.6005
R1922 VSS.n767 VSS.n766 2.6005
R1923 VSS.n765 VSS.n764 2.6005
R1924 VSS.n763 VSS.n762 2.6005
R1925 VSS.n761 VSS.n760 2.6005
R1926 VSS.n759 VSS.n758 2.6005
R1927 VSS.n757 VSS.n756 2.6005
R1928 VSS.n755 VSS.n754 2.6005
R1929 VSS.n753 VSS.n752 2.6005
R1930 VSS.n751 VSS.n750 2.6005
R1931 VSS.n749 VSS.n748 2.6005
R1932 VSS.n747 VSS.n746 2.6005
R1933 VSS.n745 VSS.n744 2.6005
R1934 VSS.n743 VSS.n742 2.6005
R1935 VSS.n741 VSS.n740 2.6005
R1936 VSS.n739 VSS.n738 2.6005
R1937 VSS.n737 VSS.n736 2.6005
R1938 VSS.n735 VSS.n734 2.6005
R1939 VSS.n733 VSS.n732 2.6005
R1940 VSS.n731 VSS.n730 2.6005
R1941 VSS.n729 VSS.n728 2.6005
R1942 VSS.n727 VSS.n726 2.6005
R1943 VSS.n725 VSS.n724 2.6005
R1944 VSS.n723 VSS.n722 2.6005
R1945 VSS.n721 VSS.n720 2.6005
R1946 VSS.n719 VSS.n718 2.6005
R1947 VSS.n717 VSS.n716 2.6005
R1948 VSS.n715 VSS.n714 2.6005
R1949 VSS.n713 VSS.n712 2.6005
R1950 VSS.n711 VSS.n710 2.6005
R1951 VSS.n709 VSS.n708 2.6005
R1952 VSS.n707 VSS.n706 2.6005
R1953 VSS.n705 VSS.n704 2.6005
R1954 VSS.n703 VSS.n702 2.6005
R1955 VSS.n701 VSS.n700 2.6005
R1956 VSS.n699 VSS.n698 2.6005
R1957 VSS.n1658 VSS.n1657 2.6005
R1958 VSS.n1660 VSS.n1659 2.6005
R1959 VSS.n1662 VSS.n1661 2.6005
R1960 VSS.n1664 VSS.n1663 2.6005
R1961 VSS.n1666 VSS.n1665 2.6005
R1962 VSS.n1668 VSS.n1667 2.6005
R1963 VSS.n1673 VSS.n1669 2.6005
R1964 VSS.n1672 VSS.n1670 2.6005
R1965 VSS.n1675 VSS.n1674 2.6005
R1966 VSS.n1677 VSS.n1676 2.6005
R1967 VSS.n1679 VSS.n1678 2.6005
R1968 VSS.n1681 VSS.n1680 2.6005
R1969 VSS.n1683 VSS.n1682 2.6005
R1970 VSS.n1685 VSS.n1684 2.6005
R1971 VSS.n1692 VSS.n1691 2.6005
R1972 VSS.n1695 VSS.n1694 2.6005
R1973 VSS.n1697 VSS.n1696 2.6005
R1974 VSS.n1699 VSS.n1698 2.6005
R1975 VSS.n1702 VSS.n1701 2.6005
R1976 VSS.n1704 VSS.n1703 2.6005
R1977 VSS.n1706 VSS.n1705 2.6005
R1978 VSS.n1708 VSS.n1707 2.6005
R1979 VSS.n1710 VSS.n1709 2.6005
R1980 VSS.n1712 VSS.n1711 2.6005
R1981 VSS.n1714 VSS.n1713 2.6005
R1982 VSS.n1716 VSS.n1715 2.6005
R1983 VSS.n1718 VSS.n1717 2.6005
R1984 VSS.n1720 VSS.n1719 2.6005
R1985 VSS.n1722 VSS.n1721 2.6005
R1986 VSS.n1724 VSS.n1723 2.6005
R1987 VSS.n1726 VSS.n1725 2.6005
R1988 VSS.n1728 VSS.n1727 2.6005
R1989 VSS.n1731 VSS.n1730 2.6005
R1990 VSS.n1734 VSS.n1733 2.6005
R1991 VSS.n1736 VSS.n1735 2.6005
R1992 VSS.n1738 VSS.n1737 2.6005
R1993 VSS.n1740 VSS.n1739 2.6005
R1994 VSS.n1742 VSS.n1741 2.6005
R1995 VSS.n1744 VSS.n1743 2.6005
R1996 VSS.n1672 VSS.n1671 2.6005
R1997 VSS.n2584 VSS.n2583 2.6005
R1998 VSS.n2587 VSS.n2586 2.6005
R1999 VSS.n2838 VSS.n2837 2.6005
R2000 VSS.n2729 VSS.n2728 2.6005
R2001 VSS.n2727 VSS.n2726 2.6005
R2002 VSS.n2725 VSS.n2724 2.6005
R2003 VSS.n2723 VSS.n2722 2.6005
R2004 VSS.n2721 VSS.n2720 2.6005
R2005 VSS.n2719 VSS.n2718 2.6005
R2006 VSS.n2717 VSS.n2716 2.6005
R2007 VSS.n2714 VSS.n2713 2.6005
R2008 VSS.n2712 VSS.n2711 2.6005
R2009 VSS.n2710 VSS.n2709 2.6005
R2010 VSS.n2707 VSS.n2706 2.6005
R2011 VSS.n2705 VSS.n2704 2.6005
R2012 VSS.n2703 VSS.n2702 2.6005
R2013 VSS.n2701 VSS.n2700 2.6005
R2014 VSS.n2699 VSS.n2698 2.6005
R2015 VSS.n2697 VSS.n2696 2.6005
R2016 VSS.n2695 VSS.n2694 2.6005
R2017 VSS.n2693 VSS.n2692 2.6005
R2018 VSS.n2691 VSS.n2690 2.6005
R2019 VSS.n2689 VSS.n2688 2.6005
R2020 VSS.n2687 VSS.n2686 2.6005
R2021 VSS.n2684 VSS.n2683 2.6005
R2022 VSS.n2682 VSS.n2681 2.6005
R2023 VSS.n2680 VSS.n2679 2.6005
R2024 VSS.n2678 VSS.n2677 2.6005
R2025 VSS.n2676 VSS.n2675 2.6005
R2026 VSS.n2674 VSS.n2673 2.6005
R2027 VSS.n2671 VSS.n2670 2.6005
R2028 VSS.n2669 VSS.n2668 2.6005
R2029 VSS.n2667 VSS.n2666 2.6005
R2030 VSS.n2665 VSS.n2664 2.6005
R2031 VSS.n2663 VSS.n2662 2.6005
R2032 VSS.n2661 VSS.n2660 2.6005
R2033 VSS.n2659 VSS.n2658 2.6005
R2034 VSS.n2657 VSS.n2656 2.6005
R2035 VSS.n2654 VSS.n2653 2.6005
R2036 VSS.n2652 VSS.n2651 2.6005
R2037 VSS.n2650 VSS.n2649 2.6005
R2038 VSS.n2648 VSS.n2647 2.6005
R2039 VSS.n2646 VSS.n2645 2.6005
R2040 VSS.n2644 VSS.n2643 2.6005
R2041 VSS.n2642 VSS.n2641 2.6005
R2042 VSS.n2639 VSS.n2638 2.6005
R2043 VSS.n2637 VSS.n2636 2.6005
R2044 VSS.n2635 VSS.n2634 2.6005
R2045 VSS.n2633 VSS.n2632 2.6005
R2046 VSS.n2631 VSS.n2630 2.6005
R2047 VSS.n2629 VSS.n2628 2.6005
R2048 VSS.n2626 VSS.n2625 2.6005
R2049 VSS.n2624 VSS.n2623 2.6005
R2050 VSS.n2622 VSS.n2621 2.6005
R2051 VSS.n2619 VSS.n2618 2.6005
R2052 VSS.n2617 VSS.n2616 2.6005
R2053 VSS.n2615 VSS.n2614 2.6005
R2054 VSS.n2612 VSS.n2611 2.6005
R2055 VSS.n2609 VSS.n2608 2.6005
R2056 VSS.n2606 VSS.n2605 2.6005
R2057 VSS.n2603 VSS.n2602 2.6005
R2058 VSS.n2836 VSS.n2835 2.6005
R2059 VSS.n2600 VSS.n2599 2.6005
R2060 VSS.n2599 VSS.n2598 2.6005
R2061 VSS.n2597 VSS.n2596 2.6005
R2062 VSS.n2596 VSS.n2595 2.6005
R2063 VSS.n2594 VSS.n2593 2.6005
R2064 VSS.n2593 VSS.n2592 2.6005
R2065 VSS.n2941 VSS.n2940 2.6005
R2066 VSS.n2940 VSS.n2939 2.6005
R2067 VSS.n2944 VSS.n2943 2.6005
R2068 VSS.n2943 VSS.n2942 2.6005
R2069 VSS.n2947 VSS.n2946 2.6005
R2070 VSS.n2946 VSS.n2945 2.6005
R2071 VSS.n2950 VSS.n2949 2.6005
R2072 VSS.n2949 VSS.n2948 2.6005
R2073 VSS.n2953 VSS.n2952 2.6005
R2074 VSS.n2952 VSS.n2951 2.6005
R2075 VSS.n2956 VSS.n2955 2.6005
R2076 VSS.n2955 VSS.n2954 2.6005
R2077 VSS.n2959 VSS.n2958 2.6005
R2078 VSS.n2958 VSS.n2957 2.6005
R2079 VSS.n2962 VSS.n2961 2.6005
R2080 VSS.n2961 VSS.n2960 2.6005
R2081 VSS.n2965 VSS.n2964 2.6005
R2082 VSS.n2964 VSS.n2963 2.6005
R2083 VSS.n2968 VSS.n2967 2.6005
R2084 VSS.n2967 VSS.n2966 2.6005
R2085 VSS.n2971 VSS.n2970 2.6005
R2086 VSS.n2970 VSS.n2969 2.6005
R2087 VSS.n2974 VSS.n2973 2.6005
R2088 VSS.n2973 VSS.n2972 2.6005
R2089 VSS.n2977 VSS.n2976 2.6005
R2090 VSS.n2976 VSS.n2975 2.6005
R2091 VSS.n2980 VSS.n2979 2.6005
R2092 VSS.n2979 VSS.n2978 2.6005
R2093 VSS.n2983 VSS.n2982 2.6005
R2094 VSS.n2982 VSS.n2981 2.6005
R2095 VSS.n2986 VSS.n2985 2.6005
R2096 VSS.n2985 VSS.n2984 2.6005
R2097 VSS.n2989 VSS.n2988 2.6005
R2098 VSS.n2988 VSS.n2987 2.6005
R2099 VSS.n2992 VSS.n2991 2.6005
R2100 VSS.n2991 VSS.n2990 2.6005
R2101 VSS.n2995 VSS.n2994 2.6005
R2102 VSS.n2994 VSS.n2993 2.6005
R2103 VSS.n2998 VSS.n2997 2.6005
R2104 VSS.n2997 VSS.n2996 2.6005
R2105 VSS.n3001 VSS.n3000 2.6005
R2106 VSS.n3000 VSS.n2999 2.6005
R2107 VSS.n3004 VSS.n3003 2.6005
R2108 VSS.n3003 VSS.n3002 2.6005
R2109 VSS.n3007 VSS.n3006 2.6005
R2110 VSS.n3006 VSS.n3005 2.6005
R2111 VSS.n3010 VSS.n3009 2.6005
R2112 VSS.n3009 VSS.n3008 2.6005
R2113 VSS.n3013 VSS.n3012 2.6005
R2114 VSS.n3012 VSS.n3011 2.6005
R2115 VSS.n3020 VSS.n3019 2.6005
R2116 VSS.n3015 VSS.n3014 2.6005
R2117 VSS.n3025 VSS.n3024 2.6005
R2118 VSS.n3027 VSS.n3026 2.6005
R2119 VSS.n3030 VSS.n3029 2.6005
R2120 VSS.n3032 VSS.n3031 2.6005
R2121 VSS.n3035 VSS.n3034 2.6005
R2122 VSS.n3039 VSS.n3038 2.6005
R2123 VSS.n3038 VSS.n3037 2.6005
R2124 VSS.n3042 VSS.n3041 2.6005
R2125 VSS.n3041 VSS.n3040 2.6005
R2126 VSS.n3046 VSS.n3045 2.6005
R2127 VSS.n3045 VSS.n3044 2.6005
R2128 VSS.n3049 VSS.n3048 2.6005
R2129 VSS.n3048 VSS.n3047 2.6005
R2130 VSS.n3052 VSS.n3051 2.6005
R2131 VSS.n3051 VSS.n3050 2.6005
R2132 VSS.n3056 VSS.n3055 2.6005
R2133 VSS.n3055 VSS.n3054 2.6005
R2134 VSS.n3059 VSS.n3058 2.6005
R2135 VSS.n3058 VSS.n3057 2.6005
R2136 VSS.n3062 VSS.n3061 2.6005
R2137 VSS.n3061 VSS.n3060 2.6005
R2138 VSS.n3065 VSS.n3064 2.6005
R2139 VSS.n3064 VSS.n3063 2.6005
R2140 VSS.n3068 VSS.n3067 2.6005
R2141 VSS.n3067 VSS.n3066 2.6005
R2142 VSS.n3071 VSS.n3070 2.6005
R2143 VSS.n3070 VSS.n3069 2.6005
R2144 VSS.n3075 VSS.n3074 2.6005
R2145 VSS.n3074 VSS.n3073 2.6005
R2146 VSS.n3078 VSS.n3077 2.6005
R2147 VSS.n3077 VSS.n3076 2.6005
R2148 VSS.n3081 VSS.n3080 2.6005
R2149 VSS.n3080 VSS.n3079 2.6005
R2150 VSS.n3084 VSS.n3083 2.6005
R2151 VSS.n3083 VSS.n3082 2.6005
R2152 VSS.n3087 VSS.n3086 2.6005
R2153 VSS.n3086 VSS.n3085 2.6005
R2154 VSS.n3090 VSS.n3089 2.6005
R2155 VSS.n3089 VSS.n3088 2.6005
R2156 VSS.n3093 VSS.n3092 2.6005
R2157 VSS.n3092 VSS.n3091 2.6005
R2158 VSS.n3097 VSS.n3096 2.6005
R2159 VSS.n3096 VSS.n3095 2.6005
R2160 VSS.n3100 VSS.n3099 2.6005
R2161 VSS.n3099 VSS.n3098 2.6005
R2162 VSS.n3103 VSS.n3102 2.6005
R2163 VSS.n3102 VSS.n3101 2.6005
R2164 VSS.n3106 VSS.n3105 2.6005
R2165 VSS.n3105 VSS.n3104 2.6005
R2166 VSS.n3109 VSS.n3108 2.6005
R2167 VSS.n3108 VSS.n3107 2.6005
R2168 VSS.n3112 VSS.n3111 2.6005
R2169 VSS.n3111 VSS.n3110 2.6005
R2170 VSS.n3115 VSS.n3114 2.6005
R2171 VSS.n3114 VSS.n3113 2.6005
R2172 VSS.n3118 VSS.n3117 2.6005
R2173 VSS.n3117 VSS.n3116 2.6005
R2174 VSS.n3122 VSS.n3121 2.6005
R2175 VSS.n3121 VSS.n3120 2.6005
R2176 VSS.n3125 VSS.n3124 2.6005
R2177 VSS.n3124 VSS.n3123 2.6005
R2178 VSS.n3128 VSS.n3127 2.6005
R2179 VSS.n3127 VSS.n3126 2.6005
R2180 VSS.n3131 VSS.n3130 2.6005
R2181 VSS.n3130 VSS.n3129 2.6005
R2182 VSS.n3134 VSS.n3133 2.6005
R2183 VSS.n3133 VSS.n3132 2.6005
R2184 VSS.n3137 VSS.n3136 2.6005
R2185 VSS.n3136 VSS.n3135 2.6005
R2186 VSS.n3141 VSS.n3140 2.6005
R2187 VSS.n3140 VSS.n3139 2.6005
R2188 VSS.n3144 VSS.n3143 2.6005
R2189 VSS.n3143 VSS.n3142 2.6005
R2190 VSS.n3147 VSS.n3146 2.6005
R2191 VSS.n3146 VSS.n3145 2.6005
R2192 VSS.n3150 VSS.n3149 2.6005
R2193 VSS.n3149 VSS.n3148 2.6005
R2194 VSS.n3153 VSS.n3152 2.6005
R2195 VSS.n3152 VSS.n3151 2.6005
R2196 VSS.n3156 VSS.n3155 2.6005
R2197 VSS.n3155 VSS.n3154 2.6005
R2198 VSS.n3159 VSS.n3158 2.6005
R2199 VSS.n3158 VSS.n3157 2.6005
R2200 VSS.n3163 VSS.n3162 2.6005
R2201 VSS.n3162 VSS.n3161 2.6005
R2202 VSS.n3167 VSS.n3166 2.6005
R2203 VSS.n3166 VSS.n3165 2.6005
R2204 VSS.n3170 VSS.n3169 2.6005
R2205 VSS.n3169 VSS.n3168 2.6005
R2206 VSS.n3174 VSS.n3173 2.6005
R2207 VSS.n3173 VSS.n3172 2.6005
R2208 VSS.n3178 VSS.n3177 2.6005
R2209 VSS.n3177 VSS.n3176 2.6005
R2210 VSS.n3181 VSS.n3180 2.6005
R2211 VSS.n3180 VSS.n3179 2.6005
R2212 VSS.n3184 VSS.n3183 2.6005
R2213 VSS.n3183 VSS.n3182 2.6005
R2214 VSS.n3188 VSS.n3187 2.6005
R2215 VSS.n3187 VSS.n3186 2.6005
R2216 VSS.n3191 VSS.n3190 2.6005
R2217 VSS.n3190 VSS.n3189 2.6005
R2218 VSS.n3194 VSS.n3193 2.6005
R2219 VSS.n3193 VSS.n3192 2.6005
R2220 VSS.n3197 VSS.n3196 2.6005
R2221 VSS.n3196 VSS.n3195 2.6005
R2222 VSS.n3200 VSS.n3199 2.6005
R2223 VSS.n3199 VSS.n3198 2.6005
R2224 VSS.n3203 VSS.n3202 2.6005
R2225 VSS.n3202 VSS.n3201 2.6005
R2226 VSS.n3206 VSS.n3205 2.6005
R2227 VSS.n3205 VSS.n3204 2.6005
R2228 VSS.n3213 VSS.n3212 2.6005
R2229 VSS.n3258 VSS.n3257 2.6005
R2230 VSS.n3218 VSS.n3217 2.6005
R2231 VSS.n3256 VSS.n3255 2.6005
R2232 VSS.n3253 VSS.n3252 2.6005
R2233 VSS.n3251 VSS.n3250 2.6005
R2234 VSS.n3248 VSS.n3247 2.6005
R2235 VSS.n3246 VSS.n3245 2.6005
R2236 VSS.n3243 VSS.n3242 2.6005
R2237 VSS.n3241 VSS.n3240 2.6005
R2238 VSS.n3238 VSS.n3237 2.6005
R2239 VSS.n3236 VSS.n3235 2.6005
R2240 VSS.n3233 VSS.n3232 2.6005
R2241 VSS.n3231 VSS.n3230 2.6005
R2242 VSS.n3228 VSS.n3227 2.6005
R2243 VSS.n3226 VSS.n3225 2.6005
R2244 VSS.n3223 VSS.n3222 2.6005
R2245 VSS.n3221 VSS.n3220 2.6005
R2246 VSS.n2517 VSS.n2516 2.6005
R2247 VSS.n2511 VSS.n2510 2.6005
R2248 VSS.n2513 VSS.n2512 2.6005
R2249 VSS.n2515 VSS.n2514 2.6005
R2250 VSS.n2526 VSS.n2525 2.6005
R2251 VSS.n2528 VSS.n2527 2.6005
R2252 VSS.n2530 VSS.n2529 2.6005
R2253 VSS.n2532 VSS.n2531 2.6005
R2254 VSS.n2534 VSS.n2533 2.6005
R2255 VSS.n2537 VSS.n2536 2.6005
R2256 VSS.n2540 VSS.n2539 2.6005
R2257 VSS.n2543 VSS.n2542 2.6005
R2258 VSS.n2550 VSS.n2548 2.6005
R2259 VSS.n2550 VSS.n2549 2.6005
R2260 VSS.n2877 VSS.n2876 2.6005
R2261 VSS.n2874 VSS.n2873 2.6005
R2262 VSS.n2872 VSS.n2871 2.6005
R2263 VSS.n2863 VSS.n2862 2.6005
R2264 VSS.n2861 VSS.n2860 2.6005
R2265 VSS.n2858 VSS.n2857 2.6005
R2266 VSS.n2856 VSS.n2855 2.6005
R2267 VSS.n2853 VSS.n2852 2.6005
R2268 VSS.n2851 VSS.n2850 2.6005
R2269 VSS.n2848 VSS.n2847 2.6005
R2270 VSS.n2846 VSS.n2845 2.6005
R2271 VSS.n2843 VSS.n2842 2.6005
R2272 VSS.n2841 VSS.n2840 2.6005
R2273 VSS.n2472 VSS.n2466 2.6005
R2274 VSS.n2508 VSS.n2507 2.6005
R2275 VSS.n2475 VSS.n2474 2.6005
R2276 VSS.n2474 VSS.n2473 2.6005
R2277 VSS.n2478 VSS.n2477 2.6005
R2278 VSS.n2477 VSS.n2476 2.6005
R2279 VSS.n2484 VSS.n2483 2.6005
R2280 VSS.n2483 VSS.n2482 2.6005
R2281 VSS.n2487 VSS.n2486 2.6005
R2282 VSS.n2486 VSS.n2485 2.6005
R2283 VSS.n2491 VSS.n2490 2.6005
R2284 VSS.n2490 VSS.n2489 2.6005
R2285 VSS.n2494 VSS.n2493 2.6005
R2286 VSS.n2493 VSS.n2492 2.6005
R2287 VSS.n2497 VSS.n2496 2.6005
R2288 VSS.n2496 VSS.n2495 2.6005
R2289 VSS.n2500 VSS.n2499 2.6005
R2290 VSS.n2499 VSS.n2498 2.6005
R2291 VSS.n2503 VSS.n2502 2.6005
R2292 VSS.n2502 VSS.n2501 2.6005
R2293 VSS.n2506 VSS.n2505 2.6005
R2294 VSS.n2505 VSS.n2504 2.6005
R2295 VSS.n2834 VSS.n2833 2.6005
R2296 VSS.n2832 VSS.n2831 2.6005
R2297 VSS.n2829 VSS.n2828 2.6005
R2298 VSS.n2827 VSS.n2826 2.6005
R2299 VSS.n2824 VSS.n2823 2.6005
R2300 VSS.n2822 VSS.n2821 2.6005
R2301 VSS.n2819 VSS.n2818 2.6005
R2302 VSS.n2816 VSS.n2815 2.6005
R2303 VSS.n2814 VSS.n2813 2.6005
R2304 VSS.n2811 VSS.n2810 2.6005
R2305 VSS.n2809 VSS.n2808 2.6005
R2306 VSS.n2806 VSS.n2805 2.6005
R2307 VSS.n2803 VSS.n2802 2.6005
R2308 VSS.n2801 VSS.n2800 2.6005
R2309 VSS.n2799 VSS.n2798 2.6005
R2310 VSS.n2797 VSS.n2796 2.6005
R2311 VSS.n2795 VSS.n2794 2.6005
R2312 VSS.n2793 VSS.n2792 2.6005
R2313 VSS.n2791 VSS.n2790 2.6005
R2314 VSS.n2789 VSS.n2788 2.6005
R2315 VSS.n2787 VSS.n2786 2.6005
R2316 VSS.n2785 VSS.n2784 2.6005
R2317 VSS.n2783 VSS.n2782 2.6005
R2318 VSS.n2781 VSS.n2780 2.6005
R2319 VSS.n2779 VSS.n2778 2.6005
R2320 VSS.n2777 VSS.n2776 2.6005
R2321 VSS.n2775 VSS.n2774 2.6005
R2322 VSS.n2773 VSS.n2772 2.6005
R2323 VSS.n2770 VSS.n2769 2.6005
R2324 VSS.n2768 VSS.n2767 2.6005
R2325 VSS.n2766 VSS.n2765 2.6005
R2326 VSS.n2764 VSS.n2763 2.6005
R2327 VSS.n2762 VSS.n2761 2.6005
R2328 VSS.n2759 VSS.n2758 2.6005
R2329 VSS.n2757 VSS.n2756 2.6005
R2330 VSS.n2755 VSS.n2754 2.6005
R2331 VSS.n3557 VSS.n3556 2.6005
R2332 VSS.n3560 VSS.n3559 2.6005
R2333 VSS.n3562 VSS.n3561 2.6005
R2334 VSS.n3564 VSS.n3563 2.6005
R2335 VSS.n3566 VSS.n3565 2.6005
R2336 VSS.n3568 VSS.n3567 2.6005
R2337 VSS.n3571 VSS.n3570 2.6005
R2338 VSS.n3573 VSS.n3572 2.6005
R2339 VSS.n3575 VSS.n3574 2.6005
R2340 VSS.n3577 VSS.n3576 2.6005
R2341 VSS.n3580 VSS.n3579 2.6005
R2342 VSS.n3582 VSS.n3581 2.6005
R2343 VSS.n3584 VSS.n3583 2.6005
R2344 VSS.n3586 VSS.n3585 2.6005
R2345 VSS.n3589 VSS.n3588 2.6005
R2346 VSS.n3591 VSS.n3590 2.6005
R2347 VSS.n3595 VSS.n3594 2.6005
R2348 VSS.n3597 VSS.n3596 2.6005
R2349 VSS.n3600 VSS.n3599 2.6005
R2350 VSS.n3675 VSS.n3674 2.6005
R2351 VSS.n3641 VSS.n3640 2.6005
R2352 VSS.n3644 VSS.n3643 2.6005
R2353 VSS.n3643 VSS.n3642 2.6005
R2354 VSS.n3647 VSS.n3646 2.6005
R2355 VSS.n3646 VSS.n3645 2.6005
R2356 VSS.n3651 VSS.n3650 2.6005
R2357 VSS.n3650 VSS.n3649 2.6005
R2358 VSS.n3654 VSS.n3653 2.6005
R2359 VSS.n3653 VSS.n3652 2.6005
R2360 VSS.n3658 VSS.n3657 2.6005
R2361 VSS.n3657 VSS.n3656 2.6005
R2362 VSS.n3661 VSS.n3660 2.6005
R2363 VSS.n3660 VSS.n3659 2.6005
R2364 VSS.n3664 VSS.n3663 2.6005
R2365 VSS.n3663 VSS.n3662 2.6005
R2366 VSS.n3667 VSS.n3666 2.6005
R2367 VSS.n3666 VSS.n3665 2.6005
R2368 VSS.n3670 VSS.n3669 2.6005
R2369 VSS.n3669 VSS.n3668 2.6005
R2370 VSS.n3673 VSS.n3672 2.6005
R2371 VSS.n3672 VSS.n3671 2.6005
R2372 VSS.n3751 VSS.n3750 2.6005
R2373 VSS.n3749 VSS.n3748 2.6005
R2374 VSS.n3746 VSS.n3745 2.6005
R2375 VSS.n3744 VSS.n3743 2.6005
R2376 VSS.n3741 VSS.n3740 2.6005
R2377 VSS.n3739 VSS.n3738 2.6005
R2378 VSS.n3736 VSS.n3735 2.6005
R2379 VSS.n3734 VSS.n3733 2.6005
R2380 VSS.n3731 VSS.n3730 2.6005
R2381 VSS.n3729 VSS.n3728 2.6005
R2382 VSS.n3726 VSS.n3725 2.6005
R2383 VSS.n3724 VSS.n3723 2.6005
R2384 VSS.n3721 VSS.n3720 2.6005
R2385 VSS.n3719 VSS.n3718 2.6005
R2386 VSS.n3716 VSS.n3715 2.6005
R2387 VSS.n3714 VSS.n3713 2.6005
R2388 VSS.n3711 VSS.n3710 2.6005
R2389 VSS.n3709 VSS.n3708 2.6005
R2390 VSS.n3707 VSS.n3706 2.6005
R2391 VSS.n3705 VSS.n3704 2.6005
R2392 VSS.n3703 VSS.n3702 2.6005
R2393 VSS.n3701 VSS.n3700 2.6005
R2394 VSS.n3699 VSS.n3698 2.6005
R2395 VSS.n3697 VSS.n3696 2.6005
R2396 VSS.n3695 VSS.n3694 2.6005
R2397 VSS.n3693 VSS.n3692 2.6005
R2398 VSS.n3691 VSS.n3690 2.6005
R2399 VSS.n3689 VSS.n3688 2.6005
R2400 VSS.n3687 VSS.n3686 2.6005
R2401 VSS.n3685 VSS.n3684 2.6005
R2402 VSS.n3683 VSS.n3682 2.6005
R2403 VSS.n3681 VSS.n3680 2.6005
R2404 VSS.n3679 VSS.n3678 2.6005
R2405 VSS.n3677 VSS.n3676 2.6005
R2406 VSS.n3764 VSS.n3763 2.6005
R2407 VSS.n3331 VSS.n3330 2.6005
R2408 VSS.n3330 VSS.n3329 2.6005
R2409 VSS.n3328 VSS.n3327 2.6005
R2410 VSS.n3327 VSS.n3326 2.6005
R2411 VSS.n3325 VSS.n3324 2.6005
R2412 VSS.n3324 VSS.n3323 2.6005
R2413 VSS.n3322 VSS.n3321 2.6005
R2414 VSS.n3321 VSS.n3320 2.6005
R2415 VSS.n3318 VSS.n3317 2.6005
R2416 VSS.n3317 VSS.n3316 2.6005
R2417 VSS.n3315 VSS.n3314 2.6005
R2418 VSS.n3314 VSS.n3313 2.6005
R2419 VSS.n3311 VSS.n3310 2.6005
R2420 VSS.n3310 VSS.n3309 2.6005
R2421 VSS.n3308 VSS.n3307 2.6005
R2422 VSS.n3307 VSS.n3306 2.6005
R2423 VSS.n3305 VSS.n3304 2.6005
R2424 VSS.n3304 VSS.n3303 2.6005
R2425 VSS.n3302 VSS.n3301 2.6005
R2426 VSS.n3301 VSS.n3300 2.6005
R2427 VSS.n3299 VSS.n3298 2.6005
R2428 VSS.n3298 VSS.n3297 2.6005
R2429 VSS.n3296 VSS.n3295 2.6005
R2430 VSS.n3295 VSS.n3294 2.6005
R2431 VSS.n3293 VSS.n3292 2.6005
R2432 VSS.n3292 VSS.n3291 2.6005
R2433 VSS.n3290 VSS.n3289 2.6005
R2434 VSS.n3289 VSS.n3288 2.6005
R2435 VSS.n3287 VSS.n3286 2.6005
R2436 VSS.n3286 VSS.n3285 2.6005
R2437 VSS.n3284 VSS.n3283 2.6005
R2438 VSS.n3283 VSS.n3282 2.6005
R2439 VSS.n3495 VSS.n3494 2.6005
R2440 VSS.n3494 VSS.n3493 2.6005
R2441 VSS.n3498 VSS.n3497 2.6005
R2442 VSS.n3497 VSS.n3496 2.6005
R2443 VSS.n3501 VSS.n3500 2.6005
R2444 VSS.n3500 VSS.n3499 2.6005
R2445 VSS.n3504 VSS.n3503 2.6005
R2446 VSS.n3503 VSS.n3502 2.6005
R2447 VSS.n3507 VSS.n3506 2.6005
R2448 VSS.n3506 VSS.n3505 2.6005
R2449 VSS.n3510 VSS.n3509 2.6005
R2450 VSS.n3509 VSS.n3508 2.6005
R2451 VSS.n3513 VSS.n3512 2.6005
R2452 VSS.n3512 VSS.n3511 2.6005
R2453 VSS.n3516 VSS.n3515 2.6005
R2454 VSS.n3515 VSS.n3514 2.6005
R2455 VSS.n3519 VSS.n3518 2.6005
R2456 VSS.n3518 VSS.n3517 2.6005
R2457 VSS.n3522 VSS.n3521 2.6005
R2458 VSS.n3521 VSS.n3520 2.6005
R2459 VSS.n3526 VSS.n3525 2.6005
R2460 VSS.n3525 VSS.n3524 2.6005
R2461 VSS.n3529 VSS.n3528 2.6005
R2462 VSS.n3528 VSS.n3527 2.6005
R2463 VSS.n3533 VSS.n3532 2.6005
R2464 VSS.n3532 VSS.n3531 2.6005
R2465 VSS.n3536 VSS.n3535 2.6005
R2466 VSS.n3535 VSS.n3534 2.6005
R2467 VSS.n3539 VSS.n3538 2.6005
R2468 VSS.n3538 VSS.n3537 2.6005
R2469 VSS.n3542 VSS.n3541 2.6005
R2470 VSS.n3541 VSS.n3540 2.6005
R2471 VSS.n3267 VSS.n3266 2.6005
R2472 VSS.n2158 VSS.n2157 2.6005
R2473 VSS.n2258 VSS.n2257 2.6005
R2474 VSS.n2094 VSS.n2093 2.6005
R2475 VSS.n2097 VSS.n2096 2.6005
R2476 VSS.n2099 VSS.n2098 2.6005
R2477 VSS.n2102 VSS.n2101 2.6005
R2478 VSS.n2104 VSS.n2103 2.6005
R2479 VSS.n2107 VSS.n2106 2.6005
R2480 VSS.n2109 VSS.n2108 2.6005
R2481 VSS.n2111 VSS.n2110 2.6005
R2482 VSS.n2113 VSS.n2112 2.6005
R2483 VSS.n2115 VSS.n2114 2.6005
R2484 VSS.n2117 VSS.n2116 2.6005
R2485 VSS.n2119 VSS.n2118 2.6005
R2486 VSS.n2121 VSS.n2120 2.6005
R2487 VSS.n2123 VSS.n2122 2.6005
R2488 VSS.n2126 VSS.n2125 2.6005
R2489 VSS.n2128 VSS.n2127 2.6005
R2490 VSS.n2130 VSS.n2129 2.6005
R2491 VSS.n2132 VSS.n2131 2.6005
R2492 VSS.n2134 VSS.n2133 2.6005
R2493 VSS.n2136 VSS.n2135 2.6005
R2494 VSS.n2138 VSS.n2137 2.6005
R2495 VSS.n2141 VSS.n2140 2.6005
R2496 VSS.n2143 VSS.n2142 2.6005
R2497 VSS.n2145 VSS.n2144 2.6005
R2498 VSS.n2147 VSS.n2146 2.6005
R2499 VSS.n2150 VSS.n2149 2.6005
R2500 VSS.n2152 VSS.n2151 2.6005
R2501 VSS.n2155 VSS.n2154 2.6005
R2502 VSS.n2164 VSS.n2163 2.6005
R2503 VSS.n2166 VSS.n2165 2.6005
R2504 VSS.n2168 VSS.n2167 2.6005
R2505 VSS.n2170 VSS.n2169 2.6005
R2506 VSS.n2172 VSS.n2171 2.6005
R2507 VSS.n2174 VSS.n2173 2.6005
R2508 VSS.n2176 VSS.n2175 2.6005
R2509 VSS.n2178 VSS.n2177 2.6005
R2510 VSS.n2180 VSS.n2179 2.6005
R2511 VSS.n2182 VSS.n2181 2.6005
R2512 VSS.n2184 VSS.n2183 2.6005
R2513 VSS.n2186 VSS.n2185 2.6005
R2514 VSS.n2188 VSS.n2187 2.6005
R2515 VSS.n2190 VSS.n2189 2.6005
R2516 VSS.n2192 VSS.n2191 2.6005
R2517 VSS.n2194 VSS.n2193 2.6005
R2518 VSS.n2196 VSS.n2195 2.6005
R2519 VSS.n2198 VSS.n2197 2.6005
R2520 VSS.n2200 VSS.n2199 2.6005
R2521 VSS.n2202 VSS.n2201 2.6005
R2522 VSS.n2204 VSS.n2203 2.6005
R2523 VSS.n2206 VSS.n2205 2.6005
R2524 VSS.n2208 VSS.n2207 2.6005
R2525 VSS.n2210 VSS.n2209 2.6005
R2526 VSS.n2212 VSS.n2211 2.6005
R2527 VSS.n2214 VSS.n2213 2.6005
R2528 VSS.n2216 VSS.n2215 2.6005
R2529 VSS.n2218 VSS.n2217 2.6005
R2530 VSS.n2221 VSS.n2220 2.6005
R2531 VSS.n2223 VSS.n2222 2.6005
R2532 VSS.n2226 VSS.n2225 2.6005
R2533 VSS.n2228 VSS.n2227 2.6005
R2534 VSS.n2231 VSS.n2230 2.6005
R2535 VSS.n2233 VSS.n2232 2.6005
R2536 VSS.n2236 VSS.n2235 2.6005
R2537 VSS.n2238 VSS.n2237 2.6005
R2538 VSS.n2241 VSS.n2240 2.6005
R2539 VSS.n2162 VSS.n2161 2.6005
R2540 VSS.n2160 VSS.n2159 2.6005
R2541 VSS.n3381 VSS.n2242 2.6005
R2542 VSS.n117 VSS.n116 2.6005
R2543 VSS.n115 VSS.n114 2.6005
R2544 VSS.n112 VSS.n111 2.6005
R2545 VSS.n109 VSS.n108 2.6005
R2546 VSS.n107 VSS.n106 2.6005
R2547 VSS.n105 VSS.n104 2.6005
R2548 VSS.n102 VSS.n101 2.6005
R2549 VSS.n100 VSS.n99 2.6005
R2550 VSS.n98 VSS.n97 2.6005
R2551 VSS.n96 VSS.n95 2.6005
R2552 VSS.n93 VSS.n92 2.6005
R2553 VSS.n91 VSS.n90 2.6005
R2554 VSS.n89 VSS.n88 2.6005
R2555 VSS.n86 VSS.n85 2.6005
R2556 VSS.n84 VSS.n83 2.6005
R2557 VSS.n82 VSS.n81 2.6005
R2558 VSS.n80 VSS.n79 2.6005
R2559 VSS.n77 VSS.n76 2.6005
R2560 VSS.n75 VSS.n74 2.6005
R2561 VSS.n73 VSS.n72 2.6005
R2562 VSS.n67 VSS.n66 2.6005
R2563 VSS.n64 VSS.n63 2.6005
R2564 VSS.n62 VSS.n61 2.6005
R2565 VSS.n3982 VSS.n3981 2.6005
R2566 VSS.n2365 VSS.n2364 2.6005
R2567 VSS.n2364 VSS.n2363 2.6005
R2568 VSS.n2369 VSS.n2368 2.6005
R2569 VSS.n2368 VSS.n2367 2.6005
R2570 VSS.n2372 VSS.n2371 2.6005
R2571 VSS.n2371 VSS.n2370 2.6005
R2572 VSS.n2382 VSS.n2381 2.6005
R2573 VSS.n2381 VSS.n2380 2.6005
R2574 VSS.n2385 VSS.n2384 2.6005
R2575 VSS.n2384 VSS.n2383 2.6005
R2576 VSS.n2388 VSS.n2387 2.6005
R2577 VSS.n2387 VSS.n2386 2.6005
R2578 VSS.n2391 VSS.n2390 2.6005
R2579 VSS.n2390 VSS.n2389 2.6005
R2580 VSS.n2394 VSS.n2393 2.6005
R2581 VSS.n2393 VSS.n2392 2.6005
R2582 VSS.n2397 VSS.n2396 2.6005
R2583 VSS.n2396 VSS.n2395 2.6005
R2584 VSS.n2400 VSS.n2399 2.6005
R2585 VSS.n2399 VSS.n2398 2.6005
R2586 VSS.n2403 VSS.n2402 2.6005
R2587 VSS.n2402 VSS.n2401 2.6005
R2588 VSS.n2406 VSS.n2405 2.6005
R2589 VSS.n2405 VSS.n2404 2.6005
R2590 VSS.n2410 VSS.n2409 2.6005
R2591 VSS.n2409 VSS.n2408 2.6005
R2592 VSS.n3337 VSS.n3336 2.6005
R2593 VSS.n3336 VSS.n3335 2.6005
R2594 VSS.n3340 VSS.n3339 2.6005
R2595 VSS.n3339 VSS.n3338 2.6005
R2596 VSS.n3343 VSS.n3342 2.6005
R2597 VSS.n3342 VSS.n3341 2.6005
R2598 VSS.n3346 VSS.n3345 2.6005
R2599 VSS.n3345 VSS.n3344 2.6005
R2600 VSS.n3349 VSS.n3348 2.6005
R2601 VSS.n3348 VSS.n3347 2.6005
R2602 VSS.n3352 VSS.n3351 2.6005
R2603 VSS.n3351 VSS.n3350 2.6005
R2604 VSS.n3355 VSS.n3354 2.6005
R2605 VSS.n3354 VSS.n3353 2.6005
R2606 VSS.n3358 VSS.n3357 2.6005
R2607 VSS.n3357 VSS.n3356 2.6005
R2608 VSS.n3361 VSS.n3360 2.6005
R2609 VSS.n3360 VSS.n3359 2.6005
R2610 VSS.n3364 VSS.n3363 2.6005
R2611 VSS.n3363 VSS.n3362 2.6005
R2612 VSS.n3367 VSS.n3366 2.6005
R2613 VSS.n3366 VSS.n3365 2.6005
R2614 VSS.n3370 VSS.n3369 2.6005
R2615 VSS.n3369 VSS.n3368 2.6005
R2616 VSS.n3374 VSS.n3373 2.6005
R2617 VSS.n3373 VSS.n3372 2.6005
R2618 VSS.n3378 VSS.n3377 2.6005
R2619 VSS.n3377 VSS.n3376 2.6005
R2620 VSS.n3424 VSS.n3380 2.6005
R2621 VSS.n3424 VSS.n3423 2.6005
R2622 VSS.n4067 VSS.n4066 2.6005
R2623 VSS.n4066 VSS.n4065 2.6005
R2624 VSS.n4064 VSS.n4063 2.6005
R2625 VSS.n4063 VSS.n4062 2.6005
R2626 VSS.n4060 VSS.n4059 2.6005
R2627 VSS.n4059 VSS.n4058 2.6005
R2628 VSS.n4050 VSS.n4049 2.6005
R2629 VSS.n4049 VSS.n4048 2.6005
R2630 VSS.n4047 VSS.n4046 2.6005
R2631 VSS.n4046 VSS.n4045 2.6005
R2632 VSS.n4044 VSS.n4043 2.6005
R2633 VSS.n4043 VSS.n4042 2.6005
R2634 VSS.n4040 VSS.n4039 2.6005
R2635 VSS.n4039 VSS.n4038 2.6005
R2636 VSS.n4037 VSS.n4036 2.6005
R2637 VSS.n4036 VSS.n4035 2.6005
R2638 VSS.n4034 VSS.n4033 2.6005
R2639 VSS.n4033 VSS.n4032 2.6005
R2640 VSS.n4031 VSS.n4030 2.6005
R2641 VSS.n4030 VSS.n4029 2.6005
R2642 VSS.n4027 VSS.n4026 2.6005
R2643 VSS.n4026 VSS.n4025 2.6005
R2644 VSS.n4024 VSS.n4023 2.6005
R2645 VSS.n4023 VSS.n4022 2.6005
R2646 VSS.n4021 VSS.n4020 2.6005
R2647 VSS.n4020 VSS.n4019 2.6005
R2648 VSS.n4017 VSS.n4016 2.6005
R2649 VSS.n4016 VSS.n4015 2.6005
R2650 VSS.n4014 VSS.n4013 2.6005
R2651 VSS.n4013 VSS.n4012 2.6005
R2652 VSS.n4011 VSS.n4010 2.6005
R2653 VSS.n4010 VSS.n4009 2.6005
R2654 VSS.n4007 VSS.n4006 2.6005
R2655 VSS.n4006 VSS.n4005 2.6005
R2656 VSS.n4002 VSS.n4001 2.6005
R2657 VSS.n4001 VSS.n4000 2.6005
R2658 VSS.n3999 VSS.n3998 2.6005
R2659 VSS.n3998 VSS.n3997 2.6005
R2660 VSS.n3996 VSS.n3995 2.6005
R2661 VSS.n3995 VSS.n3994 2.6005
R2662 VSS.n3992 VSS.n3991 2.6005
R2663 VSS.n3991 VSS.n3990 2.6005
R2664 VSS.n3988 VSS.n3987 2.6005
R2665 VSS.n3987 VSS.n3986 2.6005
R2666 VSS.n3985 VSS.n3984 2.6005
R2667 VSS.n3984 VSS.n3983 2.6005
R2668 VSS.n2362 VSS.n2361 2.6005
R2669 VSS.n2590 VSS.n2589 2.49533
R2670 VSS.n2891 VSS.n2890 2.43319
R2671 VSS.n2888 VSS.n2887 2.43319
R2672 VSS.n2885 VSS.n2884 2.43319
R2673 VSS.n2605 VSS.n2604 2.43319
R2674 VSS.n2608 VSS.n2607 2.43319
R2675 VSS.n2611 VSS.n2610 2.43319
R2676 VSS.n2539 VSS.n2538 2.43319
R2677 VSS.n2536 VSS.n2535 2.43319
R2678 VSS.n2542 VSS.n2541 2.43319
R2679 VSS.n1629 VSS.n1626 2.29321
R2680 VSS.n1497 VSS.n1494 2.29321
R2681 VSS.n1365 VSS.n1362 2.29321
R2682 VSS.n3313 VSS.t398 2.24467
R2683 VSS.n3297 VSS.t683 2.24467
R2684 VSS.n3505 VSS.t657 2.24467
R2685 VSS.n3527 VSS.t659 2.24467
R2686 VSS.n1275 VSS.n1273 2.18289
R2687 VSS.n1113 VSS.n1111 2.18289
R2688 VSS.n952 VSS.n950 2.18289
R2689 VSS.n3018 VSS.n3015 2.18289
R2690 VSS.n2590 VSS.n2587 2.18289
R2691 VSS.n2049 VSS.n2048 2.08372
R2692 VSS.n2576 VSS.n2572 2.07475
R2693 VSS.n2556 VSS.n2552 2.07475
R2694 VSS.n1630 VSS.n1629 1.9805
R2695 VSS.n1498 VSS.n1497 1.9805
R2696 VSS.n1366 VSS.n1365 1.9805
R2697 VSS.n1584 VSS.n1581 1.96158
R2698 VSS.n1604 VSS.n1601 1.96158
R2699 VSS.n1452 VSS.n1449 1.96158
R2700 VSS.n1472 VSS.n1469 1.96158
R2701 VSS.n1320 VSS.n1317 1.96158
R2702 VSS.n1340 VSS.n1337 1.96158
R2703 VSS.n1609 VSS.n1608 1.95148
R2704 VSS.n1477 VSS.n1476 1.95148
R2705 VSS.n1345 VSS.n1344 1.95148
R2706 VSS.n1640 VSS.n1639 1.91002
R2707 VSS.n1616 VSS.n1615 1.91002
R2708 VSS.n1508 VSS.n1507 1.91002
R2709 VSS.n1484 VSS.n1483 1.91002
R2710 VSS.n1376 VSS.n1375 1.91002
R2711 VSS.n1352 VSS.n1351 1.91002
R2712 VSS.n1645 VSS.n1642 1.90218
R2713 VSS.n1513 VSS.n1510 1.90218
R2714 VSS.n1381 VSS.n1378 1.90218
R2715 VSS.n1610 VSS.n1609 1.89955
R2716 VSS.n1478 VSS.n1477 1.89955
R2717 VSS.n1346 VSS.n1345 1.89955
R2718 VSS.n679 VSS.n678 1.8318
R2719 VSS.n1556 VSS.n1555 1.8318
R2720 VSS.n685 VSS.n684 1.8318
R2721 VSS.n1562 VSS.n1561 1.8318
R2722 VSS.n422 VSS.n421 1.8318
R2723 VSS.n1520 VSS.n1519 1.8318
R2724 VSS.n428 VSS.n427 1.8318
R2725 VSS.n1526 VSS.n1525 1.8318
R2726 VSS.n412 VSS.n411 1.8318
R2727 VSS.n1424 VSS.n1423 1.8318
R2728 VSS.n418 VSS.n417 1.8318
R2729 VSS.n1430 VSS.n1429 1.8318
R2730 VSS.n155 VSS.n154 1.8318
R2731 VSS.n1388 VSS.n1387 1.8318
R2732 VSS.n161 VSS.n160 1.8318
R2733 VSS.n1394 VSS.n1393 1.8318
R2734 VSS.n145 VSS.n144 1.8318
R2735 VSS.n1292 VSS.n1291 1.8318
R2736 VSS.n151 VSS.n150 1.8318
R2737 VSS.n1298 VSS.n1297 1.8318
R2738 VSS.n695 VSS.n694 1.8318
R2739 VSS.n1687 VSS.n1686 1.8318
R2740 VSS.n689 VSS.n688 1.8318
R2741 VSS.n1654 VSS.n1653 1.8318
R2742 VSS.n3375 VSS.t211 1.79583
R2743 VSS.n3288 VSS.t6 1.79583
R2744 VSS.t680 VSS.t203 1.79583
R2745 VSS.n1648 VSS.n1647 1.76495
R2746 VSS.n1516 VSS.n1515 1.76495
R2747 VSS.n1384 VSS.n1383 1.76495
R2748 VSS.n49 VSS.n48 1.68702
R2749 VSS.n48 VSS.n47 1.68702
R2750 VSS.n3791 VSS.n3790 1.68702
R2751 VSS.n3792 VSS.n3791 1.68702
R2752 VSS.n3793 VSS.n3792 1.68702
R2753 VSS.n19 VSS.n18 1.68702
R2754 VSS.n18 VSS.n17 1.68702
R2755 VSS.n3439 VSS.n3436 1.68702
R2756 VSS.n3442 VSS.n3439 1.68702
R2757 VSS.n3445 VSS.n3442 1.68702
R2758 VSS.n3448 VSS.n3445 1.68702
R2759 VSS.n28 VSS.n27 1.68702
R2760 VSS.n27 VSS.n26 1.68702
R2761 VSS.n3454 VSS.n3451 1.68702
R2762 VSS.n3457 VSS.n3454 1.68702
R2763 VSS.n3460 VSS.n3457 1.68702
R2764 VSS.n3463 VSS.n3460 1.68702
R2765 VSS.n37 VSS.n36 1.68702
R2766 VSS.n36 VSS.n35 1.68702
R2767 VSS.n3469 VSS.n3466 1.68702
R2768 VSS.n3472 VSS.n3469 1.68702
R2769 VSS.n3475 VSS.n3472 1.68702
R2770 VSS.n3478 VSS.n3475 1.68702
R2771 VSS.n2244 VSS.n2243 1.68702
R2772 VSS.n2250 VSS.n2249 1.68702
R2773 VSS.n46 VSS.n45 1.68702
R2774 VSS.n45 VSS.n44 1.68702
R2775 VSS.n3772 VSS.n3769 1.68702
R2776 VSS.n3775 VSS.n3772 1.68702
R2777 VSS.n3778 VSS.n3775 1.68702
R2778 VSS.n3781 VSS.n3778 1.68702
R2779 VSS.n2374 VSS.n2373 1.68702
R2780 VSS.n2254 VSS.n2253 1.68702
R2781 VSS.n10 VSS.n9 1.68702
R2782 VSS.n9 VSS.n8 1.68702
R2783 VSS.n4052 VSS.n4051 1.68702
R2784 VSS.n4053 VSS.n4052 1.68702
R2785 VSS.n4054 VSS.n4053 1.68702
R2786 VSS.n7 VSS.n6 1.68702
R2787 VSS.n6 VSS.n5 1.68702
R2788 VSS.n3429 VSS.n3428 1.68702
R2789 VSS.n3430 VSS.n3429 1.68702
R2790 VSS.n3431 VSS.n3430 1.68702
R2791 VSS.n70 VSS.n69 1.68702
R2792 VSS.n69 VSS.n68 1.68702
R2793 VSS.n3783 VSS.n3782 1.68702
R2794 VSS.n3784 VSS.n3783 1.68702
R2795 VSS.n3785 VSS.n3784 1.68702
R2796 VSS.n3634 VSS.n3633 1.65879
R2797 VSS.n3629 VSS.n3628 1.65879
R2798 VSS.n3624 VSS.n3623 1.65879
R2799 VSS.n3619 VSS.n3618 1.65879
R2800 VSS.n3614 VSS.n3613 1.65879
R2801 VSS.n3609 VSS.n3608 1.65879
R2802 VSS.n2462 VSS.n2461 1.65879
R2803 VSS.n2457 VSS.n2456 1.65879
R2804 VSS.n2452 VSS.n2451 1.65879
R2805 VSS.n3973 VSS.n3971 1.65879
R2806 VSS.n3970 VSS.n3968 1.65879
R2807 VSS.n3967 VSS.n3965 1.65879
R2808 VSS.n3964 VSS.n3962 1.65879
R2809 VSS.n3961 VSS.n3959 1.65879
R2810 VSS.n3958 VSS.n3956 1.65879
R2811 VSS.n3955 VSS.n3953 1.65879
R2812 VSS.n3952 VSS.n3950 1.65879
R2813 VSS.n3949 VSS.n3947 1.65879
R2814 VSS.n3946 VSS.n3945 1.65879
R2815 VSS.n2019 VSS.n2018 1.65879
R2816 VSS.n2014 VSS.n2013 1.65879
R2817 VSS.n2009 VSS.n2008 1.65879
R2818 VSS.n2004 VSS.n2003 1.65879
R2819 VSS.n1999 VSS.n1998 1.65879
R2820 VSS.n1994 VSS.n1993 1.65879
R2821 VSS.n1989 VSS.n1988 1.65879
R2822 VSS.n1984 VSS.n1983 1.65879
R2823 VSS.n1979 VSS.n1978 1.65879
R2824 VSS.n404 VSS.n403 1.65879
R2825 VSS.n399 VSS.n398 1.65879
R2826 VSS.n394 VSS.n393 1.65879
R2827 VSS.n389 VSS.n388 1.65879
R2828 VSS.n384 VSS.n383 1.65879
R2829 VSS.n379 VSS.n378 1.65879
R2830 VSS.n374 VSS.n373 1.65879
R2831 VSS.n369 VSS.n368 1.65879
R2832 VSS.n364 VSS.n363 1.65879
R2833 VSS.n359 VSS.n358 1.65879
R2834 VSS.n354 VSS.n353 1.65879
R2835 VSS.n671 VSS.n670 1.65879
R2836 VSS.n666 VSS.n665 1.65879
R2837 VSS.n661 VSS.n660 1.65879
R2838 VSS.n656 VSS.n655 1.65879
R2839 VSS.n651 VSS.n650 1.65879
R2840 VSS.n646 VSS.n645 1.65879
R2841 VSS.n641 VSS.n640 1.65879
R2842 VSS.n636 VSS.n635 1.65879
R2843 VSS.n631 VSS.n630 1.65879
R2844 VSS.n626 VSS.n625 1.65879
R2845 VSS.n621 VSS.n620 1.65879
R2846 VSS.n2742 VSS.n2740 1.65879
R2847 VSS.n3255 VSS.n3254 1.65879
R2848 VSS.n3250 VSS.n3249 1.65879
R2849 VSS.n3245 VSS.n3244 1.65879
R2850 VSS.n3240 VSS.n3239 1.65879
R2851 VSS.n3235 VSS.n3234 1.65879
R2852 VSS.n3230 VSS.n3229 1.65879
R2853 VSS.n3225 VSS.n3224 1.65879
R2854 VSS.n3220 VSS.n3219 1.65879
R2855 VSS.n3748 VSS.n3747 1.65879
R2856 VSS.n3743 VSS.n3742 1.65879
R2857 VSS.n3738 VSS.n3737 1.65879
R2858 VSS.n3733 VSS.n3732 1.65879
R2859 VSS.n3728 VSS.n3727 1.65879
R2860 VSS.n3723 VSS.n3722 1.65879
R2861 VSS.n3718 VSS.n3717 1.65879
R2862 VSS.n3713 VSS.n3712 1.65879
R2863 VSS.n2738 VSS.n2737 1.65822
R2864 VSS.n2320 VSS.n2319 1.65822
R2865 VSS.n2325 VSS.n2324 1.65822
R2866 VSS.n2330 VSS.n2329 1.65822
R2867 VSS.n2335 VSS.n2334 1.65822
R2868 VSS.n2340 VSS.n2339 1.65822
R2869 VSS.n3979 VSS.n3978 1.65822
R2870 VSS.n3920 VSS.n3919 1.65822
R2871 VSS.n3915 VSS.n3914 1.65822
R2872 VSS.n3910 VSS.n3909 1.65822
R2873 VSS.n3905 VSS.n3904 1.65822
R2874 VSS.n3900 VSS.n3899 1.65822
R2875 VSS.n3895 VSS.n3894 1.65822
R2876 VSS.n3949 VSS.n3948 1.65822
R2877 VSS.n3952 VSS.n3951 1.65822
R2878 VSS.n3955 VSS.n3954 1.65822
R2879 VSS.n3958 VSS.n3957 1.65822
R2880 VSS.n3961 VSS.n3960 1.65822
R2881 VSS.n3964 VSS.n3963 1.65822
R2882 VSS.n3967 VSS.n3966 1.65822
R2883 VSS.n3970 VSS.n3969 1.65822
R2884 VSS.n3973 VSS.n3972 1.65822
R2885 VSS.n1286 VSS.n1285 1.65822
R2886 VSS.n3034 VSS.n3033 1.65822
R2887 VSS.n3029 VSS.n3028 1.65822
R2888 VSS.n3212 VSS.n3211 1.65822
R2889 VSS.n2220 VSS.n2219 1.65811
R2890 VSS.n2225 VSS.n2224 1.65811
R2891 VSS.n2230 VSS.n2229 1.65811
R2892 VSS.n2235 VSS.n2234 1.65811
R2893 VSS.n2240 VSS.n2239 1.65811
R2894 VSS.n4 VSS.n3 1.65811
R2895 VSS.n3418 VSS.n3416 1.65811
R2896 VSS.n3415 VSS.n3413 1.65811
R2897 VSS.n3412 VSS.n3411 1.65811
R2898 VSS.n3415 VSS.n3414 1.65811
R2899 VSS.n3418 VSS.n3417 1.65811
R2900 VSS.n257 VSS.n256 1.65811
R2901 VSS.n262 VSS.n261 1.65811
R2902 VSS.n267 VSS.n266 1.65811
R2903 VSS.n272 VSS.n271 1.65811
R2904 VSS.n277 VSS.n276 1.65811
R2905 VSS.n282 VSS.n281 1.65811
R2906 VSS.n524 VSS.n523 1.65811
R2907 VSS.n529 VSS.n528 1.65811
R2908 VSS.n534 VSS.n533 1.65811
R2909 VSS.n539 VSS.n538 1.65811
R2910 VSS.n544 VSS.n543 1.65811
R2911 VSS.n549 VSS.n548 1.65811
R2912 VSS.n816 VSS.n815 1.65811
R2913 VSS.n811 VSS.n810 1.65811
R2914 VSS.n806 VSS.n805 1.65811
R2915 VSS.n801 VSS.n800 1.65811
R2916 VSS.n796 VSS.n795 1.65811
R2917 VSS.n791 VSS.n790 1.65811
R2918 VSS.n3216 VSS.n3215 1.65811
R2919 VSS.n2876 VSS.n2875 1.65811
R2920 VSS.n2860 VSS.n2859 1.65811
R2921 VSS.n2855 VSS.n2854 1.65811
R2922 VSS.n2850 VSS.n2849 1.65811
R2923 VSS.n2845 VSS.n2844 1.65811
R2924 VSS.n2744 VSS.t423 1.6385
R2925 VSS.n2412 VSS.t454 1.6385
R2926 VSS.n2412 VSS.n2411 1.6385
R2927 VSS.n2422 VSS.t614 1.6385
R2928 VSS.n2422 VSS.n2421 1.6385
R2929 VSS.n2424 VSS.t206 1.6385
R2930 VSS.n2424 VSS.n2423 1.6385
R2931 VSS.n2426 VSS.t248 1.6385
R2932 VSS.n2426 VSS.n2425 1.6385
R2933 VSS.n2428 VSS.t282 1.6385
R2934 VSS.n2428 VSS.n2427 1.6385
R2935 VSS.n2430 VSS.t204 1.6385
R2936 VSS.n2430 VSS.n2429 1.6385
R2937 VSS.n2432 VSS.t236 1.6385
R2938 VSS.n2432 VSS.n2431 1.6385
R2939 VSS.n2434 VSS.t274 1.6385
R2940 VSS.n2434 VSS.n2433 1.6385
R2941 VSS.n2436 VSS.t295 1.6385
R2942 VSS.n2436 VSS.n2435 1.6385
R2943 VSS.n2746 VSS.t523 1.6385
R2944 VSS.n2747 VSS.t483 1.6385
R2945 VSS.n2748 VSS.t578 1.6385
R2946 VSS.n2749 VSS.t530 1.6385
R2947 VSS.n2751 VSS.t387 1.6385
R2948 VSS.n2751 VSS.n2750 1.6385
R2949 VSS.n2753 VSS.t658 1.6385
R2950 VSS.n2753 VSS.n2752 1.6385
R2951 VSS.n3555 VSS.t663 1.6385
R2952 VSS.n3555 VSS.n3554 1.6385
R2953 VSS.n3553 VSS.t52 1.6385
R2954 VSS.n3553 VSS.n3552 1.6385
R2955 VSS.n3551 VSS.t50 1.6385
R2956 VSS.n3551 VSS.n3550 1.6385
R2957 VSS.n4042 VSS.t164 1.53424
R2958 VSS.n4000 VSS.t159 1.53424
R2959 VSS.n1581 VSS.n1580 1.48796
R2960 VSS.n1569 VSS.n1568 1.48796
R2961 VSS.n1601 VSS.n1600 1.48796
R2962 VSS.n1589 VSS.n1588 1.48796
R2963 VSS.n1449 VSS.n1448 1.48796
R2964 VSS.n1437 VSS.n1436 1.48796
R2965 VSS.n1469 VSS.n1468 1.48796
R2966 VSS.n1457 VSS.n1456 1.48796
R2967 VSS.n1317 VSS.n1316 1.48796
R2968 VSS.n1305 VSS.n1304 1.48796
R2969 VSS.n1337 VSS.n1336 1.48796
R2970 VSS.n1325 VSS.n1324 1.48796
R2971 VSS.n1573 VSS.n1572 1.47979
R2972 VSS.n1593 VSS.n1592 1.47979
R2973 VSS.n1613 VSS.n1612 1.47979
R2974 VSS.n1622 VSS.n1621 1.47979
R2975 VSS.n1637 VSS.n1636 1.47979
R2976 VSS.n1441 VSS.n1440 1.47979
R2977 VSS.n1481 VSS.n1480 1.47979
R2978 VSS.n1490 VSS.n1489 1.47979
R2979 VSS.n1505 VSS.n1504 1.47979
R2980 VSS.n1461 VSS.n1460 1.47979
R2981 VSS.n1309 VSS.n1308 1.47979
R2982 VSS.n1329 VSS.n1328 1.47979
R2983 VSS.n1349 VSS.n1348 1.47979
R2984 VSS.n1358 VSS.n1357 1.47979
R2985 VSS.n1373 VSS.n1372 1.47979
R2986 VSS.n3604 VSS.n3603 1.40389
R2987 VSS.n2894 VSS.n2893 1.40389
R2988 VSS.n674 VSS.n673 1.40375
R2989 VSS.n407 VSS.n406 1.40375
R2990 VSS.n1281 VSS.n1280 1.40375
R2991 VSS.n2880 VSS.n2879 1.40375
R2992 VSS.n2614 VSS.n2613 1.40375
R2993 VSS.n3021 VSS.n3020 1.40375
R2994 VSS.n2585 VSS.n2584 1.40375
R2995 VSS.n2525 VSS.n2524 1.40375
R2996 VSS.n2519 VSS.n2518 1.40375
R2997 VSS.n2510 VSS.n2509 1.40375
R2998 VSS.n2044 VSS.n2024 1.38491
R2999 VSS.n1135 VSS.n1114 1.38491
R3000 VSS.n974 VSS.n953 1.38491
R3001 VSS.n3264 VSS.n3259 1.38491
R3002 VSS.n3264 VSS.n3260 1.38491
R3003 VSS.n3264 VSS.n3261 1.38491
R3004 VSS.n3264 VSS.n3262 1.38491
R3005 VSS.n3264 VSS.n3263 1.38491
R3006 VSS.n1570 VSS.n1569 1.3649
R3007 VSS.n1590 VSS.n1589 1.3649
R3008 VSS.n1438 VSS.n1437 1.3649
R3009 VSS.n1458 VSS.n1457 1.3649
R3010 VSS.n1306 VSS.n1305 1.3649
R3011 VSS.n1326 VSS.n1325 1.3649
R3012 VSS.n3976 VSS.n3974 1.3543
R3013 VSS.n3210 VSS.n3208 1.3543
R3014 VSS.n1170 VSS.n1140 1.35379
R3015 VSS.n1009 VSS.n979 1.35379
R3016 VSS.n848 VSS.n818 1.35379
R3017 VSS.n3210 VSS.n3209 1.35379
R3018 VSS.n3640 VSS.n3639 1.35379
R3019 VSS.n3763 VSS.n3762 1.35379
R3020 VSS.n3266 VSS.n3265 1.35379
R3021 VSS.n3976 VSS.n3975 1.35379
R3022 VSS.n2361 VSS.n2360 1.35379
R3023 VSS.n3420 VSS.n3419 1.35364
R3024 VSS.n3425 VSS.n3422 1.35364
R3025 VSS.n3422 VSS.n3381 1.35364
R3026 VSS.n3057 VSS.t346 1.347
R3027 VSS.n3132 VSS.t618 1.347
R3028 VSS.n2492 VSS.t607 1.347
R3029 VSS.n3671 VSS.t330 1.347
R3030 VSS.n881 VSS.t38 1.31284
R3031 VSS.n917 VSS.t7 1.31284
R3032 VSS.n1042 VSS.t101 1.31284
R3033 VSS.n1078 VSS.t93 1.31284
R3034 VSS.n1203 VSS.t22 1.31284
R3035 VSS.n1239 VSS.t13 1.31284
R3036 VSS.n3171 VSS.n2902 1.30746
R3037 VSS.n3160 VSS.n2908 1.30746
R3038 VSS.n3094 VSS.n2925 1.30746
R3039 VSS.n3072 VSS.n2930 1.30746
R3040 VSS.n1693 VSS.n1656 1.30746
R3041 VSS.n926 VSS.n687 1.30746
R3042 VSS.n930 VSS.n683 1.30746
R3043 VSS.n1729 VSS.n1564 1.30746
R3044 VSS.n1732 VSS.n1560 1.30746
R3045 VSS.n1031 VSS.n430 1.30746
R3046 VSS.n1035 VSS.n426 1.30746
R3047 VSS.n1766 VSS.n1528 1.30746
R3048 VSS.n1769 VSS.n1524 1.30746
R3049 VSS.n1087 VSS.n420 1.30746
R3050 VSS.n1091 VSS.n416 1.30746
R3051 VSS.n1805 VSS.n1432 1.30746
R3052 VSS.n1808 VSS.n1428 1.30746
R3053 VSS.n1192 VSS.n163 1.30746
R3054 VSS.n1196 VSS.n159 1.30746
R3055 VSS.n1842 VSS.n1396 1.30746
R3056 VSS.n1845 VSS.n1392 1.30746
R3057 VSS.n1248 VSS.n153 1.30746
R3058 VSS.n1252 VSS.n149 1.30746
R3059 VSS.n1881 VSS.n1300 1.30746
R3060 VSS.n1884 VSS.n1296 1.30746
R3061 VSS.n1690 VSS.n1689 1.30746
R3062 VSS.n874 VSS.n693 1.30746
R3063 VSS.n870 VSS.n697 1.30746
R3064 VSS.n3053 VSS.n2936 1.30746
R3065 VSS.n3043 VSS.n2938 1.30746
R3066 VSS.n2620 VSS.n2582 1.30746
R3067 VSS.n2627 VSS.n2580 1.30746
R3068 VSS.n3119 VSS.n2920 1.30746
R3069 VSS.n2672 VSS.n2566 1.30746
R3070 VSS.n3138 VSS.n2914 1.30746
R3071 VSS.n2685 VSS.n2563 1.30746
R3072 VSS.n3185 VSS.n2899 1.30746
R3073 VSS.n3175 VSS.n2901 1.30746
R3074 VSS.n2708 VSS.n2560 1.30746
R3075 VSS.n2715 VSS.n2558 1.30746
R3076 VSS.n1619 VSS.n1618 1.3055
R3077 VSS.n1487 VSS.n1486 1.3055
R3078 VSS.n1355 VSS.n1354 1.3055
R3079 VSS.n1631 VSS.n1630 1.29992
R3080 VSS.n1499 VSS.n1498 1.29992
R3081 VSS.n1367 VSS.n1366 1.29992
R3082 VSS.n3333 VSS.n3332 1.20652
R3083 VSS.n3766 VSS.n3765 1.20637
R3084 VSS.n2445 VSS.n2444 1.19007
R3085 VSS.n2444 VSS.n2443 1.19007
R3086 VSS.n3334 VSS.n3333 1.12775
R3087 VSS.n4008 VSS.n3766 1.12675
R3088 VSS.n1578 VSS.n1577 1.1255
R3089 VSS.n1598 VSS.n1597 1.1255
R3090 VSS.n1618 VSS.n1617 1.1255
R3091 VSS.n1633 VSS.n1632 1.1255
R3092 VSS.n1642 VSS.n1641 1.1255
R3093 VSS.n1446 VSS.n1445 1.1255
R3094 VSS.n1486 VSS.n1485 1.1255
R3095 VSS.n1501 VSS.n1500 1.1255
R3096 VSS.n1510 VSS.n1509 1.1255
R3097 VSS.n1466 VSS.n1465 1.1255
R3098 VSS.n1314 VSS.n1313 1.1255
R3099 VSS.n1334 VSS.n1333 1.1255
R3100 VSS.n1354 VSS.n1353 1.1255
R3101 VSS.n1369 VSS.n1368 1.1255
R3102 VSS.n1378 VSS.n1377 1.1255
R3103 VSS.n65 VSS.n49 1.12354
R3104 VSS.n103 VSS.n19 1.12354
R3105 VSS.n94 VSS.n28 1.12354
R3106 VSS.n87 VSS.n37 1.12354
R3107 VSS.n78 VSS.n46 1.12354
R3108 VSS.n110 VSS.n10 1.12354
R3109 VSS.n113 VSS.n7 1.12354
R3110 VSS.n71 VSS.n70 1.12354
R3111 VSS.n4061 VSS.n3433 1.12159
R3112 VSS.n4041 VSS.n3448 1.12159
R3113 VSS.n4028 VSS.n3463 1.12159
R3114 VSS.n4018 VSS.n3478 1.12159
R3115 VSS.n4057 VSS.n4056 1.12159
R3116 VSS.n3993 VSS.n3789 1.12159
R3117 VSS.n3989 VSS.n3795 1.12159
R3118 VSS.n4004 VSS.n3781 1.10202
R3119 VSS.n952 VSS.n951 1.09195
R3120 VSS.n1113 VSS.n1112 1.09195
R3121 VSS.n1275 VSS.n1274 1.09195
R3122 VSS.n1899 VSS.n1898 1.09195
R3123 VSS.n1824 VSS.n1823 1.09195
R3124 VSS.n1748 VSS.n1747 1.09195
R3125 VSS.n3599 VSS.n3598 1.09195
R3126 VSS.n3371 VSS.n2252 1.08441
R3127 VSS.n2153 VSS.n2089 1.08441
R3128 VSS.n3379 VSS.n2248 1.08441
R3129 VSS.n2148 VSS.n2090 1.08441
R3130 VSS.n2366 VSS.n2256 1.08441
R3131 VSS.n2100 VSS.n2091 1.08441
R3132 VSS.n2379 VSS.n2378 1.08441
R3133 VSS.n2095 VSS.n2092 1.08441
R3134 VSS.n2908 VSS.n2907 1.0492
R3135 VSS.n2936 VSS.n2935 1.0492
R3136 VSS.n2938 VSS.n2937 1.0492
R3137 VSS.n2920 VSS.n2919 1.0492
R3138 VSS.n2914 VSS.n2913 1.0492
R3139 VSS.n2899 VSS.n2898 1.0492
R3140 VSS.n2901 VSS.n2900 1.0492
R3141 VSS.n3486 VSS.n3485 1.0492
R3142 VSS.n3485 VSS.n3484 1.0492
R3143 VSS.n3484 VSS.n3483 1.0492
R3144 VSS.n3492 VSS.n3491 1.0492
R3145 VSS.n3491 VSS.n3490 1.0492
R3146 VSS.n3490 VSS.n3489 1.0492
R3147 VSS.n3281 VSS.n3280 1.0492
R3148 VSS.n3280 VSS.n3279 1.0492
R3149 VSS.n3279 VSS.n3278 1.0492
R3150 VSS.n3275 VSS.n3274 1.0492
R3151 VSS.n3274 VSS.n3273 1.0492
R3152 VSS.n3273 VSS.n3272 1.0492
R3153 VSS.n1276 VSS.n1275 1.00704
R3154 VSS.n1138 VSS.n1113 1.00704
R3155 VSS.n977 VSS.n952 1.00704
R3156 VSS.n2591 VSS.n2590 1.00704
R3157 VSS.n3022 VSS.n3018 1.00704
R3158 VSS.n1609 VSS.n1606 0.95333
R3159 VSS.n1477 VSS.n1474 0.95333
R3160 VSS.n1345 VSS.n1342 0.95333
R3161 VSS.n1584 VSS.n1583 0.949983
R3162 VSS.n1604 VSS.n1603 0.949983
R3163 VSS.n1645 VSS.n1644 0.949983
R3164 VSS.n1452 VSS.n1451 0.949983
R3165 VSS.n1513 VSS.n1512 0.949983
R3166 VSS.n1472 VSS.n1471 0.949983
R3167 VSS.n1320 VSS.n1319 0.949983
R3168 VSS.n1340 VSS.n1339 0.949983
R3169 VSS.n1381 VSS.n1380 0.949983
R3170 VSS.n2572 VSS.n2571 0.890378
R3171 VSS.n2552 VSS.n2551 0.890378
R3172 VSS.n1656 VSS.n1655 0.871152
R3173 VSS.n687 VSS.n686 0.871152
R3174 VSS.n683 VSS.n682 0.871152
R3175 VSS.n682 VSS.n679 0.871152
R3176 VSS.n1559 VSS.n1556 0.871152
R3177 VSS.n686 VSS.n685 0.871152
R3178 VSS.n1563 VSS.n1562 0.871152
R3179 VSS.n1564 VSS.n1563 0.871152
R3180 VSS.n1560 VSS.n1559 0.871152
R3181 VSS.n430 VSS.n429 0.871152
R3182 VSS.n426 VSS.n425 0.871152
R3183 VSS.n425 VSS.n422 0.871152
R3184 VSS.n1523 VSS.n1520 0.871152
R3185 VSS.n429 VSS.n428 0.871152
R3186 VSS.n1527 VSS.n1526 0.871152
R3187 VSS.n1528 VSS.n1527 0.871152
R3188 VSS.n1524 VSS.n1523 0.871152
R3189 VSS.n420 VSS.n419 0.871152
R3190 VSS.n416 VSS.n415 0.871152
R3191 VSS.n415 VSS.n412 0.871152
R3192 VSS.n1427 VSS.n1424 0.871152
R3193 VSS.n419 VSS.n418 0.871152
R3194 VSS.n1431 VSS.n1430 0.871152
R3195 VSS.n1432 VSS.n1431 0.871152
R3196 VSS.n1428 VSS.n1427 0.871152
R3197 VSS.n163 VSS.n162 0.871152
R3198 VSS.n159 VSS.n158 0.871152
R3199 VSS.n158 VSS.n155 0.871152
R3200 VSS.n1391 VSS.n1388 0.871152
R3201 VSS.n162 VSS.n161 0.871152
R3202 VSS.n1395 VSS.n1394 0.871152
R3203 VSS.n1396 VSS.n1395 0.871152
R3204 VSS.n1392 VSS.n1391 0.871152
R3205 VSS.n153 VSS.n152 0.871152
R3206 VSS.n149 VSS.n148 0.871152
R3207 VSS.n148 VSS.n145 0.871152
R3208 VSS.n1295 VSS.n1292 0.871152
R3209 VSS.n152 VSS.n151 0.871152
R3210 VSS.n1299 VSS.n1298 0.871152
R3211 VSS.n1300 VSS.n1299 0.871152
R3212 VSS.n1296 VSS.n1295 0.871152
R3213 VSS.n696 VSS.n695 0.871152
R3214 VSS.n1688 VSS.n1687 0.871152
R3215 VSS.n1689 VSS.n1688 0.871152
R3216 VSS.n693 VSS.n692 0.871152
R3217 VSS.n692 VSS.n689 0.871152
R3218 VSS.n1655 VSS.n1654 0.871152
R3219 VSS.n697 VSS.n696 0.871152
R3220 VSS.n2903 VSS.t637 0.8195
R3221 VSS.n2904 VSS.t649 0.8195
R3222 VSS.n2906 VSS.t670 0.8195
R3223 VSS.n2906 VSS.n2905 0.8195
R3224 VSS.n2922 VSS.t643 0.8195
R3225 VSS.n2922 VSS.n2921 0.8195
R3226 VSS.n2924 VSS.t692 0.8195
R3227 VSS.n2924 VSS.n2923 0.8195
R3228 VSS.n2927 VSS.t642 0.8195
R3229 VSS.n2927 VSS.n2926 0.8195
R3230 VSS.n2929 VSS.t691 0.8195
R3231 VSS.n2929 VSS.n2928 0.8195
R3232 VSS.n2579 VSS.t553 0.8195
R3233 VSS.n2579 VSS.n2578 0.8195
R3234 VSS.n2934 VSS.t487 0.8195
R3235 VSS.n2934 VSS.n2933 0.8195
R3236 VSS.n2932 VSS.t443 0.8195
R3237 VSS.n2932 VSS.n2931 0.8195
R3238 VSS.n2570 VSS.t343 0.8195
R3239 VSS.n2570 VSS.n2569 0.8195
R3240 VSS.n2568 VSS.t345 0.8195
R3241 VSS.n2568 VSS.n2567 0.8195
R3242 VSS.n2565 VSS.t63 0.8195
R3243 VSS.n2565 VSS.n2564 0.8195
R3244 VSS.n2918 VSS.t623 0.8195
R3245 VSS.n2918 VSS.n2917 0.8195
R3246 VSS.n2916 VSS.t617 0.8195
R3247 VSS.n2916 VSS.n2915 0.8195
R3248 VSS.n2562 VSS.t671 0.8195
R3249 VSS.n2562 VSS.n2561 0.8195
R3250 VSS.n2912 VSS.t619 0.8195
R3251 VSS.n2912 VSS.n2911 0.8195
R3252 VSS.n2910 VSS.t646 0.8195
R3253 VSS.n2910 VSS.n2909 0.8195
R3254 VSS.n2044 VSS.n2025 0.799363
R3255 VSS.n1135 VSS.n1115 0.799363
R3256 VSS.n1136 VSS.n1135 0.799363
R3257 VSS.n974 VSS.n954 0.799363
R3258 VSS.n975 VSS.n974 0.799363
R3259 VSS.n2589 VSS.n2588 0.799363
R3260 VSS.n1276 VSS.n1272 0.799163
R3261 VSS.n1138 VSS.n1137 0.799163
R3262 VSS.n977 VSS.n976 0.799163
R3263 VSS.n2591 VSS.n2585 0.799163
R3264 VSS.n3022 VSS.n3021 0.799163
R3265 VSS.n2523 VSS.n2519 0.799163
R3266 VSS.n2523 VSS.n2522 0.799163
R3267 VSS.n3794 VSS.n3793 0.798761
R3268 VSS.n3433 VSS.n3432 0.798761
R3269 VSS.n2252 VSS.n2251 0.798761
R3270 VSS.n2247 VSS.n2244 0.798761
R3271 VSS.n2248 VSS.n2247 0.798761
R3272 VSS.n2251 VSS.n2250 0.798761
R3273 VSS.n2256 VSS.n2255 0.798761
R3274 VSS.n2377 VSS.n2374 0.798761
R3275 VSS.n2378 VSS.n2377 0.798761
R3276 VSS.n2255 VSS.n2254 0.798761
R3277 VSS.n4055 VSS.n4054 0.798761
R3278 VSS.n4056 VSS.n4055 0.798761
R3279 VSS.n3432 VSS.n3431 0.798761
R3280 VSS.n3788 VSS.n3785 0.798761
R3281 VSS.n3789 VSS.n3788 0.798761
R3282 VSS.n3795 VSS.n3794 0.798761
R3283 VSS.n2488 VSS.n2446 0.775283
R3284 VSS.n2481 VSS.n2480 0.775283
R3285 VSS.n3648 VSS.n3548 0.775283
R3286 VSS.n3655 VSS.n3546 0.775283
R3287 VSS.n4058 VSS.t413 0.767371
R3288 VSS.n3990 VSS.t404 0.767371
R3289 VSS.n3530 VSS.n3486 0.738109
R3290 VSS.n3523 VSS.n3492 0.738109
R3291 VSS.n3312 VSS.n3281 0.738109
R3292 VSS.n3319 VSS.n3275 0.738109
R3293 VSS.n2582 VSS.n2581 0.68137
R3294 VSS.n2580 VSS.n2577 0.68137
R3295 VSS.n2560 VSS.n2559 0.68137
R3296 VSS.n2558 VSS.n2557 0.68137
R3297 VSS.n871 VSS.t416 0.656668
R3298 VSS.n927 VSS.t401 0.656668
R3299 VSS.n1032 VSS.t419 0.656668
R3300 VSS.n1088 VSS.t425 0.656668
R3301 VSS.n1193 VSS.t430 0.656668
R3302 VSS.n1249 VSS.t407 0.656668
R3303 VSS.n1650 VSS.n1649 0.626587
R3304 VSS.n1649 VSS.n1648 0.626587
R3305 VSS.n1517 VSS.n1516 0.626587
R3306 VSS.n1518 VSS.n1517 0.626587
R3307 VSS.n1386 VSS.n1385 0.626587
R3308 VSS.n1385 VSS.n1384 0.626587
R3309 VSS.n2442 VSS.n2441 0.626587
R3310 VSS.n2441 VSS.n2440 0.626587
R3311 VSS.n2440 VSS.n2439 0.626587
R3312 VSS.n2439 VSS.n2438 0.626587
R3313 VSS.n2438 VSS.n2437 0.626587
R3314 VSS.n1172 VSS.n1170 0.624916
R3315 VSS.n1011 VSS.n1009 0.624916
R3316 VSS.n850 VSS.n848 0.624916
R3317 VSS.n3213 VSS.n3210 0.624916
R3318 VSS.n2469 VSS.n2468 0.624916
R3319 VSS.n3639 VSS.n3638 0.624916
R3320 VSS.n3761 VSS.n3752 0.624916
R3321 VSS.n3762 VSS.n3761 0.624916
R3322 VSS.n3265 VSS.n3264 0.624916
R3323 VSS.n2359 VSS.n2358 0.624916
R3324 VSS.n3977 VSS.n3976 0.624916
R3325 VSS.n2360 VSS.n2359 0.624916
R3326 VSS.n3421 VSS.n3420 0.62468
R3327 VSS.n1168 VSS.n1141 0.62468
R3328 VSS.n1007 VSS.n980 0.62468
R3329 VSS.n846 VSS.n819 0.62468
R3330 VSS.n3421 VSS.n3396 0.62468
R3331 VSS.n3422 VSS.n3421 0.62468
R3332 VSS.n2830 VSS.n2743 0.608978
R3333 VSS.n2825 VSS.n2745 0.608978
R3334 VSS.n3587 VSS.n3549 0.608978
R3335 VSS.n3593 VSS.n3592 0.608978
R3336 VSS.n1828 VSS.n1825 0.6035
R3337 VSS.n2480 VSS.n2479 0.57963
R3338 VSS.n3548 VSS.n3547 0.57963
R3339 VSS.n3546 VSS.n3545 0.57963
R3340 VSS.n3447 VSS.t170 0.56925
R3341 VSS.n3447 VSS.n3446 0.56925
R3342 VSS.n3444 VSS.t258 0.56925
R3343 VSS.n3444 VSS.n3443 0.56925
R3344 VSS.n3441 VSS.t277 0.56925
R3345 VSS.n3441 VSS.n3440 0.56925
R3346 VSS.n3438 VSS.t189 0.56925
R3347 VSS.n3438 VSS.n3437 0.56925
R3348 VSS.n3435 VSS.t173 0.56925
R3349 VSS.n3435 VSS.n3434 0.56925
R3350 VSS.n16 VSS.t287 0.56925
R3351 VSS.n16 VSS.n15 0.56925
R3352 VSS.n14 VSS.t183 0.56925
R3353 VSS.n14 VSS.n13 0.56925
R3354 VSS.n12 VSS.t165 0.56925
R3355 VSS.n12 VSS.n11 0.56925
R3356 VSS.n3462 VSS.t198 0.56925
R3357 VSS.n3462 VSS.n3461 0.56925
R3358 VSS.n3459 VSS.t214 0.56925
R3359 VSS.n3459 VSS.n3458 0.56925
R3360 VSS.n3456 VSS.t215 0.56925
R3361 VSS.n3456 VSS.n3455 0.56925
R3362 VSS.n3453 VSS.t283 0.56925
R3363 VSS.n3453 VSS.n3452 0.56925
R3364 VSS.n3450 VSS.t259 0.56925
R3365 VSS.n3450 VSS.n3449 0.56925
R3366 VSS.n25 VSS.t232 0.56925
R3367 VSS.n25 VSS.n24 0.56925
R3368 VSS.n23 VSS.t278 0.56925
R3369 VSS.n23 VSS.n22 0.56925
R3370 VSS.n21 VSS.t249 0.56925
R3371 VSS.n21 VSS.n20 0.56925
R3372 VSS.n3477 VSS.t210 0.56925
R3373 VSS.n3477 VSS.n3476 0.56925
R3374 VSS.n3474 VSS.t216 0.56925
R3375 VSS.n3474 VSS.n3473 0.56925
R3376 VSS.n3471 VSS.t260 0.56925
R3377 VSS.n3471 VSS.n3470 0.56925
R3378 VSS.n3468 VSS.t284 0.56925
R3379 VSS.n3468 VSS.n3467 0.56925
R3380 VSS.n3465 VSS.t261 0.56925
R3381 VSS.n3465 VSS.n3464 0.56925
R3382 VSS.n34 VSS.t237 0.56925
R3383 VSS.n34 VSS.n33 0.56925
R3384 VSS.n32 VSS.t280 0.56925
R3385 VSS.n32 VSS.n31 0.56925
R3386 VSS.n30 VSS.t250 0.56925
R3387 VSS.n30 VSS.n29 0.56925
R3388 VSS.n3780 VSS.t163 0.56925
R3389 VSS.n3780 VSS.n3779 0.56925
R3390 VSS.n3777 VSS.t279 0.56925
R3391 VSS.n3777 VSS.n3776 0.56925
R3392 VSS.n3774 VSS.t241 0.56925
R3393 VSS.n3774 VSS.n3773 0.56925
R3394 VSS.n3771 VSS.t202 0.56925
R3395 VSS.n3771 VSS.n3770 0.56925
R3396 VSS.n3768 VSS.t184 0.56925
R3397 VSS.n3768 VSS.n3767 0.56925
R3398 VSS.n43 VSS.t166 0.56925
R3399 VSS.n43 VSS.n42 0.56925
R3400 VSS.n41 VSS.t199 0.56925
R3401 VSS.n41 VSS.n40 0.56925
R3402 VSS.n39 VSS.t174 0.56925
R3403 VSS.n39 VSS.n38 0.56925
R3404 VSS.n2443 VSS.n2442 0.563978
R3405 VSS.n3218 VSS.n3213 0.556813
R3406 VSS.n1580 VSS.t381 0.5465
R3407 VSS.n1580 VSS.n1579 0.5465
R3408 VSS.n1572 VSS.t97 0.5465
R3409 VSS.n1572 VSS.n1571 0.5465
R3410 VSS.n1575 VSS.t363 0.5465
R3411 VSS.n1575 VSS.n1574 0.5465
R3412 VSS.n1568 VSS.t39 0.5465
R3413 VSS.n1568 VSS.n1567 0.5465
R3414 VSS.n1566 VSS.t323 0.5465
R3415 VSS.n1566 VSS.n1565 0.5465
R3416 VSS.n1583 VSS.t70 0.5465
R3417 VSS.n1583 VSS.n1582 0.5465
R3418 VSS.n1600 VSS.t92 0.5465
R3419 VSS.n1600 VSS.n1599 0.5465
R3420 VSS.n1592 VSS.t604 0.5465
R3421 VSS.n1592 VSS.n1591 0.5465
R3422 VSS.n1595 VSS.t395 0.5465
R3423 VSS.n1595 VSS.n1594 0.5465
R3424 VSS.n1588 VSS.t627 0.5465
R3425 VSS.n1588 VSS.n1587 0.5465
R3426 VSS.n1586 VSS.t135 0.5465
R3427 VSS.n1586 VSS.n1585 0.5465
R3428 VSS.n1603 VSS.t333 0.5465
R3429 VSS.n1603 VSS.n1602 0.5465
R3430 VSS.n1636 VSS.t124 0.5465
R3431 VSS.n1636 VSS.n1635 0.5465
R3432 VSS.n1639 VSS.t677 0.5465
R3433 VSS.n1639 VSS.n1638 0.5465
R3434 VSS.n1621 VSS.t113 0.5465
R3435 VSS.n1621 VSS.n1620 0.5465
R3436 VSS.n1624 VSS.t665 0.5465
R3437 VSS.n1624 VSS.n1623 0.5465
R3438 VSS.n1628 VSS.t356 0.5465
R3439 VSS.n1628 VSS.n1627 0.5465
R3440 VSS.n1626 VSS.t134 0.5465
R3441 VSS.n1626 VSS.n1625 0.5465
R3442 VSS.n1612 VSS.t328 0.5465
R3443 VSS.n1612 VSS.n1611 0.5465
R3444 VSS.n1615 VSS.t72 0.5465
R3445 VSS.n1615 VSS.n1614 0.5465
R3446 VSS.n1606 VSS.t629 0.5465
R3447 VSS.n1606 VSS.n1605 0.5465
R3448 VSS.n1608 VSS.t397 0.5465
R3449 VSS.n1608 VSS.n1607 0.5465
R3450 VSS.n1644 VSS.t156 0.5465
R3451 VSS.n1644 VSS.n1643 0.5465
R3452 VSS.n1647 VSS.t601 0.5465
R3453 VSS.n1647 VSS.n1646 0.5465
R3454 VSS.n1448 VSS.t674 0.5465
R3455 VSS.n1448 VSS.n1447 0.5465
R3456 VSS.n1440 VSS.t635 0.5465
R3457 VSS.n1440 VSS.n1439 0.5465
R3458 VSS.n1443 VSS.t136 0.5465
R3459 VSS.n1443 VSS.n1442 0.5465
R3460 VSS.n1436 VSS.t69 0.5465
R3461 VSS.n1436 VSS.n1435 0.5465
R3462 VSS.n1434 VSS.t383 0.5465
R3463 VSS.n1434 VSS.n1433 0.5465
R3464 VSS.n1451 VSS.t396 0.5465
R3465 VSS.n1451 VSS.n1450 0.5465
R3466 VSS.n1515 VSS.t364 0.5465
R3467 VSS.n1515 VSS.n1514 0.5465
R3468 VSS.n1504 VSS.t110 0.5465
R3469 VSS.n1504 VSS.n1503 0.5465
R3470 VSS.n1507 VSS.t304 0.5465
R3471 VSS.n1507 VSS.n1506 0.5465
R3472 VSS.n1489 VSS.t359 0.5465
R3473 VSS.n1489 VSS.n1488 0.5465
R3474 VSS.n1492 VSS.t368 0.5465
R3475 VSS.n1492 VSS.n1491 0.5465
R3476 VSS.n1496 VSS.t310 0.5465
R3477 VSS.n1496 VSS.n1495 0.5465
R3478 VSS.n1494 VSS.t111 0.5465
R3479 VSS.n1494 VSS.n1493 0.5465
R3480 VSS.n1480 VSS.t117 0.5465
R3481 VSS.n1480 VSS.n1479 0.5465
R3482 VSS.n1483 VSS.t380 0.5465
R3483 VSS.n1483 VSS.n1482 0.5465
R3484 VSS.n1474 VSS.t146 0.5465
R3485 VSS.n1474 VSS.n1473 0.5465
R3486 VSS.n1476 VSS.t102 0.5465
R3487 VSS.n1476 VSS.n1475 0.5465
R3488 VSS.n1512 VSS.t90 0.5465
R3489 VSS.n1512 VSS.n1511 0.5465
R3490 VSS.n1468 VSS.t378 0.5465
R3491 VSS.n1468 VSS.n1467 0.5465
R3492 VSS.n1460 VSS.t664 0.5465
R3493 VSS.n1460 VSS.n1459 0.5465
R3494 VSS.n1463 VSS.t675 0.5465
R3495 VSS.n1463 VSS.n1462 0.5465
R3496 VSS.n1456 VSS.t325 0.5465
R3497 VSS.n1456 VSS.n1455 0.5465
R3498 VSS.n1454 VSS.t314 0.5465
R3499 VSS.n1454 VSS.n1453 0.5465
R3500 VSS.n1471 VSS.t324 0.5465
R3501 VSS.n1471 VSS.n1470 0.5465
R3502 VSS.n1316 VSS.t43 0.5465
R3503 VSS.n1316 VSS.n1315 0.5465
R3504 VSS.n1308 VSS.t634 0.5465
R3505 VSS.n1308 VSS.n1307 0.5465
R3506 VSS.n1311 VSS.t23 0.5465
R3507 VSS.n1311 VSS.n1310 0.5465
R3508 VSS.n1304 VSS.t373 0.5465
R3509 VSS.n1304 VSS.n1303 0.5465
R3510 VSS.n1302 VSS.t27 0.5465
R3511 VSS.n1302 VSS.n1301 0.5465
R3512 VSS.n1319 VSS.t109 0.5465
R3513 VSS.n1319 VSS.n1318 0.5465
R3514 VSS.n1336 VSS.t96 0.5465
R3515 VSS.n1336 VSS.n1335 0.5465
R3516 VSS.n1328 VSS.t143 0.5465
R3517 VSS.n1328 VSS.n1327 0.5465
R3518 VSS.n1331 VSS.t80 0.5465
R3519 VSS.n1331 VSS.n1330 0.5465
R3520 VSS.n1324 VSS.t628 0.5465
R3521 VSS.n1324 VSS.n1323 0.5465
R3522 VSS.n1322 VSS.t137 0.5465
R3523 VSS.n1322 VSS.n1321 0.5465
R3524 VSS.n1339 VSS.t129 0.5465
R3525 VSS.n1339 VSS.n1338 0.5465
R3526 VSS.n1372 VSS.t329 0.5465
R3527 VSS.n1372 VSS.n1371 0.5465
R3528 VSS.n1375 VSS.t360 0.5465
R3529 VSS.n1375 VSS.n1374 0.5465
R3530 VSS.n1357 VSS.t305 0.5465
R3531 VSS.n1357 VSS.n1356 0.5465
R3532 VSS.n1360 VSS.t153 0.5465
R3533 VSS.n1360 VSS.n1359 0.5465
R3534 VSS.n1364 VSS.t334 0.5465
R3535 VSS.n1364 VSS.n1363 0.5465
R3536 VSS.n1362 VSS.t382 0.5465
R3537 VSS.n1362 VSS.n1361 0.5465
R3538 VSS.n1348 VSS.t84 0.5465
R3539 VSS.n1348 VSS.n1347 0.5465
R3540 VSS.n1351 VSS.t104 0.5465
R3541 VSS.n1351 VSS.n1350 0.5465
R3542 VSS.n1342 VSS.t676 0.5465
R3543 VSS.n1342 VSS.n1341 0.5465
R3544 VSS.n1344 VSS.t379 0.5465
R3545 VSS.n1344 VSS.n1343 0.5465
R3546 VSS.n1380 VSS.t367 0.5465
R3547 VSS.n1380 VSS.n1379 0.5465
R3548 VSS.n1383 VSS.t652 0.5465
R3549 VSS.n1383 VSS.n1382 0.5465
R3550 VSS.n1700 VSS.n1650 0.5405
R3551 VSS.n1798 VSS.n1518 0.5405
R3552 VSS.n1852 VSS.n1386 0.5405
R3553 VSS.n3488 VSS.n3487 0.479848
R3554 VSS.n3483 VSS.n3482 0.479848
R3555 VSS.n3482 VSS.n3479 0.479848
R3556 VSS.n3489 VSS.n3488 0.479848
R3557 VSS.n3271 VSS.n3268 0.479848
R3558 VSS.n3278 VSS.n3277 0.479848
R3559 VSS.n3277 VSS.n3276 0.479848
R3560 VSS.n3272 VSS.n3271 0.479848
R3561 VSS.n2468 VSS.n2467 0.472687
R3562 VSS.n3977 VSS.n3970 0.472687
R3563 VSS.n3977 VSS.n3967 0.472687
R3564 VSS.n3977 VSS.n3964 0.472687
R3565 VSS.n3977 VSS.n3961 0.472687
R3566 VSS.n3977 VSS.n3958 0.472687
R3567 VSS.n3977 VSS.n3955 0.472687
R3568 VSS.n3977 VSS.n3952 0.472687
R3569 VSS.n3977 VSS.n3949 0.472687
R3570 VSS.n3977 VSS.n3946 0.472687
R3571 VSS.n3977 VSS.n3943 0.472687
R3572 VSS.n3977 VSS.n3942 0.472687
R3573 VSS.n3977 VSS.n3941 0.472687
R3574 VSS.n3977 VSS.n3940 0.472687
R3575 VSS.n3977 VSS.n3939 0.472687
R3576 VSS.n3977 VSS.n3938 0.472687
R3577 VSS.n3977 VSS.n3937 0.472687
R3578 VSS.n3977 VSS.n3936 0.472687
R3579 VSS.n3977 VSS.n3935 0.472687
R3580 VSS.n3977 VSS.n3934 0.472687
R3581 VSS.n3977 VSS.n3933 0.472687
R3582 VSS.n3977 VSS.n3932 0.472687
R3583 VSS.n3977 VSS.n3931 0.472687
R3584 VSS.n3977 VSS.n3930 0.472687
R3585 VSS.n3977 VSS.n3929 0.472687
R3586 VSS.n3977 VSS.n3928 0.472687
R3587 VSS.n3977 VSS.n3927 0.472687
R3588 VSS.n3977 VSS.n3926 0.472687
R3589 VSS.n3977 VSS.n3925 0.472687
R3590 VSS.n3977 VSS.n3924 0.472687
R3591 VSS.n3978 VSS.n3977 0.472687
R3592 VSS.n2359 VSS.n2357 0.472687
R3593 VSS.n2359 VSS.n2356 0.472687
R3594 VSS.n2359 VSS.n2355 0.472687
R3595 VSS.n2359 VSS.n2354 0.472687
R3596 VSS.n2359 VSS.n2353 0.472687
R3597 VSS.n2359 VSS.n2352 0.472687
R3598 VSS.n2359 VSS.n2351 0.472687
R3599 VSS.n2359 VSS.n2350 0.472687
R3600 VSS.n2359 VSS.n2349 0.472687
R3601 VSS.n2359 VSS.n2348 0.472687
R3602 VSS.n2359 VSS.n2347 0.472687
R3603 VSS.n2359 VSS.n2346 0.472687
R3604 VSS.n2359 VSS.n2345 0.472687
R3605 VSS.n2359 VSS.n2344 0.472687
R3606 VSS.n3977 VSS.n3973 0.472687
R3607 VSS.n2055 VSS.n2053 0.472687
R3608 VSS.n132 VSS.n130 0.472687
R3609 VSS.n1169 VSS.n1168 0.472687
R3610 VSS.n1008 VSS.n1007 0.472687
R3611 VSS.n847 VSS.n846 0.472687
R3612 VSS.n2048 VSS.n2046 0.472687
R3613 VSS.n2045 VSS.n2044 0.472687
R3614 VSS.n2044 VSS.n2043 0.472687
R3615 VSS.n2044 VSS.n2042 0.472687
R3616 VSS.n2044 VSS.n2041 0.472687
R3617 VSS.n2044 VSS.n2040 0.472687
R3618 VSS.n2044 VSS.n2039 0.472687
R3619 VSS.n2044 VSS.n2038 0.472687
R3620 VSS.n2044 VSS.n2037 0.472687
R3621 VSS.n2044 VSS.n2036 0.472687
R3622 VSS.n2044 VSS.n2035 0.472687
R3623 VSS.n2044 VSS.n2034 0.472687
R3624 VSS.n2044 VSS.n2033 0.472687
R3625 VSS.n2044 VSS.n2032 0.472687
R3626 VSS.n2044 VSS.n2031 0.472687
R3627 VSS.n2044 VSS.n2030 0.472687
R3628 VSS.n2044 VSS.n2029 0.472687
R3629 VSS.n2044 VSS.n2028 0.472687
R3630 VSS.n2044 VSS.n2027 0.472687
R3631 VSS.n2044 VSS.n2026 0.472687
R3632 VSS.n1135 VSS.n1134 0.472687
R3633 VSS.n1135 VSS.n1133 0.472687
R3634 VSS.n1135 VSS.n1132 0.472687
R3635 VSS.n1135 VSS.n1131 0.472687
R3636 VSS.n1135 VSS.n1130 0.472687
R3637 VSS.n1135 VSS.n1129 0.472687
R3638 VSS.n1135 VSS.n1128 0.472687
R3639 VSS.n1135 VSS.n1127 0.472687
R3640 VSS.n1135 VSS.n1126 0.472687
R3641 VSS.n1135 VSS.n1125 0.472687
R3642 VSS.n1135 VSS.n1124 0.472687
R3643 VSS.n1135 VSS.n1123 0.472687
R3644 VSS.n1135 VSS.n1122 0.472687
R3645 VSS.n1135 VSS.n1121 0.472687
R3646 VSS.n1135 VSS.n1120 0.472687
R3647 VSS.n1135 VSS.n1119 0.472687
R3648 VSS.n1135 VSS.n1118 0.472687
R3649 VSS.n1135 VSS.n1117 0.472687
R3650 VSS.n1135 VSS.n1116 0.472687
R3651 VSS.n974 VSS.n973 0.472687
R3652 VSS.n974 VSS.n972 0.472687
R3653 VSS.n974 VSS.n971 0.472687
R3654 VSS.n974 VSS.n970 0.472687
R3655 VSS.n974 VSS.n969 0.472687
R3656 VSS.n974 VSS.n968 0.472687
R3657 VSS.n974 VSS.n967 0.472687
R3658 VSS.n974 VSS.n966 0.472687
R3659 VSS.n974 VSS.n965 0.472687
R3660 VSS.n974 VSS.n964 0.472687
R3661 VSS.n974 VSS.n963 0.472687
R3662 VSS.n974 VSS.n962 0.472687
R3663 VSS.n974 VSS.n961 0.472687
R3664 VSS.n974 VSS.n960 0.472687
R3665 VSS.n974 VSS.n959 0.472687
R3666 VSS.n974 VSS.n958 0.472687
R3667 VSS.n974 VSS.n957 0.472687
R3668 VSS.n974 VSS.n956 0.472687
R3669 VSS.n974 VSS.n955 0.472687
R3670 VSS.n2838 VSS.n2732 0.472687
R3671 VSS.n2836 VSS.n2742 0.472687
R3672 VSS.n3017 VSS.n3016 0.472687
R3673 VSS.n2550 VSS.n2547 0.472687
R3674 VSS.n2472 VSS.n2471 0.472687
R3675 VSS.n2869 VSS.n2865 0.472687
R3676 VSS.n2869 VSS.n2868 0.472687
R3677 VSS.n3761 VSS.n3760 0.472687
R3678 VSS.n3761 VSS.n3759 0.472687
R3679 VSS.n3761 VSS.n3758 0.472687
R3680 VSS.n3761 VSS.n3757 0.472687
R3681 VSS.n3761 VSS.n3756 0.472687
R3682 VSS.n3761 VSS.n3755 0.472687
R3683 VSS.n3761 VSS.n3754 0.472687
R3684 VSS.n3761 VSS.n3753 0.472687
R3685 VSS.n118 VSS.n4 0.472445
R3686 VSS.n3421 VSS.n3412 0.472445
R3687 VSS.n3421 VSS.n3415 0.472445
R3688 VSS.n3421 VSS.n3418 0.472445
R3689 VSS.n3421 VSS.n3407 0.472445
R3690 VSS.n3421 VSS.n3408 0.472445
R3691 VSS.n3421 VSS.n3409 0.472445
R3692 VSS.n3421 VSS.n3397 0.472445
R3693 VSS.n3421 VSS.n3398 0.472445
R3694 VSS.n3421 VSS.n3399 0.472445
R3695 VSS.n3421 VSS.n3400 0.472445
R3696 VSS.n3421 VSS.n3401 0.472445
R3697 VSS.n3421 VSS.n3402 0.472445
R3698 VSS.n3421 VSS.n3404 0.472445
R3699 VSS.n3421 VSS.n3406 0.472445
R3700 VSS.n3421 VSS.n3405 0.472445
R3701 VSS.n3421 VSS.n3410 0.472445
R3702 VSS.n1168 VSS.n1143 0.472445
R3703 VSS.n1168 VSS.n1144 0.472445
R3704 VSS.n1168 VSS.n1145 0.472445
R3705 VSS.n1168 VSS.n1146 0.472445
R3706 VSS.n1168 VSS.n1147 0.472445
R3707 VSS.n1168 VSS.n1148 0.472445
R3708 VSS.n1168 VSS.n1149 0.472445
R3709 VSS.n1168 VSS.n1150 0.472445
R3710 VSS.n1168 VSS.n1151 0.472445
R3711 VSS.n1168 VSS.n1152 0.472445
R3712 VSS.n1168 VSS.n1153 0.472445
R3713 VSS.n1168 VSS.n1154 0.472445
R3714 VSS.n1168 VSS.n1155 0.472445
R3715 VSS.n1168 VSS.n1156 0.472445
R3716 VSS.n1168 VSS.n1157 0.472445
R3717 VSS.n1168 VSS.n1158 0.472445
R3718 VSS.n1168 VSS.n1159 0.472445
R3719 VSS.n1168 VSS.n1160 0.472445
R3720 VSS.n1168 VSS.n1161 0.472445
R3721 VSS.n1168 VSS.n1162 0.472445
R3722 VSS.n1168 VSS.n1163 0.472445
R3723 VSS.n1168 VSS.n1164 0.472445
R3724 VSS.n1168 VSS.n1165 0.472445
R3725 VSS.n1168 VSS.n1166 0.472445
R3726 VSS.n1168 VSS.n1167 0.472445
R3727 VSS.n1168 VSS.n1142 0.472445
R3728 VSS.n1007 VSS.n982 0.472445
R3729 VSS.n1007 VSS.n983 0.472445
R3730 VSS.n1007 VSS.n984 0.472445
R3731 VSS.n1007 VSS.n985 0.472445
R3732 VSS.n1007 VSS.n986 0.472445
R3733 VSS.n1007 VSS.n987 0.472445
R3734 VSS.n1007 VSS.n988 0.472445
R3735 VSS.n1007 VSS.n989 0.472445
R3736 VSS.n1007 VSS.n990 0.472445
R3737 VSS.n1007 VSS.n991 0.472445
R3738 VSS.n1007 VSS.n992 0.472445
R3739 VSS.n1007 VSS.n993 0.472445
R3740 VSS.n1007 VSS.n994 0.472445
R3741 VSS.n1007 VSS.n995 0.472445
R3742 VSS.n1007 VSS.n996 0.472445
R3743 VSS.n1007 VSS.n997 0.472445
R3744 VSS.n1007 VSS.n998 0.472445
R3745 VSS.n1007 VSS.n999 0.472445
R3746 VSS.n1007 VSS.n1000 0.472445
R3747 VSS.n1007 VSS.n1001 0.472445
R3748 VSS.n1007 VSS.n1002 0.472445
R3749 VSS.n1007 VSS.n1003 0.472445
R3750 VSS.n1007 VSS.n1004 0.472445
R3751 VSS.n1007 VSS.n1005 0.472445
R3752 VSS.n1007 VSS.n1006 0.472445
R3753 VSS.n1007 VSS.n981 0.472445
R3754 VSS.n846 VSS.n845 0.472445
R3755 VSS.n846 VSS.n844 0.472445
R3756 VSS.n846 VSS.n843 0.472445
R3757 VSS.n846 VSS.n842 0.472445
R3758 VSS.n846 VSS.n841 0.472445
R3759 VSS.n846 VSS.n840 0.472445
R3760 VSS.n846 VSS.n839 0.472445
R3761 VSS.n846 VSS.n838 0.472445
R3762 VSS.n846 VSS.n837 0.472445
R3763 VSS.n846 VSS.n836 0.472445
R3764 VSS.n846 VSS.n835 0.472445
R3765 VSS.n846 VSS.n834 0.472445
R3766 VSS.n846 VSS.n833 0.472445
R3767 VSS.n846 VSS.n832 0.472445
R3768 VSS.n846 VSS.n831 0.472445
R3769 VSS.n846 VSS.n830 0.472445
R3770 VSS.n846 VSS.n829 0.472445
R3771 VSS.n846 VSS.n828 0.472445
R3772 VSS.n846 VSS.n827 0.472445
R3773 VSS.n846 VSS.n826 0.472445
R3774 VSS.n846 VSS.n825 0.472445
R3775 VSS.n846 VSS.n824 0.472445
R3776 VSS.n846 VSS.n823 0.472445
R3777 VSS.n846 VSS.n822 0.472445
R3778 VSS.n846 VSS.n821 0.472445
R3779 VSS.n846 VSS.n820 0.472445
R3780 VSS.n3218 VSS.n3216 0.472445
R3781 VSS.n2546 VSS.n2545 0.472445
R3782 VSS.n3421 VSS.n3382 0.472445
R3783 VSS.n3421 VSS.n3383 0.472445
R3784 VSS.n3421 VSS.n3384 0.472445
R3785 VSS.n3421 VSS.n3385 0.472445
R3786 VSS.n3421 VSS.n3386 0.472445
R3787 VSS.n3421 VSS.n3387 0.472445
R3788 VSS.n3421 VSS.n3388 0.472445
R3789 VSS.n3421 VSS.n3389 0.472445
R3790 VSS.n3421 VSS.n3390 0.472445
R3791 VSS.n3421 VSS.n3391 0.472445
R3792 VSS.n3421 VSS.n3392 0.472445
R3793 VSS.n3421 VSS.n3393 0.472445
R3794 VSS.n3421 VSS.n3394 0.472445
R3795 VSS.n3421 VSS.n3395 0.472445
R3796 VSS.n3421 VSS.n3403 0.459997
R3797 VSS.n3977 VSS.n3944 0.457229
R3798 VSS.n3329 VSS.t529 0.449333
R3799 VSS.n3493 VSS.t229 0.449333
R3800 VSS.t226 VSS.t477 0.449333
R3801 VSS.n1139 VSS.n1138 0.320562
R3802 VSS.n1172 VSS.n1139 0.283437
R3803 VSS.n2446 VSS.n2445 0.282239
R3804 VSS.n1752 VSS.n1749 0.270781
R3805 VSS.n2838 VSS.n2836 0.266
R3806 VSS.n1 VSS.n0 0.229438
R3807 VSS.n2050 VSS.n2049 0.229438
R3808 VSS.n128 VSS.n127 0.229438
R3809 VSS.n2445 VSS.n2420 0.207891
R3810 VSS.n2 VSS.n1 0.198781
R3811 VSS.n2051 VSS.n2050 0.198781
R3812 VSS.n129 VSS.n128 0.198781
R3813 VSS.n1650 VSS.n1584 0.190381
R3814 VSS.n1649 VSS.n1604 0.190381
R3815 VSS.n1648 VSS.n1645 0.190381
R3816 VSS.n1518 VSS.n1452 0.190381
R3817 VSS.n1516 VSS.n1513 0.190381
R3818 VSS.n1517 VSS.n1472 0.190381
R3819 VSS.n1386 VSS.n1320 0.190381
R3820 VSS.n1385 VSS.n1340 0.190381
R3821 VSS.n1384 VSS.n1381 0.190381
R3822 VSS.n119 VSS.n2 0.188375
R3823 VSS.n2056 VSS.n2051 0.188375
R3824 VSS.n133 VSS.n129 0.188375
R3825 VSS.n2247 VSS.n2246 0.157022
R3826 VSS.n682 VSS.n681 0.157022
R3827 VSS.n1559 VSS.n1558 0.157022
R3828 VSS.n425 VSS.n424 0.157022
R3829 VSS.n1523 VSS.n1522 0.157022
R3830 VSS.n415 VSS.n414 0.157022
R3831 VSS.n1427 VSS.n1426 0.157022
R3832 VSS.n158 VSS.n157 0.157022
R3833 VSS.n1391 VSS.n1390 0.157022
R3834 VSS.n148 VSS.n147 0.157022
R3835 VSS.n1295 VSS.n1294 0.157022
R3836 VSS.n1655 VSS.n1652 0.157022
R3837 VSS.n692 VSS.n691 0.157022
R3838 VSS.n2420 VSS.n2419 0.157022
R3839 VSS.n3545 VSS.n3544 0.157022
R3840 VSS.n3482 VSS.n3481 0.157022
R3841 VSS.n3271 VSS.n3270 0.157022
R3842 VSS.n2377 VSS.n2376 0.157022
R3843 VSS.n3432 VSS.n3427 0.157022
R3844 VSS.n3788 VSS.n3787 0.157022
R3845 VSS.n1139 VSS.n284 0.148156
R3846 VSS.n978 VSS.n551 0.148156
R3847 VSS.n1011 VSS.n978 0.138594
R3848 VSS.n978 VSS.n977 0.132688
R3849 VSS.n1578 VSS.n1570 0.123658
R3850 VSS.n1598 VSS.n1590 0.123658
R3851 VSS.n1618 VSS.n1610 0.123658
R3852 VSS.n1633 VSS.n1619 0.123658
R3853 VSS.n1642 VSS.n1634 0.123658
R3854 VSS.n1446 VSS.n1438 0.123658
R3855 VSS.n1486 VSS.n1478 0.123658
R3856 VSS.n1501 VSS.n1487 0.123658
R3857 VSS.n1510 VSS.n1502 0.123658
R3858 VSS.n1466 VSS.n1458 0.123658
R3859 VSS.n1314 VSS.n1306 0.123658
R3860 VSS.n1334 VSS.n1326 0.123658
R3861 VSS.n1354 VSS.n1346 0.123658
R3862 VSS.n1369 VSS.n1355 0.123658
R3863 VSS.n1378 VSS.n1370 0.123658
R3864 VSS.n1577 VSS.n1573 0.109963
R3865 VSS.n1597 VSS.n1593 0.109963
R3866 VSS.n1641 VSS.n1637 0.109963
R3867 VSS.n1632 VSS.n1622 0.109963
R3868 VSS.n1617 VSS.n1613 0.109963
R3869 VSS.n1445 VSS.n1441 0.109963
R3870 VSS.n1509 VSS.n1505 0.109963
R3871 VSS.n1500 VSS.n1490 0.109963
R3872 VSS.n1485 VSS.n1481 0.109963
R3873 VSS.n1465 VSS.n1461 0.109963
R3874 VSS.n1313 VSS.n1309 0.109963
R3875 VSS.n1333 VSS.n1329 0.109963
R3876 VSS.n1377 VSS.n1373 0.109963
R3877 VSS.n1368 VSS.n1358 0.109963
R3878 VSS.n1353 VSS.n1349 0.109963
R3879 VSS.n3811 VSS.n3809 0.0800536
R3880 VSS.n3813 VSS.n3811 0.07925
R3881 VSS.n2262 VSS.n2260 0.0760357
R3882 VSS.n2264 VSS.n2262 0.0760357
R3883 VSS.n2266 VSS.n2264 0.0760357
R3884 VSS.n2268 VSS.n2266 0.0760357
R3885 VSS.n2270 VSS.n2268 0.0760357
R3886 VSS.n2272 VSS.n2270 0.0760357
R3887 VSS.n2274 VSS.n2272 0.0760357
R3888 VSS.n2276 VSS.n2274 0.0760357
R3889 VSS.n2278 VSS.n2276 0.0760357
R3890 VSS.n2280 VSS.n2278 0.0760357
R3891 VSS.n2282 VSS.n2280 0.0760357
R3892 VSS.n2284 VSS.n2282 0.0760357
R3893 VSS.n2286 VSS.n2284 0.0760357
R3894 VSS.n2288 VSS.n2286 0.0760357
R3895 VSS.n2290 VSS.n2288 0.0760357
R3896 VSS.n2292 VSS.n2290 0.0760357
R3897 VSS.n2294 VSS.n2292 0.0760357
R3898 VSS.n2296 VSS.n2294 0.0760357
R3899 VSS.n2298 VSS.n2296 0.0760357
R3900 VSS.n2300 VSS.n2298 0.0760357
R3901 VSS.n2302 VSS.n2300 0.0760357
R3902 VSS.n2304 VSS.n2302 0.0760357
R3903 VSS.n2306 VSS.n2304 0.0760357
R3904 VSS.n2308 VSS.n2306 0.0760357
R3905 VSS.n2310 VSS.n2308 0.0760357
R3906 VSS.n2312 VSS.n2310 0.0760357
R3907 VSS.n2314 VSS.n2312 0.0760357
R3908 VSS.n2316 VSS.n2314 0.0760357
R3909 VSS.n2318 VSS.n2316 0.0760357
R3910 VSS.n2321 VSS.n2318 0.0760357
R3911 VSS.n2323 VSS.n2321 0.0760357
R3912 VSS.n2326 VSS.n2323 0.0760357
R3913 VSS.n2328 VSS.n2326 0.0760357
R3914 VSS.n2331 VSS.n2328 0.0760357
R3915 VSS.n2333 VSS.n2331 0.0760357
R3916 VSS.n2336 VSS.n2333 0.0760357
R3917 VSS.n2338 VSS.n2336 0.0760357
R3918 VSS.n2341 VSS.n2338 0.0760357
R3919 VSS.n2343 VSS.n2341 0.0760357
R3920 VSS.n59 VSS.n58 0.0760357
R3921 VSS.n58 VSS.n57 0.0760357
R3922 VSS.n57 VSS.n56 0.0760357
R3923 VSS.n56 VSS.n55 0.0760357
R3924 VSS.n55 VSS.n54 0.0760357
R3925 VSS.n54 VSS.n53 0.0760357
R3926 VSS.n53 VSS.n52 0.0760357
R3927 VSS.n52 VSS.n51 0.0760357
R3928 VSS.n51 VSS.n50 0.0760357
R3929 VSS.n3797 VSS.n3796 0.0760357
R3930 VSS.n3798 VSS.n3797 0.0760357
R3931 VSS.n3799 VSS.n3798 0.0760357
R3932 VSS.n3800 VSS.n3799 0.0760357
R3933 VSS.n3801 VSS.n3800 0.0760357
R3934 VSS.n3802 VSS.n3801 0.0760357
R3935 VSS.n3803 VSS.n3802 0.0760357
R3936 VSS.n3804 VSS.n3803 0.0760357
R3937 VSS.n3805 VSS.n3804 0.0760357
R3938 VSS.n3807 VSS.n3805 0.0760357
R3939 VSS.n3809 VSS.n3807 0.0760357
R3940 VSS.n3815 VSS.n3813 0.0760357
R3941 VSS.n3817 VSS.n3815 0.0760357
R3942 VSS.n3819 VSS.n3817 0.0760357
R3943 VSS.n3821 VSS.n3819 0.0760357
R3944 VSS.n3823 VSS.n3821 0.0760357
R3945 VSS.n3825 VSS.n3823 0.0760357
R3946 VSS.n3827 VSS.n3825 0.0760357
R3947 VSS.n3829 VSS.n3827 0.0760357
R3948 VSS.n3831 VSS.n3829 0.0760357
R3949 VSS.n3833 VSS.n3831 0.0760357
R3950 VSS.n3835 VSS.n3833 0.0760357
R3951 VSS.n3837 VSS.n3835 0.0760357
R3952 VSS.n3839 VSS.n3837 0.0760357
R3953 VSS.n3841 VSS.n3839 0.0760357
R3954 VSS.n3843 VSS.n3841 0.0760357
R3955 VSS.n3845 VSS.n3843 0.0760357
R3956 VSS.n3847 VSS.n3845 0.0760357
R3957 VSS.n3849 VSS.n3847 0.0760357
R3958 VSS.n3851 VSS.n3849 0.0760357
R3959 VSS.n3853 VSS.n3851 0.0760357
R3960 VSS.n3855 VSS.n3853 0.0760357
R3961 VSS.n3857 VSS.n3855 0.0760357
R3962 VSS.n3859 VSS.n3857 0.0760357
R3963 VSS.n3861 VSS.n3859 0.0760357
R3964 VSS.n3863 VSS.n3861 0.0760357
R3965 VSS.n3865 VSS.n3863 0.0760357
R3966 VSS.n3867 VSS.n3865 0.0760357
R3967 VSS.n3869 VSS.n3867 0.0760357
R3968 VSS.n3871 VSS.n3869 0.0760357
R3969 VSS.n3873 VSS.n3871 0.0760357
R3970 VSS.n3875 VSS.n3873 0.0760357
R3971 VSS.n3877 VSS.n3875 0.0760357
R3972 VSS.n3879 VSS.n3877 0.0760357
R3973 VSS.n3881 VSS.n3879 0.0760357
R3974 VSS.n3883 VSS.n3881 0.0760357
R3975 VSS.n3885 VSS.n3883 0.0760357
R3976 VSS.n3887 VSS.n3885 0.0760357
R3977 VSS.n3889 VSS.n3887 0.0760357
R3978 VSS.n3891 VSS.n3889 0.0760357
R3979 VSS.n3893 VSS.n3891 0.0760357
R3980 VSS.n3896 VSS.n3893 0.0760357
R3981 VSS.n3898 VSS.n3896 0.0760357
R3982 VSS.n3901 VSS.n3898 0.0760357
R3983 VSS.n3903 VSS.n3901 0.0760357
R3984 VSS.n3906 VSS.n3903 0.0760357
R3985 VSS.n3908 VSS.n3906 0.0760357
R3986 VSS.n3911 VSS.n3908 0.0760357
R3987 VSS.n3913 VSS.n3911 0.0760357
R3988 VSS.n3916 VSS.n3913 0.0760357
R3989 VSS.n3918 VSS.n3916 0.0760357
R3990 VSS.n3921 VSS.n3918 0.0760357
R3991 VSS.n3923 VSS.n3921 0.0760357
R3992 VSS.n3980 VSS.n3923 0.0760357
R3993 VSS.n2162 VSS.n2160 0.0760357
R3994 VSS.n2164 VSS.n2162 0.0760357
R3995 VSS.n2166 VSS.n2164 0.0760357
R3996 VSS.n2168 VSS.n2166 0.0760357
R3997 VSS.n2170 VSS.n2168 0.0760357
R3998 VSS.n2172 VSS.n2170 0.0760357
R3999 VSS.n2174 VSS.n2172 0.0760357
R4000 VSS.n2176 VSS.n2174 0.0760357
R4001 VSS.n2178 VSS.n2176 0.0760357
R4002 VSS.n2180 VSS.n2178 0.0760357
R4003 VSS.n2182 VSS.n2180 0.0760357
R4004 VSS.n2184 VSS.n2182 0.0760357
R4005 VSS.n2186 VSS.n2184 0.0760357
R4006 VSS.n2188 VSS.n2186 0.0760357
R4007 VSS.n2190 VSS.n2188 0.0760357
R4008 VSS.n2192 VSS.n2190 0.0760357
R4009 VSS.n2194 VSS.n2192 0.0760357
R4010 VSS.n2196 VSS.n2194 0.0760357
R4011 VSS.n2198 VSS.n2196 0.0760357
R4012 VSS.n2200 VSS.n2198 0.0760357
R4013 VSS.n2202 VSS.n2200 0.0760357
R4014 VSS.n2204 VSS.n2202 0.0760357
R4015 VSS.n2206 VSS.n2204 0.0760357
R4016 VSS.n2208 VSS.n2206 0.0760357
R4017 VSS.n2210 VSS.n2208 0.0760357
R4018 VSS.n2212 VSS.n2210 0.0760357
R4019 VSS.n2214 VSS.n2212 0.0760357
R4020 VSS.n2216 VSS.n2214 0.0760357
R4021 VSS.n2218 VSS.n2216 0.0760357
R4022 VSS.n2221 VSS.n2218 0.0760357
R4023 VSS.n2223 VSS.n2221 0.0760357
R4024 VSS.n2226 VSS.n2223 0.0760357
R4025 VSS.n2228 VSS.n2226 0.0760357
R4026 VSS.n2231 VSS.n2228 0.0760357
R4027 VSS.n2233 VSS.n2231 0.0760357
R4028 VSS.n2236 VSS.n2233 0.0760357
R4029 VSS.n2238 VSS.n2236 0.0760357
R4030 VSS.n2241 VSS.n2238 0.0760357
R4031 VSS.n2242 VSS.n2241 0.0760357
R4032 VSS.n2577 VSS.n2576 0.068
R4033 VSS.n2557 VSS.n2556 0.068
R4034 VSS.n2062 VSS.n2060 0.0561875
R4035 VSS.n2064 VSS.n2062 0.055625
R4036 VSS.n3751 VSS.n3749 0.053375
R4037 VSS.n3749 VSS.n3746 0.053375
R4038 VSS.n3746 VSS.n3744 0.053375
R4039 VSS.n3744 VSS.n3741 0.053375
R4040 VSS.n3741 VSS.n3739 0.053375
R4041 VSS.n3739 VSS.n3736 0.053375
R4042 VSS.n3736 VSS.n3734 0.053375
R4043 VSS.n3734 VSS.n3731 0.053375
R4044 VSS.n3731 VSS.n3729 0.053375
R4045 VSS.n3729 VSS.n3726 0.053375
R4046 VSS.n3726 VSS.n3724 0.053375
R4047 VSS.n3724 VSS.n3721 0.053375
R4048 VSS.n3721 VSS.n3719 0.053375
R4049 VSS.n3719 VSS.n3716 0.053375
R4050 VSS.n3716 VSS.n3714 0.053375
R4051 VSS.n3714 VSS.n3711 0.053375
R4052 VSS.n3711 VSS.n3709 0.053375
R4053 VSS.n3709 VSS.n3707 0.053375
R4054 VSS.n3707 VSS.n3705 0.053375
R4055 VSS.n3705 VSS.n3703 0.053375
R4056 VSS.n3703 VSS.n3701 0.053375
R4057 VSS.n3701 VSS.n3699 0.053375
R4058 VSS.n3699 VSS.n3697 0.053375
R4059 VSS.n3697 VSS.n3695 0.053375
R4060 VSS.n3695 VSS.n3693 0.053375
R4061 VSS.n3693 VSS.n3691 0.053375
R4062 VSS.n3691 VSS.n3689 0.053375
R4063 VSS.n3689 VSS.n3687 0.053375
R4064 VSS.n3687 VSS.n3685 0.053375
R4065 VSS.n3685 VSS.n3683 0.053375
R4066 VSS.n3683 VSS.n3681 0.053375
R4067 VSS.n3681 VSS.n3679 0.053375
R4068 VSS.n3679 VSS.n3677 0.053375
R4069 VSS.n2517 VSS.n2515 0.053375
R4070 VSS.n2515 VSS.n2513 0.053375
R4071 VSS.n2513 VSS.n2511 0.053375
R4072 VSS.n2543 VSS.n2540 0.053375
R4073 VSS.n2540 VSS.n2537 0.053375
R4074 VSS.n2537 VSS.n2534 0.053375
R4075 VSS.n2534 VSS.n2532 0.053375
R4076 VSS.n2532 VSS.n2530 0.053375
R4077 VSS.n2530 VSS.n2528 0.053375
R4078 VSS.n2528 VSS.n2526 0.053375
R4079 VSS.n2465 VSS.n2463 0.053375
R4080 VSS.n2463 VSS.n2460 0.053375
R4081 VSS.n2460 VSS.n2458 0.053375
R4082 VSS.n2458 VSS.n2455 0.053375
R4083 VSS.n2455 VSS.n2453 0.053375
R4084 VSS.n2453 VSS.n2450 0.053375
R4085 VSS.n2450 VSS.n2448 0.053375
R4086 VSS.n2736 VSS.n2734 0.053375
R4087 VSS.n2739 VSS.n2736 0.053375
R4088 VSS.n3637 VSS.n3635 0.053375
R4089 VSS.n3635 VSS.n3632 0.053375
R4090 VSS.n3632 VSS.n3630 0.053375
R4091 VSS.n3630 VSS.n3627 0.053375
R4092 VSS.n3627 VSS.n3625 0.053375
R4093 VSS.n3625 VSS.n3622 0.053375
R4094 VSS.n3622 VSS.n3620 0.053375
R4095 VSS.n3620 VSS.n3617 0.053375
R4096 VSS.n3617 VSS.n3615 0.053375
R4097 VSS.n3615 VSS.n3612 0.053375
R4098 VSS.n3612 VSS.n3610 0.053375
R4099 VSS.n3610 VSS.n3607 0.053375
R4100 VSS.n3607 VSS.n3605 0.053375
R4101 VSS.n3605 VSS.n3602 0.053375
R4102 VSS.n121 VSS.n120 0.053375
R4103 VSS.n122 VSS.n121 0.053375
R4104 VSS.n123 VSS.n122 0.053375
R4105 VSS.n124 VSS.n123 0.053375
R4106 VSS.n126 VSS.n124 0.053375
R4107 VSS.n137 VSS.n135 0.053375
R4108 VSS.n139 VSS.n137 0.053375
R4109 VSS.n141 VSS.n139 0.053375
R4110 VSS.n143 VSS.n141 0.053375
R4111 VSS.n2060 VSS.n2058 0.053375
R4112 VSS.n2066 VSS.n2064 0.053375
R4113 VSS.n2068 VSS.n2066 0.053375
R4114 VSS.n2070 VSS.n2068 0.053375
R4115 VSS.n2072 VSS.n2070 0.053375
R4116 VSS.n2074 VSS.n2072 0.053375
R4117 VSS.n2076 VSS.n2074 0.053375
R4118 VSS.n2078 VSS.n2076 0.053375
R4119 VSS.n2080 VSS.n2078 0.053375
R4120 VSS.n2082 VSS.n2080 0.053375
R4121 VSS.n2084 VSS.n2082 0.053375
R4122 VSS.n2086 VSS.n2084 0.053375
R4123 VSS.n2088 VSS.n2086 0.053375
R4124 VSS.n3258 VSS.n3256 0.053375
R4125 VSS.n3256 VSS.n3253 0.053375
R4126 VSS.n3253 VSS.n3251 0.053375
R4127 VSS.n3251 VSS.n3248 0.053375
R4128 VSS.n3248 VSS.n3246 0.053375
R4129 VSS.n3246 VSS.n3243 0.053375
R4130 VSS.n3243 VSS.n3241 0.053375
R4131 VSS.n3241 VSS.n3238 0.053375
R4132 VSS.n3238 VSS.n3236 0.053375
R4133 VSS.n3236 VSS.n3233 0.053375
R4134 VSS.n3233 VSS.n3231 0.053375
R4135 VSS.n3231 VSS.n3228 0.053375
R4136 VSS.n3228 VSS.n3226 0.053375
R4137 VSS.n3226 VSS.n3223 0.053375
R4138 VSS.n3223 VSS.n3221 0.053375
R4139 VSS.n2478 VSS.n2475 0.053375
R4140 VSS.n2487 VSS.n2484 0.053375
R4141 VSS.n2494 VSS.n2491 0.053375
R4142 VSS.n2497 VSS.n2494 0.053375
R4143 VSS.n2500 VSS.n2497 0.053375
R4144 VSS.n2503 VSS.n2500 0.053375
R4145 VSS.n2506 VSS.n2503 0.053375
R4146 VSS.n2508 VSS.n2506 0.053375
R4147 VSS.n2834 VSS.n2832 0.053375
R4148 VSS.n2829 VSS.n2827 0.053375
R4149 VSS.n2824 VSS.n2822 0.053375
R4150 VSS.n2816 VSS.n2814 0.053375
R4151 VSS.n2811 VSS.n2809 0.053375
R4152 VSS.n2803 VSS.n2801 0.053375
R4153 VSS.n2801 VSS.n2799 0.053375
R4154 VSS.n2799 VSS.n2797 0.053375
R4155 VSS.n2797 VSS.n2795 0.053375
R4156 VSS.n2795 VSS.n2793 0.053375
R4157 VSS.n2793 VSS.n2791 0.053375
R4158 VSS.n2791 VSS.n2789 0.053375
R4159 VSS.n2789 VSS.n2787 0.053375
R4160 VSS.n2787 VSS.n2785 0.053375
R4161 VSS.n2785 VSS.n2783 0.053375
R4162 VSS.n2783 VSS.n2781 0.053375
R4163 VSS.n2781 VSS.n2779 0.053375
R4164 VSS.n2779 VSS.n2777 0.053375
R4165 VSS.n2777 VSS.n2775 0.053375
R4166 VSS.n2775 VSS.n2773 0.053375
R4167 VSS.n2770 VSS.n2768 0.053375
R4168 VSS.n2768 VSS.n2766 0.053375
R4169 VSS.n2766 VSS.n2764 0.053375
R4170 VSS.n2764 VSS.n2762 0.053375
R4171 VSS.n2759 VSS.n2757 0.053375
R4172 VSS.n2757 VSS.n2755 0.053375
R4173 VSS.n3562 VSS.n3560 0.053375
R4174 VSS.n3564 VSS.n3562 0.053375
R4175 VSS.n3566 VSS.n3564 0.053375
R4176 VSS.n3568 VSS.n3566 0.053375
R4177 VSS.n3573 VSS.n3571 0.053375
R4178 VSS.n3575 VSS.n3573 0.053375
R4179 VSS.n3577 VSS.n3575 0.053375
R4180 VSS.n3582 VSS.n3580 0.053375
R4181 VSS.n3584 VSS.n3582 0.053375
R4182 VSS.n3586 VSS.n3584 0.053375
R4183 VSS.n3591 VSS.n3589 0.053375
R4184 VSS.n3597 VSS.n3595 0.053375
R4185 VSS.n3600 VSS.n3597 0.053375
R4186 VSS.n3675 VSS.n3673 0.053375
R4187 VSS.n3673 VSS.n3670 0.053375
R4188 VSS.n3670 VSS.n3667 0.053375
R4189 VSS.n3667 VSS.n3664 0.053375
R4190 VSS.n3664 VSS.n3661 0.053375
R4191 VSS.n3661 VSS.n3658 0.053375
R4192 VSS.n3654 VSS.n3651 0.053375
R4193 VSS.n3647 VSS.n3644 0.053375
R4194 VSS.n3644 VSS.n3641 0.053375
R4195 VSS.n3331 VSS.n3328 0.053375
R4196 VSS.n3328 VSS.n3325 0.053375
R4197 VSS.n3325 VSS.n3322 0.053375
R4198 VSS.n3318 VSS.n3315 0.053375
R4199 VSS.n3311 VSS.n3308 0.053375
R4200 VSS.n3308 VSS.n3305 0.053375
R4201 VSS.n3305 VSS.n3302 0.053375
R4202 VSS.n3302 VSS.n3299 0.053375
R4203 VSS.n3299 VSS.n3296 0.053375
R4204 VSS.n3296 VSS.n3293 0.053375
R4205 VSS.n3293 VSS.n3290 0.053375
R4206 VSS.n3290 VSS.n3287 0.053375
R4207 VSS.n3287 VSS.n3284 0.053375
R4208 VSS.n3498 VSS.n3495 0.053375
R4209 VSS.n3501 VSS.n3498 0.053375
R4210 VSS.n3504 VSS.n3501 0.053375
R4211 VSS.n3507 VSS.n3504 0.053375
R4212 VSS.n3510 VSS.n3507 0.053375
R4213 VSS.n3513 VSS.n3510 0.053375
R4214 VSS.n3516 VSS.n3513 0.053375
R4215 VSS.n3519 VSS.n3516 0.053375
R4216 VSS.n3522 VSS.n3519 0.053375
R4217 VSS.n3529 VSS.n3526 0.053375
R4218 VSS.n3536 VSS.n3533 0.053375
R4219 VSS.n3539 VSS.n3536 0.053375
R4220 VSS.n3542 VSS.n3539 0.053375
R4221 VSS.n2365 VSS.n2362 0.053375
R4222 VSS.n2372 VSS.n2369 0.053375
R4223 VSS.n2385 VSS.n2382 0.053375
R4224 VSS.n2388 VSS.n2385 0.053375
R4225 VSS.n2391 VSS.n2388 0.053375
R4226 VSS.n2394 VSS.n2391 0.053375
R4227 VSS.n2397 VSS.n2394 0.053375
R4228 VSS.n2400 VSS.n2397 0.053375
R4229 VSS.n2403 VSS.n2400 0.053375
R4230 VSS.n2099 VSS.n2097 0.053375
R4231 VSS.n2104 VSS.n2102 0.053375
R4232 VSS.n2109 VSS.n2107 0.053375
R4233 VSS.n2111 VSS.n2109 0.053375
R4234 VSS.n2113 VSS.n2111 0.053375
R4235 VSS.n2115 VSS.n2113 0.053375
R4236 VSS.n2117 VSS.n2115 0.053375
R4237 VSS.n2119 VSS.n2117 0.053375
R4238 VSS.n2121 VSS.n2119 0.053375
R4239 VSS.n2123 VSS.n2121 0.053375
R4240 VSS.n2128 VSS.n2126 0.053375
R4241 VSS.n2130 VSS.n2128 0.053375
R4242 VSS.n2132 VSS.n2130 0.053375
R4243 VSS.n2134 VSS.n2132 0.053375
R4244 VSS.n2136 VSS.n2134 0.053375
R4245 VSS.n2138 VSS.n2136 0.053375
R4246 VSS.n2143 VSS.n2141 0.053375
R4247 VSS.n2145 VSS.n2143 0.053375
R4248 VSS.n2147 VSS.n2145 0.053375
R4249 VSS.n2152 VSS.n2150 0.053375
R4250 VSS.n3340 VSS.n3337 0.053375
R4251 VSS.n3343 VSS.n3340 0.053375
R4252 VSS.n3346 VSS.n3343 0.053375
R4253 VSS.n3349 VSS.n3346 0.053375
R4254 VSS.n3352 VSS.n3349 0.053375
R4255 VSS.n3355 VSS.n3352 0.053375
R4256 VSS.n3358 VSS.n3355 0.053375
R4257 VSS.n3361 VSS.n3358 0.053375
R4258 VSS.n3364 VSS.n3361 0.053375
R4259 VSS.n3367 VSS.n3364 0.053375
R4260 VSS.n3370 VSS.n3367 0.053375
R4261 VSS.n3378 VSS.n3374 0.053375
R4262 VSS VSS.n3380 0.053375
R4263 VSS VSS.n4067 0.053375
R4264 VSS.n4067 VSS.n4064 0.053375
R4265 VSS.n4050 VSS.n4047 0.053375
R4266 VSS.n4047 VSS.n4044 0.053375
R4267 VSS.n4040 VSS.n4037 0.053375
R4268 VSS.n4037 VSS.n4034 0.053375
R4269 VSS.n4034 VSS.n4031 0.053375
R4270 VSS.n4027 VSS.n4024 0.053375
R4271 VSS.n4024 VSS.n4021 0.053375
R4272 VSS.n4017 VSS.n4014 0.053375
R4273 VSS.n117 VSS.n115 0.053375
R4274 VSS.n109 VSS.n107 0.053375
R4275 VSS.n107 VSS.n105 0.053375
R4276 VSS.n102 VSS.n100 0.053375
R4277 VSS.n100 VSS.n98 0.053375
R4278 VSS.n98 VSS.n96 0.053375
R4279 VSS.n93 VSS.n91 0.053375
R4280 VSS.n91 VSS.n89 0.053375
R4281 VSS.n86 VSS.n84 0.053375
R4282 VSS.n84 VSS.n82 0.053375
R4283 VSS.n82 VSS.n80 0.053375
R4284 VSS.n77 VSS.n75 0.053375
R4285 VSS.n75 VSS.n73 0.053375
R4286 VSS.n64 VSS.n62 0.053375
R4287 VSS.n62 VSS.n60 0.053375
R4288 VSS.n4002 VSS.n3999 0.053375
R4289 VSS.n3999 VSS.n3996 0.053375
R4290 VSS.n3988 VSS.n3985 0.053375
R4291 VSS.n3985 VSS.n3982 0.053375
R4292 VSS.n4014 VSS.n4011 0.0530441
R4293 VSS.n3578 VSS.n3577 0.0528125
R4294 VSS.n2406 VSS.n2403 0.05275
R4295 VSS.n2058 VSS.n2056 0.0505625
R4296 VSS.n2820 VSS.n2819 0.0505625
R4297 VSS.n3322 VSS.n3319 0.05
R4298 VSS.n3533 VSS.n3530 0.048875
R4299 VSS.n2366 VSS.n2365 0.0483125
R4300 VSS.n2095 VSS.n2094 0.0483125
R4301 VSS.n2155 VSS.n2153 0.0483125
R4302 VSS.n3380 VSS.n3379 0.0483125
R4303 VSS.n4044 VSS.n4041 0.04775
R4304 VSS.n105 VSS.n103 0.04775
R4305 VSS.n78 VSS.n77 0.04775
R4306 VSS.n4061 VSS.n4060 0.046625
R4307 VSS.n113 VSS.n112 0.046625
R4308 VSS.n67 VSS.n65 0.046625
R4309 VSS.n3992 VSS.n3989 0.046625
R4310 VSS.n2806 VSS.n2804 0.0460625
R4311 VSS.n2126 VSS.n2124 0.0460625
R4312 VSS.n2807 VSS.n2806 0.0449375
R4313 VSS.n4060 VSS.n4057 0.044375
R4314 VSS.n112 VSS.n110 0.044375
R4315 VSS.n71 VSS.n67 0.044375
R4316 VSS.n3993 VSS.n3992 0.044375
R4317 VSS.n2760 VSS.n2759 0.0426875
R4318 VSS.n3558 VSS.n3557 0.0426875
R4319 VSS.n2576 VSS.n2575 0.0410839
R4320 VSS.n2556 VSS.n2555 0.0410839
R4321 VSS.n2819 VSS.n2817 0.0404375
R4322 VSS.n2156 VSS.n2155 0.039875
R4323 VSS.n118 VSS.n117 0.037625
R4324 VSS.n4028 VSS.n4027 0.037625
R4325 VSS.n4021 VSS.n4018 0.037625
R4326 VSS.n94 VSS.n93 0.037625
R4327 VSS.n89 VSS.n87 0.037625
R4328 VSS.n4008 VSS.n4007 0.0354412
R4329 VSS.n3332 VSS.n3331 0.0349608
R4330 VSS.n3765 VSS.n3542 0.0349492
R4331 VSS.n2056 VSS.n143 0.0348125
R4332 VSS.n2481 VSS.n2478 0.0348125
R4333 VSS.n2491 VSS.n2488 0.0348125
R4334 VSS.n2832 VSS.n2830 0.0348125
R4335 VSS.n2825 VSS.n2824 0.0348125
R4336 VSS.n3587 VSS.n3586 0.0348125
R4337 VSS.n3595 VSS.n3593 0.0348125
R4338 VSS.n3658 VSS.n3655 0.0348125
R4339 VSS.n3648 VSS.n3647 0.0348125
R4340 VSS.n3315 VSS.n3312 0.03425
R4341 VSS.n2139 VSS.n2138 0.03425
R4342 VSS.n2410 VSS.n2407 0.0335
R4343 VSS.n3526 VSS.n3523 0.033125
R4344 VSS.n2773 VSS.n2771 0.0325625
R4345 VSS.n3571 VSS.n3569 0.0325625
R4346 VSS.n2379 VSS.n2372 0.0325625
R4347 VSS.n2100 VSS.n2099 0.0325625
R4348 VSS.n2150 VSS.n2148 0.0325625
R4349 VSS.n3374 VSS.n3371 0.0325625
R4350 VSS.n2836 VSS.n2834 0.030875
R4351 VSS.n2475 VSS.n2472 0.030875
R4352 VSS.n4003 VSS.n4002 0.0307426
R4353 VSS.n3337 VSS.n3334 0.029625
R4354 VSS.n2812 VSS.n2811 0.0291875
R4355 VSS.n2107 VSS.n2105 0.0280625
R4356 VSS.n851 VSS.n817 0.0269375
R4357 VSS.n817 VSS.n814 0.0269375
R4358 VSS.n814 VSS.n812 0.0269375
R4359 VSS.n812 VSS.n809 0.0269375
R4360 VSS.n809 VSS.n807 0.0269375
R4361 VSS.n807 VSS.n804 0.0269375
R4362 VSS.n804 VSS.n802 0.0269375
R4363 VSS.n802 VSS.n799 0.0269375
R4364 VSS.n799 VSS.n797 0.0269375
R4365 VSS.n797 VSS.n794 0.0269375
R4366 VSS.n794 VSS.n792 0.0269375
R4367 VSS.n792 VSS.n789 0.0269375
R4368 VSS.n789 VSS.n787 0.0269375
R4369 VSS.n787 VSS.n785 0.0269375
R4370 VSS.n785 VSS.n783 0.0269375
R4371 VSS.n783 VSS.n781 0.0269375
R4372 VSS.n781 VSS.n779 0.0269375
R4373 VSS.n779 VSS.n777 0.0269375
R4374 VSS.n777 VSS.n775 0.0269375
R4375 VSS.n775 VSS.n773 0.0269375
R4376 VSS.n773 VSS.n771 0.0269375
R4377 VSS.n771 VSS.n769 0.0269375
R4378 VSS.n769 VSS.n767 0.0269375
R4379 VSS.n767 VSS.n765 0.0269375
R4380 VSS.n765 VSS.n763 0.0269375
R4381 VSS.n763 VSS.n761 0.0269375
R4382 VSS.n761 VSS.n759 0.0269375
R4383 VSS.n759 VSS.n757 0.0269375
R4384 VSS.n757 VSS.n755 0.0269375
R4385 VSS.n755 VSS.n753 0.0269375
R4386 VSS.n753 VSS.n751 0.0269375
R4387 VSS.n751 VSS.n749 0.0269375
R4388 VSS.n749 VSS.n747 0.0269375
R4389 VSS.n747 VSS.n745 0.0269375
R4390 VSS.n745 VSS.n743 0.0269375
R4391 VSS.n743 VSS.n741 0.0269375
R4392 VSS.n741 VSS.n739 0.0269375
R4393 VSS.n739 VSS.n737 0.0269375
R4394 VSS.n737 VSS.n735 0.0269375
R4395 VSS.n735 VSS.n733 0.0269375
R4396 VSS.n733 VSS.n731 0.0269375
R4397 VSS.n731 VSS.n729 0.0269375
R4398 VSS.n729 VSS.n727 0.0269375
R4399 VSS.n727 VSS.n725 0.0269375
R4400 VSS.n725 VSS.n723 0.0269375
R4401 VSS.n723 VSS.n721 0.0269375
R4402 VSS.n721 VSS.n719 0.0269375
R4403 VSS.n719 VSS.n717 0.0269375
R4404 VSS.n717 VSS.n715 0.0269375
R4405 VSS.n715 VSS.n713 0.0269375
R4406 VSS.n713 VSS.n711 0.0269375
R4407 VSS.n711 VSS.n709 0.0269375
R4408 VSS.n709 VSS.n707 0.0269375
R4409 VSS.n707 VSS.n705 0.0269375
R4410 VSS.n705 VSS.n703 0.0269375
R4411 VSS.n703 VSS.n701 0.0269375
R4412 VSS.n701 VSS.n699 0.0269375
R4413 VSS.n1660 VSS.n1658 0.0269375
R4414 VSS.n1662 VSS.n1660 0.0269375
R4415 VSS.n1664 VSS.n1662 0.0269375
R4416 VSS.n1666 VSS.n1664 0.0269375
R4417 VSS.n1668 VSS.n1666 0.0269375
R4418 VSS.n1673 VSS.n1668 0.0269375
R4419 VSS.n949 VSS.n677 0.0269375
R4420 VSS.n677 VSS.n675 0.0269375
R4421 VSS.n675 VSS.n672 0.0269375
R4422 VSS.n672 VSS.n669 0.0269375
R4423 VSS.n669 VSS.n667 0.0269375
R4424 VSS.n667 VSS.n664 0.0269375
R4425 VSS.n664 VSS.n662 0.0269375
R4426 VSS.n662 VSS.n659 0.0269375
R4427 VSS.n659 VSS.n657 0.0269375
R4428 VSS.n657 VSS.n654 0.0269375
R4429 VSS.n654 VSS.n652 0.0269375
R4430 VSS.n652 VSS.n649 0.0269375
R4431 VSS.n649 VSS.n647 0.0269375
R4432 VSS.n647 VSS.n644 0.0269375
R4433 VSS.n644 VSS.n642 0.0269375
R4434 VSS.n642 VSS.n639 0.0269375
R4435 VSS.n639 VSS.n637 0.0269375
R4436 VSS.n637 VSS.n634 0.0269375
R4437 VSS.n634 VSS.n632 0.0269375
R4438 VSS.n632 VSS.n629 0.0269375
R4439 VSS.n629 VSS.n627 0.0269375
R4440 VSS.n627 VSS.n624 0.0269375
R4441 VSS.n624 VSS.n622 0.0269375
R4442 VSS.n622 VSS.n619 0.0269375
R4443 VSS.n619 VSS.n617 0.0269375
R4444 VSS.n617 VSS.n615 0.0269375
R4445 VSS.n615 VSS.n613 0.0269375
R4446 VSS.n613 VSS.n611 0.0269375
R4447 VSS.n611 VSS.n609 0.0269375
R4448 VSS.n609 VSS.n607 0.0269375
R4449 VSS.n607 VSS.n605 0.0269375
R4450 VSS.n605 VSS.n603 0.0269375
R4451 VSS.n603 VSS.n601 0.0269375
R4452 VSS.n601 VSS.n599 0.0269375
R4453 VSS.n599 VSS.n597 0.0269375
R4454 VSS.n597 VSS.n595 0.0269375
R4455 VSS.n595 VSS.n593 0.0269375
R4456 VSS.n593 VSS.n591 0.0269375
R4457 VSS.n591 VSS.n589 0.0269375
R4458 VSS.n589 VSS.n587 0.0269375
R4459 VSS.n587 VSS.n585 0.0269375
R4460 VSS.n585 VSS.n583 0.0269375
R4461 VSS.n583 VSS.n581 0.0269375
R4462 VSS.n581 VSS.n579 0.0269375
R4463 VSS.n579 VSS.n577 0.0269375
R4464 VSS.n577 VSS.n575 0.0269375
R4465 VSS.n575 VSS.n573 0.0269375
R4466 VSS.n573 VSS.n571 0.0269375
R4467 VSS.n571 VSS.n569 0.0269375
R4468 VSS.n569 VSS.n567 0.0269375
R4469 VSS.n567 VSS.n565 0.0269375
R4470 VSS.n565 VSS.n563 0.0269375
R4471 VSS.n563 VSS.n561 0.0269375
R4472 VSS.n561 VSS.n559 0.0269375
R4473 VSS.n559 VSS.n557 0.0269375
R4474 VSS.n557 VSS.n555 0.0269375
R4475 VSS.n555 VSS.n553 0.0269375
R4476 VSS.n1545 VSS.n1543 0.0269375
R4477 VSS.n1547 VSS.n1545 0.0269375
R4478 VSS.n1549 VSS.n1547 0.0269375
R4479 VSS.n1551 VSS.n1549 0.0269375
R4480 VSS.n1553 VSS.n1551 0.0269375
R4481 VSS.n1745 VSS.n1553 0.0269375
R4482 VSS.n1012 VSS.n550 0.0269375
R4483 VSS.n550 VSS.n547 0.0269375
R4484 VSS.n547 VSS.n545 0.0269375
R4485 VSS.n545 VSS.n542 0.0269375
R4486 VSS.n542 VSS.n540 0.0269375
R4487 VSS.n540 VSS.n537 0.0269375
R4488 VSS.n537 VSS.n535 0.0269375
R4489 VSS.n535 VSS.n532 0.0269375
R4490 VSS.n532 VSS.n530 0.0269375
R4491 VSS.n530 VSS.n527 0.0269375
R4492 VSS.n527 VSS.n525 0.0269375
R4493 VSS.n525 VSS.n522 0.0269375
R4494 VSS.n522 VSS.n520 0.0269375
R4495 VSS.n520 VSS.n518 0.0269375
R4496 VSS.n518 VSS.n516 0.0269375
R4497 VSS.n516 VSS.n514 0.0269375
R4498 VSS.n514 VSS.n512 0.0269375
R4499 VSS.n512 VSS.n510 0.0269375
R4500 VSS.n510 VSS.n508 0.0269375
R4501 VSS.n508 VSS.n506 0.0269375
R4502 VSS.n506 VSS.n504 0.0269375
R4503 VSS.n504 VSS.n502 0.0269375
R4504 VSS.n502 VSS.n500 0.0269375
R4505 VSS.n500 VSS.n498 0.0269375
R4506 VSS.n498 VSS.n496 0.0269375
R4507 VSS.n496 VSS.n494 0.0269375
R4508 VSS.n494 VSS.n492 0.0269375
R4509 VSS.n492 VSS.n490 0.0269375
R4510 VSS.n490 VSS.n488 0.0269375
R4511 VSS.n488 VSS.n486 0.0269375
R4512 VSS.n486 VSS.n484 0.0269375
R4513 VSS.n484 VSS.n482 0.0269375
R4514 VSS.n482 VSS.n480 0.0269375
R4515 VSS.n480 VSS.n478 0.0269375
R4516 VSS.n478 VSS.n476 0.0269375
R4517 VSS.n476 VSS.n474 0.0269375
R4518 VSS.n474 VSS.n472 0.0269375
R4519 VSS.n472 VSS.n470 0.0269375
R4520 VSS.n470 VSS.n468 0.0269375
R4521 VSS.n468 VSS.n466 0.0269375
R4522 VSS.n466 VSS.n464 0.0269375
R4523 VSS.n464 VSS.n462 0.0269375
R4524 VSS.n462 VSS.n460 0.0269375
R4525 VSS.n460 VSS.n458 0.0269375
R4526 VSS.n458 VSS.n456 0.0269375
R4527 VSS.n456 VSS.n454 0.0269375
R4528 VSS.n454 VSS.n452 0.0269375
R4529 VSS.n452 VSS.n450 0.0269375
R4530 VSS.n450 VSS.n448 0.0269375
R4531 VSS.n448 VSS.n446 0.0269375
R4532 VSS.n446 VSS.n444 0.0269375
R4533 VSS.n444 VSS.n442 0.0269375
R4534 VSS.n442 VSS.n440 0.0269375
R4535 VSS.n440 VSS.n438 0.0269375
R4536 VSS.n438 VSS.n436 0.0269375
R4537 VSS.n436 VSS.n434 0.0269375
R4538 VSS.n434 VSS.n432 0.0269375
R4539 VSS.n1532 VSS.n1530 0.0269375
R4540 VSS.n1534 VSS.n1532 0.0269375
R4541 VSS.n1536 VSS.n1534 0.0269375
R4542 VSS.n1538 VSS.n1536 0.0269375
R4543 VSS.n1540 VSS.n1538 0.0269375
R4544 VSS.n1753 VSS.n1540 0.0269375
R4545 VSS.n1110 VSS.n410 0.0269375
R4546 VSS.n410 VSS.n408 0.0269375
R4547 VSS.n408 VSS.n405 0.0269375
R4548 VSS.n405 VSS.n402 0.0269375
R4549 VSS.n402 VSS.n400 0.0269375
R4550 VSS.n400 VSS.n397 0.0269375
R4551 VSS.n397 VSS.n395 0.0269375
R4552 VSS.n395 VSS.n392 0.0269375
R4553 VSS.n392 VSS.n390 0.0269375
R4554 VSS.n390 VSS.n387 0.0269375
R4555 VSS.n387 VSS.n385 0.0269375
R4556 VSS.n385 VSS.n382 0.0269375
R4557 VSS.n382 VSS.n380 0.0269375
R4558 VSS.n380 VSS.n377 0.0269375
R4559 VSS.n377 VSS.n375 0.0269375
R4560 VSS.n375 VSS.n372 0.0269375
R4561 VSS.n372 VSS.n370 0.0269375
R4562 VSS.n370 VSS.n367 0.0269375
R4563 VSS.n367 VSS.n365 0.0269375
R4564 VSS.n365 VSS.n362 0.0269375
R4565 VSS.n362 VSS.n360 0.0269375
R4566 VSS.n360 VSS.n357 0.0269375
R4567 VSS.n357 VSS.n355 0.0269375
R4568 VSS.n355 VSS.n352 0.0269375
R4569 VSS.n352 VSS.n350 0.0269375
R4570 VSS.n350 VSS.n348 0.0269375
R4571 VSS.n348 VSS.n346 0.0269375
R4572 VSS.n346 VSS.n344 0.0269375
R4573 VSS.n344 VSS.n342 0.0269375
R4574 VSS.n342 VSS.n340 0.0269375
R4575 VSS.n340 VSS.n338 0.0269375
R4576 VSS.n338 VSS.n336 0.0269375
R4577 VSS.n336 VSS.n334 0.0269375
R4578 VSS.n334 VSS.n332 0.0269375
R4579 VSS.n332 VSS.n330 0.0269375
R4580 VSS.n330 VSS.n328 0.0269375
R4581 VSS.n328 VSS.n326 0.0269375
R4582 VSS.n326 VSS.n324 0.0269375
R4583 VSS.n324 VSS.n322 0.0269375
R4584 VSS.n322 VSS.n320 0.0269375
R4585 VSS.n320 VSS.n318 0.0269375
R4586 VSS.n318 VSS.n316 0.0269375
R4587 VSS.n316 VSS.n314 0.0269375
R4588 VSS.n314 VSS.n312 0.0269375
R4589 VSS.n312 VSS.n310 0.0269375
R4590 VSS.n310 VSS.n308 0.0269375
R4591 VSS.n308 VSS.n306 0.0269375
R4592 VSS.n306 VSS.n304 0.0269375
R4593 VSS.n304 VSS.n302 0.0269375
R4594 VSS.n302 VSS.n300 0.0269375
R4595 VSS.n300 VSS.n298 0.0269375
R4596 VSS.n298 VSS.n296 0.0269375
R4597 VSS.n296 VSS.n294 0.0269375
R4598 VSS.n294 VSS.n292 0.0269375
R4599 VSS.n292 VSS.n290 0.0269375
R4600 VSS.n290 VSS.n288 0.0269375
R4601 VSS.n288 VSS.n286 0.0269375
R4602 VSS.n1413 VSS.n1411 0.0269375
R4603 VSS.n1415 VSS.n1413 0.0269375
R4604 VSS.n1417 VSS.n1415 0.0269375
R4605 VSS.n1419 VSS.n1417 0.0269375
R4606 VSS.n1421 VSS.n1419 0.0269375
R4607 VSS.n1821 VSS.n1421 0.0269375
R4608 VSS.n1173 VSS.n283 0.0269375
R4609 VSS.n283 VSS.n280 0.0269375
R4610 VSS.n280 VSS.n278 0.0269375
R4611 VSS.n278 VSS.n275 0.0269375
R4612 VSS.n275 VSS.n273 0.0269375
R4613 VSS.n273 VSS.n270 0.0269375
R4614 VSS.n270 VSS.n268 0.0269375
R4615 VSS.n268 VSS.n265 0.0269375
R4616 VSS.n265 VSS.n263 0.0269375
R4617 VSS.n263 VSS.n260 0.0269375
R4618 VSS.n260 VSS.n258 0.0269375
R4619 VSS.n258 VSS.n255 0.0269375
R4620 VSS.n255 VSS.n253 0.0269375
R4621 VSS.n253 VSS.n251 0.0269375
R4622 VSS.n251 VSS.n249 0.0269375
R4623 VSS.n249 VSS.n247 0.0269375
R4624 VSS.n247 VSS.n245 0.0269375
R4625 VSS.n245 VSS.n243 0.0269375
R4626 VSS.n243 VSS.n241 0.0269375
R4627 VSS.n241 VSS.n239 0.0269375
R4628 VSS.n239 VSS.n237 0.0269375
R4629 VSS.n237 VSS.n235 0.0269375
R4630 VSS.n235 VSS.n233 0.0269375
R4631 VSS.n233 VSS.n231 0.0269375
R4632 VSS.n231 VSS.n229 0.0269375
R4633 VSS.n229 VSS.n227 0.0269375
R4634 VSS.n227 VSS.n225 0.0269375
R4635 VSS.n225 VSS.n223 0.0269375
R4636 VSS.n223 VSS.n221 0.0269375
R4637 VSS.n221 VSS.n219 0.0269375
R4638 VSS.n219 VSS.n217 0.0269375
R4639 VSS.n217 VSS.n215 0.0269375
R4640 VSS.n215 VSS.n213 0.0269375
R4641 VSS.n213 VSS.n211 0.0269375
R4642 VSS.n211 VSS.n209 0.0269375
R4643 VSS.n209 VSS.n207 0.0269375
R4644 VSS.n207 VSS.n205 0.0269375
R4645 VSS.n205 VSS.n203 0.0269375
R4646 VSS.n203 VSS.n201 0.0269375
R4647 VSS.n201 VSS.n199 0.0269375
R4648 VSS.n199 VSS.n197 0.0269375
R4649 VSS.n197 VSS.n195 0.0269375
R4650 VSS.n195 VSS.n193 0.0269375
R4651 VSS.n193 VSS.n191 0.0269375
R4652 VSS.n191 VSS.n189 0.0269375
R4653 VSS.n189 VSS.n187 0.0269375
R4654 VSS.n187 VSS.n185 0.0269375
R4655 VSS.n185 VSS.n183 0.0269375
R4656 VSS.n183 VSS.n181 0.0269375
R4657 VSS.n181 VSS.n179 0.0269375
R4658 VSS.n179 VSS.n177 0.0269375
R4659 VSS.n177 VSS.n175 0.0269375
R4660 VSS.n175 VSS.n173 0.0269375
R4661 VSS.n173 VSS.n171 0.0269375
R4662 VSS.n171 VSS.n169 0.0269375
R4663 VSS.n169 VSS.n167 0.0269375
R4664 VSS.n167 VSS.n165 0.0269375
R4665 VSS.n1400 VSS.n1398 0.0269375
R4666 VSS.n1402 VSS.n1400 0.0269375
R4667 VSS.n1404 VSS.n1402 0.0269375
R4668 VSS.n1406 VSS.n1404 0.0269375
R4669 VSS.n1408 VSS.n1406 0.0269375
R4670 VSS.n1829 VSS.n1408 0.0269375
R4671 VSS.n1279 VSS.n1277 0.0269375
R4672 VSS.n1282 VSS.n1279 0.0269375
R4673 VSS.n1284 VSS.n1282 0.0269375
R4674 VSS.n1287 VSS.n1284 0.0269375
R4675 VSS.n1289 VSS.n1287 0.0269375
R4676 VSS.n2897 VSS.n2895 0.0269375
R4677 VSS.n2895 VSS.n2892 0.0269375
R4678 VSS.n2892 VSS.n2889 0.0269375
R4679 VSS.n2889 VSS.n2886 0.0269375
R4680 VSS.n2886 VSS.n2883 0.0269375
R4681 VSS.n2883 VSS.n2881 0.0269375
R4682 VSS.n2020 VSS.n2017 0.0269375
R4683 VSS.n2017 VSS.n2015 0.0269375
R4684 VSS.n2015 VSS.n2012 0.0269375
R4685 VSS.n2012 VSS.n2010 0.0269375
R4686 VSS.n2010 VSS.n2007 0.0269375
R4687 VSS.n2007 VSS.n2005 0.0269375
R4688 VSS.n2005 VSS.n2002 0.0269375
R4689 VSS.n2002 VSS.n2000 0.0269375
R4690 VSS.n2000 VSS.n1997 0.0269375
R4691 VSS.n1997 VSS.n1995 0.0269375
R4692 VSS.n1995 VSS.n1992 0.0269375
R4693 VSS.n1992 VSS.n1990 0.0269375
R4694 VSS.n1990 VSS.n1987 0.0269375
R4695 VSS.n1987 VSS.n1985 0.0269375
R4696 VSS.n1985 VSS.n1982 0.0269375
R4697 VSS.n1982 VSS.n1980 0.0269375
R4698 VSS.n1980 VSS.n1977 0.0269375
R4699 VSS.n1977 VSS.n1975 0.0269375
R4700 VSS.n1975 VSS.n1973 0.0269375
R4701 VSS.n1973 VSS.n1971 0.0269375
R4702 VSS.n1971 VSS.n1969 0.0269375
R4703 VSS.n1969 VSS.n1967 0.0269375
R4704 VSS.n1967 VSS.n1965 0.0269375
R4705 VSS.n1965 VSS.n1963 0.0269375
R4706 VSS.n1963 VSS.n1961 0.0269375
R4707 VSS.n1961 VSS.n1959 0.0269375
R4708 VSS.n1959 VSS.n1957 0.0269375
R4709 VSS.n1957 VSS.n1955 0.0269375
R4710 VSS.n1955 VSS.n1953 0.0269375
R4711 VSS.n1953 VSS.n1951 0.0269375
R4712 VSS.n1951 VSS.n1949 0.0269375
R4713 VSS.n1949 VSS.n1947 0.0269375
R4714 VSS.n1947 VSS.n1945 0.0269375
R4715 VSS.n1945 VSS.n1943 0.0269375
R4716 VSS.n1943 VSS.n1941 0.0269375
R4717 VSS.n1941 VSS.n1939 0.0269375
R4718 VSS.n1939 VSS.n1937 0.0269375
R4719 VSS.n1937 VSS.n1935 0.0269375
R4720 VSS.n1935 VSS.n1933 0.0269375
R4721 VSS.n1933 VSS.n1931 0.0269375
R4722 VSS.n1931 VSS.n1929 0.0269375
R4723 VSS.n1929 VSS.n1927 0.0269375
R4724 VSS.n1927 VSS.n1925 0.0269375
R4725 VSS.n1925 VSS.n1923 0.0269375
R4726 VSS.n1923 VSS.n1921 0.0269375
R4727 VSS.n1921 VSS.n1919 0.0269375
R4728 VSS.n1919 VSS.n1917 0.0269375
R4729 VSS.n1917 VSS.n1915 0.0269375
R4730 VSS.n1915 VSS.n1913 0.0269375
R4731 VSS.n1913 VSS.n1911 0.0269375
R4732 VSS.n1911 VSS.n1909 0.0269375
R4733 VSS.n1909 VSS.n1907 0.0269375
R4734 VSS.n1907 VSS.n1905 0.0269375
R4735 VSS.n1905 VSS.n1903 0.0269375
R4736 VSS.n1903 VSS.n1901 0.0269375
R4737 VSS.n1677 VSS.n1675 0.0269375
R4738 VSS.n1679 VSS.n1677 0.0269375
R4739 VSS.n1681 VSS.n1679 0.0269375
R4740 VSS.n1683 VSS.n1681 0.0269375
R4741 VSS.n1685 VSS.n1683 0.0269375
R4742 VSS.n1697 VSS.n1695 0.0269375
R4743 VSS.n1699 VSS.n1697 0.0269375
R4744 VSS.n1704 VSS.n1702 0.0269375
R4745 VSS.n1706 VSS.n1704 0.0269375
R4746 VSS.n1708 VSS.n1706 0.0269375
R4747 VSS.n1710 VSS.n1708 0.0269375
R4748 VSS.n1712 VSS.n1710 0.0269375
R4749 VSS.n1714 VSS.n1712 0.0269375
R4750 VSS.n1716 VSS.n1714 0.0269375
R4751 VSS.n1718 VSS.n1716 0.0269375
R4752 VSS.n1720 VSS.n1718 0.0269375
R4753 VSS.n1722 VSS.n1720 0.0269375
R4754 VSS.n1724 VSS.n1722 0.0269375
R4755 VSS.n1726 VSS.n1724 0.0269375
R4756 VSS.n1728 VSS.n1726 0.0269375
R4757 VSS.n1736 VSS.n1734 0.0269375
R4758 VSS.n1738 VSS.n1736 0.0269375
R4759 VSS.n1740 VSS.n1738 0.0269375
R4760 VSS.n1742 VSS.n1740 0.0269375
R4761 VSS.n1744 VSS.n1742 0.0269375
R4762 VSS.n1757 VSS.n1755 0.0269375
R4763 VSS.n1759 VSS.n1757 0.0269375
R4764 VSS.n1761 VSS.n1759 0.0269375
R4765 VSS.n1763 VSS.n1761 0.0269375
R4766 VSS.n1765 VSS.n1763 0.0269375
R4767 VSS.n1773 VSS.n1771 0.0269375
R4768 VSS.n1775 VSS.n1773 0.0269375
R4769 VSS.n1777 VSS.n1775 0.0269375
R4770 VSS.n1779 VSS.n1777 0.0269375
R4771 VSS.n1781 VSS.n1779 0.0269375
R4772 VSS.n1783 VSS.n1781 0.0269375
R4773 VSS.n1785 VSS.n1783 0.0269375
R4774 VSS.n1787 VSS.n1785 0.0269375
R4775 VSS.n1789 VSS.n1787 0.0269375
R4776 VSS.n1791 VSS.n1789 0.0269375
R4777 VSS.n1793 VSS.n1791 0.0269375
R4778 VSS.n1795 VSS.n1793 0.0269375
R4779 VSS.n1797 VSS.n1795 0.0269375
R4780 VSS.n1802 VSS.n1800 0.0269375
R4781 VSS.n1804 VSS.n1802 0.0269375
R4782 VSS.n1812 VSS.n1810 0.0269375
R4783 VSS.n1814 VSS.n1812 0.0269375
R4784 VSS.n1816 VSS.n1814 0.0269375
R4785 VSS.n1818 VSS.n1816 0.0269375
R4786 VSS.n1820 VSS.n1818 0.0269375
R4787 VSS.n1833 VSS.n1831 0.0269375
R4788 VSS.n1835 VSS.n1833 0.0269375
R4789 VSS.n1837 VSS.n1835 0.0269375
R4790 VSS.n1839 VSS.n1837 0.0269375
R4791 VSS.n1841 VSS.n1839 0.0269375
R4792 VSS.n1849 VSS.n1847 0.0269375
R4793 VSS.n1851 VSS.n1849 0.0269375
R4794 VSS.n1856 VSS.n1854 0.0269375
R4795 VSS.n1858 VSS.n1856 0.0269375
R4796 VSS.n1860 VSS.n1858 0.0269375
R4797 VSS.n1862 VSS.n1860 0.0269375
R4798 VSS.n1864 VSS.n1862 0.0269375
R4799 VSS.n1866 VSS.n1864 0.0269375
R4800 VSS.n1868 VSS.n1866 0.0269375
R4801 VSS.n1870 VSS.n1868 0.0269375
R4802 VSS.n1872 VSS.n1870 0.0269375
R4803 VSS.n1874 VSS.n1872 0.0269375
R4804 VSS.n1876 VSS.n1874 0.0269375
R4805 VSS.n1878 VSS.n1876 0.0269375
R4806 VSS.n1880 VSS.n1878 0.0269375
R4807 VSS.n1888 VSS.n1886 0.0269375
R4808 VSS.n1890 VSS.n1888 0.0269375
R4809 VSS.n1892 VSS.n1890 0.0269375
R4810 VSS.n1894 VSS.n1892 0.0269375
R4811 VSS.n1896 VSS.n1894 0.0269375
R4812 VSS.n857 VSS.n854 0.0269375
R4813 VSS.n860 VSS.n857 0.0269375
R4814 VSS.n863 VSS.n860 0.0269375
R4815 VSS.n866 VSS.n863 0.0269375
R4816 VSS.n869 VSS.n866 0.0269375
R4817 VSS.n880 VSS.n877 0.0269375
R4818 VSS.n883 VSS.n880 0.0269375
R4819 VSS.n886 VSS.n883 0.0269375
R4820 VSS.n889 VSS.n886 0.0269375
R4821 VSS.n892 VSS.n889 0.0269375
R4822 VSS.n895 VSS.n892 0.0269375
R4823 VSS.n898 VSS.n895 0.0269375
R4824 VSS.n901 VSS.n898 0.0269375
R4825 VSS.n904 VSS.n901 0.0269375
R4826 VSS.n907 VSS.n904 0.0269375
R4827 VSS.n910 VSS.n907 0.0269375
R4828 VSS.n913 VSS.n910 0.0269375
R4829 VSS.n916 VSS.n913 0.0269375
R4830 VSS.n919 VSS.n916 0.0269375
R4831 VSS.n922 VSS.n919 0.0269375
R4832 VSS.n925 VSS.n922 0.0269375
R4833 VSS.n936 VSS.n933 0.0269375
R4834 VSS.n939 VSS.n936 0.0269375
R4835 VSS.n942 VSS.n939 0.0269375
R4836 VSS.n945 VSS.n942 0.0269375
R4837 VSS.n948 VSS.n945 0.0269375
R4838 VSS.n1018 VSS.n1015 0.0269375
R4839 VSS.n1021 VSS.n1018 0.0269375
R4840 VSS.n1024 VSS.n1021 0.0269375
R4841 VSS.n1027 VSS.n1024 0.0269375
R4842 VSS.n1030 VSS.n1027 0.0269375
R4843 VSS.n1041 VSS.n1038 0.0269375
R4844 VSS.n1044 VSS.n1041 0.0269375
R4845 VSS.n1047 VSS.n1044 0.0269375
R4846 VSS.n1050 VSS.n1047 0.0269375
R4847 VSS.n1053 VSS.n1050 0.0269375
R4848 VSS.n1056 VSS.n1053 0.0269375
R4849 VSS.n1059 VSS.n1056 0.0269375
R4850 VSS.n1062 VSS.n1059 0.0269375
R4851 VSS.n1065 VSS.n1062 0.0269375
R4852 VSS.n1068 VSS.n1065 0.0269375
R4853 VSS.n1071 VSS.n1068 0.0269375
R4854 VSS.n1074 VSS.n1071 0.0269375
R4855 VSS.n1077 VSS.n1074 0.0269375
R4856 VSS.n1080 VSS.n1077 0.0269375
R4857 VSS.n1083 VSS.n1080 0.0269375
R4858 VSS.n1086 VSS.n1083 0.0269375
R4859 VSS.n1097 VSS.n1094 0.0269375
R4860 VSS.n1100 VSS.n1097 0.0269375
R4861 VSS.n1103 VSS.n1100 0.0269375
R4862 VSS.n1106 VSS.n1103 0.0269375
R4863 VSS.n1109 VSS.n1106 0.0269375
R4864 VSS.n1179 VSS.n1176 0.0269375
R4865 VSS.n1182 VSS.n1179 0.0269375
R4866 VSS.n1185 VSS.n1182 0.0269375
R4867 VSS.n1188 VSS.n1185 0.0269375
R4868 VSS.n1191 VSS.n1188 0.0269375
R4869 VSS.n1202 VSS.n1199 0.0269375
R4870 VSS.n1205 VSS.n1202 0.0269375
R4871 VSS.n1208 VSS.n1205 0.0269375
R4872 VSS.n1211 VSS.n1208 0.0269375
R4873 VSS.n1214 VSS.n1211 0.0269375
R4874 VSS.n1217 VSS.n1214 0.0269375
R4875 VSS.n1220 VSS.n1217 0.0269375
R4876 VSS.n1223 VSS.n1220 0.0269375
R4877 VSS.n1226 VSS.n1223 0.0269375
R4878 VSS.n1229 VSS.n1226 0.0269375
R4879 VSS.n1232 VSS.n1229 0.0269375
R4880 VSS.n1235 VSS.n1232 0.0269375
R4881 VSS.n1238 VSS.n1235 0.0269375
R4882 VSS.n1241 VSS.n1238 0.0269375
R4883 VSS.n1244 VSS.n1241 0.0269375
R4884 VSS.n1247 VSS.n1244 0.0269375
R4885 VSS.n1258 VSS.n1255 0.0269375
R4886 VSS.n1261 VSS.n1258 0.0269375
R4887 VSS.n1264 VSS.n1261 0.0269375
R4888 VSS.n1267 VSS.n1264 0.0269375
R4889 VSS.n1270 VSS.n1267 0.0269375
R4890 VSS.n2606 VSS.n2603 0.0269375
R4891 VSS.n2609 VSS.n2606 0.0269375
R4892 VSS.n2612 VSS.n2609 0.0269375
R4893 VSS.n2615 VSS.n2612 0.0269375
R4894 VSS.n2617 VSS.n2615 0.0269375
R4895 VSS.n2619 VSS.n2617 0.0269375
R4896 VSS.n2624 VSS.n2622 0.0269375
R4897 VSS.n2626 VSS.n2624 0.0269375
R4898 VSS.n2631 VSS.n2629 0.0269375
R4899 VSS.n2633 VSS.n2631 0.0269375
R4900 VSS.n2635 VSS.n2633 0.0269375
R4901 VSS.n2637 VSS.n2635 0.0269375
R4902 VSS.n2639 VSS.n2637 0.0269375
R4903 VSS.n2644 VSS.n2642 0.0269375
R4904 VSS.n2646 VSS.n2644 0.0269375
R4905 VSS.n2648 VSS.n2646 0.0269375
R4906 VSS.n2650 VSS.n2648 0.0269375
R4907 VSS.n2652 VSS.n2650 0.0269375
R4908 VSS.n2654 VSS.n2652 0.0269375
R4909 VSS.n2659 VSS.n2657 0.0269375
R4910 VSS.n2661 VSS.n2659 0.0269375
R4911 VSS.n2663 VSS.n2661 0.0269375
R4912 VSS.n2665 VSS.n2663 0.0269375
R4913 VSS.n2667 VSS.n2665 0.0269375
R4914 VSS.n2669 VSS.n2667 0.0269375
R4915 VSS.n2671 VSS.n2669 0.0269375
R4916 VSS.n2676 VSS.n2674 0.0269375
R4917 VSS.n2678 VSS.n2676 0.0269375
R4918 VSS.n2680 VSS.n2678 0.0269375
R4919 VSS.n2682 VSS.n2680 0.0269375
R4920 VSS.n2684 VSS.n2682 0.0269375
R4921 VSS.n2689 VSS.n2687 0.0269375
R4922 VSS.n2691 VSS.n2689 0.0269375
R4923 VSS.n2693 VSS.n2691 0.0269375
R4924 VSS.n2695 VSS.n2693 0.0269375
R4925 VSS.n2697 VSS.n2695 0.0269375
R4926 VSS.n2699 VSS.n2697 0.0269375
R4927 VSS.n2701 VSS.n2699 0.0269375
R4928 VSS.n2703 VSS.n2701 0.0269375
R4929 VSS.n2705 VSS.n2703 0.0269375
R4930 VSS.n2707 VSS.n2705 0.0269375
R4931 VSS.n2712 VSS.n2710 0.0269375
R4932 VSS.n2714 VSS.n2712 0.0269375
R4933 VSS.n2719 VSS.n2717 0.0269375
R4934 VSS.n2721 VSS.n2719 0.0269375
R4935 VSS.n2723 VSS.n2721 0.0269375
R4936 VSS.n2725 VSS.n2723 0.0269375
R4937 VSS.n2727 VSS.n2725 0.0269375
R4938 VSS.n2729 VSS.n2727 0.0269375
R4939 VSS.n3013 VSS.n3010 0.0269375
R4940 VSS.n3010 VSS.n3007 0.0269375
R4941 VSS.n3007 VSS.n3004 0.0269375
R4942 VSS.n3004 VSS.n3001 0.0269375
R4943 VSS.n3001 VSS.n2998 0.0269375
R4944 VSS.n2998 VSS.n2995 0.0269375
R4945 VSS.n2995 VSS.n2992 0.0269375
R4946 VSS.n2992 VSS.n2989 0.0269375
R4947 VSS.n2989 VSS.n2986 0.0269375
R4948 VSS.n2986 VSS.n2983 0.0269375
R4949 VSS.n2983 VSS.n2980 0.0269375
R4950 VSS.n2980 VSS.n2977 0.0269375
R4951 VSS.n2977 VSS.n2974 0.0269375
R4952 VSS.n2974 VSS.n2971 0.0269375
R4953 VSS.n2971 VSS.n2968 0.0269375
R4954 VSS.n2968 VSS.n2965 0.0269375
R4955 VSS.n2965 VSS.n2962 0.0269375
R4956 VSS.n2962 VSS.n2959 0.0269375
R4957 VSS.n2959 VSS.n2956 0.0269375
R4958 VSS.n2956 VSS.n2953 0.0269375
R4959 VSS.n2953 VSS.n2950 0.0269375
R4960 VSS.n2950 VSS.n2947 0.0269375
R4961 VSS.n2947 VSS.n2944 0.0269375
R4962 VSS.n2944 VSS.n2941 0.0269375
R4963 VSS.n2597 VSS.n2594 0.0269375
R4964 VSS.n2600 VSS.n2597 0.0269375
R4965 VSS.n3027 VSS.n3025 0.0269375
R4966 VSS.n3030 VSS.n3027 0.0269375
R4967 VSS.n3032 VSS.n3030 0.0269375
R4968 VSS.n3035 VSS.n3032 0.0269375
R4969 VSS.n3039 VSS.n3035 0.0269375
R4970 VSS.n3042 VSS.n3039 0.0269375
R4971 VSS.n3049 VSS.n3046 0.0269375
R4972 VSS.n3052 VSS.n3049 0.0269375
R4973 VSS.n3059 VSS.n3056 0.0269375
R4974 VSS.n3062 VSS.n3059 0.0269375
R4975 VSS.n3065 VSS.n3062 0.0269375
R4976 VSS.n3068 VSS.n3065 0.0269375
R4977 VSS.n3071 VSS.n3068 0.0269375
R4978 VSS.n3078 VSS.n3075 0.0269375
R4979 VSS.n3081 VSS.n3078 0.0269375
R4980 VSS.n3084 VSS.n3081 0.0269375
R4981 VSS.n3087 VSS.n3084 0.0269375
R4982 VSS.n3090 VSS.n3087 0.0269375
R4983 VSS.n3093 VSS.n3090 0.0269375
R4984 VSS.n3100 VSS.n3097 0.0269375
R4985 VSS.n3103 VSS.n3100 0.0269375
R4986 VSS.n3106 VSS.n3103 0.0269375
R4987 VSS.n3109 VSS.n3106 0.0269375
R4988 VSS.n3112 VSS.n3109 0.0269375
R4989 VSS.n3115 VSS.n3112 0.0269375
R4990 VSS.n3118 VSS.n3115 0.0269375
R4991 VSS.n3125 VSS.n3122 0.0269375
R4992 VSS.n3128 VSS.n3125 0.0269375
R4993 VSS.n3131 VSS.n3128 0.0269375
R4994 VSS.n3134 VSS.n3131 0.0269375
R4995 VSS.n3137 VSS.n3134 0.0269375
R4996 VSS.n3144 VSS.n3141 0.0269375
R4997 VSS.n3147 VSS.n3144 0.0269375
R4998 VSS.n3150 VSS.n3147 0.0269375
R4999 VSS.n3153 VSS.n3150 0.0269375
R5000 VSS.n3156 VSS.n3153 0.0269375
R5001 VSS.n3159 VSS.n3156 0.0269375
R5002 VSS.n3170 VSS.n3167 0.0269375
R5003 VSS.n3181 VSS.n3178 0.0269375
R5004 VSS.n3184 VSS.n3181 0.0269375
R5005 VSS.n3191 VSS.n3188 0.0269375
R5006 VSS.n3194 VSS.n3191 0.0269375
R5007 VSS.n3197 VSS.n3194 0.0269375
R5008 VSS.n3200 VSS.n3197 0.0269375
R5009 VSS.n3203 VSS.n3200 0.0269375
R5010 VSS.n3206 VSS.n3203 0.0269375
R5011 VSS.n2877 VSS.n2874 0.0269375
R5012 VSS.n2874 VSS.n2872 0.0269375
R5013 VSS.n2863 VSS.n2861 0.0269375
R5014 VSS.n2861 VSS.n2858 0.0269375
R5015 VSS.n2858 VSS.n2856 0.0269375
R5016 VSS.n2856 VSS.n2853 0.0269375
R5017 VSS.n2853 VSS.n2851 0.0269375
R5018 VSS.n2851 VSS.n2848 0.0269375
R5019 VSS.n2848 VSS.n2846 0.0269375
R5020 VSS.n2846 VSS.n2843 0.0269375
R5021 VSS.n2843 VSS.n2841 0.0269375
R5022 VSS.n2870 VSS.n2863 0.0266563
R5023 VSS.n2878 VSS.n2877 0.0260938
R5024 VSS.n2105 VSS.n2104 0.0258125
R5025 VSS.n3163 VSS.n3160 0.0255312
R5026 VSS.n135 VSS.n133 0.0246875
R5027 VSS.n2814 VSS.n2812 0.0246875
R5028 VSS.n3207 VSS.n2897 0.0244062
R5029 VSS.n3023 VSS.n3013 0.0244062
R5030 VSS.n2601 VSS.n2600 0.0244062
R5031 VSS.n2841 VSS.n2839 0.0244062
R5032 VSS.n2472 VSS.n2465 0.024125
R5033 VSS.n2836 VSS.n2739 0.024125
R5034 VSS.n120 VSS.n119 0.024125
R5035 VSS.n1700 VSS.n1699 0.024125
R5036 VSS.n1800 VSS.n1798 0.024125
R5037 VSS.n1852 VSS.n1851 0.024125
R5038 VSS.n2622 VSS.n2620 0.0238437
R5039 VSS.n2674 VSS.n2672 0.0238437
R5040 VSS.n2715 VSS.n2714 0.0238437
R5041 VSS.n3046 VSS.n3043 0.0238437
R5042 VSS.n3122 VSS.n3119 0.0238437
R5043 VSS.n3185 VSS.n3184 0.0238437
R5044 VSS.n1692 VSS.n1690 0.0235625
R5045 VSS.n1732 VSS.n1731 0.0235625
R5046 VSS.n1768 VSS.n1766 0.0235625
R5047 VSS.n1808 VSS.n1807 0.0235625
R5048 VSS.n1844 VSS.n1842 0.0235625
R5049 VSS.n1884 VSS.n1883 0.0235625
R5050 VSS.n873 VSS.n870 0.0235625
R5051 VSS.n930 VSS.n929 0.0235625
R5052 VSS.n1034 VSS.n1031 0.0235625
R5053 VSS.n1091 VSS.n1090 0.0235625
R5054 VSS.n1195 VSS.n1192 0.0235625
R5055 VSS.n1252 VSS.n1251 0.0235625
R5056 VSS.n2523 VSS.n2517 0.023
R5057 VSS.n1693 VSS.n1692 0.0224375
R5058 VSS.n1731 VSS.n1729 0.0224375
R5059 VSS.n1769 VSS.n1768 0.0224375
R5060 VSS.n1807 VSS.n1805 0.0224375
R5061 VSS.n1845 VSS.n1844 0.0224375
R5062 VSS.n1883 VSS.n1881 0.0224375
R5063 VSS.n874 VSS.n873 0.0224375
R5064 VSS.n929 VSS.n926 0.0224375
R5065 VSS.n1035 VSS.n1034 0.0224375
R5066 VSS.n1090 VSS.n1087 0.0224375
R5067 VSS.n1196 VSS.n1195 0.0224375
R5068 VSS.n1251 VSS.n1248 0.0224375
R5069 VSS.n2640 VSS.n2639 0.0221563
R5070 VSS.n3072 VSS.n3071 0.0221563
R5071 VSS.n2771 VSS.n2770 0.0213125
R5072 VSS.n3569 VSS.n3568 0.0213125
R5073 VSS.n2382 VSS.n2379 0.0213125
R5074 VSS.n2102 VSS.n2100 0.0213125
R5075 VSS.n2148 VSS.n2147 0.0213125
R5076 VSS.n3371 VSS.n3370 0.0213125
R5077 VSS.n2575 VSS.n2574 0.0210419
R5078 VSS.n2555 VSS.n2554 0.0210419
R5079 VSS.n3523 VSS.n3522 0.02075
R5080 VSS.n3218 VSS.n2543 0.019625
R5081 VSS.n3312 VSS.n3311 0.019625
R5082 VSS.n2141 VSS.n2139 0.019625
R5083 VSS.n3334 VSS.n2410 0.0195
R5084 VSS.n2657 VSS.n2655 0.0193437
R5085 VSS.n3097 VSS.n3094 0.0193437
R5086 VSS.n3174 VSS.n3171 0.0193437
R5087 VSS.n2484 VSS.n2481 0.0190625
R5088 VSS.n2488 VSS.n2487 0.0190625
R5089 VSS.n2830 VSS.n2829 0.0190625
R5090 VSS.n2827 VSS.n2825 0.0190625
R5091 VSS.n3589 VSS.n3587 0.0190625
R5092 VSS.n3593 VSS.n3591 0.0190625
R5093 VSS.n3655 VSS.n3654 0.0190625
R5094 VSS.n3651 VSS.n3648 0.0190625
R5095 VSS.n3164 VSS.n3163 0.0182187
R5096 VSS.n2629 VSS.n2627 0.0176563
R5097 VSS.n2708 VSS.n2707 0.0176563
R5098 VSS.n3056 VSS.n3053 0.0176563
R5099 VSS.n3175 VSS.n3174 0.0176563
R5100 VSS.n2881 VSS.n2878 0.0170938
R5101 VSS.n1577 VSS.n1576 0.0167343
R5102 VSS.n1597 VSS.n1596 0.0167343
R5103 VSS.n1641 VSS.n1640 0.0167343
R5104 VSS.n1632 VSS.n1631 0.0167343
R5105 VSS.n1617 VSS.n1616 0.0167343
R5106 VSS.n1445 VSS.n1444 0.0167343
R5107 VSS.n1509 VSS.n1508 0.0167343
R5108 VSS.n1500 VSS.n1499 0.0167343
R5109 VSS.n1485 VSS.n1484 0.0167343
R5110 VSS.n1465 VSS.n1464 0.0167343
R5111 VSS.n1313 VSS.n1312 0.0167343
R5112 VSS.n1333 VSS.n1332 0.0167343
R5113 VSS.n1377 VSS.n1376 0.0167343
R5114 VSS.n1368 VSS.n1367 0.0167343
R5115 VSS.n1353 VSS.n1352 0.0167343
R5116 VSS.n2872 VSS.n2870 0.0165313
R5117 VSS.n2048 VSS.n2021 0.01625
R5118 VSS.n1673 VSS.n1672 0.01625
R5119 VSS.n1749 VSS.n1745 0.01625
R5120 VSS.n1753 VSS.n1752 0.01625
R5121 VSS.n1825 VSS.n1821 0.01625
R5122 VSS.n1829 VSS.n1828 0.01625
R5123 VSS.n1901 VSS.n1900 0.01625
R5124 VSS.n851 VSS.n850 0.01625
R5125 VSS.n977 VSS.n949 0.01625
R5126 VSS.n1012 VSS.n1011 0.01625
R5127 VSS.n1138 VSS.n1110 0.01625
R5128 VSS.n1173 VSS.n1172 0.01625
R5129 VSS.n1277 VSS.n1276 0.01625
R5130 VSS.n4031 VSS.n4028 0.01625
R5131 VSS.n4018 VSS.n4017 0.01625
R5132 VSS.n96 VSS.n94 0.01625
R5133 VSS.n87 VSS.n86 0.01625
R5134 VSS.n2685 VSS.n2684 0.0159688
R5135 VSS.n3138 VSS.n3137 0.0159688
R5136 VSS.n4011 VSS.n4008 0.0153235
R5137 VSS.n4004 VSS.n4003 0.0153235
R5138 VSS.n2407 VSS.n2406 0.0145
R5139 VSS.n2601 VSS.n2591 0.0142813
R5140 VSS.n2839 VSS.n2838 0.0142813
R5141 VSS.n3023 VSS.n3022 0.0142813
R5142 VSS.n3213 VSS.n3207 0.0142813
R5143 VSS.n2878 VSS.n2550 0.0142813
R5144 VSS.n2870 VSS.n2869 0.0142813
R5145 VSS.n3765 VSS.n3764 0.0140074
R5146 VSS.n2158 VSS.n2156 0.014
R5147 VSS.n3332 VSS.n3267 0.0139958
R5148 VSS.n2021 VSS.n2020 0.0134375
R5149 VSS.n2817 VSS.n2816 0.0134375
R5150 VSS.n2603 VSS.n2601 0.0131563
R5151 VSS.n2839 VSS.n2729 0.0131563
R5152 VSS.n3025 VSS.n3023 0.0131563
R5153 VSS.n3207 VSS.n3206 0.0131563
R5154 VSS.n3221 VSS.n3218 0.012875
R5155 VSS.n2260 VSS.n2258 0.01175
R5156 VSS.n2362 VSS.n2343 0.01175
R5157 VSS.n60 VSS.n59 0.01175
R5158 VSS.n3982 VSS.n3980 0.01175
R5159 VSS.n2160 VSS.n2158 0.01175
R5160 VSS VSS.n2242 0.01175
R5161 VSS.n2687 VSS.n2685 0.0114688
R5162 VSS.n3141 VSS.n3138 0.0114688
R5163 VSS.n1675 VSS.n1673 0.0111875
R5164 VSS.n1745 VSS.n1744 0.0111875
R5165 VSS.n1755 VSS.n1753 0.0111875
R5166 VSS.n1821 VSS.n1820 0.0111875
R5167 VSS.n1831 VSS.n1829 0.0111875
R5168 VSS.n1901 VSS.n1896 0.0111875
R5169 VSS.n854 VSS.n851 0.0111875
R5170 VSS.n949 VSS.n948 0.0111875
R5171 VSS.n1015 VSS.n1012 0.0111875
R5172 VSS.n1110 VSS.n1109 0.0111875
R5173 VSS.n1176 VSS.n1173 0.0111875
R5174 VSS.n1277 VSS.n1270 0.0111875
R5175 VSS.n2762 VSS.n2760 0.0111875
R5176 VSS.n3560 VSS.n3558 0.0111875
R5177 VSS.n2627 VSS.n2626 0.00978125
R5178 VSS.n2710 VSS.n2708 0.00978125
R5179 VSS.n3053 VSS.n3052 0.00978125
R5180 VSS.n3178 VSS.n3175 0.00978125
R5181 VSS.n2526 VSS.n2523 0.0095
R5182 VSS.n4057 VSS.n4050 0.0095
R5183 VSS.n110 VSS.n109 0.0095
R5184 VSS.n73 VSS.n71 0.0095
R5185 VSS.n3996 VSS.n3993 0.0095
R5186 VSS.n3167 VSS.n3164 0.00921875
R5187 VSS.n2809 VSS.n2807 0.0089375
R5188 VSS.n3677 VSS.n3675 0.008375
R5189 VSS.n2511 VSS.n2508 0.008375
R5190 VSS.n3641 VSS.n3637 0.008375
R5191 VSS.n3602 VSS.n3600 0.008375
R5192 VSS.n2156 VSS.n2088 0.008375
R5193 VSS.n2655 VSS.n2654 0.00809375
R5194 VSS.n3094 VSS.n3093 0.00809375
R5195 VSS.n3171 VSS.n3170 0.00809375
R5196 VSS.n133 VSS.n126 0.0078125
R5197 VSS.n2804 VSS.n2803 0.0078125
R5198 VSS.n2124 VSS.n2123 0.0078125
R5199 VSS.n119 VSS.n118 0.00725
R5200 VSS.n2056 VSS.n2055 0.00725
R5201 VSS.n133 VSS.n132 0.00725
R5202 VSS.n4064 VSS.n4061 0.00725
R5203 VSS.n115 VSS.n113 0.00725
R5204 VSS.n65 VSS.n64 0.00725
R5205 VSS.n3989 VSS.n3988 0.00725
R5206 VSS.n4041 VSS.n4040 0.006125
R5207 VSS.n103 VSS.n102 0.006125
R5208 VSS.n80 VSS.n78 0.006125
R5209 VSS.n4007 VSS.n4004 0.00579412
R5210 VSS.n2369 VSS.n2366 0.0055625
R5211 VSS.n2097 VSS.n2095 0.0055625
R5212 VSS.n2153 VSS.n2152 0.0055625
R5213 VSS.n3379 VSS.n3378 0.0055625
R5214 VSS.n2642 VSS.n2640 0.00528125
R5215 VSS.n3075 VSS.n3072 0.00528125
R5216 VSS.n1695 VSS.n1693 0.005
R5217 VSS.n1729 VSS.n1728 0.005
R5218 VSS.n1771 VSS.n1769 0.005
R5219 VSS.n1805 VSS.n1804 0.005
R5220 VSS.n1847 VSS.n1845 0.005
R5221 VSS.n1881 VSS.n1880 0.005
R5222 VSS.n877 VSS.n874 0.005
R5223 VSS.n926 VSS.n925 0.005
R5224 VSS.n1038 VSS.n1035 0.005
R5225 VSS.n1087 VSS.n1086 0.005
R5226 VSS.n1199 VSS.n1196 0.005
R5227 VSS.n1248 VSS.n1247 0.005
R5228 VSS.n3530 VSS.n3529 0.005
R5229 VSS.n1690 VSS.n1685 0.003875
R5230 VSS.n1734 VSS.n1732 0.003875
R5231 VSS.n1766 VSS.n1765 0.003875
R5232 VSS.n1810 VSS.n1808 0.003875
R5233 VSS.n1842 VSS.n1841 0.003875
R5234 VSS.n1886 VSS.n1884 0.003875
R5235 VSS.n870 VSS.n869 0.003875
R5236 VSS.n933 VSS.n930 0.003875
R5237 VSS.n1031 VSS.n1030 0.003875
R5238 VSS.n1094 VSS.n1091 0.003875
R5239 VSS.n1192 VSS.n1191 0.003875
R5240 VSS.n1255 VSS.n1252 0.003875
R5241 VSS.n3319 VSS.n3318 0.003875
R5242 VSS.n2620 VSS.n2619 0.00359375
R5243 VSS.n2672 VSS.n2671 0.00359375
R5244 VSS.n2717 VSS.n2715 0.00359375
R5245 VSS.n3043 VSS.n3042 0.00359375
R5246 VSS.n3119 VSS.n3118 0.00359375
R5247 VSS.n3188 VSS.n3185 0.00359375
R5248 VSS.n2021 VSS.n1289 0.0033125
R5249 VSS.n1702 VSS.n1700 0.0033125
R5250 VSS.n1798 VSS.n1797 0.0033125
R5251 VSS.n1854 VSS.n1852 0.0033125
R5252 VSS.n2822 VSS.n2820 0.0033125
R5253 VSS.n3764 VSS.n3751 0.00275
R5254 VSS.n3267 VSS.n3258 0.00275
R5255 VSS.n3160 VSS.n3159 0.00190625
R5256 VSS.n3580 VSS.n3578 0.0010625
R5257 VDD.t1254 VDD.t1366 147.304
R5258 VDD.t1178 VDD.t1254 147.304
R5259 VDD.t1274 VDD.t1178 147.304
R5260 VDD.t1208 VDD.t1274 147.304
R5261 VDD.t1193 VDD.t1304 147.304
R5262 VDD.t1374 VDD.t1193 147.304
R5263 VDD.t1281 VDD.t1374 147.304
R5264 VDD.t1155 VDD.t1281 147.304
R5265 VDD.t1328 VDD.t1198 135.05
R5266 VDD.t1168 VDD.t1328 135.05
R5267 VDD.t1260 VDD.t1308 135.05
R5268 VDD.t1293 VDD.t1260 135.05
R5269 VDD.t1381 VDD.t1263 135.05
R5270 VDD.t1227 VDD.t1381 135.05
R5271 VDD.t1196 VDD.t1171 135.05
R5272 VDD.t1147 VDD.t1196 135.05
R5273 VDD.t1348 VDD.t1234 118.626
R5274 VDD.t1205 VDD.t1354 118.626
R5275 VDD.n7371 VDD.t1211 103.504
R5276 VDD.n549 VDD.t1168 74.5648
R5277 VDD.n781 VDD.t1293 74.5648
R5278 VDD.n789 VDD.t1227 74.5648
R5279 VDD.n6805 VDD.t1147 74.5648
R5280 VDD.n289 VDD.t1208 72.6094
R5281 VDD.n289 VDD.t1391 72.6094
R5282 VDD.n6881 VDD.t1155 72.6094
R5283 VDD.n6881 VDD.t1267 72.6094
R5284 VDD.n2675 VDD.t1176 68.0469
R5285 VDD.n2838 VDD.t1141 68.0469
R5286 VDD.n2838 VDD.t1239 68.0469
R5287 VDD.n2675 VDD.t1330 68.0469
R5288 VDD.n3317 VDD.t1387 68.0469
R5289 VDD.n3317 VDD.t1232 68.0469
R5290 VDD.n5428 VDD.t1190 68.0469
R5291 VDD.n5428 VDD.t1244 68.0469
R5292 VDD.n3267 VDD.t1288 68.0469
R5293 VDD.n5369 VDD.t1312 68.0469
R5294 VDD.n5369 VDD.t1342 68.0469
R5295 VDD.n3267 VDD.t1187 68.0469
R5296 VDD.n3733 VDD.t1200 68.0469
R5297 VDD.n4577 VDD.t1217 68.0469
R5298 VDD.n4577 VDD.t1258 68.0469
R5299 VDD.n3733 VDD.t1316 68.0469
R5300 VDD.n3938 VDD.t1379 68.0469
R5301 VDD.n4067 VDD.t1393 68.0469
R5302 VDD.n4067 VDD.t1181 68.0469
R5303 VDD.n3938 VDD.t1332 68.0469
R5304 VDD.n2958 VDD.t1297 68.0469
R5305 VDD.n2958 VDD.t1320 68.0469
R5306 VDD.n4126 VDD.t1350 68.0469
R5307 VDD.n4126 VDD.t1246 68.0469
R5308 VDD.n2978 VDD.t1256 68.0469
R5309 VDD.n2978 VDD.t1310 68.0469
R5310 VDD.n4386 VDD.t1306 68.0469
R5311 VDD.n4386 VDD.t1236 68.0469
R5312 VDD.n3028 VDD.t1352 68.0469
R5313 VDD.n3028 VDD.t1362 68.0469
R5314 VDD.n4446 VDD.t1144 68.0469
R5315 VDD.n4446 VDD.t1161 68.0469
R5316 VDD.n3088 VDD.t1165 68.0469
R5317 VDD.n3088 VDD.t1286 68.0469
R5318 VDD.n4636 VDD.t1221 68.0469
R5319 VDD.n4636 VDD.t1265 68.0469
R5320 VDD.n3114 VDD.t1318 68.0469
R5321 VDD.n3114 VDD.t1290 68.0469
R5322 VDD.n4890 VDD.t1372 68.0469
R5323 VDD.n4890 VDD.t1322 68.0469
R5324 VDD.n3164 VDD.t1225 68.0469
R5325 VDD.n3164 VDD.t1324 68.0469
R5326 VDD.n4950 VDD.t1295 68.0469
R5327 VDD.n4950 VDD.t1184 68.0469
R5328 VDD.n3233 VDD.t1241 68.0469
R5329 VDD.n5137 VDD.t1344 68.0469
R5330 VDD.n5137 VDD.t1299 68.0469
R5331 VDD.n3233 VDD.t1272 68.0469
R5332 VDD.n3183 VDD.t1326 68.0469
R5333 VDD.n5077 VDD.t1249 68.0469
R5334 VDD.n5077 VDD.t1385 68.0469
R5335 VDD.n3183 VDD.t1276 68.0469
R5336 VDD.n2588 VDD.t1283 68.0469
R5337 VDD.n2588 VDD.t1383 68.0469
R5338 VDD.n2897 VDD.t1340 68.0469
R5339 VDD.n2897 VDD.t1336 68.0469
R5340 VDD.n387 VDD.t1205 63.8344
R5341 VDD.n398 VDD.t1214 63.8344
R5342 VDD.n7316 VDD.t1376 62.6612
R5343 VDD.n7369 VDD.t1150 62.6612
R5344 VDD.n302 VDD.t1301 62.4005
R5345 VDD.n299 VDD.t1158 62.4005
R5346 VDD.n7371 VDD.t1348 58.6612
R5347 VDD.n549 VDD.t1370 58.4005
R5348 VDD.n781 VDD.t1346 58.4005
R5349 VDD.n789 VDD.t1395 58.4005
R5350 VDD.n6805 VDD.t1219 58.4005
R5351 VDD.t1163 VDD.t1230 49.6666
R5352 VDD.t1314 VDD.t1163 49.6666
R5353 VDD.t1389 VDD.t1203 49.6666
R5354 VDD.t1173 VDD.t1389 49.6666
R5355 VDD.n1455 VDD.t1356 46.9291
R5356 VDD.n1133 VDD.t1269 46.9291
R5357 VDD.n1133 VDD.t1334 46.9291
R5358 VDD.n1455 VDD.t1338 46.9291
R5359 VDD.n1447 VDD.t1252 46.9291
R5360 VDD.n1447 VDD.t1223 46.9291
R5361 VDD.n1353 VDD.t1368 46.9291
R5362 VDD.n1107 VDD.t1278 46.9291
R5363 VDD.n1107 VDD.t1358 46.9291
R5364 VDD.n1353 VDD.t1360 46.9291
R5365 VDD.n6 VDD.t1314 24.8335
R5366 VDD.n6 VDD.t1152 24.8335
R5367 VDD.n7292 VDD.t1173 24.8335
R5368 VDD.n7292 VDD.t1364 24.8335
R5369 VDD.n370 VDD.t730 13.6237
R5370 VDD.n124 VDD.t1194 12.939
R5371 VDD.n186 VDD.t1179 12.939
R5372 VDD.t885 VDD.t581 12.7541
R5373 VDD.n7041 VDD.n7040 12.7307
R5374 VDD.n7708 VDD.t114 12.7307
R5375 VDD.n347 VDD.t212 12.4643
R5376 VDD.n7348 VDD.t792 12.4643
R5377 VDD.n137 VDD.t519 12.3639
R5378 VDD.n170 VDD.t361 12.3639
R5379 VDD.n7008 VDD.t1156 12.189
R5380 VDD.n7070 VDD.t1209 12.189
R5381 VDD.n367 VDD.t623 11.8846
R5382 VDD.n7021 VDD.t230 11.6473
R5383 VDD.n7056 VDD.t418 11.6473
R5384 VDD.n7338 VDD.t695 11.3048
R5385 VDD.n354 VDD.t790 10.7251
R5386 VDD.n351 VDD.t351 10.7251
R5387 VDD.n7258 VDD.t134 10.5639
R5388 VDD.n7554 VDD.t267 10.0222
R5389 VDD.n6863 VDD.t1148 9.91676
R5390 VDD.n1019 VDD.t1228 9.91676
R5391 VDD.n7329 VDD.t749 9.56572
R5392 VDD.n7332 VDD.t783 9.56572
R5393 VDD.n152 VDD.t107 9.48871
R5394 VDD.n155 VDD.t108 9.48871
R5395 VDD.n6850 VDD.t290 9.47604
R5396 VDD.n1007 VDD.t282 9.47604
R5397 VDD.n2488 VDD.t412 9.23695
R5398 VDD.n7037 VDD.t537 8.93874
R5399 VDD.n7041 VDD.t294 8.93874
R5400 VDD.n2118 VDD.t116 8.82644
R5401 VDD.n2429 VDD.t167 8.82644
R5402 VDD.n1062 VDD.t304 8.59459
R5403 VDD.n1083 VDD.t104 8.59459
R5404 VDD.n5608 VDD.t435 8.54751
R5405 VDD.n5628 VDD.t43 8.54751
R5406 VDD.n6079 VDD.t161 8.54751
R5407 VDD.n6099 VDD.t295 8.54751
R5408 VDD.n6226 VDD.t254 8.54751
R5409 VDD.n6246 VDD.t98 8.54751
R5410 VDD.n6381 VDD.t17 8.54751
R5411 VDD.n6401 VDD.t236 8.54751
R5412 VDD.n6540 VDD.t263 8.54751
R5413 VDD.n6560 VDD.t88 8.54751
R5414 VDD.n5777 VDD.t19 8.54751
R5415 VDD.n5797 VDD.t152 8.54751
R5416 VDD.n5924 VDD.t551 8.54751
R5417 VDD.n5944 VDD.t311 8.54751
R5418 VDD.n2109 VDD.t165 8.41594
R5419 VDD.n2449 VDD.t109 8.41594
R5420 VDD.n315 VDD.t1206 8.4063
R5421 VDD.n344 VDD.t753 8.4063
R5422 VDD.n7526 VDD.t1212 8.4063
R5423 VDD.n7288 VDD.n7287 8.2255
R5424 VDD.n7724 VDD.n7288 8.2255
R5425 VDD.n2100 VDD.t511 8.00543
R5426 VDD.n2210 VDD.t229 8.00543
R5427 VDD.n7279 VDD.t520 7.85532
R5428 VDD.n2091 VDD.t697 7.59492
R5429 VDD.n2219 VDD.t13 7.59492
R5430 VDD.n2303 VDD.t405 7.59492
R5431 VDD.n7267 VDD.t329 7.31361
R5432 VDD.n6833 VDD.t209 7.27243
R5433 VDD.n990 VDD.t105 7.27243
R5434 VDD.n1071 VDD.t309 7.27243
R5435 VDD.n1074 VDD.t103 7.27243
R5436 VDD.n370 VDD.t793 7.24688
R5437 VDD.n2183 VDD.t14 7.18441
R5438 VDD.n2291 VDD.t415 7.18441
R5439 VDD.n2471 VDD.t207 7.18441
R5440 VDD.n1464 VDD.t11 7.0395
R5441 VDD.n1463 VDD.t935 7.0395
R5442 VDD.n1936 VDD.t1072 7.0395
R5443 VDD.n1937 VDD.t420 7.0395
R5444 VDD.n5588 VDD.t86 6.91951
R5445 VDD.n5648 VDD.t179 6.91951
R5446 VDD.n6059 VDD.t567 6.91951
R5447 VDD.n6119 VDD.t158 6.91951
R5448 VDD.n6206 VDD.t52 6.91951
R5449 VDD.n6266 VDD.t508 6.91951
R5450 VDD.n6361 VDD.t125 6.91951
R5451 VDD.n6421 VDD.t376 6.91951
R5452 VDD.n6520 VDD.t645 6.91951
R5453 VDD.n6580 VDD.t445 6.91951
R5454 VDD.n5757 VDD.t492 6.91951
R5455 VDD.n5817 VDD.t577 6.91951
R5456 VDD.n5904 VDD.t5 6.91951
R5457 VDD.n5964 VDD.t127 6.91951
R5458 VDD.n2198 VDD.t573 6.7739
R5459 VDD.n2282 VDD.t35 6.7739
R5460 VDD.n2408 VDD.t320 6.7739
R5461 VDD.n2411 VDD.t574 6.7739
R5462 VDD.n344 VDD.t592 6.66717
R5463 VDD.n140 VDD.t293 6.6135
R5464 VDD.n167 VDD.t411 6.6135
R5465 VDD.n5592 VDD.t32 6.51251
R5466 VDD.n5644 VDD.t430 6.51251
R5467 VDD.n6063 VDD.t457 6.51251
R5468 VDD.n6115 VDD.t117 6.51251
R5469 VDD.n6210 VDD.t122 6.51251
R5470 VDD.n6262 VDD.t597 6.51251
R5471 VDD.n6365 VDD.t355 6.51251
R5472 VDD.n6417 VDD.t21 6.51251
R5473 VDD.n6524 VDD.t0 6.51251
R5474 VDD.n6576 VDD.t148 6.51251
R5475 VDD.n5761 VDD.t442 6.51251
R5476 VDD.n5813 VDD.t465 6.51251
R5477 VDD.n5908 VDD.t244 6.51251
R5478 VDD.n5960 VDD.t70 6.51251
R5479 VDD.n1803 VDD.t367 6.4095
R5480 VDD.n1802 VDD.t368 6.4095
R5481 VDD.n1801 VDD.t15 6.4095
R5482 VDD.n1552 VDD.t16 6.4095
R5483 VDD.n1464 VDD.t12 6.4095
R5484 VDD.n1463 VDD.t936 6.4095
R5485 VDD.n1800 VDD.t397 6.4095
R5486 VDD.n1799 VDD.t398 6.4095
R5487 VDD.n1798 VDD.t399 6.4095
R5488 VDD.n1462 VDD.t400 6.4095
R5489 VDD.n1936 VDD.t1071 6.4095
R5490 VDD.n1937 VDD.t419 6.4095
R5491 VDD.n2467 VDD.t401 6.36339
R5492 VDD VDD.n7288 6.3005
R5493 VDD VDD.n7288 6.3005
R5494 VDD.n389 VDD.t1355 6.2405
R5495 VDD.n7380 VDD.t1235 6.2405
R5496 VDD.n7025 VDD.t292 6.23019
R5497 VDD.n7053 VDD.t620 6.23019
R5498 VDD.n2130 VDD.t934 5.95288
R5499 VDD.t746 VDD.t323 5.7976
R5500 VDD.n315 VDD.t1302 5.50775
R5501 VDD.n383 VDD.t970 5.50775
R5502 VDD.n367 VDD.t1397 5.50775
R5503 VDD.n363 VDD.t788 5.50775
R5504 VDD.n7329 VDD.t750 5.50775
R5505 VDD.n7714 VDD.t137 5.14676
R5506 VDD.n7698 VDD.t1174 5.14676
R5507 VDD.n2454 VDD.t204 5.13186
R5508 VDD.n6846 VDD.t761 5.06881
R5509 VDD.n1003 VDD.t759 5.06881
R5510 VDD.n1037 VDD.t1261 5.06881
R5511 VDD.n561 VDD.t1169 5.06881
R5512 VDD.n5605 VDD.t669 4.88451
R5513 VDD.n5631 VDD.t780 4.88451
R5514 VDD.n6076 VDD.t67 4.88451
R5515 VDD.n6102 VDD.t587 4.88451
R5516 VDD.n6223 VDD.t46 4.88451
R5517 VDD.n6249 VDD.t163 4.88451
R5518 VDD.n6378 VDD.t155 4.88451
R5519 VDD.n6404 VDD.t358 4.88451
R5520 VDD.n6537 VDD.t812 4.88451
R5521 VDD.n6563 VDD.t437 4.88451
R5522 VDD.n5774 VDD.t469 4.88451
R5523 VDD.n5800 VDD.t379 4.88451
R5524 VDD.n5921 VDD.t57 4.88451
R5525 VDD.n5947 VDD.t3 4.88451
R5526 VDD.n2394 VDD.t1013 4.72135
R5527 VDD.n2425 VDD.t531 4.72135
R5528 VDD.n1444 VDD.n1443 4.64717
R5529 VDD.n5575 VDD.t252 4.4775
R5530 VDD.n5661 VDD.t483 4.4775
R5531 VDD.n6046 VDD.t374 4.4775
R5532 VDD.n6132 VDD.t216 4.4775
R5533 VDD.n6193 VDD.t214 4.4775
R5534 VDD.n6279 VDD.t494 4.4775
R5535 VDD.n6348 VDD.t433 4.4775
R5536 VDD.n6434 VDD.t666 4.4775
R5537 VDD.n6507 VDD.t275 4.4775
R5538 VDD.n6593 VDD.t317 4.4775
R5539 VDD.n5744 VDD.t385 4.4775
R5540 VDD.n5830 VDD.t60 4.4775
R5541 VDD.n5891 VDD.t50 4.4775
R5542 VDD.n5977 VDD.t38 4.4775
R5543 VDD.n322 VDD.t540 4.34833
R5544 VDD.n326 VDD.t1215 4.34833
R5545 VDD.n332 VDD.t746 4.34833
R5546 VDD.n354 VDD.t1095 4.34833
R5547 VDD.n7355 VDD.t1101 4.34833
R5548 VDD.n7366 VDD.n7365 4.31441
R5549 VDD.n2484 VDD.t364 4.31084
R5550 VDD.n396 VDD.n395 4.09528
R5551 VDD.n7082 VDD.n7079 4.09137
R5552 VDD.n7542 VDD.n7539 4.09137
R5553 VDD.n7309 VDD.n7306 4.09137
R5554 VDD.n1370 VDD.n1369 4.0405
R5555 VDD.n1381 VDD.n1380 4.0405
R5556 VDD.n1392 VDD.n1391 4.0405
R5557 VDD.n1403 VDD.n1402 4.0405
R5558 VDD.n1414 VDD.n1413 4.0405
R5559 VDD.n1425 VDD.n1424 4.0405
R5560 VDD.n791 VDD.t1396 4.02914
R5561 VDD.n6882 VDD.n6881 4.0005
R5562 VDD.n290 VDD.n289 4.0005
R5563 VDD.n7293 VDD.n7292 4.0005
R5564 VDD.n7372 VDD.n7371 4.0005
R5565 VDD.n782 VDD.n781 4.0005
R5566 VDD.n790 VDD.n789 4.0005
R5567 VDD.n6806 VDD.n6805 4.0005
R5568 VDD.n550 VDD.n549 4.0005
R5569 VDD.n3268 VDD.n3267 4.0005
R5570 VDD.n5370 VDD.n5369 4.0005
R5571 VDD.n4127 VDD.n4126 4.0005
R5572 VDD.n2959 VDD.n2958 4.0005
R5573 VDD.n4387 VDD.n4386 4.0005
R5574 VDD.n2979 VDD.n2978 4.0005
R5575 VDD.n4447 VDD.n4446 4.0005
R5576 VDD.n3029 VDD.n3028 4.0005
R5577 VDD.n3939 VDD.n3938 4.0005
R5578 VDD.n4068 VDD.n4067 4.0005
R5579 VDD.n4637 VDD.n4636 4.0005
R5580 VDD.n3089 VDD.n3088 4.0005
R5581 VDD.n4891 VDD.n4890 4.0005
R5582 VDD.n3115 VDD.n3114 4.0005
R5583 VDD.n4951 VDD.n4950 4.0005
R5584 VDD.n3165 VDD.n3164 4.0005
R5585 VDD.n3734 VDD.n3733 4.0005
R5586 VDD.n4578 VDD.n4577 4.0005
R5587 VDD.n3234 VDD.n3233 4.0005
R5588 VDD.n5138 VDD.n5137 4.0005
R5589 VDD.n3184 VDD.n3183 4.0005
R5590 VDD.n5078 VDD.n5077 4.0005
R5591 VDD.n5429 VDD.n5428 4.0005
R5592 VDD.n3318 VDD.n3317 4.0005
R5593 VDD.n2898 VDD.n2897 4.0005
R5594 VDD.n2589 VDD.n2588 4.0005
R5595 VDD.n2676 VDD.n2675 4.0005
R5596 VDD.n2839 VDD.n2838 4.0005
R5597 VDD.n1456 VDD.n1455 4.0005
R5598 VDD.n1134 VDD.n1133 4.0005
R5599 VDD.n1448 VDD.n1447 4.0005
R5600 VDD.n1354 VDD.n1353 4.0005
R5601 VDD.n1108 VDD.n1107 4.0005
R5602 VDD.n7 VDD.n6 4.0005
R5603 VDD.n399 VDD.t1216 3.9242
R5604 VDD.n7317 VDD.t1378 3.90659
R5605 VDD.n7370 VDD.t1151 3.90659
R5606 VDD.n3292 VDD.n3291 3.89963
R5607 VDD.n5392 VDD.n5391 3.89963
R5608 VDD.n5401 VDD.n5400 3.89963
R5609 VDD.n4100 VDD.n4099 3.89963
R5610 VDD.n4105 VDD.n4104 3.89963
R5611 VDD.n2942 VDD.n2941 3.89963
R5612 VDD.n4410 VDD.n4409 3.89963
R5613 VDD.n4415 VDD.n4414 3.89963
R5614 VDD.n3006 VDD.n3005 3.89963
R5615 VDD.n4610 VDD.n4609 3.89963
R5616 VDD.n4615 VDD.n4614 3.89963
R5617 VDD.n3072 VDD.n3071 3.89963
R5618 VDD.n4914 VDD.n4913 3.89963
R5619 VDD.n4919 VDD.n4918 3.89963
R5620 VDD.n3142 VDD.n3141 3.89963
R5621 VDD.n3214 VDD.n3213 3.89963
R5622 VDD.n5110 VDD.n5109 3.89963
R5623 VDD.n5119 VDD.n5118 3.89963
R5624 VDD.n2861 VDD.n2860 3.89963
R5625 VDD.n2866 VDD.n2865 3.89963
R5626 VDD.n2566 VDD.n2565 3.89963
R5627 VDD.n1449 VDD.t1224 3.88217
R5628 VDD.n7341 VDD.n7319 3.88202
R5629 VDD.n7328 VDD.n7321 3.88202
R5630 VDD.n350 VDD.n340 3.88202
R5631 VDD.n366 VDD.n338 3.88202
R5632 VDD.n379 VDD.n336 3.88202
R5633 VDD.n6546 VDD.n2878 3.83311
R5634 VDD.n6556 VDD.n2876 3.83311
R5635 VDD.n5614 VDD.n5409 3.83311
R5636 VDD.n5624 VDD.n5407 3.83311
R5637 VDD.n5930 VDD.n4931 3.83311
R5638 VDD.n5940 VDD.n4929 3.83311
R5639 VDD.n6085 VDD.n4605 3.83311
R5640 VDD.n6095 VDD.n4603 3.83311
R5641 VDD.n6232 VDD.n4427 3.83311
R5642 VDD.n6242 VDD.n4425 3.83311
R5643 VDD.n6387 VDD.n4095 3.83311
R5644 VDD.n6397 VDD.n4093 3.83311
R5645 VDD.n5783 VDD.n5105 3.83311
R5646 VDD.n5793 VDD.n5103 3.83311
R5647 VDD.n1047 VDD.t305 3.74664
R5648 VDD.n1098 VDD.t310 3.74664
R5649 VDD.n403 VDD.n402 3.6405
R5650 VDD.n2383 VDD.t843 3.48983
R5651 VDD.n2495 VDD.t130 3.48983
R5652 VDD.t970 VDD.t740 3.47876
R5653 VDD.n396 VDD.n393 3.4692
R5654 VDD.n397 VDD.n391 3.4692
R5655 VDD.n7366 VDD.n7363 3.4692
R5656 VDD.n7367 VDD.n7361 3.4692
R5657 VDD.n303 VDD.n301 3.44767
R5658 VDD.n300 VDD.n298 3.44767
R5659 VDD.n1131 VDD.n1130 3.3285
R5660 VDD.n1129 VDD.n1128 3.3285
R5661 VDD.n3292 VDD.n3289 3.27354
R5662 VDD.n5392 VDD.n5389 3.27354
R5663 VDD.n5401 VDD.n5398 3.27354
R5664 VDD.n4100 VDD.n4097 3.27354
R5665 VDD.n4105 VDD.n4102 3.27354
R5666 VDD.n2942 VDD.n2939 3.27354
R5667 VDD.n4410 VDD.n4407 3.27354
R5668 VDD.n4415 VDD.n4412 3.27354
R5669 VDD.n3006 VDD.n3003 3.27354
R5670 VDD.n4610 VDD.n4607 3.27354
R5671 VDD.n4615 VDD.n4612 3.27354
R5672 VDD.n3072 VDD.n3069 3.27354
R5673 VDD.n4914 VDD.n4911 3.27354
R5674 VDD.n4919 VDD.n4916 3.27354
R5675 VDD.n3142 VDD.n3139 3.27354
R5676 VDD.n3214 VDD.n3211 3.27354
R5677 VDD.n5110 VDD.n5107 3.27354
R5678 VDD.n5119 VDD.n5116 3.27354
R5679 VDD.n2861 VDD.n2858 3.27354
R5680 VDD.n2866 VDD.n2863 3.27354
R5681 VDD.n2566 VDD.n2563 3.27354
R5682 VDD.n5565 VDD.t1191 3.2565
R5683 VDD.n5671 VDD.t1188 3.2565
R5684 VDD.n6036 VDD.t1166 3.2565
R5685 VDD.n6142 VDD.t1201 3.2565
R5686 VDD.n6183 VDD.t1145 3.2565
R5687 VDD.n6289 VDD.t1237 3.2565
R5688 VDD.n6338 VDD.t1247 3.2565
R5689 VDD.n6444 VDD.t1182 3.2565
R5690 VDD.n6497 VDD.t1284 3.2565
R5691 VDD.n6603 VDD.t1142 3.2565
R5692 VDD.n5734 VDD.t1242 3.2565
R5693 VDD.n5840 VDD.t1250 3.2565
R5694 VDD.n5881 VDD.t1185 3.2565
R5695 VDD.n5987 VDD.t1291 3.2565
R5696 VDD.n2841 VDD.t1143 3.20717
R5697 VDD.n2837 VDD.t1240 3.20717
R5698 VDD.n2674 VDD.t1331 3.20717
R5699 VDD.n2678 VDD.t1177 3.20717
R5700 VDD.n5430 VDD.t1192 3.20717
R5701 VDD.n3316 VDD.t1233 3.20717
R5702 VDD.n5432 VDD.t1245 3.20717
R5703 VDD.n5372 VDD.t1313 3.20717
R5704 VDD.n5368 VDD.t1343 3.20717
R5705 VDD.n3266 VDD.t1189 3.20717
R5706 VDD.n3270 VDD.t1289 3.20717
R5707 VDD.n4580 VDD.t1218 3.20717
R5708 VDD.n4576 VDD.t1259 3.20717
R5709 VDD.n3732 VDD.t1317 3.20717
R5710 VDD.n3736 VDD.t1202 3.20717
R5711 VDD.n4070 VDD.t1394 3.20717
R5712 VDD.n4066 VDD.t1183 3.20717
R5713 VDD.n3937 VDD.t1333 3.20717
R5714 VDD.n3941 VDD.t1380 3.20717
R5715 VDD.n4128 VDD.t1351 3.20717
R5716 VDD.n2957 VDD.t1321 3.20717
R5717 VDD.n4130 VDD.t1248 3.20717
R5718 VDD.n2961 VDD.t1298 3.20717
R5719 VDD.n4388 VDD.t1307 3.20717
R5720 VDD.n2977 VDD.t1311 3.20717
R5721 VDD.n4390 VDD.t1238 3.20717
R5722 VDD.n2981 VDD.t1257 3.20717
R5723 VDD.n4448 VDD.t1146 3.20717
R5724 VDD.n3027 VDD.t1363 3.20717
R5725 VDD.n4450 VDD.t1162 3.20717
R5726 VDD.n3031 VDD.t1353 3.20717
R5727 VDD.n4638 VDD.t1222 3.20717
R5728 VDD.n3087 VDD.t1287 3.20717
R5729 VDD.n4640 VDD.t1266 3.20717
R5730 VDD.n3091 VDD.t1167 3.20717
R5731 VDD.n4892 VDD.t1373 3.20717
R5732 VDD.n3113 VDD.t1292 3.20717
R5733 VDD.n4894 VDD.t1323 3.20717
R5734 VDD.n3117 VDD.t1319 3.20717
R5735 VDD.n4952 VDD.t1296 3.20717
R5736 VDD.n3163 VDD.t1325 3.20717
R5737 VDD.n4954 VDD.t1186 3.20717
R5738 VDD.n3167 VDD.t1226 3.20717
R5739 VDD.n5140 VDD.t1345 3.20717
R5740 VDD.n5136 VDD.t1300 3.20717
R5741 VDD.n3232 VDD.t1273 3.20717
R5742 VDD.n3236 VDD.t1243 3.20717
R5743 VDD.n5080 VDD.t1251 3.20717
R5744 VDD.n5076 VDD.t1386 3.20717
R5745 VDD.n3182 VDD.t1277 3.20717
R5746 VDD.n3186 VDD.t1327 3.20717
R5747 VDD.n3320 VDD.t1388 3.20717
R5748 VDD.n2899 VDD.t1341 3.20717
R5749 VDD.n2587 VDD.t1384 3.20717
R5750 VDD.n2901 VDD.t1337 3.20717
R5751 VDD.n2591 VDD.t1285 3.20717
R5752 VDD.n1446 VDD.n1440 3.20717
R5753 VDD.n1445 VDD.n1441 3.20717
R5754 VDD.n1444 VDD.n1442 3.20717
R5755 VDD.n1136 VDD.t1271 3.20717
R5756 VDD.n1454 VDD.t1339 3.20717
R5757 VDD.n1132 VDD.t1335 3.20717
R5758 VDD.n1458 VDD.t1357 3.20717
R5759 VDD.n1450 VDD.t1253 3.20717
R5760 VDD.n1110 VDD.t1280 3.20717
R5761 VDD.n1352 VDD.t1361 3.20717
R5762 VDD.n1106 VDD.t1359 3.20717
R5763 VDD.n1356 VDD.t1369 3.20717
R5764 VDD.n3849 VDD.n3848 3.1914
R5765 VDD.n3644 VDD.n3643 3.1914
R5766 VDD.n3443 VDD.n3442 3.1914
R5767 VDD.n1467 VDD.n1465 3.1914
R5768 VDD.n3338 VDD.n3337 3.19093
R5769 VDD.n2349 VDD.n2348 3.19093
R5770 VDD.n2158 VDD.n2157 3.19093
R5771 VDD.n2055 VDD.n2054 3.19093
R5772 VDD.n3439 VDD.n3438 3.1908
R5773 VDD.n5708 VDD.n5707 3.1908
R5774 VDD.n2540 VDD.n2539 3.1908
R5775 VDD.n1249 VDD.n1248 3.1908
R5776 VDD.n7345 VDD.t772 3.18891
R5777 VDD.n7077 VDD.t1154 3.18197
R5778 VDD.n7302 VDD.t1365 3.18197
R5779 VDD.n552 VDD.t1371 3.18197
R5780 VDD.n548 VDD.t1170 3.18197
R5781 VDD.n547 VDD.t1329 3.18197
R5782 VDD.n571 VDD.t1199 3.18197
R5783 VDD.n784 VDD.t1347 3.18197
R5784 VDD.n780 VDD.t1294 3.18197
R5785 VDD.n779 VDD.t1262 3.18197
R5786 VDD.n572 VDD.t1309 3.18197
R5787 VDD.n792 VDD.t1229 3.18197
R5788 VDD.n793 VDD.t1382 3.18197
R5789 VDD.n794 VDD.t1264 3.18197
R5790 VDD.n6649 VDD.t1172 3.18197
R5791 VDD.n6807 VDD.t1197 3.18197
R5792 VDD.n6808 VDD.t1149 3.18197
R5793 VDD.n6810 VDD.t1220 3.18197
R5794 VDD.n7126 VDD.n7125 3.1505
R5795 VDD.n7590 VDD.n7589 3.1505
R5796 VDD.n7130 VDD.n7129 3.1505
R5797 VDD.n7132 VDD.n7131 3.1505
R5798 VDD.n7134 VDD.n7133 3.1505
R5799 VDD.n7136 VDD.n7135 3.1505
R5800 VDD.n7138 VDD.n7137 3.1505
R5801 VDD.n7140 VDD.n7139 3.1505
R5802 VDD.n7142 VDD.n7141 3.1505
R5803 VDD.n7144 VDD.n7143 3.1505
R5804 VDD.n7146 VDD.n7145 3.1505
R5805 VDD.n7148 VDD.n7147 3.1505
R5806 VDD.n7151 VDD.n7150 3.1505
R5807 VDD.n7154 VDD.n7153 3.1505
R5808 VDD.n7157 VDD.n7156 3.1505
R5809 VDD.n7160 VDD.n7159 3.1505
R5810 VDD.n7163 VDD.n7162 3.1505
R5811 VDD.n7166 VDD.n7165 3.1505
R5812 VDD.n7169 VDD.n7168 3.1505
R5813 VDD.n7172 VDD.n7171 3.1505
R5814 VDD.n7175 VDD.n7174 3.1505
R5815 VDD.n7178 VDD.n7177 3.1505
R5816 VDD.n7181 VDD.n7180 3.1505
R5817 VDD.n7184 VDD.n7183 3.1505
R5818 VDD.n7187 VDD.n7186 3.1505
R5819 VDD.n7190 VDD.n7189 3.1505
R5820 VDD.n7193 VDD.n7192 3.1505
R5821 VDD.n7196 VDD.n7195 3.1505
R5822 VDD.n7199 VDD.n7198 3.1505
R5823 VDD.n7202 VDD.n7201 3.1505
R5824 VDD.n7205 VDD.n7204 3.1505
R5825 VDD.n7208 VDD.n7207 3.1505
R5826 VDD.n7211 VDD.n7210 3.1505
R5827 VDD.n7214 VDD.n7213 3.1505
R5828 VDD.n7217 VDD.n7216 3.1505
R5829 VDD.n7220 VDD.n7219 3.1505
R5830 VDD.n7223 VDD.n7222 3.1505
R5831 VDD.n7670 VDD.n7669 3.1505
R5832 VDD.n7668 VDD.n7667 3.1505
R5833 VDD.n7665 VDD.n7664 3.1505
R5834 VDD.n7663 VDD.n7662 3.1505
R5835 VDD.n7660 VDD.n7659 3.1505
R5836 VDD.n7658 VDD.n7657 3.1505
R5837 VDD.n7655 VDD.n7654 3.1505
R5838 VDD.n7653 VDD.n7652 3.1505
R5839 VDD.n7650 VDD.n7649 3.1505
R5840 VDD.n7648 VDD.n7647 3.1505
R5841 VDD.n7645 VDD.n7644 3.1505
R5842 VDD.n7643 VDD.n7642 3.1505
R5843 VDD.n7640 VDD.n7639 3.1505
R5844 VDD.n7638 VDD.n7637 3.1505
R5845 VDD.n7635 VDD.n7634 3.1505
R5846 VDD.n7633 VDD.n7632 3.1505
R5847 VDD.n7630 VDD.n7629 3.1505
R5848 VDD.n7628 VDD.n7627 3.1505
R5849 VDD.n7626 VDD.n7625 3.1505
R5850 VDD.n7624 VDD.n7623 3.1505
R5851 VDD.n7622 VDD.n7621 3.1505
R5852 VDD.n7620 VDD.n7619 3.1505
R5853 VDD.n7618 VDD.n7617 3.1505
R5854 VDD.n7616 VDD.n7615 3.1505
R5855 VDD.n7614 VDD.n7613 3.1505
R5856 VDD.n7612 VDD.n7611 3.1505
R5857 VDD.n7610 VDD.n7609 3.1505
R5858 VDD.n7608 VDD.n7607 3.1505
R5859 VDD.n7606 VDD.n7605 3.1505
R5860 VDD.n7604 VDD.n7603 3.1505
R5861 VDD.n7602 VDD.n7601 3.1505
R5862 VDD.n7600 VDD.n7599 3.1505
R5863 VDD.n7598 VDD.n7597 3.1505
R5864 VDD.n7596 VDD.n7595 3.1505
R5865 VDD.n7594 VDD.n7593 3.1505
R5866 VDD.n7592 VDD.n7591 3.1505
R5867 VDD.n7128 VDD.n7127 3.1505
R5868 VDD.n286 VDD.n285 3.1505
R5869 VDD.n199 VDD.n198 3.1505
R5870 VDD.n201 VDD.n200 3.1505
R5871 VDD.n203 VDD.n202 3.1505
R5872 VDD.n205 VDD.n204 3.1505
R5873 VDD.n207 VDD.n206 3.1505
R5874 VDD.n209 VDD.n208 3.1505
R5875 VDD.n211 VDD.n210 3.1505
R5876 VDD.n213 VDD.n212 3.1505
R5877 VDD.n215 VDD.n214 3.1505
R5878 VDD.n217 VDD.n216 3.1505
R5879 VDD.n219 VDD.n218 3.1505
R5880 VDD.n221 VDD.n220 3.1505
R5881 VDD.n223 VDD.n222 3.1505
R5882 VDD.n225 VDD.n224 3.1505
R5883 VDD.n227 VDD.n226 3.1505
R5884 VDD.n229 VDD.n228 3.1505
R5885 VDD.n232 VDD.n231 3.1505
R5886 VDD.n234 VDD.n233 3.1505
R5887 VDD.n237 VDD.n236 3.1505
R5888 VDD.n239 VDD.n238 3.1505
R5889 VDD.n242 VDD.n241 3.1505
R5890 VDD.n244 VDD.n243 3.1505
R5891 VDD.n247 VDD.n246 3.1505
R5892 VDD.n249 VDD.n248 3.1505
R5893 VDD.n252 VDD.n251 3.1505
R5894 VDD.n254 VDD.n253 3.1505
R5895 VDD.n257 VDD.n256 3.1505
R5896 VDD.n259 VDD.n258 3.1505
R5897 VDD.n262 VDD.n261 3.1505
R5898 VDD.n264 VDD.n263 3.1505
R5899 VDD.n267 VDD.n266 3.1505
R5900 VDD.n269 VDD.n268 3.1505
R5901 VDD.n272 VDD.n271 3.1505
R5902 VDD.n274 VDD.n273 3.1505
R5903 VDD.n197 VDD.n196 3.1505
R5904 VDD.n105 VDD.n104 3.1505
R5905 VDD.n7000 VDD.n6999 3.1505
R5906 VDD.n6986 VDD.n6985 3.1505
R5907 VDD.n6983 VDD.n6982 3.1505
R5908 VDD.n6980 VDD.n6979 3.1505
R5909 VDD.n6977 VDD.n6976 3.1505
R5910 VDD.n6974 VDD.n6973 3.1505
R5911 VDD.n6971 VDD.n6970 3.1505
R5912 VDD.n6968 VDD.n6967 3.1505
R5913 VDD.n6965 VDD.n6964 3.1505
R5914 VDD.n6962 VDD.n6961 3.1505
R5915 VDD.n6959 VDD.n6958 3.1505
R5916 VDD.n6956 VDD.n6955 3.1505
R5917 VDD.n6953 VDD.n6952 3.1505
R5918 VDD.n6950 VDD.n6949 3.1505
R5919 VDD.n6947 VDD.n6946 3.1505
R5920 VDD.n6944 VDD.n6943 3.1505
R5921 VDD.n6941 VDD.n6940 3.1505
R5922 VDD.n6938 VDD.n6937 3.1505
R5923 VDD.n6935 VDD.n6934 3.1505
R5924 VDD.n6932 VDD.n6931 3.1505
R5925 VDD.n6929 VDD.n6928 3.1505
R5926 VDD.n6926 VDD.n6925 3.1505
R5927 VDD.n6923 VDD.n6922 3.1505
R5928 VDD.n6920 VDD.n6919 3.1505
R5929 VDD.n6917 VDD.n6916 3.1505
R5930 VDD.n6914 VDD.n6913 3.1505
R5931 VDD.n6911 VDD.n6910 3.1505
R5932 VDD.n6908 VDD.n6907 3.1505
R5933 VDD.n6906 VDD.n6905 3.1505
R5934 VDD.n6904 VDD.n6903 3.1505
R5935 VDD.n6902 VDD.n6901 3.1505
R5936 VDD.n6900 VDD.n6899 3.1505
R5937 VDD.n6898 VDD.n6897 3.1505
R5938 VDD.n6896 VDD.n6895 3.1505
R5939 VDD.n6894 VDD.n6893 3.1505
R5940 VDD.n6892 VDD.n6891 3.1505
R5941 VDD.n6890 VDD.n6889 3.1505
R5942 VDD.n26 VDD.n25 3.1505
R5943 VDD.n28 VDD.n27 3.1505
R5944 VDD.n30 VDD.n29 3.1505
R5945 VDD.n32 VDD.n31 3.1505
R5946 VDD.n34 VDD.n33 3.1505
R5947 VDD.n36 VDD.n35 3.1505
R5948 VDD.n38 VDD.n37 3.1505
R5949 VDD.n40 VDD.n39 3.1505
R5950 VDD.n42 VDD.n41 3.1505
R5951 VDD.n44 VDD.n43 3.1505
R5952 VDD.n46 VDD.n45 3.1505
R5953 VDD.n48 VDD.n47 3.1505
R5954 VDD.n50 VDD.n49 3.1505
R5955 VDD.n52 VDD.n51 3.1505
R5956 VDD.n54 VDD.n53 3.1505
R5957 VDD.n56 VDD.n55 3.1505
R5958 VDD.n58 VDD.n57 3.1505
R5959 VDD.n60 VDD.n59 3.1505
R5960 VDD.n62 VDD.n61 3.1505
R5961 VDD.n64 VDD.n63 3.1505
R5962 VDD.n66 VDD.n65 3.1505
R5963 VDD.n68 VDD.n67 3.1505
R5964 VDD.n71 VDD.n70 3.1505
R5965 VDD.n73 VDD.n72 3.1505
R5966 VDD.n76 VDD.n75 3.1505
R5967 VDD.n78 VDD.n77 3.1505
R5968 VDD.n81 VDD.n80 3.1505
R5969 VDD.n83 VDD.n82 3.1505
R5970 VDD.n86 VDD.n85 3.1505
R5971 VDD.n88 VDD.n87 3.1505
R5972 VDD.n91 VDD.n90 3.1505
R5973 VDD.n93 VDD.n92 3.1505
R5974 VDD.n96 VDD.n95 3.1505
R5975 VDD.n98 VDD.n97 3.1505
R5976 VDD.n101 VDD.n100 3.1505
R5977 VDD.n103 VDD.n102 3.1505
R5978 VDD.n119 VDD.n118 3.1505
R5979 VDD.n122 VDD.n121 3.1505
R5980 VDD.n121 VDD.n120 3.1505
R5981 VDD.n126 VDD.n125 3.1505
R5982 VDD.n125 VDD.n124 3.1505
R5983 VDD.n129 VDD.n128 3.1505
R5984 VDD.n128 VDD.n127 3.1505
R5985 VDD.n133 VDD.n132 3.1505
R5986 VDD.n132 VDD.n131 3.1505
R5987 VDD.n136 VDD.n135 3.1505
R5988 VDD.n135 VDD.n134 3.1505
R5989 VDD.n139 VDD.n138 3.1505
R5990 VDD.n138 VDD.n137 3.1505
R5991 VDD.n142 VDD.n141 3.1505
R5992 VDD.n141 VDD.n140 3.1505
R5993 VDD.n145 VDD.n144 3.1505
R5994 VDD.n144 VDD.n143 3.1505
R5995 VDD.n148 VDD.n147 3.1505
R5996 VDD.n147 VDD.n146 3.1505
R5997 VDD.n151 VDD.n150 3.1505
R5998 VDD.n150 VDD.n149 3.1505
R5999 VDD.n154 VDD.n153 3.1505
R6000 VDD.n153 VDD.n152 3.1505
R6001 VDD.n157 VDD.n156 3.1505
R6002 VDD.n156 VDD.n155 3.1505
R6003 VDD.n160 VDD.n159 3.1505
R6004 VDD.n159 VDD.n158 3.1505
R6005 VDD.n163 VDD.n162 3.1505
R6006 VDD.n162 VDD.n161 3.1505
R6007 VDD.n166 VDD.n165 3.1505
R6008 VDD.n165 VDD.n164 3.1505
R6009 VDD.n169 VDD.n168 3.1505
R6010 VDD.n168 VDD.n167 3.1505
R6011 VDD.n172 VDD.n171 3.1505
R6012 VDD.n171 VDD.n170 3.1505
R6013 VDD.n175 VDD.n174 3.1505
R6014 VDD.n174 VDD.n173 3.1505
R6015 VDD.n178 VDD.n177 3.1505
R6016 VDD.n177 VDD.n176 3.1505
R6017 VDD.n185 VDD.n184 3.1505
R6018 VDD.n184 VDD.n183 3.1505
R6019 VDD.n188 VDD.n187 3.1505
R6020 VDD.n187 VDD.n186 3.1505
R6021 VDD.n192 VDD.n191 3.1505
R6022 VDD.n191 VDD.n190 3.1505
R6023 VDD.n195 VDD.n194 3.1505
R6024 VDD.n534 VDD.n533 3.1505
R6025 VDD.n532 VDD.n531 3.1505
R6026 VDD.n529 VDD.n528 3.1505
R6027 VDD.n527 VDD.n526 3.1505
R6028 VDD.n524 VDD.n523 3.1505
R6029 VDD.n522 VDD.n521 3.1505
R6030 VDD.n519 VDD.n518 3.1505
R6031 VDD.n517 VDD.n516 3.1505
R6032 VDD.n514 VDD.n513 3.1505
R6033 VDD.n512 VDD.n511 3.1505
R6034 VDD.n509 VDD.n508 3.1505
R6035 VDD.n507 VDD.n506 3.1505
R6036 VDD.n504 VDD.n503 3.1505
R6037 VDD.n502 VDD.n501 3.1505
R6038 VDD.n499 VDD.n498 3.1505
R6039 VDD.n497 VDD.n496 3.1505
R6040 VDD.n494 VDD.n493 3.1505
R6041 VDD.n492 VDD.n491 3.1505
R6042 VDD.n489 VDD.n488 3.1505
R6043 VDD.n487 VDD.n486 3.1505
R6044 VDD.n484 VDD.n483 3.1505
R6045 VDD.n482 VDD.n481 3.1505
R6046 VDD.n479 VDD.n478 3.1505
R6047 VDD.n477 VDD.n476 3.1505
R6048 VDD.n475 VDD.n474 3.1505
R6049 VDD.n473 VDD.n472 3.1505
R6050 VDD.n471 VDD.n470 3.1505
R6051 VDD.n469 VDD.n468 3.1505
R6052 VDD.n467 VDD.n466 3.1505
R6053 VDD.n465 VDD.n464 3.1505
R6054 VDD.n463 VDD.n462 3.1505
R6055 VDD.n461 VDD.n460 3.1505
R6056 VDD.n459 VDD.n458 3.1505
R6057 VDD.n457 VDD.n456 3.1505
R6058 VDD.n7503 VDD.n7502 3.1505
R6059 VDD.n7426 VDD.n7425 3.1505
R6060 VDD.n7498 VDD.n7497 3.1505
R6061 VDD.n7496 VDD.n7495 3.1505
R6062 VDD.n7493 VDD.n7492 3.1505
R6063 VDD.n7491 VDD.n7490 3.1505
R6064 VDD.n7488 VDD.n7487 3.1505
R6065 VDD.n7486 VDD.n7485 3.1505
R6066 VDD.n7483 VDD.n7482 3.1505
R6067 VDD.n7481 VDD.n7480 3.1505
R6068 VDD.n7478 VDD.n7477 3.1505
R6069 VDD.n7476 VDD.n7475 3.1505
R6070 VDD.n7473 VDD.n7472 3.1505
R6071 VDD.n7471 VDD.n7470 3.1505
R6072 VDD.n7468 VDD.n7467 3.1505
R6073 VDD.n7466 VDD.n7465 3.1505
R6074 VDD.n7463 VDD.n7462 3.1505
R6075 VDD.n7461 VDD.n7460 3.1505
R6076 VDD.n7458 VDD.n7457 3.1505
R6077 VDD.n7456 VDD.n7455 3.1505
R6078 VDD.n7453 VDD.n7452 3.1505
R6079 VDD.n7451 VDD.n7450 3.1505
R6080 VDD.n7448 VDD.n7447 3.1505
R6081 VDD.n7446 VDD.n7445 3.1505
R6082 VDD.n7444 VDD.n7443 3.1505
R6083 VDD.n7442 VDD.n7441 3.1505
R6084 VDD.n7440 VDD.n7439 3.1505
R6085 VDD.n7438 VDD.n7437 3.1505
R6086 VDD.n7436 VDD.n7435 3.1505
R6087 VDD.n7434 VDD.n7433 3.1505
R6088 VDD.n7432 VDD.n7431 3.1505
R6089 VDD.n7430 VDD.n7429 3.1505
R6090 VDD.n7428 VDD.n7427 3.1505
R6091 VDD.n7501 VDD.n7500 3.1505
R6092 VDD.n7423 VDD.n7422 3.1505
R6093 VDD.n452 VDD.n451 3.1505
R6094 VDD.n450 VDD.n449 3.1505
R6095 VDD.n448 VDD.n447 3.1505
R6096 VDD.n445 VDD.n444 3.1505
R6097 VDD.n443 VDD.n442 3.1505
R6098 VDD.n440 VDD.n439 3.1505
R6099 VDD.n438 VDD.n437 3.1505
R6100 VDD.n436 VDD.n435 3.1505
R6101 VDD.n434 VDD.n433 3.1505
R6102 VDD.n432 VDD.n431 3.1505
R6103 VDD.n430 VDD.n429 3.1505
R6104 VDD.n428 VDD.n427 3.1505
R6105 VDD.n426 VDD.n425 3.1505
R6106 VDD.n424 VDD.n423 3.1505
R6107 VDD.n422 VDD.n421 3.1505
R6108 VDD.n420 VDD.n419 3.1505
R6109 VDD.n418 VDD.n417 3.1505
R6110 VDD.n416 VDD.n415 3.1505
R6111 VDD.n414 VDD.n413 3.1505
R6112 VDD.n412 VDD.n411 3.1505
R6113 VDD.n410 VDD.n409 3.1505
R6114 VDD.n408 VDD.n407 3.1505
R6115 VDD.n406 VDD.n405 3.1505
R6116 VDD.n7382 VDD.n7381 3.1505
R6117 VDD.n7384 VDD.n7383 3.1505
R6118 VDD.n7386 VDD.n7385 3.1505
R6119 VDD.n7388 VDD.n7387 3.1505
R6120 VDD.n7390 VDD.n7389 3.1505
R6121 VDD.n7392 VDD.n7391 3.1505
R6122 VDD.n7394 VDD.n7393 3.1505
R6123 VDD.n7396 VDD.n7395 3.1505
R6124 VDD.n7398 VDD.n7397 3.1505
R6125 VDD.n7400 VDD.n7399 3.1505
R6126 VDD.n7402 VDD.n7401 3.1505
R6127 VDD.n7404 VDD.n7403 3.1505
R6128 VDD.n7406 VDD.n7405 3.1505
R6129 VDD.n7408 VDD.n7407 3.1505
R6130 VDD.n7412 VDD.n7411 3.1505
R6131 VDD.n7414 VDD.n7413 3.1505
R6132 VDD.n7417 VDD.n7416 3.1505
R6133 VDD.n7419 VDD.n7418 3.1505
R6134 VDD.n7421 VDD.n7420 3.1505
R6135 VDD.n454 VDD.n453 3.1505
R6136 VDD.n7512 VDD.n7511 3.1505
R6137 VDD.n546 VDD.n542 3.1505
R6138 VDD.n545 VDD.n544 3.1505
R6139 VDD.n544 VDD.n543 3.1505
R6140 VDD.n307 VDD.n306 3.1505
R6141 VDD.n306 VDD.n305 3.1505
R6142 VDD.n310 VDD.n309 3.1505
R6143 VDD.n309 VDD.n308 3.1505
R6144 VDD.n313 VDD.n312 3.1505
R6145 VDD.n312 VDD.n311 3.1505
R6146 VDD.n317 VDD.n316 3.1505
R6147 VDD.n316 VDD.n315 3.1505
R6148 VDD.n320 VDD.n319 3.1505
R6149 VDD.n319 VDD.n318 3.1505
R6150 VDD.n324 VDD.n323 3.1505
R6151 VDD.n323 VDD.n322 3.1505
R6152 VDD.n328 VDD.n327 3.1505
R6153 VDD.n327 VDD.n326 3.1505
R6154 VDD.n331 VDD.n330 3.1505
R6155 VDD.n330 VDD.n329 3.1505
R6156 VDD.n334 VDD.n333 3.1505
R6157 VDD.n333 VDD.n332 3.1505
R6158 VDD.n385 VDD.n384 3.1505
R6159 VDD.n384 VDD.n383 3.1505
R6160 VDD.n382 VDD.n381 3.1505
R6161 VDD.n381 VDD.n380 3.1505
R6162 VDD.n378 VDD.n377 3.1505
R6163 VDD.n377 VDD.n376 3.1505
R6164 VDD.n375 VDD.n374 3.1505
R6165 VDD.n374 VDD.n373 3.1505
R6166 VDD.n372 VDD.n371 3.1505
R6167 VDD.n371 VDD.n370 3.1505
R6168 VDD.n369 VDD.n368 3.1505
R6169 VDD.n368 VDD.n367 3.1505
R6170 VDD.n365 VDD.n364 3.1505
R6171 VDD.n364 VDD.n363 3.1505
R6172 VDD.n362 VDD.n361 3.1505
R6173 VDD.n361 VDD.n360 3.1505
R6174 VDD.n359 VDD.n358 3.1505
R6175 VDD.n358 VDD.n357 3.1505
R6176 VDD.n356 VDD.n355 3.1505
R6177 VDD.n355 VDD.n354 3.1505
R6178 VDD.n353 VDD.n352 3.1505
R6179 VDD.n352 VDD.n351 3.1505
R6180 VDD.n349 VDD.n348 3.1505
R6181 VDD.n348 VDD.n347 3.1505
R6182 VDD.n346 VDD.n345 3.1505
R6183 VDD.n345 VDD.n344 3.1505
R6184 VDD.n343 VDD.n342 3.1505
R6185 VDD.n342 VDD.n341 3.1505
R6186 VDD.n7324 VDD.n7323 3.1505
R6187 VDD.n7323 VDD.n7322 3.1505
R6188 VDD.n7327 VDD.n7326 3.1505
R6189 VDD.n7326 VDD.n7325 3.1505
R6190 VDD.n7331 VDD.n7330 3.1505
R6191 VDD.n7330 VDD.n7329 3.1505
R6192 VDD.n7334 VDD.n7333 3.1505
R6193 VDD.n7333 VDD.n7332 3.1505
R6194 VDD.n7337 VDD.n7336 3.1505
R6195 VDD.n7336 VDD.n7335 3.1505
R6196 VDD.n7340 VDD.n7339 3.1505
R6197 VDD.n7339 VDD.n7338 3.1505
R6198 VDD.n7344 VDD.n7343 3.1505
R6199 VDD.n7343 VDD.n7342 3.1505
R6200 VDD.n7347 VDD.n7346 3.1505
R6201 VDD.n7346 VDD.n7345 3.1505
R6202 VDD.n7350 VDD.n7349 3.1505
R6203 VDD.n7349 VDD.n7348 3.1505
R6204 VDD.n7353 VDD.n7352 3.1505
R6205 VDD.n7352 VDD.n7351 3.1505
R6206 VDD.n7357 VDD.n7356 3.1505
R6207 VDD.n7356 VDD.n7355 3.1505
R6208 VDD.n7536 VDD.n7535 3.1505
R6209 VDD.n7535 VDD.n7534 3.1505
R6210 VDD.n7532 VDD.n7531 3.1505
R6211 VDD.n7531 VDD.n7530 3.1505
R6212 VDD.n7528 VDD.n7527 3.1505
R6213 VDD.n7527 VDD.n7526 3.1505
R6214 VDD.n7525 VDD.n7524 3.1505
R6215 VDD.n7524 VDD.n7523 3.1505
R6216 VDD.n7521 VDD.n7520 3.1505
R6217 VDD.n7520 VDD.n7519 3.1505
R6218 VDD.n7518 VDD.n7517 3.1505
R6219 VDD.n7517 VDD.n7516 3.1505
R6220 VDD.n7515 VDD.n7514 3.1505
R6221 VDD.n7514 VDD.n7513 3.1505
R6222 VDD.n971 VDD.n970 3.1505
R6223 VDD.n775 VDD.n774 3.1505
R6224 VDD.n752 VDD.n751 3.1505
R6225 VDD.n749 VDD.n748 3.1505
R6226 VDD.n746 VDD.n745 3.1505
R6227 VDD.n743 VDD.n742 3.1505
R6228 VDD.n740 VDD.n739 3.1505
R6229 VDD.n737 VDD.n736 3.1505
R6230 VDD.n734 VDD.n733 3.1505
R6231 VDD.n731 VDD.n730 3.1505
R6232 VDD.n728 VDD.n727 3.1505
R6233 VDD.n725 VDD.n724 3.1505
R6234 VDD.n722 VDD.n721 3.1505
R6235 VDD.n719 VDD.n718 3.1505
R6236 VDD.n716 VDD.n715 3.1505
R6237 VDD.n713 VDD.n712 3.1505
R6238 VDD.n710 VDD.n709 3.1505
R6239 VDD.n707 VDD.n706 3.1505
R6240 VDD.n704 VDD.n703 3.1505
R6241 VDD.n701 VDD.n700 3.1505
R6242 VDD.n698 VDD.n697 3.1505
R6243 VDD.n695 VDD.n694 3.1505
R6244 VDD.n692 VDD.n691 3.1505
R6245 VDD.n689 VDD.n688 3.1505
R6246 VDD.n686 VDD.n685 3.1505
R6247 VDD.n683 VDD.n682 3.1505
R6248 VDD.n680 VDD.n679 3.1505
R6249 VDD.n677 VDD.n676 3.1505
R6250 VDD.n674 VDD.n673 3.1505
R6251 VDD.n672 VDD.n671 3.1505
R6252 VDD.n670 VDD.n669 3.1505
R6253 VDD.n668 VDD.n667 3.1505
R6254 VDD.n666 VDD.n665 3.1505
R6255 VDD.n664 VDD.n663 3.1505
R6256 VDD.n662 VDD.n661 3.1505
R6257 VDD.n660 VDD.n659 3.1505
R6258 VDD.n658 VDD.n657 3.1505
R6259 VDD.n656 VDD.n655 3.1505
R6260 VDD.n654 VDD.n653 3.1505
R6261 VDD.n652 VDD.n651 3.1505
R6262 VDD.n650 VDD.n649 3.1505
R6263 VDD.n648 VDD.n647 3.1505
R6264 VDD.n646 VDD.n645 3.1505
R6265 VDD.n644 VDD.n643 3.1505
R6266 VDD.n642 VDD.n641 3.1505
R6267 VDD.n640 VDD.n639 3.1505
R6268 VDD.n638 VDD.n637 3.1505
R6269 VDD.n836 VDD.n835 3.1505
R6270 VDD.n946 VDD.n945 3.1505
R6271 VDD.n943 VDD.n942 3.1505
R6272 VDD.n940 VDD.n939 3.1505
R6273 VDD.n937 VDD.n936 3.1505
R6274 VDD.n934 VDD.n933 3.1505
R6275 VDD.n931 VDD.n930 3.1505
R6276 VDD.n928 VDD.n927 3.1505
R6277 VDD.n925 VDD.n924 3.1505
R6278 VDD.n922 VDD.n921 3.1505
R6279 VDD.n919 VDD.n918 3.1505
R6280 VDD.n916 VDD.n915 3.1505
R6281 VDD.n913 VDD.n912 3.1505
R6282 VDD.n910 VDD.n909 3.1505
R6283 VDD.n907 VDD.n906 3.1505
R6284 VDD.n904 VDD.n903 3.1505
R6285 VDD.n901 VDD.n900 3.1505
R6286 VDD.n898 VDD.n897 3.1505
R6287 VDD.n895 VDD.n894 3.1505
R6288 VDD.n892 VDD.n891 3.1505
R6289 VDD.n889 VDD.n888 3.1505
R6290 VDD.n886 VDD.n885 3.1505
R6291 VDD.n883 VDD.n882 3.1505
R6292 VDD.n880 VDD.n879 3.1505
R6293 VDD.n877 VDD.n876 3.1505
R6294 VDD.n874 VDD.n873 3.1505
R6295 VDD.n872 VDD.n871 3.1505
R6296 VDD.n870 VDD.n869 3.1505
R6297 VDD.n868 VDD.n867 3.1505
R6298 VDD.n866 VDD.n865 3.1505
R6299 VDD.n864 VDD.n863 3.1505
R6300 VDD.n862 VDD.n861 3.1505
R6301 VDD.n860 VDD.n859 3.1505
R6302 VDD.n858 VDD.n857 3.1505
R6303 VDD.n856 VDD.n855 3.1505
R6304 VDD.n854 VDD.n853 3.1505
R6305 VDD.n852 VDD.n851 3.1505
R6306 VDD.n850 VDD.n849 3.1505
R6307 VDD.n848 VDD.n847 3.1505
R6308 VDD.n846 VDD.n845 3.1505
R6309 VDD.n844 VDD.n843 3.1505
R6310 VDD.n842 VDD.n841 3.1505
R6311 VDD.n840 VDD.n839 3.1505
R6312 VDD.n838 VDD.n837 3.1505
R6313 VDD.n948 VDD.n947 3.1505
R6314 VDD.n6785 VDD.n6784 3.1505
R6315 VDD.n6687 VDD.n6686 3.1505
R6316 VDD.n6689 VDD.n6688 3.1505
R6317 VDD.n6691 VDD.n6690 3.1505
R6318 VDD.n6693 VDD.n6692 3.1505
R6319 VDD.n6695 VDD.n6694 3.1505
R6320 VDD.n6697 VDD.n6696 3.1505
R6321 VDD.n6699 VDD.n6698 3.1505
R6322 VDD.n6701 VDD.n6700 3.1505
R6323 VDD.n6703 VDD.n6702 3.1505
R6324 VDD.n6705 VDD.n6704 3.1505
R6325 VDD.n6707 VDD.n6706 3.1505
R6326 VDD.n6709 VDD.n6708 3.1505
R6327 VDD.n6711 VDD.n6710 3.1505
R6328 VDD.n6713 VDD.n6712 3.1505
R6329 VDD.n6715 VDD.n6714 3.1505
R6330 VDD.n6717 VDD.n6716 3.1505
R6331 VDD.n6719 VDD.n6718 3.1505
R6332 VDD.n6721 VDD.n6720 3.1505
R6333 VDD.n6723 VDD.n6722 3.1505
R6334 VDD.n6725 VDD.n6724 3.1505
R6335 VDD.n6727 VDD.n6726 3.1505
R6336 VDD.n6729 VDD.n6728 3.1505
R6337 VDD.n6731 VDD.n6730 3.1505
R6338 VDD.n6733 VDD.n6732 3.1505
R6339 VDD.n6735 VDD.n6734 3.1505
R6340 VDD.n6737 VDD.n6736 3.1505
R6341 VDD.n6739 VDD.n6738 3.1505
R6342 VDD.n6741 VDD.n6740 3.1505
R6343 VDD.n6743 VDD.n6742 3.1505
R6344 VDD.n6745 VDD.n6744 3.1505
R6345 VDD.n6748 VDD.n6747 3.1505
R6346 VDD.n6750 VDD.n6749 3.1505
R6347 VDD.n6753 VDD.n6752 3.1505
R6348 VDD.n6755 VDD.n6754 3.1505
R6349 VDD.n6758 VDD.n6757 3.1505
R6350 VDD.n6760 VDD.n6759 3.1505
R6351 VDD.n6763 VDD.n6762 3.1505
R6352 VDD.n6765 VDD.n6764 3.1505
R6353 VDD.n6768 VDD.n6767 3.1505
R6354 VDD.n6770 VDD.n6769 3.1505
R6355 VDD.n6773 VDD.n6772 3.1505
R6356 VDD.n6775 VDD.n6774 3.1505
R6357 VDD.n6778 VDD.n6777 3.1505
R6358 VDD.n6780 VDD.n6779 3.1505
R6359 VDD.n6783 VDD.n6782 3.1505
R6360 VDD.n6685 VDD.n6648 3.1505
R6361 VDD.n6684 VDD.n6683 3.1505
R6362 VDD.n6682 VDD.n6681 3.1505
R6363 VDD.n6679 VDD.n6678 3.1505
R6364 VDD.n6677 VDD.n6676 3.1505
R6365 VDD.n6674 VDD.n6673 3.1505
R6366 VDD.n6672 VDD.n6671 3.1505
R6367 VDD.n6670 VDD.n6669 3.1505
R6368 VDD.n6667 VDD.n6666 3.1505
R6369 VDD.n6665 VDD.n6664 3.1505
R6370 VDD.n6663 VDD.n6662 3.1505
R6371 VDD.n6660 VDD.n6659 3.1505
R6372 VDD.n6658 VDD.n6657 3.1505
R6373 VDD.n806 VDD.n805 3.1505
R6374 VDD.n808 VDD.n807 3.1505
R6375 VDD.n811 VDD.n810 3.1505
R6376 VDD.n813 VDD.n812 3.1505
R6377 VDD.n815 VDD.n814 3.1505
R6378 VDD.n818 VDD.n817 3.1505
R6379 VDD.n820 VDD.n819 3.1505
R6380 VDD.n822 VDD.n821 3.1505
R6381 VDD.n825 VDD.n824 3.1505
R6382 VDD.n827 VDD.n826 3.1505
R6383 VDD.n830 VDD.n829 3.1505
R6384 VDD.n832 VDD.n831 3.1505
R6385 VDD.n834 VDD.n833 3.1505
R6386 VDD.n575 VDD.n574 3.1505
R6387 VDD.n578 VDD.n577 3.1505
R6388 VDD.n580 VDD.n579 3.1505
R6389 VDD.n583 VDD.n582 3.1505
R6390 VDD.n585 VDD.n584 3.1505
R6391 VDD.n587 VDD.n586 3.1505
R6392 VDD.n589 VDD.n588 3.1505
R6393 VDD.n591 VDD.n590 3.1505
R6394 VDD.n593 VDD.n592 3.1505
R6395 VDD.n595 VDD.n594 3.1505
R6396 VDD.n597 VDD.n596 3.1505
R6397 VDD.n599 VDD.n598 3.1505
R6398 VDD.n601 VDD.n600 3.1505
R6399 VDD.n603 VDD.n602 3.1505
R6400 VDD.n605 VDD.n604 3.1505
R6401 VDD.n607 VDD.n606 3.1505
R6402 VDD.n609 VDD.n608 3.1505
R6403 VDD.n611 VDD.n610 3.1505
R6404 VDD.n613 VDD.n612 3.1505
R6405 VDD.n615 VDD.n614 3.1505
R6406 VDD.n617 VDD.n616 3.1505
R6407 VDD.n619 VDD.n618 3.1505
R6408 VDD.n621 VDD.n620 3.1505
R6409 VDD.n623 VDD.n622 3.1505
R6410 VDD.n625 VDD.n624 3.1505
R6411 VDD.n629 VDD.n628 3.1505
R6412 VDD.n631 VDD.n630 3.1505
R6413 VDD.n634 VDD.n633 3.1505
R6414 VDD.n636 VDD.n635 3.1505
R6415 VDD.n5540 VDD.n5539 3.1505
R6416 VDD.n3335 VDD.n3334 3.1505
R6417 VDD.n3333 VDD.n3332 3.1505
R6418 VDD.n3330 VDD.n3329 3.1505
R6419 VDD.n3328 VDD.n3327 3.1505
R6420 VDD.n3325 VDD.n3324 3.1505
R6421 VDD.n5434 VDD.n5433 3.1505
R6422 VDD.n5437 VDD.n5436 3.1505
R6423 VDD.n5439 VDD.n5438 3.1505
R6424 VDD.n5442 VDD.n5441 3.1505
R6425 VDD.n5444 VDD.n5443 3.1505
R6426 VDD.n5447 VDD.n5446 3.1505
R6427 VDD.n5449 VDD.n5448 3.1505
R6428 VDD.n5452 VDD.n5451 3.1505
R6429 VDD.n5454 VDD.n5453 3.1505
R6430 VDD.n5457 VDD.n5456 3.1505
R6431 VDD.n5459 VDD.n5458 3.1505
R6432 VDD.n5462 VDD.n5461 3.1505
R6433 VDD.n5464 VDD.n5463 3.1505
R6434 VDD.n5467 VDD.n5466 3.1505
R6435 VDD.n5469 VDD.n5468 3.1505
R6436 VDD.n5472 VDD.n5471 3.1505
R6437 VDD.n5474 VDD.n5473 3.1505
R6438 VDD.n5477 VDD.n5476 3.1505
R6439 VDD.n5479 VDD.n5478 3.1505
R6440 VDD.n5482 VDD.n5481 3.1505
R6441 VDD.n5484 VDD.n5483 3.1505
R6442 VDD.n5487 VDD.n5486 3.1505
R6443 VDD.n5489 VDD.n5488 3.1505
R6444 VDD.n5492 VDD.n5491 3.1505
R6445 VDD.n5494 VDD.n5493 3.1505
R6446 VDD.n5497 VDD.n5496 3.1505
R6447 VDD.n5499 VDD.n5498 3.1505
R6448 VDD.n5502 VDD.n5501 3.1505
R6449 VDD.n5504 VDD.n5503 3.1505
R6450 VDD.n5507 VDD.n5506 3.1505
R6451 VDD.n5509 VDD.n5508 3.1505
R6452 VDD.n5512 VDD.n5511 3.1505
R6453 VDD.n5514 VDD.n5513 3.1505
R6454 VDD.n5517 VDD.n5516 3.1505
R6455 VDD.n5519 VDD.n5518 3.1505
R6456 VDD.n5522 VDD.n5521 3.1505
R6457 VDD.n5524 VDD.n5523 3.1505
R6458 VDD.n5527 VDD.n5526 3.1505
R6459 VDD.n5529 VDD.n5528 3.1505
R6460 VDD.n5532 VDD.n5531 3.1505
R6461 VDD.n5535 VDD.n5534 3.1505
R6462 VDD.n5537 VDD.n5536 3.1505
R6463 VDD.n5367 VDD.n5366 3.1505
R6464 VDD.n3261 VDD.n3260 3.1505
R6465 VDD.n3259 VDD.n3258 3.1505
R6466 VDD.n3257 VDD.n3256 3.1505
R6467 VDD.n5274 VDD.n5273 3.1505
R6468 VDD.n5276 VDD.n5275 3.1505
R6469 VDD.n5278 VDD.n5277 3.1505
R6470 VDD.n5280 VDD.n5279 3.1505
R6471 VDD.n5282 VDD.n5281 3.1505
R6472 VDD.n5284 VDD.n5283 3.1505
R6473 VDD.n5286 VDD.n5285 3.1505
R6474 VDD.n5288 VDD.n5287 3.1505
R6475 VDD.n5290 VDD.n5289 3.1505
R6476 VDD.n5292 VDD.n5291 3.1505
R6477 VDD.n5294 VDD.n5293 3.1505
R6478 VDD.n5296 VDD.n5295 3.1505
R6479 VDD.n5298 VDD.n5297 3.1505
R6480 VDD.n5300 VDD.n5299 3.1505
R6481 VDD.n5302 VDD.n5301 3.1505
R6482 VDD.n5304 VDD.n5303 3.1505
R6483 VDD.n5306 VDD.n5305 3.1505
R6484 VDD.n5308 VDD.n5307 3.1505
R6485 VDD.n5310 VDD.n5309 3.1505
R6486 VDD.n5312 VDD.n5311 3.1505
R6487 VDD.n5314 VDD.n5313 3.1505
R6488 VDD.n5316 VDD.n5315 3.1505
R6489 VDD.n5318 VDD.n5317 3.1505
R6490 VDD.n5320 VDD.n5319 3.1505
R6491 VDD.n5322 VDD.n5321 3.1505
R6492 VDD.n5325 VDD.n5324 3.1505
R6493 VDD.n5327 VDD.n5326 3.1505
R6494 VDD.n5330 VDD.n5329 3.1505
R6495 VDD.n5332 VDD.n5331 3.1505
R6496 VDD.n5335 VDD.n5334 3.1505
R6497 VDD.n5337 VDD.n5336 3.1505
R6498 VDD.n5340 VDD.n5339 3.1505
R6499 VDD.n5342 VDD.n5341 3.1505
R6500 VDD.n5345 VDD.n5344 3.1505
R6501 VDD.n5347 VDD.n5346 3.1505
R6502 VDD.n5350 VDD.n5349 3.1505
R6503 VDD.n5352 VDD.n5351 3.1505
R6504 VDD.n5355 VDD.n5354 3.1505
R6505 VDD.n5357 VDD.n5356 3.1505
R6506 VDD.n5360 VDD.n5359 3.1505
R6507 VDD.n5362 VDD.n5361 3.1505
R6508 VDD.n5365 VDD.n5364 3.1505
R6509 VDD.n3263 VDD.n3262 3.1505
R6510 VDD.n3265 VDD.n3264 3.1505
R6511 VDD.n4575 VDD.n4574 3.1505
R6512 VDD.n4462 VDD.n4461 3.1505
R6513 VDD.n4465 VDD.n4464 3.1505
R6514 VDD.n4467 VDD.n4466 3.1505
R6515 VDD.n4470 VDD.n4469 3.1505
R6516 VDD.n4472 VDD.n4471 3.1505
R6517 VDD.n4475 VDD.n4474 3.1505
R6518 VDD.n4477 VDD.n4476 3.1505
R6519 VDD.n4480 VDD.n4479 3.1505
R6520 VDD.n4482 VDD.n4481 3.1505
R6521 VDD.n4485 VDD.n4484 3.1505
R6522 VDD.n4487 VDD.n4486 3.1505
R6523 VDD.n4490 VDD.n4489 3.1505
R6524 VDD.n4492 VDD.n4491 3.1505
R6525 VDD.n4495 VDD.n4494 3.1505
R6526 VDD.n4497 VDD.n4496 3.1505
R6527 VDD.n4500 VDD.n4499 3.1505
R6528 VDD.n4502 VDD.n4501 3.1505
R6529 VDD.n4505 VDD.n4504 3.1505
R6530 VDD.n4507 VDD.n4506 3.1505
R6531 VDD.n4510 VDD.n4509 3.1505
R6532 VDD.n4512 VDD.n4511 3.1505
R6533 VDD.n4515 VDD.n4514 3.1505
R6534 VDD.n4517 VDD.n4516 3.1505
R6535 VDD.n4520 VDD.n4519 3.1505
R6536 VDD.n4522 VDD.n4521 3.1505
R6537 VDD.n4525 VDD.n4524 3.1505
R6538 VDD.n4527 VDD.n4526 3.1505
R6539 VDD.n4530 VDD.n4529 3.1505
R6540 VDD.n4532 VDD.n4531 3.1505
R6541 VDD.n4535 VDD.n4534 3.1505
R6542 VDD.n4537 VDD.n4536 3.1505
R6543 VDD.n4540 VDD.n4539 3.1505
R6544 VDD.n4542 VDD.n4541 3.1505
R6545 VDD.n4545 VDD.n4544 3.1505
R6546 VDD.n4547 VDD.n4546 3.1505
R6547 VDD.n4550 VDD.n4549 3.1505
R6548 VDD.n4552 VDD.n4551 3.1505
R6549 VDD.n4555 VDD.n4554 3.1505
R6550 VDD.n4557 VDD.n4556 3.1505
R6551 VDD.n4560 VDD.n4559 3.1505
R6552 VDD.n4562 VDD.n4561 3.1505
R6553 VDD.n4565 VDD.n4564 3.1505
R6554 VDD.n4567 VDD.n4566 3.1505
R6555 VDD.n4570 VDD.n4569 3.1505
R6556 VDD.n4572 VDD.n4571 3.1505
R6557 VDD.n4460 VDD.n4459 3.1505
R6558 VDD.n4457 VDD.n4456 3.1505
R6559 VDD.n4455 VDD.n4454 3.1505
R6560 VDD.n3041 VDD.n3040 3.1505
R6561 VDD.n4385 VDD.n4384 3.1505
R6562 VDD.n4272 VDD.n4271 3.1505
R6563 VDD.n4274 VDD.n4273 3.1505
R6564 VDD.n4277 VDD.n4276 3.1505
R6565 VDD.n4279 VDD.n4278 3.1505
R6566 VDD.n4282 VDD.n4281 3.1505
R6567 VDD.n4284 VDD.n4283 3.1505
R6568 VDD.n4287 VDD.n4286 3.1505
R6569 VDD.n4289 VDD.n4288 3.1505
R6570 VDD.n4292 VDD.n4291 3.1505
R6571 VDD.n4294 VDD.n4293 3.1505
R6572 VDD.n4297 VDD.n4296 3.1505
R6573 VDD.n4299 VDD.n4298 3.1505
R6574 VDD.n4302 VDD.n4301 3.1505
R6575 VDD.n4304 VDD.n4303 3.1505
R6576 VDD.n4307 VDD.n4306 3.1505
R6577 VDD.n4309 VDD.n4308 3.1505
R6578 VDD.n4312 VDD.n4311 3.1505
R6579 VDD.n4314 VDD.n4313 3.1505
R6580 VDD.n4317 VDD.n4316 3.1505
R6581 VDD.n4319 VDD.n4318 3.1505
R6582 VDD.n4322 VDD.n4321 3.1505
R6583 VDD.n4324 VDD.n4323 3.1505
R6584 VDD.n4327 VDD.n4326 3.1505
R6585 VDD.n4329 VDD.n4328 3.1505
R6586 VDD.n4332 VDD.n4331 3.1505
R6587 VDD.n4334 VDD.n4333 3.1505
R6588 VDD.n4337 VDD.n4336 3.1505
R6589 VDD.n4339 VDD.n4338 3.1505
R6590 VDD.n4342 VDD.n4341 3.1505
R6591 VDD.n4344 VDD.n4343 3.1505
R6592 VDD.n4347 VDD.n4346 3.1505
R6593 VDD.n4349 VDD.n4348 3.1505
R6594 VDD.n4352 VDD.n4351 3.1505
R6595 VDD.n4354 VDD.n4353 3.1505
R6596 VDD.n4357 VDD.n4356 3.1505
R6597 VDD.n4359 VDD.n4358 3.1505
R6598 VDD.n4362 VDD.n4361 3.1505
R6599 VDD.n4364 VDD.n4363 3.1505
R6600 VDD.n4367 VDD.n4366 3.1505
R6601 VDD.n4369 VDD.n4368 3.1505
R6602 VDD.n4372 VDD.n4371 3.1505
R6603 VDD.n4374 VDD.n4373 3.1505
R6604 VDD.n4377 VDD.n4376 3.1505
R6605 VDD.n4380 VDD.n4379 3.1505
R6606 VDD.n4382 VDD.n4381 3.1505
R6607 VDD.n2973 VDD.n2972 3.1505
R6608 VDD.n2976 VDD.n2975 3.1505
R6609 VDD.n4065 VDD.n4064 3.1505
R6610 VDD.n4063 VDD.n4062 3.1505
R6611 VDD.n3963 VDD.n3962 3.1505
R6612 VDD.n3965 VDD.n3964 3.1505
R6613 VDD.n3967 VDD.n3966 3.1505
R6614 VDD.n3969 VDD.n3968 3.1505
R6615 VDD.n3971 VDD.n3970 3.1505
R6616 VDD.n3973 VDD.n3972 3.1505
R6617 VDD.n3975 VDD.n3974 3.1505
R6618 VDD.n3977 VDD.n3976 3.1505
R6619 VDD.n3979 VDD.n3978 3.1505
R6620 VDD.n3981 VDD.n3980 3.1505
R6621 VDD.n3983 VDD.n3982 3.1505
R6622 VDD.n3985 VDD.n3984 3.1505
R6623 VDD.n3987 VDD.n3986 3.1505
R6624 VDD.n3989 VDD.n3988 3.1505
R6625 VDD.n3991 VDD.n3990 3.1505
R6626 VDD.n3993 VDD.n3992 3.1505
R6627 VDD.n3995 VDD.n3994 3.1505
R6628 VDD.n3997 VDD.n3996 3.1505
R6629 VDD.n3999 VDD.n3998 3.1505
R6630 VDD.n4001 VDD.n4000 3.1505
R6631 VDD.n4003 VDD.n4002 3.1505
R6632 VDD.n4005 VDD.n4004 3.1505
R6633 VDD.n4007 VDD.n4006 3.1505
R6634 VDD.n4009 VDD.n4008 3.1505
R6635 VDD.n4011 VDD.n4010 3.1505
R6636 VDD.n4013 VDD.n4012 3.1505
R6637 VDD.n4015 VDD.n4014 3.1505
R6638 VDD.n4018 VDD.n4017 3.1505
R6639 VDD.n4020 VDD.n4019 3.1505
R6640 VDD.n4023 VDD.n4022 3.1505
R6641 VDD.n4025 VDD.n4024 3.1505
R6642 VDD.n4028 VDD.n4027 3.1505
R6643 VDD.n4030 VDD.n4029 3.1505
R6644 VDD.n4033 VDD.n4032 3.1505
R6645 VDD.n4035 VDD.n4034 3.1505
R6646 VDD.n4038 VDD.n4037 3.1505
R6647 VDD.n4040 VDD.n4039 3.1505
R6648 VDD.n4043 VDD.n4042 3.1505
R6649 VDD.n4045 VDD.n4044 3.1505
R6650 VDD.n4048 VDD.n4047 3.1505
R6651 VDD.n4050 VDD.n4049 3.1505
R6652 VDD.n4053 VDD.n4052 3.1505
R6653 VDD.n4055 VDD.n4054 3.1505
R6654 VDD.n4058 VDD.n4057 3.1505
R6655 VDD.n4060 VDD.n4059 3.1505
R6656 VDD.n3961 VDD.n3960 3.1505
R6657 VDD.n3959 VDD.n3958 3.1505
R6658 VDD.n3957 VDD.n3956 3.1505
R6659 VDD.n2911 VDD.n2910 3.1505
R6660 VDD.n6482 VDD.n6481 3.1505
R6661 VDD.n6461 VDD.n6460 3.1505
R6662 VDD.n6481 VDD.n6480 3.1505
R6663 VDD.n4269 VDD.n4268 3.1505
R6664 VDD.n2971 VDD.n2970 3.1505
R6665 VDD.n4264 VDD.n4263 3.1505
R6666 VDD.n4261 VDD.n4260 3.1505
R6667 VDD.n4258 VDD.n4257 3.1505
R6668 VDD.n4255 VDD.n4254 3.1505
R6669 VDD.n4252 VDD.n4251 3.1505
R6670 VDD.n4249 VDD.n4248 3.1505
R6671 VDD.n4246 VDD.n4245 3.1505
R6672 VDD.n4243 VDD.n4242 3.1505
R6673 VDD.n4240 VDD.n4239 3.1505
R6674 VDD.n4237 VDD.n4236 3.1505
R6675 VDD.n4234 VDD.n4233 3.1505
R6676 VDD.n4231 VDD.n4230 3.1505
R6677 VDD.n4228 VDD.n4227 3.1505
R6678 VDD.n4225 VDD.n4224 3.1505
R6679 VDD.n4222 VDD.n4221 3.1505
R6680 VDD.n4219 VDD.n4218 3.1505
R6681 VDD.n4216 VDD.n4215 3.1505
R6682 VDD.n4213 VDD.n4212 3.1505
R6683 VDD.n4210 VDD.n4209 3.1505
R6684 VDD.n4207 VDD.n4206 3.1505
R6685 VDD.n4204 VDD.n4203 3.1505
R6686 VDD.n4201 VDD.n4200 3.1505
R6687 VDD.n4198 VDD.n4197 3.1505
R6688 VDD.n4195 VDD.n4194 3.1505
R6689 VDD.n4192 VDD.n4191 3.1505
R6690 VDD.n4189 VDD.n4188 3.1505
R6691 VDD.n4186 VDD.n4185 3.1505
R6692 VDD.n4183 VDD.n4182 3.1505
R6693 VDD.n4180 VDD.n4179 3.1505
R6694 VDD.n4177 VDD.n4176 3.1505
R6695 VDD.n4174 VDD.n4173 3.1505
R6696 VDD.n4171 VDD.n4170 3.1505
R6697 VDD.n4168 VDD.n4167 3.1505
R6698 VDD.n4165 VDD.n4164 3.1505
R6699 VDD.n4162 VDD.n4161 3.1505
R6700 VDD.n4159 VDD.n4158 3.1505
R6701 VDD.n4156 VDD.n4155 3.1505
R6702 VDD.n4153 VDD.n4152 3.1505
R6703 VDD.n4150 VDD.n4149 3.1505
R6704 VDD.n4147 VDD.n4146 3.1505
R6705 VDD.n4144 VDD.n4143 3.1505
R6706 VDD.n4141 VDD.n4140 3.1505
R6707 VDD.n4138 VDD.n4137 3.1505
R6708 VDD.n4135 VDD.n4134 3.1505
R6709 VDD.n2969 VDD.n2968 3.1505
R6710 VDD.n4266 VDD.n4265 3.1505
R6711 VDD.n3846 VDD.n3845 3.1505
R6712 VDD.n3748 VDD.n3747 3.1505
R6713 VDD.n3750 VDD.n3749 3.1505
R6714 VDD.n3752 VDD.n3751 3.1505
R6715 VDD.n3754 VDD.n3753 3.1505
R6716 VDD.n3757 VDD.n3756 3.1505
R6717 VDD.n3759 VDD.n3758 3.1505
R6718 VDD.n3762 VDD.n3761 3.1505
R6719 VDD.n3764 VDD.n3763 3.1505
R6720 VDD.n3766 VDD.n3765 3.1505
R6721 VDD.n3769 VDD.n3768 3.1505
R6722 VDD.n3771 VDD.n3770 3.1505
R6723 VDD.n3773 VDD.n3772 3.1505
R6724 VDD.n3776 VDD.n3775 3.1505
R6725 VDD.n3778 VDD.n3777 3.1505
R6726 VDD.n3780 VDD.n3779 3.1505
R6727 VDD.n3783 VDD.n3782 3.1505
R6728 VDD.n3785 VDD.n3784 3.1505
R6729 VDD.n3787 VDD.n3786 3.1505
R6730 VDD.n3789 VDD.n3788 3.1505
R6731 VDD.n3791 VDD.n3790 3.1505
R6732 VDD.n3793 VDD.n3792 3.1505
R6733 VDD.n3795 VDD.n3794 3.1505
R6734 VDD.n3797 VDD.n3796 3.1505
R6735 VDD.n3799 VDD.n3798 3.1505
R6736 VDD.n3801 VDD.n3800 3.1505
R6737 VDD.n3803 VDD.n3802 3.1505
R6738 VDD.n3806 VDD.n3805 3.1505
R6739 VDD.n3808 VDD.n3807 3.1505
R6740 VDD.n3810 VDD.n3809 3.1505
R6741 VDD.n3813 VDD.n3812 3.1505
R6742 VDD.n3815 VDD.n3814 3.1505
R6743 VDD.n3817 VDD.n3816 3.1505
R6744 VDD.n3820 VDD.n3819 3.1505
R6745 VDD.n3822 VDD.n3821 3.1505
R6746 VDD.n3824 VDD.n3823 3.1505
R6747 VDD.n3827 VDD.n3826 3.1505
R6748 VDD.n3829 VDD.n3828 3.1505
R6749 VDD.n3832 VDD.n3831 3.1505
R6750 VDD.n3834 VDD.n3833 3.1505
R6751 VDD.n3836 VDD.n3835 3.1505
R6752 VDD.n3838 VDD.n3837 3.1505
R6753 VDD.n3840 VDD.n3839 3.1505
R6754 VDD.n3846 VDD.n3843 3.1505
R6755 VDD.n3853 VDD.n3852 3.1505
R6756 VDD.n3855 VDD.n3854 3.1505
R6757 VDD.n3857 VDD.n3856 3.1505
R6758 VDD.n3859 VDD.n3858 3.1505
R6759 VDD.n3861 VDD.n3860 3.1505
R6760 VDD.n3864 VDD.n3863 3.1505
R6761 VDD.n3866 VDD.n3865 3.1505
R6762 VDD.n3869 VDD.n3868 3.1505
R6763 VDD.n3871 VDD.n3870 3.1505
R6764 VDD.n3873 VDD.n3872 3.1505
R6765 VDD.n3876 VDD.n3875 3.1505
R6766 VDD.n3878 VDD.n3877 3.1505
R6767 VDD.n3880 VDD.n3879 3.1505
R6768 VDD.n3883 VDD.n3882 3.1505
R6769 VDD.n3885 VDD.n3884 3.1505
R6770 VDD.n3887 VDD.n3886 3.1505
R6771 VDD.n3890 VDD.n3889 3.1505
R6772 VDD.n3892 VDD.n3891 3.1505
R6773 VDD.n3894 VDD.n3893 3.1505
R6774 VDD.n3896 VDD.n3895 3.1505
R6775 VDD.n3898 VDD.n3897 3.1505
R6776 VDD.n3900 VDD.n3899 3.1505
R6777 VDD.n3902 VDD.n3901 3.1505
R6778 VDD.n3904 VDD.n3903 3.1505
R6779 VDD.n3906 VDD.n3905 3.1505
R6780 VDD.n3908 VDD.n3907 3.1505
R6781 VDD.n3910 VDD.n3909 3.1505
R6782 VDD.n3913 VDD.n3912 3.1505
R6783 VDD.n3915 VDD.n3914 3.1505
R6784 VDD.n3917 VDD.n3916 3.1505
R6785 VDD.n3920 VDD.n3919 3.1505
R6786 VDD.n3922 VDD.n3921 3.1505
R6787 VDD.n3924 VDD.n3923 3.1505
R6788 VDD.n3927 VDD.n3926 3.1505
R6789 VDD.n3929 VDD.n3928 3.1505
R6790 VDD.n3931 VDD.n3930 3.1505
R6791 VDD.n3934 VDD.n3933 3.1505
R6792 VDD.n3936 VDD.n3935 3.1505
R6793 VDD.n3944 VDD.n3943 3.1505
R6794 VDD.n3946 VDD.n3945 3.1505
R6795 VDD.n3948 VDD.n3947 3.1505
R6796 VDD.n3950 VDD.n3949 3.1505
R6797 VDD.n6319 VDD.n6318 3.1505
R6798 VDD.n6165 VDD.n6163 3.1505
R6799 VDD.n6313 VDD.n6311 3.1505
R6800 VDD.n6319 VDD.n6315 3.1505
R6801 VDD.n6459 VDD.n6458 3.1505
R6802 VDD.n6458 VDD.n6457 3.1505
R6803 VDD.n6456 VDD.n6455 3.1505
R6804 VDD.n6455 VDD.n6454 3.1505
R6805 VDD.n6453 VDD.n6452 3.1505
R6806 VDD.n6452 VDD.n6451 3.1505
R6807 VDD.n6450 VDD.n6449 3.1505
R6808 VDD.n6449 VDD.n6448 3.1505
R6809 VDD.n6446 VDD.n6445 3.1505
R6810 VDD.n6445 VDD.n6444 3.1505
R6811 VDD.n6443 VDD.n6442 3.1505
R6812 VDD.n6442 VDD.n6441 3.1505
R6813 VDD.n6439 VDD.n6438 3.1505
R6814 VDD.n6438 VDD.n6437 3.1505
R6815 VDD.n6436 VDD.n6435 3.1505
R6816 VDD.n6435 VDD.n6434 3.1505
R6817 VDD.n6433 VDD.n6432 3.1505
R6818 VDD.n6432 VDD.n6431 3.1505
R6819 VDD.n6429 VDD.n6428 3.1505
R6820 VDD.n6428 VDD.n6427 3.1505
R6821 VDD.n6426 VDD.n6425 3.1505
R6822 VDD.n6425 VDD.n6424 3.1505
R6823 VDD.n6423 VDD.n6422 3.1505
R6824 VDD.n6422 VDD.n6421 3.1505
R6825 VDD.n6419 VDD.n6418 3.1505
R6826 VDD.n6418 VDD.n6417 3.1505
R6827 VDD.n6416 VDD.n6415 3.1505
R6828 VDD.n6415 VDD.n6414 3.1505
R6829 VDD.n6413 VDD.n6412 3.1505
R6830 VDD.n6412 VDD.n6411 3.1505
R6831 VDD.n6409 VDD.n6408 3.1505
R6832 VDD.n6408 VDD.n6407 3.1505
R6833 VDD.n6406 VDD.n6405 3.1505
R6834 VDD.n6405 VDD.n6404 3.1505
R6835 VDD.n6403 VDD.n6402 3.1505
R6836 VDD.n6402 VDD.n6401 3.1505
R6837 VDD.n6400 VDD.n6399 3.1505
R6838 VDD.n6399 VDD.n6398 3.1505
R6839 VDD.n6396 VDD.n6395 3.1505
R6840 VDD.n6395 VDD.n6394 3.1505
R6841 VDD.n6393 VDD.n6392 3.1505
R6842 VDD.n6392 VDD.n6391 3.1505
R6843 VDD.n6390 VDD.n6389 3.1505
R6844 VDD.n6389 VDD.n6388 3.1505
R6845 VDD.n6386 VDD.n6385 3.1505
R6846 VDD.n6385 VDD.n6384 3.1505
R6847 VDD.n6383 VDD.n6382 3.1505
R6848 VDD.n6382 VDD.n6381 3.1505
R6849 VDD.n6380 VDD.n6379 3.1505
R6850 VDD.n6379 VDD.n6378 3.1505
R6851 VDD.n6377 VDD.n6376 3.1505
R6852 VDD.n6376 VDD.n6375 3.1505
R6853 VDD.n6373 VDD.n6372 3.1505
R6854 VDD.n6372 VDD.n6371 3.1505
R6855 VDD.n6370 VDD.n6369 3.1505
R6856 VDD.n6369 VDD.n6368 3.1505
R6857 VDD.n6367 VDD.n6366 3.1505
R6858 VDD.n6366 VDD.n6365 3.1505
R6859 VDD.n6363 VDD.n6362 3.1505
R6860 VDD.n6362 VDD.n6361 3.1505
R6861 VDD.n6360 VDD.n6359 3.1505
R6862 VDD.n6359 VDD.n6358 3.1505
R6863 VDD.n6357 VDD.n6356 3.1505
R6864 VDD.n6356 VDD.n6355 3.1505
R6865 VDD.n6353 VDD.n6352 3.1505
R6866 VDD.n6352 VDD.n6351 3.1505
R6867 VDD.n6350 VDD.n6349 3.1505
R6868 VDD.n6349 VDD.n6348 3.1505
R6869 VDD.n6347 VDD.n6346 3.1505
R6870 VDD.n6346 VDD.n6345 3.1505
R6871 VDD.n6343 VDD.n6342 3.1505
R6872 VDD.n6342 VDD.n6341 3.1505
R6873 VDD.n6340 VDD.n6339 3.1505
R6874 VDD.n6339 VDD.n6338 3.1505
R6875 VDD.n6336 VDD.n6335 3.1505
R6876 VDD.n6335 VDD.n6334 3.1505
R6877 VDD.n6333 VDD.n6332 3.1505
R6878 VDD.n6332 VDD.n6331 3.1505
R6879 VDD.n6330 VDD.n6329 3.1505
R6880 VDD.n6329 VDD.n6328 3.1505
R6881 VDD.n6327 VDD.n6326 3.1505
R6882 VDD.n6326 VDD.n6325 3.1505
R6883 VDD.n6324 VDD.n6323 3.1505
R6884 VDD.n6323 VDD.n6322 3.1505
R6885 VDD.n6160 VDD.n6159 3.1505
R6886 VDD.n6313 VDD.n6312 3.1505
R6887 VDD.n6307 VDD.n6306 3.1505
R6888 VDD.n6306 VDD.n6305 3.1505
R6889 VDD.n6304 VDD.n6303 3.1505
R6890 VDD.n6303 VDD.n6302 3.1505
R6891 VDD.n6301 VDD.n6300 3.1505
R6892 VDD.n6300 VDD.n6299 3.1505
R6893 VDD.n6298 VDD.n6297 3.1505
R6894 VDD.n6297 VDD.n6296 3.1505
R6895 VDD.n6295 VDD.n6294 3.1505
R6896 VDD.n6294 VDD.n6293 3.1505
R6897 VDD.n6291 VDD.n6290 3.1505
R6898 VDD.n6290 VDD.n6289 3.1505
R6899 VDD.n6288 VDD.n6287 3.1505
R6900 VDD.n6287 VDD.n6286 3.1505
R6901 VDD.n6284 VDD.n6283 3.1505
R6902 VDD.n6283 VDD.n6282 3.1505
R6903 VDD.n6281 VDD.n6280 3.1505
R6904 VDD.n6280 VDD.n6279 3.1505
R6905 VDD.n6278 VDD.n6277 3.1505
R6906 VDD.n6277 VDD.n6276 3.1505
R6907 VDD.n6274 VDD.n6273 3.1505
R6908 VDD.n6273 VDD.n6272 3.1505
R6909 VDD.n6271 VDD.n6270 3.1505
R6910 VDD.n6270 VDD.n6269 3.1505
R6911 VDD.n6268 VDD.n6267 3.1505
R6912 VDD.n6267 VDD.n6266 3.1505
R6913 VDD.n6264 VDD.n6263 3.1505
R6914 VDD.n6263 VDD.n6262 3.1505
R6915 VDD.n6261 VDD.n6260 3.1505
R6916 VDD.n6260 VDD.n6259 3.1505
R6917 VDD.n6258 VDD.n6257 3.1505
R6918 VDD.n6257 VDD.n6256 3.1505
R6919 VDD.n6254 VDD.n6253 3.1505
R6920 VDD.n6253 VDD.n6252 3.1505
R6921 VDD.n6251 VDD.n6250 3.1505
R6922 VDD.n6250 VDD.n6249 3.1505
R6923 VDD.n6248 VDD.n6247 3.1505
R6924 VDD.n6247 VDD.n6246 3.1505
R6925 VDD.n6245 VDD.n6244 3.1505
R6926 VDD.n6244 VDD.n6243 3.1505
R6927 VDD.n6241 VDD.n6240 3.1505
R6928 VDD.n6240 VDD.n6239 3.1505
R6929 VDD.n6238 VDD.n6237 3.1505
R6930 VDD.n6237 VDD.n6236 3.1505
R6931 VDD.n6235 VDD.n6234 3.1505
R6932 VDD.n6234 VDD.n6233 3.1505
R6933 VDD.n6231 VDD.n6230 3.1505
R6934 VDD.n6230 VDD.n6229 3.1505
R6935 VDD.n6228 VDD.n6227 3.1505
R6936 VDD.n6227 VDD.n6226 3.1505
R6937 VDD.n6225 VDD.n6224 3.1505
R6938 VDD.n6224 VDD.n6223 3.1505
R6939 VDD.n6222 VDD.n6221 3.1505
R6940 VDD.n6221 VDD.n6220 3.1505
R6941 VDD.n6218 VDD.n6217 3.1505
R6942 VDD.n6217 VDD.n6216 3.1505
R6943 VDD.n6215 VDD.n6214 3.1505
R6944 VDD.n6214 VDD.n6213 3.1505
R6945 VDD.n6212 VDD.n6211 3.1505
R6946 VDD.n6211 VDD.n6210 3.1505
R6947 VDD.n6208 VDD.n6207 3.1505
R6948 VDD.n6207 VDD.n6206 3.1505
R6949 VDD.n6205 VDD.n6204 3.1505
R6950 VDD.n6204 VDD.n6203 3.1505
R6951 VDD.n6202 VDD.n6201 3.1505
R6952 VDD.n6201 VDD.n6200 3.1505
R6953 VDD.n6198 VDD.n6197 3.1505
R6954 VDD.n6197 VDD.n6196 3.1505
R6955 VDD.n6195 VDD.n6194 3.1505
R6956 VDD.n6194 VDD.n6193 3.1505
R6957 VDD.n6192 VDD.n6191 3.1505
R6958 VDD.n6191 VDD.n6190 3.1505
R6959 VDD.n6188 VDD.n6187 3.1505
R6960 VDD.n6187 VDD.n6186 3.1505
R6961 VDD.n6185 VDD.n6184 3.1505
R6962 VDD.n6184 VDD.n6183 3.1505
R6963 VDD.n6181 VDD.n6180 3.1505
R6964 VDD.n6180 VDD.n6179 3.1505
R6965 VDD.n6178 VDD.n6177 3.1505
R6966 VDD.n6177 VDD.n6176 3.1505
R6967 VDD.n6175 VDD.n6174 3.1505
R6968 VDD.n6174 VDD.n6173 3.1505
R6969 VDD.n6172 VDD.n6171 3.1505
R6970 VDD.n6171 VDD.n6170 3.1505
R6971 VDD.n6169 VDD.n6168 3.1505
R6972 VDD.n6168 VDD.n6167 3.1505
R6973 VDD.n6165 VDD.n6164 3.1505
R6974 VDD.n6159 VDD.n6158 3.1505
R6975 VDD.n4776 VDD.n4775 3.1505
R6976 VDD.n3104 VDD.n3103 3.1505
R6977 VDD.n4771 VDD.n4770 3.1505
R6978 VDD.n4768 VDD.n4767 3.1505
R6979 VDD.n4765 VDD.n4764 3.1505
R6980 VDD.n4762 VDD.n4761 3.1505
R6981 VDD.n4759 VDD.n4758 3.1505
R6982 VDD.n4756 VDD.n4755 3.1505
R6983 VDD.n4753 VDD.n4752 3.1505
R6984 VDD.n4750 VDD.n4749 3.1505
R6985 VDD.n4747 VDD.n4746 3.1505
R6986 VDD.n4744 VDD.n4743 3.1505
R6987 VDD.n4741 VDD.n4740 3.1505
R6988 VDD.n4738 VDD.n4737 3.1505
R6989 VDD.n4735 VDD.n4734 3.1505
R6990 VDD.n4732 VDD.n4731 3.1505
R6991 VDD.n4729 VDD.n4728 3.1505
R6992 VDD.n4726 VDD.n4725 3.1505
R6993 VDD.n4723 VDD.n4722 3.1505
R6994 VDD.n4720 VDD.n4719 3.1505
R6995 VDD.n4717 VDD.n4716 3.1505
R6996 VDD.n4714 VDD.n4713 3.1505
R6997 VDD.n4711 VDD.n4710 3.1505
R6998 VDD.n4708 VDD.n4707 3.1505
R6999 VDD.n4705 VDD.n4704 3.1505
R7000 VDD.n4702 VDD.n4701 3.1505
R7001 VDD.n4699 VDD.n4698 3.1505
R7002 VDD.n4696 VDD.n4695 3.1505
R7003 VDD.n4693 VDD.n4692 3.1505
R7004 VDD.n4690 VDD.n4689 3.1505
R7005 VDD.n4687 VDD.n4686 3.1505
R7006 VDD.n4684 VDD.n4683 3.1505
R7007 VDD.n4681 VDD.n4680 3.1505
R7008 VDD.n4678 VDD.n4677 3.1505
R7009 VDD.n4675 VDD.n4674 3.1505
R7010 VDD.n4672 VDD.n4671 3.1505
R7011 VDD.n4669 VDD.n4668 3.1505
R7012 VDD.n4666 VDD.n4665 3.1505
R7013 VDD.n4663 VDD.n4662 3.1505
R7014 VDD.n4660 VDD.n4659 3.1505
R7015 VDD.n4657 VDD.n4656 3.1505
R7016 VDD.n4654 VDD.n4653 3.1505
R7017 VDD.n4651 VDD.n4650 3.1505
R7018 VDD.n4648 VDD.n4647 3.1505
R7019 VDD.n4645 VDD.n4644 3.1505
R7020 VDD.n3099 VDD.n3098 3.1505
R7021 VDD.n3102 VDD.n3101 3.1505
R7022 VDD.n4773 VDD.n4772 3.1505
R7023 VDD.n5075 VDD.n5074 3.1505
R7024 VDD.n4962 VDD.n4961 3.1505
R7025 VDD.n4965 VDD.n4964 3.1505
R7026 VDD.n4967 VDD.n4966 3.1505
R7027 VDD.n4970 VDD.n4969 3.1505
R7028 VDD.n4972 VDD.n4971 3.1505
R7029 VDD.n4975 VDD.n4974 3.1505
R7030 VDD.n4977 VDD.n4976 3.1505
R7031 VDD.n4980 VDD.n4979 3.1505
R7032 VDD.n4982 VDD.n4981 3.1505
R7033 VDD.n4985 VDD.n4984 3.1505
R7034 VDD.n4987 VDD.n4986 3.1505
R7035 VDD.n4990 VDD.n4989 3.1505
R7036 VDD.n4992 VDD.n4991 3.1505
R7037 VDD.n4995 VDD.n4994 3.1505
R7038 VDD.n4997 VDD.n4996 3.1505
R7039 VDD.n5000 VDD.n4999 3.1505
R7040 VDD.n5002 VDD.n5001 3.1505
R7041 VDD.n5005 VDD.n5004 3.1505
R7042 VDD.n5007 VDD.n5006 3.1505
R7043 VDD.n5010 VDD.n5009 3.1505
R7044 VDD.n5012 VDD.n5011 3.1505
R7045 VDD.n5015 VDD.n5014 3.1505
R7046 VDD.n5017 VDD.n5016 3.1505
R7047 VDD.n5020 VDD.n5019 3.1505
R7048 VDD.n5022 VDD.n5021 3.1505
R7049 VDD.n5025 VDD.n5024 3.1505
R7050 VDD.n5027 VDD.n5026 3.1505
R7051 VDD.n5030 VDD.n5029 3.1505
R7052 VDD.n5032 VDD.n5031 3.1505
R7053 VDD.n5035 VDD.n5034 3.1505
R7054 VDD.n5037 VDD.n5036 3.1505
R7055 VDD.n5040 VDD.n5039 3.1505
R7056 VDD.n5042 VDD.n5041 3.1505
R7057 VDD.n5045 VDD.n5044 3.1505
R7058 VDD.n5047 VDD.n5046 3.1505
R7059 VDD.n5050 VDD.n5049 3.1505
R7060 VDD.n5052 VDD.n5051 3.1505
R7061 VDD.n5055 VDD.n5054 3.1505
R7062 VDD.n5057 VDD.n5056 3.1505
R7063 VDD.n5060 VDD.n5059 3.1505
R7064 VDD.n5062 VDD.n5061 3.1505
R7065 VDD.n5065 VDD.n5064 3.1505
R7066 VDD.n5067 VDD.n5066 3.1505
R7067 VDD.n5070 VDD.n5069 3.1505
R7068 VDD.n5072 VDD.n5071 3.1505
R7069 VDD.n4960 VDD.n4959 3.1505
R7070 VDD.n3179 VDD.n3178 3.1505
R7071 VDD.n3181 VDD.n3180 3.1505
R7072 VDD.n3177 VDD.n3176 3.1505
R7073 VDD.n4889 VDD.n4888 3.1505
R7074 VDD.n3107 VDD.n3106 3.1505
R7075 VDD.n4778 VDD.n4777 3.1505
R7076 VDD.n4781 VDD.n4780 3.1505
R7077 VDD.n4783 VDD.n4782 3.1505
R7078 VDD.n4786 VDD.n4785 3.1505
R7079 VDD.n4788 VDD.n4787 3.1505
R7080 VDD.n4791 VDD.n4790 3.1505
R7081 VDD.n4793 VDD.n4792 3.1505
R7082 VDD.n4796 VDD.n4795 3.1505
R7083 VDD.n4798 VDD.n4797 3.1505
R7084 VDD.n4801 VDD.n4800 3.1505
R7085 VDD.n4803 VDD.n4802 3.1505
R7086 VDD.n4806 VDD.n4805 3.1505
R7087 VDD.n4808 VDD.n4807 3.1505
R7088 VDD.n4811 VDD.n4810 3.1505
R7089 VDD.n4813 VDD.n4812 3.1505
R7090 VDD.n4816 VDD.n4815 3.1505
R7091 VDD.n4818 VDD.n4817 3.1505
R7092 VDD.n4821 VDD.n4820 3.1505
R7093 VDD.n4823 VDD.n4822 3.1505
R7094 VDD.n4826 VDD.n4825 3.1505
R7095 VDD.n4828 VDD.n4827 3.1505
R7096 VDD.n4831 VDD.n4830 3.1505
R7097 VDD.n4833 VDD.n4832 3.1505
R7098 VDD.n4836 VDD.n4835 3.1505
R7099 VDD.n4838 VDD.n4837 3.1505
R7100 VDD.n4841 VDD.n4840 3.1505
R7101 VDD.n4843 VDD.n4842 3.1505
R7102 VDD.n4846 VDD.n4845 3.1505
R7103 VDD.n4848 VDD.n4847 3.1505
R7104 VDD.n4851 VDD.n4850 3.1505
R7105 VDD.n4853 VDD.n4852 3.1505
R7106 VDD.n4856 VDD.n4855 3.1505
R7107 VDD.n4858 VDD.n4857 3.1505
R7108 VDD.n4861 VDD.n4860 3.1505
R7109 VDD.n4863 VDD.n4862 3.1505
R7110 VDD.n4866 VDD.n4865 3.1505
R7111 VDD.n4868 VDD.n4867 3.1505
R7112 VDD.n4871 VDD.n4870 3.1505
R7113 VDD.n4873 VDD.n4872 3.1505
R7114 VDD.n4876 VDD.n4875 3.1505
R7115 VDD.n4878 VDD.n4877 3.1505
R7116 VDD.n4881 VDD.n4880 3.1505
R7117 VDD.n4884 VDD.n4883 3.1505
R7118 VDD.n4886 VDD.n4885 3.1505
R7119 VDD.n3109 VDD.n3108 3.1505
R7120 VDD.n3112 VDD.n3111 3.1505
R7121 VDD.n3641 VDD.n3640 3.1505
R7122 VDD.n3542 VDD.n3541 3.1505
R7123 VDD.n3544 VDD.n3543 3.1505
R7124 VDD.n3546 VDD.n3545 3.1505
R7125 VDD.n3548 VDD.n3547 3.1505
R7126 VDD.n3551 VDD.n3550 3.1505
R7127 VDD.n3553 VDD.n3552 3.1505
R7128 VDD.n3556 VDD.n3555 3.1505
R7129 VDD.n3558 VDD.n3557 3.1505
R7130 VDD.n3560 VDD.n3559 3.1505
R7131 VDD.n3563 VDD.n3562 3.1505
R7132 VDD.n3565 VDD.n3564 3.1505
R7133 VDD.n3567 VDD.n3566 3.1505
R7134 VDD.n3570 VDD.n3569 3.1505
R7135 VDD.n3572 VDD.n3571 3.1505
R7136 VDD.n3574 VDD.n3573 3.1505
R7137 VDD.n3577 VDD.n3576 3.1505
R7138 VDD.n3579 VDD.n3578 3.1505
R7139 VDD.n3581 VDD.n3580 3.1505
R7140 VDD.n3583 VDD.n3582 3.1505
R7141 VDD.n3585 VDD.n3584 3.1505
R7142 VDD.n3587 VDD.n3586 3.1505
R7143 VDD.n3589 VDD.n3588 3.1505
R7144 VDD.n3591 VDD.n3590 3.1505
R7145 VDD.n3593 VDD.n3592 3.1505
R7146 VDD.n3595 VDD.n3594 3.1505
R7147 VDD.n3597 VDD.n3596 3.1505
R7148 VDD.n3600 VDD.n3599 3.1505
R7149 VDD.n3602 VDD.n3601 3.1505
R7150 VDD.n3604 VDD.n3603 3.1505
R7151 VDD.n3607 VDD.n3606 3.1505
R7152 VDD.n3609 VDD.n3608 3.1505
R7153 VDD.n3611 VDD.n3610 3.1505
R7154 VDD.n3614 VDD.n3613 3.1505
R7155 VDD.n3616 VDD.n3615 3.1505
R7156 VDD.n3618 VDD.n3617 3.1505
R7157 VDD.n3621 VDD.n3620 3.1505
R7158 VDD.n3623 VDD.n3622 3.1505
R7159 VDD.n3626 VDD.n3625 3.1505
R7160 VDD.n3628 VDD.n3627 3.1505
R7161 VDD.n3630 VDD.n3629 3.1505
R7162 VDD.n3632 VDD.n3631 3.1505
R7163 VDD.n3634 VDD.n3633 3.1505
R7164 VDD.n3641 VDD.n3638 3.1505
R7165 VDD.n3648 VDD.n3647 3.1505
R7166 VDD.n3650 VDD.n3649 3.1505
R7167 VDD.n3652 VDD.n3651 3.1505
R7168 VDD.n3654 VDD.n3653 3.1505
R7169 VDD.n3656 VDD.n3655 3.1505
R7170 VDD.n3659 VDD.n3658 3.1505
R7171 VDD.n3661 VDD.n3660 3.1505
R7172 VDD.n3664 VDD.n3663 3.1505
R7173 VDD.n3666 VDD.n3665 3.1505
R7174 VDD.n3668 VDD.n3667 3.1505
R7175 VDD.n3671 VDD.n3670 3.1505
R7176 VDD.n3673 VDD.n3672 3.1505
R7177 VDD.n3675 VDD.n3674 3.1505
R7178 VDD.n3678 VDD.n3677 3.1505
R7179 VDD.n3680 VDD.n3679 3.1505
R7180 VDD.n3682 VDD.n3681 3.1505
R7181 VDD.n3685 VDD.n3684 3.1505
R7182 VDD.n3687 VDD.n3686 3.1505
R7183 VDD.n3689 VDD.n3688 3.1505
R7184 VDD.n3691 VDD.n3690 3.1505
R7185 VDD.n3693 VDD.n3692 3.1505
R7186 VDD.n3695 VDD.n3694 3.1505
R7187 VDD.n3697 VDD.n3696 3.1505
R7188 VDD.n3699 VDD.n3698 3.1505
R7189 VDD.n3701 VDD.n3700 3.1505
R7190 VDD.n3703 VDD.n3702 3.1505
R7191 VDD.n3705 VDD.n3704 3.1505
R7192 VDD.n3708 VDD.n3707 3.1505
R7193 VDD.n3710 VDD.n3709 3.1505
R7194 VDD.n3712 VDD.n3711 3.1505
R7195 VDD.n3715 VDD.n3714 3.1505
R7196 VDD.n3717 VDD.n3716 3.1505
R7197 VDD.n3719 VDD.n3718 3.1505
R7198 VDD.n3722 VDD.n3721 3.1505
R7199 VDD.n3724 VDD.n3723 3.1505
R7200 VDD.n3726 VDD.n3725 3.1505
R7201 VDD.n3729 VDD.n3728 3.1505
R7202 VDD.n3731 VDD.n3730 3.1505
R7203 VDD.n3739 VDD.n3738 3.1505
R7204 VDD.n3741 VDD.n3740 3.1505
R7205 VDD.n3743 VDD.n3742 3.1505
R7206 VDD.n3745 VDD.n3744 3.1505
R7207 VDD.n6017 VDD.n6016 3.1505
R7208 VDD.n5863 VDD.n5859 3.1505
R7209 VDD.n6011 VDD.n6009 3.1505
R7210 VDD.n6017 VDD.n6015 3.1505
R7211 VDD.n6157 VDD.n6156 3.1505
R7212 VDD.n6156 VDD.n6155 3.1505
R7213 VDD.n6154 VDD.n6153 3.1505
R7214 VDD.n6153 VDD.n6152 3.1505
R7215 VDD.n6151 VDD.n6150 3.1505
R7216 VDD.n6150 VDD.n6149 3.1505
R7217 VDD.n6148 VDD.n6147 3.1505
R7218 VDD.n6147 VDD.n6146 3.1505
R7219 VDD.n6144 VDD.n6143 3.1505
R7220 VDD.n6143 VDD.n6142 3.1505
R7221 VDD.n6141 VDD.n6140 3.1505
R7222 VDD.n6140 VDD.n6139 3.1505
R7223 VDD.n6137 VDD.n6136 3.1505
R7224 VDD.n6136 VDD.n6135 3.1505
R7225 VDD.n6134 VDD.n6133 3.1505
R7226 VDD.n6133 VDD.n6132 3.1505
R7227 VDD.n6131 VDD.n6130 3.1505
R7228 VDD.n6130 VDD.n6129 3.1505
R7229 VDD.n6127 VDD.n6126 3.1505
R7230 VDD.n6126 VDD.n6125 3.1505
R7231 VDD.n6124 VDD.n6123 3.1505
R7232 VDD.n6123 VDD.n6122 3.1505
R7233 VDD.n6121 VDD.n6120 3.1505
R7234 VDD.n6120 VDD.n6119 3.1505
R7235 VDD.n6117 VDD.n6116 3.1505
R7236 VDD.n6116 VDD.n6115 3.1505
R7237 VDD.n6114 VDD.n6113 3.1505
R7238 VDD.n6113 VDD.n6112 3.1505
R7239 VDD.n6111 VDD.n6110 3.1505
R7240 VDD.n6110 VDD.n6109 3.1505
R7241 VDD.n6107 VDD.n6106 3.1505
R7242 VDD.n6106 VDD.n6105 3.1505
R7243 VDD.n6104 VDD.n6103 3.1505
R7244 VDD.n6103 VDD.n6102 3.1505
R7245 VDD.n6101 VDD.n6100 3.1505
R7246 VDD.n6100 VDD.n6099 3.1505
R7247 VDD.n6098 VDD.n6097 3.1505
R7248 VDD.n6097 VDD.n6096 3.1505
R7249 VDD.n6094 VDD.n6093 3.1505
R7250 VDD.n6093 VDD.n6092 3.1505
R7251 VDD.n6091 VDD.n6090 3.1505
R7252 VDD.n6090 VDD.n6089 3.1505
R7253 VDD.n6088 VDD.n6087 3.1505
R7254 VDD.n6087 VDD.n6086 3.1505
R7255 VDD.n6084 VDD.n6083 3.1505
R7256 VDD.n6083 VDD.n6082 3.1505
R7257 VDD.n6081 VDD.n6080 3.1505
R7258 VDD.n6080 VDD.n6079 3.1505
R7259 VDD.n6078 VDD.n6077 3.1505
R7260 VDD.n6077 VDD.n6076 3.1505
R7261 VDD.n6075 VDD.n6074 3.1505
R7262 VDD.n6074 VDD.n6073 3.1505
R7263 VDD.n6071 VDD.n6070 3.1505
R7264 VDD.n6070 VDD.n6069 3.1505
R7265 VDD.n6068 VDD.n6067 3.1505
R7266 VDD.n6067 VDD.n6066 3.1505
R7267 VDD.n6065 VDD.n6064 3.1505
R7268 VDD.n6064 VDD.n6063 3.1505
R7269 VDD.n6061 VDD.n6060 3.1505
R7270 VDD.n6060 VDD.n6059 3.1505
R7271 VDD.n6058 VDD.n6057 3.1505
R7272 VDD.n6057 VDD.n6056 3.1505
R7273 VDD.n6055 VDD.n6054 3.1505
R7274 VDD.n6054 VDD.n6053 3.1505
R7275 VDD.n6051 VDD.n6050 3.1505
R7276 VDD.n6050 VDD.n6049 3.1505
R7277 VDD.n6048 VDD.n6047 3.1505
R7278 VDD.n6047 VDD.n6046 3.1505
R7279 VDD.n6045 VDD.n6044 3.1505
R7280 VDD.n6044 VDD.n6043 3.1505
R7281 VDD.n6041 VDD.n6040 3.1505
R7282 VDD.n6040 VDD.n6039 3.1505
R7283 VDD.n6038 VDD.n6037 3.1505
R7284 VDD.n6037 VDD.n6036 3.1505
R7285 VDD.n6034 VDD.n6033 3.1505
R7286 VDD.n6033 VDD.n6032 3.1505
R7287 VDD.n6031 VDD.n6030 3.1505
R7288 VDD.n6030 VDD.n6029 3.1505
R7289 VDD.n6028 VDD.n6027 3.1505
R7290 VDD.n6027 VDD.n6026 3.1505
R7291 VDD.n6025 VDD.n6024 3.1505
R7292 VDD.n6024 VDD.n6023 3.1505
R7293 VDD.n6022 VDD.n6021 3.1505
R7294 VDD.n6021 VDD.n6020 3.1505
R7295 VDD.n5858 VDD.n5857 3.1505
R7296 VDD.n6011 VDD.n6010 3.1505
R7297 VDD.n6005 VDD.n6004 3.1505
R7298 VDD.n6004 VDD.n6003 3.1505
R7299 VDD.n6002 VDD.n6001 3.1505
R7300 VDD.n6001 VDD.n6000 3.1505
R7301 VDD.n5999 VDD.n5998 3.1505
R7302 VDD.n5998 VDD.n5997 3.1505
R7303 VDD.n5996 VDD.n5995 3.1505
R7304 VDD.n5995 VDD.n5994 3.1505
R7305 VDD.n5993 VDD.n5992 3.1505
R7306 VDD.n5992 VDD.n5991 3.1505
R7307 VDD.n5989 VDD.n5988 3.1505
R7308 VDD.n5988 VDD.n5987 3.1505
R7309 VDD.n5986 VDD.n5985 3.1505
R7310 VDD.n5985 VDD.n5984 3.1505
R7311 VDD.n5982 VDD.n5981 3.1505
R7312 VDD.n5981 VDD.n5980 3.1505
R7313 VDD.n5979 VDD.n5978 3.1505
R7314 VDD.n5978 VDD.n5977 3.1505
R7315 VDD.n5976 VDD.n5975 3.1505
R7316 VDD.n5975 VDD.n5974 3.1505
R7317 VDD.n5972 VDD.n5971 3.1505
R7318 VDD.n5971 VDD.n5970 3.1505
R7319 VDD.n5969 VDD.n5968 3.1505
R7320 VDD.n5968 VDD.n5967 3.1505
R7321 VDD.n5966 VDD.n5965 3.1505
R7322 VDD.n5965 VDD.n5964 3.1505
R7323 VDD.n5962 VDD.n5961 3.1505
R7324 VDD.n5961 VDD.n5960 3.1505
R7325 VDD.n5959 VDD.n5958 3.1505
R7326 VDD.n5958 VDD.n5957 3.1505
R7327 VDD.n5956 VDD.n5955 3.1505
R7328 VDD.n5955 VDD.n5954 3.1505
R7329 VDD.n5952 VDD.n5951 3.1505
R7330 VDD.n5951 VDD.n5950 3.1505
R7331 VDD.n5949 VDD.n5948 3.1505
R7332 VDD.n5948 VDD.n5947 3.1505
R7333 VDD.n5946 VDD.n5945 3.1505
R7334 VDD.n5945 VDD.n5944 3.1505
R7335 VDD.n5943 VDD.n5942 3.1505
R7336 VDD.n5942 VDD.n5941 3.1505
R7337 VDD.n5939 VDD.n5938 3.1505
R7338 VDD.n5938 VDD.n5937 3.1505
R7339 VDD.n5936 VDD.n5935 3.1505
R7340 VDD.n5935 VDD.n5934 3.1505
R7341 VDD.n5933 VDD.n5932 3.1505
R7342 VDD.n5932 VDD.n5931 3.1505
R7343 VDD.n5929 VDD.n5928 3.1505
R7344 VDD.n5928 VDD.n5927 3.1505
R7345 VDD.n5926 VDD.n5925 3.1505
R7346 VDD.n5925 VDD.n5924 3.1505
R7347 VDD.n5923 VDD.n5922 3.1505
R7348 VDD.n5922 VDD.n5921 3.1505
R7349 VDD.n5920 VDD.n5919 3.1505
R7350 VDD.n5919 VDD.n5918 3.1505
R7351 VDD.n5916 VDD.n5915 3.1505
R7352 VDD.n5915 VDD.n5914 3.1505
R7353 VDD.n5913 VDD.n5912 3.1505
R7354 VDD.n5912 VDD.n5911 3.1505
R7355 VDD.n5910 VDD.n5909 3.1505
R7356 VDD.n5909 VDD.n5908 3.1505
R7357 VDD.n5906 VDD.n5905 3.1505
R7358 VDD.n5905 VDD.n5904 3.1505
R7359 VDD.n5903 VDD.n5902 3.1505
R7360 VDD.n5902 VDD.n5901 3.1505
R7361 VDD.n5900 VDD.n5899 3.1505
R7362 VDD.n5899 VDD.n5898 3.1505
R7363 VDD.n5896 VDD.n5895 3.1505
R7364 VDD.n5895 VDD.n5894 3.1505
R7365 VDD.n5893 VDD.n5892 3.1505
R7366 VDD.n5892 VDD.n5891 3.1505
R7367 VDD.n5890 VDD.n5889 3.1505
R7368 VDD.n5889 VDD.n5888 3.1505
R7369 VDD.n5886 VDD.n5885 3.1505
R7370 VDD.n5885 VDD.n5884 3.1505
R7371 VDD.n5883 VDD.n5882 3.1505
R7372 VDD.n5882 VDD.n5881 3.1505
R7373 VDD.n5879 VDD.n5878 3.1505
R7374 VDD.n5878 VDD.n5877 3.1505
R7375 VDD.n5876 VDD.n5875 3.1505
R7376 VDD.n5875 VDD.n5874 3.1505
R7377 VDD.n5873 VDD.n5872 3.1505
R7378 VDD.n5872 VDD.n5871 3.1505
R7379 VDD.n5870 VDD.n5869 3.1505
R7380 VDD.n5869 VDD.n5868 3.1505
R7381 VDD.n5867 VDD.n5866 3.1505
R7382 VDD.n5866 VDD.n5865 3.1505
R7383 VDD.n5863 VDD.n5862 3.1505
R7384 VDD.n5857 VDD.n5856 3.1505
R7385 VDD.n5271 VDD.n5270 3.1505
R7386 VDD.n3254 VDD.n3253 3.1505
R7387 VDD.n5266 VDD.n5265 3.1505
R7388 VDD.n5263 VDD.n5262 3.1505
R7389 VDD.n5260 VDD.n5259 3.1505
R7390 VDD.n5257 VDD.n5256 3.1505
R7391 VDD.n5254 VDD.n5253 3.1505
R7392 VDD.n5251 VDD.n5250 3.1505
R7393 VDD.n5248 VDD.n5247 3.1505
R7394 VDD.n5245 VDD.n5244 3.1505
R7395 VDD.n5242 VDD.n5241 3.1505
R7396 VDD.n5239 VDD.n5238 3.1505
R7397 VDD.n5236 VDD.n5235 3.1505
R7398 VDD.n5233 VDD.n5232 3.1505
R7399 VDD.n5230 VDD.n5229 3.1505
R7400 VDD.n5227 VDD.n5226 3.1505
R7401 VDD.n5224 VDD.n5223 3.1505
R7402 VDD.n5221 VDD.n5220 3.1505
R7403 VDD.n5218 VDD.n5217 3.1505
R7404 VDD.n5215 VDD.n5214 3.1505
R7405 VDD.n5212 VDD.n5211 3.1505
R7406 VDD.n5209 VDD.n5208 3.1505
R7407 VDD.n5206 VDD.n5205 3.1505
R7408 VDD.n5203 VDD.n5202 3.1505
R7409 VDD.n5200 VDD.n5199 3.1505
R7410 VDD.n5197 VDD.n5196 3.1505
R7411 VDD.n5194 VDD.n5193 3.1505
R7412 VDD.n5191 VDD.n5190 3.1505
R7413 VDD.n5188 VDD.n5187 3.1505
R7414 VDD.n5185 VDD.n5184 3.1505
R7415 VDD.n5182 VDD.n5181 3.1505
R7416 VDD.n5179 VDD.n5178 3.1505
R7417 VDD.n5176 VDD.n5175 3.1505
R7418 VDD.n5173 VDD.n5172 3.1505
R7419 VDD.n5170 VDD.n5169 3.1505
R7420 VDD.n5167 VDD.n5166 3.1505
R7421 VDD.n5164 VDD.n5163 3.1505
R7422 VDD.n5161 VDD.n5160 3.1505
R7423 VDD.n5158 VDD.n5157 3.1505
R7424 VDD.n5155 VDD.n5154 3.1505
R7425 VDD.n5152 VDD.n5151 3.1505
R7426 VDD.n5149 VDD.n5148 3.1505
R7427 VDD.n5146 VDD.n5145 3.1505
R7428 VDD.n3243 VDD.n3242 3.1505
R7429 VDD.n3246 VDD.n3245 3.1505
R7430 VDD.n3249 VDD.n3248 3.1505
R7431 VDD.n3252 VDD.n3251 3.1505
R7432 VDD.n5268 VDD.n5267 3.1505
R7433 VDD.n5715 VDD.n5714 3.1505
R7434 VDD.n5715 VDD.n5711 3.1505
R7435 VDD.n5855 VDD.n5854 3.1505
R7436 VDD.n5854 VDD.n5853 3.1505
R7437 VDD.n5852 VDD.n5851 3.1505
R7438 VDD.n5851 VDD.n5850 3.1505
R7439 VDD.n5849 VDD.n5848 3.1505
R7440 VDD.n5848 VDD.n5847 3.1505
R7441 VDD.n5846 VDD.n5845 3.1505
R7442 VDD.n5845 VDD.n5844 3.1505
R7443 VDD.n5842 VDD.n5841 3.1505
R7444 VDD.n5841 VDD.n5840 3.1505
R7445 VDD.n5839 VDD.n5838 3.1505
R7446 VDD.n5838 VDD.n5837 3.1505
R7447 VDD.n5835 VDD.n5834 3.1505
R7448 VDD.n5834 VDD.n5833 3.1505
R7449 VDD.n5832 VDD.n5831 3.1505
R7450 VDD.n5831 VDD.n5830 3.1505
R7451 VDD.n5829 VDD.n5828 3.1505
R7452 VDD.n5828 VDD.n5827 3.1505
R7453 VDD.n5825 VDD.n5824 3.1505
R7454 VDD.n5824 VDD.n5823 3.1505
R7455 VDD.n5822 VDD.n5821 3.1505
R7456 VDD.n5821 VDD.n5820 3.1505
R7457 VDD.n5819 VDD.n5818 3.1505
R7458 VDD.n5818 VDD.n5817 3.1505
R7459 VDD.n5815 VDD.n5814 3.1505
R7460 VDD.n5814 VDD.n5813 3.1505
R7461 VDD.n5812 VDD.n5811 3.1505
R7462 VDD.n5811 VDD.n5810 3.1505
R7463 VDD.n5809 VDD.n5808 3.1505
R7464 VDD.n5808 VDD.n5807 3.1505
R7465 VDD.n5805 VDD.n5804 3.1505
R7466 VDD.n5804 VDD.n5803 3.1505
R7467 VDD.n5802 VDD.n5801 3.1505
R7468 VDD.n5801 VDD.n5800 3.1505
R7469 VDD.n5799 VDD.n5798 3.1505
R7470 VDD.n5798 VDD.n5797 3.1505
R7471 VDD.n5796 VDD.n5795 3.1505
R7472 VDD.n5795 VDD.n5794 3.1505
R7473 VDD.n5792 VDD.n5791 3.1505
R7474 VDD.n5791 VDD.n5790 3.1505
R7475 VDD.n5789 VDD.n5788 3.1505
R7476 VDD.n5788 VDD.n5787 3.1505
R7477 VDD.n5786 VDD.n5785 3.1505
R7478 VDD.n5785 VDD.n5784 3.1505
R7479 VDD.n5782 VDD.n5781 3.1505
R7480 VDD.n5781 VDD.n5780 3.1505
R7481 VDD.n5779 VDD.n5778 3.1505
R7482 VDD.n5778 VDD.n5777 3.1505
R7483 VDD.n5776 VDD.n5775 3.1505
R7484 VDD.n5775 VDD.n5774 3.1505
R7485 VDD.n5773 VDD.n5772 3.1505
R7486 VDD.n5772 VDD.n5771 3.1505
R7487 VDD.n5769 VDD.n5768 3.1505
R7488 VDD.n5768 VDD.n5767 3.1505
R7489 VDD.n5766 VDD.n5765 3.1505
R7490 VDD.n5765 VDD.n5764 3.1505
R7491 VDD.n5763 VDD.n5762 3.1505
R7492 VDD.n5762 VDD.n5761 3.1505
R7493 VDD.n5759 VDD.n5758 3.1505
R7494 VDD.n5758 VDD.n5757 3.1505
R7495 VDD.n5756 VDD.n5755 3.1505
R7496 VDD.n5755 VDD.n5754 3.1505
R7497 VDD.n5753 VDD.n5752 3.1505
R7498 VDD.n5752 VDD.n5751 3.1505
R7499 VDD.n5749 VDD.n5748 3.1505
R7500 VDD.n5748 VDD.n5747 3.1505
R7501 VDD.n5746 VDD.n5745 3.1505
R7502 VDD.n5745 VDD.n5744 3.1505
R7503 VDD.n5743 VDD.n5742 3.1505
R7504 VDD.n5742 VDD.n5741 3.1505
R7505 VDD.n5739 VDD.n5738 3.1505
R7506 VDD.n5738 VDD.n5737 3.1505
R7507 VDD.n5736 VDD.n5735 3.1505
R7508 VDD.n5735 VDD.n5734 3.1505
R7509 VDD.n5732 VDD.n5731 3.1505
R7510 VDD.n5731 VDD.n5730 3.1505
R7511 VDD.n5729 VDD.n5728 3.1505
R7512 VDD.n5728 VDD.n5727 3.1505
R7513 VDD.n5726 VDD.n5725 3.1505
R7514 VDD.n5725 VDD.n5724 3.1505
R7515 VDD.n5723 VDD.n5722 3.1505
R7516 VDD.n5722 VDD.n5721 3.1505
R7517 VDD.n5719 VDD.n5718 3.1505
R7518 VDD.n5718 VDD.n5717 3.1505
R7519 VDD.n5689 VDD.n5688 3.1505
R7520 VDD.n5688 VDD.n5687 3.1505
R7521 VDD.n5686 VDD.n5685 3.1505
R7522 VDD.n5685 VDD.n5684 3.1505
R7523 VDD.n5683 VDD.n5682 3.1505
R7524 VDD.n5682 VDD.n5681 3.1505
R7525 VDD.n5680 VDD.n5679 3.1505
R7526 VDD.n5679 VDD.n5678 3.1505
R7527 VDD.n5677 VDD.n5676 3.1505
R7528 VDD.n5676 VDD.n5675 3.1505
R7529 VDD.n5673 VDD.n5672 3.1505
R7530 VDD.n5672 VDD.n5671 3.1505
R7531 VDD.n5670 VDD.n5669 3.1505
R7532 VDD.n5669 VDD.n5668 3.1505
R7533 VDD.n5666 VDD.n5665 3.1505
R7534 VDD.n5665 VDD.n5664 3.1505
R7535 VDD.n5663 VDD.n5662 3.1505
R7536 VDD.n5662 VDD.n5661 3.1505
R7537 VDD.n5660 VDD.n5659 3.1505
R7538 VDD.n5659 VDD.n5658 3.1505
R7539 VDD.n5656 VDD.n5655 3.1505
R7540 VDD.n5655 VDD.n5654 3.1505
R7541 VDD.n5653 VDD.n5652 3.1505
R7542 VDD.n5652 VDD.n5651 3.1505
R7543 VDD.n5650 VDD.n5649 3.1505
R7544 VDD.n5649 VDD.n5648 3.1505
R7545 VDD.n5646 VDD.n5645 3.1505
R7546 VDD.n5645 VDD.n5644 3.1505
R7547 VDD.n5643 VDD.n5642 3.1505
R7548 VDD.n5642 VDD.n5641 3.1505
R7549 VDD.n5640 VDD.n5639 3.1505
R7550 VDD.n5639 VDD.n5638 3.1505
R7551 VDD.n5636 VDD.n5635 3.1505
R7552 VDD.n5635 VDD.n5634 3.1505
R7553 VDD.n5633 VDD.n5632 3.1505
R7554 VDD.n5632 VDD.n5631 3.1505
R7555 VDD.n5630 VDD.n5629 3.1505
R7556 VDD.n5629 VDD.n5628 3.1505
R7557 VDD.n5627 VDD.n5626 3.1505
R7558 VDD.n5626 VDD.n5625 3.1505
R7559 VDD.n5623 VDD.n5622 3.1505
R7560 VDD.n5622 VDD.n5621 3.1505
R7561 VDD.n5620 VDD.n5619 3.1505
R7562 VDD.n5619 VDD.n5618 3.1505
R7563 VDD.n5617 VDD.n5616 3.1505
R7564 VDD.n5616 VDD.n5615 3.1505
R7565 VDD.n5613 VDD.n5612 3.1505
R7566 VDD.n5612 VDD.n5611 3.1505
R7567 VDD.n5610 VDD.n5609 3.1505
R7568 VDD.n5609 VDD.n5608 3.1505
R7569 VDD.n5607 VDD.n5606 3.1505
R7570 VDD.n5606 VDD.n5605 3.1505
R7571 VDD.n5604 VDD.n5603 3.1505
R7572 VDD.n5603 VDD.n5602 3.1505
R7573 VDD.n5600 VDD.n5599 3.1505
R7574 VDD.n5599 VDD.n5598 3.1505
R7575 VDD.n5597 VDD.n5596 3.1505
R7576 VDD.n5596 VDD.n5595 3.1505
R7577 VDD.n5594 VDD.n5593 3.1505
R7578 VDD.n5593 VDD.n5592 3.1505
R7579 VDD.n5590 VDD.n5589 3.1505
R7580 VDD.n5589 VDD.n5588 3.1505
R7581 VDD.n5587 VDD.n5586 3.1505
R7582 VDD.n5586 VDD.n5585 3.1505
R7583 VDD.n5584 VDD.n5583 3.1505
R7584 VDD.n5583 VDD.n5582 3.1505
R7585 VDD.n5580 VDD.n5579 3.1505
R7586 VDD.n5579 VDD.n5578 3.1505
R7587 VDD.n5577 VDD.n5576 3.1505
R7588 VDD.n5576 VDD.n5575 3.1505
R7589 VDD.n5574 VDD.n5573 3.1505
R7590 VDD.n5573 VDD.n5572 3.1505
R7591 VDD.n5570 VDD.n5569 3.1505
R7592 VDD.n5569 VDD.n5568 3.1505
R7593 VDD.n5567 VDD.n5566 3.1505
R7594 VDD.n5566 VDD.n5565 3.1505
R7595 VDD.n5560 VDD.n5559 3.1505
R7596 VDD.n5559 VDD.n5558 3.1505
R7597 VDD.n5557 VDD.n5556 3.1505
R7598 VDD.n5556 VDD.n5555 3.1505
R7599 VDD.n5554 VDD.n5553 3.1505
R7600 VDD.n5553 VDD.n5552 3.1505
R7601 VDD.n5551 VDD.n5550 3.1505
R7602 VDD.n5550 VDD.n5549 3.1505
R7603 VDD.n5548 VDD.n5547 3.1505
R7604 VDD.n5547 VDD.n5546 3.1505
R7605 VDD.n5543 VDD.n5542 3.1505
R7606 VDD.n3447 VDD.n3446 3.1505
R7607 VDD.n3449 VDD.n3448 3.1505
R7608 VDD.n3451 VDD.n3450 3.1505
R7609 VDD.n3453 VDD.n3452 3.1505
R7610 VDD.n3455 VDD.n3454 3.1505
R7611 VDD.n3458 VDD.n3457 3.1505
R7612 VDD.n3460 VDD.n3459 3.1505
R7613 VDD.n3463 VDD.n3462 3.1505
R7614 VDD.n3465 VDD.n3464 3.1505
R7615 VDD.n3467 VDD.n3466 3.1505
R7616 VDD.n3470 VDD.n3469 3.1505
R7617 VDD.n3472 VDD.n3471 3.1505
R7618 VDD.n3474 VDD.n3473 3.1505
R7619 VDD.n3477 VDD.n3476 3.1505
R7620 VDD.n3479 VDD.n3478 3.1505
R7621 VDD.n3481 VDD.n3480 3.1505
R7622 VDD.n3484 VDD.n3483 3.1505
R7623 VDD.n3486 VDD.n3485 3.1505
R7624 VDD.n3488 VDD.n3487 3.1505
R7625 VDD.n3490 VDD.n3489 3.1505
R7626 VDD.n3492 VDD.n3491 3.1505
R7627 VDD.n3494 VDD.n3493 3.1505
R7628 VDD.n3496 VDD.n3495 3.1505
R7629 VDD.n3498 VDD.n3497 3.1505
R7630 VDD.n3500 VDD.n3499 3.1505
R7631 VDD.n3502 VDD.n3501 3.1505
R7632 VDD.n3504 VDD.n3503 3.1505
R7633 VDD.n3507 VDD.n3506 3.1505
R7634 VDD.n3509 VDD.n3508 3.1505
R7635 VDD.n3511 VDD.n3510 3.1505
R7636 VDD.n3514 VDD.n3513 3.1505
R7637 VDD.n3516 VDD.n3515 3.1505
R7638 VDD.n3518 VDD.n3517 3.1505
R7639 VDD.n3521 VDD.n3520 3.1505
R7640 VDD.n3523 VDD.n3522 3.1505
R7641 VDD.n3525 VDD.n3524 3.1505
R7642 VDD.n3528 VDD.n3527 3.1505
R7643 VDD.n3530 VDD.n3529 3.1505
R7644 VDD.n3533 VDD.n3532 3.1505
R7645 VDD.n3535 VDD.n3534 3.1505
R7646 VDD.n3537 VDD.n3536 3.1505
R7647 VDD.n3539 VDD.n3538 3.1505
R7648 VDD.n3341 VDD.n3340 3.1505
R7649 VDD.n3343 VDD.n3342 3.1505
R7650 VDD.n3345 VDD.n3344 3.1505
R7651 VDD.n3347 VDD.n3346 3.1505
R7652 VDD.n3349 VDD.n3348 3.1505
R7653 VDD.n3352 VDD.n3351 3.1505
R7654 VDD.n3354 VDD.n3353 3.1505
R7655 VDD.n3357 VDD.n3356 3.1505
R7656 VDD.n3359 VDD.n3358 3.1505
R7657 VDD.n3361 VDD.n3360 3.1505
R7658 VDD.n3364 VDD.n3363 3.1505
R7659 VDD.n3366 VDD.n3365 3.1505
R7660 VDD.n3368 VDD.n3367 3.1505
R7661 VDD.n3371 VDD.n3370 3.1505
R7662 VDD.n3373 VDD.n3372 3.1505
R7663 VDD.n3375 VDD.n3374 3.1505
R7664 VDD.n3378 VDD.n3377 3.1505
R7665 VDD.n3380 VDD.n3379 3.1505
R7666 VDD.n3382 VDD.n3381 3.1505
R7667 VDD.n3384 VDD.n3383 3.1505
R7668 VDD.n3386 VDD.n3385 3.1505
R7669 VDD.n3388 VDD.n3387 3.1505
R7670 VDD.n3390 VDD.n3389 3.1505
R7671 VDD.n3392 VDD.n3391 3.1505
R7672 VDD.n3394 VDD.n3393 3.1505
R7673 VDD.n3396 VDD.n3395 3.1505
R7674 VDD.n3398 VDD.n3397 3.1505
R7675 VDD.n3401 VDD.n3400 3.1505
R7676 VDD.n3403 VDD.n3402 3.1505
R7677 VDD.n3405 VDD.n3404 3.1505
R7678 VDD.n3408 VDD.n3407 3.1505
R7679 VDD.n3410 VDD.n3409 3.1505
R7680 VDD.n3412 VDD.n3411 3.1505
R7681 VDD.n3415 VDD.n3414 3.1505
R7682 VDD.n3417 VDD.n3416 3.1505
R7683 VDD.n3419 VDD.n3418 3.1505
R7684 VDD.n3422 VDD.n3421 3.1505
R7685 VDD.n3424 VDD.n3423 3.1505
R7686 VDD.n3427 VDD.n3426 3.1505
R7687 VDD.n3429 VDD.n3428 3.1505
R7688 VDD.n3431 VDD.n3430 3.1505
R7689 VDD.n3433 VDD.n3432 3.1505
R7690 VDD.n3435 VDD.n3434 3.1505
R7691 VDD.n2836 VDD.n2835 3.1505
R7692 VDD.n2833 VDD.n2832 3.1505
R7693 VDD.n2830 VDD.n2829 3.1505
R7694 VDD.n2827 VDD.n2826 3.1505
R7695 VDD.n2824 VDD.n2823 3.1505
R7696 VDD.n2821 VDD.n2820 3.1505
R7697 VDD.n2818 VDD.n2817 3.1505
R7698 VDD.n2815 VDD.n2814 3.1505
R7699 VDD.n2812 VDD.n2811 3.1505
R7700 VDD.n2809 VDD.n2808 3.1505
R7701 VDD.n2806 VDD.n2805 3.1505
R7702 VDD.n2803 VDD.n2802 3.1505
R7703 VDD.n2800 VDD.n2799 3.1505
R7704 VDD.n2797 VDD.n2796 3.1505
R7705 VDD.n2794 VDD.n2793 3.1505
R7706 VDD.n2791 VDD.n2790 3.1505
R7707 VDD.n2788 VDD.n2787 3.1505
R7708 VDD.n2785 VDD.n2784 3.1505
R7709 VDD.n2782 VDD.n2781 3.1505
R7710 VDD.n2779 VDD.n2778 3.1505
R7711 VDD.n2776 VDD.n2775 3.1505
R7712 VDD.n2773 VDD.n2772 3.1505
R7713 VDD.n2770 VDD.n2769 3.1505
R7714 VDD.n2767 VDD.n2766 3.1505
R7715 VDD.n2764 VDD.n2763 3.1505
R7716 VDD.n2761 VDD.n2760 3.1505
R7717 VDD.n2758 VDD.n2757 3.1505
R7718 VDD.n2755 VDD.n2754 3.1505
R7719 VDD.n2752 VDD.n2751 3.1505
R7720 VDD.n2749 VDD.n2748 3.1505
R7721 VDD.n2746 VDD.n2745 3.1505
R7722 VDD.n2743 VDD.n2742 3.1505
R7723 VDD.n2740 VDD.n2739 3.1505
R7724 VDD.n2737 VDD.n2736 3.1505
R7725 VDD.n2734 VDD.n2733 3.1505
R7726 VDD.n2731 VDD.n2730 3.1505
R7727 VDD.n2728 VDD.n2727 3.1505
R7728 VDD.n2725 VDD.n2724 3.1505
R7729 VDD.n2722 VDD.n2721 3.1505
R7730 VDD.n2719 VDD.n2718 3.1505
R7731 VDD.n2716 VDD.n2715 3.1505
R7732 VDD.n2713 VDD.n2712 3.1505
R7733 VDD.n2710 VDD.n2709 3.1505
R7734 VDD.n2707 VDD.n2706 3.1505
R7735 VDD.n2704 VDD.n2703 3.1505
R7736 VDD.n2701 VDD.n2700 3.1505
R7737 VDD.n2698 VDD.n2697 3.1505
R7738 VDD.n2695 VDD.n2694 3.1505
R7739 VDD.n3954 VDD.n3953 3.1505
R7740 VDD.n3952 VDD.n3951 3.1505
R7741 VDD.n2596 VDD.n2595 3.1505
R7742 VDD.n2598 VDD.n2597 3.1505
R7743 VDD.n2601 VDD.n2600 3.1505
R7744 VDD.n2603 VDD.n2602 3.1505
R7745 VDD.n2606 VDD.n2605 3.1505
R7746 VDD.n2608 VDD.n2607 3.1505
R7747 VDD.n2610 VDD.n2609 3.1505
R7748 VDD.n2613 VDD.n2612 3.1505
R7749 VDD.n2615 VDD.n2614 3.1505
R7750 VDD.n2617 VDD.n2616 3.1505
R7751 VDD.n2620 VDD.n2619 3.1505
R7752 VDD.n2622 VDD.n2621 3.1505
R7753 VDD.n2624 VDD.n2623 3.1505
R7754 VDD.n2627 VDD.n2626 3.1505
R7755 VDD.n2629 VDD.n2628 3.1505
R7756 VDD.n2631 VDD.n2630 3.1505
R7757 VDD.n2633 VDD.n2632 3.1505
R7758 VDD.n2635 VDD.n2634 3.1505
R7759 VDD.n2637 VDD.n2636 3.1505
R7760 VDD.n2639 VDD.n2638 3.1505
R7761 VDD.n2641 VDD.n2640 3.1505
R7762 VDD.n2643 VDD.n2642 3.1505
R7763 VDD.n2645 VDD.n2644 3.1505
R7764 VDD.n2647 VDD.n2646 3.1505
R7765 VDD.n2650 VDD.n2649 3.1505
R7766 VDD.n2652 VDD.n2651 3.1505
R7767 VDD.n2654 VDD.n2653 3.1505
R7768 VDD.n2657 VDD.n2656 3.1505
R7769 VDD.n2659 VDD.n2658 3.1505
R7770 VDD.n2661 VDD.n2660 3.1505
R7771 VDD.n2664 VDD.n2663 3.1505
R7772 VDD.n2666 VDD.n2665 3.1505
R7773 VDD.n2668 VDD.n2667 3.1505
R7774 VDD.n2671 VDD.n2670 3.1505
R7775 VDD.n2673 VDD.n2672 3.1505
R7776 VDD.n2681 VDD.n2680 3.1505
R7777 VDD.n2683 VDD.n2682 3.1505
R7778 VDD.n2685 VDD.n2684 3.1505
R7779 VDD.n2687 VDD.n2686 3.1505
R7780 VDD.n2689 VDD.n2688 3.1505
R7781 VDD.n6626 VDD.n6622 3.1505
R7782 VDD.n6626 VDD.n6625 3.1505
R7783 VDD.n6621 VDD.n6620 3.1505
R7784 VDD.n6620 VDD.n6619 3.1505
R7785 VDD.n6618 VDD.n6617 3.1505
R7786 VDD.n6617 VDD.n6616 3.1505
R7787 VDD.n6615 VDD.n6614 3.1505
R7788 VDD.n6614 VDD.n6613 3.1505
R7789 VDD.n6612 VDD.n6611 3.1505
R7790 VDD.n6611 VDD.n6610 3.1505
R7791 VDD.n6609 VDD.n6608 3.1505
R7792 VDD.n6608 VDD.n6607 3.1505
R7793 VDD.n6605 VDD.n6604 3.1505
R7794 VDD.n6604 VDD.n6603 3.1505
R7795 VDD.n6602 VDD.n6601 3.1505
R7796 VDD.n6601 VDD.n6600 3.1505
R7797 VDD.n6598 VDD.n6597 3.1505
R7798 VDD.n6597 VDD.n6596 3.1505
R7799 VDD.n6595 VDD.n6594 3.1505
R7800 VDD.n6594 VDD.n6593 3.1505
R7801 VDD.n6592 VDD.n6591 3.1505
R7802 VDD.n6591 VDD.n6590 3.1505
R7803 VDD.n6588 VDD.n6587 3.1505
R7804 VDD.n6587 VDD.n6586 3.1505
R7805 VDD.n6585 VDD.n6584 3.1505
R7806 VDD.n6584 VDD.n6583 3.1505
R7807 VDD.n6582 VDD.n6581 3.1505
R7808 VDD.n6581 VDD.n6580 3.1505
R7809 VDD.n6578 VDD.n6577 3.1505
R7810 VDD.n6577 VDD.n6576 3.1505
R7811 VDD.n6575 VDD.n6574 3.1505
R7812 VDD.n6574 VDD.n6573 3.1505
R7813 VDD.n6572 VDD.n6571 3.1505
R7814 VDD.n6571 VDD.n6570 3.1505
R7815 VDD.n6568 VDD.n6567 3.1505
R7816 VDD.n6567 VDD.n6566 3.1505
R7817 VDD.n6565 VDD.n6564 3.1505
R7818 VDD.n6564 VDD.n6563 3.1505
R7819 VDD.n6562 VDD.n6561 3.1505
R7820 VDD.n6561 VDD.n6560 3.1505
R7821 VDD.n6559 VDD.n6558 3.1505
R7822 VDD.n6558 VDD.n6557 3.1505
R7823 VDD.n6555 VDD.n6554 3.1505
R7824 VDD.n6554 VDD.n6553 3.1505
R7825 VDD.n6552 VDD.n6551 3.1505
R7826 VDD.n6551 VDD.n6550 3.1505
R7827 VDD.n6549 VDD.n6548 3.1505
R7828 VDD.n6548 VDD.n6547 3.1505
R7829 VDD.n6545 VDD.n6544 3.1505
R7830 VDD.n6544 VDD.n6543 3.1505
R7831 VDD.n6542 VDD.n6541 3.1505
R7832 VDD.n6541 VDD.n6540 3.1505
R7833 VDD.n6539 VDD.n6538 3.1505
R7834 VDD.n6538 VDD.n6537 3.1505
R7835 VDD.n6536 VDD.n6535 3.1505
R7836 VDD.n6535 VDD.n6534 3.1505
R7837 VDD.n6532 VDD.n6531 3.1505
R7838 VDD.n6531 VDD.n6530 3.1505
R7839 VDD.n6529 VDD.n6528 3.1505
R7840 VDD.n6528 VDD.n6527 3.1505
R7841 VDD.n6526 VDD.n6525 3.1505
R7842 VDD.n6525 VDD.n6524 3.1505
R7843 VDD.n6522 VDD.n6521 3.1505
R7844 VDD.n6521 VDD.n6520 3.1505
R7845 VDD.n6519 VDD.n6518 3.1505
R7846 VDD.n6518 VDD.n6517 3.1505
R7847 VDD.n6516 VDD.n6515 3.1505
R7848 VDD.n6515 VDD.n6514 3.1505
R7849 VDD.n6512 VDD.n6511 3.1505
R7850 VDD.n6511 VDD.n6510 3.1505
R7851 VDD.n6509 VDD.n6508 3.1505
R7852 VDD.n6508 VDD.n6507 3.1505
R7853 VDD.n6506 VDD.n6505 3.1505
R7854 VDD.n6505 VDD.n6504 3.1505
R7855 VDD.n6502 VDD.n6501 3.1505
R7856 VDD.n6501 VDD.n6500 3.1505
R7857 VDD.n6499 VDD.n6498 3.1505
R7858 VDD.n6498 VDD.n6497 3.1505
R7859 VDD.n6495 VDD.n6494 3.1505
R7860 VDD.n6494 VDD.n6493 3.1505
R7861 VDD.n6492 VDD.n6491 3.1505
R7862 VDD.n6491 VDD.n6490 3.1505
R7863 VDD.n6489 VDD.n6488 3.1505
R7864 VDD.n6488 VDD.n6487 3.1505
R7865 VDD.n6486 VDD.n6485 3.1505
R7866 VDD.n6485 VDD.n6484 3.1505
R7867 VDD.n1797 VDD.n1796 3.1505
R7868 VDD.n1935 VDD.n1934 3.1505
R7869 VDD.n2039 VDD.n2038 3.1505
R7870 VDD.n1672 VDD.n1671 3.1505
R7871 VDD.n1674 VDD.n1673 3.1505
R7872 VDD.n1676 VDD.n1675 3.1505
R7873 VDD.n1678 VDD.n1677 3.1505
R7874 VDD.n1681 VDD.n1680 3.1505
R7875 VDD.n1684 VDD.n1683 3.1505
R7876 VDD.n1687 VDD.n1686 3.1505
R7877 VDD.n1690 VDD.n1689 3.1505
R7878 VDD.n1693 VDD.n1692 3.1505
R7879 VDD.n1696 VDD.n1695 3.1505
R7880 VDD.n1699 VDD.n1698 3.1505
R7881 VDD.n1702 VDD.n1701 3.1505
R7882 VDD.n1705 VDD.n1704 3.1505
R7883 VDD.n1708 VDD.n1707 3.1505
R7884 VDD.n1711 VDD.n1710 3.1505
R7885 VDD.n1714 VDD.n1713 3.1505
R7886 VDD.n1717 VDD.n1716 3.1505
R7887 VDD.n1720 VDD.n1719 3.1505
R7888 VDD.n1723 VDD.n1722 3.1505
R7889 VDD.n1726 VDD.n1725 3.1505
R7890 VDD.n1729 VDD.n1728 3.1505
R7891 VDD.n1732 VDD.n1731 3.1505
R7892 VDD.n1735 VDD.n1734 3.1505
R7893 VDD.n1738 VDD.n1737 3.1505
R7894 VDD.n1741 VDD.n1740 3.1505
R7895 VDD.n1744 VDD.n1743 3.1505
R7896 VDD.n1747 VDD.n1746 3.1505
R7897 VDD.n1750 VDD.n1749 3.1505
R7898 VDD.n1753 VDD.n1752 3.1505
R7899 VDD.n1756 VDD.n1755 3.1505
R7900 VDD.n1759 VDD.n1758 3.1505
R7901 VDD.n1762 VDD.n1761 3.1505
R7902 VDD.n1765 VDD.n1764 3.1505
R7903 VDD.n1768 VDD.n1767 3.1505
R7904 VDD.n1771 VDD.n1770 3.1505
R7905 VDD.n1774 VDD.n1773 3.1505
R7906 VDD.n1777 VDD.n1776 3.1505
R7907 VDD.n1780 VDD.n1779 3.1505
R7908 VDD.n1783 VDD.n1782 3.1505
R7909 VDD.n1786 VDD.n1785 3.1505
R7910 VDD.n1789 VDD.n1788 3.1505
R7911 VDD.n1792 VDD.n1791 3.1505
R7912 VDD.n1795 VDD.n1794 3.1505
R7913 VDD.n1669 VDD.n1668 3.1505
R7914 VDD.n1667 VDD.n1666 3.1505
R7915 VDD.n1810 VDD.n1809 3.1505
R7916 VDD.n1812 VDD.n1811 3.1505
R7917 VDD.n1814 VDD.n1813 3.1505
R7918 VDD.n1816 VDD.n1815 3.1505
R7919 VDD.n1819 VDD.n1818 3.1505
R7920 VDD.n1822 VDD.n1821 3.1505
R7921 VDD.n1825 VDD.n1824 3.1505
R7922 VDD.n1828 VDD.n1827 3.1505
R7923 VDD.n1831 VDD.n1830 3.1505
R7924 VDD.n1834 VDD.n1833 3.1505
R7925 VDD.n1837 VDD.n1836 3.1505
R7926 VDD.n1840 VDD.n1839 3.1505
R7927 VDD.n1843 VDD.n1842 3.1505
R7928 VDD.n1846 VDD.n1845 3.1505
R7929 VDD.n1849 VDD.n1848 3.1505
R7930 VDD.n1852 VDD.n1851 3.1505
R7931 VDD.n1855 VDD.n1854 3.1505
R7932 VDD.n1858 VDD.n1857 3.1505
R7933 VDD.n1861 VDD.n1860 3.1505
R7934 VDD.n1864 VDD.n1863 3.1505
R7935 VDD.n1867 VDD.n1866 3.1505
R7936 VDD.n1870 VDD.n1869 3.1505
R7937 VDD.n1873 VDD.n1872 3.1505
R7938 VDD.n1876 VDD.n1875 3.1505
R7939 VDD.n1879 VDD.n1878 3.1505
R7940 VDD.n1882 VDD.n1881 3.1505
R7941 VDD.n1885 VDD.n1884 3.1505
R7942 VDD.n1888 VDD.n1887 3.1505
R7943 VDD.n1891 VDD.n1890 3.1505
R7944 VDD.n1894 VDD.n1893 3.1505
R7945 VDD.n1897 VDD.n1896 3.1505
R7946 VDD.n1900 VDD.n1899 3.1505
R7947 VDD.n1903 VDD.n1902 3.1505
R7948 VDD.n1906 VDD.n1905 3.1505
R7949 VDD.n1909 VDD.n1908 3.1505
R7950 VDD.n1912 VDD.n1911 3.1505
R7951 VDD.n1915 VDD.n1914 3.1505
R7952 VDD.n1918 VDD.n1917 3.1505
R7953 VDD.n1921 VDD.n1920 3.1505
R7954 VDD.n1924 VDD.n1923 3.1505
R7955 VDD.n1927 VDD.n1926 3.1505
R7956 VDD.n1930 VDD.n1929 3.1505
R7957 VDD.n1933 VDD.n1932 3.1505
R7958 VDD.n1807 VDD.n1806 3.1505
R7959 VDD.n1805 VDD.n1804 3.1505
R7960 VDD.n2037 VDD.n2036 3.1505
R7961 VDD.n2034 VDD.n2033 3.1505
R7962 VDD.n2032 VDD.n2031 3.1505
R7963 VDD.n2029 VDD.n2028 3.1505
R7964 VDD.n2027 VDD.n2026 3.1505
R7965 VDD.n2024 VDD.n2023 3.1505
R7966 VDD.n2022 VDD.n2021 3.1505
R7967 VDD.n2019 VDD.n2018 3.1505
R7968 VDD.n2017 VDD.n2016 3.1505
R7969 VDD.n2014 VDD.n2013 3.1505
R7970 VDD.n2012 VDD.n2011 3.1505
R7971 VDD.n2009 VDD.n2008 3.1505
R7972 VDD.n2007 VDD.n2006 3.1505
R7973 VDD.n2004 VDD.n2003 3.1505
R7974 VDD.n2002 VDD.n2001 3.1505
R7975 VDD.n1999 VDD.n1998 3.1505
R7976 VDD.n1997 VDD.n1996 3.1505
R7977 VDD.n1994 VDD.n1993 3.1505
R7978 VDD.n1992 VDD.n1991 3.1505
R7979 VDD.n1989 VDD.n1988 3.1505
R7980 VDD.n1987 VDD.n1986 3.1505
R7981 VDD.n1985 VDD.n1984 3.1505
R7982 VDD.n1983 VDD.n1982 3.1505
R7983 VDD.n1981 VDD.n1980 3.1505
R7984 VDD.n1979 VDD.n1978 3.1505
R7985 VDD.n1977 VDD.n1976 3.1505
R7986 VDD.n1975 VDD.n1974 3.1505
R7987 VDD.n1973 VDD.n1972 3.1505
R7988 VDD.n1971 VDD.n1970 3.1505
R7989 VDD.n1969 VDD.n1968 3.1505
R7990 VDD.n1967 VDD.n1966 3.1505
R7991 VDD.n1965 VDD.n1964 3.1505
R7992 VDD.n1963 VDD.n1962 3.1505
R7993 VDD.n1961 VDD.n1960 3.1505
R7994 VDD.n1959 VDD.n1958 3.1505
R7995 VDD.n1957 VDD.n1956 3.1505
R7996 VDD.n1955 VDD.n1954 3.1505
R7997 VDD.n1953 VDD.n1952 3.1505
R7998 VDD.n1951 VDD.n1950 3.1505
R7999 VDD.n1949 VDD.n1948 3.1505
R8000 VDD.n1947 VDD.n1946 3.1505
R8001 VDD.n1945 VDD.n1944 3.1505
R8002 VDD.n1943 VDD.n1942 3.1505
R8003 VDD.n1941 VDD.n1940 3.1505
R8004 VDD.n1939 VDD.n1938 3.1505
R8005 VDD.n1351 VDD.n1105 3.1505
R8006 VDD.n1252 VDD.n1251 3.1505
R8007 VDD.n1347 VDD.n1346 3.1505
R8008 VDD.n1345 VDD.n1344 3.1505
R8009 VDD.n1342 VDD.n1341 3.1505
R8010 VDD.n1340 VDD.n1339 3.1505
R8011 VDD.n1337 VDD.n1336 3.1505
R8012 VDD.n1335 VDD.n1334 3.1505
R8013 VDD.n1332 VDD.n1331 3.1505
R8014 VDD.n1330 VDD.n1329 3.1505
R8015 VDD.n1327 VDD.n1326 3.1505
R8016 VDD.n1325 VDD.n1324 3.1505
R8017 VDD.n1322 VDD.n1321 3.1505
R8018 VDD.n1320 VDD.n1319 3.1505
R8019 VDD.n1317 VDD.n1316 3.1505
R8020 VDD.n1315 VDD.n1314 3.1505
R8021 VDD.n1312 VDD.n1311 3.1505
R8022 VDD.n1310 VDD.n1309 3.1505
R8023 VDD.n1307 VDD.n1306 3.1505
R8024 VDD.n1305 VDD.n1304 3.1505
R8025 VDD.n1302 VDD.n1301 3.1505
R8026 VDD.n1300 VDD.n1299 3.1505
R8027 VDD.n1298 VDD.n1297 3.1505
R8028 VDD.n1296 VDD.n1295 3.1505
R8029 VDD.n1294 VDD.n1293 3.1505
R8030 VDD.n1292 VDD.n1291 3.1505
R8031 VDD.n1290 VDD.n1289 3.1505
R8032 VDD.n1288 VDD.n1287 3.1505
R8033 VDD.n1286 VDD.n1285 3.1505
R8034 VDD.n1284 VDD.n1283 3.1505
R8035 VDD.n1282 VDD.n1281 3.1505
R8036 VDD.n1280 VDD.n1279 3.1505
R8037 VDD.n1278 VDD.n1277 3.1505
R8038 VDD.n1276 VDD.n1275 3.1505
R8039 VDD.n1274 VDD.n1273 3.1505
R8040 VDD.n1272 VDD.n1271 3.1505
R8041 VDD.n1270 VDD.n1269 3.1505
R8042 VDD.n1268 VDD.n1267 3.1505
R8043 VDD.n1266 VDD.n1265 3.1505
R8044 VDD.n1264 VDD.n1263 3.1505
R8045 VDD.n1262 VDD.n1261 3.1505
R8046 VDD.n1260 VDD.n1259 3.1505
R8047 VDD.n1258 VDD.n1257 3.1505
R8048 VDD.n1256 VDD.n1255 3.1505
R8049 VDD.n1254 VDD.n1253 3.1505
R8050 VDD.n1350 VDD.n1349 3.1505
R8051 VDD.n1470 VDD.n1469 3.1505
R8052 VDD.n1472 VDD.n1471 3.1505
R8053 VDD.n1474 VDD.n1473 3.1505
R8054 VDD.n1476 VDD.n1475 3.1505
R8055 VDD.n1478 VDD.n1477 3.1505
R8056 VDD.n1480 VDD.n1479 3.1505
R8057 VDD.n1483 VDD.n1482 3.1505
R8058 VDD.n1485 VDD.n1484 3.1505
R8059 VDD.n1487 VDD.n1486 3.1505
R8060 VDD.n1489 VDD.n1488 3.1505
R8061 VDD.n1491 VDD.n1490 3.1505
R8062 VDD.n1493 VDD.n1492 3.1505
R8063 VDD.n1495 VDD.n1494 3.1505
R8064 VDD.n1497 VDD.n1496 3.1505
R8065 VDD.n1499 VDD.n1498 3.1505
R8066 VDD.n1501 VDD.n1500 3.1505
R8067 VDD.n1503 VDD.n1502 3.1505
R8068 VDD.n1505 VDD.n1504 3.1505
R8069 VDD.n1507 VDD.n1506 3.1505
R8070 VDD.n1509 VDD.n1508 3.1505
R8071 VDD.n1511 VDD.n1510 3.1505
R8072 VDD.n1513 VDD.n1512 3.1505
R8073 VDD.n1515 VDD.n1514 3.1505
R8074 VDD.n1517 VDD.n1516 3.1505
R8075 VDD.n1519 VDD.n1518 3.1505
R8076 VDD.n1522 VDD.n1521 3.1505
R8077 VDD.n1524 VDD.n1523 3.1505
R8078 VDD.n1526 VDD.n1525 3.1505
R8079 VDD.n1528 VDD.n1527 3.1505
R8080 VDD.n1530 VDD.n1529 3.1505
R8081 VDD.n1532 VDD.n1531 3.1505
R8082 VDD.n1539 VDD.n1538 3.1505
R8083 VDD.n1541 VDD.n1540 3.1505
R8084 VDD.n1543 VDD.n1542 3.1505
R8085 VDD.n1545 VDD.n1544 3.1505
R8086 VDD.n1547 VDD.n1546 3.1505
R8087 VDD.n1549 VDD.n1548 3.1505
R8088 VDD.n1551 VDD.n1550 3.1505
R8089 VDD.n1555 VDD.n1554 3.1505
R8090 VDD.n1557 VDD.n1556 3.1505
R8091 VDD.n1559 VDD.n1558 3.1505
R8092 VDD.n1561 VDD.n1560 3.1505
R8093 VDD.n1563 VDD.n1562 3.1505
R8094 VDD.n1565 VDD.n1564 3.1505
R8095 VDD.n1567 VDD.n1566 3.1505
R8096 VDD.n1569 VDD.n1568 3.1505
R8097 VDD.n1571 VDD.n1570 3.1505
R8098 VDD.n1573 VDD.n1572 3.1505
R8099 VDD.n1575 VDD.n1574 3.1505
R8100 VDD.n1577 VDD.n1576 3.1505
R8101 VDD.n1579 VDD.n1578 3.1505
R8102 VDD.n1581 VDD.n1580 3.1505
R8103 VDD.n1583 VDD.n1582 3.1505
R8104 VDD.n1585 VDD.n1584 3.1505
R8105 VDD.n1587 VDD.n1586 3.1505
R8106 VDD.n1589 VDD.n1588 3.1505
R8107 VDD.n1591 VDD.n1590 3.1505
R8108 VDD.n1593 VDD.n1592 3.1505
R8109 VDD.n1595 VDD.n1594 3.1505
R8110 VDD.n1597 VDD.n1596 3.1505
R8111 VDD.n1599 VDD.n1598 3.1505
R8112 VDD.n1601 VDD.n1600 3.1505
R8113 VDD.n1603 VDD.n1602 3.1505
R8114 VDD.n1605 VDD.n1604 3.1505
R8115 VDD.n1607 VDD.n1606 3.1505
R8116 VDD.n1609 VDD.n1608 3.1505
R8117 VDD.n1611 VDD.n1610 3.1505
R8118 VDD.n1613 VDD.n1612 3.1505
R8119 VDD.n1615 VDD.n1614 3.1505
R8120 VDD.n1617 VDD.n1616 3.1505
R8121 VDD.n1619 VDD.n1618 3.1505
R8122 VDD.n1621 VDD.n1620 3.1505
R8123 VDD.n1623 VDD.n1622 3.1505
R8124 VDD.n1625 VDD.n1624 3.1505
R8125 VDD.n1627 VDD.n1626 3.1505
R8126 VDD.n1629 VDD.n1628 3.1505
R8127 VDD.n1631 VDD.n1630 3.1505
R8128 VDD.n1633 VDD.n1632 3.1505
R8129 VDD.n1635 VDD.n1634 3.1505
R8130 VDD.n1637 VDD.n1636 3.1505
R8131 VDD.n1639 VDD.n1638 3.1505
R8132 VDD.n1641 VDD.n1640 3.1505
R8133 VDD.n1643 VDD.n1642 3.1505
R8134 VDD.n1645 VDD.n1644 3.1505
R8135 VDD.n1648 VDD.n1647 3.1505
R8136 VDD.n1650 VDD.n1649 3.1505
R8137 VDD.n1652 VDD.n1651 3.1505
R8138 VDD.n1654 VDD.n1653 3.1505
R8139 VDD.n1656 VDD.n1655 3.1505
R8140 VDD.n1658 VDD.n1657 3.1505
R8141 VDD.n1660 VDD.n1659 3.1505
R8142 VDD.n1141 VDD.n1140 3.1505
R8143 VDD.n1143 VDD.n1142 3.1505
R8144 VDD.n1145 VDD.n1144 3.1505
R8145 VDD.n1147 VDD.n1146 3.1505
R8146 VDD.n1149 VDD.n1148 3.1505
R8147 VDD.n1151 VDD.n1150 3.1505
R8148 VDD.n1154 VDD.n1153 3.1505
R8149 VDD.n1157 VDD.n1156 3.1505
R8150 VDD.n1159 VDD.n1158 3.1505
R8151 VDD.n1162 VDD.n1161 3.1505
R8152 VDD.n1164 VDD.n1163 3.1505
R8153 VDD.n1166 VDD.n1165 3.1505
R8154 VDD.n1168 VDD.n1167 3.1505
R8155 VDD.n1170 VDD.n1169 3.1505
R8156 VDD.n1172 VDD.n1171 3.1505
R8157 VDD.n1175 VDD.n1174 3.1505
R8158 VDD.n1177 VDD.n1176 3.1505
R8159 VDD.n1179 VDD.n1178 3.1505
R8160 VDD.n1181 VDD.n1180 3.1505
R8161 VDD.n1184 VDD.n1183 3.1505
R8162 VDD.n1186 VDD.n1185 3.1505
R8163 VDD.n1188 VDD.n1187 3.1505
R8164 VDD.n1190 VDD.n1189 3.1505
R8165 VDD.n1192 VDD.n1191 3.1505
R8166 VDD.n1194 VDD.n1193 3.1505
R8167 VDD.n1196 VDD.n1195 3.1505
R8168 VDD.n1198 VDD.n1197 3.1505
R8169 VDD.n1200 VDD.n1199 3.1505
R8170 VDD.n1202 VDD.n1201 3.1505
R8171 VDD.n1204 VDD.n1203 3.1505
R8172 VDD.n1206 VDD.n1205 3.1505
R8173 VDD.n1208 VDD.n1207 3.1505
R8174 VDD.n1210 VDD.n1209 3.1505
R8175 VDD.n1212 VDD.n1211 3.1505
R8176 VDD.n1214 VDD.n1213 3.1505
R8177 VDD.n1216 VDD.n1215 3.1505
R8178 VDD.n1218 VDD.n1217 3.1505
R8179 VDD.n1220 VDD.n1219 3.1505
R8180 VDD.n1222 VDD.n1221 3.1505
R8181 VDD.n1224 VDD.n1223 3.1505
R8182 VDD.n1226 VDD.n1225 3.1505
R8183 VDD.n1228 VDD.n1227 3.1505
R8184 VDD.n1230 VDD.n1229 3.1505
R8185 VDD.n1233 VDD.n1232 3.1505
R8186 VDD.n1236 VDD.n1235 3.1505
R8187 VDD.n1238 VDD.n1237 3.1505
R8188 VDD.n1240 VDD.n1239 3.1505
R8189 VDD.n1242 VDD.n1241 3.1505
R8190 VDD.n1244 VDD.n1243 3.1505
R8191 VDD.n1246 VDD.n1245 3.1505
R8192 VDD.n2059 VDD.n2058 3.1505
R8193 VDD.n2058 VDD.n2057 3.1505
R8194 VDD.n2062 VDD.n2061 3.1505
R8195 VDD.n2061 VDD.n2060 3.1505
R8196 VDD.n2065 VDD.n2064 3.1505
R8197 VDD.n2064 VDD.n2063 3.1505
R8198 VDD.n2068 VDD.n2067 3.1505
R8199 VDD.n2067 VDD.n2066 3.1505
R8200 VDD.n2071 VDD.n2070 3.1505
R8201 VDD.n2070 VDD.n2069 3.1505
R8202 VDD.n2074 VDD.n2073 3.1505
R8203 VDD.n2073 VDD.n2072 3.1505
R8204 VDD.n2078 VDD.n2077 3.1505
R8205 VDD.n2077 VDD.n2076 3.1505
R8206 VDD.n2081 VDD.n2080 3.1505
R8207 VDD.n2080 VDD.n2079 3.1505
R8208 VDD.n2084 VDD.n2083 3.1505
R8209 VDD.n2083 VDD.n2082 3.1505
R8210 VDD.n2087 VDD.n2086 3.1505
R8211 VDD.n2086 VDD.n2085 3.1505
R8212 VDD.n2090 VDD.n2089 3.1505
R8213 VDD.n2089 VDD.n2088 3.1505
R8214 VDD.n2093 VDD.n2092 3.1505
R8215 VDD.n2092 VDD.n2091 3.1505
R8216 VDD.n2096 VDD.n2095 3.1505
R8217 VDD.n2095 VDD.n2094 3.1505
R8218 VDD.n2099 VDD.n2098 3.1505
R8219 VDD.n2098 VDD.n2097 3.1505
R8220 VDD.n2102 VDD.n2101 3.1505
R8221 VDD.n2101 VDD.n2100 3.1505
R8222 VDD.n2105 VDD.n2104 3.1505
R8223 VDD.n2104 VDD.n2103 3.1505
R8224 VDD.n2108 VDD.n2107 3.1505
R8225 VDD.n2107 VDD.n2106 3.1505
R8226 VDD.n2111 VDD.n2110 3.1505
R8227 VDD.n2110 VDD.n2109 3.1505
R8228 VDD.n2114 VDD.n2113 3.1505
R8229 VDD.n2113 VDD.n2112 3.1505
R8230 VDD.n2117 VDD.n2116 3.1505
R8231 VDD.n2116 VDD.n2115 3.1505
R8232 VDD.n2120 VDD.n2119 3.1505
R8233 VDD.n2119 VDD.n2118 3.1505
R8234 VDD.n2123 VDD.n2122 3.1505
R8235 VDD.n2122 VDD.n2121 3.1505
R8236 VDD.n2126 VDD.n2125 3.1505
R8237 VDD.n2125 VDD.n2124 3.1505
R8238 VDD.n2129 VDD.n2128 3.1505
R8239 VDD.n2128 VDD.n2127 3.1505
R8240 VDD.n2132 VDD.n2131 3.1505
R8241 VDD.n2131 VDD.n2130 3.1505
R8242 VDD.n2136 VDD.n2135 3.1505
R8243 VDD.n2135 VDD.n2134 3.1505
R8244 VDD.n2139 VDD.n2138 3.1505
R8245 VDD.n2138 VDD.n2137 3.1505
R8246 VDD.n2142 VDD.n2141 3.1505
R8247 VDD.n2141 VDD.n2140 3.1505
R8248 VDD.n2145 VDD.n2144 3.1505
R8249 VDD.n2144 VDD.n2143 3.1505
R8250 VDD.n2148 VDD.n2147 3.1505
R8251 VDD.n2147 VDD.n2146 3.1505
R8252 VDD.n2151 VDD.n2150 3.1505
R8253 VDD.n2150 VDD.n2149 3.1505
R8254 VDD.n2163 VDD.n2162 3.1505
R8255 VDD.n2162 VDD.n2161 3.1505
R8256 VDD.n2166 VDD.n2165 3.1505
R8257 VDD.n2165 VDD.n2164 3.1505
R8258 VDD.n2169 VDD.n2168 3.1505
R8259 VDD.n2168 VDD.n2167 3.1505
R8260 VDD.n2172 VDD.n2171 3.1505
R8261 VDD.n2171 VDD.n2170 3.1505
R8262 VDD.n2175 VDD.n2174 3.1505
R8263 VDD.n2174 VDD.n2173 3.1505
R8264 VDD.n2178 VDD.n2177 3.1505
R8265 VDD.n2177 VDD.n2176 3.1505
R8266 VDD.n2181 VDD.n2180 3.1505
R8267 VDD.n2180 VDD.n2179 3.1505
R8268 VDD.n2185 VDD.n2184 3.1505
R8269 VDD.n2184 VDD.n2183 3.1505
R8270 VDD.n2188 VDD.n2187 3.1505
R8271 VDD.n2187 VDD.n2186 3.1505
R8272 VDD.n2191 VDD.n2190 3.1505
R8273 VDD.n2190 VDD.n2189 3.1505
R8274 VDD.n2194 VDD.n2193 3.1505
R8275 VDD.n2193 VDD.n2192 3.1505
R8276 VDD.n2197 VDD.n2196 3.1505
R8277 VDD.n2196 VDD.n2195 3.1505
R8278 VDD.n2200 VDD.n2199 3.1505
R8279 VDD.n2199 VDD.n2198 3.1505
R8280 VDD.n2203 VDD.n2202 3.1505
R8281 VDD.n2202 VDD.n2201 3.1505
R8282 VDD.n2206 VDD.n2205 3.1505
R8283 VDD.n2205 VDD.n2204 3.1505
R8284 VDD.n2209 VDD.n2208 3.1505
R8285 VDD.n2208 VDD.n2207 3.1505
R8286 VDD.n2212 VDD.n2211 3.1505
R8287 VDD.n2211 VDD.n2210 3.1505
R8288 VDD.n2215 VDD.n2214 3.1505
R8289 VDD.n2214 VDD.n2213 3.1505
R8290 VDD.n2218 VDD.n2217 3.1505
R8291 VDD.n2217 VDD.n2216 3.1505
R8292 VDD.n2221 VDD.n2220 3.1505
R8293 VDD.n2220 VDD.n2219 3.1505
R8294 VDD.n2224 VDD.n2223 3.1505
R8295 VDD.n2223 VDD.n2222 3.1505
R8296 VDD.n2227 VDD.n2226 3.1505
R8297 VDD.n2226 VDD.n2225 3.1505
R8298 VDD.n2230 VDD.n2229 3.1505
R8299 VDD.n2229 VDD.n2228 3.1505
R8300 VDD.n2233 VDD.n2232 3.1505
R8301 VDD.n2232 VDD.n2231 3.1505
R8302 VDD.n2236 VDD.n2235 3.1505
R8303 VDD.n2235 VDD.n2234 3.1505
R8304 VDD.n2239 VDD.n2238 3.1505
R8305 VDD.n2238 VDD.n2237 3.1505
R8306 VDD.n2242 VDD.n2241 3.1505
R8307 VDD.n2241 VDD.n2240 3.1505
R8308 VDD.n2245 VDD.n2244 3.1505
R8309 VDD.n2244 VDD.n2243 3.1505
R8310 VDD.n2248 VDD.n2247 3.1505
R8311 VDD.n2247 VDD.n2246 3.1505
R8312 VDD.n2251 VDD.n2250 3.1505
R8313 VDD.n2250 VDD.n2249 3.1505
R8314 VDD.n2254 VDD.n2253 3.1505
R8315 VDD.n2253 VDD.n2252 3.1505
R8316 VDD.n2257 VDD.n2256 3.1505
R8317 VDD.n2256 VDD.n2255 3.1505
R8318 VDD.n2260 VDD.n2259 3.1505
R8319 VDD.n2259 VDD.n2258 3.1505
R8320 VDD.n2263 VDD.n2262 3.1505
R8321 VDD.n2262 VDD.n2261 3.1505
R8322 VDD.n2266 VDD.n2265 3.1505
R8323 VDD.n2265 VDD.n2264 3.1505
R8324 VDD.n2269 VDD.n2268 3.1505
R8325 VDD.n2268 VDD.n2267 3.1505
R8326 VDD.n2272 VDD.n2271 3.1505
R8327 VDD.n2271 VDD.n2270 3.1505
R8328 VDD.n2275 VDD.n2274 3.1505
R8329 VDD.n2274 VDD.n2273 3.1505
R8330 VDD.n2278 VDD.n2277 3.1505
R8331 VDD.n2277 VDD.n2276 3.1505
R8332 VDD.n2281 VDD.n2280 3.1505
R8333 VDD.n2280 VDD.n2279 3.1505
R8334 VDD.n2284 VDD.n2283 3.1505
R8335 VDD.n2283 VDD.n2282 3.1505
R8336 VDD.n2287 VDD.n2286 3.1505
R8337 VDD.n2286 VDD.n2285 3.1505
R8338 VDD.n2290 VDD.n2289 3.1505
R8339 VDD.n2289 VDD.n2288 3.1505
R8340 VDD.n2293 VDD.n2292 3.1505
R8341 VDD.n2292 VDD.n2291 3.1505
R8342 VDD.n2296 VDD.n2295 3.1505
R8343 VDD.n2295 VDD.n2294 3.1505
R8344 VDD.n2299 VDD.n2298 3.1505
R8345 VDD.n2298 VDD.n2297 3.1505
R8346 VDD.n2302 VDD.n2301 3.1505
R8347 VDD.n2301 VDD.n2300 3.1505
R8348 VDD.n2305 VDD.n2304 3.1505
R8349 VDD.n2304 VDD.n2303 3.1505
R8350 VDD.n2308 VDD.n2307 3.1505
R8351 VDD.n2307 VDD.n2306 3.1505
R8352 VDD.n2311 VDD.n2310 3.1505
R8353 VDD.n2310 VDD.n2309 3.1505
R8354 VDD.n2314 VDD.n2313 3.1505
R8355 VDD.n2313 VDD.n2312 3.1505
R8356 VDD.n2317 VDD.n2316 3.1505
R8357 VDD.n2316 VDD.n2315 3.1505
R8358 VDD.n2320 VDD.n2319 3.1505
R8359 VDD.n2319 VDD.n2318 3.1505
R8360 VDD.n2324 VDD.n2323 3.1505
R8361 VDD.n2323 VDD.n2322 3.1505
R8362 VDD.n2327 VDD.n2326 3.1505
R8363 VDD.n2326 VDD.n2325 3.1505
R8364 VDD.n2330 VDD.n2329 3.1505
R8365 VDD.n2329 VDD.n2328 3.1505
R8366 VDD.n2333 VDD.n2332 3.1505
R8367 VDD.n2332 VDD.n2331 3.1505
R8368 VDD.n2336 VDD.n2335 3.1505
R8369 VDD.n2335 VDD.n2334 3.1505
R8370 VDD.n2339 VDD.n2338 3.1505
R8371 VDD.n2338 VDD.n2337 3.1505
R8372 VDD.n2342 VDD.n2341 3.1505
R8373 VDD.n2341 VDD.n2340 3.1505
R8374 VDD.n2354 VDD.n2353 3.1505
R8375 VDD.n2353 VDD.n2352 3.1505
R8376 VDD.n2357 VDD.n2356 3.1505
R8377 VDD.n2356 VDD.n2355 3.1505
R8378 VDD.n2360 VDD.n2359 3.1505
R8379 VDD.n2359 VDD.n2358 3.1505
R8380 VDD.n2363 VDD.n2362 3.1505
R8381 VDD.n2362 VDD.n2361 3.1505
R8382 VDD.n2366 VDD.n2365 3.1505
R8383 VDD.n2365 VDD.n2364 3.1505
R8384 VDD.n2369 VDD.n2368 3.1505
R8385 VDD.n2368 VDD.n2367 3.1505
R8386 VDD.n2373 VDD.n2372 3.1505
R8387 VDD.n2372 VDD.n2371 3.1505
R8388 VDD.n2377 VDD.n2376 3.1505
R8389 VDD.n2376 VDD.n2375 3.1505
R8390 VDD.n2381 VDD.n2380 3.1505
R8391 VDD.n2380 VDD.n2379 3.1505
R8392 VDD.n2385 VDD.n2384 3.1505
R8393 VDD.n2384 VDD.n2383 3.1505
R8394 VDD.n2388 VDD.n2387 3.1505
R8395 VDD.n2387 VDD.n2386 3.1505
R8396 VDD.n2392 VDD.n2391 3.1505
R8397 VDD.n2391 VDD.n2390 3.1505
R8398 VDD.n2396 VDD.n2395 3.1505
R8399 VDD.n2395 VDD.n2394 3.1505
R8400 VDD.n2400 VDD.n2399 3.1505
R8401 VDD.n2399 VDD.n2398 3.1505
R8402 VDD.n2403 VDD.n2402 3.1505
R8403 VDD.n2402 VDD.n2401 3.1505
R8404 VDD.n2407 VDD.n2406 3.1505
R8405 VDD.n2406 VDD.n2405 3.1505
R8406 VDD.n2410 VDD.n2409 3.1505
R8407 VDD.n2409 VDD.n2408 3.1505
R8408 VDD.n2413 VDD.n2412 3.1505
R8409 VDD.n2412 VDD.n2411 3.1505
R8410 VDD.n2416 VDD.n2415 3.1505
R8411 VDD.n2415 VDD.n2414 3.1505
R8412 VDD.n2421 VDD.n2420 3.1505
R8413 VDD.n2420 VDD.n2419 3.1505
R8414 VDD.n2424 VDD.n2423 3.1505
R8415 VDD.n2423 VDD.n2422 3.1505
R8416 VDD.n2427 VDD.n2426 3.1505
R8417 VDD.n2426 VDD.n2425 3.1505
R8418 VDD.n2431 VDD.n2430 3.1505
R8419 VDD.n2430 VDD.n2429 3.1505
R8420 VDD.n2434 VDD.n2433 3.1505
R8421 VDD.n2433 VDD.n2432 3.1505
R8422 VDD.n2438 VDD.n2437 3.1505
R8423 VDD.n2437 VDD.n2436 3.1505
R8424 VDD.n2441 VDD.n2440 3.1505
R8425 VDD.n2440 VDD.n2439 3.1505
R8426 VDD.n2445 VDD.n2444 3.1505
R8427 VDD.n2444 VDD.n2443 3.1505
R8428 VDD.n2448 VDD.n2447 3.1505
R8429 VDD.n2447 VDD.n2446 3.1505
R8430 VDD.n2451 VDD.n2450 3.1505
R8431 VDD.n2450 VDD.n2449 3.1505
R8432 VDD.n2456 VDD.n2455 3.1505
R8433 VDD.n2455 VDD.n2454 3.1505
R8434 VDD.n2459 VDD.n2458 3.1505
R8435 VDD.n2458 VDD.n2457 3.1505
R8436 VDD.n2462 VDD.n2461 3.1505
R8437 VDD.n2461 VDD.n2460 3.1505
R8438 VDD.n2466 VDD.n2465 3.1505
R8439 VDD.n2465 VDD.n2464 3.1505
R8440 VDD.n2469 VDD.n2468 3.1505
R8441 VDD.n2468 VDD.n2467 3.1505
R8442 VDD.n2473 VDD.n2472 3.1505
R8443 VDD.n2472 VDD.n2471 3.1505
R8444 VDD.n2476 VDD.n2475 3.1505
R8445 VDD.n2475 VDD.n2474 3.1505
R8446 VDD.n2480 VDD.n2479 3.1505
R8447 VDD.n2479 VDD.n2478 3.1505
R8448 VDD.n2483 VDD.n2482 3.1505
R8449 VDD.n2482 VDD.n2481 3.1505
R8450 VDD.n2486 VDD.n2485 3.1505
R8451 VDD.n2485 VDD.n2484 3.1505
R8452 VDD.n2490 VDD.n2489 3.1505
R8453 VDD.n2489 VDD.n2488 3.1505
R8454 VDD.n2494 VDD.n2493 3.1505
R8455 VDD.n2493 VDD.n2492 3.1505
R8456 VDD.n2497 VDD.n2496 3.1505
R8457 VDD.n2496 VDD.n2495 3.1505
R8458 VDD.n2500 VDD.n2499 3.1505
R8459 VDD.n2499 VDD.n2498 3.1505
R8460 VDD.n2504 VDD.n2503 3.1505
R8461 VDD.n2503 VDD.n2502 3.1505
R8462 VDD.n2508 VDD.n2507 3.1505
R8463 VDD.n2507 VDD.n2506 3.1505
R8464 VDD.n2512 VDD.n2511 3.1505
R8465 VDD.n2511 VDD.n2510 3.1505
R8466 VDD.n2515 VDD.n2514 3.1505
R8467 VDD.n2514 VDD.n2513 3.1505
R8468 VDD.n2518 VDD.n2517 3.1505
R8469 VDD.n2517 VDD.n2516 3.1505
R8470 VDD.n2521 VDD.n2520 3.1505
R8471 VDD.n2520 VDD.n2519 3.1505
R8472 VDD.n2524 VDD.n2523 3.1505
R8473 VDD.n2523 VDD.n2522 3.1505
R8474 VDD.n6804 VDD.n6803 3.1505
R8475 VDD.n777 VDD.n776 3.1505
R8476 VDD.n570 VDD.n569 3.1505
R8477 VDD.n569 VDD.n568 3.1505
R8478 VDD.n566 VDD.n565 3.1505
R8479 VDD.n565 VDD.n564 3.1505
R8480 VDD.n563 VDD.n562 3.1505
R8481 VDD.n562 VDD.n561 3.1505
R8482 VDD.n559 VDD.n558 3.1505
R8483 VDD.n558 VDD.n557 3.1505
R8484 VDD.n1103 VDD.n1102 3.1505
R8485 VDD.n1102 VDD.n1101 3.1505
R8486 VDD.n1100 VDD.n1099 3.1505
R8487 VDD.n1099 VDD.n1098 3.1505
R8488 VDD.n1097 VDD.n1096 3.1505
R8489 VDD.n1096 VDD.n1095 3.1505
R8490 VDD.n1094 VDD.n1093 3.1505
R8491 VDD.n1093 VDD.n1092 3.1505
R8492 VDD.n1091 VDD.n1090 3.1505
R8493 VDD.n1090 VDD.n1089 3.1505
R8494 VDD.n1088 VDD.n1087 3.1505
R8495 VDD.n1087 VDD.n1086 3.1505
R8496 VDD.n1085 VDD.n1084 3.1505
R8497 VDD.n1084 VDD.n1083 3.1505
R8498 VDD.n1082 VDD.n1081 3.1505
R8499 VDD.n1081 VDD.n1080 3.1505
R8500 VDD.n1079 VDD.n1078 3.1505
R8501 VDD.n1078 VDD.n1077 3.1505
R8502 VDD.n1076 VDD.n1075 3.1505
R8503 VDD.n1075 VDD.n1074 3.1505
R8504 VDD.n1073 VDD.n1072 3.1505
R8505 VDD.n1072 VDD.n1071 3.1505
R8506 VDD.n1070 VDD.n1069 3.1505
R8507 VDD.n1069 VDD.n1068 3.1505
R8508 VDD.n1067 VDD.n1066 3.1505
R8509 VDD.n1066 VDD.n1065 3.1505
R8510 VDD.n1064 VDD.n1063 3.1505
R8511 VDD.n1063 VDD.n1062 3.1505
R8512 VDD.n1061 VDD.n1060 3.1505
R8513 VDD.n1060 VDD.n1059 3.1505
R8514 VDD.n1058 VDD.n1057 3.1505
R8515 VDD.n1057 VDD.n1056 3.1505
R8516 VDD.n1055 VDD.n1054 3.1505
R8517 VDD.n1054 VDD.n1053 3.1505
R8518 VDD.n1052 VDD.n1051 3.1505
R8519 VDD.n1051 VDD.n1050 3.1505
R8520 VDD.n1049 VDD.n1048 3.1505
R8521 VDD.n1048 VDD.n1047 3.1505
R8522 VDD.n1046 VDD.n1045 3.1505
R8523 VDD.n1045 VDD.n1044 3.1505
R8524 VDD.n1043 VDD.n1042 3.1505
R8525 VDD.n1042 VDD.n1041 3.1505
R8526 VDD.n1039 VDD.n1038 3.1505
R8527 VDD.n1038 VDD.n1037 3.1505
R8528 VDD.n1036 VDD.n1035 3.1505
R8529 VDD.n1035 VDD.n1034 3.1505
R8530 VDD.n1032 VDD.n1031 3.1505
R8531 VDD.n1031 VDD.n1030 3.1505
R8532 VDD.n1029 VDD.n1028 3.1505
R8533 VDD.n1027 VDD.n1026 3.1505
R8534 VDD.n1026 VDD.n1025 3.1505
R8535 VDD.n1024 VDD.n1023 3.1505
R8536 VDD.n1023 VDD.n1022 3.1505
R8537 VDD.n1021 VDD.n1020 3.1505
R8538 VDD.n1020 VDD.n1019 3.1505
R8539 VDD.n1018 VDD.n1017 3.1505
R8540 VDD.n1017 VDD.n1016 3.1505
R8541 VDD.n1015 VDD.n1014 3.1505
R8542 VDD.n1014 VDD.n1013 3.1505
R8543 VDD.n1012 VDD.n1011 3.1505
R8544 VDD.n1011 VDD.n1010 3.1505
R8545 VDD.n1009 VDD.n1008 3.1505
R8546 VDD.n1008 VDD.n1007 3.1505
R8547 VDD.n1005 VDD.n1004 3.1505
R8548 VDD.n1004 VDD.n1003 3.1505
R8549 VDD.n1002 VDD.n1001 3.1505
R8550 VDD.n1001 VDD.n1000 3.1505
R8551 VDD.n999 VDD.n998 3.1505
R8552 VDD.n998 VDD.n997 3.1505
R8553 VDD.n995 VDD.n994 3.1505
R8554 VDD.n994 VDD.n993 3.1505
R8555 VDD.n992 VDD.n991 3.1505
R8556 VDD.n991 VDD.n990 3.1505
R8557 VDD.n6835 VDD.n6834 3.1505
R8558 VDD.n6834 VDD.n6833 3.1505
R8559 VDD.n6838 VDD.n6837 3.1505
R8560 VDD.n6837 VDD.n6836 3.1505
R8561 VDD.n6842 VDD.n6841 3.1505
R8562 VDD.n6841 VDD.n6840 3.1505
R8563 VDD.n6845 VDD.n6844 3.1505
R8564 VDD.n6844 VDD.n6843 3.1505
R8565 VDD.n6848 VDD.n6847 3.1505
R8566 VDD.n6847 VDD.n6846 3.1505
R8567 VDD.n6852 VDD.n6851 3.1505
R8568 VDD.n6851 VDD.n6850 3.1505
R8569 VDD.n6855 VDD.n6854 3.1505
R8570 VDD.n6854 VDD.n6853 3.1505
R8571 VDD.n6858 VDD.n6857 3.1505
R8572 VDD.n6857 VDD.n6856 3.1505
R8573 VDD.n6862 VDD.n6861 3.1505
R8574 VDD.n6861 VDD.n6860 3.1505
R8575 VDD.n6865 VDD.n6864 3.1505
R8576 VDD.n6864 VDD.n6863 3.1505
R8577 VDD.n6869 VDD.n6868 3.1505
R8578 VDD.n6868 VDD.n6867 3.1505
R8579 VDD.n6872 VDD.n6871 3.1505
R8580 VDD.n6871 VDD.n6870 3.1505
R8581 VDD.n7006 VDD.n7005 3.1505
R8582 VDD.n7005 VDD.n7004 3.1505
R8583 VDD.n7010 VDD.n7009 3.1505
R8584 VDD.n7009 VDD.n7008 3.1505
R8585 VDD.n7013 VDD.n7012 3.1505
R8586 VDD.n7012 VDD.n7011 3.1505
R8587 VDD.n7017 VDD.n7016 3.1505
R8588 VDD.n7016 VDD.n7015 3.1505
R8589 VDD.n7020 VDD.n7019 3.1505
R8590 VDD.n7019 VDD.n7018 3.1505
R8591 VDD.n7023 VDD.n7022 3.1505
R8592 VDD.n7022 VDD.n7021 3.1505
R8593 VDD.n7027 VDD.n7026 3.1505
R8594 VDD.n7026 VDD.n7025 3.1505
R8595 VDD.n7030 VDD.n7029 3.1505
R8596 VDD.n7029 VDD.n7028 3.1505
R8597 VDD.n7033 VDD.n7032 3.1505
R8598 VDD.n7032 VDD.n7031 3.1505
R8599 VDD.n7036 VDD.n7035 3.1505
R8600 VDD.n7035 VDD.n7034 3.1505
R8601 VDD.n7039 VDD.n7038 3.1505
R8602 VDD.n7038 VDD.n7037 3.1505
R8603 VDD.n7043 VDD.n7042 3.1505
R8604 VDD.n7042 VDD.n7041 3.1505
R8605 VDD.n7046 VDD.n7045 3.1505
R8606 VDD.n7045 VDD.n7044 3.1505
R8607 VDD.n7049 VDD.n7048 3.1505
R8608 VDD.n7048 VDD.n7047 3.1505
R8609 VDD.n7052 VDD.n7051 3.1505
R8610 VDD.n7051 VDD.n7050 3.1505
R8611 VDD.n7055 VDD.n7054 3.1505
R8612 VDD.n7054 VDD.n7053 3.1505
R8613 VDD.n7058 VDD.n7057 3.1505
R8614 VDD.n7057 VDD.n7056 3.1505
R8615 VDD.n7062 VDD.n7061 3.1505
R8616 VDD.n7061 VDD.n7060 3.1505
R8617 VDD.n7065 VDD.n7064 3.1505
R8618 VDD.n7064 VDD.n7063 3.1505
R8619 VDD.n7069 VDD.n7068 3.1505
R8620 VDD.n7068 VDD.n7067 3.1505
R8621 VDD.n7072 VDD.n7071 3.1505
R8622 VDD.n7071 VDD.n7070 3.1505
R8623 VDD.n7076 VDD.n7075 3.1505
R8624 VDD.n7075 VDD.n7074 3.1505
R8625 VDD.n7124 VDD.n7123 3.1505
R8626 VDD.n7122 VDD.n7121 3.1505
R8627 VDD.n7120 VDD.n7119 3.1505
R8628 VDD.n7118 VDD.n7117 3.1505
R8629 VDD.n7115 VDD.n7114 3.1505
R8630 VDD.n7113 VDD.n7112 3.1505
R8631 VDD.n7111 VDD.n7110 3.1505
R8632 VDD.n7105 VDD.n7104 3.1505
R8633 VDD.n7103 VDD.n7102 3.1505
R8634 VDD.n7101 VDD.n7100 3.1505
R8635 VDD.n7099 VDD.n7098 3.1505
R8636 VDD.n7096 VDD.n7095 3.1505
R8637 VDD.n7094 VDD.n7093 3.1505
R8638 VDD.n7092 VDD.n7091 3.1505
R8639 VDD.n7090 VDD.n7089 3.1505
R8640 VDD.n7550 VDD.n7549 3.1505
R8641 VDD.n7553 VDD.n7552 3.1505
R8642 VDD.n7556 VDD.n7555 3.1505
R8643 VDD.n7555 VDD.n7554 3.1505
R8644 VDD.n7558 VDD.n7557 3.1505
R8645 VDD.n7561 VDD.n7560 3.1505
R8646 VDD.n7563 VDD.n7562 3.1505
R8647 VDD.n7566 VDD.n7565 3.1505
R8648 VDD.n7568 VDD.n7567 3.1505
R8649 VDD.n7570 VDD.n7569 3.1505
R8650 VDD.n7572 VDD.n7571 3.1505
R8651 VDD.n7575 VDD.n7574 3.1505
R8652 VDD.n7577 VDD.n7576 3.1505
R8653 VDD.n7580 VDD.n7579 3.1505
R8654 VDD.n7582 VDD.n7581 3.1505
R8655 VDD.n7584 VDD.n7583 3.1505
R8656 VDD.n7586 VDD.n7585 3.1505
R8657 VDD.n7588 VDD.n7587 3.1505
R8658 VDD.n7002 VDD.n7001 3.1505
R8659 VDD.n7237 VDD.n7236 3.1505
R8660 VDD.n7240 VDD.n7239 3.1505
R8661 VDD.n7239 VDD.n7238 3.1505
R8662 VDD.n7243 VDD.n7242 3.1505
R8663 VDD.n7242 VDD.n7241 3.1505
R8664 VDD.n7246 VDD.n7245 3.1505
R8665 VDD.n7245 VDD.n7244 3.1505
R8666 VDD.n7250 VDD.n7249 3.1505
R8667 VDD.n7249 VDD.n7248 3.1505
R8668 VDD.n7253 VDD.n7252 3.1505
R8669 VDD.n7252 VDD.n7251 3.1505
R8670 VDD.n7256 VDD.n7255 3.1505
R8671 VDD.n7255 VDD.n7254 3.1505
R8672 VDD.n7260 VDD.n7259 3.1505
R8673 VDD.n7259 VDD.n7258 3.1505
R8674 VDD.n7263 VDD.n7262 3.1505
R8675 VDD.n7262 VDD.n7261 3.1505
R8676 VDD.n7266 VDD.n7265 3.1505
R8677 VDD.n7265 VDD.n7264 3.1505
R8678 VDD.n7269 VDD.n7268 3.1505
R8679 VDD.n7268 VDD.n7267 3.1505
R8680 VDD.n7272 VDD.n7271 3.1505
R8681 VDD.n7271 VDD.n7270 3.1505
R8682 VDD.n7275 VDD.n7274 3.1505
R8683 VDD.n7274 VDD.n7273 3.1505
R8684 VDD.n7278 VDD.n7277 3.1505
R8685 VDD.n7277 VDD.n7276 3.1505
R8686 VDD.n7281 VDD.n7280 3.1505
R8687 VDD.n7280 VDD.n7279 3.1505
R8688 VDD.n7284 VDD.n7283 3.1505
R8689 VDD.n7283 VDD.n7282 3.1505
R8690 VDD.n7287 VDD.n7285 3.1505
R8691 VDD.n7287 VDD.n7286 3.1505
R8692 VDD.n7554 VDD.n7288 3.1505
R8693 VDD.n7725 VDD.n7724 3.1505
R8694 VDD.n7724 VDD.n7723 3.1505
R8695 VDD.n7722 VDD.n7721 3.1505
R8696 VDD.n7721 VDD.n7720 3.1505
R8697 VDD.n7719 VDD.n7718 3.1505
R8698 VDD.n7718 VDD.n7717 3.1505
R8699 VDD.n7716 VDD.n7715 3.1505
R8700 VDD.n7715 VDD.n7714 3.1505
R8701 VDD.n7713 VDD.n7712 3.1505
R8702 VDD.n7712 VDD.n7711 3.1505
R8703 VDD.n7710 VDD.n7709 3.1505
R8704 VDD.n7709 VDD.n7708 3.1505
R8705 VDD.n7707 VDD.n7706 3.1505
R8706 VDD.n7706 VDD.n7705 3.1505
R8707 VDD.n7703 VDD.n7702 3.1505
R8708 VDD.n7702 VDD.n7701 3.1505
R8709 VDD.n7700 VDD.n7699 3.1505
R8710 VDD.n7699 VDD.n7698 3.1505
R8711 VDD.n7696 VDD.n7695 3.1505
R8712 VDD.n7695 VDD.n7694 3.1505
R8713 VDD.n7693 VDD.n7692 3.1505
R8714 VDD.n7692 VDD.n7691 3.1505
R8715 VDD.n7690 VDD.n7689 3.1505
R8716 VDD.n7689 VDD.n7688 3.1505
R8717 VDD.n7687 VDD.n7686 3.1505
R8718 VDD.n7686 VDD.n7685 3.1505
R8719 VDD.n7684 VDD.n7683 3.1505
R8720 VDD.n292 VDD.t1392 3.08583
R8721 VDD.n288 VDD.t1210 3.08583
R8722 VDD.n287 VDD.t1275 3.08583
R8723 VDD.n16 VDD.t1180 3.08583
R8724 VDD.n17 VDD.t1255 3.08583
R8725 VDD.n18 VDD.t1367 3.08583
R8726 VDD.n6884 VDD.t1268 3.08583
R8727 VDD.n6880 VDD.t1157 3.08583
R8728 VDD.n6879 VDD.t1282 3.08583
R8729 VDD.n19 VDD.t1375 3.08583
R8730 VDD.n20 VDD.t1195 3.08583
R8731 VDD.n21 VDD.t1305 3.08583
R8732 VDD.n2076 VDD.t10 3.07932
R8733 VDD.n2234 VDD.t366 3.07932
R8734 VDD.n2318 VDD.t396 3.07932
R8735 VDD.n2436 VDD.t306 3.07932
R8736 VDD.n7359 VDD.t1349 3.0555
R8737 VDD.n388 VDD.t1207 3.0555
R8738 VDD.n7374 VDD.t1213 3.0555
R8739 VDD.n7251 VDD.t1153 2.97991
R8740 VDD.n2692 VDD.n2691 2.87353
R8741 VDD.n5615 VDD.t23 2.8495
R8742 VDD.n5621 VDD.t142 2.8495
R8743 VDD.n6086 VDD.t145 2.8495
R8744 VDD.n6092 VDD.t526 2.8495
R8745 VDD.n6233 VDD.t1107 2.8495
R8746 VDD.n6239 VDD.t202 2.8495
R8747 VDD.n6388 VDD.t7 2.8495
R8748 VDD.n6394 VDD.t171 2.8495
R8749 VDD.n6547 VDD.t199 2.8495
R8750 VDD.n6553 VDD.t336 2.8495
R8751 VDD.n5784 VDD.t515 2.8495
R8752 VDD.n5790 VDD.t195 2.8495
R8753 VDD.n5931 VDD.t173 2.8495
R8754 VDD.n5937 VDD.t140 2.8495
R8755 VDD.n2243 VDD.t183 2.66881
R8756 VDD.n2443 VDD.t331 2.66881
R8757 VDD.n322 VDD.t1159 2.6092
R8758 VDD.n329 VDD.t192 2.6092
R8759 VDD.n360 VDD.t1134 2.6092
R8760 VDD.n357 VDD.t1092 2.6092
R8761 VDD.n7082 VDD.n7081 2.6005
R8762 VDD.n7085 VDD.n7084 2.6005
R8763 VDD.n7088 VDD.n7087 2.6005
R8764 VDD.n7542 VDD.n7541 2.6005
R8765 VDD.n7545 VDD.n7544 2.6005
R8766 VDD.n7548 VDD.n7547 2.6005
R8767 VDD.n7309 VDD.n7308 2.6005
R8768 VDD.n7312 VDD.n7311 2.6005
R8769 VDD.n7315 VDD.n7314 2.6005
R8770 VDD.n7295 VDD.n7291 2.6005
R8771 VDD.n7296 VDD.n7290 2.6005
R8772 VDD.n7297 VDD.n7289 2.6005
R8773 VDD.n7304 VDD.n7303 2.6005
R8774 VDD.n404 VDD.n403 2.6005
R8775 VDD.n980 VDD.n979 2.6005
R8776 VDD.n977 VDD.n976 2.6005
R8777 VDD.n974 VDD.n973 2.6005
R8778 VDD.n801 VDD.n800 2.6005
R8779 VDD.n989 VDD.n988 2.6005
R8780 VDD.n986 VDD.n985 2.6005
R8781 VDD.n983 VDD.n982 2.6005
R8782 VDD.n804 VDD.n803 2.6005
R8783 VDD.n6832 VDD.n6831 2.6005
R8784 VDD.n6829 VDD.n6828 2.6005
R8785 VDD.n6826 VDD.n6825 2.6005
R8786 VDD.n6656 VDD.n6655 2.6005
R8787 VDD.n6823 VDD.n6822 2.6005
R8788 VDD.n6820 VDD.n6819 2.6005
R8789 VDD.n6817 VDD.n6816 2.6005
R8790 VDD.n6653 VDD.n6652 2.6005
R8791 VDD.n5427 VDD.n5426 2.6005
R8792 VDD.n5424 VDD.n5423 2.6005
R8793 VDD.n3314 VDD.n3313 2.6005
R8794 VDD.n3315 VDD.n3311 2.6005
R8795 VDD.n5421 VDD.n5420 2.6005
R8796 VDD.n5418 VDD.n5417 2.6005
R8797 VDD.n3308 VDD.n3307 2.6005
R8798 VDD.n3309 VDD.n3305 2.6005
R8799 VDD.n5415 VDD.n5414 2.6005
R8800 VDD.n5412 VDD.n5411 2.6005
R8801 VDD.n3302 VDD.n3301 2.6005
R8802 VDD.n3303 VDD.n3299 2.6005
R8803 VDD.n3297 VDD.n3287 2.6005
R8804 VDD.n3295 VDD.n3294 2.6005
R8805 VDD.n5396 VDD.n5395 2.6005
R8806 VDD.n5405 VDD.n5404 2.6005
R8807 VDD.n5387 VDD.n5386 2.6005
R8808 VDD.n5384 VDD.n5383 2.6005
R8809 VDD.n3284 VDD.n3283 2.6005
R8810 VDD.n3285 VDD.n3281 2.6005
R8811 VDD.n5381 VDD.n5380 2.6005
R8812 VDD.n5378 VDD.n5377 2.6005
R8813 VDD.n3278 VDD.n3277 2.6005
R8814 VDD.n3279 VDD.n3275 2.6005
R8815 VDD.n4079 VDD.n4078 2.6005
R8816 VDD.n4076 VDD.n4075 2.6005
R8817 VDD.n2919 VDD.n2918 2.6005
R8818 VDD.n2920 VDD.n2916 2.6005
R8819 VDD.n4085 VDD.n4084 2.6005
R8820 VDD.n4082 VDD.n4081 2.6005
R8821 VDD.n2925 VDD.n2924 2.6005
R8822 VDD.n2926 VDD.n2922 2.6005
R8823 VDD.n4091 VDD.n4090 2.6005
R8824 VDD.n4088 VDD.n4087 2.6005
R8825 VDD.n2931 VDD.n2930 2.6005
R8826 VDD.n2932 VDD.n2928 2.6005
R8827 VDD.n4113 VDD.n4112 2.6005
R8828 VDD.n4109 VDD.n4108 2.6005
R8829 VDD.n2937 VDD.n2936 2.6005
R8830 VDD.n2944 VDD.n2934 2.6005
R8831 VDD.n4119 VDD.n4118 2.6005
R8832 VDD.n4116 VDD.n4115 2.6005
R8833 VDD.n2949 VDD.n2948 2.6005
R8834 VDD.n2950 VDD.n2946 2.6005
R8835 VDD.n4125 VDD.n4124 2.6005
R8836 VDD.n4122 VDD.n4121 2.6005
R8837 VDD.n2955 VDD.n2954 2.6005
R8838 VDD.n2956 VDD.n2952 2.6005
R8839 VDD.n4399 VDD.n4398 2.6005
R8840 VDD.n4396 VDD.n4395 2.6005
R8841 VDD.n2989 VDD.n2988 2.6005
R8842 VDD.n2990 VDD.n2986 2.6005
R8843 VDD.n4405 VDD.n4404 2.6005
R8844 VDD.n4402 VDD.n4401 2.6005
R8845 VDD.n2995 VDD.n2994 2.6005
R8846 VDD.n2996 VDD.n2992 2.6005
R8847 VDD.n4423 VDD.n4422 2.6005
R8848 VDD.n4419 VDD.n4418 2.6005
R8849 VDD.n3001 VDD.n3000 2.6005
R8850 VDD.n3008 VDD.n2998 2.6005
R8851 VDD.n4433 VDD.n4432 2.6005
R8852 VDD.n4430 VDD.n4429 2.6005
R8853 VDD.n3013 VDD.n3012 2.6005
R8854 VDD.n3014 VDD.n3010 2.6005
R8855 VDD.n4439 VDD.n4438 2.6005
R8856 VDD.n4436 VDD.n4435 2.6005
R8857 VDD.n3019 VDD.n3018 2.6005
R8858 VDD.n3020 VDD.n3016 2.6005
R8859 VDD.n4445 VDD.n4444 2.6005
R8860 VDD.n4442 VDD.n4441 2.6005
R8861 VDD.n3025 VDD.n3024 2.6005
R8862 VDD.n3026 VDD.n3022 2.6005
R8863 VDD.n4589 VDD.n4588 2.6005
R8864 VDD.n4586 VDD.n4585 2.6005
R8865 VDD.n3049 VDD.n3048 2.6005
R8866 VDD.n3050 VDD.n3046 2.6005
R8867 VDD.n4595 VDD.n4594 2.6005
R8868 VDD.n4592 VDD.n4591 2.6005
R8869 VDD.n3055 VDD.n3054 2.6005
R8870 VDD.n3056 VDD.n3052 2.6005
R8871 VDD.n4601 VDD.n4600 2.6005
R8872 VDD.n4598 VDD.n4597 2.6005
R8873 VDD.n3061 VDD.n3060 2.6005
R8874 VDD.n3062 VDD.n3058 2.6005
R8875 VDD.n4623 VDD.n4622 2.6005
R8876 VDD.n4619 VDD.n4618 2.6005
R8877 VDD.n3067 VDD.n3066 2.6005
R8878 VDD.n3074 VDD.n3064 2.6005
R8879 VDD.n4629 VDD.n4628 2.6005
R8880 VDD.n4626 VDD.n4625 2.6005
R8881 VDD.n3079 VDD.n3078 2.6005
R8882 VDD.n3080 VDD.n3076 2.6005
R8883 VDD.n4635 VDD.n4634 2.6005
R8884 VDD.n4632 VDD.n4631 2.6005
R8885 VDD.n3085 VDD.n3084 2.6005
R8886 VDD.n3086 VDD.n3082 2.6005
R8887 VDD.n4903 VDD.n4902 2.6005
R8888 VDD.n4900 VDD.n4899 2.6005
R8889 VDD.n3125 VDD.n3124 2.6005
R8890 VDD.n3126 VDD.n3122 2.6005
R8891 VDD.n4909 VDD.n4908 2.6005
R8892 VDD.n4906 VDD.n4905 2.6005
R8893 VDD.n3131 VDD.n3130 2.6005
R8894 VDD.n3132 VDD.n3128 2.6005
R8895 VDD.n4927 VDD.n4926 2.6005
R8896 VDD.n4923 VDD.n4922 2.6005
R8897 VDD.n3137 VDD.n3136 2.6005
R8898 VDD.n3144 VDD.n3134 2.6005
R8899 VDD.n4937 VDD.n4936 2.6005
R8900 VDD.n4934 VDD.n4933 2.6005
R8901 VDD.n3149 VDD.n3148 2.6005
R8902 VDD.n3150 VDD.n3146 2.6005
R8903 VDD.n4943 VDD.n4942 2.6005
R8904 VDD.n4940 VDD.n4939 2.6005
R8905 VDD.n3155 VDD.n3154 2.6005
R8906 VDD.n3156 VDD.n3152 2.6005
R8907 VDD.n4949 VDD.n4948 2.6005
R8908 VDD.n4946 VDD.n4945 2.6005
R8909 VDD.n3161 VDD.n3160 2.6005
R8910 VDD.n3162 VDD.n3158 2.6005
R8911 VDD.n5135 VDD.n5134 2.6005
R8912 VDD.n5132 VDD.n5131 2.6005
R8913 VDD.n3230 VDD.n3229 2.6005
R8914 VDD.n3231 VDD.n3227 2.6005
R8915 VDD.n5129 VDD.n5128 2.6005
R8916 VDD.n5126 VDD.n5125 2.6005
R8917 VDD.n3224 VDD.n3223 2.6005
R8918 VDD.n3225 VDD.n3221 2.6005
R8919 VDD.n3219 VDD.n3209 2.6005
R8920 VDD.n3217 VDD.n3216 2.6005
R8921 VDD.n5114 VDD.n5113 2.6005
R8922 VDD.n5123 VDD.n5122 2.6005
R8923 VDD.n5101 VDD.n5100 2.6005
R8924 VDD.n5098 VDD.n5097 2.6005
R8925 VDD.n3206 VDD.n3205 2.6005
R8926 VDD.n3207 VDD.n3203 2.6005
R8927 VDD.n5095 VDD.n5094 2.6005
R8928 VDD.n5092 VDD.n5091 2.6005
R8929 VDD.n3200 VDD.n3199 2.6005
R8930 VDD.n3201 VDD.n3197 2.6005
R8931 VDD.n5089 VDD.n5088 2.6005
R8932 VDD.n5086 VDD.n5085 2.6005
R8933 VDD.n3194 VDD.n3193 2.6005
R8934 VDD.n3195 VDD.n3191 2.6005
R8935 VDD.n2850 VDD.n2849 2.6005
R8936 VDD.n2847 VDD.n2846 2.6005
R8937 VDD.n2549 VDD.n2548 2.6005
R8938 VDD.n2550 VDD.n2546 2.6005
R8939 VDD.n2856 VDD.n2855 2.6005
R8940 VDD.n2853 VDD.n2852 2.6005
R8941 VDD.n2555 VDD.n2554 2.6005
R8942 VDD.n2556 VDD.n2552 2.6005
R8943 VDD.n2874 VDD.n2873 2.6005
R8944 VDD.n2870 VDD.n2869 2.6005
R8945 VDD.n2561 VDD.n2560 2.6005
R8946 VDD.n2568 VDD.n2558 2.6005
R8947 VDD.n2884 VDD.n2883 2.6005
R8948 VDD.n2881 VDD.n2880 2.6005
R8949 VDD.n2573 VDD.n2572 2.6005
R8950 VDD.n2574 VDD.n2570 2.6005
R8951 VDD.n2890 VDD.n2889 2.6005
R8952 VDD.n2887 VDD.n2886 2.6005
R8953 VDD.n2579 VDD.n2578 2.6005
R8954 VDD.n2580 VDD.n2576 2.6005
R8955 VDD.n2896 VDD.n2895 2.6005
R8956 VDD.n2893 VDD.n2892 2.6005
R8957 VDD.n2585 VDD.n2584 2.6005
R8958 VDD.n2586 VDD.n2582 2.6005
R8959 VDD.n1370 VDD.n1367 2.6005
R8960 VDD.n1371 VDD.n1365 2.6005
R8961 VDD.n1372 VDD.n1363 2.6005
R8962 VDD.n1381 VDD.n1378 2.6005
R8963 VDD.n1382 VDD.n1376 2.6005
R8964 VDD.n1383 VDD.n1374 2.6005
R8965 VDD.n1392 VDD.n1389 2.6005
R8966 VDD.n1393 VDD.n1387 2.6005
R8967 VDD.n1394 VDD.n1385 2.6005
R8968 VDD.n1403 VDD.n1400 2.6005
R8969 VDD.n1404 VDD.n1398 2.6005
R8970 VDD.n1405 VDD.n1396 2.6005
R8971 VDD.n1414 VDD.n1411 2.6005
R8972 VDD.n1415 VDD.n1409 2.6005
R8973 VDD.n1416 VDD.n1407 2.6005
R8974 VDD.n1425 VDD.n1422 2.6005
R8975 VDD.n1426 VDD.n1420 2.6005
R8976 VDD.n1427 VDD.n1418 2.6005
R8977 VDD.n1439 VDD.n1435 2.6005
R8978 VDD.n1438 VDD.n1437 2.6005
R8979 VDD.n1124 VDD.n1123 2.6005
R8980 VDD.n1127 VDD.n1126 2.6005
R8981 VDD.n1433 VDD.n1429 2.6005
R8982 VDD.n1432 VDD.n1431 2.6005
R8983 VDD.n1118 VDD.n1117 2.6005
R8984 VDD.n1121 VDD.n1120 2.6005
R8985 VDD.n1361 VDD.n1357 2.6005
R8986 VDD.n1112 VDD.n1111 2.6005
R8987 VDD.n1359 VDD.n1358 2.6005
R8988 VDD.n1115 VDD.n1114 2.6005
R8989 VDD.n11 VDD.n1 2.6005
R8990 VDD.n10 VDD.n3 2.6005
R8991 VDD.n9 VDD.n5 2.6005
R8992 VDD.n7108 VDD.n7107 2.6005
R8993 VDD.n7222 VDD.n7221 2.48924
R8994 VDD.n7219 VDD.n7218 2.48924
R8995 VDD.n7216 VDD.n7215 2.48924
R8996 VDD.n7213 VDD.n7212 2.48924
R8997 VDD.n7210 VDD.n7209 2.48924
R8998 VDD.n7207 VDD.n7206 2.48924
R8999 VDD.n7204 VDD.n7203 2.48924
R9000 VDD.n7201 VDD.n7200 2.48924
R9001 VDD.n7198 VDD.n7197 2.48924
R9002 VDD.n7195 VDD.n7194 2.48924
R9003 VDD.n7192 VDD.n7191 2.48924
R9004 VDD.n7189 VDD.n7188 2.48924
R9005 VDD.n7186 VDD.n7185 2.48924
R9006 VDD.n7183 VDD.n7182 2.48924
R9007 VDD.n7180 VDD.n7179 2.48924
R9008 VDD.n7177 VDD.n7176 2.48924
R9009 VDD.n7174 VDD.n7173 2.48924
R9010 VDD.n7171 VDD.n7170 2.48924
R9011 VDD.n7168 VDD.n7167 2.48924
R9012 VDD.n7165 VDD.n7164 2.48924
R9013 VDD.n7162 VDD.n7161 2.48924
R9014 VDD.n7159 VDD.n7158 2.48924
R9015 VDD.n7156 VDD.n7155 2.48924
R9016 VDD.n7153 VDD.n7152 2.48924
R9017 VDD.n7150 VDD.n7149 2.48924
R9018 VDD.n6910 VDD.n6909 2.48924
R9019 VDD.n6913 VDD.n6912 2.48924
R9020 VDD.n6916 VDD.n6915 2.48924
R9021 VDD.n6919 VDD.n6918 2.48924
R9022 VDD.n6922 VDD.n6921 2.48924
R9023 VDD.n6925 VDD.n6924 2.48924
R9024 VDD.n6928 VDD.n6927 2.48924
R9025 VDD.n6931 VDD.n6930 2.48924
R9026 VDD.n6934 VDD.n6933 2.48924
R9027 VDD.n6937 VDD.n6936 2.48924
R9028 VDD.n6940 VDD.n6939 2.48924
R9029 VDD.n6943 VDD.n6942 2.48924
R9030 VDD.n6946 VDD.n6945 2.48924
R9031 VDD.n6949 VDD.n6948 2.48924
R9032 VDD.n6952 VDD.n6951 2.48924
R9033 VDD.n6955 VDD.n6954 2.48924
R9034 VDD.n6958 VDD.n6957 2.48924
R9035 VDD.n6961 VDD.n6960 2.48924
R9036 VDD.n6964 VDD.n6963 2.48924
R9037 VDD.n6967 VDD.n6966 2.48924
R9038 VDD.n6970 VDD.n6969 2.48924
R9039 VDD.n6973 VDD.n6972 2.48924
R9040 VDD.n6976 VDD.n6975 2.48924
R9041 VDD.n6979 VDD.n6978 2.48924
R9042 VDD.n6982 VDD.n6981 2.48924
R9043 VDD.n6985 VDD.n6984 2.48924
R9044 VDD.n676 VDD.n675 2.48924
R9045 VDD.n679 VDD.n678 2.48924
R9046 VDD.n682 VDD.n681 2.48924
R9047 VDD.n685 VDD.n684 2.48924
R9048 VDD.n688 VDD.n687 2.48924
R9049 VDD.n691 VDD.n690 2.48924
R9050 VDD.n694 VDD.n693 2.48924
R9051 VDD.n697 VDD.n696 2.48924
R9052 VDD.n700 VDD.n699 2.48924
R9053 VDD.n703 VDD.n702 2.48924
R9054 VDD.n706 VDD.n705 2.48924
R9055 VDD.n709 VDD.n708 2.48924
R9056 VDD.n712 VDD.n711 2.48924
R9057 VDD.n715 VDD.n714 2.48924
R9058 VDD.n718 VDD.n717 2.48924
R9059 VDD.n721 VDD.n720 2.48924
R9060 VDD.n724 VDD.n723 2.48924
R9061 VDD.n727 VDD.n726 2.48924
R9062 VDD.n730 VDD.n729 2.48924
R9063 VDD.n733 VDD.n732 2.48924
R9064 VDD.n736 VDD.n735 2.48924
R9065 VDD.n739 VDD.n738 2.48924
R9066 VDD.n742 VDD.n741 2.48924
R9067 VDD.n745 VDD.n744 2.48924
R9068 VDD.n748 VDD.n747 2.48924
R9069 VDD.n751 VDD.n750 2.48924
R9070 VDD.n876 VDD.n875 2.48924
R9071 VDD.n879 VDD.n878 2.48924
R9072 VDD.n882 VDD.n881 2.48924
R9073 VDD.n885 VDD.n884 2.48924
R9074 VDD.n888 VDD.n887 2.48924
R9075 VDD.n891 VDD.n890 2.48924
R9076 VDD.n894 VDD.n893 2.48924
R9077 VDD.n897 VDD.n896 2.48924
R9078 VDD.n900 VDD.n899 2.48924
R9079 VDD.n903 VDD.n902 2.48924
R9080 VDD.n906 VDD.n905 2.48924
R9081 VDD.n909 VDD.n908 2.48924
R9082 VDD.n912 VDD.n911 2.48924
R9083 VDD.n915 VDD.n914 2.48924
R9084 VDD.n918 VDD.n917 2.48924
R9085 VDD.n921 VDD.n920 2.48924
R9086 VDD.n924 VDD.n923 2.48924
R9087 VDD.n927 VDD.n926 2.48924
R9088 VDD.n930 VDD.n929 2.48924
R9089 VDD.n933 VDD.n932 2.48924
R9090 VDD.n936 VDD.n935 2.48924
R9091 VDD.n939 VDD.n938 2.48924
R9092 VDD.n942 VDD.n941 2.48924
R9093 VDD.n2697 VDD.n2696 2.48924
R9094 VDD.n2700 VDD.n2699 2.48924
R9095 VDD.n2703 VDD.n2702 2.48924
R9096 VDD.n2706 VDD.n2705 2.48924
R9097 VDD.n2709 VDD.n2708 2.48924
R9098 VDD.n2712 VDD.n2711 2.48924
R9099 VDD.n2715 VDD.n2714 2.48924
R9100 VDD.n2718 VDD.n2717 2.48924
R9101 VDD.n2721 VDD.n2720 2.48924
R9102 VDD.n2724 VDD.n2723 2.48924
R9103 VDD.n2727 VDD.n2726 2.48924
R9104 VDD.n2730 VDD.n2729 2.48924
R9105 VDD.n2733 VDD.n2732 2.48924
R9106 VDD.n2736 VDD.n2735 2.48924
R9107 VDD.n2739 VDD.n2738 2.48924
R9108 VDD.n2742 VDD.n2741 2.48924
R9109 VDD.n2745 VDD.n2744 2.48924
R9110 VDD.n2748 VDD.n2747 2.48924
R9111 VDD.n2751 VDD.n2750 2.48924
R9112 VDD.n2754 VDD.n2753 2.48924
R9113 VDD.n2757 VDD.n2756 2.48924
R9114 VDD.n2760 VDD.n2759 2.48924
R9115 VDD.n2763 VDD.n2762 2.48924
R9116 VDD.n2766 VDD.n2765 2.48924
R9117 VDD.n2769 VDD.n2768 2.48924
R9118 VDD.n2772 VDD.n2771 2.48924
R9119 VDD.n2775 VDD.n2774 2.48924
R9120 VDD.n2778 VDD.n2777 2.48924
R9121 VDD.n2781 VDD.n2780 2.48924
R9122 VDD.n2784 VDD.n2783 2.48924
R9123 VDD.n2787 VDD.n2786 2.48924
R9124 VDD.n2790 VDD.n2789 2.48924
R9125 VDD.n2793 VDD.n2792 2.48924
R9126 VDD.n2796 VDD.n2795 2.48924
R9127 VDD.n2799 VDD.n2798 2.48924
R9128 VDD.n2802 VDD.n2801 2.48924
R9129 VDD.n2805 VDD.n2804 2.48924
R9130 VDD.n2808 VDD.n2807 2.48924
R9131 VDD.n2811 VDD.n2810 2.48924
R9132 VDD.n2814 VDD.n2813 2.48924
R9133 VDD.n2817 VDD.n2816 2.48924
R9134 VDD.n2820 VDD.n2819 2.48924
R9135 VDD.n2823 VDD.n2822 2.48924
R9136 VDD.n2826 VDD.n2825 2.48924
R9137 VDD.n2829 VDD.n2828 2.48924
R9138 VDD.n2832 VDD.n2831 2.48924
R9139 VDD.n2975 VDD.n2974 2.48924
R9140 VDD.n4137 VDD.n4136 2.48924
R9141 VDD.n4140 VDD.n4139 2.48924
R9142 VDD.n4143 VDD.n4142 2.48924
R9143 VDD.n4146 VDD.n4145 2.48924
R9144 VDD.n4149 VDD.n4148 2.48924
R9145 VDD.n4152 VDD.n4151 2.48924
R9146 VDD.n4155 VDD.n4154 2.48924
R9147 VDD.n4158 VDD.n4157 2.48924
R9148 VDD.n4161 VDD.n4160 2.48924
R9149 VDD.n4164 VDD.n4163 2.48924
R9150 VDD.n4167 VDD.n4166 2.48924
R9151 VDD.n4170 VDD.n4169 2.48924
R9152 VDD.n4173 VDD.n4172 2.48924
R9153 VDD.n4176 VDD.n4175 2.48924
R9154 VDD.n4179 VDD.n4178 2.48924
R9155 VDD.n4182 VDD.n4181 2.48924
R9156 VDD.n4185 VDD.n4184 2.48924
R9157 VDD.n4188 VDD.n4187 2.48924
R9158 VDD.n4191 VDD.n4190 2.48924
R9159 VDD.n4194 VDD.n4193 2.48924
R9160 VDD.n4197 VDD.n4196 2.48924
R9161 VDD.n4200 VDD.n4199 2.48924
R9162 VDD.n4203 VDD.n4202 2.48924
R9163 VDD.n4206 VDD.n4205 2.48924
R9164 VDD.n4209 VDD.n4208 2.48924
R9165 VDD.n4212 VDD.n4211 2.48924
R9166 VDD.n4215 VDD.n4214 2.48924
R9167 VDD.n4218 VDD.n4217 2.48924
R9168 VDD.n4221 VDD.n4220 2.48924
R9169 VDD.n4224 VDD.n4223 2.48924
R9170 VDD.n4227 VDD.n4226 2.48924
R9171 VDD.n4230 VDD.n4229 2.48924
R9172 VDD.n4233 VDD.n4232 2.48924
R9173 VDD.n4236 VDD.n4235 2.48924
R9174 VDD.n4239 VDD.n4238 2.48924
R9175 VDD.n4242 VDD.n4241 2.48924
R9176 VDD.n4245 VDD.n4244 2.48924
R9177 VDD.n4248 VDD.n4247 2.48924
R9178 VDD.n4251 VDD.n4250 2.48924
R9179 VDD.n4254 VDD.n4253 2.48924
R9180 VDD.n4257 VDD.n4256 2.48924
R9181 VDD.n4260 VDD.n4259 2.48924
R9182 VDD.n3845 VDD.n3844 2.48924
R9183 VDD.n4647 VDD.n4646 2.48924
R9184 VDD.n4650 VDD.n4649 2.48924
R9185 VDD.n4653 VDD.n4652 2.48924
R9186 VDD.n4656 VDD.n4655 2.48924
R9187 VDD.n4659 VDD.n4658 2.48924
R9188 VDD.n4662 VDD.n4661 2.48924
R9189 VDD.n4665 VDD.n4664 2.48924
R9190 VDD.n4668 VDD.n4667 2.48924
R9191 VDD.n4671 VDD.n4670 2.48924
R9192 VDD.n4674 VDD.n4673 2.48924
R9193 VDD.n4677 VDD.n4676 2.48924
R9194 VDD.n4680 VDD.n4679 2.48924
R9195 VDD.n4683 VDD.n4682 2.48924
R9196 VDD.n4686 VDD.n4685 2.48924
R9197 VDD.n4689 VDD.n4688 2.48924
R9198 VDD.n4692 VDD.n4691 2.48924
R9199 VDD.n4695 VDD.n4694 2.48924
R9200 VDD.n4698 VDD.n4697 2.48924
R9201 VDD.n4701 VDD.n4700 2.48924
R9202 VDD.n4704 VDD.n4703 2.48924
R9203 VDD.n4707 VDD.n4706 2.48924
R9204 VDD.n4710 VDD.n4709 2.48924
R9205 VDD.n4713 VDD.n4712 2.48924
R9206 VDD.n4716 VDD.n4715 2.48924
R9207 VDD.n4719 VDD.n4718 2.48924
R9208 VDD.n4722 VDD.n4721 2.48924
R9209 VDD.n4725 VDD.n4724 2.48924
R9210 VDD.n4728 VDD.n4727 2.48924
R9211 VDD.n4731 VDD.n4730 2.48924
R9212 VDD.n4734 VDD.n4733 2.48924
R9213 VDD.n4737 VDD.n4736 2.48924
R9214 VDD.n4740 VDD.n4739 2.48924
R9215 VDD.n4743 VDD.n4742 2.48924
R9216 VDD.n4746 VDD.n4745 2.48924
R9217 VDD.n4749 VDD.n4748 2.48924
R9218 VDD.n4752 VDD.n4751 2.48924
R9219 VDD.n4755 VDD.n4754 2.48924
R9220 VDD.n4758 VDD.n4757 2.48924
R9221 VDD.n4761 VDD.n4760 2.48924
R9222 VDD.n4764 VDD.n4763 2.48924
R9223 VDD.n4767 VDD.n4766 2.48924
R9224 VDD.n3098 VDD.n3097 2.48924
R9225 VDD.n3111 VDD.n3110 2.48924
R9226 VDD.n3640 VDD.n3639 2.48924
R9227 VDD.n5148 VDD.n5147 2.48924
R9228 VDD.n5151 VDD.n5150 2.48924
R9229 VDD.n5154 VDD.n5153 2.48924
R9230 VDD.n5157 VDD.n5156 2.48924
R9231 VDD.n5160 VDD.n5159 2.48924
R9232 VDD.n5163 VDD.n5162 2.48924
R9233 VDD.n5166 VDD.n5165 2.48924
R9234 VDD.n5169 VDD.n5168 2.48924
R9235 VDD.n5172 VDD.n5171 2.48924
R9236 VDD.n5175 VDD.n5174 2.48924
R9237 VDD.n5178 VDD.n5177 2.48924
R9238 VDD.n5181 VDD.n5180 2.48924
R9239 VDD.n5184 VDD.n5183 2.48924
R9240 VDD.n5187 VDD.n5186 2.48924
R9241 VDD.n5190 VDD.n5189 2.48924
R9242 VDD.n5193 VDD.n5192 2.48924
R9243 VDD.n5196 VDD.n5195 2.48924
R9244 VDD.n5199 VDD.n5198 2.48924
R9245 VDD.n5202 VDD.n5201 2.48924
R9246 VDD.n5205 VDD.n5204 2.48924
R9247 VDD.n5208 VDD.n5207 2.48924
R9248 VDD.n5211 VDD.n5210 2.48924
R9249 VDD.n5214 VDD.n5213 2.48924
R9250 VDD.n5217 VDD.n5216 2.48924
R9251 VDD.n5220 VDD.n5219 2.48924
R9252 VDD.n5223 VDD.n5222 2.48924
R9253 VDD.n5226 VDD.n5225 2.48924
R9254 VDD.n5229 VDD.n5228 2.48924
R9255 VDD.n5232 VDD.n5231 2.48924
R9256 VDD.n5235 VDD.n5234 2.48924
R9257 VDD.n5238 VDD.n5237 2.48924
R9258 VDD.n5241 VDD.n5240 2.48924
R9259 VDD.n5244 VDD.n5243 2.48924
R9260 VDD.n5247 VDD.n5246 2.48924
R9261 VDD.n5250 VDD.n5249 2.48924
R9262 VDD.n5253 VDD.n5252 2.48924
R9263 VDD.n5256 VDD.n5255 2.48924
R9264 VDD.n5259 VDD.n5258 2.48924
R9265 VDD.n5262 VDD.n5261 2.48924
R9266 VDD.n3248 VDD.n3247 2.48924
R9267 VDD.n3245 VDD.n3244 2.48924
R9268 VDD.n3242 VDD.n3241 2.48924
R9269 VDD.n1791 VDD.n1790 2.48924
R9270 VDD.n1788 VDD.n1787 2.48924
R9271 VDD.n1785 VDD.n1784 2.48924
R9272 VDD.n1782 VDD.n1781 2.48924
R9273 VDD.n1779 VDD.n1778 2.48924
R9274 VDD.n1776 VDD.n1775 2.48924
R9275 VDD.n1773 VDD.n1772 2.48924
R9276 VDD.n1770 VDD.n1769 2.48924
R9277 VDD.n1767 VDD.n1766 2.48924
R9278 VDD.n1764 VDD.n1763 2.48924
R9279 VDD.n1761 VDD.n1760 2.48924
R9280 VDD.n1758 VDD.n1757 2.48924
R9281 VDD.n1755 VDD.n1754 2.48924
R9282 VDD.n1752 VDD.n1751 2.48924
R9283 VDD.n1749 VDD.n1748 2.48924
R9284 VDD.n1746 VDD.n1745 2.48924
R9285 VDD.n1743 VDD.n1742 2.48924
R9286 VDD.n1740 VDD.n1739 2.48924
R9287 VDD.n1737 VDD.n1736 2.48924
R9288 VDD.n1734 VDD.n1733 2.48924
R9289 VDD.n1731 VDD.n1730 2.48924
R9290 VDD.n1728 VDD.n1727 2.48924
R9291 VDD.n1725 VDD.n1724 2.48924
R9292 VDD.n1722 VDD.n1721 2.48924
R9293 VDD.n1719 VDD.n1718 2.48924
R9294 VDD.n1716 VDD.n1715 2.48924
R9295 VDD.n1713 VDD.n1712 2.48924
R9296 VDD.n1710 VDD.n1709 2.48924
R9297 VDD.n1707 VDD.n1706 2.48924
R9298 VDD.n1704 VDD.n1703 2.48924
R9299 VDD.n1701 VDD.n1700 2.48924
R9300 VDD.n1698 VDD.n1697 2.48924
R9301 VDD.n1695 VDD.n1694 2.48924
R9302 VDD.n1692 VDD.n1691 2.48924
R9303 VDD.n1689 VDD.n1688 2.48924
R9304 VDD.n1686 VDD.n1685 2.48924
R9305 VDD.n1683 VDD.n1682 2.48924
R9306 VDD.n1680 VDD.n1679 2.48924
R9307 VDD.n1929 VDD.n1928 2.48924
R9308 VDD.n1926 VDD.n1925 2.48924
R9309 VDD.n1923 VDD.n1922 2.48924
R9310 VDD.n1920 VDD.n1919 2.48924
R9311 VDD.n1917 VDD.n1916 2.48924
R9312 VDD.n1914 VDD.n1913 2.48924
R9313 VDD.n1911 VDD.n1910 2.48924
R9314 VDD.n1908 VDD.n1907 2.48924
R9315 VDD.n1905 VDD.n1904 2.48924
R9316 VDD.n1902 VDD.n1901 2.48924
R9317 VDD.n1899 VDD.n1898 2.48924
R9318 VDD.n1896 VDD.n1895 2.48924
R9319 VDD.n1893 VDD.n1892 2.48924
R9320 VDD.n1890 VDD.n1889 2.48924
R9321 VDD.n1887 VDD.n1886 2.48924
R9322 VDD.n1884 VDD.n1883 2.48924
R9323 VDD.n1881 VDD.n1880 2.48924
R9324 VDD.n1878 VDD.n1877 2.48924
R9325 VDD.n1875 VDD.n1874 2.48924
R9326 VDD.n1872 VDD.n1871 2.48924
R9327 VDD.n1869 VDD.n1868 2.48924
R9328 VDD.n1866 VDD.n1865 2.48924
R9329 VDD.n1863 VDD.n1862 2.48924
R9330 VDD.n1860 VDD.n1859 2.48924
R9331 VDD.n1857 VDD.n1856 2.48924
R9332 VDD.n1854 VDD.n1853 2.48924
R9333 VDD.n1851 VDD.n1850 2.48924
R9334 VDD.n1848 VDD.n1847 2.48924
R9335 VDD.n1845 VDD.n1844 2.48924
R9336 VDD.n1842 VDD.n1841 2.48924
R9337 VDD.n1839 VDD.n1838 2.48924
R9338 VDD.n1836 VDD.n1835 2.48924
R9339 VDD.n1833 VDD.n1832 2.48924
R9340 VDD.n1830 VDD.n1829 2.48924
R9341 VDD.n1827 VDD.n1826 2.48924
R9342 VDD.n1824 VDD.n1823 2.48924
R9343 VDD.n1821 VDD.n1820 2.48924
R9344 VDD.n1818 VDD.n1817 2.48924
R9345 VDD.n7720 VDD.t522 2.4382
R9346 VDD.n1056 VDD.t354 2.42448
R9347 VDD.n1089 VDD.t102 2.42448
R9348 VDD.t753 VDD.t1066 2.31934
R9349 VDD.t750 VDD.t767 2.31934
R9350 VDD.t695 VDD.t324 2.31934
R9351 VDD.t772 VDD.t189 2.31934
R9352 VDD.t1101 VDD.t1377 2.31934
R9353 VDD.n2267 VDD.t766 2.2583
R9354 VDD.n2371 VDD.t1270 2.2583
R9355 VDD.n2502 VDD.t1279 2.2583
R9356 VDD.n18 VDD.n17 2.21137
R9357 VDD.n17 VDD.n16 2.21137
R9358 VDD.n288 VDD.n287 2.21137
R9359 VDD.n21 VDD.n20 2.21137
R9360 VDD.n20 VDD.n19 2.21137
R9361 VDD.n6880 VDD.n6879 2.21137
R9362 VDD.n24 VDD.n23 2.21137
R9363 VDD.n23 VDD.n22 2.21137
R9364 VDD.n6886 VDD.n6885 2.21137
R9365 VDD.n181 VDD.n180 2.21137
R9366 VDD.n180 VDD.n179 2.21137
R9367 VDD.n294 VDD.n293 2.21137
R9368 VDD.n3315 VDD.n3314 2.07441
R9369 VDD.n5427 VDD.n5424 2.07441
R9370 VDD.n3309 VDD.n3308 2.07441
R9371 VDD.n5421 VDD.n5418 2.07441
R9372 VDD.n3303 VDD.n3302 2.07441
R9373 VDD.n5415 VDD.n5412 2.07441
R9374 VDD.n3285 VDD.n3284 2.07441
R9375 VDD.n5387 VDD.n5384 2.07441
R9376 VDD.n3279 VDD.n3278 2.07441
R9377 VDD.n5381 VDD.n5378 2.07441
R9378 VDD.n2920 VDD.n2919 2.07441
R9379 VDD.n4079 VDD.n4076 2.07441
R9380 VDD.n2926 VDD.n2925 2.07441
R9381 VDD.n4085 VDD.n4082 2.07441
R9382 VDD.n2932 VDD.n2931 2.07441
R9383 VDD.n4091 VDD.n4088 2.07441
R9384 VDD.n2950 VDD.n2949 2.07441
R9385 VDD.n4119 VDD.n4116 2.07441
R9386 VDD.n2956 VDD.n2955 2.07441
R9387 VDD.n4125 VDD.n4122 2.07441
R9388 VDD.n2990 VDD.n2989 2.07441
R9389 VDD.n4399 VDD.n4396 2.07441
R9390 VDD.n2996 VDD.n2995 2.07441
R9391 VDD.n4405 VDD.n4402 2.07441
R9392 VDD.n3014 VDD.n3013 2.07441
R9393 VDD.n4433 VDD.n4430 2.07441
R9394 VDD.n3020 VDD.n3019 2.07441
R9395 VDD.n4439 VDD.n4436 2.07441
R9396 VDD.n3026 VDD.n3025 2.07441
R9397 VDD.n4445 VDD.n4442 2.07441
R9398 VDD.n3050 VDD.n3049 2.07441
R9399 VDD.n4589 VDD.n4586 2.07441
R9400 VDD.n3056 VDD.n3055 2.07441
R9401 VDD.n4595 VDD.n4592 2.07441
R9402 VDD.n3062 VDD.n3061 2.07441
R9403 VDD.n4601 VDD.n4598 2.07441
R9404 VDD.n3080 VDD.n3079 2.07441
R9405 VDD.n4629 VDD.n4626 2.07441
R9406 VDD.n3086 VDD.n3085 2.07441
R9407 VDD.n4635 VDD.n4632 2.07441
R9408 VDD.n3126 VDD.n3125 2.07441
R9409 VDD.n4903 VDD.n4900 2.07441
R9410 VDD.n3132 VDD.n3131 2.07441
R9411 VDD.n4909 VDD.n4906 2.07441
R9412 VDD.n3150 VDD.n3149 2.07441
R9413 VDD.n4937 VDD.n4934 2.07441
R9414 VDD.n3156 VDD.n3155 2.07441
R9415 VDD.n4943 VDD.n4940 2.07441
R9416 VDD.n3162 VDD.n3161 2.07441
R9417 VDD.n4949 VDD.n4946 2.07441
R9418 VDD.n3231 VDD.n3230 2.07441
R9419 VDD.n5135 VDD.n5132 2.07441
R9420 VDD.n3225 VDD.n3224 2.07441
R9421 VDD.n5129 VDD.n5126 2.07441
R9422 VDD.n3207 VDD.n3206 2.07441
R9423 VDD.n5101 VDD.n5098 2.07441
R9424 VDD.n3201 VDD.n3200 2.07441
R9425 VDD.n5095 VDD.n5092 2.07441
R9426 VDD.n3195 VDD.n3194 2.07441
R9427 VDD.n5089 VDD.n5086 2.07441
R9428 VDD.n2550 VDD.n2549 2.07441
R9429 VDD.n2850 VDD.n2847 2.07441
R9430 VDD.n2556 VDD.n2555 2.07441
R9431 VDD.n2856 VDD.n2853 2.07441
R9432 VDD.n2574 VDD.n2573 2.07441
R9433 VDD.n2884 VDD.n2881 2.07441
R9434 VDD.n2580 VDD.n2579 2.07441
R9435 VDD.n2890 VDD.n2887 2.07441
R9436 VDD.n2586 VDD.n2585 2.07441
R9437 VDD.n2896 VDD.n2893 2.07441
R9438 VDD.n548 VDD.n547 2.02746
R9439 VDD.n780 VDD.n779 2.02746
R9440 VDD.n786 VDD.n785 2.02746
R9441 VDD.n794 VDD.n793 2.02746
R9442 VDD.n793 VDD.n792 2.02746
R9443 VDD.n798 VDD.n797 2.02746
R9444 VDD.n797 VDD.n796 2.02746
R9445 VDD.n977 VDD.n974 2.02746
R9446 VDD.n980 VDD.n977 2.02746
R9447 VDD.n986 VDD.n983 2.02746
R9448 VDD.n989 VDD.n986 2.02746
R9449 VDD.n6829 VDD.n6826 2.02746
R9450 VDD.n6832 VDD.n6829 2.02746
R9451 VDD.n6820 VDD.n6817 2.02746
R9452 VDD.n6823 VDD.n6820 2.02746
R9453 VDD.n6812 VDD.n6811 2.02746
R9454 VDD.n6808 VDD.n6807 2.02746
R9455 VDD.n554 VDD.n553 2.02746
R9456 VDD.n2487 VDD.n1372 1.9805
R9457 VDD.n2477 VDD.n1383 1.9805
R9458 VDD.n2463 VDD.n1394 1.9805
R9459 VDD.n2452 VDD.n1405 1.9805
R9460 VDD.n2442 VDD.n1416 1.9805
R9461 VDD.n2428 VDD.n1427 1.9805
R9462 VDD.n2393 VDD.n1446 1.9805
R9463 VDD.n2370 VDD.n1461 1.9805
R9464 VDD.n2374 VDD.n1458 1.9805
R9465 VDD.n1152 VDD.n1139 1.9805
R9466 VDD.n1155 VDD.n1136 1.9805
R9467 VDD.n2382 VDD.n1453 1.9805
R9468 VDD.n2389 VDD.n1450 1.9805
R9469 VDD.n2404 VDD.n1439 1.9805
R9470 VDD.n1173 VDD.n1127 1.9805
R9471 VDD.n2418 VDD.n1433 1.9805
R9472 VDD.n1182 VDD.n1121 1.9805
R9473 VDD.n2501 VDD.n1361 1.9805
R9474 VDD.n2505 VDD.n1356 1.9805
R9475 VDD.n1231 VDD.n1115 1.9805
R9476 VDD.n1234 VDD.n1110 1.9805
R9477 VDD.n7234 VDD.n7226 1.90688
R9478 VDD.n7234 VDD.n7227 1.90688
R9479 VDD.n7234 VDD.n7228 1.90688
R9480 VDD.n7234 VDD.n7229 1.90688
R9481 VDD.n7234 VDD.n7230 1.90688
R9482 VDD.n7234 VDD.n7231 1.90688
R9483 VDD.n7234 VDD.n7232 1.90688
R9484 VDD.n7234 VDD.n7233 1.90688
R9485 VDD.n6997 VDD.n6987 1.90688
R9486 VDD.n6997 VDD.n6988 1.90688
R9487 VDD.n6997 VDD.n6989 1.90688
R9488 VDD.n6997 VDD.n6990 1.90688
R9489 VDD.n6997 VDD.n6991 1.90688
R9490 VDD.n6997 VDD.n6992 1.90688
R9491 VDD.n6997 VDD.n6993 1.90688
R9492 VDD.n6997 VDD.n6994 1.90688
R9493 VDD.n6997 VDD.n6995 1.90688
R9494 VDD.n772 VDD.n753 1.90688
R9495 VDD.n772 VDD.n754 1.90688
R9496 VDD.n772 VDD.n755 1.90688
R9497 VDD.n772 VDD.n756 1.90688
R9498 VDD.n772 VDD.n757 1.90688
R9499 VDD.n772 VDD.n758 1.90688
R9500 VDD.n772 VDD.n759 1.90688
R9501 VDD.n772 VDD.n760 1.90688
R9502 VDD.n772 VDD.n761 1.90688
R9503 VDD.n772 VDD.n762 1.90688
R9504 VDD.n772 VDD.n763 1.90688
R9505 VDD.n772 VDD.n764 1.90688
R9506 VDD.n772 VDD.n765 1.90688
R9507 VDD.n772 VDD.n766 1.90688
R9508 VDD.n772 VDD.n767 1.90688
R9509 VDD.n772 VDD.n768 1.90688
R9510 VDD.n772 VDD.n769 1.90688
R9511 VDD.n772 VDD.n770 1.90688
R9512 VDD.n968 VDD.n949 1.90688
R9513 VDD.n968 VDD.n950 1.90688
R9514 VDD.n968 VDD.n951 1.90688
R9515 VDD.n968 VDD.n952 1.90688
R9516 VDD.n968 VDD.n953 1.90688
R9517 VDD.n968 VDD.n954 1.90688
R9518 VDD.n968 VDD.n955 1.90688
R9519 VDD.n968 VDD.n956 1.90688
R9520 VDD.n968 VDD.n957 1.90688
R9521 VDD.n968 VDD.n958 1.90688
R9522 VDD.n968 VDD.n959 1.90688
R9523 VDD.n968 VDD.n960 1.90688
R9524 VDD.n968 VDD.n961 1.90688
R9525 VDD.n968 VDD.n962 1.90688
R9526 VDD.n968 VDD.n963 1.90688
R9527 VDD.n968 VDD.n964 1.90688
R9528 VDD.n968 VDD.n965 1.90688
R9529 VDD.n2347 VDD.n2345 1.90688
R9530 VDD.n2347 VDD.n2346 1.90688
R9531 VDD.n2156 VDD.n2154 1.90688
R9532 VDD.n2156 VDD.n2155 1.90688
R9533 VDD.n1160 VDD.n1131 1.88267
R9534 VDD.n2258 VDD.t580 1.84779
R9535 VDD.n7667 VDD.n7666 1.7854
R9536 VDD.n7662 VDD.n7661 1.7854
R9537 VDD.n7657 VDD.n7656 1.7854
R9538 VDD.n7652 VDD.n7651 1.7854
R9539 VDD.n7647 VDD.n7646 1.7854
R9540 VDD.n7642 VDD.n7641 1.7854
R9541 VDD.n7637 VDD.n7636 1.7854
R9542 VDD.n7632 VDD.n7631 1.7854
R9543 VDD.n285 VDD.n284 1.7854
R9544 VDD.n531 VDD.n530 1.7854
R9545 VDD.n526 VDD.n525 1.7854
R9546 VDD.n521 VDD.n520 1.7854
R9547 VDD.n516 VDD.n515 1.7854
R9548 VDD.n511 VDD.n510 1.7854
R9549 VDD.n506 VDD.n505 1.7854
R9550 VDD.n501 VDD.n500 1.7854
R9551 VDD.n496 VDD.n495 1.7854
R9552 VDD.n491 VDD.n490 1.7854
R9553 VDD.n486 VDD.n485 1.7854
R9554 VDD.n481 VDD.n480 1.7854
R9555 VDD.n970 VDD.n969 1.7854
R9556 VDD.n3332 VDD.n3331 1.7854
R9557 VDD.n3327 VDD.n3326 1.7854
R9558 VDD.n2909 VDD.n2907 1.7854
R9559 VDD.n4268 VDD.n4267 1.7854
R9560 VDD.n4775 VDD.n4774 1.7854
R9561 VDD.n5270 VDD.n5269 1.7854
R9562 VDD.n2036 VDD.n2035 1.7854
R9563 VDD.n2031 VDD.n2030 1.7854
R9564 VDD.n2026 VDD.n2025 1.7854
R9565 VDD.n2021 VDD.n2020 1.7854
R9566 VDD.n2016 VDD.n2015 1.7854
R9567 VDD.n2011 VDD.n2010 1.7854
R9568 VDD.n2006 VDD.n2005 1.7854
R9569 VDD.n2001 VDD.n2000 1.7854
R9570 VDD.n1996 VDD.n1995 1.7854
R9571 VDD.n1991 VDD.n1990 1.7854
R9572 VDD.n271 VDD.n270 1.78487
R9573 VDD.n266 VDD.n265 1.78487
R9574 VDD.n261 VDD.n260 1.78487
R9575 VDD.n256 VDD.n255 1.78487
R9576 VDD.n251 VDD.n250 1.78487
R9577 VDD.n246 VDD.n245 1.78487
R9578 VDD.n241 VDD.n240 1.78487
R9579 VDD.n236 VDD.n235 1.78487
R9580 VDD.n231 VDD.n230 1.78487
R9581 VDD.n5436 VDD.n5435 1.78487
R9582 VDD.n5441 VDD.n5440 1.78487
R9583 VDD.n5446 VDD.n5445 1.78487
R9584 VDD.n5451 VDD.n5450 1.78487
R9585 VDD.n5456 VDD.n5455 1.78487
R9586 VDD.n5461 VDD.n5460 1.78487
R9587 VDD.n5466 VDD.n5465 1.78487
R9588 VDD.n5471 VDD.n5470 1.78487
R9589 VDD.n5476 VDD.n5475 1.78487
R9590 VDD.n5481 VDD.n5480 1.78487
R9591 VDD.n5486 VDD.n5485 1.78487
R9592 VDD.n5491 VDD.n5490 1.78487
R9593 VDD.n5496 VDD.n5495 1.78487
R9594 VDD.n5501 VDD.n5500 1.78487
R9595 VDD.n5506 VDD.n5505 1.78487
R9596 VDD.n5511 VDD.n5510 1.78487
R9597 VDD.n5516 VDD.n5515 1.78487
R9598 VDD.n5521 VDD.n5520 1.78487
R9599 VDD.n5526 VDD.n5525 1.78487
R9600 VDD.n5531 VDD.n5530 1.78487
R9601 VDD.n4376 VDD.n4375 1.78487
R9602 VDD.n4371 VDD.n4370 1.78487
R9603 VDD.n4366 VDD.n4365 1.78487
R9604 VDD.n4361 VDD.n4360 1.78487
R9605 VDD.n4356 VDD.n4355 1.78487
R9606 VDD.n4351 VDD.n4350 1.78487
R9607 VDD.n4346 VDD.n4345 1.78487
R9608 VDD.n4341 VDD.n4340 1.78487
R9609 VDD.n4336 VDD.n4335 1.78487
R9610 VDD.n4331 VDD.n4330 1.78487
R9611 VDD.n4326 VDD.n4325 1.78487
R9612 VDD.n4321 VDD.n4320 1.78487
R9613 VDD.n4316 VDD.n4315 1.78487
R9614 VDD.n4311 VDD.n4310 1.78487
R9615 VDD.n4306 VDD.n4305 1.78487
R9616 VDD.n4301 VDD.n4300 1.78487
R9617 VDD.n4296 VDD.n4295 1.78487
R9618 VDD.n4291 VDD.n4290 1.78487
R9619 VDD.n4286 VDD.n4285 1.78487
R9620 VDD.n4281 VDD.n4280 1.78487
R9621 VDD.n4276 VDD.n4275 1.78487
R9622 VDD.n2909 VDD.n2908 1.78487
R9623 VDD.n4880 VDD.n4879 1.78487
R9624 VDD.n4875 VDD.n4874 1.78487
R9625 VDD.n4870 VDD.n4869 1.78487
R9626 VDD.n4865 VDD.n4864 1.78487
R9627 VDD.n4860 VDD.n4859 1.78487
R9628 VDD.n4855 VDD.n4854 1.78487
R9629 VDD.n4850 VDD.n4849 1.78487
R9630 VDD.n4845 VDD.n4844 1.78487
R9631 VDD.n4840 VDD.n4839 1.78487
R9632 VDD.n4835 VDD.n4834 1.78487
R9633 VDD.n4830 VDD.n4829 1.78487
R9634 VDD.n4825 VDD.n4824 1.78487
R9635 VDD.n4820 VDD.n4819 1.78487
R9636 VDD.n4815 VDD.n4814 1.78487
R9637 VDD.n4810 VDD.n4809 1.78487
R9638 VDD.n4805 VDD.n4804 1.78487
R9639 VDD.n4800 VDD.n4799 1.78487
R9640 VDD.n4795 VDD.n4794 1.78487
R9641 VDD.n4790 VDD.n4789 1.78487
R9642 VDD.n4785 VDD.n4784 1.78487
R9643 VDD.n4780 VDD.n4779 1.78487
R9644 VDD.n100 VDD.n99 1.78473
R9645 VDD.n95 VDD.n94 1.78473
R9646 VDD.n90 VDD.n89 1.78473
R9647 VDD.n85 VDD.n84 1.78473
R9648 VDD.n80 VDD.n79 1.78473
R9649 VDD.n75 VDD.n74 1.78473
R9650 VDD.n70 VDD.n69 1.78473
R9651 VDD.n7450 VDD.n7449 1.78473
R9652 VDD.n7455 VDD.n7454 1.78473
R9653 VDD.n7460 VDD.n7459 1.78473
R9654 VDD.n7465 VDD.n7464 1.78473
R9655 VDD.n7470 VDD.n7469 1.78473
R9656 VDD.n7475 VDD.n7474 1.78473
R9657 VDD.n7480 VDD.n7479 1.78473
R9658 VDD.n7485 VDD.n7484 1.78473
R9659 VDD.n7490 VDD.n7489 1.78473
R9660 VDD.n7495 VDD.n7494 1.78473
R9661 VDD.n7500 VDD.n7499 1.78473
R9662 VDD.n6747 VDD.n6746 1.78473
R9663 VDD.n6752 VDD.n6751 1.78473
R9664 VDD.n6757 VDD.n6756 1.78473
R9665 VDD.n6762 VDD.n6761 1.78473
R9666 VDD.n6767 VDD.n6766 1.78473
R9667 VDD.n6772 VDD.n6771 1.78473
R9668 VDD.n6777 VDD.n6776 1.78473
R9669 VDD.n6782 VDD.n6781 1.78473
R9670 VDD.n5364 VDD.n5363 1.78473
R9671 VDD.n5359 VDD.n5358 1.78473
R9672 VDD.n5354 VDD.n5353 1.78473
R9673 VDD.n5349 VDD.n5348 1.78473
R9674 VDD.n5344 VDD.n5343 1.78473
R9675 VDD.n5339 VDD.n5338 1.78473
R9676 VDD.n5334 VDD.n5333 1.78473
R9677 VDD.n5329 VDD.n5328 1.78473
R9678 VDD.n5324 VDD.n5323 1.78473
R9679 VDD.n4574 VDD.n4573 1.78473
R9680 VDD.n4569 VDD.n4568 1.78473
R9681 VDD.n4564 VDD.n4563 1.78473
R9682 VDD.n4559 VDD.n4558 1.78473
R9683 VDD.n4554 VDD.n4553 1.78473
R9684 VDD.n4549 VDD.n4548 1.78473
R9685 VDD.n4544 VDD.n4543 1.78473
R9686 VDD.n4539 VDD.n4538 1.78473
R9687 VDD.n4534 VDD.n4533 1.78473
R9688 VDD.n4529 VDD.n4528 1.78473
R9689 VDD.n4524 VDD.n4523 1.78473
R9690 VDD.n4519 VDD.n4518 1.78473
R9691 VDD.n4514 VDD.n4513 1.78473
R9692 VDD.n4509 VDD.n4508 1.78473
R9693 VDD.n4504 VDD.n4503 1.78473
R9694 VDD.n4499 VDD.n4498 1.78473
R9695 VDD.n4494 VDD.n4493 1.78473
R9696 VDD.n4489 VDD.n4488 1.78473
R9697 VDD.n4484 VDD.n4483 1.78473
R9698 VDD.n4479 VDD.n4478 1.78473
R9699 VDD.n4474 VDD.n4473 1.78473
R9700 VDD.n4469 VDD.n4468 1.78473
R9701 VDD.n4464 VDD.n4463 1.78473
R9702 VDD.n4459 VDD.n4458 1.78473
R9703 VDD.n3039 VDD.n3036 1.78473
R9704 VDD.n3039 VDD.n3038 1.78473
R9705 VDD.n4062 VDD.n4061 1.78473
R9706 VDD.n4057 VDD.n4056 1.78473
R9707 VDD.n4052 VDD.n4051 1.78473
R9708 VDD.n4047 VDD.n4046 1.78473
R9709 VDD.n4042 VDD.n4041 1.78473
R9710 VDD.n4037 VDD.n4036 1.78473
R9711 VDD.n4032 VDD.n4031 1.78473
R9712 VDD.n4027 VDD.n4026 1.78473
R9713 VDD.n4022 VDD.n4021 1.78473
R9714 VDD.n4017 VDD.n4016 1.78473
R9715 VDD.n6479 VDD.n6461 1.78473
R9716 VDD.n6479 VDD.n6478 1.78473
R9717 VDD.n5074 VDD.n5073 1.78473
R9718 VDD.n5069 VDD.n5068 1.78473
R9719 VDD.n5064 VDD.n5063 1.78473
R9720 VDD.n5059 VDD.n5058 1.78473
R9721 VDD.n5054 VDD.n5053 1.78473
R9722 VDD.n5049 VDD.n5048 1.78473
R9723 VDD.n5044 VDD.n5043 1.78473
R9724 VDD.n5039 VDD.n5038 1.78473
R9725 VDD.n5034 VDD.n5033 1.78473
R9726 VDD.n5029 VDD.n5028 1.78473
R9727 VDD.n5024 VDD.n5023 1.78473
R9728 VDD.n5019 VDD.n5018 1.78473
R9729 VDD.n5014 VDD.n5013 1.78473
R9730 VDD.n5009 VDD.n5008 1.78473
R9731 VDD.n5004 VDD.n5003 1.78473
R9732 VDD.n4999 VDD.n4998 1.78473
R9733 VDD.n4994 VDD.n4993 1.78473
R9734 VDD.n4989 VDD.n4988 1.78473
R9735 VDD.n4984 VDD.n4983 1.78473
R9736 VDD.n4979 VDD.n4978 1.78473
R9737 VDD.n4974 VDD.n4973 1.78473
R9738 VDD.n4969 VDD.n4968 1.78473
R9739 VDD.n4964 VDD.n4963 1.78473
R9740 VDD.n4959 VDD.n4958 1.78473
R9741 VDD.n3175 VDD.n3172 1.78473
R9742 VDD.n3175 VDD.n3174 1.78473
R9743 VDD.n1304 VDD.n1303 1.78473
R9744 VDD.n1309 VDD.n1308 1.78473
R9745 VDD.n1314 VDD.n1313 1.78473
R9746 VDD.n1319 VDD.n1318 1.78473
R9747 VDD.n1324 VDD.n1323 1.78473
R9748 VDD.n1329 VDD.n1328 1.78473
R9749 VDD.n1334 VDD.n1333 1.78473
R9750 VDD.n1339 VDD.n1338 1.78473
R9751 VDD.n1344 VDD.n1343 1.78473
R9752 VDD.n1349 VDD.n1348 1.78473
R9753 VDD.n389 VDD.n388 1.78093
R9754 VDD.n404 VDD.n401 1.78093
R9755 VDD.n6638 VDD.n6637 1.61319
R9756 VDD.n7368 VDD.n7367 1.54224
R9757 VDD.n7374 VDD.n7373 1.52463
R9758 VDD.n7378 VDD.n7377 1.52463
R9759 VDD.n7085 VDD.n7082 1.49137
R9760 VDD.n7088 VDD.n7085 1.49137
R9761 VDD.n7545 VDD.n7542 1.49137
R9762 VDD.n7548 VDD.n7545 1.49137
R9763 VDD.n7312 VDD.n7309 1.49137
R9764 VDD.n7315 VDD.n7312 1.49137
R9765 VDD.n7301 VDD.n7300 1.49137
R9766 VDD.n7300 VDD.n7299 1.49137
R9767 VDD.n7297 VDD.n7296 1.49137
R9768 VDD.n7296 VDD.n7295 1.49137
R9769 VDD.n11 VDD.n10 1.49137
R9770 VDD.n10 VDD.n9 1.49137
R9771 VDD.n15 VDD.n14 1.49137
R9772 VDD.n14 VDD.n13 1.49137
R9773 VDD.n2968 VDD.n2967 1.467
R9774 VDD.n3101 VDD.n3100 1.467
R9775 VDD.n3251 VDD.n3250 1.467
R9776 VDD.n1794 VDD.n1793 1.467
R9777 VDD.n1932 VDD.n1931 1.467
R9778 VDD.n6999 VDD.n6998 1.46684
R9779 VDD.n774 VDD.n773 1.46684
R9780 VDD.n945 VDD.n944 1.46684
R9781 VDD.n2835 VDD.n2834 1.46684
R9782 VDD.n5534 VDD.n5533 1.46684
R9783 VDD.n5539 VDD.n5538 1.46684
R9784 VDD.n4271 VDD.n4270 1.46684
R9785 VDD.n4379 VDD.n4378 1.46684
R9786 VDD.n4384 VDD.n4383 1.46684
R9787 VDD.n4263 VDD.n4262 1.46684
R9788 VDD.n4770 VDD.n4769 1.46684
R9789 VDD.n3106 VDD.n3105 1.46684
R9790 VDD.n4883 VDD.n4882 1.46684
R9791 VDD.n4888 VDD.n4887 1.46684
R9792 VDD.n5265 VDD.n5264 1.46684
R9793 VDD.n1809 VDD.n1808 1.46684
R9794 VDD.n1671 VDD.n1670 1.46684
R9795 VDD.n7338 VDD.t652 1.44978
R9796 VDD.n1372 VDD.n1371 1.4405
R9797 VDD.n1371 VDD.n1370 1.4405
R9798 VDD.n1383 VDD.n1382 1.4405
R9799 VDD.n1382 VDD.n1381 1.4405
R9800 VDD.n1394 VDD.n1393 1.4405
R9801 VDD.n1393 VDD.n1392 1.4405
R9802 VDD.n1405 VDD.n1404 1.4405
R9803 VDD.n1404 VDD.n1403 1.4405
R9804 VDD.n1416 VDD.n1415 1.4405
R9805 VDD.n1415 VDD.n1414 1.4405
R9806 VDD.n1427 VDD.n1426 1.4405
R9807 VDD.n1426 VDD.n1425 1.4405
R9808 VDD.n1446 VDD.n1445 1.4405
R9809 VDD.n1445 VDD.n1444 1.4405
R9810 VDD.n1131 VDD.n1129 1.4405
R9811 VDD.n1439 VDD.n1438 1.4405
R9812 VDD.n1127 VDD.n1124 1.4405
R9813 VDD.n1433 VDD.n1432 1.4405
R9814 VDD.n1121 VDD.n1118 1.4405
R9815 VDD.n146 VDD.t353 1.43811
R9816 VDD.n161 VDD.t166 1.43811
R9817 VDD.n2478 VDD.t186 1.43728
R9818 VDD.n456 VDD.n455 1.40703
R9819 VDD.n5708 VDD.n5691 1.40703
R9820 VDD.n6318 VDD.n6317 1.40703
R9821 VDD.n5544 VDD.n5541 1.40703
R9822 VDD.n5714 VDD.n5713 1.40703
R9823 VDD.n3338 VDD.n3336 1.40703
R9824 VDD.n3439 VDD.n3437 1.40703
R9825 VDD.n1249 VDD.n1247 1.40703
R9826 VDD.n1663 VDD.n1661 1.40703
R9827 VDD.n1535 VDD.n1533 1.40703
R9828 VDD.n2349 VDD.n2343 1.40703
R9829 VDD.n2158 VDD.n2152 1.40703
R9830 VDD.n2055 VDD.n2040 1.40703
R9831 VDD.n2540 VDD.n2525 1.40703
R9832 VDD.n542 VDD.n541 1.40656
R9833 VDD.n3849 VDD.n3847 1.40656
R9834 VDD.n3644 VDD.n3642 1.40656
R9835 VDD.n6015 VDD.n6014 1.40656
R9836 VDD.n5544 VDD.n5543 1.40656
R9837 VDD.n3443 VDD.n3441 1.40656
R9838 VDD.n2692 VDD.n2690 1.40656
R9839 VDD.n1535 VDD.n1534 1.40656
R9840 VDD.n1663 VDD.n1662 1.40656
R9841 VDD.n1467 VDD.n1466 1.40656
R9842 VDD.n7683 VDD.n7682 1.40656
R9843 VDD.n118 VDD.n117 1.40638
R9844 VDD.n7511 VDD.n7510 1.40638
R9845 VDD.n7425 VDD.n7424 1.40638
R9846 VDD.n6803 VDD.n6802 1.40638
R9847 VDD.n6625 VDD.n6624 1.40638
R9848 VDD.n3038 VDD.n3037 1.40638
R9849 VDD.n2907 VDD.n2906 1.40638
R9850 VDD.n6478 VDD.n6477 1.40638
R9851 VDD.n6163 VDD.n6162 1.40638
R9852 VDD.n6311 VDD.n6310 1.40638
R9853 VDD.n3174 VDD.n3173 1.40638
R9854 VDD.n5862 VDD.n5861 1.40638
R9855 VDD.n6009 VDD.n6008 1.40638
R9856 VDD.n772 VDD.n771 1.36744
R9857 VDD.n7235 VDD.n7234 1.36744
R9858 VDD.n7031 VDD.t37 1.35478
R9859 VDD.n7047 VDD.t530 1.35478
R9860 VDD.n7059 VDD.n386 1.33475
R9861 VDD.n7559 VDD.n7537 1.33475
R9862 VDD.n3296 VDD.n3295 1.31137
R9863 VDD.n5396 VDD.n5393 1.31137
R9864 VDD.n5405 VDD.n5402 1.31137
R9865 VDD.n4113 VDD.n4110 1.31137
R9866 VDD.n4109 VDD.n4106 1.31137
R9867 VDD.n2943 VDD.n2937 1.31137
R9868 VDD.n4423 VDD.n4420 1.31137
R9869 VDD.n4419 VDD.n4416 1.31137
R9870 VDD.n3007 VDD.n3001 1.31137
R9871 VDD.n4623 VDD.n4620 1.31137
R9872 VDD.n4619 VDD.n4616 1.31137
R9873 VDD.n3073 VDD.n3067 1.31137
R9874 VDD.n4927 VDD.n4924 1.31137
R9875 VDD.n4923 VDD.n4920 1.31137
R9876 VDD.n3143 VDD.n3137 1.31137
R9877 VDD.n3218 VDD.n3217 1.31137
R9878 VDD.n5114 VDD.n5111 1.31137
R9879 VDD.n5123 VDD.n5120 1.31137
R9880 VDD.n2874 VDD.n2871 1.31137
R9881 VDD.n2870 VDD.n2867 1.31137
R9882 VDD.n2567 VDD.n2561 1.31137
R9883 VDD.n6875 VDD.n6874 1.30325
R9884 VDD.n189 VDD.n18 1.23311
R9885 VDD.n130 VDD.n21 1.23311
R9886 VDD.n123 VDD.n24 1.23311
R9887 VDD.n182 VDD.n181 1.23311
R9888 VDD.n5571 VDD.n5432 1.23311
R9889 VDD.n3362 VDD.n3315 1.23311
R9890 VDD.n5581 VDD.n5427 1.23311
R9891 VDD.n3369 VDD.n3309 1.23311
R9892 VDD.n5591 VDD.n5421 1.23311
R9893 VDD.n3376 VDD.n3303 1.23311
R9894 VDD.n5601 VDD.n5415 1.23311
R9895 VDD.n3399 VDD.n3297 1.23311
R9896 VDD.n5637 VDD.n5405 1.23311
R9897 VDD.n3406 VDD.n3285 1.23311
R9898 VDD.n5647 VDD.n5387 1.23311
R9899 VDD.n3413 VDD.n3279 1.23311
R9900 VDD.n5657 VDD.n5381 1.23311
R9901 VDD.n3420 VDD.n3273 1.23311
R9902 VDD.n3425 VDD.n3270 1.23311
R9903 VDD.n5667 VDD.n5375 1.23311
R9904 VDD.n5674 VDD.n5372 1.23311
R9905 VDD.n3932 VDD.n2914 1.23311
R9906 VDD.n3925 VDD.n2920 1.23311
R9907 VDD.n6430 VDD.n4079 1.23311
R9908 VDD.n3918 VDD.n2926 1.23311
R9909 VDD.n6420 VDD.n4085 1.23311
R9910 VDD.n3911 VDD.n2932 1.23311
R9911 VDD.n6410 VDD.n4091 1.23311
R9912 VDD.n6374 VDD.n4113 1.23311
R9913 VDD.n3888 VDD.n2944 1.23311
R9914 VDD.n3881 VDD.n2950 1.23311
R9915 VDD.n6364 VDD.n4119 1.23311
R9916 VDD.n3874 VDD.n2956 1.23311
R9917 VDD.n6354 VDD.n4125 1.23311
R9918 VDD.n6344 VDD.n4130 1.23311
R9919 VDD.n6337 VDD.n4133 1.23311
R9920 VDD.n3867 VDD.n2961 1.23311
R9921 VDD.n3862 VDD.n2964 1.23311
R9922 VDD.n6292 VDD.n4390 1.23311
R9923 VDD.n6285 VDD.n4393 1.23311
R9924 VDD.n3830 VDD.n2981 1.23311
R9925 VDD.n3825 VDD.n2984 1.23311
R9926 VDD.n3818 VDD.n2990 1.23311
R9927 VDD.n6275 VDD.n4399 1.23311
R9928 VDD.n3811 VDD.n2996 1.23311
R9929 VDD.n6265 VDD.n4405 1.23311
R9930 VDD.n6255 VDD.n4423 1.23311
R9931 VDD.n3804 VDD.n3008 1.23311
R9932 VDD.n3781 VDD.n3014 1.23311
R9933 VDD.n6219 VDD.n4433 1.23311
R9934 VDD.n3774 VDD.n3020 1.23311
R9935 VDD.n6209 VDD.n4439 1.23311
R9936 VDD.n3767 VDD.n3026 1.23311
R9937 VDD.n6199 VDD.n4445 1.23311
R9938 VDD.n6189 VDD.n4450 1.23311
R9939 VDD.n6182 VDD.n4453 1.23311
R9940 VDD.n3760 VDD.n3031 1.23311
R9941 VDD.n3755 VDD.n3034 1.23311
R9942 VDD.n3942 VDD.n3941 1.23311
R9943 VDD.n6440 VDD.n4073 1.23311
R9944 VDD.n6447 VDD.n4070 1.23311
R9945 VDD.n3727 VDD.n3044 1.23311
R9946 VDD.n3720 VDD.n3050 1.23311
R9947 VDD.n6128 VDD.n4589 1.23311
R9948 VDD.n3713 VDD.n3056 1.23311
R9949 VDD.n6118 VDD.n4595 1.23311
R9950 VDD.n3706 VDD.n3062 1.23311
R9951 VDD.n6108 VDD.n4601 1.23311
R9952 VDD.n6072 VDD.n4623 1.23311
R9953 VDD.n3683 VDD.n3074 1.23311
R9954 VDD.n3676 VDD.n3080 1.23311
R9955 VDD.n6062 VDD.n4629 1.23311
R9956 VDD.n3669 VDD.n3086 1.23311
R9957 VDD.n6052 VDD.n4635 1.23311
R9958 VDD.n6042 VDD.n4640 1.23311
R9959 VDD.n6035 VDD.n4643 1.23311
R9960 VDD.n3662 VDD.n3091 1.23311
R9961 VDD.n3657 VDD.n3094 1.23311
R9962 VDD.n5990 VDD.n4894 1.23311
R9963 VDD.n5983 VDD.n4897 1.23311
R9964 VDD.n3624 VDD.n3117 1.23311
R9965 VDD.n3619 VDD.n3120 1.23311
R9966 VDD.n3612 VDD.n3126 1.23311
R9967 VDD.n5973 VDD.n4903 1.23311
R9968 VDD.n3605 VDD.n3132 1.23311
R9969 VDD.n5963 VDD.n4909 1.23311
R9970 VDD.n5953 VDD.n4927 1.23311
R9971 VDD.n3598 VDD.n3144 1.23311
R9972 VDD.n3575 VDD.n3150 1.23311
R9973 VDD.n5917 VDD.n4937 1.23311
R9974 VDD.n3568 VDD.n3156 1.23311
R9975 VDD.n5907 VDD.n4943 1.23311
R9976 VDD.n3561 VDD.n3162 1.23311
R9977 VDD.n5897 VDD.n4949 1.23311
R9978 VDD.n5887 VDD.n4954 1.23311
R9979 VDD.n5880 VDD.n4957 1.23311
R9980 VDD.n3554 VDD.n3167 1.23311
R9981 VDD.n3549 VDD.n3170 1.23311
R9982 VDD.n3737 VDD.n3736 1.23311
R9983 VDD.n6138 VDD.n4583 1.23311
R9984 VDD.n6145 VDD.n4580 1.23311
R9985 VDD.n3456 VDD.n3239 1.23311
R9986 VDD.n3461 VDD.n3236 1.23311
R9987 VDD.n5733 VDD.n5143 1.23311
R9988 VDD.n5740 VDD.n5140 1.23311
R9989 VDD.n3468 VDD.n3231 1.23311
R9990 VDD.n5750 VDD.n5135 1.23311
R9991 VDD.n3475 VDD.n3225 1.23311
R9992 VDD.n5760 VDD.n5129 1.23311
R9993 VDD.n3482 VDD.n3219 1.23311
R9994 VDD.n5770 VDD.n5123 1.23311
R9995 VDD.n3505 VDD.n3207 1.23311
R9996 VDD.n5806 VDD.n5101 1.23311
R9997 VDD.n3512 VDD.n3201 1.23311
R9998 VDD.n5816 VDD.n5095 1.23311
R9999 VDD.n3519 VDD.n3195 1.23311
R10000 VDD.n5826 VDD.n5089 1.23311
R10001 VDD.n3526 VDD.n3189 1.23311
R10002 VDD.n3531 VDD.n3186 1.23311
R10003 VDD.n5836 VDD.n5083 1.23311
R10004 VDD.n5843 VDD.n5080 1.23311
R10005 VDD.n5564 VDD.n5563 1.23311
R10006 VDD.n3355 VDD.n3320 1.23311
R10007 VDD.n3350 VDD.n3323 1.23311
R10008 VDD.n2669 VDD.n2544 1.23311
R10009 VDD.n2662 VDD.n2550 1.23311
R10010 VDD.n6589 VDD.n2850 1.23311
R10011 VDD.n2655 VDD.n2556 1.23311
R10012 VDD.n6579 VDD.n2856 1.23311
R10013 VDD.n6569 VDD.n2874 1.23311
R10014 VDD.n2648 VDD.n2568 1.23311
R10015 VDD.n2625 VDD.n2574 1.23311
R10016 VDD.n6533 VDD.n2884 1.23311
R10017 VDD.n2618 VDD.n2580 1.23311
R10018 VDD.n6523 VDD.n2890 1.23311
R10019 VDD.n2611 VDD.n2586 1.23311
R10020 VDD.n6513 VDD.n2896 1.23311
R10021 VDD.n6503 VDD.n2901 1.23311
R10022 VDD.n6496 VDD.n2904 1.23311
R10023 VDD.n2604 VDD.n2591 1.23311
R10024 VDD.n2599 VDD.n2594 1.23311
R10025 VDD.n2679 VDD.n2678 1.23311
R10026 VDD.n6599 VDD.n2844 1.23311
R10027 VDD.n6606 VDD.n2841 1.23311
R10028 VDD.n5582 VDD.t314 1.2215
R10029 VDD.n5654 VDD.t96 1.2215
R10030 VDD.n6053 VDD.t28 1.2215
R10031 VDD.n6125 VDD.t301 1.2215
R10032 VDD.n6200 VDD.t91 1.2215
R10033 VDD.n6272 VDD.t256 1.2215
R10034 VDD.n6355 VDD.t74 1.2215
R10035 VDD.n6427 VDD.t94 1.2215
R10036 VDD.n6514 VDD.t54 1.2215
R10037 VDD.n6586 VDD.t461 1.2215
R10038 VDD.n5751 VDD.t77 1.2215
R10039 VDD.n5823 VDD.t227 1.2215
R10040 VDD.n5898 VDD.t241 1.2215
R10041 VDD.n5970 VDD.t81 1.2215
R10042 VDD.n7007 VDD.n6888 1.21354
R10043 VDD.n7014 VDD.n6884 1.21354
R10044 VDD.n7066 VDD.n296 1.21354
R10045 VDD.n7073 VDD.n292 1.21354
R10046 VDD.t1134 VDD.t886 1.15992
R10047 VDD.t36 VDD.t1069 1.15992
R10048 VDD.t621 VDD.t36 1.15992
R10049 VDD.t189 VDD.t591 1.15992
R10050 VDD.n6629 VDD.n6628 1.15363
R10051 VDD.n6631 VDD.n6630 1.15363
R10052 VDD.n6632 VDD.n6631 1.15363
R10053 VDD.n6634 VDD.n6633 1.15363
R10054 VDD.n6635 VDD.n6634 1.15363
R10055 VDD.n6877 VDD.n6876 1.14664
R10056 VDD.n7116 VDD.n7077 1.13137
R10057 VDD.n7097 VDD.n7088 1.13137
R10058 VDD.n7551 VDD.n7548 1.13137
R10059 VDD.n7564 VDD.n7315 1.13137
R10060 VDD.n7573 VDD.n7304 1.13137
R10061 VDD.n7578 VDD.n7302 1.13137
R10062 VDD.n7109 VDD.n7108 1.13137
R10063 VDD.n632 VDD.n571 1.1255
R10064 VDD.n1033 VDD.n788 1.1255
R10065 VDD.n581 VDD.n572 1.1255
R10066 VDD.n1040 VDD.n784 1.1255
R10067 VDD.n576 VDD.n573 1.1255
R10068 VDD.n828 VDD.n794 1.1255
R10069 VDD.n823 VDD.n798 1.1255
R10070 VDD.n816 VDD.n801 1.1255
R10071 VDD.n1006 VDD.n980 1.1255
R10072 VDD.n809 VDD.n804 1.1255
R10073 VDD.n996 VDD.n989 1.1255
R10074 VDD.n6661 VDD.n6656 1.1255
R10075 VDD.n6839 VDD.n6832 1.1255
R10076 VDD.n6668 VDD.n6653 1.1255
R10077 VDD.n6849 VDD.n6823 1.1255
R10078 VDD.n6866 VDD.n6810 1.1255
R10079 VDD.n6675 VDD.n6650 1.1255
R10080 VDD.n6859 VDD.n6814 1.1255
R10081 VDD.n6680 VDD.n6649 1.1255
R10082 VDD.n627 VDD.n626 1.1255
R10083 VDD.n560 VDD.n556 1.1255
R10084 VDD.n567 VDD.n552 1.1255
R10085 VDD.n6997 VDD.n6996 1.12396
R10086 VDD.n968 VDD.n966 1.12396
R10087 VDD.n7234 VDD.n7225 1.12377
R10088 VDD.n283 VDD.n282 1.12377
R10089 VDD.n6998 VDD.n6997 1.12377
R10090 VDD.n773 VDD.n772 1.12377
R10091 VDD.n6840 VDD.t770 1.10231
R10092 VDD.n997 VDD.t285 1.10231
R10093 VDD.n194 VDD.n193 1.1018
R10094 VDD.n7236 VDD.n7235 1.1018
R10095 VDD.n3843 VDD.n3842 1.1016
R10096 VDD.n3638 VDD.n3637 1.1016
R10097 VDD.n397 VDD.n396 1.09615
R10098 VDD.n551 VDD.n548 1.09028
R10099 VDD.n783 VDD.n780 1.09028
R10100 VDD.n787 VDD.n786 1.09028
R10101 VDD.n792 VDD.n791 1.09028
R10102 VDD.n796 VDD.n795 1.09028
R10103 VDD.n6813 VDD.n6812 1.09028
R10104 VDD.n6809 VDD.n6808 1.09028
R10105 VDD.n555 VDD.n554 1.09028
R10106 VDD.n7697 VDD.n7301 1.07267
R10107 VDD.n7704 VDD.n7297 1.07267
R10108 VDD.n7257 VDD.n11 1.07267
R10109 VDD.n7247 VDD.n15 1.07267
R10110 VDD.n291 VDD.n288 1.06093
R10111 VDD.n6888 VDD.n6887 1.06093
R10112 VDD.n6883 VDD.n6880 1.06093
R10113 VDD.n6884 VDD.n6883 1.06093
R10114 VDD.n6887 VDD.n6886 1.06093
R10115 VDD.n295 VDD.n294 1.06093
R10116 VDD.n296 VDD.n295 1.06093
R10117 VDD.n292 VDD.n291 1.06093
R10118 VDD.n2401 VDD.t895 1.02677
R10119 VDD.n2419 VDD.t406 1.02677
R10120 VDD.n388 VDD.n387 1.02572
R10121 VDD.n7369 VDD.n7368 1.00811
R10122 VDD.n5432 VDD.n5431 0.992457
R10123 VDD.n3273 VDD.n3272 0.992457
R10124 VDD.n3270 VDD.n3269 0.992457
R10125 VDD.n3269 VDD.n3266 0.992457
R10126 VDD.n5371 VDD.n5368 0.992457
R10127 VDD.n3272 VDD.n3271 0.992457
R10128 VDD.n5374 VDD.n5373 0.992457
R10129 VDD.n5375 VDD.n5374 0.992457
R10130 VDD.n5372 VDD.n5371 0.992457
R10131 VDD.n2914 VDD.n2913 0.992457
R10132 VDD.n4130 VDD.n4129 0.992457
R10133 VDD.n2963 VDD.n2962 0.992457
R10134 VDD.n4132 VDD.n4131 0.992457
R10135 VDD.n4133 VDD.n4132 0.992457
R10136 VDD.n2961 VDD.n2960 0.992457
R10137 VDD.n2960 VDD.n2957 0.992457
R10138 VDD.n4129 VDD.n4128 0.992457
R10139 VDD.n2964 VDD.n2963 0.992457
R10140 VDD.n4390 VDD.n4389 0.992457
R10141 VDD.n2983 VDD.n2982 0.992457
R10142 VDD.n4392 VDD.n4391 0.992457
R10143 VDD.n4393 VDD.n4392 0.992457
R10144 VDD.n2981 VDD.n2980 0.992457
R10145 VDD.n2980 VDD.n2977 0.992457
R10146 VDD.n4389 VDD.n4388 0.992457
R10147 VDD.n2984 VDD.n2983 0.992457
R10148 VDD.n4450 VDD.n4449 0.992457
R10149 VDD.n3033 VDD.n3032 0.992457
R10150 VDD.n4452 VDD.n4451 0.992457
R10151 VDD.n4453 VDD.n4452 0.992457
R10152 VDD.n3031 VDD.n3030 0.992457
R10153 VDD.n3030 VDD.n3027 0.992457
R10154 VDD.n4449 VDD.n4448 0.992457
R10155 VDD.n3034 VDD.n3033 0.992457
R10156 VDD.n3941 VDD.n3940 0.992457
R10157 VDD.n3940 VDD.n3937 0.992457
R10158 VDD.n4069 VDD.n4066 0.992457
R10159 VDD.n2913 VDD.n2912 0.992457
R10160 VDD.n4072 VDD.n4071 0.992457
R10161 VDD.n4073 VDD.n4072 0.992457
R10162 VDD.n4070 VDD.n4069 0.992457
R10163 VDD.n3044 VDD.n3043 0.992457
R10164 VDD.n4640 VDD.n4639 0.992457
R10165 VDD.n3093 VDD.n3092 0.992457
R10166 VDD.n4642 VDD.n4641 0.992457
R10167 VDD.n4643 VDD.n4642 0.992457
R10168 VDD.n3091 VDD.n3090 0.992457
R10169 VDD.n3090 VDD.n3087 0.992457
R10170 VDD.n4639 VDD.n4638 0.992457
R10171 VDD.n3094 VDD.n3093 0.992457
R10172 VDD.n4894 VDD.n4893 0.992457
R10173 VDD.n3119 VDD.n3118 0.992457
R10174 VDD.n4896 VDD.n4895 0.992457
R10175 VDD.n4897 VDD.n4896 0.992457
R10176 VDD.n3117 VDD.n3116 0.992457
R10177 VDD.n3116 VDD.n3113 0.992457
R10178 VDD.n4893 VDD.n4892 0.992457
R10179 VDD.n3120 VDD.n3119 0.992457
R10180 VDD.n4954 VDD.n4953 0.992457
R10181 VDD.n3169 VDD.n3168 0.992457
R10182 VDD.n4956 VDD.n4955 0.992457
R10183 VDD.n4957 VDD.n4956 0.992457
R10184 VDD.n3167 VDD.n3166 0.992457
R10185 VDD.n3166 VDD.n3163 0.992457
R10186 VDD.n4953 VDD.n4952 0.992457
R10187 VDD.n3170 VDD.n3169 0.992457
R10188 VDD.n3736 VDD.n3735 0.992457
R10189 VDD.n3735 VDD.n3732 0.992457
R10190 VDD.n4579 VDD.n4576 0.992457
R10191 VDD.n3043 VDD.n3042 0.992457
R10192 VDD.n4582 VDD.n4581 0.992457
R10193 VDD.n4583 VDD.n4582 0.992457
R10194 VDD.n4580 VDD.n4579 0.992457
R10195 VDD.n3239 VDD.n3238 0.992457
R10196 VDD.n3236 VDD.n3235 0.992457
R10197 VDD.n3235 VDD.n3232 0.992457
R10198 VDD.n5139 VDD.n5136 0.992457
R10199 VDD.n3238 VDD.n3237 0.992457
R10200 VDD.n5142 VDD.n5141 0.992457
R10201 VDD.n5143 VDD.n5142 0.992457
R10202 VDD.n5140 VDD.n5139 0.992457
R10203 VDD.n3189 VDD.n3188 0.992457
R10204 VDD.n3186 VDD.n3185 0.992457
R10205 VDD.n3185 VDD.n3182 0.992457
R10206 VDD.n5079 VDD.n5076 0.992457
R10207 VDD.n3188 VDD.n3187 0.992457
R10208 VDD.n5082 VDD.n5081 0.992457
R10209 VDD.n5083 VDD.n5082 0.992457
R10210 VDD.n5080 VDD.n5079 0.992457
R10211 VDD.n3322 VDD.n3321 0.992457
R10212 VDD.n5562 VDD.n5561 0.992457
R10213 VDD.n5563 VDD.n5562 0.992457
R10214 VDD.n3320 VDD.n3319 0.992457
R10215 VDD.n3319 VDD.n3316 0.992457
R10216 VDD.n5431 VDD.n5430 0.992457
R10217 VDD.n3323 VDD.n3322 0.992457
R10218 VDD.n2544 VDD.n2543 0.992457
R10219 VDD.n2901 VDD.n2900 0.992457
R10220 VDD.n2593 VDD.n2592 0.992457
R10221 VDD.n2903 VDD.n2902 0.992457
R10222 VDD.n2904 VDD.n2903 0.992457
R10223 VDD.n2591 VDD.n2590 0.992457
R10224 VDD.n2590 VDD.n2587 0.992457
R10225 VDD.n2900 VDD.n2899 0.992457
R10226 VDD.n2594 VDD.n2593 0.992457
R10227 VDD.n2678 VDD.n2677 0.992457
R10228 VDD.n2677 VDD.n2674 0.992457
R10229 VDD.n2840 VDD.n2837 0.992457
R10230 VDD.n2543 VDD.n2542 0.992457
R10231 VDD.n2843 VDD.n2842 0.992457
R10232 VDD.n2844 VDD.n2843 0.992457
R10233 VDD.n2841 VDD.n2840 0.992457
R10234 VDD.n6878 VDD.n546 0.932563
R10235 VDD.n5545 VDD.n5544 0.878601
R10236 VDD.n3339 VDD.n3338 0.878601
R10237 VDD.n2693 VDD.n2692 0.878601
R10238 VDD.n1468 VDD.n1467 0.875507
R10239 VDD.n1250 VDD.n1249 0.875507
R10240 VDD.n2541 VDD.n2540 0.875507
R10241 VDD.n2056 VDD.n2055 0.875507
R10242 VDD.n541 VDD.n540 0.873539
R10243 VDD.n968 VDD.n967 0.873539
R10244 VDD.n3850 VDD.n3849 0.873539
R10245 VDD.n6317 VDD.n6316 0.873539
R10246 VDD.n3645 VDD.n3644 0.873539
R10247 VDD.n6014 VDD.n6013 0.873539
R10248 VDD.n5709 VDD.n5708 0.873539
R10249 VDD.n5713 VDD.n5712 0.873539
R10250 VDD.n3440 VDD.n3439 0.873539
R10251 VDD.n3444 VDD.n3443 0.873539
R10252 VDD.n1664 VDD.n1663 0.873539
R10253 VDD.n1536 VDD.n1535 0.873539
R10254 VDD.n2159 VDD.n2158 0.873539
R10255 VDD.n2350 VDD.n2349 0.873539
R10256 VDD.n7682 VDD.n7681 0.873539
R10257 VDD.n117 VDD.n116 0.873308
R10258 VDD.n7510 VDD.n7509 0.873308
R10259 VDD.n6801 VDD.n6786 0.873308
R10260 VDD.n6477 VDD.n6476 0.873308
R10261 VDD.n6162 VDD.n6161 0.873308
R10262 VDD.n6310 VDD.n6309 0.873308
R10263 VDD.n5861 VDD.n5860 0.873308
R10264 VDD.n6008 VDD.n6007 0.873308
R10265 VDD.n6624 VDD.n6623 0.873308
R10266 VDD.n6802 VDD.n6801 0.873308
R10267 VDD.n376 VDD.t885 0.870065
R10268 VDD.n401 VDD.n400 0.869196
R10269 VDD.n7377 VDD.n7376 0.851587
R10270 VDD.n7375 VDD.n7374 0.851587
R10271 VDD.n7373 VDD.n7359 0.851587
R10272 VDD.n7379 VDD.n7378 0.851587
R10273 VDD.n788 VDD.n787 0.847674
R10274 VDD.n784 VDD.n783 0.847674
R10275 VDD.n6810 VDD.n6809 0.847674
R10276 VDD.n6814 VDD.n6813 0.847674
R10277 VDD.n556 VDD.n555 0.847674
R10278 VDD.n552 VDD.n551 0.847674
R10279 VDD.n6637 VDD.n6636 0.8465
R10280 VDD.n7367 VDD.n7366 0.845717
R10281 VDD.n5598 VDD.t261 0.814501
R10282 VDD.n5638 VDD.t83 0.814501
R10283 VDD.n6069 VDD.t72 0.814501
R10284 VDD.n6109 VDD.t675 0.814501
R10285 VDD.n6216 VDD.t41 0.814501
R10286 VDD.n6256 VDD.t119 0.814501
R10287 VDD.n6371 VDD.t150 0.814501
R10288 VDD.n6411 VDD.t221 0.814501
R10289 VDD.n6530 VDD.t63 0.814501
R10290 VDD.n6570 VDD.t224 0.814501
R10291 VDD.n5767 VDD.t454 0.814501
R10292 VDD.n5807 VDD.t176 0.814501
R10293 VDD.n5914 VDD.t389 0.814501
R10294 VDD.n5954 VDD.t624 0.814501
R10295 VDD.n7299 VDD.n7298 0.700935
R10296 VDD.n7295 VDD.n7294 0.700935
R10297 VDD.n9 VDD.n8 0.700935
R10298 VDD.n13 VDD.n12 0.700935
R10299 VDD.n2348 VDD.n2347 0.684371
R10300 VDD.n2157 VDD.n2156 0.684371
R10301 VDD.n2054 VDD.n2053 0.684371
R10302 VDD.n7681 VDD.n7680 0.684371
R10303 VDD.n7681 VDD.n7679 0.684371
R10304 VDD.n7681 VDD.n7678 0.684371
R10305 VDD.n7681 VDD.n7677 0.684371
R10306 VDD.n7681 VDD.n7676 0.684371
R10307 VDD.n7681 VDD.n7675 0.684371
R10308 VDD.n7681 VDD.n7674 0.684371
R10309 VDD.n7681 VDD.n7673 0.684371
R10310 VDD.n7681 VDD.n7672 0.684371
R10311 VDD.n7681 VDD.n7671 0.684371
R10312 VDD.n7234 VDD.n7224 0.684371
R10313 VDD.n283 VDD.n281 0.684371
R10314 VDD.n283 VDD.n280 0.684371
R10315 VDD.n283 VDD.n279 0.684371
R10316 VDD.n283 VDD.n278 0.684371
R10317 VDD.n283 VDD.n277 0.684371
R10318 VDD.n283 VDD.n276 0.684371
R10319 VDD.n283 VDD.n275 0.684371
R10320 VDD.n284 VDD.n283 0.684371
R10321 VDD.n540 VDD.n539 0.684371
R10322 VDD.n540 VDD.n538 0.684371
R10323 VDD.n540 VDD.n537 0.684371
R10324 VDD.n540 VDD.n536 0.684371
R10325 VDD.n540 VDD.n535 0.684371
R10326 VDD.n969 VDD.n968 0.684371
R10327 VDD.n2911 VDD.n2909 0.684371
R10328 VDD.n2347 VDD.n2344 0.684371
R10329 VDD.n2156 VDD.n2153 0.684371
R10330 VDD.n2053 VDD.n2052 0.684371
R10331 VDD.n2053 VDD.n2051 0.684371
R10332 VDD.n2053 VDD.n2050 0.684371
R10333 VDD.n2053 VDD.n2049 0.684371
R10334 VDD.n2053 VDD.n2048 0.684371
R10335 VDD.n2053 VDD.n2047 0.684371
R10336 VDD.n2053 VDD.n2046 0.684371
R10337 VDD.n2053 VDD.n2045 0.684371
R10338 VDD.n2053 VDD.n2044 0.684371
R10339 VDD.n2053 VDD.n2043 0.684371
R10340 VDD.n2053 VDD.n2042 0.684371
R10341 VDD.n2053 VDD.n2041 0.684371
R10342 VDD.n116 VDD.n115 0.684132
R10343 VDD.n116 VDD.n114 0.684132
R10344 VDD.n116 VDD.n113 0.684132
R10345 VDD.n116 VDD.n112 0.684132
R10346 VDD.n116 VDD.n111 0.684132
R10347 VDD.n116 VDD.n110 0.684132
R10348 VDD.n116 VDD.n109 0.684132
R10349 VDD.n116 VDD.n108 0.684132
R10350 VDD.n116 VDD.n107 0.684132
R10351 VDD.n116 VDD.n106 0.684132
R10352 VDD.n7509 VDD.n7504 0.684132
R10353 VDD.n7509 VDD.n7505 0.684132
R10354 VDD.n7509 VDD.n7506 0.684132
R10355 VDD.n7509 VDD.n7507 0.684132
R10356 VDD.n7509 VDD.n7508 0.684132
R10357 VDD.n6801 VDD.n6787 0.684132
R10358 VDD.n6801 VDD.n6788 0.684132
R10359 VDD.n6801 VDD.n6789 0.684132
R10360 VDD.n6801 VDD.n6790 0.684132
R10361 VDD.n6801 VDD.n6791 0.684132
R10362 VDD.n6801 VDD.n6792 0.684132
R10363 VDD.n6801 VDD.n6793 0.684132
R10364 VDD.n6801 VDD.n6794 0.684132
R10365 VDD.n6801 VDD.n6795 0.684132
R10366 VDD.n6801 VDD.n6796 0.684132
R10367 VDD.n6801 VDD.n6797 0.684132
R10368 VDD.n6801 VDD.n6798 0.684132
R10369 VDD.n6801 VDD.n6799 0.684132
R10370 VDD.n6801 VDD.n6800 0.684132
R10371 VDD.n5706 VDD.n5705 0.684132
R10372 VDD.n5706 VDD.n5704 0.684132
R10373 VDD.n5706 VDD.n5703 0.684132
R10374 VDD.n5706 VDD.n5702 0.684132
R10375 VDD.n5706 VDD.n5701 0.684132
R10376 VDD.n5706 VDD.n5700 0.684132
R10377 VDD.n5706 VDD.n5699 0.684132
R10378 VDD.n5706 VDD.n5698 0.684132
R10379 VDD.n5706 VDD.n5697 0.684132
R10380 VDD.n5706 VDD.n5696 0.684132
R10381 VDD.n5706 VDD.n5695 0.684132
R10382 VDD.n5706 VDD.n5694 0.684132
R10383 VDD.n5706 VDD.n5693 0.684132
R10384 VDD.n5706 VDD.n5692 0.684132
R10385 VDD.n3041 VDD.n3039 0.684132
R10386 VDD.n6476 VDD.n6462 0.684132
R10387 VDD.n6476 VDD.n6475 0.684132
R10388 VDD.n6476 VDD.n6474 0.684132
R10389 VDD.n6476 VDD.n6473 0.684132
R10390 VDD.n6476 VDD.n6472 0.684132
R10391 VDD.n6476 VDD.n6471 0.684132
R10392 VDD.n6476 VDD.n6470 0.684132
R10393 VDD.n6476 VDD.n6469 0.684132
R10394 VDD.n6476 VDD.n6468 0.684132
R10395 VDD.n6476 VDD.n6467 0.684132
R10396 VDD.n6476 VDD.n6466 0.684132
R10397 VDD.n6476 VDD.n6465 0.684132
R10398 VDD.n6476 VDD.n6464 0.684132
R10399 VDD.n6476 VDD.n6463 0.684132
R10400 VDD.n6482 VDD.n6479 0.684132
R10401 VDD.n3177 VDD.n3175 0.684132
R10402 VDD.n5707 VDD.n5706 0.684132
R10403 VDD.n2538 VDD.n2526 0.684132
R10404 VDD.n2538 VDD.n2527 0.684132
R10405 VDD.n2538 VDD.n2528 0.684132
R10406 VDD.n2538 VDD.n2529 0.684132
R10407 VDD.n2538 VDD.n2530 0.684132
R10408 VDD.n2538 VDD.n2531 0.684132
R10409 VDD.n2538 VDD.n2532 0.684132
R10410 VDD.n2538 VDD.n2533 0.684132
R10411 VDD.n2538 VDD.n2534 0.684132
R10412 VDD.n2538 VDD.n2535 0.684132
R10413 VDD.n2538 VDD.n2536 0.684132
R10414 VDD.n2538 VDD.n2537 0.684132
R10415 VDD.n2539 VDD.n2538 0.684132
R10416 VDD.n1461 VDD.n1460 0.6755
R10417 VDD.n1458 VDD.n1457 0.6755
R10418 VDD.n1457 VDD.n1454 0.6755
R10419 VDD.n1135 VDD.n1132 0.6755
R10420 VDD.n1460 VDD.n1459 0.6755
R10421 VDD.n1138 VDD.n1137 0.6755
R10422 VDD.n1139 VDD.n1138 0.6755
R10423 VDD.n1136 VDD.n1135 0.6755
R10424 VDD.n1453 VDD.n1452 0.6755
R10425 VDD.n1450 VDD.n1449 0.6755
R10426 VDD.n1452 VDD.n1451 0.6755
R10427 VDD.n1361 VDD.n1360 0.6755
R10428 VDD.n1356 VDD.n1355 0.6755
R10429 VDD.n1355 VDD.n1352 0.6755
R10430 VDD.n1109 VDD.n1106 0.6755
R10431 VDD.n1360 VDD.n1359 0.6755
R10432 VDD.n1113 VDD.n1112 0.6755
R10433 VDD.n1115 VDD.n1113 0.6755
R10434 VDD.n1110 VDD.n1109 0.6755
R10435 VDD.n3297 VDD.n3296 0.673543
R10436 VDD.n5402 VDD.n5396 0.673543
R10437 VDD.n4110 VDD.n4109 0.673543
R10438 VDD.n2944 VDD.n2943 0.673543
R10439 VDD.n4420 VDD.n4419 0.673543
R10440 VDD.n3008 VDD.n3007 0.673543
R10441 VDD.n4620 VDD.n4619 0.673543
R10442 VDD.n3074 VDD.n3073 0.673543
R10443 VDD.n4924 VDD.n4923 0.673543
R10444 VDD.n3144 VDD.n3143 0.673543
R10445 VDD.n3219 VDD.n3218 0.673543
R10446 VDD.n5120 VDD.n5114 0.673543
R10447 VDD.n2871 VDD.n2870 0.673543
R10448 VDD.n2568 VDD.n2567 0.673543
R10449 VDD.n3296 VDD.n3292 0.626587
R10450 VDD.n5393 VDD.n5392 0.626587
R10451 VDD.n5402 VDD.n5401 0.626587
R10452 VDD.n4110 VDD.n4100 0.626587
R10453 VDD.n4106 VDD.n4105 0.626587
R10454 VDD.n2943 VDD.n2942 0.626587
R10455 VDD.n4420 VDD.n4410 0.626587
R10456 VDD.n4416 VDD.n4415 0.626587
R10457 VDD.n3007 VDD.n3006 0.626587
R10458 VDD.n4620 VDD.n4610 0.626587
R10459 VDD.n4616 VDD.n4615 0.626587
R10460 VDD.n3073 VDD.n3072 0.626587
R10461 VDD.n4924 VDD.n4914 0.626587
R10462 VDD.n4920 VDD.n4919 0.626587
R10463 VDD.n3143 VDD.n3142 0.626587
R10464 VDD.n3218 VDD.n3214 0.626587
R10465 VDD.n5111 VDD.n5110 0.626587
R10466 VDD.n5120 VDD.n5119 0.626587
R10467 VDD.n2871 VDD.n2861 0.626587
R10468 VDD.n2867 VDD.n2866 0.626587
R10469 VDD.n2567 VDD.n2566 0.626587
R10470 VDD.n2460 VDD.t184 0.616264
R10471 VDD.n2878 VDD.t264 0.607167
R10472 VDD.n2878 VDD.n2877 0.607167
R10473 VDD.n2876 VDD.t1125 0.607167
R10474 VDD.n2876 VDD.n2875 0.607167
R10475 VDD.n3311 VDD.t904 0.607167
R10476 VDD.n3311 VDD.n3310 0.607167
R10477 VDD.n3313 VDD.t253 0.607167
R10478 VDD.n3313 VDD.n3312 0.607167
R10479 VDD.n5423 VDD.t876 0.607167
R10480 VDD.n5423 VDD.n5422 0.607167
R10481 VDD.n5426 VDD.t260 0.607167
R10482 VDD.n5426 VDD.n5425 0.607167
R10483 VDD.n3305 VDD.t87 0.607167
R10484 VDD.n3305 VDD.n3304 0.607167
R10485 VDD.n3307 VDD.t182 0.607167
R10486 VDD.n3307 VDD.n3306 0.607167
R10487 VDD.n5417 VDD.t1025 0.607167
R10488 VDD.n5417 VDD.n5416 0.607167
R10489 VDD.n5420 VDD.t855 0.607167
R10490 VDD.n5420 VDD.n5419 0.607167
R10491 VDD.n3299 VDD.t925 0.607167
R10492 VDD.n3299 VDD.n3298 0.607167
R10493 VDD.n3301 VDD.t649 0.607167
R10494 VDD.n3301 VDD.n3300 0.607167
R10495 VDD.n5411 VDD.t262 0.607167
R10496 VDD.n5411 VDD.n5410 0.607167
R10497 VDD.n5414 VDD.t562 0.607167
R10498 VDD.n5414 VDD.n5413 0.607167
R10499 VDD.n5409 VDD.t710 0.607167
R10500 VDD.n5409 VDD.n5408 0.607167
R10501 VDD.n5407 VDD.t143 0.607167
R10502 VDD.n5407 VDD.n5406 0.607167
R10503 VDD.n5404 VDD.t912 0.607167
R10504 VDD.n5404 VDD.n5403 0.607167
R10505 VDD.n5395 VDD.t887 0.607167
R10506 VDD.n5395 VDD.n5394 0.607167
R10507 VDD.n3294 VDD.t781 0.607167
R10508 VDD.n3294 VDD.n3293 0.607167
R10509 VDD.n3287 VDD.t822 0.607167
R10510 VDD.n3287 VDD.n3286 0.607167
R10511 VDD.n3291 VDD.t436 0.607167
R10512 VDD.n3291 VDD.n3290 0.607167
R10513 VDD.n3289 VDD.t915 0.607167
R10514 VDD.n3289 VDD.n3288 0.607167
R10515 VDD.n5391 VDD.t456 0.607167
R10516 VDD.n5391 VDD.n5390 0.607167
R10517 VDD.n5389 VDD.t144 0.607167
R10518 VDD.n5389 VDD.n5388 0.607167
R10519 VDD.n5400 VDD.t543 0.607167
R10520 VDD.n5400 VDD.n5399 0.607167
R10521 VDD.n5398 VDD.t757 0.607167
R10522 VDD.n5398 VDD.n5397 0.607167
R10523 VDD.n3281 VDD.t634 0.607167
R10524 VDD.n3281 VDD.n3280 0.607167
R10525 VDD.n3283 VDD.t431 0.607167
R10526 VDD.n3283 VDD.n3282 0.607167
R10527 VDD.n5383 VDD.t930 0.607167
R10528 VDD.n5383 VDD.n5382 0.607167
R10529 VDD.n5386 VDD.t836 0.607167
R10530 VDD.n5386 VDD.n5385 0.607167
R10531 VDD.n3275 VDD.t475 0.607167
R10532 VDD.n3275 VDD.n3274 0.607167
R10533 VDD.n3277 VDD.t383 0.607167
R10534 VDD.n3277 VDD.n3276 0.607167
R10535 VDD.n5377 VDD.t715 0.607167
R10536 VDD.n5377 VDD.n5376 0.607167
R10537 VDD.n5380 VDD.t97 0.607167
R10538 VDD.n5380 VDD.n5379 0.607167
R10539 VDD.n4931 VDD.t552 0.607167
R10540 VDD.n4931 VDD.n4930 0.607167
R10541 VDD.n4929 VDD.t427 0.607167
R10542 VDD.n4929 VDD.n4928 0.607167
R10543 VDD.n4605 VDD.t1055 0.607167
R10544 VDD.n4605 VDD.n4604 0.607167
R10545 VDD.n4603 VDD.t1075 0.607167
R10546 VDD.n4603 VDD.n4602 0.607167
R10547 VDD.n4427 VDD.t911 0.607167
R10548 VDD.n4427 VDD.n4426 0.607167
R10549 VDD.n4425 VDD.t1116 0.607167
R10550 VDD.n4425 VDD.n4424 0.607167
R10551 VDD.n4095 VDD.t31 0.607167
R10552 VDD.n4095 VDD.n4094 0.607167
R10553 VDD.n4093 VDD.t785 0.607167
R10554 VDD.n4093 VDD.n4092 0.607167
R10555 VDD.n2916 VDD.t488 0.607167
R10556 VDD.n2916 VDD.n2915 0.607167
R10557 VDD.n2918 VDD.t951 0.607167
R10558 VDD.n2918 VDD.n2917 0.607167
R10559 VDD.n4075 VDD.t615 0.607167
R10560 VDD.n4075 VDD.n4074 0.607167
R10561 VDD.n4078 VDD.t95 0.607167
R10562 VDD.n4078 VDD.n4077 0.607167
R10563 VDD.n2922 VDD.t739 0.607167
R10564 VDD.n2922 VDD.n2921 0.607167
R10565 VDD.n2924 VDD.t22 0.607167
R10566 VDD.n2924 VDD.n2923 0.607167
R10567 VDD.n4081 VDD.t233 0.607167
R10568 VDD.n4081 VDD.n4080 0.607167
R10569 VDD.n4084 VDD.t997 0.607167
R10570 VDD.n4084 VDD.n4083 0.607167
R10571 VDD.n2928 VDD.t956 0.607167
R10572 VDD.n2928 VDD.n2927 0.607167
R10573 VDD.n2930 VDD.t714 0.607167
R10574 VDD.n2930 VDD.n2929 0.607167
R10575 VDD.n4087 VDD.t507 0.607167
R10576 VDD.n4087 VDD.n4086 0.607167
R10577 VDD.n4090 VDD.t359 0.607167
R10578 VDD.n4090 VDD.n4089 0.607167
R10579 VDD.n2934 VDD.t868 0.607167
R10580 VDD.n2934 VDD.n2933 0.607167
R10581 VDD.n2936 VDD.t544 0.607167
R10582 VDD.n2936 VDD.n2935 0.607167
R10583 VDD.n4108 VDD.t953 0.607167
R10584 VDD.n4108 VDD.n4107 0.607167
R10585 VDD.n4112 VDD.t151 0.607167
R10586 VDD.n4112 VDD.n4111 0.607167
R10587 VDD.n4097 VDD.t18 0.607167
R10588 VDD.n4097 VDD.n4096 0.607167
R10589 VDD.n4099 VDD.t525 0.607167
R10590 VDD.n4099 VDD.n4098 0.607167
R10591 VDD.n4102 VDD.t643 0.607167
R10592 VDD.n4102 VDD.n4101 0.607167
R10593 VDD.n4104 VDD.t172 0.607167
R10594 VDD.n4104 VDD.n4103 0.607167
R10595 VDD.n2939 VDD.t49 0.607167
R10596 VDD.n2939 VDD.n2938 0.607167
R10597 VDD.n2941 VDD.t426 0.607167
R10598 VDD.n2941 VDD.n2940 0.607167
R10599 VDD.n2946 VDD.t983 0.607167
R10600 VDD.n2946 VDD.n2945 0.607167
R10601 VDD.n2948 VDD.t977 0.607167
R10602 VDD.n2948 VDD.n2947 0.607167
R10603 VDD.n4115 VDD.t711 0.607167
R10604 VDD.n4115 VDD.n4114 0.607167
R10605 VDD.n4118 VDD.t126 0.607167
R10606 VDD.n4118 VDD.n4117 0.607167
R10607 VDD.n2952 VDD.t434 0.607167
R10608 VDD.n2952 VDD.n2951 0.607167
R10609 VDD.n2954 VDD.t689 0.607167
R10610 VDD.n2954 VDD.n2953 0.607167
R10611 VDD.n4121 VDD.t482 0.607167
R10612 VDD.n4121 VDD.n4120 0.607167
R10613 VDD.n4124 VDD.t561 0.607167
R10614 VDD.n4124 VDD.n4123 0.607167
R10615 VDD.n2986 VDD.t257 0.607167
R10616 VDD.n2986 VDD.n2985 0.607167
R10617 VDD.n2988 VDD.t635 0.607167
R10618 VDD.n2988 VDD.n2987 0.607167
R10619 VDD.n4395 VDD.t725 0.607167
R10620 VDD.n4395 VDD.n4394 0.607167
R10621 VDD.n4398 VDD.t884 0.607167
R10622 VDD.n4398 VDD.n4397 0.607167
R10623 VDD.n2992 VDD.t871 0.607167
R10624 VDD.n2992 VDD.n2991 0.607167
R10625 VDD.n2994 VDD.t650 0.607167
R10626 VDD.n2994 VDD.n2993 0.607167
R10627 VDD.n4401 VDD.t598 0.607167
R10628 VDD.n4401 VDD.n4400 0.607167
R10629 VDD.n4404 VDD.t890 0.607167
R10630 VDD.n4404 VDD.n4403 0.607167
R10631 VDD.n2998 VDD.t682 0.607167
R10632 VDD.n2998 VDD.n2997 0.607167
R10633 VDD.n3000 VDD.t164 0.607167
R10634 VDD.n3000 VDD.n2999 0.607167
R10635 VDD.n4418 VDD.t692 0.607167
R10636 VDD.n4418 VDD.n4417 0.607167
R10637 VDD.n4422 VDD.t604 0.607167
R10638 VDD.n4422 VDD.n4421 0.607167
R10639 VDD.n4409 VDD.t636 0.607167
R10640 VDD.n4409 VDD.n4408 0.607167
R10641 VDD.n4407 VDD.t797 0.607167
R10642 VDD.n4407 VDD.n4406 0.607167
R10643 VDD.n4414 VDD.t255 0.607167
R10644 VDD.n4414 VDD.n4413 0.607167
R10645 VDD.n4412 VDD.t203 0.607167
R10646 VDD.n4412 VDD.n4411 0.607167
R10647 VDD.n3005 VDD.t384 0.607167
R10648 VDD.n3005 VDD.n3004 0.607167
R10649 VDD.n3003 VDD.t756 0.607167
R10650 VDD.n3003 VDD.n3002 0.607167
R10651 VDD.n3010 VDD.t860 0.607167
R10652 VDD.n3010 VDD.n3009 0.607167
R10653 VDD.n3012 VDD.t42 0.607167
R10654 VDD.n3012 VDD.n3011 0.607167
R10655 VDD.n4429 VDD.t491 0.607167
R10656 VDD.n4429 VDD.n4428 0.607167
R10657 VDD.n4432 VDD.t554 0.607167
R10658 VDD.n4432 VDD.n4431 0.607167
R10659 VDD.n3016 VDD.t1412 0.607167
R10660 VDD.n3016 VDD.n3015 0.607167
R10661 VDD.n3018 VDD.t66 0.607167
R10662 VDD.n3018 VDD.n3017 0.607167
R10663 VDD.n4435 VDD.t460 0.607167
R10664 VDD.n4435 VDD.n4434 0.607167
R10665 VDD.n4438 VDD.t53 0.607167
R10666 VDD.n4438 VDD.n4437 0.607167
R10667 VDD.n3022 VDD.t894 0.607167
R10668 VDD.n3022 VDD.n3021 0.607167
R10669 VDD.n3024 VDD.t596 0.607167
R10670 VDD.n3024 VDD.n3023 0.607167
R10671 VDD.n4441 VDD.t215 0.607167
R10672 VDD.n4441 VDD.n4440 0.607167
R10673 VDD.n4444 VDD.t982 0.607167
R10674 VDD.n4444 VDD.n4443 0.607167
R10675 VDD.n3046 VDD.t441 0.607167
R10676 VDD.n3046 VDD.n3045 0.607167
R10677 VDD.n3048 VDD.t955 0.607167
R10678 VDD.n3048 VDD.n3047 0.607167
R10679 VDD.n4585 VDD.t698 0.607167
R10680 VDD.n4585 VDD.n4584 0.607167
R10681 VDD.n4588 VDD.t302 0.607167
R10682 VDD.n4588 VDD.n4587 0.607167
R10683 VDD.n3052 VDD.t674 0.607167
R10684 VDD.n3052 VDD.n3051 0.607167
R10685 VDD.n3054 VDD.t612 0.607167
R10686 VDD.n3054 VDD.n3053 0.607167
R10687 VDD.n4591 VDD.t118 0.607167
R10688 VDD.n4591 VDD.n4590 0.607167
R10689 VDD.n4594 VDD.t859 0.607167
R10690 VDD.n4594 VDD.n4593 0.607167
R10691 VDD.n3058 VDD.t659 0.607167
R10692 VDD.n3058 VDD.n3057 0.607167
R10693 VDD.n3060 VDD.t873 0.607167
R10694 VDD.n3060 VDD.n3059 0.607167
R10695 VDD.n4597 VDD.t588 0.607167
R10696 VDD.n4597 VDD.n4596 0.607167
R10697 VDD.n4600 VDD.t913 0.607167
R10698 VDD.n4600 VDD.n4599 0.607167
R10699 VDD.n3064 VDD.t1041 0.607167
R10700 VDD.n3064 VDD.n3063 0.607167
R10701 VDD.n3066 VDD.t73 0.607167
R10702 VDD.n3066 VDD.n3065 0.607167
R10703 VDD.n4618 VDD.t741 0.607167
R10704 VDD.n4618 VDD.n4617 0.607167
R10705 VDD.n4622 VDD.t815 0.607167
R10706 VDD.n4622 VDD.n4621 0.607167
R10707 VDD.n4607 VDD.t1010 0.607167
R10708 VDD.n4607 VDD.n4606 0.607167
R10709 VDD.n4609 VDD.t1409 0.607167
R10710 VDD.n4609 VDD.n4608 0.607167
R10711 VDD.n4612 VDD.t867 0.607167
R10712 VDD.n4612 VDD.n4611 0.607167
R10713 VDD.n4614 VDD.t527 0.607167
R10714 VDD.n4614 VDD.n4613 0.607167
R10715 VDD.n3069 VDD.t162 0.607167
R10716 VDD.n3069 VDD.n3068 0.607167
R10717 VDD.n3071 VDD.t758 0.607167
R10718 VDD.n3071 VDD.n3070 0.607167
R10719 VDD.n3076 VDD.t576 0.607167
R10720 VDD.n3076 VDD.n3075 0.607167
R10721 VDD.n3078 VDD.t568 0.607167
R10722 VDD.n3078 VDD.n3077 0.607167
R10723 VDD.n4625 VDD.t724 0.607167
R10724 VDD.n4625 VDD.n4624 0.607167
R10725 VDD.n4628 VDD.t893 0.607167
R10726 VDD.n4628 VDD.n4627 0.607167
R10727 VDD.n3082 VDD.t856 0.607167
R10728 VDD.n3082 VDD.n3081 0.607167
R10729 VDD.n3084 VDD.t637 0.607167
R10730 VDD.n3084 VDD.n3083 0.607167
R10731 VDD.n4631 VDD.t375 0.607167
R10732 VDD.n4631 VDD.n4630 0.607167
R10733 VDD.n4634 VDD.t564 0.607167
R10734 VDD.n4634 VDD.n4633 0.607167
R10735 VDD.n3122 VDD.t968 0.607167
R10736 VDD.n3122 VDD.n3121 0.607167
R10737 VDD.n3124 VDD.t872 0.607167
R10738 VDD.n3124 VDD.n3123 0.607167
R10739 VDD.n4899 VDD.t82 0.607167
R10740 VDD.n4899 VDD.n4898 0.607167
R10741 VDD.n4902 VDD.t719 0.607167
R10742 VDD.n4902 VDD.n4901 0.607167
R10743 VDD.n3128 VDD.t553 0.607167
R10744 VDD.n3128 VDD.n3127 0.607167
R10745 VDD.n3130 VDD.t464 0.607167
R10746 VDD.n3130 VDD.n3129 0.607167
R10747 VDD.n4905 VDD.t954 0.607167
R10748 VDD.n4905 VDD.n4904 0.607167
R10749 VDD.n4908 VDD.t71 0.607167
R10750 VDD.n4908 VDD.n4907 0.607167
R10751 VDD.n3134 VDD.t270 0.607167
R10752 VDD.n3134 VDD.n3133 0.607167
R10753 VDD.n3136 VDD.t718 0.607167
R10754 VDD.n3136 VDD.n3135 0.607167
R10755 VDD.n4922 VDD.t4 0.607167
R10756 VDD.n4922 VDD.n4921 0.607167
R10757 VDD.n4926 VDD.t854 0.607167
R10758 VDD.n4926 VDD.n4925 0.607167
R10759 VDD.n4913 VDD.t883 0.607167
R10760 VDD.n4913 VDD.n4912 0.607167
R10761 VDD.n4911 VDD.t335 0.607167
R10762 VDD.n4911 VDD.n4910 0.607167
R10763 VDD.n4918 VDD.t1090 0.607167
R10764 VDD.n4918 VDD.n4917 0.607167
R10765 VDD.n4916 VDD.t1405 0.607167
R10766 VDD.n4916 VDD.n4915 0.607167
R10767 VDD.n3141 VDD.t572 0.607167
R10768 VDD.n3141 VDD.n3140 0.607167
R10769 VDD.n3139 VDD.t141 0.607167
R10770 VDD.n3139 VDD.n3138 0.607167
R10771 VDD.n3146 VDD.t931 0.607167
R10772 VDD.n3146 VDD.n3145 0.607167
R10773 VDD.n3148 VDD.t601 0.607167
R10774 VDD.n3148 VDD.n3147 0.607167
R10775 VDD.n4933 VDD.t914 0.607167
R10776 VDD.n4933 VDD.n4932 0.607167
R10777 VDD.n4936 VDD.t390 0.607167
R10778 VDD.n4936 VDD.n4935 0.607167
R10779 VDD.n3152 VDD.t6 0.607167
R10780 VDD.n3152 VDD.n3151 0.607167
R10781 VDD.n3154 VDD.t303 0.607167
R10782 VDD.n3154 VDD.n3153 0.607167
R10783 VDD.n4939 VDD.t432 0.607167
R10784 VDD.n4939 VDD.n4938 0.607167
R10785 VDD.n4942 VDD.t65 0.607167
R10786 VDD.n4942 VDD.n4941 0.607167
R10787 VDD.n3158 VDD.t51 0.607167
R10788 VDD.n3158 VDD.n3157 0.607167
R10789 VDD.n3160 VDD.t644 0.607167
R10790 VDD.n3160 VDD.n3159 0.607167
R10791 VDD.n4945 VDD.t277 0.607167
R10792 VDD.n4945 VDD.n4944 0.607167
R10793 VDD.n4948 VDD.t1042 0.607167
R10794 VDD.n4948 VDD.n4947 0.607167
R10795 VDD.n3227 VDD.t487 0.607167
R10796 VDD.n3227 VDD.n3226 0.607167
R10797 VDD.n3229 VDD.t957 0.607167
R10798 VDD.n3229 VDD.n3228 0.607167
R10799 VDD.n5131 VDD.t565 0.607167
R10800 VDD.n5131 VDD.n5130 0.607167
R10801 VDD.n5134 VDD.t386 0.607167
R10802 VDD.n5134 VDD.n5133 0.607167
R10803 VDD.n3221 VDD.t642 0.607167
R10804 VDD.n3221 VDD.n3220 0.607167
R10805 VDD.n3223 VDD.t493 0.607167
R10806 VDD.n3223 VDD.n3222 0.607167
R10807 VDD.n5125 VDD.t864 0.607167
R10808 VDD.n5125 VDD.n5124 0.607167
R10809 VDD.n5128 VDD.t1123 0.607167
R10810 VDD.n5128 VDD.n5127 0.607167
R10811 VDD.n5122 VDD.t775 0.607167
R10812 VDD.n5122 VDD.n5121 0.607167
R10813 VDD.n5113 VDD.t1000 0.607167
R10814 VDD.n5113 VDD.n5112 0.607167
R10815 VDD.n3216 VDD.t1047 0.607167
R10816 VDD.n3216 VDD.n3215 0.607167
R10817 VDD.n3209 VDD.t455 0.607167
R10818 VDD.n3209 VDD.n3208 0.607167
R10819 VDD.n3211 VDD.t967 0.607167
R10820 VDD.n3211 VDD.n3210 0.607167
R10821 VDD.n3213 VDD.t1399 0.607167
R10822 VDD.n3213 VDD.n3212 0.607167
R10823 VDD.n5107 VDD.t20 0.607167
R10824 VDD.n5107 VDD.n5106 0.607167
R10825 VDD.n5109 VDD.t1400 0.607167
R10826 VDD.n5109 VDD.n5108 0.607167
R10827 VDD.n5116 VDD.t80 0.607167
R10828 VDD.n5116 VDD.n5115 0.607167
R10829 VDD.n5118 VDD.t196 0.607167
R10830 VDD.n5118 VDD.n5117 0.607167
R10831 VDD.n5105 VDD.t101 0.607167
R10832 VDD.n5105 VDD.n5104 0.607167
R10833 VDD.n5103 VDD.t425 0.607167
R10834 VDD.n5103 VDD.n5102 0.607167
R10835 VDD.n3203 VDD.t380 0.607167
R10836 VDD.n3203 VDD.n3202 0.607167
R10837 VDD.n3205 VDD.t474 0.607167
R10838 VDD.n3205 VDD.n3204 0.607167
R10839 VDD.n5097 VDD.t1124 0.607167
R10840 VDD.n5097 VDD.n5096 0.607167
R10841 VDD.n5100 VDD.t502 0.607167
R10842 VDD.n5100 VDD.n5099 0.607167
R10843 VDD.n3197 VDD.t962 0.607167
R10844 VDD.n3197 VDD.n3196 0.607167
R10845 VDD.n3199 VDD.t466 0.607167
R10846 VDD.n3199 VDD.n3198 0.607167
R10847 VDD.n5091 VDD.t651 0.607167
R10848 VDD.n5091 VDD.n5090 0.607167
R10849 VDD.n5094 VDD.t733 0.607167
R10850 VDD.n5094 VDD.n5093 0.607167
R10851 VDD.n3191 VDD.t501 0.607167
R10852 VDD.n3191 VDD.n3190 0.607167
R10853 VDD.n3193 VDD.t251 0.607167
R10854 VDD.n3193 VDD.n3192 0.607167
R10855 VDD.n5085 VDD.t736 0.607167
R10856 VDD.n5085 VDD.n5084 0.607167
R10857 VDD.n5088 VDD.t228 0.607167
R10858 VDD.n5088 VDD.n5087 0.607167
R10859 VDD.n2546 VDD.t463 0.607167
R10860 VDD.n2546 VDD.n2545 0.607167
R10861 VDD.n2548 VDD.t631 0.607167
R10862 VDD.n2548 VDD.n2547 0.607167
R10863 VDD.n2846 VDD.t1088 0.607167
R10864 VDD.n2846 VDD.n2845 0.607167
R10865 VDD.n2849 VDD.t462 0.607167
R10866 VDD.n2849 VDD.n2848 0.607167
R10867 VDD.n2552 VDD.t300 0.607167
R10868 VDD.n2552 VDD.n2551 0.607167
R10869 VDD.n2554 VDD.t1052 0.607167
R10870 VDD.n2554 VDD.n2553 0.607167
R10871 VDD.n2852 VDD.t149 0.607167
R10872 VDD.n2852 VDD.n2851 0.607167
R10873 VDD.n2855 VDD.t569 0.607167
R10874 VDD.n2855 VDD.n2854 0.607167
R10875 VDD.n2558 VDD.t505 0.607167
R10876 VDD.n2558 VDD.n2557 0.607167
R10877 VDD.n2560 VDD.t438 0.607167
R10878 VDD.n2560 VDD.n2559 0.607167
R10879 VDD.n2869 VDD.t566 0.607167
R10880 VDD.n2869 VDD.n2868 0.607167
R10881 VDD.n2873 VDD.t586 0.607167
R10882 VDD.n2873 VDD.n2872 0.607167
R10883 VDD.n2860 VDD.t371 0.607167
R10884 VDD.n2860 VDD.n2859 0.607167
R10885 VDD.n2858 VDD.t518 0.607167
R10886 VDD.n2858 VDD.n2857 0.607167
R10887 VDD.n2865 VDD.t607 0.607167
R10888 VDD.n2865 VDD.n2864 0.607167
R10889 VDD.n2863 VDD.t337 0.607167
R10890 VDD.n2863 VDD.n2862 0.607167
R10891 VDD.n2565 VDD.t1089 0.607167
R10892 VDD.n2565 VDD.n2564 0.607167
R10893 VDD.n2563 VDD.t524 0.607167
R10894 VDD.n2563 VDD.n2562 0.607167
R10895 VDD.n2570 VDD.t563 0.607167
R10896 VDD.n2570 VDD.n2569 0.607167
R10897 VDD.n2572 VDD.t64 0.607167
R10898 VDD.n2572 VDD.n2571 0.607167
R10899 VDD.n2880 VDD.t707 0.607167
R10900 VDD.n2880 VDD.n2879 0.607167
R10901 VDD.n2883 VDD.t863 0.607167
R10902 VDD.n2883 VDD.n2882 0.607167
R10903 VDD.n2576 VDD.t646 0.607167
R10904 VDD.n2576 VDD.n2575 0.607167
R10905 VDD.n2578 VDD.t1038 0.607167
R10906 VDD.n2578 VDD.n2577 0.607167
R10907 VDD.n2886 VDD.t1009 0.607167
R10908 VDD.n2886 VDD.n2885 0.607167
R10909 VDD.n2889 VDD.t952 0.607167
R10910 VDD.n2889 VDD.n2888 0.607167
R10911 VDD.n2582 VDD.t486 0.607167
R10912 VDD.n2582 VDD.n2581 0.607167
R10913 VDD.n2584 VDD.t506 0.607167
R10914 VDD.n2584 VDD.n2583 0.607167
R10915 VDD.n2892 VDD.t1020 0.607167
R10916 VDD.n2892 VDD.n2891 0.607167
R10917 VDD.n2895 VDD.t276 0.607167
R10918 VDD.n2895 VDD.n2894 0.607167
R10919 VDD.n1363 VDD.t1091 0.607167
R10920 VDD.n1363 VDD.n1362 0.607167
R10921 VDD.n1365 VDD.t365 0.607167
R10922 VDD.n1365 VDD.n1364 0.607167
R10923 VDD.n1367 VDD.t1078 0.607167
R10924 VDD.n1367 VDD.n1366 0.607167
R10925 VDD.n1369 VDD.t514 0.607167
R10926 VDD.n1369 VDD.n1368 0.607167
R10927 VDD.n1374 VDD.t208 0.607167
R10928 VDD.n1374 VDD.n1373 0.607167
R10929 VDD.n1376 VDD.t1085 0.607167
R10930 VDD.n1376 VDD.n1375 0.607167
R10931 VDD.n1378 VDD.t1106 0.607167
R10932 VDD.n1378 VDD.n1377 0.607167
R10933 VDD.n1380 VDD.t334 0.607167
R10934 VDD.n1380 VDD.n1379 0.607167
R10935 VDD.n1385 VDD.t185 0.607167
R10936 VDD.n1385 VDD.n1384 0.607167
R10937 VDD.n1387 VDD.t363 0.607167
R10938 VDD.n1387 VDD.n1386 0.607167
R10939 VDD.n1389 VDD.t920 0.607167
R10940 VDD.n1389 VDD.n1388 0.607167
R10941 VDD.n1391 VDD.t946 0.607167
R10942 VDD.n1391 VDD.n1390 0.607167
R10943 VDD.n1396 VDD.t170 0.607167
R10944 VDD.n1396 VDD.n1395 0.607167
R10945 VDD.n1398 VDD.t360 0.607167
R10946 VDD.n1398 VDD.n1397 0.607167
R10947 VDD.n1400 VDD.t110 0.607167
R10948 VDD.n1400 VDD.n1399 0.607167
R10949 VDD.n1402 VDD.t534 0.607167
R10950 VDD.n1402 VDD.n1401 0.607167
R10951 VDD.n1407 VDD.t943 0.607167
R10952 VDD.n1407 VDD.n1406 0.607167
R10953 VDD.n1409 VDD.t307 0.607167
R10954 VDD.n1409 VDD.n1408 0.607167
R10955 VDD.n1411 VDD.t308 0.607167
R10956 VDD.n1411 VDD.n1410 0.607167
R10957 VDD.n1413 VDD.t807 0.607167
R10958 VDD.n1413 VDD.n1412 0.607167
R10959 VDD.n1418 VDD.t794 0.607167
R10960 VDD.n1418 VDD.n1417 0.607167
R10961 VDD.n1420 VDD.t532 0.607167
R10962 VDD.n1420 VDD.n1419 0.607167
R10963 VDD.n1422 VDD.t533 0.607167
R10964 VDD.n1422 VDD.n1421 0.607167
R10965 VDD.n1424 VDD.t539 0.607167
R10966 VDD.n1424 VDD.n1423 0.607167
R10967 VDD.n1126 VDD.t897 0.607167
R10968 VDD.n1126 VDD.n1125 0.607167
R10969 VDD.n1123 VDD.t896 0.607167
R10970 VDD.n1123 VDD.n1122 0.607167
R10971 VDD.n1437 VDD.t1017 0.607167
R10972 VDD.n1437 VDD.n1436 0.607167
R10973 VDD.n1435 VDD.t1016 0.607167
R10974 VDD.n1435 VDD.n1434 0.607167
R10975 VDD.n1120 VDD.t593 0.607167
R10976 VDD.n1120 VDD.n1119 0.607167
R10977 VDD.n1117 VDD.t1132 0.607167
R10978 VDD.n1117 VDD.n1116 0.607167
R10979 VDD.n1431 VDD.t831 0.607167
R10980 VDD.n1431 VDD.n1430 0.607167
R10981 VDD.n1429 VDD.t575 0.607167
R10982 VDD.n1429 VDD.n1428 0.607167
R10983 VDD.n1114 VDD.t213 0.607167
R10984 VDD.n1358 VDD.t131 0.607167
R10985 VDD.n1111 VDD.t132 0.607167
R10986 VDD.n1357 VDD.t362 0.607167
R10987 VDD.n446 VDD.n389 0.597239
R10988 VDD.n441 VDD.n404 0.597239
R10989 VDD.n7415 VDD.n7380 0.597239
R10990 VDD.n7410 VDD.n7409 0.597239
R10991 VDD.n7107 VDD.n7106 0.58197
R10992 VDD.n7087 VDD.t1137 0.58197
R10993 VDD.n7087 VDD.n7086 0.58197
R10994 VDD.n7084 VDD.t346 0.58197
R10995 VDD.n7084 VDD.n7083 0.58197
R10996 VDD.n7081 VDD.t395 0.58197
R10997 VDD.n7081 VDD.n7080 0.58197
R10998 VDD.n7079 VDD.t330 0.58197
R10999 VDD.n7079 VDD.n7078 0.58197
R11000 VDD.n7547 VDD.t1102 0.58197
R11001 VDD.n7547 VDD.n7546 0.58197
R11002 VDD.n7544 VDD.t521 0.58197
R11003 VDD.n7544 VDD.n7543 0.58197
R11004 VDD.n7541 VDD.t1098 0.58197
R11005 VDD.n7541 VDD.n7540 0.58197
R11006 VDD.n7539 VDD.t1074 0.58197
R11007 VDD.n7539 VDD.n7538 0.58197
R11008 VDD.n7314 VDD.t523 0.58197
R11009 VDD.n7314 VDD.n7313 0.58197
R11010 VDD.n7311 VDD.t1103 0.58197
R11011 VDD.n7311 VDD.n7310 0.58197
R11012 VDD.n7308 VDD.t1073 0.58197
R11013 VDD.n7308 VDD.n7307 0.58197
R11014 VDD.n7306 VDD.t655 0.58197
R11015 VDD.n7306 VDD.n7305 0.58197
R11016 VDD.n7303 VDD.t115 0.58197
R11017 VDD.n7289 VDD.t326 0.58197
R11018 VDD.n7289 VDD.t1204 0.58197
R11019 VDD.n7290 VDD.t656 0.58197
R11020 VDD.n7290 VDD.t1390 0.58197
R11021 VDD.n7291 VDD.t972 0.58197
R11022 VDD.n7291 VDD.t1175 0.58197
R11023 VDD.n800 VDD.t1140 0.58197
R11024 VDD.n800 VDD.n799 0.58197
R11025 VDD.n973 VDD.t760 0.58197
R11026 VDD.n973 VDD.n972 0.58197
R11027 VDD.n976 VDD.t969 0.58197
R11028 VDD.n976 VDD.n975 0.58197
R11029 VDD.n979 VDD.t782 0.58197
R11030 VDD.n979 VDD.n978 0.58197
R11031 VDD.n803 VDD.t538 0.58197
R11032 VDD.n803 VDD.n802 0.58197
R11033 VDD.n982 VDD.t940 0.58197
R11034 VDD.n982 VDD.n981 0.58197
R11035 VDD.n985 VDD.t133 0.58197
R11036 VDD.n985 VDD.n984 0.58197
R11037 VDD.n988 VDD.t106 0.58197
R11038 VDD.n988 VDD.n987 0.58197
R11039 VDD.n6655 VDD.t1133 0.58197
R11040 VDD.n6655 VDD.n6654 0.58197
R11041 VDD.n6825 VDD.t771 0.58197
R11042 VDD.n6825 VDD.n6824 0.58197
R11043 VDD.n6828 VDD.t1406 0.58197
R11044 VDD.n6828 VDD.n6827 0.58197
R11045 VDD.n6831 VDD.t802 0.58197
R11046 VDD.n6831 VDD.n6830 0.58197
R11047 VDD.n6652 VDD.t291 0.58197
R11048 VDD.n6652 VDD.n6651 0.58197
R11049 VDD.n6816 VDD.t404 0.58197
R11050 VDD.n6816 VDD.n6815 0.58197
R11051 VDD.n6819 VDD.t937 0.58197
R11052 VDD.n6819 VDD.n6818 0.58197
R11053 VDD.n6822 VDD.t994 0.58197
R11054 VDD.n6822 VDD.n6821 0.58197
R11055 VDD.n5 VDD.t1315 0.58197
R11056 VDD.n5 VDD.n4 0.58197
R11057 VDD.n3 VDD.t1164 0.58197
R11058 VDD.n3 VDD.n2 0.58197
R11059 VDD.n1 VDD.t1231 0.58197
R11060 VDD.n1 VDD.n0 0.58197
R11061 VDD.n1800 VDD.n1799 0.520296
R11062 VDD.n1803 VDD.n1802 0.520296
R11063 VDD.n3041 VDD.n3035 0.480464
R11064 VDD.n2911 VDD.n2905 0.480464
R11065 VDD.n3177 VDD.n3171 0.480464
R11066 VDD.n395 VDD.t789 0.4555
R11067 VDD.n395 VDD.n394 0.4555
R11068 VDD.n393 VDD.t784 0.4555
R11069 VDD.n393 VDD.n392 0.4555
R11070 VDD.n391 VDD.n390 0.4555
R11071 VDD.n7365 VDD.t352 0.4555
R11072 VDD.n7365 VDD.n7364 0.4555
R11073 VDD.n7363 VDD.t1070 0.4555
R11074 VDD.n7363 VDD.n7362 0.4555
R11075 VDD.n7361 VDD.t325 0.4555
R11076 VDD.n7361 VDD.n7360 0.4555
R11077 VDD.n7319 VDD.t696 0.4555
R11078 VDD.n7319 VDD.n7318 0.4555
R11079 VDD.n7321 VDD.t622 0.4555
R11080 VDD.n7321 VDD.n7320 0.4555
R11081 VDD.n340 VDD.t791 0.4555
R11082 VDD.n340 VDD.n339 0.4555
R11083 VDD.n338 VDD.t1398 0.4555
R11084 VDD.n338 VDD.n337 0.4555
R11085 VDD.n336 VDD.t971 0.4555
R11086 VDD.n336 VDD.n335 0.4555
R11087 VDD.n301 VDD.t1303 0.4555
R11088 VDD.n298 VDD.t1160 0.4555
R11089 VDD.n298 VDD.n297 0.4555
R11090 VDD.n3436 VDD.n3255 0.444312
R11091 VDD.n3445 VDD.n3240 0.444312
R11092 VDD.n3851 VDD.n2966 0.444312
R11093 VDD.n3646 VDD.n3096 0.444312
R11094 VDD.n3096 VDD.n3095 0.42125
R11095 VDD.n2966 VDD.n2965 0.411125
R11096 VDD.n6630 VDD.n6629 0.411125
R11097 VDD.n6633 VDD.n6632 0.411125
R11098 VDD.n3850 VDD.n3846 0.401
R11099 VDD.n3645 VDD.n3641 0.401
R11100 VDD.n3444 VDD.n3440 0.401
R11101 VDD.n6319 VDD.n6314 0.395938
R11102 VDD.n1799 VDD.n1798 0.386214
R11103 VDD.n1802 VDD.n1801 0.386214
R11104 VDD.n6017 VDD.n6012 0.385812
R11105 VDD.n5715 VDD.n5710 0.375687
R11106 VDD.n6874 VDD.n6647 0.354031
R11107 VDD.n321 VDD.n303 0.344848
R11108 VDD.n325 VDD.n300 0.344848
R11109 VDD.n314 VDD.n304 0.344848
R11110 VDD.n7533 VDD.n7358 0.340935
R11111 VDD.n7529 VDD.n7375 0.340935
R11112 VDD.n7522 VDD.n7379 0.340935
R11113 VDD.n7354 VDD.n7317 0.340935
R11114 VDD.n7322 VDD.t621 0.290355
R11115 VDD.n2321 VDD.n1800 0.279684
R11116 VDD.n2182 VDD.n1803 0.279684
R11117 VDD.n7273 VDD.t111 0.271356
R11118 VDD.n400 VDD.n399 0.266587
R11119 VDD.n7373 VDD.n7370 0.266587
R11120 VDD.n6636 VDD.n6635 0.257
R11121 VDD.n1646 VDD.n1462 0.239276
R11122 VDD.n1553 VDD.n1552 0.239276
R11123 VDD.n6875 VDD.n1104 0.222688
R11124 VDD.n6874 VDD.n6873 0.222688
R11125 VDD.n6639 VDD.n6638 0.219875
R11126 VDD.n7024 VDD.n6878 0.203563
R11127 VDD.n6647 VDD.n2541 0.195969
R11128 VDD.n1481 VDD.n1464 0.195194
R11129 VDD.n1520 VDD.n1463 0.195194
R11130 VDD.n2133 VDD.n1936 0.195194
R11131 VDD.n2075 VDD.n1937 0.195194
R11132 VDD.n7294 VDD.n7293 0.190283
R11133 VDD.n8 VDD.n7 0.190283
R11134 VDD.n6883 VDD.n6882 0.157022
R11135 VDD.n291 VDD.n290 0.157022
R11136 VDD.n399 VDD.n398 0.157022
R11137 VDD.n398 VDD.n397 0.157022
R11138 VDD.n7370 VDD.n7369 0.157022
R11139 VDD.n7373 VDD.n7372 0.157022
R11140 VDD.n7317 VDD.n7316 0.157022
R11141 VDD.n303 VDD.n302 0.157022
R11142 VDD.n300 VDD.n299 0.157022
R11143 VDD.n783 VDD.n782 0.157022
R11144 VDD.n791 VDD.n790 0.157022
R11145 VDD.n6809 VDD.n6806 0.157022
R11146 VDD.n551 VDD.n550 0.157022
R11147 VDD.n3269 VDD.n3268 0.157022
R11148 VDD.n5371 VDD.n5370 0.157022
R11149 VDD.n4129 VDD.n4127 0.157022
R11150 VDD.n2960 VDD.n2959 0.157022
R11151 VDD.n4389 VDD.n4387 0.157022
R11152 VDD.n2980 VDD.n2979 0.157022
R11153 VDD.n4449 VDD.n4447 0.157022
R11154 VDD.n3030 VDD.n3029 0.157022
R11155 VDD.n3940 VDD.n3939 0.157022
R11156 VDD.n4069 VDD.n4068 0.157022
R11157 VDD.n4639 VDD.n4637 0.157022
R11158 VDD.n3090 VDD.n3089 0.157022
R11159 VDD.n4893 VDD.n4891 0.157022
R11160 VDD.n3116 VDD.n3115 0.157022
R11161 VDD.n4953 VDD.n4951 0.157022
R11162 VDD.n3166 VDD.n3165 0.157022
R11163 VDD.n3735 VDD.n3734 0.157022
R11164 VDD.n4579 VDD.n4578 0.157022
R11165 VDD.n3235 VDD.n3234 0.157022
R11166 VDD.n5139 VDD.n5138 0.157022
R11167 VDD.n3185 VDD.n3184 0.157022
R11168 VDD.n5079 VDD.n5078 0.157022
R11169 VDD.n5431 VDD.n5429 0.157022
R11170 VDD.n3319 VDD.n3318 0.157022
R11171 VDD.n2900 VDD.n2898 0.157022
R11172 VDD.n2590 VDD.n2589 0.157022
R11173 VDD.n2677 VDD.n2676 0.157022
R11174 VDD.n2840 VDD.n2839 0.157022
R11175 VDD.n1457 VDD.n1456 0.157022
R11176 VDD.n1135 VDD.n1134 0.157022
R11177 VDD.n1449 VDD.n1448 0.157022
R11178 VDD.n1355 VDD.n1354 0.157022
R11179 VDD.n1109 VDD.n1108 0.157022
R11180 VDD.n6878 VDD.n6877 0.149958
R11181 VDD.n6640 VDD.n6639 0.141125
R11182 VDD.n6641 VDD.n6640 0.141125
R11183 VDD.n6642 VDD.n6641 0.141125
R11184 VDD.n6643 VDD.n6642 0.141125
R11185 VDD.n6644 VDD.n6643 0.141125
R11186 VDD.n6645 VDD.n6644 0.141125
R11187 VDD.n6646 VDD.n6645 0.141125
R11188 VDD.n6647 VDD.n6646 0.141125
R11189 VDD.n6876 VDD.n778 0.122562
R11190 VDD.n5720 VDD.n5144 0.122281
R11191 VDD.n5710 VDD.n5272 0.122281
R11192 VDD.n6635 VDD.n6627 0.122281
R11193 VDD.n6876 VDD.n6875 0.104958
R11194 VDD.n199 VDD.n197 0.0760357
R11195 VDD.n201 VDD.n199 0.0760357
R11196 VDD.n203 VDD.n201 0.0760357
R11197 VDD.n205 VDD.n203 0.0760357
R11198 VDD.n207 VDD.n205 0.0760357
R11199 VDD.n209 VDD.n207 0.0760357
R11200 VDD.n211 VDD.n209 0.0760357
R11201 VDD.n213 VDD.n211 0.0760357
R11202 VDD.n215 VDD.n213 0.0760357
R11203 VDD.n217 VDD.n215 0.0760357
R11204 VDD.n219 VDD.n217 0.0760357
R11205 VDD.n221 VDD.n219 0.0760357
R11206 VDD.n223 VDD.n221 0.0760357
R11207 VDD.n225 VDD.n223 0.0760357
R11208 VDD.n227 VDD.n225 0.0760357
R11209 VDD.n229 VDD.n227 0.0760357
R11210 VDD.n232 VDD.n229 0.0760357
R11211 VDD.n234 VDD.n232 0.0760357
R11212 VDD.n237 VDD.n234 0.0760357
R11213 VDD.n239 VDD.n237 0.0760357
R11214 VDD.n242 VDD.n239 0.0760357
R11215 VDD.n244 VDD.n242 0.0760357
R11216 VDD.n247 VDD.n244 0.0760357
R11217 VDD.n249 VDD.n247 0.0760357
R11218 VDD.n252 VDD.n249 0.0760357
R11219 VDD.n254 VDD.n252 0.0760357
R11220 VDD.n257 VDD.n254 0.0760357
R11221 VDD.n259 VDD.n257 0.0760357
R11222 VDD.n262 VDD.n259 0.0760357
R11223 VDD.n264 VDD.n262 0.0760357
R11224 VDD.n267 VDD.n264 0.0760357
R11225 VDD.n269 VDD.n267 0.0760357
R11226 VDD.n272 VDD.n269 0.0760357
R11227 VDD.n274 VDD.n272 0.0760357
R11228 VDD.n286 VDD.n274 0.0760357
R11229 VDD.n7670 VDD.n7668 0.0760357
R11230 VDD.n7668 VDD.n7665 0.0760357
R11231 VDD.n7665 VDD.n7663 0.0760357
R11232 VDD.n7663 VDD.n7660 0.0760357
R11233 VDD.n7660 VDD.n7658 0.0760357
R11234 VDD.n7658 VDD.n7655 0.0760357
R11235 VDD.n7655 VDD.n7653 0.0760357
R11236 VDD.n7653 VDD.n7650 0.0760357
R11237 VDD.n7650 VDD.n7648 0.0760357
R11238 VDD.n7648 VDD.n7645 0.0760357
R11239 VDD.n7645 VDD.n7643 0.0760357
R11240 VDD.n7643 VDD.n7640 0.0760357
R11241 VDD.n7640 VDD.n7638 0.0760357
R11242 VDD.n7638 VDD.n7635 0.0760357
R11243 VDD.n7635 VDD.n7633 0.0760357
R11244 VDD.n7633 VDD.n7630 0.0760357
R11245 VDD.n7630 VDD.n7628 0.0760357
R11246 VDD.n7628 VDD.n7626 0.0760357
R11247 VDD.n7626 VDD.n7624 0.0760357
R11248 VDD.n7624 VDD.n7622 0.0760357
R11249 VDD.n7622 VDD.n7620 0.0760357
R11250 VDD.n7620 VDD.n7618 0.0760357
R11251 VDD.n7618 VDD.n7616 0.0760357
R11252 VDD.n7616 VDD.n7614 0.0760357
R11253 VDD.n7614 VDD.n7612 0.0760357
R11254 VDD.n7612 VDD.n7610 0.0760357
R11255 VDD.n7610 VDD.n7608 0.0760357
R11256 VDD.n7608 VDD.n7606 0.0760357
R11257 VDD.n7606 VDD.n7604 0.0760357
R11258 VDD.n7604 VDD.n7602 0.0760357
R11259 VDD.n7602 VDD.n7600 0.0760357
R11260 VDD.n7600 VDD.n7598 0.0760357
R11261 VDD.n7598 VDD.n7596 0.0760357
R11262 VDD.n7596 VDD.n7594 0.0760357
R11263 VDD.n7594 VDD.n7592 0.0760357
R11264 VDD.n7592 VDD.n7590 0.0760357
R11265 VDD.n7223 VDD.n7220 0.0760357
R11266 VDD.n7220 VDD.n7217 0.0760357
R11267 VDD.n7217 VDD.n7214 0.0760357
R11268 VDD.n7214 VDD.n7211 0.0760357
R11269 VDD.n7211 VDD.n7208 0.0760357
R11270 VDD.n7208 VDD.n7205 0.0760357
R11271 VDD.n7205 VDD.n7202 0.0760357
R11272 VDD.n7202 VDD.n7199 0.0760357
R11273 VDD.n7199 VDD.n7196 0.0760357
R11274 VDD.n7196 VDD.n7193 0.0760357
R11275 VDD.n7193 VDD.n7190 0.0760357
R11276 VDD.n7190 VDD.n7187 0.0760357
R11277 VDD.n7187 VDD.n7184 0.0760357
R11278 VDD.n7184 VDD.n7181 0.0760357
R11279 VDD.n7181 VDD.n7178 0.0760357
R11280 VDD.n7178 VDD.n7175 0.0760357
R11281 VDD.n7175 VDD.n7172 0.0760357
R11282 VDD.n7172 VDD.n7169 0.0760357
R11283 VDD.n7169 VDD.n7166 0.0760357
R11284 VDD.n7166 VDD.n7163 0.0760357
R11285 VDD.n7163 VDD.n7160 0.0760357
R11286 VDD.n7160 VDD.n7157 0.0760357
R11287 VDD.n7157 VDD.n7154 0.0760357
R11288 VDD.n7154 VDD.n7151 0.0760357
R11289 VDD.n7151 VDD.n7148 0.0760357
R11290 VDD.n7148 VDD.n7146 0.0760357
R11291 VDD.n7146 VDD.n7144 0.0760357
R11292 VDD.n7144 VDD.n7142 0.0760357
R11293 VDD.n7142 VDD.n7140 0.0760357
R11294 VDD.n7140 VDD.n7138 0.0760357
R11295 VDD.n7138 VDD.n7136 0.0760357
R11296 VDD.n7136 VDD.n7134 0.0760357
R11297 VDD.n7134 VDD.n7132 0.0760357
R11298 VDD.n7132 VDD.n7130 0.0760357
R11299 VDD.n7130 VDD.n7128 0.0760357
R11300 VDD.n7128 VDD.n7126 0.0760357
R11301 VDD.n105 VDD.n103 0.0760357
R11302 VDD.n103 VDD.n101 0.0760357
R11303 VDD.n101 VDD.n98 0.0760357
R11304 VDD.n98 VDD.n96 0.0760357
R11305 VDD.n96 VDD.n93 0.0760357
R11306 VDD.n93 VDD.n91 0.0760357
R11307 VDD.n91 VDD.n88 0.0760357
R11308 VDD.n88 VDD.n86 0.0760357
R11309 VDD.n86 VDD.n83 0.0760357
R11310 VDD.n83 VDD.n81 0.0760357
R11311 VDD.n81 VDD.n78 0.0760357
R11312 VDD.n78 VDD.n76 0.0760357
R11313 VDD.n76 VDD.n73 0.0760357
R11314 VDD.n73 VDD.n71 0.0760357
R11315 VDD.n71 VDD.n68 0.0760357
R11316 VDD.n68 VDD.n66 0.0760357
R11317 VDD.n66 VDD.n64 0.0760357
R11318 VDD.n64 VDD.n62 0.0760357
R11319 VDD.n62 VDD.n60 0.0760357
R11320 VDD.n60 VDD.n58 0.0760357
R11321 VDD.n58 VDD.n56 0.0760357
R11322 VDD.n56 VDD.n54 0.0760357
R11323 VDD.n54 VDD.n52 0.0760357
R11324 VDD.n52 VDD.n50 0.0760357
R11325 VDD.n50 VDD.n48 0.0760357
R11326 VDD.n48 VDD.n46 0.0760357
R11327 VDD.n46 VDD.n44 0.0760357
R11328 VDD.n44 VDD.n42 0.0760357
R11329 VDD.n42 VDD.n40 0.0760357
R11330 VDD.n40 VDD.n38 0.0760357
R11331 VDD.n38 VDD.n36 0.0760357
R11332 VDD.n36 VDD.n34 0.0760357
R11333 VDD.n34 VDD.n32 0.0760357
R11334 VDD.n32 VDD.n30 0.0760357
R11335 VDD.n30 VDD.n28 0.0760357
R11336 VDD.n28 VDD.n26 0.0760357
R11337 VDD.n6892 VDD.n6890 0.0760357
R11338 VDD.n6894 VDD.n6892 0.0760357
R11339 VDD.n6896 VDD.n6894 0.0760357
R11340 VDD.n6898 VDD.n6896 0.0760357
R11341 VDD.n6900 VDD.n6898 0.0760357
R11342 VDD.n6902 VDD.n6900 0.0760357
R11343 VDD.n6904 VDD.n6902 0.0760357
R11344 VDD.n6906 VDD.n6904 0.0760357
R11345 VDD.n6908 VDD.n6906 0.0760357
R11346 VDD.n6911 VDD.n6908 0.0760357
R11347 VDD.n6914 VDD.n6911 0.0760357
R11348 VDD.n6917 VDD.n6914 0.0760357
R11349 VDD.n6920 VDD.n6917 0.0760357
R11350 VDD.n6923 VDD.n6920 0.0760357
R11351 VDD.n6926 VDD.n6923 0.0760357
R11352 VDD.n6929 VDD.n6926 0.0760357
R11353 VDD.n6932 VDD.n6929 0.0760357
R11354 VDD.n6935 VDD.n6932 0.0760357
R11355 VDD.n6938 VDD.n6935 0.0760357
R11356 VDD.n6941 VDD.n6938 0.0760357
R11357 VDD.n6944 VDD.n6941 0.0760357
R11358 VDD.n6947 VDD.n6944 0.0760357
R11359 VDD.n6950 VDD.n6947 0.0760357
R11360 VDD.n6953 VDD.n6950 0.0760357
R11361 VDD.n6956 VDD.n6953 0.0760357
R11362 VDD.n6959 VDD.n6956 0.0760357
R11363 VDD.n6962 VDD.n6959 0.0760357
R11364 VDD.n6965 VDD.n6962 0.0760357
R11365 VDD.n6968 VDD.n6965 0.0760357
R11366 VDD.n6971 VDD.n6968 0.0760357
R11367 VDD.n6974 VDD.n6971 0.0760357
R11368 VDD.n6977 VDD.n6974 0.0760357
R11369 VDD.n6980 VDD.n6977 0.0760357
R11370 VDD.n6983 VDD.n6980 0.0760357
R11371 VDD.n6986 VDD.n6983 0.0760357
R11372 VDD.n7000 VDD.n6986 0.0760357
R11373 VDD.n640 VDD.n638 0.0760357
R11374 VDD.n642 VDD.n640 0.0760357
R11375 VDD.n644 VDD.n642 0.0760357
R11376 VDD.n646 VDD.n644 0.0760357
R11377 VDD.n648 VDD.n646 0.0760357
R11378 VDD.n650 VDD.n648 0.0760357
R11379 VDD.n652 VDD.n650 0.0760357
R11380 VDD.n654 VDD.n652 0.0760357
R11381 VDD.n656 VDD.n654 0.0760357
R11382 VDD.n658 VDD.n656 0.0760357
R11383 VDD.n660 VDD.n658 0.0760357
R11384 VDD.n662 VDD.n660 0.0760357
R11385 VDD.n664 VDD.n662 0.0760357
R11386 VDD.n666 VDD.n664 0.0760357
R11387 VDD.n668 VDD.n666 0.0760357
R11388 VDD.n670 VDD.n668 0.0760357
R11389 VDD.n672 VDD.n670 0.0760357
R11390 VDD.n674 VDD.n672 0.0760357
R11391 VDD.n677 VDD.n674 0.0760357
R11392 VDD.n680 VDD.n677 0.0760357
R11393 VDD.n683 VDD.n680 0.0760357
R11394 VDD.n686 VDD.n683 0.0760357
R11395 VDD.n689 VDD.n686 0.0760357
R11396 VDD.n692 VDD.n689 0.0760357
R11397 VDD.n695 VDD.n692 0.0760357
R11398 VDD.n698 VDD.n695 0.0760357
R11399 VDD.n701 VDD.n698 0.0760357
R11400 VDD.n704 VDD.n701 0.0760357
R11401 VDD.n707 VDD.n704 0.0760357
R11402 VDD.n710 VDD.n707 0.0760357
R11403 VDD.n713 VDD.n710 0.0760357
R11404 VDD.n716 VDD.n713 0.0760357
R11405 VDD.n719 VDD.n716 0.0760357
R11406 VDD.n722 VDD.n719 0.0760357
R11407 VDD.n725 VDD.n722 0.0760357
R11408 VDD.n728 VDD.n725 0.0760357
R11409 VDD.n731 VDD.n728 0.0760357
R11410 VDD.n734 VDD.n731 0.0760357
R11411 VDD.n737 VDD.n734 0.0760357
R11412 VDD.n740 VDD.n737 0.0760357
R11413 VDD.n743 VDD.n740 0.0760357
R11414 VDD.n746 VDD.n743 0.0760357
R11415 VDD.n749 VDD.n746 0.0760357
R11416 VDD.n752 VDD.n749 0.0760357
R11417 VDD.n775 VDD.n752 0.0760357
R11418 VDD.n838 VDD.n836 0.0760357
R11419 VDD.n840 VDD.n838 0.0760357
R11420 VDD.n842 VDD.n840 0.0760357
R11421 VDD.n844 VDD.n842 0.0760357
R11422 VDD.n846 VDD.n844 0.0760357
R11423 VDD.n848 VDD.n846 0.0760357
R11424 VDD.n850 VDD.n848 0.0760357
R11425 VDD.n852 VDD.n850 0.0760357
R11426 VDD.n854 VDD.n852 0.0760357
R11427 VDD.n856 VDD.n854 0.0760357
R11428 VDD.n858 VDD.n856 0.0760357
R11429 VDD.n860 VDD.n858 0.0760357
R11430 VDD.n862 VDD.n860 0.0760357
R11431 VDD.n864 VDD.n862 0.0760357
R11432 VDD.n866 VDD.n864 0.0760357
R11433 VDD.n868 VDD.n866 0.0760357
R11434 VDD.n870 VDD.n868 0.0760357
R11435 VDD.n872 VDD.n870 0.0760357
R11436 VDD.n874 VDD.n872 0.0760357
R11437 VDD.n877 VDD.n874 0.0760357
R11438 VDD.n880 VDD.n877 0.0760357
R11439 VDD.n883 VDD.n880 0.0760357
R11440 VDD.n886 VDD.n883 0.0760357
R11441 VDD.n889 VDD.n886 0.0760357
R11442 VDD.n892 VDD.n889 0.0760357
R11443 VDD.n895 VDD.n892 0.0760357
R11444 VDD.n898 VDD.n895 0.0760357
R11445 VDD.n901 VDD.n898 0.0760357
R11446 VDD.n904 VDD.n901 0.0760357
R11447 VDD.n907 VDD.n904 0.0760357
R11448 VDD.n910 VDD.n907 0.0760357
R11449 VDD.n913 VDD.n910 0.0760357
R11450 VDD.n916 VDD.n913 0.0760357
R11451 VDD.n919 VDD.n916 0.0760357
R11452 VDD.n922 VDD.n919 0.0760357
R11453 VDD.n925 VDD.n922 0.0760357
R11454 VDD.n928 VDD.n925 0.0760357
R11455 VDD.n931 VDD.n928 0.0760357
R11456 VDD.n934 VDD.n931 0.0760357
R11457 VDD.n937 VDD.n934 0.0760357
R11458 VDD.n940 VDD.n937 0.0760357
R11459 VDD.n943 VDD.n940 0.0760357
R11460 VDD.n946 VDD.n943 0.0760357
R11461 VDD.n948 VDD.n946 0.0760357
R11462 VDD.n971 VDD.n948 0.0760357
R11463 VDD.n6689 VDD.n6687 0.0760357
R11464 VDD.n6691 VDD.n6689 0.0760357
R11465 VDD.n6693 VDD.n6691 0.0760357
R11466 VDD.n6695 VDD.n6693 0.0760357
R11467 VDD.n6697 VDD.n6695 0.0760357
R11468 VDD.n6699 VDD.n6697 0.0760357
R11469 VDD.n6701 VDD.n6699 0.0760357
R11470 VDD.n6703 VDD.n6701 0.0760357
R11471 VDD.n6705 VDD.n6703 0.0760357
R11472 VDD.n6707 VDD.n6705 0.0760357
R11473 VDD.n6709 VDD.n6707 0.0760357
R11474 VDD.n6711 VDD.n6709 0.0760357
R11475 VDD.n6713 VDD.n6711 0.0760357
R11476 VDD.n6715 VDD.n6713 0.0760357
R11477 VDD.n6717 VDD.n6715 0.0760357
R11478 VDD.n6719 VDD.n6717 0.0760357
R11479 VDD.n6721 VDD.n6719 0.0760357
R11480 VDD.n6723 VDD.n6721 0.0760357
R11481 VDD.n6725 VDD.n6723 0.0760357
R11482 VDD.n6727 VDD.n6725 0.0760357
R11483 VDD.n6729 VDD.n6727 0.0760357
R11484 VDD.n6731 VDD.n6729 0.0760357
R11485 VDD.n6733 VDD.n6731 0.0760357
R11486 VDD.n6735 VDD.n6733 0.0760357
R11487 VDD.n6737 VDD.n6735 0.0760357
R11488 VDD.n6739 VDD.n6737 0.0760357
R11489 VDD.n6741 VDD.n6739 0.0760357
R11490 VDD.n6743 VDD.n6741 0.0760357
R11491 VDD.n6745 VDD.n6743 0.0760357
R11492 VDD.n6748 VDD.n6745 0.0760357
R11493 VDD.n6750 VDD.n6748 0.0760357
R11494 VDD.n6753 VDD.n6750 0.0760357
R11495 VDD.n6755 VDD.n6753 0.0760357
R11496 VDD.n6758 VDD.n6755 0.0760357
R11497 VDD.n6760 VDD.n6758 0.0760357
R11498 VDD.n6763 VDD.n6760 0.0760357
R11499 VDD.n6765 VDD.n6763 0.0760357
R11500 VDD.n6768 VDD.n6765 0.0760357
R11501 VDD.n6770 VDD.n6768 0.0760357
R11502 VDD.n6773 VDD.n6770 0.0760357
R11503 VDD.n6775 VDD.n6773 0.0760357
R11504 VDD.n6778 VDD.n6775 0.0760357
R11505 VDD.n6780 VDD.n6778 0.0760357
R11506 VDD.n6783 VDD.n6780 0.0745948
R11507 VDD.n6785 VDD.n6783 0.073431
R11508 VDD.n122 VDD.n119 0.053375
R11509 VDD.n129 VDD.n126 0.053375
R11510 VDD.n136 VDD.n133 0.053375
R11511 VDD.n139 VDD.n136 0.053375
R11512 VDD.n142 VDD.n139 0.053375
R11513 VDD.n145 VDD.n142 0.053375
R11514 VDD.n148 VDD.n145 0.053375
R11515 VDD.n151 VDD.n148 0.053375
R11516 VDD.n154 VDD.n151 0.053375
R11517 VDD.n157 VDD.n154 0.053375
R11518 VDD.n160 VDD.n157 0.053375
R11519 VDD.n163 VDD.n160 0.053375
R11520 VDD.n166 VDD.n163 0.053375
R11521 VDD.n169 VDD.n166 0.053375
R11522 VDD.n172 VDD.n169 0.053375
R11523 VDD.n175 VDD.n172 0.053375
R11524 VDD.n178 VDD.n175 0.053375
R11525 VDD.n188 VDD.n185 0.053375
R11526 VDD.n195 VDD.n192 0.053375
R11527 VDD.n534 VDD.n532 0.053375
R11528 VDD.n532 VDD.n529 0.053375
R11529 VDD.n529 VDD.n527 0.053375
R11530 VDD.n527 VDD.n524 0.053375
R11531 VDD.n524 VDD.n522 0.053375
R11532 VDD.n522 VDD.n519 0.053375
R11533 VDD.n519 VDD.n517 0.053375
R11534 VDD.n517 VDD.n514 0.053375
R11535 VDD.n514 VDD.n512 0.053375
R11536 VDD.n512 VDD.n509 0.053375
R11537 VDD.n509 VDD.n507 0.053375
R11538 VDD.n507 VDD.n504 0.053375
R11539 VDD.n504 VDD.n502 0.053375
R11540 VDD.n502 VDD.n499 0.053375
R11541 VDD.n499 VDD.n497 0.053375
R11542 VDD.n497 VDD.n494 0.053375
R11543 VDD.n494 VDD.n492 0.053375
R11544 VDD.n492 VDD.n489 0.053375
R11545 VDD.n489 VDD.n487 0.053375
R11546 VDD.n487 VDD.n484 0.053375
R11547 VDD.n484 VDD.n482 0.053375
R11548 VDD.n482 VDD.n479 0.053375
R11549 VDD.n479 VDD.n477 0.053375
R11550 VDD.n477 VDD.n475 0.053375
R11551 VDD.n475 VDD.n473 0.053375
R11552 VDD.n473 VDD.n471 0.053375
R11553 VDD.n471 VDD.n469 0.053375
R11554 VDD.n469 VDD.n467 0.053375
R11555 VDD.n467 VDD.n465 0.053375
R11556 VDD.n465 VDD.n463 0.053375
R11557 VDD.n463 VDD.n461 0.053375
R11558 VDD.n461 VDD.n459 0.053375
R11559 VDD.n459 VDD.n457 0.053375
R11560 VDD.n7503 VDD.n7501 0.053375
R11561 VDD.n7501 VDD.n7498 0.053375
R11562 VDD.n7498 VDD.n7496 0.053375
R11563 VDD.n7496 VDD.n7493 0.053375
R11564 VDD.n7493 VDD.n7491 0.053375
R11565 VDD.n7491 VDD.n7488 0.053375
R11566 VDD.n7488 VDD.n7486 0.053375
R11567 VDD.n7486 VDD.n7483 0.053375
R11568 VDD.n7483 VDD.n7481 0.053375
R11569 VDD.n7481 VDD.n7478 0.053375
R11570 VDD.n7478 VDD.n7476 0.053375
R11571 VDD.n7476 VDD.n7473 0.053375
R11572 VDD.n7473 VDD.n7471 0.053375
R11573 VDD.n7471 VDD.n7468 0.053375
R11574 VDD.n7468 VDD.n7466 0.053375
R11575 VDD.n7466 VDD.n7463 0.053375
R11576 VDD.n7463 VDD.n7461 0.053375
R11577 VDD.n7461 VDD.n7458 0.053375
R11578 VDD.n7458 VDD.n7456 0.053375
R11579 VDD.n7456 VDD.n7453 0.053375
R11580 VDD.n7453 VDD.n7451 0.053375
R11581 VDD.n7451 VDD.n7448 0.053375
R11582 VDD.n7448 VDD.n7446 0.053375
R11583 VDD.n7446 VDD.n7444 0.053375
R11584 VDD.n7444 VDD.n7442 0.053375
R11585 VDD.n7442 VDD.n7440 0.053375
R11586 VDD.n7440 VDD.n7438 0.053375
R11587 VDD.n7438 VDD.n7436 0.053375
R11588 VDD.n7436 VDD.n7434 0.053375
R11589 VDD.n7434 VDD.n7432 0.053375
R11590 VDD.n7432 VDD.n7430 0.053375
R11591 VDD.n7430 VDD.n7428 0.053375
R11592 VDD.n7428 VDD.n7426 0.053375
R11593 VDD.n454 VDD.n452 0.053375
R11594 VDD.n452 VDD.n450 0.053375
R11595 VDD.n450 VDD.n448 0.053375
R11596 VDD.n445 VDD.n443 0.053375
R11597 VDD.n440 VDD.n438 0.053375
R11598 VDD.n438 VDD.n436 0.053375
R11599 VDD.n436 VDD.n434 0.053375
R11600 VDD.n434 VDD.n432 0.053375
R11601 VDD.n432 VDD.n430 0.053375
R11602 VDD.n430 VDD.n428 0.053375
R11603 VDD.n428 VDD.n426 0.053375
R11604 VDD.n426 VDD.n424 0.053375
R11605 VDD.n424 VDD.n422 0.053375
R11606 VDD.n422 VDD.n420 0.053375
R11607 VDD.n420 VDD.n418 0.053375
R11608 VDD.n418 VDD.n416 0.053375
R11609 VDD.n416 VDD.n414 0.053375
R11610 VDD.n414 VDD.n412 0.053375
R11611 VDD.n412 VDD.n410 0.053375
R11612 VDD.n410 VDD.n408 0.053375
R11613 VDD.n408 VDD.n406 0.053375
R11614 VDD.n7384 VDD.n7382 0.053375
R11615 VDD.n7386 VDD.n7384 0.053375
R11616 VDD.n7388 VDD.n7386 0.053375
R11617 VDD.n7390 VDD.n7388 0.053375
R11618 VDD.n7392 VDD.n7390 0.053375
R11619 VDD.n7394 VDD.n7392 0.053375
R11620 VDD.n7396 VDD.n7394 0.053375
R11621 VDD.n7398 VDD.n7396 0.053375
R11622 VDD.n7400 VDD.n7398 0.053375
R11623 VDD.n7402 VDD.n7400 0.053375
R11624 VDD.n7404 VDD.n7402 0.053375
R11625 VDD.n7406 VDD.n7404 0.053375
R11626 VDD.n7408 VDD.n7406 0.053375
R11627 VDD.n7414 VDD.n7412 0.053375
R11628 VDD.n7419 VDD.n7417 0.053375
R11629 VDD.n7421 VDD.n7419 0.053375
R11630 VDD.n7423 VDD.n7421 0.053375
R11631 VDD.n546 VDD.n545 0.053375
R11632 VDD.n310 VDD.n307 0.053375
R11633 VDD.n313 VDD.n310 0.053375
R11634 VDD.n320 VDD.n317 0.053375
R11635 VDD.n331 VDD.n328 0.053375
R11636 VDD.n334 VDD.n331 0.053375
R11637 VDD.n385 VDD.n382 0.053375
R11638 VDD.n378 VDD.n375 0.053375
R11639 VDD.n375 VDD.n372 0.053375
R11640 VDD.n372 VDD.n369 0.053375
R11641 VDD.n365 VDD.n362 0.053375
R11642 VDD.n362 VDD.n359 0.053375
R11643 VDD.n359 VDD.n356 0.053375
R11644 VDD.n356 VDD.n353 0.053375
R11645 VDD.n349 VDD.n346 0.053375
R11646 VDD.n346 VDD.n343 0.053375
R11647 VDD.n7327 VDD.n7324 0.053375
R11648 VDD.n7334 VDD.n7331 0.053375
R11649 VDD.n7337 VDD.n7334 0.053375
R11650 VDD.n7340 VDD.n7337 0.053375
R11651 VDD.n7347 VDD.n7344 0.053375
R11652 VDD.n7350 VDD.n7347 0.053375
R11653 VDD.n7353 VDD.n7350 0.053375
R11654 VDD.n7528 VDD.n7525 0.053375
R11655 VDD.n7521 VDD.n7518 0.053375
R11656 VDD.n7518 VDD.n7515 0.053375
R11657 VDD.n7515 VDD.n7512 0.053375
R11658 VDD.n6685 VDD.n6684 0.053375
R11659 VDD.n6684 VDD.n6682 0.053375
R11660 VDD.n6679 VDD.n6677 0.053375
R11661 VDD.n6674 VDD.n6672 0.053375
R11662 VDD.n6672 VDD.n6670 0.053375
R11663 VDD.n6667 VDD.n6665 0.053375
R11664 VDD.n6665 VDD.n6663 0.053375
R11665 VDD.n6660 VDD.n6658 0.053375
R11666 VDD.n808 VDD.n806 0.053375
R11667 VDD.n813 VDD.n811 0.053375
R11668 VDD.n815 VDD.n813 0.053375
R11669 VDD.n820 VDD.n818 0.053375
R11670 VDD.n822 VDD.n820 0.053375
R11671 VDD.n827 VDD.n825 0.053375
R11672 VDD.n832 VDD.n830 0.053375
R11673 VDD.n834 VDD.n832 0.053375
R11674 VDD.n580 VDD.n578 0.053375
R11675 VDD.n585 VDD.n583 0.053375
R11676 VDD.n587 VDD.n585 0.053375
R11677 VDD.n589 VDD.n587 0.053375
R11678 VDD.n591 VDD.n589 0.053375
R11679 VDD.n593 VDD.n591 0.053375
R11680 VDD.n595 VDD.n593 0.053375
R11681 VDD.n597 VDD.n595 0.053375
R11682 VDD.n599 VDD.n597 0.053375
R11683 VDD.n601 VDD.n599 0.053375
R11684 VDD.n603 VDD.n601 0.053375
R11685 VDD.n605 VDD.n603 0.053375
R11686 VDD.n607 VDD.n605 0.053375
R11687 VDD.n609 VDD.n607 0.053375
R11688 VDD.n611 VDD.n609 0.053375
R11689 VDD.n613 VDD.n611 0.053375
R11690 VDD.n615 VDD.n613 0.053375
R11691 VDD.n617 VDD.n615 0.053375
R11692 VDD.n619 VDD.n617 0.053375
R11693 VDD.n621 VDD.n619 0.053375
R11694 VDD.n623 VDD.n621 0.053375
R11695 VDD.n625 VDD.n623 0.053375
R11696 VDD.n631 VDD.n629 0.053375
R11697 VDD.n636 VDD.n634 0.053375
R11698 VDD.n6872 VDD.n6869 0.053375
R11699 VDD.n6865 VDD.n6862 0.053375
R11700 VDD.n6858 VDD.n6855 0.053375
R11701 VDD.n6855 VDD.n6852 0.053375
R11702 VDD.n6848 VDD.n6845 0.053375
R11703 VDD.n6845 VDD.n6842 0.053375
R11704 VDD.n6838 VDD.n6835 0.053375
R11705 VDD.n995 VDD.n992 0.053375
R11706 VDD.n1002 VDD.n999 0.053375
R11707 VDD.n1005 VDD.n1002 0.053375
R11708 VDD.n1012 VDD.n1009 0.053375
R11709 VDD.n1015 VDD.n1012 0.053375
R11710 VDD.n1018 VDD.n1015 0.053375
R11711 VDD.n1021 VDD.n1018 0.053375
R11712 VDD.n1024 VDD.n1021 0.053375
R11713 VDD.n1027 VDD.n1024 0.053375
R11714 VDD.n1029 VDD.n1027 0.053375
R11715 VDD.n1032 VDD.n1029 0.053375
R11716 VDD.n1039 VDD.n1036 0.053375
R11717 VDD.n1046 VDD.n1043 0.053375
R11718 VDD.n1049 VDD.n1046 0.053375
R11719 VDD.n1052 VDD.n1049 0.053375
R11720 VDD.n1055 VDD.n1052 0.053375
R11721 VDD.n1058 VDD.n1055 0.053375
R11722 VDD.n1061 VDD.n1058 0.053375
R11723 VDD.n1064 VDD.n1061 0.053375
R11724 VDD.n1067 VDD.n1064 0.053375
R11725 VDD.n1070 VDD.n1067 0.053375
R11726 VDD.n1073 VDD.n1070 0.053375
R11727 VDD.n1076 VDD.n1073 0.053375
R11728 VDD.n1079 VDD.n1076 0.053375
R11729 VDD.n1082 VDD.n1079 0.053375
R11730 VDD.n1085 VDD.n1082 0.053375
R11731 VDD.n1088 VDD.n1085 0.053375
R11732 VDD.n1091 VDD.n1088 0.053375
R11733 VDD.n1094 VDD.n1091 0.053375
R11734 VDD.n1097 VDD.n1094 0.053375
R11735 VDD.n1100 VDD.n1097 0.053375
R11736 VDD.n1103 VDD.n1100 0.053375
R11737 VDD.n566 VDD.n563 0.053375
R11738 VDD.n7013 VDD.n7010 0.053375
R11739 VDD.n7020 VDD.n7017 0.053375
R11740 VDD.n7023 VDD.n7020 0.053375
R11741 VDD.n7030 VDD.n7027 0.053375
R11742 VDD.n7033 VDD.n7030 0.053375
R11743 VDD.n7036 VDD.n7033 0.053375
R11744 VDD.n7039 VDD.n7036 0.053375
R11745 VDD.n7043 VDD.n7039 0.053375
R11746 VDD.n7046 VDD.n7043 0.053375
R11747 VDD.n7049 VDD.n7046 0.053375
R11748 VDD.n7052 VDD.n7049 0.053375
R11749 VDD.n7055 VDD.n7052 0.053375
R11750 VDD.n7058 VDD.n7055 0.053375
R11751 VDD.n7065 VDD.n7062 0.053375
R11752 VDD.n7072 VDD.n7069 0.053375
R11753 VDD.n7124 VDD.n7076 0.053375
R11754 VDD.n7124 VDD.n7122 0.053375
R11755 VDD.n7122 VDD.n7120 0.053375
R11756 VDD.n7120 VDD.n7118 0.053375
R11757 VDD.n7115 VDD.n7113 0.053375
R11758 VDD.n7113 VDD.n7111 0.053375
R11759 VDD.n7105 VDD.n7103 0.053375
R11760 VDD.n7103 VDD.n7101 0.053375
R11761 VDD.n7101 VDD.n7099 0.053375
R11762 VDD.n7096 VDD.n7094 0.053375
R11763 VDD.n7094 VDD.n7092 0.053375
R11764 VDD.n7092 VDD.n7090 0.053375
R11765 VDD.n7556 VDD.n7553 0.053375
R11766 VDD.n7558 VDD.n7556 0.053375
R11767 VDD.n7563 VDD.n7561 0.053375
R11768 VDD.n7568 VDD.n7566 0.053375
R11769 VDD.n7570 VDD.n7568 0.053375
R11770 VDD.n7572 VDD.n7570 0.053375
R11771 VDD.n7577 VDD.n7575 0.053375
R11772 VDD.n7582 VDD.n7580 0.053375
R11773 VDD.n7584 VDD.n7582 0.053375
R11774 VDD.n7586 VDD.n7584 0.053375
R11775 VDD.n7588 VDD.n7586 0.053375
R11776 VDD.n7240 VDD.n7237 0.053375
R11777 VDD.n7243 VDD.n7240 0.053375
R11778 VDD.n7246 VDD.n7243 0.053375
R11779 VDD.n7253 VDD.n7250 0.053375
R11780 VDD.n7256 VDD.n7253 0.053375
R11781 VDD.n7263 VDD.n7260 0.053375
R11782 VDD.n7266 VDD.n7263 0.053375
R11783 VDD.n7269 VDD.n7266 0.053375
R11784 VDD.n7272 VDD.n7269 0.053375
R11785 VDD.n7275 VDD.n7272 0.053375
R11786 VDD.n7278 VDD.n7275 0.053375
R11787 VDD.n7281 VDD.n7278 0.053375
R11788 VDD.n7284 VDD.n7281 0.053375
R11789 VDD.n7285 VDD.n7284 0.053375
R11790 VDD VDD.n7285 0.053375
R11791 VDD VDD.n7725 0.053375
R11792 VDD.n7725 VDD.n7722 0.053375
R11793 VDD.n7722 VDD.n7719 0.053375
R11794 VDD.n7719 VDD.n7716 0.053375
R11795 VDD.n7716 VDD.n7713 0.053375
R11796 VDD.n7713 VDD.n7710 0.053375
R11797 VDD.n7710 VDD.n7707 0.053375
R11798 VDD.n7703 VDD.n7700 0.053375
R11799 VDD.n7696 VDD.n7693 0.053375
R11800 VDD.n7693 VDD.n7690 0.053375
R11801 VDD.n7690 VDD.n7687 0.053375
R11802 VDD.n7687 VDD.n7684 0.053375
R11803 VDD.n7537 VDD.n7536 0.0528125
R11804 VDD.n7118 VDD.n7116 0.0516875
R11805 VDD.n7247 VDD.n7246 0.0516875
R11806 VDD.n324 VDD.n321 0.0505625
R11807 VDD.n369 VDD.n366 0.0505625
R11808 VDD.n7566 VDD.n7564 0.0505625
R11809 VDD.n7578 VDD.n7577 0.0505625
R11810 VDD.n7700 VDD.n7697 0.0505625
R11811 VDD.n7533 VDD.n7532 0.0483125
R11812 VDD.n576 VDD.n575 0.0483125
R11813 VDD.n634 VDD.n632 0.0483125
R11814 VDD.n1033 VDD.n1032 0.0483125
R11815 VDD.n570 VDD.n567 0.0483125
R11816 VDD.n7331 VDD.n7328 0.0460625
R11817 VDD.n7099 VDD.n7097 0.0460625
R11818 VDD.n448 VDD.n446 0.0449375
R11819 VDD.n7417 VDD.n7415 0.0449375
R11820 VDD.n7522 VDD.n7521 0.0449375
R11821 VDD.n6663 VDD.n6661 0.0426875
R11822 VDD.n811 VDD.n809 0.0426875
R11823 VDD.n6842 VDD.n6839 0.0426875
R11824 VDD.n999 VDD.n996 0.0426875
R11825 VDD.n6873 VDD.n6872 0.042125
R11826 VDD.n7559 VDD.n7558 0.041
R11827 VDD.n325 VDD.n324 0.0404375
R11828 VDD.n7024 VDD.n7023 0.0404375
R11829 VDD.n778 VDD.n570 0.039875
R11830 VDD.n7006 VDD.n7003 0.039875
R11831 VDD.n7341 VDD.n7340 0.0393125
R11832 VDD.n7109 VDD.n7105 0.0393125
R11833 VDD.n7260 VDD.n7257 0.0393125
R11834 VDD.n7062 VDD.n7059 0.03875
R11835 VDD.n133 VDD.n130 0.0359375
R11836 VDD.n182 VDD.n178 0.0359375
R11837 VDD.n6675 VDD.n6674 0.0359375
R11838 VDD.n823 VDD.n822 0.0359375
R11839 VDD.n6859 VDD.n6858 0.0359375
R11840 VDD.n7017 VDD.n7014 0.0359375
R11841 VDD.n7066 VDD.n7065 0.0359375
R11842 VDD.n317 VDD.n314 0.0348125
R11843 VDD.n379 VDD.n378 0.0348125
R11844 VDD.n7573 VDD.n7572 0.0348125
R11845 VDD.n7707 VDD.n7704 0.0348125
R11846 VDD.n123 VDD.n122 0.0336875
R11847 VDD.n192 VDD.n189 0.0336875
R11848 VDD.n6682 VDD.n6680 0.0336875
R11849 VDD.n830 VDD.n828 0.0336875
R11850 VDD.n6869 VDD.n6866 0.0336875
R11851 VDD.n7007 VDD.n7006 0.0336875
R11852 VDD.n7076 VDD.n7073 0.0336875
R11853 VDD.n7357 VDD.n7354 0.0325625
R11854 VDD.n6668 VDD.n6667 0.0325625
R11855 VDD.n816 VDD.n815 0.0325625
R11856 VDD.n581 VDD.n580 0.0325625
R11857 VDD.n629 VDD.n627 0.0325625
R11858 VDD.n6849 VDD.n6848 0.0325625
R11859 VDD.n1006 VDD.n1005 0.0325625
R11860 VDD.n1040 VDD.n1039 0.0325625
R11861 VDD.n563 VDD.n560 0.0325625
R11862 VDD.n443 VDD.n441 0.0291875
R11863 VDD.n7412 VDD.n7410 0.0291875
R11864 VDD.n353 VDD.n350 0.0291875
R11865 VDD.n7529 VDD.n7528 0.0291875
R11866 VDD.n7553 VDD.n7551 0.0291875
R11867 VDD.n386 VDD.n334 0.0280625
R11868 VDD.n3335 VDD.n3333 0.0269375
R11869 VDD.n3333 VDD.n3330 0.0269375
R11870 VDD.n3330 VDD.n3328 0.0269375
R11871 VDD.n3328 VDD.n3325 0.0269375
R11872 VDD.n5437 VDD.n5434 0.0269375
R11873 VDD.n5439 VDD.n5437 0.0269375
R11874 VDD.n5442 VDD.n5439 0.0269375
R11875 VDD.n5444 VDD.n5442 0.0269375
R11876 VDD.n5447 VDD.n5444 0.0269375
R11877 VDD.n5449 VDD.n5447 0.0269375
R11878 VDD.n5452 VDD.n5449 0.0269375
R11879 VDD.n5454 VDD.n5452 0.0269375
R11880 VDD.n5457 VDD.n5454 0.0269375
R11881 VDD.n5459 VDD.n5457 0.0269375
R11882 VDD.n5462 VDD.n5459 0.0269375
R11883 VDD.n5464 VDD.n5462 0.0269375
R11884 VDD.n5467 VDD.n5464 0.0269375
R11885 VDD.n5469 VDD.n5467 0.0269375
R11886 VDD.n5472 VDD.n5469 0.0269375
R11887 VDD.n5474 VDD.n5472 0.0269375
R11888 VDD.n5477 VDD.n5474 0.0269375
R11889 VDD.n5479 VDD.n5477 0.0269375
R11890 VDD.n5482 VDD.n5479 0.0269375
R11891 VDD.n5484 VDD.n5482 0.0269375
R11892 VDD.n5487 VDD.n5484 0.0269375
R11893 VDD.n5489 VDD.n5487 0.0269375
R11894 VDD.n5492 VDD.n5489 0.0269375
R11895 VDD.n5494 VDD.n5492 0.0269375
R11896 VDD.n5497 VDD.n5494 0.0269375
R11897 VDD.n5499 VDD.n5497 0.0269375
R11898 VDD.n5502 VDD.n5499 0.0269375
R11899 VDD.n5504 VDD.n5502 0.0269375
R11900 VDD.n5507 VDD.n5504 0.0269375
R11901 VDD.n5509 VDD.n5507 0.0269375
R11902 VDD.n5512 VDD.n5509 0.0269375
R11903 VDD.n5514 VDD.n5512 0.0269375
R11904 VDD.n5517 VDD.n5514 0.0269375
R11905 VDD.n5519 VDD.n5517 0.0269375
R11906 VDD.n5522 VDD.n5519 0.0269375
R11907 VDD.n5524 VDD.n5522 0.0269375
R11908 VDD.n5527 VDD.n5524 0.0269375
R11909 VDD.n5529 VDD.n5527 0.0269375
R11910 VDD.n5532 VDD.n5529 0.0269375
R11911 VDD.n5535 VDD.n5532 0.0269375
R11912 VDD.n5537 VDD.n5535 0.0269375
R11913 VDD.n5540 VDD.n5537 0.0269375
R11914 VDD.n3265 VDD.n3263 0.0269375
R11915 VDD.n3263 VDD.n3261 0.0269375
R11916 VDD.n3261 VDD.n3259 0.0269375
R11917 VDD.n3259 VDD.n3257 0.0269375
R11918 VDD.n5276 VDD.n5274 0.0269375
R11919 VDD.n5278 VDD.n5276 0.0269375
R11920 VDD.n5280 VDD.n5278 0.0269375
R11921 VDD.n5282 VDD.n5280 0.0269375
R11922 VDD.n5284 VDD.n5282 0.0269375
R11923 VDD.n5286 VDD.n5284 0.0269375
R11924 VDD.n5288 VDD.n5286 0.0269375
R11925 VDD.n5290 VDD.n5288 0.0269375
R11926 VDD.n5292 VDD.n5290 0.0269375
R11927 VDD.n5294 VDD.n5292 0.0269375
R11928 VDD.n5296 VDD.n5294 0.0269375
R11929 VDD.n5298 VDD.n5296 0.0269375
R11930 VDD.n5300 VDD.n5298 0.0269375
R11931 VDD.n5302 VDD.n5300 0.0269375
R11932 VDD.n5304 VDD.n5302 0.0269375
R11933 VDD.n5306 VDD.n5304 0.0269375
R11934 VDD.n5308 VDD.n5306 0.0269375
R11935 VDD.n5310 VDD.n5308 0.0269375
R11936 VDD.n5312 VDD.n5310 0.0269375
R11937 VDD.n5314 VDD.n5312 0.0269375
R11938 VDD.n5316 VDD.n5314 0.0269375
R11939 VDD.n5318 VDD.n5316 0.0269375
R11940 VDD.n5320 VDD.n5318 0.0269375
R11941 VDD.n5322 VDD.n5320 0.0269375
R11942 VDD.n5325 VDD.n5322 0.0269375
R11943 VDD.n5327 VDD.n5325 0.0269375
R11944 VDD.n5330 VDD.n5327 0.0269375
R11945 VDD.n5332 VDD.n5330 0.0269375
R11946 VDD.n5335 VDD.n5332 0.0269375
R11947 VDD.n5337 VDD.n5335 0.0269375
R11948 VDD.n5340 VDD.n5337 0.0269375
R11949 VDD.n5342 VDD.n5340 0.0269375
R11950 VDD.n5345 VDD.n5342 0.0269375
R11951 VDD.n5347 VDD.n5345 0.0269375
R11952 VDD.n5350 VDD.n5347 0.0269375
R11953 VDD.n5352 VDD.n5350 0.0269375
R11954 VDD.n5355 VDD.n5352 0.0269375
R11955 VDD.n5357 VDD.n5355 0.0269375
R11956 VDD.n5360 VDD.n5357 0.0269375
R11957 VDD.n5362 VDD.n5360 0.0269375
R11958 VDD.n5365 VDD.n5362 0.0269375
R11959 VDD.n5367 VDD.n5365 0.0269375
R11960 VDD.n2976 VDD.n2973 0.0269375
R11961 VDD.n4274 VDD.n4272 0.0269375
R11962 VDD.n4277 VDD.n4274 0.0269375
R11963 VDD.n4279 VDD.n4277 0.0269375
R11964 VDD.n4282 VDD.n4279 0.0269375
R11965 VDD.n4284 VDD.n4282 0.0269375
R11966 VDD.n4287 VDD.n4284 0.0269375
R11967 VDD.n4289 VDD.n4287 0.0269375
R11968 VDD.n4292 VDD.n4289 0.0269375
R11969 VDD.n4294 VDD.n4292 0.0269375
R11970 VDD.n4297 VDD.n4294 0.0269375
R11971 VDD.n4299 VDD.n4297 0.0269375
R11972 VDD.n4302 VDD.n4299 0.0269375
R11973 VDD.n4304 VDD.n4302 0.0269375
R11974 VDD.n4307 VDD.n4304 0.0269375
R11975 VDD.n4309 VDD.n4307 0.0269375
R11976 VDD.n4312 VDD.n4309 0.0269375
R11977 VDD.n4314 VDD.n4312 0.0269375
R11978 VDD.n4317 VDD.n4314 0.0269375
R11979 VDD.n4319 VDD.n4317 0.0269375
R11980 VDD.n4322 VDD.n4319 0.0269375
R11981 VDD.n4324 VDD.n4322 0.0269375
R11982 VDD.n4327 VDD.n4324 0.0269375
R11983 VDD.n4329 VDD.n4327 0.0269375
R11984 VDD.n4332 VDD.n4329 0.0269375
R11985 VDD.n4334 VDD.n4332 0.0269375
R11986 VDD.n4337 VDD.n4334 0.0269375
R11987 VDD.n4339 VDD.n4337 0.0269375
R11988 VDD.n4342 VDD.n4339 0.0269375
R11989 VDD.n4344 VDD.n4342 0.0269375
R11990 VDD.n4347 VDD.n4344 0.0269375
R11991 VDD.n4349 VDD.n4347 0.0269375
R11992 VDD.n4352 VDD.n4349 0.0269375
R11993 VDD.n4354 VDD.n4352 0.0269375
R11994 VDD.n4357 VDD.n4354 0.0269375
R11995 VDD.n4359 VDD.n4357 0.0269375
R11996 VDD.n4362 VDD.n4359 0.0269375
R11997 VDD.n4364 VDD.n4362 0.0269375
R11998 VDD.n4367 VDD.n4364 0.0269375
R11999 VDD.n4369 VDD.n4367 0.0269375
R12000 VDD.n4372 VDD.n4369 0.0269375
R12001 VDD.n4374 VDD.n4372 0.0269375
R12002 VDD.n4377 VDD.n4374 0.0269375
R12003 VDD.n4380 VDD.n4377 0.0269375
R12004 VDD.n4382 VDD.n4380 0.0269375
R12005 VDD.n4385 VDD.n4382 0.0269375
R12006 VDD.n2971 VDD.n2969 0.0269375
R12007 VDD.n4138 VDD.n4135 0.0269375
R12008 VDD.n4141 VDD.n4138 0.0269375
R12009 VDD.n4144 VDD.n4141 0.0269375
R12010 VDD.n4147 VDD.n4144 0.0269375
R12011 VDD.n4150 VDD.n4147 0.0269375
R12012 VDD.n4153 VDD.n4150 0.0269375
R12013 VDD.n4156 VDD.n4153 0.0269375
R12014 VDD.n4159 VDD.n4156 0.0269375
R12015 VDD.n4162 VDD.n4159 0.0269375
R12016 VDD.n4165 VDD.n4162 0.0269375
R12017 VDD.n4168 VDD.n4165 0.0269375
R12018 VDD.n4171 VDD.n4168 0.0269375
R12019 VDD.n4174 VDD.n4171 0.0269375
R12020 VDD.n4177 VDD.n4174 0.0269375
R12021 VDD.n4180 VDD.n4177 0.0269375
R12022 VDD.n4183 VDD.n4180 0.0269375
R12023 VDD.n4186 VDD.n4183 0.0269375
R12024 VDD.n4189 VDD.n4186 0.0269375
R12025 VDD.n4192 VDD.n4189 0.0269375
R12026 VDD.n4195 VDD.n4192 0.0269375
R12027 VDD.n4198 VDD.n4195 0.0269375
R12028 VDD.n4201 VDD.n4198 0.0269375
R12029 VDD.n4204 VDD.n4201 0.0269375
R12030 VDD.n4207 VDD.n4204 0.0269375
R12031 VDD.n4210 VDD.n4207 0.0269375
R12032 VDD.n4213 VDD.n4210 0.0269375
R12033 VDD.n4216 VDD.n4213 0.0269375
R12034 VDD.n4219 VDD.n4216 0.0269375
R12035 VDD.n4222 VDD.n4219 0.0269375
R12036 VDD.n4225 VDD.n4222 0.0269375
R12037 VDD.n4228 VDD.n4225 0.0269375
R12038 VDD.n4231 VDD.n4228 0.0269375
R12039 VDD.n4234 VDD.n4231 0.0269375
R12040 VDD.n4237 VDD.n4234 0.0269375
R12041 VDD.n4240 VDD.n4237 0.0269375
R12042 VDD.n4243 VDD.n4240 0.0269375
R12043 VDD.n4246 VDD.n4243 0.0269375
R12044 VDD.n4249 VDD.n4246 0.0269375
R12045 VDD.n4252 VDD.n4249 0.0269375
R12046 VDD.n4255 VDD.n4252 0.0269375
R12047 VDD.n4258 VDD.n4255 0.0269375
R12048 VDD.n4261 VDD.n4258 0.0269375
R12049 VDD.n4264 VDD.n4261 0.0269375
R12050 VDD.n4266 VDD.n4264 0.0269375
R12051 VDD.n4269 VDD.n4266 0.0269375
R12052 VDD.n3750 VDD.n3748 0.0269375
R12053 VDD.n3752 VDD.n3750 0.0269375
R12054 VDD.n3754 VDD.n3752 0.0269375
R12055 VDD.n3759 VDD.n3757 0.0269375
R12056 VDD.n3764 VDD.n3762 0.0269375
R12057 VDD.n3766 VDD.n3764 0.0269375
R12058 VDD.n3771 VDD.n3769 0.0269375
R12059 VDD.n3773 VDD.n3771 0.0269375
R12060 VDD.n3778 VDD.n3776 0.0269375
R12061 VDD.n3780 VDD.n3778 0.0269375
R12062 VDD.n3785 VDD.n3783 0.0269375
R12063 VDD.n3787 VDD.n3785 0.0269375
R12064 VDD.n3789 VDD.n3787 0.0269375
R12065 VDD.n3791 VDD.n3789 0.0269375
R12066 VDD.n3793 VDD.n3791 0.0269375
R12067 VDD.n3795 VDD.n3793 0.0269375
R12068 VDD.n3797 VDD.n3795 0.0269375
R12069 VDD.n3799 VDD.n3797 0.0269375
R12070 VDD.n3801 VDD.n3799 0.0269375
R12071 VDD.n3803 VDD.n3801 0.0269375
R12072 VDD.n3808 VDD.n3806 0.0269375
R12073 VDD.n3810 VDD.n3808 0.0269375
R12074 VDD.n3815 VDD.n3813 0.0269375
R12075 VDD.n3817 VDD.n3815 0.0269375
R12076 VDD.n3822 VDD.n3820 0.0269375
R12077 VDD.n3824 VDD.n3822 0.0269375
R12078 VDD.n3829 VDD.n3827 0.0269375
R12079 VDD.n3834 VDD.n3832 0.0269375
R12080 VDD.n3836 VDD.n3834 0.0269375
R12081 VDD.n3838 VDD.n3836 0.0269375
R12082 VDD.n3840 VDD.n3838 0.0269375
R12083 VDD.n3855 VDD.n3853 0.0269375
R12084 VDD.n3857 VDD.n3855 0.0269375
R12085 VDD.n3859 VDD.n3857 0.0269375
R12086 VDD.n3861 VDD.n3859 0.0269375
R12087 VDD.n3866 VDD.n3864 0.0269375
R12088 VDD.n3871 VDD.n3869 0.0269375
R12089 VDD.n3873 VDD.n3871 0.0269375
R12090 VDD.n3878 VDD.n3876 0.0269375
R12091 VDD.n3880 VDD.n3878 0.0269375
R12092 VDD.n3885 VDD.n3883 0.0269375
R12093 VDD.n3887 VDD.n3885 0.0269375
R12094 VDD.n3892 VDD.n3890 0.0269375
R12095 VDD.n3894 VDD.n3892 0.0269375
R12096 VDD.n3896 VDD.n3894 0.0269375
R12097 VDD.n3898 VDD.n3896 0.0269375
R12098 VDD.n3900 VDD.n3898 0.0269375
R12099 VDD.n3902 VDD.n3900 0.0269375
R12100 VDD.n3904 VDD.n3902 0.0269375
R12101 VDD.n3906 VDD.n3904 0.0269375
R12102 VDD.n3908 VDD.n3906 0.0269375
R12103 VDD.n3910 VDD.n3908 0.0269375
R12104 VDD.n3915 VDD.n3913 0.0269375
R12105 VDD.n3917 VDD.n3915 0.0269375
R12106 VDD.n3922 VDD.n3920 0.0269375
R12107 VDD.n3924 VDD.n3922 0.0269375
R12108 VDD.n3929 VDD.n3927 0.0269375
R12109 VDD.n3931 VDD.n3929 0.0269375
R12110 VDD.n3936 VDD.n3934 0.0269375
R12111 VDD.n3946 VDD.n3944 0.0269375
R12112 VDD.n3948 VDD.n3946 0.0269375
R12113 VDD.n3950 VDD.n3948 0.0269375
R12114 VDD.n6160 VDD.n6157 0.0269375
R12115 VDD.n6165 VDD.n6160 0.0269375
R12116 VDD.n6172 VDD.n6169 0.0269375
R12117 VDD.n6175 VDD.n6172 0.0269375
R12118 VDD.n6178 VDD.n6175 0.0269375
R12119 VDD.n6181 VDD.n6178 0.0269375
R12120 VDD.n6188 VDD.n6185 0.0269375
R12121 VDD.n6195 VDD.n6192 0.0269375
R12122 VDD.n6198 VDD.n6195 0.0269375
R12123 VDD.n6205 VDD.n6202 0.0269375
R12124 VDD.n6208 VDD.n6205 0.0269375
R12125 VDD.n6215 VDD.n6212 0.0269375
R12126 VDD.n6218 VDD.n6215 0.0269375
R12127 VDD.n6225 VDD.n6222 0.0269375
R12128 VDD.n6228 VDD.n6225 0.0269375
R12129 VDD.n6231 VDD.n6228 0.0269375
R12130 VDD.n6238 VDD.n6235 0.0269375
R12131 VDD.n6241 VDD.n6238 0.0269375
R12132 VDD.n6248 VDD.n6245 0.0269375
R12133 VDD.n6251 VDD.n6248 0.0269375
R12134 VDD.n6254 VDD.n6251 0.0269375
R12135 VDD.n6261 VDD.n6258 0.0269375
R12136 VDD.n6264 VDD.n6261 0.0269375
R12137 VDD.n6271 VDD.n6268 0.0269375
R12138 VDD.n6274 VDD.n6271 0.0269375
R12139 VDD.n6281 VDD.n6278 0.0269375
R12140 VDD.n6284 VDD.n6281 0.0269375
R12141 VDD.n6291 VDD.n6288 0.0269375
R12142 VDD.n6298 VDD.n6295 0.0269375
R12143 VDD.n6301 VDD.n6298 0.0269375
R12144 VDD.n6304 VDD.n6301 0.0269375
R12145 VDD.n6307 VDD.n6304 0.0269375
R12146 VDD.n6327 VDD.n6324 0.0269375
R12147 VDD.n6330 VDD.n6327 0.0269375
R12148 VDD.n6333 VDD.n6330 0.0269375
R12149 VDD.n6336 VDD.n6333 0.0269375
R12150 VDD.n6343 VDD.n6340 0.0269375
R12151 VDD.n6350 VDD.n6347 0.0269375
R12152 VDD.n6353 VDD.n6350 0.0269375
R12153 VDD.n6360 VDD.n6357 0.0269375
R12154 VDD.n6363 VDD.n6360 0.0269375
R12155 VDD.n6370 VDD.n6367 0.0269375
R12156 VDD.n6373 VDD.n6370 0.0269375
R12157 VDD.n6380 VDD.n6377 0.0269375
R12158 VDD.n6383 VDD.n6380 0.0269375
R12159 VDD.n6386 VDD.n6383 0.0269375
R12160 VDD.n6393 VDD.n6390 0.0269375
R12161 VDD.n6396 VDD.n6393 0.0269375
R12162 VDD.n6403 VDD.n6400 0.0269375
R12163 VDD.n6406 VDD.n6403 0.0269375
R12164 VDD.n6409 VDD.n6406 0.0269375
R12165 VDD.n6416 VDD.n6413 0.0269375
R12166 VDD.n6419 VDD.n6416 0.0269375
R12167 VDD.n6426 VDD.n6423 0.0269375
R12168 VDD.n6429 VDD.n6426 0.0269375
R12169 VDD.n6436 VDD.n6433 0.0269375
R12170 VDD.n6439 VDD.n6436 0.0269375
R12171 VDD.n6446 VDD.n6443 0.0269375
R12172 VDD.n6453 VDD.n6450 0.0269375
R12173 VDD.n6456 VDD.n6453 0.0269375
R12174 VDD.n6459 VDD.n6456 0.0269375
R12175 VDD.n3104 VDD.n3102 0.0269375
R12176 VDD.n3102 VDD.n3099 0.0269375
R12177 VDD.n4648 VDD.n4645 0.0269375
R12178 VDD.n4651 VDD.n4648 0.0269375
R12179 VDD.n4654 VDD.n4651 0.0269375
R12180 VDD.n4657 VDD.n4654 0.0269375
R12181 VDD.n4660 VDD.n4657 0.0269375
R12182 VDD.n4663 VDD.n4660 0.0269375
R12183 VDD.n4666 VDD.n4663 0.0269375
R12184 VDD.n4669 VDD.n4666 0.0269375
R12185 VDD.n4672 VDD.n4669 0.0269375
R12186 VDD.n4675 VDD.n4672 0.0269375
R12187 VDD.n4678 VDD.n4675 0.0269375
R12188 VDD.n4681 VDD.n4678 0.0269375
R12189 VDD.n4684 VDD.n4681 0.0269375
R12190 VDD.n4687 VDD.n4684 0.0269375
R12191 VDD.n4690 VDD.n4687 0.0269375
R12192 VDD.n4693 VDD.n4690 0.0269375
R12193 VDD.n4696 VDD.n4693 0.0269375
R12194 VDD.n4699 VDD.n4696 0.0269375
R12195 VDD.n4702 VDD.n4699 0.0269375
R12196 VDD.n4705 VDD.n4702 0.0269375
R12197 VDD.n4708 VDD.n4705 0.0269375
R12198 VDD.n4711 VDD.n4708 0.0269375
R12199 VDD.n4714 VDD.n4711 0.0269375
R12200 VDD.n4717 VDD.n4714 0.0269375
R12201 VDD.n4720 VDD.n4717 0.0269375
R12202 VDD.n4723 VDD.n4720 0.0269375
R12203 VDD.n4726 VDD.n4723 0.0269375
R12204 VDD.n4729 VDD.n4726 0.0269375
R12205 VDD.n4732 VDD.n4729 0.0269375
R12206 VDD.n4735 VDD.n4732 0.0269375
R12207 VDD.n4738 VDD.n4735 0.0269375
R12208 VDD.n4741 VDD.n4738 0.0269375
R12209 VDD.n4744 VDD.n4741 0.0269375
R12210 VDD.n4747 VDD.n4744 0.0269375
R12211 VDD.n4750 VDD.n4747 0.0269375
R12212 VDD.n4753 VDD.n4750 0.0269375
R12213 VDD.n4756 VDD.n4753 0.0269375
R12214 VDD.n4759 VDD.n4756 0.0269375
R12215 VDD.n4762 VDD.n4759 0.0269375
R12216 VDD.n4765 VDD.n4762 0.0269375
R12217 VDD.n4768 VDD.n4765 0.0269375
R12218 VDD.n4771 VDD.n4768 0.0269375
R12219 VDD.n4773 VDD.n4771 0.0269375
R12220 VDD.n4776 VDD.n4773 0.0269375
R12221 VDD.n3112 VDD.n3109 0.0269375
R12222 VDD.n3109 VDD.n3107 0.0269375
R12223 VDD.n4781 VDD.n4778 0.0269375
R12224 VDD.n4783 VDD.n4781 0.0269375
R12225 VDD.n4786 VDD.n4783 0.0269375
R12226 VDD.n4788 VDD.n4786 0.0269375
R12227 VDD.n4791 VDD.n4788 0.0269375
R12228 VDD.n4793 VDD.n4791 0.0269375
R12229 VDD.n4796 VDD.n4793 0.0269375
R12230 VDD.n4798 VDD.n4796 0.0269375
R12231 VDD.n4801 VDD.n4798 0.0269375
R12232 VDD.n4803 VDD.n4801 0.0269375
R12233 VDD.n4806 VDD.n4803 0.0269375
R12234 VDD.n4808 VDD.n4806 0.0269375
R12235 VDD.n4811 VDD.n4808 0.0269375
R12236 VDD.n4813 VDD.n4811 0.0269375
R12237 VDD.n4816 VDD.n4813 0.0269375
R12238 VDD.n4818 VDD.n4816 0.0269375
R12239 VDD.n4821 VDD.n4818 0.0269375
R12240 VDD.n4823 VDD.n4821 0.0269375
R12241 VDD.n4826 VDD.n4823 0.0269375
R12242 VDD.n4828 VDD.n4826 0.0269375
R12243 VDD.n4831 VDD.n4828 0.0269375
R12244 VDD.n4833 VDD.n4831 0.0269375
R12245 VDD.n4836 VDD.n4833 0.0269375
R12246 VDD.n4838 VDD.n4836 0.0269375
R12247 VDD.n4841 VDD.n4838 0.0269375
R12248 VDD.n4843 VDD.n4841 0.0269375
R12249 VDD.n4846 VDD.n4843 0.0269375
R12250 VDD.n4848 VDD.n4846 0.0269375
R12251 VDD.n4851 VDD.n4848 0.0269375
R12252 VDD.n4853 VDD.n4851 0.0269375
R12253 VDD.n4856 VDD.n4853 0.0269375
R12254 VDD.n4858 VDD.n4856 0.0269375
R12255 VDD.n4861 VDD.n4858 0.0269375
R12256 VDD.n4863 VDD.n4861 0.0269375
R12257 VDD.n4866 VDD.n4863 0.0269375
R12258 VDD.n4868 VDD.n4866 0.0269375
R12259 VDD.n4871 VDD.n4868 0.0269375
R12260 VDD.n4873 VDD.n4871 0.0269375
R12261 VDD.n4876 VDD.n4873 0.0269375
R12262 VDD.n4878 VDD.n4876 0.0269375
R12263 VDD.n4881 VDD.n4878 0.0269375
R12264 VDD.n4884 VDD.n4881 0.0269375
R12265 VDD.n4886 VDD.n4884 0.0269375
R12266 VDD.n4889 VDD.n4886 0.0269375
R12267 VDD.n3544 VDD.n3542 0.0269375
R12268 VDD.n3546 VDD.n3544 0.0269375
R12269 VDD.n3548 VDD.n3546 0.0269375
R12270 VDD.n3553 VDD.n3551 0.0269375
R12271 VDD.n3558 VDD.n3556 0.0269375
R12272 VDD.n3560 VDD.n3558 0.0269375
R12273 VDD.n3565 VDD.n3563 0.0269375
R12274 VDD.n3567 VDD.n3565 0.0269375
R12275 VDD.n3572 VDD.n3570 0.0269375
R12276 VDD.n3574 VDD.n3572 0.0269375
R12277 VDD.n3579 VDD.n3577 0.0269375
R12278 VDD.n3581 VDD.n3579 0.0269375
R12279 VDD.n3583 VDD.n3581 0.0269375
R12280 VDD.n3585 VDD.n3583 0.0269375
R12281 VDD.n3587 VDD.n3585 0.0269375
R12282 VDD.n3589 VDD.n3587 0.0269375
R12283 VDD.n3591 VDD.n3589 0.0269375
R12284 VDD.n3593 VDD.n3591 0.0269375
R12285 VDD.n3595 VDD.n3593 0.0269375
R12286 VDD.n3597 VDD.n3595 0.0269375
R12287 VDD.n3602 VDD.n3600 0.0269375
R12288 VDD.n3604 VDD.n3602 0.0269375
R12289 VDD.n3609 VDD.n3607 0.0269375
R12290 VDD.n3611 VDD.n3609 0.0269375
R12291 VDD.n3616 VDD.n3614 0.0269375
R12292 VDD.n3618 VDD.n3616 0.0269375
R12293 VDD.n3623 VDD.n3621 0.0269375
R12294 VDD.n3628 VDD.n3626 0.0269375
R12295 VDD.n3630 VDD.n3628 0.0269375
R12296 VDD.n3632 VDD.n3630 0.0269375
R12297 VDD.n3634 VDD.n3632 0.0269375
R12298 VDD.n3650 VDD.n3648 0.0269375
R12299 VDD.n3652 VDD.n3650 0.0269375
R12300 VDD.n3654 VDD.n3652 0.0269375
R12301 VDD.n3656 VDD.n3654 0.0269375
R12302 VDD.n3661 VDD.n3659 0.0269375
R12303 VDD.n3666 VDD.n3664 0.0269375
R12304 VDD.n3668 VDD.n3666 0.0269375
R12305 VDD.n3673 VDD.n3671 0.0269375
R12306 VDD.n3675 VDD.n3673 0.0269375
R12307 VDD.n3680 VDD.n3678 0.0269375
R12308 VDD.n3682 VDD.n3680 0.0269375
R12309 VDD.n3687 VDD.n3685 0.0269375
R12310 VDD.n3689 VDD.n3687 0.0269375
R12311 VDD.n3691 VDD.n3689 0.0269375
R12312 VDD.n3693 VDD.n3691 0.0269375
R12313 VDD.n3695 VDD.n3693 0.0269375
R12314 VDD.n3697 VDD.n3695 0.0269375
R12315 VDD.n3699 VDD.n3697 0.0269375
R12316 VDD.n3701 VDD.n3699 0.0269375
R12317 VDD.n3703 VDD.n3701 0.0269375
R12318 VDD.n3705 VDD.n3703 0.0269375
R12319 VDD.n3710 VDD.n3708 0.0269375
R12320 VDD.n3712 VDD.n3710 0.0269375
R12321 VDD.n3717 VDD.n3715 0.0269375
R12322 VDD.n3719 VDD.n3717 0.0269375
R12323 VDD.n3724 VDD.n3722 0.0269375
R12324 VDD.n3726 VDD.n3724 0.0269375
R12325 VDD.n3731 VDD.n3729 0.0269375
R12326 VDD.n3741 VDD.n3739 0.0269375
R12327 VDD.n3743 VDD.n3741 0.0269375
R12328 VDD.n3745 VDD.n3743 0.0269375
R12329 VDD.n5858 VDD.n5855 0.0269375
R12330 VDD.n5863 VDD.n5858 0.0269375
R12331 VDD.n5870 VDD.n5867 0.0269375
R12332 VDD.n5873 VDD.n5870 0.0269375
R12333 VDD.n5876 VDD.n5873 0.0269375
R12334 VDD.n5879 VDD.n5876 0.0269375
R12335 VDD.n5886 VDD.n5883 0.0269375
R12336 VDD.n5893 VDD.n5890 0.0269375
R12337 VDD.n5896 VDD.n5893 0.0269375
R12338 VDD.n5903 VDD.n5900 0.0269375
R12339 VDD.n5906 VDD.n5903 0.0269375
R12340 VDD.n5913 VDD.n5910 0.0269375
R12341 VDD.n5916 VDD.n5913 0.0269375
R12342 VDD.n5923 VDD.n5920 0.0269375
R12343 VDD.n5926 VDD.n5923 0.0269375
R12344 VDD.n5929 VDD.n5926 0.0269375
R12345 VDD.n5936 VDD.n5933 0.0269375
R12346 VDD.n5939 VDD.n5936 0.0269375
R12347 VDD.n5946 VDD.n5943 0.0269375
R12348 VDD.n5949 VDD.n5946 0.0269375
R12349 VDD.n5952 VDD.n5949 0.0269375
R12350 VDD.n5959 VDD.n5956 0.0269375
R12351 VDD.n5962 VDD.n5959 0.0269375
R12352 VDD.n5969 VDD.n5966 0.0269375
R12353 VDD.n5972 VDD.n5969 0.0269375
R12354 VDD.n5979 VDD.n5976 0.0269375
R12355 VDD.n5982 VDD.n5979 0.0269375
R12356 VDD.n5989 VDD.n5986 0.0269375
R12357 VDD.n5996 VDD.n5993 0.0269375
R12358 VDD.n5999 VDD.n5996 0.0269375
R12359 VDD.n6002 VDD.n5999 0.0269375
R12360 VDD.n6005 VDD.n6002 0.0269375
R12361 VDD.n6025 VDD.n6022 0.0269375
R12362 VDD.n6028 VDD.n6025 0.0269375
R12363 VDD.n6031 VDD.n6028 0.0269375
R12364 VDD.n6034 VDD.n6031 0.0269375
R12365 VDD.n6041 VDD.n6038 0.0269375
R12366 VDD.n6048 VDD.n6045 0.0269375
R12367 VDD.n6051 VDD.n6048 0.0269375
R12368 VDD.n6058 VDD.n6055 0.0269375
R12369 VDD.n6061 VDD.n6058 0.0269375
R12370 VDD.n6068 VDD.n6065 0.0269375
R12371 VDD.n6071 VDD.n6068 0.0269375
R12372 VDD.n6078 VDD.n6075 0.0269375
R12373 VDD.n6081 VDD.n6078 0.0269375
R12374 VDD.n6084 VDD.n6081 0.0269375
R12375 VDD.n6091 VDD.n6088 0.0269375
R12376 VDD.n6094 VDD.n6091 0.0269375
R12377 VDD.n6101 VDD.n6098 0.0269375
R12378 VDD.n6104 VDD.n6101 0.0269375
R12379 VDD.n6107 VDD.n6104 0.0269375
R12380 VDD.n6114 VDD.n6111 0.0269375
R12381 VDD.n6117 VDD.n6114 0.0269375
R12382 VDD.n6124 VDD.n6121 0.0269375
R12383 VDD.n6127 VDD.n6124 0.0269375
R12384 VDD.n6134 VDD.n6131 0.0269375
R12385 VDD.n6137 VDD.n6134 0.0269375
R12386 VDD.n6144 VDD.n6141 0.0269375
R12387 VDD.n6151 VDD.n6148 0.0269375
R12388 VDD.n6154 VDD.n6151 0.0269375
R12389 VDD.n6157 VDD.n6154 0.0269375
R12390 VDD.n3254 VDD.n3252 0.0269375
R12391 VDD.n3252 VDD.n3249 0.0269375
R12392 VDD.n3249 VDD.n3246 0.0269375
R12393 VDD.n3246 VDD.n3243 0.0269375
R12394 VDD.n5149 VDD.n5146 0.0269375
R12395 VDD.n5152 VDD.n5149 0.0269375
R12396 VDD.n5155 VDD.n5152 0.0269375
R12397 VDD.n5158 VDD.n5155 0.0269375
R12398 VDD.n5161 VDD.n5158 0.0269375
R12399 VDD.n5164 VDD.n5161 0.0269375
R12400 VDD.n5167 VDD.n5164 0.0269375
R12401 VDD.n5170 VDD.n5167 0.0269375
R12402 VDD.n5173 VDD.n5170 0.0269375
R12403 VDD.n5176 VDD.n5173 0.0269375
R12404 VDD.n5179 VDD.n5176 0.0269375
R12405 VDD.n5182 VDD.n5179 0.0269375
R12406 VDD.n5185 VDD.n5182 0.0269375
R12407 VDD.n5188 VDD.n5185 0.0269375
R12408 VDD.n5191 VDD.n5188 0.0269375
R12409 VDD.n5194 VDD.n5191 0.0269375
R12410 VDD.n5197 VDD.n5194 0.0269375
R12411 VDD.n5200 VDD.n5197 0.0269375
R12412 VDD.n5203 VDD.n5200 0.0269375
R12413 VDD.n5206 VDD.n5203 0.0269375
R12414 VDD.n5209 VDD.n5206 0.0269375
R12415 VDD.n5212 VDD.n5209 0.0269375
R12416 VDD.n5215 VDD.n5212 0.0269375
R12417 VDD.n5218 VDD.n5215 0.0269375
R12418 VDD.n5221 VDD.n5218 0.0269375
R12419 VDD.n5224 VDD.n5221 0.0269375
R12420 VDD.n5227 VDD.n5224 0.0269375
R12421 VDD.n5230 VDD.n5227 0.0269375
R12422 VDD.n5233 VDD.n5230 0.0269375
R12423 VDD.n5236 VDD.n5233 0.0269375
R12424 VDD.n5239 VDD.n5236 0.0269375
R12425 VDD.n5242 VDD.n5239 0.0269375
R12426 VDD.n5245 VDD.n5242 0.0269375
R12427 VDD.n5248 VDD.n5245 0.0269375
R12428 VDD.n5251 VDD.n5248 0.0269375
R12429 VDD.n5254 VDD.n5251 0.0269375
R12430 VDD.n5257 VDD.n5254 0.0269375
R12431 VDD.n5260 VDD.n5257 0.0269375
R12432 VDD.n5263 VDD.n5260 0.0269375
R12433 VDD.n5266 VDD.n5263 0.0269375
R12434 VDD.n5268 VDD.n5266 0.0269375
R12435 VDD.n5271 VDD.n5268 0.0269375
R12436 VDD.n5551 VDD.n5548 0.0269375
R12437 VDD.n5554 VDD.n5551 0.0269375
R12438 VDD.n5557 VDD.n5554 0.0269375
R12439 VDD.n5560 VDD.n5557 0.0269375
R12440 VDD.n5570 VDD.n5567 0.0269375
R12441 VDD.n5577 VDD.n5574 0.0269375
R12442 VDD.n5580 VDD.n5577 0.0269375
R12443 VDD.n5587 VDD.n5584 0.0269375
R12444 VDD.n5590 VDD.n5587 0.0269375
R12445 VDD.n5597 VDD.n5594 0.0269375
R12446 VDD.n5600 VDD.n5597 0.0269375
R12447 VDD.n5607 VDD.n5604 0.0269375
R12448 VDD.n5610 VDD.n5607 0.0269375
R12449 VDD.n5613 VDD.n5610 0.0269375
R12450 VDD.n5620 VDD.n5617 0.0269375
R12451 VDD.n5623 VDD.n5620 0.0269375
R12452 VDD.n5630 VDD.n5627 0.0269375
R12453 VDD.n5633 VDD.n5630 0.0269375
R12454 VDD.n5636 VDD.n5633 0.0269375
R12455 VDD.n5643 VDD.n5640 0.0269375
R12456 VDD.n5646 VDD.n5643 0.0269375
R12457 VDD.n5653 VDD.n5650 0.0269375
R12458 VDD.n5656 VDD.n5653 0.0269375
R12459 VDD.n5663 VDD.n5660 0.0269375
R12460 VDD.n5666 VDD.n5663 0.0269375
R12461 VDD.n5673 VDD.n5670 0.0269375
R12462 VDD.n5680 VDD.n5677 0.0269375
R12463 VDD.n5683 VDD.n5680 0.0269375
R12464 VDD.n5686 VDD.n5683 0.0269375
R12465 VDD.n5689 VDD.n5686 0.0269375
R12466 VDD.n5726 VDD.n5723 0.0269375
R12467 VDD.n5729 VDD.n5726 0.0269375
R12468 VDD.n5732 VDD.n5729 0.0269375
R12469 VDD.n5739 VDD.n5736 0.0269375
R12470 VDD.n5746 VDD.n5743 0.0269375
R12471 VDD.n5749 VDD.n5746 0.0269375
R12472 VDD.n5756 VDD.n5753 0.0269375
R12473 VDD.n5759 VDD.n5756 0.0269375
R12474 VDD.n5766 VDD.n5763 0.0269375
R12475 VDD.n5769 VDD.n5766 0.0269375
R12476 VDD.n5776 VDD.n5773 0.0269375
R12477 VDD.n5779 VDD.n5776 0.0269375
R12478 VDD.n5782 VDD.n5779 0.0269375
R12479 VDD.n5789 VDD.n5786 0.0269375
R12480 VDD.n5792 VDD.n5789 0.0269375
R12481 VDD.n5799 VDD.n5796 0.0269375
R12482 VDD.n5802 VDD.n5799 0.0269375
R12483 VDD.n5805 VDD.n5802 0.0269375
R12484 VDD.n5812 VDD.n5809 0.0269375
R12485 VDD.n5815 VDD.n5812 0.0269375
R12486 VDD.n5822 VDD.n5819 0.0269375
R12487 VDD.n5825 VDD.n5822 0.0269375
R12488 VDD.n5832 VDD.n5829 0.0269375
R12489 VDD.n5835 VDD.n5832 0.0269375
R12490 VDD.n5842 VDD.n5839 0.0269375
R12491 VDD.n5849 VDD.n5846 0.0269375
R12492 VDD.n5852 VDD.n5849 0.0269375
R12493 VDD.n5855 VDD.n5852 0.0269375
R12494 VDD.n3343 VDD.n3341 0.0269375
R12495 VDD.n3345 VDD.n3343 0.0269375
R12496 VDD.n3347 VDD.n3345 0.0269375
R12497 VDD.n3349 VDD.n3347 0.0269375
R12498 VDD.n3354 VDD.n3352 0.0269375
R12499 VDD.n3359 VDD.n3357 0.0269375
R12500 VDD.n3361 VDD.n3359 0.0269375
R12501 VDD.n3366 VDD.n3364 0.0269375
R12502 VDD.n3368 VDD.n3366 0.0269375
R12503 VDD.n3373 VDD.n3371 0.0269375
R12504 VDD.n3375 VDD.n3373 0.0269375
R12505 VDD.n3380 VDD.n3378 0.0269375
R12506 VDD.n3382 VDD.n3380 0.0269375
R12507 VDD.n3384 VDD.n3382 0.0269375
R12508 VDD.n3386 VDD.n3384 0.0269375
R12509 VDD.n3388 VDD.n3386 0.0269375
R12510 VDD.n3390 VDD.n3388 0.0269375
R12511 VDD.n3392 VDD.n3390 0.0269375
R12512 VDD.n3394 VDD.n3392 0.0269375
R12513 VDD.n3396 VDD.n3394 0.0269375
R12514 VDD.n3398 VDD.n3396 0.0269375
R12515 VDD.n3403 VDD.n3401 0.0269375
R12516 VDD.n3405 VDD.n3403 0.0269375
R12517 VDD.n3410 VDD.n3408 0.0269375
R12518 VDD.n3412 VDD.n3410 0.0269375
R12519 VDD.n3417 VDD.n3415 0.0269375
R12520 VDD.n3419 VDD.n3417 0.0269375
R12521 VDD.n3424 VDD.n3422 0.0269375
R12522 VDD.n3429 VDD.n3427 0.0269375
R12523 VDD.n3431 VDD.n3429 0.0269375
R12524 VDD.n3433 VDD.n3431 0.0269375
R12525 VDD.n3435 VDD.n3433 0.0269375
R12526 VDD.n3449 VDD.n3447 0.0269375
R12527 VDD.n3451 VDD.n3449 0.0269375
R12528 VDD.n3453 VDD.n3451 0.0269375
R12529 VDD.n3455 VDD.n3453 0.0269375
R12530 VDD.n3460 VDD.n3458 0.0269375
R12531 VDD.n3465 VDD.n3463 0.0269375
R12532 VDD.n3467 VDD.n3465 0.0269375
R12533 VDD.n3472 VDD.n3470 0.0269375
R12534 VDD.n3474 VDD.n3472 0.0269375
R12535 VDD.n3479 VDD.n3477 0.0269375
R12536 VDD.n3481 VDD.n3479 0.0269375
R12537 VDD.n3486 VDD.n3484 0.0269375
R12538 VDD.n3488 VDD.n3486 0.0269375
R12539 VDD.n3490 VDD.n3488 0.0269375
R12540 VDD.n3492 VDD.n3490 0.0269375
R12541 VDD.n3494 VDD.n3492 0.0269375
R12542 VDD.n3496 VDD.n3494 0.0269375
R12543 VDD.n3498 VDD.n3496 0.0269375
R12544 VDD.n3500 VDD.n3498 0.0269375
R12545 VDD.n3502 VDD.n3500 0.0269375
R12546 VDD.n3504 VDD.n3502 0.0269375
R12547 VDD.n3509 VDD.n3507 0.0269375
R12548 VDD.n3511 VDD.n3509 0.0269375
R12549 VDD.n3516 VDD.n3514 0.0269375
R12550 VDD.n3518 VDD.n3516 0.0269375
R12551 VDD.n3523 VDD.n3521 0.0269375
R12552 VDD.n3525 VDD.n3523 0.0269375
R12553 VDD.n3530 VDD.n3528 0.0269375
R12554 VDD.n3535 VDD.n3533 0.0269375
R12555 VDD.n3537 VDD.n3535 0.0269375
R12556 VDD.n3539 VDD.n3537 0.0269375
R12557 VDD.n2698 VDD.n2695 0.0269375
R12558 VDD.n2701 VDD.n2698 0.0269375
R12559 VDD.n2704 VDD.n2701 0.0269375
R12560 VDD.n2707 VDD.n2704 0.0269375
R12561 VDD.n2710 VDD.n2707 0.0269375
R12562 VDD.n2713 VDD.n2710 0.0269375
R12563 VDD.n2716 VDD.n2713 0.0269375
R12564 VDD.n2719 VDD.n2716 0.0269375
R12565 VDD.n2722 VDD.n2719 0.0269375
R12566 VDD.n2725 VDD.n2722 0.0269375
R12567 VDD.n2728 VDD.n2725 0.0269375
R12568 VDD.n2731 VDD.n2728 0.0269375
R12569 VDD.n2734 VDD.n2731 0.0269375
R12570 VDD.n2737 VDD.n2734 0.0269375
R12571 VDD.n2740 VDD.n2737 0.0269375
R12572 VDD.n2743 VDD.n2740 0.0269375
R12573 VDD.n2746 VDD.n2743 0.0269375
R12574 VDD.n2749 VDD.n2746 0.0269375
R12575 VDD.n2752 VDD.n2749 0.0269375
R12576 VDD.n2755 VDD.n2752 0.0269375
R12577 VDD.n2758 VDD.n2755 0.0269375
R12578 VDD.n2761 VDD.n2758 0.0269375
R12579 VDD.n2764 VDD.n2761 0.0269375
R12580 VDD.n2767 VDD.n2764 0.0269375
R12581 VDD.n2770 VDD.n2767 0.0269375
R12582 VDD.n2773 VDD.n2770 0.0269375
R12583 VDD.n2776 VDD.n2773 0.0269375
R12584 VDD.n2779 VDD.n2776 0.0269375
R12585 VDD.n2782 VDD.n2779 0.0269375
R12586 VDD.n2785 VDD.n2782 0.0269375
R12587 VDD.n2788 VDD.n2785 0.0269375
R12588 VDD.n2791 VDD.n2788 0.0269375
R12589 VDD.n2794 VDD.n2791 0.0269375
R12590 VDD.n2797 VDD.n2794 0.0269375
R12591 VDD.n2800 VDD.n2797 0.0269375
R12592 VDD.n2803 VDD.n2800 0.0269375
R12593 VDD.n2806 VDD.n2803 0.0269375
R12594 VDD.n2809 VDD.n2806 0.0269375
R12595 VDD.n2812 VDD.n2809 0.0269375
R12596 VDD.n2815 VDD.n2812 0.0269375
R12597 VDD.n2818 VDD.n2815 0.0269375
R12598 VDD.n2821 VDD.n2818 0.0269375
R12599 VDD.n2824 VDD.n2821 0.0269375
R12600 VDD.n2827 VDD.n2824 0.0269375
R12601 VDD.n2830 VDD.n2827 0.0269375
R12602 VDD.n2833 VDD.n2830 0.0269375
R12603 VDD.n2836 VDD.n2833 0.0269375
R12604 VDD.n3954 VDD.n3952 0.0269375
R12605 VDD.n2598 VDD.n2596 0.0269375
R12606 VDD.n2603 VDD.n2601 0.0269375
R12607 VDD.n2608 VDD.n2606 0.0269375
R12608 VDD.n2610 VDD.n2608 0.0269375
R12609 VDD.n2615 VDD.n2613 0.0269375
R12610 VDD.n2617 VDD.n2615 0.0269375
R12611 VDD.n2622 VDD.n2620 0.0269375
R12612 VDD.n2624 VDD.n2622 0.0269375
R12613 VDD.n2629 VDD.n2627 0.0269375
R12614 VDD.n2631 VDD.n2629 0.0269375
R12615 VDD.n2633 VDD.n2631 0.0269375
R12616 VDD.n2635 VDD.n2633 0.0269375
R12617 VDD.n2637 VDD.n2635 0.0269375
R12618 VDD.n2639 VDD.n2637 0.0269375
R12619 VDD.n2641 VDD.n2639 0.0269375
R12620 VDD.n2643 VDD.n2641 0.0269375
R12621 VDD.n2645 VDD.n2643 0.0269375
R12622 VDD.n2647 VDD.n2645 0.0269375
R12623 VDD.n2652 VDD.n2650 0.0269375
R12624 VDD.n2654 VDD.n2652 0.0269375
R12625 VDD.n2659 VDD.n2657 0.0269375
R12626 VDD.n2661 VDD.n2659 0.0269375
R12627 VDD.n2666 VDD.n2664 0.0269375
R12628 VDD.n2668 VDD.n2666 0.0269375
R12629 VDD.n2673 VDD.n2671 0.0269375
R12630 VDD.n2683 VDD.n2681 0.0269375
R12631 VDD.n2685 VDD.n2683 0.0269375
R12632 VDD.n2687 VDD.n2685 0.0269375
R12633 VDD.n2689 VDD.n2687 0.0269375
R12634 VDD.n6489 VDD.n6486 0.0269375
R12635 VDD.n6492 VDD.n6489 0.0269375
R12636 VDD.n6495 VDD.n6492 0.0269375
R12637 VDD.n6502 VDD.n6499 0.0269375
R12638 VDD.n6509 VDD.n6506 0.0269375
R12639 VDD.n6512 VDD.n6509 0.0269375
R12640 VDD.n6519 VDD.n6516 0.0269375
R12641 VDD.n6522 VDD.n6519 0.0269375
R12642 VDD.n6529 VDD.n6526 0.0269375
R12643 VDD.n6532 VDD.n6529 0.0269375
R12644 VDD.n6539 VDD.n6536 0.0269375
R12645 VDD.n6542 VDD.n6539 0.0269375
R12646 VDD.n6545 VDD.n6542 0.0269375
R12647 VDD.n6552 VDD.n6549 0.0269375
R12648 VDD.n6555 VDD.n6552 0.0269375
R12649 VDD.n6562 VDD.n6559 0.0269375
R12650 VDD.n6565 VDD.n6562 0.0269375
R12651 VDD.n6568 VDD.n6565 0.0269375
R12652 VDD.n6575 VDD.n6572 0.0269375
R12653 VDD.n6578 VDD.n6575 0.0269375
R12654 VDD.n6585 VDD.n6582 0.0269375
R12655 VDD.n6588 VDD.n6585 0.0269375
R12656 VDD.n6595 VDD.n6592 0.0269375
R12657 VDD.n6598 VDD.n6595 0.0269375
R12658 VDD.n6605 VDD.n6602 0.0269375
R12659 VDD.n6612 VDD.n6609 0.0269375
R12660 VDD.n6615 VDD.n6612 0.0269375
R12661 VDD.n6618 VDD.n6615 0.0269375
R12662 VDD.n6621 VDD.n6618 0.0269375
R12663 VDD.n2039 VDD.n2037 0.0269375
R12664 VDD.n2037 VDD.n2034 0.0269375
R12665 VDD.n2034 VDD.n2032 0.0269375
R12666 VDD.n2032 VDD.n2029 0.0269375
R12667 VDD.n2029 VDD.n2027 0.0269375
R12668 VDD.n2027 VDD.n2024 0.0269375
R12669 VDD.n2024 VDD.n2022 0.0269375
R12670 VDD.n2022 VDD.n2019 0.0269375
R12671 VDD.n2019 VDD.n2017 0.0269375
R12672 VDD.n2017 VDD.n2014 0.0269375
R12673 VDD.n2014 VDD.n2012 0.0269375
R12674 VDD.n2012 VDD.n2009 0.0269375
R12675 VDD.n2009 VDD.n2007 0.0269375
R12676 VDD.n2007 VDD.n2004 0.0269375
R12677 VDD.n2004 VDD.n2002 0.0269375
R12678 VDD.n2002 VDD.n1999 0.0269375
R12679 VDD.n1999 VDD.n1997 0.0269375
R12680 VDD.n1997 VDD.n1994 0.0269375
R12681 VDD.n1994 VDD.n1992 0.0269375
R12682 VDD.n1992 VDD.n1989 0.0269375
R12683 VDD.n1989 VDD.n1987 0.0269375
R12684 VDD.n1987 VDD.n1985 0.0269375
R12685 VDD.n1985 VDD.n1983 0.0269375
R12686 VDD.n1983 VDD.n1981 0.0269375
R12687 VDD.n1981 VDD.n1979 0.0269375
R12688 VDD.n1979 VDD.n1977 0.0269375
R12689 VDD.n1977 VDD.n1975 0.0269375
R12690 VDD.n1975 VDD.n1973 0.0269375
R12691 VDD.n1973 VDD.n1971 0.0269375
R12692 VDD.n1971 VDD.n1969 0.0269375
R12693 VDD.n1969 VDD.n1967 0.0269375
R12694 VDD.n1967 VDD.n1965 0.0269375
R12695 VDD.n1965 VDD.n1963 0.0269375
R12696 VDD.n1963 VDD.n1961 0.0269375
R12697 VDD.n1961 VDD.n1959 0.0269375
R12698 VDD.n1959 VDD.n1957 0.0269375
R12699 VDD.n1957 VDD.n1955 0.0269375
R12700 VDD.n1955 VDD.n1953 0.0269375
R12701 VDD.n1953 VDD.n1951 0.0269375
R12702 VDD.n1951 VDD.n1949 0.0269375
R12703 VDD.n1949 VDD.n1947 0.0269375
R12704 VDD.n1947 VDD.n1945 0.0269375
R12705 VDD.n1945 VDD.n1943 0.0269375
R12706 VDD.n1943 VDD.n1941 0.0269375
R12707 VDD.n1941 VDD.n1939 0.0269375
R12708 VDD.n1935 VDD.n1933 0.0269375
R12709 VDD.n1933 VDD.n1930 0.0269375
R12710 VDD.n1930 VDD.n1927 0.0269375
R12711 VDD.n1927 VDD.n1924 0.0269375
R12712 VDD.n1924 VDD.n1921 0.0269375
R12713 VDD.n1921 VDD.n1918 0.0269375
R12714 VDD.n1918 VDD.n1915 0.0269375
R12715 VDD.n1915 VDD.n1912 0.0269375
R12716 VDD.n1912 VDD.n1909 0.0269375
R12717 VDD.n1909 VDD.n1906 0.0269375
R12718 VDD.n1906 VDD.n1903 0.0269375
R12719 VDD.n1903 VDD.n1900 0.0269375
R12720 VDD.n1900 VDD.n1897 0.0269375
R12721 VDD.n1897 VDD.n1894 0.0269375
R12722 VDD.n1894 VDD.n1891 0.0269375
R12723 VDD.n1891 VDD.n1888 0.0269375
R12724 VDD.n1888 VDD.n1885 0.0269375
R12725 VDD.n1885 VDD.n1882 0.0269375
R12726 VDD.n1882 VDD.n1879 0.0269375
R12727 VDD.n1879 VDD.n1876 0.0269375
R12728 VDD.n1876 VDD.n1873 0.0269375
R12729 VDD.n1873 VDD.n1870 0.0269375
R12730 VDD.n1870 VDD.n1867 0.0269375
R12731 VDD.n1867 VDD.n1864 0.0269375
R12732 VDD.n1864 VDD.n1861 0.0269375
R12733 VDD.n1861 VDD.n1858 0.0269375
R12734 VDD.n1858 VDD.n1855 0.0269375
R12735 VDD.n1855 VDD.n1852 0.0269375
R12736 VDD.n1852 VDD.n1849 0.0269375
R12737 VDD.n1849 VDD.n1846 0.0269375
R12738 VDD.n1846 VDD.n1843 0.0269375
R12739 VDD.n1843 VDD.n1840 0.0269375
R12740 VDD.n1840 VDD.n1837 0.0269375
R12741 VDD.n1837 VDD.n1834 0.0269375
R12742 VDD.n1834 VDD.n1831 0.0269375
R12743 VDD.n1831 VDD.n1828 0.0269375
R12744 VDD.n1828 VDD.n1825 0.0269375
R12745 VDD.n1825 VDD.n1822 0.0269375
R12746 VDD.n1822 VDD.n1819 0.0269375
R12747 VDD.n1819 VDD.n1816 0.0269375
R12748 VDD.n1816 VDD.n1814 0.0269375
R12749 VDD.n1814 VDD.n1812 0.0269375
R12750 VDD.n1812 VDD.n1810 0.0269375
R12751 VDD.n1810 VDD.n1807 0.0269375
R12752 VDD.n1807 VDD.n1805 0.0269375
R12753 VDD.n1797 VDD.n1795 0.0269375
R12754 VDD.n1795 VDD.n1792 0.0269375
R12755 VDD.n1792 VDD.n1789 0.0269375
R12756 VDD.n1789 VDD.n1786 0.0269375
R12757 VDD.n1786 VDD.n1783 0.0269375
R12758 VDD.n1783 VDD.n1780 0.0269375
R12759 VDD.n1780 VDD.n1777 0.0269375
R12760 VDD.n1777 VDD.n1774 0.0269375
R12761 VDD.n1774 VDD.n1771 0.0269375
R12762 VDD.n1771 VDD.n1768 0.0269375
R12763 VDD.n1768 VDD.n1765 0.0269375
R12764 VDD.n1765 VDD.n1762 0.0269375
R12765 VDD.n1762 VDD.n1759 0.0269375
R12766 VDD.n1759 VDD.n1756 0.0269375
R12767 VDD.n1756 VDD.n1753 0.0269375
R12768 VDD.n1753 VDD.n1750 0.0269375
R12769 VDD.n1750 VDD.n1747 0.0269375
R12770 VDD.n1747 VDD.n1744 0.0269375
R12771 VDD.n1744 VDD.n1741 0.0269375
R12772 VDD.n1741 VDD.n1738 0.0269375
R12773 VDD.n1738 VDD.n1735 0.0269375
R12774 VDD.n1735 VDD.n1732 0.0269375
R12775 VDD.n1732 VDD.n1729 0.0269375
R12776 VDD.n1729 VDD.n1726 0.0269375
R12777 VDD.n1726 VDD.n1723 0.0269375
R12778 VDD.n1723 VDD.n1720 0.0269375
R12779 VDD.n1720 VDD.n1717 0.0269375
R12780 VDD.n1717 VDD.n1714 0.0269375
R12781 VDD.n1714 VDD.n1711 0.0269375
R12782 VDD.n1711 VDD.n1708 0.0269375
R12783 VDD.n1708 VDD.n1705 0.0269375
R12784 VDD.n1705 VDD.n1702 0.0269375
R12785 VDD.n1702 VDD.n1699 0.0269375
R12786 VDD.n1699 VDD.n1696 0.0269375
R12787 VDD.n1696 VDD.n1693 0.0269375
R12788 VDD.n1693 VDD.n1690 0.0269375
R12789 VDD.n1690 VDD.n1687 0.0269375
R12790 VDD.n1687 VDD.n1684 0.0269375
R12791 VDD.n1684 VDD.n1681 0.0269375
R12792 VDD.n1681 VDD.n1678 0.0269375
R12793 VDD.n1678 VDD.n1676 0.0269375
R12794 VDD.n1676 VDD.n1674 0.0269375
R12795 VDD.n1674 VDD.n1672 0.0269375
R12796 VDD.n1672 VDD.n1669 0.0269375
R12797 VDD.n1669 VDD.n1667 0.0269375
R12798 VDD.n1351 VDD.n1350 0.0269375
R12799 VDD.n1350 VDD.n1347 0.0269375
R12800 VDD.n1347 VDD.n1345 0.0269375
R12801 VDD.n1345 VDD.n1342 0.0269375
R12802 VDD.n1342 VDD.n1340 0.0269375
R12803 VDD.n1340 VDD.n1337 0.0269375
R12804 VDD.n1337 VDD.n1335 0.0269375
R12805 VDD.n1335 VDD.n1332 0.0269375
R12806 VDD.n1332 VDD.n1330 0.0269375
R12807 VDD.n1330 VDD.n1327 0.0269375
R12808 VDD.n1327 VDD.n1325 0.0269375
R12809 VDD.n1325 VDD.n1322 0.0269375
R12810 VDD.n1322 VDD.n1320 0.0269375
R12811 VDD.n1320 VDD.n1317 0.0269375
R12812 VDD.n1317 VDD.n1315 0.0269375
R12813 VDD.n1315 VDD.n1312 0.0269375
R12814 VDD.n1312 VDD.n1310 0.0269375
R12815 VDD.n1310 VDD.n1307 0.0269375
R12816 VDD.n1307 VDD.n1305 0.0269375
R12817 VDD.n1305 VDD.n1302 0.0269375
R12818 VDD.n1302 VDD.n1300 0.0269375
R12819 VDD.n1300 VDD.n1298 0.0269375
R12820 VDD.n1298 VDD.n1296 0.0269375
R12821 VDD.n1296 VDD.n1294 0.0269375
R12822 VDD.n1294 VDD.n1292 0.0269375
R12823 VDD.n1292 VDD.n1290 0.0269375
R12824 VDD.n1290 VDD.n1288 0.0269375
R12825 VDD.n1288 VDD.n1286 0.0269375
R12826 VDD.n1286 VDD.n1284 0.0269375
R12827 VDD.n1284 VDD.n1282 0.0269375
R12828 VDD.n1282 VDD.n1280 0.0269375
R12829 VDD.n1280 VDD.n1278 0.0269375
R12830 VDD.n1278 VDD.n1276 0.0269375
R12831 VDD.n1276 VDD.n1274 0.0269375
R12832 VDD.n1274 VDD.n1272 0.0269375
R12833 VDD.n1272 VDD.n1270 0.0269375
R12834 VDD.n1270 VDD.n1268 0.0269375
R12835 VDD.n1268 VDD.n1266 0.0269375
R12836 VDD.n1266 VDD.n1264 0.0269375
R12837 VDD.n1264 VDD.n1262 0.0269375
R12838 VDD.n1262 VDD.n1260 0.0269375
R12839 VDD.n1260 VDD.n1258 0.0269375
R12840 VDD.n1258 VDD.n1256 0.0269375
R12841 VDD.n1256 VDD.n1254 0.0269375
R12842 VDD.n1254 VDD.n1252 0.0269375
R12843 VDD.n1472 VDD.n1470 0.0269375
R12844 VDD.n1474 VDD.n1472 0.0269375
R12845 VDD.n1476 VDD.n1474 0.0269375
R12846 VDD.n1478 VDD.n1476 0.0269375
R12847 VDD.n1480 VDD.n1478 0.0269375
R12848 VDD.n1485 VDD.n1483 0.0269375
R12849 VDD.n1487 VDD.n1485 0.0269375
R12850 VDD.n1489 VDD.n1487 0.0269375
R12851 VDD.n1491 VDD.n1489 0.0269375
R12852 VDD.n1493 VDD.n1491 0.0269375
R12853 VDD.n1495 VDD.n1493 0.0269375
R12854 VDD.n1497 VDD.n1495 0.0269375
R12855 VDD.n1499 VDD.n1497 0.0269375
R12856 VDD.n1501 VDD.n1499 0.0269375
R12857 VDD.n1503 VDD.n1501 0.0269375
R12858 VDD.n1505 VDD.n1503 0.0269375
R12859 VDD.n1507 VDD.n1505 0.0269375
R12860 VDD.n1509 VDD.n1507 0.0269375
R12861 VDD.n1511 VDD.n1509 0.0269375
R12862 VDD.n1513 VDD.n1511 0.0269375
R12863 VDD.n1515 VDD.n1513 0.0269375
R12864 VDD.n1517 VDD.n1515 0.0269375
R12865 VDD.n1519 VDD.n1517 0.0269375
R12866 VDD.n1524 VDD.n1522 0.0269375
R12867 VDD.n1526 VDD.n1524 0.0269375
R12868 VDD.n1528 VDD.n1526 0.0269375
R12869 VDD.n1530 VDD.n1528 0.0269375
R12870 VDD.n1532 VDD.n1530 0.0269375
R12871 VDD.n1536 VDD.n1532 0.0269375
R12872 VDD.n1541 VDD.n1539 0.0269375
R12873 VDD.n1543 VDD.n1541 0.0269375
R12874 VDD.n1545 VDD.n1543 0.0269375
R12875 VDD.n1547 VDD.n1545 0.0269375
R12876 VDD.n1549 VDD.n1547 0.0269375
R12877 VDD.n1551 VDD.n1549 0.0269375
R12878 VDD.n1557 VDD.n1555 0.0269375
R12879 VDD.n1559 VDD.n1557 0.0269375
R12880 VDD.n1561 VDD.n1559 0.0269375
R12881 VDD.n1563 VDD.n1561 0.0269375
R12882 VDD.n1565 VDD.n1563 0.0269375
R12883 VDD.n1567 VDD.n1565 0.0269375
R12884 VDD.n1569 VDD.n1567 0.0269375
R12885 VDD.n1571 VDD.n1569 0.0269375
R12886 VDD.n1573 VDD.n1571 0.0269375
R12887 VDD.n1575 VDD.n1573 0.0269375
R12888 VDD.n1577 VDD.n1575 0.0269375
R12889 VDD.n1579 VDD.n1577 0.0269375
R12890 VDD.n1581 VDD.n1579 0.0269375
R12891 VDD.n1583 VDD.n1581 0.0269375
R12892 VDD.n1585 VDD.n1583 0.0269375
R12893 VDD.n1587 VDD.n1585 0.0269375
R12894 VDD.n1589 VDD.n1587 0.0269375
R12895 VDD.n1591 VDD.n1589 0.0269375
R12896 VDD.n1593 VDD.n1591 0.0269375
R12897 VDD.n1595 VDD.n1593 0.0269375
R12898 VDD.n1597 VDD.n1595 0.0269375
R12899 VDD.n1599 VDD.n1597 0.0269375
R12900 VDD.n1601 VDD.n1599 0.0269375
R12901 VDD.n1603 VDD.n1601 0.0269375
R12902 VDD.n1605 VDD.n1603 0.0269375
R12903 VDD.n1607 VDD.n1605 0.0269375
R12904 VDD.n1609 VDD.n1607 0.0269375
R12905 VDD.n1611 VDD.n1609 0.0269375
R12906 VDD.n1613 VDD.n1611 0.0269375
R12907 VDD.n1615 VDD.n1613 0.0269375
R12908 VDD.n1617 VDD.n1615 0.0269375
R12909 VDD.n1619 VDD.n1617 0.0269375
R12910 VDD.n1621 VDD.n1619 0.0269375
R12911 VDD.n1623 VDD.n1621 0.0269375
R12912 VDD.n1625 VDD.n1623 0.0269375
R12913 VDD.n1627 VDD.n1625 0.0269375
R12914 VDD.n1629 VDD.n1627 0.0269375
R12915 VDD.n1631 VDD.n1629 0.0269375
R12916 VDD.n1633 VDD.n1631 0.0269375
R12917 VDD.n1635 VDD.n1633 0.0269375
R12918 VDD.n1637 VDD.n1635 0.0269375
R12919 VDD.n1639 VDD.n1637 0.0269375
R12920 VDD.n1641 VDD.n1639 0.0269375
R12921 VDD.n1643 VDD.n1641 0.0269375
R12922 VDD.n1645 VDD.n1643 0.0269375
R12923 VDD.n1650 VDD.n1648 0.0269375
R12924 VDD.n1652 VDD.n1650 0.0269375
R12925 VDD.n1654 VDD.n1652 0.0269375
R12926 VDD.n1656 VDD.n1654 0.0269375
R12927 VDD.n1658 VDD.n1656 0.0269375
R12928 VDD.n1660 VDD.n1658 0.0269375
R12929 VDD.n1664 VDD.n1660 0.0269375
R12930 VDD.n1143 VDD.n1141 0.0269375
R12931 VDD.n1145 VDD.n1143 0.0269375
R12932 VDD.n1147 VDD.n1145 0.0269375
R12933 VDD.n1149 VDD.n1147 0.0269375
R12934 VDD.n1151 VDD.n1149 0.0269375
R12935 VDD.n1159 VDD.n1157 0.0269375
R12936 VDD.n1164 VDD.n1162 0.0269375
R12937 VDD.n1166 VDD.n1164 0.0269375
R12938 VDD.n1168 VDD.n1166 0.0269375
R12939 VDD.n1170 VDD.n1168 0.0269375
R12940 VDD.n1172 VDD.n1170 0.0269375
R12941 VDD.n1177 VDD.n1175 0.0269375
R12942 VDD.n1179 VDD.n1177 0.0269375
R12943 VDD.n1181 VDD.n1179 0.0269375
R12944 VDD.n1186 VDD.n1184 0.0269375
R12945 VDD.n1188 VDD.n1186 0.0269375
R12946 VDD.n1190 VDD.n1188 0.0269375
R12947 VDD.n1192 VDD.n1190 0.0269375
R12948 VDD.n1194 VDD.n1192 0.0269375
R12949 VDD.n1196 VDD.n1194 0.0269375
R12950 VDD.n1198 VDD.n1196 0.0269375
R12951 VDD.n1200 VDD.n1198 0.0269375
R12952 VDD.n1202 VDD.n1200 0.0269375
R12953 VDD.n1204 VDD.n1202 0.0269375
R12954 VDD.n1206 VDD.n1204 0.0269375
R12955 VDD.n1208 VDD.n1206 0.0269375
R12956 VDD.n1210 VDD.n1208 0.0269375
R12957 VDD.n1212 VDD.n1210 0.0269375
R12958 VDD.n1214 VDD.n1212 0.0269375
R12959 VDD.n1216 VDD.n1214 0.0269375
R12960 VDD.n1218 VDD.n1216 0.0269375
R12961 VDD.n1220 VDD.n1218 0.0269375
R12962 VDD.n1222 VDD.n1220 0.0269375
R12963 VDD.n1224 VDD.n1222 0.0269375
R12964 VDD.n1226 VDD.n1224 0.0269375
R12965 VDD.n1228 VDD.n1226 0.0269375
R12966 VDD.n1230 VDD.n1228 0.0269375
R12967 VDD.n1238 VDD.n1236 0.0269375
R12968 VDD.n1240 VDD.n1238 0.0269375
R12969 VDD.n1242 VDD.n1240 0.0269375
R12970 VDD.n1244 VDD.n1242 0.0269375
R12971 VDD.n1246 VDD.n1244 0.0269375
R12972 VDD.n2062 VDD.n2059 0.0269375
R12973 VDD.n2065 VDD.n2062 0.0269375
R12974 VDD.n2068 VDD.n2065 0.0269375
R12975 VDD.n2071 VDD.n2068 0.0269375
R12976 VDD.n2074 VDD.n2071 0.0269375
R12977 VDD.n2081 VDD.n2078 0.0269375
R12978 VDD.n2084 VDD.n2081 0.0269375
R12979 VDD.n2087 VDD.n2084 0.0269375
R12980 VDD.n2090 VDD.n2087 0.0269375
R12981 VDD.n2093 VDD.n2090 0.0269375
R12982 VDD.n2096 VDD.n2093 0.0269375
R12983 VDD.n2099 VDD.n2096 0.0269375
R12984 VDD.n2102 VDD.n2099 0.0269375
R12985 VDD.n2105 VDD.n2102 0.0269375
R12986 VDD.n2108 VDD.n2105 0.0269375
R12987 VDD.n2111 VDD.n2108 0.0269375
R12988 VDD.n2114 VDD.n2111 0.0269375
R12989 VDD.n2117 VDD.n2114 0.0269375
R12990 VDD.n2120 VDD.n2117 0.0269375
R12991 VDD.n2123 VDD.n2120 0.0269375
R12992 VDD.n2126 VDD.n2123 0.0269375
R12993 VDD.n2129 VDD.n2126 0.0269375
R12994 VDD.n2132 VDD.n2129 0.0269375
R12995 VDD.n2139 VDD.n2136 0.0269375
R12996 VDD.n2142 VDD.n2139 0.0269375
R12997 VDD.n2145 VDD.n2142 0.0269375
R12998 VDD.n2148 VDD.n2145 0.0269375
R12999 VDD.n2151 VDD.n2148 0.0269375
R13000 VDD.n2159 VDD.n2151 0.0269375
R13001 VDD.n2166 VDD.n2163 0.0269375
R13002 VDD.n2169 VDD.n2166 0.0269375
R13003 VDD.n2172 VDD.n2169 0.0269375
R13004 VDD.n2175 VDD.n2172 0.0269375
R13005 VDD.n2178 VDD.n2175 0.0269375
R13006 VDD.n2181 VDD.n2178 0.0269375
R13007 VDD.n2188 VDD.n2185 0.0269375
R13008 VDD.n2191 VDD.n2188 0.0269375
R13009 VDD.n2194 VDD.n2191 0.0269375
R13010 VDD.n2197 VDD.n2194 0.0269375
R13011 VDD.n2200 VDD.n2197 0.0269375
R13012 VDD.n2203 VDD.n2200 0.0269375
R13013 VDD.n2206 VDD.n2203 0.0269375
R13014 VDD.n2209 VDD.n2206 0.0269375
R13015 VDD.n2212 VDD.n2209 0.0269375
R13016 VDD.n2215 VDD.n2212 0.0269375
R13017 VDD.n2218 VDD.n2215 0.0269375
R13018 VDD.n2221 VDD.n2218 0.0269375
R13019 VDD.n2224 VDD.n2221 0.0269375
R13020 VDD.n2227 VDD.n2224 0.0269375
R13021 VDD.n2230 VDD.n2227 0.0269375
R13022 VDD.n2233 VDD.n2230 0.0269375
R13023 VDD.n2236 VDD.n2233 0.0269375
R13024 VDD.n2239 VDD.n2236 0.0269375
R13025 VDD.n2242 VDD.n2239 0.0269375
R13026 VDD.n2245 VDD.n2242 0.0269375
R13027 VDD.n2248 VDD.n2245 0.0269375
R13028 VDD.n2251 VDD.n2248 0.0269375
R13029 VDD.n2254 VDD.n2251 0.0269375
R13030 VDD.n2257 VDD.n2254 0.0269375
R13031 VDD.n2260 VDD.n2257 0.0269375
R13032 VDD.n2263 VDD.n2260 0.0269375
R13033 VDD.n2266 VDD.n2263 0.0269375
R13034 VDD.n2269 VDD.n2266 0.0269375
R13035 VDD.n2272 VDD.n2269 0.0269375
R13036 VDD.n2275 VDD.n2272 0.0269375
R13037 VDD.n2278 VDD.n2275 0.0269375
R13038 VDD.n2281 VDD.n2278 0.0269375
R13039 VDD.n2284 VDD.n2281 0.0269375
R13040 VDD.n2287 VDD.n2284 0.0269375
R13041 VDD.n2290 VDD.n2287 0.0269375
R13042 VDD.n2293 VDD.n2290 0.0269375
R13043 VDD.n2296 VDD.n2293 0.0269375
R13044 VDD.n2299 VDD.n2296 0.0269375
R13045 VDD.n2302 VDD.n2299 0.0269375
R13046 VDD.n2305 VDD.n2302 0.0269375
R13047 VDD.n2308 VDD.n2305 0.0269375
R13048 VDD.n2311 VDD.n2308 0.0269375
R13049 VDD.n2314 VDD.n2311 0.0269375
R13050 VDD.n2317 VDD.n2314 0.0269375
R13051 VDD.n2320 VDD.n2317 0.0269375
R13052 VDD.n2327 VDD.n2324 0.0269375
R13053 VDD.n2330 VDD.n2327 0.0269375
R13054 VDD.n2333 VDD.n2330 0.0269375
R13055 VDD.n2336 VDD.n2333 0.0269375
R13056 VDD.n2339 VDD.n2336 0.0269375
R13057 VDD.n2342 VDD.n2339 0.0269375
R13058 VDD.n2350 VDD.n2342 0.0269375
R13059 VDD.n2357 VDD.n2354 0.0269375
R13060 VDD.n2360 VDD.n2357 0.0269375
R13061 VDD.n2363 VDD.n2360 0.0269375
R13062 VDD.n2366 VDD.n2363 0.0269375
R13063 VDD.n2369 VDD.n2366 0.0269375
R13064 VDD.n2388 VDD.n2385 0.0269375
R13065 VDD.n2403 VDD.n2400 0.0269375
R13066 VDD.n2410 VDD.n2407 0.0269375
R13067 VDD.n2413 VDD.n2410 0.0269375
R13068 VDD.n2416 VDD.n2413 0.0269375
R13069 VDD.n2424 VDD.n2421 0.0269375
R13070 VDD.n2427 VDD.n2424 0.0269375
R13071 VDD.n2434 VDD.n2431 0.0269375
R13072 VDD.n2441 VDD.n2438 0.0269375
R13073 VDD.n2448 VDD.n2445 0.0269375
R13074 VDD.n2451 VDD.n2448 0.0269375
R13075 VDD.n2459 VDD.n2456 0.0269375
R13076 VDD.n2462 VDD.n2459 0.0269375
R13077 VDD.n2469 VDD.n2466 0.0269375
R13078 VDD.n2476 VDD.n2473 0.0269375
R13079 VDD.n2483 VDD.n2480 0.0269375
R13080 VDD.n2486 VDD.n2483 0.0269375
R13081 VDD.n2497 VDD.n2494 0.0269375
R13082 VDD.n2500 VDD.n2497 0.0269375
R13083 VDD.n2515 VDD.n2512 0.0269375
R13084 VDD.n2518 VDD.n2515 0.0269375
R13085 VDD.n2521 VDD.n2518 0.0269375
R13086 VDD.n2524 VDD.n2521 0.0269375
R13087 VDD.n2445 VDD.n2442 0.0266563
R13088 VDD.n3762 VDD.n3760 0.026375
R13089 VDD.n3825 VDD.n3824 0.026375
R13090 VDD.n3869 VDD.n3867 0.026375
R13091 VDD.n3932 VDD.n3931 0.026375
R13092 VDD.n6192 VDD.n6189 0.026375
R13093 VDD.n6285 VDD.n6284 0.026375
R13094 VDD.n6347 VDD.n6344 0.026375
R13095 VDD.n6440 VDD.n6439 0.026375
R13096 VDD.n3556 VDD.n3554 0.026375
R13097 VDD.n3619 VDD.n3618 0.026375
R13098 VDD.n3664 VDD.n3662 0.026375
R13099 VDD.n3727 VDD.n3726 0.026375
R13100 VDD.n5890 VDD.n5887 0.026375
R13101 VDD.n5983 VDD.n5982 0.026375
R13102 VDD.n6045 VDD.n6042 0.026375
R13103 VDD.n6138 VDD.n6137 0.026375
R13104 VDD.n5574 VDD.n5571 0.026375
R13105 VDD.n5667 VDD.n5666 0.026375
R13106 VDD.n5743 VDD.n5740 0.026375
R13107 VDD.n5836 VDD.n5835 0.026375
R13108 VDD.n3357 VDD.n3355 0.026375
R13109 VDD.n3420 VDD.n3419 0.026375
R13110 VDD.n3463 VDD.n3461 0.026375
R13111 VDD.n3526 VDD.n3525 0.026375
R13112 VDD.n2606 VDD.n2604 0.026375
R13113 VDD.n2669 VDD.n2668 0.026375
R13114 VDD.n6506 VDD.n6503 0.026375
R13115 VDD.n6599 VDD.n6598 0.026375
R13116 VDD.n1104 VDD.n1103 0.026375
R13117 VDD.n1155 VDD.n1154 0.0260938
R13118 VDD.n1233 VDD.n1231 0.0260938
R13119 VDD.n2374 VDD.n2373 0.0260938
R13120 VDD.n2392 VDD.n2389 0.0260938
R13121 VDD.n2470 VDD.n2469 0.0260938
R13122 VDD.n2504 VDD.n2501 0.0260938
R13123 VDD.n386 VDD.n385 0.0258125
R13124 VDD.n5864 VDD.n5863 0.0258125
R13125 VDD.n5710 VDD.n5709 0.0258125
R13126 VDD.n1470 VDD.n1468 0.0249687
R13127 VDD.n1539 VDD.n1537 0.0249687
R13128 VDD.n1250 VDD.n1246 0.0249687
R13129 VDD.n2059 VDD.n2056 0.0249687
R13130 VDD.n2163 VDD.n2160 0.0249687
R13131 VDD.n2354 VDD.n2351 0.0249687
R13132 VDD.n2541 VDD.n2524 0.0249687
R13133 VDD.n441 VDD.n440 0.0246875
R13134 VDD.n7410 VDD.n7408 0.0246875
R13135 VDD.n350 VDD.n349 0.0246875
R13136 VDD.n7532 VDD.n7529 0.0246875
R13137 VDD.n3769 VDD.n3767 0.0246875
R13138 VDD.n3818 VDD.n3817 0.0246875
R13139 VDD.n3876 VDD.n3874 0.0246875
R13140 VDD.n3925 VDD.n3924 0.0246875
R13141 VDD.n6202 VDD.n6199 0.0246875
R13142 VDD.n6275 VDD.n6274 0.0246875
R13143 VDD.n6357 VDD.n6354 0.0246875
R13144 VDD.n6430 VDD.n6429 0.0246875
R13145 VDD.n3563 VDD.n3561 0.0246875
R13146 VDD.n3612 VDD.n3611 0.0246875
R13147 VDD.n3671 VDD.n3669 0.0246875
R13148 VDD.n3720 VDD.n3719 0.0246875
R13149 VDD.n5900 VDD.n5897 0.0246875
R13150 VDD.n5973 VDD.n5972 0.0246875
R13151 VDD.n6055 VDD.n6052 0.0246875
R13152 VDD.n6128 VDD.n6127 0.0246875
R13153 VDD.n5584 VDD.n5581 0.0246875
R13154 VDD.n5657 VDD.n5656 0.0246875
R13155 VDD.n5753 VDD.n5750 0.0246875
R13156 VDD.n5826 VDD.n5825 0.0246875
R13157 VDD.n3364 VDD.n3362 0.0246875
R13158 VDD.n3413 VDD.n3412 0.0246875
R13159 VDD.n3470 VDD.n3468 0.0246875
R13160 VDD.n3519 VDD.n3518 0.0246875
R13161 VDD.n2613 VDD.n2611 0.0246875
R13162 VDD.n2662 VDD.n2661 0.0246875
R13163 VDD.n6516 VDD.n6513 0.0246875
R13164 VDD.n6589 VDD.n6588 0.0246875
R13165 VDD.n7551 VDD.n7550 0.0246875
R13166 VDD.n4457 VDD.n4455 0.024264
R13167 VDD.n4460 VDD.n4457 0.024264
R13168 VDD.n4462 VDD.n4460 0.024264
R13169 VDD.n4465 VDD.n4462 0.024264
R13170 VDD.n4467 VDD.n4465 0.024264
R13171 VDD.n4470 VDD.n4467 0.024264
R13172 VDD.n4472 VDD.n4470 0.024264
R13173 VDD.n4475 VDD.n4472 0.024264
R13174 VDD.n4477 VDD.n4475 0.024264
R13175 VDD.n4480 VDD.n4477 0.024264
R13176 VDD.n4482 VDD.n4480 0.024264
R13177 VDD.n4485 VDD.n4482 0.024264
R13178 VDD.n4487 VDD.n4485 0.024264
R13179 VDD.n4490 VDD.n4487 0.024264
R13180 VDD.n4492 VDD.n4490 0.024264
R13181 VDD.n4495 VDD.n4492 0.024264
R13182 VDD.n4497 VDD.n4495 0.024264
R13183 VDD.n4500 VDD.n4497 0.024264
R13184 VDD.n4502 VDD.n4500 0.024264
R13185 VDD.n4505 VDD.n4502 0.024264
R13186 VDD.n4507 VDD.n4505 0.024264
R13187 VDD.n4510 VDD.n4507 0.024264
R13188 VDD.n4512 VDD.n4510 0.024264
R13189 VDD.n4515 VDD.n4512 0.024264
R13190 VDD.n4517 VDD.n4515 0.024264
R13191 VDD.n4520 VDD.n4517 0.024264
R13192 VDD.n4522 VDD.n4520 0.024264
R13193 VDD.n4525 VDD.n4522 0.024264
R13194 VDD.n4527 VDD.n4525 0.024264
R13195 VDD.n4530 VDD.n4527 0.024264
R13196 VDD.n4532 VDD.n4530 0.024264
R13197 VDD.n4535 VDD.n4532 0.024264
R13198 VDD.n4537 VDD.n4535 0.024264
R13199 VDD.n4540 VDD.n4537 0.024264
R13200 VDD.n4542 VDD.n4540 0.024264
R13201 VDD.n4545 VDD.n4542 0.024264
R13202 VDD.n4547 VDD.n4545 0.024264
R13203 VDD.n4550 VDD.n4547 0.024264
R13204 VDD.n4552 VDD.n4550 0.024264
R13205 VDD.n4555 VDD.n4552 0.024264
R13206 VDD.n4557 VDD.n4555 0.024264
R13207 VDD.n4560 VDD.n4557 0.024264
R13208 VDD.n4562 VDD.n4560 0.024264
R13209 VDD.n4565 VDD.n4562 0.024264
R13210 VDD.n4567 VDD.n4565 0.024264
R13211 VDD.n4570 VDD.n4567 0.024264
R13212 VDD.n4572 VDD.n4570 0.024264
R13213 VDD.n4575 VDD.n4572 0.024264
R13214 VDD.n3959 VDD.n3957 0.024264
R13215 VDD.n3961 VDD.n3959 0.024264
R13216 VDD.n3963 VDD.n3961 0.024264
R13217 VDD.n3965 VDD.n3963 0.024264
R13218 VDD.n3967 VDD.n3965 0.024264
R13219 VDD.n3969 VDD.n3967 0.024264
R13220 VDD.n3971 VDD.n3969 0.024264
R13221 VDD.n3973 VDD.n3971 0.024264
R13222 VDD.n3975 VDD.n3973 0.024264
R13223 VDD.n3977 VDD.n3975 0.024264
R13224 VDD.n3979 VDD.n3977 0.024264
R13225 VDD.n3981 VDD.n3979 0.024264
R13226 VDD.n3983 VDD.n3981 0.024264
R13227 VDD.n3985 VDD.n3983 0.024264
R13228 VDD.n3987 VDD.n3985 0.024264
R13229 VDD.n3989 VDD.n3987 0.024264
R13230 VDD.n3991 VDD.n3989 0.024264
R13231 VDD.n3993 VDD.n3991 0.024264
R13232 VDD.n3995 VDD.n3993 0.024264
R13233 VDD.n3997 VDD.n3995 0.024264
R13234 VDD.n3999 VDD.n3997 0.024264
R13235 VDD.n4001 VDD.n3999 0.024264
R13236 VDD.n4003 VDD.n4001 0.024264
R13237 VDD.n4005 VDD.n4003 0.024264
R13238 VDD.n4007 VDD.n4005 0.024264
R13239 VDD.n4009 VDD.n4007 0.024264
R13240 VDD.n4011 VDD.n4009 0.024264
R13241 VDD.n4013 VDD.n4011 0.024264
R13242 VDD.n4015 VDD.n4013 0.024264
R13243 VDD.n4018 VDD.n4015 0.024264
R13244 VDD.n4020 VDD.n4018 0.024264
R13245 VDD.n4023 VDD.n4020 0.024264
R13246 VDD.n4025 VDD.n4023 0.024264
R13247 VDD.n4028 VDD.n4025 0.024264
R13248 VDD.n4030 VDD.n4028 0.024264
R13249 VDD.n4033 VDD.n4030 0.024264
R13250 VDD.n4035 VDD.n4033 0.024264
R13251 VDD.n4038 VDD.n4035 0.024264
R13252 VDD.n4040 VDD.n4038 0.024264
R13253 VDD.n4043 VDD.n4040 0.024264
R13254 VDD.n4045 VDD.n4043 0.024264
R13255 VDD.n4048 VDD.n4045 0.024264
R13256 VDD.n4050 VDD.n4048 0.024264
R13257 VDD.n4053 VDD.n4050 0.024264
R13258 VDD.n4055 VDD.n4053 0.024264
R13259 VDD.n4058 VDD.n4055 0.024264
R13260 VDD.n4060 VDD.n4058 0.024264
R13261 VDD.n4063 VDD.n4060 0.024264
R13262 VDD.n4065 VDD.n4063 0.024264
R13263 VDD.n3181 VDD.n3179 0.024264
R13264 VDD.n4962 VDD.n4960 0.024264
R13265 VDD.n4965 VDD.n4962 0.024264
R13266 VDD.n4967 VDD.n4965 0.024264
R13267 VDD.n4970 VDD.n4967 0.024264
R13268 VDD.n4972 VDD.n4970 0.024264
R13269 VDD.n4975 VDD.n4972 0.024264
R13270 VDD.n4977 VDD.n4975 0.024264
R13271 VDD.n4980 VDD.n4977 0.024264
R13272 VDD.n4982 VDD.n4980 0.024264
R13273 VDD.n4985 VDD.n4982 0.024264
R13274 VDD.n4987 VDD.n4985 0.024264
R13275 VDD.n4990 VDD.n4987 0.024264
R13276 VDD.n4992 VDD.n4990 0.024264
R13277 VDD.n4995 VDD.n4992 0.024264
R13278 VDD.n4997 VDD.n4995 0.024264
R13279 VDD.n5000 VDD.n4997 0.024264
R13280 VDD.n5002 VDD.n5000 0.024264
R13281 VDD.n5005 VDD.n5002 0.024264
R13282 VDD.n5007 VDD.n5005 0.024264
R13283 VDD.n5010 VDD.n5007 0.024264
R13284 VDD.n5012 VDD.n5010 0.024264
R13285 VDD.n5015 VDD.n5012 0.024264
R13286 VDD.n5017 VDD.n5015 0.024264
R13287 VDD.n5020 VDD.n5017 0.024264
R13288 VDD.n5022 VDD.n5020 0.024264
R13289 VDD.n5025 VDD.n5022 0.024264
R13290 VDD.n5027 VDD.n5025 0.024264
R13291 VDD.n5030 VDD.n5027 0.024264
R13292 VDD.n5032 VDD.n5030 0.024264
R13293 VDD.n5035 VDD.n5032 0.024264
R13294 VDD.n5037 VDD.n5035 0.024264
R13295 VDD.n5040 VDD.n5037 0.024264
R13296 VDD.n5042 VDD.n5040 0.024264
R13297 VDD.n5045 VDD.n5042 0.024264
R13298 VDD.n5047 VDD.n5045 0.024264
R13299 VDD.n5050 VDD.n5047 0.024264
R13300 VDD.n5052 VDD.n5050 0.024264
R13301 VDD.n5055 VDD.n5052 0.024264
R13302 VDD.n5057 VDD.n5055 0.024264
R13303 VDD.n5060 VDD.n5057 0.024264
R13304 VDD.n5062 VDD.n5060 0.024264
R13305 VDD.n5065 VDD.n5062 0.024264
R13306 VDD.n5067 VDD.n5065 0.024264
R13307 VDD.n5070 VDD.n5067 0.024264
R13308 VDD.n5072 VDD.n5070 0.024264
R13309 VDD.n5075 VDD.n5072 0.024264
R13310 VDD.n3781 VDD.n3780 0.024125
R13311 VDD.n3806 VDD.n3804 0.024125
R13312 VDD.n3888 VDD.n3887 0.024125
R13313 VDD.n3913 VDD.n3911 0.024125
R13314 VDD.n6219 VDD.n6218 0.024125
R13315 VDD.n6258 VDD.n6255 0.024125
R13316 VDD.n6374 VDD.n6373 0.024125
R13317 VDD.n6413 VDD.n6410 0.024125
R13318 VDD.n3575 VDD.n3574 0.024125
R13319 VDD.n3600 VDD.n3598 0.024125
R13320 VDD.n3683 VDD.n3682 0.024125
R13321 VDD.n3708 VDD.n3706 0.024125
R13322 VDD.n5917 VDD.n5916 0.024125
R13323 VDD.n5956 VDD.n5953 0.024125
R13324 VDD.n6072 VDD.n6071 0.024125
R13325 VDD.n6111 VDD.n6108 0.024125
R13326 VDD.n5601 VDD.n5600 0.024125
R13327 VDD.n5640 VDD.n5637 0.024125
R13328 VDD.n5770 VDD.n5769 0.024125
R13329 VDD.n5809 VDD.n5806 0.024125
R13330 VDD.n3376 VDD.n3375 0.024125
R13331 VDD.n3401 VDD.n3399 0.024125
R13332 VDD.n3482 VDD.n3481 0.024125
R13333 VDD.n3507 VDD.n3505 0.024125
R13334 VDD.n2625 VDD.n2624 0.024125
R13335 VDD.n2650 VDD.n2648 0.024125
R13336 VDD.n6533 VDD.n6532 0.024125
R13337 VDD.n6572 VDD.n6569 0.024125
R13338 VDD.n1481 VDD.n1480 0.0227188
R13339 VDD.n1648 VDD.n1646 0.0227188
R13340 VDD.n2075 VDD.n2074 0.0227188
R13341 VDD.n2324 VDD.n2321 0.0227188
R13342 VDD.n2463 VDD.n2462 0.0221563
R13343 VDD.n3841 VDD.n3840 0.021875
R13344 VDD.n3853 VDD.n3851 0.021875
R13345 VDD.n6308 VDD.n6307 0.021875
R13346 VDD.n3648 VDD.n3646 0.021875
R13347 VDD.n6006 VDD.n6005 0.021875
R13348 VDD.n5548 VDD.n5545 0.021875
R13349 VDD.n5690 VDD.n5689 0.021875
R13350 VDD.n5719 VDD.n5716 0.021875
R13351 VDD.n3341 VDD.n3339 0.021875
R13352 VDD.n3436 VDD.n3435 0.021875
R13353 VDD.n3447 VDD.n3445 0.021875
R13354 VDD.n2693 VDD.n2689 0.021875
R13355 VDD.n6627 VDD.n6621 0.021875
R13356 VDD.n1173 VDD.n1172 0.0215938
R13357 VDD.n1184 VDD.n1182 0.0215938
R13358 VDD.n2404 VDD.n2403 0.0215938
R13359 VDD.n2421 VDD.n2418 0.0215938
R13360 VDD.n7354 VDD.n7353 0.0213125
R13361 VDD.n6670 VDD.n6668 0.0213125
R13362 VDD.n818 VDD.n816 0.0213125
R13363 VDD.n583 VDD.n581 0.0213125
R13364 VDD.n627 VDD.n625 0.0213125
R13365 VDD.n6852 VDD.n6849 0.0213125
R13366 VDD.n1009 VDD.n1006 0.0213125
R13367 VDD.n1043 VDD.n1040 0.0213125
R13368 VDD.n560 VDD.n559 0.0213125
R13369 VDD.n2480 VDD.n2477 0.0210313
R13370 VDD.n6019 VDD.n6018 0.02075
R13371 VDD.n126 VDD.n123 0.0201875
R13372 VDD.n189 VDD.n188 0.0201875
R13373 VDD.n6680 VDD.n6679 0.0201875
R13374 VDD.n828 VDD.n827 0.0201875
R13375 VDD.n6866 VDD.n6865 0.0201875
R13376 VDD.n7010 VDD.n7007 0.0201875
R13377 VDD.n7073 VDD.n7072 0.0201875
R13378 VDD.n3957 VDD.n3955 0.0199663
R13379 VDD.n6483 VDD.n4065 0.0199663
R13380 VDD.n3540 VDD.n3181 0.0199663
R13381 VDD.n1154 VDD.n1152 0.0199062
R13382 VDD.n1234 VDD.n1233 0.0199062
R13383 VDD.n2373 VDD.n2370 0.0199062
R13384 VDD.n2505 VDD.n2504 0.0199062
R13385 VDD.n197 VDD.n195 0.0197857
R13386 VDD.n119 VDD.n105 0.0197857
R13387 VDD.n2494 VDD.n2491 0.0193437
R13388 VDD.n314 VDD.n313 0.0190625
R13389 VDD.n382 VDD.n379 0.0190625
R13390 VDD.n6235 VDD.n6232 0.0190625
R13391 VDD.n6242 VDD.n6241 0.0190625
R13392 VDD.n6390 VDD.n6387 0.0190625
R13393 VDD.n6397 VDD.n6396 0.0190625
R13394 VDD.n5933 VDD.n5930 0.0190625
R13395 VDD.n5940 VDD.n5939 0.0190625
R13396 VDD.n6088 VDD.n6085 0.0190625
R13397 VDD.n6095 VDD.n6094 0.0190625
R13398 VDD.n5617 VDD.n5614 0.0190625
R13399 VDD.n5624 VDD.n5623 0.0190625
R13400 VDD.n5786 VDD.n5783 0.0190625
R13401 VDD.n5793 VDD.n5792 0.0190625
R13402 VDD.n6549 VDD.n6546 0.0190625
R13403 VDD.n6556 VDD.n6555 0.0190625
R13404 VDD.n7575 VDD.n7573 0.0190625
R13405 VDD.n7704 VDD.n7703 0.0190625
R13406 VDD.n1522 VDD.n1520 0.0187812
R13407 VDD.n2136 VDD.n2133 0.0187812
R13408 VDD.n2397 VDD.n2396 0.0187812
R13409 VDD.n3757 VDD.n3755 0.0185
R13410 VDD.n3830 VDD.n3829 0.0185
R13411 VDD.n3864 VDD.n3862 0.0185
R13412 VDD.n3942 VDD.n3936 0.0185
R13413 VDD.n6185 VDD.n6182 0.0185
R13414 VDD.n6292 VDD.n6291 0.0185
R13415 VDD.n6340 VDD.n6337 0.0185
R13416 VDD.n6447 VDD.n6446 0.0185
R13417 VDD.n3551 VDD.n3549 0.0185
R13418 VDD.n3624 VDD.n3623 0.0185
R13419 VDD.n3659 VDD.n3657 0.0185
R13420 VDD.n3737 VDD.n3731 0.0185
R13421 VDD.n5883 VDD.n5880 0.0185
R13422 VDD.n5990 VDD.n5989 0.0185
R13423 VDD.n6038 VDD.n6035 0.0185
R13424 VDD.n6145 VDD.n6144 0.0185
R13425 VDD.n5567 VDD.n5564 0.0185
R13426 VDD.n5674 VDD.n5673 0.0185
R13427 VDD.n5736 VDD.n5733 0.0185
R13428 VDD.n5843 VDD.n5842 0.0185
R13429 VDD.n3352 VDD.n3350 0.0185
R13430 VDD.n3425 VDD.n3424 0.0185
R13431 VDD.n3458 VDD.n3456 0.0185
R13432 VDD.n3531 VDD.n3530 0.0185
R13433 VDD.n2601 VDD.n2599 0.0185
R13434 VDD.n2679 VDD.n2673 0.0185
R13435 VDD.n6499 VDD.n6496 0.0185
R13436 VDD.n6606 VDD.n6605 0.0185
R13437 VDD.n1162 VDD.n1160 0.0182187
R13438 VDD.n2385 VDD.n2382 0.0182187
R13439 VDD.n2438 VDD.n2435 0.0182187
R13440 VDD.n130 VDD.n129 0.0179375
R13441 VDD.n185 VDD.n182 0.0179375
R13442 VDD.n6677 VDD.n6675 0.0179375
R13443 VDD.n825 VDD.n823 0.0179375
R13444 VDD.n5723 VDD.n5720 0.0179375
R13445 VDD.n6862 VDD.n6859 0.0179375
R13446 VDD.n7014 VDD.n7013 0.0179375
R13447 VDD.n7069 VDD.n7066 0.0179375
R13448 VDD.n1553 VDD.n1551 0.0170938
R13449 VDD.n2182 VDD.n2181 0.0170938
R13450 VDD.n2381 VDD.n2378 0.0170938
R13451 VDD.n2487 VDD.n2486 0.0170938
R13452 VDD.n2396 VDD.n2393 0.0165313
R13453 VDD.n2428 VDD.n2427 0.0165313
R13454 VDD.n2509 VDD.n2508 0.0165313
R13455 VDD.n6166 VDD.n6165 0.0156875
R13456 VDD.n6012 VDD.n6011 0.0156875
R13457 VDD.n7059 VDD.n7058 0.015125
R13458 VDD.n7344 VDD.n7341 0.0145625
R13459 VDD.n7111 VDD.n7109 0.0145625
R13460 VDD.n7257 VDD.n7256 0.0145625
R13461 VDD.n3776 VDD.n3774 0.014
R13462 VDD.n3811 VDD.n3810 0.014
R13463 VDD.n3883 VDD.n3881 0.014
R13464 VDD.n3918 VDD.n3917 0.014
R13465 VDD.n6212 VDD.n6209 0.014
R13466 VDD.n6265 VDD.n6264 0.014
R13467 VDD.n6367 VDD.n6364 0.014
R13468 VDD.n6420 VDD.n6419 0.014
R13469 VDD.n3570 VDD.n3568 0.014
R13470 VDD.n3605 VDD.n3604 0.014
R13471 VDD.n3678 VDD.n3676 0.014
R13472 VDD.n3713 VDD.n3712 0.014
R13473 VDD.n5910 VDD.n5907 0.014
R13474 VDD.n5963 VDD.n5962 0.014
R13475 VDD.n6065 VDD.n6062 0.014
R13476 VDD.n6118 VDD.n6117 0.014
R13477 VDD.n5594 VDD.n5591 0.014
R13478 VDD.n5647 VDD.n5646 0.014
R13479 VDD.n5763 VDD.n5760 0.014
R13480 VDD.n5816 VDD.n5815 0.014
R13481 VDD.n3371 VDD.n3369 0.014
R13482 VDD.n3406 VDD.n3405 0.014
R13483 VDD.n3477 VDD.n3475 0.014
R13484 VDD.n3512 VDD.n3511 0.014
R13485 VDD.n2620 VDD.n2618 0.014
R13486 VDD.n2655 VDD.n2654 0.014
R13487 VDD.n6526 VDD.n6523 0.014
R13488 VDD.n6579 VDD.n6578 0.014
R13489 VDD.n778 VDD.n777 0.014
R13490 VDD.n7003 VDD.n7002 0.014
R13491 VDD.n328 VDD.n325 0.0134375
R13492 VDD.n3774 VDD.n3773 0.0134375
R13493 VDD.n3813 VDD.n3811 0.0134375
R13494 VDD.n3881 VDD.n3880 0.0134375
R13495 VDD.n3920 VDD.n3918 0.0134375
R13496 VDD.n6209 VDD.n6208 0.0134375
R13497 VDD.n6268 VDD.n6265 0.0134375
R13498 VDD.n6364 VDD.n6363 0.0134375
R13499 VDD.n6423 VDD.n6420 0.0134375
R13500 VDD.n3568 VDD.n3567 0.0134375
R13501 VDD.n3607 VDD.n3605 0.0134375
R13502 VDD.n3676 VDD.n3675 0.0134375
R13503 VDD.n3715 VDD.n3713 0.0134375
R13504 VDD.n5907 VDD.n5906 0.0134375
R13505 VDD.n5966 VDD.n5963 0.0134375
R13506 VDD.n6062 VDD.n6061 0.0134375
R13507 VDD.n6121 VDD.n6118 0.0134375
R13508 VDD.n5591 VDD.n5590 0.0134375
R13509 VDD.n5650 VDD.n5647 0.0134375
R13510 VDD.n5760 VDD.n5759 0.0134375
R13511 VDD.n5819 VDD.n5816 0.0134375
R13512 VDD.n3369 VDD.n3368 0.0134375
R13513 VDD.n3408 VDD.n3406 0.0134375
R13514 VDD.n3475 VDD.n3474 0.0134375
R13515 VDD.n3514 VDD.n3512 0.0134375
R13516 VDD.n2618 VDD.n2617 0.0134375
R13517 VDD.n2657 VDD.n2655 0.0134375
R13518 VDD.n6523 VDD.n6522 0.0134375
R13519 VDD.n6582 VDD.n6579 0.0134375
R13520 VDD.n7027 VDD.n7024 0.0134375
R13521 VDD.n7561 VDD.n7559 0.012875
R13522 VDD.n6804 VDD.n6785 0.0124871
R13523 VDD.n7237 VDD.n286 0.01175
R13524 VDD.n7684 VDD.n7670 0.01175
R13525 VDD.n7590 VDD.n7588 0.01175
R13526 VDD.n7237 VDD.n7223 0.01175
R13527 VDD.n7126 VDD.n7124 0.01175
R13528 VDD.n7002 VDD.n7000 0.01175
R13529 VDD.n638 VDD.n636 0.01175
R13530 VDD.n777 VDD.n775 0.01175
R13531 VDD.n836 VDD.n834 0.01175
R13532 VDD.n1029 VDD.n971 0.01175
R13533 VDD.n6687 VDD.n6685 0.01175
R13534 VDD.n6169 VDD.n6166 0.01175
R13535 VDD.n6324 VDD.n6321 0.01175
R13536 VDD.n3635 VDD.n3634 0.01175
R13537 VDD.n6873 VDD.n6804 0.01175
R13538 VDD.n2452 VDD.n2451 0.0114688
R13539 VDD.n6661 VDD.n6660 0.0111875
R13540 VDD.n809 VDD.n808 0.0111875
R13541 VDD.n6839 VDD.n6838 0.0111875
R13542 VDD.n996 VDD.n995 0.0111875
R13543 VDD.n2393 VDD.n2392 0.0109063
R13544 VDD.n2431 VDD.n2428 0.0109063
R13545 VDD.n2512 VDD.n2509 0.0109063
R13546 VDD.n6321 VDD.n6320 0.010625
R13547 VDD.n3636 VDD.n3635 0.010625
R13548 VDD.n1555 VDD.n1553 0.0103438
R13549 VDD.n2185 VDD.n2182 0.0103438
R13550 VDD.n2378 VDD.n2377 0.0103438
R13551 VDD.n2490 VDD.n2487 0.0103438
R13552 VDD.n2456 VDD.n2453 0.00978125
R13553 VDD.n5720 VDD.n5719 0.0095
R13554 VDD.n1160 VDD.n1159 0.00921875
R13555 VDD.n2382 VDD.n2381 0.00921875
R13556 VDD.n2435 VDD.n2434 0.00921875
R13557 VDD.n446 VDD.n445 0.0089375
R13558 VDD.n7415 VDD.n7414 0.0089375
R13559 VDD.n7525 VDD.n7522 0.0089375
R13560 VDD.n3755 VDD.n3754 0.0089375
R13561 VDD.n3832 VDD.n3830 0.0089375
R13562 VDD.n3862 VDD.n3861 0.0089375
R13563 VDD.n3944 VDD.n3942 0.0089375
R13564 VDD.n6182 VDD.n6181 0.0089375
R13565 VDD.n6295 VDD.n6292 0.0089375
R13566 VDD.n6337 VDD.n6336 0.0089375
R13567 VDD.n6450 VDD.n6447 0.0089375
R13568 VDD.n3549 VDD.n3548 0.0089375
R13569 VDD.n3626 VDD.n3624 0.0089375
R13570 VDD.n3657 VDD.n3656 0.0089375
R13571 VDD.n3739 VDD.n3737 0.0089375
R13572 VDD.n5880 VDD.n5879 0.0089375
R13573 VDD.n5993 VDD.n5990 0.0089375
R13574 VDD.n6035 VDD.n6034 0.0089375
R13575 VDD.n6148 VDD.n6145 0.0089375
R13576 VDD.n5564 VDD.n5560 0.0089375
R13577 VDD.n5677 VDD.n5674 0.0089375
R13578 VDD.n5733 VDD.n5732 0.0089375
R13579 VDD.n5846 VDD.n5843 0.0089375
R13580 VDD.n3350 VDD.n3349 0.0089375
R13581 VDD.n3427 VDD.n3425 0.0089375
R13582 VDD.n3456 VDD.n3455 0.0089375
R13583 VDD.n3533 VDD.n3531 0.0089375
R13584 VDD.n2599 VDD.n2598 0.0089375
R13585 VDD.n2681 VDD.n2679 0.0089375
R13586 VDD.n6496 VDD.n6495 0.0089375
R13587 VDD.n6609 VDD.n6606 0.0089375
R13588 VDD.n1520 VDD.n1519 0.00865625
R13589 VDD.n2133 VDD.n2132 0.00865625
R13590 VDD.n2400 VDD.n2397 0.00865625
R13591 VDD.n546 VDD.n534 0.008375
R13592 VDD.n457 VDD.n454 0.008375
R13593 VDD.n7512 VDD.n7503 0.008375
R13594 VDD.n7426 VDD.n7423 0.008375
R13595 VDD.n6232 VDD.n6231 0.008375
R13596 VDD.n6245 VDD.n6242 0.008375
R13597 VDD.n6387 VDD.n6386 0.008375
R13598 VDD.n6400 VDD.n6397 0.008375
R13599 VDD.n5930 VDD.n5929 0.008375
R13600 VDD.n5943 VDD.n5940 0.008375
R13601 VDD.n6085 VDD.n6084 0.008375
R13602 VDD.n6098 VDD.n6095 0.008375
R13603 VDD.n5614 VDD.n5613 0.008375
R13604 VDD.n5627 VDD.n5624 0.008375
R13605 VDD.n5783 VDD.n5782 0.008375
R13606 VDD.n5796 VDD.n5793 0.008375
R13607 VDD.n6546 VDD.n6545 0.008375
R13608 VDD.n6559 VDD.n6556 0.008375
R13609 VDD.n2491 VDD.n2490 0.00809375
R13610 VDD.n7328 VDD.n7327 0.0078125
R13611 VDD.n7097 VDD.n7096 0.0078125
R13612 VDD.n1152 VDD.n1151 0.00753125
R13613 VDD.n1236 VDD.n1234 0.00753125
R13614 VDD.n2370 VDD.n2369 0.00753125
R13615 VDD.n2508 VDD.n2505 0.00753125
R13616 VDD.n2453 VDD.n2452 0.0066875
R13617 VDD.n2477 VDD.n2476 0.00640625
R13618 VDD.n1175 VDD.n1173 0.00584375
R13619 VDD.n1182 VDD.n1181 0.00584375
R13620 VDD.n2407 VDD.n2404 0.00584375
R13621 VDD.n7536 VDD.n7533 0.0055625
R13622 VDD.n578 VDD.n576 0.0055625
R13623 VDD.n632 VDD.n631 0.0055625
R13624 VDD.n3846 VDD.n3841 0.0055625
R13625 VDD.n3851 VDD.n3850 0.0055625
R13626 VDD.n6313 VDD.n6308 0.0055625
R13627 VDD.n6314 VDD.n6313 0.0055625
R13628 VDD.n6320 VDD.n6319 0.0055625
R13629 VDD.n3641 VDD.n3636 0.0055625
R13630 VDD.n3646 VDD.n3645 0.0055625
R13631 VDD.n6011 VDD.n6006 0.0055625
R13632 VDD.n6018 VDD.n6017 0.0055625
R13633 VDD.n5709 VDD.n5690 0.0055625
R13634 VDD.n5716 VDD.n5715 0.0055625
R13635 VDD.n3440 VDD.n3436 0.0055625
R13636 VDD.n3445 VDD.n3444 0.0055625
R13637 VDD.n6627 VDD.n6626 0.0055625
R13638 VDD.n2418 VDD.n2417 0.0055625
R13639 VDD.n1036 VDD.n1033 0.0055625
R13640 VDD.n567 VDD.n566 0.0055625
R13641 VDD.n2466 VDD.n2463 0.00528125
R13642 VDD.n3746 VDD.n3041 0.00479775
R13643 VDD.n3955 VDD.n2911 0.00479775
R13644 VDD.n6483 VDD.n6482 0.00479775
R13645 VDD.n3540 VDD.n3177 0.00479775
R13646 VDD.n1483 VDD.n1481 0.00471875
R13647 VDD.n1646 VDD.n1645 0.00471875
R13648 VDD.n2078 VDD.n2075 0.00471875
R13649 VDD.n2321 VDD.n2320 0.00471875
R13650 VDD.n3339 VDD.n3335 0.00359375
R13651 VDD.n5545 VDD.n5540 0.00359375
R13652 VDD.n3436 VDD.n3265 0.00359375
R13653 VDD.n5690 VDD.n5367 0.00359375
R13654 VDD.n3841 VDD.n2976 0.00359375
R13655 VDD.n6308 VDD.n4385 0.00359375
R13656 VDD.n3851 VDD.n2971 0.00359375
R13657 VDD.n6320 VDD.n4269 0.00359375
R13658 VDD.n3646 VDD.n3104 0.00359375
R13659 VDD.n6018 VDD.n4776 0.00359375
R13660 VDD.n3636 VDD.n3112 0.00359375
R13661 VDD.n6006 VDD.n4889 0.00359375
R13662 VDD.n3445 VDD.n3254 0.00359375
R13663 VDD.n5716 VDD.n5271 0.00359375
R13664 VDD.n2695 VDD.n2693 0.00359375
R13665 VDD.n6627 VDD.n2836 0.00359375
R13666 VDD.n321 VDD.n320 0.0033125
R13667 VDD.n366 VDD.n365 0.0033125
R13668 VDD.n3748 VDD.n3746 0.0033125
R13669 VDD.n3783 VDD.n3781 0.0033125
R13670 VDD.n3804 VDD.n3803 0.0033125
R13671 VDD.n3890 VDD.n3888 0.0033125
R13672 VDD.n3911 VDD.n3910 0.0033125
R13673 VDD.n3955 VDD.n3950 0.0033125
R13674 VDD.n6222 VDD.n6219 0.0033125
R13675 VDD.n6255 VDD.n6254 0.0033125
R13676 VDD.n6377 VDD.n6374 0.0033125
R13677 VDD.n6410 VDD.n6409 0.0033125
R13678 VDD.n6483 VDD.n6459 0.0033125
R13679 VDD.n3542 VDD.n3540 0.0033125
R13680 VDD.n3577 VDD.n3575 0.0033125
R13681 VDD.n3598 VDD.n3597 0.0033125
R13682 VDD.n3685 VDD.n3683 0.0033125
R13683 VDD.n3706 VDD.n3705 0.0033125
R13684 VDD.n3746 VDD.n3745 0.0033125
R13685 VDD.n5920 VDD.n5917 0.0033125
R13686 VDD.n5953 VDD.n5952 0.0033125
R13687 VDD.n6075 VDD.n6072 0.0033125
R13688 VDD.n6108 VDD.n6107 0.0033125
R13689 VDD.n5604 VDD.n5601 0.0033125
R13690 VDD.n5637 VDD.n5636 0.0033125
R13691 VDD.n5773 VDD.n5770 0.0033125
R13692 VDD.n5806 VDD.n5805 0.0033125
R13693 VDD.n3378 VDD.n3376 0.0033125
R13694 VDD.n3399 VDD.n3398 0.0033125
R13695 VDD.n3484 VDD.n3482 0.0033125
R13696 VDD.n3505 VDD.n3504 0.0033125
R13697 VDD.n3540 VDD.n3539 0.0033125
R13698 VDD.n3955 VDD.n3954 0.0033125
R13699 VDD.n2627 VDD.n2625 0.0033125
R13700 VDD.n2648 VDD.n2647 0.0033125
R13701 VDD.n6486 VDD.n6483 0.0033125
R13702 VDD.n6536 VDD.n6533 0.0033125
R13703 VDD.n6569 VDD.n6568 0.0033125
R13704 VDD.n7564 VDD.n7563 0.0033125
R13705 VDD.n7580 VDD.n7578 0.0033125
R13706 VDD.n7697 VDD.n7696 0.0033125
R13707 VDD.n6165 VDD.n4575 0.0032809
R13708 VDD.n5863 VDD.n5075 0.0032809
R13709 VDD.n3767 VDD.n3766 0.00275
R13710 VDD.n3820 VDD.n3818 0.00275
R13711 VDD.n3874 VDD.n3873 0.00275
R13712 VDD.n3927 VDD.n3925 0.00275
R13713 VDD.n6199 VDD.n6198 0.00275
R13714 VDD.n6278 VDD.n6275 0.00275
R13715 VDD.n6354 VDD.n6353 0.00275
R13716 VDD.n6433 VDD.n6430 0.00275
R13717 VDD.n3561 VDD.n3560 0.00275
R13718 VDD.n3614 VDD.n3612 0.00275
R13719 VDD.n3669 VDD.n3668 0.00275
R13720 VDD.n3722 VDD.n3720 0.00275
R13721 VDD.n5897 VDD.n5896 0.00275
R13722 VDD.n5976 VDD.n5973 0.00275
R13723 VDD.n6052 VDD.n6051 0.00275
R13724 VDD.n6131 VDD.n6128 0.00275
R13725 VDD.n5581 VDD.n5580 0.00275
R13726 VDD.n5660 VDD.n5657 0.00275
R13727 VDD.n5750 VDD.n5749 0.00275
R13728 VDD.n5829 VDD.n5826 0.00275
R13729 VDD.n3362 VDD.n3361 0.00275
R13730 VDD.n3415 VDD.n3413 0.00275
R13731 VDD.n3468 VDD.n3467 0.00275
R13732 VDD.n3521 VDD.n3519 0.00275
R13733 VDD.n2611 VDD.n2610 0.00275
R13734 VDD.n2664 VDD.n2662 0.00275
R13735 VDD.n6513 VDD.n6512 0.00275
R13736 VDD.n6592 VDD.n6589 0.00275
R13737 VDD.n1537 VDD.n1536 0.00246875
R13738 VDD.n1665 VDD.n1664 0.00246875
R13739 VDD.n2160 VDD.n2159 0.00246875
R13740 VDD.n2351 VDD.n2350 0.00246875
R13741 VDD.n7116 VDD.n7115 0.0021875
R13742 VDD.n7250 VDD.n7247 0.0021875
R13743 VDD.n5867 VDD.n5864 0.001625
R13744 VDD.n6022 VDD.n6019 0.001625
R13745 VDD.n1157 VDD.n1155 0.00134375
R13746 VDD.n1231 VDD.n1230 0.00134375
R13747 VDD.n2377 VDD.n2374 0.00134375
R13748 VDD.n2389 VDD.n2388 0.00134375
R13749 VDD.n2473 VDD.n2470 0.00134375
R13750 VDD.n2501 VDD.n2500 0.00134375
R13751 VDD.n7537 VDD.n7357 0.0010625
R13752 VDD.n3760 VDD.n3759 0.0010625
R13753 VDD.n3827 VDD.n3825 0.0010625
R13754 VDD.n3867 VDD.n3866 0.0010625
R13755 VDD.n3934 VDD.n3932 0.0010625
R13756 VDD.n6189 VDD.n6188 0.0010625
R13757 VDD.n6288 VDD.n6285 0.0010625
R13758 VDD.n6344 VDD.n6343 0.0010625
R13759 VDD.n6443 VDD.n6440 0.0010625
R13760 VDD.n3554 VDD.n3553 0.0010625
R13761 VDD.n3621 VDD.n3619 0.0010625
R13762 VDD.n3662 VDD.n3661 0.0010625
R13763 VDD.n3729 VDD.n3727 0.0010625
R13764 VDD.n5887 VDD.n5886 0.0010625
R13765 VDD.n5986 VDD.n5983 0.0010625
R13766 VDD.n6042 VDD.n6041 0.0010625
R13767 VDD.n6141 VDD.n6138 0.0010625
R13768 VDD.n5571 VDD.n5570 0.0010625
R13769 VDD.n5670 VDD.n5667 0.0010625
R13770 VDD.n5740 VDD.n5739 0.0010625
R13771 VDD.n5839 VDD.n5836 0.0010625
R13772 VDD.n3355 VDD.n3354 0.0010625
R13773 VDD.n3422 VDD.n3420 0.0010625
R13774 VDD.n3461 VDD.n3460 0.0010625
R13775 VDD.n3528 VDD.n3526 0.0010625
R13776 VDD.n2604 VDD.n2603 0.0010625
R13777 VDD.n2671 VDD.n2669 0.0010625
R13778 VDD.n6503 VDD.n6502 0.0010625
R13779 VDD.n6602 VDD.n6599 0.0010625
R13780 VDD.n2056 VDD.n2039 0.00078125
R13781 VDD.n2160 VDD.n1935 0.00078125
R13782 VDD.n2351 VDD.n1797 0.00078125
R13783 VDD.n1667 VDD.n1665 0.00078125
R13784 VDD.n2541 VDD.n1351 0.00078125
R13785 VDD.n1252 VDD.n1250 0.00078125
R13786 VDD.n2417 VDD.n2416 0.00078125
R13787 VDD.n2442 VDD.n2441 0.00078125
R13788 IBIAS2.n214 IBIAS2.t264 81.7344
R13789 IBIAS2.n215 IBIAS2.t388 81.7344
R13790 IBIAS2.n216 IBIAS2.t405 81.7344
R13791 IBIAS2.n217 IBIAS2.t528 81.7344
R13792 IBIAS2.n218 IBIAS2.t399 81.7344
R13793 IBIAS2.n219 IBIAS2.t521 81.7344
R13794 IBIAS2.n220 IBIAS2.t221 81.7344
R13795 IBIAS2.n231 IBIAS2.t373 81.7344
R13796 IBIAS2.n230 IBIAS2.t353 81.7344
R13797 IBIAS2.n229 IBIAS2.t480 81.7344
R13798 IBIAS2.n228 IBIAS2.t498 81.7344
R13799 IBIAS2.n227 IBIAS2.t193 81.7344
R13800 IBIAS2.n226 IBIAS2.t211 81.7344
R13801 IBIAS2.n225 IBIAS2.t331 81.7344
R13802 IBIAS2.n317 IBIAS2.t484 81.7344
R13803 IBIAS2.n318 IBIAS2.t461 81.7344
R13804 IBIAS2.n319 IBIAS2.t160 81.7344
R13805 IBIAS2.n320 IBIAS2.t183 81.7344
R13806 IBIAS2.n321 IBIAS2.t304 81.7344
R13807 IBIAS2.n322 IBIAS2.t316 81.7344
R13808 IBIAS2.n323 IBIAS2.t439 81.7344
R13809 IBIAS2.n334 IBIAS2.t138 81.7344
R13810 IBIAS2.n333 IBIAS2.t151 81.7344
R13811 IBIAS2.n332 IBIAS2.t267 81.7344
R13812 IBIAS2.n331 IBIAS2.t393 81.7344
R13813 IBIAS2.n330 IBIAS2.t406 81.7344
R13814 IBIAS2.n329 IBIAS2.t387 81.7344
R13815 IBIAS2.n328 IBIAS2.t403 81.7344
R13816 IBIAS2.n420 IBIAS2.t467 81.7344
R13817 IBIAS2.n421 IBIAS2.t168 81.7344
R13818 IBIAS2.n422 IBIAS2.t462 81.7344
R13819 IBIAS2.n423 IBIAS2.t161 81.7344
R13820 IBIAS2.n424 IBIAS2.t281 81.7344
R13821 IBIAS2.n425 IBIAS2.t302 81.7344
R13822 IBIAS2.n426 IBIAS2.t420 81.7344
R13823 IBIAS2.n437 IBIAS2.t538 81.7344
R13824 IBIAS2.n436 IBIAS2.t136 81.7344
R13825 IBIAS2.n435 IBIAS2.t248 81.7344
R13826 IBIAS2.n434 IBIAS2.t268 81.7344
R13827 IBIAS2.n433 IBIAS2.t391 81.7344
R13828 IBIAS2.n432 IBIAS2.t368 81.7344
R13829 IBIAS2.n431 IBIAS2.t385 81.7344
R13830 IBIAS2.n523 IBIAS2.t222 81.7344
R13831 IBIAS2.n524 IBIAS2.t235 81.7344
R13832 IBIAS2.n525 IBIAS2.t356 81.7344
R13833 IBIAS2.n526 IBIAS2.t372 81.7344
R13834 IBIAS2.n527 IBIAS2.t501 81.7344
R13835 IBIAS2.n528 IBIAS2.t481 81.7344
R13836 IBIAS2.n529 IBIAS2.t496 81.7344
R13837 IBIAS2.n540 IBIAS2.t332 81.7344
R13838 IBIAS2.n539 IBIAS2.t454 81.7344
R13839 IBIAS2.n538 IBIAS2.t475 81.7344
R13840 IBIAS2.n537 IBIAS2.t447 81.7344
R13841 IBIAS2.n536 IBIAS2.t465 81.7344
R13842 IBIAS2.n535 IBIAS2.t167 81.7344
R13843 IBIAS2.n534 IBIAS2.t286 81.7344
R13844 IBIAS2.n626 IBIAS2.t210 81.7344
R13845 IBIAS2.n627 IBIAS2.t329 81.7344
R13846 IBIAS2.n628 IBIAS2.t345 81.7344
R13847 IBIAS2.n629 IBIAS2.t476 81.7344
R13848 IBIAS2.n630 IBIAS2.t175 81.7344
R13849 IBIAS2.n631 IBIAS2.t189 81.7344
R13850 IBIAS2.n632 IBIAS2.t166 81.7344
R13851 IBIAS2.n643 IBIAS2.t423 81.7344
R13852 IBIAS2.n642 IBIAS2.t440 81.7344
R13853 IBIAS2.n641 IBIAS2.t141 81.7344
R13854 IBIAS2.n640 IBIAS2.t157 81.7344
R13855 IBIAS2.n639 IBIAS2.t140 81.7344
R13856 IBIAS2.n638 IBIAS2.t253 81.7344
R13857 IBIAS2.n637 IBIAS2.t271 81.7344
R13858 IBIAS2.n729 IBIAS2.t530 81.7344
R13859 IBIAS2.n730 IBIAS2.t124 81.7344
R13860 IBIAS2.n731 IBIAS2.t242 81.7344
R13861 IBIAS2.n732 IBIAS2.t259 81.7344
R13862 IBIAS2.n733 IBIAS2.t240 81.7344
R13863 IBIAS2.n734 IBIAS2.t358 81.7344
R13864 IBIAS2.n735 IBIAS2.t378 81.7344
R13865 IBIAS2.n746 IBIAS2.t219 81.7344
R13866 IBIAS2.n745 IBIAS2.t197 81.7344
R13867 IBIAS2.n744 IBIAS2.t213 81.7344
R13868 IBIAS2.n743 IBIAS2.t336 81.7344
R13869 IBIAS2.n742 IBIAS2.t348 81.7344
R13870 IBIAS2.n741 IBIAS2.t478 81.7344
R13871 IBIAS2.n740 IBIAS2.t179 81.7344
R13872 IBIAS2.n116 IBIAS2.t180 81.7344
R13873 IBIAS2.n117 IBIAS2.t293 81.7344
R13874 IBIAS2.n118 IBIAS2.t417 81.7344
R13875 IBIAS2.n119 IBIAS2.t288 81.7344
R13876 IBIAS2.n120 IBIAS2.t412 81.7344
R13877 IBIAS2.n121 IBIAS2.t428 81.7344
R13878 IBIAS2.n122 IBIAS2.t133 81.7344
R13879 IBIAS2.n133 IBIAS2.t243 81.7344
R13880 IBIAS2.n132 IBIAS2.t260 81.7344
R13881 IBIAS2.n131 IBIAS2.t382 81.7344
R13882 IBIAS2.n130 IBIAS2.t512 81.7344
R13883 IBIAS2.n129 IBIAS2.t522 81.7344
R13884 IBIAS2.n128 IBIAS2.t223 81.7344
R13885 IBIAS2.n127 IBIAS2.t236 81.7344
R13886 IBIAS2.n155 IBIAS2.t50 53.5894
R13887 IBIAS2.n152 IBIAS2.t88 53.5894
R13888 IBIAS2.n258 IBIAS2.t26 53.5894
R13889 IBIAS2.n255 IBIAS2.t32 53.5894
R13890 IBIAS2.n361 IBIAS2.t30 53.5894
R13891 IBIAS2.n358 IBIAS2.t24 53.5894
R13892 IBIAS2.n464 IBIAS2.t92 53.5894
R13893 IBIAS2.n461 IBIAS2.t98 53.5894
R13894 IBIAS2.n567 IBIAS2.t70 53.5894
R13895 IBIAS2.n564 IBIAS2.t100 53.5894
R13896 IBIAS2.n670 IBIAS2.t10 53.5894
R13897 IBIAS2.n667 IBIAS2.t16 53.5894
R13898 IBIAS2.n16 IBIAS2.t78 53.5894
R13899 IBIAS2.n11 IBIAS2.t84 53.5894
R13900 IBIAS2.n176 IBIAS2.t18 47.0594
R13901 IBIAS2.n204 IBIAS2.t80 47.0594
R13902 IBIAS2.n232 IBIAS2.t6 47.0594
R13903 IBIAS2.n165 IBIAS2.t40 47.0594
R13904 IBIAS2.n193 IBIAS2.t110 47.0594
R13905 IBIAS2.n221 IBIAS2.t74 47.0594
R13906 IBIAS2.n214 IBIAS2.t250 47.0594
R13907 IBIAS2.n215 IBIAS2.t500 47.0594
R13908 IBIAS2.n216 IBIAS2.t426 47.0594
R13909 IBIAS2.n217 IBIAS2.t245 47.0594
R13910 IBIAS2.n218 IBIAS2.t285 47.0594
R13911 IBIAS2.n219 IBIAS2.t529 47.0594
R13912 IBIAS2.n220 IBIAS2.t346 47.0594
R13913 IBIAS2.n231 IBIAS2.t450 47.0594
R13914 IBIAS2.n230 IBIAS2.t375 47.0594
R13915 IBIAS2.n229 IBIAS2.t198 47.0594
R13916 IBIAS2.n228 IBIAS2.t131 47.0594
R13917 IBIAS2.n227 IBIAS2.t367 47.0594
R13918 IBIAS2.n170 IBIAS2.t227 47.0594
R13919 IBIAS2.n158 IBIAS2.t146 47.0594
R13920 IBIAS2.n186 IBIAS2.t177 47.0594
R13921 IBIAS2.n159 IBIAS2.t230 47.0594
R13922 IBIAS2.n187 IBIAS2.t291 47.0594
R13923 IBIAS2.n160 IBIAS2.t464 47.0594
R13924 IBIAS2.n188 IBIAS2.t313 47.0594
R13925 IBIAS2.n161 IBIAS2.t135 47.0594
R13926 IBIAS2.n189 IBIAS2.t430 47.0594
R13927 IBIAS2.n162 IBIAS2.t410 47.0594
R13928 IBIAS2.n190 IBIAS2.t310 47.0594
R13929 IBIAS2.n163 IBIAS2.t502 47.0594
R13930 IBIAS2.n191 IBIAS2.t424 47.0594
R13931 IBIAS2.n164 IBIAS2.t169 47.0594
R13932 IBIAS2.n192 IBIAS2.t129 47.0594
R13933 IBIAS2.n175 IBIAS2.t294 47.0594
R13934 IBIAS2.n203 IBIAS2.t280 47.0594
R13935 IBIAS2.n174 IBIAS2.t431 47.0594
R13936 IBIAS2.n202 IBIAS2.t255 47.0594
R13937 IBIAS2.n173 IBIAS2.t520 47.0594
R13938 IBIAS2.n201 IBIAS2.t381 47.0594
R13939 IBIAS2.n172 IBIAS2.t328 47.0594
R13940 IBIAS2.n200 IBIAS2.t396 47.0594
R13941 IBIAS2.n171 IBIAS2.t418 47.0594
R13942 IBIAS2.n199 IBIAS2.t517 47.0594
R13943 IBIAS2.n169 IBIAS2.t317 47.0594
R13944 IBIAS2.n197 IBIAS2.t234 47.0594
R13945 IBIAS2.n198 IBIAS2.t537 47.0594
R13946 IBIAS2.n226 IBIAS2.t306 47.0594
R13947 IBIAS2.n225 IBIAS2.t541 47.0594
R13948 IBIAS2.n279 IBIAS2.t42 47.0594
R13949 IBIAS2.n307 IBIAS2.t58 47.0594
R13950 IBIAS2.n335 IBIAS2.t86 47.0594
R13951 IBIAS2.n268 IBIAS2.t108 47.0594
R13952 IBIAS2.n296 IBIAS2.t62 47.0594
R13953 IBIAS2.n324 IBIAS2.t66 47.0594
R13954 IBIAS2.n317 IBIAS2.t299 47.0594
R13955 IBIAS2.n318 IBIAS2.t226 47.0594
R13956 IBIAS2.n319 IBIAS2.t472 47.0594
R13957 IBIAS2.n320 IBIAS2.t395 47.0594
R13958 IBIAS2.n321 IBIAS2.t218 47.0594
R13959 IBIAS2.n322 IBIAS2.t152 47.0594
R13960 IBIAS2.n323 IBIAS2.t390 47.0594
R13961 IBIAS2.n334 IBIAS2.t492 47.0594
R13962 IBIAS2.n333 IBIAS2.t421 47.0594
R13963 IBIAS2.n332 IBIAS2.t239 47.0594
R13964 IBIAS2.n331 IBIAS2.t485 47.0594
R13965 IBIAS2.n330 IBIAS2.t415 47.0594
R13966 IBIAS2.n273 IBIAS2.t398 47.0594
R13967 IBIAS2.n261 IBIAS2.t408 47.0594
R13968 IBIAS2.n289 IBIAS2.t384 47.0594
R13969 IBIAS2.n262 IBIAS2.t126 47.0594
R13970 IBIAS2.n290 IBIAS2.t362 47.0594
R13971 IBIAS2.n263 IBIAS2.t214 47.0594
R13972 IBIAS2.n291 IBIAS2.t489 47.0594
R13973 IBIAS2.n264 IBIAS2.t445 47.0594
R13974 IBIAS2.n292 IBIAS2.t511 47.0594
R13975 IBIAS2.n265 IBIAS2.t532 47.0594
R13976 IBIAS2.n293 IBIAS2.t205 47.0594
R13977 IBIAS2.n266 IBIAS2.t340 47.0594
R13978 IBIAS2.n294 IBIAS2.t220 47.0594
R13979 IBIAS2.n267 IBIAS2.t432 47.0594
R13980 IBIAS2.n295 IBIAS2.t339 47.0594
R13981 IBIAS2.n278 IBIAS2.t468 47.0594
R13982 IBIAS2.n306 IBIAS2.t459 47.0594
R13983 IBIAS2.n277 IBIAS2.t274 47.0594
R13984 IBIAS2.n305 IBIAS2.t479 47.0594
R13985 IBIAS2.n276 IBIAS2.t359 47.0594
R13986 IBIAS2.n304 IBIAS2.t182 47.0594
R13987 IBIAS2.n275 IBIAS2.t452 47.0594
R13988 IBIAS2.n303 IBIAS2.t300 47.0594
R13989 IBIAS2.n274 IBIAS2.t257 47.0594
R13990 IBIAS2.n302 IBIAS2.t315 47.0594
R13991 IBIAS2.n272 IBIAS2.t209 47.0594
R13992 IBIAS2.n300 IBIAS2.t311 47.0594
R13993 IBIAS2.n301 IBIAS2.t290 47.0594
R13994 IBIAS2.n329 IBIAS2.t338 47.0594
R13995 IBIAS2.n328 IBIAS2.t269 47.0594
R13996 IBIAS2.n382 IBIAS2.t14 47.0594
R13997 IBIAS2.n410 IBIAS2.t64 47.0594
R13998 IBIAS2.n438 IBIAS2.t82 47.0594
R13999 IBIAS2.n371 IBIAS2.t46 47.0594
R14000 IBIAS2.n399 IBIAS2.t56 47.0594
R14001 IBIAS2.n427 IBIAS2.t60 47.0594
R14002 IBIAS2.n420 IBIAS2.t314 47.0594
R14003 IBIAS2.n421 IBIAS2.t137 47.0594
R14004 IBIAS2.n422 IBIAS2.t172 47.0594
R14005 IBIAS2.n423 IBIAS2.t407 47.0594
R14006 IBIAS2.n424 IBIAS2.t229 47.0594
R14007 IBIAS2.n425 IBIAS2.t163 47.0594
R14008 IBIAS2.n426 IBIAS2.t404 47.0594
R14009 IBIAS2.n437 IBIAS2.t510 47.0594
R14010 IBIAS2.n436 IBIAS2.t435 47.0594
R14011 IBIAS2.n435 IBIAS2.t249 47.0594
R14012 IBIAS2.n434 IBIAS2.t188 47.0594
R14013 IBIAS2.n433 IBIAS2.t425 47.0594
R14014 IBIAS2.n376 IBIAS2.t524 47.0594
R14015 IBIAS2.n364 IBIAS2.t534 47.0594
R14016 IBIAS2.n392 IBIAS2.t366 47.0594
R14017 IBIAS2.n365 IBIAS2.t203 47.0594
R14018 IBIAS2.n393 IBIAS2.t495 47.0594
R14019 IBIAS2.n366 IBIAS2.t483 47.0594
R14020 IBIAS2.n394 IBIAS2.t361 47.0594
R14021 IBIAS2.n367 IBIAS2.t150 47.0594
R14022 IBIAS2.n395 IBIAS2.t488 47.0594
R14023 IBIAS2.n368 IBIAS2.t232 47.0594
R14024 IBIAS2.n396 IBIAS2.t190 47.0594
R14025 IBIAS2.n369 IBIAS2.t473 47.0594
R14026 IBIAS2.n397 IBIAS2.t204 47.0594
R14027 IBIAS2.n370 IBIAS2.t139 47.0594
R14028 IBIAS2.n398 IBIAS2.t325 47.0594
R14029 IBIAS2.n381 IBIAS2.t174 47.0594
R14030 IBIAS2.n409 IBIAS2.t442 47.0594
R14031 IBIAS2.n380 IBIAS2.t401 47.0594
R14032 IBIAS2.n408 IBIAS2.t460 47.0594
R14033 IBIAS2.n379 IBIAS2.t491 47.0594
R14034 IBIAS2.n407 IBIAS2.t158 47.0594
R14035 IBIAS2.n378 IBIAS2.t303 47.0594
R14036 IBIAS2.n406 IBIAS2.t181 47.0594
R14037 IBIAS2.n377 IBIAS2.t386 47.0594
R14038 IBIAS2.n405 IBIAS2.t296 47.0594
R14039 IBIAS2.n375 IBIAS2.t334 47.0594
R14040 IBIAS2.n403 IBIAS2.t289 47.0594
R14041 IBIAS2.n404 IBIAS2.t275 47.0594
R14042 IBIAS2.n432 IBIAS2.t352 47.0594
R14043 IBIAS2.n431 IBIAS2.t283 47.0594
R14044 IBIAS2.n485 IBIAS2.t52 47.0594
R14045 IBIAS2.n513 IBIAS2.t2 47.0594
R14046 IBIAS2.n541 IBIAS2.t68 47.0594
R14047 IBIAS2.n474 IBIAS2.t0 47.0594
R14048 IBIAS2.n502 IBIAS2.t8 47.0594
R14049 IBIAS2.n530 IBIAS2.t44 47.0594
R14050 IBIAS2.n523 IBIAS2.t347 47.0594
R14051 IBIAS2.n524 IBIAS2.t278 47.0594
R14052 IBIAS2.n525 IBIAS2.t525 47.0594
R14053 IBIAS2.n526 IBIAS2.t455 47.0594
R14054 IBIAS2.n527 IBIAS2.t272 47.0594
R14055 IBIAS2.n528 IBIAS2.t199 47.0594
R14056 IBIAS2.n529 IBIAS2.t134 47.0594
R14057 IBIAS2.n540 IBIAS2.t123 47.0594
R14058 IBIAS2.n539 IBIAS2.t363 47.0594
R14059 IBIAS2.n538 IBIAS2.t297 47.0594
R14060 IBIAS2.n537 IBIAS2.t224 47.0594
R14061 IBIAS2.n536 IBIAS2.t156 47.0594
R14062 IBIAS2.n479 IBIAS2.t364 47.0594
R14063 IBIAS2.n467 IBIAS2.t282 47.0594
R14064 IBIAS2.n495 IBIAS2.t128 47.0594
R14065 IBIAS2.n468 IBIAS2.t515 47.0594
R14066 IBIAS2.n496 IBIAS2.t144 47.0594
R14067 IBIAS2.n469 IBIAS2.t186 47.0594
R14068 IBIAS2.n497 IBIAS2.t262 47.0594
R14069 IBIAS2.n470 IBIAS2.t413 47.0594
R14070 IBIAS2.n498 IBIAS2.t279 47.0594
R14071 IBIAS2.n471 IBIAS2.t507 47.0594
R14072 IBIAS2.n499 IBIAS2.t402 47.0594
R14073 IBIAS2.n472 IBIAS2.t216 47.0594
R14074 IBIAS2.n500 IBIAS2.t380 47.0594
R14075 IBIAS2.n473 IBIAS2.t446 47.0594
R14076 IBIAS2.n501 IBIAS2.t397 47.0594
R14077 IBIAS2.n484 IBIAS2.t436 47.0594
R14078 IBIAS2.n512 IBIAS2.t233 47.0594
R14079 IBIAS2.n483 IBIAS2.t523 47.0594
R14080 IBIAS2.n511 IBIAS2.t355 47.0594
R14081 IBIAS2.n482 IBIAS2.t333 47.0594
R14082 IBIAS2.n510 IBIAS2.t371 47.0594
R14083 IBIAS2.n481 IBIAS2.t474 47.0594
R14084 IBIAS2.n509 IBIAS2.t351 47.0594
R14085 IBIAS2.n480 IBIAS2.t277 47.0594
R14086 IBIAS2.n508 IBIAS2.t365 47.0594
R14087 IBIAS2.n478 IBIAS2.t456 47.0594
R14088 IBIAS2.n506 IBIAS2.t191 47.0594
R14089 IBIAS2.n507 IBIAS2.t494 47.0594
R14090 IBIAS2.n535 IBIAS2.t394 47.0594
R14091 IBIAS2.n534 IBIAS2.t217 47.0594
R14092 IBIAS2.n588 IBIAS2.t48 47.0594
R14093 IBIAS2.n616 IBIAS2.t96 47.0594
R14094 IBIAS2.n644 IBIAS2.t72 47.0594
R14095 IBIAS2.n577 IBIAS2.t76 47.0594
R14096 IBIAS2.n605 IBIAS2.t12 47.0594
R14097 IBIAS2.n633 IBIAS2.t20 47.0594
R14098 IBIAS2.n626 IBIAS2.t458 47.0594
R14099 IBIAS2.n627 IBIAS2.t276 47.0594
R14100 IBIAS2.n628 IBIAS2.t206 47.0594
R14101 IBIAS2.n629 IBIAS2.t448 47.0594
R14102 IBIAS2.n630 IBIAS2.t270 47.0594
R14103 IBIAS2.n631 IBIAS2.t200 47.0594
R14104 IBIAS2.n632 IBIAS2.t130 47.0594
R14105 IBIAS2.n643 IBIAS2.t540 47.0594
R14106 IBIAS2.n642 IBIAS2.t477 47.0594
R14107 IBIAS2.n641 IBIAS2.t292 47.0594
R14108 IBIAS2.n640 IBIAS2.t225 47.0594
R14109 IBIAS2.n639 IBIAS2.t153 47.0594
R14110 IBIAS2.n582 IBIAS2.t383 47.0594
R14111 IBIAS2.n570 IBIAS2.t444 47.0594
R14112 IBIAS2.n598 IBIAS2.t535 47.0594
R14113 IBIAS2.n571 IBIAS2.t533 47.0594
R14114 IBIAS2.n599 IBIAS2.t231 47.0594
R14115 IBIAS2.n572 IBIAS2.t341 47.0594
R14116 IBIAS2.n600 IBIAS2.t247 47.0594
R14117 IBIAS2.n573 IBIAS2.t429 47.0594
R14118 IBIAS2.n601 IBIAS2.t369 47.0594
R14119 IBIAS2.n574 IBIAS2.t518 47.0594
R14120 IBIAS2.n602 IBIAS2.t499 47.0594
R14121 IBIAS2.n575 IBIAS2.t327 47.0594
R14122 IBIAS2.n603 IBIAS2.t513 47.0594
R14123 IBIAS2.n576 IBIAS2.t469 47.0594
R14124 IBIAS2.n604 IBIAS2.t493 47.0594
R14125 IBIAS2.n587 IBIAS2.t453 47.0594
R14126 IBIAS2.n615 IBIAS2.t326 47.0594
R14127 IBIAS2.n586 IBIAS2.t258 47.0594
R14128 IBIAS2.n614 IBIAS2.t343 47.0594
R14129 IBIAS2.n585 IBIAS2.t350 47.0594
R14130 IBIAS2.n613 IBIAS2.t470 47.0594
R14131 IBIAS2.n584 IBIAS2.t162 47.0594
R14132 IBIAS2.n612 IBIAS2.t486 47.0594
R14133 IBIAS2.n583 IBIAS2.t298 47.0594
R14134 IBIAS2.n611 IBIAS2.t463 47.0594
R14135 IBIAS2.n581 IBIAS2.t195 47.0594
R14136 IBIAS2.n609 IBIAS2.t184 47.0594
R14137 IBIAS2.n610 IBIAS2.t164 47.0594
R14138 IBIAS2.n638 IBIAS2.t392 47.0594
R14139 IBIAS2.n637 IBIAS2.t323 47.0594
R14140 IBIAS2.n691 IBIAS2.t94 47.0594
R14141 IBIAS2.n719 IBIAS2.t28 47.0594
R14142 IBIAS2.n747 IBIAS2.t54 47.0594
R14143 IBIAS2.n680 IBIAS2.t38 47.0594
R14144 IBIAS2.n708 IBIAS2.t36 47.0594
R14145 IBIAS2.n736 IBIAS2.t34 47.0594
R14146 IBIAS2.n729 IBIAS2.t389 47.0594
R14147 IBIAS2.n730 IBIAS2.t320 47.0594
R14148 IBIAS2.n731 IBIAS2.t143 47.0594
R14149 IBIAS2.n732 IBIAS2.t497 47.0594
R14150 IBIAS2.n733 IBIAS2.t419 47.0594
R14151 IBIAS2.n734 IBIAS2.t238 47.0594
R14152 IBIAS2.n735 IBIAS2.t176 47.0594
R14153 IBIAS2.n746 IBIAS2.t165 47.0594
R14154 IBIAS2.n745 IBIAS2.t514 47.0594
R14155 IBIAS2.n744 IBIAS2.t441 47.0594
R14156 IBIAS2.n743 IBIAS2.t261 47.0594
R14157 IBIAS2.n742 IBIAS2.t192 47.0594
R14158 IBIAS2.n685 IBIAS2.t228 47.0594
R14159 IBIAS2.n673 IBIAS2.t147 47.0594
R14160 IBIAS2.n701 IBIAS2.t437 47.0594
R14161 IBIAS2.n674 IBIAS2.t374 47.0594
R14162 IBIAS2.n702 IBIAS2.t451 47.0594
R14163 IBIAS2.n675 IBIAS2.t466 47.0594
R14164 IBIAS2.n703 IBIAS2.t154 47.0594
R14165 IBIAS2.n676 IBIAS2.t273 47.0594
R14166 IBIAS2.n704 IBIAS2.t170 47.0594
R14167 IBIAS2.n677 IBIAS2.t411 47.0594
R14168 IBIAS2.n705 IBIAS2.t148 47.0594
R14169 IBIAS2.n678 IBIAS2.t503 47.0594
R14170 IBIAS2.n706 IBIAS2.t266 47.0594
R14171 IBIAS2.n679 IBIAS2.t312 47.0594
R14172 IBIAS2.n707 IBIAS2.t284 47.0594
R14173 IBIAS2.n690 IBIAS2.t295 47.0594
R14174 IBIAS2.n718 IBIAS2.t122 47.0594
R14175 IBIAS2.n689 IBIAS2.t433 47.0594
R14176 IBIAS2.n717 IBIAS2.t526 47.0594
R14177 IBIAS2.n688 IBIAS2.t241 47.0594
R14178 IBIAS2.n716 IBIAS2.t539 47.0594
R14179 IBIAS2.n687 IBIAS2.t330 47.0594
R14180 IBIAS2.n715 IBIAS2.t237 47.0594
R14181 IBIAS2.n686 IBIAS2.t142 47.0594
R14182 IBIAS2.n714 IBIAS2.t251 47.0594
R14183 IBIAS2.n684 IBIAS2.t318 47.0594
R14184 IBIAS2.n712 IBIAS2.t504 47.0594
R14185 IBIAS2.n713 IBIAS2.t377 47.0594
R14186 IBIAS2.n741 IBIAS2.t438 47.0594
R14187 IBIAS2.n740 IBIAS2.t252 47.0594
R14188 IBIAS2.n27 IBIAS2.t90 47.0594
R14189 IBIAS2.n38 IBIAS2.t22 47.0594
R14190 IBIAS2.n96 IBIAS2.t106 47.0594
R14191 IBIAS2.n107 IBIAS2.t102 47.0594
R14192 IBIAS2.n134 IBIAS2.t4 47.0594
R14193 IBIAS2.n123 IBIAS2.t104 47.0594
R14194 IBIAS2.n116 IBIAS2.t254 47.0594
R14195 IBIAS2.n117 IBIAS2.t505 47.0594
R14196 IBIAS2.n118 IBIAS2.t322 47.0594
R14197 IBIAS2.n119 IBIAS2.t354 47.0594
R14198 IBIAS2.n120 IBIAS2.t185 47.0594
R14199 IBIAS2.n121 IBIAS2.t531 47.0594
R14200 IBIAS2.n122 IBIAS2.t349 47.0594
R14201 IBIAS2.n133 IBIAS2.t449 47.0594
R14202 IBIAS2.n132 IBIAS2.t379 47.0594
R14203 IBIAS2.n131 IBIAS2.t201 47.0594
R14204 IBIAS2.n130 IBIAS2.t443 47.0594
R14205 IBIAS2.n129 IBIAS2.t370 47.0594
R14206 IBIAS2.n32 IBIAS2.t490 47.0594
R14207 IBIAS2.n20 IBIAS2.t127 47.0594
R14208 IBIAS2.n89 IBIAS2.t506 47.0594
R14209 IBIAS2.n21 IBIAS2.t215 47.0594
R14210 IBIAS2.n90 IBIAS2.t202 47.0594
R14211 IBIAS2.n22 IBIAS2.t308 47.0594
R14212 IBIAS2.n91 IBIAS2.t324 47.0594
R14213 IBIAS2.n23 IBIAS2.t159 47.0594
R14214 IBIAS2.n92 IBIAS2.t196 47.0594
R14215 IBIAS2.n24 IBIAS2.t246 47.0594
R14216 IBIAS2.n93 IBIAS2.t319 47.0594
R14217 IBIAS2.n25 IBIAS2.t482 47.0594
R14218 IBIAS2.n94 IBIAS2.t335 47.0594
R14219 IBIAS2.n26 IBIAS2.t149 47.0594
R14220 IBIAS2.n95 IBIAS2.t457 47.0594
R14221 IBIAS2.n37 IBIAS2.t187 47.0594
R14222 IBIAS2.n106 IBIAS2.t155 47.0594
R14223 IBIAS2.n36 IBIAS2.t414 47.0594
R14224 IBIAS2.n105 IBIAS2.t171 47.0594
R14225 IBIAS2.n35 IBIAS2.t508 47.0594
R14226 IBIAS2.n104 IBIAS2.t287 47.0594
R14227 IBIAS2.n34 IBIAS2.t173 47.0594
R14228 IBIAS2.n103 IBIAS2.t409 47.0594
R14229 IBIAS2.n33 IBIAS2.t400 47.0594
R14230 IBIAS2.n102 IBIAS2.t427 47.0594
R14231 IBIAS2.n31 IBIAS2.t301 47.0594
R14232 IBIAS2.n100 IBIAS2.t145 47.0594
R14233 IBIAS2.n101 IBIAS2.t132 47.0594
R14234 IBIAS2.n128 IBIAS2.t194 47.0594
R14235 IBIAS2.n127 IBIAS2.t125 47.0594
R14236 IBIAS2.n159 IBIAS2.n158 16.2227
R14237 IBIAS2.n160 IBIAS2.n159 16.2227
R14238 IBIAS2.n161 IBIAS2.n160 16.2227
R14239 IBIAS2.n162 IBIAS2.n161 16.2227
R14240 IBIAS2.n163 IBIAS2.n162 16.2227
R14241 IBIAS2.n164 IBIAS2.n163 16.2227
R14242 IBIAS2.n165 IBIAS2.n164 16.2227
R14243 IBIAS2.n176 IBIAS2.n175 16.2227
R14244 IBIAS2.n175 IBIAS2.n174 16.2227
R14245 IBIAS2.n174 IBIAS2.n173 16.2227
R14246 IBIAS2.n173 IBIAS2.n172 16.2227
R14247 IBIAS2.n172 IBIAS2.n171 16.2227
R14248 IBIAS2.n171 IBIAS2.n170 16.2227
R14249 IBIAS2.n170 IBIAS2.n169 16.2227
R14250 IBIAS2.n187 IBIAS2.n186 16.2227
R14251 IBIAS2.n188 IBIAS2.n187 16.2227
R14252 IBIAS2.n189 IBIAS2.n188 16.2227
R14253 IBIAS2.n190 IBIAS2.n189 16.2227
R14254 IBIAS2.n191 IBIAS2.n190 16.2227
R14255 IBIAS2.n192 IBIAS2.n191 16.2227
R14256 IBIAS2.n193 IBIAS2.n192 16.2227
R14257 IBIAS2.n204 IBIAS2.n203 16.2227
R14258 IBIAS2.n203 IBIAS2.n202 16.2227
R14259 IBIAS2.n202 IBIAS2.n201 16.2227
R14260 IBIAS2.n201 IBIAS2.n200 16.2227
R14261 IBIAS2.n200 IBIAS2.n199 16.2227
R14262 IBIAS2.n199 IBIAS2.n198 16.2227
R14263 IBIAS2.n198 IBIAS2.n197 16.2227
R14264 IBIAS2.n215 IBIAS2.n214 16.2227
R14265 IBIAS2.n216 IBIAS2.n215 16.2227
R14266 IBIAS2.n217 IBIAS2.n216 16.2227
R14267 IBIAS2.n218 IBIAS2.n217 16.2227
R14268 IBIAS2.n219 IBIAS2.n218 16.2227
R14269 IBIAS2.n220 IBIAS2.n219 16.2227
R14270 IBIAS2.n221 IBIAS2.n220 16.2227
R14271 IBIAS2.n232 IBIAS2.n231 16.2227
R14272 IBIAS2.n231 IBIAS2.n230 16.2227
R14273 IBIAS2.n230 IBIAS2.n229 16.2227
R14274 IBIAS2.n229 IBIAS2.n228 16.2227
R14275 IBIAS2.n228 IBIAS2.n227 16.2227
R14276 IBIAS2.n227 IBIAS2.n226 16.2227
R14277 IBIAS2.n226 IBIAS2.n225 16.2227
R14278 IBIAS2.n262 IBIAS2.n261 16.2227
R14279 IBIAS2.n263 IBIAS2.n262 16.2227
R14280 IBIAS2.n264 IBIAS2.n263 16.2227
R14281 IBIAS2.n265 IBIAS2.n264 16.2227
R14282 IBIAS2.n266 IBIAS2.n265 16.2227
R14283 IBIAS2.n267 IBIAS2.n266 16.2227
R14284 IBIAS2.n268 IBIAS2.n267 16.2227
R14285 IBIAS2.n279 IBIAS2.n278 16.2227
R14286 IBIAS2.n278 IBIAS2.n277 16.2227
R14287 IBIAS2.n277 IBIAS2.n276 16.2227
R14288 IBIAS2.n276 IBIAS2.n275 16.2227
R14289 IBIAS2.n275 IBIAS2.n274 16.2227
R14290 IBIAS2.n274 IBIAS2.n273 16.2227
R14291 IBIAS2.n273 IBIAS2.n272 16.2227
R14292 IBIAS2.n290 IBIAS2.n289 16.2227
R14293 IBIAS2.n291 IBIAS2.n290 16.2227
R14294 IBIAS2.n292 IBIAS2.n291 16.2227
R14295 IBIAS2.n293 IBIAS2.n292 16.2227
R14296 IBIAS2.n294 IBIAS2.n293 16.2227
R14297 IBIAS2.n295 IBIAS2.n294 16.2227
R14298 IBIAS2.n296 IBIAS2.n295 16.2227
R14299 IBIAS2.n307 IBIAS2.n306 16.2227
R14300 IBIAS2.n306 IBIAS2.n305 16.2227
R14301 IBIAS2.n305 IBIAS2.n304 16.2227
R14302 IBIAS2.n304 IBIAS2.n303 16.2227
R14303 IBIAS2.n303 IBIAS2.n302 16.2227
R14304 IBIAS2.n302 IBIAS2.n301 16.2227
R14305 IBIAS2.n301 IBIAS2.n300 16.2227
R14306 IBIAS2.n318 IBIAS2.n317 16.2227
R14307 IBIAS2.n319 IBIAS2.n318 16.2227
R14308 IBIAS2.n320 IBIAS2.n319 16.2227
R14309 IBIAS2.n321 IBIAS2.n320 16.2227
R14310 IBIAS2.n322 IBIAS2.n321 16.2227
R14311 IBIAS2.n323 IBIAS2.n322 16.2227
R14312 IBIAS2.n324 IBIAS2.n323 16.2227
R14313 IBIAS2.n335 IBIAS2.n334 16.2227
R14314 IBIAS2.n334 IBIAS2.n333 16.2227
R14315 IBIAS2.n333 IBIAS2.n332 16.2227
R14316 IBIAS2.n332 IBIAS2.n331 16.2227
R14317 IBIAS2.n331 IBIAS2.n330 16.2227
R14318 IBIAS2.n330 IBIAS2.n329 16.2227
R14319 IBIAS2.n329 IBIAS2.n328 16.2227
R14320 IBIAS2.n365 IBIAS2.n364 16.2227
R14321 IBIAS2.n366 IBIAS2.n365 16.2227
R14322 IBIAS2.n367 IBIAS2.n366 16.2227
R14323 IBIAS2.n368 IBIAS2.n367 16.2227
R14324 IBIAS2.n369 IBIAS2.n368 16.2227
R14325 IBIAS2.n370 IBIAS2.n369 16.2227
R14326 IBIAS2.n371 IBIAS2.n370 16.2227
R14327 IBIAS2.n382 IBIAS2.n381 16.2227
R14328 IBIAS2.n381 IBIAS2.n380 16.2227
R14329 IBIAS2.n380 IBIAS2.n379 16.2227
R14330 IBIAS2.n379 IBIAS2.n378 16.2227
R14331 IBIAS2.n378 IBIAS2.n377 16.2227
R14332 IBIAS2.n377 IBIAS2.n376 16.2227
R14333 IBIAS2.n376 IBIAS2.n375 16.2227
R14334 IBIAS2.n393 IBIAS2.n392 16.2227
R14335 IBIAS2.n394 IBIAS2.n393 16.2227
R14336 IBIAS2.n395 IBIAS2.n394 16.2227
R14337 IBIAS2.n396 IBIAS2.n395 16.2227
R14338 IBIAS2.n397 IBIAS2.n396 16.2227
R14339 IBIAS2.n398 IBIAS2.n397 16.2227
R14340 IBIAS2.n399 IBIAS2.n398 16.2227
R14341 IBIAS2.n410 IBIAS2.n409 16.2227
R14342 IBIAS2.n409 IBIAS2.n408 16.2227
R14343 IBIAS2.n408 IBIAS2.n407 16.2227
R14344 IBIAS2.n407 IBIAS2.n406 16.2227
R14345 IBIAS2.n406 IBIAS2.n405 16.2227
R14346 IBIAS2.n405 IBIAS2.n404 16.2227
R14347 IBIAS2.n404 IBIAS2.n403 16.2227
R14348 IBIAS2.n421 IBIAS2.n420 16.2227
R14349 IBIAS2.n422 IBIAS2.n421 16.2227
R14350 IBIAS2.n423 IBIAS2.n422 16.2227
R14351 IBIAS2.n424 IBIAS2.n423 16.2227
R14352 IBIAS2.n425 IBIAS2.n424 16.2227
R14353 IBIAS2.n426 IBIAS2.n425 16.2227
R14354 IBIAS2.n427 IBIAS2.n426 16.2227
R14355 IBIAS2.n438 IBIAS2.n437 16.2227
R14356 IBIAS2.n437 IBIAS2.n436 16.2227
R14357 IBIAS2.n436 IBIAS2.n435 16.2227
R14358 IBIAS2.n435 IBIAS2.n434 16.2227
R14359 IBIAS2.n434 IBIAS2.n433 16.2227
R14360 IBIAS2.n433 IBIAS2.n432 16.2227
R14361 IBIAS2.n432 IBIAS2.n431 16.2227
R14362 IBIAS2.n468 IBIAS2.n467 16.2227
R14363 IBIAS2.n469 IBIAS2.n468 16.2227
R14364 IBIAS2.n470 IBIAS2.n469 16.2227
R14365 IBIAS2.n471 IBIAS2.n470 16.2227
R14366 IBIAS2.n472 IBIAS2.n471 16.2227
R14367 IBIAS2.n473 IBIAS2.n472 16.2227
R14368 IBIAS2.n474 IBIAS2.n473 16.2227
R14369 IBIAS2.n485 IBIAS2.n484 16.2227
R14370 IBIAS2.n484 IBIAS2.n483 16.2227
R14371 IBIAS2.n483 IBIAS2.n482 16.2227
R14372 IBIAS2.n482 IBIAS2.n481 16.2227
R14373 IBIAS2.n481 IBIAS2.n480 16.2227
R14374 IBIAS2.n480 IBIAS2.n479 16.2227
R14375 IBIAS2.n479 IBIAS2.n478 16.2227
R14376 IBIAS2.n496 IBIAS2.n495 16.2227
R14377 IBIAS2.n497 IBIAS2.n496 16.2227
R14378 IBIAS2.n498 IBIAS2.n497 16.2227
R14379 IBIAS2.n499 IBIAS2.n498 16.2227
R14380 IBIAS2.n500 IBIAS2.n499 16.2227
R14381 IBIAS2.n501 IBIAS2.n500 16.2227
R14382 IBIAS2.n502 IBIAS2.n501 16.2227
R14383 IBIAS2.n513 IBIAS2.n512 16.2227
R14384 IBIAS2.n512 IBIAS2.n511 16.2227
R14385 IBIAS2.n511 IBIAS2.n510 16.2227
R14386 IBIAS2.n510 IBIAS2.n509 16.2227
R14387 IBIAS2.n509 IBIAS2.n508 16.2227
R14388 IBIAS2.n508 IBIAS2.n507 16.2227
R14389 IBIAS2.n507 IBIAS2.n506 16.2227
R14390 IBIAS2.n524 IBIAS2.n523 16.2227
R14391 IBIAS2.n525 IBIAS2.n524 16.2227
R14392 IBIAS2.n526 IBIAS2.n525 16.2227
R14393 IBIAS2.n527 IBIAS2.n526 16.2227
R14394 IBIAS2.n528 IBIAS2.n527 16.2227
R14395 IBIAS2.n529 IBIAS2.n528 16.2227
R14396 IBIAS2.n530 IBIAS2.n529 16.2227
R14397 IBIAS2.n541 IBIAS2.n540 16.2227
R14398 IBIAS2.n540 IBIAS2.n539 16.2227
R14399 IBIAS2.n539 IBIAS2.n538 16.2227
R14400 IBIAS2.n538 IBIAS2.n537 16.2227
R14401 IBIAS2.n537 IBIAS2.n536 16.2227
R14402 IBIAS2.n536 IBIAS2.n535 16.2227
R14403 IBIAS2.n535 IBIAS2.n534 16.2227
R14404 IBIAS2.n571 IBIAS2.n570 16.2227
R14405 IBIAS2.n572 IBIAS2.n571 16.2227
R14406 IBIAS2.n573 IBIAS2.n572 16.2227
R14407 IBIAS2.n574 IBIAS2.n573 16.2227
R14408 IBIAS2.n575 IBIAS2.n574 16.2227
R14409 IBIAS2.n576 IBIAS2.n575 16.2227
R14410 IBIAS2.n577 IBIAS2.n576 16.2227
R14411 IBIAS2.n588 IBIAS2.n587 16.2227
R14412 IBIAS2.n587 IBIAS2.n586 16.2227
R14413 IBIAS2.n586 IBIAS2.n585 16.2227
R14414 IBIAS2.n585 IBIAS2.n584 16.2227
R14415 IBIAS2.n584 IBIAS2.n583 16.2227
R14416 IBIAS2.n583 IBIAS2.n582 16.2227
R14417 IBIAS2.n582 IBIAS2.n581 16.2227
R14418 IBIAS2.n599 IBIAS2.n598 16.2227
R14419 IBIAS2.n600 IBIAS2.n599 16.2227
R14420 IBIAS2.n601 IBIAS2.n600 16.2227
R14421 IBIAS2.n602 IBIAS2.n601 16.2227
R14422 IBIAS2.n603 IBIAS2.n602 16.2227
R14423 IBIAS2.n604 IBIAS2.n603 16.2227
R14424 IBIAS2.n605 IBIAS2.n604 16.2227
R14425 IBIAS2.n616 IBIAS2.n615 16.2227
R14426 IBIAS2.n615 IBIAS2.n614 16.2227
R14427 IBIAS2.n614 IBIAS2.n613 16.2227
R14428 IBIAS2.n613 IBIAS2.n612 16.2227
R14429 IBIAS2.n612 IBIAS2.n611 16.2227
R14430 IBIAS2.n611 IBIAS2.n610 16.2227
R14431 IBIAS2.n610 IBIAS2.n609 16.2227
R14432 IBIAS2.n627 IBIAS2.n626 16.2227
R14433 IBIAS2.n628 IBIAS2.n627 16.2227
R14434 IBIAS2.n629 IBIAS2.n628 16.2227
R14435 IBIAS2.n630 IBIAS2.n629 16.2227
R14436 IBIAS2.n631 IBIAS2.n630 16.2227
R14437 IBIAS2.n632 IBIAS2.n631 16.2227
R14438 IBIAS2.n633 IBIAS2.n632 16.2227
R14439 IBIAS2.n644 IBIAS2.n643 16.2227
R14440 IBIAS2.n643 IBIAS2.n642 16.2227
R14441 IBIAS2.n642 IBIAS2.n641 16.2227
R14442 IBIAS2.n641 IBIAS2.n640 16.2227
R14443 IBIAS2.n640 IBIAS2.n639 16.2227
R14444 IBIAS2.n639 IBIAS2.n638 16.2227
R14445 IBIAS2.n638 IBIAS2.n637 16.2227
R14446 IBIAS2.n674 IBIAS2.n673 16.2227
R14447 IBIAS2.n675 IBIAS2.n674 16.2227
R14448 IBIAS2.n676 IBIAS2.n675 16.2227
R14449 IBIAS2.n677 IBIAS2.n676 16.2227
R14450 IBIAS2.n678 IBIAS2.n677 16.2227
R14451 IBIAS2.n679 IBIAS2.n678 16.2227
R14452 IBIAS2.n680 IBIAS2.n679 16.2227
R14453 IBIAS2.n691 IBIAS2.n690 16.2227
R14454 IBIAS2.n690 IBIAS2.n689 16.2227
R14455 IBIAS2.n689 IBIAS2.n688 16.2227
R14456 IBIAS2.n688 IBIAS2.n687 16.2227
R14457 IBIAS2.n687 IBIAS2.n686 16.2227
R14458 IBIAS2.n686 IBIAS2.n685 16.2227
R14459 IBIAS2.n685 IBIAS2.n684 16.2227
R14460 IBIAS2.n702 IBIAS2.n701 16.2227
R14461 IBIAS2.n703 IBIAS2.n702 16.2227
R14462 IBIAS2.n704 IBIAS2.n703 16.2227
R14463 IBIAS2.n705 IBIAS2.n704 16.2227
R14464 IBIAS2.n706 IBIAS2.n705 16.2227
R14465 IBIAS2.n707 IBIAS2.n706 16.2227
R14466 IBIAS2.n708 IBIAS2.n707 16.2227
R14467 IBIAS2.n719 IBIAS2.n718 16.2227
R14468 IBIAS2.n718 IBIAS2.n717 16.2227
R14469 IBIAS2.n717 IBIAS2.n716 16.2227
R14470 IBIAS2.n716 IBIAS2.n715 16.2227
R14471 IBIAS2.n715 IBIAS2.n714 16.2227
R14472 IBIAS2.n714 IBIAS2.n713 16.2227
R14473 IBIAS2.n713 IBIAS2.n712 16.2227
R14474 IBIAS2.n730 IBIAS2.n729 16.2227
R14475 IBIAS2.n731 IBIAS2.n730 16.2227
R14476 IBIAS2.n732 IBIAS2.n731 16.2227
R14477 IBIAS2.n733 IBIAS2.n732 16.2227
R14478 IBIAS2.n734 IBIAS2.n733 16.2227
R14479 IBIAS2.n735 IBIAS2.n734 16.2227
R14480 IBIAS2.n736 IBIAS2.n735 16.2227
R14481 IBIAS2.n747 IBIAS2.n746 16.2227
R14482 IBIAS2.n746 IBIAS2.n745 16.2227
R14483 IBIAS2.n745 IBIAS2.n744 16.2227
R14484 IBIAS2.n744 IBIAS2.n743 16.2227
R14485 IBIAS2.n743 IBIAS2.n742 16.2227
R14486 IBIAS2.n742 IBIAS2.n741 16.2227
R14487 IBIAS2.n741 IBIAS2.n740 16.2227
R14488 IBIAS2.n21 IBIAS2.n20 16.2227
R14489 IBIAS2.n22 IBIAS2.n21 16.2227
R14490 IBIAS2.n23 IBIAS2.n22 16.2227
R14491 IBIAS2.n24 IBIAS2.n23 16.2227
R14492 IBIAS2.n25 IBIAS2.n24 16.2227
R14493 IBIAS2.n26 IBIAS2.n25 16.2227
R14494 IBIAS2.n27 IBIAS2.n26 16.2227
R14495 IBIAS2.n38 IBIAS2.n37 16.2227
R14496 IBIAS2.n37 IBIAS2.n36 16.2227
R14497 IBIAS2.n36 IBIAS2.n35 16.2227
R14498 IBIAS2.n35 IBIAS2.n34 16.2227
R14499 IBIAS2.n34 IBIAS2.n33 16.2227
R14500 IBIAS2.n33 IBIAS2.n32 16.2227
R14501 IBIAS2.n32 IBIAS2.n31 16.2227
R14502 IBIAS2.n90 IBIAS2.n89 16.2227
R14503 IBIAS2.n91 IBIAS2.n90 16.2227
R14504 IBIAS2.n92 IBIAS2.n91 16.2227
R14505 IBIAS2.n93 IBIAS2.n92 16.2227
R14506 IBIAS2.n94 IBIAS2.n93 16.2227
R14507 IBIAS2.n95 IBIAS2.n94 16.2227
R14508 IBIAS2.n96 IBIAS2.n95 16.2227
R14509 IBIAS2.n107 IBIAS2.n106 16.2227
R14510 IBIAS2.n106 IBIAS2.n105 16.2227
R14511 IBIAS2.n105 IBIAS2.n104 16.2227
R14512 IBIAS2.n104 IBIAS2.n103 16.2227
R14513 IBIAS2.n103 IBIAS2.n102 16.2227
R14514 IBIAS2.n102 IBIAS2.n101 16.2227
R14515 IBIAS2.n101 IBIAS2.n100 16.2227
R14516 IBIAS2.n117 IBIAS2.n116 16.2227
R14517 IBIAS2.n118 IBIAS2.n117 16.2227
R14518 IBIAS2.n119 IBIAS2.n118 16.2227
R14519 IBIAS2.n120 IBIAS2.n119 16.2227
R14520 IBIAS2.n121 IBIAS2.n120 16.2227
R14521 IBIAS2.n122 IBIAS2.n121 16.2227
R14522 IBIAS2.n123 IBIAS2.n122 16.2227
R14523 IBIAS2.n134 IBIAS2.n133 16.2227
R14524 IBIAS2.n133 IBIAS2.n132 16.2227
R14525 IBIAS2.n132 IBIAS2.n131 16.2227
R14526 IBIAS2.n131 IBIAS2.n130 16.2227
R14527 IBIAS2.n130 IBIAS2.n129 16.2227
R14528 IBIAS2.n129 IBIAS2.n128 16.2227
R14529 IBIAS2.n128 IBIAS2.n127 16.2227
R14530 IBIAS2.n82 IBIAS2.n81 11.6793
R14531 IBIAS2.n44 IBIAS2.t117 4.65943
R14532 IBIAS2.n56 IBIAS2.n55 3.86296
R14533 IBIAS2.n71 IBIAS2.n70 3.86296
R14534 IBIAS2.n235 IBIAS2.n224 3.30289
R14535 IBIAS2.n207 IBIAS2.n196 3.30289
R14536 IBIAS2.n179 IBIAS2.n168 3.30289
R14537 IBIAS2.n154 IBIAS2.n151 3.30289
R14538 IBIAS2.n338 IBIAS2.n327 3.30289
R14539 IBIAS2.n310 IBIAS2.n299 3.30289
R14540 IBIAS2.n282 IBIAS2.n271 3.30289
R14541 IBIAS2.n257 IBIAS2.n254 3.30289
R14542 IBIAS2.n441 IBIAS2.n430 3.30289
R14543 IBIAS2.n413 IBIAS2.n402 3.30289
R14544 IBIAS2.n385 IBIAS2.n374 3.30289
R14545 IBIAS2.n360 IBIAS2.n357 3.30289
R14546 IBIAS2.n544 IBIAS2.n533 3.30289
R14547 IBIAS2.n516 IBIAS2.n505 3.30289
R14548 IBIAS2.n488 IBIAS2.n477 3.30289
R14549 IBIAS2.n463 IBIAS2.n460 3.30289
R14550 IBIAS2.n647 IBIAS2.n636 3.30289
R14551 IBIAS2.n619 IBIAS2.n608 3.30289
R14552 IBIAS2.n591 IBIAS2.n580 3.30289
R14553 IBIAS2.n566 IBIAS2.n563 3.30289
R14554 IBIAS2.n750 IBIAS2.n739 3.30289
R14555 IBIAS2.n722 IBIAS2.n711 3.30289
R14556 IBIAS2.n694 IBIAS2.n683 3.30289
R14557 IBIAS2.n669 IBIAS2.n666 3.30289
R14558 IBIAS2.n126 IBIAS2.n115 3.30289
R14559 IBIAS2.n99 IBIAS2.n88 3.30289
R14560 IBIAS2.n30 IBIAS2.n19 3.30289
R14561 IBIAS2.n15 IBIAS2.n14 3.30289
R14562 IBIAS2.n166 IBIAS2.n165 2.8805
R14563 IBIAS2.n194 IBIAS2.n193 2.8805
R14564 IBIAS2.n222 IBIAS2.n221 2.8805
R14565 IBIAS2.n205 IBIAS2.n204 2.8805
R14566 IBIAS2.n233 IBIAS2.n232 2.8805
R14567 IBIAS2.n177 IBIAS2.n176 2.8805
R14568 IBIAS2.n269 IBIAS2.n268 2.8805
R14569 IBIAS2.n297 IBIAS2.n296 2.8805
R14570 IBIAS2.n325 IBIAS2.n324 2.8805
R14571 IBIAS2.n308 IBIAS2.n307 2.8805
R14572 IBIAS2.n336 IBIAS2.n335 2.8805
R14573 IBIAS2.n280 IBIAS2.n279 2.8805
R14574 IBIAS2.n372 IBIAS2.n371 2.8805
R14575 IBIAS2.n400 IBIAS2.n399 2.8805
R14576 IBIAS2.n428 IBIAS2.n427 2.8805
R14577 IBIAS2.n411 IBIAS2.n410 2.8805
R14578 IBIAS2.n439 IBIAS2.n438 2.8805
R14579 IBIAS2.n383 IBIAS2.n382 2.8805
R14580 IBIAS2.n475 IBIAS2.n474 2.8805
R14581 IBIAS2.n503 IBIAS2.n502 2.8805
R14582 IBIAS2.n531 IBIAS2.n530 2.8805
R14583 IBIAS2.n514 IBIAS2.n513 2.8805
R14584 IBIAS2.n542 IBIAS2.n541 2.8805
R14585 IBIAS2.n486 IBIAS2.n485 2.8805
R14586 IBIAS2.n578 IBIAS2.n577 2.8805
R14587 IBIAS2.n606 IBIAS2.n605 2.8805
R14588 IBIAS2.n634 IBIAS2.n633 2.8805
R14589 IBIAS2.n617 IBIAS2.n616 2.8805
R14590 IBIAS2.n645 IBIAS2.n644 2.8805
R14591 IBIAS2.n589 IBIAS2.n588 2.8805
R14592 IBIAS2.n681 IBIAS2.n680 2.8805
R14593 IBIAS2.n709 IBIAS2.n708 2.8805
R14594 IBIAS2.n737 IBIAS2.n736 2.8805
R14595 IBIAS2.n720 IBIAS2.n719 2.8805
R14596 IBIAS2.n748 IBIAS2.n747 2.8805
R14597 IBIAS2.n692 IBIAS2.n691 2.8805
R14598 IBIAS2.n39 IBIAS2.n38 2.8805
R14599 IBIAS2.n108 IBIAS2.n107 2.8805
R14600 IBIAS2.n135 IBIAS2.n134 2.8805
R14601 IBIAS2.n124 IBIAS2.n123 2.8805
R14602 IBIAS2.n97 IBIAS2.n96 2.8805
R14603 IBIAS2.n28 IBIAS2.n27 2.8805
R14604 IBIAS2.n661 IBIAS2.n660 1.69656
R14605 IBIAS2.n455 IBIAS2.n454 1.69656
R14606 IBIAS2.n249 IBIAS2.n248 1.69656
R14607 IBIAS2.n61 IBIAS2.n60 1.44217
R14608 IBIAS2.n76 IBIAS2.n75 1.44217
R14609 IBIAS2.n558 IBIAS2.n557 1.24529
R14610 IBIAS2.n352 IBIAS2.n351 1.24529
R14611 IBIAS2.n146 IBIAS2.n145 1.24529
R14612 IBIAS2.n43 IBIAS2.n42 1.16617
R14613 IBIAS2.n62 IBIAS2.n61 1.14036
R14614 IBIAS2.n77 IBIAS2.n76 1.14036
R14615 IBIAS2.n46 IBIAS2.n45 1.1255
R14616 IBIAS2.n58 IBIAS2.n57 1.1255
R14617 IBIAS2.n73 IBIAS2.n72 1.1255
R14618 IBIAS2.n237 IBIAS2.n236 1.1228
R14619 IBIAS2.n209 IBIAS2.n208 1.1228
R14620 IBIAS2.n181 IBIAS2.n180 1.1228
R14621 IBIAS2.n340 IBIAS2.n339 1.1228
R14622 IBIAS2.n312 IBIAS2.n311 1.1228
R14623 IBIAS2.n284 IBIAS2.n283 1.1228
R14624 IBIAS2.n443 IBIAS2.n442 1.1228
R14625 IBIAS2.n415 IBIAS2.n414 1.1228
R14626 IBIAS2.n387 IBIAS2.n386 1.1228
R14627 IBIAS2.n546 IBIAS2.n545 1.1228
R14628 IBIAS2.n518 IBIAS2.n517 1.1228
R14629 IBIAS2.n490 IBIAS2.n489 1.1228
R14630 IBIAS2.n649 IBIAS2.n648 1.1228
R14631 IBIAS2.n621 IBIAS2.n620 1.1228
R14632 IBIAS2.n593 IBIAS2.n592 1.1228
R14633 IBIAS2.n752 IBIAS2.n751 1.1228
R14634 IBIAS2.n724 IBIAS2.n723 1.1228
R14635 IBIAS2.n696 IBIAS2.n695 1.1228
R14636 IBIAS2.n241 IBIAS2.n156 1.12272
R14637 IBIAS2.n344 IBIAS2.n259 1.12272
R14638 IBIAS2.n447 IBIAS2.n362 1.12272
R14639 IBIAS2.n550 IBIAS2.n465 1.12272
R14640 IBIAS2.n653 IBIAS2.n568 1.12272
R14641 IBIAS2.n756 IBIAS2.n671 1.12272
R14642 IBIAS2.n137 IBIAS2.n136 1.12272
R14643 IBIAS2.n110 IBIAS2.n109 1.12272
R14644 IBIAS2.n83 IBIAS2.n40 1.12272
R14645 IBIAS2.n141 IBIAS2.n17 1.12272
R14646 IBIAS2.n141 IBIAS2.n12 1.12243
R14647 IBIAS2.n248 IBIAS2.n247 1.11801
R14648 IBIAS2.n763 IBIAS2.n762 1.11801
R14649 IBIAS2.n660 IBIAS2.n659 1.11801
R14650 IBIAS2.n557 IBIAS2.n556 1.11801
R14651 IBIAS2.n454 IBIAS2.n453 1.11801
R14652 IBIAS2.n351 IBIAS2.n350 1.11801
R14653 IBIAS2.n144 IBIAS2.n143 1.11782
R14654 IBIAS2.n760 IBIAS2.n759 1.11782
R14655 IBIAS2.n657 IBIAS2.n656 1.11782
R14656 IBIAS2.n554 IBIAS2.n553 1.11782
R14657 IBIAS2.n451 IBIAS2.n450 1.11782
R14658 IBIAS2.n348 IBIAS2.n347 1.11782
R14659 IBIAS2.n245 IBIAS2.n244 1.11782
R14660 IBIAS2.n42 IBIAS2.n41 1.07327
R14661 IBIAS2.n764 IBIAS2.n763 0.962646
R14662 IBIAS2.n41 IBIAS2.t121 0.8195
R14663 IBIAS2.n60 IBIAS2.t118 0.8195
R14664 IBIAS2.n60 IBIAS2.n59 0.8195
R14665 IBIAS2.n55 IBIAS2.t115 0.8195
R14666 IBIAS2.n55 IBIAS2.n54 0.8195
R14667 IBIAS2.n75 IBIAS2.t116 0.8195
R14668 IBIAS2.n75 IBIAS2.n74 0.8195
R14669 IBIAS2.n70 IBIAS2.t112 0.8195
R14670 IBIAS2.n70 IBIAS2.n69 0.8195
R14671 IBIAS2.n768 IBIAS2.n767 0.767554
R14672 IBIAS2.n4 IBIAS2.n3 0.7505
R14673 IBIAS2.n64 IBIAS2.n63 0.727916
R14674 IBIAS2.n79 IBIAS2.n78 0.727916
R14675 IBIAS2.n49 IBIAS2.n47 0.616779
R14676 IBIAS2.n224 IBIAS2.t75 0.607167
R14677 IBIAS2.n224 IBIAS2.n223 0.607167
R14678 IBIAS2.n196 IBIAS2.t111 0.607167
R14679 IBIAS2.n196 IBIAS2.n195 0.607167
R14680 IBIAS2.n168 IBIAS2.t41 0.607167
R14681 IBIAS2.n168 IBIAS2.n167 0.607167
R14682 IBIAS2.n151 IBIAS2.t89 0.607167
R14683 IBIAS2.n151 IBIAS2.n150 0.607167
R14684 IBIAS2.n327 IBIAS2.t67 0.607167
R14685 IBIAS2.n327 IBIAS2.n326 0.607167
R14686 IBIAS2.n299 IBIAS2.t63 0.607167
R14687 IBIAS2.n299 IBIAS2.n298 0.607167
R14688 IBIAS2.n271 IBIAS2.t109 0.607167
R14689 IBIAS2.n271 IBIAS2.n270 0.607167
R14690 IBIAS2.n254 IBIAS2.t33 0.607167
R14691 IBIAS2.n254 IBIAS2.n253 0.607167
R14692 IBIAS2.n430 IBIAS2.t61 0.607167
R14693 IBIAS2.n430 IBIAS2.n429 0.607167
R14694 IBIAS2.n402 IBIAS2.t57 0.607167
R14695 IBIAS2.n402 IBIAS2.n401 0.607167
R14696 IBIAS2.n374 IBIAS2.t47 0.607167
R14697 IBIAS2.n374 IBIAS2.n373 0.607167
R14698 IBIAS2.n357 IBIAS2.t25 0.607167
R14699 IBIAS2.n357 IBIAS2.n356 0.607167
R14700 IBIAS2.n533 IBIAS2.t45 0.607167
R14701 IBIAS2.n533 IBIAS2.n532 0.607167
R14702 IBIAS2.n505 IBIAS2.t9 0.607167
R14703 IBIAS2.n505 IBIAS2.n504 0.607167
R14704 IBIAS2.n477 IBIAS2.t1 0.607167
R14705 IBIAS2.n477 IBIAS2.n476 0.607167
R14706 IBIAS2.n460 IBIAS2.t99 0.607167
R14707 IBIAS2.n460 IBIAS2.n459 0.607167
R14708 IBIAS2.n636 IBIAS2.t21 0.607167
R14709 IBIAS2.n636 IBIAS2.n635 0.607167
R14710 IBIAS2.n608 IBIAS2.t13 0.607167
R14711 IBIAS2.n608 IBIAS2.n607 0.607167
R14712 IBIAS2.n580 IBIAS2.t77 0.607167
R14713 IBIAS2.n580 IBIAS2.n579 0.607167
R14714 IBIAS2.n563 IBIAS2.t101 0.607167
R14715 IBIAS2.n563 IBIAS2.n562 0.607167
R14716 IBIAS2.n739 IBIAS2.t35 0.607167
R14717 IBIAS2.n739 IBIAS2.n738 0.607167
R14718 IBIAS2.n711 IBIAS2.t37 0.607167
R14719 IBIAS2.n711 IBIAS2.n710 0.607167
R14720 IBIAS2.n683 IBIAS2.t39 0.607167
R14721 IBIAS2.n683 IBIAS2.n682 0.607167
R14722 IBIAS2.n666 IBIAS2.t17 0.607167
R14723 IBIAS2.n666 IBIAS2.n665 0.607167
R14724 IBIAS2.n115 IBIAS2.t105 0.607167
R14725 IBIAS2.n115 IBIAS2.n114 0.607167
R14726 IBIAS2.n88 IBIAS2.t107 0.607167
R14727 IBIAS2.n88 IBIAS2.n87 0.607167
R14728 IBIAS2.n19 IBIAS2.t91 0.607167
R14729 IBIAS2.n19 IBIAS2.n18 0.607167
R14730 IBIAS2.n14 IBIAS2.t85 0.607167
R14731 IBIAS2.n14 IBIAS2.n13 0.607167
R14732 IBIAS2.n240 IBIAS2.n239 0.386051
R14733 IBIAS2.n212 IBIAS2.n211 0.386051
R14734 IBIAS2.n184 IBIAS2.n183 0.386051
R14735 IBIAS2.n343 IBIAS2.n342 0.386051
R14736 IBIAS2.n315 IBIAS2.n314 0.386051
R14737 IBIAS2.n287 IBIAS2.n286 0.386051
R14738 IBIAS2.n446 IBIAS2.n445 0.386051
R14739 IBIAS2.n418 IBIAS2.n417 0.386051
R14740 IBIAS2.n390 IBIAS2.n389 0.386051
R14741 IBIAS2.n549 IBIAS2.n548 0.386051
R14742 IBIAS2.n521 IBIAS2.n520 0.386051
R14743 IBIAS2.n493 IBIAS2.n492 0.386051
R14744 IBIAS2.n652 IBIAS2.n651 0.386051
R14745 IBIAS2.n624 IBIAS2.n623 0.386051
R14746 IBIAS2.n596 IBIAS2.n595 0.386051
R14747 IBIAS2.n755 IBIAS2.n754 0.386051
R14748 IBIAS2.n727 IBIAS2.n726 0.386051
R14749 IBIAS2.n699 IBIAS2.n698 0.386051
R14750 IBIAS2.n140 IBIAS2.n139 0.386051
R14751 IBIAS2.n113 IBIAS2.n112 0.386051
R14752 IBIAS2.n86 IBIAS2.n85 0.386051
R14753 IBIAS2.n244 IBIAS2.n243 0.380932
R14754 IBIAS2.n347 IBIAS2.n346 0.380932
R14755 IBIAS2.n450 IBIAS2.n449 0.380932
R14756 IBIAS2.n553 IBIAS2.n552 0.380932
R14757 IBIAS2.n656 IBIAS2.n655 0.380932
R14758 IBIAS2.n759 IBIAS2.n758 0.380932
R14759 IBIAS2.n143 IBIAS2.n142 0.380932
R14760 IBIAS2.n67 IBIAS2.n66 0.2775
R14761 IBIAS2.n52 IBIAS2.n51 0.2775
R14762 IBIAS2.n767 IBIAS2.n766 0.147906
R14763 IBIAS2.n156 IBIAS2.n154 0.101374
R14764 IBIAS2.n259 IBIAS2.n257 0.101374
R14765 IBIAS2.n362 IBIAS2.n360 0.101374
R14766 IBIAS2.n465 IBIAS2.n463 0.101374
R14767 IBIAS2.n568 IBIAS2.n566 0.101374
R14768 IBIAS2.n671 IBIAS2.n669 0.101374
R14769 IBIAS2.n136 IBIAS2.n126 0.101374
R14770 IBIAS2.n109 IBIAS2.n99 0.101374
R14771 IBIAS2.n40 IBIAS2.n30 0.101374
R14772 IBIAS2.n17 IBIAS2.n15 0.101374
R14773 IBIAS2.n236 IBIAS2.n235 0.100442
R14774 IBIAS2.n208 IBIAS2.n207 0.100442
R14775 IBIAS2.n180 IBIAS2.n179 0.100442
R14776 IBIAS2.n339 IBIAS2.n338 0.100442
R14777 IBIAS2.n311 IBIAS2.n310 0.100442
R14778 IBIAS2.n283 IBIAS2.n282 0.100442
R14779 IBIAS2.n442 IBIAS2.n441 0.100442
R14780 IBIAS2.n414 IBIAS2.n413 0.100442
R14781 IBIAS2.n386 IBIAS2.n385 0.100442
R14782 IBIAS2.n545 IBIAS2.n544 0.100442
R14783 IBIAS2.n517 IBIAS2.n516 0.100442
R14784 IBIAS2.n489 IBIAS2.n488 0.100442
R14785 IBIAS2.n648 IBIAS2.n647 0.100442
R14786 IBIAS2.n620 IBIAS2.n619 0.100442
R14787 IBIAS2.n592 IBIAS2.n591 0.100442
R14788 IBIAS2.n751 IBIAS2.n750 0.100442
R14789 IBIAS2.n723 IBIAS2.n722 0.100442
R14790 IBIAS2.n695 IBIAS2.n694 0.100442
R14791 IBIAS2.n154 IBIAS2.n153 0.0986789
R14792 IBIAS2.n257 IBIAS2.n256 0.0986789
R14793 IBIAS2.n360 IBIAS2.n359 0.0986789
R14794 IBIAS2.n463 IBIAS2.n462 0.0986789
R14795 IBIAS2.n566 IBIAS2.n565 0.0986789
R14796 IBIAS2.n669 IBIAS2.n668 0.0986789
R14797 IBIAS2.n99 IBIAS2.n98 0.0986789
R14798 IBIAS2.n126 IBIAS2.n125 0.0986789
R14799 IBIAS2.n30 IBIAS2.n29 0.0986789
R14800 IBIAS2.n235 IBIAS2.n234 0.0937119
R14801 IBIAS2.n207 IBIAS2.n206 0.0937119
R14802 IBIAS2.n179 IBIAS2.n178 0.0937119
R14803 IBIAS2.n338 IBIAS2.n337 0.0937119
R14804 IBIAS2.n310 IBIAS2.n309 0.0937119
R14805 IBIAS2.n282 IBIAS2.n281 0.0937119
R14806 IBIAS2.n441 IBIAS2.n440 0.0937119
R14807 IBIAS2.n413 IBIAS2.n412 0.0937119
R14808 IBIAS2.n385 IBIAS2.n384 0.0937119
R14809 IBIAS2.n544 IBIAS2.n543 0.0937119
R14810 IBIAS2.n516 IBIAS2.n515 0.0937119
R14811 IBIAS2.n488 IBIAS2.n487 0.0937119
R14812 IBIAS2.n647 IBIAS2.n646 0.0937119
R14813 IBIAS2.n619 IBIAS2.n618 0.0937119
R14814 IBIAS2.n591 IBIAS2.n590 0.0937119
R14815 IBIAS2.n750 IBIAS2.n749 0.0937119
R14816 IBIAS2.n722 IBIAS2.n721 0.0937119
R14817 IBIAS2.n694 IBIAS2.n693 0.0937119
R14818 IBIAS2.n63 IBIAS2.n62 0.0826464
R14819 IBIAS2.n78 IBIAS2.n77 0.0826464
R14820 IBIAS2 IBIAS2.n768 0.0822606
R14821 IBIAS2.n47 IBIAS2.n43 0.0712285
R14822 IBIAS2.n47 IBIAS2.n46 0.0534597
R14823 IBIAS2.n63 IBIAS2.n58 0.0423164
R14824 IBIAS2.n78 IBIAS2.n73 0.0423164
R14825 IBIAS2.n45 IBIAS2.n44 0.0383947
R14826 IBIAS2.n768 IBIAS2.n4 0.0334577
R14827 IBIAS2.n6 IBIAS2.n5 0.0235313
R14828 IBIAS2.n8 IBIAS2.n7 0.0228651
R14829 IBIAS2.n143 IBIAS2.n10 0.0179841
R14830 IBIAS2.n759 IBIAS2.n664 0.0179841
R14831 IBIAS2.n656 IBIAS2.n561 0.0179841
R14832 IBIAS2.n553 IBIAS2.n458 0.0179841
R14833 IBIAS2.n450 IBIAS2.n355 0.0179841
R14834 IBIAS2.n347 IBIAS2.n252 0.0179841
R14835 IBIAS2.n244 IBIAS2.n149 0.0179841
R14836 IBIAS2.n762 IBIAS2.n761 0.0179841
R14837 IBIAS2.n663 IBIAS2.n662 0.0179841
R14838 IBIAS2.n659 IBIAS2.n658 0.0179841
R14839 IBIAS2.n560 IBIAS2.n559 0.0179841
R14840 IBIAS2.n556 IBIAS2.n555 0.0179841
R14841 IBIAS2.n457 IBIAS2.n456 0.0179841
R14842 IBIAS2.n453 IBIAS2.n452 0.0179841
R14843 IBIAS2.n354 IBIAS2.n353 0.0179841
R14844 IBIAS2.n350 IBIAS2.n349 0.0179841
R14845 IBIAS2.n251 IBIAS2.n250 0.0179841
R14846 IBIAS2.n247 IBIAS2.n246 0.0179841
R14847 IBIAS2.n148 IBIAS2.n147 0.0179841
R14848 IBIAS2.n10 IBIAS2.n9 0.0177304
R14849 IBIAS2.n662 IBIAS2.n661 0.0177304
R14850 IBIAS2.n559 IBIAS2.n558 0.0177304
R14851 IBIAS2.n456 IBIAS2.n455 0.0177304
R14852 IBIAS2.n353 IBIAS2.n352 0.0177304
R14853 IBIAS2.n250 IBIAS2.n249 0.0177304
R14854 IBIAS2.n147 IBIAS2.n146 0.0177304
R14855 IBIAS2.n760 IBIAS2.n663 0.0173591
R14856 IBIAS2.n657 IBIAS2.n560 0.0173591
R14857 IBIAS2.n554 IBIAS2.n457 0.0173591
R14858 IBIAS2.n451 IBIAS2.n354 0.0173591
R14859 IBIAS2.n348 IBIAS2.n251 0.0173591
R14860 IBIAS2.n245 IBIAS2.n148 0.0173591
R14861 IBIAS2.n144 IBIAS2.n6 0.0173591
R14862 IBIAS2.n145 IBIAS2.n144 0.0173591
R14863 IBIAS2.n763 IBIAS2.n760 0.0173591
R14864 IBIAS2.n660 IBIAS2.n657 0.0173591
R14865 IBIAS2.n557 IBIAS2.n554 0.0173591
R14866 IBIAS2.n454 IBIAS2.n451 0.0173591
R14867 IBIAS2.n351 IBIAS2.n348 0.0173591
R14868 IBIAS2.n248 IBIAS2.n245 0.0173591
R14869 IBIAS2.n57 IBIAS2.n56 0.0167343
R14870 IBIAS2.n72 IBIAS2.n71 0.0167343
R14871 IBIAS2.n2 IBIAS2.n1 0.0163451
R14872 IBIAS2.n766 IBIAS2.n765 0.0163451
R14873 IBIAS2.n178 IBIAS2.n177 0.0151658
R14874 IBIAS2.n206 IBIAS2.n205 0.0151658
R14875 IBIAS2.n234 IBIAS2.n233 0.0151658
R14876 IBIAS2.n281 IBIAS2.n280 0.0151658
R14877 IBIAS2.n309 IBIAS2.n308 0.0151658
R14878 IBIAS2.n337 IBIAS2.n336 0.0151658
R14879 IBIAS2.n384 IBIAS2.n383 0.0151658
R14880 IBIAS2.n412 IBIAS2.n411 0.0151658
R14881 IBIAS2.n440 IBIAS2.n439 0.0151658
R14882 IBIAS2.n487 IBIAS2.n486 0.0151658
R14883 IBIAS2.n515 IBIAS2.n514 0.0151658
R14884 IBIAS2.n543 IBIAS2.n542 0.0151658
R14885 IBIAS2.n590 IBIAS2.n589 0.0151658
R14886 IBIAS2.n618 IBIAS2.n617 0.0151658
R14887 IBIAS2.n646 IBIAS2.n645 0.0151658
R14888 IBIAS2.n693 IBIAS2.n692 0.0151658
R14889 IBIAS2.n721 IBIAS2.n720 0.0151658
R14890 IBIAS2.n749 IBIAS2.n748 0.0151658
R14891 IBIAS2.n49 IBIAS2.n48 0.014
R14892 IBIAS2.n9 IBIAS2.n8 0.0119325
R14893 IBIAS2.n765 IBIAS2.n764 0.0112521
R14894 IBIAS2.n153 IBIAS2.n152 0.0111568
R14895 IBIAS2.n256 IBIAS2.n255 0.0111568
R14896 IBIAS2.n359 IBIAS2.n358 0.0111568
R14897 IBIAS2.n462 IBIAS2.n461 0.0111568
R14898 IBIAS2.n565 IBIAS2.n564 0.0111568
R14899 IBIAS2.n668 IBIAS2.n667 0.0111568
R14900 IBIAS2.n98 IBIAS2.n97 0.0111568
R14901 IBIAS2.n125 IBIAS2.n124 0.0111568
R14902 IBIAS2.n29 IBIAS2.n28 0.0111568
R14903 IBIAS2.n241 IBIAS2.n240 0.0100339
R14904 IBIAS2.n181 IBIAS2.n157 0.0100339
R14905 IBIAS2.n344 IBIAS2.n343 0.0100339
R14906 IBIAS2.n284 IBIAS2.n260 0.0100339
R14907 IBIAS2.n447 IBIAS2.n446 0.0100339
R14908 IBIAS2.n387 IBIAS2.n363 0.0100339
R14909 IBIAS2.n550 IBIAS2.n549 0.0100339
R14910 IBIAS2.n490 IBIAS2.n466 0.0100339
R14911 IBIAS2.n653 IBIAS2.n652 0.0100339
R14912 IBIAS2.n593 IBIAS2.n569 0.0100339
R14913 IBIAS2.n756 IBIAS2.n755 0.0100339
R14914 IBIAS2.n696 IBIAS2.n672 0.0100339
R14915 IBIAS2.n141 IBIAS2.n140 0.0100339
R14916 IBIAS2.n137 IBIAS2.n113 0.0100339
R14917 IBIAS2.n110 IBIAS2.n86 0.0100339
R14918 IBIAS2.n83 IBIAS2.n82 0.0100339
R14919 IBIAS2.n142 IBIAS2.n141 0.00965254
R14920 IBIAS2.n3 IBIAS2.n2 0.00905634
R14921 IBIAS2.n1 IBIAS2.n0 0.00905634
R14922 IBIAS2.n12 IBIAS2.n11 0.00899732
R14923 IBIAS2.n156 IBIAS2.n155 0.00845754
R14924 IBIAS2.n259 IBIAS2.n258 0.00845754
R14925 IBIAS2.n362 IBIAS2.n361 0.00845754
R14926 IBIAS2.n465 IBIAS2.n464 0.00845754
R14927 IBIAS2.n568 IBIAS2.n567 0.00845754
R14928 IBIAS2.n671 IBIAS2.n670 0.00845754
R14929 IBIAS2.n136 IBIAS2.n135 0.00845754
R14930 IBIAS2.n109 IBIAS2.n108 0.00845754
R14931 IBIAS2.n40 IBIAS2.n39 0.00845754
R14932 IBIAS2.n17 IBIAS2.n16 0.00845754
R14933 IBIAS2.n236 IBIAS2.n222 0.00838025
R14934 IBIAS2.n208 IBIAS2.n194 0.00838025
R14935 IBIAS2.n180 IBIAS2.n166 0.00838025
R14936 IBIAS2.n339 IBIAS2.n325 0.00838025
R14937 IBIAS2.n311 IBIAS2.n297 0.00838025
R14938 IBIAS2.n283 IBIAS2.n269 0.00838025
R14939 IBIAS2.n442 IBIAS2.n428 0.00838025
R14940 IBIAS2.n414 IBIAS2.n400 0.00838025
R14941 IBIAS2.n386 IBIAS2.n372 0.00838025
R14942 IBIAS2.n545 IBIAS2.n531 0.00838025
R14943 IBIAS2.n517 IBIAS2.n503 0.00838025
R14944 IBIAS2.n489 IBIAS2.n475 0.00838025
R14945 IBIAS2.n648 IBIAS2.n634 0.00838025
R14946 IBIAS2.n620 IBIAS2.n606 0.00838025
R14947 IBIAS2.n592 IBIAS2.n578 0.00838025
R14948 IBIAS2.n751 IBIAS2.n737 0.00838025
R14949 IBIAS2.n723 IBIAS2.n709 0.00838025
R14950 IBIAS2.n695 IBIAS2.n681 0.00838025
R14951 IBIAS2.n50 IBIAS2.n49 0.00776379
R14952 IBIAS2.n183 IBIAS2.n182 0.00775263
R14953 IBIAS2.n286 IBIAS2.n285 0.00775263
R14954 IBIAS2.n389 IBIAS2.n388 0.00775263
R14955 IBIAS2.n492 IBIAS2.n491 0.00775263
R14956 IBIAS2.n595 IBIAS2.n594 0.00775263
R14957 IBIAS2.n698 IBIAS2.n697 0.00775263
R14958 IBIAS2.n80 IBIAS2.n79 0.00773989
R14959 IBIAS2.n68 IBIAS2.n67 0.00773989
R14960 IBIAS2.n65 IBIAS2.n64 0.00773989
R14961 IBIAS2.n53 IBIAS2.n52 0.00773989
R14962 IBIAS2.n81 IBIAS2.n80 0.00773989
R14963 IBIAS2.n79 IBIAS2.n68 0.00773989
R14964 IBIAS2.n66 IBIAS2.n65 0.00773989
R14965 IBIAS2.n64 IBIAS2.n53 0.00773989
R14966 IBIAS2.n51 IBIAS2.n50 0.00771607
R14967 IBIAS2.n237 IBIAS2.n213 0.00577753
R14968 IBIAS2.n209 IBIAS2.n185 0.00577753
R14969 IBIAS2.n340 IBIAS2.n316 0.00577753
R14970 IBIAS2.n312 IBIAS2.n288 0.00577753
R14971 IBIAS2.n443 IBIAS2.n419 0.00577753
R14972 IBIAS2.n415 IBIAS2.n391 0.00577753
R14973 IBIAS2.n546 IBIAS2.n522 0.00577753
R14974 IBIAS2.n518 IBIAS2.n494 0.00577753
R14975 IBIAS2.n649 IBIAS2.n625 0.00577753
R14976 IBIAS2.n621 IBIAS2.n597 0.00577753
R14977 IBIAS2.n752 IBIAS2.n728 0.00577753
R14978 IBIAS2.n724 IBIAS2.n700 0.00577753
R14979 IBIAS2.n213 IBIAS2.n212 0.00574631
R14980 IBIAS2.n185 IBIAS2.n184 0.00574631
R14981 IBIAS2.n316 IBIAS2.n315 0.00574631
R14982 IBIAS2.n288 IBIAS2.n287 0.00574631
R14983 IBIAS2.n419 IBIAS2.n418 0.00574631
R14984 IBIAS2.n391 IBIAS2.n390 0.00574631
R14985 IBIAS2.n522 IBIAS2.n521 0.00574631
R14986 IBIAS2.n494 IBIAS2.n493 0.00574631
R14987 IBIAS2.n625 IBIAS2.n624 0.00574631
R14988 IBIAS2.n597 IBIAS2.n596 0.00574631
R14989 IBIAS2.n728 IBIAS2.n727 0.00574631
R14990 IBIAS2.n700 IBIAS2.n699 0.00574631
R14991 IBIAS2.n242 IBIAS2.n241 0.00558603
R14992 IBIAS2.n345 IBIAS2.n344 0.00558603
R14993 IBIAS2.n448 IBIAS2.n447 0.00558603
R14994 IBIAS2.n551 IBIAS2.n550 0.00558603
R14995 IBIAS2.n654 IBIAS2.n653 0.00558603
R14996 IBIAS2.n757 IBIAS2.n756 0.00558603
R14997 IBIAS2.n138 IBIAS2.n137 0.00558603
R14998 IBIAS2.n111 IBIAS2.n110 0.00558603
R14999 IBIAS2.n84 IBIAS2.n83 0.00558603
R15000 IBIAS2.n238 IBIAS2.n237 0.00557162
R15001 IBIAS2.n210 IBIAS2.n209 0.00557162
R15002 IBIAS2.n211 IBIAS2.n210 0.00557162
R15003 IBIAS2.n239 IBIAS2.n238 0.00557162
R15004 IBIAS2.n341 IBIAS2.n340 0.00557162
R15005 IBIAS2.n313 IBIAS2.n312 0.00557162
R15006 IBIAS2.n314 IBIAS2.n313 0.00557162
R15007 IBIAS2.n342 IBIAS2.n341 0.00557162
R15008 IBIAS2.n444 IBIAS2.n443 0.00557162
R15009 IBIAS2.n416 IBIAS2.n415 0.00557162
R15010 IBIAS2.n417 IBIAS2.n416 0.00557162
R15011 IBIAS2.n445 IBIAS2.n444 0.00557162
R15012 IBIAS2.n547 IBIAS2.n546 0.00557162
R15013 IBIAS2.n519 IBIAS2.n518 0.00557162
R15014 IBIAS2.n520 IBIAS2.n519 0.00557162
R15015 IBIAS2.n548 IBIAS2.n547 0.00557162
R15016 IBIAS2.n650 IBIAS2.n649 0.00557162
R15017 IBIAS2.n622 IBIAS2.n621 0.00557162
R15018 IBIAS2.n623 IBIAS2.n622 0.00557162
R15019 IBIAS2.n651 IBIAS2.n650 0.00557162
R15020 IBIAS2.n753 IBIAS2.n752 0.00557162
R15021 IBIAS2.n725 IBIAS2.n724 0.00557162
R15022 IBIAS2.n726 IBIAS2.n725 0.00557162
R15023 IBIAS2.n754 IBIAS2.n753 0.00557162
R15024 IBIAS2.n243 IBIAS2.n242 0.00555725
R15025 IBIAS2.n346 IBIAS2.n345 0.00555725
R15026 IBIAS2.n449 IBIAS2.n448 0.00555725
R15027 IBIAS2.n552 IBIAS2.n551 0.00555725
R15028 IBIAS2.n655 IBIAS2.n654 0.00555725
R15029 IBIAS2.n758 IBIAS2.n757 0.00555725
R15030 IBIAS2.n139 IBIAS2.n138 0.00555725
R15031 IBIAS2.n112 IBIAS2.n111 0.00555725
R15032 IBIAS2.n85 IBIAS2.n84 0.00555725
R15033 IBIAS2.n182 IBIAS2.n181 0.00438682
R15034 IBIAS2.n285 IBIAS2.n284 0.00438682
R15035 IBIAS2.n388 IBIAS2.n387 0.00438682
R15036 IBIAS2.n491 IBIAS2.n490 0.00438682
R15037 IBIAS2.n594 IBIAS2.n593 0.00438682
R15038 IBIAS2.n697 IBIAS2.n696 0.00438682
R15039 OUT_N.n176 OUT_N.t244 7.30465
R15040 OUT_N.n170 OUT_N.n169 4.07744
R15041 OUT_N.n179 OUT_N.n178 2.40958
R15042 OUT_N.n1909 OUT_N.n1908 1.84464
R15043 OUT_N.n1896 OUT_N.n1895 1.84464
R15044 OUT_N.n169 OUT_N.n168 1.52554
R15045 OUT_N.n2150 OUT_N.n2149 1.50509
R15046 OUT_N.n2156 OUT_N.n2155 1.50275
R15047 OUT_N.n145 OUT_N.n144 1.50001
R15048 OUT_N.n127 OUT_N.n126 1.50001
R15049 OUT_N.n167 OUT_N.n166 1.50001
R15050 OUT_N.n66 OUT_N.n65 1.50001
R15051 OUT_N.n92 OUT_N.n91 1.50001
R15052 OUT_N.n104 OUT_N.n103 1.4999
R15053 OUT_N.n2047 OUT_N.n2046 1.49371
R15054 OUT_N.n2170 OUT_N.n2169 1.49371
R15055 OUT_N.n1631 OUT_N.n1349 1.49371
R15056 OUT_N.n1630 OUT_N.n1351 1.49371
R15057 OUT_N.n2201 OUT_N.n2200 1.49371
R15058 OUT_N.n1672 OUT_N.n1671 1.49371
R15059 OUT_N.n1300 OUT_N.n1299 1.49371
R15060 OUT_N.n942 OUT_N.n941 1.49371
R15061 OUT_N.n2151 OUT_N.n2146 1.48107
R15062 OUT_N.n1939 OUT_N.n1938 1.47979
R15063 OUT_N.n2143 OUT_N.n2142 1.47979
R15064 OUT_N.n1708 OUT_N.n1707 1.47979
R15065 OUT_N.n551 OUT_N.t39 1.46987
R15066 OUT_N.n541 OUT_N.n540 1.46987
R15067 OUT_N.n532 OUT_N.t33 1.46987
R15068 OUT_N.n522 OUT_N.n521 1.46987
R15069 OUT_N.n517 OUT_N.t263 1.46987
R15070 OUT_N.n507 OUT_N.n506 1.46987
R15071 OUT_N.n1823 OUT_N.n1822 1.46987
R15072 OUT_N.n1833 OUT_N.t0 1.46987
R15073 OUT_N.n1838 OUT_N.n1837 1.46987
R15074 OUT_N.n1848 OUT_N.t19 1.46987
R15075 OUT_N.n2011 OUT_N.n2010 1.46987
R15076 OUT_N.n2022 OUT_N.t2 1.46959
R15077 OUT_N.n326 OUT_N.n325 1.43193
R15078 OUT_N.n1454 OUT_N.n1453 1.43193
R15079 OUT_N.n1437 OUT_N.t211 1.43193
R15080 OUT_N.n1433 OUT_N.n1432 1.43193
R15081 OUT_N.n1416 OUT_N.t176 1.43193
R15082 OUT_N.n1412 OUT_N.n1411 1.43193
R15083 OUT_N.n1395 OUT_N.t167 1.43193
R15084 OUT_N.n1391 OUT_N.n1390 1.43193
R15085 OUT_N.n1374 OUT_N.t121 1.43193
R15086 OUT_N.n1370 OUT_N.n1369 1.43193
R15087 OUT_N.n1306 OUT_N.t191 1.43193
R15088 OUT_N.n1323 OUT_N.n1322 1.43193
R15089 OUT_N.n1327 OUT_N.t147 1.43193
R15090 OUT_N.n1344 OUT_N.n1343 1.43193
R15091 OUT_N.n1353 OUT_N.t114 1.43193
R15092 OUT_N.n309 OUT_N.t155 1.43193
R15093 OUT_N.n305 OUT_N.n304 1.43193
R15094 OUT_N.n288 OUT_N.t206 1.43193
R15095 OUT_N.n284 OUT_N.n283 1.43193
R15096 OUT_N.n267 OUT_N.t90 1.43193
R15097 OUT_N.n263 OUT_N.n262 1.43193
R15098 OUT_N.n246 OUT_N.t145 1.43193
R15099 OUT_N.n242 OUT_N.n241 1.43193
R15100 OUT_N.n225 OUT_N.t200 1.43193
R15101 OUT_N.n221 OUT_N.n220 1.43193
R15102 OUT_N.n204 OUT_N.t156 1.43193
R15103 OUT_N.n200 OUT_N.n199 1.43193
R15104 OUT_N.n183 OUT_N.t162 1.43193
R15105 OUT_N.n1903 OUT_N.n1902 1.28777
R15106 OUT_N.n2065 OUT_N.n2064 1.28777
R15107 OUT_N.n2058 OUT_N.n2057 1.28777
R15108 OUT_N.n2075 OUT_N.n2074 1.28777
R15109 OUT_N.n1778 OUT_N.n1777 1.28777
R15110 OUT_N.n1786 OUT_N.n1785 1.28777
R15111 OUT_N.n1770 OUT_N.n1769 1.28777
R15112 OUT_N.n2178 OUT_N.n2175 1.1949
R15113 OUT_N.n2188 OUT_N.n2187 1.1949
R15114 OUT_N.n1981 OUT_N.n1980 1.1949
R15115 OUT_N.n1988 OUT_N.n1985 1.1949
R15116 OUT_N.n11 OUT_N.n10 1.1949
R15117 OUT_N.n18 OUT_N.n15 1.1949
R15118 OUT_N.n1740 OUT_N.n1739 1.1949
R15119 OUT_N.n1747 OUT_N.n1744 1.1949
R15120 OUT_N.n783 OUT_N.n782 1.1948
R15121 OUT_N.n771 OUT_N.n770 1.1948
R15122 OUT_N.n759 OUT_N.n758 1.1948
R15123 OUT_N.n747 OUT_N.n746 1.1948
R15124 OUT_N.n735 OUT_N.n734 1.1948
R15125 OUT_N.n723 OUT_N.n722 1.1948
R15126 OUT_N.n627 OUT_N.n626 1.1948
R15127 OUT_N.n639 OUT_N.n638 1.1948
R15128 OUT_N.n651 OUT_N.n650 1.1948
R15129 OUT_N.n663 OUT_N.n662 1.1948
R15130 OUT_N.n675 OUT_N.n674 1.1948
R15131 OUT_N.n687 OUT_N.n686 1.1948
R15132 OUT_N.n699 OUT_N.n698 1.1948
R15133 OUT_N.n711 OUT_N.n710 1.1948
R15134 OUT_N.n1118 OUT_N.n1117 1.1948
R15135 OUT_N.n1106 OUT_N.n1105 1.1948
R15136 OUT_N.n1094 OUT_N.n1093 1.1948
R15137 OUT_N.n1082 OUT_N.n1081 1.1948
R15138 OUT_N.n1070 OUT_N.n1069 1.1948
R15139 OUT_N.n1058 OUT_N.n1057 1.1948
R15140 OUT_N.n1046 OUT_N.n1045 1.1948
R15141 OUT_N.n1034 OUT_N.n1033 1.1948
R15142 OUT_N.n1022 OUT_N.n1021 1.1948
R15143 OUT_N.n1010 OUT_N.n1009 1.1948
R15144 OUT_N.n956 OUT_N.n955 1.1948
R15145 OUT_N.n968 OUT_N.n967 1.1948
R15146 OUT_N.n980 OUT_N.n979 1.1948
R15147 OUT_N.n992 OUT_N.n991 1.1948
R15148 OUT_N.n1438 OUT_N.n1437 1.19473
R15149 OUT_N.n1417 OUT_N.n1416 1.19473
R15150 OUT_N.n1396 OUT_N.n1395 1.19473
R15151 OUT_N.n1375 OUT_N.n1374 1.19473
R15152 OUT_N.n1307 OUT_N.n1306 1.19473
R15153 OUT_N.n1328 OUT_N.n1327 1.19473
R15154 OUT_N.n1354 OUT_N.n1353 1.19473
R15155 OUT_N.n310 OUT_N.n309 1.19473
R15156 OUT_N.n289 OUT_N.n288 1.19473
R15157 OUT_N.n268 OUT_N.n267 1.19473
R15158 OUT_N.n247 OUT_N.n246 1.19473
R15159 OUT_N.n226 OUT_N.n225 1.19473
R15160 OUT_N.n205 OUT_N.n204 1.19473
R15161 OUT_N.n184 OUT_N.n183 1.19473
R15162 OUT_N.n2106 OUT_N.n2105 1.19461
R15163 OUT_N.n1866 OUT_N.n1865 1.19461
R15164 OUT_N.n552 OUT_N.n551 1.19458
R15165 OUT_N.n542 OUT_N.n541 1.19458
R15166 OUT_N.n518 OUT_N.n517 1.19458
R15167 OUT_N.n508 OUT_N.n507 1.19458
R15168 OUT_N.n1839 OUT_N.n1838 1.19458
R15169 OUT_N.n1849 OUT_N.n1848 1.19458
R15170 OUT_N.n322 OUT_N.n321 1.19445
R15171 OUT_N.n1450 OUT_N.n1449 1.19445
R15172 OUT_N.n1429 OUT_N.n1428 1.19445
R15173 OUT_N.n1408 OUT_N.n1407 1.19445
R15174 OUT_N.n1387 OUT_N.n1386 1.19445
R15175 OUT_N.n1366 OUT_N.n1365 1.19445
R15176 OUT_N.n1319 OUT_N.n1318 1.19445
R15177 OUT_N.n1340 OUT_N.n1339 1.19445
R15178 OUT_N.n301 OUT_N.n300 1.19445
R15179 OUT_N.n280 OUT_N.n279 1.19445
R15180 OUT_N.n259 OUT_N.n258 1.19445
R15181 OUT_N.n238 OUT_N.n237 1.19445
R15182 OUT_N.n217 OUT_N.n216 1.19445
R15183 OUT_N.n196 OUT_N.n195 1.19445
R15184 OUT_N.n529 OUT_N.n528 1.19426
R15185 OUT_N.n1830 OUT_N.n1829 1.19426
R15186 OUT_N.n2018 OUT_N.n2017 1.19426
R15187 OUT_N.n548 OUT_N.n547 1.17959
R15188 OUT_N.n514 OUT_N.n513 1.17959
R15189 OUT_N.n1845 OUT_N.n1844 1.17959
R15190 OUT_N.n533 OUT_N.n532 1.1793
R15191 OUT_N.n523 OUT_N.n522 1.1793
R15192 OUT_N.n1824 OUT_N.n1823 1.1793
R15193 OUT_N.n1834 OUT_N.n1833 1.1793
R15194 OUT_N.n2012 OUT_N.n2011 1.1793
R15195 OUT_N.n316 OUT_N.n315 1.1791
R15196 OUT_N.n1444 OUT_N.n1443 1.1791
R15197 OUT_N.n1423 OUT_N.n1422 1.1791
R15198 OUT_N.n1402 OUT_N.n1401 1.1791
R15199 OUT_N.n1381 OUT_N.n1380 1.1791
R15200 OUT_N.n1360 OUT_N.n1359 1.1791
R15201 OUT_N.n1313 OUT_N.n1312 1.1791
R15202 OUT_N.n1334 OUT_N.n1333 1.1791
R15203 OUT_N.n295 OUT_N.n294 1.1791
R15204 OUT_N.n274 OUT_N.n273 1.1791
R15205 OUT_N.n253 OUT_N.n252 1.1791
R15206 OUT_N.n232 OUT_N.n231 1.1791
R15207 OUT_N.n211 OUT_N.n210 1.1791
R15208 OUT_N.n190 OUT_N.n189 1.1791
R15209 OUT_N.n1872 OUT_N.n1871 1.17896
R15210 OUT_N.n2100 OUT_N.n2099 1.17896
R15211 OUT_N.n2023 OUT_N.n2022 1.17896
R15212 OUT_N.n327 OUT_N.n326 1.17884
R15213 OUT_N.n1455 OUT_N.n1454 1.17884
R15214 OUT_N.n1434 OUT_N.n1433 1.17884
R15215 OUT_N.n1413 OUT_N.n1412 1.17884
R15216 OUT_N.n1392 OUT_N.n1391 1.17884
R15217 OUT_N.n1371 OUT_N.n1370 1.17884
R15218 OUT_N.n1324 OUT_N.n1323 1.17884
R15219 OUT_N.n1345 OUT_N.n1344 1.17884
R15220 OUT_N.n306 OUT_N.n305 1.17884
R15221 OUT_N.n285 OUT_N.n284 1.17884
R15222 OUT_N.n264 OUT_N.n263 1.17884
R15223 OUT_N.n243 OUT_N.n242 1.17884
R15224 OUT_N.n222 OUT_N.n221 1.17884
R15225 OUT_N.n201 OUT_N.n200 1.17884
R15226 OUT_N.n777 OUT_N.n776 1.17849
R15227 OUT_N.n765 OUT_N.n764 1.17849
R15228 OUT_N.n753 OUT_N.n752 1.17849
R15229 OUT_N.n741 OUT_N.n740 1.17849
R15230 OUT_N.n729 OUT_N.n728 1.17849
R15231 OUT_N.n621 OUT_N.n620 1.17849
R15232 OUT_N.n633 OUT_N.n632 1.17849
R15233 OUT_N.n645 OUT_N.n644 1.17849
R15234 OUT_N.n657 OUT_N.n656 1.17849
R15235 OUT_N.n669 OUT_N.n668 1.17849
R15236 OUT_N.n681 OUT_N.n680 1.17849
R15237 OUT_N.n693 OUT_N.n692 1.17849
R15238 OUT_N.n705 OUT_N.n704 1.17849
R15239 OUT_N.n717 OUT_N.n716 1.17849
R15240 OUT_N.n1112 OUT_N.n1111 1.17849
R15241 OUT_N.n1100 OUT_N.n1099 1.17849
R15242 OUT_N.n1088 OUT_N.n1087 1.17849
R15243 OUT_N.n1076 OUT_N.n1075 1.17849
R15244 OUT_N.n1064 OUT_N.n1063 1.17849
R15245 OUT_N.n1052 OUT_N.n1051 1.17849
R15246 OUT_N.n1040 OUT_N.n1039 1.17849
R15247 OUT_N.n1028 OUT_N.n1027 1.17849
R15248 OUT_N.n1016 OUT_N.n1015 1.17849
R15249 OUT_N.n950 OUT_N.n949 1.17849
R15250 OUT_N.n962 OUT_N.n961 1.17849
R15251 OUT_N.n974 OUT_N.n973 1.17849
R15252 OUT_N.n986 OUT_N.n985 1.17849
R15253 OUT_N.n1004 OUT_N.n1003 1.17849
R15254 OUT_N.n2059 OUT_N.n2058 1.1742
R15255 OUT_N.n2076 OUT_N.n2075 1.1742
R15256 OUT_N.n2155 OUT_N.n2154 1.16696
R15257 OUT_N.n1944 OUT_N.n1943 1.16696
R15258 OUT_N.n1966 OUT_N.n1965 1.16696
R15259 OUT_N.n2136 OUT_N.n2135 1.16696
R15260 OUT_N.n1699 OUT_N.n1698 1.16696
R15261 OUT_N.n1720 OUT_N.n1719 1.16696
R15262 OUT_N.n1897 OUT_N.n1896 1.14437
R15263 OUT_N.n1940 OUT_N.n1939 1.14073
R15264 OUT_N.n2144 OUT_N.n2143 1.14073
R15265 OUT_N.n1709 OUT_N.n1708 1.14073
R15266 OUT_N.n1686 OUT_N.n1685 1.1353
R15267 OUT_N.n1734 OUT_N.n1733 1.12925
R15268 OUT_N.n1764 OUT_N.n1763 1.12925
R15269 OUT_N.n2179 OUT_N.n2178 1.12829
R15270 OUT_N.n1914 OUT_N.n1913 1.12829
R15271 OUT_N.n1700 OUT_N.n1699 1.12829
R15272 OUT_N.n1989 OUT_N.n1988 1.12795
R15273 OUT_N.n19 OUT_N.n18 1.12795
R15274 OUT_N.n1789 OUT_N.n1788 1.12795
R15275 OUT_N.n1748 OUT_N.n1747 1.12795
R15276 OUT_N.n2024 OUT_N.n2023 1.12758
R15277 OUT_N.n1710 OUT_N.n1709 1.12695
R15278 OUT_N.n1947 OUT_N.n1946 1.1255
R15279 OUT_N.n1913 OUT_N.n1910 1.1255
R15280 OUT_N.n1962 OUT_N.n1961 1.1255
R15281 OUT_N.n1893 OUT_N.n1892 1.1255
R15282 OUT_N.n1905 OUT_N.n1904 1.1255
R15283 OUT_N.n2067 OUT_N.n2066 1.1255
R15284 OUT_N.n2056 OUT_N.n2055 1.1255
R15285 OUT_N.n2072 OUT_N.n2071 1.1255
R15286 OUT_N.n2149 OUT_N.n2148 1.1255
R15287 OUT_N.n2140 OUT_N.n2139 1.1255
R15288 OUT_N.n2133 OUT_N.n2132 1.1255
R15289 OUT_N.n1936 OUT_N.n1935 1.1255
R15290 OUT_N.n1780 OUT_N.n1779 1.1255
R15291 OUT_N.n1691 OUT_N.n1690 1.1255
R15292 OUT_N.n1788 OUT_N.n1787 1.1255
R15293 OUT_N.n1716 OUT_N.n1715 1.1255
R15294 OUT_N.n1772 OUT_N.n1771 1.1255
R15295 OUT_N.n2000 OUT_N.n1999 1.11801
R15296 OUT_N.n1928 OUT_N.n1927 1.11801
R15297 OUT_N.n1884 OUT_N.n1883 1.11801
R15298 OUT_N.n2126 OUT_N.n2092 1.11801
R15299 OUT_N.n2196 OUT_N.n2053 1.11801
R15300 OUT_N.n1244 OUT_N.n999 1.11801
R15301 OUT_N.n1540 OUT_N.n1539 1.11801
R15302 OUT_N.n1620 OUT_N.n1619 1.11801
R15303 OUT_N.n1628 OUT_N.n1627 1.11801
R15304 OUT_N.n1579 OUT_N.n1578 1.11801
R15305 OUT_N.n1559 OUT_N.n1558 1.11801
R15306 OUT_N.n1147 OUT_N.n1146 1.11801
R15307 OUT_N.n1499 OUT_N.n1498 1.11801
R15308 OUT_N.n1158 OUT_N.n1157 1.11801
R15309 OUT_N.n574 OUT_N.n538 1.11801
R15310 OUT_N.n575 OUT_N.n536 1.11801
R15311 OUT_N.n466 OUT_N.n465 1.11801
R15312 OUT_N.n454 OUT_N.n453 1.11801
R15313 OUT_N.n413 OUT_N.n412 1.11801
R15314 OUT_N.n410 OUT_N.n409 1.11801
R15315 OUT_N.n364 OUT_N.n363 1.11801
R15316 OUT_N.n355 OUT_N.n354 1.11801
R15317 OUT_N.n457 OUT_N.n456 1.11801
R15318 OUT_N.n1759 OUT_N.n1758 1.11801
R15319 OUT_N.n1810 OUT_N.n1725 1.11801
R15320 OUT_N.n2044 OUT_N.n2043 1.11801
R15321 OUT_N.n2236 OUT_N.n2235 1.11801
R15322 OUT_N.n2233 OUT_N.n1820 1.11801
R15323 OUT_N.n2040 OUT_N.n2008 1.11801
R15324 OUT_N.n611 OUT_N.n610 1.11801
R15325 OUT_N.n1678 OUT_N.n33 1.11801
R15326 OUT_N.n178 OUT_N.n171 1.11801
R15327 OUT_N.n1976 OUT_N.n1975 1.11782
R15328 OUT_N.n1971 OUT_N.n1970 1.11782
R15329 OUT_N.n2004 OUT_N.n2003 1.11782
R15330 OUT_N.n1885 OUT_N.n1854 1.11782
R15331 OUT_N.n2118 OUT_N.n2117 1.11782
R15332 OUT_N.n2122 OUT_N.n2121 1.11782
R15333 OUT_N.n2195 OUT_N.n2194 1.11782
R15334 OUT_N.n1257 OUT_N.n1256 1.11782
R15335 OUT_N.n1486 OUT_N.n1485 1.11782
R15336 OUT_N.n361 OUT_N.n360 1.11782
R15337 OUT_N.n463 OUT_N.n462 1.11782
R15338 OUT_N.n1805 OUT_N.n1804 1.11782
R15339 OUT_N.n1809 OUT_N.n1808 1.11782
R15340 OUT_N.n2239 OUT_N.n2238 1.11782
R15341 OUT_N.n1677 OUT_N.n1676 1.11782
R15342 OUT_N.n177 OUT_N.n176 1.11782
R15343 OUT_N.n2241 OUT_N.n2240 1.11782
R15344 OUT_N.n1705 OUT_N.n1692 1.10737
R15345 OUT_N.n1943 OUT_N.n1942 1.09451
R15346 OUT_N.n1965 OUT_N.n1964 1.09451
R15347 OUT_N.n2135 OUT_N.n2134 1.09451
R15348 OUT_N.n2154 OUT_N.n2153 1.09451
R15349 OUT_N.n1698 OUT_N.n1695 1.09451
R15350 OUT_N.n1719 OUT_N.n1718 1.09451
R15351 OUT_N.n2105 OUT_N.n2104 0.923611
R15352 OUT_N.n1865 OUT_N.n1864 0.923611
R15353 OUT_N.n1871 OUT_N.n1870 0.923589
R15354 OUT_N.n2099 OUT_N.n2098 0.923589
R15355 OUT_N.n2175 OUT_N.n2174 0.923589
R15356 OUT_N.n2187 OUT_N.n2186 0.923589
R15357 OUT_N.n1980 OUT_N.n1979 0.923589
R15358 OUT_N.n1985 OUT_N.n1984 0.923589
R15359 OUT_N.n10 OUT_N.n9 0.923589
R15360 OUT_N.n15 OUT_N.n14 0.923589
R15361 OUT_N.n1739 OUT_N.n1738 0.923589
R15362 OUT_N.n1744 OUT_N.n1743 0.923589
R15363 OUT_N.n547 OUT_N.n546 0.923538
R15364 OUT_N.n528 OUT_N.n527 0.923538
R15365 OUT_N.n513 OUT_N.n512 0.923538
R15366 OUT_N.n1829 OUT_N.n1828 0.923538
R15367 OUT_N.n1844 OUT_N.n1843 0.923538
R15368 OUT_N.n2017 OUT_N.n2016 0.923538
R15369 OUT_N.n1995 OUT_N.n1982 0.885703
R15370 OUT_N.n2190 OUT_N.n2189 0.885703
R15371 OUT_N.n25 OUT_N.n12 0.885703
R15372 OUT_N.n1722 OUT_N.n1721 0.885703
R15373 OUT_N.n1754 OUT_N.n1741 0.885703
R15374 OUT_N.n590 OUT_N.n589 0.835535
R15375 OUT_N.n2216 OUT_N.n2215 0.835535
R15376 OUT_N.n782 OUT_N.n781 0.824999
R15377 OUT_N.n770 OUT_N.n769 0.824999
R15378 OUT_N.n758 OUT_N.n757 0.824999
R15379 OUT_N.n746 OUT_N.n745 0.824999
R15380 OUT_N.n734 OUT_N.n733 0.824999
R15381 OUT_N.n722 OUT_N.n721 0.824999
R15382 OUT_N.n626 OUT_N.n625 0.824999
R15383 OUT_N.n638 OUT_N.n637 0.824999
R15384 OUT_N.n650 OUT_N.n649 0.824999
R15385 OUT_N.n662 OUT_N.n661 0.824999
R15386 OUT_N.n674 OUT_N.n673 0.824999
R15387 OUT_N.n686 OUT_N.n685 0.824999
R15388 OUT_N.n698 OUT_N.n697 0.824999
R15389 OUT_N.n710 OUT_N.n709 0.824999
R15390 OUT_N.n1117 OUT_N.n1116 0.824999
R15391 OUT_N.n1105 OUT_N.n1104 0.824999
R15392 OUT_N.n1093 OUT_N.n1092 0.824999
R15393 OUT_N.n1081 OUT_N.n1080 0.824999
R15394 OUT_N.n1069 OUT_N.n1068 0.824999
R15395 OUT_N.n1057 OUT_N.n1056 0.824999
R15396 OUT_N.n1045 OUT_N.n1044 0.824999
R15397 OUT_N.n1033 OUT_N.n1032 0.824999
R15398 OUT_N.n1021 OUT_N.n1020 0.824999
R15399 OUT_N.n1009 OUT_N.n1008 0.824999
R15400 OUT_N.n955 OUT_N.n954 0.824999
R15401 OUT_N.n967 OUT_N.n966 0.824999
R15402 OUT_N.n979 OUT_N.n978 0.824999
R15403 OUT_N.n991 OUT_N.n990 0.824999
R15404 OUT_N.n776 OUT_N.n775 0.824997
R15405 OUT_N.n764 OUT_N.n763 0.824997
R15406 OUT_N.n752 OUT_N.n751 0.824997
R15407 OUT_N.n740 OUT_N.n739 0.824997
R15408 OUT_N.n728 OUT_N.n727 0.824997
R15409 OUT_N.n620 OUT_N.n619 0.824997
R15410 OUT_N.n632 OUT_N.n631 0.824997
R15411 OUT_N.n644 OUT_N.n643 0.824997
R15412 OUT_N.n656 OUT_N.n655 0.824997
R15413 OUT_N.n668 OUT_N.n667 0.824997
R15414 OUT_N.n680 OUT_N.n679 0.824997
R15415 OUT_N.n692 OUT_N.n691 0.824997
R15416 OUT_N.n704 OUT_N.n703 0.824997
R15417 OUT_N.n716 OUT_N.n715 0.824997
R15418 OUT_N.n1111 OUT_N.n1110 0.824997
R15419 OUT_N.n1099 OUT_N.n1098 0.824997
R15420 OUT_N.n1087 OUT_N.n1086 0.824997
R15421 OUT_N.n1075 OUT_N.n1074 0.824997
R15422 OUT_N.n1063 OUT_N.n1062 0.824997
R15423 OUT_N.n1051 OUT_N.n1050 0.824997
R15424 OUT_N.n1039 OUT_N.n1038 0.824997
R15425 OUT_N.n1027 OUT_N.n1026 0.824997
R15426 OUT_N.n1015 OUT_N.n1014 0.824997
R15427 OUT_N.n949 OUT_N.n948 0.824997
R15428 OUT_N.n961 OUT_N.n960 0.824997
R15429 OUT_N.n973 OUT_N.n972 0.824997
R15430 OUT_N.n985 OUT_N.n984 0.824997
R15431 OUT_N.n1003 OUT_N.n1002 0.824997
R15432 OUT_N.n321 OUT_N.n320 0.82495
R15433 OUT_N.n315 OUT_N.n314 0.82495
R15434 OUT_N.n1449 OUT_N.n1448 0.82495
R15435 OUT_N.n1443 OUT_N.n1442 0.82495
R15436 OUT_N.n1428 OUT_N.n1427 0.82495
R15437 OUT_N.n1422 OUT_N.n1421 0.82495
R15438 OUT_N.n1407 OUT_N.n1406 0.82495
R15439 OUT_N.n1401 OUT_N.n1400 0.82495
R15440 OUT_N.n1386 OUT_N.n1385 0.82495
R15441 OUT_N.n1380 OUT_N.n1379 0.82495
R15442 OUT_N.n1365 OUT_N.n1364 0.82495
R15443 OUT_N.n1359 OUT_N.n1358 0.82495
R15444 OUT_N.n1312 OUT_N.n1311 0.82495
R15445 OUT_N.n1318 OUT_N.n1317 0.82495
R15446 OUT_N.n1333 OUT_N.n1332 0.82495
R15447 OUT_N.n1339 OUT_N.n1338 0.82495
R15448 OUT_N.n300 OUT_N.n299 0.82495
R15449 OUT_N.n294 OUT_N.n293 0.82495
R15450 OUT_N.n279 OUT_N.n278 0.82495
R15451 OUT_N.n273 OUT_N.n272 0.82495
R15452 OUT_N.n258 OUT_N.n257 0.82495
R15453 OUT_N.n252 OUT_N.n251 0.82495
R15454 OUT_N.n237 OUT_N.n236 0.82495
R15455 OUT_N.n231 OUT_N.n230 0.82495
R15456 OUT_N.n216 OUT_N.n215 0.82495
R15457 OUT_N.n210 OUT_N.n209 0.82495
R15458 OUT_N.n195 OUT_N.n194 0.82495
R15459 OUT_N.n189 OUT_N.n188 0.82495
R15460 OUT_N.n102 OUT_N.n101 0.736598
R15461 OUT_N.n2082 OUT_N.n2068 0.727104
R15462 OUT_N.n2160 OUT_N.n2145 0.727104
R15463 OUT_N.n2165 OUT_N.n2137 0.727104
R15464 OUT_N.n1955 OUT_N.n1941 0.727104
R15465 OUT_N.n1880 OUT_N.n1867 0.727104
R15466 OUT_N.n2109 OUT_N.n2107 0.727104
R15467 OUT_N.n1290 OUT_N.n957 0.727104
R15468 OUT_N.n1281 OUT_N.n969 0.727104
R15469 OUT_N.n1272 OUT_N.n981 0.727104
R15470 OUT_N.n1263 OUT_N.n993 0.727104
R15471 OUT_N.n1121 OUT_N.n1119 0.727104
R15472 OUT_N.n1130 OUT_N.n1107 0.727104
R15473 OUT_N.n1161 OUT_N.n1095 0.727104
R15474 OUT_N.n1170 OUT_N.n1083 0.727104
R15475 OUT_N.n1179 OUT_N.n1071 0.727104
R15476 OUT_N.n1188 OUT_N.n1059 0.727104
R15477 OUT_N.n1207 OUT_N.n1047 0.727104
R15478 OUT_N.n1216 OUT_N.n1035 0.727104
R15479 OUT_N.n1225 OUT_N.n1023 0.727104
R15480 OUT_N.n1234 OUT_N.n1011 0.727104
R15481 OUT_N.n1662 OUT_N.n1314 0.727104
R15482 OUT_N.n1653 OUT_N.n1325 0.727104
R15483 OUT_N.n1644 OUT_N.n1335 0.727104
R15484 OUT_N.n1635 OUT_N.n1346 0.727104
R15485 OUT_N.n1458 OUT_N.n1456 0.727104
R15486 OUT_N.n1467 OUT_N.n1445 0.727104
R15487 OUT_N.n1502 OUT_N.n1435 0.727104
R15488 OUT_N.n1511 OUT_N.n1424 0.727104
R15489 OUT_N.n1520 OUT_N.n1414 0.727104
R15490 OUT_N.n1529 OUT_N.n1403 0.727104
R15491 OUT_N.n1582 OUT_N.n1393 0.727104
R15492 OUT_N.n1591 OUT_N.n1382 0.727104
R15493 OUT_N.n1600 OUT_N.n1372 0.727104
R15494 OUT_N.n1609 OUT_N.n1361 0.727104
R15495 OUT_N.n931 OUT_N.n628 0.727104
R15496 OUT_N.n922 OUT_N.n640 0.727104
R15497 OUT_N.n913 OUT_N.n652 0.727104
R15498 OUT_N.n904 OUT_N.n664 0.727104
R15499 OUT_N.n885 OUT_N.n676 0.727104
R15500 OUT_N.n876 OUT_N.n688 0.727104
R15501 OUT_N.n867 OUT_N.n700 0.727104
R15502 OUT_N.n858 OUT_N.n712 0.727104
R15503 OUT_N.n786 OUT_N.n784 0.727104
R15504 OUT_N.n795 OUT_N.n772 0.727104
R15505 OUT_N.n814 OUT_N.n760 0.727104
R15506 OUT_N.n823 OUT_N.n748 0.727104
R15507 OUT_N.n832 OUT_N.n736 0.727104
R15508 OUT_N.n841 OUT_N.n724 0.727104
R15509 OUT_N.n560 OUT_N.n549 0.727104
R15510 OUT_N.n578 OUT_N.n534 0.727104
R15511 OUT_N.n587 OUT_N.n524 0.727104
R15512 OUT_N.n596 OUT_N.n515 0.727104
R15513 OUT_N.n330 OUT_N.n328 0.727104
R15514 OUT_N.n339 OUT_N.n317 0.727104
R15515 OUT_N.n367 OUT_N.n307 0.727104
R15516 OUT_N.n376 OUT_N.n296 0.727104
R15517 OUT_N.n385 OUT_N.n286 0.727104
R15518 OUT_N.n394 OUT_N.n275 0.727104
R15519 OUT_N.n416 OUT_N.n265 0.727104
R15520 OUT_N.n425 OUT_N.n254 0.727104
R15521 OUT_N.n434 OUT_N.n244 0.727104
R15522 OUT_N.n443 OUT_N.n233 0.727104
R15523 OUT_N.n469 OUT_N.n223 0.727104
R15524 OUT_N.n478 OUT_N.n212 0.727104
R15525 OUT_N.n487 OUT_N.n202 0.727104
R15526 OUT_N.n496 OUT_N.n191 0.727104
R15527 OUT_N.n1795 OUT_N.n1781 0.727104
R15528 OUT_N.n2227 OUT_N.n1825 0.727104
R15529 OUT_N.n2218 OUT_N.n1835 0.727104
R15530 OUT_N.n2209 OUT_N.n1846 0.727104
R15531 OUT_N.n2034 OUT_N.n2013 0.727104
R15532 OUT_N.n1919 OUT_N.n1906 0.726858
R15533 OUT_N.n1800 OUT_N.n1773 0.726858
R15534 OUT_N.n1177 OUT_N.n1176 0.685007
R15535 OUT_N.n1223 OUT_N.n1222 0.685007
R15536 OUT_N.n1279 OUT_N.n1278 0.685007
R15537 OUT_N.n830 OUT_N.n829 0.685007
R15538 OUT_N.n874 OUT_N.n873 0.685007
R15539 OUT_N.n920 OUT_N.n919 0.685007
R15540 OUT_N.n2240 OUT_N.n2239 0.659441
R15541 OUT_N.n1968 OUT_N.n1967 0.617177
R15542 OUT_N.n335 OUT_N.n323 0.616779
R15543 OUT_N.n555 OUT_N.n553 0.616779
R15544 OUT_N.n564 OUT_N.n543 0.616779
R15545 OUT_N.n1875 OUT_N.n1873 0.616779
R15546 OUT_N.n2114 OUT_N.n2101 0.616779
R15547 OUT_N.n1950 OUT_N.n1948 0.616779
R15548 OUT_N.n1923 OUT_N.n1898 0.616779
R15549 OUT_N.n2078 OUT_N.n2077 0.616779
R15550 OUT_N.n2087 OUT_N.n2060 0.616779
R15551 OUT_N.n582 OUT_N.n530 0.616779
R15552 OUT_N.n591 OUT_N.n519 0.616779
R15553 OUT_N.n600 OUT_N.n509 0.616779
R15554 OUT_N.n791 OUT_N.n778 0.616779
R15555 OUT_N.n800 OUT_N.n766 0.616779
R15556 OUT_N.n819 OUT_N.n754 0.616779
R15557 OUT_N.n828 OUT_N.n742 0.616779
R15558 OUT_N.n837 OUT_N.n730 0.616779
R15559 OUT_N.n936 OUT_N.n622 0.616779
R15560 OUT_N.n927 OUT_N.n634 0.616779
R15561 OUT_N.n918 OUT_N.n646 0.616779
R15562 OUT_N.n909 OUT_N.n658 0.616779
R15563 OUT_N.n890 OUT_N.n670 0.616779
R15564 OUT_N.n881 OUT_N.n682 0.616779
R15565 OUT_N.n872 OUT_N.n694 0.616779
R15566 OUT_N.n863 OUT_N.n706 0.616779
R15567 OUT_N.n846 OUT_N.n718 0.616779
R15568 OUT_N.n1463 OUT_N.n1451 0.616779
R15569 OUT_N.n1472 OUT_N.n1439 0.616779
R15570 OUT_N.n1507 OUT_N.n1430 0.616779
R15571 OUT_N.n1516 OUT_N.n1418 0.616779
R15572 OUT_N.n1525 OUT_N.n1409 0.616779
R15573 OUT_N.n1534 OUT_N.n1397 0.616779
R15574 OUT_N.n1587 OUT_N.n1388 0.616779
R15575 OUT_N.n1596 OUT_N.n1376 0.616779
R15576 OUT_N.n1605 OUT_N.n1367 0.616779
R15577 OUT_N.n1667 OUT_N.n1308 0.616779
R15578 OUT_N.n1658 OUT_N.n1320 0.616779
R15579 OUT_N.n1649 OUT_N.n1329 0.616779
R15580 OUT_N.n1640 OUT_N.n1341 0.616779
R15581 OUT_N.n1614 OUT_N.n1355 0.616779
R15582 OUT_N.n1126 OUT_N.n1113 0.616779
R15583 OUT_N.n1135 OUT_N.n1101 0.616779
R15584 OUT_N.n1166 OUT_N.n1089 0.616779
R15585 OUT_N.n1175 OUT_N.n1077 0.616779
R15586 OUT_N.n1184 OUT_N.n1065 0.616779
R15587 OUT_N.n1193 OUT_N.n1053 0.616779
R15588 OUT_N.n1212 OUT_N.n1041 0.616779
R15589 OUT_N.n1221 OUT_N.n1029 0.616779
R15590 OUT_N.n1230 OUT_N.n1017 0.616779
R15591 OUT_N.n1295 OUT_N.n951 0.616779
R15592 OUT_N.n1286 OUT_N.n963 0.616779
R15593 OUT_N.n1277 OUT_N.n975 0.616779
R15594 OUT_N.n1268 OUT_N.n987 0.616779
R15595 OUT_N.n1239 OUT_N.n1005 0.616779
R15596 OUT_N.n344 OUT_N.n311 0.616779
R15597 OUT_N.n372 OUT_N.n302 0.616779
R15598 OUT_N.n381 OUT_N.n290 0.616779
R15599 OUT_N.n390 OUT_N.n281 0.616779
R15600 OUT_N.n399 OUT_N.n269 0.616779
R15601 OUT_N.n421 OUT_N.n260 0.616779
R15602 OUT_N.n430 OUT_N.n248 0.616779
R15603 OUT_N.n439 OUT_N.n239 0.616779
R15604 OUT_N.n448 OUT_N.n227 0.616779
R15605 OUT_N.n474 OUT_N.n218 0.616779
R15606 OUT_N.n483 OUT_N.n206 0.616779
R15607 OUT_N.n492 OUT_N.n197 0.616779
R15608 OUT_N.n501 OUT_N.n185 0.616779
R15609 OUT_N.n2222 OUT_N.n1831 0.616779
R15610 OUT_N.n2213 OUT_N.n1840 0.616779
R15611 OUT_N.n2204 OUT_N.n1850 0.616779
R15612 OUT_N.n2029 OUT_N.n2019 0.616779
R15613 OUT_N.n320 OUT_N.t175 0.607167
R15614 OUT_N.n320 OUT_N.n319 0.607167
R15615 OUT_N.n314 OUT_N.t188 0.607167
R15616 OUT_N.n314 OUT_N.n313 0.607167
R15617 OUT_N.n781 OUT_N.t92 0.607167
R15618 OUT_N.n781 OUT_N.n780 0.607167
R15619 OUT_N.n775 OUT_N.t179 0.607167
R15620 OUT_N.n775 OUT_N.n774 0.607167
R15621 OUT_N.n769 OUT_N.t243 0.607167
R15622 OUT_N.n769 OUT_N.n768 0.607167
R15623 OUT_N.n763 OUT_N.t184 0.607167
R15624 OUT_N.n763 OUT_N.n762 0.607167
R15625 OUT_N.n757 OUT_N.t194 0.607167
R15626 OUT_N.n757 OUT_N.n756 0.607167
R15627 OUT_N.n751 OUT_N.t62 0.607167
R15628 OUT_N.n751 OUT_N.n750 0.607167
R15629 OUT_N.n745 OUT_N.t150 0.607167
R15630 OUT_N.n745 OUT_N.n744 0.607167
R15631 OUT_N.n739 OUT_N.t86 0.607167
R15632 OUT_N.n739 OUT_N.n738 0.607167
R15633 OUT_N.n733 OUT_N.t232 0.607167
R15634 OUT_N.n733 OUT_N.n732 0.607167
R15635 OUT_N.n727 OUT_N.t123 0.607167
R15636 OUT_N.n727 OUT_N.n726 0.607167
R15637 OUT_N.n721 OUT_N.t192 0.607167
R15638 OUT_N.n721 OUT_N.n720 0.607167
R15639 OUT_N.n619 OUT_N.t102 0.607167
R15640 OUT_N.n619 OUT_N.n618 0.607167
R15641 OUT_N.n625 OUT_N.t225 0.607167
R15642 OUT_N.n625 OUT_N.n624 0.607167
R15643 OUT_N.n631 OUT_N.t144 0.607167
R15644 OUT_N.n631 OUT_N.n630 0.607167
R15645 OUT_N.n637 OUT_N.t203 0.607167
R15646 OUT_N.n637 OUT_N.n636 0.607167
R15647 OUT_N.n643 OUT_N.t60 0.607167
R15648 OUT_N.n643 OUT_N.n642 0.607167
R15649 OUT_N.n649 OUT_N.t171 0.607167
R15650 OUT_N.n649 OUT_N.n648 0.607167
R15651 OUT_N.n655 OUT_N.t105 0.607167
R15652 OUT_N.n655 OUT_N.n654 0.607167
R15653 OUT_N.n661 OUT_N.t164 0.607167
R15654 OUT_N.n661 OUT_N.n660 0.607167
R15655 OUT_N.n667 OUT_N.t157 0.607167
R15656 OUT_N.n667 OUT_N.n666 0.607167
R15657 OUT_N.n673 OUT_N.t88 0.607167
R15658 OUT_N.n673 OUT_N.n672 0.607167
R15659 OUT_N.n679 OUT_N.t197 0.607167
R15660 OUT_N.n679 OUT_N.n678 0.607167
R15661 OUT_N.n685 OUT_N.t132 0.607167
R15662 OUT_N.n685 OUT_N.n684 0.607167
R15663 OUT_N.n691 OUT_N.t163 0.607167
R15664 OUT_N.n691 OUT_N.n690 0.607167
R15665 OUT_N.n697 OUT_N.t98 0.607167
R15666 OUT_N.n697 OUT_N.n696 0.607167
R15667 OUT_N.n703 OUT_N.t202 0.607167
R15668 OUT_N.n703 OUT_N.n702 0.607167
R15669 OUT_N.n709 OUT_N.t71 0.607167
R15670 OUT_N.n709 OUT_N.n708 0.607167
R15671 OUT_N.n715 OUT_N.t130 0.607167
R15672 OUT_N.n715 OUT_N.n714 0.607167
R15673 OUT_N.n1448 OUT_N.t182 0.607167
R15674 OUT_N.n1448 OUT_N.n1447 0.607167
R15675 OUT_N.n1442 OUT_N.t198 0.607167
R15676 OUT_N.n1442 OUT_N.n1441 0.607167
R15677 OUT_N.n1427 OUT_N.t81 0.607167
R15678 OUT_N.n1427 OUT_N.n1426 0.607167
R15679 OUT_N.n1421 OUT_N.t234 0.607167
R15680 OUT_N.n1421 OUT_N.n1420 0.607167
R15681 OUT_N.n1406 OUT_N.t127 0.607167
R15682 OUT_N.n1406 OUT_N.n1405 0.607167
R15683 OUT_N.n1400 OUT_N.t82 0.607167
R15684 OUT_N.n1400 OUT_N.n1399 0.607167
R15685 OUT_N.n1385 OUT_N.t221 0.607167
R15686 OUT_N.n1385 OUT_N.n1384 0.607167
R15687 OUT_N.n1379 OUT_N.t185 0.607167
R15688 OUT_N.n1379 OUT_N.n1378 0.607167
R15689 OUT_N.n1364 OUT_N.t209 0.607167
R15690 OUT_N.n1364 OUT_N.n1363 0.607167
R15691 OUT_N.n1358 OUT_N.t178 0.607167
R15692 OUT_N.n1358 OUT_N.n1357 0.607167
R15693 OUT_N.n1311 OUT_N.t122 0.607167
R15694 OUT_N.n1311 OUT_N.n1310 0.607167
R15695 OUT_N.n1317 OUT_N.t166 0.607167
R15696 OUT_N.n1317 OUT_N.n1316 0.607167
R15697 OUT_N.n1332 OUT_N.t78 0.607167
R15698 OUT_N.n1332 OUT_N.n1331 0.607167
R15699 OUT_N.n1338 OUT_N.t55 0.607167
R15700 OUT_N.n1338 OUT_N.n1337 0.607167
R15701 OUT_N.n1116 OUT_N.t154 0.607167
R15702 OUT_N.n1116 OUT_N.n1115 0.607167
R15703 OUT_N.n1110 OUT_N.t190 0.607167
R15704 OUT_N.n1110 OUT_N.n1109 0.607167
R15705 OUT_N.n1104 OUT_N.t217 0.607167
R15706 OUT_N.n1104 OUT_N.n1103 0.607167
R15707 OUT_N.n1098 OUT_N.t208 0.607167
R15708 OUT_N.n1098 OUT_N.n1097 0.607167
R15709 OUT_N.n1092 OUT_N.t173 0.607167
R15710 OUT_N.n1092 OUT_N.n1091 0.607167
R15711 OUT_N.n1086 OUT_N.t204 0.607167
R15712 OUT_N.n1086 OUT_N.n1085 0.607167
R15713 OUT_N.n1080 OUT_N.t48 0.607167
R15714 OUT_N.n1080 OUT_N.n1079 0.607167
R15715 OUT_N.n1074 OUT_N.t227 0.607167
R15716 OUT_N.n1074 OUT_N.n1073 0.607167
R15717 OUT_N.n1068 OUT_N.t172 0.607167
R15718 OUT_N.n1068 OUT_N.n1067 0.607167
R15719 OUT_N.n1062 OUT_N.t205 0.607167
R15720 OUT_N.n1062 OUT_N.n1061 0.607167
R15721 OUT_N.n1056 OUT_N.t242 0.607167
R15722 OUT_N.n1056 OUT_N.n1055 0.607167
R15723 OUT_N.n1050 OUT_N.t224 0.607167
R15724 OUT_N.n1050 OUT_N.n1049 0.607167
R15725 OUT_N.n1044 OUT_N.t235 0.607167
R15726 OUT_N.n1044 OUT_N.n1043 0.607167
R15727 OUT_N.n1038 OUT_N.t219 0.607167
R15728 OUT_N.n1038 OUT_N.n1037 0.607167
R15729 OUT_N.n1032 OUT_N.t64 0.607167
R15730 OUT_N.n1032 OUT_N.n1031 0.607167
R15731 OUT_N.n1026 OUT_N.t104 0.607167
R15732 OUT_N.n1026 OUT_N.n1025 0.607167
R15733 OUT_N.n1020 OUT_N.t195 0.607167
R15734 OUT_N.n1020 OUT_N.n1019 0.607167
R15735 OUT_N.n1014 OUT_N.t228 0.607167
R15736 OUT_N.n1014 OUT_N.n1013 0.607167
R15737 OUT_N.n1008 OUT_N.t74 0.607167
R15738 OUT_N.n1008 OUT_N.n1007 0.607167
R15739 OUT_N.n948 OUT_N.t128 0.607167
R15740 OUT_N.n948 OUT_N.n947 0.607167
R15741 OUT_N.n954 OUT_N.t94 0.607167
R15742 OUT_N.n954 OUT_N.n953 0.607167
R15743 OUT_N.n960 OUT_N.t52 0.607167
R15744 OUT_N.n960 OUT_N.n959 0.607167
R15745 OUT_N.n966 OUT_N.t67 0.607167
R15746 OUT_N.n966 OUT_N.n965 0.607167
R15747 OUT_N.n972 OUT_N.t129 0.607167
R15748 OUT_N.n972 OUT_N.n971 0.607167
R15749 OUT_N.n978 OUT_N.t93 0.607167
R15750 OUT_N.n978 OUT_N.n977 0.607167
R15751 OUT_N.n984 OUT_N.t54 0.607167
R15752 OUT_N.n984 OUT_N.n983 0.607167
R15753 OUT_N.n990 OUT_N.t69 0.607167
R15754 OUT_N.n990 OUT_N.n989 0.607167
R15755 OUT_N.n1002 OUT_N.t107 0.607167
R15756 OUT_N.n1002 OUT_N.n1001 0.607167
R15757 OUT_N.n299 OUT_N.t101 0.607167
R15758 OUT_N.n299 OUT_N.n298 0.607167
R15759 OUT_N.n293 OUT_N.t137 0.607167
R15760 OUT_N.n293 OUT_N.n292 0.607167
R15761 OUT_N.n278 OUT_N.t108 0.607167
R15762 OUT_N.n278 OUT_N.n277 0.607167
R15763 OUT_N.n272 OUT_N.t146 0.607167
R15764 OUT_N.n272 OUT_N.n271 0.607167
R15765 OUT_N.n257 OUT_N.t229 0.607167
R15766 OUT_N.n257 OUT_N.n256 0.607167
R15767 OUT_N.n251 OUT_N.t75 0.607167
R15768 OUT_N.n251 OUT_N.n250 0.607167
R15769 OUT_N.n236 OUT_N.t96 0.607167
R15770 OUT_N.n236 OUT_N.n235 0.607167
R15771 OUT_N.n230 OUT_N.t134 0.607167
R15772 OUT_N.n230 OUT_N.n229 0.607167
R15773 OUT_N.n215 OUT_N.t236 0.607167
R15774 OUT_N.n215 OUT_N.n214 0.607167
R15775 OUT_N.n209 OUT_N.t58 0.607167
R15776 OUT_N.n209 OUT_N.n208 0.607167
R15777 OUT_N.n194 OUT_N.t222 0.607167
R15778 OUT_N.n194 OUT_N.n193 0.607167
R15779 OUT_N.n188 OUT_N.t65 0.607167
R15780 OUT_N.n188 OUT_N.n187 0.607167
R15781 OUT_N.n546 OUT_N.t25 0.5465
R15782 OUT_N.n546 OUT_N.n545 0.5465
R15783 OUT_N.n2104 OUT_N.t264 0.5465
R15784 OUT_N.n2104 OUT_N.n2103 0.5465
R15785 OUT_N.n1870 OUT_N.t22 0.5465
R15786 OUT_N.n1870 OUT_N.n1869 0.5465
R15787 OUT_N.n1864 OUT_N.t46 0.5465
R15788 OUT_N.n1864 OUT_N.n1863 0.5465
R15789 OUT_N.n2098 OUT_N.t1 0.5465
R15790 OUT_N.n2098 OUT_N.n2097 0.5465
R15791 OUT_N.n2153 OUT_N.n2152 0.5465
R15792 OUT_N.n2074 OUT_N.n2073 0.5465
R15793 OUT_N.n1908 OUT_N.t9 0.5465
R15794 OUT_N.n1942 OUT_N.t35 0.5465
R15795 OUT_N.n1895 OUT_N.n1894 0.5465
R15796 OUT_N.n1964 OUT_N.n1963 0.5465
R15797 OUT_N.n1902 OUT_N.t3 0.5465
R15798 OUT_N.n1902 OUT_N.n1901 0.5465
R15799 OUT_N.n1938 OUT_N.t37 0.5465
R15800 OUT_N.n1938 OUT_N.n1937 0.5465
R15801 OUT_N.n2064 OUT_N.t43 0.5465
R15802 OUT_N.n2064 OUT_N.n2063 0.5465
R15803 OUT_N.n2142 OUT_N.t4 0.5465
R15804 OUT_N.n2142 OUT_N.n2141 0.5465
R15805 OUT_N.n2057 OUT_N.t258 0.5465
R15806 OUT_N.n2134 OUT_N.t26 0.5465
R15807 OUT_N.n2174 OUT_N.t10 0.5465
R15808 OUT_N.n2174 OUT_N.n2173 0.5465
R15809 OUT_N.n2186 OUT_N.t270 0.5465
R15810 OUT_N.n2186 OUT_N.n2185 0.5465
R15811 OUT_N.n1979 OUT_N.t41 0.5465
R15812 OUT_N.n1979 OUT_N.n1978 0.5465
R15813 OUT_N.n1984 OUT_N.t259 0.5465
R15814 OUT_N.n1984 OUT_N.n1983 0.5465
R15815 OUT_N.n527 OUT_N.t248 0.5465
R15816 OUT_N.n527 OUT_N.n526 0.5465
R15817 OUT_N.n512 OUT_N.t13 0.5465
R15818 OUT_N.n512 OUT_N.n511 0.5465
R15819 OUT_N.n9 OUT_N.t44 0.5465
R15820 OUT_N.n9 OUT_N.n8 0.5465
R15821 OUT_N.n14 OUT_N.t251 0.5465
R15822 OUT_N.n14 OUT_N.n13 0.5465
R15823 OUT_N.n1769 OUT_N.n1768 0.5465
R15824 OUT_N.n1707 OUT_N.t8 0.5465
R15825 OUT_N.n1707 OUT_N.n1706 0.5465
R15826 OUT_N.n1777 OUT_N.t17 0.5465
R15827 OUT_N.n1777 OUT_N.n1776 0.5465
R15828 OUT_N.n1695 OUT_N.t34 0.5465
R15829 OUT_N.n1785 OUT_N.t36 0.5465
R15830 OUT_N.n1718 OUT_N.n1717 0.5465
R15831 OUT_N.n1738 OUT_N.t31 0.5465
R15832 OUT_N.n1738 OUT_N.n1737 0.5465
R15833 OUT_N.n1743 OUT_N.t6 0.5465
R15834 OUT_N.n1743 OUT_N.n1742 0.5465
R15835 OUT_N.n1828 OUT_N.t265 0.5465
R15836 OUT_N.n1828 OUT_N.n1827 0.5465
R15837 OUT_N.n1843 OUT_N.t11 0.5465
R15838 OUT_N.n1843 OUT_N.n1842 0.5465
R15839 OUT_N.n2016 OUT_N.t12 0.5465
R15840 OUT_N.n2016 OUT_N.n2015 0.5465
R15841 OUT_N.n1518 OUT_N.n1517 0.482824
R15842 OUT_N.n1598 OUT_N.n1597 0.482824
R15843 OUT_N.n1651 OUT_N.n1650 0.482824
R15844 OUT_N.n383 OUT_N.n382 0.482824
R15845 OUT_N.n432 OUT_N.n431 0.482824
R15846 OUT_N.n485 OUT_N.n484 0.482824
R15847 OUT_N.n151 OUT_N.n150 0.469524
R15848 OUT_N.n92 OUT_N.n71 0.469524
R15849 OUT_N.n2193 OUT_N.n2192 0.468246
R15850 OUT_N.n1998 OUT_N.n1997 0.468246
R15851 OUT_N.n2117 OUT_N.n2115 0.468246
R15852 OUT_N.n1883 OUT_N.n1882 0.468246
R15853 OUT_N.n28 OUT_N.n27 0.468246
R15854 OUT_N.n1757 OUT_N.n1756 0.468246
R15855 OUT_N.n103 OUT_N.n102 0.4505
R15856 OUT_N.n84 OUT_N.n75 0.4505
R15857 OUT_N.n90 OUT_N.n74 0.4505
R15858 OUT_N.n65 OUT_N.n62 0.4505
R15859 OUT_N.n1297 OUT_N.n1296 0.43212
R15860 OUT_N.n938 OUT_N.n937 0.43212
R15861 OUT_N.n1195 OUT_N.n1194 0.431486
R15862 OUT_N.n848 OUT_N.n847 0.431486
R15863 OUT_N.n1241 OUT_N.n1240 0.428951
R15864 OUT_N.n892 OUT_N.n891 0.428951
R15865 OUT_N.n608 OUT_N.n607 0.428
R15866 OUT_N.n33 OUT_N.n32 0.428
R15867 OUT_N.n2237 OUT_N.n2236 0.428
R15868 OUT_N.n1137 OUT_N.n1136 0.415007
R15869 OUT_N.n1159 OUT_N.n1158 0.415007
R15870 OUT_N.n1261 OUT_N.n1260 0.415007
R15871 OUT_N.n802 OUT_N.n801 0.415007
R15872 OUT_N.n812 OUT_N.n811 0.415007
R15873 OUT_N.n902 OUT_N.n901 0.415007
R15874 OUT_N.n1205 OUT_N.n1204 0.408669
R15875 OUT_N.n856 OUT_N.n855 0.408669
R15876 OUT_N.n1547 OUT_N.n1546 0.395359
R15877 OUT_N.n613 OUT_N.n612 0.395359
R15878 OUT_N.n1465 OUT_N.n1464 0.389021
R15879 OUT_N.n1509 OUT_N.n1508 0.389021
R15880 OUT_N.n1527 OUT_N.n1526 0.389021
R15881 OUT_N.n1589 OUT_N.n1588 0.389021
R15882 OUT_N.n1607 OUT_N.n1606 0.389021
R15883 OUT_N.n1642 OUT_N.n1641 0.389021
R15884 OUT_N.n1660 OUT_N.n1659 0.389021
R15885 OUT_N.n337 OUT_N.n336 0.389021
R15886 OUT_N.n374 OUT_N.n373 0.389021
R15887 OUT_N.n392 OUT_N.n391 0.389021
R15888 OUT_N.n423 OUT_N.n422 0.389021
R15889 OUT_N.n441 OUT_N.n440 0.389021
R15890 OUT_N.n476 OUT_N.n475 0.389021
R15891 OUT_N.n494 OUT_N.n493 0.389021
R15892 OUT_N.n2089 OUT_N.n2088 0.366838
R15893 OUT_N.n1926 OUT_N.n1925 0.366838
R15894 OUT_N.n2168 OUT_N.n2167 0.366838
R15895 OUT_N.n1970 OUT_N.n1969 0.366838
R15896 OUT_N.n603 OUT_N.n602 0.366838
R15897 OUT_N.n576 OUT_N.n575 0.366838
R15898 OUT_N.n567 OUT_N.n566 0.366838
R15899 OUT_N.n1725 OUT_N.n1724 0.366838
R15900 OUT_N.n1803 OUT_N.n1802 0.366838
R15901 OUT_N.n2230 OUT_N.n2229 0.366838
R15902 OUT_N.n2203 OUT_N.n2202 0.366838
R15903 OUT_N.n2037 OUT_N.n2036 0.366838
R15904 OUT_N.n2000 OUT_N.n1976 0.356063
R15905 OUT_N.n1859 OUT_N.n1858 0.356063
R15906 OUT_N.n2195 OUT_N.n2171 0.356063
R15907 OUT_N.n1814 OUT_N.n1813 0.356063
R15908 OUT_N.n1730 OUT_N.n1729 0.356063
R15909 OUT_N.n1974 OUT_N.n1973 0.345923
R15910 OUT_N.n572 OUT_N.n571 0.345923
R15911 OUT_N.n2045 OUT_N.n2044 0.345923
R15912 OUT_N.n1904 OUT_N.n1900 0.336464
R15913 OUT_N.n2066 OUT_N.n2062 0.336464
R15914 OUT_N.n2055 OUT_N.n2054 0.336464
R15915 OUT_N.n2071 OUT_N.n2070 0.336464
R15916 OUT_N.n1779 OUT_N.n1775 0.336464
R15917 OUT_N.n1787 OUT_N.n1784 0.336464
R15918 OUT_N.n1771 OUT_N.n1767 0.336464
R15919 OUT_N.n1669 OUT_N.n1668 0.330394
R15920 OUT_N.n503 OUT_N.n502 0.330394
R15921 OUT_N.n1536 OUT_N.n1535 0.329761
R15922 OUT_N.n401 OUT_N.n400 0.329761
R15923 OUT_N.n1616 OUT_N.n1615 0.327225
R15924 OUT_N.n450 OUT_N.n449 0.327225
R15925 OUT_N.n1474 OUT_N.n1473 0.313282
R15926 OUT_N.n1500 OUT_N.n1499 0.313282
R15927 OUT_N.n1633 OUT_N.n1632 0.313282
R15928 OUT_N.n346 OUT_N.n345 0.313282
R15929 OUT_N.n365 OUT_N.n364 0.313282
R15930 OUT_N.n467 OUT_N.n466 0.313282
R15931 OUT_N.n1580 OUT_N.n1579 0.306944
R15932 OUT_N.n414 OUT_N.n413 0.306944
R15933 OUT_N.n999 OUT_N.n998 0.2705
R15934 OUT_N.n1256 OUT_N.n1255 0.2705
R15935 OUT_N.n1552 OUT_N.n1551 0.2705
R15936 OUT_N.n1569 OUT_N.n1568 0.2705
R15937 OUT_N.n1145 OUT_N.n1144 0.2705
R15938 OUT_N.n1156 OUT_N.n1155 0.2705
R15939 OUT_N.n943 OUT_N.n942 0.2705
R15940 OUT_N.n1677 OUT_N.n1673 0.238176
R15941 OUT_N.n1930 OUT_N.n1929 0.231204
R15942 OUT_N.n2128 OUT_N.n2127 0.231204
R15943 OUT_N.n1809 OUT_N.n1805 0.231204
R15944 OUT_N.n1910 OUT_N.n1907 0.191654
R15945 OUT_N.n1892 OUT_N.n1891 0.191654
R15946 OUT_N.n2080 OUT_N.n2079 0.186204
R15947 OUT_N.n2085 OUT_N.n2084 0.186204
R15948 OUT_N.n1922 OUT_N.n1921 0.186204
R15949 OUT_N.n1917 OUT_N.n1916 0.186204
R15950 OUT_N.n2158 OUT_N.n2157 0.186204
R15951 OUT_N.n2163 OUT_N.n2162 0.186204
R15952 OUT_N.n1958 OUT_N.n1957 0.186204
R15953 OUT_N.n1953 OUT_N.n1952 0.186204
R15954 OUT_N.n2182 OUT_N.n2181 0.186204
R15955 OUT_N.n1993 OUT_N.n1992 0.186204
R15956 OUT_N.n2112 OUT_N.n2111 0.186204
R15957 OUT_N.n1878 OUT_N.n1877 0.186204
R15958 OUT_N.n1124 OUT_N.n1123 0.186204
R15959 OUT_N.n1128 OUT_N.n1127 0.186204
R15960 OUT_N.n1133 OUT_N.n1132 0.186204
R15961 OUT_N.n1164 OUT_N.n1163 0.186204
R15962 OUT_N.n1168 OUT_N.n1167 0.186204
R15963 OUT_N.n1173 OUT_N.n1172 0.186204
R15964 OUT_N.n1182 OUT_N.n1181 0.186204
R15965 OUT_N.n1186 OUT_N.n1185 0.186204
R15966 OUT_N.n1191 OUT_N.n1190 0.186204
R15967 OUT_N.n1210 OUT_N.n1209 0.186204
R15968 OUT_N.n1214 OUT_N.n1213 0.186204
R15969 OUT_N.n1219 OUT_N.n1218 0.186204
R15970 OUT_N.n1228 OUT_N.n1227 0.186204
R15971 OUT_N.n1232 OUT_N.n1231 0.186204
R15972 OUT_N.n1237 OUT_N.n1236 0.186204
R15973 OUT_N.n1266 OUT_N.n1265 0.186204
R15974 OUT_N.n1270 OUT_N.n1269 0.186204
R15975 OUT_N.n1275 OUT_N.n1274 0.186204
R15976 OUT_N.n1284 OUT_N.n1283 0.186204
R15977 OUT_N.n1288 OUT_N.n1287 0.186204
R15978 OUT_N.n1293 OUT_N.n1292 0.186204
R15979 OUT_N.n1461 OUT_N.n1460 0.186204
R15980 OUT_N.n1470 OUT_N.n1469 0.186204
R15981 OUT_N.n1505 OUT_N.n1504 0.186204
R15982 OUT_N.n1514 OUT_N.n1513 0.186204
R15983 OUT_N.n1523 OUT_N.n1522 0.186204
R15984 OUT_N.n1532 OUT_N.n1531 0.186204
R15985 OUT_N.n1585 OUT_N.n1584 0.186204
R15986 OUT_N.n1594 OUT_N.n1593 0.186204
R15987 OUT_N.n1603 OUT_N.n1602 0.186204
R15988 OUT_N.n1612 OUT_N.n1611 0.186204
R15989 OUT_N.n1638 OUT_N.n1637 0.186204
R15990 OUT_N.n1647 OUT_N.n1646 0.186204
R15991 OUT_N.n1656 OUT_N.n1655 0.186204
R15992 OUT_N.n1665 OUT_N.n1664 0.186204
R15993 OUT_N.n789 OUT_N.n788 0.186204
R15994 OUT_N.n793 OUT_N.n792 0.186204
R15995 OUT_N.n798 OUT_N.n797 0.186204
R15996 OUT_N.n817 OUT_N.n816 0.186204
R15997 OUT_N.n821 OUT_N.n820 0.186204
R15998 OUT_N.n826 OUT_N.n825 0.186204
R15999 OUT_N.n835 OUT_N.n834 0.186204
R16000 OUT_N.n839 OUT_N.n838 0.186204
R16001 OUT_N.n844 OUT_N.n843 0.186204
R16002 OUT_N.n861 OUT_N.n860 0.186204
R16003 OUT_N.n865 OUT_N.n864 0.186204
R16004 OUT_N.n870 OUT_N.n869 0.186204
R16005 OUT_N.n879 OUT_N.n878 0.186204
R16006 OUT_N.n883 OUT_N.n882 0.186204
R16007 OUT_N.n888 OUT_N.n887 0.186204
R16008 OUT_N.n907 OUT_N.n906 0.186204
R16009 OUT_N.n911 OUT_N.n910 0.186204
R16010 OUT_N.n916 OUT_N.n915 0.186204
R16011 OUT_N.n925 OUT_N.n924 0.186204
R16012 OUT_N.n929 OUT_N.n928 0.186204
R16013 OUT_N.n934 OUT_N.n933 0.186204
R16014 OUT_N.n333 OUT_N.n332 0.186204
R16015 OUT_N.n342 OUT_N.n341 0.186204
R16016 OUT_N.n370 OUT_N.n369 0.186204
R16017 OUT_N.n379 OUT_N.n378 0.186204
R16018 OUT_N.n388 OUT_N.n387 0.186204
R16019 OUT_N.n397 OUT_N.n396 0.186204
R16020 OUT_N.n419 OUT_N.n418 0.186204
R16021 OUT_N.n428 OUT_N.n427 0.186204
R16022 OUT_N.n437 OUT_N.n436 0.186204
R16023 OUT_N.n446 OUT_N.n445 0.186204
R16024 OUT_N.n472 OUT_N.n471 0.186204
R16025 OUT_N.n481 OUT_N.n480 0.186204
R16026 OUT_N.n490 OUT_N.n489 0.186204
R16027 OUT_N.n499 OUT_N.n498 0.186204
R16028 OUT_N.n599 OUT_N.n598 0.186204
R16029 OUT_N.n594 OUT_N.n593 0.186204
R16030 OUT_N.n585 OUT_N.n584 0.186204
R16031 OUT_N.n581 OUT_N.n580 0.186204
R16032 OUT_N.n563 OUT_N.n562 0.186204
R16033 OUT_N.n558 OUT_N.n557 0.186204
R16034 OUT_N.n23 OUT_N.n22 0.186204
R16035 OUT_N.n1712 OUT_N.n1711 0.186204
R16036 OUT_N.n1703 OUT_N.n1702 0.186204
R16037 OUT_N.n1798 OUT_N.n1797 0.186204
R16038 OUT_N.n1793 OUT_N.n1792 0.186204
R16039 OUT_N.n1752 OUT_N.n1751 0.186204
R16040 OUT_N.n2225 OUT_N.n2224 0.186204
R16041 OUT_N.n2221 OUT_N.n2220 0.186204
R16042 OUT_N.n2212 OUT_N.n2211 0.186204
R16043 OUT_N.n2207 OUT_N.n2206 0.186204
R16044 OUT_N.n2032 OUT_N.n2031 0.186204
R16045 OUT_N.n2028 OUT_N.n2027 0.186204
R16046 OUT_N.n1148 OUT_N.n1147 0.176697
R16047 OUT_N.n1487 OUT_N.n1486 0.176697
R16048 OUT_N.n807 OUT_N.n806 0.176697
R16049 OUT_N.n356 OUT_N.n355 0.176697
R16050 OUT_N.n1200 OUT_N.n1199 0.166556
R16051 OUT_N.n1560 OUT_N.n1559 0.166556
R16052 OUT_N.n853 OUT_N.n852 0.166556
R16053 OUT_N.n406 OUT_N.n405 0.166556
R16054 OUT_N.n1246 OUT_N.n1245 0.162754
R16055 OUT_N.n1629 OUT_N.n1628 0.162754
R16056 OUT_N.n897 OUT_N.n896 0.162754
R16057 OUT_N.n458 OUT_N.n457 0.162754
R16058 OUT_N.n1626 OUT_N.n1625 0.145641
R16059 OUT_N.n1557 OUT_N.n1556 0.145641
R16060 OUT_N.n1574 OUT_N.n1573 0.145641
R16061 OUT_N.n1481 OUT_N.n1480 0.145641
R16062 OUT_N.n1497 OUT_N.n1496 0.145641
R16063 OUT_N.n1302 OUT_N.n1301 0.145641
R16064 OUT_N.n1910 OUT_N.n1909 0.106363
R16065 OUT_N.n2008 OUT_N.n2007 0.106345
R16066 OUT_N.n1886 OUT_N.n1885 0.106345
R16067 OUT_N.n2200 OUT_N.n2199 0.106345
R16068 OUT_N.n2123 OUT_N.n2122 0.106345
R16069 OUT_N.n1820 OUT_N.n1818 0.106345
R16070 OUT_N.n1760 OUT_N.n1759 0.106345
R16071 OUT_N.n1682 OUT_N.n1681 0.106345
R16072 OUT_N.n169 OUT_N.n105 0.105505
R16073 OUT_N.n2189 OUT_N.n2184 0.0992756
R16074 OUT_N.n1982 OUT_N.n1977 0.0992756
R16075 OUT_N.n12 OUT_N.n7 0.0992756
R16076 OUT_N.n1721 OUT_N.n1716 0.0992756
R16077 OUT_N.n1741 OUT_N.n1736 0.0992756
R16078 OUT_N OUT_N.n2242 0.0835282
R16079 OUT_N.n1913 OUT_N.n1912 0.0832399
R16080 OUT_N.n1699 OUT_N.n1694 0.0832399
R16081 OUT_N.n2023 OUT_N.n2021 0.0832399
R16082 OUT_N.n2178 OUT_N.n2177 0.0831446
R16083 OUT_N.n1906 OUT_N.n1899 0.0824117
R16084 OUT_N.n1773 OUT_N.n1766 0.0824117
R16085 OUT_N.n328 OUT_N.n324 0.0823987
R16086 OUT_N.n317 OUT_N.n312 0.0823987
R16087 OUT_N.n549 OUT_N.n544 0.0823987
R16088 OUT_N.n2107 OUT_N.n2102 0.0823987
R16089 OUT_N.n1867 OUT_N.n1862 0.0823987
R16090 OUT_N.n1941 OUT_N.n1936 0.0823987
R16091 OUT_N.n2145 OUT_N.n2140 0.0823987
R16092 OUT_N.n2068 OUT_N.n2061 0.0823987
R16093 OUT_N.n2137 OUT_N.n2133 0.0823987
R16094 OUT_N.n534 OUT_N.n531 0.0823987
R16095 OUT_N.n524 OUT_N.n520 0.0823987
R16096 OUT_N.n515 OUT_N.n510 0.0823987
R16097 OUT_N.n784 OUT_N.n779 0.0823987
R16098 OUT_N.n772 OUT_N.n767 0.0823987
R16099 OUT_N.n760 OUT_N.n755 0.0823987
R16100 OUT_N.n748 OUT_N.n743 0.0823987
R16101 OUT_N.n736 OUT_N.n731 0.0823987
R16102 OUT_N.n724 OUT_N.n719 0.0823987
R16103 OUT_N.n628 OUT_N.n623 0.0823987
R16104 OUT_N.n640 OUT_N.n635 0.0823987
R16105 OUT_N.n652 OUT_N.n647 0.0823987
R16106 OUT_N.n664 OUT_N.n659 0.0823987
R16107 OUT_N.n676 OUT_N.n671 0.0823987
R16108 OUT_N.n688 OUT_N.n683 0.0823987
R16109 OUT_N.n700 OUT_N.n695 0.0823987
R16110 OUT_N.n712 OUT_N.n707 0.0823987
R16111 OUT_N.n1456 OUT_N.n1452 0.0823987
R16112 OUT_N.n1445 OUT_N.n1440 0.0823987
R16113 OUT_N.n1435 OUT_N.n1431 0.0823987
R16114 OUT_N.n1424 OUT_N.n1419 0.0823987
R16115 OUT_N.n1414 OUT_N.n1410 0.0823987
R16116 OUT_N.n1403 OUT_N.n1398 0.0823987
R16117 OUT_N.n1393 OUT_N.n1389 0.0823987
R16118 OUT_N.n1382 OUT_N.n1377 0.0823987
R16119 OUT_N.n1372 OUT_N.n1368 0.0823987
R16120 OUT_N.n1361 OUT_N.n1356 0.0823987
R16121 OUT_N.n1314 OUT_N.n1309 0.0823987
R16122 OUT_N.n1325 OUT_N.n1321 0.0823987
R16123 OUT_N.n1335 OUT_N.n1330 0.0823987
R16124 OUT_N.n1346 OUT_N.n1342 0.0823987
R16125 OUT_N.n1119 OUT_N.n1114 0.0823987
R16126 OUT_N.n1107 OUT_N.n1102 0.0823987
R16127 OUT_N.n1095 OUT_N.n1090 0.0823987
R16128 OUT_N.n1083 OUT_N.n1078 0.0823987
R16129 OUT_N.n1071 OUT_N.n1066 0.0823987
R16130 OUT_N.n1059 OUT_N.n1054 0.0823987
R16131 OUT_N.n1047 OUT_N.n1042 0.0823987
R16132 OUT_N.n1035 OUT_N.n1030 0.0823987
R16133 OUT_N.n1023 OUT_N.n1018 0.0823987
R16134 OUT_N.n1011 OUT_N.n1006 0.0823987
R16135 OUT_N.n957 OUT_N.n952 0.0823987
R16136 OUT_N.n969 OUT_N.n964 0.0823987
R16137 OUT_N.n981 OUT_N.n976 0.0823987
R16138 OUT_N.n993 OUT_N.n988 0.0823987
R16139 OUT_N.n307 OUT_N.n303 0.0823987
R16140 OUT_N.n296 OUT_N.n291 0.0823987
R16141 OUT_N.n286 OUT_N.n282 0.0823987
R16142 OUT_N.n275 OUT_N.n270 0.0823987
R16143 OUT_N.n265 OUT_N.n261 0.0823987
R16144 OUT_N.n254 OUT_N.n249 0.0823987
R16145 OUT_N.n244 OUT_N.n240 0.0823987
R16146 OUT_N.n233 OUT_N.n228 0.0823987
R16147 OUT_N.n223 OUT_N.n219 0.0823987
R16148 OUT_N.n212 OUT_N.n207 0.0823987
R16149 OUT_N.n202 OUT_N.n198 0.0823987
R16150 OUT_N.n191 OUT_N.n186 0.0823987
R16151 OUT_N.n1781 OUT_N.n1774 0.0823987
R16152 OUT_N.n1825 OUT_N.n1821 0.0823987
R16153 OUT_N.n1835 OUT_N.n1832 0.0823987
R16154 OUT_N.n1846 OUT_N.n1841 0.0823987
R16155 OUT_N.n2013 OUT_N.n2009 0.0823987
R16156 OUT_N.n1698 OUT_N.n1697 0.0817926
R16157 OUT_N.n1904 OUT_N.n1903 0.0748144
R16158 OUT_N.n2066 OUT_N.n2065 0.0748144
R16159 OUT_N.n1779 OUT_N.n1778 0.0748144
R16160 OUT_N.n1787 OUT_N.n1786 0.0748144
R16161 OUT_N.n1771 OUT_N.n1770 0.0748144
R16162 OUT_N.n2060 OUT_N.n2056 0.0712285
R16163 OUT_N.n1898 OUT_N.n1893 0.0712285
R16164 OUT_N.n2077 OUT_N.n2072 0.0712285
R16165 OUT_N.n1948 OUT_N.n1944 0.0712285
R16166 OUT_N.n2101 OUT_N.n2096 0.0712285
R16167 OUT_N.n1873 OUT_N.n1868 0.0712285
R16168 OUT_N.n1005 OUT_N.n1000 0.0712285
R16169 OUT_N.n987 OUT_N.n982 0.0712285
R16170 OUT_N.n975 OUT_N.n970 0.0712285
R16171 OUT_N.n963 OUT_N.n958 0.0712285
R16172 OUT_N.n951 OUT_N.n946 0.0712285
R16173 OUT_N.n1017 OUT_N.n1012 0.0712285
R16174 OUT_N.n1029 OUT_N.n1024 0.0712285
R16175 OUT_N.n1041 OUT_N.n1036 0.0712285
R16176 OUT_N.n1053 OUT_N.n1048 0.0712285
R16177 OUT_N.n1065 OUT_N.n1060 0.0712285
R16178 OUT_N.n1077 OUT_N.n1072 0.0712285
R16179 OUT_N.n1089 OUT_N.n1084 0.0712285
R16180 OUT_N.n1101 OUT_N.n1096 0.0712285
R16181 OUT_N.n1113 OUT_N.n1108 0.0712285
R16182 OUT_N.n1355 OUT_N.n1352 0.0712285
R16183 OUT_N.n1341 OUT_N.n1336 0.0712285
R16184 OUT_N.n1329 OUT_N.n1326 0.0712285
R16185 OUT_N.n1320 OUT_N.n1315 0.0712285
R16186 OUT_N.n1308 OUT_N.n1305 0.0712285
R16187 OUT_N.n1367 OUT_N.n1362 0.0712285
R16188 OUT_N.n1376 OUT_N.n1373 0.0712285
R16189 OUT_N.n1388 OUT_N.n1383 0.0712285
R16190 OUT_N.n1397 OUT_N.n1394 0.0712285
R16191 OUT_N.n1409 OUT_N.n1404 0.0712285
R16192 OUT_N.n1418 OUT_N.n1415 0.0712285
R16193 OUT_N.n1430 OUT_N.n1425 0.0712285
R16194 OUT_N.n1439 OUT_N.n1436 0.0712285
R16195 OUT_N.n1451 OUT_N.n1446 0.0712285
R16196 OUT_N.n718 OUT_N.n713 0.0712285
R16197 OUT_N.n706 OUT_N.n701 0.0712285
R16198 OUT_N.n694 OUT_N.n689 0.0712285
R16199 OUT_N.n682 OUT_N.n677 0.0712285
R16200 OUT_N.n670 OUT_N.n665 0.0712285
R16201 OUT_N.n658 OUT_N.n653 0.0712285
R16202 OUT_N.n646 OUT_N.n641 0.0712285
R16203 OUT_N.n634 OUT_N.n629 0.0712285
R16204 OUT_N.n622 OUT_N.n617 0.0712285
R16205 OUT_N.n730 OUT_N.n725 0.0712285
R16206 OUT_N.n742 OUT_N.n737 0.0712285
R16207 OUT_N.n754 OUT_N.n749 0.0712285
R16208 OUT_N.n766 OUT_N.n761 0.0712285
R16209 OUT_N.n778 OUT_N.n773 0.0712285
R16210 OUT_N.n185 OUT_N.n182 0.0712285
R16211 OUT_N.n197 OUT_N.n192 0.0712285
R16212 OUT_N.n206 OUT_N.n203 0.0712285
R16213 OUT_N.n218 OUT_N.n213 0.0712285
R16214 OUT_N.n227 OUT_N.n224 0.0712285
R16215 OUT_N.n239 OUT_N.n234 0.0712285
R16216 OUT_N.n248 OUT_N.n245 0.0712285
R16217 OUT_N.n260 OUT_N.n255 0.0712285
R16218 OUT_N.n269 OUT_N.n266 0.0712285
R16219 OUT_N.n281 OUT_N.n276 0.0712285
R16220 OUT_N.n290 OUT_N.n287 0.0712285
R16221 OUT_N.n302 OUT_N.n297 0.0712285
R16222 OUT_N.n311 OUT_N.n308 0.0712285
R16223 OUT_N.n509 OUT_N.n505 0.0712285
R16224 OUT_N.n519 OUT_N.n516 0.0712285
R16225 OUT_N.n530 OUT_N.n525 0.0712285
R16226 OUT_N.n543 OUT_N.n539 0.0712285
R16227 OUT_N.n553 OUT_N.n550 0.0712285
R16228 OUT_N.n323 OUT_N.n318 0.0712285
R16229 OUT_N.n2019 OUT_N.n2014 0.0712285
R16230 OUT_N.n1850 OUT_N.n1847 0.0712285
R16231 OUT_N.n1840 OUT_N.n1836 0.0712285
R16232 OUT_N.n1831 OUT_N.n1826 0.0712285
R16233 OUT_N.n1967 OUT_N.n1966 0.0709833
R16234 OUT_N.n147 OUT_N.n146 0.0707439
R16235 OUT_N.n68 OUT_N.n67 0.0707439
R16236 OUT_N.n1988 OUT_N.n1987 0.0623855
R16237 OUT_N.n1987 OUT_N.n1986 0.0623855
R16238 OUT_N.n18 OUT_N.n17 0.0623855
R16239 OUT_N.n17 OUT_N.n16 0.0623855
R16240 OUT_N.n1788 OUT_N.n1783 0.0623855
R16241 OUT_N.n1783 OUT_N.n1782 0.0623855
R16242 OUT_N.n1747 OUT_N.n1746 0.0623855
R16243 OUT_N.n1746 OUT_N.n1745 0.0623855
R16244 OUT_N.n1967 OUT_N.n1962 0.0536862
R16245 OUT_N.n1898 OUT_N.n1897 0.0534597
R16246 OUT_N.n2077 OUT_N.n2076 0.0534597
R16247 OUT_N.n2060 OUT_N.n2059 0.0534597
R16248 OUT_N.n1948 OUT_N.n1947 0.0534597
R16249 OUT_N.n1873 OUT_N.n1872 0.0534597
R16250 OUT_N.n2101 OUT_N.n2100 0.0534597
R16251 OUT_N.n951 OUT_N.n950 0.0534597
R16252 OUT_N.n963 OUT_N.n962 0.0534597
R16253 OUT_N.n975 OUT_N.n974 0.0534597
R16254 OUT_N.n987 OUT_N.n986 0.0534597
R16255 OUT_N.n1113 OUT_N.n1112 0.0534597
R16256 OUT_N.n1101 OUT_N.n1100 0.0534597
R16257 OUT_N.n1089 OUT_N.n1088 0.0534597
R16258 OUT_N.n1077 OUT_N.n1076 0.0534597
R16259 OUT_N.n1065 OUT_N.n1064 0.0534597
R16260 OUT_N.n1053 OUT_N.n1052 0.0534597
R16261 OUT_N.n1041 OUT_N.n1040 0.0534597
R16262 OUT_N.n1029 OUT_N.n1028 0.0534597
R16263 OUT_N.n1017 OUT_N.n1016 0.0534597
R16264 OUT_N.n1005 OUT_N.n1004 0.0534597
R16265 OUT_N.n1308 OUT_N.n1307 0.0534597
R16266 OUT_N.n1320 OUT_N.n1319 0.0534597
R16267 OUT_N.n1329 OUT_N.n1328 0.0534597
R16268 OUT_N.n1341 OUT_N.n1340 0.0534597
R16269 OUT_N.n1451 OUT_N.n1450 0.0534597
R16270 OUT_N.n1439 OUT_N.n1438 0.0534597
R16271 OUT_N.n1430 OUT_N.n1429 0.0534597
R16272 OUT_N.n1418 OUT_N.n1417 0.0534597
R16273 OUT_N.n1409 OUT_N.n1408 0.0534597
R16274 OUT_N.n1397 OUT_N.n1396 0.0534597
R16275 OUT_N.n1388 OUT_N.n1387 0.0534597
R16276 OUT_N.n1376 OUT_N.n1375 0.0534597
R16277 OUT_N.n1367 OUT_N.n1366 0.0534597
R16278 OUT_N.n1355 OUT_N.n1354 0.0534597
R16279 OUT_N.n622 OUT_N.n621 0.0534597
R16280 OUT_N.n634 OUT_N.n633 0.0534597
R16281 OUT_N.n646 OUT_N.n645 0.0534597
R16282 OUT_N.n658 OUT_N.n657 0.0534597
R16283 OUT_N.n670 OUT_N.n669 0.0534597
R16284 OUT_N.n682 OUT_N.n681 0.0534597
R16285 OUT_N.n694 OUT_N.n693 0.0534597
R16286 OUT_N.n706 OUT_N.n705 0.0534597
R16287 OUT_N.n778 OUT_N.n777 0.0534597
R16288 OUT_N.n766 OUT_N.n765 0.0534597
R16289 OUT_N.n754 OUT_N.n753 0.0534597
R16290 OUT_N.n742 OUT_N.n741 0.0534597
R16291 OUT_N.n730 OUT_N.n729 0.0534597
R16292 OUT_N.n718 OUT_N.n717 0.0534597
R16293 OUT_N.n553 OUT_N.n552 0.0534597
R16294 OUT_N.n543 OUT_N.n542 0.0534597
R16295 OUT_N.n530 OUT_N.n529 0.0534597
R16296 OUT_N.n519 OUT_N.n518 0.0534597
R16297 OUT_N.n509 OUT_N.n508 0.0534597
R16298 OUT_N.n323 OUT_N.n322 0.0534597
R16299 OUT_N.n311 OUT_N.n310 0.0534597
R16300 OUT_N.n302 OUT_N.n301 0.0534597
R16301 OUT_N.n290 OUT_N.n289 0.0534597
R16302 OUT_N.n281 OUT_N.n280 0.0534597
R16303 OUT_N.n269 OUT_N.n268 0.0534597
R16304 OUT_N.n260 OUT_N.n259 0.0534597
R16305 OUT_N.n248 OUT_N.n247 0.0534597
R16306 OUT_N.n239 OUT_N.n238 0.0534597
R16307 OUT_N.n227 OUT_N.n226 0.0534597
R16308 OUT_N.n218 OUT_N.n217 0.0534597
R16309 OUT_N.n206 OUT_N.n205 0.0534597
R16310 OUT_N.n197 OUT_N.n196 0.0534597
R16311 OUT_N.n185 OUT_N.n184 0.0534597
R16312 OUT_N.n1831 OUT_N.n1830 0.0534597
R16313 OUT_N.n1840 OUT_N.n1839 0.0534597
R16314 OUT_N.n1850 OUT_N.n1849 0.0534597
R16315 OUT_N.n2019 OUT_N.n2018 0.0534597
R16316 OUT_N.n2177 OUT_N.n2176 0.0420655
R16317 OUT_N.n1912 OUT_N.n1911 0.0419676
R16318 OUT_N.n1694 OUT_N.n1693 0.0419676
R16319 OUT_N.n2021 OUT_N.n2020 0.0419676
R16320 OUT_N.n2068 OUT_N.n2067 0.0415773
R16321 OUT_N.n1941 OUT_N.n1940 0.0415773
R16322 OUT_N.n2145 OUT_N.n2144 0.0415773
R16323 OUT_N.n2137 OUT_N.n2136 0.0415773
R16324 OUT_N.n1867 OUT_N.n1866 0.0415773
R16325 OUT_N.n2107 OUT_N.n2106 0.0415773
R16326 OUT_N.n993 OUT_N.n992 0.0415773
R16327 OUT_N.n981 OUT_N.n980 0.0415773
R16328 OUT_N.n969 OUT_N.n968 0.0415773
R16329 OUT_N.n957 OUT_N.n956 0.0415773
R16330 OUT_N.n1011 OUT_N.n1010 0.0415773
R16331 OUT_N.n1023 OUT_N.n1022 0.0415773
R16332 OUT_N.n1035 OUT_N.n1034 0.0415773
R16333 OUT_N.n1047 OUT_N.n1046 0.0415773
R16334 OUT_N.n1059 OUT_N.n1058 0.0415773
R16335 OUT_N.n1071 OUT_N.n1070 0.0415773
R16336 OUT_N.n1083 OUT_N.n1082 0.0415773
R16337 OUT_N.n1095 OUT_N.n1094 0.0415773
R16338 OUT_N.n1107 OUT_N.n1106 0.0415773
R16339 OUT_N.n1119 OUT_N.n1118 0.0415773
R16340 OUT_N.n1346 OUT_N.n1345 0.0415773
R16341 OUT_N.n1335 OUT_N.n1334 0.0415773
R16342 OUT_N.n1325 OUT_N.n1324 0.0415773
R16343 OUT_N.n1314 OUT_N.n1313 0.0415773
R16344 OUT_N.n1361 OUT_N.n1360 0.0415773
R16345 OUT_N.n1372 OUT_N.n1371 0.0415773
R16346 OUT_N.n1382 OUT_N.n1381 0.0415773
R16347 OUT_N.n1393 OUT_N.n1392 0.0415773
R16348 OUT_N.n1403 OUT_N.n1402 0.0415773
R16349 OUT_N.n1414 OUT_N.n1413 0.0415773
R16350 OUT_N.n1424 OUT_N.n1423 0.0415773
R16351 OUT_N.n1435 OUT_N.n1434 0.0415773
R16352 OUT_N.n1445 OUT_N.n1444 0.0415773
R16353 OUT_N.n1456 OUT_N.n1455 0.0415773
R16354 OUT_N.n712 OUT_N.n711 0.0415773
R16355 OUT_N.n700 OUT_N.n699 0.0415773
R16356 OUT_N.n688 OUT_N.n687 0.0415773
R16357 OUT_N.n676 OUT_N.n675 0.0415773
R16358 OUT_N.n664 OUT_N.n663 0.0415773
R16359 OUT_N.n652 OUT_N.n651 0.0415773
R16360 OUT_N.n640 OUT_N.n639 0.0415773
R16361 OUT_N.n628 OUT_N.n627 0.0415773
R16362 OUT_N.n724 OUT_N.n723 0.0415773
R16363 OUT_N.n736 OUT_N.n735 0.0415773
R16364 OUT_N.n748 OUT_N.n747 0.0415773
R16365 OUT_N.n760 OUT_N.n759 0.0415773
R16366 OUT_N.n772 OUT_N.n771 0.0415773
R16367 OUT_N.n784 OUT_N.n783 0.0415773
R16368 OUT_N.n191 OUT_N.n190 0.0415773
R16369 OUT_N.n202 OUT_N.n201 0.0415773
R16370 OUT_N.n212 OUT_N.n211 0.0415773
R16371 OUT_N.n223 OUT_N.n222 0.0415773
R16372 OUT_N.n233 OUT_N.n232 0.0415773
R16373 OUT_N.n244 OUT_N.n243 0.0415773
R16374 OUT_N.n254 OUT_N.n253 0.0415773
R16375 OUT_N.n265 OUT_N.n264 0.0415773
R16376 OUT_N.n275 OUT_N.n274 0.0415773
R16377 OUT_N.n286 OUT_N.n285 0.0415773
R16378 OUT_N.n296 OUT_N.n295 0.0415773
R16379 OUT_N.n307 OUT_N.n306 0.0415773
R16380 OUT_N.n515 OUT_N.n514 0.0415773
R16381 OUT_N.n524 OUT_N.n523 0.0415773
R16382 OUT_N.n534 OUT_N.n533 0.0415773
R16383 OUT_N.n549 OUT_N.n548 0.0415773
R16384 OUT_N.n317 OUT_N.n316 0.0415773
R16385 OUT_N.n328 OUT_N.n327 0.0415773
R16386 OUT_N.n1781 OUT_N.n1780 0.0415773
R16387 OUT_N.n2013 OUT_N.n2012 0.0415773
R16388 OUT_N.n1846 OUT_N.n1845 0.0415773
R16389 OUT_N.n1835 OUT_N.n1834 0.0415773
R16390 OUT_N.n1825 OUT_N.n1824 0.0415773
R16391 OUT_N.n1906 OUT_N.n1905 0.0415636
R16392 OUT_N.n1773 OUT_N.n1772 0.0415636
R16393 OUT_N.n1946 OUT_N.n1945 0.0383947
R16394 OUT_N.n1961 OUT_N.n1960 0.0383947
R16395 OUT_N.n2132 OUT_N.n2131 0.0383947
R16396 OUT_N.n2148 OUT_N.n2147 0.0383947
R16397 OUT_N.n1697 OUT_N.n1696 0.0383947
R16398 OUT_N.n1715 OUT_N.n1714 0.0383947
R16399 OUT_N.n2092 OUT_N.n2089 0.0334577
R16400 OUT_N.n1927 OUT_N.n1926 0.0334577
R16401 OUT_N.n2169 OUT_N.n2168 0.0334577
R16402 OUT_N.n1147 OUT_N.n1139 0.0334577
R16403 OUT_N.n1158 OUT_N.n1150 0.0334577
R16404 OUT_N.n1299 OUT_N.n1297 0.0334577
R16405 OUT_N.n1299 OUT_N.n1298 0.0334577
R16406 OUT_N.n1559 OUT_N.n1540 0.0334577
R16407 OUT_N.n1628 OUT_N.n1620 0.0334577
R16408 OUT_N.n1632 OUT_N.n1631 0.0334577
R16409 OUT_N.n1671 OUT_N.n1669 0.0334577
R16410 OUT_N.n1671 OUT_N.n1670 0.0334577
R16411 OUT_N.n854 OUT_N.n853 0.0334577
R16412 OUT_N.n855 OUT_N.n854 0.0334577
R16413 OUT_N.n939 OUT_N.n938 0.0334577
R16414 OUT_N.n413 OUT_N.n410 0.0334577
R16415 OUT_N.n457 OUT_N.n454 0.0334577
R16416 OUT_N.n575 OUT_N.n574 0.0334577
R16417 OUT_N.n1727 OUT_N.n1726 0.0334577
R16418 OUT_N.n1692 OUT_N.n1691 0.0319869
R16419 OUT_N.n67 OUT_N.t253 0.0306947
R16420 OUT_N.n146 OUT_N.t254 0.0285465
R16421 OUT_N.n1982 OUT_N.n1981 0.0254881
R16422 OUT_N.n2189 OUT_N.n2188 0.0254881
R16423 OUT_N.n12 OUT_N.n11 0.0254881
R16424 OUT_N.n1721 OUT_N.n1720 0.0254881
R16425 OUT_N.n1741 OUT_N.n1740 0.0254881
R16426 OUT_N.n1931 OUT_N.n1930 0.0235313
R16427 OUT_N.n1198 OUT_N.n1197 0.0235313
R16428 OUT_N.n1563 OUT_N.n1562 0.0235313
R16429 OUT_N.n805 OUT_N.n804 0.0235313
R16430 OUT_N.n998 OUT_N.n997 0.0235313
R16431 OUT_N.n1490 OUT_N.n1489 0.0235313
R16432 OUT_N.n349 OUT_N.n348 0.0235313
R16433 OUT_N.n1 OUT_N.n0 0.0235313
R16434 OUT_N.n405 OUT_N.n404 0.0228651
R16435 OUT_N.n2047 OUT_N.n2045 0.0228651
R16436 OUT_N.n2007 OUT_N.n2006 0.0228651
R16437 OUT_N.n2002 OUT_N.n2001 0.0228651
R16438 OUT_N.n2170 OUT_N.n2130 0.0228651
R16439 OUT_N.n2199 OUT_N.n2198 0.0228651
R16440 OUT_N.n2130 OUT_N.n2129 0.0228651
R16441 OUT_N.n2094 OUT_N.n2093 0.0228651
R16442 OUT_N.n1250 OUT_N.n1249 0.0228651
R16443 OUT_N.n1249 OUT_N.n1248 0.0228651
R16444 OUT_N.n1553 OUT_N.n1552 0.0228651
R16445 OUT_N.n1202 OUT_N.n1201 0.0228651
R16446 OUT_N.n1570 OUT_N.n1569 0.0228651
R16447 OUT_N.n1576 OUT_N.n1575 0.0228651
R16448 OUT_N.n1349 OUT_N.n1347 0.0228651
R16449 OUT_N.n1631 OUT_N.n1630 0.0228651
R16450 OUT_N.n1477 OUT_N.n1476 0.0228651
R16451 OUT_N.n1483 OUT_N.n1482 0.0228651
R16452 OUT_N.n1566 OUT_N.n1565 0.0228651
R16453 OUT_N.n895 OUT_N.n894 0.0228651
R16454 OUT_N.n996 OUT_N.n995 0.0228651
R16455 OUT_N.n1255 OUT_N.n1254 0.0228651
R16456 OUT_N.n900 OUT_N.n899 0.0228651
R16457 OUT_N.n893 OUT_N.n892 0.0228651
R16458 OUT_N.n851 OUT_N.n850 0.0228651
R16459 OUT_N.n1567 OUT_N.n1566 0.0228651
R16460 OUT_N.n1141 OUT_N.n1140 0.0228651
R16461 OUT_N.n1548 OUT_N.n1547 0.0228651
R16462 OUT_N.n809 OUT_N.n808 0.0228651
R16463 OUT_N.n1492 OUT_N.n1491 0.0228651
R16464 OUT_N.n1152 OUT_N.n1151 0.0228651
R16465 OUT_N.n1546 OUT_N.n1545 0.0228651
R16466 OUT_N.n352 OUT_N.n351 0.0228651
R16467 OUT_N.n1543 OUT_N.n1542 0.0228651
R16468 OUT_N.n403 OUT_N.n402 0.0228651
R16469 OUT_N.n1731 OUT_N.n1730 0.0228651
R16470 OUT_N.n1813 OUT_N.n1812 0.0228651
R16471 OUT_N.n1761 OUT_N.n1760 0.0228651
R16472 OUT_N.n1815 OUT_N.n1814 0.0228651
R16473 OUT_N.n31 OUT_N.n30 0.0228651
R16474 OUT_N.n2200 OUT_N.n2051 0.0228651
R16475 OUT_N.n2201 OUT_N.n2048 0.0228651
R16476 OUT_N.n1304 OUT_N.n1303 0.0228651
R16477 OUT_N.n945 OUT_N.n944 0.0228651
R16478 OUT_N.n941 OUT_N.n939 0.0228651
R16479 OUT_N.n1681 OUT_N.n1680 0.0228651
R16480 OUT_N.n610 OUT_N.n609 0.0228651
R16481 OUT_N.n615 OUT_N.n614 0.0228651
R16482 OUT_N.n1672 OUT_N.n1304 0.0228651
R16483 OUT_N.n1300 OUT_N.n945 0.0228651
R16484 OUT_N.n180 OUT_N.n179 0.0228651
R16485 OUT_N.n173 OUT_N.n172 0.0228651
R16486 OUT_N.n3 OUT_N.n2 0.0228651
R16487 OUT_N.n99 OUT_N.n98 0.0195244
R16488 OUT_N.n100 OUT_N.n99 0.0195244
R16489 OUT_N.n101 OUT_N.n100 0.0195244
R16490 OUT_N.n148 OUT_N.n147 0.0195244
R16491 OUT_N.n149 OUT_N.n148 0.0195244
R16492 OUT_N.n150 OUT_N.n149 0.0195244
R16493 OUT_N.n69 OUT_N.n68 0.0195244
R16494 OUT_N.n70 OUT_N.n69 0.0195244
R16495 OUT_N.n71 OUT_N.n70 0.0195244
R16496 OUT_N.n1927 OUT_N.n1890 0.0179841
R16497 OUT_N.n1929 OUT_N.n1928 0.0179841
R16498 OUT_N.n1885 OUT_N.n1884 0.0179841
R16499 OUT_N.n1861 OUT_N.n1860 0.0179841
R16500 OUT_N.n2125 OUT_N.n2124 0.0179841
R16501 OUT_N.n2127 OUT_N.n2126 0.0179841
R16502 OUT_N.n2197 OUT_N.n2196 0.0179841
R16503 OUT_N.n2092 OUT_N.n2091 0.0179841
R16504 OUT_N.n456 OUT_N.n455 0.0179841
R16505 OUT_N.n1556 OUT_N.n1555 0.0179841
R16506 OUT_N.n1625 OUT_N.n1624 0.0179841
R16507 OUT_N.n1245 OUT_N.n1244 0.0179841
R16508 OUT_N.n1623 OUT_N.n1622 0.0179841
R16509 OUT_N.n1578 OUT_N.n1574 0.0179841
R16510 OUT_N.n1627 OUT_N.n1621 0.0179841
R16511 OUT_N.n1558 OUT_N.n1541 0.0179841
R16512 OUT_N.n1480 OUT_N.n1479 0.0179841
R16513 OUT_N.n1138 OUT_N.n1137 0.0179841
R16514 OUT_N.n1144 OUT_N.n1143 0.0179841
R16515 OUT_N.n1252 OUT_N.n1251 0.0179841
R16516 OUT_N.n1551 OUT_N.n1550 0.0179841
R16517 OUT_N.n1496 OUT_N.n1495 0.0179841
R16518 OUT_N.n1498 OUT_N.n1493 0.0179841
R16519 OUT_N.n1149 OUT_N.n1148 0.0179841
R16520 OUT_N.n605 OUT_N.n604 0.0179841
R16521 OUT_N.n360 OUT_N.n359 0.0179841
R16522 OUT_N.n409 OUT_N.n408 0.0179841
R16523 OUT_N.n453 OUT_N.n452 0.0179841
R16524 OUT_N.n538 OUT_N.n537 0.0179841
R16525 OUT_N.n1858 OUT_N.n1857 0.0179841
R16526 OUT_N.n569 OUT_N.n568 0.0179841
R16527 OUT_N.n1856 OUT_N.n1855 0.0179841
R16528 OUT_N.n462 OUT_N.n461 0.0179841
R16529 OUT_N.n354 OUT_N.n350 0.0179841
R16530 OUT_N.n357 OUT_N.n356 0.0179841
R16531 OUT_N.n363 OUT_N.n362 0.0179841
R16532 OUT_N.n407 OUT_N.n406 0.0179841
R16533 OUT_N.n412 OUT_N.n411 0.0179841
R16534 OUT_N.n451 OUT_N.n450 0.0179841
R16535 OUT_N.n459 OUT_N.n458 0.0179841
R16536 OUT_N.n465 OUT_N.n464 0.0179841
R16537 OUT_N.n1758 OUT_N.n1735 0.0179841
R16538 OUT_N.n1811 OUT_N.n1810 0.0179841
R16539 OUT_N.n30 OUT_N.n29 0.0179841
R16540 OUT_N.n606 OUT_N.n605 0.0179841
R16541 OUT_N.n1728 OUT_N.n1727 0.0179841
R16542 OUT_N.n2236 OUT_N.n2233 0.0179841
R16543 OUT_N.n2044 OUT_N.n2040 0.0179841
R16544 OUT_N.n2042 OUT_N.n2041 0.0179841
R16545 OUT_N.n611 OUT_N.n181 0.0179841
R16546 OUT_N.n1679 OUT_N.n1678 0.0179841
R16547 OUT_N.n171 OUT_N.n34 0.0179841
R16548 OUT_N.n1684 OUT_N.n1683 0.0179841
R16549 OUT_N.n2240 OUT_N.n5 0.0179841
R16550 OUT_N.n2043 OUT_N.n2042 0.0177304
R16551 OUT_N.n1857 OUT_N.n1856 0.0177304
R16552 OUT_N.n1999 OUT_N.n1998 0.0177304
R16553 OUT_N.n1928 OUT_N.n1888 0.0177304
R16554 OUT_N.n1890 OUT_N.n1889 0.0177304
R16555 OUT_N.n1853 OUT_N.n1852 0.0177304
R16556 OUT_N.n1884 OUT_N.n1861 0.0177304
R16557 OUT_N.n1860 OUT_N.n1859 0.0177304
R16558 OUT_N.n2091 OUT_N.n2090 0.0177304
R16559 OUT_N.n2196 OUT_N.n2195 0.0177304
R16560 OUT_N.n2126 OUT_N.n2125 0.0177304
R16561 OUT_N.n2124 OUT_N.n2123 0.0177304
R16562 OUT_N.n1555 OUT_N.n1554 0.0177304
R16563 OUT_N.n1244 OUT_N.n1243 0.0177304
R16564 OUT_N.n1624 OUT_N.n1623 0.0177304
R16565 OUT_N.n1578 OUT_N.n1577 0.0177304
R16566 OUT_N.n1558 OUT_N.n1557 0.0177304
R16567 OUT_N.n1627 OUT_N.n1626 0.0177304
R16568 OUT_N.n1619 OUT_N.n1618 0.0177304
R16569 OUT_N.n1539 OUT_N.n1538 0.0177304
R16570 OUT_N.n354 OUT_N.n353 0.0177304
R16571 OUT_N.n1139 OUT_N.n1138 0.0177304
R16572 OUT_N.n1479 OUT_N.n1478 0.0177304
R16573 OUT_N.n1146 OUT_N.n1145 0.0177304
R16574 OUT_N.n1143 OUT_N.n1142 0.0177304
R16575 OUT_N.n1550 OUT_N.n1549 0.0177304
R16576 OUT_N.n1253 OUT_N.n1252 0.0177304
R16577 OUT_N.n1150 OUT_N.n1149 0.0177304
R16578 OUT_N.n1498 OUT_N.n1497 0.0177304
R16579 OUT_N.n1495 OUT_N.n1494 0.0177304
R16580 OUT_N.n1157 OUT_N.n1156 0.0177304
R16581 OUT_N.n536 OUT_N.n535 0.0177304
R16582 OUT_N.n568 OUT_N.n567 0.0177304
R16583 OUT_N.n358 OUT_N.n357 0.0177304
R16584 OUT_N.n410 OUT_N.n407 0.0177304
R16585 OUT_N.n454 OUT_N.n451 0.0177304
R16586 OUT_N.n460 OUT_N.n459 0.0177304
R16587 OUT_N.n2235 OUT_N.n2234 0.0177304
R16588 OUT_N.n1758 OUT_N.n1757 0.0177304
R16589 OUT_N.n1810 OUT_N.n1809 0.0177304
R16590 OUT_N.n29 OUT_N.n28 0.0177304
R16591 OUT_N.n604 OUT_N.n603 0.0177304
R16592 OUT_N.n607 OUT_N.n606 0.0177304
R16593 OUT_N.n1729 OUT_N.n1728 0.0177304
R16594 OUT_N.n2233 OUT_N.n2232 0.0177304
R16595 OUT_N.n1820 OUT_N.n1819 0.0177304
R16596 OUT_N.n2040 OUT_N.n2039 0.0177304
R16597 OUT_N.n1678 OUT_N.n1677 0.0177304
R16598 OUT_N.n612 OUT_N.n611 0.0177304
R16599 OUT_N.n171 OUT_N.n170 0.0177304
R16600 OUT_N.n1683 OUT_N.n1682 0.0177304
R16601 OUT_N.n5 OUT_N.n4 0.0177304
R16602 OUT_N.n1260 OUT_N.n1259 0.0174187
R16603 OUT_N.n1259 OUT_N.n1258 0.0174187
R16604 OUT_N.n1351 OUT_N.n1350 0.0174187
R16605 OUT_N.n850 OUT_N.n849 0.0174187
R16606 OUT_N.n899 OUT_N.n898 0.0174187
R16607 OUT_N.n898 OUT_N.n897 0.0174187
R16608 OUT_N.n849 OUT_N.n848 0.0174187
R16609 OUT_N.n610 OUT_N.n504 0.0174187
R16610 OUT_N.n616 OUT_N.n615 0.0174187
R16611 OUT_N.n942 OUT_N.n616 0.0174187
R16612 OUT_N.n504 OUT_N.n503 0.0174187
R16613 OUT_N.n1975 OUT_N.n1972 0.0173591
R16614 OUT_N.n2194 OUT_N.n2172 0.0173591
R16615 OUT_N.n2004 OUT_N.n2000 0.0173591
R16616 OUT_N.n1971 OUT_N.n1932 0.0173591
R16617 OUT_N.n1887 OUT_N.n1886 0.0173591
R16618 OUT_N.n2005 OUT_N.n2004 0.0173591
R16619 OUT_N.n1976 OUT_N.n1971 0.0173591
R16620 OUT_N.n1975 OUT_N.n1974 0.0173591
R16621 OUT_N.n1888 OUT_N.n1887 0.0173591
R16622 OUT_N.n2121 OUT_N.n2119 0.0173591
R16623 OUT_N.n1854 OUT_N.n1851 0.0173591
R16624 OUT_N.n1854 OUT_N.n1853 0.0173591
R16625 OUT_N.n2122 OUT_N.n2118 0.0173591
R16626 OUT_N.n2118 OUT_N.n2095 0.0173591
R16627 OUT_N.n2121 OUT_N.n2120 0.0173591
R16628 OUT_N.n2194 OUT_N.n2193 0.0173591
R16629 OUT_N.n1196 OUT_N.n1195 0.0173591
R16630 OUT_N.n1203 OUT_N.n1202 0.0173591
R16631 OUT_N.n1242 OUT_N.n1241 0.0173591
R16632 OUT_N.n1258 OUT_N.n1257 0.0173591
R16633 OUT_N.n1197 OUT_N.n1196 0.0173591
R16634 OUT_N.n1257 OUT_N.n1246 0.0173591
R16635 OUT_N.n1243 OUT_N.n1242 0.0173591
R16636 OUT_N.n1573 OUT_N.n1572 0.0173591
R16637 OUT_N.n1572 OUT_N.n1571 0.0173591
R16638 OUT_N.n1204 OUT_N.n1203 0.0173591
R16639 OUT_N.n1476 OUT_N.n1475 0.0173591
R16640 OUT_N.n1489 OUT_N.n1488 0.0173591
R16641 OUT_N.n1540 OUT_N.n1537 0.0173591
R16642 OUT_N.n1562 OUT_N.n1561 0.0173591
R16643 OUT_N.n1620 OUT_N.n1617 0.0173591
R16644 OUT_N.n1561 OUT_N.n1560 0.0173591
R16645 OUT_N.n1537 OUT_N.n1536 0.0173591
R16646 OUT_N.n1617 OUT_N.n1616 0.0173591
R16647 OUT_N.n1485 OUT_N.n1481 0.0173591
R16648 OUT_N.n1485 OUT_N.n1484 0.0173591
R16649 OUT_N.n1475 OUT_N.n1474 0.0173591
R16650 OUT_N.n803 OUT_N.n802 0.0173591
R16651 OUT_N.n810 OUT_N.n809 0.0173591
R16652 OUT_N.n804 OUT_N.n803 0.0173591
R16653 OUT_N.n1155 OUT_N.n1154 0.0173591
R16654 OUT_N.n1154 OUT_N.n1153 0.0173591
R16655 OUT_N.n1488 OUT_N.n1487 0.0173591
R16656 OUT_N.n811 OUT_N.n810 0.0173591
R16657 OUT_N.n348 OUT_N.n347 0.0173591
R16658 OUT_N.n364 OUT_N.n361 0.0173591
R16659 OUT_N.n463 OUT_N.n460 0.0173591
R16660 OUT_N.n573 OUT_N.n572 0.0173591
R16661 OUT_N.n570 OUT_N.n569 0.0173591
R16662 OUT_N.n361 OUT_N.n358 0.0173591
R16663 OUT_N.n574 OUT_N.n573 0.0173591
R16664 OUT_N.n571 OUT_N.n570 0.0173591
R16665 OUT_N.n466 OUT_N.n463 0.0173591
R16666 OUT_N.n347 OUT_N.n346 0.0173591
R16667 OUT_N.n1676 OUT_N.n1674 0.0173591
R16668 OUT_N.n1808 OUT_N.n1806 0.0173591
R16669 OUT_N.n1804 OUT_N.n1765 0.0173591
R16670 OUT_N.n1818 OUT_N.n1817 0.0173591
R16671 OUT_N.n1805 OUT_N.n1764 0.0173591
R16672 OUT_N.n1759 OUT_N.n1734 0.0173591
R16673 OUT_N.n1734 OUT_N.n1732 0.0173591
R16674 OUT_N.n1764 OUT_N.n1762 0.0173591
R16675 OUT_N.n1804 OUT_N.n1803 0.0173591
R16676 OUT_N.n1808 OUT_N.n1807 0.0173591
R16677 OUT_N.n1817 OUT_N.n1816 0.0173591
R16678 OUT_N.n2238 OUT_N.n1687 0.0173591
R16679 OUT_N.n2231 OUT_N.n2230 0.0173591
R16680 OUT_N.n2039 OUT_N.n2038 0.0173591
R16681 OUT_N.n2232 OUT_N.n2231 0.0173591
R16682 OUT_N.n2038 OUT_N.n2037 0.0173591
R16683 OUT_N.n2239 OUT_N.n1686 0.0173591
R16684 OUT_N.n177 OUT_N.n174 0.0173591
R16685 OUT_N.n1686 OUT_N.n1684 0.0173591
R16686 OUT_N.n2238 OUT_N.n2237 0.0173591
R16687 OUT_N.n1676 OUT_N.n1675 0.0173591
R16688 OUT_N.n178 OUT_N.n177 0.0173591
R16689 OUT_N.n2241 OUT_N.n1 0.0173591
R16690 OUT_N.n2242 OUT_N.n2241 0.0173591
R16691 OUT_N.n1935 OUT_N.n1934 0.0167343
R16692 OUT_N.n2139 OUT_N.n2138 0.0167343
R16693 OUT_N.n1690 OUT_N.n1689 0.0167343
R16694 OUT_N.n1932 OUT_N.n1931 0.0122638
R16695 OUT_N.n2053 OUT_N.n2052 0.0122638
R16696 OUT_N.n1199 OUT_N.n1198 0.0122638
R16697 OUT_N.n1579 OUT_N.n1563 0.0122638
R16698 OUT_N.n806 OUT_N.n805 0.0122638
R16699 OUT_N.n997 OUT_N.n996 0.0122638
R16700 OUT_N.n1499 OUT_N.n1490 0.0122638
R16701 OUT_N.n355 OUT_N.n349 0.0122638
R16702 OUT_N.n33 OUT_N.n6 0.0122638
R16703 OUT_N.n1725 OUT_N.n1688 0.0122638
R16704 OUT_N.n404 OUT_N.n403 0.0119325
R16705 OUT_N.n2048 OUT_N.n2047 0.0119325
R16706 OUT_N.n176 OUT_N.n175 0.0119325
R16707 OUT_N.n1970 OUT_N.n1933 0.0119325
R16708 OUT_N.n2003 OUT_N.n2002 0.0119325
R16709 OUT_N.n2006 OUT_N.n2005 0.0119325
R16710 OUT_N.n2117 OUT_N.n2116 0.0119325
R16711 OUT_N.n2050 OUT_N.n2049 0.0119325
R16712 OUT_N.n2051 OUT_N.n2050 0.0119325
R16713 OUT_N.n2198 OUT_N.n2197 0.0119325
R16714 OUT_N.n2171 OUT_N.n2170 0.0119325
R16715 OUT_N.n2129 OUT_N.n2128 0.0119325
R16716 OUT_N.n2095 OUT_N.n2094 0.0119325
R16717 OUT_N.n995 OUT_N.n994 0.0119325
R16718 OUT_N.n1349 OUT_N.n1348 0.0119325
R16719 OUT_N.n1248 OUT_N.n1247 0.0119325
R16720 OUT_N.n1256 OUT_N.n1250 0.0119325
R16721 OUT_N.n1254 OUT_N.n1253 0.0119325
R16722 OUT_N.n1554 OUT_N.n1553 0.0119325
R16723 OUT_N.n1549 OUT_N.n1548 0.0119325
R16724 OUT_N.n1545 OUT_N.n1544 0.0119325
R16725 OUT_N.n1544 OUT_N.n1543 0.0119325
R16726 OUT_N.n1201 OUT_N.n1200 0.0119325
R16727 OUT_N.n1577 OUT_N.n1576 0.0119325
R16728 OUT_N.n1571 OUT_N.n1570 0.0119325
R16729 OUT_N.n1568 OUT_N.n1567 0.0119325
R16730 OUT_N.n1565 OUT_N.n1564 0.0119325
R16731 OUT_N.n1486 OUT_N.n1477 0.0119325
R16732 OUT_N.n1630 OUT_N.n1629 0.0119325
R16733 OUT_N.n1484 OUT_N.n1483 0.0119325
R16734 OUT_N.n1142 OUT_N.n1141 0.0119325
R16735 OUT_N.n353 OUT_N.n352 0.0119325
R16736 OUT_N.n808 OUT_N.n807 0.0119325
R16737 OUT_N.n852 OUT_N.n851 0.0119325
R16738 OUT_N.n894 OUT_N.n893 0.0119325
R16739 OUT_N.n896 OUT_N.n895 0.0119325
R16740 OUT_N.n901 OUT_N.n900 0.0119325
R16741 OUT_N.n941 OUT_N.n940 0.0119325
R16742 OUT_N.n1493 OUT_N.n1492 0.0119325
R16743 OUT_N.n1153 OUT_N.n1152 0.0119325
R16744 OUT_N.n402 OUT_N.n401 0.0119325
R16745 OUT_N.n609 OUT_N.n608 0.0119325
R16746 OUT_N.n32 OUT_N.n31 0.0119325
R16747 OUT_N.n1816 OUT_N.n1815 0.0119325
R16748 OUT_N.n1812 OUT_N.n1811 0.0119325
R16749 OUT_N.n1762 OUT_N.n1761 0.0119325
R16750 OUT_N.n1732 OUT_N.n1731 0.0119325
R16751 OUT_N.n2202 OUT_N.n2201 0.0119325
R16752 OUT_N.n1680 OUT_N.n1679 0.0119325
R16753 OUT_N.n1673 OUT_N.n1672 0.0119325
R16754 OUT_N.n1303 OUT_N.n1302 0.0119325
R16755 OUT_N.n1301 OUT_N.n1300 0.0119325
R16756 OUT_N.n944 OUT_N.n943 0.0119325
R16757 OUT_N.n614 OUT_N.n613 0.0119325
R16758 OUT_N.n181 OUT_N.n180 0.0119325
R16759 OUT_N.n174 OUT_N.n173 0.0119325
R16760 OUT_N.n4 OUT_N.n3 0.0119325
R16761 OUT_N.n2079 OUT_N.n2078 0.00905634
R16762 OUT_N.n2088 OUT_N.n2087 0.00905634
R16763 OUT_N.n1923 OUT_N.n1922 0.00905634
R16764 OUT_N.n1916 OUT_N.n1915 0.00905634
R16765 OUT_N.n1969 OUT_N.n1968 0.00905634
R16766 OUT_N.n1950 OUT_N.n1949 0.00905634
R16767 OUT_N.n2181 OUT_N.n2180 0.00905634
R16768 OUT_N.n2115 OUT_N.n2114 0.00905634
R16769 OUT_N.n1875 OUT_N.n1874 0.00905634
R16770 OUT_N.n1127 OUT_N.n1126 0.00905634
R16771 OUT_N.n1136 OUT_N.n1135 0.00905634
R16772 OUT_N.n1167 OUT_N.n1166 0.00905634
R16773 OUT_N.n1176 OUT_N.n1175 0.00905634
R16774 OUT_N.n1185 OUT_N.n1184 0.00905634
R16775 OUT_N.n1194 OUT_N.n1193 0.00905634
R16776 OUT_N.n1213 OUT_N.n1212 0.00905634
R16777 OUT_N.n1222 OUT_N.n1221 0.00905634
R16778 OUT_N.n1231 OUT_N.n1230 0.00905634
R16779 OUT_N.n1240 OUT_N.n1239 0.00905634
R16780 OUT_N.n1269 OUT_N.n1268 0.00905634
R16781 OUT_N.n1278 OUT_N.n1277 0.00905634
R16782 OUT_N.n1287 OUT_N.n1286 0.00905634
R16783 OUT_N.n1296 OUT_N.n1295 0.00905634
R16784 OUT_N.n1464 OUT_N.n1463 0.00905634
R16785 OUT_N.n1473 OUT_N.n1472 0.00905634
R16786 OUT_N.n1508 OUT_N.n1507 0.00905634
R16787 OUT_N.n1517 OUT_N.n1516 0.00905634
R16788 OUT_N.n1526 OUT_N.n1525 0.00905634
R16789 OUT_N.n1535 OUT_N.n1534 0.00905634
R16790 OUT_N.n1588 OUT_N.n1587 0.00905634
R16791 OUT_N.n1597 OUT_N.n1596 0.00905634
R16792 OUT_N.n1606 OUT_N.n1605 0.00905634
R16793 OUT_N.n1615 OUT_N.n1614 0.00905634
R16794 OUT_N.n1641 OUT_N.n1640 0.00905634
R16795 OUT_N.n1650 OUT_N.n1649 0.00905634
R16796 OUT_N.n1659 OUT_N.n1658 0.00905634
R16797 OUT_N.n1668 OUT_N.n1667 0.00905634
R16798 OUT_N.n792 OUT_N.n791 0.00905634
R16799 OUT_N.n801 OUT_N.n800 0.00905634
R16800 OUT_N.n820 OUT_N.n819 0.00905634
R16801 OUT_N.n829 OUT_N.n828 0.00905634
R16802 OUT_N.n838 OUT_N.n837 0.00905634
R16803 OUT_N.n847 OUT_N.n846 0.00905634
R16804 OUT_N.n864 OUT_N.n863 0.00905634
R16805 OUT_N.n873 OUT_N.n872 0.00905634
R16806 OUT_N.n882 OUT_N.n881 0.00905634
R16807 OUT_N.n891 OUT_N.n890 0.00905634
R16808 OUT_N.n910 OUT_N.n909 0.00905634
R16809 OUT_N.n919 OUT_N.n918 0.00905634
R16810 OUT_N.n928 OUT_N.n927 0.00905634
R16811 OUT_N.n937 OUT_N.n936 0.00905634
R16812 OUT_N.n336 OUT_N.n335 0.00905634
R16813 OUT_N.n345 OUT_N.n344 0.00905634
R16814 OUT_N.n373 OUT_N.n372 0.00905634
R16815 OUT_N.n382 OUT_N.n381 0.00905634
R16816 OUT_N.n391 OUT_N.n390 0.00905634
R16817 OUT_N.n400 OUT_N.n399 0.00905634
R16818 OUT_N.n422 OUT_N.n421 0.00905634
R16819 OUT_N.n431 OUT_N.n430 0.00905634
R16820 OUT_N.n440 OUT_N.n439 0.00905634
R16821 OUT_N.n449 OUT_N.n448 0.00905634
R16822 OUT_N.n475 OUT_N.n474 0.00905634
R16823 OUT_N.n484 OUT_N.n483 0.00905634
R16824 OUT_N.n493 OUT_N.n492 0.00905634
R16825 OUT_N.n502 OUT_N.n501 0.00905634
R16826 OUT_N.n600 OUT_N.n599 0.00905634
R16827 OUT_N.n591 OUT_N.n590 0.00905634
R16828 OUT_N.n582 OUT_N.n581 0.00905634
R16829 OUT_N.n564 OUT_N.n563 0.00905634
R16830 OUT_N.n555 OUT_N.n554 0.00905634
R16831 OUT_N.n1702 OUT_N.n1701 0.00905634
R16832 OUT_N.n2222 OUT_N.n2221 0.00905634
R16833 OUT_N.n2213 OUT_N.n2212 0.00905634
R16834 OUT_N.n2204 OUT_N.n2203 0.00905634
R16835 OUT_N.n2029 OUT_N.n2028 0.00905634
R16836 OUT_N.n1711 OUT_N.n1710 0.00740328
R16837 OUT_N.n2157 OUT_N.n2156 0.00735609
R16838 OUT_N.n1992 OUT_N.n1991 0.00735609
R16839 OUT_N.n1997 OUT_N.n1996 0.00735609
R16840 OUT_N.n2183 OUT_N.n2182 0.00735609
R16841 OUT_N.n22 OUT_N.n21 0.00735609
R16842 OUT_N.n27 OUT_N.n26 0.00735609
R16843 OUT_N.n1724 OUT_N.n1723 0.00735609
R16844 OUT_N.n1792 OUT_N.n1791 0.00735609
R16845 OUT_N.n1751 OUT_N.n1750 0.00735609
R16846 OUT_N.n1756 OUT_N.n1755 0.00735609
R16847 OUT_N.n73 OUT_N.n72 0.00556853
R16848 OUT_N.n87 OUT_N.n86 0.00556853
R16849 OUT_N.n81 OUT_N.n80 0.00556853
R16850 OUT_N.n158 OUT_N.n157 0.00556853
R16851 OUT_N.n163 OUT_N.n162 0.00556853
R16852 OUT_N.n134 OUT_N.n133 0.00556853
R16853 OUT_N.n141 OUT_N.n140 0.00556853
R16854 OUT_N.n112 OUT_N.n111 0.00556853
R16855 OUT_N.n118 OUT_N.n117 0.00556853
R16856 OUT_N.n124 OUT_N.n123 0.00556853
R16857 OUT_N.n131 OUT_N.n130 0.00556853
R16858 OUT_N.n130 OUT_N.n129 0.00556853
R16859 OUT_N.n157 OUT_N.n156 0.00556853
R16860 OUT_N.n117 OUT_N.n116 0.00556853
R16861 OUT_N.n142 OUT_N.n141 0.00556853
R16862 OUT_N.n123 OUT_N.n122 0.00556853
R16863 OUT_N.n164 OUT_N.n163 0.00556853
R16864 OUT_N.n133 OUT_N.n132 0.00556853
R16865 OUT_N.n111 OUT_N.n110 0.00556853
R16866 OUT_N.n41 OUT_N.n40 0.00556853
R16867 OUT_N.n46 OUT_N.n45 0.00556853
R16868 OUT_N.n53 OUT_N.n52 0.00556853
R16869 OUT_N.n59 OUT_N.n58 0.00556853
R16870 OUT_N.n58 OUT_N.n57 0.00556853
R16871 OUT_N.n47 OUT_N.n46 0.00556853
R16872 OUT_N.n52 OUT_N.n51 0.00556853
R16873 OUT_N.n40 OUT_N.n39 0.00556853
R16874 OUT_N.n82 OUT_N.n81 0.00556853
R16875 OUT_N.n96 OUT_N.n95 0.00556853
R16876 OUT_N.n88 OUT_N.n87 0.00556853
R16877 OUT_N.n331 OUT_N.n330 0.00528925
R16878 OUT_N.n335 OUT_N.n334 0.00528925
R16879 OUT_N.n340 OUT_N.n339 0.00528925
R16880 OUT_N.n556 OUT_N.n555 0.00528925
R16881 OUT_N.n560 OUT_N.n559 0.00528925
R16882 OUT_N.n565 OUT_N.n564 0.00528925
R16883 OUT_N.n2110 OUT_N.n2109 0.00528925
R16884 OUT_N.n1876 OUT_N.n1875 0.00528925
R16885 OUT_N.n1880 OUT_N.n1879 0.00528925
R16886 OUT_N.n2114 OUT_N.n2113 0.00528925
R16887 OUT_N.n1951 OUT_N.n1950 0.00528925
R16888 OUT_N.n1924 OUT_N.n1923 0.00528925
R16889 OUT_N.n1956 OUT_N.n1955 0.00528925
R16890 OUT_N.n2078 OUT_N.n2069 0.00528925
R16891 OUT_N.n2160 OUT_N.n2159 0.00528925
R16892 OUT_N.n2083 OUT_N.n2082 0.00528925
R16893 OUT_N.n2165 OUT_N.n2164 0.00528925
R16894 OUT_N.n2087 OUT_N.n2086 0.00528925
R16895 OUT_N.n1920 OUT_N.n1919 0.00528925
R16896 OUT_N.n578 OUT_N.n577 0.00528925
R16897 OUT_N.n583 OUT_N.n582 0.00528925
R16898 OUT_N.n587 OUT_N.n586 0.00528925
R16899 OUT_N.n592 OUT_N.n591 0.00528925
R16900 OUT_N.n596 OUT_N.n595 0.00528925
R16901 OUT_N.n601 OUT_N.n600 0.00528925
R16902 OUT_N.n787 OUT_N.n786 0.00528925
R16903 OUT_N.n791 OUT_N.n790 0.00528925
R16904 OUT_N.n796 OUT_N.n795 0.00528925
R16905 OUT_N.n800 OUT_N.n799 0.00528925
R16906 OUT_N.n815 OUT_N.n814 0.00528925
R16907 OUT_N.n819 OUT_N.n818 0.00528925
R16908 OUT_N.n824 OUT_N.n823 0.00528925
R16909 OUT_N.n828 OUT_N.n827 0.00528925
R16910 OUT_N.n833 OUT_N.n832 0.00528925
R16911 OUT_N.n837 OUT_N.n836 0.00528925
R16912 OUT_N.n842 OUT_N.n841 0.00528925
R16913 OUT_N.n936 OUT_N.n935 0.00528925
R16914 OUT_N.n932 OUT_N.n931 0.00528925
R16915 OUT_N.n927 OUT_N.n926 0.00528925
R16916 OUT_N.n923 OUT_N.n922 0.00528925
R16917 OUT_N.n918 OUT_N.n917 0.00528925
R16918 OUT_N.n914 OUT_N.n913 0.00528925
R16919 OUT_N.n909 OUT_N.n908 0.00528925
R16920 OUT_N.n905 OUT_N.n904 0.00528925
R16921 OUT_N.n890 OUT_N.n889 0.00528925
R16922 OUT_N.n886 OUT_N.n885 0.00528925
R16923 OUT_N.n881 OUT_N.n880 0.00528925
R16924 OUT_N.n877 OUT_N.n876 0.00528925
R16925 OUT_N.n872 OUT_N.n871 0.00528925
R16926 OUT_N.n868 OUT_N.n867 0.00528925
R16927 OUT_N.n863 OUT_N.n862 0.00528925
R16928 OUT_N.n859 OUT_N.n858 0.00528925
R16929 OUT_N.n846 OUT_N.n845 0.00528925
R16930 OUT_N.n1459 OUT_N.n1458 0.00528925
R16931 OUT_N.n1463 OUT_N.n1462 0.00528925
R16932 OUT_N.n1468 OUT_N.n1467 0.00528925
R16933 OUT_N.n1472 OUT_N.n1471 0.00528925
R16934 OUT_N.n1503 OUT_N.n1502 0.00528925
R16935 OUT_N.n1507 OUT_N.n1506 0.00528925
R16936 OUT_N.n1512 OUT_N.n1511 0.00528925
R16937 OUT_N.n1516 OUT_N.n1515 0.00528925
R16938 OUT_N.n1521 OUT_N.n1520 0.00528925
R16939 OUT_N.n1525 OUT_N.n1524 0.00528925
R16940 OUT_N.n1530 OUT_N.n1529 0.00528925
R16941 OUT_N.n1534 OUT_N.n1533 0.00528925
R16942 OUT_N.n1583 OUT_N.n1582 0.00528925
R16943 OUT_N.n1587 OUT_N.n1586 0.00528925
R16944 OUT_N.n1592 OUT_N.n1591 0.00528925
R16945 OUT_N.n1596 OUT_N.n1595 0.00528925
R16946 OUT_N.n1601 OUT_N.n1600 0.00528925
R16947 OUT_N.n1605 OUT_N.n1604 0.00528925
R16948 OUT_N.n1610 OUT_N.n1609 0.00528925
R16949 OUT_N.n1667 OUT_N.n1666 0.00528925
R16950 OUT_N.n1663 OUT_N.n1662 0.00528925
R16951 OUT_N.n1658 OUT_N.n1657 0.00528925
R16952 OUT_N.n1654 OUT_N.n1653 0.00528925
R16953 OUT_N.n1649 OUT_N.n1648 0.00528925
R16954 OUT_N.n1645 OUT_N.n1644 0.00528925
R16955 OUT_N.n1640 OUT_N.n1639 0.00528925
R16956 OUT_N.n1636 OUT_N.n1635 0.00528925
R16957 OUT_N.n1614 OUT_N.n1613 0.00528925
R16958 OUT_N.n1122 OUT_N.n1121 0.00528925
R16959 OUT_N.n1126 OUT_N.n1125 0.00528925
R16960 OUT_N.n1131 OUT_N.n1130 0.00528925
R16961 OUT_N.n1135 OUT_N.n1134 0.00528925
R16962 OUT_N.n1162 OUT_N.n1161 0.00528925
R16963 OUT_N.n1166 OUT_N.n1165 0.00528925
R16964 OUT_N.n1171 OUT_N.n1170 0.00528925
R16965 OUT_N.n1175 OUT_N.n1174 0.00528925
R16966 OUT_N.n1180 OUT_N.n1179 0.00528925
R16967 OUT_N.n1184 OUT_N.n1183 0.00528925
R16968 OUT_N.n1189 OUT_N.n1188 0.00528925
R16969 OUT_N.n1193 OUT_N.n1192 0.00528925
R16970 OUT_N.n1208 OUT_N.n1207 0.00528925
R16971 OUT_N.n1212 OUT_N.n1211 0.00528925
R16972 OUT_N.n1217 OUT_N.n1216 0.00528925
R16973 OUT_N.n1221 OUT_N.n1220 0.00528925
R16974 OUT_N.n1226 OUT_N.n1225 0.00528925
R16975 OUT_N.n1230 OUT_N.n1229 0.00528925
R16976 OUT_N.n1235 OUT_N.n1234 0.00528925
R16977 OUT_N.n1295 OUT_N.n1294 0.00528925
R16978 OUT_N.n1291 OUT_N.n1290 0.00528925
R16979 OUT_N.n1286 OUT_N.n1285 0.00528925
R16980 OUT_N.n1282 OUT_N.n1281 0.00528925
R16981 OUT_N.n1277 OUT_N.n1276 0.00528925
R16982 OUT_N.n1273 OUT_N.n1272 0.00528925
R16983 OUT_N.n1268 OUT_N.n1267 0.00528925
R16984 OUT_N.n1264 OUT_N.n1263 0.00528925
R16985 OUT_N.n1239 OUT_N.n1238 0.00528925
R16986 OUT_N.n344 OUT_N.n343 0.00528925
R16987 OUT_N.n368 OUT_N.n367 0.00528925
R16988 OUT_N.n372 OUT_N.n371 0.00528925
R16989 OUT_N.n377 OUT_N.n376 0.00528925
R16990 OUT_N.n381 OUT_N.n380 0.00528925
R16991 OUT_N.n386 OUT_N.n385 0.00528925
R16992 OUT_N.n390 OUT_N.n389 0.00528925
R16993 OUT_N.n395 OUT_N.n394 0.00528925
R16994 OUT_N.n399 OUT_N.n398 0.00528925
R16995 OUT_N.n417 OUT_N.n416 0.00528925
R16996 OUT_N.n421 OUT_N.n420 0.00528925
R16997 OUT_N.n426 OUT_N.n425 0.00528925
R16998 OUT_N.n430 OUT_N.n429 0.00528925
R16999 OUT_N.n435 OUT_N.n434 0.00528925
R17000 OUT_N.n439 OUT_N.n438 0.00528925
R17001 OUT_N.n444 OUT_N.n443 0.00528925
R17002 OUT_N.n448 OUT_N.n447 0.00528925
R17003 OUT_N.n470 OUT_N.n469 0.00528925
R17004 OUT_N.n474 OUT_N.n473 0.00528925
R17005 OUT_N.n479 OUT_N.n478 0.00528925
R17006 OUT_N.n483 OUT_N.n482 0.00528925
R17007 OUT_N.n488 OUT_N.n487 0.00528925
R17008 OUT_N.n492 OUT_N.n491 0.00528925
R17009 OUT_N.n497 OUT_N.n496 0.00528925
R17010 OUT_N.n501 OUT_N.n500 0.00528925
R17011 OUT_N.n1796 OUT_N.n1795 0.00528925
R17012 OUT_N.n1705 OUT_N.n1704 0.00528925
R17013 OUT_N.n1801 OUT_N.n1800 0.00528925
R17014 OUT_N.n2227 OUT_N.n2226 0.00528925
R17015 OUT_N.n2223 OUT_N.n2222 0.00528925
R17016 OUT_N.n2218 OUT_N.n2217 0.00528925
R17017 OUT_N.n2214 OUT_N.n2213 0.00528925
R17018 OUT_N.n2209 OUT_N.n2208 0.00528925
R17019 OUT_N.n2205 OUT_N.n2204 0.00528925
R17020 OUT_N.n2034 OUT_N.n2033 0.00528925
R17021 OUT_N.n2030 OUT_N.n2029 0.00528925
R17022 OUT_N.n2026 OUT_N.n2025 0.00528925
R17023 OUT_N.n2081 OUT_N.n2080 0.00527411
R17024 OUT_N.n1918 OUT_N.n1917 0.00527411
R17025 OUT_N.n2082 OUT_N.n2081 0.00527411
R17026 OUT_N.n1919 OUT_N.n1918 0.00527411
R17027 OUT_N.n2162 OUT_N.n2161 0.00527411
R17028 OUT_N.n2167 OUT_N.n2166 0.00527411
R17029 OUT_N.n1959 OUT_N.n1958 0.00527411
R17030 OUT_N.n1954 OUT_N.n1953 0.00527411
R17031 OUT_N.n2161 OUT_N.n2160 0.00527411
R17032 OUT_N.n2166 OUT_N.n2165 0.00527411
R17033 OUT_N.n1955 OUT_N.n1954 0.00527411
R17034 OUT_N.n1968 OUT_N.n1959 0.00527411
R17035 OUT_N.n2192 OUT_N.n2191 0.00527411
R17036 OUT_N.n1994 OUT_N.n1993 0.00527411
R17037 OUT_N.n1995 OUT_N.n1994 0.00527411
R17038 OUT_N.n2191 OUT_N.n2190 0.00527411
R17039 OUT_N.n1882 OUT_N.n1881 0.00527411
R17040 OUT_N.n1881 OUT_N.n1880 0.00527411
R17041 OUT_N.n2109 OUT_N.n2108 0.00527411
R17042 OUT_N.n1129 OUT_N.n1128 0.00527411
R17043 OUT_N.n1160 OUT_N.n1159 0.00527411
R17044 OUT_N.n1169 OUT_N.n1168 0.00527411
R17045 OUT_N.n1178 OUT_N.n1177 0.00527411
R17046 OUT_N.n1187 OUT_N.n1186 0.00527411
R17047 OUT_N.n1206 OUT_N.n1205 0.00527411
R17048 OUT_N.n1215 OUT_N.n1214 0.00527411
R17049 OUT_N.n1224 OUT_N.n1223 0.00527411
R17050 OUT_N.n1233 OUT_N.n1232 0.00527411
R17051 OUT_N.n1262 OUT_N.n1261 0.00527411
R17052 OUT_N.n1271 OUT_N.n1270 0.00527411
R17053 OUT_N.n1280 OUT_N.n1279 0.00527411
R17054 OUT_N.n1289 OUT_N.n1288 0.00527411
R17055 OUT_N.n1263 OUT_N.n1262 0.00527411
R17056 OUT_N.n1272 OUT_N.n1271 0.00527411
R17057 OUT_N.n1281 OUT_N.n1280 0.00527411
R17058 OUT_N.n1290 OUT_N.n1289 0.00527411
R17059 OUT_N.n1234 OUT_N.n1233 0.00527411
R17060 OUT_N.n1225 OUT_N.n1224 0.00527411
R17061 OUT_N.n1216 OUT_N.n1215 0.00527411
R17062 OUT_N.n1207 OUT_N.n1206 0.00527411
R17063 OUT_N.n1188 OUT_N.n1187 0.00527411
R17064 OUT_N.n1179 OUT_N.n1178 0.00527411
R17065 OUT_N.n1170 OUT_N.n1169 0.00527411
R17066 OUT_N.n1161 OUT_N.n1160 0.00527411
R17067 OUT_N.n1130 OUT_N.n1129 0.00527411
R17068 OUT_N.n1121 OUT_N.n1120 0.00527411
R17069 OUT_N.n1466 OUT_N.n1465 0.00527411
R17070 OUT_N.n1501 OUT_N.n1500 0.00527411
R17071 OUT_N.n1510 OUT_N.n1509 0.00527411
R17072 OUT_N.n1519 OUT_N.n1518 0.00527411
R17073 OUT_N.n1528 OUT_N.n1527 0.00527411
R17074 OUT_N.n1581 OUT_N.n1580 0.00527411
R17075 OUT_N.n1590 OUT_N.n1589 0.00527411
R17076 OUT_N.n1599 OUT_N.n1598 0.00527411
R17077 OUT_N.n1608 OUT_N.n1607 0.00527411
R17078 OUT_N.n1634 OUT_N.n1633 0.00527411
R17079 OUT_N.n1643 OUT_N.n1642 0.00527411
R17080 OUT_N.n1652 OUT_N.n1651 0.00527411
R17081 OUT_N.n1661 OUT_N.n1660 0.00527411
R17082 OUT_N.n1635 OUT_N.n1634 0.00527411
R17083 OUT_N.n1644 OUT_N.n1643 0.00527411
R17084 OUT_N.n1653 OUT_N.n1652 0.00527411
R17085 OUT_N.n1662 OUT_N.n1661 0.00527411
R17086 OUT_N.n1609 OUT_N.n1608 0.00527411
R17087 OUT_N.n1600 OUT_N.n1599 0.00527411
R17088 OUT_N.n1591 OUT_N.n1590 0.00527411
R17089 OUT_N.n1582 OUT_N.n1581 0.00527411
R17090 OUT_N.n1529 OUT_N.n1528 0.00527411
R17091 OUT_N.n1520 OUT_N.n1519 0.00527411
R17092 OUT_N.n1511 OUT_N.n1510 0.00527411
R17093 OUT_N.n1502 OUT_N.n1501 0.00527411
R17094 OUT_N.n1467 OUT_N.n1466 0.00527411
R17095 OUT_N.n1458 OUT_N.n1457 0.00527411
R17096 OUT_N.n794 OUT_N.n793 0.00527411
R17097 OUT_N.n813 OUT_N.n812 0.00527411
R17098 OUT_N.n822 OUT_N.n821 0.00527411
R17099 OUT_N.n831 OUT_N.n830 0.00527411
R17100 OUT_N.n840 OUT_N.n839 0.00527411
R17101 OUT_N.n857 OUT_N.n856 0.00527411
R17102 OUT_N.n866 OUT_N.n865 0.00527411
R17103 OUT_N.n875 OUT_N.n874 0.00527411
R17104 OUT_N.n884 OUT_N.n883 0.00527411
R17105 OUT_N.n903 OUT_N.n902 0.00527411
R17106 OUT_N.n912 OUT_N.n911 0.00527411
R17107 OUT_N.n921 OUT_N.n920 0.00527411
R17108 OUT_N.n930 OUT_N.n929 0.00527411
R17109 OUT_N.n858 OUT_N.n857 0.00527411
R17110 OUT_N.n867 OUT_N.n866 0.00527411
R17111 OUT_N.n876 OUT_N.n875 0.00527411
R17112 OUT_N.n885 OUT_N.n884 0.00527411
R17113 OUT_N.n904 OUT_N.n903 0.00527411
R17114 OUT_N.n913 OUT_N.n912 0.00527411
R17115 OUT_N.n922 OUT_N.n921 0.00527411
R17116 OUT_N.n931 OUT_N.n930 0.00527411
R17117 OUT_N.n841 OUT_N.n840 0.00527411
R17118 OUT_N.n832 OUT_N.n831 0.00527411
R17119 OUT_N.n823 OUT_N.n822 0.00527411
R17120 OUT_N.n814 OUT_N.n813 0.00527411
R17121 OUT_N.n795 OUT_N.n794 0.00527411
R17122 OUT_N.n786 OUT_N.n785 0.00527411
R17123 OUT_N.n338 OUT_N.n337 0.00527411
R17124 OUT_N.n366 OUT_N.n365 0.00527411
R17125 OUT_N.n375 OUT_N.n374 0.00527411
R17126 OUT_N.n384 OUT_N.n383 0.00527411
R17127 OUT_N.n393 OUT_N.n392 0.00527411
R17128 OUT_N.n415 OUT_N.n414 0.00527411
R17129 OUT_N.n424 OUT_N.n423 0.00527411
R17130 OUT_N.n433 OUT_N.n432 0.00527411
R17131 OUT_N.n442 OUT_N.n441 0.00527411
R17132 OUT_N.n468 OUT_N.n467 0.00527411
R17133 OUT_N.n477 OUT_N.n476 0.00527411
R17134 OUT_N.n486 OUT_N.n485 0.00527411
R17135 OUT_N.n495 OUT_N.n494 0.00527411
R17136 OUT_N.n598 OUT_N.n597 0.00527411
R17137 OUT_N.n589 OUT_N.n588 0.00527411
R17138 OUT_N.n580 OUT_N.n579 0.00527411
R17139 OUT_N.n562 OUT_N.n561 0.00527411
R17140 OUT_N.n496 OUT_N.n495 0.00527411
R17141 OUT_N.n487 OUT_N.n486 0.00527411
R17142 OUT_N.n478 OUT_N.n477 0.00527411
R17143 OUT_N.n469 OUT_N.n468 0.00527411
R17144 OUT_N.n443 OUT_N.n442 0.00527411
R17145 OUT_N.n434 OUT_N.n433 0.00527411
R17146 OUT_N.n425 OUT_N.n424 0.00527411
R17147 OUT_N.n416 OUT_N.n415 0.00527411
R17148 OUT_N.n394 OUT_N.n393 0.00527411
R17149 OUT_N.n385 OUT_N.n384 0.00527411
R17150 OUT_N.n376 OUT_N.n375 0.00527411
R17151 OUT_N.n367 OUT_N.n366 0.00527411
R17152 OUT_N.n597 OUT_N.n596 0.00527411
R17153 OUT_N.n588 OUT_N.n587 0.00527411
R17154 OUT_N.n579 OUT_N.n578 0.00527411
R17155 OUT_N.n561 OUT_N.n560 0.00527411
R17156 OUT_N.n339 OUT_N.n338 0.00527411
R17157 OUT_N.n330 OUT_N.n329 0.00527411
R17158 OUT_N.n24 OUT_N.n23 0.00527411
R17159 OUT_N.n25 OUT_N.n24 0.00527411
R17160 OUT_N.n1713 OUT_N.n1712 0.00527411
R17161 OUT_N.n1722 OUT_N.n1713 0.00527411
R17162 OUT_N.n1799 OUT_N.n1798 0.00527411
R17163 OUT_N.n1794 OUT_N.n1793 0.00527411
R17164 OUT_N.n1795 OUT_N.n1794 0.00527411
R17165 OUT_N.n1800 OUT_N.n1799 0.00527411
R17166 OUT_N.n1753 OUT_N.n1752 0.00527411
R17167 OUT_N.n1754 OUT_N.n1753 0.00527411
R17168 OUT_N.n2229 OUT_N.n2228 0.00527411
R17169 OUT_N.n2220 OUT_N.n2219 0.00527411
R17170 OUT_N.n2211 OUT_N.n2210 0.00527411
R17171 OUT_N.n2036 OUT_N.n2035 0.00527411
R17172 OUT_N.n2035 OUT_N.n2034 0.00527411
R17173 OUT_N.n2210 OUT_N.n2209 0.00527411
R17174 OUT_N.n2219 OUT_N.n2218 0.00527411
R17175 OUT_N.n2228 OUT_N.n2227 0.00527411
R17176 OUT_N.n2084 OUT_N.n2083 0.00525899
R17177 OUT_N.n2086 OUT_N.n2085 0.00525899
R17178 OUT_N.n1925 OUT_N.n1924 0.00525899
R17179 OUT_N.n1921 OUT_N.n1920 0.00525899
R17180 OUT_N.n2159 OUT_N.n2158 0.00525899
R17181 OUT_N.n2164 OUT_N.n2163 0.00525899
R17182 OUT_N.n1957 OUT_N.n1956 0.00525899
R17183 OUT_N.n1952 OUT_N.n1951 0.00525899
R17184 OUT_N.n2111 OUT_N.n2110 0.00525899
R17185 OUT_N.n2113 OUT_N.n2112 0.00525899
R17186 OUT_N.n1879 OUT_N.n1878 0.00525899
R17187 OUT_N.n1877 OUT_N.n1876 0.00525899
R17188 OUT_N.n1123 OUT_N.n1122 0.00525899
R17189 OUT_N.n1125 OUT_N.n1124 0.00525899
R17190 OUT_N.n1132 OUT_N.n1131 0.00525899
R17191 OUT_N.n1134 OUT_N.n1133 0.00525899
R17192 OUT_N.n1163 OUT_N.n1162 0.00525899
R17193 OUT_N.n1165 OUT_N.n1164 0.00525899
R17194 OUT_N.n1172 OUT_N.n1171 0.00525899
R17195 OUT_N.n1174 OUT_N.n1173 0.00525899
R17196 OUT_N.n1181 OUT_N.n1180 0.00525899
R17197 OUT_N.n1183 OUT_N.n1182 0.00525899
R17198 OUT_N.n1190 OUT_N.n1189 0.00525899
R17199 OUT_N.n1192 OUT_N.n1191 0.00525899
R17200 OUT_N.n1209 OUT_N.n1208 0.00525899
R17201 OUT_N.n1211 OUT_N.n1210 0.00525899
R17202 OUT_N.n1218 OUT_N.n1217 0.00525899
R17203 OUT_N.n1220 OUT_N.n1219 0.00525899
R17204 OUT_N.n1227 OUT_N.n1226 0.00525899
R17205 OUT_N.n1229 OUT_N.n1228 0.00525899
R17206 OUT_N.n1236 OUT_N.n1235 0.00525899
R17207 OUT_N.n1238 OUT_N.n1237 0.00525899
R17208 OUT_N.n1265 OUT_N.n1264 0.00525899
R17209 OUT_N.n1267 OUT_N.n1266 0.00525899
R17210 OUT_N.n1274 OUT_N.n1273 0.00525899
R17211 OUT_N.n1276 OUT_N.n1275 0.00525899
R17212 OUT_N.n1283 OUT_N.n1282 0.00525899
R17213 OUT_N.n1285 OUT_N.n1284 0.00525899
R17214 OUT_N.n1292 OUT_N.n1291 0.00525899
R17215 OUT_N.n1294 OUT_N.n1293 0.00525899
R17216 OUT_N.n1460 OUT_N.n1459 0.00525899
R17217 OUT_N.n1462 OUT_N.n1461 0.00525899
R17218 OUT_N.n1469 OUT_N.n1468 0.00525899
R17219 OUT_N.n1471 OUT_N.n1470 0.00525899
R17220 OUT_N.n1504 OUT_N.n1503 0.00525899
R17221 OUT_N.n1506 OUT_N.n1505 0.00525899
R17222 OUT_N.n1513 OUT_N.n1512 0.00525899
R17223 OUT_N.n1515 OUT_N.n1514 0.00525899
R17224 OUT_N.n1522 OUT_N.n1521 0.00525899
R17225 OUT_N.n1524 OUT_N.n1523 0.00525899
R17226 OUT_N.n1531 OUT_N.n1530 0.00525899
R17227 OUT_N.n1533 OUT_N.n1532 0.00525899
R17228 OUT_N.n1584 OUT_N.n1583 0.00525899
R17229 OUT_N.n1586 OUT_N.n1585 0.00525899
R17230 OUT_N.n1593 OUT_N.n1592 0.00525899
R17231 OUT_N.n1595 OUT_N.n1594 0.00525899
R17232 OUT_N.n1602 OUT_N.n1601 0.00525899
R17233 OUT_N.n1604 OUT_N.n1603 0.00525899
R17234 OUT_N.n1611 OUT_N.n1610 0.00525899
R17235 OUT_N.n1613 OUT_N.n1612 0.00525899
R17236 OUT_N.n1637 OUT_N.n1636 0.00525899
R17237 OUT_N.n1639 OUT_N.n1638 0.00525899
R17238 OUT_N.n1646 OUT_N.n1645 0.00525899
R17239 OUT_N.n1648 OUT_N.n1647 0.00525899
R17240 OUT_N.n1655 OUT_N.n1654 0.00525899
R17241 OUT_N.n1657 OUT_N.n1656 0.00525899
R17242 OUT_N.n1664 OUT_N.n1663 0.00525899
R17243 OUT_N.n1666 OUT_N.n1665 0.00525899
R17244 OUT_N.n788 OUT_N.n787 0.00525899
R17245 OUT_N.n790 OUT_N.n789 0.00525899
R17246 OUT_N.n797 OUT_N.n796 0.00525899
R17247 OUT_N.n799 OUT_N.n798 0.00525899
R17248 OUT_N.n816 OUT_N.n815 0.00525899
R17249 OUT_N.n818 OUT_N.n817 0.00525899
R17250 OUT_N.n825 OUT_N.n824 0.00525899
R17251 OUT_N.n827 OUT_N.n826 0.00525899
R17252 OUT_N.n834 OUT_N.n833 0.00525899
R17253 OUT_N.n836 OUT_N.n835 0.00525899
R17254 OUT_N.n843 OUT_N.n842 0.00525899
R17255 OUT_N.n845 OUT_N.n844 0.00525899
R17256 OUT_N.n860 OUT_N.n859 0.00525899
R17257 OUT_N.n862 OUT_N.n861 0.00525899
R17258 OUT_N.n869 OUT_N.n868 0.00525899
R17259 OUT_N.n871 OUT_N.n870 0.00525899
R17260 OUT_N.n878 OUT_N.n877 0.00525899
R17261 OUT_N.n880 OUT_N.n879 0.00525899
R17262 OUT_N.n887 OUT_N.n886 0.00525899
R17263 OUT_N.n889 OUT_N.n888 0.00525899
R17264 OUT_N.n906 OUT_N.n905 0.00525899
R17265 OUT_N.n908 OUT_N.n907 0.00525899
R17266 OUT_N.n915 OUT_N.n914 0.00525899
R17267 OUT_N.n917 OUT_N.n916 0.00525899
R17268 OUT_N.n924 OUT_N.n923 0.00525899
R17269 OUT_N.n926 OUT_N.n925 0.00525899
R17270 OUT_N.n933 OUT_N.n932 0.00525899
R17271 OUT_N.n935 OUT_N.n934 0.00525899
R17272 OUT_N.n332 OUT_N.n331 0.00525899
R17273 OUT_N.n334 OUT_N.n333 0.00525899
R17274 OUT_N.n341 OUT_N.n340 0.00525899
R17275 OUT_N.n343 OUT_N.n342 0.00525899
R17276 OUT_N.n369 OUT_N.n368 0.00525899
R17277 OUT_N.n371 OUT_N.n370 0.00525899
R17278 OUT_N.n378 OUT_N.n377 0.00525899
R17279 OUT_N.n380 OUT_N.n379 0.00525899
R17280 OUT_N.n387 OUT_N.n386 0.00525899
R17281 OUT_N.n389 OUT_N.n388 0.00525899
R17282 OUT_N.n396 OUT_N.n395 0.00525899
R17283 OUT_N.n398 OUT_N.n397 0.00525899
R17284 OUT_N.n418 OUT_N.n417 0.00525899
R17285 OUT_N.n420 OUT_N.n419 0.00525899
R17286 OUT_N.n427 OUT_N.n426 0.00525899
R17287 OUT_N.n429 OUT_N.n428 0.00525899
R17288 OUT_N.n436 OUT_N.n435 0.00525899
R17289 OUT_N.n438 OUT_N.n437 0.00525899
R17290 OUT_N.n445 OUT_N.n444 0.00525899
R17291 OUT_N.n447 OUT_N.n446 0.00525899
R17292 OUT_N.n471 OUT_N.n470 0.00525899
R17293 OUT_N.n473 OUT_N.n472 0.00525899
R17294 OUT_N.n480 OUT_N.n479 0.00525899
R17295 OUT_N.n482 OUT_N.n481 0.00525899
R17296 OUT_N.n489 OUT_N.n488 0.00525899
R17297 OUT_N.n491 OUT_N.n490 0.00525899
R17298 OUT_N.n498 OUT_N.n497 0.00525899
R17299 OUT_N.n500 OUT_N.n499 0.00525899
R17300 OUT_N.n602 OUT_N.n601 0.00525899
R17301 OUT_N.n595 OUT_N.n594 0.00525899
R17302 OUT_N.n593 OUT_N.n592 0.00525899
R17303 OUT_N.n586 OUT_N.n585 0.00525899
R17304 OUT_N.n584 OUT_N.n583 0.00525899
R17305 OUT_N.n577 OUT_N.n576 0.00525899
R17306 OUT_N.n566 OUT_N.n565 0.00525899
R17307 OUT_N.n559 OUT_N.n558 0.00525899
R17308 OUT_N.n557 OUT_N.n556 0.00525899
R17309 OUT_N.n1704 OUT_N.n1703 0.00525899
R17310 OUT_N.n1797 OUT_N.n1796 0.00525899
R17311 OUT_N.n1802 OUT_N.n1801 0.00525899
R17312 OUT_N.n2226 OUT_N.n2225 0.00525899
R17313 OUT_N.n2224 OUT_N.n2223 0.00525899
R17314 OUT_N.n2217 OUT_N.n2216 0.00525899
R17315 OUT_N.n2215 OUT_N.n2214 0.00525899
R17316 OUT_N.n2208 OUT_N.n2207 0.00525899
R17317 OUT_N.n2206 OUT_N.n2205 0.00525899
R17318 OUT_N.n2033 OUT_N.n2032 0.00525899
R17319 OUT_N.n2031 OUT_N.n2030 0.00525899
R17320 OUT_N.n2027 OUT_N.n2026 0.00525899
R17321 OUT_N.n153 OUT_N.n152 0.00495689
R17322 OUT_N.n159 OUT_N.n158 0.00495689
R17323 OUT_N.n162 OUT_N.n161 0.00495689
R17324 OUT_N.n140 OUT_N.n139 0.00495689
R17325 OUT_N.n145 OUT_N.n131 0.00495689
R17326 OUT_N.n168 OUT_N.n167 0.00495689
R17327 OUT_N.n156 OUT_N.n155 0.00495689
R17328 OUT_N.n137 OUT_N.n136 0.00495689
R17329 OUT_N.n54 OUT_N.n53 0.00495689
R17330 OUT_N.n66 OUT_N.n59 0.00495689
R17331 OUT_N.n116 OUT_N.n115 0.00495689
R17332 OUT_N.n110 OUT_N.n109 0.00495689
R17333 OUT_N.n113 OUT_N.n112 0.00495689
R17334 OUT_N.n91 OUT_N.n73 0.00495689
R17335 OUT_N.n97 OUT_N.n96 0.00429028
R17336 OUT_N.n105 OUT_N.n104 0.00429028
R17337 OUT_N.n94 OUT_N.n93 0.00429028
R17338 OUT_N.n2156 OUT_N.n2151 0.00418876
R17339 OUT_N.n2190 OUT_N.n2183 0.00418876
R17340 OUT_N.n1996 OUT_N.n1995 0.00418876
R17341 OUT_N.n1991 OUT_N.n1990 0.00418876
R17342 OUT_N.n26 OUT_N.n25 0.00418876
R17343 OUT_N.n21 OUT_N.n20 0.00418876
R17344 OUT_N.n1723 OUT_N.n1722 0.00418876
R17345 OUT_N.n1791 OUT_N.n1790 0.00418876
R17346 OUT_N.n1755 OUT_N.n1754 0.00418876
R17347 OUT_N.n1750 OUT_N.n1749 0.00418876
R17348 OUT_N.n65 OUT_N.n61 0.00346816
R17349 OUT_N.n64 OUT_N.n63 0.00346816
R17350 OUT_N.n89 OUT_N.n88 0.00346816
R17351 OUT_N.n85 OUT_N.n84 0.00346816
R17352 OUT_N.n83 OUT_N.n82 0.00346816
R17353 OUT_N.n79 OUT_N.n78 0.00346816
R17354 OUT_N.n77 OUT_N.n76 0.00346816
R17355 OUT_N.n165 OUT_N.n164 0.00346816
R17356 OUT_N.n144 OUT_N.n135 0.00346816
R17357 OUT_N.n143 OUT_N.n142 0.00346816
R17358 OUT_N.n108 OUT_N.n107 0.00346816
R17359 OUT_N.n120 OUT_N.n119 0.00346816
R17360 OUT_N.n122 OUT_N.n121 0.00346816
R17361 OUT_N.n127 OUT_N.n125 0.00346816
R17362 OUT_N.n129 OUT_N.n128 0.00346816
R17363 OUT_N.n135 OUT_N.n134 0.00346816
R17364 OUT_N.n107 OUT_N.n106 0.00346816
R17365 OUT_N.n119 OUT_N.n118 0.00346816
R17366 OUT_N.n125 OUT_N.n124 0.00346816
R17367 OUT_N.n121 OUT_N.n120 0.00346816
R17368 OUT_N.n166 OUT_N.n165 0.00346816
R17369 OUT_N.n144 OUT_N.n143 0.00346816
R17370 OUT_N.n128 OUT_N.n127 0.00346816
R17371 OUT_N.n37 OUT_N.n36 0.00346816
R17372 OUT_N.n39 OUT_N.n38 0.00346816
R17373 OUT_N.n43 OUT_N.n42 0.00346816
R17374 OUT_N.n45 OUT_N.n44 0.00346816
R17375 OUT_N.n49 OUT_N.n48 0.00346816
R17376 OUT_N.n51 OUT_N.n50 0.00346816
R17377 OUT_N.n57 OUT_N.n56 0.00346816
R17378 OUT_N.n84 OUT_N.n83 0.00346816
R17379 OUT_N.n50 OUT_N.n49 0.00346816
R17380 OUT_N.n90 OUT_N.n89 0.00346816
R17381 OUT_N.n44 OUT_N.n43 0.00346816
R17382 OUT_N.n38 OUT_N.n37 0.00346816
R17383 OUT_N.n36 OUT_N.n35 0.00346816
R17384 OUT_N.n86 OUT_N.n85 0.00346816
R17385 OUT_N.n42 OUT_N.n41 0.00346816
R17386 OUT_N.n65 OUT_N.n64 0.00346816
R17387 OUT_N.n61 OUT_N.n60 0.00346816
R17388 OUT_N.n78 OUT_N.n77 0.00346816
R17389 OUT_N.n80 OUT_N.n79 0.00346816
R17390 OUT_N.n48 OUT_N.n47 0.00346816
R17391 OUT_N.n56 OUT_N.n55 0.00346816
R17392 OUT_N.n1710 OUT_N.n1705 0.00314088
R17393 OUT_N.n114 OUT_N.n113 0.00297812
R17394 OUT_N.n161 OUT_N.n160 0.00297812
R17395 OUT_N.n166 OUT_N.n159 0.00297812
R17396 OUT_N.n151 OUT_N.n145 0.00297812
R17397 OUT_N.n154 OUT_N.n153 0.00297812
R17398 OUT_N.n155 OUT_N.n154 0.00297812
R17399 OUT_N.n115 OUT_N.n114 0.00297812
R17400 OUT_N.n138 OUT_N.n137 0.00297812
R17401 OUT_N.n109 OUT_N.n108 0.00297812
R17402 OUT_N.n139 OUT_N.n138 0.00297812
R17403 OUT_N.n167 OUT_N.n151 0.00297812
R17404 OUT_N.n92 OUT_N.n66 0.00297812
R17405 OUT_N.n55 OUT_N.n54 0.00297812
R17406 OUT_N.n91 OUT_N.n90 0.00297812
R17407 OUT_N.n2151 OUT_N.n2150 0.00284163
R17408 OUT_N.n2025 OUT_N.n2024 0.00281899
R17409 OUT_N.n103 OUT_N.n94 0.00264514
R17410 OUT_N.n104 OUT_N.n92 0.00264514
R17411 OUT_N.n103 OUT_N.n97 0.00264514
R17412 OUT_N.n1990 OUT_N.n1989 0.00219433
R17413 OUT_N.n20 OUT_N.n19 0.00219433
R17414 OUT_N.n1790 OUT_N.n1789 0.00219433
R17415 OUT_N.n1749 OUT_N.n1748 0.00219433
R17416 OUT_N.n1915 OUT_N.n1914 0.00192237
R17417 OUT_N.n1701 OUT_N.n1700 0.00192237
R17418 OUT_N.n2180 OUT_N.n2179 0.00192078
R17419 OUT_P.n1101 OUT_P.t231 6.959
R17420 OUT_P.n1104 OUT_P.n1103 2.40737
R17421 OUT_P.n549 OUT_P.n546 1.84464
R17422 OUT_P.n928 OUT_P.n927 1.76234
R17423 OUT_P.n943 OUT_P.n942 1.76234
R17424 OUT_P.n537 OUT_P.n196 1.49643
R17425 OUT_P.n446 OUT_P.n199 1.49371
R17426 OUT_P.n445 OUT_P.n201 1.49371
R17427 OUT_P.n538 OUT_P.n194 1.49371
R17428 OUT_P.n971 OUT_P.n934 1.49371
R17429 OUT_P.n1921 OUT_P.n541 1.49371
R17430 OUT_P.n958 OUT_P.n957 1.47979
R17431 OUT_P.n922 OUT_P.n921 1.47979
R17432 OUT_P.n937 OUT_P.n936 1.47979
R17433 OUT_P.n982 OUT_P.n981 1.47979
R17434 OUT_P.n914 OUT_P.n913 1.47979
R17435 OUT_P.n906 OUT_P.n905 1.47979
R17436 OUT_P.n1458 OUT_P.n1457 1.46987
R17437 OUT_P.n1468 OUT_P.t13 1.46987
R17438 OUT_P.n1473 OUT_P.n1472 1.46987
R17439 OUT_P.n1497 OUT_P.t14 1.46987
R17440 OUT_P.n1488 OUT_P.n1487 1.46987
R17441 OUT_P.n1483 OUT_P.t28 1.46987
R17442 OUT_P.n6 OUT_P.t263 1.46987
R17443 OUT_P.n27 OUT_P.n26 1.46987
R17444 OUT_P.n132 OUT_P.t242 1.46987
R17445 OUT_P.n153 OUT_P.n152 1.46987
R17446 OUT_P.n162 OUT_P.t261 1.46987
R17447 OUT_P.n183 OUT_P.n182 1.46987
R17448 OUT_P.n1705 OUT_P.n1704 1.43193
R17449 OUT_P.n1688 OUT_P.t47 1.43193
R17450 OUT_P.n1684 OUT_P.n1683 1.43193
R17451 OUT_P.n1667 OUT_P.t204 1.43193
R17452 OUT_P.n1663 OUT_P.n1662 1.43193
R17453 OUT_P.n1646 OUT_P.t197 1.43193
R17454 OUT_P.n1642 OUT_P.n1641 1.43193
R17455 OUT_P.n1625 OUT_P.t149 1.43193
R17456 OUT_P.n1621 OUT_P.n1620 1.43193
R17457 OUT_P.n1891 OUT_P.t219 1.43193
R17458 OUT_P.n1860 OUT_P.n1859 1.43193
R17459 OUT_P.n1850 OUT_P.t174 1.43193
R17460 OUT_P.n1819 OUT_P.n1818 1.43193
R17461 OUT_P.n1604 OUT_P.t137 1.43193
R17462 OUT_P.n712 OUT_P.n711 1.43193
R17463 OUT_P.n695 OUT_P.t165 1.43193
R17464 OUT_P.n691 OUT_P.n690 1.43193
R17465 OUT_P.n674 OUT_P.t132 1.43193
R17466 OUT_P.n670 OUT_P.n669 1.43193
R17467 OUT_P.n653 OUT_P.t185 1.43193
R17468 OUT_P.n649 OUT_P.n648 1.43193
R17469 OUT_P.n632 OUT_P.t152 1.43193
R17470 OUT_P.n628 OUT_P.n627 1.43193
R17471 OUT_P.n611 OUT_P.t158 1.43193
R17472 OUT_P.n607 OUT_P.n606 1.43193
R17473 OUT_P.n590 OUT_P.t35 1.43193
R17474 OUT_P.n586 OUT_P.n585 1.43193
R17475 OUT_P.n569 OUT_P.t229 1.43193
R17476 OUT_P.n929 OUT_P.n928 1.3488
R17477 OUT_P.n944 OUT_P.n943 1.3488
R17478 OUT_P.n952 OUT_P.n951 1.28777
R17479 OUT_P.n986 OUT_P.n985 1.28777
R17480 OUT_P.n561 OUT_P.n560 1.28752
R17481 OUT_P.n1070 OUT_P.n1063 1.26239
R17482 OUT_P.n955 OUT_P.n954 1.21718
R17483 OUT_P.n992 OUT_P.n991 1.21718
R17484 OUT_P.n207 OUT_P.n204 1.19506
R17485 OUT_P.n217 OUT_P.n216 1.19506
R17486 OUT_P.n228 OUT_P.n227 1.19506
R17487 OUT_P.n239 OUT_P.n238 1.19506
R17488 OUT_P.n265 OUT_P.n264 1.19506
R17489 OUT_P.n276 OUT_P.n275 1.19506
R17490 OUT_P.n287 OUT_P.n286 1.19506
R17491 OUT_P.n298 OUT_P.n297 1.19506
R17492 OUT_P.n309 OUT_P.n308 1.19506
R17493 OUT_P.n320 OUT_P.n319 1.19506
R17494 OUT_P.n331 OUT_P.n330 1.19506
R17495 OUT_P.n342 OUT_P.n341 1.19506
R17496 OUT_P.n362 OUT_P.n361 1.19506
R17497 OUT_P.n373 OUT_P.n372 1.19506
R17498 OUT_P.n384 OUT_P.n383 1.19506
R17499 OUT_P.n395 OUT_P.n394 1.19506
R17500 OUT_P.n406 OUT_P.n405 1.19506
R17501 OUT_P.n417 OUT_P.n416 1.19506
R17502 OUT_P.n428 OUT_P.n427 1.19506
R17503 OUT_P.n439 OUT_P.n438 1.19506
R17504 OUT_P.n454 OUT_P.n453 1.19506
R17505 OUT_P.n465 OUT_P.n464 1.19506
R17506 OUT_P.n476 OUT_P.n475 1.19506
R17507 OUT_P.n487 OUT_P.n486 1.19506
R17508 OUT_P.n498 OUT_P.n497 1.19506
R17509 OUT_P.n509 OUT_P.n508 1.19506
R17510 OUT_P.n520 OUT_P.n519 1.19506
R17511 OUT_P.n531 OUT_P.n530 1.19506
R17512 OUT_P.n1932 OUT_P.n1931 1.1949
R17513 OUT_P.n1939 OUT_P.n1936 1.1949
R17514 OUT_P.n1298 OUT_P.n1297 1.1948
R17515 OUT_P.n1286 OUT_P.n1285 1.1948
R17516 OUT_P.n1274 OUT_P.n1273 1.1948
R17517 OUT_P.n1262 OUT_P.n1261 1.1948
R17518 OUT_P.n1250 OUT_P.n1249 1.1948
R17519 OUT_P.n1238 OUT_P.n1237 1.1948
R17520 OUT_P.n1226 OUT_P.n1225 1.1948
R17521 OUT_P.n1214 OUT_P.n1213 1.1948
R17522 OUT_P.n1202 OUT_P.n1201 1.1948
R17523 OUT_P.n1190 OUT_P.n1189 1.1948
R17524 OUT_P.n1178 OUT_P.n1177 1.1948
R17525 OUT_P.n1166 OUT_P.n1165 1.1948
R17526 OUT_P.n1154 OUT_P.n1153 1.1948
R17527 OUT_P.n1142 OUT_P.n1141 1.1948
R17528 OUT_P.n1689 OUT_P.n1688 1.19473
R17529 OUT_P.n1668 OUT_P.n1667 1.19473
R17530 OUT_P.n1647 OUT_P.n1646 1.19473
R17531 OUT_P.n1626 OUT_P.n1625 1.19473
R17532 OUT_P.n1605 OUT_P.n1604 1.19473
R17533 OUT_P.n713 OUT_P.n712 1.19473
R17534 OUT_P.n692 OUT_P.n691 1.19473
R17535 OUT_P.n671 OUT_P.n670 1.19473
R17536 OUT_P.n650 OUT_P.n649 1.19473
R17537 OUT_P.n629 OUT_P.n628 1.19473
R17538 OUT_P.n608 OUT_P.n607 1.19473
R17539 OUT_P.n587 OUT_P.n586 1.19473
R17540 OUT_P.n1112 OUT_P.n1111 1.19461
R17541 OUT_P.n1553 OUT_P.n1552 1.19461
R17542 OUT_P.n1523 OUT_P.n1522 1.19461
R17543 OUT_P.n43 OUT_P.n42 1.19461
R17544 OUT_P.n1474 OUT_P.n1473 1.19458
R17545 OUT_P.n1484 OUT_P.n1483 1.19458
R17546 OUT_P.n7 OUT_P.n6 1.19458
R17547 OUT_P.n28 OUT_P.n27 1.19458
R17548 OUT_P.n133 OUT_P.n132 1.19458
R17549 OUT_P.n154 OUT_P.n153 1.19458
R17550 OUT_P.n163 OUT_P.n162 1.19458
R17551 OUT_P.n184 OUT_P.n183 1.19458
R17552 OUT_P.n74 OUT_P.n73 1.19458
R17553 OUT_P.n1701 OUT_P.n1700 1.19445
R17554 OUT_P.n1680 OUT_P.n1679 1.19445
R17555 OUT_P.n1659 OUT_P.n1658 1.19445
R17556 OUT_P.n1638 OUT_P.n1637 1.19445
R17557 OUT_P.n1617 OUT_P.n1616 1.19445
R17558 OUT_P.n702 OUT_P.n701 1.19445
R17559 OUT_P.n681 OUT_P.n680 1.19445
R17560 OUT_P.n660 OUT_P.n659 1.19445
R17561 OUT_P.n639 OUT_P.n638 1.19445
R17562 OUT_P.n618 OUT_P.n617 1.19445
R17563 OUT_P.n597 OUT_P.n596 1.19445
R17564 OUT_P.n576 OUT_P.n575 1.19445
R17565 OUT_P.n1465 OUT_P.n1464 1.19426
R17566 OUT_P.n1495 OUT_P.n1494 1.19426
R17567 OUT_P.n18 OUT_P.n17 1.19426
R17568 OUT_P.n144 OUT_P.n143 1.19426
R17569 OUT_P.n174 OUT_P.n173 1.19426
R17570 OUT_P.n1095 OUT_P.n1094 1.18729
R17571 OUT_P.n1480 OUT_P.n1479 1.17959
R17572 OUT_P.n1459 OUT_P.n1458 1.1793
R17573 OUT_P.n1469 OUT_P.n1468 1.1793
R17574 OUT_P.n1500 OUT_P.n1497 1.1793
R17575 OUT_P.n1489 OUT_P.n1488 1.1793
R17576 OUT_P.n1695 OUT_P.n1694 1.1791
R17577 OUT_P.n1674 OUT_P.n1673 1.1791
R17578 OUT_P.n1653 OUT_P.n1652 1.1791
R17579 OUT_P.n1632 OUT_P.n1631 1.1791
R17580 OUT_P.n1611 OUT_P.n1610 1.1791
R17581 OUT_P.n1883 OUT_P.n1882 1.1791
R17582 OUT_P.n1872 OUT_P.n1871 1.1791
R17583 OUT_P.n1842 OUT_P.n1841 1.1791
R17584 OUT_P.n1831 OUT_P.n1830 1.1791
R17585 OUT_P.n708 OUT_P.n707 1.1791
R17586 OUT_P.n687 OUT_P.n686 1.1791
R17587 OUT_P.n666 OUT_P.n665 1.1791
R17588 OUT_P.n645 OUT_P.n644 1.1791
R17589 OUT_P.n624 OUT_P.n623 1.1791
R17590 OUT_P.n603 OUT_P.n602 1.1791
R17591 OUT_P.n582 OUT_P.n581 1.1791
R17592 OUT_P.n1118 OUT_P.n1117 1.17896
R17593 OUT_P.n1529 OUT_P.n1528 1.17896
R17594 OUT_P.n1547 OUT_P.n1546 1.17896
R17595 OUT_P.n49 OUT_P.n48 1.17896
R17596 OUT_P.n67 OUT_P.n66 1.17896
R17597 OUT_P.n1706 OUT_P.n1705 1.17884
R17598 OUT_P.n1685 OUT_P.n1684 1.17884
R17599 OUT_P.n1664 OUT_P.n1663 1.17884
R17600 OUT_P.n1643 OUT_P.n1642 1.17884
R17601 OUT_P.n1622 OUT_P.n1621 1.17884
R17602 OUT_P.n1892 OUT_P.n1891 1.17884
R17603 OUT_P.n1861 OUT_P.n1860 1.17884
R17604 OUT_P.n1851 OUT_P.n1850 1.17884
R17605 OUT_P.n1820 OUT_P.n1819 1.17884
R17606 OUT_P.n696 OUT_P.n695 1.17884
R17607 OUT_P.n675 OUT_P.n674 1.17884
R17608 OUT_P.n654 OUT_P.n653 1.17884
R17609 OUT_P.n633 OUT_P.n632 1.17884
R17610 OUT_P.n612 OUT_P.n611 1.17884
R17611 OUT_P.n591 OUT_P.n590 1.17884
R17612 OUT_P.n570 OUT_P.n569 1.17884
R17613 OUT_P.n1292 OUT_P.n1291 1.17849
R17614 OUT_P.n1280 OUT_P.n1279 1.17849
R17615 OUT_P.n1268 OUT_P.n1267 1.17849
R17616 OUT_P.n1256 OUT_P.n1255 1.17849
R17617 OUT_P.n1244 OUT_P.n1243 1.17849
R17618 OUT_P.n1232 OUT_P.n1231 1.17849
R17619 OUT_P.n1220 OUT_P.n1219 1.17849
R17620 OUT_P.n1208 OUT_P.n1207 1.17849
R17621 OUT_P.n1196 OUT_P.n1195 1.17849
R17622 OUT_P.n1184 OUT_P.n1183 1.17849
R17623 OUT_P.n1172 OUT_P.n1171 1.17849
R17624 OUT_P.n1160 OUT_P.n1159 1.17849
R17625 OUT_P.n1148 OUT_P.n1147 1.17849
R17626 OUT_P.n1136 OUT_P.n1135 1.17849
R17627 OUT_P.n562 OUT_P.n561 1.17419
R17628 OUT_P.n550 OUT_P.n549 1.14437
R17629 OUT_P.n923 OUT_P.n922 1.14073
R17630 OUT_P.n938 OUT_P.n937 1.14073
R17631 OUT_P.n983 OUT_P.n982 1.14073
R17632 OUT_P.n915 OUT_P.n914 1.14073
R17633 OUT_P.n907 OUT_P.n906 1.14073
R17634 OUT_P.n354 OUT_P.n353 1.1353
R17635 OUT_P.n1926 OUT_P.n1925 1.12925
R17636 OUT_P.n208 OUT_P.n207 1.12829
R17637 OUT_P.n105 OUT_P.n104 1.12829
R17638 OUT_P.n551 OUT_P.n550 1.12829
R17639 OUT_P.n1501 OUT_P.n1500 1.12829
R17640 OUT_P.n1940 OUT_P.n1939 1.12795
R17641 OUT_P.n961 OUT_P.n960 1.12795
R17642 OUT_P.n75 OUT_P.n74 1.12758
R17643 OUT_P.n960 OUT_P.n959 1.1255
R17644 OUT_P.n931 OUT_P.n930 1.1255
R17645 OUT_P.n946 OUT_P.n945 1.1255
R17646 OUT_P.n990 OUT_P.n989 1.1255
R17647 OUT_P.n994 OUT_P.n993 1.1255
R17648 OUT_P.n918 OUT_P.n917 1.1255
R17649 OUT_P.n558 OUT_P.n557 1.1255
R17650 OUT_P.n910 OUT_P.n909 1.1255
R17651 OUT_P.n1062 OUT_P.n1061 1.12145
R17652 OUT_P.n1062 OUT_P.n1057 1.12145
R17653 OUT_P.n1052 OUT_P.n1049 1.12145
R17654 OUT_P.n1052 OUT_P.n1051 1.12145
R17655 OUT_P.n1093 OUT_P.n1092 1.12145
R17656 OUT_P.n1086 OUT_P.n1085 1.12145
R17657 OUT_P.n902 OUT_P.n901 1.11801
R17658 OUT_P.n842 OUT_P.n841 1.11801
R17659 OUT_P.n845 OUT_P.n844 1.11801
R17660 OUT_P.n121 OUT_P.n114 1.11801
R17661 OUT_P.n258 OUT_P.n257 1.11801
R17662 OUT_P.n1325 OUT_P.n1324 1.11801
R17663 OUT_P.n1907 OUT_P.n1010 1.11801
R17664 OUT_P.n1913 OUT_P.n567 1.11801
R17665 OUT_P.n1951 OUT_P.n1950 1.11801
R17666 OUT_P.n1601 OUT_P.n1600 1.11801
R17667 OUT_P.n1103 OUT_P.n1096 1.11801
R17668 OUT_P.n791 OUT_P.n790 1.11782
R17669 OUT_P.n85 OUT_P.n84 1.11782
R17670 OUT_P.n128 OUT_P.n127 1.11782
R17671 OUT_P.n1565 OUT_P.n1564 1.11782
R17672 OUT_P.n1541 OUT_P.n1540 1.11782
R17673 OUT_P.n61 OUT_P.n60 1.11782
R17674 OUT_P.n1571 OUT_P.n1570 1.11782
R17675 OUT_P.n1733 OUT_P.n1732 1.11782
R17676 OUT_P.n1322 OUT_P.n1321 1.11782
R17677 OUT_P.n1451 OUT_P.n1450 1.11782
R17678 OUT_P.n1130 OUT_P.n1129 1.11782
R17679 OUT_P.n1912 OUT_P.n1911 1.11782
R17680 OUT_P.n1903 OUT_P.n1902 1.11782
R17681 OUT_P.n1102 OUT_P.n1101 1.11782
R17682 OUT_P.n1953 OUT_P.n1952 1.11782
R17683 OUT_P.n998 OUT_P.n997 1.03835
R17684 OUT_P.n73 OUT_P.n72 0.923874
R17685 OUT_P.n1111 OUT_P.n1110 0.923611
R17686 OUT_P.n1552 OUT_P.n1551 0.923611
R17687 OUT_P.n1522 OUT_P.n1521 0.923611
R17688 OUT_P.n42 OUT_P.n41 0.923611
R17689 OUT_P.n1931 OUT_P.n1930 0.923589
R17690 OUT_P.n1936 OUT_P.n1935 0.923589
R17691 OUT_P.n1117 OUT_P.n1116 0.923589
R17692 OUT_P.n1528 OUT_P.n1527 0.923589
R17693 OUT_P.n1546 OUT_P.n1545 0.923589
R17694 OUT_P.n48 OUT_P.n47 0.923589
R17695 OUT_P.n66 OUT_P.n65 0.923589
R17696 OUT_P.n1464 OUT_P.n1463 0.923538
R17697 OUT_P.n1479 OUT_P.n1478 0.923538
R17698 OUT_P.n1494 OUT_P.n1493 0.923538
R17699 OUT_P.n17 OUT_P.n16 0.923538
R17700 OUT_P.n143 OUT_P.n142 0.923538
R17701 OUT_P.n173 OUT_P.n172 0.923538
R17702 OUT_P.n1946 OUT_P.n1933 0.885703
R17703 OUT_P.n564 OUT_P.n563 0.885703
R17704 OUT_P.n533 OUT_P.n532 0.885703
R17705 OUT_P.n522 OUT_P.n521 0.885703
R17706 OUT_P.n511 OUT_P.n510 0.885703
R17707 OUT_P.n500 OUT_P.n499 0.885703
R17708 OUT_P.n489 OUT_P.n488 0.885703
R17709 OUT_P.n478 OUT_P.n477 0.885703
R17710 OUT_P.n467 OUT_P.n466 0.885703
R17711 OUT_P.n456 OUT_P.n455 0.885703
R17712 OUT_P.n441 OUT_P.n440 0.885703
R17713 OUT_P.n430 OUT_P.n429 0.885703
R17714 OUT_P.n419 OUT_P.n418 0.885703
R17715 OUT_P.n408 OUT_P.n407 0.885703
R17716 OUT_P.n397 OUT_P.n396 0.885703
R17717 OUT_P.n386 OUT_P.n385 0.885703
R17718 OUT_P.n375 OUT_P.n374 0.885703
R17719 OUT_P.n364 OUT_P.n363 0.885703
R17720 OUT_P.n344 OUT_P.n343 0.885703
R17721 OUT_P.n333 OUT_P.n332 0.885703
R17722 OUT_P.n322 OUT_P.n321 0.885703
R17723 OUT_P.n311 OUT_P.n310 0.885703
R17724 OUT_P.n300 OUT_P.n299 0.885703
R17725 OUT_P.n289 OUT_P.n288 0.885703
R17726 OUT_P.n278 OUT_P.n277 0.885703
R17727 OUT_P.n267 OUT_P.n266 0.885703
R17728 OUT_P.n241 OUT_P.n240 0.885703
R17729 OUT_P.n230 OUT_P.n229 0.885703
R17730 OUT_P.n219 OUT_P.n218 0.885703
R17731 OUT_P.n1822 OUT_P.n1821 0.885703
R17732 OUT_P.n1833 OUT_P.n1832 0.885703
R17733 OUT_P.n1844 OUT_P.n1843 0.885703
R17734 OUT_P.n1853 OUT_P.n1852 0.885703
R17735 OUT_P.n1863 OUT_P.n1862 0.885703
R17736 OUT_P.n1874 OUT_P.n1873 0.885703
R17737 OUT_P.n1885 OUT_P.n1884 0.885703
R17738 OUT_P.n1894 OUT_P.n1893 0.885703
R17739 OUT_P.n160 OUT_P.n159 0.835535
R17740 OUT_P.n1586 OUT_P.n1585 0.835535
R17741 OUT_P.n1297 OUT_P.n1296 0.824999
R17742 OUT_P.n1285 OUT_P.n1284 0.824999
R17743 OUT_P.n1273 OUT_P.n1272 0.824999
R17744 OUT_P.n1261 OUT_P.n1260 0.824999
R17745 OUT_P.n1249 OUT_P.n1248 0.824999
R17746 OUT_P.n1237 OUT_P.n1236 0.824999
R17747 OUT_P.n1225 OUT_P.n1224 0.824999
R17748 OUT_P.n1213 OUT_P.n1212 0.824999
R17749 OUT_P.n1201 OUT_P.n1200 0.824999
R17750 OUT_P.n1189 OUT_P.n1188 0.824999
R17751 OUT_P.n1177 OUT_P.n1176 0.824999
R17752 OUT_P.n1165 OUT_P.n1164 0.824999
R17753 OUT_P.n1153 OUT_P.n1152 0.824999
R17754 OUT_P.n1141 OUT_P.n1140 0.824999
R17755 OUT_P.n1291 OUT_P.n1290 0.824997
R17756 OUT_P.n204 OUT_P.n203 0.824997
R17757 OUT_P.n216 OUT_P.n215 0.824997
R17758 OUT_P.n227 OUT_P.n226 0.824997
R17759 OUT_P.n238 OUT_P.n237 0.824997
R17760 OUT_P.n264 OUT_P.n263 0.824997
R17761 OUT_P.n275 OUT_P.n274 0.824997
R17762 OUT_P.n286 OUT_P.n285 0.824997
R17763 OUT_P.n297 OUT_P.n296 0.824997
R17764 OUT_P.n308 OUT_P.n307 0.824997
R17765 OUT_P.n319 OUT_P.n318 0.824997
R17766 OUT_P.n330 OUT_P.n329 0.824997
R17767 OUT_P.n341 OUT_P.n340 0.824997
R17768 OUT_P.n361 OUT_P.n360 0.824997
R17769 OUT_P.n372 OUT_P.n371 0.824997
R17770 OUT_P.n383 OUT_P.n382 0.824997
R17771 OUT_P.n394 OUT_P.n393 0.824997
R17772 OUT_P.n405 OUT_P.n404 0.824997
R17773 OUT_P.n416 OUT_P.n415 0.824997
R17774 OUT_P.n427 OUT_P.n426 0.824997
R17775 OUT_P.n438 OUT_P.n437 0.824997
R17776 OUT_P.n453 OUT_P.n452 0.824997
R17777 OUT_P.n464 OUT_P.n463 0.824997
R17778 OUT_P.n475 OUT_P.n474 0.824997
R17779 OUT_P.n486 OUT_P.n485 0.824997
R17780 OUT_P.n497 OUT_P.n496 0.824997
R17781 OUT_P.n508 OUT_P.n507 0.824997
R17782 OUT_P.n519 OUT_P.n518 0.824997
R17783 OUT_P.n530 OUT_P.n529 0.824997
R17784 OUT_P.n1279 OUT_P.n1278 0.824997
R17785 OUT_P.n1267 OUT_P.n1266 0.824997
R17786 OUT_P.n1255 OUT_P.n1254 0.824997
R17787 OUT_P.n1243 OUT_P.n1242 0.824997
R17788 OUT_P.n1231 OUT_P.n1230 0.824997
R17789 OUT_P.n1219 OUT_P.n1218 0.824997
R17790 OUT_P.n1207 OUT_P.n1206 0.824997
R17791 OUT_P.n1195 OUT_P.n1194 0.824997
R17792 OUT_P.n1183 OUT_P.n1182 0.824997
R17793 OUT_P.n1171 OUT_P.n1170 0.824997
R17794 OUT_P.n1159 OUT_P.n1158 0.824997
R17795 OUT_P.n1147 OUT_P.n1146 0.824997
R17796 OUT_P.n1135 OUT_P.n1134 0.824997
R17797 OUT_P.n1700 OUT_P.n1699 0.82495
R17798 OUT_P.n1694 OUT_P.n1693 0.82495
R17799 OUT_P.n1679 OUT_P.n1678 0.82495
R17800 OUT_P.n1673 OUT_P.n1672 0.82495
R17801 OUT_P.n1658 OUT_P.n1657 0.82495
R17802 OUT_P.n1652 OUT_P.n1651 0.82495
R17803 OUT_P.n1637 OUT_P.n1636 0.82495
R17804 OUT_P.n1631 OUT_P.n1630 0.82495
R17805 OUT_P.n1616 OUT_P.n1615 0.82495
R17806 OUT_P.n1610 OUT_P.n1609 0.82495
R17807 OUT_P.n1882 OUT_P.n1881 0.82495
R17808 OUT_P.n1871 OUT_P.n1870 0.82495
R17809 OUT_P.n1841 OUT_P.n1840 0.82495
R17810 OUT_P.n1830 OUT_P.n1829 0.82495
R17811 OUT_P.n707 OUT_P.n706 0.82495
R17812 OUT_P.n701 OUT_P.n700 0.82495
R17813 OUT_P.n686 OUT_P.n685 0.82495
R17814 OUT_P.n680 OUT_P.n679 0.82495
R17815 OUT_P.n665 OUT_P.n664 0.82495
R17816 OUT_P.n659 OUT_P.n658 0.82495
R17817 OUT_P.n644 OUT_P.n643 0.82495
R17818 OUT_P.n638 OUT_P.n637 0.82495
R17819 OUT_P.n623 OUT_P.n622 0.82495
R17820 OUT_P.n617 OUT_P.n616 0.82495
R17821 OUT_P.n602 OUT_P.n601 0.82495
R17822 OUT_P.n596 OUT_P.n595 0.82495
R17823 OUT_P.n581 OUT_P.n580 0.82495
R17824 OUT_P.n575 OUT_P.n574 0.82495
R17825 OUT_P.n1068 OUT_P.n1067 0.736598
R17826 OUT_P.n11 OUT_P.n9 0.727916
R17827 OUT_P.n21 OUT_P.n20 0.727916
R17828 OUT_P.n31 OUT_P.n30 0.727916
R17829 OUT_P.n136 OUT_P.n135 0.727916
R17830 OUT_P.n147 OUT_P.n146 0.727916
R17831 OUT_P.n157 OUT_P.n156 0.727916
R17832 OUT_P.n166 OUT_P.n165 0.727916
R17833 OUT_P.n177 OUT_P.n176 0.727916
R17834 OUT_P.n187 OUT_P.n186 0.727916
R17835 OUT_P.n1537 OUT_P.n1524 0.727104
R17836 OUT_P.n1556 OUT_P.n1554 0.727104
R17837 OUT_P.n975 OUT_P.n932 0.727104
R17838 OUT_P.n1000 OUT_P.n919 0.727104
R17839 OUT_P.n967 OUT_P.n947 0.727104
R17840 OUT_P.n720 OUT_P.n709 0.727104
R17841 OUT_P.n729 OUT_P.n697 0.727104
R17842 OUT_P.n742 OUT_P.n688 0.727104
R17843 OUT_P.n751 OUT_P.n676 0.727104
R17844 OUT_P.n760 OUT_P.n667 0.727104
R17845 OUT_P.n769 OUT_P.n655 0.727104
R17846 OUT_P.n798 OUT_P.n646 0.727104
R17847 OUT_P.n807 OUT_P.n634 0.727104
R17848 OUT_P.n816 OUT_P.n625 0.727104
R17849 OUT_P.n825 OUT_P.n613 0.727104
R17850 OUT_P.n853 OUT_P.n604 0.727104
R17851 OUT_P.n862 OUT_P.n592 0.727104
R17852 OUT_P.n871 OUT_P.n583 0.727104
R17853 OUT_P.n880 OUT_P.n571 0.727104
R17854 OUT_P.n56 OUT_P.n44 0.727104
R17855 OUT_P.n1510 OUT_P.n1490 0.727104
R17856 OUT_P.n1597 OUT_P.n1460 0.727104
R17857 OUT_P.n1588 OUT_P.n1470 0.727104
R17858 OUT_P.n1579 OUT_P.n1481 0.727104
R17859 OUT_P.n1709 OUT_P.n1707 0.727104
R17860 OUT_P.n1718 OUT_P.n1696 0.727104
R17861 OUT_P.n1737 OUT_P.n1686 0.727104
R17862 OUT_P.n1746 OUT_P.n1675 0.727104
R17863 OUT_P.n1755 OUT_P.n1665 0.727104
R17864 OUT_P.n1764 OUT_P.n1654 0.727104
R17865 OUT_P.n1777 OUT_P.n1644 0.727104
R17866 OUT_P.n1786 OUT_P.n1633 0.727104
R17867 OUT_P.n1795 OUT_P.n1623 0.727104
R17868 OUT_P.n1804 OUT_P.n1612 0.727104
R17869 OUT_P.n1126 OUT_P.n1113 0.727104
R17870 OUT_P.n1301 OUT_P.n1299 0.727104
R17871 OUT_P.n1310 OUT_P.n1287 0.727104
R17872 OUT_P.n1328 OUT_P.n1275 0.727104
R17873 OUT_P.n1337 OUT_P.n1263 0.727104
R17874 OUT_P.n1346 OUT_P.n1251 0.727104
R17875 OUT_P.n1355 OUT_P.n1239 0.727104
R17876 OUT_P.n1369 OUT_P.n1227 0.727104
R17877 OUT_P.n1378 OUT_P.n1215 0.727104
R17878 OUT_P.n1387 OUT_P.n1203 0.727104
R17879 OUT_P.n1396 OUT_P.n1191 0.727104
R17880 OUT_P.n1410 OUT_P.n1179 0.727104
R17881 OUT_P.n1419 OUT_P.n1167 0.727104
R17882 OUT_P.n1428 OUT_P.n1155 0.727104
R17883 OUT_P.n1437 OUT_P.n1143 0.727104
R17884 OUT_P.n110 OUT_P.n101 0.726858
R17885 OUT_P.n1005 OUT_P.n911 0.726858
R17886 OUT_P.n1952 OUT_P.n1951 0.706873
R17887 OUT_P.n303 OUT_P.n302 0.685007
R17888 OUT_P.n400 OUT_P.n399 0.685007
R17889 OUT_P.n492 OUT_P.n491 0.685007
R17890 OUT_P.n1344 OUT_P.n1343 0.685007
R17891 OUT_P.n1385 OUT_P.n1384 0.685007
R17892 OUT_P.n1426 OUT_P.n1425 0.685007
R17893 OUT_P.n1949 OUT_P.n1948 0.673915
R17894 OUT_P.n1563 OUT_P.n1562 0.673915
R17895 OUT_P.n1540 OUT_P.n1539 0.673915
R17896 OUT_P.n97 OUT_P.n96 0.673915
R17897 OUT_P.n113 OUT_P.n112 0.673915
R17898 OUT_P.n567 OUT_P.n566 0.673915
R17899 OUT_P.n1008 OUT_P.n1007 0.673915
R17900 OUT_P.n973 OUT_P.n972 0.673915
R17901 OUT_P.n970 OUT_P.n969 0.673915
R17902 OUT_P.n60 OUT_P.n58 0.673915
R17903 OUT_P.n83 OUT_P.n82 0.673915
R17904 OUT_P.n1129 OUT_P.n1128 0.673915
R17905 OUT_P.n996 OUT_P.n995 0.617177
R17906 OUT_P.n1306 OUT_P.n1293 0.616779
R17907 OUT_P.n1121 OUT_P.n1119 0.616779
R17908 OUT_P.n1714 OUT_P.n1702 0.616779
R17909 OUT_P.n1723 OUT_P.n1690 0.616779
R17910 OUT_P.n1742 OUT_P.n1681 0.616779
R17911 OUT_P.n1751 OUT_P.n1669 0.616779
R17912 OUT_P.n1760 OUT_P.n1660 0.616779
R17913 OUT_P.n1769 OUT_P.n1648 0.616779
R17914 OUT_P.n1782 OUT_P.n1639 0.616779
R17915 OUT_P.n1791 OUT_P.n1627 0.616779
R17916 OUT_P.n1800 OUT_P.n1618 0.616779
R17917 OUT_P.n1809 OUT_P.n1606 0.616779
R17918 OUT_P.n1592 OUT_P.n1466 0.616779
R17919 OUT_P.n1583 OUT_P.n1475 0.616779
R17920 OUT_P.n1505 OUT_P.n1496 0.616779
R17921 OUT_P.n1574 OUT_P.n1485 0.616779
R17922 OUT_P.n1532 OUT_P.n1530 0.616779
R17923 OUT_P.n1561 OUT_P.n1548 0.616779
R17924 OUT_P.n716 OUT_P.n714 0.616779
R17925 OUT_P.n725 OUT_P.n703 0.616779
R17926 OUT_P.n738 OUT_P.n693 0.616779
R17927 OUT_P.n747 OUT_P.n682 0.616779
R17928 OUT_P.n756 OUT_P.n672 0.616779
R17929 OUT_P.n765 OUT_P.n661 0.616779
R17930 OUT_P.n794 OUT_P.n651 0.616779
R17931 OUT_P.n803 OUT_P.n640 0.616779
R17932 OUT_P.n812 OUT_P.n630 0.616779
R17933 OUT_P.n821 OUT_P.n619 0.616779
R17934 OUT_P.n849 OUT_P.n609 0.616779
R17935 OUT_P.n858 OUT_P.n598 0.616779
R17936 OUT_P.n867 OUT_P.n588 0.616779
R17937 OUT_P.n876 OUT_P.n577 0.616779
R17938 OUT_P.n95 OUT_P.n88 0.616779
R17939 OUT_P.n52 OUT_P.n50 0.616779
R17940 OUT_P.n80 OUT_P.n68 0.616779
R17941 OUT_P.n1315 OUT_P.n1281 0.616779
R17942 OUT_P.n1333 OUT_P.n1269 0.616779
R17943 OUT_P.n1342 OUT_P.n1257 0.616779
R17944 OUT_P.n1351 OUT_P.n1245 0.616779
R17945 OUT_P.n1360 OUT_P.n1233 0.616779
R17946 OUT_P.n1374 OUT_P.n1221 0.616779
R17947 OUT_P.n1383 OUT_P.n1209 0.616779
R17948 OUT_P.n1392 OUT_P.n1197 0.616779
R17949 OUT_P.n1401 OUT_P.n1185 0.616779
R17950 OUT_P.n1415 OUT_P.n1173 0.616779
R17951 OUT_P.n1424 OUT_P.n1161 0.616779
R17952 OUT_P.n1433 OUT_P.n1149 0.616779
R17953 OUT_P.n1442 OUT_P.n1137 0.616779
R17954 OUT_P.n1296 OUT_P.t112 0.607167
R17955 OUT_P.n1296 OUT_P.n1295 0.607167
R17956 OUT_P.n1290 OUT_P.t48 0.607167
R17957 OUT_P.n1290 OUT_P.n1289 0.607167
R17958 OUT_P.n1284 OUT_P.t145 0.607167
R17959 OUT_P.n1284 OUT_P.n1283 0.607167
R17960 OUT_P.n1699 OUT_P.t209 0.607167
R17961 OUT_P.n1699 OUT_P.n1698 0.607167
R17962 OUT_P.n1693 OUT_P.t36 0.607167
R17963 OUT_P.n1693 OUT_P.n1692 0.607167
R17964 OUT_P.n1678 OUT_P.t115 0.607167
R17965 OUT_P.n1678 OUT_P.n1677 0.607167
R17966 OUT_P.n1672 OUT_P.t62 0.607167
R17967 OUT_P.n1672 OUT_P.n1671 0.607167
R17968 OUT_P.n1657 OUT_P.t153 0.607167
R17969 OUT_P.n1657 OUT_P.n1656 0.607167
R17970 OUT_P.n1651 OUT_P.t114 0.607167
R17971 OUT_P.n1651 OUT_P.n1650 0.607167
R17972 OUT_P.n1636 OUT_P.t54 0.607167
R17973 OUT_P.n1636 OUT_P.n1635 0.607167
R17974 OUT_P.n1630 OUT_P.t215 0.607167
R17975 OUT_P.n1630 OUT_P.n1629 0.607167
R17976 OUT_P.n1615 OUT_P.t45 0.607167
R17977 OUT_P.n1615 OUT_P.n1614 0.607167
R17978 OUT_P.n1609 OUT_P.t205 0.607167
R17979 OUT_P.n1609 OUT_P.n1608 0.607167
R17980 OUT_P.n1881 OUT_P.t150 0.607167
R17981 OUT_P.n1881 OUT_P.n1880 0.607167
R17982 OUT_P.n1870 OUT_P.t195 0.607167
R17983 OUT_P.n1870 OUT_P.n1869 0.607167
R17984 OUT_P.n1840 OUT_P.t110 0.607167
R17985 OUT_P.n1840 OUT_P.n1839 0.607167
R17986 OUT_P.n1829 OUT_P.t85 0.607167
R17987 OUT_P.n1829 OUT_P.n1828 0.607167
R17988 OUT_P.n203 OUT_P.t230 0.607167
R17989 OUT_P.n203 OUT_P.n202 0.607167
R17990 OUT_P.n215 OUT_P.t119 0.607167
R17991 OUT_P.n215 OUT_P.n214 0.607167
R17992 OUT_P.n226 OUT_P.t183 0.607167
R17993 OUT_P.n226 OUT_P.n225 0.607167
R17994 OUT_P.n237 OUT_P.t124 0.607167
R17995 OUT_P.n237 OUT_P.n236 0.607167
R17996 OUT_P.n263 OUT_P.t130 0.607167
R17997 OUT_P.n263 OUT_P.n262 0.607167
R17998 OUT_P.n274 OUT_P.t199 0.607167
R17999 OUT_P.n274 OUT_P.n273 0.607167
R18000 OUT_P.n285 OUT_P.t87 0.607167
R18001 OUT_P.n285 OUT_P.n284 0.607167
R18002 OUT_P.n296 OUT_P.t221 0.607167
R18003 OUT_P.n296 OUT_P.n295 0.607167
R18004 OUT_P.n307 OUT_P.t173 0.607167
R18005 OUT_P.n307 OUT_P.n306 0.607167
R18006 OUT_P.n318 OUT_P.t59 0.607167
R18007 OUT_P.n318 OUT_P.n317 0.607167
R18008 OUT_P.n329 OUT_P.t129 0.607167
R18009 OUT_P.n329 OUT_P.n328 0.607167
R18010 OUT_P.n340 OUT_P.t66 0.607167
R18011 OUT_P.n340 OUT_P.n339 0.607167
R18012 OUT_P.n360 OUT_P.t211 0.607167
R18013 OUT_P.n360 OUT_P.n359 0.607167
R18014 OUT_P.n371 OUT_P.t140 0.607167
R18015 OUT_P.n371 OUT_P.n370 0.607167
R18016 OUT_P.n382 OUT_P.t37 0.607167
R18017 OUT_P.n382 OUT_P.n381 0.607167
R18018 OUT_P.n393 OUT_P.t103 0.607167
R18019 OUT_P.n393 OUT_P.n392 0.607167
R18020 OUT_P.n404 OUT_P.t69 0.607167
R18021 OUT_P.n404 OUT_P.n403 0.607167
R18022 OUT_P.n415 OUT_P.t134 0.607167
R18023 OUT_P.n415 OUT_P.n414 0.607167
R18024 OUT_P.n426 OUT_P.t223 0.607167
R18025 OUT_P.n426 OUT_P.n425 0.607167
R18026 OUT_P.n437 OUT_P.t95 0.607167
R18027 OUT_P.n437 OUT_P.n436 0.607167
R18028 OUT_P.n452 OUT_P.t105 0.607167
R18029 OUT_P.n452 OUT_P.n451 0.607167
R18030 OUT_P.n463 OUT_P.t43 0.607167
R18031 OUT_P.n463 OUT_P.n462 0.607167
R18032 OUT_P.n474 OUT_P.t113 0.607167
R18033 OUT_P.n474 OUT_P.n473 0.607167
R18034 OUT_P.n485 OUT_P.t196 0.607167
R18035 OUT_P.n485 OUT_P.n484 0.607167
R18036 OUT_P.n496 OUT_P.t147 0.607167
R18037 OUT_P.n496 OUT_P.n495 0.607167
R18038 OUT_P.n507 OUT_P.t86 0.607167
R18039 OUT_P.n507 OUT_P.n506 0.607167
R18040 OUT_P.n518 OUT_P.t169 0.607167
R18041 OUT_P.n518 OUT_P.n517 0.607167
R18042 OUT_P.n529 OUT_P.t42 0.607167
R18043 OUT_P.n529 OUT_P.n528 0.607167
R18044 OUT_P.n706 OUT_P.t51 0.607167
R18045 OUT_P.n706 OUT_P.n705 0.607167
R18046 OUT_P.n700 OUT_P.t77 0.607167
R18047 OUT_P.n700 OUT_P.n699 0.607167
R18048 OUT_P.n685 OUT_P.t74 0.607167
R18049 OUT_P.n685 OUT_P.n684 0.607167
R18050 OUT_P.n679 OUT_P.t148 0.607167
R18051 OUT_P.n679 OUT_P.n678 0.607167
R18052 OUT_P.n664 OUT_P.t71 0.607167
R18053 OUT_P.n664 OUT_P.n663 0.607167
R18054 OUT_P.n658 OUT_P.t144 0.607167
R18055 OUT_P.n658 OUT_P.n657 0.607167
R18056 OUT_P.n643 OUT_P.t94 0.607167
R18057 OUT_P.n643 OUT_P.n642 0.607167
R18058 OUT_P.n637 OUT_P.t167 0.607167
R18059 OUT_P.n637 OUT_P.n636 0.607167
R18060 OUT_P.n622 OUT_P.t102 0.607167
R18061 OUT_P.n622 OUT_P.n621 0.607167
R18062 OUT_P.n616 OUT_P.t171 0.607167
R18063 OUT_P.n616 OUT_P.n615 0.607167
R18064 OUT_P.n601 OUT_P.t168 0.607167
R18065 OUT_P.n601 OUT_P.n600 0.607167
R18066 OUT_P.n595 OUT_P.t193 0.607167
R18067 OUT_P.n595 OUT_P.n594 0.607167
R18068 OUT_P.n580 OUT_P.t121 0.607167
R18069 OUT_P.n580 OUT_P.n579 0.607167
R18070 OUT_P.n574 OUT_P.t192 0.607167
R18071 OUT_P.n574 OUT_P.n573 0.607167
R18072 OUT_P.n1278 OUT_P.t220 0.607167
R18073 OUT_P.n1278 OUT_P.n1277 0.607167
R18074 OUT_P.n1272 OUT_P.t39 0.607167
R18075 OUT_P.n1272 OUT_P.n1271 0.607167
R18076 OUT_P.n1266 OUT_P.t131 0.607167
R18077 OUT_P.n1266 OUT_P.n1265 0.607167
R18078 OUT_P.n1260 OUT_P.t73 0.607167
R18079 OUT_P.n1260 OUT_P.n1259 0.607167
R18080 OUT_P.n1254 OUT_P.t143 0.607167
R18081 OUT_P.n1254 OUT_P.n1253 0.607167
R18082 OUT_P.n1248 OUT_P.t44 0.607167
R18083 OUT_P.n1248 OUT_P.n1247 0.607167
R18084 OUT_P.n1242 OUT_P.t186 0.607167
R18085 OUT_P.n1242 OUT_P.n1241 0.607167
R18086 OUT_P.n1236 OUT_P.t81 0.607167
R18087 OUT_P.n1236 OUT_P.n1235 0.607167
R18088 OUT_P.n1230 OUT_P.t154 0.607167
R18089 OUT_P.n1230 OUT_P.n1229 0.607167
R18090 OUT_P.n1224 OUT_P.t191 0.607167
R18091 OUT_P.n1224 OUT_P.n1223 0.607167
R18092 OUT_P.n1218 OUT_P.t61 0.607167
R18093 OUT_P.n1218 OUT_P.n1217 0.607167
R18094 OUT_P.n1212 OUT_P.t208 0.607167
R18095 OUT_P.n1212 OUT_P.n1211 0.607167
R18096 OUT_P.n1206 OUT_P.t107 0.607167
R18097 OUT_P.n1206 OUT_P.n1205 0.607167
R18098 OUT_P.n1200 OUT_P.t228 0.607167
R18099 OUT_P.n1200 OUT_P.n1199 0.607167
R18100 OUT_P.n1194 OUT_P.t128 0.607167
R18101 OUT_P.n1194 OUT_P.n1193 0.607167
R18102 OUT_P.n1188 OUT_P.t64 0.607167
R18103 OUT_P.n1188 OUT_P.n1187 0.607167
R18104 OUT_P.n1182 OUT_P.t162 0.607167
R18105 OUT_P.n1182 OUT_P.n1181 0.607167
R18106 OUT_P.n1176 OUT_P.t175 0.607167
R18107 OUT_P.n1176 OUT_P.n1175 0.607167
R18108 OUT_P.n1170 OUT_P.t49 0.607167
R18109 OUT_P.n1170 OUT_P.n1169 0.607167
R18110 OUT_P.n1164 OUT_P.t146 0.607167
R18111 OUT_P.n1164 OUT_P.n1163 0.607167
R18112 OUT_P.n1158 OUT_P.t90 0.607167
R18113 OUT_P.n1158 OUT_P.n1157 0.607167
R18114 OUT_P.n1152 OUT_P.t187 0.607167
R18115 OUT_P.n1152 OUT_P.n1151 0.607167
R18116 OUT_P.n1146 OUT_P.t58 0.607167
R18117 OUT_P.n1146 OUT_P.n1145 0.607167
R18118 OUT_P.n1140 OUT_P.t201 0.607167
R18119 OUT_P.n1140 OUT_P.n1139 0.607167
R18120 OUT_P.n1134 OUT_P.t99 0.607167
R18121 OUT_P.n1134 OUT_P.n1133 0.607167
R18122 OUT_P.n190 OUT_P.n189 0.572507
R18123 OUT_P.n130 OUT_P.n129 0.572507
R18124 OUT_P.n34 OUT_P.n33 0.572507
R18125 OUT_P.n1600 OUT_P.n1599 0.572507
R18126 OUT_P.n1573 OUT_P.n1572 0.572507
R18127 OUT_P.n1513 OUT_P.n1512 0.572507
R18128 OUT_P.n347 OUT_P.n346 0.555711
R18129 OUT_P.n1362 OUT_P.n1361 0.555711
R18130 OUT_P.n1444 OUT_P.n1443 0.552542
R18131 OUT_P.n536 OUT_P.n535 0.548033
R18132 OUT_P.n1930 OUT_P.t245 0.5465
R18133 OUT_P.n1930 OUT_P.n1929 0.5465
R18134 OUT_P.n1935 OUT_P.t29 0.5465
R18135 OUT_P.n1935 OUT_P.n1934 0.5465
R18136 OUT_P.n1116 OUT_P.t31 0.5465
R18137 OUT_P.n1116 OUT_P.n1115 0.5465
R18138 OUT_P.n1110 OUT_P.t249 0.5465
R18139 OUT_P.n1110 OUT_P.n1109 0.5465
R18140 OUT_P.n1463 OUT_P.t268 0.5465
R18141 OUT_P.n1463 OUT_P.n1462 0.5465
R18142 OUT_P.n1478 OUT_P.t3 0.5465
R18143 OUT_P.n1478 OUT_P.n1477 0.5465
R18144 OUT_P.n1493 OUT_P.t34 0.5465
R18145 OUT_P.n1493 OUT_P.n1492 0.5465
R18146 OUT_P.n1551 OUT_P.t16 0.5465
R18147 OUT_P.n1551 OUT_P.n1550 0.5465
R18148 OUT_P.n1527 OUT_P.t33 0.5465
R18149 OUT_P.n1527 OUT_P.n1526 0.5465
R18150 OUT_P.n1521 OUT_P.t26 0.5465
R18151 OUT_P.n1521 OUT_P.n1520 0.5465
R18152 OUT_P.n1545 OUT_P.t239 0.5465
R18153 OUT_P.n1545 OUT_P.n1544 0.5465
R18154 OUT_P.n16 OUT_P.t27 0.5465
R18155 OUT_P.n16 OUT_P.n15 0.5465
R18156 OUT_P.n142 OUT_P.t265 0.5465
R18157 OUT_P.n142 OUT_P.n141 0.5465
R18158 OUT_P.n172 OUT_P.t32 0.5465
R18159 OUT_P.n172 OUT_P.n171 0.5465
R18160 OUT_P.n985 OUT_P.t267 0.5465
R18161 OUT_P.n985 OUT_P.n984 0.5465
R18162 OUT_P.n951 OUT_P.t24 0.5465
R18163 OUT_P.n951 OUT_P.n950 0.5465
R18164 OUT_P.n957 OUT_P.t248 0.5465
R18165 OUT_P.n957 OUT_P.n956 0.5465
R18166 OUT_P.n927 OUT_P.t246 0.5465
R18167 OUT_P.n927 OUT_P.n926 0.5465
R18168 OUT_P.n921 OUT_P.t10 0.5465
R18169 OUT_P.n921 OUT_P.n920 0.5465
R18170 OUT_P.n942 OUT_P.t238 0.5465
R18171 OUT_P.n942 OUT_P.n941 0.5465
R18172 OUT_P.n936 OUT_P.t1 0.5465
R18173 OUT_P.n936 OUT_P.n935 0.5465
R18174 OUT_P.n981 OUT_P.t240 0.5465
R18175 OUT_P.n981 OUT_P.n980 0.5465
R18176 OUT_P.n560 OUT_P.t233 0.5465
R18177 OUT_P.n560 OUT_P.n559 0.5465
R18178 OUT_P.n546 OUT_P.t5 0.5465
R18179 OUT_P.n546 OUT_P.n545 0.5465
R18180 OUT_P.n913 OUT_P.t256 0.5465
R18181 OUT_P.n913 OUT_P.n912 0.5465
R18182 OUT_P.n905 OUT_P.t17 0.5465
R18183 OUT_P.n905 OUT_P.n904 0.5465
R18184 OUT_P.n47 OUT_P.t9 0.5465
R18185 OUT_P.n47 OUT_P.n46 0.5465
R18186 OUT_P.n41 OUT_P.t7 0.5465
R18187 OUT_P.n41 OUT_P.n40 0.5465
R18188 OUT_P.n65 OUT_P.t4 0.5465
R18189 OUT_P.n65 OUT_P.n64 0.5465
R18190 OUT_P.n72 OUT_P.t22 0.5465
R18191 OUT_P.n72 OUT_P.n71 0.5465
R18192 OUT_P.n259 OUT_P.n258 0.543352
R18193 OUT_P.n1326 OUT_P.n1325 0.543352
R18194 OUT_P.n444 OUT_P.n443 0.542718
R18195 OUT_P.n1403 OUT_P.n1402 0.542718
R18196 OUT_P.n448 OUT_P.n447 0.529408
R18197 OUT_P.n1408 OUT_P.n1407 0.529408
R18198 OUT_P.n244 OUT_P.n243 0.528775
R18199 OUT_P.n1317 OUT_P.n1316 0.528775
R18200 OUT_P.n356 OUT_P.n355 0.516415
R18201 OUT_P.n1367 OUT_P.n1366 0.516415
R18202 OUT_P.n754 OUT_P.n753 0.482824
R18203 OUT_P.n810 OUT_P.n809 0.482824
R18204 OUT_P.n865 OUT_P.n864 0.482824
R18205 OUT_P.n1753 OUT_P.n1752 0.482824
R18206 OUT_P.n1793 OUT_P.n1792 0.482824
R18207 OUT_P.n1856 OUT_P.n1855 0.482824
R18208 OUT_P.n772 OUT_P.n771 0.453986
R18209 OUT_P.n1771 OUT_P.n1770 0.453986
R18210 OUT_P.n1023 OUT_P.n1022 0.4505
R18211 OUT_P.n1015 OUT_P.n1014 0.4505
R18212 OUT_P.n1069 OUT_P.n1068 0.4505
R18213 OUT_P.n1019 OUT_P.n1018 0.4505
R18214 OUT_P.n1897 OUT_P.n1896 0.447157
R18215 OUT_P.n883 OUT_P.n882 0.446728
R18216 OUT_P.n736 OUT_P.n735 0.441627
R18217 OUT_P.n1735 OUT_P.n1734 0.441627
R18218 OUT_P.n828 OUT_P.n827 0.440993
R18219 OUT_P.n1811 OUT_P.n1810 0.440993
R18220 OUT_P.n847 OUT_P.n846 0.427683
R18221 OUT_P.n1815 OUT_P.n1814 0.427683
R18222 OUT_P.n732 OUT_P.n731 0.427049
R18223 OUT_P.n1725 OUT_P.n1724 0.427049
R18224 OUT_P.n792 OUT_P.n791 0.41469
R18225 OUT_P.n1775 OUT_P.n1774 0.41469
R18226 OUT_P.n256 OUT_P.n255 0.395359
R18227 OUT_P.n723 OUT_P.n722 0.389021
R18228 OUT_P.n745 OUT_P.n744 0.389021
R18229 OUT_P.n763 OUT_P.n762 0.389021
R18230 OUT_P.n801 OUT_P.n800 0.389021
R18231 OUT_P.n819 OUT_P.n818 0.389021
R18232 OUT_P.n856 OUT_P.n855 0.389021
R18233 OUT_P.n874 OUT_P.n873 0.389021
R18234 OUT_P.n1716 OUT_P.n1715 0.389021
R18235 OUT_P.n1744 OUT_P.n1743 0.389021
R18236 OUT_P.n1762 OUT_P.n1761 0.389021
R18237 OUT_P.n1784 OUT_P.n1783 0.389021
R18238 OUT_P.n1802 OUT_P.n1801 0.389021
R18239 OUT_P.n1836 OUT_P.n1835 0.389021
R18240 OUT_P.n1877 OUT_P.n1876 0.389021
R18241 OUT_P.n127 OUT_P.n85 0.356063
R18242 OUT_P.n1922 OUT_P.n1921 0.356063
R18243 OUT_P.n1904 OUT_P.n1903 0.356063
R18244 OUT_P.n954 OUT_P.n953 0.336464
R18245 OUT_P.n991 OUT_P.n990 0.336464
R18246 OUT_P.n557 OUT_P.n556 0.336464
R18247 OUT_P.n840 OUT_P.n839 0.2705
R18248 OUT_P.n897 OUT_P.n896 0.2705
R18249 OUT_P.n786 OUT_P.n785 0.2705
R18250 OUT_P.n118 OUT_P.n117 0.231204
R18251 OUT_P.n1912 OUT_P.n1908 0.231204
R18252 OUT_P.n928 OUT_P.n925 0.191654
R18253 OUT_P.n943 OUT_P.n940 0.191654
R18254 OUT_P.n548 OUT_P.n547 0.191654
R18255 OUT_P.n1040 OUT_P.n1039 0.187374
R18256 OUT_P.n1944 OUT_P.n1943 0.186204
R18257 OUT_P.n1559 OUT_P.n1558 0.186204
R18258 OUT_P.n1535 OUT_P.n1534 0.186204
R18259 OUT_P.n93 OUT_P.n92 0.186204
R18260 OUT_P.n108 OUT_P.n107 0.186204
R18261 OUT_P.n554 OUT_P.n553 0.186204
R18262 OUT_P.n1003 OUT_P.n1002 0.186204
R18263 OUT_P.n978 OUT_P.n977 0.186204
R18264 OUT_P.n965 OUT_P.n964 0.186204
R18265 OUT_P.n718 OUT_P.n717 0.186204
R18266 OUT_P.n727 OUT_P.n726 0.186204
R18267 OUT_P.n740 OUT_P.n739 0.186204
R18268 OUT_P.n749 OUT_P.n748 0.186204
R18269 OUT_P.n758 OUT_P.n757 0.186204
R18270 OUT_P.n767 OUT_P.n766 0.186204
R18271 OUT_P.n796 OUT_P.n795 0.186204
R18272 OUT_P.n805 OUT_P.n804 0.186204
R18273 OUT_P.n814 OUT_P.n813 0.186204
R18274 OUT_P.n823 OUT_P.n822 0.186204
R18275 OUT_P.n851 OUT_P.n850 0.186204
R18276 OUT_P.n860 OUT_P.n859 0.186204
R18277 OUT_P.n869 OUT_P.n868 0.186204
R18278 OUT_P.n878 OUT_P.n877 0.186204
R18279 OUT_P.n211 OUT_P.n210 0.186204
R18280 OUT_P.n222 OUT_P.n221 0.186204
R18281 OUT_P.n233 OUT_P.n232 0.186204
R18282 OUT_P.n270 OUT_P.n269 0.186204
R18283 OUT_P.n281 OUT_P.n280 0.186204
R18284 OUT_P.n292 OUT_P.n291 0.186204
R18285 OUT_P.n314 OUT_P.n313 0.186204
R18286 OUT_P.n325 OUT_P.n324 0.186204
R18287 OUT_P.n336 OUT_P.n335 0.186204
R18288 OUT_P.n367 OUT_P.n366 0.186204
R18289 OUT_P.n378 OUT_P.n377 0.186204
R18290 OUT_P.n389 OUT_P.n388 0.186204
R18291 OUT_P.n411 OUT_P.n410 0.186204
R18292 OUT_P.n422 OUT_P.n421 0.186204
R18293 OUT_P.n433 OUT_P.n432 0.186204
R18294 OUT_P.n459 OUT_P.n458 0.186204
R18295 OUT_P.n470 OUT_P.n469 0.186204
R18296 OUT_P.n481 OUT_P.n480 0.186204
R18297 OUT_P.n503 OUT_P.n502 0.186204
R18298 OUT_P.n514 OUT_P.n513 0.186204
R18299 OUT_P.n525 OUT_P.n524 0.186204
R18300 OUT_P.n180 OUT_P.n179 0.186204
R18301 OUT_P.n169 OUT_P.n168 0.186204
R18302 OUT_P.n150 OUT_P.n149 0.186204
R18303 OUT_P.n139 OUT_P.n138 0.186204
R18304 OUT_P.n24 OUT_P.n23 0.186204
R18305 OUT_P.n13 OUT_P.n12 0.186204
R18306 OUT_P.n54 OUT_P.n53 0.186204
R18307 OUT_P.n79 OUT_P.n78 0.186204
R18308 OUT_P.n1595 OUT_P.n1594 0.186204
R18309 OUT_P.n1591 OUT_P.n1590 0.186204
R18310 OUT_P.n1582 OUT_P.n1581 0.186204
R18311 OUT_P.n1577 OUT_P.n1576 0.186204
R18312 OUT_P.n1508 OUT_P.n1507 0.186204
R18313 OUT_P.n1504 OUT_P.n1503 0.186204
R18314 OUT_P.n1712 OUT_P.n1711 0.186204
R18315 OUT_P.n1721 OUT_P.n1720 0.186204
R18316 OUT_P.n1740 OUT_P.n1739 0.186204
R18317 OUT_P.n1749 OUT_P.n1748 0.186204
R18318 OUT_P.n1758 OUT_P.n1757 0.186204
R18319 OUT_P.n1767 OUT_P.n1766 0.186204
R18320 OUT_P.n1780 OUT_P.n1779 0.186204
R18321 OUT_P.n1789 OUT_P.n1788 0.186204
R18322 OUT_P.n1798 OUT_P.n1797 0.186204
R18323 OUT_P.n1807 OUT_P.n1806 0.186204
R18324 OUT_P.n1825 OUT_P.n1824 0.186204
R18325 OUT_P.n1847 OUT_P.n1846 0.186204
R18326 OUT_P.n1866 OUT_P.n1865 0.186204
R18327 OUT_P.n1888 OUT_P.n1887 0.186204
R18328 OUT_P.n1304 OUT_P.n1303 0.186204
R18329 OUT_P.n1308 OUT_P.n1307 0.186204
R18330 OUT_P.n1313 OUT_P.n1312 0.186204
R18331 OUT_P.n1331 OUT_P.n1330 0.186204
R18332 OUT_P.n1335 OUT_P.n1334 0.186204
R18333 OUT_P.n1340 OUT_P.n1339 0.186204
R18334 OUT_P.n1349 OUT_P.n1348 0.186204
R18335 OUT_P.n1353 OUT_P.n1352 0.186204
R18336 OUT_P.n1358 OUT_P.n1357 0.186204
R18337 OUT_P.n1372 OUT_P.n1371 0.186204
R18338 OUT_P.n1376 OUT_P.n1375 0.186204
R18339 OUT_P.n1381 OUT_P.n1380 0.186204
R18340 OUT_P.n1390 OUT_P.n1389 0.186204
R18341 OUT_P.n1394 OUT_P.n1393 0.186204
R18342 OUT_P.n1399 OUT_P.n1398 0.186204
R18343 OUT_P.n1413 OUT_P.n1412 0.186204
R18344 OUT_P.n1417 OUT_P.n1416 0.186204
R18345 OUT_P.n1422 OUT_P.n1421 0.186204
R18346 OUT_P.n1431 OUT_P.n1430 0.186204
R18347 OUT_P.n1435 OUT_P.n1434 0.186204
R18348 OUT_P.n1440 OUT_P.n1439 0.186204
R18349 OUT_P.n1124 OUT_P.n1123 0.186204
R18350 OUT_P.n1070 OUT_P.n1069 0.180553
R18351 OUT_P.n1063 OUT_P.n1038 0.180553
R18352 OUT_P.n1094 OUT_P.n1026 0.180553
R18353 OUT_P.n835 OUT_P.n834 0.145641
R18354 OUT_P.n892 OUT_P.n891 0.145641
R18355 OUT_P.n781 OUT_P.n780 0.145641
R18356 OUT_P.n959 OUT_P.n958 0.109963
R18357 OUT_P.n925 OUT_P.n924 0.106363
R18358 OUT_P.n940 OUT_P.n939 0.106363
R18359 OUT_P.n549 OUT_P.n548 0.106363
R18360 OUT_P.n123 OUT_P.n122 0.106345
R18361 OUT_P.n1566 OUT_P.n1565 0.106345
R18362 OUT_P.n1917 OUT_P.n1916 0.106345
R18363 OUT_P.n1452 OUT_P.n1451 0.106345
R18364 OUT_P.n1449 OUT_P.n1448 0.101908
R18365 OUT_P.n1933 OUT_P.n1928 0.0992756
R18366 OUT_P.n1893 OUT_P.n1890 0.0992756
R18367 OUT_P.n1884 OUT_P.n1879 0.0992756
R18368 OUT_P.n1873 OUT_P.n1868 0.0992756
R18369 OUT_P.n1862 OUT_P.n1858 0.0992756
R18370 OUT_P.n1852 OUT_P.n1849 0.0992756
R18371 OUT_P.n1843 OUT_P.n1838 0.0992756
R18372 OUT_P.n1832 OUT_P.n1827 0.0992756
R18373 OUT_P.n1821 OUT_P.n1817 0.0992756
R18374 OUT_P.n218 OUT_P.n213 0.0992756
R18375 OUT_P.n229 OUT_P.n224 0.0992756
R18376 OUT_P.n240 OUT_P.n235 0.0992756
R18377 OUT_P.n266 OUT_P.n261 0.0992756
R18378 OUT_P.n277 OUT_P.n272 0.0992756
R18379 OUT_P.n288 OUT_P.n283 0.0992756
R18380 OUT_P.n299 OUT_P.n294 0.0992756
R18381 OUT_P.n310 OUT_P.n305 0.0992756
R18382 OUT_P.n321 OUT_P.n316 0.0992756
R18383 OUT_P.n332 OUT_P.n327 0.0992756
R18384 OUT_P.n343 OUT_P.n338 0.0992756
R18385 OUT_P.n363 OUT_P.n358 0.0992756
R18386 OUT_P.n374 OUT_P.n369 0.0992756
R18387 OUT_P.n385 OUT_P.n380 0.0992756
R18388 OUT_P.n396 OUT_P.n391 0.0992756
R18389 OUT_P.n407 OUT_P.n402 0.0992756
R18390 OUT_P.n418 OUT_P.n413 0.0992756
R18391 OUT_P.n429 OUT_P.n424 0.0992756
R18392 OUT_P.n440 OUT_P.n435 0.0992756
R18393 OUT_P.n455 OUT_P.n450 0.0992756
R18394 OUT_P.n466 OUT_P.n461 0.0992756
R18395 OUT_P.n477 OUT_P.n472 0.0992756
R18396 OUT_P.n488 OUT_P.n483 0.0992756
R18397 OUT_P.n499 OUT_P.n494 0.0992756
R18398 OUT_P.n510 OUT_P.n505 0.0992756
R18399 OUT_P.n521 OUT_P.n516 0.0992756
R18400 OUT_P.n532 OUT_P.n527 0.0992756
R18401 OUT_P.n563 OUT_P.n558 0.0992756
R18402 OUT_P.n1901 OUT_P.n1900 0.0982485
R18403 OUT_P.n903 OUT_P.n902 0.0978197
R18404 OUT_P.n540 OUT_P.n539 0.0973992
R18405 OUT_P.n1091 OUT_P.n1090 0.0890366
R18406 OUT_P.n1060 OUT_P.n1059 0.0890366
R18407 OUT_P.n1500 OUT_P.n1499 0.0832399
R18408 OUT_P.n104 OUT_P.n103 0.0832399
R18409 OUT_P.n550 OUT_P.n544 0.0832399
R18410 OUT_P.n74 OUT_P.n70 0.0832399
R18411 OUT_P.n207 OUT_P.n206 0.0831446
R18412 OUT_P.n9 OUT_P.n8 0.0826464
R18413 OUT_P.n20 OUT_P.n19 0.0826464
R18414 OUT_P.n30 OUT_P.n29 0.0826464
R18415 OUT_P.n135 OUT_P.n134 0.0826464
R18416 OUT_P.n146 OUT_P.n145 0.0826464
R18417 OUT_P.n156 OUT_P.n155 0.0826464
R18418 OUT_P.n165 OUT_P.n164 0.0826464
R18419 OUT_P.n176 OUT_P.n175 0.0826464
R18420 OUT_P.n186 OUT_P.n185 0.0826464
R18421 OUT_P.n101 OUT_P.n99 0.0824117
R18422 OUT_P.n911 OUT_P.n907 0.0824117
R18423 OUT_P.n1299 OUT_P.n1294 0.0823987
R18424 OUT_P.n1287 OUT_P.n1282 0.0823987
R18425 OUT_P.n1113 OUT_P.n1108 0.0823987
R18426 OUT_P.n1707 OUT_P.n1703 0.0823987
R18427 OUT_P.n1696 OUT_P.n1691 0.0823987
R18428 OUT_P.n1686 OUT_P.n1682 0.0823987
R18429 OUT_P.n1675 OUT_P.n1670 0.0823987
R18430 OUT_P.n1665 OUT_P.n1661 0.0823987
R18431 OUT_P.n1654 OUT_P.n1649 0.0823987
R18432 OUT_P.n1644 OUT_P.n1640 0.0823987
R18433 OUT_P.n1633 OUT_P.n1628 0.0823987
R18434 OUT_P.n1623 OUT_P.n1619 0.0823987
R18435 OUT_P.n1612 OUT_P.n1607 0.0823987
R18436 OUT_P.n1460 OUT_P.n1456 0.0823987
R18437 OUT_P.n1470 OUT_P.n1467 0.0823987
R18438 OUT_P.n1481 OUT_P.n1476 0.0823987
R18439 OUT_P.n1490 OUT_P.n1486 0.0823987
R18440 OUT_P.n1554 OUT_P.n1549 0.0823987
R18441 OUT_P.n1524 OUT_P.n1519 0.0823987
R18442 OUT_P.n709 OUT_P.n704 0.0823987
R18443 OUT_P.n697 OUT_P.n694 0.0823987
R18444 OUT_P.n688 OUT_P.n683 0.0823987
R18445 OUT_P.n676 OUT_P.n673 0.0823987
R18446 OUT_P.n667 OUT_P.n662 0.0823987
R18447 OUT_P.n655 OUT_P.n652 0.0823987
R18448 OUT_P.n646 OUT_P.n641 0.0823987
R18449 OUT_P.n634 OUT_P.n631 0.0823987
R18450 OUT_P.n625 OUT_P.n620 0.0823987
R18451 OUT_P.n613 OUT_P.n610 0.0823987
R18452 OUT_P.n604 OUT_P.n599 0.0823987
R18453 OUT_P.n592 OUT_P.n589 0.0823987
R18454 OUT_P.n583 OUT_P.n578 0.0823987
R18455 OUT_P.n571 OUT_P.n568 0.0823987
R18456 OUT_P.n989 OUT_P.n988 0.0823987
R18457 OUT_P.n932 OUT_P.n923 0.0823987
R18458 OUT_P.n947 OUT_P.n938 0.0823987
R18459 OUT_P.n919 OUT_P.n915 0.0823987
R18460 OUT_P.n44 OUT_P.n39 0.0823987
R18461 OUT_P.n1275 OUT_P.n1270 0.0823987
R18462 OUT_P.n1263 OUT_P.n1258 0.0823987
R18463 OUT_P.n1251 OUT_P.n1246 0.0823987
R18464 OUT_P.n1239 OUT_P.n1234 0.0823987
R18465 OUT_P.n1227 OUT_P.n1222 0.0823987
R18466 OUT_P.n1215 OUT_P.n1210 0.0823987
R18467 OUT_P.n1203 OUT_P.n1198 0.0823987
R18468 OUT_P.n1191 OUT_P.n1186 0.0823987
R18469 OUT_P.n1179 OUT_P.n1174 0.0823987
R18470 OUT_P.n1167 OUT_P.n1162 0.0823987
R18471 OUT_P.n1155 OUT_P.n1150 0.0823987
R18472 OUT_P.n1143 OUT_P.n1138 0.0823987
R18473 OUT_P.n953 OUT_P.n952 0.0748144
R18474 OUT_P.n990 OUT_P.n986 0.0748144
R18475 OUT_P.n1548 OUT_P.n1543 0.0712285
R18476 OUT_P.n1530 OUT_P.n1525 0.0712285
R18477 OUT_P.n88 OUT_P.n86 0.0712285
R18478 OUT_P.n577 OUT_P.n572 0.0712285
R18479 OUT_P.n588 OUT_P.n584 0.0712285
R18480 OUT_P.n598 OUT_P.n593 0.0712285
R18481 OUT_P.n609 OUT_P.n605 0.0712285
R18482 OUT_P.n619 OUT_P.n614 0.0712285
R18483 OUT_P.n630 OUT_P.n626 0.0712285
R18484 OUT_P.n640 OUT_P.n635 0.0712285
R18485 OUT_P.n651 OUT_P.n647 0.0712285
R18486 OUT_P.n661 OUT_P.n656 0.0712285
R18487 OUT_P.n672 OUT_P.n668 0.0712285
R18488 OUT_P.n682 OUT_P.n677 0.0712285
R18489 OUT_P.n693 OUT_P.n689 0.0712285
R18490 OUT_P.n703 OUT_P.n698 0.0712285
R18491 OUT_P.n714 OUT_P.n710 0.0712285
R18492 OUT_P.n68 OUT_P.n63 0.0712285
R18493 OUT_P.n50 OUT_P.n45 0.0712285
R18494 OUT_P.n1485 OUT_P.n1482 0.0712285
R18495 OUT_P.n1496 OUT_P.n1491 0.0712285
R18496 OUT_P.n1475 OUT_P.n1471 0.0712285
R18497 OUT_P.n1466 OUT_P.n1461 0.0712285
R18498 OUT_P.n1606 OUT_P.n1603 0.0712285
R18499 OUT_P.n1618 OUT_P.n1613 0.0712285
R18500 OUT_P.n1627 OUT_P.n1624 0.0712285
R18501 OUT_P.n1639 OUT_P.n1634 0.0712285
R18502 OUT_P.n1648 OUT_P.n1645 0.0712285
R18503 OUT_P.n1660 OUT_P.n1655 0.0712285
R18504 OUT_P.n1669 OUT_P.n1666 0.0712285
R18505 OUT_P.n1681 OUT_P.n1676 0.0712285
R18506 OUT_P.n1690 OUT_P.n1687 0.0712285
R18507 OUT_P.n1702 OUT_P.n1697 0.0712285
R18508 OUT_P.n1137 OUT_P.n1132 0.0712285
R18509 OUT_P.n1149 OUT_P.n1144 0.0712285
R18510 OUT_P.n1161 OUT_P.n1156 0.0712285
R18511 OUT_P.n1173 OUT_P.n1168 0.0712285
R18512 OUT_P.n1185 OUT_P.n1180 0.0712285
R18513 OUT_P.n1197 OUT_P.n1192 0.0712285
R18514 OUT_P.n1209 OUT_P.n1204 0.0712285
R18515 OUT_P.n1221 OUT_P.n1216 0.0712285
R18516 OUT_P.n1233 OUT_P.n1228 0.0712285
R18517 OUT_P.n1245 OUT_P.n1240 0.0712285
R18518 OUT_P.n1257 OUT_P.n1252 0.0712285
R18519 OUT_P.n1269 OUT_P.n1264 0.0712285
R18520 OUT_P.n1281 OUT_P.n1276 0.0712285
R18521 OUT_P.n1119 OUT_P.n1114 0.0712285
R18522 OUT_P.n1293 OUT_P.n1288 0.0712285
R18523 OUT_P.n995 OUT_P.n994 0.0709833
R18524 OUT_P OUT_P.n1954 0.0683169
R18525 OUT_P.n1939 OUT_P.n1938 0.0623855
R18526 OUT_P.n1938 OUT_P.n1937 0.0623855
R18527 OUT_P.n960 OUT_P.n949 0.0623855
R18528 OUT_P.n949 OUT_P.n948 0.0623855
R18529 OUT_P.n995 OUT_P.n983 0.0536862
R18530 OUT_P.n1530 OUT_P.n1529 0.0534597
R18531 OUT_P.n1548 OUT_P.n1547 0.0534597
R18532 OUT_P.n88 OUT_P.n87 0.0534597
R18533 OUT_P.n714 OUT_P.n713 0.0534597
R18534 OUT_P.n703 OUT_P.n702 0.0534597
R18535 OUT_P.n693 OUT_P.n692 0.0534597
R18536 OUT_P.n682 OUT_P.n681 0.0534597
R18537 OUT_P.n672 OUT_P.n671 0.0534597
R18538 OUT_P.n661 OUT_P.n660 0.0534597
R18539 OUT_P.n651 OUT_P.n650 0.0534597
R18540 OUT_P.n640 OUT_P.n639 0.0534597
R18541 OUT_P.n630 OUT_P.n629 0.0534597
R18542 OUT_P.n619 OUT_P.n618 0.0534597
R18543 OUT_P.n609 OUT_P.n608 0.0534597
R18544 OUT_P.n598 OUT_P.n597 0.0534597
R18545 OUT_P.n588 OUT_P.n587 0.0534597
R18546 OUT_P.n577 OUT_P.n576 0.0534597
R18547 OUT_P.n50 OUT_P.n49 0.0534597
R18548 OUT_P.n68 OUT_P.n67 0.0534597
R18549 OUT_P.n1496 OUT_P.n1495 0.0534597
R18550 OUT_P.n1466 OUT_P.n1465 0.0534597
R18551 OUT_P.n1475 OUT_P.n1474 0.0534597
R18552 OUT_P.n1485 OUT_P.n1484 0.0534597
R18553 OUT_P.n1702 OUT_P.n1701 0.0534597
R18554 OUT_P.n1690 OUT_P.n1689 0.0534597
R18555 OUT_P.n1681 OUT_P.n1680 0.0534597
R18556 OUT_P.n1669 OUT_P.n1668 0.0534597
R18557 OUT_P.n1660 OUT_P.n1659 0.0534597
R18558 OUT_P.n1648 OUT_P.n1647 0.0534597
R18559 OUT_P.n1639 OUT_P.n1638 0.0534597
R18560 OUT_P.n1627 OUT_P.n1626 0.0534597
R18561 OUT_P.n1618 OUT_P.n1617 0.0534597
R18562 OUT_P.n1606 OUT_P.n1605 0.0534597
R18563 OUT_P.n1119 OUT_P.n1118 0.0534597
R18564 OUT_P.n1293 OUT_P.n1292 0.0534597
R18565 OUT_P.n1281 OUT_P.n1280 0.0534597
R18566 OUT_P.n1269 OUT_P.n1268 0.0534597
R18567 OUT_P.n1257 OUT_P.n1256 0.0534597
R18568 OUT_P.n1245 OUT_P.n1244 0.0534597
R18569 OUT_P.n1233 OUT_P.n1232 0.0534597
R18570 OUT_P.n1221 OUT_P.n1220 0.0534597
R18571 OUT_P.n1209 OUT_P.n1208 0.0534597
R18572 OUT_P.n1197 OUT_P.n1196 0.0534597
R18573 OUT_P.n1185 OUT_P.n1184 0.0534597
R18574 OUT_P.n1173 OUT_P.n1172 0.0534597
R18575 OUT_P.n1161 OUT_P.n1160 0.0534597
R18576 OUT_P.n1149 OUT_P.n1148 0.0534597
R18577 OUT_P.n1137 OUT_P.n1136 0.0534597
R18578 OUT_P.n9 OUT_P.n7 0.0423164
R18579 OUT_P.n20 OUT_P.n18 0.0423164
R18580 OUT_P.n30 OUT_P.n28 0.0423164
R18581 OUT_P.n135 OUT_P.n133 0.0423164
R18582 OUT_P.n146 OUT_P.n144 0.0423164
R18583 OUT_P.n156 OUT_P.n154 0.0423164
R18584 OUT_P.n165 OUT_P.n163 0.0423164
R18585 OUT_P.n176 OUT_P.n174 0.0423164
R18586 OUT_P.n186 OUT_P.n184 0.0423164
R18587 OUT_P.n206 OUT_P.n205 0.0420655
R18588 OUT_P.n1499 OUT_P.n1498 0.0419676
R18589 OUT_P.n103 OUT_P.n102 0.0419676
R18590 OUT_P.n544 OUT_P.n543 0.0419676
R18591 OUT_P.n70 OUT_P.n69 0.0419676
R18592 OUT_P.n1524 OUT_P.n1523 0.0415773
R18593 OUT_P.n1554 OUT_P.n1553 0.0415773
R18594 OUT_P.n988 OUT_P.n987 0.0415773
R18595 OUT_P.n947 OUT_P.n946 0.0415773
R18596 OUT_P.n932 OUT_P.n931 0.0415773
R18597 OUT_P.n919 OUT_P.n918 0.0415773
R18598 OUT_P.n571 OUT_P.n570 0.0415773
R18599 OUT_P.n583 OUT_P.n582 0.0415773
R18600 OUT_P.n592 OUT_P.n591 0.0415773
R18601 OUT_P.n604 OUT_P.n603 0.0415773
R18602 OUT_P.n613 OUT_P.n612 0.0415773
R18603 OUT_P.n625 OUT_P.n624 0.0415773
R18604 OUT_P.n634 OUT_P.n633 0.0415773
R18605 OUT_P.n646 OUT_P.n645 0.0415773
R18606 OUT_P.n655 OUT_P.n654 0.0415773
R18607 OUT_P.n667 OUT_P.n666 0.0415773
R18608 OUT_P.n676 OUT_P.n675 0.0415773
R18609 OUT_P.n688 OUT_P.n687 0.0415773
R18610 OUT_P.n697 OUT_P.n696 0.0415773
R18611 OUT_P.n709 OUT_P.n708 0.0415773
R18612 OUT_P.n44 OUT_P.n43 0.0415773
R18613 OUT_P.n1490 OUT_P.n1489 0.0415773
R18614 OUT_P.n1481 OUT_P.n1480 0.0415773
R18615 OUT_P.n1470 OUT_P.n1469 0.0415773
R18616 OUT_P.n1460 OUT_P.n1459 0.0415773
R18617 OUT_P.n1612 OUT_P.n1611 0.0415773
R18618 OUT_P.n1623 OUT_P.n1622 0.0415773
R18619 OUT_P.n1633 OUT_P.n1632 0.0415773
R18620 OUT_P.n1644 OUT_P.n1643 0.0415773
R18621 OUT_P.n1654 OUT_P.n1653 0.0415773
R18622 OUT_P.n1665 OUT_P.n1664 0.0415773
R18623 OUT_P.n1675 OUT_P.n1674 0.0415773
R18624 OUT_P.n1686 OUT_P.n1685 0.0415773
R18625 OUT_P.n1696 OUT_P.n1695 0.0415773
R18626 OUT_P.n1707 OUT_P.n1706 0.0415773
R18627 OUT_P.n1143 OUT_P.n1142 0.0415773
R18628 OUT_P.n1155 OUT_P.n1154 0.0415773
R18629 OUT_P.n1167 OUT_P.n1166 0.0415773
R18630 OUT_P.n1179 OUT_P.n1178 0.0415773
R18631 OUT_P.n1191 OUT_P.n1190 0.0415773
R18632 OUT_P.n1203 OUT_P.n1202 0.0415773
R18633 OUT_P.n1215 OUT_P.n1214 0.0415773
R18634 OUT_P.n1227 OUT_P.n1226 0.0415773
R18635 OUT_P.n1239 OUT_P.n1238 0.0415773
R18636 OUT_P.n1251 OUT_P.n1250 0.0415773
R18637 OUT_P.n1263 OUT_P.n1262 0.0415773
R18638 OUT_P.n1275 OUT_P.n1274 0.0415773
R18639 OUT_P.n1113 OUT_P.n1112 0.0415773
R18640 OUT_P.n1287 OUT_P.n1286 0.0415773
R18641 OUT_P.n1299 OUT_P.n1298 0.0415773
R18642 OUT_P.n101 OUT_P.n100 0.0415636
R18643 OUT_P.n911 OUT_P.n910 0.0415636
R18644 OUT_P.n114 OUT_P.n113 0.0334577
R18645 OUT_P.n1010 OUT_P.n903 0.0334577
R18646 OUT_P.n972 OUT_P.n971 0.0334577
R18647 OUT_P.n971 OUT_P.n970 0.0334577
R18648 OUT_P.n735 OUT_P.n734 0.0334577
R18649 OUT_P.n842 OUT_P.n828 0.0334577
R18650 OUT_P.n447 OUT_P.n446 0.0334577
R18651 OUT_P.n191 OUT_P.n190 0.0334577
R18652 OUT_P.n1774 OUT_P.n1773 0.0334577
R18653 OUT_P.n1814 OUT_P.n1813 0.0334577
R18654 OUT_P.n1090 OUT_P.t269 0.0306947
R18655 OUT_P.n1059 OUT_P.t270 0.0285465
R18656 OUT_P.n1933 OUT_P.n1932 0.0254881
R18657 OUT_P.n563 OUT_P.n562 0.0254881
R18658 OUT_P.n532 OUT_P.n531 0.0254881
R18659 OUT_P.n521 OUT_P.n520 0.0254881
R18660 OUT_P.n510 OUT_P.n509 0.0254881
R18661 OUT_P.n499 OUT_P.n498 0.0254881
R18662 OUT_P.n488 OUT_P.n487 0.0254881
R18663 OUT_P.n477 OUT_P.n476 0.0254881
R18664 OUT_P.n466 OUT_P.n465 0.0254881
R18665 OUT_P.n455 OUT_P.n454 0.0254881
R18666 OUT_P.n440 OUT_P.n439 0.0254881
R18667 OUT_P.n429 OUT_P.n428 0.0254881
R18668 OUT_P.n418 OUT_P.n417 0.0254881
R18669 OUT_P.n407 OUT_P.n406 0.0254881
R18670 OUT_P.n396 OUT_P.n395 0.0254881
R18671 OUT_P.n385 OUT_P.n384 0.0254881
R18672 OUT_P.n374 OUT_P.n373 0.0254881
R18673 OUT_P.n363 OUT_P.n362 0.0254881
R18674 OUT_P.n343 OUT_P.n342 0.0254881
R18675 OUT_P.n332 OUT_P.n331 0.0254881
R18676 OUT_P.n321 OUT_P.n320 0.0254881
R18677 OUT_P.n310 OUT_P.n309 0.0254881
R18678 OUT_P.n299 OUT_P.n298 0.0254881
R18679 OUT_P.n288 OUT_P.n287 0.0254881
R18680 OUT_P.n277 OUT_P.n276 0.0254881
R18681 OUT_P.n266 OUT_P.n265 0.0254881
R18682 OUT_P.n240 OUT_P.n239 0.0254881
R18683 OUT_P.n229 OUT_P.n228 0.0254881
R18684 OUT_P.n218 OUT_P.n217 0.0254881
R18685 OUT_P.n1821 OUT_P.n1820 0.0254881
R18686 OUT_P.n1832 OUT_P.n1831 0.0254881
R18687 OUT_P.n1843 OUT_P.n1842 0.0254881
R18688 OUT_P.n1852 OUT_P.n1851 0.0254881
R18689 OUT_P.n1862 OUT_P.n1861 0.0254881
R18690 OUT_P.n1873 OUT_P.n1872 0.0254881
R18691 OUT_P.n1884 OUT_P.n1883 0.0254881
R18692 OUT_P.n1893 OUT_P.n1892 0.0254881
R18693 OUT_P.n787 OUT_P.n786 0.0235313
R18694 OUT_P.n349 OUT_P.n348 0.0235313
R18695 OUT_P.n124 OUT_P.n123 0.0235313
R18696 OUT_P.n247 OUT_P.n246 0.0235313
R18697 OUT_P.n1365 OUT_P.n1364 0.0235313
R18698 OUT_P.n1406 OUT_P.n1405 0.0235313
R18699 OUT_P.n1447 OUT_P.n1446 0.0235313
R18700 OUT_P.n1 OUT_P.n0 0.0235313
R18701 OUT_P.n1898 OUT_P.n1897 0.0234412
R18702 OUT_P.n899 OUT_P.n898 0.0228651
R18703 OUT_P.n775 OUT_P.n774 0.0228651
R18704 OUT_P.n446 OUT_P.n445 0.0228651
R18705 OUT_P.n351 OUT_P.n350 0.0228651
R18706 OUT_P.n199 OUT_P.n197 0.0228651
R18707 OUT_P.n194 OUT_P.n192 0.0228651
R18708 OUT_P.n36 OUT_P.n35 0.0228651
R18709 OUT_P.n116 OUT_P.n115 0.0228651
R18710 OUT_P.n1515 OUT_P.n1514 0.0228651
R18711 OUT_P.n1567 OUT_P.n1566 0.0228651
R18712 OUT_P.n836 OUT_P.n835 0.0228651
R18713 OUT_P.n1812 OUT_P.n1811 0.0228651
R18714 OUT_P.n1727 OUT_P.n1726 0.0228651
R18715 OUT_P.n734 OUT_P.n733 0.0228651
R18716 OUT_P.n249 OUT_P.n248 0.0228651
R18717 OUT_P.n253 OUT_P.n252 0.0228651
R18718 OUT_P.n1729 OUT_P.n1728 0.0228651
R18719 OUT_P.n777 OUT_P.n776 0.0228651
R18720 OUT_P.n831 OUT_P.n830 0.0228651
R18721 OUT_P.n888 OUT_P.n887 0.0228651
R18722 OUT_P.n1916 OUT_P.n1915 0.0228651
R18723 OUT_P.n1919 OUT_P.n1918 0.0228651
R18724 OUT_P.n541 OUT_P.n191 0.0228651
R18725 OUT_P.n1923 OUT_P.n1922 0.0228651
R18726 OUT_P.n1098 OUT_P.n1097 0.0228651
R18727 OUT_P.n1453 OUT_P.n1452 0.0228651
R18728 OUT_P.n3 OUT_P.n2 0.0228651
R18729 OUT_P.n539 OUT_P.n538 0.0211167
R18730 OUT_P.n1065 OUT_P.n1064 0.0195244
R18731 OUT_P.n1066 OUT_P.n1065 0.0195244
R18732 OUT_P.n1067 OUT_P.n1066 0.0195244
R18733 OUT_P.n901 OUT_P.n897 0.0179841
R18734 OUT_P.n841 OUT_P.n829 0.0179841
R18735 OUT_P.n845 OUT_P.n842 0.0179841
R18736 OUT_P.n773 OUT_P.n772 0.0179841
R18737 OUT_P.n60 OUT_P.n59 0.0179841
R18738 OUT_P.n122 OUT_P.n121 0.0179841
R18739 OUT_P.n120 OUT_P.n119 0.0179841
R18740 OUT_P.n98 OUT_P.n97 0.0179841
R18741 OUT_P.n1540 OUT_P.n1518 0.0179841
R18742 OUT_P.n1517 OUT_P.n1516 0.0179841
R18743 OUT_P.n1570 OUT_P.n1569 0.0179841
R18744 OUT_P.n894 OUT_P.n893 0.0179841
R18745 OUT_P.n896 OUT_P.n895 0.0179841
R18746 OUT_P.n785 OUT_P.n784 0.0179841
R18747 OUT_P.n783 OUT_P.n782 0.0179841
R18748 OUT_P.n839 OUT_P.n838 0.0179841
R18749 OUT_P.n1772 OUT_P.n1771 0.0179841
R18750 OUT_P.n257 OUT_P.n250 0.0179841
R18751 OUT_P.n1321 OUT_P.n1320 0.0179841
R18752 OUT_P.n890 OUT_P.n889 0.0179841
R18753 OUT_P.n833 OUT_P.n832 0.0179841
R18754 OUT_P.n780 OUT_P.n779 0.0179841
R18755 OUT_P.n1318 OUT_P.n1317 0.0179841
R18756 OUT_P.n1324 OUT_P.n1323 0.0179841
R18757 OUT_P.n1129 OUT_P.n1107 0.0179841
R18758 OUT_P.n1906 OUT_P.n1905 0.0179841
R18759 OUT_P.n1908 OUT_P.n1907 0.0179841
R18760 OUT_P.n1914 OUT_P.n1913 0.0179841
R18761 OUT_P.n1010 OUT_P.n1009 0.0179841
R18762 OUT_P.n1950 OUT_P.n1927 0.0179841
R18763 OUT_P.n1601 OUT_P.n1454 0.0179841
R18764 OUT_P.n1106 OUT_P.n1105 0.0179841
R18765 OUT_P.n1096 OUT_P.n1011 0.0179841
R18766 OUT_P.n1952 OUT_P.n5 0.0179841
R18767 OUT_P.n841 OUT_P.n840 0.0177304
R18768 OUT_P.n901 OUT_P.n900 0.0177304
R18769 OUT_P.n844 OUT_P.n843 0.0177304
R18770 OUT_P.n846 OUT_P.n845 0.0177304
R18771 OUT_P.n779 OUT_P.n778 0.0177304
R18772 OUT_P.n774 OUT_P.n773 0.0177304
R18773 OUT_P.n353 OUT_P.n352 0.0177304
R18774 OUT_P.n114 OUT_P.n98 0.0177304
R18775 OUT_P.n121 OUT_P.n120 0.0177304
R18776 OUT_P.n119 OUT_P.n118 0.0177304
R18777 OUT_P.n38 OUT_P.n37 0.0177304
R18778 OUT_P.n1569 OUT_P.n1568 0.0177304
R18779 OUT_P.n895 OUT_P.n894 0.0177304
R18780 OUT_P.n893 OUT_P.n892 0.0177304
R18781 OUT_P.n1773 OUT_P.n1772 0.0177304
R18782 OUT_P.n838 OUT_P.n837 0.0177304
R18783 OUT_P.n784 OUT_P.n783 0.0177304
R18784 OUT_P.n782 OUT_P.n781 0.0177304
R18785 OUT_P.n257 OUT_P.n256 0.0177304
R18786 OUT_P.n891 OUT_P.n890 0.0177304
R18787 OUT_P.n834 OUT_P.n833 0.0177304
R18788 OUT_P.n1319 OUT_P.n1318 0.0177304
R18789 OUT_P.n1009 OUT_P.n1008 0.0177304
R18790 OUT_P.n1913 OUT_P.n1912 0.0177304
R18791 OUT_P.n1907 OUT_P.n1906 0.0177304
R18792 OUT_P.n1905 OUT_P.n1904 0.0177304
R18793 OUT_P.n1950 OUT_P.n1949 0.0177304
R18794 OUT_P.n1903 OUT_P.n1601 0.0177304
R18795 OUT_P.n1105 OUT_P.n1104 0.0177304
R18796 OUT_P.n1096 OUT_P.n1095 0.0177304
R18797 OUT_P.n5 OUT_P.n4 0.0177304
R18798 OUT_P.n201 OUT_P.n200 0.0174187
R18799 OUT_P.n196 OUT_P.n195 0.0174187
R18800 OUT_P.n254 OUT_P.n253 0.0174187
R18801 OUT_P.n255 OUT_P.n254 0.0174187
R18802 OUT_P.n1920 OUT_P.n1919 0.0174187
R18803 OUT_P.n1921 OUT_P.n1920 0.0174187
R18804 OUT_P.n1564 OUT_P.n1542 0.0173591
R18805 OUT_P.n1911 OUT_P.n1909 0.0173591
R18806 OUT_P.n790 OUT_P.n788 0.0173591
R18807 OUT_P.n790 OUT_P.n789 0.0173591
R18808 OUT_P.n246 OUT_P.n245 0.0173591
R18809 OUT_P.n355 OUT_P.n354 0.0173591
R18810 OUT_P.n354 OUT_P.n349 0.0173591
R18811 OUT_P.n128 OUT_P.n36 0.0173591
R18812 OUT_P.n84 OUT_P.n62 0.0173591
R18813 OUT_P.n61 OUT_P.n38 0.0173591
R18814 OUT_P.n126 OUT_P.n125 0.0173591
R18815 OUT_P.n1541 OUT_P.n1517 0.0173591
R18816 OUT_P.n84 OUT_P.n83 0.0173591
R18817 OUT_P.n127 OUT_P.n126 0.0173591
R18818 OUT_P.n129 OUT_P.n128 0.0173591
R18819 OUT_P.n1565 OUT_P.n1541 0.0173591
R18820 OUT_P.n1564 OUT_P.n1563 0.0173591
R18821 OUT_P.n85 OUT_P.n61 0.0173591
R18822 OUT_P.n1902 OUT_P.n1602 0.0173591
R18823 OUT_P.n1572 OUT_P.n1571 0.0173591
R18824 OUT_P.n1571 OUT_P.n1515 0.0173591
R18825 OUT_P.n1733 OUT_P.n1727 0.0173591
R18826 OUT_P.n1732 OUT_P.n1731 0.0173591
R18827 OUT_P.n1731 OUT_P.n1730 0.0173591
R18828 OUT_P.n1734 OUT_P.n1733 0.0173591
R18829 OUT_P.n245 OUT_P.n244 0.0173591
R18830 OUT_P.n1325 OUT_P.n1322 0.0173591
R18831 OUT_P.n1364 OUT_P.n1363 0.0173591
R18832 OUT_P.n1405 OUT_P.n1404 0.0173591
R18833 OUT_P.n1446 OUT_P.n1445 0.0173591
R18834 OUT_P.n1450 OUT_P.n1131 0.0173591
R18835 OUT_P.n1322 OUT_P.n1319 0.0173591
R18836 OUT_P.n1445 OUT_P.n1444 0.0173591
R18837 OUT_P.n1404 OUT_P.n1403 0.0173591
R18838 OUT_P.n1363 OUT_P.n1362 0.0173591
R18839 OUT_P.n1951 OUT_P.n1926 0.0173591
R18840 OUT_P.n1130 OUT_P.n1106 0.0173591
R18841 OUT_P.n1102 OUT_P.n1099 0.0173591
R18842 OUT_P.n1451 OUT_P.n1130 0.0173591
R18843 OUT_P.n1911 OUT_P.n1910 0.0173591
R18844 OUT_P.n1926 OUT_P.n1924 0.0173591
R18845 OUT_P.n1902 OUT_P.n1901 0.0173591
R18846 OUT_P.n1450 OUT_P.n1449 0.0173591
R18847 OUT_P.n1103 OUT_P.n1102 0.0173591
R18848 OUT_P.n1953 OUT_P.n1 0.0173591
R18849 OUT_P.n1954 OUT_P.n1953 0.0173591
R18850 OUT_P.n959 OUT_P.n955 0.0167343
R18851 OUT_P.n930 OUT_P.n929 0.0167343
R18852 OUT_P.n945 OUT_P.n944 0.0167343
R18853 OUT_P.n993 OUT_P.n992 0.0167343
R18854 OUT_P.n917 OUT_P.n916 0.0167343
R18855 OUT_P.n909 OUT_P.n908 0.0167343
R18856 OUT_P.n886 OUT_P.n885 0.0161314
R18857 OUT_P.n538 OUT_P.n537 0.0147026
R18858 OUT_P.n1083 OUT_P.n1082 0.0136473
R18859 OUT_P.n1082 OUT_P.n1081 0.0136473
R18860 OUT_P.n1899 OUT_P.n1898 0.0130374
R18861 OUT_P.n1900 OUT_P.n1899 0.0127848
R18862 OUT_P.n788 OUT_P.n787 0.0122638
R18863 OUT_P.n348 OUT_P.n347 0.0122638
R18864 OUT_P.n125 OUT_P.n124 0.0122638
R18865 OUT_P.n258 OUT_P.n247 0.0122638
R18866 OUT_P.n1366 OUT_P.n1365 0.0122638
R18867 OUT_P.n1407 OUT_P.n1406 0.0122638
R18868 OUT_P.n1448 OUT_P.n1447 0.0122638
R18869 OUT_P.n567 OUT_P.n542 0.0122638
R18870 OUT_P.n1600 OUT_P.n1455 0.0122638
R18871 OUT_P.n1101 OUT_P.n1100 0.0119325
R18872 OUT_P.n199 OUT_P.n198 0.0119325
R18873 OUT_P.n837 OUT_P.n836 0.0119325
R18874 OUT_P.n832 OUT_P.n831 0.0119325
R18875 OUT_P.n194 OUT_P.n193 0.0119325
R18876 OUT_P.n900 OUT_P.n899 0.0119325
R18877 OUT_P.n889 OUT_P.n888 0.0119325
R18878 OUT_P.n733 OUT_P.n732 0.0119325
R18879 OUT_P.n791 OUT_P.n775 0.0119325
R18880 OUT_P.n352 OUT_P.n351 0.0119325
R18881 OUT_P.n778 OUT_P.n777 0.0119325
R18882 OUT_P.n445 OUT_P.n444 0.0119325
R18883 OUT_P.n541 OUT_P.n540 0.0119325
R18884 OUT_P.n35 OUT_P.n34 0.0119325
R18885 OUT_P.n117 OUT_P.n116 0.0119325
R18886 OUT_P.n934 OUT_P.n933 0.0119325
R18887 OUT_P.n1568 OUT_P.n1567 0.0119325
R18888 OUT_P.n1514 OUT_P.n1513 0.0119325
R18889 OUT_P.n1726 OUT_P.n1725 0.0119325
R18890 OUT_P.n1813 OUT_P.n1812 0.0119325
R18891 OUT_P.n250 OUT_P.n249 0.0119325
R18892 OUT_P.n252 OUT_P.n251 0.0119325
R18893 OUT_P.n1730 OUT_P.n1729 0.0119325
R18894 OUT_P.n4 OUT_P.n3 0.0119325
R18895 OUT_P.n1924 OUT_P.n1923 0.0119325
R18896 OUT_P.n1918 OUT_P.n1917 0.0119325
R18897 OUT_P.n1915 OUT_P.n1914 0.0119325
R18898 OUT_P.n1454 OUT_P.n1453 0.0119325
R18899 OUT_P.n1099 OUT_P.n1098 0.0119325
R18900 OUT_P.n885 OUT_P.n884 0.0118313
R18901 OUT_P.n884 OUT_P.n883 0.0118313
R18902 OUT_P.n1057 OUT_P.n1055 0.0110972
R18903 OUT_P.n1061 OUT_P.n1058 0.0110972
R18904 OUT_P.n1092 OUT_P.n1089 0.0110972
R18905 OUT_P.n1061 OUT_P.n1060 0.010845
R18906 OUT_P.n1057 OUT_P.n1056 0.010845
R18907 OUT_P.n1051 OUT_P.n1050 0.010845
R18908 OUT_P.n1092 OUT_P.n1091 0.010845
R18909 OUT_P.n1085 OUT_P.n1084 0.010845
R18910 OUT_P.n1013 OUT_P.n1012 0.00964634
R18911 OUT_P.n1017 OUT_P.n1016 0.00964634
R18912 OUT_P.n1021 OUT_P.n1020 0.00964634
R18913 OUT_P.n1025 OUT_P.n1024 0.00964634
R18914 OUT_P.n1028 OUT_P.n1027 0.00964634
R18915 OUT_P.n1031 OUT_P.n1030 0.00964634
R18916 OUT_P.n1034 OUT_P.n1033 0.00964634
R18917 OUT_P.n1037 OUT_P.n1036 0.00964634
R18918 OUT_P.n1562 OUT_P.n1561 0.00905634
R18919 OUT_P.n1532 OUT_P.n1531 0.00905634
R18920 OUT_P.n96 OUT_P.n95 0.00905634
R18921 OUT_P.n107 OUT_P.n106 0.00905634
R18922 OUT_P.n553 OUT_P.n552 0.00905634
R18923 OUT_P.n997 OUT_P.n996 0.00905634
R18924 OUT_P.n717 OUT_P.n716 0.00905634
R18925 OUT_P.n726 OUT_P.n725 0.00905634
R18926 OUT_P.n739 OUT_P.n738 0.00905634
R18927 OUT_P.n748 OUT_P.n747 0.00905634
R18928 OUT_P.n757 OUT_P.n756 0.00905634
R18929 OUT_P.n766 OUT_P.n765 0.00905634
R18930 OUT_P.n795 OUT_P.n794 0.00905634
R18931 OUT_P.n804 OUT_P.n803 0.00905634
R18932 OUT_P.n813 OUT_P.n812 0.00905634
R18933 OUT_P.n822 OUT_P.n821 0.00905634
R18934 OUT_P.n850 OUT_P.n849 0.00905634
R18935 OUT_P.n859 OUT_P.n858 0.00905634
R18936 OUT_P.n868 OUT_P.n867 0.00905634
R18937 OUT_P.n877 OUT_P.n876 0.00905634
R18938 OUT_P.n210 OUT_P.n209 0.00905634
R18939 OUT_P.n12 OUT_P.n11 0.00905634
R18940 OUT_P.n53 OUT_P.n52 0.00905634
R18941 OUT_P.n80 OUT_P.n79 0.00905634
R18942 OUT_P.n1592 OUT_P.n1591 0.00905634
R18943 OUT_P.n1583 OUT_P.n1582 0.00905634
R18944 OUT_P.n1574 OUT_P.n1573 0.00905634
R18945 OUT_P.n1505 OUT_P.n1504 0.00905634
R18946 OUT_P.n1503 OUT_P.n1502 0.00905634
R18947 OUT_P.n1715 OUT_P.n1714 0.00905634
R18948 OUT_P.n1724 OUT_P.n1723 0.00905634
R18949 OUT_P.n1743 OUT_P.n1742 0.00905634
R18950 OUT_P.n1752 OUT_P.n1751 0.00905634
R18951 OUT_P.n1761 OUT_P.n1760 0.00905634
R18952 OUT_P.n1770 OUT_P.n1769 0.00905634
R18953 OUT_P.n1783 OUT_P.n1782 0.00905634
R18954 OUT_P.n1792 OUT_P.n1791 0.00905634
R18955 OUT_P.n1801 OUT_P.n1800 0.00905634
R18956 OUT_P.n1810 OUT_P.n1809 0.00905634
R18957 OUT_P.n1307 OUT_P.n1306 0.00905634
R18958 OUT_P.n1316 OUT_P.n1315 0.00905634
R18959 OUT_P.n1334 OUT_P.n1333 0.00905634
R18960 OUT_P.n1343 OUT_P.n1342 0.00905634
R18961 OUT_P.n1352 OUT_P.n1351 0.00905634
R18962 OUT_P.n1361 OUT_P.n1360 0.00905634
R18963 OUT_P.n1375 OUT_P.n1374 0.00905634
R18964 OUT_P.n1384 OUT_P.n1383 0.00905634
R18965 OUT_P.n1393 OUT_P.n1392 0.00905634
R18966 OUT_P.n1402 OUT_P.n1401 0.00905634
R18967 OUT_P.n1416 OUT_P.n1415 0.00905634
R18968 OUT_P.n1425 OUT_P.n1424 0.00905634
R18969 OUT_P.n1434 OUT_P.n1433 0.00905634
R18970 OUT_P.n1443 OUT_P.n1442 0.00905634
R18971 OUT_P.n1121 OUT_P.n1120 0.00905634
R18972 OUT_P.n902 OUT_P.n886 0.00856444
R18973 OUT_P.n1042 OUT_P.n1041 0.008
R18974 OUT_P.n1045 OUT_P.n1044 0.008
R18975 OUT_P.n1048 OUT_P.n1047 0.008
R18976 OUT_P.n1054 OUT_P.n1053 0.008
R18977 OUT_P.n1073 OUT_P.n1072 0.008
R18978 OUT_P.n1076 OUT_P.n1075 0.008
R18979 OUT_P.n1079 OUT_P.n1078 0.008
R18980 OUT_P.n1088 OUT_P.n1087 0.008
R18981 OUT_P.n537 OUT_P.n536 0.00785132
R18982 OUT_P.n1943 OUT_P.n1942 0.00735609
R18983 OUT_P.n1948 OUT_P.n1947 0.00735609
R18984 OUT_P.n566 OUT_P.n565 0.00735609
R18985 OUT_P.n964 OUT_P.n963 0.00735609
R18986 OUT_P.n526 OUT_P.n525 0.00735609
R18987 OUT_P.n515 OUT_P.n514 0.00735609
R18988 OUT_P.n504 OUT_P.n503 0.00735609
R18989 OUT_P.n493 OUT_P.n492 0.00735609
R18990 OUT_P.n482 OUT_P.n481 0.00735609
R18991 OUT_P.n471 OUT_P.n470 0.00735609
R18992 OUT_P.n460 OUT_P.n459 0.00735609
R18993 OUT_P.n449 OUT_P.n448 0.00735609
R18994 OUT_P.n434 OUT_P.n433 0.00735609
R18995 OUT_P.n423 OUT_P.n422 0.00735609
R18996 OUT_P.n412 OUT_P.n411 0.00735609
R18997 OUT_P.n401 OUT_P.n400 0.00735609
R18998 OUT_P.n390 OUT_P.n389 0.00735609
R18999 OUT_P.n379 OUT_P.n378 0.00735609
R19000 OUT_P.n368 OUT_P.n367 0.00735609
R19001 OUT_P.n357 OUT_P.n356 0.00735609
R19002 OUT_P.n337 OUT_P.n336 0.00735609
R19003 OUT_P.n326 OUT_P.n325 0.00735609
R19004 OUT_P.n315 OUT_P.n314 0.00735609
R19005 OUT_P.n304 OUT_P.n303 0.00735609
R19006 OUT_P.n293 OUT_P.n292 0.00735609
R19007 OUT_P.n282 OUT_P.n281 0.00735609
R19008 OUT_P.n271 OUT_P.n270 0.00735609
R19009 OUT_P.n260 OUT_P.n259 0.00735609
R19010 OUT_P.n234 OUT_P.n233 0.00735609
R19011 OUT_P.n223 OUT_P.n222 0.00735609
R19012 OUT_P.n212 OUT_P.n211 0.00735609
R19013 OUT_P.n1816 OUT_P.n1815 0.00735609
R19014 OUT_P.n1826 OUT_P.n1825 0.00735609
R19015 OUT_P.n1837 OUT_P.n1836 0.00735609
R19016 OUT_P.n1848 OUT_P.n1847 0.00735609
R19017 OUT_P.n1857 OUT_P.n1856 0.00735609
R19018 OUT_P.n1867 OUT_P.n1866 0.00735609
R19019 OUT_P.n1878 OUT_P.n1877 0.00735609
R19020 OUT_P.n1889 OUT_P.n1888 0.00735609
R19021 OUT_P.n1084 OUT_P.n1083 0.00732364
R19022 OUT_P.n1081 OUT_P.n1080 0.00732364
R19023 OUT_P.n1015 OUT_P.n1013 0.00543902
R19024 OUT_P.n1016 OUT_P.n1015 0.00543902
R19025 OUT_P.n1019 OUT_P.n1017 0.00543902
R19026 OUT_P.n1020 OUT_P.n1019 0.00543902
R19027 OUT_P.n1023 OUT_P.n1021 0.00543902
R19028 OUT_P.n1024 OUT_P.n1023 0.00543902
R19029 OUT_P.n1026 OUT_P.n1025 0.00543902
R19030 OUT_P.n1029 OUT_P.n1028 0.00543902
R19031 OUT_P.n1030 OUT_P.n1029 0.00543902
R19032 OUT_P.n1032 OUT_P.n1031 0.00543902
R19033 OUT_P.n1033 OUT_P.n1032 0.00543902
R19034 OUT_P.n1035 OUT_P.n1034 0.00543902
R19035 OUT_P.n1036 OUT_P.n1035 0.00543902
R19036 OUT_P.n1038 OUT_P.n1037 0.00543902
R19037 OUT_P.n1302 OUT_P.n1301 0.00528925
R19038 OUT_P.n1306 OUT_P.n1305 0.00528925
R19039 OUT_P.n1311 OUT_P.n1310 0.00528925
R19040 OUT_P.n1122 OUT_P.n1121 0.00528925
R19041 OUT_P.n1126 OUT_P.n1125 0.00528925
R19042 OUT_P.n1710 OUT_P.n1709 0.00528925
R19043 OUT_P.n1714 OUT_P.n1713 0.00528925
R19044 OUT_P.n1719 OUT_P.n1718 0.00528925
R19045 OUT_P.n1723 OUT_P.n1722 0.00528925
R19046 OUT_P.n1738 OUT_P.n1737 0.00528925
R19047 OUT_P.n1742 OUT_P.n1741 0.00528925
R19048 OUT_P.n1747 OUT_P.n1746 0.00528925
R19049 OUT_P.n1751 OUT_P.n1750 0.00528925
R19050 OUT_P.n1756 OUT_P.n1755 0.00528925
R19051 OUT_P.n1760 OUT_P.n1759 0.00528925
R19052 OUT_P.n1765 OUT_P.n1764 0.00528925
R19053 OUT_P.n1769 OUT_P.n1768 0.00528925
R19054 OUT_P.n1778 OUT_P.n1777 0.00528925
R19055 OUT_P.n1782 OUT_P.n1781 0.00528925
R19056 OUT_P.n1787 OUT_P.n1786 0.00528925
R19057 OUT_P.n1791 OUT_P.n1790 0.00528925
R19058 OUT_P.n1796 OUT_P.n1795 0.00528925
R19059 OUT_P.n1800 OUT_P.n1799 0.00528925
R19060 OUT_P.n1805 OUT_P.n1804 0.00528925
R19061 OUT_P.n1809 OUT_P.n1808 0.00528925
R19062 OUT_P.n1597 OUT_P.n1596 0.00528925
R19063 OUT_P.n1593 OUT_P.n1592 0.00528925
R19064 OUT_P.n1588 OUT_P.n1587 0.00528925
R19065 OUT_P.n1584 OUT_P.n1583 0.00528925
R19066 OUT_P.n1579 OUT_P.n1578 0.00528925
R19067 OUT_P.n1506 OUT_P.n1505 0.00528925
R19068 OUT_P.n1510 OUT_P.n1509 0.00528925
R19069 OUT_P.n1575 OUT_P.n1574 0.00528925
R19070 OUT_P.n1557 OUT_P.n1556 0.00528925
R19071 OUT_P.n1533 OUT_P.n1532 0.00528925
R19072 OUT_P.n1537 OUT_P.n1536 0.00528925
R19073 OUT_P.n1561 OUT_P.n1560 0.00528925
R19074 OUT_P.n716 OUT_P.n715 0.00528925
R19075 OUT_P.n721 OUT_P.n720 0.00528925
R19076 OUT_P.n725 OUT_P.n724 0.00528925
R19077 OUT_P.n730 OUT_P.n729 0.00528925
R19078 OUT_P.n738 OUT_P.n737 0.00528925
R19079 OUT_P.n743 OUT_P.n742 0.00528925
R19080 OUT_P.n747 OUT_P.n746 0.00528925
R19081 OUT_P.n752 OUT_P.n751 0.00528925
R19082 OUT_P.n756 OUT_P.n755 0.00528925
R19083 OUT_P.n761 OUT_P.n760 0.00528925
R19084 OUT_P.n765 OUT_P.n764 0.00528925
R19085 OUT_P.n770 OUT_P.n769 0.00528925
R19086 OUT_P.n794 OUT_P.n793 0.00528925
R19087 OUT_P.n799 OUT_P.n798 0.00528925
R19088 OUT_P.n803 OUT_P.n802 0.00528925
R19089 OUT_P.n808 OUT_P.n807 0.00528925
R19090 OUT_P.n812 OUT_P.n811 0.00528925
R19091 OUT_P.n817 OUT_P.n816 0.00528925
R19092 OUT_P.n821 OUT_P.n820 0.00528925
R19093 OUT_P.n826 OUT_P.n825 0.00528925
R19094 OUT_P.n849 OUT_P.n848 0.00528925
R19095 OUT_P.n854 OUT_P.n853 0.00528925
R19096 OUT_P.n858 OUT_P.n857 0.00528925
R19097 OUT_P.n863 OUT_P.n862 0.00528925
R19098 OUT_P.n867 OUT_P.n866 0.00528925
R19099 OUT_P.n872 OUT_P.n871 0.00528925
R19100 OUT_P.n876 OUT_P.n875 0.00528925
R19101 OUT_P.n881 OUT_P.n880 0.00528925
R19102 OUT_P.n91 OUT_P.n90 0.00528925
R19103 OUT_P.n976 OUT_P.n975 0.00528925
R19104 OUT_P.n95 OUT_P.n94 0.00528925
R19105 OUT_P.n968 OUT_P.n967 0.00528925
R19106 OUT_P.n111 OUT_P.n110 0.00528925
R19107 OUT_P.n1001 OUT_P.n1000 0.00528925
R19108 OUT_P.n1006 OUT_P.n1005 0.00528925
R19109 OUT_P.n52 OUT_P.n51 0.00528925
R19110 OUT_P.n57 OUT_P.n56 0.00528925
R19111 OUT_P.n81 OUT_P.n80 0.00528925
R19112 OUT_P.n77 OUT_P.n76 0.00528925
R19113 OUT_P.n1315 OUT_P.n1314 0.00528925
R19114 OUT_P.n1329 OUT_P.n1328 0.00528925
R19115 OUT_P.n1333 OUT_P.n1332 0.00528925
R19116 OUT_P.n1338 OUT_P.n1337 0.00528925
R19117 OUT_P.n1342 OUT_P.n1341 0.00528925
R19118 OUT_P.n1347 OUT_P.n1346 0.00528925
R19119 OUT_P.n1351 OUT_P.n1350 0.00528925
R19120 OUT_P.n1356 OUT_P.n1355 0.00528925
R19121 OUT_P.n1360 OUT_P.n1359 0.00528925
R19122 OUT_P.n1370 OUT_P.n1369 0.00528925
R19123 OUT_P.n1374 OUT_P.n1373 0.00528925
R19124 OUT_P.n1379 OUT_P.n1378 0.00528925
R19125 OUT_P.n1383 OUT_P.n1382 0.00528925
R19126 OUT_P.n1388 OUT_P.n1387 0.00528925
R19127 OUT_P.n1392 OUT_P.n1391 0.00528925
R19128 OUT_P.n1397 OUT_P.n1396 0.00528925
R19129 OUT_P.n1401 OUT_P.n1400 0.00528925
R19130 OUT_P.n1411 OUT_P.n1410 0.00528925
R19131 OUT_P.n1415 OUT_P.n1414 0.00528925
R19132 OUT_P.n1420 OUT_P.n1419 0.00528925
R19133 OUT_P.n1424 OUT_P.n1423 0.00528925
R19134 OUT_P.n1429 OUT_P.n1428 0.00528925
R19135 OUT_P.n1433 OUT_P.n1432 0.00528925
R19136 OUT_P.n1438 OUT_P.n1437 0.00528925
R19137 OUT_P.n1442 OUT_P.n1441 0.00528925
R19138 OUT_P.n1945 OUT_P.n1944 0.00527411
R19139 OUT_P.n1946 OUT_P.n1945 0.00527411
R19140 OUT_P.n1539 OUT_P.n1538 0.00527411
R19141 OUT_P.n1538 OUT_P.n1537 0.00527411
R19142 OUT_P.n1556 OUT_P.n1555 0.00527411
R19143 OUT_P.n109 OUT_P.n108 0.00527411
R19144 OUT_P.n90 OUT_P.n89 0.00527411
R19145 OUT_P.n110 OUT_P.n109 0.00527411
R19146 OUT_P.n555 OUT_P.n554 0.00527411
R19147 OUT_P.n564 OUT_P.n555 0.00527411
R19148 OUT_P.n1004 OUT_P.n1003 0.00527411
R19149 OUT_P.n999 OUT_P.n998 0.00527411
R19150 OUT_P.n979 OUT_P.n978 0.00527411
R19151 OUT_P.n974 OUT_P.n973 0.00527411
R19152 OUT_P.n966 OUT_P.n965 0.00527411
R19153 OUT_P.n1000 OUT_P.n999 0.00527411
R19154 OUT_P.n975 OUT_P.n974 0.00527411
R19155 OUT_P.n967 OUT_P.n966 0.00527411
R19156 OUT_P.n996 OUT_P.n979 0.00527411
R19157 OUT_P.n1005 OUT_P.n1004 0.00527411
R19158 OUT_P.n719 OUT_P.n718 0.00527411
R19159 OUT_P.n728 OUT_P.n727 0.00527411
R19160 OUT_P.n741 OUT_P.n740 0.00527411
R19161 OUT_P.n750 OUT_P.n749 0.00527411
R19162 OUT_P.n759 OUT_P.n758 0.00527411
R19163 OUT_P.n768 OUT_P.n767 0.00527411
R19164 OUT_P.n797 OUT_P.n796 0.00527411
R19165 OUT_P.n806 OUT_P.n805 0.00527411
R19166 OUT_P.n815 OUT_P.n814 0.00527411
R19167 OUT_P.n824 OUT_P.n823 0.00527411
R19168 OUT_P.n852 OUT_P.n851 0.00527411
R19169 OUT_P.n861 OUT_P.n860 0.00527411
R19170 OUT_P.n870 OUT_P.n869 0.00527411
R19171 OUT_P.n879 OUT_P.n878 0.00527411
R19172 OUT_P.n880 OUT_P.n879 0.00527411
R19173 OUT_P.n871 OUT_P.n870 0.00527411
R19174 OUT_P.n862 OUT_P.n861 0.00527411
R19175 OUT_P.n853 OUT_P.n852 0.00527411
R19176 OUT_P.n825 OUT_P.n824 0.00527411
R19177 OUT_P.n816 OUT_P.n815 0.00527411
R19178 OUT_P.n807 OUT_P.n806 0.00527411
R19179 OUT_P.n798 OUT_P.n797 0.00527411
R19180 OUT_P.n769 OUT_P.n768 0.00527411
R19181 OUT_P.n760 OUT_P.n759 0.00527411
R19182 OUT_P.n751 OUT_P.n750 0.00527411
R19183 OUT_P.n742 OUT_P.n741 0.00527411
R19184 OUT_P.n729 OUT_P.n728 0.00527411
R19185 OUT_P.n720 OUT_P.n719 0.00527411
R19186 OUT_P.n221 OUT_P.n220 0.00527411
R19187 OUT_P.n232 OUT_P.n231 0.00527411
R19188 OUT_P.n243 OUT_P.n242 0.00527411
R19189 OUT_P.n269 OUT_P.n268 0.00527411
R19190 OUT_P.n280 OUT_P.n279 0.00527411
R19191 OUT_P.n291 OUT_P.n290 0.00527411
R19192 OUT_P.n302 OUT_P.n301 0.00527411
R19193 OUT_P.n313 OUT_P.n312 0.00527411
R19194 OUT_P.n324 OUT_P.n323 0.00527411
R19195 OUT_P.n335 OUT_P.n334 0.00527411
R19196 OUT_P.n346 OUT_P.n345 0.00527411
R19197 OUT_P.n366 OUT_P.n365 0.00527411
R19198 OUT_P.n377 OUT_P.n376 0.00527411
R19199 OUT_P.n388 OUT_P.n387 0.00527411
R19200 OUT_P.n399 OUT_P.n398 0.00527411
R19201 OUT_P.n410 OUT_P.n409 0.00527411
R19202 OUT_P.n421 OUT_P.n420 0.00527411
R19203 OUT_P.n432 OUT_P.n431 0.00527411
R19204 OUT_P.n443 OUT_P.n442 0.00527411
R19205 OUT_P.n458 OUT_P.n457 0.00527411
R19206 OUT_P.n469 OUT_P.n468 0.00527411
R19207 OUT_P.n480 OUT_P.n479 0.00527411
R19208 OUT_P.n491 OUT_P.n490 0.00527411
R19209 OUT_P.n502 OUT_P.n501 0.00527411
R19210 OUT_P.n513 OUT_P.n512 0.00527411
R19211 OUT_P.n524 OUT_P.n523 0.00527411
R19212 OUT_P.n535 OUT_P.n534 0.00527411
R19213 OUT_P.n534 OUT_P.n533 0.00527411
R19214 OUT_P.n523 OUT_P.n522 0.00527411
R19215 OUT_P.n512 OUT_P.n511 0.00527411
R19216 OUT_P.n501 OUT_P.n500 0.00527411
R19217 OUT_P.n490 OUT_P.n489 0.00527411
R19218 OUT_P.n479 OUT_P.n478 0.00527411
R19219 OUT_P.n468 OUT_P.n467 0.00527411
R19220 OUT_P.n457 OUT_P.n456 0.00527411
R19221 OUT_P.n442 OUT_P.n441 0.00527411
R19222 OUT_P.n431 OUT_P.n430 0.00527411
R19223 OUT_P.n420 OUT_P.n419 0.00527411
R19224 OUT_P.n409 OUT_P.n408 0.00527411
R19225 OUT_P.n398 OUT_P.n397 0.00527411
R19226 OUT_P.n387 OUT_P.n386 0.00527411
R19227 OUT_P.n376 OUT_P.n375 0.00527411
R19228 OUT_P.n365 OUT_P.n364 0.00527411
R19229 OUT_P.n345 OUT_P.n344 0.00527411
R19230 OUT_P.n334 OUT_P.n333 0.00527411
R19231 OUT_P.n323 OUT_P.n322 0.00527411
R19232 OUT_P.n312 OUT_P.n311 0.00527411
R19233 OUT_P.n301 OUT_P.n300 0.00527411
R19234 OUT_P.n290 OUT_P.n289 0.00527411
R19235 OUT_P.n279 OUT_P.n278 0.00527411
R19236 OUT_P.n268 OUT_P.n267 0.00527411
R19237 OUT_P.n242 OUT_P.n241 0.00527411
R19238 OUT_P.n231 OUT_P.n230 0.00527411
R19239 OUT_P.n220 OUT_P.n219 0.00527411
R19240 OUT_P.n188 OUT_P.n187 0.00527411
R19241 OUT_P.n181 OUT_P.n180 0.00527411
R19242 OUT_P.n178 OUT_P.n177 0.00527411
R19243 OUT_P.n170 OUT_P.n169 0.00527411
R19244 OUT_P.n167 OUT_P.n166 0.00527411
R19245 OUT_P.n161 OUT_P.n160 0.00527411
R19246 OUT_P.n158 OUT_P.n157 0.00527411
R19247 OUT_P.n151 OUT_P.n150 0.00527411
R19248 OUT_P.n148 OUT_P.n147 0.00527411
R19249 OUT_P.n140 OUT_P.n139 0.00527411
R19250 OUT_P.n137 OUT_P.n136 0.00527411
R19251 OUT_P.n131 OUT_P.n130 0.00527411
R19252 OUT_P.n32 OUT_P.n31 0.00527411
R19253 OUT_P.n25 OUT_P.n24 0.00527411
R19254 OUT_P.n22 OUT_P.n21 0.00527411
R19255 OUT_P.n14 OUT_P.n13 0.00527411
R19256 OUT_P.n23 OUT_P.n22 0.00527411
R19257 OUT_P.n21 OUT_P.n14 0.00527411
R19258 OUT_P.n33 OUT_P.n32 0.00527411
R19259 OUT_P.n31 OUT_P.n25 0.00527411
R19260 OUT_P.n138 OUT_P.n137 0.00527411
R19261 OUT_P.n136 OUT_P.n131 0.00527411
R19262 OUT_P.n149 OUT_P.n148 0.00527411
R19263 OUT_P.n147 OUT_P.n140 0.00527411
R19264 OUT_P.n159 OUT_P.n158 0.00527411
R19265 OUT_P.n157 OUT_P.n151 0.00527411
R19266 OUT_P.n168 OUT_P.n167 0.00527411
R19267 OUT_P.n166 OUT_P.n161 0.00527411
R19268 OUT_P.n179 OUT_P.n178 0.00527411
R19269 OUT_P.n177 OUT_P.n170 0.00527411
R19270 OUT_P.n189 OUT_P.n188 0.00527411
R19271 OUT_P.n187 OUT_P.n181 0.00527411
R19272 OUT_P.n55 OUT_P.n54 0.00527411
R19273 OUT_P.n56 OUT_P.n55 0.00527411
R19274 OUT_P.n1599 OUT_P.n1598 0.00527411
R19275 OUT_P.n1590 OUT_P.n1589 0.00527411
R19276 OUT_P.n1581 OUT_P.n1580 0.00527411
R19277 OUT_P.n1512 OUT_P.n1511 0.00527411
R19278 OUT_P.n1511 OUT_P.n1510 0.00527411
R19279 OUT_P.n1580 OUT_P.n1579 0.00527411
R19280 OUT_P.n1589 OUT_P.n1588 0.00527411
R19281 OUT_P.n1598 OUT_P.n1597 0.00527411
R19282 OUT_P.n1717 OUT_P.n1716 0.00527411
R19283 OUT_P.n1736 OUT_P.n1735 0.00527411
R19284 OUT_P.n1745 OUT_P.n1744 0.00527411
R19285 OUT_P.n1754 OUT_P.n1753 0.00527411
R19286 OUT_P.n1763 OUT_P.n1762 0.00527411
R19287 OUT_P.n1776 OUT_P.n1775 0.00527411
R19288 OUT_P.n1785 OUT_P.n1784 0.00527411
R19289 OUT_P.n1794 OUT_P.n1793 0.00527411
R19290 OUT_P.n1803 OUT_P.n1802 0.00527411
R19291 OUT_P.n1824 OUT_P.n1823 0.00527411
R19292 OUT_P.n1835 OUT_P.n1834 0.00527411
R19293 OUT_P.n1846 OUT_P.n1845 0.00527411
R19294 OUT_P.n1855 OUT_P.n1854 0.00527411
R19295 OUT_P.n1865 OUT_P.n1864 0.00527411
R19296 OUT_P.n1876 OUT_P.n1875 0.00527411
R19297 OUT_P.n1887 OUT_P.n1886 0.00527411
R19298 OUT_P.n1896 OUT_P.n1895 0.00527411
R19299 OUT_P.n1823 OUT_P.n1822 0.00527411
R19300 OUT_P.n1834 OUT_P.n1833 0.00527411
R19301 OUT_P.n1845 OUT_P.n1844 0.00527411
R19302 OUT_P.n1854 OUT_P.n1853 0.00527411
R19303 OUT_P.n1864 OUT_P.n1863 0.00527411
R19304 OUT_P.n1875 OUT_P.n1874 0.00527411
R19305 OUT_P.n1886 OUT_P.n1885 0.00527411
R19306 OUT_P.n1895 OUT_P.n1894 0.00527411
R19307 OUT_P.n1804 OUT_P.n1803 0.00527411
R19308 OUT_P.n1795 OUT_P.n1794 0.00527411
R19309 OUT_P.n1786 OUT_P.n1785 0.00527411
R19310 OUT_P.n1777 OUT_P.n1776 0.00527411
R19311 OUT_P.n1764 OUT_P.n1763 0.00527411
R19312 OUT_P.n1755 OUT_P.n1754 0.00527411
R19313 OUT_P.n1746 OUT_P.n1745 0.00527411
R19314 OUT_P.n1737 OUT_P.n1736 0.00527411
R19315 OUT_P.n1718 OUT_P.n1717 0.00527411
R19316 OUT_P.n1709 OUT_P.n1708 0.00527411
R19317 OUT_P.n1309 OUT_P.n1308 0.00527411
R19318 OUT_P.n1327 OUT_P.n1326 0.00527411
R19319 OUT_P.n1336 OUT_P.n1335 0.00527411
R19320 OUT_P.n1345 OUT_P.n1344 0.00527411
R19321 OUT_P.n1354 OUT_P.n1353 0.00527411
R19322 OUT_P.n1368 OUT_P.n1367 0.00527411
R19323 OUT_P.n1377 OUT_P.n1376 0.00527411
R19324 OUT_P.n1386 OUT_P.n1385 0.00527411
R19325 OUT_P.n1395 OUT_P.n1394 0.00527411
R19326 OUT_P.n1409 OUT_P.n1408 0.00527411
R19327 OUT_P.n1418 OUT_P.n1417 0.00527411
R19328 OUT_P.n1427 OUT_P.n1426 0.00527411
R19329 OUT_P.n1436 OUT_P.n1435 0.00527411
R19330 OUT_P.n1128 OUT_P.n1127 0.00527411
R19331 OUT_P.n1437 OUT_P.n1436 0.00527411
R19332 OUT_P.n1428 OUT_P.n1427 0.00527411
R19333 OUT_P.n1419 OUT_P.n1418 0.00527411
R19334 OUT_P.n1410 OUT_P.n1409 0.00527411
R19335 OUT_P.n1396 OUT_P.n1395 0.00527411
R19336 OUT_P.n1387 OUT_P.n1386 0.00527411
R19337 OUT_P.n1378 OUT_P.n1377 0.00527411
R19338 OUT_P.n1369 OUT_P.n1368 0.00527411
R19339 OUT_P.n1355 OUT_P.n1354 0.00527411
R19340 OUT_P.n1346 OUT_P.n1345 0.00527411
R19341 OUT_P.n1337 OUT_P.n1336 0.00527411
R19342 OUT_P.n1328 OUT_P.n1327 0.00527411
R19343 OUT_P.n1127 OUT_P.n1126 0.00527411
R19344 OUT_P.n1310 OUT_P.n1309 0.00527411
R19345 OUT_P.n1301 OUT_P.n1300 0.00527411
R19346 OUT_P.n1558 OUT_P.n1557 0.00525899
R19347 OUT_P.n1560 OUT_P.n1559 0.00525899
R19348 OUT_P.n1536 OUT_P.n1535 0.00525899
R19349 OUT_P.n1534 OUT_P.n1533 0.00525899
R19350 OUT_P.n92 OUT_P.n91 0.00525899
R19351 OUT_P.n94 OUT_P.n93 0.00525899
R19352 OUT_P.n112 OUT_P.n111 0.00525899
R19353 OUT_P.n1002 OUT_P.n1001 0.00525899
R19354 OUT_P.n977 OUT_P.n976 0.00525899
R19355 OUT_P.n969 OUT_P.n968 0.00525899
R19356 OUT_P.n1007 OUT_P.n1006 0.00525899
R19357 OUT_P.n722 OUT_P.n721 0.00525899
R19358 OUT_P.n724 OUT_P.n723 0.00525899
R19359 OUT_P.n731 OUT_P.n730 0.00525899
R19360 OUT_P.n737 OUT_P.n736 0.00525899
R19361 OUT_P.n744 OUT_P.n743 0.00525899
R19362 OUT_P.n746 OUT_P.n745 0.00525899
R19363 OUT_P.n753 OUT_P.n752 0.00525899
R19364 OUT_P.n755 OUT_P.n754 0.00525899
R19365 OUT_P.n762 OUT_P.n761 0.00525899
R19366 OUT_P.n764 OUT_P.n763 0.00525899
R19367 OUT_P.n771 OUT_P.n770 0.00525899
R19368 OUT_P.n793 OUT_P.n792 0.00525899
R19369 OUT_P.n800 OUT_P.n799 0.00525899
R19370 OUT_P.n802 OUT_P.n801 0.00525899
R19371 OUT_P.n809 OUT_P.n808 0.00525899
R19372 OUT_P.n811 OUT_P.n810 0.00525899
R19373 OUT_P.n818 OUT_P.n817 0.00525899
R19374 OUT_P.n820 OUT_P.n819 0.00525899
R19375 OUT_P.n827 OUT_P.n826 0.00525899
R19376 OUT_P.n848 OUT_P.n847 0.00525899
R19377 OUT_P.n855 OUT_P.n854 0.00525899
R19378 OUT_P.n857 OUT_P.n856 0.00525899
R19379 OUT_P.n864 OUT_P.n863 0.00525899
R19380 OUT_P.n866 OUT_P.n865 0.00525899
R19381 OUT_P.n873 OUT_P.n872 0.00525899
R19382 OUT_P.n875 OUT_P.n874 0.00525899
R19383 OUT_P.n882 OUT_P.n881 0.00525899
R19384 OUT_P.n58 OUT_P.n57 0.00525899
R19385 OUT_P.n82 OUT_P.n81 0.00525899
R19386 OUT_P.n78 OUT_P.n77 0.00525899
R19387 OUT_P.n1596 OUT_P.n1595 0.00525899
R19388 OUT_P.n1594 OUT_P.n1593 0.00525899
R19389 OUT_P.n1587 OUT_P.n1586 0.00525899
R19390 OUT_P.n1585 OUT_P.n1584 0.00525899
R19391 OUT_P.n1578 OUT_P.n1577 0.00525899
R19392 OUT_P.n1576 OUT_P.n1575 0.00525899
R19393 OUT_P.n1509 OUT_P.n1508 0.00525899
R19394 OUT_P.n1507 OUT_P.n1506 0.00525899
R19395 OUT_P.n1711 OUT_P.n1710 0.00525899
R19396 OUT_P.n1713 OUT_P.n1712 0.00525899
R19397 OUT_P.n1720 OUT_P.n1719 0.00525899
R19398 OUT_P.n1722 OUT_P.n1721 0.00525899
R19399 OUT_P.n1739 OUT_P.n1738 0.00525899
R19400 OUT_P.n1741 OUT_P.n1740 0.00525899
R19401 OUT_P.n1748 OUT_P.n1747 0.00525899
R19402 OUT_P.n1750 OUT_P.n1749 0.00525899
R19403 OUT_P.n1757 OUT_P.n1756 0.00525899
R19404 OUT_P.n1759 OUT_P.n1758 0.00525899
R19405 OUT_P.n1766 OUT_P.n1765 0.00525899
R19406 OUT_P.n1768 OUT_P.n1767 0.00525899
R19407 OUT_P.n1779 OUT_P.n1778 0.00525899
R19408 OUT_P.n1781 OUT_P.n1780 0.00525899
R19409 OUT_P.n1788 OUT_P.n1787 0.00525899
R19410 OUT_P.n1790 OUT_P.n1789 0.00525899
R19411 OUT_P.n1797 OUT_P.n1796 0.00525899
R19412 OUT_P.n1799 OUT_P.n1798 0.00525899
R19413 OUT_P.n1806 OUT_P.n1805 0.00525899
R19414 OUT_P.n1808 OUT_P.n1807 0.00525899
R19415 OUT_P.n1303 OUT_P.n1302 0.00525899
R19416 OUT_P.n1305 OUT_P.n1304 0.00525899
R19417 OUT_P.n1312 OUT_P.n1311 0.00525899
R19418 OUT_P.n1314 OUT_P.n1313 0.00525899
R19419 OUT_P.n1330 OUT_P.n1329 0.00525899
R19420 OUT_P.n1332 OUT_P.n1331 0.00525899
R19421 OUT_P.n1339 OUT_P.n1338 0.00525899
R19422 OUT_P.n1341 OUT_P.n1340 0.00525899
R19423 OUT_P.n1348 OUT_P.n1347 0.00525899
R19424 OUT_P.n1350 OUT_P.n1349 0.00525899
R19425 OUT_P.n1357 OUT_P.n1356 0.00525899
R19426 OUT_P.n1359 OUT_P.n1358 0.00525899
R19427 OUT_P.n1371 OUT_P.n1370 0.00525899
R19428 OUT_P.n1373 OUT_P.n1372 0.00525899
R19429 OUT_P.n1380 OUT_P.n1379 0.00525899
R19430 OUT_P.n1382 OUT_P.n1381 0.00525899
R19431 OUT_P.n1389 OUT_P.n1388 0.00525899
R19432 OUT_P.n1391 OUT_P.n1390 0.00525899
R19433 OUT_P.n1398 OUT_P.n1397 0.00525899
R19434 OUT_P.n1400 OUT_P.n1399 0.00525899
R19435 OUT_P.n1412 OUT_P.n1411 0.00525899
R19436 OUT_P.n1414 OUT_P.n1413 0.00525899
R19437 OUT_P.n1421 OUT_P.n1420 0.00525899
R19438 OUT_P.n1423 OUT_P.n1422 0.00525899
R19439 OUT_P.n1430 OUT_P.n1429 0.00525899
R19440 OUT_P.n1432 OUT_P.n1431 0.00525899
R19441 OUT_P.n1439 OUT_P.n1438 0.00525899
R19442 OUT_P.n1441 OUT_P.n1440 0.00525899
R19443 OUT_P.n1125 OUT_P.n1124 0.00525899
R19444 OUT_P.n1123 OUT_P.n1122 0.00525899
R19445 OUT_P.n1041 OUT_P.n1040 0.00455
R19446 OUT_P.n1043 OUT_P.n1042 0.00455
R19447 OUT_P.n1044 OUT_P.n1043 0.00455
R19448 OUT_P.n1046 OUT_P.n1045 0.00455
R19449 OUT_P.n1047 OUT_P.n1046 0.00455
R19450 OUT_P.n1052 OUT_P.n1048 0.00455
R19451 OUT_P.n1053 OUT_P.n1052 0.00455
R19452 OUT_P.n1062 OUT_P.n1054 0.00455
R19453 OUT_P.n1072 OUT_P.n1071 0.00455
R19454 OUT_P.n1074 OUT_P.n1073 0.00455
R19455 OUT_P.n1075 OUT_P.n1074 0.00455
R19456 OUT_P.n1077 OUT_P.n1076 0.00455
R19457 OUT_P.n1078 OUT_P.n1077 0.00455
R19458 OUT_P.n1086 OUT_P.n1079 0.00455
R19459 OUT_P.n1087 OUT_P.n1086 0.00455
R19460 OUT_P.n1093 OUT_P.n1088 0.00455
R19461 OUT_P.n1947 OUT_P.n1946 0.00418876
R19462 OUT_P.n1942 OUT_P.n1941 0.00418876
R19463 OUT_P.n565 OUT_P.n564 0.00418876
R19464 OUT_P.n963 OUT_P.n962 0.00418876
R19465 OUT_P.n219 OUT_P.n212 0.00418876
R19466 OUT_P.n230 OUT_P.n223 0.00418876
R19467 OUT_P.n241 OUT_P.n234 0.00418876
R19468 OUT_P.n267 OUT_P.n260 0.00418876
R19469 OUT_P.n278 OUT_P.n271 0.00418876
R19470 OUT_P.n289 OUT_P.n282 0.00418876
R19471 OUT_P.n300 OUT_P.n293 0.00418876
R19472 OUT_P.n311 OUT_P.n304 0.00418876
R19473 OUT_P.n322 OUT_P.n315 0.00418876
R19474 OUT_P.n333 OUT_P.n326 0.00418876
R19475 OUT_P.n344 OUT_P.n337 0.00418876
R19476 OUT_P.n364 OUT_P.n357 0.00418876
R19477 OUT_P.n375 OUT_P.n368 0.00418876
R19478 OUT_P.n386 OUT_P.n379 0.00418876
R19479 OUT_P.n397 OUT_P.n390 0.00418876
R19480 OUT_P.n408 OUT_P.n401 0.00418876
R19481 OUT_P.n419 OUT_P.n412 0.00418876
R19482 OUT_P.n430 OUT_P.n423 0.00418876
R19483 OUT_P.n441 OUT_P.n434 0.00418876
R19484 OUT_P.n456 OUT_P.n449 0.00418876
R19485 OUT_P.n467 OUT_P.n460 0.00418876
R19486 OUT_P.n478 OUT_P.n471 0.00418876
R19487 OUT_P.n489 OUT_P.n482 0.00418876
R19488 OUT_P.n500 OUT_P.n493 0.00418876
R19489 OUT_P.n511 OUT_P.n504 0.00418876
R19490 OUT_P.n522 OUT_P.n515 0.00418876
R19491 OUT_P.n533 OUT_P.n526 0.00418876
R19492 OUT_P.n1822 OUT_P.n1816 0.00418876
R19493 OUT_P.n1833 OUT_P.n1826 0.00418876
R19494 OUT_P.n1844 OUT_P.n1837 0.00418876
R19495 OUT_P.n1853 OUT_P.n1848 0.00418876
R19496 OUT_P.n1863 OUT_P.n1857 0.00418876
R19497 OUT_P.n1874 OUT_P.n1867 0.00418876
R19498 OUT_P.n1885 OUT_P.n1878 0.00418876
R19499 OUT_P.n1894 OUT_P.n1889 0.00418876
R19500 OUT_P.n11 OUT_P.n10 0.00418126
R19501 OUT_P.n76 OUT_P.n75 0.00281899
R19502 OUT_P.n1941 OUT_P.n1940 0.00219433
R19503 OUT_P.n962 OUT_P.n961 0.00219433
R19504 OUT_P.n106 OUT_P.n105 0.00192237
R19505 OUT_P.n552 OUT_P.n551 0.00192237
R19506 OUT_P.n1502 OUT_P.n1501 0.00192237
R19507 OUT_P.n209 OUT_P.n208 0.00192078
R19508 OUT_P.n1063 OUT_P.n1062 0.00180358
R19509 OUT_P.n1094 OUT_P.n1093 0.00180358
R19510 OUT_P.n1071 OUT_P.n1070 0.00180358
R19511 VCM.n2 VCM.t24 43.4933
R19512 VCM.n37 VCM.t27 39.2493
R19513 VCM.n18 VCM.t13 38.9885
R19514 VCM.n24 VCM.t12 38.877
R19515 VCM.n43 VCM.t25 38.6755
R19516 VCM.n1 VCM.t22 37.5555
R19517 VCM.n16 VCM.t0 36.7612
R19518 VCM.n17 VCM.t2 36.7612
R19519 VCM.n29 VCM.t16 36.5005
R19520 VCM.n27 VCM.t18 36.5005
R19521 VCM.n35 VCM.t5 36.5005
R19522 VCM.n36 VCM.t6 36.5005
R19523 VCM.n39 VCM.t17 36.2398
R19524 VCM.n40 VCM.t3 36.2398
R19525 VCM.n21 VCM.t20 35.9791
R19526 VCM.n38 VCM.t29 34.9362
R19527 VCM.n41 VCM.t23 34.9362
R19528 VCM.n22 VCM.t11 34.6755
R19529 VCM.n20 VCM.t9 32.0684
R19530 VCM.n3 VCM.t14 31.938
R19531 VCM.n4 VCM.t1 31.938
R19532 VCM.n19 VCM.t15 31.0255
R19533 VCM.n5 VCM.t19 31.0255
R19534 VCM.n2 VCM.t26 31.0255
R19535 VCM.n4 VCM.n3 20.8576
R19536 VCM.n20 VCM.n19 19.8148
R19537 VCM.n3 VCM.n2 19.8148
R19538 VCM.n5 VCM.n4 19.8148
R19539 VCM.n21 VCM.n20 18.5368
R19540 VCM.n16 VCM.t4 15.9041
R19541 VCM.n17 VCM.t10 15.9041
R19542 VCM.n28 VCM.n27 15.7269
R19543 VCM.n29 VCM.t28 15.6434
R19544 VCM.n27 VCM.t7 15.6434
R19545 VCM.n35 VCM.t8 15.6434
R19546 VCM.n36 VCM.t21 15.6434
R19547 VCM.n40 VCM.n39 14.8868
R19548 VCM.n22 VCM.n21 13.9445
R19549 VCM.n39 VCM.n38 13.9445
R19550 VCM.n41 VCM.n40 13.9445
R19551 VCM.n23 VCM.n16 13.9076
R19552 VCM.n18 VCM.n17 13.9076
R19553 VCM.n42 VCM.n35 13.9076
R19554 VCM.n37 VCM.n36 13.9076
R19555 VCM.n30 VCM.n29 11.2018
R19556 VCM.n45 VCM.n24 5.43841
R19557 VCM.n6 VCM.n5 4.8863
R19558 VCM.n19 VCM.n18 4.62659
R19559 VCM.n38 VCM.n37 4.62659
R19560 VCM.n23 VCM.n22 4.31354
R19561 VCM.n42 VCM.n41 4.31354
R19562 VCM.n44 VCM.n43 3.38239
R19563 VCM.n44 VCM.n34 2.39553
R19564 VCM.n32 VCM.n30 1.50178
R19565 VCM.n55 VCM.n52 1.50106
R19566 VCM.n15 VCM.n14 1.49801
R19567 VCM.n7 VCM.n6 1.49456
R19568 VCM.n45 VCM.n44 1.24481
R19569 VCM.n56 VCM.n47 1.12675
R19570 VCM.n56 VCM.n55 1.126
R19571 VCM.n34 VCM.n33 1.12411
R19572 VCM.n9 VCM.n8 1.12176
R19573 VCM.n43 VCM.n42 0.623652
R19574 VCM.n46 VCM.n45 0.582814
R19575 VCM.n11 VCM.n10 0.582
R19576 VCM.n24 VCM.n23 0.36637
R19577 VCM VCM.n56 0.0998882
R19578 VCM.n30 VCM.n28 0.0301053
R19579 VCM.n33 VCM.n26 0.0206316
R19580 VCM.n10 VCM.n9 0.0156875
R19581 VCM.n7 VCM.n0 0.0152105
R19582 VCM.n55 VCM.n48 0.014
R19583 VCM.n55 VCM.n54 0.014
R19584 VCM.n47 VCM.n46 0.014
R19585 VCM.n51 VCM.n50 0.014
R19586 VCM.n50 VCM.n49 0.0134654
R19587 VCM.n54 VCM.n53 0.0134654
R19588 VCM.n6 VCM.n1 0.0111568
R19589 VCM.n8 VCM.n7 0.00898969
R19590 VCM.n33 VCM.n32 0.00808664
R19591 VCM.n12 VCM.n11 0.00773989
R19592 VCM.n14 VCM.n13 0.00773989
R19593 VCM.n14 VCM.n12 0.00773989
R19594 VCM.n47 VCM.n15 0.00549102
R19595 VCM.n34 VCM.n25 0.00503958
R19596 VCM.n32 VCM.n31 0.00455447
R19597 VCM.n52 VCM.n51 0.00299297
R19598 VBM.n6 VBM.t0 63.68
R19599 VBM.n6 VBM.t2 63.68
R19600 VBM.n24 VBM.n23 6.32241
R19601 VBM.n16 VBM.n15 6.32241
R19602 VBM.n49 VBM.t11 6.32241
R19603 VBM.n46 VBM.n45 6.32241
R19604 VBM.n42 VBM.n41 5.47432
R19605 VBM.n7 VBM.n6 5.14084
R19606 VBM.n32 VBM.n31 4.38115
R19607 VBM.n53 VBM.n52 4.38115
R19608 VBM.n8 VBM.n7 3.74876
R19609 VBM.n25 VBM.n20 3.43224
R19610 VBM.n24 VBM.n22 3.43224
R19611 VBM.n28 VBM.n18 3.43224
R19612 VBM.n16 VBM.n14 3.43224
R19613 VBM.n49 VBM.n48 3.43224
R19614 VBM.n46 VBM.n44 3.43224
R19615 VBM.n27 VBM.n26 2.72313
R19616 VBM.n69 VBM.n68 2.69081
R19617 VBM.n27 VBM.t19 2.56499
R19618 VBM.n26 VBM.t12 2.56298
R19619 VBM.n56 VBM.n42 2.12306
R19620 VBM.n64 VBM.t24 1.6385
R19621 VBM.n64 VBM.n63 1.6385
R19622 VBM.n31 VBM.t25 1.6385
R19623 VBM.n31 VBM.n30 1.6385
R19624 VBM.n20 VBM.t18 1.6385
R19625 VBM.n20 VBM.n19 1.6385
R19626 VBM.n22 VBM.t14 1.6385
R19627 VBM.n22 VBM.n21 1.6385
R19628 VBM.n18 VBM.t21 1.6385
R19629 VBM.n18 VBM.n17 1.6385
R19630 VBM.n14 VBM.t20 1.6385
R19631 VBM.n14 VBM.n13 1.6385
R19632 VBM.n36 VBM.t22 1.6385
R19633 VBM.n36 VBM.n35 1.6385
R19634 VBM.n52 VBM.t23 1.6385
R19635 VBM.n52 VBM.n51 1.6385
R19636 VBM.n48 VBM.t16 1.6385
R19637 VBM.n48 VBM.n47 1.6385
R19638 VBM.n44 VBM.t13 1.6385
R19639 VBM.n44 VBM.n43 1.6385
R19640 VBM.n39 VBM.t15 1.6385
R19641 VBM.n39 VBM.n38 1.6385
R19642 VBM.n41 VBM.t17 1.6385
R19643 VBM.n41 VBM.n40 1.6385
R19644 VBM.n58 VBM.n57 1.50853
R19645 VBM.n67 VBM.n66 1.50128
R19646 VBM.n74 VBM.n3 1.49812
R19647 VBM.n74 VBM.n73 1.49812
R19648 VBM.n62 VBM.n60 1.48107
R19649 VBM.n26 VBM.n25 1.44185
R19650 VBM.n28 VBM.n27 1.43911
R19651 VBM.n37 VBM.n36 1.42054
R19652 VBM.n66 VBM.n65 1.17622
R19653 VBM.n57 VBM.n37 1.15277
R19654 VBM.n56 VBM.n55 1.1255
R19655 VBM.n59 VBM.n34 1.1255
R19656 VBM.n75 VBM.n74 1.1255
R19657 VBM.n65 VBM.n64 1.0626
R19658 VBM.n54 VBM.n53 1.05315
R19659 VBM.n33 VBM.n32 1.03406
R19660 VBM.n42 VBM.n39 0.926316
R19661 VBM.n7 VBM.n5 0.715901
R19662 VBM.n25 VBM.n24 0.626587
R19663 VBM.n5 VBM.t3 0.4555
R19664 VBM.n5 VBM.n4 0.4555
R19665 VBM.n29 VBM.n16 0.323326
R19666 VBM.n50 VBM.n46 0.323326
R19667 VBM.n32 VBM.n29 0.305717
R19668 VBM.n53 VBM.n50 0.305717
R19669 VBM.n29 VBM.n28 0.303761
R19670 VBM.n50 VBM.n49 0.303761
R19671 VBM.n57 VBM.n56 0.123658
R19672 VBM VBM.n75 0.09825
R19673 VBM.n60 VBM.n59 0.0419676
R19674 VBM.n34 VBM.n33 0.0324737
R19675 VBM.n73 VBM.n72 0.0236139
R19676 VBM.n11 VBM.n10 0.0229474
R19677 VBM.n59 VBM.n58 0.0169302
R19678 VBM.n55 VBM.n54 0.014283
R19679 VBM.n74 VBM.n0 0.014
R19680 VBM.n74 VBM.n12 0.014
R19681 VBM.n9 VBM.n8 0.014
R19682 VBM.n2 VBM.n1 0.014
R19683 VBM.n12 VBM.n11 0.0134654
R19684 VBM.n68 VBM.n67 0.0117561
R19685 VBM.n70 VBM.n69 0.00998204
R19686 VBM.n62 VBM.n61 0.00858096
R19687 VBM.n67 VBM.n62 0.00639619
R19688 VBM.n73 VBM.n71 0.00582347
R19689 VBM.n3 VBM.n2 0.00582347
R19690 VBM.n10 VBM.n9 0.00549102
R19691 VBM.n71 VBM.n70 0.00549102
R19692 VCD.n227 VCD.n226 4.27746
R19693 VCD.n227 VCD.n224 3.43224
R19694 VCD.n229 VCD.n228 2.39976
R19695 VCD.n9 VCD.n6 2.24691
R19696 VCD.n22 VCD.n19 2.24691
R19697 VCD.n41 VCD.n38 2.24691
R19698 VCD.n54 VCD.n51 2.24691
R19699 VCD.n69 VCD.n66 2.24691
R19700 VCD.n173 VCD.n172 2.15529
R19701 VCD.n222 VCD.t5 1.6385
R19702 VCD.n222 VCD.n221 1.6385
R19703 VCD.n224 VCD.t53 1.6385
R19704 VCD.n224 VCD.n223 1.6385
R19705 VCD.n226 VCD.t4 1.6385
R19706 VCD.n226 VCD.n225 1.6385
R19707 VCD.n3 VCD.t11 1.6385
R19708 VCD.n3 VCD.n2 1.6385
R19709 VCD.n8 VCD.t17 1.6385
R19710 VCD.n8 VCD.n7 1.6385
R19711 VCD.n6 VCD.t43 1.6385
R19712 VCD.n6 VCD.n5 1.6385
R19713 VCD.n26 VCD.t34 1.6385
R19714 VCD.n26 VCD.n25 1.6385
R19715 VCD.n21 VCD.t48 1.6385
R19716 VCD.n21 VCD.n20 1.6385
R19717 VCD.n19 VCD.t14 1.6385
R19718 VCD.n19 VCD.n18 1.6385
R19719 VCD.n35 VCD.t0 1.6385
R19720 VCD.n35 VCD.n34 1.6385
R19721 VCD.n40 VCD.t39 1.6385
R19722 VCD.n40 VCD.n39 1.6385
R19723 VCD.n38 VCD.t46 1.6385
R19724 VCD.n38 VCD.n37 1.6385
R19725 VCD.n58 VCD.t55 1.6385
R19726 VCD.n58 VCD.n57 1.6385
R19727 VCD.n53 VCD.t13 1.6385
R19728 VCD.n53 VCD.n52 1.6385
R19729 VCD.n51 VCD.t60 1.6385
R19730 VCD.n51 VCD.n50 1.6385
R19731 VCD.n72 VCD.t21 1.6385
R19732 VCD.n72 VCD.n71 1.6385
R19733 VCD.n212 VCD.t61 1.6385
R19734 VCD.n212 VCD.n211 1.6385
R19735 VCD.n135 VCD.t30 1.6385
R19736 VCD.n135 VCD.n134 1.6385
R19737 VCD.n129 VCD.t7 1.6385
R19738 VCD.n129 VCD.n128 1.6385
R19739 VCD.n123 VCD.t22 1.6385
R19740 VCD.n123 VCD.n122 1.6385
R19741 VCD.n200 VCD.t27 1.6385
R19742 VCD.n200 VCD.n199 1.6385
R19743 VCD.n156 VCD.t65 1.6385
R19744 VCD.n156 VCD.n155 1.6385
R19745 VCD.n176 VCD.t63 1.6385
R19746 VCD.n176 VCD.n175 1.6385
R19747 VCD.n172 VCD.t20 1.6385
R19748 VCD.n172 VCD.n171 1.6385
R19749 VCD.n166 VCD.t38 1.6385
R19750 VCD.n166 VCD.n165 1.6385
R19751 VCD.n160 VCD.t10 1.6385
R19752 VCD.n160 VCD.n159 1.6385
R19753 VCD.n117 VCD.t32 1.6385
R19754 VCD.n117 VCD.n116 1.6385
R19755 VCD.n89 VCD.t59 1.6385
R19756 VCD.n89 VCD.n88 1.6385
R19757 VCD.n83 VCD.t41 1.6385
R19758 VCD.n83 VCD.n82 1.6385
R19759 VCD.n77 VCD.t16 1.6385
R19760 VCD.n77 VCD.n76 1.6385
R19761 VCD.n112 VCD.t51 1.6385
R19762 VCD.n112 VCD.n111 1.6385
R19763 VCD.n68 VCD.t57 1.6385
R19764 VCD.n68 VCD.n67 1.6385
R19765 VCD.n66 VCD.t35 1.6385
R19766 VCD.n66 VCD.n65 1.6385
R19767 VCD.n195 VCD.n194 1.49763
R19768 VCD.n9 VCD.n8 1.46669
R19769 VCD.n22 VCD.n21 1.46669
R19770 VCD.n41 VCD.n40 1.46669
R19771 VCD.n54 VCD.n53 1.46669
R19772 VCD.n69 VCD.n68 1.46669
R19773 VCD.n118 VCD.n117 1.46648
R19774 VCD.n74 VCD.n73 1.18861
R19775 VCD.n214 VCD.n213 1.18861
R19776 VCD.n195 VCD.n157 1.1885
R19777 VCD.n114 VCD.n113 1.1885
R19778 VCD.n131 VCD.n130 1.18813
R19779 VCD.n202 VCD.n201 1.18813
R19780 VCD.n178 VCD.n177 1.18813
R19781 VCD.n162 VCD.n161 1.18813
R19782 VCD.n91 VCD.n90 1.18813
R19783 VCD.n79 VCD.n78 1.18813
R19784 VCD.n13 VCD.n4 1.18665
R19785 VCD.n45 VCD.n36 1.18665
R19786 VCD.n137 VCD.n136 1.18665
R19787 VCD.n125 VCD.n124 1.18665
R19788 VCD.n168 VCD.n167 1.18665
R19789 VCD.n85 VCD.n84 1.18665
R19790 VCD.n28 VCD.n27 1.18614
R19791 VCD.n60 VCD.n59 1.18614
R19792 VCD.n46 VCD.n45 1.12572
R19793 VCD.n14 VCD.n13 1.12572
R19794 VCD.n210 VCD.n209 1.10736
R19795 VCD.n228 VCD.n227 1.02906
R19796 VCD VCD.n229 1.01357
R19797 VCD.n228 VCD.n222 0.927451
R19798 VCD.n4 VCD.n3 0.901687
R19799 VCD.n36 VCD.n35 0.901687
R19800 VCD.n73 VCD.n72 0.901687
R19801 VCD.n213 VCD.n212 0.901687
R19802 VCD.n136 VCD.n135 0.901687
R19803 VCD.n124 VCD.n123 0.901687
R19804 VCD.n167 VCD.n166 0.901687
R19805 VCD.n84 VCD.n83 0.901687
R19806 VCD.n157 VCD.n156 0.90147
R19807 VCD.n113 VCD.n112 0.90147
R19808 VCD.n27 VCD.n26 0.90147
R19809 VCD.n59 VCD.n58 0.90147
R19810 VCD.n130 VCD.n129 0.90147
R19811 VCD.n201 VCD.n200 0.90147
R19812 VCD.n177 VCD.n176 0.90147
R19813 VCD.n161 VCD.n160 0.90147
R19814 VCD.n90 VCD.n89 0.90147
R19815 VCD.n78 VCD.n77 0.90147
R19816 VCD.n110 VCD.n108 0.88565
R19817 VCD.n219 VCD.n218 0.874917
R19818 VCD.n184 VCD.n169 0.727104
R19819 VCD.n140 VCD.n138 0.727104
R19820 VCD.n149 VCD.n126 0.727104
R19821 VCD.n98 VCD.n86 0.727104
R19822 VCD.n62 VCD.n61 0.722779
R19823 VCD.n30 VCD.n29 0.722779
R19824 VCD.n10 VCD.n9 0.693301
R19825 VCD.n42 VCD.n41 0.693301
R19826 VCD.n119 VCD.n118 0.68976
R19827 VCD.n118 VCD.n115 0.689663
R19828 VCD.n23 VCD.n22 0.676871
R19829 VCD.n55 VCD.n54 0.676871
R19830 VCD.n70 VCD.n69 0.676871
R19831 VCD.n145 VCD.n132 0.616779
R19832 VCD.n180 VCD.n179 0.616779
R19833 VCD.n189 VCD.n163 0.616779
R19834 VCD.n204 VCD.n203 0.616779
R19835 VCD.n94 VCD.n92 0.616779
R19836 VCD.n103 VCD.n80 0.616779
R19837 VCD.n216 VCD.n215 0.615126
R19838 VCD.n197 VCD.n196 0.598695
R19839 VCD.n229 VCD.n220 0.499954
R19840 VCD.n182 VCD.n181 0.150125
R19841 VCD.n187 VCD.n186 0.150125
R19842 VCD.n191 VCD.n190 0.150125
R19843 VCD.n143 VCD.n142 0.150125
R19844 VCD.n147 VCD.n146 0.150125
R19845 VCD.n152 VCD.n151 0.150125
R19846 VCD.n206 VCD.n205 0.150125
R19847 VCD.n96 VCD.n95 0.150125
R19848 VCD.n101 VCD.n100 0.150125
R19849 VCD.n105 VCD.n104 0.150125
R19850 VCD.n16 VCD.n15 0.149196
R19851 VCD.n32 VCD.n31 0.149196
R19852 VCD.n48 VCD.n47 0.149196
R19853 VCD.n64 VCD.n63 0.149196
R19854 VCD.n114 VCD.n110 0.0995747
R19855 VCD.n214 VCD.n210 0.0929251
R19856 VCD.n13 VCD.n12 0.0832399
R19857 VCD.n45 VCD.n44 0.0832399
R19858 VCD.n195 VCD.n154 0.0831446
R19859 VCD.n138 VCD.n133 0.0823987
R19860 VCD.n126 VCD.n121 0.0823987
R19861 VCD.n169 VCD.n164 0.0823987
R19862 VCD.n86 VCD.n81 0.0823987
R19863 VCD.n218 VCD.n217 0.0754039
R19864 VCD.n163 VCD.n158 0.0712285
R19865 VCD.n179 VCD.n174 0.0712285
R19866 VCD.n203 VCD.n198 0.0712285
R19867 VCD.n132 VCD.n127 0.0712285
R19868 VCD.n80 VCD.n75 0.0712285
R19869 VCD.n92 VCD.n87 0.0712285
R19870 VCD.n61 VCD.n60 0.0623678
R19871 VCD.n29 VCD.n28 0.0623678
R19872 VCD.n29 VCD.n24 0.0620327
R19873 VCD.n61 VCD.n56 0.0620327
R19874 VCD.n179 VCD.n178 0.0534597
R19875 VCD.n163 VCD.n162 0.0534597
R19876 VCD.n132 VCD.n131 0.0534597
R19877 VCD.n203 VCD.n202 0.0534597
R19878 VCD.n92 VCD.n91 0.0534597
R19879 VCD.n80 VCD.n79 0.0534597
R19880 VCD.n218 VCD.n74 0.0500104
R19881 VCD.n154 VCD.n153 0.0420655
R19882 VCD.n12 VCD.n11 0.0419676
R19883 VCD.n44 VCD.n43 0.0419676
R19884 VCD.n169 VCD.n168 0.0415773
R19885 VCD.n126 VCD.n125 0.0415773
R19886 VCD.n138 VCD.n137 0.0415773
R19887 VCD.n86 VCD.n85 0.0415773
R19888 VCD.n24 VCD.n23 0.0324737
R19889 VCD.n56 VCD.n55 0.0324737
R19890 VCD.n174 VCD.n173 0.0324737
R19891 VCD.n196 VCD.n195 0.0324737
R19892 VCD.n198 VCD.n197 0.0324737
R19893 VCD.n115 VCD.n114 0.0324737
R19894 VCD.n120 VCD.n119 0.0324737
R19895 VCD.n215 VCD.n214 0.0324737
R19896 VCD.n74 VCD.n70 0.0324737
R19897 VCD.n210 VCD.n120 0.0320039
R19898 VCD.n110 VCD.n109 0.0261793
R19899 VCD.n217 VCD.n216 0.0169302
R19900 VCD.n43 VCD.n42 0.0169302
R19901 VCD.n11 VCD.n10 0.0169302
R19902 VCD.n180 VCD.n170 0.0156875
R19903 VCD.n181 VCD.n180 0.0156875
R19904 VCD.n190 VCD.n189 0.0156875
R19905 VCD.n146 VCD.n145 0.0156875
R19906 VCD.n204 VCD.n152 0.0156875
R19907 VCD.n205 VCD.n204 0.0156875
R19908 VCD.n209 VCD.n208 0.0156875
R19909 VCD.n95 VCD.n94 0.0156875
R19910 VCD.n104 VCD.n103 0.0156875
R19911 VCD.n108 VCD.n107 0.0156875
R19912 VCD.n1 VCD.n0 0.0155932
R19913 VCD.n31 VCD.n30 0.0155932
R19914 VCD.n33 VCD.n32 0.0155932
R19915 VCD.n63 VCD.n62 0.0155932
R19916 VCD.n219 VCD.n64 0.0155932
R19917 VCD.n220 VCD.n219 0.0155932
R19918 VCD.n47 VCD.n46 0.012283
R19919 VCD.n15 VCD.n14 0.012283
R19920 VCD.n192 VCD.n191 0.0111023
R19921 VCD.n106 VCD.n105 0.0111023
R19922 VCD.n207 VCD.n206 0.0111023
R19923 VCD.n141 VCD.n140 0.00860784
R19924 VCD.n145 VCD.n144 0.00860784
R19925 VCD.n150 VCD.n149 0.00860784
R19926 VCD.n185 VCD.n184 0.00860784
R19927 VCD.n189 VCD.n188 0.00860784
R19928 VCD.n94 VCD.n93 0.00860784
R19929 VCD.n99 VCD.n98 0.00860784
R19930 VCD.n103 VCD.n102 0.00860784
R19931 VCD.n183 VCD.n182 0.00858096
R19932 VCD.n184 VCD.n183 0.00858096
R19933 VCD.n148 VCD.n147 0.00858096
R19934 VCD.n149 VCD.n148 0.00858096
R19935 VCD.n140 VCD.n139 0.00858096
R19936 VCD.n97 VCD.n96 0.00858096
R19937 VCD.n98 VCD.n97 0.00858096
R19938 VCD.n30 VCD.n17 0.00856066
R19939 VCD.n62 VCD.n49 0.00856066
R19940 VCD.n186 VCD.n185 0.00855417
R19941 VCD.n188 VCD.n187 0.00855417
R19942 VCD.n142 VCD.n141 0.00855417
R19943 VCD.n144 VCD.n143 0.00855417
R19944 VCD.n151 VCD.n150 0.00855417
R19945 VCD.n100 VCD.n99 0.00855417
R19946 VCD.n102 VCD.n101 0.00855417
R19947 VCD.n17 VCD.n16 0.00850732
R19948 VCD.n49 VCD.n48 0.00850732
R19949 VCD.n193 VCD.n192 0.00605114
R19950 VCD.n194 VCD.n193 0.00605114
R19951 VCD.n209 VCD.n207 0.00605114
R19952 VCD.n108 VCD.n106 0.00605114
R19953 VCD.n14 VCD.n1 0.00477236
R19954 VCD.n46 VCD.n33 0.00477236
R19955 IN_N.t6 IN_N.t14 147.304
R19956 IN_N.t8 IN_N.t19 147.304
R19957 IN_N.t0 IN_N.t11 147.304
R19958 IN_N.t22 IN_N.t13 147.304
R19959 IN_N.n13 IN_N.t4 75.2545
R19960 IN_N.n24 IN_N.t23 75.1498
R19961 IN_N.n43 IN_N.t0 75.0919
R19962 IN_N.n30 IN_N.t15 73.4037
R19963 IN_N.n49 IN_N.t22 73.3458
R19964 IN_N.n14 IN_N.t3 72.8823
R19965 IN_N.n46 IN_N.t7 72.3487
R19966 IN_N.n44 IN_N.t8 72.3487
R19967 IN_N.n42 IN_N.t20 72.3487
R19968 IN_N.n27 IN_N.t10 72.3487
R19969 IN_N.n25 IN_N.t5 72.3487
R19970 IN_N.n23 IN_N.t21 72.3487
R19971 IN_N.n12 IN_N.t18 72.3487
R19972 IN_N.n46 IN_N.t9 51.4916
R19973 IN_N.n44 IN_N.t6 51.4916
R19974 IN_N.n42 IN_N.t1 51.4916
R19975 IN_N.n27 IN_N.t12 51.4916
R19976 IN_N.n25 IN_N.t17 51.4916
R19977 IN_N.n23 IN_N.t2 51.4916
R19978 IN_N.n12 IN_N.t16 51.4916
R19979 IN_N.n47 IN_N.n46 19.9041
R19980 IN_N.n43 IN_N.n42 19.9041
R19981 IN_N.n28 IN_N.n27 19.9041
R19982 IN_N.n24 IN_N.n23 19.9041
R19983 IN_N.n45 IN_N.n44 15.6747
R19984 IN_N.n26 IN_N.n25 15.6747
R19985 IN_N.n13 IN_N.n12 15.2112
R19986 IN_N.n57 IN_N.n38 2.82762
R19987 IN_N.n50 IN_N.n49 1.5005
R19988 IN_N.n9 IN_N.n3 1.49812
R19989 IN_N.n9 IN_N.n8 1.49812
R19990 IN_N.n59 IN_N.n21 1.49801
R19991 IN_N.n58 IN_N.n57 1.21977
R19992 IN_N.n18 IN_N.n17 1.14692
R19993 IN_N.n60 IN_N.n59 1.12675
R19994 IN_N.n60 IN_N.n9 1.126
R19995 IN_N.n16 IN_N.n15 1.12272
R19996 IN_N.n54 IN_N.n53 1.1073
R19997 IN_N.n36 IN_N.n35 1.1073
R19998 IN_N.n57 IN_N.n56 0.933295
R19999 IN_N.n15 IN_N.n13 0.90419
R20000 IN_N.n31 IN_N.n30 0.897484
R20001 IN_N.n45 IN_N.n43 0.626587
R20002 IN_N.n47 IN_N.n45 0.626587
R20003 IN_N.n26 IN_N.n24 0.626587
R20004 IN_N.n28 IN_N.n26 0.626587
R20005 IN_N.n20 IN_N.n19 0.366019
R20006 IN_N.n49 IN_N.n47 0.239196
R20007 IN_N.n30 IN_N.n28 0.239196
R20008 IN_N IN_N.n60 0.112826
R20009 IN_N.n35 IN_N.n33 0.0649899
R20010 IN_N.n53 IN_N.n51 0.0638057
R20011 IN_N.n53 IN_N.n52 0.032498
R20012 IN_N.n35 IN_N.n34 0.032498
R20013 IN_N.n16 IN_N.n11 0.0301053
R20014 IN_N.n30 IN_N.n29 0.0289211
R20015 IN_N.n33 IN_N.n32 0.0289211
R20016 IN_N.n49 IN_N.n48 0.0277368
R20017 IN_N.n51 IN_N.n50 0.0277368
R20018 IN_N.n8 IN_N.n7 0.0236139
R20019 IN_N.n17 IN_N.n16 0.0220754
R20020 IN_N.n41 IN_N.n40 0.0151213
R20021 IN_N.n9 IN_N.n0 0.014
R20022 IN_N.n9 IN_N.n5 0.014
R20023 IN_N.n59 IN_N.n58 0.014
R20024 IN_N.n2 IN_N.n1 0.014
R20025 IN_N.n5 IN_N.n4 0.0134654
R20026 IN_N.n56 IN_N.n55 0.0111023
R20027 IN_N.n38 IN_N.n37 0.0111023
R20028 IN_N.n21 IN_N.n20 0.00998204
R20029 IN_N.n54 IN_N.n39 0.00860784
R20030 IN_N.n36 IN_N.n22 0.00860784
R20031 IN_N.n15 IN_N.n14 0.00845754
R20032 IN_N.n32 IN_N.n31 0.00685938
R20033 IN_N.n19 IN_N.n18 0.00638348
R20034 IN_N.n55 IN_N.n54 0.00605114
R20035 IN_N.n37 IN_N.n36 0.00605114
R20036 IN_N.n8 IN_N.n6 0.00582347
R20037 IN_N.n3 IN_N.n2 0.00582347
R20038 IN_N.n59 IN_N.n10 0.00549102
R20039 IN_N.n50 IN_N.n41 0.00286842
R20040 BD.n106 BD.n105 4.81137
R20041 BD.n111 BD.n110 4.81137
R20042 BD.n116 BD.n115 4.81137
R20043 BD.n179 BD.n178 4.09137
R20044 BD.n168 BD.n167 4.09137
R20045 BD.n157 BD.n156 4.09137
R20046 BD.n195 BD.n194 4.04637
R20047 BD.n79 BD.n78 4.04637
R20048 BD.n43 BD.n42 4.04637
R20049 BD.n24 BD.n23 4.04637
R20050 BD.n196 BD.n190 3.42028
R20051 BD.n195 BD.n192 3.42028
R20052 BD.n80 BD.n74 3.42028
R20053 BD.n79 BD.n76 3.42028
R20054 BD.n44 BD.n38 3.42028
R20055 BD.n43 BD.n40 3.42028
R20056 BD.n25 BD.n19 3.42028
R20057 BD.n24 BD.n21 3.42028
R20058 BD.n179 BD.n176 2.6005
R20059 BD.n180 BD.n174 2.6005
R20060 BD.n181 BD.n172 2.6005
R20061 BD.n168 BD.n165 2.6005
R20062 BD.n169 BD.n163 2.6005
R20063 BD.n170 BD.n161 2.6005
R20064 BD.n157 BD.n154 2.6005
R20065 BD.n158 BD.n152 2.6005
R20066 BD.n159 BD.n150 2.6005
R20067 BD.n68 BD.n36 2.6005
R20068 BD.n106 BD.n103 2.6005
R20069 BD.n111 BD.n108 2.6005
R20070 BD.n116 BD.n113 2.6005
R20071 BD.n121 BD.n120 2.6005
R20072 BD.n122 BD.n121 1.79659
R20073 BD.n148 BD.n147 1.64287
R20074 BD.n182 BD.n181 1.5442
R20075 BD.n72 BD.n34 1.54399
R20076 BD.n16 BD.n15 1.50472
R20077 BD.n29 BD.n28 1.50128
R20078 BD.n138 BD.n136 1.49812
R20079 BD.n9 BD.n3 1.49812
R20080 BD.n9 BD.n8 1.49812
R20081 BD.n145 BD.n144 1.49801
R20082 BD.n210 BD.n32 1.49801
R20083 BD.n181 BD.n180 1.49137
R20084 BD.n180 BD.n179 1.49137
R20085 BD.n170 BD.n169 1.49137
R20086 BD.n169 BD.n168 1.49137
R20087 BD.n159 BD.n158 1.49137
R20088 BD.n158 BD.n157 1.49137
R20089 BD.n17 BD.n11 1.48107
R20090 BD.n117 BD.n116 1.44637
R20091 BD.n121 BD.n118 1.44637
R20092 BD.n208 BD.n188 1.36943
R20093 BD.n208 BD.n207 1.33886
R20094 BD.n184 BD.n183 1.28649
R20095 BD.n65 BD.n64 1.26677
R20096 BD.n128 BD.n127 1.17988
R20097 BD.n51 BD.n50 1.16583
R20098 BD.n203 BD.n202 1.1658
R20099 BD.n87 BD.n86 1.1658
R20100 BD.n15 BD.n14 1.1658
R20101 BD.n211 BD.n210 1.12675
R20102 BD.n211 BD.n9 1.126
R20103 BD.n199 BD.n198 1.1255
R20104 BD.n83 BD.n82 1.1255
R20105 BD.n47 BD.n46 1.1255
R20106 BD.n66 BD.n62 1.1255
R20107 BD.n98 BD.n97 1.1255
R20108 BD.n71 BD.n70 1.1255
R20109 BD.n124 BD.n123 1.1255
R20110 BD.n28 BD.n27 1.1255
R20111 BD.n68 BD.n67 1.11357
R20112 BD.n96 BD.n95 1.10736
R20113 BD.n61 BD.n59 1.10736
R20114 BD.n69 BD.n68 1.01985
R20115 BD.n202 BD.n201 1.00677
R20116 BD.n86 BD.n85 1.00677
R20117 BD.n14 BD.n13 1.00677
R20118 BD.n100 BD.n99 0.984698
R20119 BD.n45 BD.n44 0.968978
R20120 BD.n50 BD.n49 0.966825
R20121 BD.n127 BD.n126 0.963628
R20122 BD.n183 BD.n182 0.845717
R20123 BD.n118 BD.n106 0.820283
R20124 BD.n117 BD.n111 0.820283
R20125 BD.n197 BD.n196 0.773326
R20126 BD.n81 BD.n80 0.773326
R20127 BD.n26 BD.n25 0.773326
R20128 BD.n92 BD.n91 0.761
R20129 BD.n56 BD.n55 0.761
R20130 BD.n133 BD.n132 0.760312
R20131 BD.n31 BD.n30 0.760312
R20132 BD.n186 BD.n185 0.7505
R20133 BD.n138 BD.n101 0.7505
R20134 BD.n182 BD.n170 0.698978
R20135 BD.n183 BD.n159 0.698978
R20136 BD.n196 BD.n195 0.626587
R20137 BD.n80 BD.n79 0.626587
R20138 BD.n44 BD.n43 0.626587
R20139 BD.n118 BD.n117 0.626587
R20140 BD.n25 BD.n24 0.626587
R20141 BD.n206 BD.n204 0.616779
R20142 BD.n90 BD.n88 0.616779
R20143 BD.n54 BD.n52 0.616779
R20144 BD.n131 BD.n129 0.616779
R20145 BD.n209 BD.n208 0.585272
R20146 BD.n172 BD.t7 0.58197
R20147 BD.n172 BD.n171 0.58197
R20148 BD.n174 BD.t69 0.58197
R20149 BD.n174 BD.n173 0.58197
R20150 BD.n176 BD.t70 0.58197
R20151 BD.n176 BD.n175 0.58197
R20152 BD.n178 BD.t3 0.58197
R20153 BD.n178 BD.n177 0.58197
R20154 BD.n161 BD.t79 0.58197
R20155 BD.n161 BD.n160 0.58197
R20156 BD.n163 BD.t75 0.58197
R20157 BD.n163 BD.n162 0.58197
R20158 BD.n165 BD.t5 0.58197
R20159 BD.n165 BD.n164 0.58197
R20160 BD.n167 BD.t68 0.58197
R20161 BD.n167 BD.n166 0.58197
R20162 BD.n150 BD.t4 0.58197
R20163 BD.n150 BD.n149 0.58197
R20164 BD.n152 BD.t65 0.58197
R20165 BD.n152 BD.n151 0.58197
R20166 BD.n154 BD.t9 0.58197
R20167 BD.n154 BD.n153 0.58197
R20168 BD.n156 BD.t0 0.58197
R20169 BD.n156 BD.n155 0.58197
R20170 BD.n147 BD.t11 0.58197
R20171 BD.n147 BD.n146 0.58197
R20172 BD.n34 BD.t73 0.58197
R20173 BD.n34 BD.n33 0.58197
R20174 BD.n36 BD.t66 0.58197
R20175 BD.n36 BD.n35 0.58197
R20176 BD.n64 BD.t2 0.58197
R20177 BD.n64 BD.n63 0.58197
R20178 BD.n190 BD.t26 0.485833
R20179 BD.n190 BD.n189 0.485833
R20180 BD.n192 BD.t57 0.485833
R20181 BD.n192 BD.n191 0.485833
R20182 BD.n194 BD.t24 0.485833
R20183 BD.n194 BD.n193 0.485833
R20184 BD.n201 BD.t49 0.485833
R20185 BD.n201 BD.n200 0.485833
R20186 BD.n74 BD.t20 0.485833
R20187 BD.n74 BD.n73 0.485833
R20188 BD.n76 BD.t56 0.485833
R20189 BD.n76 BD.n75 0.485833
R20190 BD.n78 BD.t34 0.485833
R20191 BD.n78 BD.n77 0.485833
R20192 BD.n85 BD.t46 0.485833
R20193 BD.n85 BD.n84 0.485833
R20194 BD.n38 BD.t41 0.485833
R20195 BD.n38 BD.n37 0.485833
R20196 BD.n40 BD.t23 0.485833
R20197 BD.n40 BD.n39 0.485833
R20198 BD.n42 BD.t35 0.485833
R20199 BD.n42 BD.n41 0.485833
R20200 BD.n49 BD.t60 0.485833
R20201 BD.n49 BD.n48 0.485833
R20202 BD.n120 BD.t17 0.485833
R20203 BD.n120 BD.n119 0.485833
R20204 BD.n103 BD.t52 0.485833
R20205 BD.n103 BD.n102 0.485833
R20206 BD.n105 BD.t44 0.485833
R20207 BD.n105 BD.n104 0.485833
R20208 BD.n108 BD.t59 0.485833
R20209 BD.n108 BD.n107 0.485833
R20210 BD.n110 BD.t29 0.485833
R20211 BD.n110 BD.n109 0.485833
R20212 BD.n113 BD.t58 0.485833
R20213 BD.n113 BD.n112 0.485833
R20214 BD.n115 BD.t47 0.485833
R20215 BD.n115 BD.n114 0.485833
R20216 BD.n126 BD.t21 0.485833
R20217 BD.n126 BD.n125 0.485833
R20218 BD.n19 BD.t42 0.485833
R20219 BD.n19 BD.n18 0.485833
R20220 BD.n21 BD.t16 0.485833
R20221 BD.n21 BD.n20 0.485833
R20222 BD.n23 BD.t54 0.485833
R20223 BD.n23 BD.n22 0.485833
R20224 BD.n13 BD.t31 0.485833
R20225 BD.n13 BD.n12 0.485833
R20226 BD.n123 BD.n122 0.3155
R20227 BD.n46 BD.n45 0.252891
R20228 BD.n101 BD.n100 0.213196
R20229 BD.n99 BD.n98 0.204046
R20230 BD.n71 BD.n69 0.137457
R20231 BD.n66 BD.n65 0.109357
R20232 BD.n185 BD.n184 0.097556
R20233 BD.n61 BD.n60 0.0929251
R20234 BD BD.n211 0.0903257
R20235 BD.n204 BD.n199 0.0712285
R20236 BD.n88 BD.n83 0.0712285
R20237 BD.n52 BD.n47 0.0712285
R20238 BD.n129 BD.n124 0.0712285
R20239 BD.n67 BD.n66 0.0698213
R20240 BD.n72 BD.n71 0.0624212
R20241 BD.n98 BD.n72 0.0620608
R20242 BD.n198 BD.n197 0.0572391
R20243 BD.n82 BD.n81 0.0572391
R20244 BD.n27 BD.n26 0.0572391
R20245 BD.n204 BD.n203 0.0534597
R20246 BD.n88 BD.n87 0.0534597
R20247 BD.n52 BD.n51 0.0534597
R20248 BD.n129 BD.n128 0.0534597
R20249 BD.n185 BD.n148 0.0364864
R20250 BD.n97 BD.n96 0.0320039
R20251 BD.n62 BD.n61 0.0320039
R20252 BD.n8 BD.n7 0.0236139
R20253 BD.n142 BD.n141 0.0229474
R20254 BD.n145 BD.n140 0.0229474
R20255 BD.n207 BD.n206 0.0156875
R20256 BD.n91 BD.n90 0.0156875
R20257 BD.n55 BD.n54 0.0156875
R20258 BD.n132 BD.n131 0.0156875
R20259 BD.n144 BD.n143 0.014
R20260 BD.n139 BD.n138 0.014
R20261 BD.n138 BD.n137 0.014
R20262 BD.n9 BD.n0 0.014
R20263 BD.n9 BD.n5 0.014
R20264 BD.n210 BD.n209 0.014
R20265 BD.n2 BD.n1 0.014
R20266 BD.n140 BD.n139 0.0134654
R20267 BD.n5 BD.n4 0.0134654
R20268 BD.n30 BD.n29 0.0117561
R20269 BD.n93 BD.n92 0.0111023
R20270 BD.n57 BD.n56 0.0111023
R20271 BD.n32 BD.n31 0.00998204
R20272 BD.n206 BD.n205 0.00860784
R20273 BD.n90 BD.n89 0.00860784
R20274 BD.n54 BD.n53 0.00860784
R20275 BD.n131 BD.n130 0.00860784
R20276 BD.n135 BD.n134 0.00773989
R20277 BD.n188 BD.n187 0.00773989
R20278 BD.n134 BD.n133 0.00773989
R20279 BD.n187 BD.n186 0.00773989
R20280 BD.n29 BD.n17 0.00639619
R20281 BD.n95 BD.n93 0.00605114
R20282 BD.n59 BD.n57 0.00605114
R20283 BD.n136 BD.n135 0.00582347
R20284 BD.n8 BD.n6 0.00582347
R20285 BD.n3 BD.n2 0.00582347
R20286 BD.n144 BD.n142 0.00549102
R20287 BD.n186 BD.n145 0.00549102
R20288 BD.n210 BD.n10 0.00549102
R20289 BD.n95 BD.n94 0.005061
R20290 BD.n59 BD.n58 0.005061
R20291 BD.n17 BD.n16 0.0039419
R20292 IBIAS3.t80 IBIAS3.t40 95.9434
R20293 IBIAS3.t79 IBIAS3.t80 95.9434
R20294 IBIAS3.t73 IBIAS3.t79 95.9434
R20295 IBIAS3.t66 IBIAS3.t24 95.9434
R20296 IBIAS3.t65 IBIAS3.t66 95.9434
R20297 IBIAS3.t60 IBIAS3.t65 95.9434
R20298 IBIAS3.t36 IBIAS3.t52 95.9434
R20299 IBIAS3.t35 IBIAS3.t36 95.9434
R20300 IBIAS3.t29 IBIAS3.t35 95.9434
R20301 IBIAS3.t72 IBIAS3.t33 95.9434
R20302 IBIAS3.t70 IBIAS3.t72 95.9434
R20303 IBIAS3.t68 IBIAS3.t70 95.9434
R20304 IBIAS3.t43 IBIAS3.t56 95.9434
R20305 IBIAS3.t42 IBIAS3.t43 95.9434
R20306 IBIAS3.t39 IBIAS3.t42 95.9434
R20307 IBIAS3.t28 IBIAS3.t46 95.9434
R20308 IBIAS3.t26 IBIAS3.t28 95.9434
R20309 IBIAS3.t23 IBIAS3.t26 95.9434
R20310 IBIAS3.t76 IBIAS3.t37 95.9434
R20311 IBIAS3.t74 IBIAS3.t76 95.9434
R20312 IBIAS3.t69 IBIAS3.t74 95.9434
R20313 IBIAS3.t45 IBIAS3.t58 95.9434
R20314 IBIAS3.t44 IBIAS3.t45 95.9434
R20315 IBIAS3.t41 IBIAS3.t44 95.9434
R20316 IBIAS3.t31 IBIAS3.t48 95.9434
R20317 IBIAS3.t30 IBIAS3.t31 95.9434
R20318 IBIAS3.t25 IBIAS3.t30 95.9434
R20319 IBIAS3.t55 IBIAS3.t75 95.9434
R20320 IBIAS3.t54 IBIAS3.t55 95.9434
R20321 IBIAS3.t53 IBIAS3.t54 95.9434
R20322 IBIAS3.t62 IBIAS3.t21 95.9434
R20323 IBIAS3.t61 IBIAS3.t62 95.9434
R20324 IBIAS3.t57 IBIAS3.t61 95.9434
R20325 IBIAS3.t51 IBIAS3.t67 95.9434
R20326 IBIAS3.t49 IBIAS3.t51 95.9434
R20327 IBIAS3.t47 IBIAS3.t49 95.9434
R20328 IBIAS3.t78 IBIAS3.t38 95.9434
R20329 IBIAS3.t77 IBIAS3.t78 95.9434
R20330 IBIAS3.t71 IBIAS3.t77 95.9434
R20331 IBIAS3.t64 IBIAS3.t22 95.9434
R20332 IBIAS3.t63 IBIAS3.t64 95.9434
R20333 IBIAS3.t59 IBIAS3.t63 95.9434
R20334 IBIAS3.t15 IBIAS3.t11 95.9434
R20335 IBIAS3.t17 IBIAS3.t15 95.9434
R20336 IBIAS3.t19 IBIAS3.t17 95.9434
R20337 IBIAS3.t5 IBIAS3.t13 95.9434
R20338 IBIAS3.t7 IBIAS3.t5 95.9434
R20339 IBIAS3.t9 IBIAS3.t7 95.9434
R20340 IBIAS3.n14 IBIAS3.t73 65.3674
R20341 IBIAS3.n37 IBIAS3.t9 57.2563
R20342 IBIAS3.n14 IBIAS3.t60 49.1451
R20343 IBIAS3.n15 IBIAS3.t29 49.1451
R20344 IBIAS3.n16 IBIAS3.t68 49.1451
R20345 IBIAS3.n17 IBIAS3.t39 49.1451
R20346 IBIAS3.n18 IBIAS3.t23 49.1451
R20347 IBIAS3.n19 IBIAS3.t69 49.1451
R20348 IBIAS3.n20 IBIAS3.t41 49.1451
R20349 IBIAS3.n21 IBIAS3.t25 49.1451
R20350 IBIAS3.n22 IBIAS3.t53 49.1451
R20351 IBIAS3.n23 IBIAS3.t57 49.1451
R20352 IBIAS3.n41 IBIAS3.t47 49.1451
R20353 IBIAS3.n40 IBIAS3.t71 49.1451
R20354 IBIAS3.n39 IBIAS3.t59 49.1451
R20355 IBIAS3.n38 IBIAS3.t19 49.1451
R20356 IBIAS3.n39 IBIAS3.n38 16.2227
R20357 IBIAS3.n40 IBIAS3.n39 16.2227
R20358 IBIAS3.n41 IBIAS3.n40 16.2227
R20359 IBIAS3.n23 IBIAS3.n22 16.2227
R20360 IBIAS3.n22 IBIAS3.n21 16.2227
R20361 IBIAS3.n21 IBIAS3.n20 16.2227
R20362 IBIAS3.n20 IBIAS3.n19 16.2227
R20363 IBIAS3.n19 IBIAS3.n18 16.2227
R20364 IBIAS3.n18 IBIAS3.n17 16.2227
R20365 IBIAS3.n17 IBIAS3.n16 16.2227
R20366 IBIAS3.n16 IBIAS3.n15 16.2227
R20367 IBIAS3.n15 IBIAS3.n14 16.2227
R20368 IBIAS3.n38 IBIAS3.n37 8.11161
R20369 IBIAS3.n4 IBIAS3.t0 5.63646
R20370 IBIAS3.n4 IBIAS3.n3 4.81746
R20371 IBIAS3.n37 IBIAS3.n36 4.80854
R20372 IBIAS3.n34 IBIAS3.n33 4.0405
R20373 IBIAS3.n42 IBIAS3.n41 2.94078
R20374 IBIAS3.n43 IBIAS3.n42 2.8805
R20375 IBIAS3.n25 IBIAS3.n24 2.8805
R20376 IBIAS3.n24 IBIAS3.n23 2.738
R20377 IBIAS3.n34 IBIAS3.n31 2.6005
R20378 IBIAS3.n35 IBIAS3.n29 2.6005
R20379 IBIAS3.n36 IBIAS3.n27 2.6005
R20380 IBIAS3.n55 IBIAS3.n52 1.52353
R20381 IBIAS3.n36 IBIAS3.n35 1.4405
R20382 IBIAS3.n35 IBIAS3.n34 1.4405
R20383 IBIAS3.n66 IBIAS3.n65 1.28809
R20384 IBIAS3.n72 IBIAS3.n71 1.14402
R20385 IBIAS3.n56 IBIAS3.n8 1.13468
R20386 IBIAS3.n68 IBIAS3.n67 1.1255
R20387 IBIAS3.n61 IBIAS3.n6 1.1255
R20388 IBIAS3.n52 IBIAS3.n51 1.11801
R20389 IBIAS3.n56 IBIAS3.n55 1.11782
R20390 IBIAS3.n84 IBIAS3.n83 1.11782
R20391 IBIAS3.n65 IBIAS3.t4 0.8195
R20392 IBIAS3.n65 IBIAS3.n64 0.8195
R20393 IBIAS3.n3 IBIAS3.t3 0.8195
R20394 IBIAS3.n3 IBIAS3.n2 0.8195
R20395 IBIAS3.n27 IBIAS3.t10 0.607167
R20396 IBIAS3.n27 IBIAS3.n26 0.607167
R20397 IBIAS3.n29 IBIAS3.t8 0.607167
R20398 IBIAS3.n29 IBIAS3.n28 0.607167
R20399 IBIAS3.n31 IBIAS3.t6 0.607167
R20400 IBIAS3.n31 IBIAS3.n30 0.607167
R20401 IBIAS3.n33 IBIAS3.t14 0.607167
R20402 IBIAS3.n33 IBIAS3.n32 0.607167
R20403 IBIAS3.n83 IBIAS3.n78 0.574897
R20404 IBIAS3.n47 IBIAS3.n46 0.549056
R20405 IBIAS3.n45 IBIAS3.n44 0.5355
R20406 IBIAS3.n78 IBIAS3.n77 0.508819
R20407 IBIAS3.n5 IBIAS3.n4 0.211804
R20408 IBIAS3.n60 IBIAS3.n59 0.209193
R20409 IBIAS3.n6 IBIAS3.n5 0.121804
R20410 IBIAS3 IBIAS3.n85 0.0917676
R20411 IBIAS3.n44 IBIAS3.n43 0.062564
R20412 IBIAS3.n44 IBIAS3.n25 0.0620381
R20413 IBIAS3.n67 IBIAS3.n66 0.061035
R20414 IBIAS3.n12 IBIAS3.n11 0.0235313
R20415 IBIAS3.n1 IBIAS3.n0 0.0235313
R20416 IBIAS3.n49 IBIAS3.n48 0.0228651
R20417 IBIAS3.n54 IBIAS3.n53 0.0228651
R20418 IBIAS3.n59 IBIAS3.n58 0.0228651
R20419 IBIAS3.n80 IBIAS3.n79 0.0228651
R20420 IBIAS3.n51 IBIAS3.n47 0.0179841
R20421 IBIAS3.n83 IBIAS3.n82 0.0179841
R20422 IBIAS3.n51 IBIAS3.n50 0.0177304
R20423 IBIAS3.n82 IBIAS3.n81 0.0177304
R20424 IBIAS3.n10 IBIAS3.n9 0.0173591
R20425 IBIAS3.n11 IBIAS3.n10 0.0173591
R20426 IBIAS3.n57 IBIAS3.n56 0.0173591
R20427 IBIAS3.n8 IBIAS3.n7 0.0173591
R20428 IBIAS3.n85 IBIAS3.n84 0.0173591
R20429 IBIAS3.n84 IBIAS3.n1 0.0173591
R20430 IBIAS3.n74 IBIAS3.n73 0.0163451
R20431 IBIAS3.n77 IBIAS3.n76 0.0163451
R20432 IBIAS3.n63 IBIAS3.n62 0.0163451
R20433 IBIAS3.n70 IBIAS3.n69 0.0163451
R20434 IBIAS3.n52 IBIAS3.n12 0.0122638
R20435 IBIAS3.n50 IBIAS3.n49 0.0119325
R20436 IBIAS3.n55 IBIAS3.n54 0.0119325
R20437 IBIAS3.n58 IBIAS3.n57 0.0119325
R20438 IBIAS3.n81 IBIAS3.n80 0.0119325
R20439 IBIAS3.n75 IBIAS3.n74 0.00905634
R20440 IBIAS3.n76 IBIAS3.n75 0.00905634
R20441 IBIAS3.n62 IBIAS3.n61 0.00905634
R20442 IBIAS3.n68 IBIAS3.n63 0.00905634
R20443 IBIAS3.n69 IBIAS3.n68 0.00905634
R20444 IBIAS3.n72 IBIAS3.n70 0.00905634
R20445 IBIAS3.n46 IBIAS3.n45 0.00842254
R20446 IBIAS3.n45 IBIAS3.n13 0.00810563
R20447 IBIAS3.n61 IBIAS3.n60 0.0019475
R20448 IBIAS3.n78 IBIAS3.n72 0.0019475
R20449 IVS.t77 IVS.t82 19.5645
R20450 IVS.t88 IVS.t78 19.5645
R20451 IVS.t81 IVS.t86 19.5645
R20452 IVS.t89 IVS.t79 19.5645
R20453 IVS.t84 IVS.t91 19.5645
R20454 IVS.t68 IVS.t62 19.5645
R20455 IVS.t58 IVS.t70 19.5645
R20456 IVS.t64 IVS.t56 19.5645
R20457 IVS.t74 IVS.t66 19.5645
R20458 IVS.t60 IVS.t72 19.5645
R20459 IVS.n211 IVS.t60 13.4946
R20460 IVS.n229 IVS.n228 11.0965
R20461 IVS.n228 IVS.n227 11.0965
R20462 IVS.n227 IVS.n226 11.0965
R20463 IVS.n221 IVS.n220 11.0965
R20464 IVS.n213 IVS.n212 11.0965
R20465 IVS.n240 IVS.t77 10.987
R20466 IVS.n229 IVS.t88 9.4905
R20467 IVS.n228 IVS.t81 9.4905
R20468 IVS.n227 IVS.t89 9.4905
R20469 IVS.n226 IVS.t84 9.4905
R20470 IVS.n221 IVS.t68 9.4905
R20471 IVS.n220 IVS.t58 9.4905
R20472 IVS.n213 IVS.t64 9.4905
R20473 IVS.n212 IVS.t74 9.4905
R20474 IVS.n226 IVS.n225 8.67515
R20475 IVS.n224 IVS.n222 5.0182
R20476 IVS.n218 IVS.n215 4.1992
R20477 IVS.n210 IVS.n207 4.1992
R20478 IVS.n175 IVS.n172 4.0405
R20479 IVS.n75 IVS.n72 4.0405
R20480 IVS.n106 IVS.n103 4.0405
R20481 IVS.n52 IVS.n49 4.0405
R20482 IVS.n29 IVS.n26 4.0405
R20483 IVS.n150 IVS.n147 4.0405
R20484 IVS.n4 IVS.n1 4.0405
R20485 IVS.n225 IVS.n221 4.00459
R20486 IVS.n219 IVS.n213 4.00459
R20487 IVS.n220 IVS.n219 4.00315
R20488 IVS.n212 IVS.n211 4.00315
R20489 IVS.n224 IVS.n223 3.9695
R20490 IVS.n218 IVS.n217 3.1505
R20491 IVS.n210 IVS.n209 3.1505
R20492 IVS.n178 IVS.n177 2.6005
R20493 IVS.n175 IVS.n174 2.6005
R20494 IVS.n75 IVS.n74 2.6005
R20495 IVS.n78 IVS.n77 2.6005
R20496 IVS.n106 IVS.n105 2.6005
R20497 IVS.n109 IVS.n108 2.6005
R20498 IVS.n52 IVS.n51 2.6005
R20499 IVS.n55 IVS.n54 2.6005
R20500 IVS.n29 IVS.n28 2.6005
R20501 IVS.n32 IVS.n31 2.6005
R20502 IVS.n150 IVS.n149 2.6005
R20503 IVS.n153 IVS.n152 2.6005
R20504 IVS.n4 IVS.n3 2.6005
R20505 IVS.n7 IVS.n6 2.6005
R20506 IVS.n87 IVS.n86 2.40398
R20507 IVS.n65 IVS.n64 2.40398
R20508 IVS.n42 IVS.n41 2.40398
R20509 IVS.n139 IVS.n138 2.40398
R20510 IVS.n19 IVS.n18 2.40398
R20511 IVS.n187 IVS.n186 2.40398
R20512 IVS.n230 IVS.n229 2.008
R20513 IVS.n110 IVS.n101 1.58214
R20514 IVS.n242 IVS.n241 1.49924
R20515 IVS.n233 IVS.n232 1.49862
R20516 IVS.n178 IVS.n175 1.4405
R20517 IVS.n78 IVS.n75 1.4405
R20518 IVS.n109 IVS.n106 1.4405
R20519 IVS.n55 IVS.n52 1.4405
R20520 IVS.n32 IVS.n29 1.4405
R20521 IVS.n153 IVS.n150 1.4405
R20522 IVS.n7 IVS.n4 1.4405
R20523 IVS.n236 IVS.n235 1.4405
R20524 IVS.n241 IVS.n240 1.4405
R20525 IVS.n231 IVS.n230 1.4405
R20526 IVS.n110 IVS.n109 1.36839
R20527 IVS.n179 IVS.n178 1.30464
R20528 IVS.n79 IVS.n78 1.30464
R20529 IVS.n56 IVS.n55 1.30464
R20530 IVS.n33 IVS.n32 1.30464
R20531 IVS.n154 IVS.n153 1.30464
R20532 IVS.n8 IVS.n7 1.30464
R20533 IVS.n225 IVS.n224 1.24943
R20534 IVS.n219 IVS.n218 1.24943
R20535 IVS.n211 IVS.n210 1.24943
R20536 IVS.n247 IVS.n195 1.13468
R20537 IVS.n89 IVS.n88 1.1255
R20538 IVS.n67 IVS.n66 1.1255
R20539 IVS.n44 IVS.n43 1.1255
R20540 IVS.n141 IVS.n140 1.1255
R20541 IVS.n21 IVS.n20 1.1255
R20542 IVS.n15 IVS.n14 1.1255
R20543 IVS.n145 IVS.n144 1.1255
R20544 IVS.n157 IVS.n156 1.1255
R20545 IVS.n61 IVS.n60 1.1255
R20546 IVS.n114 IVS.n113 1.1255
R20547 IVS.n84 IVS.n83 1.1255
R20548 IVS.n38 IVS.n37 1.1255
R20549 IVS.n183 IVS.n182 1.1255
R20550 IVS.n10 IVS.n9 1.1255
R20551 IVS.n119 IVS.n118 1.1255
R20552 IVS.n189 IVS.n188 1.1255
R20553 IVS.n247 IVS.n246 1.11782
R20554 IVS.n159 IVS.n142 0.885646
R20555 IVS.n191 IVS.n190 0.885413
R20556 IVS.n121 IVS.n120 0.885412
R20557 IVS.n159 IVS.n158 0.874835
R20558 IVS.n217 IVS.t59 0.8195
R20559 IVS.n217 IVS.n216 0.8195
R20560 IVS.n215 IVS.t71 0.8195
R20561 IVS.n215 IVS.n214 0.8195
R20562 IVS.n209 IVS.t75 0.8195
R20563 IVS.n209 IVS.n208 0.8195
R20564 IVS.n207 IVS.t67 0.8195
R20565 IVS.n207 IVS.n206 0.8195
R20566 IVS.n93 IVS.n90 0.727165
R20567 IVS.n131 IVS.n45 0.727165
R20568 IVS.n126 IVS.n68 0.616779
R20569 IVS.n164 IVS.n22 0.616779
R20570 IVS.n172 IVS.t20 0.607167
R20571 IVS.n172 IVS.n171 0.607167
R20572 IVS.n174 IVS.t15 0.607167
R20573 IVS.n174 IVS.n173 0.607167
R20574 IVS.n177 IVS.t14 0.607167
R20575 IVS.n177 IVS.n176 0.607167
R20576 IVS.n186 IVS.t52 0.607167
R20577 IVS.n186 IVS.n185 0.607167
R20578 IVS.n86 IVS.t54 0.607167
R20579 IVS.n86 IVS.n85 0.607167
R20580 IVS.n77 IVS.t16 0.607167
R20581 IVS.n77 IVS.n76 0.607167
R20582 IVS.n74 IVS.t17 0.607167
R20583 IVS.n74 IVS.n73 0.607167
R20584 IVS.n72 IVS.t21 0.607167
R20585 IVS.n72 IVS.n71 0.607167
R20586 IVS.n101 IVS.t13 0.607167
R20587 IVS.n101 IVS.n100 0.607167
R20588 IVS.n108 IVS.t29 0.607167
R20589 IVS.n108 IVS.n107 0.607167
R20590 IVS.n105 IVS.t30 0.607167
R20591 IVS.n105 IVS.n104 0.607167
R20592 IVS.n103 IVS.t32 0.607167
R20593 IVS.n103 IVS.n102 0.607167
R20594 IVS.n64 IVS.t5 0.607167
R20595 IVS.n64 IVS.n63 0.607167
R20596 IVS.n54 IVS.t25 0.607167
R20597 IVS.n54 IVS.n53 0.607167
R20598 IVS.n51 IVS.t26 0.607167
R20599 IVS.n51 IVS.n50 0.607167
R20600 IVS.n49 IVS.t27 0.607167
R20601 IVS.n49 IVS.n48 0.607167
R20602 IVS.n41 IVS.t22 0.607167
R20603 IVS.n41 IVS.n40 0.607167
R20604 IVS.n31 IVS.t34 0.607167
R20605 IVS.n31 IVS.n30 0.607167
R20606 IVS.n28 IVS.t35 0.607167
R20607 IVS.n28 IVS.n27 0.607167
R20608 IVS.n26 IVS.t38 0.607167
R20609 IVS.n26 IVS.n25 0.607167
R20610 IVS.n138 IVS.t33 0.607167
R20611 IVS.n138 IVS.n137 0.607167
R20612 IVS.n152 IVS.t49 0.607167
R20613 IVS.n152 IVS.n151 0.607167
R20614 IVS.n149 IVS.t50 0.607167
R20615 IVS.n149 IVS.n148 0.607167
R20616 IVS.n147 IVS.t53 0.607167
R20617 IVS.n147 IVS.n146 0.607167
R20618 IVS.n18 IVS.t45 0.607167
R20619 IVS.n18 IVS.n17 0.607167
R20620 IVS.n6 IVS.t8 0.607167
R20621 IVS.n6 IVS.n5 0.607167
R20622 IVS.n3 IVS.t10 0.607167
R20623 IVS.n3 IVS.n2 0.607167
R20624 IVS.n1 IVS.t12 0.607167
R20625 IVS.n1 IVS.n0 0.607167
R20626 IVS IVS.n250 0.451768
R20627 IVS IVS.n193 0.402965
R20628 IVS.n117 IVS.n116 0.198558
R20629 IVS.n65 IVS.n62 0.198558
R20630 IVS.n42 IVS.n39 0.198558
R20631 IVS.n139 IVS.n136 0.198558
R20632 IVS.n19 IVS.n16 0.198558
R20633 IVS.n180 IVS.n179 0.181594
R20634 IVS.n80 IVS.n79 0.181594
R20635 IVS.n57 IVS.n56 0.181594
R20636 IVS.n34 IVS.n33 0.181594
R20637 IVS.n156 IVS.n154 0.181594
R20638 IVS.n9 IVS.n8 0.181594
R20639 IVS.n246 IVS.n243 0.120289
R20640 IVS.n111 IVS.n110 0.114284
R20641 IVS.n190 IVS.n183 0.0999822
R20642 IVS.n120 IVS.n114 0.0999822
R20643 IVS.n83 IVS.n81 0.0953821
R20644 IVS.n112 IVS.n111 0.0953821
R20645 IVS.n60 IVS.n58 0.0953821
R20646 IVS.n37 IVS.n35 0.0953821
R20647 IVS.n14 IVS.n12 0.0953821
R20648 IVS.n182 IVS.n181 0.0953821
R20649 IVS.n188 IVS.n184 0.0953821
R20650 IVS.n170 IVS.n169 0.0939351
R20651 IVS.n96 IVS.n95 0.0847958
R20652 IVS.n124 IVS.n123 0.0847958
R20653 IVS.n129 IVS.n128 0.0847958
R20654 IVS.n134 IVS.n133 0.0847958
R20655 IVS.n162 IVS.n161 0.0847958
R20656 IVS.n167 IVS.n166 0.0847958
R20657 IVS.n45 IVS.n38 0.082822
R20658 IVS.n90 IVS.n84 0.082822
R20659 IVS.n158 IVS.n145 0.0743545
R20660 IVS.n22 IVS.n15 0.0712285
R20661 IVS.n68 IVS.n61 0.0712285
R20662 IVS.n84 IVS.n70 0.0625655
R20663 IVS.n38 IVS.n24 0.0625655
R20664 IVS.n70 IVS.n69 0.0625188
R20665 IVS.n24 IVS.n23 0.0625188
R20666 IVS.n99 IVS.n98 0.0623855
R20667 IVS.n114 IVS.n99 0.0623855
R20668 IVS.n47 IVS.n46 0.0623855
R20669 IVS.n61 IVS.n47 0.0623855
R20670 IVS.n11 IVS.n10 0.0623855
R20671 IVS.n15 IVS.n11 0.0623855
R20672 IVS.n118 IVS.n115 0.0620789
R20673 IVS.n68 IVS.n67 0.0534597
R20674 IVS.n22 IVS.n21 0.0534597
R20675 IVS.n158 IVS.n157 0.05104
R20676 IVS.n90 IVS.n89 0.0421496
R20677 IVS.n45 IVS.n44 0.0421496
R20678 IVS.n183 IVS.n170 0.0319869
R20679 IVS.n83 IVS.n82 0.0293873
R20680 IVS.n81 IVS.n80 0.0293873
R20681 IVS.n113 IVS.n112 0.0293873
R20682 IVS.n60 IVS.n59 0.0293873
R20683 IVS.n58 IVS.n57 0.0293873
R20684 IVS.n37 IVS.n36 0.0293873
R20685 IVS.n35 IVS.n34 0.0293873
R20686 IVS.n156 IVS.n155 0.0293873
R20687 IVS.n144 IVS.n143 0.0293873
R20688 IVS.n14 IVS.n13 0.0293873
R20689 IVS.n181 IVS.n180 0.0293873
R20690 IVS.n142 IVS.n141 0.0263867
R20691 IVS.n190 IVS.n189 0.0257704
R20692 IVS.n120 IVS.n119 0.0257704
R20693 IVS.n245 IVS.n244 0.0228651
R20694 IVS.n250 IVS.n249 0.0228651
R20695 IVS.n205 IVS.n204 0.0216961
R20696 IVS.n204 IVS.n203 0.019459
R20697 IVS.n238 IVS.n237 0.0192346
R20698 IVS.n88 IVS.n87 0.0185116
R20699 IVS.n118 IVS.n117 0.0185116
R20700 IVS.n66 IVS.n65 0.0185116
R20701 IVS.n43 IVS.n42 0.0185116
R20702 IVS.n140 IVS.n139 0.0185116
R20703 IVS.n20 IVS.n19 0.0185116
R20704 IVS.n188 IVS.n187 0.0185116
R20705 IVS.n248 IVS.n247 0.0173591
R20706 IVS.n195 IVS.n194 0.0173591
R20707 IVS.n239 IVS.n238 0.0133411
R20708 IVS.n246 IVS.n245 0.0119325
R20709 IVS.n249 IVS.n248 0.0119325
R20710 IVS.n241 IVS.n239 0.01175
R20711 IVS.n200 IVS.n199 0.00969794
R20712 IVS.n201 IVS.n200 0.00969794
R20713 IVS.n199 IVS.n198 0.00842254
R20714 IVS.n97 IVS.n96 0.00740328
R20715 IVS.n123 IVS.n122 0.00736358
R20716 IVS.n193 IVS.n192 0.00735609
R20717 IVS.n128 IVS.n127 0.0066903
R20718 IVS.n166 IVS.n165 0.0066903
R20719 IVS.n237 IVS.n236 0.00639353
R20720 IVS.n243 IVS.n242 0.0062755
R20721 IVS.n159 IVS.n135 0.00528925
R20722 IVS.n92 IVS.n91 0.00527411
R20723 IVS.n95 IVS.n94 0.00527411
R20724 IVS.n125 IVS.n124 0.00527411
R20725 IVS.n130 IVS.n129 0.00527411
R20726 IVS.n133 IVS.n132 0.00527411
R20727 IVS.n161 IVS.n160 0.00527411
R20728 IVS.n163 IVS.n162 0.00527411
R20729 IVS.n191 IVS.n168 0.00527411
R20730 IVS.n160 IVS.n159 0.00527411
R20731 IVS.n132 IVS.n131 0.00527411
R20732 IVS.n94 IVS.n93 0.00527411
R20733 IVS.n126 IVS.n125 0.00527411
R20734 IVS.n168 IVS.n167 0.00527411
R20735 IVS.n164 IVS.n163 0.00527411
R20736 IVS.n93 IVS.n92 0.00527411
R20737 IVS.n131 IVS.n130 0.00527411
R20738 IVS.n135 IVS.n134 0.00525899
R20739 IVS.n232 IVS.n231 0.00507635
R20740 IVS.n231 IVS.n205 0.00492687
R20741 IVS.n198 IVS.n197 0.00479961
R20742 IVS.n233 IVS.n202 0.00479961
R20743 IVS.n197 IVS.n196 0.00479961
R20744 IVS.n202 IVS.n201 0.00479961
R20745 IVS.n241 IVS.n234 0.00459425
R20746 IVS.n192 IVS.n191 0.00418876
R20747 IVS.n122 IVS.n121 0.00418126
R20748 IVS.n127 IVS.n126 0.00385522
R20749 IVS.n165 IVS.n164 0.00385522
R20750 IVS.n242 IVS.n233 0.00363775
R20751 IVS.n121 IVS.n97 0.00314088
R20752 VB1.n16 VB1.t4 63.68
R20753 VB1.n16 VB1.t2 63.68
R20754 VB1.n83 VB1.t41 61.7898
R20755 VB1.n90 VB1.t56 61.7898
R20756 VB1.n86 VB1.t60 61.7898
R20757 VB1.n87 VB1.t36 61.7898
R20758 VB1.n88 VB1.t40 61.7898
R20759 VB1.n89 VB1.t43 61.7898
R20760 VB1.n85 VB1.t54 61.7898
R20761 VB1.n84 VB1.t53 61.7898
R20762 VB1.n99 VB1.t61 61.5291
R20763 VB1.n100 VB1.t62 61.5291
R20764 VB1.n101 VB1.t38 61.5291
R20765 VB1.n102 VB1.t44 61.5291
R20766 VB1.n103 VB1.t48 61.5291
R20767 VB1.n104 VB1.t59 61.5291
R20768 VB1.n105 VB1.t47 61.5291
R20769 VB1.n91 VB1.t35 60.6166
R20770 VB1.n92 VB1.t64 60.6166
R20771 VB1.n93 VB1.t46 60.6166
R20772 VB1.n94 VB1.t34 60.6166
R20773 VB1.n95 VB1.t63 60.6166
R20774 VB1.n96 VB1.t45 60.6166
R20775 VB1.n98 VB1.t37 60.6166
R20776 VB1.n97 VB1.t50 60.6166
R20777 VB1.t57 VB1.n98 58.7916
R20778 VB1.n99 VB1.t66 57.8791
R20779 VB1.n100 VB1.t51 57.8791
R20780 VB1.n101 VB1.t58 57.8791
R20781 VB1.n102 VB1.t65 57.8791
R20782 VB1.n103 VB1.t49 57.8791
R20783 VB1.n104 VB1.t55 57.8791
R20784 VB1.n105 VB1.t42 57.8791
R20785 VB1.n106 VB1.t52 57.8791
R20786 VB1.t35 VB1.n90 57.6184
R20787 VB1.t63 VB1.n89 57.6184
R20788 VB1.t45 VB1.n85 57.6184
R20789 VB1.t37 VB1.n84 57.6184
R20790 VB1.n108 VB1.t57 56.0585
R20791 VB1.n87 VB1.n86 9.73383
R20792 VB1.n88 VB1.n87 9.73383
R20793 VB1.n89 VB1.n88 9.73383
R20794 VB1.n84 VB1.n83 9.73383
R20795 VB1.n92 VB1.n91 9.73383
R20796 VB1.n93 VB1.n92 9.73383
R20797 VB1.n94 VB1.n93 9.73383
R20798 VB1.n95 VB1.n94 9.73383
R20799 VB1.n96 VB1.n95 9.73383
R20800 VB1.n97 VB1.n96 9.73383
R20801 VB1.n98 VB1.n97 9.73383
R20802 VB1.n100 VB1.n99 9.73383
R20803 VB1.n101 VB1.n100 9.73383
R20804 VB1.n102 VB1.n101 9.73383
R20805 VB1.n103 VB1.n102 9.73383
R20806 VB1.n104 VB1.n103 9.73383
R20807 VB1.n105 VB1.n104 9.73383
R20808 VB1.n106 VB1.n105 9.73383
R20809 VB1.n60 VB1.t22 6.32241
R20810 VB1.n57 VB1.n56 6.32241
R20811 VB1.n44 VB1.t24 6.32241
R20812 VB1.n41 VB1.n40 6.32241
R20813 VB1.n27 VB1.t14 6.32241
R20814 VB1.n24 VB1.n23 6.32241
R20815 VB1.n17 VB1.n16 5.14084
R20816 VB1.n18 VB1.n17 4.52144
R20817 VB1.n64 VB1.n63 4.39485
R20818 VB1.n48 VB1.n47 4.36159
R20819 VB1.n31 VB1.n30 4.36159
R20820 VB1.n60 VB1.n59 3.43224
R20821 VB1.n57 VB1.n55 3.43224
R20822 VB1.n44 VB1.n43 3.43224
R20823 VB1.n41 VB1.n39 3.43224
R20824 VB1.n27 VB1.n26 3.43224
R20825 VB1.n24 VB1.n22 3.43224
R20826 VB1.n77 VB1.n76 3.1965
R20827 VB1.n112 VB1.n108 2.8805
R20828 VB1.n123 VB1.n122 2.32081
R20829 VB1.n107 VB1.n106 1.88633
R20830 VB1.n69 VB1.t30 1.6385
R20831 VB1.n69 VB1.n68 1.6385
R20832 VB1.n63 VB1.t6 1.6385
R20833 VB1.n63 VB1.n62 1.6385
R20834 VB1.n59 VB1.t19 1.6385
R20835 VB1.n59 VB1.n58 1.6385
R20836 VB1.n55 VB1.t1 1.6385
R20837 VB1.n55 VB1.n54 1.6385
R20838 VB1.n8 VB1.t26 1.6385
R20839 VB1.n8 VB1.n7 1.6385
R20840 VB1.n47 VB1.t15 1.6385
R20841 VB1.n47 VB1.n46 1.6385
R20842 VB1.n43 VB1.t8 1.6385
R20843 VB1.n43 VB1.n42 1.6385
R20844 VB1.n39 VB1.t12 1.6385
R20845 VB1.n39 VB1.n38 1.6385
R20846 VB1.n11 VB1.t17 1.6385
R20847 VB1.n11 VB1.n10 1.6385
R20848 VB1.n30 VB1.t9 1.6385
R20849 VB1.n30 VB1.n29 1.6385
R20850 VB1.n26 VB1.t32 1.6385
R20851 VB1.n26 VB1.n25 1.6385
R20852 VB1.n22 VB1.t20 1.6385
R20853 VB1.n22 VB1.n21 1.6385
R20854 VB1.n120 VB1.n119 1.50393
R20855 VB1.n80 VB1.n79 1.49812
R20856 VB1.n51 VB1.n37 1.49167
R20857 VB1.n53 VB1.n52 1.49167
R20858 VB1.n9 VB1.n8 1.42054
R20859 VB1.n12 VB1.n11 1.42054
R20860 VB1.n70 VB1.n69 1.42034
R20861 VB1.n108 VB1.n107 1.36152
R20862 VB1.n52 VB1.n9 1.15277
R20863 VB1.n36 VB1.n12 1.15277
R20864 VB1.n71 VB1.n70 1.15212
R20865 VB1.n127 VB1.n126 1.12675
R20866 VB1.n127 VB1.n81 1.126
R20867 VB1.n34 VB1.n33 1.1255
R20868 VB1.n51 VB1.n50 1.1255
R20869 VB1.n67 VB1.n66 1.1255
R20870 VB1.n35 VB1.n20 1.10736
R20871 VB1.n49 VB1.n48 1.07272
R20872 VB1.n32 VB1.n31 1.07272
R20873 VB1.n65 VB1.n64 1.03946
R20874 VB1.n119 VB1.n112 0.901294
R20875 VB1.n74 VB1.n72 0.722779
R20876 VB1.n17 VB1.n15 0.715901
R20877 VB1.n15 VB1.t3 0.4555
R20878 VB1.n15 VB1.n14 0.4555
R20879 VB1.n61 VB1.n60 0.337022
R20880 VB1.n45 VB1.n41 0.323326
R20881 VB1.n28 VB1.n24 0.323326
R20882 VB1.n64 VB1.n61 0.305717
R20883 VB1.n48 VB1.n45 0.305717
R20884 VB1.n31 VB1.n28 0.305717
R20885 VB1.n45 VB1.n44 0.303761
R20886 VB1.n28 VB1.n27 0.303761
R20887 VB1.n61 VB1.n57 0.290065
R20888 VB1.n52 VB1.n51 0.123658
R20889 VB1 VB1.n127 0.110576
R20890 VB1.n35 VB1.n34 0.0929251
R20891 VB1.n111 VB1.n110 0.0656316
R20892 VB1.n72 VB1.n71 0.0623678
R20893 VB1.n72 VB1.n67 0.0620327
R20894 VB1.n116 VB1.n115 0.0339644
R20895 VB1.n117 VB1.n116 0.0327802
R20896 VB1.n37 VB1.n36 0.0324737
R20897 VB1.n67 VB1.n53 0.0324737
R20898 VB1.n36 VB1.n35 0.0320039
R20899 VB1.n112 VB1.n111 0.0301053
R20900 VB1.n118 VB1.n117 0.0301053
R20901 VB1.n110 VB1.n109 0.0289211
R20902 VB1.n115 VB1.n114 0.0289211
R20903 VB1.n6 VB1.n5 0.0207053
R20904 VB1.n1 VB1.n0 0.0207053
R20905 VB1.n74 VB1.n73 0.0156875
R20906 VB1.n66 VB1.n65 0.014283
R20907 VB1.n50 VB1.n49 0.014283
R20908 VB1.n33 VB1.n32 0.014283
R20909 VB1.n4 VB1.n3 0.014
R20910 VB1.n5 VB1.n4 0.0134654
R20911 VB1.n20 VB1.n19 0.00860784
R20912 VB1.n75 VB1.n74 0.00860784
R20913 VB1.n122 VB1.n121 0.00858096
R20914 VB1.n120 VB1.n82 0.00858096
R20915 VB1.n121 VB1.n120 0.00858096
R20916 VB1.n19 VB1.n18 0.00855417
R20917 VB1.n76 VB1.n75 0.00855417
R20918 VB1.n126 VB1.n124 0.00773989
R20919 VB1.n78 VB1.n77 0.00773989
R20920 VB1.n124 VB1.n123 0.00773989
R20921 VB1.n79 VB1.n78 0.00773989
R20922 VB1.n3 VB1.n2 0.00773989
R20923 VB1.n126 VB1.n125 0.00773989
R20924 VB1.n79 VB1.n6 0.00773989
R20925 VB1.n81 VB1.n1 0.00773989
R20926 VB1.n114 VB1.n113 0.00685938
R20927 VB1.n20 VB1.n13 0.00605114
R20928 VB1.n81 VB1.n80 0.00582347
R20929 VB1.n119 VB1.n118 0.0030309
R20930 VPD.n82 VPD.t27 5.22731
R20931 VPD.n76 VPD.n75 5.20893
R20932 VPD.n73 VPD.t0 5.20893
R20933 VPD.n72 VPD.n71 5.20893
R20934 VPD.n42 VPD.n41 5.11385
R20935 VPD.n59 VPD.t5 5.11385
R20936 VPD.n67 VPD.t23 4.55153
R20937 VPD.n5 VPD.t31 4.55153
R20938 VPD.n48 VPD.n47 4.53238
R20939 VPD.n69 VPD.n65 3.92545
R20940 VPD.n68 VPD.t17 3.92545
R20941 VPD.n67 VPD.n66 3.92545
R20942 VPD.n6 VPD.t28 3.92545
R20943 VPD.n5 VPD.n4 3.92545
R20944 VPD.n76 VPD.n74 3.18197
R20945 VPD.n73 VPD.t22 3.18197
R20946 VPD.n72 VPD.n70 3.18197
R20947 VPD.n104 VPD.n36 2.26197
R20948 VPD.n141 VPD.n137 2.24763
R20949 VPD.n141 VPD.n112 2.24763
R20950 VPD.n77 VPD.n76 1.87093
R20951 VPD.n82 VPD.n81 1.55818
R20952 VPD.n7 VPD.n6 1.276
R20953 VPD.n117 VPD.n116 1.19453
R20954 VPD.n128 VPD.n127 1.19453
R20955 VPD.n39 VPD.n38 1.18339
R20956 VPD.n53 VPD.n52 1.18339
R20957 VPD.n57 VPD.n56 1.18339
R20958 VPD.n2 VPD.n1 1.18328
R20959 VPD.n20 VPD.n19 1.17867
R20960 VPD.n31 VPD.n30 1.17867
R20961 VPD.n142 VPD.n107 1.1775
R20962 VPD.n40 VPD.n39 1.17279
R20963 VPD.n54 VPD.n53 1.17279
R20964 VPD.n58 VPD.n57 1.17279
R20965 VPD.n3 VPD.n2 1.17279
R20966 VPD.n68 VPD.n67 1.12746
R20967 VPD.n6 VPD.n5 1.12746
R20968 VPD.n87 VPD.n86 1.12717
R20969 VPD.n44 VPD.n43 1.1255
R20970 VPD.n61 VPD.n60 1.1255
R20971 VPD.n86 VPD.n85 1.1255
R20972 VPD.n50 VPD.n49 1.1255
R20973 VPD.n9 VPD.n8 1.1255
R20974 VPD.n142 VPD.n141 1.1255
R20975 VPD.n104 VPD.n103 0.927211
R20976 VPD.n79 VPD.n78 0.877022
R20977 VPD.n15 VPD.n14 0.87575
R20978 VPD.n19 VPD.n18 0.824494
R20979 VPD.n30 VPD.n29 0.824494
R20980 VPD.n116 VPD.n115 0.824332
R20981 VPD.n127 VPD.n126 0.824332
R20982 VPD.n77 VPD.n73 0.743978
R20983 VPD.n78 VPD.n72 0.743978
R20984 VPD.n23 VPD.n22 0.727916
R20985 VPD.n34 VPD.n33 0.727916
R20986 VPD.n131 VPD.n130 0.727916
R20987 VPD.n97 VPD.n55 0.727104
R20988 VPD.n69 VPD.n68 0.626587
R20989 VPD.n78 VPD.n77 0.626587
R20990 VPD.n91 VPD.n90 0.62375
R20991 VPD.n101 VPD.n45 0.616779
R20992 VPD.n92 VPD.n62 0.616779
R20993 VPD.n12 VPD.n10 0.616779
R20994 VPD.n120 VPD.n118 0.616779
R20995 VPD.n38 VPD.n37 0.58197
R20996 VPD.n52 VPD.t16 0.58197
R20997 VPD.n52 VPD.n51 0.58197
R20998 VPD.n47 VPD.t10 0.58197
R20999 VPD.n47 VPD.n46 0.58197
R21000 VPD.n56 VPD.t13 0.58197
R21001 VPD.n81 VPD.t18 0.58197
R21002 VPD.n1 VPD.n0 0.58197
R21003 VPD.n18 VPD.t6 0.58197
R21004 VPD.n18 VPD.n17 0.58197
R21005 VPD.n29 VPD.t8 0.58197
R21006 VPD.n29 VPD.n28 0.58197
R21007 VPD.n115 VPD.t7 0.58197
R21008 VPD.n115 VPD.n114 0.58197
R21009 VPD.n126 VPD.t3 0.58197
R21010 VPD.n126 VPD.n125 0.58197
R21011 VPD.n134 VPD.n133 0.53025
R21012 VPD.n80 VPD.n79 0.442674
R21013 VPD.n79 VPD.n69 0.3605
R21014 VPD.n8 VPD.n7 0.330999
R21015 VPD.n100 VPD.n99 0.330125
R21016 VPD.n95 VPD.n94 0.330125
R21017 VPD.n26 VPD.n25 0.330125
R21018 VPD.n123 VPD.n122 0.330125
R21019 VPD.n43 VPD.n42 0.32803
R21020 VPD.n49 VPD.n48 0.32803
R21021 VPD.n60 VPD.n59 0.32803
R21022 VPD.n105 VPD.n104 0.321971
R21023 VPD VPD.n142 0.29625
R21024 VPD.n83 VPD.n82 0.201042
R21025 VPD.n84 VPD.n83 0.0953821
R21026 VPD.n86 VPD.n64 0.0832399
R21027 VPD.n22 VPD.n21 0.0826464
R21028 VPD.n33 VPD.n32 0.0826464
R21029 VPD.n130 VPD.n129 0.0826464
R21030 VPD.n55 VPD.n50 0.0823987
R21031 VPD.n62 VPD.n58 0.0712285
R21032 VPD.n45 VPD.n40 0.0712285
R21033 VPD.n10 VPD.n3 0.0712285
R21034 VPD.n118 VPD.n113 0.0712285
R21035 VPD.n85 VPD.n80 0.0552826
R21036 VPD.n45 VPD.n44 0.0534597
R21037 VPD.n62 VPD.n61 0.0534597
R21038 VPD.n10 VPD.n9 0.0534597
R21039 VPD.n118 VPD.n117 0.0534597
R21040 VPD.n22 VPD.n20 0.0423164
R21041 VPD.n33 VPD.n31 0.0423164
R21042 VPD.n130 VPD.n128 0.0423164
R21043 VPD.n64 VPD.n63 0.0419676
R21044 VPD.n55 VPD.n54 0.0415773
R21045 VPD.n85 VPD.n84 0.0293873
R21046 VPD.n139 VPD.n138 0.0207053
R21047 VPD.n112 VPD.n111 0.0207053
R21048 VPD.n101 VPD.n100 0.0156875
R21049 VPD.n92 VPD.n91 0.0156875
R21050 VPD.n12 VPD.n11 0.0156875
R21051 VPD.n120 VPD.n119 0.0156875
R21052 VPD.n141 VPD.n140 0.014
R21053 VPD.n140 VPD.n139 0.0134654
R21054 VPD.n102 VPD.n101 0.00860784
R21055 VPD.n97 VPD.n96 0.00860784
R21056 VPD.n93 VPD.n92 0.00860784
R21057 VPD.n89 VPD.n88 0.00860784
R21058 VPD.n13 VPD.n12 0.00860784
R21059 VPD.n121 VPD.n120 0.00860784
R21060 VPD.n99 VPD.n98 0.00858096
R21061 VPD.n98 VPD.n97 0.00858096
R21062 VPD.n35 VPD.n34 0.00858096
R21063 VPD.n27 VPD.n26 0.00858096
R21064 VPD.n24 VPD.n23 0.00858096
R21065 VPD.n16 VPD.n15 0.00858096
R21066 VPD.n36 VPD.n35 0.00858096
R21067 VPD.n34 VPD.n27 0.00858096
R21068 VPD.n25 VPD.n24 0.00858096
R21069 VPD.n23 VPD.n16 0.00858096
R21070 VPD.n132 VPD.n131 0.00858096
R21071 VPD.n124 VPD.n123 0.00858096
R21072 VPD.n133 VPD.n132 0.00858096
R21073 VPD.n131 VPD.n124 0.00858096
R21074 VPD.n103 VPD.n102 0.00855417
R21075 VPD.n96 VPD.n95 0.00855417
R21076 VPD.n94 VPD.n93 0.00855417
R21077 VPD.n90 VPD.n89 0.00855417
R21078 VPD.n14 VPD.n13 0.00855417
R21079 VPD.n122 VPD.n121 0.00855417
R21080 VPD.n106 VPD.n105 0.00773989
R21081 VPD.n135 VPD.n134 0.00773989
R21082 VPD.n110 VPD.n109 0.00773989
R21083 VPD.n136 VPD.n135 0.00773989
R21084 VPD.n107 VPD.n106 0.00773989
R21085 VPD.n137 VPD.n136 0.00773989
R21086 VPD.n112 VPD.n110 0.00773989
R21087 VPD.n141 VPD.n108 0.00461413
R21088 VPD.n88 VPD.n87 0.00364318
R21089 OUT1.t45 OUT1.t85 122.014
R21090 OUT1.t88 OUT1.t72 122.014
R21091 OUT1.t71 OUT1.t103 122.014
R21092 OUT1.t99 OUT1.t105 122.014
R21093 OUT1.t44 OUT1.t70 122.014
R21094 OUT1.t40 OUT1.t37 122.014
R21095 OUT1.t84 OUT1.t63 122.014
R21096 OUT1.t49 OUT1.t66 122.014
R21097 OUT1.t57 OUT1.t91 122.014
R21098 OUT1.t104 OUT1.t89 122.014
R21099 OUT1.t36 OUT1.t78 122.014
R21100 OUT1.t54 OUT1.t97 122.014
R21101 OUT1.n34 OUT1.t106 68.0848
R21102 OUT1.n68 OUT1.t51 65.7181
R21103 OUT1.n72 OUT1.t83 65.7181
R21104 OUT1.n35 OUT1.t100 65.7179
R21105 OUT1.n71 OUT1.t47 65.7179
R21106 OUT1.n75 OUT1.t102 65.7179
R21107 OUT1.n84 OUT1.t55 63.548
R21108 OUT1.n77 OUT1.t99 63.548
R21109 OUT1.n52 OUT1.t61 63.548
R21110 OUT1.n61 OUT1.t43 63.548
R21111 OUT1.n37 OUT1.t49 63.548
R21112 OUT1.n46 OUT1.t54 63.548
R21113 OUT1.n87 OUT1.t50 62.5719
R21114 OUT1.n85 OUT1.t53 62.5719
R21115 OUT1.n83 OUT1.t92 62.5719
R21116 OUT1.n80 OUT1.t98 62.5719
R21117 OUT1.n78 OUT1.t71 62.5719
R21118 OUT1.n76 OUT1.t75 62.5719
R21119 OUT1.n73 OUT1.t58 62.5719
R21120 OUT1.n69 OUT1.t93 62.5719
R21121 OUT1.n55 OUT1.t82 62.5719
R21122 OUT1.n53 OUT1.t59 62.5719
R21123 OUT1.n51 OUT1.t41 62.5719
R21124 OUT1.n58 OUT1.t56 62.5719
R21125 OUT1.n59 OUT1.t107 62.5719
R21126 OUT1.n60 OUT1.t77 62.5719
R21127 OUT1.n40 OUT1.t68 62.5719
R21128 OUT1.n38 OUT1.t84 62.5719
R21129 OUT1.n36 OUT1.t90 62.5719
R21130 OUT1.n43 OUT1.t42 62.5719
R21131 OUT1.n44 OUT1.t36 62.5719
R21132 OUT1.n45 OUT1.t60 62.5719
R21133 OUT1.n33 OUT1.t76 62.5719
R21134 OUT1.n64 OUT1.t67 61.8074
R21135 OUT1.n49 OUT1.t57 61.8074
R21136 OUT1.n89 OUT1.t73 61.8072
R21137 OUT1.n82 OUT1.t45 61.8072
R21138 OUT1.n57 OUT1.t38 61.8072
R21139 OUT1.n42 OUT1.t44 61.8072
R21140 OUT1.n87 OUT1.t64 41.7148
R21141 OUT1.n85 OUT1.t69 41.7148
R21142 OUT1.n83 OUT1.t48 41.7148
R21143 OUT1.n80 OUT1.t52 41.7148
R21144 OUT1.n78 OUT1.t88 41.7148
R21145 OUT1.n76 OUT1.t95 41.7148
R21146 OUT1.n73 OUT1.t79 41.7148
R21147 OUT1.n69 OUT1.t87 41.7148
R21148 OUT1.n55 OUT1.t80 41.7148
R21149 OUT1.n53 OUT1.t74 41.7148
R21150 OUT1.n51 OUT1.t46 41.7148
R21151 OUT1.n58 OUT1.t39 41.7148
R21152 OUT1.n59 OUT1.t65 41.7148
R21153 OUT1.n60 OUT1.t101 41.7148
R21154 OUT1.n40 OUT1.t62 41.7148
R21155 OUT1.n38 OUT1.t40 41.7148
R21156 OUT1.n36 OUT1.t94 41.7148
R21157 OUT1.n43 OUT1.t86 41.7148
R21158 OUT1.n44 OUT1.t104 41.7148
R21159 OUT1.n45 OUT1.t81 41.7148
R21160 OUT1.n33 OUT1.t96 41.7148
R21161 OUT1.n74 OUT1.n73 17.8184
R21162 OUT1.n70 OUT1.n69 17.8184
R21163 OUT1.n34 OUT1.n33 17.8184
R21164 OUT1.n88 OUT1.n87 15.9934
R21165 OUT1.n84 OUT1.n83 15.9934
R21166 OUT1.n81 OUT1.n80 15.9934
R21167 OUT1.n77 OUT1.n76 15.9934
R21168 OUT1.n56 OUT1.n55 15.9934
R21169 OUT1.n52 OUT1.n51 15.9934
R21170 OUT1.n63 OUT1.n58 15.9934
R21171 OUT1.n61 OUT1.n60 15.9934
R21172 OUT1.n41 OUT1.n40 15.9934
R21173 OUT1.n37 OUT1.n36 15.9934
R21174 OUT1.n48 OUT1.n43 15.9934
R21175 OUT1.n46 OUT1.n45 15.9934
R21176 OUT1.n86 OUT1.n85 13.9076
R21177 OUT1.n79 OUT1.n78 13.9076
R21178 OUT1.n54 OUT1.n53 13.9076
R21179 OUT1.n62 OUT1.n59 13.9076
R21180 OUT1.n39 OUT1.n38 13.9076
R21181 OUT1.n47 OUT1.n44 13.9076
R21182 OUT1.n92 OUT1.n91 8.881
R21183 OUT1.n90 OUT1.n89 8.79758
R21184 OUT1.n165 OUT1.n164 8.0005
R21185 OUT1.n155 OUT1.n152 8.0005
R21186 OUT1.n72 OUT1.n71 7.75675
R21187 OUT1.n156 OUT1.t20 6.49823
R21188 OUT1.n156 OUT1.t22 6.4095
R21189 OUT1.n66 OUT1.n65 5.6201
R21190 OUT1.n120 OUT1.n119 5.52316
R21191 OUT1.n101 OUT1.n100 5.49577
R21192 OUT1.n90 OUT1.n82 5.42798
R21193 OUT1.n123 OUT1.t13 5.40577
R21194 OUT1.n126 OUT1.n124 5.40577
R21195 OUT1.n127 OUT1.t15 5.40577
R21196 OUT1.n116 OUT1.n115 5.31701
R21197 OUT1.n241 OUT1.n240 4.67186
R21198 OUT1.n122 OUT1.t12 4.64664
R21199 OUT1.n229 OUT1.n226 4.54551
R21200 OUT1.n91 OUT1.n90 4.5329
R21201 OUT1.n67 OUT1.n66 4.5329
R21202 OUT1.n233 OUT1.n232 4.50858
R21203 OUT1.n198 OUT1.n197 4.50855
R21204 OUT1.n13 OUT1.n12 4.50855
R21205 OUT1.n111 OUT1.n97 4.5005
R21206 OUT1.n108 OUT1.n97 4.5005
R21207 OUT1.n109 OUT1.n108 4.5005
R21208 OUT1.n235 OUT1.n220 4.5005
R21209 OUT1.n246 OUT1.n220 4.5005
R21210 OUT1.n234 OUT1.n233 4.5005
R21211 OUT1.n246 OUT1.n245 4.5005
R21212 OUT1.n140 OUT1.n113 4.5005
R21213 OUT1.n137 OUT1.n113 4.5005
R21214 OUT1.n138 OUT1.n137 4.5005
R21215 OUT1.n210 OUT1.n190 4.5005
R21216 OUT1.n215 OUT1.n190 4.5005
R21217 OUT1.n208 OUT1.n207 4.5005
R21218 OUT1.n209 OUT1.n208 4.5005
R21219 OUT1.n203 OUT1.n197 4.5005
R21220 OUT1.n203 OUT1.n202 4.5005
R21221 OUT1.n215 OUT1.n214 4.5005
R21222 OUT1.n159 OUT1.n151 4.5005
R21223 OUT1.n163 OUT1.n159 4.5005
R21224 OUT1.n172 OUT1.n151 4.5005
R21225 OUT1.n168 OUT1.n157 4.5005
R21226 OUT1.n172 OUT1.n149 4.5005
R21227 OUT1.n172 OUT1.n171 4.5005
R21228 OUT1.n25 OUT1.n5 4.5005
R21229 OUT1.n30 OUT1.n5 4.5005
R21230 OUT1.n23 OUT1.n22 4.5005
R21231 OUT1.n24 OUT1.n23 4.5005
R21232 OUT1.n18 OUT1.n12 4.5005
R21233 OUT1.n18 OUT1.n17 4.5005
R21234 OUT1.n30 OUT1.n29 4.5005
R21235 OUT1.n252 OUT1.n92 4.5005
R21236 OUT1.n255 OUT1.n31 4.5005
R21237 OUT1.n251 OUT1.n96 4.5005
R21238 OUT1.n255 OUT1.n32 4.5005
R21239 OUT1.n252 OUT1.n251 4.5005
R21240 OUT1.n120 OUT1.t16 4.39621
R21241 OUT1.n121 OUT1.n118 4.39621
R21242 OUT1.n101 OUT1.t34 4.36882
R21243 OUT1.n102 OUT1.n99 4.36882
R21244 OUT1.n182 OUT1.n181 3.79067
R21245 OUT1.n123 OUT1.t21 3.71925
R21246 OUT1.n126 OUT1.n125 3.71925
R21247 OUT1.n127 OUT1.t18 3.71925
R21248 OUT1.n216 OUT1.n188 3.19194
R21249 OUT1.n65 OUT1.n57 3.17917
R21250 OUT1.n50 OUT1.n42 3.17917
R21251 OUT1.n67 OUT1.n35 3.17917
R21252 OUT1.n65 OUT1.n64 3.17779
R21253 OUT1.n50 OUT1.n49 3.17779
R21254 OUT1.n91 OUT1.n75 3.17736
R21255 OUT1.n68 OUT1.n67 3.17716
R21256 OUT1.n133 OUT1.n116 3.10759
R21257 OUT1.n133 OUT1.n131 2.61464
R21258 OUT1.n134 OUT1.n133 2.61112
R21259 OUT1.n229 OUT1.n228 2.56103
R21260 OUT1.n155 OUT1.t4 2.4095
R21261 OUT1.n165 OUT1.t24 2.4095
R21262 OUT1.n110 OUT1.n109 2.25517
R21263 OUT1.n245 OUT1.n236 2.25517
R21264 OUT1.n231 OUT1.n221 2.25517
R21265 OUT1.n139 OUT1.n138 2.25517
R21266 OUT1.n214 OUT1.n211 2.25517
R21267 OUT1.n205 OUT1.n191 2.25517
R21268 OUT1.n202 OUT1.n198 2.25517
R21269 OUT1.n29 OUT1.n26 2.25517
R21270 OUT1.n20 OUT1.n6 2.25517
R21271 OUT1.n17 OUT1.n13 2.25517
R21272 OUT1.n255 OUT1.n3 2.25362
R21273 OUT1.n168 OUT1.n167 2.25068
R21274 OUT1.n66 OUT1.n50 2.2505
R21275 OUT1.n163 OUT1.n161 2.2505
R21276 OUT1.n162 OUT1.n149 2.2505
R21277 OUT1.n161 OUT1.n151 2.2505
R21278 OUT1.n161 OUT1.n158 2.2505
R21279 OUT1.n168 OUT1.n158 2.2505
R21280 OUT1.n163 OUT1.n162 2.2505
R21281 OUT1.n162 OUT1.n158 2.2505
R21282 OUT1.n162 OUT1.n151 2.2505
R21283 OUT1.n147 OUT1.n145 2.2505
R21284 OUT1.n179 OUT1.n147 2.2505
R21285 OUT1.n179 OUT1.n178 2.2505
R21286 OUT1.n176 OUT1.n175 2.2505
R21287 OUT1.n96 OUT1.n2 2.24763
R21288 OUT1.n96 OUT1.n95 2.24763
R21289 OUT1.n94 OUT1.n0 2.24763
R21290 OUT1.n255 OUT1.n254 2.24763
R21291 OUT1.n96 OUT1.n1 2.24763
R21292 OUT1.n232 OUT1.n231 2.24721
R21293 OUT1.n206 OUT1.n205 2.24721
R21294 OUT1.n21 OUT1.n20 2.24721
R21295 OUT1.n252 OUT1.n93 2.24477
R21296 OUT1.n253 OUT1.n0 2.24477
R21297 OUT1.n105 OUT1.n104 1.84515
R21298 OUT1.n103 OUT1.n102 1.80781
R21299 OUT1.n104 OUT1.n103 1.76998
R21300 OUT1.n243 OUT1.n238 1.63933
R21301 OUT1.n241 OUT1.n238 1.55253
R21302 OUT1.n169 OUT1.n168 1.50171
R21303 OUT1.n184 OUT1.n143 1.5005
R21304 OUT1.n186 OUT1.n185 1.5005
R21305 OUT1.n3 OUT1.n0 1.50031
R21306 OUT1.n163 OUT1.n150 1.50014
R21307 OUT1.n171 OUT1.n153 1.5001
R21308 OUT1.n160 OUT1.n149 1.4978
R21309 OUT1.n173 OUT1.n148 1.49678
R21310 OUT1.n175 OUT1.n174 1.49371
R21311 OUT1.n166 OUT1.n165 1.43397
R21312 OUT1.n170 OUT1.n155 1.4339
R21313 OUT1.n200 OUT1.n199 1.40904
R21314 OUT1.n212 OUT1.t7 1.40904
R21315 OUT1.n15 OUT1.n14 1.40609
R21316 OUT1.n27 OUT1.t11 1.40609
R21317 OUT1.n128 OUT1.n127 1.27615
R21318 OUT1.n71 OUT1.n70 1.21895
R21319 OUT1.n74 OUT1.n72 1.21875
R21320 OUT1.n217 OUT1.n140 1.20171
R21321 OUT1.n200 OUT1.n197 1.19459
R21322 OUT1.n212 OUT1.n190 1.19459
R21323 OUT1.n20 OUT1.n10 1.19453
R21324 OUT1.n15 OUT1.n12 1.19451
R21325 OUT1.n27 OUT1.n5 1.19451
R21326 OUT1.n205 OUT1.n195 1.19431
R21327 OUT1.n228 OUT1.n223 1.18237
R21328 OUT1.n208 OUT1.n195 1.17925
R21329 OUT1.n23 OUT1.n10 1.17901
R21330 OUT1.n202 OUT1.n200 1.17899
R21331 OUT1.n214 OUT1.n212 1.17899
R21332 OUT1.n17 OUT1.n15 1.17808
R21333 OUT1.n29 OUT1.n27 1.17808
R21334 OUT1.n256 OUT1.n0 1.1775
R21335 OUT1.n233 OUT1.n223 1.17275
R21336 OUT1.n250 OUT1.n112 1.1515
R21337 OUT1.n247 OUT1.n218 1.1515
R21338 OUT1.n245 OUT1.n243 1.14574
R21339 OUT1.n105 OUT1.n97 1.14438
R21340 OUT1.n129 OUT1.n128 1.12746
R21341 OUT1.n109 OUT1.n106 1.1255
R21342 OUT1.n242 OUT1.n220 1.1255
R21343 OUT1.n231 OUT1.n230 1.1255
R21344 OUT1.n138 OUT1.n135 1.1255
R21345 OUT1.n117 OUT1.n113 1.1255
R21346 OUT1.n249 OUT1.n248 1.1255
R21347 OUT1.n256 OUT1.n255 1.1255
R21348 OUT1.n171 OUT1.n154 1.12145
R21349 OUT1.n181 OUT1.n180 1.12145
R21350 OUT1.n175 OUT1.n144 1.11801
R21351 OUT1.n177 OUT1.n145 1.11782
R21352 OUT1.n179 OUT1.n146 1.11782
R21353 OUT1.n75 OUT1.n74 0.905911
R21354 OUT1.n35 OUT1.n34 0.90591
R21355 OUT1.n70 OUT1.n68 0.905703
R21356 OUT1.n216 OUT1.n215 0.890545
R21357 OUT1.n122 OUT1.n121 0.877022
R21358 OUT1.n218 OUT1.n217 0.873064
R21359 OUT1.n195 OUT1.n194 0.827253
R21360 OUT1.n10 OUT1.n9 0.824332
R21361 OUT1.n183 OUT1.n141 0.783458
R21362 OUT1.n188 OUT1.n187 0.767554
R21363 OUT1.n142 OUT1.n141 0.7505
R21364 OUT1.n224 OUT1.n222 0.727104
R21365 OUT1.n204 OUT1.n192 0.727104
R21366 OUT1.n19 OUT1.n7 0.727104
R21367 OUT1.n129 OUT1.n123 0.650065
R21368 OUT1.n128 OUT1.n126 0.650065
R21369 OUT1.n86 OUT1.n84 0.626587
R21370 OUT1.n88 OUT1.n86 0.626587
R21371 OUT1.n79 OUT1.n77 0.626587
R21372 OUT1.n81 OUT1.n79 0.626587
R21373 OUT1.n54 OUT1.n52 0.626587
R21374 OUT1.n56 OUT1.n54 0.626587
R21375 OUT1.n63 OUT1.n62 0.626587
R21376 OUT1.n62 OUT1.n61 0.626587
R21377 OUT1.n39 OUT1.n37 0.626587
R21378 OUT1.n41 OUT1.n39 0.626587
R21379 OUT1.n48 OUT1.n47 0.626587
R21380 OUT1.n47 OUT1.n46 0.626587
R21381 OUT1.n102 OUT1.n101 0.626587
R21382 OUT1.n121 OUT1.n120 0.626587
R21383 OUT1.n130 OUT1.n129 0.626587
R21384 OUT1.n107 OUT1.n98 0.616779
R21385 OUT1.n244 OUT1.n219 0.616779
R21386 OUT1.n136 OUT1.n114 0.616779
R21387 OUT1.n201 OUT1.n196 0.616779
R21388 OUT1.n213 OUT1.n189 0.616779
R21389 OUT1.n16 OUT1.n11 0.616779
R21390 OUT1.n28 OUT1.n4 0.616779
R21391 OUT1.n228 OUT1.t10 0.58197
R21392 OUT1.n228 OUT1.n227 0.58197
R21393 OUT1.n226 OUT1.t8 0.58197
R21394 OUT1.n226 OUT1.n225 0.58197
R21395 OUT1.n238 OUT1.t2 0.58197
R21396 OUT1.n238 OUT1.n237 0.58197
R21397 OUT1.n240 OUT1.t30 0.58197
R21398 OUT1.n240 OUT1.n239 0.58197
R21399 OUT1.n194 OUT1.t27 0.58197
R21400 OUT1.n194 OUT1.n193 0.58197
R21401 OUT1.n9 OUT1.t26 0.58197
R21402 OUT1.n9 OUT1.n8 0.58197
R21403 OUT1.n104 OUT1.t3 0.56925
R21404 OUT1.n133 OUT1.n132 0.56925
R21405 OUT1.n247 OUT1.n246 0.5585
R21406 OUT1.n112 OUT1.n111 0.54725
R21407 OUT1.n175 OUT1.n172 0.50922
R21408 OUT1.n217 OUT1.n216 0.485118
R21409 OUT1.n235 OUT1.n234 0.474125
R21410 OUT1.n207 OUT1.n203 0.474125
R21411 OUT1.n210 OUT1.n209 0.474125
R21412 OUT1.n22 OUT1.n18 0.474125
R21413 OUT1.n25 OUT1.n24 0.474125
R21414 OUT1.n230 OUT1.n229 0.366599
R21415 OUT1.n31 OUT1.n30 0.312
R21416 OUT1.n183 OUT1.n182 0.299983
R21417 OUT1.n135 OUT1.n116 0.293265
R21418 OUT1.n89 OUT1.n88 0.279823
R21419 OUT1.n82 OUT1.n81 0.279823
R21420 OUT1.n57 OUT1.n56 0.279823
R21421 OUT1.n42 OUT1.n41 0.279823
R21422 OUT1.n64 OUT1.n63 0.279615
R21423 OUT1.n49 OUT1.n48 0.279615
R21424 OUT1.n242 OUT1.n241 0.223214
R21425 OUT1.n251 OUT1.n250 0.221875
R21426 OUT1.n130 OUT1.n122 0.1805
R21427 OUT1.n106 OUT1.n103 0.171378
R21428 OUT1.n131 OUT1.n130 0.163273
R21429 OUT1.n187 OUT1.n186 0.147906
R21430 OUT1.n106 OUT1.n105 0.106358
R21431 OUT1.n243 OUT1.n242 0.104922
R21432 OUT1.n134 OUT1.n117 0.0982964
R21433 OUT1.n231 OUT1.n222 0.0823987
R21434 OUT1.n205 OUT1.n192 0.0823987
R21435 OUT1.n20 OUT1.n7 0.0823987
R21436 OUT1.n230 OUT1.n223 0.076187
R21437 OUT1.n109 OUT1.n107 0.0712285
R21438 OUT1.n245 OUT1.n244 0.0712285
R21439 OUT1.n138 OUT1.n136 0.0712285
R21440 OUT1.n214 OUT1.n213 0.0712285
R21441 OUT1.n202 OUT1.n201 0.0712285
R21442 OUT1.n29 OUT1.n28 0.0712285
R21443 OUT1.n17 OUT1.n16 0.0712285
R21444 OUT1.n157 OUT1.n156 0.0607113
R21445 OUT1.n107 OUT1.n97 0.0534597
R21446 OUT1.n244 OUT1.n220 0.0534597
R21447 OUT1.n136 OUT1.n113 0.0534597
R21448 OUT1.n201 OUT1.n197 0.0534597
R21449 OUT1.n213 OUT1.n190 0.0534597
R21450 OUT1.n16 OUT1.n12 0.0534597
R21451 OUT1.n28 OUT1.n5 0.0534597
R21452 OUT1.n250 OUT1.n249 0.0525
R21453 OUT1.n249 OUT1.n218 0.0525
R21454 OUT1.n233 OUT1.n222 0.0415773
R21455 OUT1.n208 OUT1.n192 0.0415773
R21456 OUT1.n23 OUT1.n7 0.0415773
R21457 OUT1.n188 OUT1.n141 0.0334577
R21458 OUT1.n135 OUT1.n134 0.0265124
R21459 OUT1.n248 OUT1.n112 0.0265
R21460 OUT1.n248 OUT1.n247 0.0265
R21461 OUT1.n174 OUT1.n173 0.0228651
R21462 OUT1.n158 OUT1.n152 0.0214155
R21463 OUT1.n164 OUT1.n158 0.0210986
R21464 OUT1.n93 OUT1.n2 0.0207053
R21465 OUT1.n254 OUT1.n253 0.0207053
R21466 OUT1.n95 OUT1.n93 0.0207053
R21467 OUT1.n131 OUT1.n117 0.0204805
R21468 OUT1.n170 OUT1.n169 0.0204798
R21469 OUT1.n167 OUT1.n166 0.0195995
R21470 OUT1.n178 OUT1.n144 0.0179841
R21471 OUT1.n187 OUT1.n142 0.0177783
R21472 OUT1.n181 OUT1.n144 0.0177304
R21473 OUT1.n176 OUT1.n146 0.0173591
R21474 OUT1.n178 OUT1.n177 0.0173591
R21475 OUT1.n177 OUT1.n176 0.0173591
R21476 OUT1.n173 OUT1.n146 0.0173591
R21477 OUT1.n171 OUT1.n170 0.0172037
R21478 OUT1.n166 OUT1.n163 0.0171032
R21479 OUT1.n185 OUT1.n184 0.0163451
R21480 OUT1.n186 OUT1.n143 0.0163451
R21481 OUT1.n108 OUT1.n98 0.0156875
R21482 OUT1.n246 OUT1.n219 0.0156875
R21483 OUT1.n137 OUT1.n114 0.0156875
R21484 OUT1.n203 OUT1.n196 0.0156875
R21485 OUT1.n215 OUT1.n189 0.0156875
R21486 OUT1.n18 OUT1.n11 0.0156875
R21487 OUT1.n30 OUT1.n4 0.0156875
R21488 OUT1.n251 OUT1.n0 0.014
R21489 OUT1.n96 OUT1.n32 0.014
R21490 OUT1.n175 OUT1.n148 0.0136473
R21491 OUT1 OUT1.n256 0.0135
R21492 OUT1.n253 OUT1.n32 0.0134654
R21493 OUT1.n164 OUT1.n163 0.0128592
R21494 OUT1.n171 OUT1.n152 0.0125423
R21495 OUT1.n174 OUT1.n147 0.0119325
R21496 OUT1.n182 OUT1.n143 0.0112521
R21497 OUT1.n161 OUT1.n154 0.0110972
R21498 OUT1.n180 OUT1.n145 0.0110972
R21499 OUT1.n162 OUT1.n154 0.010845
R21500 OUT1.n180 OUT1.n179 0.010845
R21501 OUT1.n160 OUT1.n159 0.0106136
R21502 OUT1.n184 OUT1.n183 0.00905634
R21503 OUT1.n185 OUT1.n142 0.00905634
R21504 OUT1.n110 OUT1.n98 0.00860784
R21505 OUT1.n224 OUT1.n221 0.00860784
R21506 OUT1.n236 OUT1.n219 0.00860784
R21507 OUT1.n139 OUT1.n114 0.00860784
R21508 OUT1.n198 OUT1.n196 0.00860784
R21509 OUT1.n204 OUT1.n191 0.00860784
R21510 OUT1.n211 OUT1.n189 0.00860784
R21511 OUT1.n13 OUT1.n11 0.00860784
R21512 OUT1.n19 OUT1.n6 0.00860784
R21513 OUT1.n26 OUT1.n4 0.00860784
R21514 OUT1.n232 OUT1.n224 0.00858096
R21515 OUT1.n207 OUT1.n206 0.00858096
R21516 OUT1.n206 OUT1.n204 0.00858096
R21517 OUT1.n22 OUT1.n21 0.00858096
R21518 OUT1.n21 OUT1.n19 0.00858096
R21519 OUT1.n111 OUT1.n110 0.00855417
R21520 OUT1.n234 OUT1.n221 0.00855417
R21521 OUT1.n236 OUT1.n235 0.00855417
R21522 OUT1.n140 OUT1.n139 0.00855417
R21523 OUT1.n209 OUT1.n191 0.00855417
R21524 OUT1.n211 OUT1.n210 0.00855417
R21525 OUT1.n24 OUT1.n6 0.00855417
R21526 OUT1.n26 OUT1.n25 0.00855417
R21527 OUT1.n255 OUT1.n1 0.00773989
R21528 OUT1.n94 OUT1.n31 0.00773989
R21529 OUT1.n92 OUT1.n1 0.00773989
R21530 OUT1.n96 OUT1.n94 0.00773989
R21531 OUT1.n255 OUT1.n2 0.00773989
R21532 OUT1.n254 OUT1.n252 0.00773989
R21533 OUT1.n95 OUT1.n0 0.00773989
R21534 OUT1.n157 OUT1.n151 0.00747183
R21535 OUT1.n148 OUT1.n145 0.00732364
R21536 OUT1.n161 OUT1.n160 0.00580678
R21537 OUT1.n159 OUT1.n153 0.00471334
R21538 OUT1.n172 OUT1.n150 0.00459155
R21539 OUT1.n252 OUT1.n3 0.00374088
R21540 OUT1.n168 OUT1.n153 0.00285636
R21541 OUT1.n168 OUT1.n150 0.00279548
R21542 OUT1.n169 OUT1.n149 0.00165043
R21543 OUT1.n167 OUT1.n151 0.00163371
R21544 a_29248_n7510.t0 a_29248_n7510.t1 6.46072
R21545 a_29248_n7510.t1 a_29248_n7510.t2 6.4095
R21546 a_29248_n7510.n0 a_29248_n7510.t4 2.38861
R21547 a_29248_n7510.n0 a_29248_n7510.t3 2.2505
R21548 a_29248_n7510.t1 a_29248_n7510.n0 5.52236
R21549 IBIAS.t45 IBIAS.t26 49.6666
R21550 IBIAS.t23 IBIAS.t45 49.6666
R21551 IBIAS.t24 IBIAS.t23 49.6666
R21552 IBIAS.t27 IBIAS.t20 49.6666
R21553 IBIAS.t38 IBIAS.t27 49.6666
R21554 IBIAS.t35 IBIAS.t38 49.6666
R21555 IBIAS.t21 IBIAS.t15 49.6666
R21556 IBIAS.t37 IBIAS.t21 49.6666
R21557 IBIAS.t43 IBIAS.t37 49.6666
R21558 IBIAS.t39 IBIAS.t42 49.6666
R21559 IBIAS.t13 IBIAS.t39 49.6666
R21560 IBIAS.t17 IBIAS.t13 49.6666
R21561 IBIAS.t40 IBIAS.t36 49.6666
R21562 IBIAS.t16 IBIAS.t40 49.6666
R21563 IBIAS.t33 IBIAS.t16 49.6666
R21564 IBIAS.t41 IBIAS.t30 49.6666
R21565 IBIAS.t18 IBIAS.t41 49.6666
R21566 IBIAS.t14 IBIAS.t18 49.6666
R21567 IBIAS.t28 IBIAS.t19 49.6666
R21568 IBIAS.t29 IBIAS.t28 49.6666
R21569 IBIAS.t25 IBIAS.t29 49.6666
R21570 IBIAS.t31 IBIAS.t12 49.6666
R21571 IBIAS.t32 IBIAS.t31 49.6666
R21572 IBIAS.t44 IBIAS.t32 49.6666
R21573 IBIAS.n27 IBIAS.t8 45.8862
R21574 IBIAS.n16 IBIAS.t6 39.6291
R21575 IBIAS.n4 IBIAS.t24 35.7835
R21576 IBIAS.n24 IBIAS.t2 31.8076
R21577 IBIAS.n18 IBIAS.t10 31.8076
R21578 IBIAS.n27 IBIAS.t4 31.8076
R21579 IBIAS.n2 IBIAS.t44 22.1612
R21580 IBIAS.n4 IBIAS.t35 21.705
R21581 IBIAS.n5 IBIAS.t43 21.705
R21582 IBIAS.n6 IBIAS.t17 21.705
R21583 IBIAS.n7 IBIAS.t33 21.705
R21584 IBIAS.n8 IBIAS.t14 21.705
R21585 IBIAS.n9 IBIAS.t25 21.705
R21586 IBIAS.n5 IBIAS.n4 14.0791
R21587 IBIAS.n6 IBIAS.n5 14.0791
R21588 IBIAS.n7 IBIAS.n6 14.0791
R21589 IBIAS.n8 IBIAS.n7 14.0791
R21590 IBIAS.n9 IBIAS.n8 14.0791
R21591 IBIAS.n10 IBIAS.n9 6.84425
R21592 IBIAS.n40 IBIAS.n39 6.27404
R21593 IBIAS.n17 IBIAS.t7 4.52093
R21594 IBIAS.n26 IBIAS.n13 4.0005
R21595 IBIAS.n25 IBIAS.n24 4.0005
R21596 IBIAS.n23 IBIAS.n22 4.0005
R21597 IBIAS.n20 IBIAS.n19 4.0005
R21598 IBIAS.n17 IBIAS.n16 4.0005
R21599 IBIAS.n29 IBIAS.n28 4.0005
R21600 IBIAS.n44 IBIAS.n43 3.78325
R21601 IBIAS.n21 IBIAS.n15 3.61985
R21602 IBIAS.n11 IBIAS.n10 2.8805
R21603 IBIAS.n3 IBIAS.n2 2.8805
R21604 IBIAS.n39 IBIAS.t1 1.6385
R21605 IBIAS.n39 IBIAS.n38 1.6385
R21606 IBIAS IBIAS.n52 1.35703
R21607 IBIAS.n36 IBIAS.n35 1.16629
R21608 IBIAS.n32 IBIAS.n31 1.1255
R21609 IBIAS.n35 IBIAS.n34 1.01901
R21610 IBIAS.n50 IBIAS.n48 0.894307
R21611 IBIAS.n42 IBIAS.n37 0.616779
R21612 IBIAS.n48 IBIAS.n12 0.5355
R21613 IBIAS.n28 IBIAS.n27 0.521929
R21614 IBIAS.n19 IBIAS.n18 0.521929
R21615 IBIAS.n30 IBIAS.n29 0.483092
R21616 IBIAS.n15 IBIAS.t3 0.4555
R21617 IBIAS.n15 IBIAS.n14 0.4555
R21618 IBIAS.n34 IBIAS.t9 0.4555
R21619 IBIAS.n34 IBIAS.n33 0.4555
R21620 IBIAS.n29 IBIAS.n26 0.203978
R21621 IBIAS.n26 IBIAS.n25 0.203978
R21622 IBIAS.n25 IBIAS.n23 0.203978
R21623 IBIAS.n20 IBIAS.n17 0.203978
R21624 IBIAS.n21 IBIAS.n20 0.196152
R21625 IBIAS.n37 IBIAS.n32 0.0712285
R21626 IBIAS.n12 IBIAS.n11 0.062564
R21627 IBIAS.n12 IBIAS.n3 0.0620381
R21628 IBIAS.n37 IBIAS.n36 0.0534597
R21629 IBIAS.n51 IBIAS.n50 0.0432108
R21630 IBIAS.n31 IBIAS.n30 0.0324737
R21631 IBIAS.n46 IBIAS.n45 0.0265211
R21632 IBIAS.n43 IBIAS.n42 0.0156875
R21633 IBIAS.n45 IBIAS.n44 0.0137606
R21634 IBIAS.n48 IBIAS.n47 0.013
R21635 IBIAS.n48 IBIAS.n1 0.0125
R21636 IBIAS.n50 IBIAS.n49 0.0115343
R21637 IBIAS.n42 IBIAS.n41 0.00860784
R21638 IBIAS.n41 IBIAS.n40 0.00855417
R21639 IBIAS.n23 IBIAS.n21 0.00832609
R21640 IBIAS.n52 IBIAS.n51 0.00582347
R21641 IBIAS.n1 IBIAS.n0 0.002
R21642 IBIAS.n47 IBIAS.n46 0.0015
R21643 VOUT.n8 VOUT.t4 39.2493
R21644 VOUT.n17 VOUT.t18 39.2493
R21645 VOUT.n23 VOUT.t17 38.6755
R21646 VOUT.n28 VOUT.t9 38.3255
R21647 VOUT.n27 VOUT.t5 38.3255
R21648 VOUT.n14 VOUT.t3 37.8216
R21649 VOUT.n29 VOUT.t26 37.0332
R21650 VOUT.n35 VOUT.t25 36.7201
R21651 VOUT.n6 VOUT.t28 36.5005
R21652 VOUT.n7 VOUT.t30 36.5005
R21653 VOUT.n15 VOUT.t8 36.5005
R21654 VOUT.n16 VOUT.t10 36.5005
R21655 VOUT.n10 VOUT.t29 36.2398
R21656 VOUT.n11 VOUT.t11 36.2398
R21657 VOUT.n19 VOUT.t14 36.2398
R21658 VOUT.n20 VOUT.t22 36.2398
R21659 VOUT.n9 VOUT.t7 34.9362
R21660 VOUT.n12 VOUT.t2 34.9362
R21661 VOUT.n18 VOUT.t19 34.9362
R21662 VOUT.n21 VOUT.t16 34.9362
R21663 VOUT.n31 VOUT.t20 30.113
R21664 VOUT.n32 VOUT.t31 30.113
R21665 VOUT.n33 VOUT.t24 29.0701
R21666 VOUT.n30 VOUT.t27 29.0701
R21667 VOUT.n32 VOUT.n31 20.8576
R21668 VOUT.n31 VOUT.n30 19.8148
R21669 VOUT.n33 VOUT.n32 19.8148
R21670 VOUT.n28 VOUT.t21 17.4684
R21671 VOUT.n27 VOUT.t12 17.4684
R21672 VOUT.n6 VOUT.t6 15.6434
R21673 VOUT.n7 VOUT.t15 15.6434
R21674 VOUT.n15 VOUT.t13 15.6434
R21675 VOUT.n16 VOUT.t23 15.6434
R21676 VOUT.n11 VOUT.n10 14.8868
R21677 VOUT.n20 VOUT.n19 14.8868
R21678 VOUT.n29 VOUT.n28 14.2987
R21679 VOUT.n34 VOUT.n27 14.2987
R21680 VOUT.n10 VOUT.n9 13.9445
R21681 VOUT.n12 VOUT.n11 13.9445
R21682 VOUT.n19 VOUT.n18 13.9445
R21683 VOUT.n21 VOUT.n20 13.9445
R21684 VOUT.n13 VOUT.n6 13.9076
R21685 VOUT.n8 VOUT.n7 13.9076
R21686 VOUT.n22 VOUT.n15 13.9076
R21687 VOUT.n17 VOUT.n16 13.9076
R21688 VOUT VOUT.n0 9.36069
R21689 VOUT.n0 VOUT.t1 7.14109
R21690 VOUT.n36 VOUT.n35 5.09856
R21691 VOUT.n24 VOUT.n23 4.77125
R21692 VOUT.n9 VOUT.n8 4.62659
R21693 VOUT.n18 VOUT.n17 4.62659
R21694 VOUT.n30 VOUT.n29 4.62659
R21695 VOUT.n13 VOUT.n12 4.31354
R21696 VOUT.n22 VOUT.n21 4.31354
R21697 VOUT.n34 VOUT.n33 4.31354
R21698 VOUT.n24 VOUT.n14 4.17447
R21699 VOUT.n0 VOUT.t0 3.4687
R21700 VOUT.n26 VOUT.n5 1.49812
R21701 VOUT.n40 VOUT.n39 1.49801
R21702 VOUT.n43 VOUT.n41 1.49801
R21703 VOUT.n44 VOUT.n43 1.12675
R21704 VOUT.n44 VOUT.n26 1.126
R21705 VOUT.n35 VOUT.n34 0.626587
R21706 VOUT.n23 VOUT.n22 0.623815
R21707 VOUT.n14 VOUT.n13 0.592658
R21708 VOUT.n25 VOUT.n24 0.546814
R21709 VOUT VOUT.n44 0.111701
R21710 VOUT.n5 VOUT.n4 0.0236139
R21711 VOUT.n43 VOUT.n42 0.014
R21712 VOUT.n26 VOUT.n2 0.014
R21713 VOUT.n26 VOUT.n25 0.014
R21714 VOUT.n2 VOUT.n1 0.0134654
R21715 VOUT.n37 VOUT.n36 0.00773989
R21716 VOUT.n39 VOUT.n37 0.00773989
R21717 VOUT.n39 VOUT.n38 0.00773989
R21718 VOUT.n5 VOUT.n3 0.00582347
R21719 VOUT.n43 VOUT.n40 0.00549102
R21720 OUT2.t88 OUT2.t38 122.014
R21721 OUT2.t99 OUT2.t40 122.014
R21722 OUT2.t100 OUT2.t73 122.014
R21723 OUT2.t37 OUT2.t68 122.014
R21724 OUT2.t87 OUT2.t65 122.014
R21725 OUT2.t55 OUT2.t90 122.014
R21726 OUT2.t53 OUT2.t57 122.014
R21727 OUT2.t60 OUT2.t107 122.014
R21728 OUT2.t48 OUT2.t97 122.014
R21729 OUT2.t83 OUT2.t76 122.014
R21730 OUT2.t41 OUT2.t75 122.014
R21731 OUT2.t80 OUT2.t49 122.014
R21732 OUT2.n30 OUT2.t96 63.548
R21733 OUT2.n50 OUT2.t104 63.548
R21734 OUT2.n22 OUT2.t79 63.548
R21735 OUT2.n42 OUT2.t89 63.548
R21736 OUT2.n8 OUT2.t81 63.548
R21737 OUT2.n1 OUT2.t58 63.548
R21738 OUT2.n14 OUT2.t45 62.5719
R21739 OUT2.n15 OUT2.t78 62.5719
R21740 OUT2.n16 OUT2.t101 62.5719
R21741 OUT2.n17 OUT2.t54 62.5719
R21742 OUT2.n33 OUT2.t99 62.5719
R21743 OUT2.n31 OUT2.t66 62.5719
R21744 OUT2.n29 OUT2.t37 62.5719
R21745 OUT2.n47 OUT2.t55 62.5719
R21746 OUT2.n48 OUT2.t85 62.5719
R21747 OUT2.n49 OUT2.t60 62.5719
R21748 OUT2.n25 OUT2.t105 62.5719
R21749 OUT2.n23 OUT2.t44 62.5719
R21750 OUT2.n21 OUT2.t56 62.5719
R21751 OUT2.n39 OUT2.t77 62.5719
R21752 OUT2.n40 OUT2.t67 62.5719
R21753 OUT2.n41 OUT2.t98 62.5719
R21754 OUT2.n18 OUT2.t43 62.5719
R21755 OUT2.n19 OUT2.t84 62.5719
R21756 OUT2.n11 OUT2.t83 62.5719
R21757 OUT2.n9 OUT2.t46 62.5719
R21758 OUT2.n7 OUT2.t80 62.5719
R21759 OUT2.n4 OUT2.t62 62.5719
R21760 OUT2.n2 OUT2.t103 62.5719
R21761 OUT2.n0 OUT2.t39 62.5719
R21762 OUT2.n53 OUT2.t106 61.8074
R21763 OUT2.n45 OUT2.t95 61.8074
R21764 OUT2.n35 OUT2.t92 61.8072
R21765 OUT2.n27 OUT2.t72 61.8072
R21766 OUT2.n13 OUT2.t93 61.8072
R21767 OUT2.n6 OUT2.t74 61.8072
R21768 OUT2.n14 OUT2.t64 41.7148
R21769 OUT2.n15 OUT2.t94 41.7148
R21770 OUT2.n16 OUT2.t50 41.7148
R21771 OUT2.n17 OUT2.t36 41.7148
R21772 OUT2.n33 OUT2.t88 41.7148
R21773 OUT2.n31 OUT2.t91 41.7148
R21774 OUT2.n29 OUT2.t100 41.7148
R21775 OUT2.n47 OUT2.t87 41.7148
R21776 OUT2.n48 OUT2.t82 41.7148
R21777 OUT2.n49 OUT2.t53 41.7148
R21778 OUT2.n25 OUT2.t102 41.7148
R21779 OUT2.n23 OUT2.t69 41.7148
R21780 OUT2.n21 OUT2.t59 41.7148
R21781 OUT2.n39 OUT2.t52 41.7148
R21782 OUT2.n40 OUT2.t63 41.7148
R21783 OUT2.n41 OUT2.t42 41.7148
R21784 OUT2.n18 OUT2.t71 41.7148
R21785 OUT2.n19 OUT2.t47 41.7148
R21786 OUT2.n11 OUT2.t48 41.7148
R21787 OUT2.n9 OUT2.t70 41.7148
R21788 OUT2.n7 OUT2.t41 41.7148
R21789 OUT2.n4 OUT2.t86 41.7148
R21790 OUT2.n2 OUT2.t51 41.7148
R21791 OUT2.n0 OUT2.t61 41.7148
R21792 OUT2.n20 OUT2.n19 17.2118
R21793 OUT2.n34 OUT2.n33 15.9934
R21794 OUT2.n30 OUT2.n29 15.9934
R21795 OUT2.n52 OUT2.n47 15.9934
R21796 OUT2.n50 OUT2.n49 15.9934
R21797 OUT2.n26 OUT2.n25 15.9934
R21798 OUT2.n22 OUT2.n21 15.9934
R21799 OUT2.n44 OUT2.n39 15.9934
R21800 OUT2.n42 OUT2.n41 15.9934
R21801 OUT2.n12 OUT2.n11 15.9934
R21802 OUT2.n8 OUT2.n7 15.9934
R21803 OUT2.n5 OUT2.n4 15.9934
R21804 OUT2.n1 OUT2.n0 15.9934
R21805 OUT2.n57 OUT2.n17 14.8788
R21806 OUT2.n59 OUT2.n15 14.8788
R21807 OUT2.n20 OUT2.n18 14.8786
R21808 OUT2.n58 OUT2.n16 14.8786
R21809 OUT2.n60 OUT2.n14 14.8786
R21810 OUT2.n32 OUT2.n31 13.9076
R21811 OUT2.n51 OUT2.n48 13.9076
R21812 OUT2.n24 OUT2.n23 13.9076
R21813 OUT2.n43 OUT2.n40 13.9076
R21814 OUT2.n10 OUT2.n9 13.9076
R21815 OUT2.n3 OUT2.n2 13.9076
R21816 OUT2 OUT2.n62 8.55615
R21817 OUT2.n59 OUT2.n58 8.51465
R21818 OUT2.n61 OUT2.n60 7.59746
R21819 OUT2.n154 OUT2.t26 6.49823
R21820 OUT2.n154 OUT2.t2 6.4095
R21821 OUT2.n55 OUT2.n46 5.57576
R21822 OUT2.n37 OUT2.n28 5.57576
R21823 OUT2.n62 OUT2.n61 5.57576
R21824 OUT2.n104 OUT2.n103 5.40577
R21825 OUT2.n101 OUT2.t12 5.40577
R21826 OUT2.n100 OUT2.n99 5.40577
R21827 OUT2.n61 OUT2.n13 5.19114
R21828 OUT2.n113 OUT2.t22 5.08295
R21829 OUT2.n95 OUT2.t18 4.9949
R21830 OUT2.n127 OUT2.t1 4.9949
R21831 OUT2.n230 OUT2.n229 4.66184
R21832 OUT2.n212 OUT2.t32 4.66184
R21833 OUT2.n56 OUT2.n55 4.46734
R21834 OUT2.n38 OUT2.n37 4.46734
R21835 OUT2.n97 OUT2.n93 4.36882
R21836 OUT2.n96 OUT2.t17 4.36882
R21837 OUT2.n95 OUT2.n94 4.36882
R21838 OUT2.n128 OUT2.t34 4.36882
R21839 OUT2.n127 OUT2.n126 4.36882
R21840 OUT2.n183 OUT2.n182 4.10662
R21841 OUT2.n225 OUT2.n224 4.08037
R21842 OUT2.n104 OUT2.n102 3.71925
R21843 OUT2.n101 OUT2.t35 3.71925
R21844 OUT2.n100 OUT2.n98 3.71925
R21845 OUT2.n188 OUT2.n187 3.14508
R21846 OUT2.n38 OUT2.n20 3.13062
R21847 OUT2.n57 OUT2.n56 3.12979
R21848 OUT2.n28 OUT2.n27 2.94114
R21849 OUT2.n36 OUT2.n35 2.94114
R21850 OUT2.n46 OUT2.n45 2.94095
R21851 OUT2.n54 OUT2.n53 2.94095
R21852 OUT2.n62 OUT2.n6 2.94051
R21853 OUT2.n153 OUT2.t10 2.4095
R21854 OUT2.n159 OUT2.t24 2.4095
R21855 OUT2.n55 OUT2.n54 2.2505
R21856 OUT2.n37 OUT2.n36 2.2505
R21857 OUT2.n158 OUT2.n153 2.11382
R21858 OUT2.n105 OUT2.n104 1.77702
R21859 OUT2.n129 OUT2.n125 1.76122
R21860 OUT2.n135 OUT2.n131 1.50459
R21861 OUT2.n135 OUT2.n134 1.5025
R21862 OUT2.n253 OUT2.n92 1.49812
R21863 OUT2.n259 OUT2.n258 1.49801
R21864 OUT2.n188 OUT2.n139 1.48953
R21865 OUT2.n210 OUT2.n209 1.48953
R21866 OUT2.n136 OUT2.n121 1.48107
R21867 OUT2.n162 OUT2.n159 1.43397
R21868 OUT2.n129 OUT2.n128 1.34243
R21869 OUT2.n235 OUT2.n234 1.30811
R21870 OUT2.n221 OUT2.n220 1.30811
R21871 OUT2.n216 OUT2.n215 1.30811
R21872 OUT2.n112 OUT2.n111 1.28725
R21873 OUT2.n199 OUT2.n198 1.19489
R21874 OUT2.n58 OUT2.n57 1.18503
R21875 OUT2.n60 OUT2.n59 1.18503
R21876 OUT2.n193 OUT2.n192 1.17841
R21877 OUT2.n72 OUT2.n71 1.16484
R21878 OUT2.n85 OUT2.n84 1.1643
R21879 OUT2.n236 OUT2.n235 1.14175
R21880 OUT2.n222 OUT2.n221 1.14175
R21881 OUT2.n217 OUT2.n216 1.14175
R21882 OUT2.n96 OUT2.n95 1.12746
R21883 OUT2.n128 OUT2.n127 1.12746
R21884 OUT2.n110 OUT2.n109 1.1255
R21885 OUT2.n115 OUT2.n114 1.1255
R21886 OUT2.n232 OUT2.n231 1.1255
R21887 OUT2.n227 OUT2.n226 1.1255
R21888 OUT2.n214 OUT2.n213 1.1255
R21889 OUT2.n131 OUT2.n130 1.1255
R21890 OUT2.n168 OUT2.n167 1.12145
R21891 OUT2.n182 OUT2.n181 1.12145
R21892 OUT2.n177 OUT2.n176 1.11801
R21893 OUT2.n74 OUT2.n73 1.10737
R21894 OUT2.n250 OUT2.n249 1.04129
R21895 OUT2.n84 OUT2.n83 1.00262
R21896 OUT2.n71 OUT2.n70 1.00232
R21897 OUT2.n251 OUT2.n120 0.978961
R21898 OUT2.n260 OUT2.n63 0.917563
R21899 OUT2.n87 OUT2.n86 0.88565
R21900 OUT2.n107 OUT2.n106 0.877022
R21901 OUT2.n252 OUT2.n251 0.857314
R21902 OUT2.n198 OUT2.n197 0.824494
R21903 OUT2.n192 OUT2.n191 0.824494
R21904 OUT2.n187 OUT2.n186 0.767554
R21905 OUT2.n144 OUT2.n143 0.7505
R21906 OUT2.n209 OUT2.n208 0.72825
R21907 OUT2.n243 OUT2.n228 0.727104
R21908 OUT2.n202 OUT2.n200 0.727104
R21909 OUT2.n89 OUT2.n88 0.71475
R21910 OUT2.n105 OUT2.n101 0.650065
R21911 OUT2.n106 OUT2.n100 0.650065
R21912 OUT2.n32 OUT2.n30 0.626587
R21913 OUT2.n34 OUT2.n32 0.626587
R21914 OUT2.n52 OUT2.n51 0.626587
R21915 OUT2.n51 OUT2.n50 0.626587
R21916 OUT2.n24 OUT2.n22 0.626587
R21917 OUT2.n26 OUT2.n24 0.626587
R21918 OUT2.n44 OUT2.n43 0.626587
R21919 OUT2.n43 OUT2.n42 0.626587
R21920 OUT2.n10 OUT2.n8 0.626587
R21921 OUT2.n12 OUT2.n10 0.626587
R21922 OUT2.n3 OUT2.n1 0.626587
R21923 OUT2.n5 OUT2.n3 0.626587
R21924 OUT2.n97 OUT2.n96 0.626587
R21925 OUT2.n106 OUT2.n105 0.626587
R21926 OUT2.n118 OUT2.n116 0.616779
R21927 OUT2.n239 OUT2.n237 0.616779
R21928 OUT2.n248 OUT2.n218 0.616779
R21929 OUT2.n207 OUT2.n194 0.616779
R21930 OUT2.n70 OUT2.t31 0.58197
R21931 OUT2.n70 OUT2.n69 0.58197
R21932 OUT2.n83 OUT2.t25 0.58197
R21933 OUT2.n83 OUT2.n82 0.58197
R21934 OUT2.n234 OUT2.n233 0.58197
R21935 OUT2.n224 OUT2.t5 0.58197
R21936 OUT2.n224 OUT2.n223 0.58197
R21937 OUT2.n220 OUT2.t6 0.58197
R21938 OUT2.n220 OUT2.n219 0.58197
R21939 OUT2.n215 OUT2.t28 0.58197
R21940 OUT2.n197 OUT2.t7 0.58197
R21941 OUT2.n197 OUT2.n196 0.58197
R21942 OUT2.n191 OUT2.t27 0.58197
R21943 OUT2.n191 OUT2.n190 0.58197
R21944 OUT2.n111 OUT2.t21 0.56925
R21945 OUT2.n125 OUT2.n124 0.56925
R21946 OUT2.n250 OUT2.n211 0.553805
R21947 OUT2.n108 OUT2.n107 0.532674
R21948 OUT2.n138 OUT2.n137 0.4875
R21949 OUT2.n56 OUT2.n38 0.475368
R21950 OUT2.n77 OUT2.n76 0.474125
R21951 OUT2.n241 OUT2.n240 0.474125
R21952 OUT2.n246 OUT2.n245 0.474125
R21953 OUT2.n205 OUT2.n204 0.474125
R21954 OUT2.n6 OUT2.n5 0.279824
R21955 OUT2.n35 OUT2.n34 0.279823
R21956 OUT2.n27 OUT2.n26 0.279823
R21957 OUT2.n13 OUT2.n12 0.279823
R21958 OUT2.n53 OUT2.n52 0.279615
R21959 OUT2.n45 OUT2.n44 0.279615
R21960 OUT2.n251 OUT2.n250 0.264618
R21961 OUT2.n114 OUT2.n113 0.239196
R21962 OUT2.n107 OUT2.n97 0.207891
R21963 OUT2.n176 OUT2.n175 0.203732
R21964 OUT2.n130 OUT2.n129 0.19908
R21965 OUT2.n109 OUT2.n108 0.190283
R21966 OUT2.n186 OUT2.n185 0.147906
R21967 OUT2 OUT2.n262 0.0999375
R21968 OUT2.n86 OUT2.n80 0.0936537
R21969 OUT2.n130 OUT2.n123 0.0935118
R21970 OUT2.n73 OUT2.n67 0.0880141
R21971 OUT2.n228 OUT2.n222 0.0823987
R21972 OUT2.n200 OUT2.n195 0.0823987
R21973 OUT2.n71 OUT2.n68 0.0790912
R21974 OUT2.n84 OUT2.n81 0.0786471
R21975 OUT2.n116 OUT2.n110 0.0712285
R21976 OUT2.n218 OUT2.n214 0.0712285
R21977 OUT2.n237 OUT2.n232 0.0712285
R21978 OUT2.n194 OUT2.n189 0.0712285
R21979 OUT2.n155 OUT2.n154 0.0603944
R21980 OUT2.n114 OUT2.n112 0.0568678
R21981 OUT2.n116 OUT2.n115 0.0534597
R21982 OUT2.n237 OUT2.n236 0.0534597
R21983 OUT2.n218 OUT2.n217 0.0534597
R21984 OUT2.n194 OUT2.n193 0.0534597
R21985 OUT2.n228 OUT2.n227 0.0415773
R21986 OUT2.n200 OUT2.n199 0.0415773
R21987 OUT2.n210 OUT2.n188 0.0354016
R21988 OUT2.n187 OUT2.n144 0.0334577
R21989 OUT2.n73 OUT2.n72 0.0319869
R21990 OUT2.n166 OUT2.n165 0.0296151
R21991 OUT2.n86 OUT2.n85 0.0261793
R21992 OUT2.n167 OUT2.n158 0.0241583
R21993 OUT2.n123 OUT2.n122 0.0230949
R21994 OUT2.n257 OUT2.n256 0.0229474
R21995 OUT2.n259 OUT2.n255 0.0229474
R21996 OUT2.n147 OUT2.n146 0.0228651
R21997 OUT2.n165 OUT2.n164 0.0210986
R21998 OUT2.n231 OUT2.n230 0.0201463
R21999 OUT2.n226 OUT2.n225 0.0201463
R22000 OUT2.n213 OUT2.n212 0.0201463
R22001 OUT2.n162 OUT2.n161 0.0195995
R22002 OUT2.n139 OUT2.n138 0.0182008
R22003 OUT2.n211 OUT2.n210 0.0182008
R22004 OUT2.n177 OUT2.n151 0.0179841
R22005 OUT2.n182 OUT2.n177 0.0177304
R22006 OUT2.n149 OUT2.n148 0.0173591
R22007 OUT2.n151 OUT2.n150 0.0173591
R22008 OUT2.n150 OUT2.n149 0.0173591
R22009 OUT2.n148 OUT2.n147 0.0173591
R22010 OUT2.n163 OUT2.n162 0.0171032
R22011 OUT2.n142 OUT2.n141 0.0163451
R22012 OUT2.n185 OUT2.n184 0.0163451
R22013 OUT2.n87 OUT2.n77 0.0156875
R22014 OUT2.n88 OUT2.n87 0.0156875
R22015 OUT2.n118 OUT2.n117 0.0156875
R22016 OUT2.n240 OUT2.n239 0.0156875
R22017 OUT2.n249 OUT2.n248 0.0156875
R22018 OUT2.n137 OUT2.n136 0.0156875
R22019 OUT2.n208 OUT2.n207 0.0156875
R22020 OUT2.n254 OUT2.n253 0.014
R22021 OUT2.n253 OUT2.n252 0.014
R22022 OUT2.n255 OUT2.n254 0.0134654
R22023 OUT2.n66 OUT2.n65 0.0133659
R22024 OUT2.n164 OUT2.n163 0.0128592
R22025 OUT2.n134 OUT2.n132 0.012194
R22026 OUT2.n146 OUT2.n145 0.0119325
R22027 OUT2.n158 OUT2.n157 0.011782
R22028 OUT2.n184 OUT2.n183 0.0112521
R22029 OUT2.n76 OUT2.n75 0.0111023
R22030 OUT2.n169 OUT2.n168 0.0110972
R22031 OUT2.n181 OUT2.n179 0.0110972
R22032 OUT2.n168 OUT2.n152 0.010845
R22033 OUT2.n181 OUT2.n180 0.010845
R22034 OUT2.n171 OUT2.n170 0.0106136
R22035 OUT2.n141 OUT2.n140 0.00905634
R22036 OUT2.n143 OUT2.n142 0.00905634
R22037 OUT2.n134 OUT2.n133 0.00878947
R22038 OUT2.n74 OUT2.n64 0.00860784
R22039 OUT2.n119 OUT2.n118 0.00860784
R22040 OUT2.n239 OUT2.n238 0.00860784
R22041 OUT2.n244 OUT2.n243 0.00860784
R22042 OUT2.n248 OUT2.n247 0.00860784
R22043 OUT2.n203 OUT2.n202 0.00860784
R22044 OUT2.n207 OUT2.n206 0.00860784
R22045 OUT2.n242 OUT2.n241 0.00858096
R22046 OUT2.n243 OUT2.n242 0.00858096
R22047 OUT2.n202 OUT2.n201 0.00858096
R22048 OUT2.n120 OUT2.n119 0.00855417
R22049 OUT2.n245 OUT2.n244 0.00855417
R22050 OUT2.n247 OUT2.n246 0.00855417
R22051 OUT2.n204 OUT2.n203 0.00855417
R22052 OUT2.n206 OUT2.n205 0.00855417
R22053 OUT2.n156 OUT2.n155 0.00778873
R22054 OUT2.n91 OUT2.n90 0.00773989
R22055 OUT2.n262 OUT2.n261 0.00773989
R22056 OUT2.n90 OUT2.n89 0.00773989
R22057 OUT2.n261 OUT2.n260 0.00773989
R22058 OUT2.n179 OUT2.n178 0.00732364
R22059 OUT2.n67 OUT2.n66 0.00642105
R22060 OUT2.n80 OUT2.n79 0.00642105
R22061 OUT2.n75 OUT2.n74 0.00605114
R22062 OUT2.n92 OUT2.n91 0.00582347
R22063 OUT2.n170 OUT2.n169 0.00580678
R22064 OUT2.n79 OUT2.n78 0.00551512
R22065 OUT2.n258 OUT2.n257 0.00549102
R22066 OUT2.n260 OUT2.n259 0.00549102
R22067 OUT2.n167 OUT2.n166 0.00533104
R22068 OUT2.n172 OUT2.n171 0.00471334
R22069 OUT2.n174 OUT2.n173 0.00319575
R22070 OUT2.n175 OUT2.n174 0.00319235
R22071 OUT2.n136 OUT2.n135 0.00318273
R22072 OUT2.n173 OUT2.n172 0.00285636
R22073 OUT2.n161 OUT2.n160 0.00163371
R22074 OUT2.n157 OUT2.n156 0.0014753
R22075 IBS.n2 IBS.t9 15.4765
R22076 IBS.n3 IBS.n2 11.0965
R22077 IBS IBS.n26 7.19841
R22078 IBS.n1 IBS.t2 7.191
R22079 IBS.n14 IBS.t8 4.76941
R22080 IBS.n4 IBS.n3 4.49
R22081 IBS.n2 IBS.t10 4.3805
R22082 IBS.n3 IBS.t0 4.3805
R22083 IBS.n14 IBS.n13 3.4692
R22084 IBS.n8 IBS.n7 3.42896
R22085 IBS.n15 IBS.n14 1.82057
R22086 IBS.n21 IBS.n20 1.63898
R22087 IBS.n7 IBS.t3 1.6385
R22088 IBS.n7 IBS.n6 1.6385
R22089 IBS IBS.n11 1.61193
R22090 IBS.n22 IBS.n21 1.14573
R22091 IBS.n5 IBS.n4 1.14565
R22092 IBS.n5 IBS.n1 1.14531
R22093 IBS.n23 IBS.n22 1.12717
R22094 IBS.n17 IBS.n16 1.1255
R22095 IBS.n9 IBS.n5 0.869271
R22096 IBS.n20 IBS.t6 0.4555
R22097 IBS.n20 IBS.n19 0.4555
R22098 IBS.n13 IBS.t7 0.4555
R22099 IBS.n13 IBS.n12 0.4555
R22100 IBS.n16 IBS.n15 0.324453
R22101 IBS.n11 IBS.n10 0.220997
R22102 IBS.n22 IBS.n18 0.0832399
R22103 IBS.n18 IBS.n17 0.0419676
R22104 IBS.n10 IBS.n9 0.0269958
R22105 IBS.n10 IBS.n0 0.0263488
R22106 IBS.n9 IBS.n8 0.013
R22107 IBS.n25 IBS.n24 0.00860784
R22108 IBS.n26 IBS.n25 0.00855417
R22109 IBS.n24 IBS.n23 0.00364318
R22110 IPD.n355 IPD.n354 5.29686
R22111 IPD.n336 IPD.t12 5.29686
R22112 IPD.n221 IPD.n220 4.97729
R22113 IPD.n202 IPD.t48 4.97729
R22114 IPD.n91 IPD.n90 4.86858
R22115 IPD.n342 IPD.n341 4.72811
R22116 IPD.n106 IPD.n105 4.71629
R22117 IPD.n208 IPD.n207 4.40854
R22118 IPD.n331 IPD.n330 2.41042
R22119 IPD.n405 IPD.n403 1.6654
R22120 IPD.n430 IPD.t10 1.6654
R22121 IPD.n87 IPD.n86 1.64142
R22122 IPD.n53 IPD.n49 1.49801
R22123 IPD.n25 IPD.n24 1.49801
R22124 IPD.n283 IPD.n282 1.48953
R22125 IPD.n375 IPD.n84 1.48953
R22126 IPD.n397 IPD.n396 1.48953
R22127 IPD.n196 IPD.n195 1.47785
R22128 IPD.n185 IPD.t27 1.47785
R22129 IPD.n257 IPD.t59 1.31982
R22130 IPD.n253 IPD.n252 1.31982
R22131 IPD.n60 IPD.t45 1.30711
R22132 IPD.n56 IPD.n55 1.30711
R22133 IPD.n352 IPD.n351 1.28973
R22134 IPD.n347 IPD.n346 1.28973
R22135 IPD.n334 IPD.n333 1.28973
R22136 IPD.n192 IPD.n191 1.19571
R22137 IPD.n386 IPD.n385 1.19534
R22138 IPD.n38 IPD.n37 1.19519
R22139 IPD.n72 IPD.n71 1.19509
R22140 IPD.n61 IPD.n60 1.19506
R22141 IPD.n125 IPD.n124 1.19466
R22142 IPD.n13 IPD.n12 1.19457
R22143 IPD.n315 IPD.n314 1.19444
R22144 IPD.n269 IPD.n268 1.19395
R22145 IPD.n258 IPD.n257 1.19393
R22146 IPD.n103 IPD.n102 1.18349
R22147 IPD.n321 IPD.n320 1.17941
R22148 IPD.n176 IPD.n175 1.17929
R22149 IPD.n165 IPD.n164 1.17902
R22150 IPD.n6 IPD.n5 1.17902
R22151 IPD.n119 IPD.n118 1.17891
R22152 IPD.n254 IPD.n253 1.1787
R22153 IPD.n380 IPD.n379 1.1782
R22154 IPD.n197 IPD.n196 1.17812
R22155 IPD.n186 IPD.n185 1.17812
R22156 IPD.n32 IPD.n31 1.17768
R22157 IPD.n57 IPD.n56 1.17753
R22158 IPD.n439 IPD.n438 1.1775
R22159 IPD.n353 IPD.n352 1.17428
R22160 IPD.n348 IPD.n347 1.17428
R22161 IPD.n335 IPD.n334 1.17428
R22162 IPD.n421 IPD.n420 1.16675
R22163 IPD.n219 IPD.n218 1.16619
R22164 IPD.n214 IPD.n213 1.16619
R22165 IPD.n201 IPD.n200 1.16619
R22166 IPD.n293 IPD.n292 1.16617
R22167 IPD.n406 IPD.n405 1.16588
R22168 IPD.n431 IPD.n430 1.16588
R22169 IPD.n135 IPD.n134 1.16562
R22170 IPD.n306 IPD.n305 1.1656
R22171 IPD.n148 IPD.n147 1.16506
R22172 IPD.n374 IPD.n114 1.1515
R22173 IPD.n88 IPD.n87 1.14576
R22174 IPD.n14 IPD.n13 1.12717
R22175 IPD.n422 IPD.n421 1.1257
R22176 IPD.n93 IPD.n92 1.1255
R22177 IPD.n108 IPD.n107 1.1255
R22178 IPD.n357 IPD.n356 1.1255
R22179 IPD.n338 IPD.n337 1.1255
R22180 IPD.n344 IPD.n343 1.1255
R22181 IPD.n223 IPD.n222 1.1255
R22182 IPD.n210 IPD.n209 1.1255
R22183 IPD.n204 IPD.n203 1.1255
R22184 IPD.n373 IPD.n372 1.1255
R22185 IPD.n439 IPD.n53 1.1255
R22186 IPD.n295 IPD.n294 1.10737
R22187 IPD.n137 IPD.n136 1.10737
R22188 IPD.n408 IPD.n407 1.1073
R22189 IPD.n433 IPD.n432 1.1073
R22190 IPD.n147 IPD.n146 1.09806
R22191 IPD.n134 IPD.n133 1.09777
R22192 IPD.n305 IPD.n304 1.09692
R22193 IPD.n292 IPD.n291 1.09663
R22194 IPD.n420 IPD.n418 1.09644
R22195 IPD.n310 IPD.n309 1.08123
R22196 IPD.n218 IPD.n217 1.07378
R22197 IPD.n213 IPD.n212 1.07378
R22198 IPD.n200 IPD.n199 1.07378
R22199 IPD.n152 IPD.n151 0.939312
R22200 IPD.n124 IPD.n123 0.922529
R22201 IPD.n118 IPD.n117 0.922508
R22202 IPD.n320 IPD.n319 0.920678
R22203 IPD.n314 IPD.n313 0.920678
R22204 IPD.n385 IPD.n384 0.913532
R22205 IPD.n379 IPD.n378 0.913527
R22206 IPD.n37 IPD.n36 0.911021
R22207 IPD.n31 IPD.n30 0.911021
R22208 IPD.n191 IPD.n190 0.909101
R22209 IPD.n436 IPD.n435 0.901232
R22210 IPD.n308 IPD.n307 0.88565
R22211 IPD.n150 IPD.n149 0.88565
R22212 IPD.n175 IPD.n174 0.834379
R22213 IPD.n164 IPD.n163 0.834365
R22214 IPD.n5 IPD.n4 0.834365
R22215 IPD.n12 IPD.n11 0.834365
R22216 IPD.n268 IPD.n267 0.834193
R22217 IPD.n71 IPD.n70 0.821487
R22218 IPD.n75 IPD.n74 0.727916
R22219 IPD.n111 IPD.n110 0.727916
R22220 IPD.n272 IPD.n271 0.727916
R22221 IPD.n179 IPD.n178 0.727916
R22222 IPD.n80 IPD.n58 0.727104
R22223 IPD.n389 IPD.n387 0.727104
R22224 IPD.n364 IPD.n349 0.727104
R22225 IPD.n324 IPD.n322 0.727104
R22226 IPD.n277 IPD.n255 0.727104
R22227 IPD.n226 IPD.n224 0.727104
R22228 IPD.n235 IPD.n205 0.727104
R22229 IPD.n244 IPD.n193 0.727104
R22230 IPD.n154 IPD.n126 0.727104
R22231 IPD.n45 IPD.n33 0.727104
R22232 IPD.n183 IPD.n182 0.691748
R22233 IPD.n182 IPD.n181 0.648341
R22234 IPD.n332 IPD.n331 0.632522
R22235 IPD.n22 IPD.n21 0.628687
R22236 IPD.n114 IPD.n113 0.623188
R22237 IPD.n64 IPD.n62 0.616779
R22238 IPD.n394 IPD.n381 0.616779
R22239 IPD.n96 IPD.n94 0.616779
R22240 IPD.n360 IPD.n358 0.616779
R22241 IPD.n369 IPD.n339 0.616779
R22242 IPD.n329 IPD.n316 0.616779
R22243 IPD.n261 IPD.n259 0.616779
R22244 IPD.n231 IPD.n215 0.616779
R22245 IPD.n240 IPD.n198 0.616779
R22246 IPD.n249 IPD.n187 0.616779
R22247 IPD.n168 IPD.n166 0.616779
R22248 IPD.n159 IPD.n120 0.616779
R22249 IPD.n19 IPD.n7 0.616779
R22250 IPD.n41 IPD.n39 0.616779
R22251 IPD.n418 IPD.t31 0.56925
R22252 IPD.n418 IPD.n417 0.56925
R22253 IPD.n384 IPD.t20 0.56925
R22254 IPD.n384 IPD.n383 0.56925
R22255 IPD.n378 IPD.t14 0.56925
R22256 IPD.n378 IPD.n377 0.56925
R22257 IPD.n351 IPD.n350 0.56925
R22258 IPD.n346 IPD.t26 0.56925
R22259 IPD.n346 IPD.n345 0.56925
R22260 IPD.n341 IPD.t32 0.56925
R22261 IPD.n341 IPD.n340 0.56925
R22262 IPD.n333 IPD.t5 0.56925
R22263 IPD.n319 IPD.t56 0.56925
R22264 IPD.n319 IPD.n318 0.56925
R22265 IPD.n313 IPD.t42 0.56925
R22266 IPD.n313 IPD.n312 0.56925
R22267 IPD.n291 IPD.t11 0.56925
R22268 IPD.n291 IPD.n290 0.56925
R22269 IPD.n304 IPD.t7 0.56925
R22270 IPD.n304 IPD.n303 0.56925
R22271 IPD.n217 IPD.n216 0.56925
R22272 IPD.n207 IPD.t38 0.56925
R22273 IPD.n207 IPD.n206 0.56925
R22274 IPD.n212 IPD.t36 0.56925
R22275 IPD.n212 IPD.n211 0.56925
R22276 IPD.n199 IPD.t57 0.56925
R22277 IPD.n190 IPD.t18 0.56925
R22278 IPD.n190 IPD.n189 0.56925
R22279 IPD.n133 IPD.t43 0.56925
R22280 IPD.n133 IPD.n132 0.56925
R22281 IPD.n146 IPD.t69 0.56925
R22282 IPD.n146 IPD.n145 0.56925
R22283 IPD.n123 IPD.t28 0.56925
R22284 IPD.n123 IPD.n122 0.56925
R22285 IPD.n117 IPD.t8 0.56925
R22286 IPD.n117 IPD.n116 0.56925
R22287 IPD.n36 IPD.t23 0.56925
R22288 IPD.n36 IPD.n35 0.56925
R22289 IPD.n30 IPD.t15 0.56925
R22290 IPD.n30 IPD.n29 0.56925
R22291 IPD.n310 IPD.n284 0.526243
R22292 IPD.n182 IPD.n160 0.524913
R22293 IPD.n396 IPD.n395 0.516188
R22294 IPD.n238 IPD.n237 0.507313
R22295 IPD.n48 IPD.n47 0.502687
R22296 IPD.n437 IPD.n436 0.500334
R22297 IPD.n70 IPD.t39 0.485833
R22298 IPD.n70 IPD.n69 0.485833
R22299 IPD.n86 IPD.t33 0.485833
R22300 IPD.n86 IPD.n85 0.485833
R22301 IPD.n90 IPD.t40 0.485833
R22302 IPD.n90 IPD.n89 0.485833
R22303 IPD.n102 IPD.t51 0.485833
R22304 IPD.n102 IPD.n101 0.485833
R22305 IPD.n105 IPD.t66 0.485833
R22306 IPD.n105 IPD.n104 0.485833
R22307 IPD.n267 IPD.t65 0.485833
R22308 IPD.n267 IPD.n266 0.485833
R22309 IPD.n163 IPD.t60 0.485833
R22310 IPD.n163 IPD.n162 0.485833
R22311 IPD.n174 IPD.t64 0.485833
R22312 IPD.n174 IPD.n173 0.485833
R22313 IPD.n4 IPD.t67 0.485833
R22314 IPD.n4 IPD.n3 0.485833
R22315 IPD.n11 IPD.t54 0.485833
R22316 IPD.n11 IPD.n10 0.485833
R22317 IPD.n327 IPD.n326 0.474125
R22318 IPD.n229 IPD.n228 0.474125
R22319 IPD.n233 IPD.n232 0.474125
R22320 IPD.n140 IPD.n139 0.474125
R22321 IPD.n83 IPD.n82 0.46275
R22322 IPD.n280 IPD.n279 0.46275
R22323 IPD.n107 IPD.n106 0.447377
R22324 IPD.n375 IPD.n374 0.352375
R22325 IPD.n282 IPD.n250 0.336187
R22326 IPD.n99 IPD.n98 0.330687
R22327 IPD.n171 IPD.n170 0.330687
R22328 IPD.n18 IPD.n17 0.330687
R22329 IPD.n411 IPD.n410 0.330125
R22330 IPD.n424 IPD.n423 0.330125
R22331 IPD.n78 IPD.n77 0.330125
R22332 IPD.n67 IPD.n66 0.330125
R22333 IPD.n392 IPD.n391 0.330125
R22334 IPD.n362 IPD.n361 0.330125
R22335 IPD.n367 IPD.n366 0.330125
R22336 IPD.n298 IPD.n297 0.330125
R22337 IPD.n275 IPD.n274 0.330125
R22338 IPD.n264 IPD.n263 0.330125
R22339 IPD.n242 IPD.n241 0.330125
R22340 IPD.n247 IPD.n246 0.330125
R22341 IPD.n157 IPD.n156 0.330125
R22342 IPD.n43 IPD.n42 0.330125
R22343 IPD.n371 IPD.n370 0.317187
R22344 IPD.n92 IPD.n91 0.269474
R22345 IPD.n436 IPD.n398 0.268618
R22346 IPD.n331 IPD.n310 0.248389
R22347 IPD IPD.n439 0.241687
R22348 IPD.n356 IPD.n355 0.235932
R22349 IPD.n343 IPD.n342 0.235932
R22350 IPD.n337 IPD.n336 0.235932
R22351 IPD.n222 IPD.n221 0.12963
R22352 IPD.n209 IPD.n208 0.12963
R22353 IPD.n203 IPD.n202 0.12963
R22354 IPD.n307 IPD.n301 0.0936537
R22355 IPD.n149 IPD.n143 0.0912853
R22356 IPD.n407 IPD.n402 0.0886741
R22357 IPD.n432 IPD.n428 0.0886741
R22358 IPD.n294 IPD.n288 0.0880141
R22359 IPD.n136 IPD.n130 0.0856456
R22360 IPD.n13 IPD.n9 0.0832399
R22361 IPD.n74 IPD.n73 0.0826464
R22362 IPD.n110 IPD.n109 0.0826464
R22363 IPD.n271 IPD.n270 0.0826464
R22364 IPD.n178 IPD.n177 0.0826464
R22365 IPD.n58 IPD.n54 0.0823987
R22366 IPD.n387 IPD.n382 0.0823987
R22367 IPD.n349 IPD.n344 0.0823987
R22368 IPD.n322 IPD.n317 0.0823987
R22369 IPD.n255 IPD.n251 0.0823987
R22370 IPD.n224 IPD.n219 0.0823987
R22371 IPD.n205 IPD.n201 0.0823987
R22372 IPD.n193 IPD.n188 0.0823987
R22373 IPD.n126 IPD.n121 0.0823987
R22374 IPD.n33 IPD.n28 0.0823987
R22375 IPD.n420 IPD.n419 0.0784141
R22376 IPD.n405 IPD.n404 0.0783056
R22377 IPD.n430 IPD.n429 0.0783056
R22378 IPD.n292 IPD.n289 0.0778549
R22379 IPD.n305 IPD.n302 0.0774429
R22380 IPD.n107 IPD.n103 0.0761444
R22381 IPD.n134 IPD.n131 0.0761073
R22382 IPD.n147 IPD.n144 0.0756955
R22383 IPD.n62 IPD.n59 0.0712285
R22384 IPD.n381 IPD.n376 0.0712285
R22385 IPD.n94 IPD.n88 0.0712285
R22386 IPD.n339 IPD.n335 0.0712285
R22387 IPD.n358 IPD.n353 0.0712285
R22388 IPD.n316 IPD.n311 0.0712285
R22389 IPD.n259 IPD.n256 0.0712285
R22390 IPD.n187 IPD.n184 0.0712285
R22391 IPD.n198 IPD.n194 0.0712285
R22392 IPD.n215 IPD.n210 0.0712285
R22393 IPD.n166 IPD.n161 0.0712285
R22394 IPD.n120 IPD.n115 0.0712285
R22395 IPD.n7 IPD.n2 0.0712285
R22396 IPD.n39 IPD.n34 0.0712285
R22397 IPD.n421 IPD.n416 0.0623855
R22398 IPD.n416 IPD.n415 0.0576486
R22399 IPD.n62 IPD.n61 0.0534597
R22400 IPD.n381 IPD.n380 0.0534597
R22401 IPD.n94 IPD.n93 0.0534597
R22402 IPD.n358 IPD.n357 0.0534597
R22403 IPD.n339 IPD.n338 0.0534597
R22404 IPD.n316 IPD.n315 0.0534597
R22405 IPD.n259 IPD.n258 0.0534597
R22406 IPD.n215 IPD.n214 0.0534597
R22407 IPD.n198 IPD.n197 0.0534597
R22408 IPD.n187 IPD.n186 0.0534597
R22409 IPD.n166 IPD.n165 0.0534597
R22410 IPD.n120 IPD.n119 0.0534597
R22411 IPD.n7 IPD.n6 0.0534597
R22412 IPD.n39 IPD.n38 0.0534597
R22413 IPD.n374 IPD.n373 0.0525
R22414 IPD.n373 IPD.n332 0.0525
R22415 IPD.n74 IPD.n72 0.0423164
R22416 IPD.n110 IPD.n108 0.0423164
R22417 IPD.n271 IPD.n269 0.0423164
R22418 IPD.n178 IPD.n176 0.0423164
R22419 IPD.n9 IPD.n8 0.0419676
R22420 IPD.n58 IPD.n57 0.0415773
R22421 IPD.n387 IPD.n386 0.0415773
R22422 IPD.n349 IPD.n348 0.0415773
R22423 IPD.n322 IPD.n321 0.0415773
R22424 IPD.n255 IPD.n254 0.0415773
R22425 IPD.n193 IPD.n192 0.0415773
R22426 IPD.n205 IPD.n204 0.0415773
R22427 IPD.n224 IPD.n223 0.0415773
R22428 IPD.n126 IPD.n125 0.0415773
R22429 IPD.n33 IPD.n32 0.0415773
R22430 IPD.n282 IPD.n281 0.0354016
R22431 IPD.n283 IPD.n183 0.0354016
R22432 IPD.n397 IPD.n375 0.0354016
R22433 IPD.n432 IPD.n431 0.032498
R22434 IPD.n407 IPD.n406 0.032498
R22435 IPD.n294 IPD.n293 0.0319869
R22436 IPD.n136 IPD.n135 0.0319869
R22437 IPD.n372 IPD.n371 0.0265
R22438 IPD.n307 IPD.n306 0.0261793
R22439 IPD.n149 IPD.n148 0.0261793
R22440 IPD.n51 IPD.n50 0.0207053
R22441 IPD.n1 IPD.n0 0.0207053
R22442 IPD.n84 IPD.n83 0.0182008
R22443 IPD.n281 IPD.n280 0.0182008
R22444 IPD.n284 IPD.n283 0.0182008
R22445 IPD.n398 IPD.n397 0.0182008
R22446 IPD.n412 IPD.n411 0.0156875
R22447 IPD.n64 IPD.n63 0.0156875
R22448 IPD.n395 IPD.n394 0.0156875
R22449 IPD.n96 IPD.n95 0.0156875
R22450 IPD.n361 IPD.n360 0.0156875
R22451 IPD.n370 IPD.n369 0.0156875
R22452 IPD.n330 IPD.n329 0.0156875
R22453 IPD.n308 IPD.n298 0.0156875
R22454 IPD.n309 IPD.n308 0.0156875
R22455 IPD.n261 IPD.n260 0.0156875
R22456 IPD.n232 IPD.n231 0.0156875
R22457 IPD.n241 IPD.n240 0.0156875
R22458 IPD.n250 IPD.n249 0.0156875
R22459 IPD.n168 IPD.n167 0.0156875
R22460 IPD.n150 IPD.n140 0.0156875
R22461 IPD.n151 IPD.n150 0.0156875
R22462 IPD.n160 IPD.n159 0.0156875
R22463 IPD.n19 IPD.n18 0.0156875
R22464 IPD.n42 IPD.n41 0.0156875
R22465 IPD.n53 IPD.n52 0.014
R22466 IPD.n438 IPD.n437 0.014
R22467 IPD.n427 IPD.n426 0.0139513
R22468 IPD.n401 IPD.n400 0.0139513
R22469 IPD.n52 IPD.n51 0.0134654
R22470 IPD.n287 IPD.n286 0.0133659
R22471 IPD.n423 IPD.n422 0.0123533
R22472 IPD.n129 IPD.n128 0.012194
R22473 IPD.n410 IPD.n409 0.0111023
R22474 IPD.n435 IPD.n434 0.0111023
R22475 IPD.n297 IPD.n296 0.0111023
R22476 IPD.n139 IPD.n138 0.0111023
R22477 IPD.n49 IPD.n48 0.00998204
R22478 IPD.n130 IPD.n129 0.00878947
R22479 IPD.n143 IPD.n142 0.00878947
R22480 IPD.n408 IPD.n399 0.00860784
R22481 IPD.n433 IPD.n425 0.00860784
R22482 IPD.n65 IPD.n64 0.00860784
R22483 IPD.n80 IPD.n79 0.00860784
R22484 IPD.n390 IPD.n389 0.00860784
R22485 IPD.n394 IPD.n393 0.00860784
R22486 IPD.n97 IPD.n96 0.00860784
R22487 IPD.n360 IPD.n359 0.00860784
R22488 IPD.n365 IPD.n364 0.00860784
R22489 IPD.n369 IPD.n368 0.00860784
R22490 IPD.n325 IPD.n324 0.00860784
R22491 IPD.n329 IPD.n328 0.00860784
R22492 IPD.n295 IPD.n285 0.00860784
R22493 IPD.n262 IPD.n261 0.00860784
R22494 IPD.n277 IPD.n276 0.00860784
R22495 IPD.n227 IPD.n226 0.00860784
R22496 IPD.n231 IPD.n230 0.00860784
R22497 IPD.n236 IPD.n235 0.00860784
R22498 IPD.n240 IPD.n239 0.00860784
R22499 IPD.n245 IPD.n244 0.00860784
R22500 IPD.n249 IPD.n248 0.00860784
R22501 IPD.n169 IPD.n168 0.00860784
R22502 IPD.n137 IPD.n127 0.00860784
R22503 IPD.n155 IPD.n154 0.00860784
R22504 IPD.n159 IPD.n158 0.00860784
R22505 IPD.n20 IPD.n19 0.00860784
R22506 IPD.n16 IPD.n15 0.00860784
R22507 IPD.n41 IPD.n40 0.00860784
R22508 IPD.n46 IPD.n45 0.00860784
R22509 IPD.n82 IPD.n81 0.00858096
R22510 IPD.n76 IPD.n75 0.00858096
R22511 IPD.n68 IPD.n67 0.00858096
R22512 IPD.n81 IPD.n80 0.00858096
R22513 IPD.n77 IPD.n76 0.00858096
R22514 IPD.n75 IPD.n68 0.00858096
R22515 IPD.n389 IPD.n388 0.00858096
R22516 IPD.n112 IPD.n111 0.00858096
R22517 IPD.n100 IPD.n99 0.00858096
R22518 IPD.n113 IPD.n112 0.00858096
R22519 IPD.n111 IPD.n100 0.00858096
R22520 IPD.n363 IPD.n362 0.00858096
R22521 IPD.n364 IPD.n363 0.00858096
R22522 IPD.n324 IPD.n323 0.00858096
R22523 IPD.n279 IPD.n278 0.00858096
R22524 IPD.n273 IPD.n272 0.00858096
R22525 IPD.n265 IPD.n264 0.00858096
R22526 IPD.n278 IPD.n277 0.00858096
R22527 IPD.n274 IPD.n273 0.00858096
R22528 IPD.n272 IPD.n265 0.00858096
R22529 IPD.n234 IPD.n233 0.00858096
R22530 IPD.n243 IPD.n242 0.00858096
R22531 IPD.n244 IPD.n243 0.00858096
R22532 IPD.n235 IPD.n234 0.00858096
R22533 IPD.n226 IPD.n225 0.00858096
R22534 IPD.n180 IPD.n179 0.00858096
R22535 IPD.n172 IPD.n171 0.00858096
R22536 IPD.n181 IPD.n180 0.00858096
R22537 IPD.n179 IPD.n172 0.00858096
R22538 IPD.n153 IPD.n152 0.00858096
R22539 IPD.n154 IPD.n153 0.00858096
R22540 IPD.n44 IPD.n43 0.00858096
R22541 IPD.n45 IPD.n44 0.00858096
R22542 IPD.n425 IPD.n424 0.00855417
R22543 IPD.n79 IPD.n78 0.00855417
R22544 IPD.n66 IPD.n65 0.00855417
R22545 IPD.n391 IPD.n390 0.00855417
R22546 IPD.n393 IPD.n392 0.00855417
R22547 IPD.n98 IPD.n97 0.00855417
R22548 IPD.n366 IPD.n365 0.00855417
R22549 IPD.n368 IPD.n367 0.00855417
R22550 IPD.n326 IPD.n325 0.00855417
R22551 IPD.n328 IPD.n327 0.00855417
R22552 IPD.n276 IPD.n275 0.00855417
R22553 IPD.n263 IPD.n262 0.00855417
R22554 IPD.n228 IPD.n227 0.00855417
R22555 IPD.n230 IPD.n229 0.00855417
R22556 IPD.n237 IPD.n236 0.00855417
R22557 IPD.n239 IPD.n238 0.00855417
R22558 IPD.n246 IPD.n245 0.00855417
R22559 IPD.n248 IPD.n247 0.00855417
R22560 IPD.n170 IPD.n169 0.00855417
R22561 IPD.n156 IPD.n155 0.00855417
R22562 IPD.n158 IPD.n157 0.00855417
R22563 IPD.n21 IPD.n20 0.00855417
R22564 IPD.n17 IPD.n16 0.00855417
R22565 IPD.n47 IPD.n46 0.00855417
R22566 IPD.n23 IPD.n22 0.00773989
R22567 IPD.n24 IPD.n23 0.00773989
R22568 IPD.n24 IPD.n1 0.00773989
R22569 IPD.n27 IPD.n26 0.00773989
R22570 IPD.n288 IPD.n287 0.00642105
R22571 IPD.n301 IPD.n300 0.00642105
R22572 IPD.n434 IPD.n433 0.00605114
R22573 IPD.n409 IPD.n408 0.00605114
R22574 IPD.n296 IPD.n295 0.00605114
R22575 IPD.n138 IPD.n137 0.00605114
R22576 IPD.n414 IPD.n413 0.00570918
R22577 IPD.n300 IPD.n299 0.00551512
R22578 IPD.n53 IPD.n25 0.00549102
R22579 IPD.n49 IPD.n27 0.00549102
R22580 IPD.n402 IPD.n401 0.00523684
R22581 IPD.n415 IPD.n414 0.00523684
R22582 IPD.n428 IPD.n427 0.00523684
R22583 IPD.n142 IPD.n141 0.0051267
R22584 IPD.n422 IPD.n412 0.00479588
R22585 IPD.n15 IPD.n14 0.00364318
R22586 VB2.n87 VB2.t50 62.1809
R22587 VB2.n88 VB2.t46 62.1809
R22588 VB2.n89 VB2.t60 62.1809
R22589 VB2.n90 VB2.t39 62.1809
R22590 VB2.n91 VB2.t55 62.1809
R22591 VB2.n92 VB2.t36 62.1809
R22592 VB2.n93 VB2.t54 62.1809
R22593 VB2.n78 VB2.t61 61.6594
R22594 VB2.n79 VB2.t67 61.6594
R22595 VB2.n80 VB2.t51 61.6594
R22596 VB2.n81 VB2.t63 61.6594
R22597 VB2.n82 VB2.t42 61.6594
R22598 VB2.n83 VB2.t56 61.6594
R22599 VB2.n85 VB2.t45 61.6594
R22600 VB2.n84 VB2.t34 61.6594
R22601 VB2.n72 VB2.t47 59.8344
R22602 VB2.n76 VB2.t44 59.8344
R22603 VB2.n77 VB2.t43 59.8344
R22604 VB2.n74 VB2.t57 59.8344
R22605 VB2.n75 VB2.t35 59.8344
R22606 VB2.n70 VB2.t49 59.8344
R22607 VB2.n71 VB2.t33 59.8344
R22608 VB2.n73 VB2.t69 59.8344
R22609 VB2.t67 VB2.n77 59.5737
R22610 VB2.t63 VB2.n75 59.5737
R22611 VB2.t45 VB2.n73 59.5737
R22612 VB2.t73 VB2.n85 57.7487
R22613 VB2.n87 VB2.t64 57.2273
R22614 VB2.n88 VB2.t40 57.2273
R22615 VB2.n89 VB2.t53 57.2273
R22616 VB2.n90 VB2.t71 57.2273
R22617 VB2.n91 VB2.t38 57.2273
R22618 VB2.n92 VB2.t70 57.2273
R22619 VB2.n93 VB2.t37 57.2273
R22620 VB2.n94 VB2.t65 57.2273
R22621 VB2.n86 VB2.t73 56.8812
R22622 VB2.n28 VB2.t10 31.4166
R22623 VB2.n38 VB2.t66 26.7169
R22624 VB2.n39 VB2.n38 20.8576
R22625 VB2.n40 VB2.n39 20.8576
R22626 VB2.n41 VB2.n40 20.8576
R22627 VB2.n42 VB2.n41 20.8576
R22628 VB2.n43 VB2.n42 20.8576
R22629 VB2.n45 VB2.n44 20.8576
R22630 VB2.n31 VB2.n30 19.8148
R22631 VB2.n21 VB2.n20 19.8148
R22632 VB2.n46 VB2.n43 19.8148
R22633 VB2.n46 VB2.n45 19.8148
R22634 VB2.n21 VB2.n19 19.8148
R22635 VB2.n77 VB2.n76 17.5205
R22636 VB2.n75 VB2.n74 17.5205
R22637 VB2.n71 VB2.n70 17.5205
R22638 VB2.n73 VB2.n72 17.5205
R22639 VB2.n79 VB2.n78 17.5205
R22640 VB2.n81 VB2.n80 17.5205
R22641 VB2.n83 VB2.n82 17.5205
R22642 VB2.n85 VB2.n84 17.5205
R22643 VB2.n88 VB2.n87 17.5205
R22644 VB2.n90 VB2.n89 17.5205
R22645 VB2.n92 VB2.n91 17.5205
R22646 VB2.n94 VB2.n93 17.5205
R22647 VB2.n20 VB2.t14 11.6023
R22648 VB2.n30 VB2.t26 11.6023
R22649 VB2.n38 VB2.t16 11.6023
R22650 VB2.n39 VB2.t8 11.6023
R22651 VB2.n40 VB2.t20 11.6023
R22652 VB2.n41 VB2.t0 11.6023
R22653 VB2.n42 VB2.t24 11.6023
R22654 VB2.n43 VB2.t2 11.6023
R22655 VB2.n45 VB2.t6 11.6023
R22656 VB2.n44 VB2.t18 11.6023
R22657 VB2.n19 VB2.t12 11.6023
R22658 VB2.n46 VB2.t28 10.5594
R22659 VB2.n28 VB2.t30 10.5594
R22660 VB2.n31 VB2.t4 10.5594
R22661 VB2.n21 VB2.t22 10.5594
R22662 VB2.n72 VB2.n71 9.73383
R22663 VB2.n80 VB2.n79 9.73383
R22664 VB2.n82 VB2.n81 9.73383
R22665 VB2.n84 VB2.n83 9.73383
R22666 VB2.n89 VB2.n88 9.73383
R22667 VB2.n91 VB2.n90 9.73383
R22668 VB2.n93 VB2.n92 9.73383
R22669 VB2.n110 VB2.n109 4.829
R22670 VB2.n64 VB2.n63 4.46943
R22671 VB2.n35 VB2.n21 4.0005
R22672 VB2.n32 VB2.n31 4.0005
R22673 VB2.n29 VB2.n28 4.0005
R22674 VB2.n47 VB2.n46 4.0005
R22675 VB2.n96 VB2.n95 3.91467
R22676 VB2.n12 VB2.t21 3.6405
R22677 VB2.n12 VB2.n11 3.6405
R22678 VB2.n14 VB2.t25 3.6405
R22679 VB2.n14 VB2.n13 3.6405
R22680 VB2.n16 VB2.t29 3.6405
R22681 VB2.n16 VB2.n15 3.6405
R22682 VB2.n18 VB2.t19 3.6405
R22683 VB2.n18 VB2.n17 3.6405
R22684 VB2.n23 VB2.t23 3.6405
R22685 VB2.n23 VB2.n22 3.6405
R22686 VB2.n25 VB2.t27 3.6405
R22687 VB2.n25 VB2.n24 3.6405
R22688 VB2.n27 VB2.t31 3.6405
R22689 VB2.n27 VB2.n26 3.6405
R22690 VB2.n51 VB2.t17 3.6405
R22691 VB2.n51 VB2.n50 3.6405
R22692 VB2.n29 VB2.n27 2.94093
R22693 VB2.n99 VB2.n86 2.8805
R22694 VB2.n52 VB2.n51 2.80007
R22695 VB2.n49 VB2.n12 2.78441
R22696 VB2.n48 VB2.n14 2.78441
R22697 VB2.n37 VB2.n16 2.78441
R22698 VB2.n36 VB2.n18 2.78441
R22699 VB2.n34 VB2.n23 2.78441
R22700 VB2.n33 VB2.n25 2.78441
R22701 VB2.n9 VB2.t32 2.53976
R22702 VB2.n53 VB2.n52 2.2505
R22703 VB2.n95 VB2.n94 1.643
R22704 VB2.n107 VB2.n106 1.50393
R22705 VB2.n67 VB2.n66 1.49812
R22706 VB2.n62 VB2.n61 1.49763
R22707 VB2.n58 VB2.n57 1.34881
R22708 VB2.n62 VB2.n9 1.18731
R22709 VB2.n114 VB2.n113 1.12675
R22710 VB2.n114 VB2.n68 1.126
R22711 VB2.n106 VB2.n99 0.901294
R22712 VB2.n56 VB2.n54 0.727916
R22713 VB2.n49 VB2.n48 0.626587
R22714 VB2.n37 VB2.n36 0.626587
R22715 VB2.n34 VB2.n33 0.626587
R22716 VB2.n52 VB2.n49 0.552239
R22717 VB2.n48 VB2.n47 0.470065
R22718 VB2.n36 VB2.n35 0.470065
R22719 VB2.n32 VB2.n29 0.313543
R22720 VB2.n47 VB2.n37 0.157022
R22721 VB2.n35 VB2.n34 0.157022
R22722 VB2.n33 VB2.n32 0.157022
R22723 VB2 VB2.n114 0.110576
R22724 VB2.n62 VB2.n8 0.0831446
R22725 VB2.n54 VB2.n53 0.0826464
R22726 VB2.n98 VB2.n97 0.0656316
R22727 VB2.n54 VB2.n10 0.0423164
R22728 VB2.n8 VB2.n7 0.0420655
R22729 VB2.n103 VB2.n102 0.0339644
R22730 VB2.n104 VB2.n103 0.0327802
R22731 VB2.n63 VB2.n62 0.0324737
R22732 VB2.n99 VB2.n98 0.0301053
R22733 VB2.n105 VB2.n104 0.0301053
R22734 VB2.n97 VB2.n96 0.0289211
R22735 VB2.n102 VB2.n101 0.0289211
R22736 VB2.n6 VB2.n5 0.0207053
R22737 VB2.n1 VB2.n0 0.0207053
R22738 VB2.n57 VB2.n56 0.0156875
R22739 VB2.n4 VB2.n3 0.014
R22740 VB2.n5 VB2.n4 0.0134654
R22741 VB2.n61 VB2.n58 0.0111023
R22742 VB2.n109 VB2.n108 0.00858096
R22743 VB2.n107 VB2.n69 0.00858096
R22744 VB2.n108 VB2.n107 0.00858096
R22745 VB2.n113 VB2.n111 0.00773989
R22746 VB2.n65 VB2.n64 0.00773989
R22747 VB2.n111 VB2.n110 0.00773989
R22748 VB2.n66 VB2.n65 0.00773989
R22749 VB2.n3 VB2.n2 0.00773989
R22750 VB2.n113 VB2.n112 0.00773989
R22751 VB2.n66 VB2.n6 0.00773989
R22752 VB2.n68 VB2.n1 0.00773989
R22753 VB2.n101 VB2.n100 0.00685938
R22754 VB2.n56 VB2.n55 0.00638348
R22755 VB2.n60 VB2.n59 0.00605114
R22756 VB2.n61 VB2.n60 0.00605114
R22757 VB2.n68 VB2.n67 0.00582347
R22758 VB2.n106 VB2.n105 0.0030309
R22759 IBIAS1.t13 IBIAS1.t0 82.1255
R22760 IBIAS1.n3 IBIAS1.t3 49.4342
R22761 IBIAS1.n0 IBIAS1.t11 42.7576
R22762 IBIAS1.n4 IBIAS1.t7 42.7576
R22763 IBIAS1.t0 IBIAS1.n3 29.7219
R22764 IBIAS1.n0 IBIAS1.t4 28.6791
R22765 IBIAS1.n11 IBIAS1.t14 28.6791
R22766 IBIAS1.n10 IBIAS1.t12 28.6791
R22767 IBIAS1.n9 IBIAS1.t8 28.6791
R22768 IBIAS1.n8 IBIAS1.t2 28.6791
R22769 IBIAS1.n7 IBIAS1.t10 28.6791
R22770 IBIAS1.n6 IBIAS1.t6 28.6791
R22771 IBIAS1.n5 IBIAS1.t13 28.6791
R22772 IBIAS1.n4 IBIAS1.t9 28.6791
R22773 IBIAS1.n5 IBIAS1.n4 14.0791
R22774 IBIAS1.n6 IBIAS1.n5 14.0791
R22775 IBIAS1.n7 IBIAS1.n6 14.0791
R22776 IBIAS1.n8 IBIAS1.n7 14.0791
R22777 IBIAS1.n9 IBIAS1.n8 14.0791
R22778 IBIAS1.n10 IBIAS1.n9 14.0791
R22779 IBIAS1.n11 IBIAS1.n10 14.0791
R22780 IBIAS1.n3 IBIAS1.n2 8.09246
R22781 IBIAS1.n12 IBIAS1.n11 7.3005
R22782 IBIAS1.n13 IBIAS1.n12 2.8805
R22783 IBIAS1.n1 IBIAS1.n0 2.8805
R22784 IBIAS1 IBIAS1.n17 1.03603
R22785 IBIAS1.n16 IBIAS1.n14 0.5355
R22786 IBIAS1.n14 IBIAS1.n13 0.062564
R22787 IBIAS1.n14 IBIAS1.n1 0.0620381
R22788 IBIAS1.n16 IBIAS1.n15 0.0145625
R22789 IBIAS1.n17 IBIAS1.n16 0.014
R22790 IB5.n18 IB5.t8 37.9344
R22791 IB5.n16 IB5.t6 37.9344
R22792 IB5.n18 IB5.t10 17.0773
R22793 IB5.n16 IB5.t4 17.0773
R22794 IB5.n6 IB5.n5 4.4194
R22795 IB5.n17 IB5.n16 4.0005
R22796 IB5.n19 IB5.n18 4.0005
R22797 IB5.n17 IB5.n15 3.58876
R22798 IB5 IB5.n30 1.8225
R22799 IB5 IB5.n13 1.68241
R22800 IB5.n24 IB5.t11 1.6385
R22801 IB5.n24 IB5.n23 1.6385
R22802 IB5.n15 IB5.t7 1.6385
R22803 IB5.n15 IB5.n14 1.6385
R22804 IB5.n26 IB5.n25 1.17795
R22805 IB5.n9 IB5.n8 1.16629
R22806 IB5.n10 IB5.n9 1.12717
R22807 IB5.n22 IB5.n21 1.1255
R22808 IB5.n25 IB5.n24 1.06216
R22809 IB5.n8 IB5.n3 1.01901
R22810 IB5.n29 IB5.n27 0.616779
R22811 IB5.n3 IB5.t0 0.4555
R22812 IB5.n3 IB5.n2 0.4555
R22813 IB5.n5 IB5.t1 0.4555
R22814 IB5.n5 IB5.n4 0.4555
R22815 IB5.n19 IB5.n17 0.313543
R22816 IB5.n20 IB5.n19 0.281106
R22817 IB5.n9 IB5.n1 0.0832399
R22818 IB5.n8 IB5.n7 0.0824054
R22819 IB5.n27 IB5.n22 0.0712285
R22820 IB5.n27 IB5.n26 0.0534597
R22821 IB5.n1 IB5.n0 0.0419676
R22822 IB5.n21 IB5.n20 0.0407632
R22823 IB5.n7 IB5.n6 0.0324737
R22824 IB5.n30 IB5.n29 0.0156875
R22825 IB5.n12 IB5.n11 0.00860784
R22826 IB5.n29 IB5.n28 0.00860784
R22827 IB5.n13 IB5.n12 0.00855417
R22828 IB5.n11 IB5.n10 0.00364318
R22829 VND.n73 VND.t8 5.20893
R22830 VND.n76 VND.n74 5.20893
R22831 VND.n77 VND.t15 5.20893
R22832 VND.n64 VND.n63 5.11992
R22833 VND.n70 VND.n69 5.0524
R22834 VND.n17 VND.n16 5.0524
R22835 VND.n99 VND.n98 4.53845
R22836 VND.n114 VND.n113 4.53845
R22837 VND.n72 VND.t4 4.17588
R22838 VND.n70 VND.t12 3.92545
R22839 VND.n71 VND.n68 3.92545
R22840 VND.n17 VND.t9 3.92545
R22841 VND.n18 VND.n15 3.92545
R22842 VND.n73 VND.t5 3.18197
R22843 VND.n76 VND.n75 3.18197
R22844 VND.n77 VND.t7 3.18197
R22845 VND.n83 VND.n82 2.40175
R22846 VND.n150 VND.n149 1.65012
R22847 VND.n54 VND.n53 1.58409
R22848 VND.n38 VND.t22 1.58409
R22849 VND.n22 VND.t11 1.58402
R22850 VND.n156 VND.n5 1.50106
R22851 VND.n153 VND.n62 1.49801
R22852 VND.n29 VND.n28 1.4964
R22853 VND.n29 VND.n24 1.48461
R22854 VND.n122 VND.t23 1.40773
R22855 VND.n143 VND.n142 1.40773
R22856 VND.n78 VND.n77 1.37007
R22857 VND.n151 VND.n150 1.35681
R22858 VND.n19 VND.n18 1.26302
R22859 VND.n150 VND.n120 1.25459
R22860 VND.n123 VND.n122 1.19469
R22861 VND.n144 VND.n143 1.19469
R22862 VND.n134 VND.n133 1.19441
R22863 VND.n95 VND.n94 1.18273
R22864 VND.n110 VND.n109 1.18273
R22865 VND.n96 VND.n95 1.17276
R22866 VND.n111 VND.n110 1.17276
R22867 VND.n55 VND.n54 1.1643
R22868 VND.n13 VND.n12 1.1643
R22869 VND.n39 VND.n38 1.1643
R22870 VND.n23 VND.n22 1.1643
R22871 VND.n79 VND.n78 1.12746
R22872 VND.n67 VND.n66 1.1255
R22873 VND.n85 VND.n84 1.1255
R22874 VND.n101 VND.n100 1.1255
R22875 VND.n116 VND.n115 1.1255
R22876 VND.n157 VND.n156 1.1255
R22877 VND.n41 VND.n40 1.10737
R22878 VND.n57 VND.n56 1.10737
R22879 VND.n12 VND.n11 1.00262
R22880 VND.n45 VND.n14 0.88565
R22881 VND.n72 VND.n71 0.877022
R22882 VND.n91 VND.n90 0.87575
R22883 VND.n133 VND.n132 0.825944
R22884 VND.n79 VND.n73 0.743978
R22885 VND.n78 VND.n76 0.743978
R22886 VND.n103 VND.n102 0.727916
R22887 VND.n118 VND.n117 0.727916
R22888 VND.n137 VND.n136 0.727916
R22889 VND.n147 VND.n146 0.727916
R22890 VND.n71 VND.n70 0.626587
R22891 VND.n80 VND.n79 0.626587
R22892 VND.n18 VND.n17 0.626587
R22893 VND.n32 VND.n31 0.62375
R22894 VND.n88 VND.n86 0.616779
R22895 VND.n126 VND.n124 0.616779
R22896 VND.n82 VND.n81 0.58197
R22897 VND.n98 VND.t28 0.58197
R22898 VND.n98 VND.n97 0.58197
R22899 VND.n94 VND.t20 0.58197
R22900 VND.n94 VND.n93 0.58197
R22901 VND.n113 VND.t18 0.58197
R22902 VND.n113 VND.n112 0.58197
R22903 VND.n109 VND.t19 0.58197
R22904 VND.n109 VND.n108 0.58197
R22905 VND.n132 VND.t17 0.58197
R22906 VND.n132 VND.n131 0.58197
R22907 VND.n11 VND.t30 0.58197
R22908 VND.n11 VND.n10 0.58197
R22909 VND.n60 VND.n59 0.497625
R22910 VND.n80 VND.n72 0.3605
R22911 VND.n66 VND.n64 0.341925
R22912 VND.n100 VND.n99 0.341925
R22913 VND.n115 VND.n114 0.341925
R22914 VND.n106 VND.n105 0.330125
R22915 VND.n140 VND.n139 0.330125
R22916 VND.n129 VND.n128 0.330125
R22917 VND.n47 VND.n46 0.330125
R22918 VND.n44 VND.n43 0.330125
R22919 VND.n83 VND.n80 0.206051
R22920 VND VND.n157 0.09825
R22921 VND.n14 VND.n8 0.0936537
R22922 VND.n56 VND.n51 0.0880141
R22923 VND.n40 VND.n36 0.0880141
R22924 VND.n102 VND.n101 0.0826464
R22925 VND.n117 VND.n116 0.0826464
R22926 VND.n136 VND.n135 0.0826464
R22927 VND.n146 VND.n145 0.0826464
R22928 VND.n22 VND.n21 0.0786497
R22929 VND.n54 VND.n52 0.0786471
R22930 VND.n12 VND.n9 0.0786471
R22931 VND.n38 VND.n37 0.0786471
R22932 VND.n86 VND.n67 0.0712285
R22933 VND.n124 VND.n121 0.0712285
R22934 VND.n86 VND.n85 0.0534597
R22935 VND.n124 VND.n123 0.0534597
R22936 VND.n102 VND.n96 0.0423164
R22937 VND.n117 VND.n111 0.0423164
R22938 VND.n136 VND.n134 0.0423164
R22939 VND.n146 VND.n144 0.0423164
R22940 VND.n24 VND.n23 0.0420655
R22941 VND.n56 VND.n55 0.0319869
R22942 VND.n40 VND.n39 0.0319869
R22943 VND.n66 VND.n65 0.0293873
R22944 VND.n14 VND.n13 0.0261793
R22945 VND.n20 VND.n19 0.0253684
R22946 VND.n154 VND.n153 0.0229474
R22947 VND.n84 VND.n83 0.022679
R22948 VND.n2 VND.n1 0.0207053
R22949 VND.n88 VND.n87 0.0156875
R22950 VND.n126 VND.n125 0.0156875
R22951 VND.n46 VND.n45 0.0156875
R22952 VND.n45 VND.n44 0.0156875
R22953 VND.n156 VND.n0 0.014
R22954 VND.n156 VND.n155 0.014
R22955 VND.n152 VND.n151 0.014
R22956 VND.n4 VND.n3 0.014
R22957 VND.n3 VND.n2 0.0134654
R22958 VND.n155 VND.n154 0.0134654
R22959 VND.n50 VND.n49 0.0133659
R22960 VND.n35 VND.n34 0.0133659
R22961 VND.n48 VND.n47 0.0111023
R22962 VND.n33 VND.n32 0.0111023
R22963 VND.n28 VND.n27 0.00958206
R22964 VND.n89 VND.n88 0.00860784
R22965 VND.n127 VND.n126 0.00860784
R22966 VND.n58 VND.n57 0.00860784
R22967 VND.n42 VND.n41 0.00860784
R22968 VND.n119 VND.n118 0.00858096
R22969 VND.n107 VND.n106 0.00858096
R22970 VND.n104 VND.n103 0.00858096
R22971 VND.n92 VND.n91 0.00858096
R22972 VND.n120 VND.n119 0.00858096
R22973 VND.n118 VND.n107 0.00858096
R22974 VND.n105 VND.n104 0.00858096
R22975 VND.n103 VND.n92 0.00858096
R22976 VND.n148 VND.n147 0.00858096
R22977 VND.n141 VND.n140 0.00858096
R22978 VND.n138 VND.n137 0.00858096
R22979 VND.n130 VND.n129 0.00858096
R22980 VND.n149 VND.n148 0.00858096
R22981 VND.n147 VND.n141 0.00858096
R22982 VND.n139 VND.n138 0.00858096
R22983 VND.n137 VND.n130 0.00858096
R22984 VND.n31 VND.n30 0.00858096
R22985 VND.n30 VND.n29 0.00858096
R22986 VND.n29 VND.n25 0.00858096
R22987 VND.n90 VND.n89 0.00855417
R22988 VND.n128 VND.n127 0.00855417
R22989 VND.n59 VND.n58 0.00855417
R22990 VND.n43 VND.n42 0.00855417
R22991 VND.n61 VND.n60 0.00773989
R22992 VND.n62 VND.n61 0.00773989
R22993 VND.n51 VND.n50 0.00642105
R22994 VND.n8 VND.n7 0.00642105
R22995 VND.n36 VND.n35 0.00642105
R22996 VND.n21 VND.n20 0.00642105
R22997 VND.n27 VND.n26 0.00642105
R22998 VND.n41 VND.n33 0.00605114
R22999 VND.n57 VND.n48 0.00605114
R23000 VND.n7 VND.n6 0.00551512
R23001 VND.n153 VND.n152 0.00549102
R23002 VND.n5 VND.n4 0.00299297
R23003 IBIAS4.t1 IBIAS4.t3 95.9434
R23004 IBIAS4.t6 IBIAS4.t5 95.9434
R23005 IBIAS4.t7 IBIAS4.t6 95.9434
R23006 IBIAS4.t8 IBIAS4.t7 95.9434
R23007 IBIAS4.t10 IBIAS4.t9 95.9434
R23008 IBIAS4.t11 IBIAS4.t10 95.9434
R23009 IBIAS4.t12 IBIAS4.t11 95.9434
R23010 IBIAS4.n11 IBIAS4.t12 51.7088
R23011 IBIAS4.n4 IBIAS4.t1 48.1313
R23012 IBIAS4.n8 IBIAS4.t8 46.538
R23013 IBIAS4.n5 IBIAS4.n4 11.0519
R23014 IBIAS4.n3 IBIAS4.t4 4.7685
R23015 IBIAS4.n4 IBIAS4.n3 4.67159
R23016 IBIAS4.n3 IBIAS4.t2 3.3285
R23017 IBIAS4.n10 IBIAS4.n9 2.8805
R23018 IBIAS4.n6 IBIAS4.n5 2.8805
R23019 IBIAS4.n12 IBIAS4.n11 2.8805
R23020 IBIAS4.n65 IBIAS4.n64 2.06258
R23021 IBIAS4.n81 IBIAS4.n79 1.4991
R23022 IBIAS4.n81 IBIAS4.n73 1.4991
R23023 IBIAS4.n68 IBIAS4.n67 1.4991
R23024 IBIAS4.n48 IBIAS4.n47 1.1785
R23025 IBIAS4.n44 IBIAS4.n43 1.14437
R23026 IBIAS4.n42 IBIAS4.n41 1.1255
R23027 IBIAS4.n57 IBIAS4.n56 1.11801
R23028 IBIAS4.n58 IBIAS4.n38 1.11801
R23029 IBIAS4.n64 IBIAS4.n63 1.11801
R23030 IBIAS4.n61 IBIAS4.n60 1.11782
R23031 IBIAS4.n26 IBIAS4.n25 1.11782
R23032 IBIAS4.n82 IBIAS4.n81 1.11782
R23033 IBIAS4.n47 IBIAS4.n46 1.06459
R23034 IBIAS4.n52 IBIAS4.n49 0.885535
R23035 IBIAS4.n52 IBIAS4.n45 0.885413
R23036 IBIAS4.n14 IBIAS4.n13 0.884809
R23037 IBIAS4.n46 IBIAS4.t0 0.8195
R23038 IBIAS4.n56 IBIAS4.n54 0.55888
R23039 IBIAS4.n9 IBIAS4.n8 0.507444
R23040 IBIAS4.n60 IBIAS4.n58 0.416908
R23041 IBIAS4.n17 IBIAS4.n16 0.342754
R23042 IBIAS4.n13 IBIAS4.n10 0.10277
R23043 IBIAS4 IBIAS4.n83 0.101275
R23044 IBIAS4.n45 IBIAS4.n42 0.0999822
R23045 IBIAS4.n7 IBIAS4.n6 0.0857741
R23046 IBIAS4.n10 IBIAS4.n7 0.042637
R23047 IBIAS4.n49 IBIAS4.n48 0.0265722
R23048 IBIAS4.n13 IBIAS4.n12 0.0261711
R23049 IBIAS4.n45 IBIAS4.n44 0.0257704
R23050 IBIAS4.n57 IBIAS4.n40 0.0179841
R23051 IBIAS4.n60 IBIAS4.n59 0.0179841
R23052 IBIAS4.n63 IBIAS4.n62 0.0179841
R23053 IBIAS4.n38 IBIAS4.n37 0.0177304
R23054 IBIAS4.n58 IBIAS4.n57 0.0177304
R23055 IBIAS4.n36 IBIAS4.n35 0.0177304
R23056 IBIAS4.n40 IBIAS4.n39 0.0173591
R23057 IBIAS4.n56 IBIAS4.n55 0.0173591
R23058 IBIAS4.n64 IBIAS4.n61 0.0173591
R23059 IBIAS4.n61 IBIAS4.n36 0.0173591
R23060 IBIAS4.n83 IBIAS4.n82 0.0173591
R23061 IBIAS4.n26 IBIAS4.n0 0.0173591
R23062 IBIAS4.n82 IBIAS4.n27 0.0173591
R23063 IBIAS4.n27 IBIAS4.n26 0.0173591
R23064 IBIAS4.n81 IBIAS4.n80 0.00905634
R23065 IBIAS4.n33 IBIAS4.n32 0.00890861
R23066 IBIAS4.n23 IBIAS4.n22 0.00890861
R23067 IBIAS4.n30 IBIAS4.n29 0.00890861
R23068 IBIAS4.n78 IBIAS4.n77 0.00890861
R23069 IBIAS4.n22 IBIAS4.n21 0.00890861
R23070 IBIAS4.n31 IBIAS4.n30 0.00890861
R23071 IBIAS4.n75 IBIAS4.n74 0.00736358
R23072 IBIAS4.n21 IBIAS4.n20 0.00736358
R23073 IBIAS4.n16 IBIAS4.n15 0.00692989
R23074 IBIAS4.n73 IBIAS4.n72 0.006697
R23075 IBIAS4.n79 IBIAS4.n78 0.006697
R23076 IBIAS4.n68 IBIAS4.n31 0.006697
R23077 IBIAS4.n19 IBIAS4.n18 0.00527411
R23078 IBIAS4.n24 IBIAS4.n23 0.00527411
R23079 IBIAS4.n29 IBIAS4.n28 0.00527411
R23080 IBIAS4.n53 IBIAS4.n52 0.00527411
R23081 IBIAS4.n51 IBIAS4.n50 0.00527411
R23082 IBIAS4.n54 IBIAS4.n53 0.00527411
R23083 IBIAS4.n52 IBIAS4.n51 0.00527411
R23084 IBIAS4.n70 IBIAS4.n69 0.00527411
R23085 IBIAS4.n67 IBIAS4.n34 0.00527411
R23086 IBIAS4.n66 IBIAS4.n65 0.00527411
R23087 IBIAS4.n34 IBIAS4.n33 0.00527411
R23088 IBIAS4.n18 IBIAS4.n17 0.00527411
R23089 IBIAS4.n67 IBIAS4.n66 0.00527411
R23090 IBIAS4.n71 IBIAS4.n70 0.00527411
R23091 IBIAS4.n25 IBIAS4.n24 0.00527411
R23092 IBIAS4.n14 IBIAS4.n2 0.00479961
R23093 IBIAS4.n2 IBIAS4.n1 0.00479961
R23094 IBIAS4.n20 IBIAS4.n19 0.00418126
R23095 IBIAS4.n76 IBIAS4.n75 0.00418126
R23096 IBIAS4.n79 IBIAS4.n76 0.0038485
R23097 IBIAS4.n73 IBIAS4.n71 0.0038485
R23098 IBIAS4.n81 IBIAS4.n68 0.0038485
R23099 IBIAS4.n15 IBIAS4.n14 0.0029822
R23100 IB4.n40 IB4.t23 22.0465
R23101 IB4.n33 IB4.t6 14.9532
R23102 IB4.n41 IB4.n40 11.0965
R23103 IB4.n42 IB4.n41 11.0965
R23104 IB4.n43 IB4.n42 11.0965
R23105 IB4.n47 IB4.n46 11.0965
R23106 IB4.n35 IB4.n34 11.0965
R23107 IB4.n40 IB4.t21 10.9505
R23108 IB4.n41 IB4.t25 10.9505
R23109 IB4.n42 IB4.t22 10.9505
R23110 IB4.n43 IB4.t19 10.9505
R23111 IB4.n46 IB4.t0 10.9505
R23112 IB4.n47 IB4.t4 10.9505
R23113 IB4.n35 IB4.t8 10.9505
R23114 IB4.n34 IB4.t2 10.9505
R23115 IB4.n45 IB4.n43 8.67659
R23116 IB4.n45 IB4.n44 5.29669
R23117 IB4.n33 IB4.n32 4.47769
R23118 IB4.n16 IB4.n15 4.0405
R23119 IB4.n34 IB4.n33 4.00459
R23120 IB4.n46 IB4.n45 4.00315
R23121 IB4.n52 IB4.n39 3.85876
R23122 IB4.n37 IB4.n36 2.8805
R23123 IB4.n49 IB4.n48 2.8805
R23124 IB4.n52 IB4.n51 2.8805
R23125 IB4.n16 IB4.n13 2.6005
R23126 IB4.n17 IB4.n11 2.6005
R23127 IB4.n48 IB4.n47 1.7525
R23128 IB4.n36 IB4.n35 1.7525
R23129 IB4.n17 IB4.n16 1.4405
R23130 IB4.n6 IB4.n5 1.26725
R23131 IB4 IB4.n24 1.20885
R23132 IB4.n20 IB4.n19 1.1255
R23133 IB4.n8 IB4.n7 1.1255
R23134 IB4.n29 IB4.n27 1.11801
R23135 IB4.n58 IB4.n57 1.11782
R23136 IB4 IB4.n59 1.07796
R23137 IB4.n18 IB4.n17 0.906819
R23138 IB4.n22 IB4.n21 0.885413
R23139 IB4.n39 IB4.t5 0.8195
R23140 IB4.n39 IB4.n38 0.8195
R23141 IB4.n32 IB4.t3 0.8195
R23142 IB4.n32 IB4.n31 0.8195
R23143 IB4.n57 IB4.n56 0.760113
R23144 IB4.n55 IB4.n53 0.61639
R23145 IB4.n5 IB4.t17 0.607167
R23146 IB4.n5 IB4.n4 0.607167
R23147 IB4.n11 IB4.t16 0.607167
R23148 IB4.n11 IB4.n10 0.607167
R23149 IB4.n13 IB4.t15 0.607167
R23150 IB4.n13 IB4.n12 0.607167
R23151 IB4.n15 IB4.t14 0.607167
R23152 IB4.n15 IB4.n14 0.607167
R23153 IB4.n7 IB4.n6 0.109351
R23154 IB4.n21 IB4.n8 0.0999822
R23155 IB4.n52 IB4.n50 0.0996189
R23156 IB4.n19 IB4.n9 0.0953821
R23157 IB4.n3 IB4.n2 0.0939351
R23158 IB4.n53 IB4.n52 0.0710322
R23159 IB4.n53 IB4.n37 0.0535557
R23160 IB4.n29 IB4.n28 0.0334577
R23161 IB4.n8 IB4.n3 0.0319869
R23162 IB4.n50 IB4.n49 0.0269989
R23163 IB4.n21 IB4.n20 0.0257704
R23164 IB4.n19 IB4.n18 0.0185116
R23165 IB4.n27 IB4.n25 0.0179841
R23166 IB4.n57 IB4.n30 0.0179841
R23167 IB4.n27 IB4.n26 0.0177304
R23168 IB4.n58 IB4.n29 0.0173591
R23169 IB4.n59 IB4.n58 0.0173591
R23170 IB4.n55 IB4.n54 0.00842254
R23171 IB4.n56 IB4.n55 0.00810563
R23172 IB4.n24 IB4.n23 0.00735609
R23173 IB4.n22 IB4.n1 0.00527411
R23174 IB4.n1 IB4.n0 0.00527411
R23175 IB4.n23 IB4.n22 0.00418876
R23176 IN_P.t23 IN_P.t13 147.304
R23177 IN_P.t3 IN_P.t11 147.304
R23178 IN_P.t20 IN_P.t8 147.304
R23179 IN_P.t6 IN_P.t0 147.304
R23180 IN_P.n41 IN_P.t19 75.0919
R23181 IN_P.n14 IN_P.t16 74.8891
R23182 IN_P.n47 IN_P.t17 73.3458
R23183 IN_P.n20 IN_P.t14 73.143
R23184 IN_P.n44 IN_P.t3 72.3487
R23185 IN_P.n42 IN_P.t5 72.3487
R23186 IN_P.n40 IN_P.t6 72.3487
R23187 IN_P.n34 IN_P.t18 72.3487
R23188 IN_P.n30 IN_P.t10 72.3487
R23189 IN_P.n17 IN_P.t21 72.3487
R23190 IN_P.n15 IN_P.t2 72.3487
R23191 IN_P.n13 IN_P.t7 72.3487
R23192 IN_P.n44 IN_P.t23 51.4916
R23193 IN_P.n42 IN_P.t4 51.4916
R23194 IN_P.n40 IN_P.t20 51.4916
R23195 IN_P.n34 IN_P.t9 51.4916
R23196 IN_P.n30 IN_P.t15 51.4916
R23197 IN_P.n17 IN_P.t22 51.4916
R23198 IN_P.n15 IN_P.t1 51.4916
R23199 IN_P.n13 IN_P.t12 51.4916
R23200 IN_P.n18 IN_P.n17 20.1648
R23201 IN_P.n14 IN_P.n13 20.1648
R23202 IN_P.n45 IN_P.n44 19.9041
R23203 IN_P.n41 IN_P.n40 19.9041
R23204 IN_P.n43 IN_P.n42 15.6747
R23205 IN_P.n16 IN_P.n15 15.4719
R23206 IN_P.n31 IN_P.n30 15.1167
R23207 IN_P.n35 IN_P.n34 12.7876
R23208 IN_P.n56 IN_P.n38 2.48131
R23209 IN_P.n36 IN_P.n35 2.26226
R23210 IN_P.n33 IN_P.n31 2.24392
R23211 IN_P.n57 IN_P.n56 1.8554
R23212 IN_P.n22 IN_P.n21 1.50595
R23213 IN_P.n25 IN_P.n24 1.50128
R23214 IN_P.n37 IN_P.n36 1.49987
R23215 IN_P.n6 IN_P.n1 1.49812
R23216 IN_P.n6 IN_P.n5 1.49812
R23217 IN_P.n58 IN_P.n29 1.49801
R23218 IN_P.n9 IN_P.n8 1.49801
R23219 IN_P.n59 IN_P.n58 1.12675
R23220 IN_P.n59 IN_P.n6 1.126
R23221 IN_P.n53 IN_P.n52 1.1073
R23222 IN_P.n56 IN_P.n55 1.09079
R23223 IN_P.n21 IN_P.n20 0.901569
R23224 IN_P.n48 IN_P.n47 0.897484
R23225 IN_P.n43 IN_P.n41 0.626587
R23226 IN_P.n45 IN_P.n43 0.626587
R23227 IN_P.n16 IN_P.n14 0.626587
R23228 IN_P.n18 IN_P.n16 0.626587
R23229 IN_P.n27 IN_P.n26 0.51225
R23230 IN_P.n47 IN_P.n45 0.239196
R23231 IN_P.n20 IN_P.n18 0.239196
R23232 IN_P IN_P.n59 0.128013
R23233 IN_P.n52 IN_P.n50 0.0649899
R23234 IN_P.n24 IN_P.n23 0.0623855
R23235 IN_P.n52 IN_P.n51 0.032498
R23236 IN_P.n47 IN_P.n46 0.0289211
R23237 IN_P.n50 IN_P.n49 0.0289211
R23238 IN_P.n20 IN_P.n19 0.0289211
R23239 IN_P.n12 IN_P.n11 0.0289211
R23240 IN_P.n5 IN_P.n4 0.0236139
R23241 IN_P.n33 IN_P.n32 0.0157541
R23242 IN_P.n6 IN_P.n0 0.014
R23243 IN_P.n6 IN_P.n3 0.014
R23244 IN_P.n58 IN_P.n57 0.014
R23245 IN_P.n8 IN_P.n7 0.014
R23246 IN_P.n3 IN_P.n2 0.0134654
R23247 IN_P.n26 IN_P.n25 0.0117561
R23248 IN_P.n55 IN_P.n54 0.0111023
R23249 IN_P.n29 IN_P.n27 0.00998204
R23250 IN_P.n53 IN_P.n39 0.00860784
R23251 IN_P.n38 IN_P.n37 0.00859375
R23252 IN_P.n22 IN_P.n10 0.00858096
R23253 IN_P.n49 IN_P.n48 0.00685938
R23254 IN_P.n25 IN_P.n22 0.00639619
R23255 IN_P.n36 IN_P.n33 0.00621251
R23256 IN_P.n54 IN_P.n53 0.00605114
R23257 IN_P.n58 IN_P.n9 0.00549102
R23258 IN_P.n29 IN_P.n28 0.00549102
R23259 IN_P.n21 IN_P.n12 0.00400424
R23260 VB3.n88 VB3.t36 51.5034
R23261 VB3.n87 VB3.t25 50.3184
R23262 VB3.n86 VB3.t32 50.3184
R23263 VB3.n85 VB3.t38 50.3184
R23264 VB3.n84 VB3.t23 50.3184
R23265 VB3.n83 VB3.t37 50.3184
R23266 VB3.n82 VB3.t49 50.3184
R23267 VB3.n81 VB3.t31 50.3184
R23268 VB3.n74 VB3.t20 50.3184
R23269 VB3.n66 VB3.t41 50.3184
R23270 VB3.n65 VB3.t52 50.3184
R23271 VB3.n70 VB3.t51 50.3184
R23272 VB3.n69 VB3.t45 50.3184
R23273 VB3.n71 VB3.t35 50.3184
R23274 VB3.n68 VB3.t17 50.3184
R23275 VB3.n72 VB3.t34 50.3184
R23276 VB3.n67 VB3.t26 50.3184
R23277 VB3.n77 VB3.t29 50.3184
R23278 VB3.n76 VB3.t27 50.3184
R23279 VB3.n80 VB3.t28 50.3184
R23280 VB3.n75 VB3.t24 50.3184
R23281 VB3.n78 VB3.t21 50.3184
R23282 VB3.n73 VB3.t18 50.3184
R23283 VB3.n79 VB3.t22 50.3184
R23284 VB3.n88 VB3.t48 48.2728
R23285 VB3.t36 VB3.n66 46.4076
R23286 VB3.n87 VB3.t30 46.4076
R23287 VB3.t30 VB3.n70 46.4076
R23288 VB3.n86 VB3.t39 46.4076
R23289 VB3.t39 VB3.n71 46.4076
R23290 VB3.n85 VB3.t46 46.4076
R23291 VB3.t46 VB3.n72 46.4076
R23292 VB3.n84 VB3.t47 46.4076
R23293 VB3.t47 VB3.n77 46.4076
R23294 VB3.n83 VB3.t44 46.4076
R23295 VB3.t44 VB3.n80 46.4076
R23296 VB3.n82 VB3.t43 46.4076
R23297 VB3.t41 VB3.n65 46.4076
R23298 VB3.t51 VB3.n69 46.4076
R23299 VB3.t29 VB3.n76 46.4076
R23300 VB3.n81 VB3.t40 46.4076
R23301 VB3.n45 VB3.t10 20.6621
R23302 VB3.n18 VB3.t33 20.0755
R23303 VB3.n88 VB3.n87 18.9805
R23304 VB3.n68 VB3.n67 17.5205
R23305 VB3.n76 VB3.n75 17.5205
R23306 VB3.n74 VB3.n73 17.5205
R23307 VB3.n79 VB3.n78 17.5205
R23308 VB3.n86 VB3.n85 17.5205
R23309 VB3.n84 VB3.n83 17.5205
R23310 VB3.n82 VB3.n81 17.5205
R23311 VB3.n18 VB3.t12 15.6434
R23312 VB3.n21 VB3.t0 15.6434
R23313 VB3.n24 VB3.t6 15.6434
R23314 VB3.n27 VB3.t4 15.6434
R23315 VB3.n32 VB3.t8 15.6434
R23316 VB3.n48 VB3.t2 15.6434
R23317 VB3.n69 VB3.n68 9.73383
R23318 VB3.n75 VB3.n74 9.73383
R23319 VB3.n80 VB3.n79 9.73383
R23320 VB3.n87 VB3.n86 9.73383
R23321 VB3.n85 VB3.n84 9.73383
R23322 VB3.n83 VB3.n82 9.73383
R23323 VB3.n10 VB3.n9 6.30365
R23324 VB3.n44 VB3.n43 5.31813
R23325 VB3.n28 VB3.n27 5.21479
R23326 VB3.n25 VB3.n24 5.21479
R23327 VB3.n22 VB3.n21 5.21479
R23328 VB3.n19 VB3.n18 5.21479
R23329 VB3.n101 VB3.n100 4.81124
R23330 VB3.n50 VB3.n49 4.5005
R23331 VB3.n33 VB3.n32 4.04157
R23332 VB3.n29 VB3.n28 4.0005
R23333 VB3.n26 VB3.n25 4.0005
R23334 VB3.n23 VB3.n22 4.0005
R23335 VB3.n20 VB3.n19 4.0005
R23336 VB3.n47 VB3.n46 4.0005
R23337 VB3.n35 VB3.n34 4.0005
R23338 VB3.n49 VB3.n48 3.91121
R23339 VB3.n35 VB3.n13 3.43224
R23340 VB3.n20 VB3.n17 3.43224
R23341 VB3.n26 VB3.n15 3.43224
R23342 VB3.n90 VB3.n89 2.8805
R23343 VB3.n13 VB3.t3 1.6385
R23344 VB3.n13 VB3.n12 1.6385
R23345 VB3.n17 VB3.t1 1.6385
R23346 VB3.n17 VB3.n16 1.6385
R23347 VB3.n15 VB3.t5 1.6385
R23348 VB3.n15 VB3.n14 1.6385
R23349 VB3.n98 VB3.n97 1.50393
R23350 VB3.n5 VB3.n2 1.19078
R23351 VB3.n34 VB3.n33 1.17371
R23352 VB3.n6 VB3.n5 1.12754
R23353 VB3.n58 VB3.n53 1.1255
R23354 VB3.n38 VB3.n37 1.1255
R23355 VB3 VB3.n101 1.05692
R23356 VB3.n89 VB3.n88 0.973833
R23357 VB3.n97 VB3.n90 0.901294
R23358 VB3.n2 VB3.n1 0.813065
R23359 VB3.n101 VB3.n60 0.806689
R23360 VB3.n39 VB3.n38 0.563
R23361 VB3.n59 VB3.n58 0.563
R23362 VB3.n1 VB3.t15 0.4555
R23363 VB3.n1 VB3.n0 0.4555
R23364 VB3.n34 VB3.n31 0.326393
R23365 VB3.n29 VB3.n26 0.253132
R23366 VB3.n26 VB3.n23 0.253132
R23367 VB3.n23 VB3.n20 0.253132
R23368 VB3.n30 VB3.n29 0.218237
R23369 VB3.n46 VB3.n45 0.196036
R23370 VB3.n64 VB3.n63 0.0656316
R23371 VB3.n5 VB3.n4 0.0623855
R23372 VB3.n4 VB3.n3 0.0623855
R23373 VB3.n52 VB3.n51 0.042
R23374 VB3.n94 VB3.n93 0.0339644
R23375 VB3.n95 VB3.n94 0.0327802
R23376 VB3.n90 VB3.n64 0.0301053
R23377 VB3.n96 VB3.n95 0.0301053
R23378 VB3.n63 VB3.n62 0.0289211
R23379 VB3.n93 VB3.n92 0.0289211
R23380 VB3.n56 VB3.n55 0.0255
R23381 VB3.n41 VB3.n40 0.0255
R23382 VB3.n50 VB3.n47 0.0148158
R23383 VB3.n60 VB3.n59 0.014
R23384 VB3.n59 VB3.n41 0.014
R23385 VB3.n40 VB3.n39 0.014
R23386 VB3.n39 VB3.n10 0.014
R23387 VB3.n57 VB3.n56 0.012
R23388 VB3.n9 VB3.n8 0.0117561
R23389 VB3.n53 VB3.n50 0.0115
R23390 VB3.n58 VB3.n42 0.0115
R23391 VB3.n35 VB3.n30 0.0095
R23392 VB3.n100 VB3.n99 0.00858096
R23393 VB3.n99 VB3.n98 0.00858096
R23394 VB3.n98 VB3.n61 0.00858096
R23395 VB3.n92 VB3.n91 0.00685938
R23396 VB3.n8 VB3.n7 0.00639619
R23397 VB3.n55 VB3.n54 0.0055
R23398 VB3.n47 VB3.n44 0.00523684
R23399 VB3.n37 VB3.n36 0.005
R23400 VB3.n38 VB3.n11 0.005
R23401 VB3.n97 VB3.n96 0.0030309
R23402 VB3.n7 VB3.n6 0.00301938
R23403 VB3.n36 VB3.n35 0.003
R23404 VB3.n53 VB3.n52 0.0025
R23405 VB3.n58 VB3.n57 0.0025
R23406 IB3.n4 IB3.n3 4.05833
R23407 IB3.n9 IB3.n8 4.05833
R23408 IB3.n4 IB3.n1 3.43224
R23409 IB3.n9 IB3.n6 3.43224
R23410 IB3.n3 IB3.t6 1.6385
R23411 IB3.n3 IB3.n2 1.6385
R23412 IB3.n1 IB3.t0 1.6385
R23413 IB3.n1 IB3.n0 1.6385
R23414 IB3.n6 IB3.t2 1.6385
R23415 IB3.n6 IB3.n5 1.6385
R23416 IB3.n8 IB3.t5 1.6385
R23417 IB3.n8 IB3.n7 1.6385
R23418 IB3 IB3.n4 0.313543
R23419 IB3 IB3.n9 0.313543
R23420 VBIASN.n7 VBIASN.t7 15.7407
R23421 VBIASN.n25 VBIASN.n24 14.0791
R23422 VBIASN.n26 VBIASN.n25 14.0791
R23423 VBIASN.n27 VBIASN.n26 14.0791
R23424 VBIASN.n28 VBIASN.n27 14.0791
R23425 VBIASN.n29 VBIASN.n28 14.0791
R23426 VBIASN.n30 VBIASN.n29 14.0791
R23427 VBIASN.n23 VBIASN.t1 11.2226
R23428 VBIASN.n31 VBIASN.n30 8.47371
R23429 VBIASN.n37 VBIASN.t12 7.82193
R23430 VBIASN.n30 VBIASN.t8 7.82193
R23431 VBIASN.n29 VBIASN.t13 7.82193
R23432 VBIASN.n28 VBIASN.t10 7.82193
R23433 VBIASN.n27 VBIASN.t5 7.82193
R23434 VBIASN.n26 VBIASN.t6 7.82193
R23435 VBIASN.n25 VBIASN.t11 7.82193
R23436 VBIASN.n24 VBIASN.t3 7.82193
R23437 VBIASN.n43 VBIASN.n15 6.50674
R23438 VBIASN.n38 VBIASN.n37 4.05371
R23439 VBIASN.n23 VBIASN.n22 3.82142
R23440 VBIASN.n24 VBIASN.n23 3.3996
R23441 VBIASN.n32 VBIASN.n31 2.8805
R23442 VBIASN VBIASN.n52 2.30347
R23443 VBIASN.n22 VBIASN.t2 1.6385
R23444 VBIASN.n22 VBIASN.n21 1.6385
R23445 VBIASN.n14 VBIASN.n13 1.49823
R23446 VBIASN.n46 VBIASN.t0 1.4744
R23447 VBIASN.n13 VBIASN.n7 1.44232
R23448 VBIASN.n43 VBIASN.n42 1.25829
R23449 VBIASN.n52 VBIASN.n51 1.23398
R23450 VBIASN.n47 VBIASN.n46 1.1663
R23451 VBIASN.n48 VBIASN.n47 1.12717
R23452 VBIASN.n33 VBIASN.n32 0.902051
R23453 VBIASN.n39 VBIASN.n38 0.90016
R23454 VBIASN.n41 VBIASN.n40 0.7505
R23455 VBIASN.n34 VBIASN.n33 0.660817
R23456 VBIASN.n52 VBIASN.n43 0.287827
R23457 VBIASN.n47 VBIASN.n45 0.0832399
R23458 VBIASN.n45 VBIASN.n44 0.0419676
R23459 VBIASN.n32 VBIASN.n20 0.0293462
R23460 VBIASN.n38 VBIASN.n36 0.0281923
R23461 VBIASN.n18 VBIASN.n17 0.0255
R23462 VBIASN.n35 VBIASN.n34 0.0255
R23463 VBIASN.n11 VBIASN.n10 0.0212001
R23464 VBIASN.n4 VBIASN.n3 0.0212001
R23465 VBIASN.n3 VBIASN.n2 0.0147081
R23466 VBIASN.n12 VBIASN.n11 0.0147081
R23467 VBIASN.n33 VBIASN.n19 0.0144191
R23468 VBIASN.n41 VBIASN.n35 0.014
R23469 VBIASN.n42 VBIASN.n41 0.014
R23470 VBIASN.n13 VBIASN.n12 0.013
R23471 VBIASN.n9 VBIASN.n8 0.013
R23472 VBIASN.n2 VBIASN.n1 0.013
R23473 VBIASN.n15 VBIASN.n14 0.00931793
R23474 VBIASN.n50 VBIASN.n49 0.00860784
R23475 VBIASN.n51 VBIASN.n50 0.00855417
R23476 VBIASN.n10 VBIASN.n9 0.00699201
R23477 VBIASN.n5 VBIASN.n4 0.00699201
R23478 VBIASN.n1 VBIASN.n0 0.00532545
R23479 VBIASN.n14 VBIASN.n5 0.00515896
R23480 VBIASN.n13 VBIASN.n6 0.0049929
R23481 VBIASN.n49 VBIASN.n48 0.00364318
R23482 VBIASN.n40 VBIASN.n39 0.00348176
R23483 VBIASN.n17 VBIASN.n16 0.002
R23484 VBIASN.n19 VBIASN.n18 0.0015
R23485 a_29248_n5498.t1 a_29248_n5498.t2 6.46072
R23486 a_29248_n5498.t0 a_29248_n5498.t1 6.4095
R23487 IB2.n18 IB2.t11 7.0505
R23488 IB2.n17 IB2.t6 3.6405
R23489 IB2.n17 IB2.n16 3.6405
R23490 IB2.n15 IB2.t14 3.6405
R23491 IB2.n15 IB2.n14 3.6405
R23492 IB2.n13 IB2.t13 3.6405
R23493 IB2.n13 IB2.n12 3.6405
R23494 IB2.n11 IB2.t8 3.6405
R23495 IB2.n11 IB2.n10 3.6405
R23496 IB2.n9 IB2.t2 3.6405
R23497 IB2.n9 IB2.n8 3.6405
R23498 IB2.n1 IB2.t1 3.6405
R23499 IB2.n1 IB2.n0 3.6405
R23500 IB2.n3 IB2.t9 3.6405
R23501 IB2.n3 IB2.n2 3.6405
R23502 IB2.n5 IB2.t16 3.6405
R23503 IB2.n5 IB2.n4 3.6405
R23504 IB2.n6 IB2.n5 3.4105
R23505 IB2.n18 IB2.n17 2.78441
R23506 IB2.n19 IB2.n15 2.78441
R23507 IB2.n20 IB2.n13 2.78441
R23508 IB2.n21 IB2.n11 2.78441
R23509 IB2.n22 IB2.n9 2.78441
R23510 IB2.n7 IB2.n1 2.78441
R23511 IB2.n6 IB2.n3 2.78441
R23512 IB2.n7 IB2.n6 0.626587
R23513 IB2.n22 IB2.n21 0.626587
R23514 IB2.n21 IB2.n20 0.626587
R23515 IB2.n20 IB2.n19 0.626587
R23516 IB2.n19 IB2.n18 0.626587
R23517 IB2 IB2.n7 0.503326
R23518 IB2 IB2.n22 0.123761
C0 OUT2 IBIAS3 0.00232f
C1 VB2 IBS 1.95f
C2 VB1 VOUT 6.79f
C3 VB3 IBIAS1 0.0776f
C4 a_24070_n5442# VOUT 0.00744f
C5 a_25806_n7414# VDD 1.11f
C6 VDD VB4 0.72f
C7 IN_N IBIAS 0.00717f
C8 IN_P IPD 0.59f
C9 IND BD 9.48f
C10 a_24798_n7414# OUT_P 0.00312f
C11 VOUT IB4 0.376f
C12 IBIAS1 IB2 0.0416f
C13 a_24350_n7414# a_25078_n6312# 0.00757f
C14 VDD IBIAS1 4.43f
C15 OUT1 VND 6.12f
C16 OUT2 VB3 1.58f
C17 IBIAS VB1 1.84f
C18 a_25078_n5442# a_26254_n4340# 0.00743f
C19 a_25526_n5442# a_25806_n4340# 0.00743f
C20 a_23622_n5442# VOUT 0.0181f
C21 a_24350_n7414# a_24798_n7414# 0.281f
C22 a_24798_n4340# OUT1 0.0033f
C23 a_26254_n7414# IBIAS2 5.5e-19
C24 a_24350_n7414# OUT_P 0.0246f
C25 VB2 VBIASN 1.23f
C26 VB1 VCD 7.56f
C27 VCM VOUT 2.44f
C28 VB3 IB5 0.562f
C29 a_25526_n6312# VDD 0.299f
C30 BD IPD 9.31f
C31 VDD OUT2 12.2f
C32 IND IBIAS 0.00217f
C33 a_25078_n5442# a_25806_n4340# 0.00757f
C34 VBIASN IBIAS4 0.155f
C35 IB5 IB2 0.00262f
C36 a_24350_n4340# OUT1 0.0251f
C37 a_25806_n7414# IBIAS2 5.3e-19
C38 a_25078_n5442# a_25526_n5442# 0.281f
C39 VDD IB5 1.28f
C40 OUT1 VB1 0.656f
C41 OUT2 VPD 5.35f
C42 OUT_N VND 0.0017f
C43 IBIAS VCM 0.572f
C44 a_25078_n6312# VDD 0.747f
C45 a_23622_n6312# a_25078_n6312# 0.199f
C46 a_24798_n7414# VDD 0.302f
C47 OUT1 IB4 0.0172f
C48 VB2 IBIAS4 0.0154f
C49 VCM VCD 0.982f
C50 VB1 IBS 0.292f
C51 VOUT VBM 0.542f
C52 a_23622_n5442# a_26534_n5442# 2.06e-20
C53 a_23622_n6312# a_24798_n7414# 0.00743f
C54 a_24070_n6312# a_24350_n7414# 0.00743f
C55 IPD IBIAS 0.0029f
C56 VDD OUT_P 87f
C57 IND OUT1 4.85f
C58 a_25526_n6312# IBIAS2 0.00495f
C59 a_23622_n6312# OUT_P 0.00905f
C60 a_24350_n7414# VDD 1.05f
C61 VB2 VND 0.998f
C62 OUT2 IBIAS2 5.16e-19
C63 VB4 VOUT 0.0409f
C64 OUT1 VCM 0.00957f
C65 VDD IBIAS3 9.66f
C66 IBIAS VBM 0.235f
C67 a_24350_n4340# a_25806_n4340# 0.199f
C68 a_26534_n6312# a_26254_n7414# 0.00743f
C69 a_23622_n6312# a_24350_n7414# 0.00757f
C70 VB2 IVS 0.0083f
C71 VB1 VBIASN 0.128f
C72 VBM VCD 7.59f
C73 VCM IBS 0.108f
C74 a_25078_n6312# IBIAS2 0.0642f
C75 a_24798_n4340# a_25078_n5442# 0.00743f
C76 a_24350_n4340# a_25526_n5442# 0.00743f
C77 IPD OUT1 0.874f
C78 IBIAS VB4 0.185f
C79 VDD VB3 0.946f
C80 a_24798_n7414# IBIAS2 5.5e-19
C81 IBIAS4 IVS 0.393f
C82 VBIASN IB4 0.0856f
C83 a_26534_n6312# a_25806_n7414# 0.00659f
C84 a_24070_n6312# VDD 0.299f
C85 VB2 VB1 0.191f
C86 VB4 VCD 0.772f
C87 IBIAS IBIAS1 0.196f
C88 VDD IB2 0.845f
C89 OUT_P IBIAS2 16.4f
C90 OUT2 VOUT 0.0466f
C91 a_24350_n4340# a_25078_n5442# 0.00757f
C92 a_23622_n6312# a_24070_n6312# 0.281f
C93 a_24350_n7414# IBIAS2 5.3e-19
C94 VBM IBS 0.409f
C95 VB2 IB4 0.00218f
C96 VB3 IB3 1.09f
C97 IBIAS2 IBIAS3 1.68f
C98 a_26534_n5442# a_25806_n7414# 0.0101f
C99 a_23622_n6312# VDD 0.836f
C100 VB4 OUT1 0.00709f
C101 IND VB2 2.07e-20
C102 VDD VPD 10.7f
C103 IBIAS4 IB4 0.949f
C104 a_26254_n7414# OUT_N 5.58e-19
C105 a_24350_n4340# a_24798_n4340# 0.281f
C106 a_23622_n5442# a_25078_n5442# 0.199f
C107 IBIAS IB5 0.178f
C108 VB2 VCM 5.28e-19
C109 VND VB1 0.78f
C110 VB4 IBS 0.029f
C111 VDD IN_P 6.67f
C112 a_24070_n6312# IBIAS2 0.00495f
C113 a_26534_n6312# a_25078_n6312# 0.199f
C114 a_26534_n5442# a_25526_n6312# 0.0015f
C115 VBM VBIASN 0.174f
C116 VCD IB5 0.124f
C117 IBIAS1 IBS 0.361f
C118 VOUT IBIAS3 0.063f
C119 a_25806_n7414# OUT_N 7.77e-19
C120 OUT1 OUT2 30.7f
C121 VDD IBIAS2 0.142p
C122 IPD VB2 8.26e-20
C123 IVS IB4 1.15f
C124 a_23622_n6312# IBIAS2 0.0642f
C125 a_23622_n5442# a_24798_n4340# 0.00743f
C126 a_24070_n5442# a_24350_n4340# 0.00743f
C127 a_26534_n5442# a_25078_n6312# 0.00886f
C128 VB2 VBM 0.00633f
C129 VB4 VBIASN 0.108f
C130 VB3 VOUT 0.594f
C131 VDD BD 8.89f
C132 IN_N IND 0.716f
C133 a_26254_n4340# OUT2 6.86e-19
C134 IBS IB5 0.854f
C135 VB1 IB4 0.0425f
C136 IBIAS1 VBIASN 0.559f
C137 a_23622_n5442# a_24350_n4340# 0.00757f
C138 IBIAS VB3 0.656f
C139 OUT1 OUT_P 5.73f
C140 VDD VOUT 2.29f
C141 OUT2 OUT_N 5.36f
C142 VB4 VB2 0.0126f
C143 a_23622_n5442# a_24070_n5442# 0.281f
C144 a_25806_n4340# OUT2 6.86e-19
C145 OUT1 IBIAS3 0.00364f
C146 VB1 VCM 1.05f
C147 VB2 IBIAS1 0.0175f
C148 VB3 VCD 0.713f
C149 IBIAS IB2 0.0141f
C150 a_25526_n5442# a_25526_n6312# 0.00586f
C151 IN_N IPD 0.486f
C152 VDD IBIAS 9.74f
C153 IN_P BD 4.78f
C154 a_24798_n7414# OUT_N 0.00274f
C155 IB5 VBIASN 1.08f
C156 VOUT IB3 1.55e-19
C157 a_26534_n6312# VDD 0.859f
C158 OUT_N OUT_P 0.109p
C159 VDD VCD 0.0275f
C160 OUT2 VB2 1.03f
C161 OUT1 VB3 1.2f
C162 a_25078_n5442# a_25526_n6312# 0.00229f
C163 a_25526_n5442# a_25078_n6312# 0.00229f
C164 a_24350_n7414# OUT_N 0.153f
C165 VB3 IBS 1.14f
C166 VB2 IB5 0.004f
C167 VB1 VBM 2.6f
C168 IBIAS2 VOUT 0.00234f
C169 a_26534_n5442# VDD 0.951f
C170 VDD OUT1 8.72f
C171 IND IPD 14.3f
C172 IN_P IBIAS 0.216f
C173 a_25078_n5442# a_25078_n6312# 0.276f
C174 VCD IB3 5.9e-19
C175 VB4 VB1 0.193f
C176 IPD VCM 3.16e-20
C177 VDD IBS 2.11f
C178 OUT1 VPD 0.748f
C179 OUT2 VND 1.17f
C180 a_24798_n4340# OUT2 6.86e-19
C181 a_26534_n6312# IBIAS2 0.0606f
C182 a_24070_n6312# OUT_N 0.00833f
C183 VB3 VBIASN 0.285f
C184 VB1 IBIAS1 0.0893f
C185 VCM VBM 6.03f
C186 a_26254_n4340# VDD 0.303f
C187 VDD OUT_N 90.8f
C188 BD IBIAS 0.95f
C189 IND VB4 1.39f
C190 IBIAS3 IBIAS4 0.739f
C191 VBIASN IB2 0.0176f
C192 IBS IB3 0.00347f
C193 a_24350_n4340# OUT2 6.86e-19
C194 a_23622_n6312# OUT_N 5.3e-19
C195 a_26534_n5442# IBIAS2 0.205f
C196 a_25806_n4340# VDD 1.05f
C197 OUT_P VND 0.00173f
C198 VB4 VCM 0.412f
C199 IBIAS VOUT 0.352f
C200 VB2 VB3 0.619f
C201 OUT1 IBIAS2 0.431f
C202 VDD VBIASN 1.45f
C203 OUT2 VB1 0.3f
C204 a_25526_n5442# VDD 0.299f
C205 VB1 IB5 0.53f
C206 VOUT VCD 0.929f
C207 VB2 IB2 2.01f
C208 VDD VB2 12.7f
C209 IPD VB4 1.68f
C210 IND OUT2 0.655f
C211 a_26254_n4340# IBIAS2 0.00167f
C212 VBIASN IB3 3.45e-20
C213 IBIAS3 IVS 2.78f
C214 a_25806_n7414# a_26254_n7414# 0.281f
C215 a_25078_n5442# VDD 0.774f
C216 OUT2 VCM 0.00142f
C217 OUT1 VOUT 1.63f
C218 VB2 VPD 0.982f
C219 IBIAS VCD 0.515f
C220 VB4 VBM 0.561f
C221 OUT_N IBIAS2 14.4f
C222 VDD IBIAS4 3.94f
C223 VB3 VND 2.36e-19
C224 a_25806_n4340# IBIAS2 0.00769f
C225 VB2 IB3 0.0152f
C226 VBM IBIAS1 0.243f
C227 VOUT IBS 0.0174f
C228 VDD VND 9.42f
C229 IPD OUT2 5.04f
C230 a_25526_n5442# IBIAS2 0.00751f
C231 a_26534_n5442# a_26534_n6312# 0.372f
C232 IBIAS3 IB4 1.33f
C233 a_24798_n4340# VDD 0.302f
C234 VDD IVS 17.6f
C235 IBIAS IBS 0.597f
C236 VND VPD 10.7f
C237 VB3 VB1 0.553f
C238 VDD IN_N 7.53f
C239 a_25078_n5442# IBIAS2 0.142f
C240 a_24070_n5442# a_24070_n6312# 0.00586f
C241 IBIAS2 IBIAS4 0.0575f
C242 VBM IB5 0.101f
C243 a_25526_n6312# a_25806_n7414# 0.00743f
C244 a_25078_n6312# a_26254_n7414# 0.00743f
C245 VCD IBS 0.0309f
C246 VB1 IB2 0.0224f
C247 a_24350_n4340# VDD 1.01f
C248 a_26534_n5442# OUT1 0.00111f
C249 IND VB3 0.576f
C250 VDD VB1 9.95f
C251 VB4 OUT2 0.00296f
C252 a_24070_n5442# VDD 0.299f
C253 a_26254_n7414# OUT_P 0.00312f
C254 a_24070_n5442# a_23622_n6312# 0.00229f
C255 a_23622_n5442# a_24070_n6312# 0.00229f
C256 a_25078_n6312# a_25806_n7414# 0.00757f
C257 VB4 IB5 0.719f
C258 VB2 VOUT 0.149f
C259 VB3 VCM 0.267f
C260 VDD IB4 2.94f
C261 VPD VB1 0.946f
C262 IBIAS VBIASN 0.317f
C263 a_24798_n4340# IBIAS2 0.00167f
C264 a_26254_n4340# a_26534_n5442# 0.0146f
C265 a_25806_n4340# a_26534_n6312# 2.39e-19
C266 IN_N IN_P 2.38f
C267 VDD IND 7.04f
C268 a_23622_n5442# VDD 0.834f
C269 IBIAS1 IB5 0.186f
C270 IBIAS2 IVS 1.2f
C271 a_26254_n4340# OUT1 0.0033f
C272 VCD VBIASN 0.391f
C273 VOUT IBIAS4 0.0051f
C274 a_23622_n5442# a_23622_n6312# 0.276f
C275 a_25806_n7414# OUT_P 0.0232f
C276 OUT1 OUT_N 3.09f
C277 IBIAS VB2 0.0347f
C278 VDD VCM 0.101f
C279 IPD VB3 0.53f
C280 a_24350_n4340# IBIAS2 0.00769f
C281 a_25806_n4340# a_26534_n5442# 0.0341f
C282 a_24350_n7414# a_25806_n7414# 0.199f
C283 a_25078_n6312# a_25526_n6312# 0.281f
C284 a_25806_n4340# OUT1 0.0251f
C285 VB2 VCD 0.0792f
C286 VB3 VBM 0.0534f
C287 a_24070_n5442# IBIAS2 0.00751f
C288 a_25078_n5442# a_26534_n6312# 0.0223f
C289 a_25526_n5442# a_26534_n5442# 0.00199f
C290 a_24798_n4340# VOUT 8.94e-19
C291 IN_P IND 0.571f
C292 VDD IPD 2.94f
C293 IN_N BD 4.42f
C294 VBM IB2 0.0221f
C295 VCM IB3 6.71e-19
C296 VOUT IVS 0.0183f
C297 IBIAS2 IB4 0.725f
C298 IBS VBIASN 1.95f
C299 a_26254_n7414# VDD 0.303f
C300 VDD VBM 1.61f
C301 VB4 VB3 0.388f
C302 OUT2 OUT_P 4.06f
C303 OUT1 VB2 1.45f
C304 a_23622_n5442# IBIAS2 0.139f
C305 a_25806_n4340# a_26254_n4340# 0.281f
C306 a_25078_n5442# a_26534_n5442# 0.0543f
C307 a_24350_n4340# VOUT 0.0607f
C308 a_24350_n7414# a_25526_n6312# 0.00743f
C309 a_24798_n7414# a_25078_n6312# 0.00743f
.ends

