magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -1968 -1968 12576 14320
<< psubdiff >>
rect 32 12298 368 12320
rect 32 12252 54 12298
rect 100 12252 168 12298
rect 214 12252 368 12298
rect 32 12184 368 12252
rect 32 12138 54 12184
rect 100 12138 168 12184
rect 214 12138 368 12184
rect 32 12116 368 12138
rect 32 12070 236 12116
rect 32 12024 54 12070
rect 100 12024 168 12070
rect 214 12024 236 12070
rect 32 11500 236 12024
rect 32 11454 54 11500
rect 100 11454 168 11500
rect 214 11454 236 11500
rect 32 11386 236 11454
rect 32 11340 54 11386
rect 100 11340 168 11386
rect 214 11340 236 11386
rect 32 11272 236 11340
rect 32 11226 54 11272
rect 100 11226 168 11272
rect 214 11226 236 11272
rect 32 11158 236 11226
rect 32 11112 54 11158
rect 100 11112 168 11158
rect 214 11112 236 11158
rect 32 11044 236 11112
rect 32 10998 54 11044
rect 100 10998 168 11044
rect 214 10998 236 11044
rect 32 10930 236 10998
rect 32 10884 54 10930
rect 100 10884 168 10930
rect 214 10884 236 10930
rect 32 10816 236 10884
rect 32 10770 54 10816
rect 100 10770 168 10816
rect 214 10770 236 10816
rect 32 10702 236 10770
rect 32 10656 54 10702
rect 100 10656 168 10702
rect 214 10656 236 10702
rect 32 10588 236 10656
rect 32 10542 54 10588
rect 100 10542 168 10588
rect 214 10542 236 10588
rect 32 10474 236 10542
rect 32 10428 54 10474
rect 100 10428 168 10474
rect 214 10428 236 10474
rect 32 10360 236 10428
rect 32 10314 54 10360
rect 100 10314 168 10360
rect 214 10314 236 10360
rect 32 10246 236 10314
rect 32 10200 54 10246
rect 100 10200 168 10246
rect 214 10200 236 10246
rect 32 10132 236 10200
rect 32 10086 54 10132
rect 100 10086 168 10132
rect 214 10086 236 10132
rect 32 10018 236 10086
rect 32 9972 54 10018
rect 100 9972 168 10018
rect 214 9972 236 10018
rect 32 9904 236 9972
rect 32 9858 54 9904
rect 100 9858 168 9904
rect 214 9858 236 9904
rect 32 9790 236 9858
rect 32 9744 54 9790
rect 100 9744 168 9790
rect 214 9744 236 9790
rect 32 9676 236 9744
rect 32 9630 54 9676
rect 100 9630 168 9676
rect 214 9630 236 9676
rect 32 9562 236 9630
rect 32 9516 54 9562
rect 100 9516 168 9562
rect 214 9516 236 9562
rect 32 9448 236 9516
rect 32 9402 54 9448
rect 100 9402 168 9448
rect 214 9402 236 9448
rect 32 9334 236 9402
rect 32 9288 54 9334
rect 100 9288 168 9334
rect 214 9288 236 9334
rect 32 9220 236 9288
rect 32 9174 54 9220
rect 100 9174 168 9220
rect 214 9174 236 9220
rect 32 9106 236 9174
rect 32 9060 54 9106
rect 100 9060 168 9106
rect 214 9060 236 9106
rect 32 8992 236 9060
rect 32 8946 54 8992
rect 100 8946 168 8992
rect 214 8946 236 8992
rect 32 8878 236 8946
rect 32 8832 54 8878
rect 100 8832 168 8878
rect 214 8832 236 8878
rect 32 8764 236 8832
rect 32 8718 54 8764
rect 100 8718 168 8764
rect 214 8718 236 8764
rect 32 8650 236 8718
rect 32 8604 54 8650
rect 100 8604 168 8650
rect 214 8604 236 8650
rect 32 8536 236 8604
rect 32 8490 54 8536
rect 100 8490 168 8536
rect 214 8490 236 8536
rect 32 8422 236 8490
rect 32 8376 54 8422
rect 100 8376 168 8422
rect 214 8376 236 8422
rect 32 8308 236 8376
rect 32 8262 54 8308
rect 100 8262 168 8308
rect 214 8262 236 8308
rect 32 8194 236 8262
rect 32 8148 54 8194
rect 100 8148 168 8194
rect 214 8148 236 8194
rect 32 8080 236 8148
rect 32 8034 54 8080
rect 100 8034 168 8080
rect 214 8034 236 8080
rect 32 7966 236 8034
rect 32 7920 54 7966
rect 100 7920 168 7966
rect 214 7920 236 7966
rect 32 7852 236 7920
rect 32 7806 54 7852
rect 100 7806 168 7852
rect 214 7806 236 7852
rect 32 7738 236 7806
rect 32 7692 54 7738
rect 100 7692 168 7738
rect 214 7692 236 7738
rect 32 7624 236 7692
rect 32 7578 54 7624
rect 100 7578 168 7624
rect 214 7578 236 7624
rect 32 7510 236 7578
rect 32 7464 54 7510
rect 100 7464 168 7510
rect 214 7464 236 7510
rect 32 7396 236 7464
rect 32 7350 54 7396
rect 100 7350 168 7396
rect 214 7350 236 7396
rect 32 7282 236 7350
rect 32 7236 54 7282
rect 100 7236 168 7282
rect 214 7236 236 7282
rect 32 7168 236 7236
rect 32 7122 54 7168
rect 100 7122 168 7168
rect 214 7122 236 7168
rect 32 7054 236 7122
rect 32 7008 54 7054
rect 100 7008 168 7054
rect 214 7008 236 7054
rect 32 6940 236 7008
rect 32 6894 54 6940
rect 100 6894 168 6940
rect 214 6894 236 6940
rect 32 6826 236 6894
rect 32 6780 54 6826
rect 100 6780 168 6826
rect 214 6780 236 6826
rect 32 6712 236 6780
rect 32 6666 54 6712
rect 100 6666 168 6712
rect 214 6666 236 6712
rect 32 6598 236 6666
rect 32 6552 54 6598
rect 100 6552 168 6598
rect 214 6552 236 6598
rect 32 6484 236 6552
rect 32 6438 54 6484
rect 100 6438 168 6484
rect 214 6438 236 6484
rect 32 6370 236 6438
rect 32 6324 54 6370
rect 100 6324 168 6370
rect 214 6324 236 6370
rect 32 6256 236 6324
rect 32 6210 54 6256
rect 100 6210 168 6256
rect 214 6229 236 6256
rect 214 6210 300 6229
rect 32 6142 300 6210
rect 32 6096 54 6142
rect 100 6096 168 6142
rect 214 6096 300 6142
rect 32 6028 300 6096
rect 32 5982 54 6028
rect 100 5982 168 6028
rect 214 6025 300 6028
rect 214 5982 236 6025
rect 32 5914 236 5982
rect 32 5868 54 5914
rect 100 5868 168 5914
rect 214 5868 236 5914
rect 32 5800 236 5868
rect 32 5754 54 5800
rect 100 5754 168 5800
rect 214 5754 236 5800
rect 32 5686 236 5754
rect 32 5640 54 5686
rect 100 5640 168 5686
rect 214 5640 236 5686
rect 32 5572 236 5640
rect 32 5526 54 5572
rect 100 5526 168 5572
rect 214 5526 236 5572
rect 32 5458 236 5526
rect 32 5412 54 5458
rect 100 5412 168 5458
rect 214 5412 236 5458
rect 32 5344 236 5412
rect 32 5298 54 5344
rect 100 5298 168 5344
rect 214 5298 236 5344
rect 32 5230 236 5298
rect 32 5184 54 5230
rect 100 5184 168 5230
rect 214 5184 236 5230
rect 32 5116 236 5184
rect 32 5070 54 5116
rect 100 5070 168 5116
rect 214 5070 236 5116
rect 32 5002 236 5070
rect 32 4956 54 5002
rect 100 4956 168 5002
rect 214 4956 236 5002
rect 32 4888 236 4956
rect 32 4842 54 4888
rect 100 4842 168 4888
rect 214 4842 236 4888
rect 32 4774 236 4842
rect 32 4728 54 4774
rect 100 4728 168 4774
rect 214 4728 236 4774
rect 32 4660 236 4728
rect 32 4614 54 4660
rect 100 4614 168 4660
rect 214 4614 236 4660
rect 32 4546 236 4614
rect 32 4500 54 4546
rect 100 4500 168 4546
rect 214 4500 236 4546
rect 32 4432 236 4500
rect 32 4386 54 4432
rect 100 4386 168 4432
rect 214 4386 236 4432
rect 32 4318 236 4386
rect 32 4272 54 4318
rect 100 4272 168 4318
rect 214 4272 236 4318
rect 32 4204 236 4272
rect 32 4158 54 4204
rect 100 4158 168 4204
rect 214 4158 236 4204
rect 32 4090 236 4158
rect 32 4044 54 4090
rect 100 4044 168 4090
rect 214 4044 236 4090
rect 32 3976 236 4044
rect 32 3930 54 3976
rect 100 3930 168 3976
rect 214 3930 236 3976
rect 32 3862 236 3930
rect 32 3816 54 3862
rect 100 3816 168 3862
rect 214 3816 236 3862
rect 32 3748 236 3816
rect 32 3702 54 3748
rect 100 3702 168 3748
rect 214 3702 236 3748
rect 32 3634 236 3702
rect 32 3588 54 3634
rect 100 3588 168 3634
rect 214 3588 236 3634
rect 32 3520 236 3588
rect 32 3474 54 3520
rect 100 3474 168 3520
rect 214 3474 236 3520
rect 32 3406 236 3474
rect 32 3360 54 3406
rect 100 3360 168 3406
rect 214 3360 236 3406
rect 32 3292 236 3360
rect 32 3246 54 3292
rect 100 3246 168 3292
rect 214 3246 236 3292
rect 32 3178 236 3246
rect 32 3132 54 3178
rect 100 3132 168 3178
rect 214 3132 236 3178
rect 32 3064 236 3132
rect 32 3018 54 3064
rect 100 3018 168 3064
rect 214 3018 236 3064
rect 32 2950 236 3018
rect 32 2904 54 2950
rect 100 2904 168 2950
rect 214 2904 236 2950
rect 32 2836 236 2904
rect 32 2790 54 2836
rect 100 2790 168 2836
rect 214 2790 236 2836
rect 32 2722 236 2790
rect 32 2676 54 2722
rect 100 2676 168 2722
rect 214 2676 236 2722
rect 32 2608 236 2676
rect 32 2562 54 2608
rect 100 2562 168 2608
rect 214 2562 236 2608
rect 32 2494 236 2562
rect 32 2448 54 2494
rect 100 2448 168 2494
rect 214 2448 236 2494
rect 32 2380 236 2448
rect 32 2334 54 2380
rect 100 2334 168 2380
rect 214 2334 236 2380
rect 32 2266 236 2334
rect 32 2220 54 2266
rect 100 2220 168 2266
rect 214 2220 236 2266
rect 32 2152 236 2220
rect 32 2106 54 2152
rect 100 2106 168 2152
rect 214 2106 236 2152
rect 32 2038 236 2106
rect 32 1992 54 2038
rect 100 1992 168 2038
rect 214 1992 236 2038
rect 32 1924 236 1992
rect 32 1878 54 1924
rect 100 1878 168 1924
rect 214 1878 236 1924
rect 32 1810 236 1878
rect 32 1764 54 1810
rect 100 1764 168 1810
rect 214 1764 236 1810
rect 32 1696 236 1764
rect 32 1650 54 1696
rect 100 1650 168 1696
rect 214 1650 236 1696
rect 32 1582 236 1650
rect 32 1536 54 1582
rect 100 1536 168 1582
rect 214 1536 236 1582
rect 32 1468 236 1536
rect 32 1422 54 1468
rect 100 1422 168 1468
rect 214 1422 236 1468
rect 32 1354 236 1422
rect 32 1308 54 1354
rect 100 1308 168 1354
rect 214 1308 236 1354
rect 32 1240 236 1308
rect 32 1194 54 1240
rect 100 1194 168 1240
rect 214 1194 236 1240
rect 32 1126 236 1194
rect 32 1080 54 1126
rect 100 1080 168 1126
rect 214 1080 236 1126
rect 32 1012 236 1080
rect 32 966 54 1012
rect 100 966 168 1012
rect 214 966 236 1012
rect 32 898 236 966
rect 32 852 54 898
rect 100 852 168 898
rect 214 852 236 898
rect 32 784 236 852
rect 32 738 54 784
rect 100 738 168 784
rect 214 738 236 784
rect 32 328 236 738
rect 32 282 54 328
rect 100 282 168 328
rect 214 282 236 328
rect 32 236 236 282
rect 32 214 368 236
rect 32 168 54 214
rect 100 168 168 214
rect 214 168 368 214
rect 32 100 368 168
rect 32 54 54 100
rect 100 54 168 100
rect 214 54 368 100
rect 32 32 368 54
<< psubdiffcont >>
rect 54 12252 100 12298
rect 168 12252 214 12298
rect 54 12138 100 12184
rect 168 12138 214 12184
rect 54 12024 100 12070
rect 168 12024 214 12070
rect 54 11454 100 11500
rect 168 11454 214 11500
rect 54 11340 100 11386
rect 168 11340 214 11386
rect 54 11226 100 11272
rect 168 11226 214 11272
rect 54 11112 100 11158
rect 168 11112 214 11158
rect 54 10998 100 11044
rect 168 10998 214 11044
rect 54 10884 100 10930
rect 168 10884 214 10930
rect 54 10770 100 10816
rect 168 10770 214 10816
rect 54 10656 100 10702
rect 168 10656 214 10702
rect 54 10542 100 10588
rect 168 10542 214 10588
rect 54 10428 100 10474
rect 168 10428 214 10474
rect 54 10314 100 10360
rect 168 10314 214 10360
rect 54 10200 100 10246
rect 168 10200 214 10246
rect 54 10086 100 10132
rect 168 10086 214 10132
rect 54 9972 100 10018
rect 168 9972 214 10018
rect 54 9858 100 9904
rect 168 9858 214 9904
rect 54 9744 100 9790
rect 168 9744 214 9790
rect 54 9630 100 9676
rect 168 9630 214 9676
rect 54 9516 100 9562
rect 168 9516 214 9562
rect 54 9402 100 9448
rect 168 9402 214 9448
rect 54 9288 100 9334
rect 168 9288 214 9334
rect 54 9174 100 9220
rect 168 9174 214 9220
rect 54 9060 100 9106
rect 168 9060 214 9106
rect 54 8946 100 8992
rect 168 8946 214 8992
rect 54 8832 100 8878
rect 168 8832 214 8878
rect 54 8718 100 8764
rect 168 8718 214 8764
rect 54 8604 100 8650
rect 168 8604 214 8650
rect 54 8490 100 8536
rect 168 8490 214 8536
rect 54 8376 100 8422
rect 168 8376 214 8422
rect 54 8262 100 8308
rect 168 8262 214 8308
rect 54 8148 100 8194
rect 168 8148 214 8194
rect 54 8034 100 8080
rect 168 8034 214 8080
rect 54 7920 100 7966
rect 168 7920 214 7966
rect 54 7806 100 7852
rect 168 7806 214 7852
rect 54 7692 100 7738
rect 168 7692 214 7738
rect 54 7578 100 7624
rect 168 7578 214 7624
rect 54 7464 100 7510
rect 168 7464 214 7510
rect 54 7350 100 7396
rect 168 7350 214 7396
rect 54 7236 100 7282
rect 168 7236 214 7282
rect 54 7122 100 7168
rect 168 7122 214 7168
rect 54 7008 100 7054
rect 168 7008 214 7054
rect 54 6894 100 6940
rect 168 6894 214 6940
rect 54 6780 100 6826
rect 168 6780 214 6826
rect 54 6666 100 6712
rect 168 6666 214 6712
rect 54 6552 100 6598
rect 168 6552 214 6598
rect 54 6438 100 6484
rect 168 6438 214 6484
rect 54 6324 100 6370
rect 168 6324 214 6370
rect 54 6210 100 6256
rect 168 6210 214 6256
rect 54 6096 100 6142
rect 168 6096 214 6142
rect 54 5982 100 6028
rect 168 5982 214 6028
rect 54 5868 100 5914
rect 168 5868 214 5914
rect 54 5754 100 5800
rect 168 5754 214 5800
rect 54 5640 100 5686
rect 168 5640 214 5686
rect 54 5526 100 5572
rect 168 5526 214 5572
rect 54 5412 100 5458
rect 168 5412 214 5458
rect 54 5298 100 5344
rect 168 5298 214 5344
rect 54 5184 100 5230
rect 168 5184 214 5230
rect 54 5070 100 5116
rect 168 5070 214 5116
rect 54 4956 100 5002
rect 168 4956 214 5002
rect 54 4842 100 4888
rect 168 4842 214 4888
rect 54 4728 100 4774
rect 168 4728 214 4774
rect 54 4614 100 4660
rect 168 4614 214 4660
rect 54 4500 100 4546
rect 168 4500 214 4546
rect 54 4386 100 4432
rect 168 4386 214 4432
rect 54 4272 100 4318
rect 168 4272 214 4318
rect 54 4158 100 4204
rect 168 4158 214 4204
rect 54 4044 100 4090
rect 168 4044 214 4090
rect 54 3930 100 3976
rect 168 3930 214 3976
rect 54 3816 100 3862
rect 168 3816 214 3862
rect 54 3702 100 3748
rect 168 3702 214 3748
rect 54 3588 100 3634
rect 168 3588 214 3634
rect 54 3474 100 3520
rect 168 3474 214 3520
rect 54 3360 100 3406
rect 168 3360 214 3406
rect 54 3246 100 3292
rect 168 3246 214 3292
rect 54 3132 100 3178
rect 168 3132 214 3178
rect 54 3018 100 3064
rect 168 3018 214 3064
rect 54 2904 100 2950
rect 168 2904 214 2950
rect 54 2790 100 2836
rect 168 2790 214 2836
rect 54 2676 100 2722
rect 168 2676 214 2722
rect 54 2562 100 2608
rect 168 2562 214 2608
rect 54 2448 100 2494
rect 168 2448 214 2494
rect 54 2334 100 2380
rect 168 2334 214 2380
rect 54 2220 100 2266
rect 168 2220 214 2266
rect 54 2106 100 2152
rect 168 2106 214 2152
rect 54 1992 100 2038
rect 168 1992 214 2038
rect 54 1878 100 1924
rect 168 1878 214 1924
rect 54 1764 100 1810
rect 168 1764 214 1810
rect 54 1650 100 1696
rect 168 1650 214 1696
rect 54 1536 100 1582
rect 168 1536 214 1582
rect 54 1422 100 1468
rect 168 1422 214 1468
rect 54 1308 100 1354
rect 168 1308 214 1354
rect 54 1194 100 1240
rect 168 1194 214 1240
rect 54 1080 100 1126
rect 168 1080 214 1126
rect 54 966 100 1012
rect 168 966 214 1012
rect 54 852 100 898
rect 168 852 214 898
rect 54 738 100 784
rect 168 738 214 784
rect 54 282 100 328
rect 168 282 214 328
rect 54 168 100 214
rect 168 168 214 214
rect 54 54 100 100
rect 168 54 214 100
<< metal1 >>
rect 43 12298 10565 12310
rect 43 12252 54 12298
rect 100 12252 168 12298
rect 214 12252 10565 12298
rect 43 12184 10565 12252
rect 43 12138 54 12184
rect 100 12138 168 12184
rect 214 12138 10565 12184
rect 43 12126 10565 12138
rect 43 12070 225 12126
rect 43 12024 54 12070
rect 100 12024 168 12070
rect 214 12024 225 12070
rect 43 11633 225 12024
rect 689 11723 9913 11855
rect 689 11655 2605 11723
rect 3125 11655 5041 11723
rect 5561 11655 7477 11723
rect 7997 11655 9913 11723
rect 43 11500 429 11633
rect 43 11454 54 11500
rect 100 11454 168 11500
rect 214 11454 429 11500
rect 43 11386 429 11454
rect 43 11340 54 11386
rect 100 11340 168 11386
rect 214 11340 429 11386
rect 43 11272 429 11340
rect 43 11226 54 11272
rect 100 11226 168 11272
rect 214 11226 429 11272
rect 43 11158 429 11226
rect 43 11112 54 11158
rect 100 11112 168 11158
rect 214 11112 429 11158
rect 43 11044 429 11112
rect 43 10998 54 11044
rect 100 10998 168 11044
rect 214 10998 429 11044
rect 43 10930 429 10998
rect 43 10884 54 10930
rect 100 10884 168 10930
rect 214 10884 429 10930
rect 43 10816 429 10884
rect 43 10770 54 10816
rect 100 10770 168 10816
rect 214 10770 429 10816
rect 43 10702 429 10770
rect 43 10656 54 10702
rect 100 10656 168 10702
rect 214 10656 429 10702
rect 43 10588 429 10656
rect 43 10542 54 10588
rect 100 10542 168 10588
rect 214 10542 429 10588
rect 43 10474 429 10542
rect 43 10428 54 10474
rect 100 10428 168 10474
rect 214 10428 429 10474
rect 43 10360 429 10428
rect 43 10314 54 10360
rect 100 10314 168 10360
rect 214 10314 429 10360
rect 43 10246 429 10314
rect 43 10200 54 10246
rect 100 10200 168 10246
rect 214 10200 429 10246
rect 43 10132 429 10200
rect 43 10086 54 10132
rect 100 10086 168 10132
rect 214 10086 429 10132
rect 43 10018 429 10086
rect 43 9972 54 10018
rect 100 9972 168 10018
rect 214 9972 429 10018
rect 43 9904 429 9972
rect 43 9858 54 9904
rect 100 9858 168 9904
rect 214 9858 429 9904
rect 43 9790 429 9858
rect 43 9744 54 9790
rect 100 9744 168 9790
rect 214 9744 429 9790
rect 43 9676 429 9744
rect 43 9630 54 9676
rect 100 9630 168 9676
rect 214 9630 429 9676
rect 43 9562 429 9630
rect 43 9516 54 9562
rect 100 9516 168 9562
rect 214 9516 429 9562
rect 43 9448 429 9516
rect 43 9402 54 9448
rect 100 9402 168 9448
rect 214 9402 429 9448
rect 43 9334 429 9402
rect 43 9288 54 9334
rect 100 9288 168 9334
rect 214 9288 429 9334
rect 43 9220 429 9288
rect 43 9174 54 9220
rect 100 9174 168 9220
rect 214 9174 429 9220
rect 43 9106 429 9174
rect 43 9060 54 9106
rect 100 9060 168 9106
rect 214 9060 429 9106
rect 43 8992 429 9060
rect 43 8946 54 8992
rect 100 8946 168 8992
rect 214 8946 429 8992
rect 43 8878 429 8946
rect 43 8832 54 8878
rect 100 8832 168 8878
rect 214 8832 429 8878
rect 43 8764 429 8832
rect 43 8718 54 8764
rect 100 8718 168 8764
rect 214 8718 429 8764
rect 43 8650 429 8718
rect 43 8604 54 8650
rect 100 8604 168 8650
rect 214 8604 429 8650
rect 43 8536 429 8604
rect 43 8490 54 8536
rect 100 8490 168 8536
rect 214 8490 429 8536
rect 43 8422 429 8490
rect 43 8376 54 8422
rect 100 8376 168 8422
rect 214 8376 429 8422
rect 43 8308 429 8376
rect 43 8262 54 8308
rect 100 8262 168 8308
rect 214 8262 429 8308
rect 43 8194 429 8262
rect 43 8148 54 8194
rect 100 8148 168 8194
rect 214 8148 429 8194
rect 43 8080 429 8148
rect 43 8034 54 8080
rect 100 8034 168 8080
rect 214 8034 429 8080
rect 43 7966 429 8034
rect 43 7920 54 7966
rect 100 7920 168 7966
rect 214 7920 429 7966
rect 43 7852 429 7920
rect 43 7806 54 7852
rect 100 7806 168 7852
rect 214 7806 429 7852
rect 43 7738 429 7806
rect 43 7692 54 7738
rect 100 7692 168 7738
rect 214 7692 429 7738
rect 43 7624 429 7692
rect 43 7578 54 7624
rect 100 7578 168 7624
rect 214 7578 429 7624
rect 43 7510 429 7578
rect 43 7464 54 7510
rect 100 7464 168 7510
rect 214 7464 429 7510
rect 43 7396 429 7464
rect 43 7350 54 7396
rect 100 7350 168 7396
rect 214 7350 429 7396
rect 43 7282 429 7350
rect 43 7236 54 7282
rect 100 7236 168 7282
rect 214 7236 429 7282
rect 43 7168 429 7236
rect 43 7122 54 7168
rect 100 7122 168 7168
rect 214 7122 429 7168
rect 43 7054 429 7122
rect 43 7008 54 7054
rect 100 7008 168 7054
rect 214 7008 429 7054
rect 43 6940 429 7008
rect 43 6894 54 6940
rect 100 6894 168 6940
rect 214 6894 429 6940
rect 43 6826 429 6894
rect 43 6780 54 6826
rect 100 6780 168 6826
rect 214 6780 429 6826
rect 43 6712 429 6780
rect 43 6666 54 6712
rect 100 6666 168 6712
rect 214 6666 429 6712
rect 43 6598 429 6666
rect 43 6552 54 6598
rect 100 6552 168 6598
rect 214 6552 429 6598
rect 43 6484 429 6552
rect 43 6438 54 6484
rect 100 6438 168 6484
rect 214 6483 429 6484
rect 10173 6483 10383 11633
rect 214 6438 10383 6483
rect 43 6370 10383 6438
rect 43 6324 54 6370
rect 100 6324 168 6370
rect 214 6324 10383 6370
rect 43 6256 10383 6324
rect 43 6210 54 6256
rect 100 6210 168 6256
rect 214 6210 10383 6256
rect 43 6142 10383 6210
rect 43 6096 54 6142
rect 100 6096 168 6142
rect 214 6096 10383 6142
rect 43 6028 10383 6096
rect 43 5982 54 6028
rect 100 5982 168 6028
rect 214 5982 10383 6028
rect 43 5914 10383 5982
rect 43 5868 54 5914
rect 100 5868 168 5914
rect 214 5868 10383 5914
rect 43 5800 10383 5868
rect 43 5754 54 5800
rect 100 5754 168 5800
rect 214 5771 10383 5800
rect 214 5754 429 5771
rect 43 5686 429 5754
rect 43 5640 54 5686
rect 100 5640 168 5686
rect 214 5640 429 5686
rect 43 5572 429 5640
rect 43 5526 54 5572
rect 100 5526 168 5572
rect 214 5526 429 5572
rect 43 5458 429 5526
rect 43 5412 54 5458
rect 100 5412 168 5458
rect 214 5412 429 5458
rect 43 5344 429 5412
rect 43 5298 54 5344
rect 100 5298 168 5344
rect 214 5298 429 5344
rect 43 5230 429 5298
rect 43 5184 54 5230
rect 100 5184 168 5230
rect 214 5184 429 5230
rect 43 5116 429 5184
rect 43 5070 54 5116
rect 100 5070 168 5116
rect 214 5070 429 5116
rect 43 5002 429 5070
rect 43 4956 54 5002
rect 100 4956 168 5002
rect 214 4956 429 5002
rect 43 4888 429 4956
rect 43 4842 54 4888
rect 100 4842 168 4888
rect 214 4842 429 4888
rect 43 4774 429 4842
rect 43 4728 54 4774
rect 100 4728 168 4774
rect 214 4728 429 4774
rect 43 4660 429 4728
rect 43 4614 54 4660
rect 100 4614 168 4660
rect 214 4614 429 4660
rect 43 4546 429 4614
rect 43 4500 54 4546
rect 100 4500 168 4546
rect 214 4500 429 4546
rect 43 4432 429 4500
rect 43 4386 54 4432
rect 100 4386 168 4432
rect 214 4386 429 4432
rect 43 4318 429 4386
rect 43 4272 54 4318
rect 100 4272 168 4318
rect 214 4272 429 4318
rect 43 4204 429 4272
rect 43 4158 54 4204
rect 100 4158 168 4204
rect 214 4158 429 4204
rect 43 4090 429 4158
rect 43 4044 54 4090
rect 100 4044 168 4090
rect 214 4044 429 4090
rect 43 3976 429 4044
rect 43 3930 54 3976
rect 100 3930 168 3976
rect 214 3930 429 3976
rect 43 3862 429 3930
rect 43 3816 54 3862
rect 100 3816 168 3862
rect 214 3816 429 3862
rect 43 3748 429 3816
rect 43 3702 54 3748
rect 100 3702 168 3748
rect 214 3702 429 3748
rect 43 3634 429 3702
rect 43 3588 54 3634
rect 100 3588 168 3634
rect 214 3588 429 3634
rect 43 3520 429 3588
rect 43 3474 54 3520
rect 100 3474 168 3520
rect 214 3474 429 3520
rect 43 3406 429 3474
rect 43 3360 54 3406
rect 100 3360 168 3406
rect 214 3360 429 3406
rect 43 3292 429 3360
rect 43 3246 54 3292
rect 100 3246 168 3292
rect 214 3246 429 3292
rect 43 3178 429 3246
rect 43 3132 54 3178
rect 100 3132 168 3178
rect 214 3132 429 3178
rect 43 3064 429 3132
rect 43 3018 54 3064
rect 100 3018 168 3064
rect 214 3018 429 3064
rect 43 2950 429 3018
rect 43 2904 54 2950
rect 100 2904 168 2950
rect 214 2904 429 2950
rect 43 2836 429 2904
rect 43 2790 54 2836
rect 100 2790 168 2836
rect 214 2790 429 2836
rect 43 2722 429 2790
rect 43 2676 54 2722
rect 100 2676 168 2722
rect 214 2676 429 2722
rect 43 2608 429 2676
rect 43 2562 54 2608
rect 100 2562 168 2608
rect 214 2562 429 2608
rect 43 2494 429 2562
rect 43 2448 54 2494
rect 100 2448 168 2494
rect 214 2448 429 2494
rect 43 2380 429 2448
rect 43 2334 54 2380
rect 100 2334 168 2380
rect 214 2334 429 2380
rect 43 2266 429 2334
rect 43 2220 54 2266
rect 100 2220 168 2266
rect 214 2220 429 2266
rect 43 2152 429 2220
rect 43 2106 54 2152
rect 100 2106 168 2152
rect 214 2106 429 2152
rect 43 2038 429 2106
rect 43 1992 54 2038
rect 100 1992 168 2038
rect 214 1992 429 2038
rect 43 1924 429 1992
rect 43 1878 54 1924
rect 100 1878 168 1924
rect 214 1878 429 1924
rect 43 1810 429 1878
rect 43 1764 54 1810
rect 100 1764 168 1810
rect 214 1764 429 1810
rect 43 1696 429 1764
rect 43 1650 54 1696
rect 100 1650 168 1696
rect 214 1650 429 1696
rect 43 1582 429 1650
rect 43 1536 54 1582
rect 100 1536 168 1582
rect 214 1536 429 1582
rect 43 1468 429 1536
rect 43 1422 54 1468
rect 100 1422 168 1468
rect 214 1422 429 1468
rect 43 1354 429 1422
rect 43 1308 54 1354
rect 100 1308 168 1354
rect 214 1308 429 1354
rect 43 1240 429 1308
rect 43 1194 54 1240
rect 100 1194 168 1240
rect 214 1194 429 1240
rect 43 1126 429 1194
rect 43 1080 54 1126
rect 100 1080 168 1126
rect 214 1080 429 1126
rect 43 1012 429 1080
rect 43 966 54 1012
rect 100 966 168 1012
rect 214 966 429 1012
rect 43 898 429 966
rect 43 852 54 898
rect 100 852 168 898
rect 214 852 429 898
rect 43 784 429 852
rect 43 738 54 784
rect 100 738 168 784
rect 214 738 429 784
rect 43 621 429 738
rect 10173 621 10383 5771
rect 43 328 225 621
rect 689 531 2605 599
rect 3125 531 5041 599
rect 5561 531 7477 599
rect 7997 531 9913 599
rect 689 399 9913 531
rect 43 282 54 328
rect 100 282 168 328
rect 214 282 225 328
rect 43 226 225 282
rect 43 214 10565 226
rect 43 168 54 214
rect 100 168 168 214
rect 214 168 10565 214
rect 43 100 10565 168
rect 43 54 54 100
rect 100 54 168 100
rect 214 54 10565 100
rect 43 42 10565 54
use M1_PSUB_CDNS_69033583165350  M1_PSUB_CDNS_69033583165350_0
timestamp 1713338890
transform 0 -1 5304 1 0 134
box -102 -5004 102 5004
use M1_PSUB_CDNS_69033583165350  M1_PSUB_CDNS_69033583165350_1
timestamp 1713338890
transform 0 -1 5304 1 0 6127
box -102 -5004 102 5004
use M1_PSUB_CDNS_69033583165350  M1_PSUB_CDNS_69033583165350_2
timestamp 1713338890
transform 0 -1 5304 1 0 12218
box -102 -5004 102 5004
use M1_PSUB_CDNS_69033583165351  M1_PSUB_CDNS_69033583165351_0
timestamp 1713338890
transform 1 0 10474 0 1 6176
box -102 -6144 102 6144
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_0
timestamp 1713338890
transform 1 0 647 0 -1 5621
box -218 -350 2218 5092
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_1
timestamp 1713338890
transform 1 0 3083 0 -1 5621
box -218 -350 2218 5092
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_2
timestamp 1713338890
transform 1 0 5519 0 -1 5621
box -218 -350 2218 5092
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_3
timestamp 1713338890
transform 1 0 7955 0 -1 5621
box -218 -350 2218 5092
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_4
timestamp 1713338890
transform 1 0 647 0 1 6633
box -218 -350 2218 5092
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_5
timestamp 1713338890
transform 1 0 3083 0 1 6633
box -218 -350 2218 5092
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_6
timestamp 1713338890
transform 1 0 5519 0 1 6633
box -218 -350 2218 5092
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_7
timestamp 1713338890
transform 1 0 7955 0 1 6633
box -218 -350 2218 5092
<< labels >>
rlabel metal1 s 5302 6126 5302 6126 4 VMINUS
port 1 nsew
<< end >>
