magic
tech gf180mcuD
magscale 1 10
timestamp 1713277963
<< checkpaint >>
rect -8012 -10693 3961 -1553
<< nwell >>
rect -5337 -3607 -5228 -3605
rect -5440 -3684 -5228 -3607
rect -5440 -3685 -5333 -3684
rect -2396 -4661 -1957 -3581
rect -2396 -4731 -2395 -4661
rect -1958 -4731 -1957 -4661
rect -2456 -7640 -2396 -7390
rect -2456 -8317 -1959 -7640
rect -2396 -8567 -1959 -8317
<< nsubdiff >>
rect -5337 -3607 -5228 -3605
rect -5440 -3622 -5228 -3607
rect -5440 -3668 -5305 -3622
rect -5259 -3668 -5228 -3622
rect -5440 -3684 -5228 -3668
rect -5440 -3685 -5333 -3684
<< nsubdiffcont >>
rect -5305 -3668 -5259 -3622
<< metal1 >>
rect -5337 -3607 -5228 -3604
rect -5440 -3622 -5228 -3607
rect -5440 -3668 -5305 -3622
rect -5259 -3668 -5228 -3622
rect -5440 -3684 -5228 -3668
rect -5190 -3684 -4936 -3604
rect -2407 -3683 -1883 -3623
rect 12 -3636 126 -3608
rect -5440 -3685 -5333 -3684
rect 12 -3688 38 -3636
rect 90 -3688 126 -3636
rect 12 -3720 126 -3688
rect -2178 -4272 -2093 -4270
rect -2178 -4286 -2082 -4272
rect -2178 -4338 -2155 -4286
rect -2103 -4325 -2082 -4286
rect 164 -4308 192 -4229
rect -2103 -4338 -2093 -4325
rect -2178 -4352 -2093 -4338
rect -6012 -8622 -5965 -4457
rect -5056 -4562 -4943 -4482
rect -2150 -4710 -2095 -4652
rect -2150 -4781 -2017 -4710
rect 302 -4735 554 -4689
rect -2137 -4782 -2017 -4781
rect -5771 -5820 -5678 -5019
rect -5530 -5820 -5437 -5015
rect -2117 -5020 -2037 -5013
rect -2128 -5033 -2033 -5020
rect -2128 -5085 -2107 -5033
rect -2055 -5085 -2033 -5033
rect -2128 -5092 -2033 -5085
rect -5102 -5669 -5024 -5665
rect -5138 -5678 -5024 -5669
rect -5138 -5730 -5088 -5678
rect -5036 -5730 -5024 -5678
rect -5138 -5743 -5024 -5730
rect -5138 -5744 -5073 -5743
rect -5771 -5855 -5437 -5820
rect -5771 -5909 -5268 -5855
rect -5771 -5913 -5437 -5909
rect -5573 -5914 -5437 -5913
rect -5830 -6291 -5272 -6244
rect -5830 -7129 -5769 -6291
rect -5659 -6293 -5272 -6291
rect -5659 -7140 -5568 -6293
rect -3472 -6296 -3378 -5884
rect -5058 -6473 -5046 -6424
rect -2533 -6491 -2455 -6473
rect -2533 -6543 -2515 -6491
rect -2463 -6543 -2455 -6491
rect -2533 -6559 -2455 -6543
rect -2117 -7448 -2037 -5092
rect -687 -5300 -632 -5299
rect -687 -5352 -686 -5300
rect -634 -5352 -632 -5300
rect -687 -5353 -632 -5352
rect 508 -5819 554 -4735
rect -1075 -5865 554 -5819
rect -1075 -6059 -1006 -5865
rect -1088 -6076 -1006 -6059
rect -1088 -6128 -1074 -6076
rect -1022 -6081 -1006 -6076
rect -1022 -6128 -1007 -6081
rect -1088 -6141 -1007 -6128
rect -685 -6245 -630 -6244
rect -685 -6297 -684 -6245
rect -632 -6297 -630 -6245
rect -685 -6298 -630 -6297
rect -1205 -6424 -1134 -6413
rect -1205 -6426 -1057 -6424
rect -1205 -6478 -1191 -6426
rect -1139 -6473 -1057 -6426
rect -1139 -6478 -1134 -6473
rect -1205 -6491 -1134 -6478
rect -1841 -7093 -1771 -7089
rect -1841 -7145 -1831 -7093
rect -1779 -7145 -1771 -7093
rect -1841 -7151 -1771 -7145
rect -2192 -7495 -2037 -7448
rect 1810 -7495 1844 -7448
rect -2117 -7497 -2037 -7495
rect -1079 -7612 -1015 -7597
rect -5064 -7667 -5037 -7618
rect -2190 -7678 -1942 -7626
rect -1079 -7664 -1074 -7612
rect -1022 -7664 -1015 -7612
rect -1079 -7678 -1015 -7664
rect -2190 -8340 -2138 -7678
rect -2204 -8354 -2126 -8340
rect -2204 -8406 -2190 -8354
rect -2138 -8406 -2126 -8354
rect -2204 -8417 -2126 -8406
rect -2421 -8531 -1841 -8478
rect -2206 -8622 -2127 -8617
rect -6012 -8625 -2127 -8622
rect -6012 -8669 -2192 -8625
rect -2206 -8677 -2192 -8669
rect -2140 -8677 -2127 -8625
rect -2206 -8693 -2127 -8677
<< via1 >>
rect 38 -3688 90 -3636
rect -2155 -4338 -2103 -4286
rect -2107 -5085 -2055 -5033
rect -5088 -5730 -5036 -5678
rect -2515 -6543 -2463 -6491
rect -686 -5352 -634 -5300
rect -1074 -6128 -1022 -6076
rect -684 -6297 -632 -6245
rect -1191 -6478 -1139 -6426
rect -1831 -7145 -1779 -7093
rect -1074 -7664 -1022 -7612
rect -2190 -8406 -2138 -8354
rect -2192 -8677 -2140 -8625
<< metal2 >>
rect 8 -3636 126 -3608
rect 8 -3688 38 -3636
rect 90 -3688 126 -3636
rect 8 -3720 126 -3688
rect -2178 -4271 -2093 -4270
rect -2178 -4286 -2087 -4271
rect -2178 -4338 -2155 -4286
rect -2103 -4338 -2087 -4286
rect -2178 -4352 -2087 -4338
rect -2160 -4957 -2087 -4352
rect -2162 -5020 -2071 -4957
rect -2162 -5033 -2033 -5020
rect -2162 -5045 -2107 -5033
rect -2128 -5085 -2107 -5045
rect -2055 -5085 -2033 -5033
rect -2128 -5092 -2033 -5085
rect -700 -5300 -618 -5292
rect -700 -5352 -686 -5300
rect -634 -5352 -618 -5300
rect -5102 -5678 -5024 -5665
rect -5102 -5730 -5088 -5678
rect -5036 -5730 -5024 -5678
rect -5102 -5743 -5024 -5730
rect -5090 -5998 -5034 -5743
rect -5090 -6054 -1217 -5998
rect -1273 -6413 -1217 -6054
rect -1088 -6076 -1007 -6059
rect -1088 -6128 -1074 -6076
rect -1022 -6128 -1007 -6076
rect -1088 -6141 -1007 -6128
rect -1273 -6426 -1134 -6413
rect -2533 -6488 -2455 -6473
rect -1273 -6478 -1191 -6426
rect -1139 -6478 -1134 -6426
rect -1273 -6480 -1134 -6478
rect -2533 -6489 -2401 -6488
rect -2533 -6491 -1776 -6489
rect -1205 -6491 -1134 -6480
rect -2533 -6543 -2515 -6491
rect -2463 -6543 -1776 -6491
rect -2533 -6546 -1776 -6543
rect -2533 -6559 -2455 -6546
rect -1833 -7086 -1776 -6546
rect -1846 -7093 -1764 -7086
rect -1846 -7145 -1831 -7093
rect -1779 -7145 -1764 -7093
rect -1846 -7161 -1764 -7145
rect -1077 -7598 -1016 -6141
rect -694 -6236 -623 -5352
rect -169 -5610 -97 -5601
rect 28 -5610 100 -3720
rect -169 -5682 104 -5610
rect -697 -6245 -618 -6236
rect -697 -6297 -684 -6245
rect -632 -6297 -618 -6245
rect -697 -6304 -618 -6297
rect -169 -7213 -97 -5682
rect -957 -7285 -97 -7213
rect -957 -7336 -885 -7285
rect -1079 -7612 -1015 -7598
rect -1079 -7664 -1074 -7612
rect -1022 -7664 -1015 -7612
rect -1079 -7678 -1015 -7664
rect -2204 -8354 -2126 -8340
rect -2204 -8406 -2190 -8354
rect -2138 -8406 -2126 -8354
rect -2204 -8417 -2126 -8406
rect -2193 -8617 -2137 -8417
rect -2206 -8625 -2127 -8617
rect -2206 -8677 -2192 -8625
rect -2140 -8677 -2127 -8625
rect -2206 -8693 -2127 -8677
use mux_magic  mux_magic_0
timestamp 1713277963
transform 1 0 -4332 0 1 -5117
box -1637 -810 2187 1564
use mux_magic  mux_magic_2
timestamp 1713277963
transform 1 0 -356 0 -1 -7031
box -1637 -810 2187 1564
use mux_magic  mux_magic_3
timestamp 1713277963
transform 1 0 -4332 0 -1 -7031
box -1637 -810 2187 1564
use tspc2_magic  tspc2_magic_0
timestamp 1713185578
transform 1 0 -2109 0 1 -4247
box 9 -1127 2457 666
<< labels >>
flabel nsubdiffcont -5282 -3643 -5282 -3643 0 FreeSans 750 0 0 0 VDD
flabel metal1 s -5991 -6620 -5991 -6620 0 FreeSans 750 0 0 0 LD
port 1 nsew
flabel metal1 s 1833 -7471 1833 -7471 0 FreeSans 750 0 0 0 Q
port 2 nsew
flabel metal1 s 181 -4262 181 -4262 0 FreeSans 750 0 0 0 QB
port 3 nsew
flabel metal1 s -5125 -5711 -5125 -5711 0 FreeSans 750 0 0 0 DATA
port 4 nsew
flabel metal1 s -5014 -4550 -5014 -4550 0 FreeSans 750 0 0 0 D1
port 5 nsew
flabel metal1 s -5052 -6451 -5052 -6451 0 FreeSans 750 0 0 0 G-CLK
port 6 nsew
flabel metal1 s -5050 -7640 -5050 -7640 0 FreeSans 750 0 0 0 CLK
port 7 nsew
flabel metal1 s -5622 -5877 -5622 -5877 0 FreeSans 1250 0 0 0 VSS
port 8 nsew
<< end >>
