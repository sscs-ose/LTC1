magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2747 -2051 15709 48134
<< nwell >>
rect 2170 27755 10792 29293
<< psubdiff >>
rect 2253 27417 10709 27507
rect 2253 27178 2343 27417
rect 10619 27178 10709 27417
rect 2253 25802 2343 25866
rect 10619 25802 10709 25866
rect 2253 25780 10709 25802
rect 2253 25734 2275 25780
rect 6739 25734 6975 25780
rect 7209 25734 7445 25780
rect 7679 25734 8009 25780
rect 10687 25734 10709 25780
rect 2253 25712 10709 25734
<< psubdiffcont >>
rect 2275 25734 6739 25780
rect 6975 25734 7209 25780
rect 7445 25734 7679 25780
rect 8009 25734 10687 25780
<< polysilicon >>
rect 2665 27729 2805 27873
rect 2909 27729 3049 27873
rect 3153 27729 3293 27873
rect 3397 27729 3537 27873
rect 2665 27645 3537 27729
rect 3641 27729 3781 27873
rect 3885 27729 4025 27873
rect 4129 27729 4269 27873
rect 3641 27645 4269 27729
rect 4545 27729 4685 27873
rect 4789 27729 4929 27873
rect 5033 27729 5173 27873
rect 4545 27645 5173 27729
rect 5277 27729 5417 27873
rect 5521 27729 5661 27873
rect 5765 27729 5905 27873
rect 5277 27645 5905 27729
rect 6009 27729 6149 27873
rect 6253 27729 6393 27873
rect 6497 27729 6637 27873
rect 6009 27645 6637 27729
rect 6741 27729 6881 27873
rect 6985 27729 7125 27873
rect 7229 27729 7369 27873
rect 6741 27645 7369 27729
rect 7473 27729 7613 27873
rect 7717 27729 7857 27873
rect 7961 27729 8101 27873
rect 7473 27645 8101 27729
rect 8205 27729 8345 27873
rect 8449 27729 8589 27873
rect 8693 27729 8833 27873
rect 8205 27645 8833 27729
rect 8937 27729 9077 27873
rect 9181 27729 9321 27873
rect 9425 27729 9565 27873
rect 8937 27645 9565 27729
rect 9669 27729 9809 27873
rect 9913 27729 10053 27873
rect 10157 27729 10297 27873
rect 9669 27645 10297 27729
rect 5191 27194 5819 27278
rect 4129 27050 4269 27150
rect 5191 27050 5331 27194
rect 5435 27050 5575 27194
rect 5679 27050 5819 27194
rect 5923 27194 6551 27278
rect 5923 27050 6063 27194
rect 6167 27050 6307 27194
rect 6411 27050 6551 27194
rect 6655 27194 7283 27278
rect 6655 27050 6795 27194
rect 6899 27050 7039 27194
rect 7143 27050 7283 27194
rect 7387 27194 8015 27278
rect 7387 27050 7527 27194
rect 7631 27050 7771 27194
rect 7875 27050 8015 27194
<< metal1 >>
rect -50 27721 110 30038
rect 1473 29123 2332 29199
rect 2264 29045 2332 29123
rect 2575 27917 2651 29199
rect 2819 27857 2895 28917
rect 3063 27917 3139 29199
rect 3307 27857 3383 28917
rect 3551 27917 3627 29199
rect 4033 29123 4115 29199
rect 3795 27857 3871 28917
rect 4039 27917 4115 29123
rect 4283 27857 4359 28917
rect 4455 27917 4531 29199
rect 2819 27781 3627 27857
rect 3795 27781 4359 27857
rect 4699 27857 4775 28917
rect 4943 27917 5019 29199
rect 5187 27857 5263 28917
rect 5431 27917 5507 29199
rect 5675 27857 5751 28917
rect 5919 27917 5995 29199
rect 6163 27857 6239 28917
rect 6407 27917 6483 29199
rect 6651 27857 6727 28917
rect 6895 27917 6971 29199
rect 7139 27857 7215 28917
rect 7383 27917 7459 29199
rect 7627 27857 7703 28917
rect 7871 27917 7947 29199
rect 8115 27857 8191 28917
rect 8359 27917 8435 29199
rect 8847 29123 8929 29199
rect 8603 27857 8679 28917
rect 8847 27917 8923 29123
rect 9091 27857 9167 28917
rect 9335 27917 9411 29199
rect 9579 27857 9655 28917
rect 9823 27917 9899 29199
rect 10067 27857 10143 28917
rect 10311 27917 10387 29199
rect 10630 29123 11489 29199
rect 10630 29045 10698 29123
rect 4699 27781 10433 27857
rect 3551 27725 3627 27781
rect -50 27521 3464 27721
rect 3388 27146 3464 27521
rect 3551 27649 4224 27725
rect 4283 27721 4359 27781
rect 3551 27274 3627 27649
rect 4283 27645 10275 27721
rect 3551 27198 6516 27274
rect 3388 27070 4223 27146
rect 2264 25791 2332 25877
rect 4039 25799 4115 27006
rect 4283 26006 4359 27198
rect 6652 27142 6728 27645
rect 10357 27142 10433 27781
rect 5345 27066 6728 27142
rect 6809 27066 10433 27142
rect 4033 25791 4115 25799
rect 5101 25791 5177 27006
rect 5345 26006 5421 27066
rect 5589 25791 5665 27006
rect 5833 26006 5909 27066
rect 6077 25791 6153 27006
rect 6321 26006 6397 27066
rect 6565 25791 6641 27006
rect 2264 25780 6759 25791
rect 2264 25734 2275 25780
rect 6739 25734 6759 25780
rect 2264 25723 6759 25734
rect 6809 25617 6885 27066
rect 7053 25791 7129 27006
rect 7297 25916 7373 27066
rect 7541 25791 7617 27006
rect 7785 25916 7861 27066
rect 8029 25791 8105 27006
rect 10630 25791 10698 25877
rect 6935 25780 10698 25791
rect 6935 25734 6975 25780
rect 7209 25734 7445 25780
rect 7679 25734 8009 25780
rect 10687 25734 10698 25780
rect 6935 25723 10698 25734
rect 1213 25417 11749 25617
<< metal2 >>
rect -747 25617 1153 46134
rect 1473 25617 1673 46134
rect 1733 25617 3783 46134
rect 3843 25617 4043 46134
rect 4103 25617 6153 46134
rect 6213 25617 6749 46134
rect 6809 25617 8859 46134
rect 8919 25617 9119 46134
rect 9179 25617 11229 46134
rect 11289 25617 11489 46134
rect 11809 25617 13709 46134
use comp018green_esd_rc_v5p0  comp018green_esd_rc_v5p0_0
timestamp 1713338890
transform 1 0 -356 0 -1 46507
box -51 491 13725 17038
use M1_NWELL_CDNS_40661953145107  M1_NWELL_CDNS_40661953145107_0
timestamp 1713338890
transform 1 0 6481 0 1 29165
box -4311 -128 4311 128
use M1_NWELL_CDNS_40661953145111  M1_NWELL_CDNS_40661953145111_0
timestamp 1713338890
transform 1 0 2298 0 1 28447
box -128 -692 128 692
use M1_NWELL_CDNS_40661953145111  M1_NWELL_CDNS_40661953145111_1
timestamp 1713338890
transform 1 0 10664 0 1 28447
box -128 -692 128 692
use M1_POLY2_CDNS_69033583165343  M1_POLY2_CDNS_69033583165343_0
timestamp 1713338890
transform 1 0 7421 0 1 27687
box -2862 -42 2862 42
use M1_POLY2_CDNS_69033583165344  M1_POLY2_CDNS_69033583165344_0
timestamp 1713338890
transform 1 0 5871 0 1 27236
box -653 -42 653 42
use M1_POLY2_CDNS_69033583165344  M1_POLY2_CDNS_69033583165344_1
timestamp 1713338890
transform 1 0 7335 0 1 27236
box -653 -42 653 42
use M1_POLY2_CDNS_69033583165345  M1_POLY2_CDNS_69033583165345_0
timestamp 1713338890
transform 1 0 3955 0 1 27687
box -277 -42 277 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_0
timestamp 1713338890
transform 1 0 4142 0 1 27108
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165347  M1_POLY2_CDNS_69033583165347_0
timestamp 1713338890
transform 1 0 3101 0 1 27687
box -371 -42 371 42
use M1_PSUB_CDNS_69033583165349  M1_PSUB_CDNS_69033583165349_0
timestamp 1713338890
transform 1 0 2298 0 -1 26522
box -45 -656 45 656
use M1_PSUB_CDNS_69033583165349  M1_PSUB_CDNS_69033583165349_1
timestamp 1713338890
transform 1 0 10664 0 -1 26522
box -45 -656 45 656
use M1_PSUB_CDNS_69033583165519  M1_PSUB_CDNS_69033583165519_0
timestamp 1713338890
transform 1 0 8557 0 1 27462
box -1690 -45 1690 45
use M1_PSUB_CDNS_69033583165520  M1_PSUB_CDNS_69033583165520_0
timestamp 1713338890
transform 1 0 5134 0 1 27462
box -1408 -45 1408 45
use M2_M1_CDNS_69033583165348  M2_M1_CDNS_69033583165348_0
timestamp 1713338890
transform 1 0 1313 0 1 25517
box -92 -92 92 92
use M2_M1_CDNS_69033583165348  M2_M1_CDNS_69033583165348_1
timestamp 1713338890
transform 1 0 11649 0 1 25517
box -92 -92 92 92
use M2_M1_CDNS_69033583165506  M2_M1_CDNS_69033583165506_0
timestamp 1713338890
transform 1 0 2758 0 1 29571
box -1010 -92 1010 92
use M2_M1_CDNS_69033583165506  M2_M1_CDNS_69033583165506_1
timestamp 1713338890
transform 1 0 7834 0 1 29571
box -1010 -92 1010 92
use M2_M1_CDNS_69033583165506  M2_M1_CDNS_69033583165506_2
timestamp 1713338890
transform 1 0 10204 0 1 29571
box -1010 -92 1010 92
use M2_M1_CDNS_69033583165506  M2_M1_CDNS_69033583165506_3
timestamp 1713338890
transform 1 0 5128 0 1 29571
box -1010 -92 1010 92
use M2_M1_CDNS_69033583165506  M2_M1_CDNS_69033583165506_4
timestamp 1713338890
transform 1 0 2758 0 1 41655
box -1010 -92 1010 92
use M2_M1_CDNS_69033583165506  M2_M1_CDNS_69033583165506_5
timestamp 1713338890
transform 1 0 5128 0 1 41655
box -1010 -92 1010 92
use M2_M1_CDNS_69033583165506  M2_M1_CDNS_69033583165506_6
timestamp 1713338890
transform 1 0 7834 0 1 41655
box -1010 -92 1010 92
use M2_M1_CDNS_69033583165506  M2_M1_CDNS_69033583165506_7
timestamp 1713338890
transform 1 0 10204 0 1 41655
box -1010 -92 1010 92
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_0
timestamp 1713338890
transform 1 0 1573 0 1 42148
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_1
timestamp 1713338890
transform 1 0 3943 0 1 42148
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_2
timestamp 1713338890
transform 1 0 11389 0 1 42148
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_3
timestamp 1713338890
transform 1 0 9019 0 1 42148
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_4
timestamp 1713338890
transform 1 0 1573 0 1 45888
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_5
timestamp 1713338890
transform 1 0 3943 0 1 45888
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_6
timestamp 1713338890
transform 1 0 11389 0 1 45888
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_7
timestamp 1713338890
transform 1 0 9019 0 1 45888
box -92 -38 92 38
use M2_M1_CDNS_69033583165515  M2_M1_CDNS_69033583165515_0
timestamp 1713338890
transform 1 0 9730 0 1 27458
box -506 -38 506 38
use M2_M1_CDNS_69033583165516  M2_M1_CDNS_69033583165516_0
timestamp 1713338890
transform 1 0 2758 0 1 35662
box -968 -348 968 348
use M2_M1_CDNS_69033583165516  M2_M1_CDNS_69033583165516_1
timestamp 1713338890
transform 1 0 5128 0 1 35662
box -968 -348 968 348
use M2_M1_CDNS_69033583165516  M2_M1_CDNS_69033583165516_2
timestamp 1713338890
transform 1 0 7834 0 1 35662
box -968 -348 968 348
use M2_M1_CDNS_69033583165516  M2_M1_CDNS_69033583165516_3
timestamp 1713338890
transform 1 0 10204 0 1 35662
box -968 -348 968 348
use M2_M1_CDNS_69033583165517  M2_M1_CDNS_69033583165517_0
timestamp 1713338890
transform 1 0 2978 0 1 25753
box -714 -38 714 38
use M2_M1_CDNS_69033583165517  M2_M1_CDNS_69033583165517_1
timestamp 1713338890
transform -1 0 9984 0 1 25753
box -714 -38 714 38
use M2_M1_CDNS_69033583165518  M2_M1_CDNS_69033583165518_0
timestamp 1713338890
transform 1 0 7089 0 1 25753
box -142 -38 142 38
use M2_M1_CDNS_69033583165518  M2_M1_CDNS_69033583165518_1
timestamp 1713338890
transform 1 0 7578 0 1 25753
box -142 -38 142 38
use M2_M1_CDNS_69033583165521  M2_M1_CDNS_69033583165521_0
timestamp 1713338890
transform 1 0 2302 0 1 26557
box -38 -610 38 610
use M2_M1_CDNS_69033583165521  M2_M1_CDNS_69033583165521_1
timestamp 1713338890
transform -1 0 10660 0 1 26557
box -38 -610 38 610
use M2_M1_CDNS_69033583165522  M2_M1_CDNS_69033583165522_0
timestamp 1713338890
transform 1 0 5128 0 1 25753
box -974 -38 974 38
use M2_M1_CDNS_69033583165522  M2_M1_CDNS_69033583165522_1
timestamp 1713338890
transform 1 0 5128 0 1 27458
box -974 -38 974 38
use M2_M1_CDNS_69033583165522  M2_M1_CDNS_69033583165522_2
timestamp 1713338890
transform 1 0 7834 0 1 27458
box -974 -38 974 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_0
timestamp 1713338890
transform 1 0 1573 0 1 29161
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_1
timestamp 1713338890
transform -1 0 11389 0 1 29161
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_2
timestamp 1713338890
transform -1 0 9019 0 1 29161
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_3
timestamp 1713338890
transform -1 0 3943 0 1 29161
box -90 -38 90 38
use M2_M1_CDNS_69033583165524  M2_M1_CDNS_69033583165524_0
timestamp 1713338890
transform 1 0 8405 0 1 25753
box -454 -38 454 38
use M2_M1_CDNS_69033583165525  M2_M1_CDNS_69033583165525_0
timestamp 1713338890
transform -1 0 6481 0 1 29161
box -246 -38 246 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_0
timestamp 1713338890
transform 1 0 6481 0 1 42148
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_1
timestamp 1713338890
transform 1 0 6481 0 1 45888
box -254 -38 254 38
use nmos_6p0_CDNS_406619531458  nmos_6p0_CDNS_406619531458_0
timestamp 1713338890
transform 1 0 5191 0 1 26006
box -88 -44 1448 1044
use nmos_6p0_CDNS_406619531458  nmos_6p0_CDNS_406619531458_1
timestamp 1713338890
transform 1 0 6655 0 1 26006
box -88 -44 1448 1044
use nmos_6p0_CDNS_406619531459  nmos_6p0_CDNS_406619531459_0
timestamp 1713338890
transform 1 0 4129 0 1 26006
box -88 -44 228 1044
use nmos_clamp_20_50_4_DVSS  nmos_clamp_20_50_4_DVSS_0
timestamp 1713338890
transform 1 0 0 0 1 0
box -747 -51 13709 25617
use pmos_6p0_CDNS_406619531452  pmos_6p0_CDNS_406619531452_0
timestamp 1713338890
transform 1 0 2665 0 1 27917
box -208 -120 1080 1120
use pmos_6p0_CDNS_406619531455  pmos_6p0_CDNS_406619531455_0
timestamp 1713338890
transform 1 0 4545 0 1 27917
box -208 -120 5960 1120
use pmos_6p0_CDNS_406619531456  pmos_6p0_CDNS_406619531456_0
timestamp 1713338890
transform 1 0 3641 0 1 27917
box -208 -120 836 1120
<< end >>
