magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -14941 -2097 14941 2097
<< psubdiff >>
rect -12941 75 12941 97
rect -12941 29 -12919 75
rect -12873 29 -12815 75
rect -12769 29 -12711 75
rect -12665 29 -12607 75
rect -12561 29 -12503 75
rect -12457 29 -12399 75
rect -12353 29 -12295 75
rect -12249 29 -12191 75
rect -12145 29 -12087 75
rect -12041 29 -11983 75
rect -11937 29 -11879 75
rect -11833 29 -11775 75
rect -11729 29 -11671 75
rect -11625 29 -11567 75
rect -11521 29 -11463 75
rect -11417 29 -11359 75
rect -11313 29 -11255 75
rect -11209 29 -11151 75
rect -11105 29 -11047 75
rect -11001 29 -10943 75
rect -10897 29 -10839 75
rect -10793 29 -10735 75
rect -10689 29 -10631 75
rect -10585 29 -10527 75
rect -10481 29 -10423 75
rect -10377 29 -10319 75
rect -10273 29 -10215 75
rect -10169 29 -10111 75
rect -10065 29 -10007 75
rect -9961 29 -9903 75
rect -9857 29 -9799 75
rect -9753 29 -9695 75
rect -9649 29 -9591 75
rect -9545 29 -9487 75
rect -9441 29 -9383 75
rect -9337 29 -9279 75
rect -9233 29 -9175 75
rect -9129 29 -9071 75
rect -9025 29 -8967 75
rect -8921 29 -8863 75
rect -8817 29 -8759 75
rect -8713 29 -8655 75
rect -8609 29 -8551 75
rect -8505 29 -8447 75
rect -8401 29 -8343 75
rect -8297 29 -8239 75
rect -8193 29 -8135 75
rect -8089 29 -8031 75
rect -7985 29 -7927 75
rect -7881 29 -7823 75
rect -7777 29 -7719 75
rect -7673 29 -7615 75
rect -7569 29 -7511 75
rect -7465 29 -7407 75
rect -7361 29 -7303 75
rect -7257 29 -7199 75
rect -7153 29 -7095 75
rect -7049 29 -6991 75
rect -6945 29 -6887 75
rect -6841 29 -6783 75
rect -6737 29 -6679 75
rect -6633 29 -6575 75
rect -6529 29 -6471 75
rect -6425 29 -6367 75
rect -6321 29 -6263 75
rect -6217 29 -6159 75
rect -6113 29 -6055 75
rect -6009 29 -5951 75
rect -5905 29 -5847 75
rect -5801 29 -5743 75
rect -5697 29 -5639 75
rect -5593 29 -5535 75
rect -5489 29 -5431 75
rect -5385 29 -5327 75
rect -5281 29 -5223 75
rect -5177 29 -5119 75
rect -5073 29 -5015 75
rect -4969 29 -4911 75
rect -4865 29 -4807 75
rect -4761 29 -4703 75
rect -4657 29 -4599 75
rect -4553 29 -4495 75
rect -4449 29 -4391 75
rect -4345 29 -4287 75
rect -4241 29 -4183 75
rect -4137 29 -4079 75
rect -4033 29 -3975 75
rect -3929 29 -3871 75
rect -3825 29 -3767 75
rect -3721 29 -3663 75
rect -3617 29 -3559 75
rect -3513 29 -3455 75
rect -3409 29 -3351 75
rect -3305 29 -3247 75
rect -3201 29 -3143 75
rect -3097 29 -3039 75
rect -2993 29 -2935 75
rect -2889 29 -2831 75
rect -2785 29 -2727 75
rect -2681 29 -2623 75
rect -2577 29 -2519 75
rect -2473 29 -2415 75
rect -2369 29 -2311 75
rect -2265 29 -2207 75
rect -2161 29 -2103 75
rect -2057 29 -1999 75
rect -1953 29 -1895 75
rect -1849 29 -1791 75
rect -1745 29 -1687 75
rect -1641 29 -1583 75
rect -1537 29 -1479 75
rect -1433 29 -1375 75
rect -1329 29 -1271 75
rect -1225 29 -1167 75
rect -1121 29 -1063 75
rect -1017 29 -959 75
rect -913 29 -855 75
rect -809 29 -751 75
rect -705 29 -647 75
rect -601 29 -543 75
rect -497 29 -439 75
rect -393 29 -335 75
rect -289 29 -231 75
rect -185 29 -127 75
rect -81 29 -23 75
rect 23 29 81 75
rect 127 29 185 75
rect 231 29 289 75
rect 335 29 393 75
rect 439 29 497 75
rect 543 29 601 75
rect 647 29 705 75
rect 751 29 809 75
rect 855 29 913 75
rect 959 29 1017 75
rect 1063 29 1121 75
rect 1167 29 1225 75
rect 1271 29 1329 75
rect 1375 29 1433 75
rect 1479 29 1537 75
rect 1583 29 1641 75
rect 1687 29 1745 75
rect 1791 29 1849 75
rect 1895 29 1953 75
rect 1999 29 2057 75
rect 2103 29 2161 75
rect 2207 29 2265 75
rect 2311 29 2369 75
rect 2415 29 2473 75
rect 2519 29 2577 75
rect 2623 29 2681 75
rect 2727 29 2785 75
rect 2831 29 2889 75
rect 2935 29 2993 75
rect 3039 29 3097 75
rect 3143 29 3201 75
rect 3247 29 3305 75
rect 3351 29 3409 75
rect 3455 29 3513 75
rect 3559 29 3617 75
rect 3663 29 3721 75
rect 3767 29 3825 75
rect 3871 29 3929 75
rect 3975 29 4033 75
rect 4079 29 4137 75
rect 4183 29 4241 75
rect 4287 29 4345 75
rect 4391 29 4449 75
rect 4495 29 4553 75
rect 4599 29 4657 75
rect 4703 29 4761 75
rect 4807 29 4865 75
rect 4911 29 4969 75
rect 5015 29 5073 75
rect 5119 29 5177 75
rect 5223 29 5281 75
rect 5327 29 5385 75
rect 5431 29 5489 75
rect 5535 29 5593 75
rect 5639 29 5697 75
rect 5743 29 5801 75
rect 5847 29 5905 75
rect 5951 29 6009 75
rect 6055 29 6113 75
rect 6159 29 6217 75
rect 6263 29 6321 75
rect 6367 29 6425 75
rect 6471 29 6529 75
rect 6575 29 6633 75
rect 6679 29 6737 75
rect 6783 29 6841 75
rect 6887 29 6945 75
rect 6991 29 7049 75
rect 7095 29 7153 75
rect 7199 29 7257 75
rect 7303 29 7361 75
rect 7407 29 7465 75
rect 7511 29 7569 75
rect 7615 29 7673 75
rect 7719 29 7777 75
rect 7823 29 7881 75
rect 7927 29 7985 75
rect 8031 29 8089 75
rect 8135 29 8193 75
rect 8239 29 8297 75
rect 8343 29 8401 75
rect 8447 29 8505 75
rect 8551 29 8609 75
rect 8655 29 8713 75
rect 8759 29 8817 75
rect 8863 29 8921 75
rect 8967 29 9025 75
rect 9071 29 9129 75
rect 9175 29 9233 75
rect 9279 29 9337 75
rect 9383 29 9441 75
rect 9487 29 9545 75
rect 9591 29 9649 75
rect 9695 29 9753 75
rect 9799 29 9857 75
rect 9903 29 9961 75
rect 10007 29 10065 75
rect 10111 29 10169 75
rect 10215 29 10273 75
rect 10319 29 10377 75
rect 10423 29 10481 75
rect 10527 29 10585 75
rect 10631 29 10689 75
rect 10735 29 10793 75
rect 10839 29 10897 75
rect 10943 29 11001 75
rect 11047 29 11105 75
rect 11151 29 11209 75
rect 11255 29 11313 75
rect 11359 29 11417 75
rect 11463 29 11521 75
rect 11567 29 11625 75
rect 11671 29 11729 75
rect 11775 29 11833 75
rect 11879 29 11937 75
rect 11983 29 12041 75
rect 12087 29 12145 75
rect 12191 29 12249 75
rect 12295 29 12353 75
rect 12399 29 12457 75
rect 12503 29 12561 75
rect 12607 29 12665 75
rect 12711 29 12769 75
rect 12815 29 12873 75
rect 12919 29 12941 75
rect -12941 -29 12941 29
rect -12941 -75 -12919 -29
rect -12873 -75 -12815 -29
rect -12769 -75 -12711 -29
rect -12665 -75 -12607 -29
rect -12561 -75 -12503 -29
rect -12457 -75 -12399 -29
rect -12353 -75 -12295 -29
rect -12249 -75 -12191 -29
rect -12145 -75 -12087 -29
rect -12041 -75 -11983 -29
rect -11937 -75 -11879 -29
rect -11833 -75 -11775 -29
rect -11729 -75 -11671 -29
rect -11625 -75 -11567 -29
rect -11521 -75 -11463 -29
rect -11417 -75 -11359 -29
rect -11313 -75 -11255 -29
rect -11209 -75 -11151 -29
rect -11105 -75 -11047 -29
rect -11001 -75 -10943 -29
rect -10897 -75 -10839 -29
rect -10793 -75 -10735 -29
rect -10689 -75 -10631 -29
rect -10585 -75 -10527 -29
rect -10481 -75 -10423 -29
rect -10377 -75 -10319 -29
rect -10273 -75 -10215 -29
rect -10169 -75 -10111 -29
rect -10065 -75 -10007 -29
rect -9961 -75 -9903 -29
rect -9857 -75 -9799 -29
rect -9753 -75 -9695 -29
rect -9649 -75 -9591 -29
rect -9545 -75 -9487 -29
rect -9441 -75 -9383 -29
rect -9337 -75 -9279 -29
rect -9233 -75 -9175 -29
rect -9129 -75 -9071 -29
rect -9025 -75 -8967 -29
rect -8921 -75 -8863 -29
rect -8817 -75 -8759 -29
rect -8713 -75 -8655 -29
rect -8609 -75 -8551 -29
rect -8505 -75 -8447 -29
rect -8401 -75 -8343 -29
rect -8297 -75 -8239 -29
rect -8193 -75 -8135 -29
rect -8089 -75 -8031 -29
rect -7985 -75 -7927 -29
rect -7881 -75 -7823 -29
rect -7777 -75 -7719 -29
rect -7673 -75 -7615 -29
rect -7569 -75 -7511 -29
rect -7465 -75 -7407 -29
rect -7361 -75 -7303 -29
rect -7257 -75 -7199 -29
rect -7153 -75 -7095 -29
rect -7049 -75 -6991 -29
rect -6945 -75 -6887 -29
rect -6841 -75 -6783 -29
rect -6737 -75 -6679 -29
rect -6633 -75 -6575 -29
rect -6529 -75 -6471 -29
rect -6425 -75 -6367 -29
rect -6321 -75 -6263 -29
rect -6217 -75 -6159 -29
rect -6113 -75 -6055 -29
rect -6009 -75 -5951 -29
rect -5905 -75 -5847 -29
rect -5801 -75 -5743 -29
rect -5697 -75 -5639 -29
rect -5593 -75 -5535 -29
rect -5489 -75 -5431 -29
rect -5385 -75 -5327 -29
rect -5281 -75 -5223 -29
rect -5177 -75 -5119 -29
rect -5073 -75 -5015 -29
rect -4969 -75 -4911 -29
rect -4865 -75 -4807 -29
rect -4761 -75 -4703 -29
rect -4657 -75 -4599 -29
rect -4553 -75 -4495 -29
rect -4449 -75 -4391 -29
rect -4345 -75 -4287 -29
rect -4241 -75 -4183 -29
rect -4137 -75 -4079 -29
rect -4033 -75 -3975 -29
rect -3929 -75 -3871 -29
rect -3825 -75 -3767 -29
rect -3721 -75 -3663 -29
rect -3617 -75 -3559 -29
rect -3513 -75 -3455 -29
rect -3409 -75 -3351 -29
rect -3305 -75 -3247 -29
rect -3201 -75 -3143 -29
rect -3097 -75 -3039 -29
rect -2993 -75 -2935 -29
rect -2889 -75 -2831 -29
rect -2785 -75 -2727 -29
rect -2681 -75 -2623 -29
rect -2577 -75 -2519 -29
rect -2473 -75 -2415 -29
rect -2369 -75 -2311 -29
rect -2265 -75 -2207 -29
rect -2161 -75 -2103 -29
rect -2057 -75 -1999 -29
rect -1953 -75 -1895 -29
rect -1849 -75 -1791 -29
rect -1745 -75 -1687 -29
rect -1641 -75 -1583 -29
rect -1537 -75 -1479 -29
rect -1433 -75 -1375 -29
rect -1329 -75 -1271 -29
rect -1225 -75 -1167 -29
rect -1121 -75 -1063 -29
rect -1017 -75 -959 -29
rect -913 -75 -855 -29
rect -809 -75 -751 -29
rect -705 -75 -647 -29
rect -601 -75 -543 -29
rect -497 -75 -439 -29
rect -393 -75 -335 -29
rect -289 -75 -231 -29
rect -185 -75 -127 -29
rect -81 -75 -23 -29
rect 23 -75 81 -29
rect 127 -75 185 -29
rect 231 -75 289 -29
rect 335 -75 393 -29
rect 439 -75 497 -29
rect 543 -75 601 -29
rect 647 -75 705 -29
rect 751 -75 809 -29
rect 855 -75 913 -29
rect 959 -75 1017 -29
rect 1063 -75 1121 -29
rect 1167 -75 1225 -29
rect 1271 -75 1329 -29
rect 1375 -75 1433 -29
rect 1479 -75 1537 -29
rect 1583 -75 1641 -29
rect 1687 -75 1745 -29
rect 1791 -75 1849 -29
rect 1895 -75 1953 -29
rect 1999 -75 2057 -29
rect 2103 -75 2161 -29
rect 2207 -75 2265 -29
rect 2311 -75 2369 -29
rect 2415 -75 2473 -29
rect 2519 -75 2577 -29
rect 2623 -75 2681 -29
rect 2727 -75 2785 -29
rect 2831 -75 2889 -29
rect 2935 -75 2993 -29
rect 3039 -75 3097 -29
rect 3143 -75 3201 -29
rect 3247 -75 3305 -29
rect 3351 -75 3409 -29
rect 3455 -75 3513 -29
rect 3559 -75 3617 -29
rect 3663 -75 3721 -29
rect 3767 -75 3825 -29
rect 3871 -75 3929 -29
rect 3975 -75 4033 -29
rect 4079 -75 4137 -29
rect 4183 -75 4241 -29
rect 4287 -75 4345 -29
rect 4391 -75 4449 -29
rect 4495 -75 4553 -29
rect 4599 -75 4657 -29
rect 4703 -75 4761 -29
rect 4807 -75 4865 -29
rect 4911 -75 4969 -29
rect 5015 -75 5073 -29
rect 5119 -75 5177 -29
rect 5223 -75 5281 -29
rect 5327 -75 5385 -29
rect 5431 -75 5489 -29
rect 5535 -75 5593 -29
rect 5639 -75 5697 -29
rect 5743 -75 5801 -29
rect 5847 -75 5905 -29
rect 5951 -75 6009 -29
rect 6055 -75 6113 -29
rect 6159 -75 6217 -29
rect 6263 -75 6321 -29
rect 6367 -75 6425 -29
rect 6471 -75 6529 -29
rect 6575 -75 6633 -29
rect 6679 -75 6737 -29
rect 6783 -75 6841 -29
rect 6887 -75 6945 -29
rect 6991 -75 7049 -29
rect 7095 -75 7153 -29
rect 7199 -75 7257 -29
rect 7303 -75 7361 -29
rect 7407 -75 7465 -29
rect 7511 -75 7569 -29
rect 7615 -75 7673 -29
rect 7719 -75 7777 -29
rect 7823 -75 7881 -29
rect 7927 -75 7985 -29
rect 8031 -75 8089 -29
rect 8135 -75 8193 -29
rect 8239 -75 8297 -29
rect 8343 -75 8401 -29
rect 8447 -75 8505 -29
rect 8551 -75 8609 -29
rect 8655 -75 8713 -29
rect 8759 -75 8817 -29
rect 8863 -75 8921 -29
rect 8967 -75 9025 -29
rect 9071 -75 9129 -29
rect 9175 -75 9233 -29
rect 9279 -75 9337 -29
rect 9383 -75 9441 -29
rect 9487 -75 9545 -29
rect 9591 -75 9649 -29
rect 9695 -75 9753 -29
rect 9799 -75 9857 -29
rect 9903 -75 9961 -29
rect 10007 -75 10065 -29
rect 10111 -75 10169 -29
rect 10215 -75 10273 -29
rect 10319 -75 10377 -29
rect 10423 -75 10481 -29
rect 10527 -75 10585 -29
rect 10631 -75 10689 -29
rect 10735 -75 10793 -29
rect 10839 -75 10897 -29
rect 10943 -75 11001 -29
rect 11047 -75 11105 -29
rect 11151 -75 11209 -29
rect 11255 -75 11313 -29
rect 11359 -75 11417 -29
rect 11463 -75 11521 -29
rect 11567 -75 11625 -29
rect 11671 -75 11729 -29
rect 11775 -75 11833 -29
rect 11879 -75 11937 -29
rect 11983 -75 12041 -29
rect 12087 -75 12145 -29
rect 12191 -75 12249 -29
rect 12295 -75 12353 -29
rect 12399 -75 12457 -29
rect 12503 -75 12561 -29
rect 12607 -75 12665 -29
rect 12711 -75 12769 -29
rect 12815 -75 12873 -29
rect 12919 -75 12941 -29
rect -12941 -97 12941 -75
<< psubdiffcont >>
rect -12919 29 -12873 75
rect -12815 29 -12769 75
rect -12711 29 -12665 75
rect -12607 29 -12561 75
rect -12503 29 -12457 75
rect -12399 29 -12353 75
rect -12295 29 -12249 75
rect -12191 29 -12145 75
rect -12087 29 -12041 75
rect -11983 29 -11937 75
rect -11879 29 -11833 75
rect -11775 29 -11729 75
rect -11671 29 -11625 75
rect -11567 29 -11521 75
rect -11463 29 -11417 75
rect -11359 29 -11313 75
rect -11255 29 -11209 75
rect -11151 29 -11105 75
rect -11047 29 -11001 75
rect -10943 29 -10897 75
rect -10839 29 -10793 75
rect -10735 29 -10689 75
rect -10631 29 -10585 75
rect -10527 29 -10481 75
rect -10423 29 -10377 75
rect -10319 29 -10273 75
rect -10215 29 -10169 75
rect -10111 29 -10065 75
rect -10007 29 -9961 75
rect -9903 29 -9857 75
rect -9799 29 -9753 75
rect -9695 29 -9649 75
rect -9591 29 -9545 75
rect -9487 29 -9441 75
rect -9383 29 -9337 75
rect -9279 29 -9233 75
rect -9175 29 -9129 75
rect -9071 29 -9025 75
rect -8967 29 -8921 75
rect -8863 29 -8817 75
rect -8759 29 -8713 75
rect -8655 29 -8609 75
rect -8551 29 -8505 75
rect -8447 29 -8401 75
rect -8343 29 -8297 75
rect -8239 29 -8193 75
rect -8135 29 -8089 75
rect -8031 29 -7985 75
rect -7927 29 -7881 75
rect -7823 29 -7777 75
rect -7719 29 -7673 75
rect -7615 29 -7569 75
rect -7511 29 -7465 75
rect -7407 29 -7361 75
rect -7303 29 -7257 75
rect -7199 29 -7153 75
rect -7095 29 -7049 75
rect -6991 29 -6945 75
rect -6887 29 -6841 75
rect -6783 29 -6737 75
rect -6679 29 -6633 75
rect -6575 29 -6529 75
rect -6471 29 -6425 75
rect -6367 29 -6321 75
rect -6263 29 -6217 75
rect -6159 29 -6113 75
rect -6055 29 -6009 75
rect -5951 29 -5905 75
rect -5847 29 -5801 75
rect -5743 29 -5697 75
rect -5639 29 -5593 75
rect -5535 29 -5489 75
rect -5431 29 -5385 75
rect -5327 29 -5281 75
rect -5223 29 -5177 75
rect -5119 29 -5073 75
rect -5015 29 -4969 75
rect -4911 29 -4865 75
rect -4807 29 -4761 75
rect -4703 29 -4657 75
rect -4599 29 -4553 75
rect -4495 29 -4449 75
rect -4391 29 -4345 75
rect -4287 29 -4241 75
rect -4183 29 -4137 75
rect -4079 29 -4033 75
rect -3975 29 -3929 75
rect -3871 29 -3825 75
rect -3767 29 -3721 75
rect -3663 29 -3617 75
rect -3559 29 -3513 75
rect -3455 29 -3409 75
rect -3351 29 -3305 75
rect -3247 29 -3201 75
rect -3143 29 -3097 75
rect -3039 29 -2993 75
rect -2935 29 -2889 75
rect -2831 29 -2785 75
rect -2727 29 -2681 75
rect -2623 29 -2577 75
rect -2519 29 -2473 75
rect -2415 29 -2369 75
rect -2311 29 -2265 75
rect -2207 29 -2161 75
rect -2103 29 -2057 75
rect -1999 29 -1953 75
rect -1895 29 -1849 75
rect -1791 29 -1745 75
rect -1687 29 -1641 75
rect -1583 29 -1537 75
rect -1479 29 -1433 75
rect -1375 29 -1329 75
rect -1271 29 -1225 75
rect -1167 29 -1121 75
rect -1063 29 -1017 75
rect -959 29 -913 75
rect -855 29 -809 75
rect -751 29 -705 75
rect -647 29 -601 75
rect -543 29 -497 75
rect -439 29 -393 75
rect -335 29 -289 75
rect -231 29 -185 75
rect -127 29 -81 75
rect -23 29 23 75
rect 81 29 127 75
rect 185 29 231 75
rect 289 29 335 75
rect 393 29 439 75
rect 497 29 543 75
rect 601 29 647 75
rect 705 29 751 75
rect 809 29 855 75
rect 913 29 959 75
rect 1017 29 1063 75
rect 1121 29 1167 75
rect 1225 29 1271 75
rect 1329 29 1375 75
rect 1433 29 1479 75
rect 1537 29 1583 75
rect 1641 29 1687 75
rect 1745 29 1791 75
rect 1849 29 1895 75
rect 1953 29 1999 75
rect 2057 29 2103 75
rect 2161 29 2207 75
rect 2265 29 2311 75
rect 2369 29 2415 75
rect 2473 29 2519 75
rect 2577 29 2623 75
rect 2681 29 2727 75
rect 2785 29 2831 75
rect 2889 29 2935 75
rect 2993 29 3039 75
rect 3097 29 3143 75
rect 3201 29 3247 75
rect 3305 29 3351 75
rect 3409 29 3455 75
rect 3513 29 3559 75
rect 3617 29 3663 75
rect 3721 29 3767 75
rect 3825 29 3871 75
rect 3929 29 3975 75
rect 4033 29 4079 75
rect 4137 29 4183 75
rect 4241 29 4287 75
rect 4345 29 4391 75
rect 4449 29 4495 75
rect 4553 29 4599 75
rect 4657 29 4703 75
rect 4761 29 4807 75
rect 4865 29 4911 75
rect 4969 29 5015 75
rect 5073 29 5119 75
rect 5177 29 5223 75
rect 5281 29 5327 75
rect 5385 29 5431 75
rect 5489 29 5535 75
rect 5593 29 5639 75
rect 5697 29 5743 75
rect 5801 29 5847 75
rect 5905 29 5951 75
rect 6009 29 6055 75
rect 6113 29 6159 75
rect 6217 29 6263 75
rect 6321 29 6367 75
rect 6425 29 6471 75
rect 6529 29 6575 75
rect 6633 29 6679 75
rect 6737 29 6783 75
rect 6841 29 6887 75
rect 6945 29 6991 75
rect 7049 29 7095 75
rect 7153 29 7199 75
rect 7257 29 7303 75
rect 7361 29 7407 75
rect 7465 29 7511 75
rect 7569 29 7615 75
rect 7673 29 7719 75
rect 7777 29 7823 75
rect 7881 29 7927 75
rect 7985 29 8031 75
rect 8089 29 8135 75
rect 8193 29 8239 75
rect 8297 29 8343 75
rect 8401 29 8447 75
rect 8505 29 8551 75
rect 8609 29 8655 75
rect 8713 29 8759 75
rect 8817 29 8863 75
rect 8921 29 8967 75
rect 9025 29 9071 75
rect 9129 29 9175 75
rect 9233 29 9279 75
rect 9337 29 9383 75
rect 9441 29 9487 75
rect 9545 29 9591 75
rect 9649 29 9695 75
rect 9753 29 9799 75
rect 9857 29 9903 75
rect 9961 29 10007 75
rect 10065 29 10111 75
rect 10169 29 10215 75
rect 10273 29 10319 75
rect 10377 29 10423 75
rect 10481 29 10527 75
rect 10585 29 10631 75
rect 10689 29 10735 75
rect 10793 29 10839 75
rect 10897 29 10943 75
rect 11001 29 11047 75
rect 11105 29 11151 75
rect 11209 29 11255 75
rect 11313 29 11359 75
rect 11417 29 11463 75
rect 11521 29 11567 75
rect 11625 29 11671 75
rect 11729 29 11775 75
rect 11833 29 11879 75
rect 11937 29 11983 75
rect 12041 29 12087 75
rect 12145 29 12191 75
rect 12249 29 12295 75
rect 12353 29 12399 75
rect 12457 29 12503 75
rect 12561 29 12607 75
rect 12665 29 12711 75
rect 12769 29 12815 75
rect 12873 29 12919 75
rect -12919 -75 -12873 -29
rect -12815 -75 -12769 -29
rect -12711 -75 -12665 -29
rect -12607 -75 -12561 -29
rect -12503 -75 -12457 -29
rect -12399 -75 -12353 -29
rect -12295 -75 -12249 -29
rect -12191 -75 -12145 -29
rect -12087 -75 -12041 -29
rect -11983 -75 -11937 -29
rect -11879 -75 -11833 -29
rect -11775 -75 -11729 -29
rect -11671 -75 -11625 -29
rect -11567 -75 -11521 -29
rect -11463 -75 -11417 -29
rect -11359 -75 -11313 -29
rect -11255 -75 -11209 -29
rect -11151 -75 -11105 -29
rect -11047 -75 -11001 -29
rect -10943 -75 -10897 -29
rect -10839 -75 -10793 -29
rect -10735 -75 -10689 -29
rect -10631 -75 -10585 -29
rect -10527 -75 -10481 -29
rect -10423 -75 -10377 -29
rect -10319 -75 -10273 -29
rect -10215 -75 -10169 -29
rect -10111 -75 -10065 -29
rect -10007 -75 -9961 -29
rect -9903 -75 -9857 -29
rect -9799 -75 -9753 -29
rect -9695 -75 -9649 -29
rect -9591 -75 -9545 -29
rect -9487 -75 -9441 -29
rect -9383 -75 -9337 -29
rect -9279 -75 -9233 -29
rect -9175 -75 -9129 -29
rect -9071 -75 -9025 -29
rect -8967 -75 -8921 -29
rect -8863 -75 -8817 -29
rect -8759 -75 -8713 -29
rect -8655 -75 -8609 -29
rect -8551 -75 -8505 -29
rect -8447 -75 -8401 -29
rect -8343 -75 -8297 -29
rect -8239 -75 -8193 -29
rect -8135 -75 -8089 -29
rect -8031 -75 -7985 -29
rect -7927 -75 -7881 -29
rect -7823 -75 -7777 -29
rect -7719 -75 -7673 -29
rect -7615 -75 -7569 -29
rect -7511 -75 -7465 -29
rect -7407 -75 -7361 -29
rect -7303 -75 -7257 -29
rect -7199 -75 -7153 -29
rect -7095 -75 -7049 -29
rect -6991 -75 -6945 -29
rect -6887 -75 -6841 -29
rect -6783 -75 -6737 -29
rect -6679 -75 -6633 -29
rect -6575 -75 -6529 -29
rect -6471 -75 -6425 -29
rect -6367 -75 -6321 -29
rect -6263 -75 -6217 -29
rect -6159 -75 -6113 -29
rect -6055 -75 -6009 -29
rect -5951 -75 -5905 -29
rect -5847 -75 -5801 -29
rect -5743 -75 -5697 -29
rect -5639 -75 -5593 -29
rect -5535 -75 -5489 -29
rect -5431 -75 -5385 -29
rect -5327 -75 -5281 -29
rect -5223 -75 -5177 -29
rect -5119 -75 -5073 -29
rect -5015 -75 -4969 -29
rect -4911 -75 -4865 -29
rect -4807 -75 -4761 -29
rect -4703 -75 -4657 -29
rect -4599 -75 -4553 -29
rect -4495 -75 -4449 -29
rect -4391 -75 -4345 -29
rect -4287 -75 -4241 -29
rect -4183 -75 -4137 -29
rect -4079 -75 -4033 -29
rect -3975 -75 -3929 -29
rect -3871 -75 -3825 -29
rect -3767 -75 -3721 -29
rect -3663 -75 -3617 -29
rect -3559 -75 -3513 -29
rect -3455 -75 -3409 -29
rect -3351 -75 -3305 -29
rect -3247 -75 -3201 -29
rect -3143 -75 -3097 -29
rect -3039 -75 -2993 -29
rect -2935 -75 -2889 -29
rect -2831 -75 -2785 -29
rect -2727 -75 -2681 -29
rect -2623 -75 -2577 -29
rect -2519 -75 -2473 -29
rect -2415 -75 -2369 -29
rect -2311 -75 -2265 -29
rect -2207 -75 -2161 -29
rect -2103 -75 -2057 -29
rect -1999 -75 -1953 -29
rect -1895 -75 -1849 -29
rect -1791 -75 -1745 -29
rect -1687 -75 -1641 -29
rect -1583 -75 -1537 -29
rect -1479 -75 -1433 -29
rect -1375 -75 -1329 -29
rect -1271 -75 -1225 -29
rect -1167 -75 -1121 -29
rect -1063 -75 -1017 -29
rect -959 -75 -913 -29
rect -855 -75 -809 -29
rect -751 -75 -705 -29
rect -647 -75 -601 -29
rect -543 -75 -497 -29
rect -439 -75 -393 -29
rect -335 -75 -289 -29
rect -231 -75 -185 -29
rect -127 -75 -81 -29
rect -23 -75 23 -29
rect 81 -75 127 -29
rect 185 -75 231 -29
rect 289 -75 335 -29
rect 393 -75 439 -29
rect 497 -75 543 -29
rect 601 -75 647 -29
rect 705 -75 751 -29
rect 809 -75 855 -29
rect 913 -75 959 -29
rect 1017 -75 1063 -29
rect 1121 -75 1167 -29
rect 1225 -75 1271 -29
rect 1329 -75 1375 -29
rect 1433 -75 1479 -29
rect 1537 -75 1583 -29
rect 1641 -75 1687 -29
rect 1745 -75 1791 -29
rect 1849 -75 1895 -29
rect 1953 -75 1999 -29
rect 2057 -75 2103 -29
rect 2161 -75 2207 -29
rect 2265 -75 2311 -29
rect 2369 -75 2415 -29
rect 2473 -75 2519 -29
rect 2577 -75 2623 -29
rect 2681 -75 2727 -29
rect 2785 -75 2831 -29
rect 2889 -75 2935 -29
rect 2993 -75 3039 -29
rect 3097 -75 3143 -29
rect 3201 -75 3247 -29
rect 3305 -75 3351 -29
rect 3409 -75 3455 -29
rect 3513 -75 3559 -29
rect 3617 -75 3663 -29
rect 3721 -75 3767 -29
rect 3825 -75 3871 -29
rect 3929 -75 3975 -29
rect 4033 -75 4079 -29
rect 4137 -75 4183 -29
rect 4241 -75 4287 -29
rect 4345 -75 4391 -29
rect 4449 -75 4495 -29
rect 4553 -75 4599 -29
rect 4657 -75 4703 -29
rect 4761 -75 4807 -29
rect 4865 -75 4911 -29
rect 4969 -75 5015 -29
rect 5073 -75 5119 -29
rect 5177 -75 5223 -29
rect 5281 -75 5327 -29
rect 5385 -75 5431 -29
rect 5489 -75 5535 -29
rect 5593 -75 5639 -29
rect 5697 -75 5743 -29
rect 5801 -75 5847 -29
rect 5905 -75 5951 -29
rect 6009 -75 6055 -29
rect 6113 -75 6159 -29
rect 6217 -75 6263 -29
rect 6321 -75 6367 -29
rect 6425 -75 6471 -29
rect 6529 -75 6575 -29
rect 6633 -75 6679 -29
rect 6737 -75 6783 -29
rect 6841 -75 6887 -29
rect 6945 -75 6991 -29
rect 7049 -75 7095 -29
rect 7153 -75 7199 -29
rect 7257 -75 7303 -29
rect 7361 -75 7407 -29
rect 7465 -75 7511 -29
rect 7569 -75 7615 -29
rect 7673 -75 7719 -29
rect 7777 -75 7823 -29
rect 7881 -75 7927 -29
rect 7985 -75 8031 -29
rect 8089 -75 8135 -29
rect 8193 -75 8239 -29
rect 8297 -75 8343 -29
rect 8401 -75 8447 -29
rect 8505 -75 8551 -29
rect 8609 -75 8655 -29
rect 8713 -75 8759 -29
rect 8817 -75 8863 -29
rect 8921 -75 8967 -29
rect 9025 -75 9071 -29
rect 9129 -75 9175 -29
rect 9233 -75 9279 -29
rect 9337 -75 9383 -29
rect 9441 -75 9487 -29
rect 9545 -75 9591 -29
rect 9649 -75 9695 -29
rect 9753 -75 9799 -29
rect 9857 -75 9903 -29
rect 9961 -75 10007 -29
rect 10065 -75 10111 -29
rect 10169 -75 10215 -29
rect 10273 -75 10319 -29
rect 10377 -75 10423 -29
rect 10481 -75 10527 -29
rect 10585 -75 10631 -29
rect 10689 -75 10735 -29
rect 10793 -75 10839 -29
rect 10897 -75 10943 -29
rect 11001 -75 11047 -29
rect 11105 -75 11151 -29
rect 11209 -75 11255 -29
rect 11313 -75 11359 -29
rect 11417 -75 11463 -29
rect 11521 -75 11567 -29
rect 11625 -75 11671 -29
rect 11729 -75 11775 -29
rect 11833 -75 11879 -29
rect 11937 -75 11983 -29
rect 12041 -75 12087 -29
rect 12145 -75 12191 -29
rect 12249 -75 12295 -29
rect 12353 -75 12399 -29
rect 12457 -75 12503 -29
rect 12561 -75 12607 -29
rect 12665 -75 12711 -29
rect 12769 -75 12815 -29
rect 12873 -75 12919 -29
<< metal1 >>
rect -12930 75 12930 86
rect -12930 29 -12919 75
rect -12873 29 -12815 75
rect -12769 29 -12711 75
rect -12665 29 -12607 75
rect -12561 29 -12503 75
rect -12457 29 -12399 75
rect -12353 29 -12295 75
rect -12249 29 -12191 75
rect -12145 29 -12087 75
rect -12041 29 -11983 75
rect -11937 29 -11879 75
rect -11833 29 -11775 75
rect -11729 29 -11671 75
rect -11625 29 -11567 75
rect -11521 29 -11463 75
rect -11417 29 -11359 75
rect -11313 29 -11255 75
rect -11209 29 -11151 75
rect -11105 29 -11047 75
rect -11001 29 -10943 75
rect -10897 29 -10839 75
rect -10793 29 -10735 75
rect -10689 29 -10631 75
rect -10585 29 -10527 75
rect -10481 29 -10423 75
rect -10377 29 -10319 75
rect -10273 29 -10215 75
rect -10169 29 -10111 75
rect -10065 29 -10007 75
rect -9961 29 -9903 75
rect -9857 29 -9799 75
rect -9753 29 -9695 75
rect -9649 29 -9591 75
rect -9545 29 -9487 75
rect -9441 29 -9383 75
rect -9337 29 -9279 75
rect -9233 29 -9175 75
rect -9129 29 -9071 75
rect -9025 29 -8967 75
rect -8921 29 -8863 75
rect -8817 29 -8759 75
rect -8713 29 -8655 75
rect -8609 29 -8551 75
rect -8505 29 -8447 75
rect -8401 29 -8343 75
rect -8297 29 -8239 75
rect -8193 29 -8135 75
rect -8089 29 -8031 75
rect -7985 29 -7927 75
rect -7881 29 -7823 75
rect -7777 29 -7719 75
rect -7673 29 -7615 75
rect -7569 29 -7511 75
rect -7465 29 -7407 75
rect -7361 29 -7303 75
rect -7257 29 -7199 75
rect -7153 29 -7095 75
rect -7049 29 -6991 75
rect -6945 29 -6887 75
rect -6841 29 -6783 75
rect -6737 29 -6679 75
rect -6633 29 -6575 75
rect -6529 29 -6471 75
rect -6425 29 -6367 75
rect -6321 29 -6263 75
rect -6217 29 -6159 75
rect -6113 29 -6055 75
rect -6009 29 -5951 75
rect -5905 29 -5847 75
rect -5801 29 -5743 75
rect -5697 29 -5639 75
rect -5593 29 -5535 75
rect -5489 29 -5431 75
rect -5385 29 -5327 75
rect -5281 29 -5223 75
rect -5177 29 -5119 75
rect -5073 29 -5015 75
rect -4969 29 -4911 75
rect -4865 29 -4807 75
rect -4761 29 -4703 75
rect -4657 29 -4599 75
rect -4553 29 -4495 75
rect -4449 29 -4391 75
rect -4345 29 -4287 75
rect -4241 29 -4183 75
rect -4137 29 -4079 75
rect -4033 29 -3975 75
rect -3929 29 -3871 75
rect -3825 29 -3767 75
rect -3721 29 -3663 75
rect -3617 29 -3559 75
rect -3513 29 -3455 75
rect -3409 29 -3351 75
rect -3305 29 -3247 75
rect -3201 29 -3143 75
rect -3097 29 -3039 75
rect -2993 29 -2935 75
rect -2889 29 -2831 75
rect -2785 29 -2727 75
rect -2681 29 -2623 75
rect -2577 29 -2519 75
rect -2473 29 -2415 75
rect -2369 29 -2311 75
rect -2265 29 -2207 75
rect -2161 29 -2103 75
rect -2057 29 -1999 75
rect -1953 29 -1895 75
rect -1849 29 -1791 75
rect -1745 29 -1687 75
rect -1641 29 -1583 75
rect -1537 29 -1479 75
rect -1433 29 -1375 75
rect -1329 29 -1271 75
rect -1225 29 -1167 75
rect -1121 29 -1063 75
rect -1017 29 -959 75
rect -913 29 -855 75
rect -809 29 -751 75
rect -705 29 -647 75
rect -601 29 -543 75
rect -497 29 -439 75
rect -393 29 -335 75
rect -289 29 -231 75
rect -185 29 -127 75
rect -81 29 -23 75
rect 23 29 81 75
rect 127 29 185 75
rect 231 29 289 75
rect 335 29 393 75
rect 439 29 497 75
rect 543 29 601 75
rect 647 29 705 75
rect 751 29 809 75
rect 855 29 913 75
rect 959 29 1017 75
rect 1063 29 1121 75
rect 1167 29 1225 75
rect 1271 29 1329 75
rect 1375 29 1433 75
rect 1479 29 1537 75
rect 1583 29 1641 75
rect 1687 29 1745 75
rect 1791 29 1849 75
rect 1895 29 1953 75
rect 1999 29 2057 75
rect 2103 29 2161 75
rect 2207 29 2265 75
rect 2311 29 2369 75
rect 2415 29 2473 75
rect 2519 29 2577 75
rect 2623 29 2681 75
rect 2727 29 2785 75
rect 2831 29 2889 75
rect 2935 29 2993 75
rect 3039 29 3097 75
rect 3143 29 3201 75
rect 3247 29 3305 75
rect 3351 29 3409 75
rect 3455 29 3513 75
rect 3559 29 3617 75
rect 3663 29 3721 75
rect 3767 29 3825 75
rect 3871 29 3929 75
rect 3975 29 4033 75
rect 4079 29 4137 75
rect 4183 29 4241 75
rect 4287 29 4345 75
rect 4391 29 4449 75
rect 4495 29 4553 75
rect 4599 29 4657 75
rect 4703 29 4761 75
rect 4807 29 4865 75
rect 4911 29 4969 75
rect 5015 29 5073 75
rect 5119 29 5177 75
rect 5223 29 5281 75
rect 5327 29 5385 75
rect 5431 29 5489 75
rect 5535 29 5593 75
rect 5639 29 5697 75
rect 5743 29 5801 75
rect 5847 29 5905 75
rect 5951 29 6009 75
rect 6055 29 6113 75
rect 6159 29 6217 75
rect 6263 29 6321 75
rect 6367 29 6425 75
rect 6471 29 6529 75
rect 6575 29 6633 75
rect 6679 29 6737 75
rect 6783 29 6841 75
rect 6887 29 6945 75
rect 6991 29 7049 75
rect 7095 29 7153 75
rect 7199 29 7257 75
rect 7303 29 7361 75
rect 7407 29 7465 75
rect 7511 29 7569 75
rect 7615 29 7673 75
rect 7719 29 7777 75
rect 7823 29 7881 75
rect 7927 29 7985 75
rect 8031 29 8089 75
rect 8135 29 8193 75
rect 8239 29 8297 75
rect 8343 29 8401 75
rect 8447 29 8505 75
rect 8551 29 8609 75
rect 8655 29 8713 75
rect 8759 29 8817 75
rect 8863 29 8921 75
rect 8967 29 9025 75
rect 9071 29 9129 75
rect 9175 29 9233 75
rect 9279 29 9337 75
rect 9383 29 9441 75
rect 9487 29 9545 75
rect 9591 29 9649 75
rect 9695 29 9753 75
rect 9799 29 9857 75
rect 9903 29 9961 75
rect 10007 29 10065 75
rect 10111 29 10169 75
rect 10215 29 10273 75
rect 10319 29 10377 75
rect 10423 29 10481 75
rect 10527 29 10585 75
rect 10631 29 10689 75
rect 10735 29 10793 75
rect 10839 29 10897 75
rect 10943 29 11001 75
rect 11047 29 11105 75
rect 11151 29 11209 75
rect 11255 29 11313 75
rect 11359 29 11417 75
rect 11463 29 11521 75
rect 11567 29 11625 75
rect 11671 29 11729 75
rect 11775 29 11833 75
rect 11879 29 11937 75
rect 11983 29 12041 75
rect 12087 29 12145 75
rect 12191 29 12249 75
rect 12295 29 12353 75
rect 12399 29 12457 75
rect 12503 29 12561 75
rect 12607 29 12665 75
rect 12711 29 12769 75
rect 12815 29 12873 75
rect 12919 29 12930 75
rect -12930 -29 12930 29
rect -12930 -75 -12919 -29
rect -12873 -75 -12815 -29
rect -12769 -75 -12711 -29
rect -12665 -75 -12607 -29
rect -12561 -75 -12503 -29
rect -12457 -75 -12399 -29
rect -12353 -75 -12295 -29
rect -12249 -75 -12191 -29
rect -12145 -75 -12087 -29
rect -12041 -75 -11983 -29
rect -11937 -75 -11879 -29
rect -11833 -75 -11775 -29
rect -11729 -75 -11671 -29
rect -11625 -75 -11567 -29
rect -11521 -75 -11463 -29
rect -11417 -75 -11359 -29
rect -11313 -75 -11255 -29
rect -11209 -75 -11151 -29
rect -11105 -75 -11047 -29
rect -11001 -75 -10943 -29
rect -10897 -75 -10839 -29
rect -10793 -75 -10735 -29
rect -10689 -75 -10631 -29
rect -10585 -75 -10527 -29
rect -10481 -75 -10423 -29
rect -10377 -75 -10319 -29
rect -10273 -75 -10215 -29
rect -10169 -75 -10111 -29
rect -10065 -75 -10007 -29
rect -9961 -75 -9903 -29
rect -9857 -75 -9799 -29
rect -9753 -75 -9695 -29
rect -9649 -75 -9591 -29
rect -9545 -75 -9487 -29
rect -9441 -75 -9383 -29
rect -9337 -75 -9279 -29
rect -9233 -75 -9175 -29
rect -9129 -75 -9071 -29
rect -9025 -75 -8967 -29
rect -8921 -75 -8863 -29
rect -8817 -75 -8759 -29
rect -8713 -75 -8655 -29
rect -8609 -75 -8551 -29
rect -8505 -75 -8447 -29
rect -8401 -75 -8343 -29
rect -8297 -75 -8239 -29
rect -8193 -75 -8135 -29
rect -8089 -75 -8031 -29
rect -7985 -75 -7927 -29
rect -7881 -75 -7823 -29
rect -7777 -75 -7719 -29
rect -7673 -75 -7615 -29
rect -7569 -75 -7511 -29
rect -7465 -75 -7407 -29
rect -7361 -75 -7303 -29
rect -7257 -75 -7199 -29
rect -7153 -75 -7095 -29
rect -7049 -75 -6991 -29
rect -6945 -75 -6887 -29
rect -6841 -75 -6783 -29
rect -6737 -75 -6679 -29
rect -6633 -75 -6575 -29
rect -6529 -75 -6471 -29
rect -6425 -75 -6367 -29
rect -6321 -75 -6263 -29
rect -6217 -75 -6159 -29
rect -6113 -75 -6055 -29
rect -6009 -75 -5951 -29
rect -5905 -75 -5847 -29
rect -5801 -75 -5743 -29
rect -5697 -75 -5639 -29
rect -5593 -75 -5535 -29
rect -5489 -75 -5431 -29
rect -5385 -75 -5327 -29
rect -5281 -75 -5223 -29
rect -5177 -75 -5119 -29
rect -5073 -75 -5015 -29
rect -4969 -75 -4911 -29
rect -4865 -75 -4807 -29
rect -4761 -75 -4703 -29
rect -4657 -75 -4599 -29
rect -4553 -75 -4495 -29
rect -4449 -75 -4391 -29
rect -4345 -75 -4287 -29
rect -4241 -75 -4183 -29
rect -4137 -75 -4079 -29
rect -4033 -75 -3975 -29
rect -3929 -75 -3871 -29
rect -3825 -75 -3767 -29
rect -3721 -75 -3663 -29
rect -3617 -75 -3559 -29
rect -3513 -75 -3455 -29
rect -3409 -75 -3351 -29
rect -3305 -75 -3247 -29
rect -3201 -75 -3143 -29
rect -3097 -75 -3039 -29
rect -2993 -75 -2935 -29
rect -2889 -75 -2831 -29
rect -2785 -75 -2727 -29
rect -2681 -75 -2623 -29
rect -2577 -75 -2519 -29
rect -2473 -75 -2415 -29
rect -2369 -75 -2311 -29
rect -2265 -75 -2207 -29
rect -2161 -75 -2103 -29
rect -2057 -75 -1999 -29
rect -1953 -75 -1895 -29
rect -1849 -75 -1791 -29
rect -1745 -75 -1687 -29
rect -1641 -75 -1583 -29
rect -1537 -75 -1479 -29
rect -1433 -75 -1375 -29
rect -1329 -75 -1271 -29
rect -1225 -75 -1167 -29
rect -1121 -75 -1063 -29
rect -1017 -75 -959 -29
rect -913 -75 -855 -29
rect -809 -75 -751 -29
rect -705 -75 -647 -29
rect -601 -75 -543 -29
rect -497 -75 -439 -29
rect -393 -75 -335 -29
rect -289 -75 -231 -29
rect -185 -75 -127 -29
rect -81 -75 -23 -29
rect 23 -75 81 -29
rect 127 -75 185 -29
rect 231 -75 289 -29
rect 335 -75 393 -29
rect 439 -75 497 -29
rect 543 -75 601 -29
rect 647 -75 705 -29
rect 751 -75 809 -29
rect 855 -75 913 -29
rect 959 -75 1017 -29
rect 1063 -75 1121 -29
rect 1167 -75 1225 -29
rect 1271 -75 1329 -29
rect 1375 -75 1433 -29
rect 1479 -75 1537 -29
rect 1583 -75 1641 -29
rect 1687 -75 1745 -29
rect 1791 -75 1849 -29
rect 1895 -75 1953 -29
rect 1999 -75 2057 -29
rect 2103 -75 2161 -29
rect 2207 -75 2265 -29
rect 2311 -75 2369 -29
rect 2415 -75 2473 -29
rect 2519 -75 2577 -29
rect 2623 -75 2681 -29
rect 2727 -75 2785 -29
rect 2831 -75 2889 -29
rect 2935 -75 2993 -29
rect 3039 -75 3097 -29
rect 3143 -75 3201 -29
rect 3247 -75 3305 -29
rect 3351 -75 3409 -29
rect 3455 -75 3513 -29
rect 3559 -75 3617 -29
rect 3663 -75 3721 -29
rect 3767 -75 3825 -29
rect 3871 -75 3929 -29
rect 3975 -75 4033 -29
rect 4079 -75 4137 -29
rect 4183 -75 4241 -29
rect 4287 -75 4345 -29
rect 4391 -75 4449 -29
rect 4495 -75 4553 -29
rect 4599 -75 4657 -29
rect 4703 -75 4761 -29
rect 4807 -75 4865 -29
rect 4911 -75 4969 -29
rect 5015 -75 5073 -29
rect 5119 -75 5177 -29
rect 5223 -75 5281 -29
rect 5327 -75 5385 -29
rect 5431 -75 5489 -29
rect 5535 -75 5593 -29
rect 5639 -75 5697 -29
rect 5743 -75 5801 -29
rect 5847 -75 5905 -29
rect 5951 -75 6009 -29
rect 6055 -75 6113 -29
rect 6159 -75 6217 -29
rect 6263 -75 6321 -29
rect 6367 -75 6425 -29
rect 6471 -75 6529 -29
rect 6575 -75 6633 -29
rect 6679 -75 6737 -29
rect 6783 -75 6841 -29
rect 6887 -75 6945 -29
rect 6991 -75 7049 -29
rect 7095 -75 7153 -29
rect 7199 -75 7257 -29
rect 7303 -75 7361 -29
rect 7407 -75 7465 -29
rect 7511 -75 7569 -29
rect 7615 -75 7673 -29
rect 7719 -75 7777 -29
rect 7823 -75 7881 -29
rect 7927 -75 7985 -29
rect 8031 -75 8089 -29
rect 8135 -75 8193 -29
rect 8239 -75 8297 -29
rect 8343 -75 8401 -29
rect 8447 -75 8505 -29
rect 8551 -75 8609 -29
rect 8655 -75 8713 -29
rect 8759 -75 8817 -29
rect 8863 -75 8921 -29
rect 8967 -75 9025 -29
rect 9071 -75 9129 -29
rect 9175 -75 9233 -29
rect 9279 -75 9337 -29
rect 9383 -75 9441 -29
rect 9487 -75 9545 -29
rect 9591 -75 9649 -29
rect 9695 -75 9753 -29
rect 9799 -75 9857 -29
rect 9903 -75 9961 -29
rect 10007 -75 10065 -29
rect 10111 -75 10169 -29
rect 10215 -75 10273 -29
rect 10319 -75 10377 -29
rect 10423 -75 10481 -29
rect 10527 -75 10585 -29
rect 10631 -75 10689 -29
rect 10735 -75 10793 -29
rect 10839 -75 10897 -29
rect 10943 -75 11001 -29
rect 11047 -75 11105 -29
rect 11151 -75 11209 -29
rect 11255 -75 11313 -29
rect 11359 -75 11417 -29
rect 11463 -75 11521 -29
rect 11567 -75 11625 -29
rect 11671 -75 11729 -29
rect 11775 -75 11833 -29
rect 11879 -75 11937 -29
rect 11983 -75 12041 -29
rect 12087 -75 12145 -29
rect 12191 -75 12249 -29
rect 12295 -75 12353 -29
rect 12399 -75 12457 -29
rect 12503 -75 12561 -29
rect 12607 -75 12665 -29
rect 12711 -75 12769 -29
rect 12815 -75 12873 -29
rect 12919 -75 12930 -29
rect -12930 -86 12930 -75
<< end >>
