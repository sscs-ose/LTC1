magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2045 -2327 2045 2327
<< ndiff >>
rect -45 305 45 327
rect -45 -305 -23 305
rect 23 -305 45 305
rect -45 -327 45 -305
<< ndiffc >>
rect -23 -305 23 305
<< metal1 >>
rect -34 305 34 316
rect -34 -305 -23 305
rect 23 -305 34 305
rect -34 -316 34 -305
<< end >>
