magic
tech gf180mcuC
magscale 1 10
timestamp 1699111554
<< nwell >>
rect -3024 -1086 3024 1086
<< nsubdiff >>
rect -3000 990 3000 1062
rect -3000 -990 -2928 990
rect 2928 -990 3000 990
rect -3000 -1062 3000 -990
<< polysilicon >>
rect -2840 889 -2440 902
rect -2840 843 -2827 889
rect -2453 843 -2440 889
rect -2840 800 -2440 843
rect -2840 -843 -2440 -800
rect -2840 -889 -2827 -843
rect -2453 -889 -2440 -843
rect -2840 -902 -2440 -889
rect -2360 889 -1960 902
rect -2360 843 -2347 889
rect -1973 843 -1960 889
rect -2360 800 -1960 843
rect -2360 -843 -1960 -800
rect -2360 -889 -2347 -843
rect -1973 -889 -1960 -843
rect -2360 -902 -1960 -889
rect -1880 889 -1480 902
rect -1880 843 -1867 889
rect -1493 843 -1480 889
rect -1880 800 -1480 843
rect -1880 -843 -1480 -800
rect -1880 -889 -1867 -843
rect -1493 -889 -1480 -843
rect -1880 -902 -1480 -889
rect -1400 889 -1000 902
rect -1400 843 -1387 889
rect -1013 843 -1000 889
rect -1400 800 -1000 843
rect -1400 -843 -1000 -800
rect -1400 -889 -1387 -843
rect -1013 -889 -1000 -843
rect -1400 -902 -1000 -889
rect -920 889 -520 902
rect -920 843 -907 889
rect -533 843 -520 889
rect -920 800 -520 843
rect -920 -843 -520 -800
rect -920 -889 -907 -843
rect -533 -889 -520 -843
rect -920 -902 -520 -889
rect -440 889 -40 902
rect -440 843 -427 889
rect -53 843 -40 889
rect -440 800 -40 843
rect -440 -843 -40 -800
rect -440 -889 -427 -843
rect -53 -889 -40 -843
rect -440 -902 -40 -889
rect 40 889 440 902
rect 40 843 53 889
rect 427 843 440 889
rect 40 800 440 843
rect 40 -843 440 -800
rect 40 -889 53 -843
rect 427 -889 440 -843
rect 40 -902 440 -889
rect 520 889 920 902
rect 520 843 533 889
rect 907 843 920 889
rect 520 800 920 843
rect 520 -843 920 -800
rect 520 -889 533 -843
rect 907 -889 920 -843
rect 520 -902 920 -889
rect 1000 889 1400 902
rect 1000 843 1013 889
rect 1387 843 1400 889
rect 1000 800 1400 843
rect 1000 -843 1400 -800
rect 1000 -889 1013 -843
rect 1387 -889 1400 -843
rect 1000 -902 1400 -889
rect 1480 889 1880 902
rect 1480 843 1493 889
rect 1867 843 1880 889
rect 1480 800 1880 843
rect 1480 -843 1880 -800
rect 1480 -889 1493 -843
rect 1867 -889 1880 -843
rect 1480 -902 1880 -889
rect 1960 889 2360 902
rect 1960 843 1973 889
rect 2347 843 2360 889
rect 1960 800 2360 843
rect 1960 -843 2360 -800
rect 1960 -889 1973 -843
rect 2347 -889 2360 -843
rect 1960 -902 2360 -889
rect 2440 889 2840 902
rect 2440 843 2453 889
rect 2827 843 2840 889
rect 2440 800 2840 843
rect 2440 -843 2840 -800
rect 2440 -889 2453 -843
rect 2827 -889 2840 -843
rect 2440 -902 2840 -889
<< polycontact >>
rect -2827 843 -2453 889
rect -2827 -889 -2453 -843
rect -2347 843 -1973 889
rect -2347 -889 -1973 -843
rect -1867 843 -1493 889
rect -1867 -889 -1493 -843
rect -1387 843 -1013 889
rect -1387 -889 -1013 -843
rect -907 843 -533 889
rect -907 -889 -533 -843
rect -427 843 -53 889
rect -427 -889 -53 -843
rect 53 843 427 889
rect 53 -889 427 -843
rect 533 843 907 889
rect 533 -889 907 -843
rect 1013 843 1387 889
rect 1013 -889 1387 -843
rect 1493 843 1867 889
rect 1493 -889 1867 -843
rect 1973 843 2347 889
rect 1973 -889 2347 -843
rect 2453 843 2827 889
rect 2453 -889 2827 -843
<< ppolyres >>
rect -2840 -800 -2440 800
rect -2360 -800 -1960 800
rect -1880 -800 -1480 800
rect -1400 -800 -1000 800
rect -920 -800 -520 800
rect -440 -800 -40 800
rect 40 -800 440 800
rect 520 -800 920 800
rect 1000 -800 1400 800
rect 1480 -800 1880 800
rect 1960 -800 2360 800
rect 2440 -800 2840 800
<< metal1 >>
rect -2838 843 -2827 889
rect -2453 843 -2442 889
rect -2358 843 -2347 889
rect -1973 843 -1962 889
rect -1878 843 -1867 889
rect -1493 843 -1482 889
rect -1398 843 -1387 889
rect -1013 843 -1002 889
rect -918 843 -907 889
rect -533 843 -522 889
rect -438 843 -427 889
rect -53 843 -42 889
rect 42 843 53 889
rect 427 843 438 889
rect 522 843 533 889
rect 907 843 918 889
rect 1002 843 1013 889
rect 1387 843 1398 889
rect 1482 843 1493 889
rect 1867 843 1878 889
rect 1962 843 1973 889
rect 2347 843 2358 889
rect 2442 843 2453 889
rect 2827 843 2838 889
rect -2838 -889 -2827 -843
rect -2453 -889 -2442 -843
rect -2358 -889 -2347 -843
rect -1973 -889 -1962 -843
rect -1878 -889 -1867 -843
rect -1493 -889 -1482 -843
rect -1398 -889 -1387 -843
rect -1013 -889 -1002 -843
rect -918 -889 -907 -843
rect -533 -889 -522 -843
rect -438 -889 -427 -843
rect -53 -889 -42 -843
rect 42 -889 53 -843
rect 427 -889 438 -843
rect 522 -889 533 -843
rect 907 -889 918 -843
rect 1002 -889 1013 -843
rect 1387 -889 1398 -843
rect 1482 -889 1493 -843
rect 1867 -889 1878 -843
rect 1962 -889 1973 -843
rect 2347 -889 2358 -843
rect 2442 -889 2453 -843
rect 2827 -889 2838 -843
<< properties >>
string FIXED_BBOX -2964 -1026 2964 1026
string gencell ppolyf_u
string library gf180mcu
string parameters w 2.0 l 8.0 m 1 nx 12 wmin 0.80 lmin 1.00 rho 315 val 1.305k dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 0 grc 0 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 0
<< end >>
