magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1298 -1019 1298 1019
<< metal1 >>
rect -298 13 298 19
rect -298 -13 -292 13
rect -266 -13 -230 13
rect -204 -13 -168 13
rect -142 -13 -106 13
rect -80 -13 -44 13
rect -18 -13 18 13
rect 44 -13 80 13
rect 106 -13 142 13
rect 168 -13 204 13
rect 230 -13 266 13
rect 292 -13 298 13
rect -298 -19 298 -13
<< via1 >>
rect -292 -13 -266 13
rect -230 -13 -204 13
rect -168 -13 -142 13
rect -106 -13 -80 13
rect -44 -13 -18 13
rect 18 -13 44 13
rect 80 -13 106 13
rect 142 -13 168 13
rect 204 -13 230 13
rect 266 -13 292 13
<< metal2 >>
rect -298 13 298 19
rect -298 -13 -292 13
rect -266 -13 -230 13
rect -204 -13 -168 13
rect -142 -13 -106 13
rect -80 -13 -44 13
rect -18 -13 18 13
rect 44 -13 80 13
rect 106 -13 142 13
rect 168 -13 204 13
rect 230 -13 266 13
rect 292 -13 298 13
rect -298 -19 298 -13
<< end >>
