magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -1979 -2485 3081 2648
<< nwell >>
rect 21 513 1081 648
rect 21 507 166 513
rect 168 507 525 508
rect 528 507 1081 513
rect 371 470 907 483
rect 321 180 324 242
<< psubdiff >>
rect 38 -385 1061 -372
rect 38 -431 51 -385
rect 1037 -431 1061 -385
rect 38 -444 1061 -431
<< nsubdiff >>
rect 47 604 1002 617
rect 47 558 66 604
rect 958 558 1002 604
rect 47 545 1002 558
<< psubdiffcont >>
rect 51 -431 1037 -385
<< nsubdiffcont >>
rect 66 558 958 604
<< polysilicon >>
rect 195 417 907 483
rect 195 180 907 242
rect 194 -40 295 9
rect 194 -86 208 -40
rect 254 -83 295 -40
rect 399 -83 499 3
rect 603 -83 703 3
rect 807 -83 907 3
rect 254 -86 907 -83
rect 194 -131 907 -86
<< polycontact >>
rect 208 -86 254 -40
<< metal1 >>
rect 21 604 1081 648
rect 21 558 66 604
rect 958 558 1081 604
rect 21 525 1081 558
rect 21 524 574 525
rect 40 381 106 524
rect 40 295 166 381
rect 120 135 166 295
rect 324 141 370 381
rect 528 372 574 524
rect 936 372 982 525
rect 528 140 574 302
rect 732 142 778 290
rect 936 134 982 298
rect 324 2 370 53
rect 732 2 778 50
rect 35 -40 266 -27
rect 35 -86 208 -40
rect 254 -86 266 -40
rect 35 -99 266 -86
rect 324 -44 1071 2
rect 324 -189 370 -44
rect 732 -182 778 -44
rect 120 -342 166 -256
rect 528 -342 574 -253
rect 936 -342 982 -252
rect 22 -385 1080 -342
rect 22 -431 51 -385
rect 1037 -431 1080 -385
rect 22 -485 1080 -431
use nmos_3p3_6FEA4B  nmos_3p3_6FEA4B_0
timestamp 1713185578
transform 1 0 551 0 1 -225
box -468 -118 468 118
use pmos_3p3_KYEELV  pmos_3p3_KYEELV_0
timestamp 1713185578
transform 1 0 551 0 1 215
box -530 -298 530 298
<< labels >>
flabel nsubdiffcont 559 581 559 581 0 FreeSans 1250 0 0 0 VDD
flabel psubdiffcont 544 -408 544 -408 0 FreeSans 1250 0 0 0 VSS
flabel metal1 s 53 -64 53 -64 0 FreeSans 1250 0 0 0 IN
port 1 nsew
flabel metal1 s 1042 -23 1042 -23 0 FreeSans 1250 0 0 0 OUT
port 2 nsew
<< end >>
