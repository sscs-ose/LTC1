magic
tech gf180mcuC
magscale 1 10
timestamp 1692949102
<< error_p >>
rect -3352 -3116 -3074 -3084
rect -3282 -3140 -3206 -3116
rect -1306 -3140 -1230 -3116
rect -3306 -3164 -3182 -3140
rect -1330 -3164 -1206 -3140
<< nwell >>
rect -3327 -3140 -1192 -2523
rect -3130 -3190 -1330 -3140
<< nsubdiff >>
rect -3282 -2593 -1230 -2578
rect -3282 -2640 -3267 -2593
rect -3220 -2639 -3172 -2593
rect -3126 -2639 -3078 -2593
rect -3032 -2639 -2984 -2593
rect -2938 -2639 -2890 -2593
rect -2844 -2639 -2796 -2593
rect -2750 -2639 -2702 -2593
rect -2656 -2639 -2608 -2593
rect -2562 -2639 -2514 -2593
rect -2468 -2639 -2420 -2593
rect -2374 -2639 -2326 -2593
rect -2280 -2639 -2232 -2593
rect -2186 -2639 -2138 -2593
rect -2092 -2639 -2044 -2593
rect -1998 -2639 -1950 -2593
rect -1904 -2639 -1856 -2593
rect -1810 -2639 -1762 -2593
rect -1716 -2639 -1668 -2593
rect -1622 -2639 -1574 -2593
rect -1528 -2639 -1480 -2593
rect -1434 -2639 -1386 -2593
rect -1340 -2639 -1292 -2593
rect -3220 -2640 -1292 -2639
rect -1245 -2640 -1230 -2593
rect -3282 -2654 -1230 -2640
rect -3282 -2688 -3206 -2654
rect -3282 -2734 -3267 -2688
rect -3221 -2734 -3206 -2688
rect -1306 -2688 -1230 -2654
rect -3282 -2782 -3206 -2734
rect -3282 -2828 -3267 -2782
rect -3221 -2828 -3206 -2782
rect -3282 -2876 -3206 -2828
rect -1306 -2734 -1291 -2688
rect -1245 -2734 -1230 -2688
rect -1306 -2782 -1230 -2734
rect -1306 -2828 -1291 -2782
rect -1245 -2828 -1230 -2782
rect -3282 -2922 -3267 -2876
rect -3221 -2922 -3206 -2876
rect -3282 -2970 -3206 -2922
rect -3282 -3016 -3267 -2970
rect -3221 -3016 -3206 -2970
rect -3282 -3064 -3206 -3016
rect -3282 -3110 -3267 -3064
rect -3221 -3110 -3206 -3064
rect -3282 -3140 -3206 -3110
rect -1306 -2876 -1230 -2828
rect -1306 -2922 -1291 -2876
rect -1245 -2922 -1230 -2876
rect -1306 -2970 -1230 -2922
rect -1306 -3016 -1291 -2970
rect -1245 -3016 -1230 -2970
rect -1306 -3064 -1230 -3016
rect -1306 -3110 -1291 -3064
rect -1245 -3110 -1230 -3064
rect -1306 -3140 -1230 -3110
<< nsubdiffcont >>
rect -3267 -2640 -3220 -2593
rect -3172 -2639 -3126 -2593
rect -3078 -2639 -3032 -2593
rect -2984 -2639 -2938 -2593
rect -2890 -2639 -2844 -2593
rect -2796 -2639 -2750 -2593
rect -2702 -2639 -2656 -2593
rect -2608 -2639 -2562 -2593
rect -2514 -2639 -2468 -2593
rect -2420 -2639 -2374 -2593
rect -2326 -2639 -2280 -2593
rect -2232 -2639 -2186 -2593
rect -2138 -2639 -2092 -2593
rect -2044 -2639 -1998 -2593
rect -1950 -2639 -1904 -2593
rect -1856 -2639 -1810 -2593
rect -1762 -2639 -1716 -2593
rect -1668 -2639 -1622 -2593
rect -1574 -2639 -1528 -2593
rect -1480 -2639 -1434 -2593
rect -1386 -2639 -1340 -2593
rect -1292 -2640 -1245 -2593
rect -3267 -2734 -3221 -2688
rect -3267 -2828 -3221 -2782
rect -1291 -2734 -1245 -2688
rect -1291 -2828 -1245 -2782
rect -3267 -2922 -3221 -2876
rect -3267 -3016 -3221 -2970
rect -3267 -3110 -3221 -3064
rect -1291 -2922 -1245 -2876
rect -1291 -3016 -1245 -2970
rect -1291 -3110 -1245 -3064
<< polysilicon >>
rect -2849 -2747 -2762 -2733
rect -2849 -2793 -2828 -2747
rect -2782 -2793 -2762 -2747
rect -2849 -2813 -2762 -2793
rect -2370 -2747 -2283 -2731
rect -2370 -2793 -2348 -2747
rect -2302 -2793 -2283 -2747
rect -2370 -2811 -2283 -2793
rect -2207 -2747 -2120 -2731
rect -2207 -2793 -2188 -2747
rect -2142 -2793 -2120 -2747
rect -2207 -2811 -2120 -2793
rect -1728 -2747 -1642 -2733
rect -1728 -2793 -1708 -2747
rect -1662 -2793 -1642 -2747
rect -2833 -2865 -2777 -2813
rect -2353 -2821 -2297 -2811
rect -2193 -2821 -2137 -2811
rect -1728 -2813 -1642 -2793
rect -1713 -2865 -1657 -2813
<< polycontact >>
rect -2828 -2793 -2782 -2747
rect -2348 -2793 -2302 -2747
rect -2188 -2793 -2142 -2747
rect -1708 -2793 -1662 -2747
<< metal1 >>
rect -1536 -2567 -1372 -2500
rect -3293 -2593 -1219 -2567
rect -3293 -2640 -3267 -2593
rect -3220 -2639 -3172 -2593
rect -3126 -2639 -3078 -2593
rect -3032 -2639 -2984 -2593
rect -2938 -2639 -2890 -2593
rect -2844 -2639 -2796 -2593
rect -2750 -2639 -2702 -2593
rect -2656 -2639 -2608 -2593
rect -2562 -2639 -2514 -2593
rect -2468 -2639 -2420 -2593
rect -2374 -2639 -2326 -2593
rect -2280 -2639 -2232 -2593
rect -2186 -2639 -2138 -2593
rect -2092 -2639 -2044 -2593
rect -1998 -2639 -1950 -2593
rect -1904 -2639 -1856 -2593
rect -1810 -2639 -1762 -2593
rect -1716 -2639 -1668 -2593
rect -1622 -2639 -1574 -2593
rect -1528 -2639 -1480 -2593
rect -1434 -2639 -1386 -2593
rect -1340 -2639 -1292 -2593
rect -3220 -2640 -1292 -2639
rect -1245 -2640 -1219 -2593
rect -3293 -2654 -1219 -2640
rect -3293 -2665 -1120 -2654
rect -3293 -2688 -3195 -2665
rect -3293 -2734 -3267 -2688
rect -3221 -2734 -3195 -2688
rect -1317 -2688 -1120 -2665
rect -3293 -2782 -3195 -2734
rect -1743 -2743 -1642 -2723
rect -3293 -2828 -3267 -2782
rect -3221 -2828 -3195 -2782
rect -2849 -2744 -1642 -2743
rect -2849 -2747 -1722 -2744
rect -1666 -2747 -1642 -2744
rect -2849 -2793 -2828 -2747
rect -2782 -2793 -2348 -2747
rect -2302 -2793 -2188 -2747
rect -2142 -2793 -1722 -2747
rect -1662 -2793 -1642 -2747
rect -2849 -2799 -1722 -2793
rect -1743 -2800 -1722 -2799
rect -1666 -2800 -1642 -2793
rect -1743 -2820 -1642 -2800
rect -1317 -2734 -1291 -2688
rect -1245 -2734 -1120 -2688
rect -1317 -2782 -1120 -2734
rect -3293 -2876 -3195 -2828
rect -3293 -2922 -3267 -2876
rect -3221 -2922 -3195 -2876
rect -3293 -2970 -3195 -2922
rect -1317 -2828 -1291 -2782
rect -1245 -2793 -1120 -2782
rect -1245 -2828 -1219 -2793
rect -1317 -2876 -1219 -2828
rect -1317 -2922 -1291 -2876
rect -1245 -2922 -1219 -2876
rect -3293 -3016 -3267 -2970
rect -3221 -3016 -3195 -2970
rect -3293 -3064 -3195 -3016
rect -2607 -2967 -2524 -2953
rect -2607 -3023 -2593 -2967
rect -2537 -3023 -2524 -2967
rect -2607 -3035 -2524 -3023
rect -1965 -2967 -1882 -2952
rect -1965 -3023 -1952 -2967
rect -1896 -3023 -1882 -2967
rect -1965 -3036 -1882 -3023
rect -1317 -2970 -1219 -2922
rect -1317 -3016 -1291 -2970
rect -1245 -3016 -1219 -2970
rect -3293 -3110 -3267 -3064
rect -3221 -3110 -3195 -3064
rect -1317 -3064 -1219 -3016
rect -3293 -3140 -3195 -3110
rect -2766 -3119 -2683 -3105
rect -2766 -3175 -2752 -3119
rect -2696 -3175 -2683 -3119
rect -2766 -3187 -2683 -3175
rect -2447 -3118 -2364 -3104
rect -2447 -3174 -2433 -3118
rect -2377 -3174 -2364 -3118
rect -2447 -3186 -2364 -3174
rect -2125 -3118 -2042 -3104
rect -2125 -3174 -2111 -3118
rect -2055 -3174 -2042 -3118
rect -2125 -3186 -2042 -3174
rect -1810 -3118 -1727 -3104
rect -1810 -3174 -1796 -3118
rect -1740 -3174 -1727 -3118
rect -1317 -3110 -1291 -3064
rect -1245 -3110 -1219 -3064
rect -1317 -3140 -1219 -3110
rect -1810 -3186 -1727 -3174
<< via1 >>
rect -1722 -2747 -1666 -2744
rect -1722 -2793 -1708 -2747
rect -1708 -2793 -1666 -2747
rect -1722 -2800 -1666 -2793
rect -2593 -3023 -2537 -2967
rect -1952 -3023 -1896 -2967
rect -2752 -3175 -2696 -3119
rect -2433 -3174 -2377 -3118
rect -2111 -3174 -2055 -3118
rect -1796 -3174 -1740 -3118
<< metal2 >>
rect -3472 -3116 -3352 -2500
rect -1743 -2744 -1642 -2723
rect -1743 -2800 -1722 -2744
rect -1666 -2800 -1642 -2744
rect -1743 -2820 -1642 -2800
rect -2607 -2965 -2524 -2953
rect -2156 -2965 -1882 -2952
rect -2607 -2967 -2142 -2965
rect -2607 -3023 -2593 -2967
rect -2537 -3021 -2142 -2967
rect -2086 -3021 -2032 -2965
rect -1976 -2967 -1882 -2965
rect -1976 -3021 -1952 -2967
rect -2537 -3023 -1952 -3021
rect -1896 -3023 -1882 -2967
rect -2607 -3025 -1882 -3023
rect -2607 -3035 -2524 -3025
rect -2156 -3036 -1882 -3025
rect -2766 -3116 -2683 -3105
rect -2447 -3116 -2364 -3104
rect -2125 -3116 -2042 -3104
rect -1810 -3116 -1727 -3104
rect -3472 -3118 -1727 -3116
rect -3472 -3119 -2433 -3118
rect -3472 -3140 -2752 -3119
rect -3472 -3177 -3350 -3140
rect -3130 -3175 -2752 -3140
rect -2696 -3174 -2433 -3119
rect -2377 -3174 -2111 -3118
rect -2055 -3174 -1796 -3118
rect -1740 -3174 -1727 -3118
rect -2696 -3175 -1727 -3174
rect -3130 -3177 -1727 -3175
rect -3472 -3190 -3352 -3177
rect -2766 -3187 -2683 -3177
rect -2447 -3186 -2364 -3177
rect -2125 -3186 -2042 -3177
rect -1810 -3186 -1727 -3177
<< via2 >>
rect -1722 -2800 -1666 -2744
rect -2142 -3021 -2086 -2965
rect -2032 -3021 -1976 -2965
<< metal3 >>
rect -3500 -2572 -1660 -2506
rect -1726 -2723 -1660 -2572
rect -3500 -2804 -2767 -2738
rect -2833 -3190 -2767 -2804
rect -1743 -2744 -1642 -2723
rect -1743 -2800 -1722 -2744
rect -1666 -2800 -1642 -2744
rect -1743 -2820 -1642 -2800
rect -2156 -2965 -1964 -2952
rect -2156 -3021 -2142 -2965
rect -2086 -3021 -2032 -2965
rect -1976 -3021 -1964 -2965
rect -2156 -3036 -1964 -3021
rect -2097 -3190 -2031 -3036
rect -1726 -3190 -1660 -2820
<< end >>
