magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -9351 -2677 9351 2677
<< metal3 >>
rect -7351 667 7351 677
rect -7351 611 -7341 667
rect -7285 611 -7199 667
rect -7143 611 -7057 667
rect -7001 611 -6915 667
rect -6859 611 -6773 667
rect -6717 611 -6631 667
rect -6575 611 -6489 667
rect -6433 611 -6347 667
rect -6291 611 -6205 667
rect -6149 611 -6063 667
rect -6007 611 -5921 667
rect -5865 611 -5779 667
rect -5723 611 -5637 667
rect -5581 611 -5495 667
rect -5439 611 -5353 667
rect -5297 611 -5211 667
rect -5155 611 -5069 667
rect -5013 611 -4927 667
rect -4871 611 -4785 667
rect -4729 611 -4643 667
rect -4587 611 -4501 667
rect -4445 611 -4359 667
rect -4303 611 -4217 667
rect -4161 611 -4075 667
rect -4019 611 -3933 667
rect -3877 611 -3791 667
rect -3735 611 -3649 667
rect -3593 611 -3507 667
rect -3451 611 -3365 667
rect -3309 611 -3223 667
rect -3167 611 -3081 667
rect -3025 611 -2939 667
rect -2883 611 -2797 667
rect -2741 611 -2655 667
rect -2599 611 -2513 667
rect -2457 611 -2371 667
rect -2315 611 -2229 667
rect -2173 611 -2087 667
rect -2031 611 -1945 667
rect -1889 611 -1803 667
rect -1747 611 -1661 667
rect -1605 611 -1519 667
rect -1463 611 -1377 667
rect -1321 611 -1235 667
rect -1179 611 -1093 667
rect -1037 611 -951 667
rect -895 611 -809 667
rect -753 611 -667 667
rect -611 611 -525 667
rect -469 611 -383 667
rect -327 611 -241 667
rect -185 611 -99 667
rect -43 611 43 667
rect 99 611 185 667
rect 241 611 327 667
rect 383 611 469 667
rect 525 611 611 667
rect 667 611 753 667
rect 809 611 895 667
rect 951 611 1037 667
rect 1093 611 1179 667
rect 1235 611 1321 667
rect 1377 611 1463 667
rect 1519 611 1605 667
rect 1661 611 1747 667
rect 1803 611 1889 667
rect 1945 611 2031 667
rect 2087 611 2173 667
rect 2229 611 2315 667
rect 2371 611 2457 667
rect 2513 611 2599 667
rect 2655 611 2741 667
rect 2797 611 2883 667
rect 2939 611 3025 667
rect 3081 611 3167 667
rect 3223 611 3309 667
rect 3365 611 3451 667
rect 3507 611 3593 667
rect 3649 611 3735 667
rect 3791 611 3877 667
rect 3933 611 4019 667
rect 4075 611 4161 667
rect 4217 611 4303 667
rect 4359 611 4445 667
rect 4501 611 4587 667
rect 4643 611 4729 667
rect 4785 611 4871 667
rect 4927 611 5013 667
rect 5069 611 5155 667
rect 5211 611 5297 667
rect 5353 611 5439 667
rect 5495 611 5581 667
rect 5637 611 5723 667
rect 5779 611 5865 667
rect 5921 611 6007 667
rect 6063 611 6149 667
rect 6205 611 6291 667
rect 6347 611 6433 667
rect 6489 611 6575 667
rect 6631 611 6717 667
rect 6773 611 6859 667
rect 6915 611 7001 667
rect 7057 611 7143 667
rect 7199 611 7285 667
rect 7341 611 7351 667
rect -7351 525 7351 611
rect -7351 469 -7341 525
rect -7285 469 -7199 525
rect -7143 469 -7057 525
rect -7001 469 -6915 525
rect -6859 469 -6773 525
rect -6717 469 -6631 525
rect -6575 469 -6489 525
rect -6433 469 -6347 525
rect -6291 469 -6205 525
rect -6149 469 -6063 525
rect -6007 469 -5921 525
rect -5865 469 -5779 525
rect -5723 469 -5637 525
rect -5581 469 -5495 525
rect -5439 469 -5353 525
rect -5297 469 -5211 525
rect -5155 469 -5069 525
rect -5013 469 -4927 525
rect -4871 469 -4785 525
rect -4729 469 -4643 525
rect -4587 469 -4501 525
rect -4445 469 -4359 525
rect -4303 469 -4217 525
rect -4161 469 -4075 525
rect -4019 469 -3933 525
rect -3877 469 -3791 525
rect -3735 469 -3649 525
rect -3593 469 -3507 525
rect -3451 469 -3365 525
rect -3309 469 -3223 525
rect -3167 469 -3081 525
rect -3025 469 -2939 525
rect -2883 469 -2797 525
rect -2741 469 -2655 525
rect -2599 469 -2513 525
rect -2457 469 -2371 525
rect -2315 469 -2229 525
rect -2173 469 -2087 525
rect -2031 469 -1945 525
rect -1889 469 -1803 525
rect -1747 469 -1661 525
rect -1605 469 -1519 525
rect -1463 469 -1377 525
rect -1321 469 -1235 525
rect -1179 469 -1093 525
rect -1037 469 -951 525
rect -895 469 -809 525
rect -753 469 -667 525
rect -611 469 -525 525
rect -469 469 -383 525
rect -327 469 -241 525
rect -185 469 -99 525
rect -43 469 43 525
rect 99 469 185 525
rect 241 469 327 525
rect 383 469 469 525
rect 525 469 611 525
rect 667 469 753 525
rect 809 469 895 525
rect 951 469 1037 525
rect 1093 469 1179 525
rect 1235 469 1321 525
rect 1377 469 1463 525
rect 1519 469 1605 525
rect 1661 469 1747 525
rect 1803 469 1889 525
rect 1945 469 2031 525
rect 2087 469 2173 525
rect 2229 469 2315 525
rect 2371 469 2457 525
rect 2513 469 2599 525
rect 2655 469 2741 525
rect 2797 469 2883 525
rect 2939 469 3025 525
rect 3081 469 3167 525
rect 3223 469 3309 525
rect 3365 469 3451 525
rect 3507 469 3593 525
rect 3649 469 3735 525
rect 3791 469 3877 525
rect 3933 469 4019 525
rect 4075 469 4161 525
rect 4217 469 4303 525
rect 4359 469 4445 525
rect 4501 469 4587 525
rect 4643 469 4729 525
rect 4785 469 4871 525
rect 4927 469 5013 525
rect 5069 469 5155 525
rect 5211 469 5297 525
rect 5353 469 5439 525
rect 5495 469 5581 525
rect 5637 469 5723 525
rect 5779 469 5865 525
rect 5921 469 6007 525
rect 6063 469 6149 525
rect 6205 469 6291 525
rect 6347 469 6433 525
rect 6489 469 6575 525
rect 6631 469 6717 525
rect 6773 469 6859 525
rect 6915 469 7001 525
rect 7057 469 7143 525
rect 7199 469 7285 525
rect 7341 469 7351 525
rect -7351 383 7351 469
rect -7351 327 -7341 383
rect -7285 327 -7199 383
rect -7143 327 -7057 383
rect -7001 327 -6915 383
rect -6859 327 -6773 383
rect -6717 327 -6631 383
rect -6575 327 -6489 383
rect -6433 327 -6347 383
rect -6291 327 -6205 383
rect -6149 327 -6063 383
rect -6007 327 -5921 383
rect -5865 327 -5779 383
rect -5723 327 -5637 383
rect -5581 327 -5495 383
rect -5439 327 -5353 383
rect -5297 327 -5211 383
rect -5155 327 -5069 383
rect -5013 327 -4927 383
rect -4871 327 -4785 383
rect -4729 327 -4643 383
rect -4587 327 -4501 383
rect -4445 327 -4359 383
rect -4303 327 -4217 383
rect -4161 327 -4075 383
rect -4019 327 -3933 383
rect -3877 327 -3791 383
rect -3735 327 -3649 383
rect -3593 327 -3507 383
rect -3451 327 -3365 383
rect -3309 327 -3223 383
rect -3167 327 -3081 383
rect -3025 327 -2939 383
rect -2883 327 -2797 383
rect -2741 327 -2655 383
rect -2599 327 -2513 383
rect -2457 327 -2371 383
rect -2315 327 -2229 383
rect -2173 327 -2087 383
rect -2031 327 -1945 383
rect -1889 327 -1803 383
rect -1747 327 -1661 383
rect -1605 327 -1519 383
rect -1463 327 -1377 383
rect -1321 327 -1235 383
rect -1179 327 -1093 383
rect -1037 327 -951 383
rect -895 327 -809 383
rect -753 327 -667 383
rect -611 327 -525 383
rect -469 327 -383 383
rect -327 327 -241 383
rect -185 327 -99 383
rect -43 327 43 383
rect 99 327 185 383
rect 241 327 327 383
rect 383 327 469 383
rect 525 327 611 383
rect 667 327 753 383
rect 809 327 895 383
rect 951 327 1037 383
rect 1093 327 1179 383
rect 1235 327 1321 383
rect 1377 327 1463 383
rect 1519 327 1605 383
rect 1661 327 1747 383
rect 1803 327 1889 383
rect 1945 327 2031 383
rect 2087 327 2173 383
rect 2229 327 2315 383
rect 2371 327 2457 383
rect 2513 327 2599 383
rect 2655 327 2741 383
rect 2797 327 2883 383
rect 2939 327 3025 383
rect 3081 327 3167 383
rect 3223 327 3309 383
rect 3365 327 3451 383
rect 3507 327 3593 383
rect 3649 327 3735 383
rect 3791 327 3877 383
rect 3933 327 4019 383
rect 4075 327 4161 383
rect 4217 327 4303 383
rect 4359 327 4445 383
rect 4501 327 4587 383
rect 4643 327 4729 383
rect 4785 327 4871 383
rect 4927 327 5013 383
rect 5069 327 5155 383
rect 5211 327 5297 383
rect 5353 327 5439 383
rect 5495 327 5581 383
rect 5637 327 5723 383
rect 5779 327 5865 383
rect 5921 327 6007 383
rect 6063 327 6149 383
rect 6205 327 6291 383
rect 6347 327 6433 383
rect 6489 327 6575 383
rect 6631 327 6717 383
rect 6773 327 6859 383
rect 6915 327 7001 383
rect 7057 327 7143 383
rect 7199 327 7285 383
rect 7341 327 7351 383
rect -7351 241 7351 327
rect -7351 185 -7341 241
rect -7285 185 -7199 241
rect -7143 185 -7057 241
rect -7001 185 -6915 241
rect -6859 185 -6773 241
rect -6717 185 -6631 241
rect -6575 185 -6489 241
rect -6433 185 -6347 241
rect -6291 185 -6205 241
rect -6149 185 -6063 241
rect -6007 185 -5921 241
rect -5865 185 -5779 241
rect -5723 185 -5637 241
rect -5581 185 -5495 241
rect -5439 185 -5353 241
rect -5297 185 -5211 241
rect -5155 185 -5069 241
rect -5013 185 -4927 241
rect -4871 185 -4785 241
rect -4729 185 -4643 241
rect -4587 185 -4501 241
rect -4445 185 -4359 241
rect -4303 185 -4217 241
rect -4161 185 -4075 241
rect -4019 185 -3933 241
rect -3877 185 -3791 241
rect -3735 185 -3649 241
rect -3593 185 -3507 241
rect -3451 185 -3365 241
rect -3309 185 -3223 241
rect -3167 185 -3081 241
rect -3025 185 -2939 241
rect -2883 185 -2797 241
rect -2741 185 -2655 241
rect -2599 185 -2513 241
rect -2457 185 -2371 241
rect -2315 185 -2229 241
rect -2173 185 -2087 241
rect -2031 185 -1945 241
rect -1889 185 -1803 241
rect -1747 185 -1661 241
rect -1605 185 -1519 241
rect -1463 185 -1377 241
rect -1321 185 -1235 241
rect -1179 185 -1093 241
rect -1037 185 -951 241
rect -895 185 -809 241
rect -753 185 -667 241
rect -611 185 -525 241
rect -469 185 -383 241
rect -327 185 -241 241
rect -185 185 -99 241
rect -43 185 43 241
rect 99 185 185 241
rect 241 185 327 241
rect 383 185 469 241
rect 525 185 611 241
rect 667 185 753 241
rect 809 185 895 241
rect 951 185 1037 241
rect 1093 185 1179 241
rect 1235 185 1321 241
rect 1377 185 1463 241
rect 1519 185 1605 241
rect 1661 185 1747 241
rect 1803 185 1889 241
rect 1945 185 2031 241
rect 2087 185 2173 241
rect 2229 185 2315 241
rect 2371 185 2457 241
rect 2513 185 2599 241
rect 2655 185 2741 241
rect 2797 185 2883 241
rect 2939 185 3025 241
rect 3081 185 3167 241
rect 3223 185 3309 241
rect 3365 185 3451 241
rect 3507 185 3593 241
rect 3649 185 3735 241
rect 3791 185 3877 241
rect 3933 185 4019 241
rect 4075 185 4161 241
rect 4217 185 4303 241
rect 4359 185 4445 241
rect 4501 185 4587 241
rect 4643 185 4729 241
rect 4785 185 4871 241
rect 4927 185 5013 241
rect 5069 185 5155 241
rect 5211 185 5297 241
rect 5353 185 5439 241
rect 5495 185 5581 241
rect 5637 185 5723 241
rect 5779 185 5865 241
rect 5921 185 6007 241
rect 6063 185 6149 241
rect 6205 185 6291 241
rect 6347 185 6433 241
rect 6489 185 6575 241
rect 6631 185 6717 241
rect 6773 185 6859 241
rect 6915 185 7001 241
rect 7057 185 7143 241
rect 7199 185 7285 241
rect 7341 185 7351 241
rect -7351 99 7351 185
rect -7351 43 -7341 99
rect -7285 43 -7199 99
rect -7143 43 -7057 99
rect -7001 43 -6915 99
rect -6859 43 -6773 99
rect -6717 43 -6631 99
rect -6575 43 -6489 99
rect -6433 43 -6347 99
rect -6291 43 -6205 99
rect -6149 43 -6063 99
rect -6007 43 -5921 99
rect -5865 43 -5779 99
rect -5723 43 -5637 99
rect -5581 43 -5495 99
rect -5439 43 -5353 99
rect -5297 43 -5211 99
rect -5155 43 -5069 99
rect -5013 43 -4927 99
rect -4871 43 -4785 99
rect -4729 43 -4643 99
rect -4587 43 -4501 99
rect -4445 43 -4359 99
rect -4303 43 -4217 99
rect -4161 43 -4075 99
rect -4019 43 -3933 99
rect -3877 43 -3791 99
rect -3735 43 -3649 99
rect -3593 43 -3507 99
rect -3451 43 -3365 99
rect -3309 43 -3223 99
rect -3167 43 -3081 99
rect -3025 43 -2939 99
rect -2883 43 -2797 99
rect -2741 43 -2655 99
rect -2599 43 -2513 99
rect -2457 43 -2371 99
rect -2315 43 -2229 99
rect -2173 43 -2087 99
rect -2031 43 -1945 99
rect -1889 43 -1803 99
rect -1747 43 -1661 99
rect -1605 43 -1519 99
rect -1463 43 -1377 99
rect -1321 43 -1235 99
rect -1179 43 -1093 99
rect -1037 43 -951 99
rect -895 43 -809 99
rect -753 43 -667 99
rect -611 43 -525 99
rect -469 43 -383 99
rect -327 43 -241 99
rect -185 43 -99 99
rect -43 43 43 99
rect 99 43 185 99
rect 241 43 327 99
rect 383 43 469 99
rect 525 43 611 99
rect 667 43 753 99
rect 809 43 895 99
rect 951 43 1037 99
rect 1093 43 1179 99
rect 1235 43 1321 99
rect 1377 43 1463 99
rect 1519 43 1605 99
rect 1661 43 1747 99
rect 1803 43 1889 99
rect 1945 43 2031 99
rect 2087 43 2173 99
rect 2229 43 2315 99
rect 2371 43 2457 99
rect 2513 43 2599 99
rect 2655 43 2741 99
rect 2797 43 2883 99
rect 2939 43 3025 99
rect 3081 43 3167 99
rect 3223 43 3309 99
rect 3365 43 3451 99
rect 3507 43 3593 99
rect 3649 43 3735 99
rect 3791 43 3877 99
rect 3933 43 4019 99
rect 4075 43 4161 99
rect 4217 43 4303 99
rect 4359 43 4445 99
rect 4501 43 4587 99
rect 4643 43 4729 99
rect 4785 43 4871 99
rect 4927 43 5013 99
rect 5069 43 5155 99
rect 5211 43 5297 99
rect 5353 43 5439 99
rect 5495 43 5581 99
rect 5637 43 5723 99
rect 5779 43 5865 99
rect 5921 43 6007 99
rect 6063 43 6149 99
rect 6205 43 6291 99
rect 6347 43 6433 99
rect 6489 43 6575 99
rect 6631 43 6717 99
rect 6773 43 6859 99
rect 6915 43 7001 99
rect 7057 43 7143 99
rect 7199 43 7285 99
rect 7341 43 7351 99
rect -7351 -43 7351 43
rect -7351 -99 -7341 -43
rect -7285 -99 -7199 -43
rect -7143 -99 -7057 -43
rect -7001 -99 -6915 -43
rect -6859 -99 -6773 -43
rect -6717 -99 -6631 -43
rect -6575 -99 -6489 -43
rect -6433 -99 -6347 -43
rect -6291 -99 -6205 -43
rect -6149 -99 -6063 -43
rect -6007 -99 -5921 -43
rect -5865 -99 -5779 -43
rect -5723 -99 -5637 -43
rect -5581 -99 -5495 -43
rect -5439 -99 -5353 -43
rect -5297 -99 -5211 -43
rect -5155 -99 -5069 -43
rect -5013 -99 -4927 -43
rect -4871 -99 -4785 -43
rect -4729 -99 -4643 -43
rect -4587 -99 -4501 -43
rect -4445 -99 -4359 -43
rect -4303 -99 -4217 -43
rect -4161 -99 -4075 -43
rect -4019 -99 -3933 -43
rect -3877 -99 -3791 -43
rect -3735 -99 -3649 -43
rect -3593 -99 -3507 -43
rect -3451 -99 -3365 -43
rect -3309 -99 -3223 -43
rect -3167 -99 -3081 -43
rect -3025 -99 -2939 -43
rect -2883 -99 -2797 -43
rect -2741 -99 -2655 -43
rect -2599 -99 -2513 -43
rect -2457 -99 -2371 -43
rect -2315 -99 -2229 -43
rect -2173 -99 -2087 -43
rect -2031 -99 -1945 -43
rect -1889 -99 -1803 -43
rect -1747 -99 -1661 -43
rect -1605 -99 -1519 -43
rect -1463 -99 -1377 -43
rect -1321 -99 -1235 -43
rect -1179 -99 -1093 -43
rect -1037 -99 -951 -43
rect -895 -99 -809 -43
rect -753 -99 -667 -43
rect -611 -99 -525 -43
rect -469 -99 -383 -43
rect -327 -99 -241 -43
rect -185 -99 -99 -43
rect -43 -99 43 -43
rect 99 -99 185 -43
rect 241 -99 327 -43
rect 383 -99 469 -43
rect 525 -99 611 -43
rect 667 -99 753 -43
rect 809 -99 895 -43
rect 951 -99 1037 -43
rect 1093 -99 1179 -43
rect 1235 -99 1321 -43
rect 1377 -99 1463 -43
rect 1519 -99 1605 -43
rect 1661 -99 1747 -43
rect 1803 -99 1889 -43
rect 1945 -99 2031 -43
rect 2087 -99 2173 -43
rect 2229 -99 2315 -43
rect 2371 -99 2457 -43
rect 2513 -99 2599 -43
rect 2655 -99 2741 -43
rect 2797 -99 2883 -43
rect 2939 -99 3025 -43
rect 3081 -99 3167 -43
rect 3223 -99 3309 -43
rect 3365 -99 3451 -43
rect 3507 -99 3593 -43
rect 3649 -99 3735 -43
rect 3791 -99 3877 -43
rect 3933 -99 4019 -43
rect 4075 -99 4161 -43
rect 4217 -99 4303 -43
rect 4359 -99 4445 -43
rect 4501 -99 4587 -43
rect 4643 -99 4729 -43
rect 4785 -99 4871 -43
rect 4927 -99 5013 -43
rect 5069 -99 5155 -43
rect 5211 -99 5297 -43
rect 5353 -99 5439 -43
rect 5495 -99 5581 -43
rect 5637 -99 5723 -43
rect 5779 -99 5865 -43
rect 5921 -99 6007 -43
rect 6063 -99 6149 -43
rect 6205 -99 6291 -43
rect 6347 -99 6433 -43
rect 6489 -99 6575 -43
rect 6631 -99 6717 -43
rect 6773 -99 6859 -43
rect 6915 -99 7001 -43
rect 7057 -99 7143 -43
rect 7199 -99 7285 -43
rect 7341 -99 7351 -43
rect -7351 -185 7351 -99
rect -7351 -241 -7341 -185
rect -7285 -241 -7199 -185
rect -7143 -241 -7057 -185
rect -7001 -241 -6915 -185
rect -6859 -241 -6773 -185
rect -6717 -241 -6631 -185
rect -6575 -241 -6489 -185
rect -6433 -241 -6347 -185
rect -6291 -241 -6205 -185
rect -6149 -241 -6063 -185
rect -6007 -241 -5921 -185
rect -5865 -241 -5779 -185
rect -5723 -241 -5637 -185
rect -5581 -241 -5495 -185
rect -5439 -241 -5353 -185
rect -5297 -241 -5211 -185
rect -5155 -241 -5069 -185
rect -5013 -241 -4927 -185
rect -4871 -241 -4785 -185
rect -4729 -241 -4643 -185
rect -4587 -241 -4501 -185
rect -4445 -241 -4359 -185
rect -4303 -241 -4217 -185
rect -4161 -241 -4075 -185
rect -4019 -241 -3933 -185
rect -3877 -241 -3791 -185
rect -3735 -241 -3649 -185
rect -3593 -241 -3507 -185
rect -3451 -241 -3365 -185
rect -3309 -241 -3223 -185
rect -3167 -241 -3081 -185
rect -3025 -241 -2939 -185
rect -2883 -241 -2797 -185
rect -2741 -241 -2655 -185
rect -2599 -241 -2513 -185
rect -2457 -241 -2371 -185
rect -2315 -241 -2229 -185
rect -2173 -241 -2087 -185
rect -2031 -241 -1945 -185
rect -1889 -241 -1803 -185
rect -1747 -241 -1661 -185
rect -1605 -241 -1519 -185
rect -1463 -241 -1377 -185
rect -1321 -241 -1235 -185
rect -1179 -241 -1093 -185
rect -1037 -241 -951 -185
rect -895 -241 -809 -185
rect -753 -241 -667 -185
rect -611 -241 -525 -185
rect -469 -241 -383 -185
rect -327 -241 -241 -185
rect -185 -241 -99 -185
rect -43 -241 43 -185
rect 99 -241 185 -185
rect 241 -241 327 -185
rect 383 -241 469 -185
rect 525 -241 611 -185
rect 667 -241 753 -185
rect 809 -241 895 -185
rect 951 -241 1037 -185
rect 1093 -241 1179 -185
rect 1235 -241 1321 -185
rect 1377 -241 1463 -185
rect 1519 -241 1605 -185
rect 1661 -241 1747 -185
rect 1803 -241 1889 -185
rect 1945 -241 2031 -185
rect 2087 -241 2173 -185
rect 2229 -241 2315 -185
rect 2371 -241 2457 -185
rect 2513 -241 2599 -185
rect 2655 -241 2741 -185
rect 2797 -241 2883 -185
rect 2939 -241 3025 -185
rect 3081 -241 3167 -185
rect 3223 -241 3309 -185
rect 3365 -241 3451 -185
rect 3507 -241 3593 -185
rect 3649 -241 3735 -185
rect 3791 -241 3877 -185
rect 3933 -241 4019 -185
rect 4075 -241 4161 -185
rect 4217 -241 4303 -185
rect 4359 -241 4445 -185
rect 4501 -241 4587 -185
rect 4643 -241 4729 -185
rect 4785 -241 4871 -185
rect 4927 -241 5013 -185
rect 5069 -241 5155 -185
rect 5211 -241 5297 -185
rect 5353 -241 5439 -185
rect 5495 -241 5581 -185
rect 5637 -241 5723 -185
rect 5779 -241 5865 -185
rect 5921 -241 6007 -185
rect 6063 -241 6149 -185
rect 6205 -241 6291 -185
rect 6347 -241 6433 -185
rect 6489 -241 6575 -185
rect 6631 -241 6717 -185
rect 6773 -241 6859 -185
rect 6915 -241 7001 -185
rect 7057 -241 7143 -185
rect 7199 -241 7285 -185
rect 7341 -241 7351 -185
rect -7351 -327 7351 -241
rect -7351 -383 -7341 -327
rect -7285 -383 -7199 -327
rect -7143 -383 -7057 -327
rect -7001 -383 -6915 -327
rect -6859 -383 -6773 -327
rect -6717 -383 -6631 -327
rect -6575 -383 -6489 -327
rect -6433 -383 -6347 -327
rect -6291 -383 -6205 -327
rect -6149 -383 -6063 -327
rect -6007 -383 -5921 -327
rect -5865 -383 -5779 -327
rect -5723 -383 -5637 -327
rect -5581 -383 -5495 -327
rect -5439 -383 -5353 -327
rect -5297 -383 -5211 -327
rect -5155 -383 -5069 -327
rect -5013 -383 -4927 -327
rect -4871 -383 -4785 -327
rect -4729 -383 -4643 -327
rect -4587 -383 -4501 -327
rect -4445 -383 -4359 -327
rect -4303 -383 -4217 -327
rect -4161 -383 -4075 -327
rect -4019 -383 -3933 -327
rect -3877 -383 -3791 -327
rect -3735 -383 -3649 -327
rect -3593 -383 -3507 -327
rect -3451 -383 -3365 -327
rect -3309 -383 -3223 -327
rect -3167 -383 -3081 -327
rect -3025 -383 -2939 -327
rect -2883 -383 -2797 -327
rect -2741 -383 -2655 -327
rect -2599 -383 -2513 -327
rect -2457 -383 -2371 -327
rect -2315 -383 -2229 -327
rect -2173 -383 -2087 -327
rect -2031 -383 -1945 -327
rect -1889 -383 -1803 -327
rect -1747 -383 -1661 -327
rect -1605 -383 -1519 -327
rect -1463 -383 -1377 -327
rect -1321 -383 -1235 -327
rect -1179 -383 -1093 -327
rect -1037 -383 -951 -327
rect -895 -383 -809 -327
rect -753 -383 -667 -327
rect -611 -383 -525 -327
rect -469 -383 -383 -327
rect -327 -383 -241 -327
rect -185 -383 -99 -327
rect -43 -383 43 -327
rect 99 -383 185 -327
rect 241 -383 327 -327
rect 383 -383 469 -327
rect 525 -383 611 -327
rect 667 -383 753 -327
rect 809 -383 895 -327
rect 951 -383 1037 -327
rect 1093 -383 1179 -327
rect 1235 -383 1321 -327
rect 1377 -383 1463 -327
rect 1519 -383 1605 -327
rect 1661 -383 1747 -327
rect 1803 -383 1889 -327
rect 1945 -383 2031 -327
rect 2087 -383 2173 -327
rect 2229 -383 2315 -327
rect 2371 -383 2457 -327
rect 2513 -383 2599 -327
rect 2655 -383 2741 -327
rect 2797 -383 2883 -327
rect 2939 -383 3025 -327
rect 3081 -383 3167 -327
rect 3223 -383 3309 -327
rect 3365 -383 3451 -327
rect 3507 -383 3593 -327
rect 3649 -383 3735 -327
rect 3791 -383 3877 -327
rect 3933 -383 4019 -327
rect 4075 -383 4161 -327
rect 4217 -383 4303 -327
rect 4359 -383 4445 -327
rect 4501 -383 4587 -327
rect 4643 -383 4729 -327
rect 4785 -383 4871 -327
rect 4927 -383 5013 -327
rect 5069 -383 5155 -327
rect 5211 -383 5297 -327
rect 5353 -383 5439 -327
rect 5495 -383 5581 -327
rect 5637 -383 5723 -327
rect 5779 -383 5865 -327
rect 5921 -383 6007 -327
rect 6063 -383 6149 -327
rect 6205 -383 6291 -327
rect 6347 -383 6433 -327
rect 6489 -383 6575 -327
rect 6631 -383 6717 -327
rect 6773 -383 6859 -327
rect 6915 -383 7001 -327
rect 7057 -383 7143 -327
rect 7199 -383 7285 -327
rect 7341 -383 7351 -327
rect -7351 -469 7351 -383
rect -7351 -525 -7341 -469
rect -7285 -525 -7199 -469
rect -7143 -525 -7057 -469
rect -7001 -525 -6915 -469
rect -6859 -525 -6773 -469
rect -6717 -525 -6631 -469
rect -6575 -525 -6489 -469
rect -6433 -525 -6347 -469
rect -6291 -525 -6205 -469
rect -6149 -525 -6063 -469
rect -6007 -525 -5921 -469
rect -5865 -525 -5779 -469
rect -5723 -525 -5637 -469
rect -5581 -525 -5495 -469
rect -5439 -525 -5353 -469
rect -5297 -525 -5211 -469
rect -5155 -525 -5069 -469
rect -5013 -525 -4927 -469
rect -4871 -525 -4785 -469
rect -4729 -525 -4643 -469
rect -4587 -525 -4501 -469
rect -4445 -525 -4359 -469
rect -4303 -525 -4217 -469
rect -4161 -525 -4075 -469
rect -4019 -525 -3933 -469
rect -3877 -525 -3791 -469
rect -3735 -525 -3649 -469
rect -3593 -525 -3507 -469
rect -3451 -525 -3365 -469
rect -3309 -525 -3223 -469
rect -3167 -525 -3081 -469
rect -3025 -525 -2939 -469
rect -2883 -525 -2797 -469
rect -2741 -525 -2655 -469
rect -2599 -525 -2513 -469
rect -2457 -525 -2371 -469
rect -2315 -525 -2229 -469
rect -2173 -525 -2087 -469
rect -2031 -525 -1945 -469
rect -1889 -525 -1803 -469
rect -1747 -525 -1661 -469
rect -1605 -525 -1519 -469
rect -1463 -525 -1377 -469
rect -1321 -525 -1235 -469
rect -1179 -525 -1093 -469
rect -1037 -525 -951 -469
rect -895 -525 -809 -469
rect -753 -525 -667 -469
rect -611 -525 -525 -469
rect -469 -525 -383 -469
rect -327 -525 -241 -469
rect -185 -525 -99 -469
rect -43 -525 43 -469
rect 99 -525 185 -469
rect 241 -525 327 -469
rect 383 -525 469 -469
rect 525 -525 611 -469
rect 667 -525 753 -469
rect 809 -525 895 -469
rect 951 -525 1037 -469
rect 1093 -525 1179 -469
rect 1235 -525 1321 -469
rect 1377 -525 1463 -469
rect 1519 -525 1605 -469
rect 1661 -525 1747 -469
rect 1803 -525 1889 -469
rect 1945 -525 2031 -469
rect 2087 -525 2173 -469
rect 2229 -525 2315 -469
rect 2371 -525 2457 -469
rect 2513 -525 2599 -469
rect 2655 -525 2741 -469
rect 2797 -525 2883 -469
rect 2939 -525 3025 -469
rect 3081 -525 3167 -469
rect 3223 -525 3309 -469
rect 3365 -525 3451 -469
rect 3507 -525 3593 -469
rect 3649 -525 3735 -469
rect 3791 -525 3877 -469
rect 3933 -525 4019 -469
rect 4075 -525 4161 -469
rect 4217 -525 4303 -469
rect 4359 -525 4445 -469
rect 4501 -525 4587 -469
rect 4643 -525 4729 -469
rect 4785 -525 4871 -469
rect 4927 -525 5013 -469
rect 5069 -525 5155 -469
rect 5211 -525 5297 -469
rect 5353 -525 5439 -469
rect 5495 -525 5581 -469
rect 5637 -525 5723 -469
rect 5779 -525 5865 -469
rect 5921 -525 6007 -469
rect 6063 -525 6149 -469
rect 6205 -525 6291 -469
rect 6347 -525 6433 -469
rect 6489 -525 6575 -469
rect 6631 -525 6717 -469
rect 6773 -525 6859 -469
rect 6915 -525 7001 -469
rect 7057 -525 7143 -469
rect 7199 -525 7285 -469
rect 7341 -525 7351 -469
rect -7351 -611 7351 -525
rect -7351 -667 -7341 -611
rect -7285 -667 -7199 -611
rect -7143 -667 -7057 -611
rect -7001 -667 -6915 -611
rect -6859 -667 -6773 -611
rect -6717 -667 -6631 -611
rect -6575 -667 -6489 -611
rect -6433 -667 -6347 -611
rect -6291 -667 -6205 -611
rect -6149 -667 -6063 -611
rect -6007 -667 -5921 -611
rect -5865 -667 -5779 -611
rect -5723 -667 -5637 -611
rect -5581 -667 -5495 -611
rect -5439 -667 -5353 -611
rect -5297 -667 -5211 -611
rect -5155 -667 -5069 -611
rect -5013 -667 -4927 -611
rect -4871 -667 -4785 -611
rect -4729 -667 -4643 -611
rect -4587 -667 -4501 -611
rect -4445 -667 -4359 -611
rect -4303 -667 -4217 -611
rect -4161 -667 -4075 -611
rect -4019 -667 -3933 -611
rect -3877 -667 -3791 -611
rect -3735 -667 -3649 -611
rect -3593 -667 -3507 -611
rect -3451 -667 -3365 -611
rect -3309 -667 -3223 -611
rect -3167 -667 -3081 -611
rect -3025 -667 -2939 -611
rect -2883 -667 -2797 -611
rect -2741 -667 -2655 -611
rect -2599 -667 -2513 -611
rect -2457 -667 -2371 -611
rect -2315 -667 -2229 -611
rect -2173 -667 -2087 -611
rect -2031 -667 -1945 -611
rect -1889 -667 -1803 -611
rect -1747 -667 -1661 -611
rect -1605 -667 -1519 -611
rect -1463 -667 -1377 -611
rect -1321 -667 -1235 -611
rect -1179 -667 -1093 -611
rect -1037 -667 -951 -611
rect -895 -667 -809 -611
rect -753 -667 -667 -611
rect -611 -667 -525 -611
rect -469 -667 -383 -611
rect -327 -667 -241 -611
rect -185 -667 -99 -611
rect -43 -667 43 -611
rect 99 -667 185 -611
rect 241 -667 327 -611
rect 383 -667 469 -611
rect 525 -667 611 -611
rect 667 -667 753 -611
rect 809 -667 895 -611
rect 951 -667 1037 -611
rect 1093 -667 1179 -611
rect 1235 -667 1321 -611
rect 1377 -667 1463 -611
rect 1519 -667 1605 -611
rect 1661 -667 1747 -611
rect 1803 -667 1889 -611
rect 1945 -667 2031 -611
rect 2087 -667 2173 -611
rect 2229 -667 2315 -611
rect 2371 -667 2457 -611
rect 2513 -667 2599 -611
rect 2655 -667 2741 -611
rect 2797 -667 2883 -611
rect 2939 -667 3025 -611
rect 3081 -667 3167 -611
rect 3223 -667 3309 -611
rect 3365 -667 3451 -611
rect 3507 -667 3593 -611
rect 3649 -667 3735 -611
rect 3791 -667 3877 -611
rect 3933 -667 4019 -611
rect 4075 -667 4161 -611
rect 4217 -667 4303 -611
rect 4359 -667 4445 -611
rect 4501 -667 4587 -611
rect 4643 -667 4729 -611
rect 4785 -667 4871 -611
rect 4927 -667 5013 -611
rect 5069 -667 5155 -611
rect 5211 -667 5297 -611
rect 5353 -667 5439 -611
rect 5495 -667 5581 -611
rect 5637 -667 5723 -611
rect 5779 -667 5865 -611
rect 5921 -667 6007 -611
rect 6063 -667 6149 -611
rect 6205 -667 6291 -611
rect 6347 -667 6433 -611
rect 6489 -667 6575 -611
rect 6631 -667 6717 -611
rect 6773 -667 6859 -611
rect 6915 -667 7001 -611
rect 7057 -667 7143 -611
rect 7199 -667 7285 -611
rect 7341 -667 7351 -611
rect -7351 -677 7351 -667
<< via3 >>
rect -7341 611 -7285 667
rect -7199 611 -7143 667
rect -7057 611 -7001 667
rect -6915 611 -6859 667
rect -6773 611 -6717 667
rect -6631 611 -6575 667
rect -6489 611 -6433 667
rect -6347 611 -6291 667
rect -6205 611 -6149 667
rect -6063 611 -6007 667
rect -5921 611 -5865 667
rect -5779 611 -5723 667
rect -5637 611 -5581 667
rect -5495 611 -5439 667
rect -5353 611 -5297 667
rect -5211 611 -5155 667
rect -5069 611 -5013 667
rect -4927 611 -4871 667
rect -4785 611 -4729 667
rect -4643 611 -4587 667
rect -4501 611 -4445 667
rect -4359 611 -4303 667
rect -4217 611 -4161 667
rect -4075 611 -4019 667
rect -3933 611 -3877 667
rect -3791 611 -3735 667
rect -3649 611 -3593 667
rect -3507 611 -3451 667
rect -3365 611 -3309 667
rect -3223 611 -3167 667
rect -3081 611 -3025 667
rect -2939 611 -2883 667
rect -2797 611 -2741 667
rect -2655 611 -2599 667
rect -2513 611 -2457 667
rect -2371 611 -2315 667
rect -2229 611 -2173 667
rect -2087 611 -2031 667
rect -1945 611 -1889 667
rect -1803 611 -1747 667
rect -1661 611 -1605 667
rect -1519 611 -1463 667
rect -1377 611 -1321 667
rect -1235 611 -1179 667
rect -1093 611 -1037 667
rect -951 611 -895 667
rect -809 611 -753 667
rect -667 611 -611 667
rect -525 611 -469 667
rect -383 611 -327 667
rect -241 611 -185 667
rect -99 611 -43 667
rect 43 611 99 667
rect 185 611 241 667
rect 327 611 383 667
rect 469 611 525 667
rect 611 611 667 667
rect 753 611 809 667
rect 895 611 951 667
rect 1037 611 1093 667
rect 1179 611 1235 667
rect 1321 611 1377 667
rect 1463 611 1519 667
rect 1605 611 1661 667
rect 1747 611 1803 667
rect 1889 611 1945 667
rect 2031 611 2087 667
rect 2173 611 2229 667
rect 2315 611 2371 667
rect 2457 611 2513 667
rect 2599 611 2655 667
rect 2741 611 2797 667
rect 2883 611 2939 667
rect 3025 611 3081 667
rect 3167 611 3223 667
rect 3309 611 3365 667
rect 3451 611 3507 667
rect 3593 611 3649 667
rect 3735 611 3791 667
rect 3877 611 3933 667
rect 4019 611 4075 667
rect 4161 611 4217 667
rect 4303 611 4359 667
rect 4445 611 4501 667
rect 4587 611 4643 667
rect 4729 611 4785 667
rect 4871 611 4927 667
rect 5013 611 5069 667
rect 5155 611 5211 667
rect 5297 611 5353 667
rect 5439 611 5495 667
rect 5581 611 5637 667
rect 5723 611 5779 667
rect 5865 611 5921 667
rect 6007 611 6063 667
rect 6149 611 6205 667
rect 6291 611 6347 667
rect 6433 611 6489 667
rect 6575 611 6631 667
rect 6717 611 6773 667
rect 6859 611 6915 667
rect 7001 611 7057 667
rect 7143 611 7199 667
rect 7285 611 7341 667
rect -7341 469 -7285 525
rect -7199 469 -7143 525
rect -7057 469 -7001 525
rect -6915 469 -6859 525
rect -6773 469 -6717 525
rect -6631 469 -6575 525
rect -6489 469 -6433 525
rect -6347 469 -6291 525
rect -6205 469 -6149 525
rect -6063 469 -6007 525
rect -5921 469 -5865 525
rect -5779 469 -5723 525
rect -5637 469 -5581 525
rect -5495 469 -5439 525
rect -5353 469 -5297 525
rect -5211 469 -5155 525
rect -5069 469 -5013 525
rect -4927 469 -4871 525
rect -4785 469 -4729 525
rect -4643 469 -4587 525
rect -4501 469 -4445 525
rect -4359 469 -4303 525
rect -4217 469 -4161 525
rect -4075 469 -4019 525
rect -3933 469 -3877 525
rect -3791 469 -3735 525
rect -3649 469 -3593 525
rect -3507 469 -3451 525
rect -3365 469 -3309 525
rect -3223 469 -3167 525
rect -3081 469 -3025 525
rect -2939 469 -2883 525
rect -2797 469 -2741 525
rect -2655 469 -2599 525
rect -2513 469 -2457 525
rect -2371 469 -2315 525
rect -2229 469 -2173 525
rect -2087 469 -2031 525
rect -1945 469 -1889 525
rect -1803 469 -1747 525
rect -1661 469 -1605 525
rect -1519 469 -1463 525
rect -1377 469 -1321 525
rect -1235 469 -1179 525
rect -1093 469 -1037 525
rect -951 469 -895 525
rect -809 469 -753 525
rect -667 469 -611 525
rect -525 469 -469 525
rect -383 469 -327 525
rect -241 469 -185 525
rect -99 469 -43 525
rect 43 469 99 525
rect 185 469 241 525
rect 327 469 383 525
rect 469 469 525 525
rect 611 469 667 525
rect 753 469 809 525
rect 895 469 951 525
rect 1037 469 1093 525
rect 1179 469 1235 525
rect 1321 469 1377 525
rect 1463 469 1519 525
rect 1605 469 1661 525
rect 1747 469 1803 525
rect 1889 469 1945 525
rect 2031 469 2087 525
rect 2173 469 2229 525
rect 2315 469 2371 525
rect 2457 469 2513 525
rect 2599 469 2655 525
rect 2741 469 2797 525
rect 2883 469 2939 525
rect 3025 469 3081 525
rect 3167 469 3223 525
rect 3309 469 3365 525
rect 3451 469 3507 525
rect 3593 469 3649 525
rect 3735 469 3791 525
rect 3877 469 3933 525
rect 4019 469 4075 525
rect 4161 469 4217 525
rect 4303 469 4359 525
rect 4445 469 4501 525
rect 4587 469 4643 525
rect 4729 469 4785 525
rect 4871 469 4927 525
rect 5013 469 5069 525
rect 5155 469 5211 525
rect 5297 469 5353 525
rect 5439 469 5495 525
rect 5581 469 5637 525
rect 5723 469 5779 525
rect 5865 469 5921 525
rect 6007 469 6063 525
rect 6149 469 6205 525
rect 6291 469 6347 525
rect 6433 469 6489 525
rect 6575 469 6631 525
rect 6717 469 6773 525
rect 6859 469 6915 525
rect 7001 469 7057 525
rect 7143 469 7199 525
rect 7285 469 7341 525
rect -7341 327 -7285 383
rect -7199 327 -7143 383
rect -7057 327 -7001 383
rect -6915 327 -6859 383
rect -6773 327 -6717 383
rect -6631 327 -6575 383
rect -6489 327 -6433 383
rect -6347 327 -6291 383
rect -6205 327 -6149 383
rect -6063 327 -6007 383
rect -5921 327 -5865 383
rect -5779 327 -5723 383
rect -5637 327 -5581 383
rect -5495 327 -5439 383
rect -5353 327 -5297 383
rect -5211 327 -5155 383
rect -5069 327 -5013 383
rect -4927 327 -4871 383
rect -4785 327 -4729 383
rect -4643 327 -4587 383
rect -4501 327 -4445 383
rect -4359 327 -4303 383
rect -4217 327 -4161 383
rect -4075 327 -4019 383
rect -3933 327 -3877 383
rect -3791 327 -3735 383
rect -3649 327 -3593 383
rect -3507 327 -3451 383
rect -3365 327 -3309 383
rect -3223 327 -3167 383
rect -3081 327 -3025 383
rect -2939 327 -2883 383
rect -2797 327 -2741 383
rect -2655 327 -2599 383
rect -2513 327 -2457 383
rect -2371 327 -2315 383
rect -2229 327 -2173 383
rect -2087 327 -2031 383
rect -1945 327 -1889 383
rect -1803 327 -1747 383
rect -1661 327 -1605 383
rect -1519 327 -1463 383
rect -1377 327 -1321 383
rect -1235 327 -1179 383
rect -1093 327 -1037 383
rect -951 327 -895 383
rect -809 327 -753 383
rect -667 327 -611 383
rect -525 327 -469 383
rect -383 327 -327 383
rect -241 327 -185 383
rect -99 327 -43 383
rect 43 327 99 383
rect 185 327 241 383
rect 327 327 383 383
rect 469 327 525 383
rect 611 327 667 383
rect 753 327 809 383
rect 895 327 951 383
rect 1037 327 1093 383
rect 1179 327 1235 383
rect 1321 327 1377 383
rect 1463 327 1519 383
rect 1605 327 1661 383
rect 1747 327 1803 383
rect 1889 327 1945 383
rect 2031 327 2087 383
rect 2173 327 2229 383
rect 2315 327 2371 383
rect 2457 327 2513 383
rect 2599 327 2655 383
rect 2741 327 2797 383
rect 2883 327 2939 383
rect 3025 327 3081 383
rect 3167 327 3223 383
rect 3309 327 3365 383
rect 3451 327 3507 383
rect 3593 327 3649 383
rect 3735 327 3791 383
rect 3877 327 3933 383
rect 4019 327 4075 383
rect 4161 327 4217 383
rect 4303 327 4359 383
rect 4445 327 4501 383
rect 4587 327 4643 383
rect 4729 327 4785 383
rect 4871 327 4927 383
rect 5013 327 5069 383
rect 5155 327 5211 383
rect 5297 327 5353 383
rect 5439 327 5495 383
rect 5581 327 5637 383
rect 5723 327 5779 383
rect 5865 327 5921 383
rect 6007 327 6063 383
rect 6149 327 6205 383
rect 6291 327 6347 383
rect 6433 327 6489 383
rect 6575 327 6631 383
rect 6717 327 6773 383
rect 6859 327 6915 383
rect 7001 327 7057 383
rect 7143 327 7199 383
rect 7285 327 7341 383
rect -7341 185 -7285 241
rect -7199 185 -7143 241
rect -7057 185 -7001 241
rect -6915 185 -6859 241
rect -6773 185 -6717 241
rect -6631 185 -6575 241
rect -6489 185 -6433 241
rect -6347 185 -6291 241
rect -6205 185 -6149 241
rect -6063 185 -6007 241
rect -5921 185 -5865 241
rect -5779 185 -5723 241
rect -5637 185 -5581 241
rect -5495 185 -5439 241
rect -5353 185 -5297 241
rect -5211 185 -5155 241
rect -5069 185 -5013 241
rect -4927 185 -4871 241
rect -4785 185 -4729 241
rect -4643 185 -4587 241
rect -4501 185 -4445 241
rect -4359 185 -4303 241
rect -4217 185 -4161 241
rect -4075 185 -4019 241
rect -3933 185 -3877 241
rect -3791 185 -3735 241
rect -3649 185 -3593 241
rect -3507 185 -3451 241
rect -3365 185 -3309 241
rect -3223 185 -3167 241
rect -3081 185 -3025 241
rect -2939 185 -2883 241
rect -2797 185 -2741 241
rect -2655 185 -2599 241
rect -2513 185 -2457 241
rect -2371 185 -2315 241
rect -2229 185 -2173 241
rect -2087 185 -2031 241
rect -1945 185 -1889 241
rect -1803 185 -1747 241
rect -1661 185 -1605 241
rect -1519 185 -1463 241
rect -1377 185 -1321 241
rect -1235 185 -1179 241
rect -1093 185 -1037 241
rect -951 185 -895 241
rect -809 185 -753 241
rect -667 185 -611 241
rect -525 185 -469 241
rect -383 185 -327 241
rect -241 185 -185 241
rect -99 185 -43 241
rect 43 185 99 241
rect 185 185 241 241
rect 327 185 383 241
rect 469 185 525 241
rect 611 185 667 241
rect 753 185 809 241
rect 895 185 951 241
rect 1037 185 1093 241
rect 1179 185 1235 241
rect 1321 185 1377 241
rect 1463 185 1519 241
rect 1605 185 1661 241
rect 1747 185 1803 241
rect 1889 185 1945 241
rect 2031 185 2087 241
rect 2173 185 2229 241
rect 2315 185 2371 241
rect 2457 185 2513 241
rect 2599 185 2655 241
rect 2741 185 2797 241
rect 2883 185 2939 241
rect 3025 185 3081 241
rect 3167 185 3223 241
rect 3309 185 3365 241
rect 3451 185 3507 241
rect 3593 185 3649 241
rect 3735 185 3791 241
rect 3877 185 3933 241
rect 4019 185 4075 241
rect 4161 185 4217 241
rect 4303 185 4359 241
rect 4445 185 4501 241
rect 4587 185 4643 241
rect 4729 185 4785 241
rect 4871 185 4927 241
rect 5013 185 5069 241
rect 5155 185 5211 241
rect 5297 185 5353 241
rect 5439 185 5495 241
rect 5581 185 5637 241
rect 5723 185 5779 241
rect 5865 185 5921 241
rect 6007 185 6063 241
rect 6149 185 6205 241
rect 6291 185 6347 241
rect 6433 185 6489 241
rect 6575 185 6631 241
rect 6717 185 6773 241
rect 6859 185 6915 241
rect 7001 185 7057 241
rect 7143 185 7199 241
rect 7285 185 7341 241
rect -7341 43 -7285 99
rect -7199 43 -7143 99
rect -7057 43 -7001 99
rect -6915 43 -6859 99
rect -6773 43 -6717 99
rect -6631 43 -6575 99
rect -6489 43 -6433 99
rect -6347 43 -6291 99
rect -6205 43 -6149 99
rect -6063 43 -6007 99
rect -5921 43 -5865 99
rect -5779 43 -5723 99
rect -5637 43 -5581 99
rect -5495 43 -5439 99
rect -5353 43 -5297 99
rect -5211 43 -5155 99
rect -5069 43 -5013 99
rect -4927 43 -4871 99
rect -4785 43 -4729 99
rect -4643 43 -4587 99
rect -4501 43 -4445 99
rect -4359 43 -4303 99
rect -4217 43 -4161 99
rect -4075 43 -4019 99
rect -3933 43 -3877 99
rect -3791 43 -3735 99
rect -3649 43 -3593 99
rect -3507 43 -3451 99
rect -3365 43 -3309 99
rect -3223 43 -3167 99
rect -3081 43 -3025 99
rect -2939 43 -2883 99
rect -2797 43 -2741 99
rect -2655 43 -2599 99
rect -2513 43 -2457 99
rect -2371 43 -2315 99
rect -2229 43 -2173 99
rect -2087 43 -2031 99
rect -1945 43 -1889 99
rect -1803 43 -1747 99
rect -1661 43 -1605 99
rect -1519 43 -1463 99
rect -1377 43 -1321 99
rect -1235 43 -1179 99
rect -1093 43 -1037 99
rect -951 43 -895 99
rect -809 43 -753 99
rect -667 43 -611 99
rect -525 43 -469 99
rect -383 43 -327 99
rect -241 43 -185 99
rect -99 43 -43 99
rect 43 43 99 99
rect 185 43 241 99
rect 327 43 383 99
rect 469 43 525 99
rect 611 43 667 99
rect 753 43 809 99
rect 895 43 951 99
rect 1037 43 1093 99
rect 1179 43 1235 99
rect 1321 43 1377 99
rect 1463 43 1519 99
rect 1605 43 1661 99
rect 1747 43 1803 99
rect 1889 43 1945 99
rect 2031 43 2087 99
rect 2173 43 2229 99
rect 2315 43 2371 99
rect 2457 43 2513 99
rect 2599 43 2655 99
rect 2741 43 2797 99
rect 2883 43 2939 99
rect 3025 43 3081 99
rect 3167 43 3223 99
rect 3309 43 3365 99
rect 3451 43 3507 99
rect 3593 43 3649 99
rect 3735 43 3791 99
rect 3877 43 3933 99
rect 4019 43 4075 99
rect 4161 43 4217 99
rect 4303 43 4359 99
rect 4445 43 4501 99
rect 4587 43 4643 99
rect 4729 43 4785 99
rect 4871 43 4927 99
rect 5013 43 5069 99
rect 5155 43 5211 99
rect 5297 43 5353 99
rect 5439 43 5495 99
rect 5581 43 5637 99
rect 5723 43 5779 99
rect 5865 43 5921 99
rect 6007 43 6063 99
rect 6149 43 6205 99
rect 6291 43 6347 99
rect 6433 43 6489 99
rect 6575 43 6631 99
rect 6717 43 6773 99
rect 6859 43 6915 99
rect 7001 43 7057 99
rect 7143 43 7199 99
rect 7285 43 7341 99
rect -7341 -99 -7285 -43
rect -7199 -99 -7143 -43
rect -7057 -99 -7001 -43
rect -6915 -99 -6859 -43
rect -6773 -99 -6717 -43
rect -6631 -99 -6575 -43
rect -6489 -99 -6433 -43
rect -6347 -99 -6291 -43
rect -6205 -99 -6149 -43
rect -6063 -99 -6007 -43
rect -5921 -99 -5865 -43
rect -5779 -99 -5723 -43
rect -5637 -99 -5581 -43
rect -5495 -99 -5439 -43
rect -5353 -99 -5297 -43
rect -5211 -99 -5155 -43
rect -5069 -99 -5013 -43
rect -4927 -99 -4871 -43
rect -4785 -99 -4729 -43
rect -4643 -99 -4587 -43
rect -4501 -99 -4445 -43
rect -4359 -99 -4303 -43
rect -4217 -99 -4161 -43
rect -4075 -99 -4019 -43
rect -3933 -99 -3877 -43
rect -3791 -99 -3735 -43
rect -3649 -99 -3593 -43
rect -3507 -99 -3451 -43
rect -3365 -99 -3309 -43
rect -3223 -99 -3167 -43
rect -3081 -99 -3025 -43
rect -2939 -99 -2883 -43
rect -2797 -99 -2741 -43
rect -2655 -99 -2599 -43
rect -2513 -99 -2457 -43
rect -2371 -99 -2315 -43
rect -2229 -99 -2173 -43
rect -2087 -99 -2031 -43
rect -1945 -99 -1889 -43
rect -1803 -99 -1747 -43
rect -1661 -99 -1605 -43
rect -1519 -99 -1463 -43
rect -1377 -99 -1321 -43
rect -1235 -99 -1179 -43
rect -1093 -99 -1037 -43
rect -951 -99 -895 -43
rect -809 -99 -753 -43
rect -667 -99 -611 -43
rect -525 -99 -469 -43
rect -383 -99 -327 -43
rect -241 -99 -185 -43
rect -99 -99 -43 -43
rect 43 -99 99 -43
rect 185 -99 241 -43
rect 327 -99 383 -43
rect 469 -99 525 -43
rect 611 -99 667 -43
rect 753 -99 809 -43
rect 895 -99 951 -43
rect 1037 -99 1093 -43
rect 1179 -99 1235 -43
rect 1321 -99 1377 -43
rect 1463 -99 1519 -43
rect 1605 -99 1661 -43
rect 1747 -99 1803 -43
rect 1889 -99 1945 -43
rect 2031 -99 2087 -43
rect 2173 -99 2229 -43
rect 2315 -99 2371 -43
rect 2457 -99 2513 -43
rect 2599 -99 2655 -43
rect 2741 -99 2797 -43
rect 2883 -99 2939 -43
rect 3025 -99 3081 -43
rect 3167 -99 3223 -43
rect 3309 -99 3365 -43
rect 3451 -99 3507 -43
rect 3593 -99 3649 -43
rect 3735 -99 3791 -43
rect 3877 -99 3933 -43
rect 4019 -99 4075 -43
rect 4161 -99 4217 -43
rect 4303 -99 4359 -43
rect 4445 -99 4501 -43
rect 4587 -99 4643 -43
rect 4729 -99 4785 -43
rect 4871 -99 4927 -43
rect 5013 -99 5069 -43
rect 5155 -99 5211 -43
rect 5297 -99 5353 -43
rect 5439 -99 5495 -43
rect 5581 -99 5637 -43
rect 5723 -99 5779 -43
rect 5865 -99 5921 -43
rect 6007 -99 6063 -43
rect 6149 -99 6205 -43
rect 6291 -99 6347 -43
rect 6433 -99 6489 -43
rect 6575 -99 6631 -43
rect 6717 -99 6773 -43
rect 6859 -99 6915 -43
rect 7001 -99 7057 -43
rect 7143 -99 7199 -43
rect 7285 -99 7341 -43
rect -7341 -241 -7285 -185
rect -7199 -241 -7143 -185
rect -7057 -241 -7001 -185
rect -6915 -241 -6859 -185
rect -6773 -241 -6717 -185
rect -6631 -241 -6575 -185
rect -6489 -241 -6433 -185
rect -6347 -241 -6291 -185
rect -6205 -241 -6149 -185
rect -6063 -241 -6007 -185
rect -5921 -241 -5865 -185
rect -5779 -241 -5723 -185
rect -5637 -241 -5581 -185
rect -5495 -241 -5439 -185
rect -5353 -241 -5297 -185
rect -5211 -241 -5155 -185
rect -5069 -241 -5013 -185
rect -4927 -241 -4871 -185
rect -4785 -241 -4729 -185
rect -4643 -241 -4587 -185
rect -4501 -241 -4445 -185
rect -4359 -241 -4303 -185
rect -4217 -241 -4161 -185
rect -4075 -241 -4019 -185
rect -3933 -241 -3877 -185
rect -3791 -241 -3735 -185
rect -3649 -241 -3593 -185
rect -3507 -241 -3451 -185
rect -3365 -241 -3309 -185
rect -3223 -241 -3167 -185
rect -3081 -241 -3025 -185
rect -2939 -241 -2883 -185
rect -2797 -241 -2741 -185
rect -2655 -241 -2599 -185
rect -2513 -241 -2457 -185
rect -2371 -241 -2315 -185
rect -2229 -241 -2173 -185
rect -2087 -241 -2031 -185
rect -1945 -241 -1889 -185
rect -1803 -241 -1747 -185
rect -1661 -241 -1605 -185
rect -1519 -241 -1463 -185
rect -1377 -241 -1321 -185
rect -1235 -241 -1179 -185
rect -1093 -241 -1037 -185
rect -951 -241 -895 -185
rect -809 -241 -753 -185
rect -667 -241 -611 -185
rect -525 -241 -469 -185
rect -383 -241 -327 -185
rect -241 -241 -185 -185
rect -99 -241 -43 -185
rect 43 -241 99 -185
rect 185 -241 241 -185
rect 327 -241 383 -185
rect 469 -241 525 -185
rect 611 -241 667 -185
rect 753 -241 809 -185
rect 895 -241 951 -185
rect 1037 -241 1093 -185
rect 1179 -241 1235 -185
rect 1321 -241 1377 -185
rect 1463 -241 1519 -185
rect 1605 -241 1661 -185
rect 1747 -241 1803 -185
rect 1889 -241 1945 -185
rect 2031 -241 2087 -185
rect 2173 -241 2229 -185
rect 2315 -241 2371 -185
rect 2457 -241 2513 -185
rect 2599 -241 2655 -185
rect 2741 -241 2797 -185
rect 2883 -241 2939 -185
rect 3025 -241 3081 -185
rect 3167 -241 3223 -185
rect 3309 -241 3365 -185
rect 3451 -241 3507 -185
rect 3593 -241 3649 -185
rect 3735 -241 3791 -185
rect 3877 -241 3933 -185
rect 4019 -241 4075 -185
rect 4161 -241 4217 -185
rect 4303 -241 4359 -185
rect 4445 -241 4501 -185
rect 4587 -241 4643 -185
rect 4729 -241 4785 -185
rect 4871 -241 4927 -185
rect 5013 -241 5069 -185
rect 5155 -241 5211 -185
rect 5297 -241 5353 -185
rect 5439 -241 5495 -185
rect 5581 -241 5637 -185
rect 5723 -241 5779 -185
rect 5865 -241 5921 -185
rect 6007 -241 6063 -185
rect 6149 -241 6205 -185
rect 6291 -241 6347 -185
rect 6433 -241 6489 -185
rect 6575 -241 6631 -185
rect 6717 -241 6773 -185
rect 6859 -241 6915 -185
rect 7001 -241 7057 -185
rect 7143 -241 7199 -185
rect 7285 -241 7341 -185
rect -7341 -383 -7285 -327
rect -7199 -383 -7143 -327
rect -7057 -383 -7001 -327
rect -6915 -383 -6859 -327
rect -6773 -383 -6717 -327
rect -6631 -383 -6575 -327
rect -6489 -383 -6433 -327
rect -6347 -383 -6291 -327
rect -6205 -383 -6149 -327
rect -6063 -383 -6007 -327
rect -5921 -383 -5865 -327
rect -5779 -383 -5723 -327
rect -5637 -383 -5581 -327
rect -5495 -383 -5439 -327
rect -5353 -383 -5297 -327
rect -5211 -383 -5155 -327
rect -5069 -383 -5013 -327
rect -4927 -383 -4871 -327
rect -4785 -383 -4729 -327
rect -4643 -383 -4587 -327
rect -4501 -383 -4445 -327
rect -4359 -383 -4303 -327
rect -4217 -383 -4161 -327
rect -4075 -383 -4019 -327
rect -3933 -383 -3877 -327
rect -3791 -383 -3735 -327
rect -3649 -383 -3593 -327
rect -3507 -383 -3451 -327
rect -3365 -383 -3309 -327
rect -3223 -383 -3167 -327
rect -3081 -383 -3025 -327
rect -2939 -383 -2883 -327
rect -2797 -383 -2741 -327
rect -2655 -383 -2599 -327
rect -2513 -383 -2457 -327
rect -2371 -383 -2315 -327
rect -2229 -383 -2173 -327
rect -2087 -383 -2031 -327
rect -1945 -383 -1889 -327
rect -1803 -383 -1747 -327
rect -1661 -383 -1605 -327
rect -1519 -383 -1463 -327
rect -1377 -383 -1321 -327
rect -1235 -383 -1179 -327
rect -1093 -383 -1037 -327
rect -951 -383 -895 -327
rect -809 -383 -753 -327
rect -667 -383 -611 -327
rect -525 -383 -469 -327
rect -383 -383 -327 -327
rect -241 -383 -185 -327
rect -99 -383 -43 -327
rect 43 -383 99 -327
rect 185 -383 241 -327
rect 327 -383 383 -327
rect 469 -383 525 -327
rect 611 -383 667 -327
rect 753 -383 809 -327
rect 895 -383 951 -327
rect 1037 -383 1093 -327
rect 1179 -383 1235 -327
rect 1321 -383 1377 -327
rect 1463 -383 1519 -327
rect 1605 -383 1661 -327
rect 1747 -383 1803 -327
rect 1889 -383 1945 -327
rect 2031 -383 2087 -327
rect 2173 -383 2229 -327
rect 2315 -383 2371 -327
rect 2457 -383 2513 -327
rect 2599 -383 2655 -327
rect 2741 -383 2797 -327
rect 2883 -383 2939 -327
rect 3025 -383 3081 -327
rect 3167 -383 3223 -327
rect 3309 -383 3365 -327
rect 3451 -383 3507 -327
rect 3593 -383 3649 -327
rect 3735 -383 3791 -327
rect 3877 -383 3933 -327
rect 4019 -383 4075 -327
rect 4161 -383 4217 -327
rect 4303 -383 4359 -327
rect 4445 -383 4501 -327
rect 4587 -383 4643 -327
rect 4729 -383 4785 -327
rect 4871 -383 4927 -327
rect 5013 -383 5069 -327
rect 5155 -383 5211 -327
rect 5297 -383 5353 -327
rect 5439 -383 5495 -327
rect 5581 -383 5637 -327
rect 5723 -383 5779 -327
rect 5865 -383 5921 -327
rect 6007 -383 6063 -327
rect 6149 -383 6205 -327
rect 6291 -383 6347 -327
rect 6433 -383 6489 -327
rect 6575 -383 6631 -327
rect 6717 -383 6773 -327
rect 6859 -383 6915 -327
rect 7001 -383 7057 -327
rect 7143 -383 7199 -327
rect 7285 -383 7341 -327
rect -7341 -525 -7285 -469
rect -7199 -525 -7143 -469
rect -7057 -525 -7001 -469
rect -6915 -525 -6859 -469
rect -6773 -525 -6717 -469
rect -6631 -525 -6575 -469
rect -6489 -525 -6433 -469
rect -6347 -525 -6291 -469
rect -6205 -525 -6149 -469
rect -6063 -525 -6007 -469
rect -5921 -525 -5865 -469
rect -5779 -525 -5723 -469
rect -5637 -525 -5581 -469
rect -5495 -525 -5439 -469
rect -5353 -525 -5297 -469
rect -5211 -525 -5155 -469
rect -5069 -525 -5013 -469
rect -4927 -525 -4871 -469
rect -4785 -525 -4729 -469
rect -4643 -525 -4587 -469
rect -4501 -525 -4445 -469
rect -4359 -525 -4303 -469
rect -4217 -525 -4161 -469
rect -4075 -525 -4019 -469
rect -3933 -525 -3877 -469
rect -3791 -525 -3735 -469
rect -3649 -525 -3593 -469
rect -3507 -525 -3451 -469
rect -3365 -525 -3309 -469
rect -3223 -525 -3167 -469
rect -3081 -525 -3025 -469
rect -2939 -525 -2883 -469
rect -2797 -525 -2741 -469
rect -2655 -525 -2599 -469
rect -2513 -525 -2457 -469
rect -2371 -525 -2315 -469
rect -2229 -525 -2173 -469
rect -2087 -525 -2031 -469
rect -1945 -525 -1889 -469
rect -1803 -525 -1747 -469
rect -1661 -525 -1605 -469
rect -1519 -525 -1463 -469
rect -1377 -525 -1321 -469
rect -1235 -525 -1179 -469
rect -1093 -525 -1037 -469
rect -951 -525 -895 -469
rect -809 -525 -753 -469
rect -667 -525 -611 -469
rect -525 -525 -469 -469
rect -383 -525 -327 -469
rect -241 -525 -185 -469
rect -99 -525 -43 -469
rect 43 -525 99 -469
rect 185 -525 241 -469
rect 327 -525 383 -469
rect 469 -525 525 -469
rect 611 -525 667 -469
rect 753 -525 809 -469
rect 895 -525 951 -469
rect 1037 -525 1093 -469
rect 1179 -525 1235 -469
rect 1321 -525 1377 -469
rect 1463 -525 1519 -469
rect 1605 -525 1661 -469
rect 1747 -525 1803 -469
rect 1889 -525 1945 -469
rect 2031 -525 2087 -469
rect 2173 -525 2229 -469
rect 2315 -525 2371 -469
rect 2457 -525 2513 -469
rect 2599 -525 2655 -469
rect 2741 -525 2797 -469
rect 2883 -525 2939 -469
rect 3025 -525 3081 -469
rect 3167 -525 3223 -469
rect 3309 -525 3365 -469
rect 3451 -525 3507 -469
rect 3593 -525 3649 -469
rect 3735 -525 3791 -469
rect 3877 -525 3933 -469
rect 4019 -525 4075 -469
rect 4161 -525 4217 -469
rect 4303 -525 4359 -469
rect 4445 -525 4501 -469
rect 4587 -525 4643 -469
rect 4729 -525 4785 -469
rect 4871 -525 4927 -469
rect 5013 -525 5069 -469
rect 5155 -525 5211 -469
rect 5297 -525 5353 -469
rect 5439 -525 5495 -469
rect 5581 -525 5637 -469
rect 5723 -525 5779 -469
rect 5865 -525 5921 -469
rect 6007 -525 6063 -469
rect 6149 -525 6205 -469
rect 6291 -525 6347 -469
rect 6433 -525 6489 -469
rect 6575 -525 6631 -469
rect 6717 -525 6773 -469
rect 6859 -525 6915 -469
rect 7001 -525 7057 -469
rect 7143 -525 7199 -469
rect 7285 -525 7341 -469
rect -7341 -667 -7285 -611
rect -7199 -667 -7143 -611
rect -7057 -667 -7001 -611
rect -6915 -667 -6859 -611
rect -6773 -667 -6717 -611
rect -6631 -667 -6575 -611
rect -6489 -667 -6433 -611
rect -6347 -667 -6291 -611
rect -6205 -667 -6149 -611
rect -6063 -667 -6007 -611
rect -5921 -667 -5865 -611
rect -5779 -667 -5723 -611
rect -5637 -667 -5581 -611
rect -5495 -667 -5439 -611
rect -5353 -667 -5297 -611
rect -5211 -667 -5155 -611
rect -5069 -667 -5013 -611
rect -4927 -667 -4871 -611
rect -4785 -667 -4729 -611
rect -4643 -667 -4587 -611
rect -4501 -667 -4445 -611
rect -4359 -667 -4303 -611
rect -4217 -667 -4161 -611
rect -4075 -667 -4019 -611
rect -3933 -667 -3877 -611
rect -3791 -667 -3735 -611
rect -3649 -667 -3593 -611
rect -3507 -667 -3451 -611
rect -3365 -667 -3309 -611
rect -3223 -667 -3167 -611
rect -3081 -667 -3025 -611
rect -2939 -667 -2883 -611
rect -2797 -667 -2741 -611
rect -2655 -667 -2599 -611
rect -2513 -667 -2457 -611
rect -2371 -667 -2315 -611
rect -2229 -667 -2173 -611
rect -2087 -667 -2031 -611
rect -1945 -667 -1889 -611
rect -1803 -667 -1747 -611
rect -1661 -667 -1605 -611
rect -1519 -667 -1463 -611
rect -1377 -667 -1321 -611
rect -1235 -667 -1179 -611
rect -1093 -667 -1037 -611
rect -951 -667 -895 -611
rect -809 -667 -753 -611
rect -667 -667 -611 -611
rect -525 -667 -469 -611
rect -383 -667 -327 -611
rect -241 -667 -185 -611
rect -99 -667 -43 -611
rect 43 -667 99 -611
rect 185 -667 241 -611
rect 327 -667 383 -611
rect 469 -667 525 -611
rect 611 -667 667 -611
rect 753 -667 809 -611
rect 895 -667 951 -611
rect 1037 -667 1093 -611
rect 1179 -667 1235 -611
rect 1321 -667 1377 -611
rect 1463 -667 1519 -611
rect 1605 -667 1661 -611
rect 1747 -667 1803 -611
rect 1889 -667 1945 -611
rect 2031 -667 2087 -611
rect 2173 -667 2229 -611
rect 2315 -667 2371 -611
rect 2457 -667 2513 -611
rect 2599 -667 2655 -611
rect 2741 -667 2797 -611
rect 2883 -667 2939 -611
rect 3025 -667 3081 -611
rect 3167 -667 3223 -611
rect 3309 -667 3365 -611
rect 3451 -667 3507 -611
rect 3593 -667 3649 -611
rect 3735 -667 3791 -611
rect 3877 -667 3933 -611
rect 4019 -667 4075 -611
rect 4161 -667 4217 -611
rect 4303 -667 4359 -611
rect 4445 -667 4501 -611
rect 4587 -667 4643 -611
rect 4729 -667 4785 -611
rect 4871 -667 4927 -611
rect 5013 -667 5069 -611
rect 5155 -667 5211 -611
rect 5297 -667 5353 -611
rect 5439 -667 5495 -611
rect 5581 -667 5637 -611
rect 5723 -667 5779 -611
rect 5865 -667 5921 -611
rect 6007 -667 6063 -611
rect 6149 -667 6205 -611
rect 6291 -667 6347 -611
rect 6433 -667 6489 -611
rect 6575 -667 6631 -611
rect 6717 -667 6773 -611
rect 6859 -667 6915 -611
rect 7001 -667 7057 -611
rect 7143 -667 7199 -611
rect 7285 -667 7341 -611
<< metal4 >>
rect -7351 667 7351 677
rect -7351 611 -7341 667
rect -7285 611 -7199 667
rect -7143 611 -7057 667
rect -7001 611 -6915 667
rect -6859 611 -6773 667
rect -6717 611 -6631 667
rect -6575 611 -6489 667
rect -6433 611 -6347 667
rect -6291 611 -6205 667
rect -6149 611 -6063 667
rect -6007 611 -5921 667
rect -5865 611 -5779 667
rect -5723 611 -5637 667
rect -5581 611 -5495 667
rect -5439 611 -5353 667
rect -5297 611 -5211 667
rect -5155 611 -5069 667
rect -5013 611 -4927 667
rect -4871 611 -4785 667
rect -4729 611 -4643 667
rect -4587 611 -4501 667
rect -4445 611 -4359 667
rect -4303 611 -4217 667
rect -4161 611 -4075 667
rect -4019 611 -3933 667
rect -3877 611 -3791 667
rect -3735 611 -3649 667
rect -3593 611 -3507 667
rect -3451 611 -3365 667
rect -3309 611 -3223 667
rect -3167 611 -3081 667
rect -3025 611 -2939 667
rect -2883 611 -2797 667
rect -2741 611 -2655 667
rect -2599 611 -2513 667
rect -2457 611 -2371 667
rect -2315 611 -2229 667
rect -2173 611 -2087 667
rect -2031 611 -1945 667
rect -1889 611 -1803 667
rect -1747 611 -1661 667
rect -1605 611 -1519 667
rect -1463 611 -1377 667
rect -1321 611 -1235 667
rect -1179 611 -1093 667
rect -1037 611 -951 667
rect -895 611 -809 667
rect -753 611 -667 667
rect -611 611 -525 667
rect -469 611 -383 667
rect -327 611 -241 667
rect -185 611 -99 667
rect -43 611 43 667
rect 99 611 185 667
rect 241 611 327 667
rect 383 611 469 667
rect 525 611 611 667
rect 667 611 753 667
rect 809 611 895 667
rect 951 611 1037 667
rect 1093 611 1179 667
rect 1235 611 1321 667
rect 1377 611 1463 667
rect 1519 611 1605 667
rect 1661 611 1747 667
rect 1803 611 1889 667
rect 1945 611 2031 667
rect 2087 611 2173 667
rect 2229 611 2315 667
rect 2371 611 2457 667
rect 2513 611 2599 667
rect 2655 611 2741 667
rect 2797 611 2883 667
rect 2939 611 3025 667
rect 3081 611 3167 667
rect 3223 611 3309 667
rect 3365 611 3451 667
rect 3507 611 3593 667
rect 3649 611 3735 667
rect 3791 611 3877 667
rect 3933 611 4019 667
rect 4075 611 4161 667
rect 4217 611 4303 667
rect 4359 611 4445 667
rect 4501 611 4587 667
rect 4643 611 4729 667
rect 4785 611 4871 667
rect 4927 611 5013 667
rect 5069 611 5155 667
rect 5211 611 5297 667
rect 5353 611 5439 667
rect 5495 611 5581 667
rect 5637 611 5723 667
rect 5779 611 5865 667
rect 5921 611 6007 667
rect 6063 611 6149 667
rect 6205 611 6291 667
rect 6347 611 6433 667
rect 6489 611 6575 667
rect 6631 611 6717 667
rect 6773 611 6859 667
rect 6915 611 7001 667
rect 7057 611 7143 667
rect 7199 611 7285 667
rect 7341 611 7351 667
rect -7351 525 7351 611
rect -7351 469 -7341 525
rect -7285 469 -7199 525
rect -7143 469 -7057 525
rect -7001 469 -6915 525
rect -6859 469 -6773 525
rect -6717 469 -6631 525
rect -6575 469 -6489 525
rect -6433 469 -6347 525
rect -6291 469 -6205 525
rect -6149 469 -6063 525
rect -6007 469 -5921 525
rect -5865 469 -5779 525
rect -5723 469 -5637 525
rect -5581 469 -5495 525
rect -5439 469 -5353 525
rect -5297 469 -5211 525
rect -5155 469 -5069 525
rect -5013 469 -4927 525
rect -4871 469 -4785 525
rect -4729 469 -4643 525
rect -4587 469 -4501 525
rect -4445 469 -4359 525
rect -4303 469 -4217 525
rect -4161 469 -4075 525
rect -4019 469 -3933 525
rect -3877 469 -3791 525
rect -3735 469 -3649 525
rect -3593 469 -3507 525
rect -3451 469 -3365 525
rect -3309 469 -3223 525
rect -3167 469 -3081 525
rect -3025 469 -2939 525
rect -2883 469 -2797 525
rect -2741 469 -2655 525
rect -2599 469 -2513 525
rect -2457 469 -2371 525
rect -2315 469 -2229 525
rect -2173 469 -2087 525
rect -2031 469 -1945 525
rect -1889 469 -1803 525
rect -1747 469 -1661 525
rect -1605 469 -1519 525
rect -1463 469 -1377 525
rect -1321 469 -1235 525
rect -1179 469 -1093 525
rect -1037 469 -951 525
rect -895 469 -809 525
rect -753 469 -667 525
rect -611 469 -525 525
rect -469 469 -383 525
rect -327 469 -241 525
rect -185 469 -99 525
rect -43 469 43 525
rect 99 469 185 525
rect 241 469 327 525
rect 383 469 469 525
rect 525 469 611 525
rect 667 469 753 525
rect 809 469 895 525
rect 951 469 1037 525
rect 1093 469 1179 525
rect 1235 469 1321 525
rect 1377 469 1463 525
rect 1519 469 1605 525
rect 1661 469 1747 525
rect 1803 469 1889 525
rect 1945 469 2031 525
rect 2087 469 2173 525
rect 2229 469 2315 525
rect 2371 469 2457 525
rect 2513 469 2599 525
rect 2655 469 2741 525
rect 2797 469 2883 525
rect 2939 469 3025 525
rect 3081 469 3167 525
rect 3223 469 3309 525
rect 3365 469 3451 525
rect 3507 469 3593 525
rect 3649 469 3735 525
rect 3791 469 3877 525
rect 3933 469 4019 525
rect 4075 469 4161 525
rect 4217 469 4303 525
rect 4359 469 4445 525
rect 4501 469 4587 525
rect 4643 469 4729 525
rect 4785 469 4871 525
rect 4927 469 5013 525
rect 5069 469 5155 525
rect 5211 469 5297 525
rect 5353 469 5439 525
rect 5495 469 5581 525
rect 5637 469 5723 525
rect 5779 469 5865 525
rect 5921 469 6007 525
rect 6063 469 6149 525
rect 6205 469 6291 525
rect 6347 469 6433 525
rect 6489 469 6575 525
rect 6631 469 6717 525
rect 6773 469 6859 525
rect 6915 469 7001 525
rect 7057 469 7143 525
rect 7199 469 7285 525
rect 7341 469 7351 525
rect -7351 383 7351 469
rect -7351 327 -7341 383
rect -7285 327 -7199 383
rect -7143 327 -7057 383
rect -7001 327 -6915 383
rect -6859 327 -6773 383
rect -6717 327 -6631 383
rect -6575 327 -6489 383
rect -6433 327 -6347 383
rect -6291 327 -6205 383
rect -6149 327 -6063 383
rect -6007 327 -5921 383
rect -5865 327 -5779 383
rect -5723 327 -5637 383
rect -5581 327 -5495 383
rect -5439 327 -5353 383
rect -5297 327 -5211 383
rect -5155 327 -5069 383
rect -5013 327 -4927 383
rect -4871 327 -4785 383
rect -4729 327 -4643 383
rect -4587 327 -4501 383
rect -4445 327 -4359 383
rect -4303 327 -4217 383
rect -4161 327 -4075 383
rect -4019 327 -3933 383
rect -3877 327 -3791 383
rect -3735 327 -3649 383
rect -3593 327 -3507 383
rect -3451 327 -3365 383
rect -3309 327 -3223 383
rect -3167 327 -3081 383
rect -3025 327 -2939 383
rect -2883 327 -2797 383
rect -2741 327 -2655 383
rect -2599 327 -2513 383
rect -2457 327 -2371 383
rect -2315 327 -2229 383
rect -2173 327 -2087 383
rect -2031 327 -1945 383
rect -1889 327 -1803 383
rect -1747 327 -1661 383
rect -1605 327 -1519 383
rect -1463 327 -1377 383
rect -1321 327 -1235 383
rect -1179 327 -1093 383
rect -1037 327 -951 383
rect -895 327 -809 383
rect -753 327 -667 383
rect -611 327 -525 383
rect -469 327 -383 383
rect -327 327 -241 383
rect -185 327 -99 383
rect -43 327 43 383
rect 99 327 185 383
rect 241 327 327 383
rect 383 327 469 383
rect 525 327 611 383
rect 667 327 753 383
rect 809 327 895 383
rect 951 327 1037 383
rect 1093 327 1179 383
rect 1235 327 1321 383
rect 1377 327 1463 383
rect 1519 327 1605 383
rect 1661 327 1747 383
rect 1803 327 1889 383
rect 1945 327 2031 383
rect 2087 327 2173 383
rect 2229 327 2315 383
rect 2371 327 2457 383
rect 2513 327 2599 383
rect 2655 327 2741 383
rect 2797 327 2883 383
rect 2939 327 3025 383
rect 3081 327 3167 383
rect 3223 327 3309 383
rect 3365 327 3451 383
rect 3507 327 3593 383
rect 3649 327 3735 383
rect 3791 327 3877 383
rect 3933 327 4019 383
rect 4075 327 4161 383
rect 4217 327 4303 383
rect 4359 327 4445 383
rect 4501 327 4587 383
rect 4643 327 4729 383
rect 4785 327 4871 383
rect 4927 327 5013 383
rect 5069 327 5155 383
rect 5211 327 5297 383
rect 5353 327 5439 383
rect 5495 327 5581 383
rect 5637 327 5723 383
rect 5779 327 5865 383
rect 5921 327 6007 383
rect 6063 327 6149 383
rect 6205 327 6291 383
rect 6347 327 6433 383
rect 6489 327 6575 383
rect 6631 327 6717 383
rect 6773 327 6859 383
rect 6915 327 7001 383
rect 7057 327 7143 383
rect 7199 327 7285 383
rect 7341 327 7351 383
rect -7351 241 7351 327
rect -7351 185 -7341 241
rect -7285 185 -7199 241
rect -7143 185 -7057 241
rect -7001 185 -6915 241
rect -6859 185 -6773 241
rect -6717 185 -6631 241
rect -6575 185 -6489 241
rect -6433 185 -6347 241
rect -6291 185 -6205 241
rect -6149 185 -6063 241
rect -6007 185 -5921 241
rect -5865 185 -5779 241
rect -5723 185 -5637 241
rect -5581 185 -5495 241
rect -5439 185 -5353 241
rect -5297 185 -5211 241
rect -5155 185 -5069 241
rect -5013 185 -4927 241
rect -4871 185 -4785 241
rect -4729 185 -4643 241
rect -4587 185 -4501 241
rect -4445 185 -4359 241
rect -4303 185 -4217 241
rect -4161 185 -4075 241
rect -4019 185 -3933 241
rect -3877 185 -3791 241
rect -3735 185 -3649 241
rect -3593 185 -3507 241
rect -3451 185 -3365 241
rect -3309 185 -3223 241
rect -3167 185 -3081 241
rect -3025 185 -2939 241
rect -2883 185 -2797 241
rect -2741 185 -2655 241
rect -2599 185 -2513 241
rect -2457 185 -2371 241
rect -2315 185 -2229 241
rect -2173 185 -2087 241
rect -2031 185 -1945 241
rect -1889 185 -1803 241
rect -1747 185 -1661 241
rect -1605 185 -1519 241
rect -1463 185 -1377 241
rect -1321 185 -1235 241
rect -1179 185 -1093 241
rect -1037 185 -951 241
rect -895 185 -809 241
rect -753 185 -667 241
rect -611 185 -525 241
rect -469 185 -383 241
rect -327 185 -241 241
rect -185 185 -99 241
rect -43 185 43 241
rect 99 185 185 241
rect 241 185 327 241
rect 383 185 469 241
rect 525 185 611 241
rect 667 185 753 241
rect 809 185 895 241
rect 951 185 1037 241
rect 1093 185 1179 241
rect 1235 185 1321 241
rect 1377 185 1463 241
rect 1519 185 1605 241
rect 1661 185 1747 241
rect 1803 185 1889 241
rect 1945 185 2031 241
rect 2087 185 2173 241
rect 2229 185 2315 241
rect 2371 185 2457 241
rect 2513 185 2599 241
rect 2655 185 2741 241
rect 2797 185 2883 241
rect 2939 185 3025 241
rect 3081 185 3167 241
rect 3223 185 3309 241
rect 3365 185 3451 241
rect 3507 185 3593 241
rect 3649 185 3735 241
rect 3791 185 3877 241
rect 3933 185 4019 241
rect 4075 185 4161 241
rect 4217 185 4303 241
rect 4359 185 4445 241
rect 4501 185 4587 241
rect 4643 185 4729 241
rect 4785 185 4871 241
rect 4927 185 5013 241
rect 5069 185 5155 241
rect 5211 185 5297 241
rect 5353 185 5439 241
rect 5495 185 5581 241
rect 5637 185 5723 241
rect 5779 185 5865 241
rect 5921 185 6007 241
rect 6063 185 6149 241
rect 6205 185 6291 241
rect 6347 185 6433 241
rect 6489 185 6575 241
rect 6631 185 6717 241
rect 6773 185 6859 241
rect 6915 185 7001 241
rect 7057 185 7143 241
rect 7199 185 7285 241
rect 7341 185 7351 241
rect -7351 99 7351 185
rect -7351 43 -7341 99
rect -7285 43 -7199 99
rect -7143 43 -7057 99
rect -7001 43 -6915 99
rect -6859 43 -6773 99
rect -6717 43 -6631 99
rect -6575 43 -6489 99
rect -6433 43 -6347 99
rect -6291 43 -6205 99
rect -6149 43 -6063 99
rect -6007 43 -5921 99
rect -5865 43 -5779 99
rect -5723 43 -5637 99
rect -5581 43 -5495 99
rect -5439 43 -5353 99
rect -5297 43 -5211 99
rect -5155 43 -5069 99
rect -5013 43 -4927 99
rect -4871 43 -4785 99
rect -4729 43 -4643 99
rect -4587 43 -4501 99
rect -4445 43 -4359 99
rect -4303 43 -4217 99
rect -4161 43 -4075 99
rect -4019 43 -3933 99
rect -3877 43 -3791 99
rect -3735 43 -3649 99
rect -3593 43 -3507 99
rect -3451 43 -3365 99
rect -3309 43 -3223 99
rect -3167 43 -3081 99
rect -3025 43 -2939 99
rect -2883 43 -2797 99
rect -2741 43 -2655 99
rect -2599 43 -2513 99
rect -2457 43 -2371 99
rect -2315 43 -2229 99
rect -2173 43 -2087 99
rect -2031 43 -1945 99
rect -1889 43 -1803 99
rect -1747 43 -1661 99
rect -1605 43 -1519 99
rect -1463 43 -1377 99
rect -1321 43 -1235 99
rect -1179 43 -1093 99
rect -1037 43 -951 99
rect -895 43 -809 99
rect -753 43 -667 99
rect -611 43 -525 99
rect -469 43 -383 99
rect -327 43 -241 99
rect -185 43 -99 99
rect -43 43 43 99
rect 99 43 185 99
rect 241 43 327 99
rect 383 43 469 99
rect 525 43 611 99
rect 667 43 753 99
rect 809 43 895 99
rect 951 43 1037 99
rect 1093 43 1179 99
rect 1235 43 1321 99
rect 1377 43 1463 99
rect 1519 43 1605 99
rect 1661 43 1747 99
rect 1803 43 1889 99
rect 1945 43 2031 99
rect 2087 43 2173 99
rect 2229 43 2315 99
rect 2371 43 2457 99
rect 2513 43 2599 99
rect 2655 43 2741 99
rect 2797 43 2883 99
rect 2939 43 3025 99
rect 3081 43 3167 99
rect 3223 43 3309 99
rect 3365 43 3451 99
rect 3507 43 3593 99
rect 3649 43 3735 99
rect 3791 43 3877 99
rect 3933 43 4019 99
rect 4075 43 4161 99
rect 4217 43 4303 99
rect 4359 43 4445 99
rect 4501 43 4587 99
rect 4643 43 4729 99
rect 4785 43 4871 99
rect 4927 43 5013 99
rect 5069 43 5155 99
rect 5211 43 5297 99
rect 5353 43 5439 99
rect 5495 43 5581 99
rect 5637 43 5723 99
rect 5779 43 5865 99
rect 5921 43 6007 99
rect 6063 43 6149 99
rect 6205 43 6291 99
rect 6347 43 6433 99
rect 6489 43 6575 99
rect 6631 43 6717 99
rect 6773 43 6859 99
rect 6915 43 7001 99
rect 7057 43 7143 99
rect 7199 43 7285 99
rect 7341 43 7351 99
rect -7351 -43 7351 43
rect -7351 -99 -7341 -43
rect -7285 -99 -7199 -43
rect -7143 -99 -7057 -43
rect -7001 -99 -6915 -43
rect -6859 -99 -6773 -43
rect -6717 -99 -6631 -43
rect -6575 -99 -6489 -43
rect -6433 -99 -6347 -43
rect -6291 -99 -6205 -43
rect -6149 -99 -6063 -43
rect -6007 -99 -5921 -43
rect -5865 -99 -5779 -43
rect -5723 -99 -5637 -43
rect -5581 -99 -5495 -43
rect -5439 -99 -5353 -43
rect -5297 -99 -5211 -43
rect -5155 -99 -5069 -43
rect -5013 -99 -4927 -43
rect -4871 -99 -4785 -43
rect -4729 -99 -4643 -43
rect -4587 -99 -4501 -43
rect -4445 -99 -4359 -43
rect -4303 -99 -4217 -43
rect -4161 -99 -4075 -43
rect -4019 -99 -3933 -43
rect -3877 -99 -3791 -43
rect -3735 -99 -3649 -43
rect -3593 -99 -3507 -43
rect -3451 -99 -3365 -43
rect -3309 -99 -3223 -43
rect -3167 -99 -3081 -43
rect -3025 -99 -2939 -43
rect -2883 -99 -2797 -43
rect -2741 -99 -2655 -43
rect -2599 -99 -2513 -43
rect -2457 -99 -2371 -43
rect -2315 -99 -2229 -43
rect -2173 -99 -2087 -43
rect -2031 -99 -1945 -43
rect -1889 -99 -1803 -43
rect -1747 -99 -1661 -43
rect -1605 -99 -1519 -43
rect -1463 -99 -1377 -43
rect -1321 -99 -1235 -43
rect -1179 -99 -1093 -43
rect -1037 -99 -951 -43
rect -895 -99 -809 -43
rect -753 -99 -667 -43
rect -611 -99 -525 -43
rect -469 -99 -383 -43
rect -327 -99 -241 -43
rect -185 -99 -99 -43
rect -43 -99 43 -43
rect 99 -99 185 -43
rect 241 -99 327 -43
rect 383 -99 469 -43
rect 525 -99 611 -43
rect 667 -99 753 -43
rect 809 -99 895 -43
rect 951 -99 1037 -43
rect 1093 -99 1179 -43
rect 1235 -99 1321 -43
rect 1377 -99 1463 -43
rect 1519 -99 1605 -43
rect 1661 -99 1747 -43
rect 1803 -99 1889 -43
rect 1945 -99 2031 -43
rect 2087 -99 2173 -43
rect 2229 -99 2315 -43
rect 2371 -99 2457 -43
rect 2513 -99 2599 -43
rect 2655 -99 2741 -43
rect 2797 -99 2883 -43
rect 2939 -99 3025 -43
rect 3081 -99 3167 -43
rect 3223 -99 3309 -43
rect 3365 -99 3451 -43
rect 3507 -99 3593 -43
rect 3649 -99 3735 -43
rect 3791 -99 3877 -43
rect 3933 -99 4019 -43
rect 4075 -99 4161 -43
rect 4217 -99 4303 -43
rect 4359 -99 4445 -43
rect 4501 -99 4587 -43
rect 4643 -99 4729 -43
rect 4785 -99 4871 -43
rect 4927 -99 5013 -43
rect 5069 -99 5155 -43
rect 5211 -99 5297 -43
rect 5353 -99 5439 -43
rect 5495 -99 5581 -43
rect 5637 -99 5723 -43
rect 5779 -99 5865 -43
rect 5921 -99 6007 -43
rect 6063 -99 6149 -43
rect 6205 -99 6291 -43
rect 6347 -99 6433 -43
rect 6489 -99 6575 -43
rect 6631 -99 6717 -43
rect 6773 -99 6859 -43
rect 6915 -99 7001 -43
rect 7057 -99 7143 -43
rect 7199 -99 7285 -43
rect 7341 -99 7351 -43
rect -7351 -185 7351 -99
rect -7351 -241 -7341 -185
rect -7285 -241 -7199 -185
rect -7143 -241 -7057 -185
rect -7001 -241 -6915 -185
rect -6859 -241 -6773 -185
rect -6717 -241 -6631 -185
rect -6575 -241 -6489 -185
rect -6433 -241 -6347 -185
rect -6291 -241 -6205 -185
rect -6149 -241 -6063 -185
rect -6007 -241 -5921 -185
rect -5865 -241 -5779 -185
rect -5723 -241 -5637 -185
rect -5581 -241 -5495 -185
rect -5439 -241 -5353 -185
rect -5297 -241 -5211 -185
rect -5155 -241 -5069 -185
rect -5013 -241 -4927 -185
rect -4871 -241 -4785 -185
rect -4729 -241 -4643 -185
rect -4587 -241 -4501 -185
rect -4445 -241 -4359 -185
rect -4303 -241 -4217 -185
rect -4161 -241 -4075 -185
rect -4019 -241 -3933 -185
rect -3877 -241 -3791 -185
rect -3735 -241 -3649 -185
rect -3593 -241 -3507 -185
rect -3451 -241 -3365 -185
rect -3309 -241 -3223 -185
rect -3167 -241 -3081 -185
rect -3025 -241 -2939 -185
rect -2883 -241 -2797 -185
rect -2741 -241 -2655 -185
rect -2599 -241 -2513 -185
rect -2457 -241 -2371 -185
rect -2315 -241 -2229 -185
rect -2173 -241 -2087 -185
rect -2031 -241 -1945 -185
rect -1889 -241 -1803 -185
rect -1747 -241 -1661 -185
rect -1605 -241 -1519 -185
rect -1463 -241 -1377 -185
rect -1321 -241 -1235 -185
rect -1179 -241 -1093 -185
rect -1037 -241 -951 -185
rect -895 -241 -809 -185
rect -753 -241 -667 -185
rect -611 -241 -525 -185
rect -469 -241 -383 -185
rect -327 -241 -241 -185
rect -185 -241 -99 -185
rect -43 -241 43 -185
rect 99 -241 185 -185
rect 241 -241 327 -185
rect 383 -241 469 -185
rect 525 -241 611 -185
rect 667 -241 753 -185
rect 809 -241 895 -185
rect 951 -241 1037 -185
rect 1093 -241 1179 -185
rect 1235 -241 1321 -185
rect 1377 -241 1463 -185
rect 1519 -241 1605 -185
rect 1661 -241 1747 -185
rect 1803 -241 1889 -185
rect 1945 -241 2031 -185
rect 2087 -241 2173 -185
rect 2229 -241 2315 -185
rect 2371 -241 2457 -185
rect 2513 -241 2599 -185
rect 2655 -241 2741 -185
rect 2797 -241 2883 -185
rect 2939 -241 3025 -185
rect 3081 -241 3167 -185
rect 3223 -241 3309 -185
rect 3365 -241 3451 -185
rect 3507 -241 3593 -185
rect 3649 -241 3735 -185
rect 3791 -241 3877 -185
rect 3933 -241 4019 -185
rect 4075 -241 4161 -185
rect 4217 -241 4303 -185
rect 4359 -241 4445 -185
rect 4501 -241 4587 -185
rect 4643 -241 4729 -185
rect 4785 -241 4871 -185
rect 4927 -241 5013 -185
rect 5069 -241 5155 -185
rect 5211 -241 5297 -185
rect 5353 -241 5439 -185
rect 5495 -241 5581 -185
rect 5637 -241 5723 -185
rect 5779 -241 5865 -185
rect 5921 -241 6007 -185
rect 6063 -241 6149 -185
rect 6205 -241 6291 -185
rect 6347 -241 6433 -185
rect 6489 -241 6575 -185
rect 6631 -241 6717 -185
rect 6773 -241 6859 -185
rect 6915 -241 7001 -185
rect 7057 -241 7143 -185
rect 7199 -241 7285 -185
rect 7341 -241 7351 -185
rect -7351 -327 7351 -241
rect -7351 -383 -7341 -327
rect -7285 -383 -7199 -327
rect -7143 -383 -7057 -327
rect -7001 -383 -6915 -327
rect -6859 -383 -6773 -327
rect -6717 -383 -6631 -327
rect -6575 -383 -6489 -327
rect -6433 -383 -6347 -327
rect -6291 -383 -6205 -327
rect -6149 -383 -6063 -327
rect -6007 -383 -5921 -327
rect -5865 -383 -5779 -327
rect -5723 -383 -5637 -327
rect -5581 -383 -5495 -327
rect -5439 -383 -5353 -327
rect -5297 -383 -5211 -327
rect -5155 -383 -5069 -327
rect -5013 -383 -4927 -327
rect -4871 -383 -4785 -327
rect -4729 -383 -4643 -327
rect -4587 -383 -4501 -327
rect -4445 -383 -4359 -327
rect -4303 -383 -4217 -327
rect -4161 -383 -4075 -327
rect -4019 -383 -3933 -327
rect -3877 -383 -3791 -327
rect -3735 -383 -3649 -327
rect -3593 -383 -3507 -327
rect -3451 -383 -3365 -327
rect -3309 -383 -3223 -327
rect -3167 -383 -3081 -327
rect -3025 -383 -2939 -327
rect -2883 -383 -2797 -327
rect -2741 -383 -2655 -327
rect -2599 -383 -2513 -327
rect -2457 -383 -2371 -327
rect -2315 -383 -2229 -327
rect -2173 -383 -2087 -327
rect -2031 -383 -1945 -327
rect -1889 -383 -1803 -327
rect -1747 -383 -1661 -327
rect -1605 -383 -1519 -327
rect -1463 -383 -1377 -327
rect -1321 -383 -1235 -327
rect -1179 -383 -1093 -327
rect -1037 -383 -951 -327
rect -895 -383 -809 -327
rect -753 -383 -667 -327
rect -611 -383 -525 -327
rect -469 -383 -383 -327
rect -327 -383 -241 -327
rect -185 -383 -99 -327
rect -43 -383 43 -327
rect 99 -383 185 -327
rect 241 -383 327 -327
rect 383 -383 469 -327
rect 525 -383 611 -327
rect 667 -383 753 -327
rect 809 -383 895 -327
rect 951 -383 1037 -327
rect 1093 -383 1179 -327
rect 1235 -383 1321 -327
rect 1377 -383 1463 -327
rect 1519 -383 1605 -327
rect 1661 -383 1747 -327
rect 1803 -383 1889 -327
rect 1945 -383 2031 -327
rect 2087 -383 2173 -327
rect 2229 -383 2315 -327
rect 2371 -383 2457 -327
rect 2513 -383 2599 -327
rect 2655 -383 2741 -327
rect 2797 -383 2883 -327
rect 2939 -383 3025 -327
rect 3081 -383 3167 -327
rect 3223 -383 3309 -327
rect 3365 -383 3451 -327
rect 3507 -383 3593 -327
rect 3649 -383 3735 -327
rect 3791 -383 3877 -327
rect 3933 -383 4019 -327
rect 4075 -383 4161 -327
rect 4217 -383 4303 -327
rect 4359 -383 4445 -327
rect 4501 -383 4587 -327
rect 4643 -383 4729 -327
rect 4785 -383 4871 -327
rect 4927 -383 5013 -327
rect 5069 -383 5155 -327
rect 5211 -383 5297 -327
rect 5353 -383 5439 -327
rect 5495 -383 5581 -327
rect 5637 -383 5723 -327
rect 5779 -383 5865 -327
rect 5921 -383 6007 -327
rect 6063 -383 6149 -327
rect 6205 -383 6291 -327
rect 6347 -383 6433 -327
rect 6489 -383 6575 -327
rect 6631 -383 6717 -327
rect 6773 -383 6859 -327
rect 6915 -383 7001 -327
rect 7057 -383 7143 -327
rect 7199 -383 7285 -327
rect 7341 -383 7351 -327
rect -7351 -469 7351 -383
rect -7351 -525 -7341 -469
rect -7285 -525 -7199 -469
rect -7143 -525 -7057 -469
rect -7001 -525 -6915 -469
rect -6859 -525 -6773 -469
rect -6717 -525 -6631 -469
rect -6575 -525 -6489 -469
rect -6433 -525 -6347 -469
rect -6291 -525 -6205 -469
rect -6149 -525 -6063 -469
rect -6007 -525 -5921 -469
rect -5865 -525 -5779 -469
rect -5723 -525 -5637 -469
rect -5581 -525 -5495 -469
rect -5439 -525 -5353 -469
rect -5297 -525 -5211 -469
rect -5155 -525 -5069 -469
rect -5013 -525 -4927 -469
rect -4871 -525 -4785 -469
rect -4729 -525 -4643 -469
rect -4587 -525 -4501 -469
rect -4445 -525 -4359 -469
rect -4303 -525 -4217 -469
rect -4161 -525 -4075 -469
rect -4019 -525 -3933 -469
rect -3877 -525 -3791 -469
rect -3735 -525 -3649 -469
rect -3593 -525 -3507 -469
rect -3451 -525 -3365 -469
rect -3309 -525 -3223 -469
rect -3167 -525 -3081 -469
rect -3025 -525 -2939 -469
rect -2883 -525 -2797 -469
rect -2741 -525 -2655 -469
rect -2599 -525 -2513 -469
rect -2457 -525 -2371 -469
rect -2315 -525 -2229 -469
rect -2173 -525 -2087 -469
rect -2031 -525 -1945 -469
rect -1889 -525 -1803 -469
rect -1747 -525 -1661 -469
rect -1605 -525 -1519 -469
rect -1463 -525 -1377 -469
rect -1321 -525 -1235 -469
rect -1179 -525 -1093 -469
rect -1037 -525 -951 -469
rect -895 -525 -809 -469
rect -753 -525 -667 -469
rect -611 -525 -525 -469
rect -469 -525 -383 -469
rect -327 -525 -241 -469
rect -185 -525 -99 -469
rect -43 -525 43 -469
rect 99 -525 185 -469
rect 241 -525 327 -469
rect 383 -525 469 -469
rect 525 -525 611 -469
rect 667 -525 753 -469
rect 809 -525 895 -469
rect 951 -525 1037 -469
rect 1093 -525 1179 -469
rect 1235 -525 1321 -469
rect 1377 -525 1463 -469
rect 1519 -525 1605 -469
rect 1661 -525 1747 -469
rect 1803 -525 1889 -469
rect 1945 -525 2031 -469
rect 2087 -525 2173 -469
rect 2229 -525 2315 -469
rect 2371 -525 2457 -469
rect 2513 -525 2599 -469
rect 2655 -525 2741 -469
rect 2797 -525 2883 -469
rect 2939 -525 3025 -469
rect 3081 -525 3167 -469
rect 3223 -525 3309 -469
rect 3365 -525 3451 -469
rect 3507 -525 3593 -469
rect 3649 -525 3735 -469
rect 3791 -525 3877 -469
rect 3933 -525 4019 -469
rect 4075 -525 4161 -469
rect 4217 -525 4303 -469
rect 4359 -525 4445 -469
rect 4501 -525 4587 -469
rect 4643 -525 4729 -469
rect 4785 -525 4871 -469
rect 4927 -525 5013 -469
rect 5069 -525 5155 -469
rect 5211 -525 5297 -469
rect 5353 -525 5439 -469
rect 5495 -525 5581 -469
rect 5637 -525 5723 -469
rect 5779 -525 5865 -469
rect 5921 -525 6007 -469
rect 6063 -525 6149 -469
rect 6205 -525 6291 -469
rect 6347 -525 6433 -469
rect 6489 -525 6575 -469
rect 6631 -525 6717 -469
rect 6773 -525 6859 -469
rect 6915 -525 7001 -469
rect 7057 -525 7143 -469
rect 7199 -525 7285 -469
rect 7341 -525 7351 -469
rect -7351 -611 7351 -525
rect -7351 -667 -7341 -611
rect -7285 -667 -7199 -611
rect -7143 -667 -7057 -611
rect -7001 -667 -6915 -611
rect -6859 -667 -6773 -611
rect -6717 -667 -6631 -611
rect -6575 -667 -6489 -611
rect -6433 -667 -6347 -611
rect -6291 -667 -6205 -611
rect -6149 -667 -6063 -611
rect -6007 -667 -5921 -611
rect -5865 -667 -5779 -611
rect -5723 -667 -5637 -611
rect -5581 -667 -5495 -611
rect -5439 -667 -5353 -611
rect -5297 -667 -5211 -611
rect -5155 -667 -5069 -611
rect -5013 -667 -4927 -611
rect -4871 -667 -4785 -611
rect -4729 -667 -4643 -611
rect -4587 -667 -4501 -611
rect -4445 -667 -4359 -611
rect -4303 -667 -4217 -611
rect -4161 -667 -4075 -611
rect -4019 -667 -3933 -611
rect -3877 -667 -3791 -611
rect -3735 -667 -3649 -611
rect -3593 -667 -3507 -611
rect -3451 -667 -3365 -611
rect -3309 -667 -3223 -611
rect -3167 -667 -3081 -611
rect -3025 -667 -2939 -611
rect -2883 -667 -2797 -611
rect -2741 -667 -2655 -611
rect -2599 -667 -2513 -611
rect -2457 -667 -2371 -611
rect -2315 -667 -2229 -611
rect -2173 -667 -2087 -611
rect -2031 -667 -1945 -611
rect -1889 -667 -1803 -611
rect -1747 -667 -1661 -611
rect -1605 -667 -1519 -611
rect -1463 -667 -1377 -611
rect -1321 -667 -1235 -611
rect -1179 -667 -1093 -611
rect -1037 -667 -951 -611
rect -895 -667 -809 -611
rect -753 -667 -667 -611
rect -611 -667 -525 -611
rect -469 -667 -383 -611
rect -327 -667 -241 -611
rect -185 -667 -99 -611
rect -43 -667 43 -611
rect 99 -667 185 -611
rect 241 -667 327 -611
rect 383 -667 469 -611
rect 525 -667 611 -611
rect 667 -667 753 -611
rect 809 -667 895 -611
rect 951 -667 1037 -611
rect 1093 -667 1179 -611
rect 1235 -667 1321 -611
rect 1377 -667 1463 -611
rect 1519 -667 1605 -611
rect 1661 -667 1747 -611
rect 1803 -667 1889 -611
rect 1945 -667 2031 -611
rect 2087 -667 2173 -611
rect 2229 -667 2315 -611
rect 2371 -667 2457 -611
rect 2513 -667 2599 -611
rect 2655 -667 2741 -611
rect 2797 -667 2883 -611
rect 2939 -667 3025 -611
rect 3081 -667 3167 -611
rect 3223 -667 3309 -611
rect 3365 -667 3451 -611
rect 3507 -667 3593 -611
rect 3649 -667 3735 -611
rect 3791 -667 3877 -611
rect 3933 -667 4019 -611
rect 4075 -667 4161 -611
rect 4217 -667 4303 -611
rect 4359 -667 4445 -611
rect 4501 -667 4587 -611
rect 4643 -667 4729 -611
rect 4785 -667 4871 -611
rect 4927 -667 5013 -611
rect 5069 -667 5155 -611
rect 5211 -667 5297 -611
rect 5353 -667 5439 -611
rect 5495 -667 5581 -611
rect 5637 -667 5723 -611
rect 5779 -667 5865 -611
rect 5921 -667 6007 -611
rect 6063 -667 6149 -611
rect 6205 -667 6291 -611
rect 6347 -667 6433 -611
rect 6489 -667 6575 -611
rect 6631 -667 6717 -611
rect 6773 -667 6859 -611
rect 6915 -667 7001 -611
rect 7057 -667 7143 -611
rect 7199 -667 7285 -611
rect 7341 -667 7351 -611
rect -7351 -677 7351 -667
<< end >>
