magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect 11097 11097 73000 73000
use GF_NI_COR_BASE  GF_NI_COR_BASE_0
timestamp 1713338890
transform 1 0 12 0 1 0
box 13436 13361 70889 70890
use POWER_RAIL_COR  POWER_RAIL_COR_0
timestamp 1713338890
transform 1 0 0 0 1 0
box 13097 13097 71000 71000
<< labels >>
rlabel metal5 s 67482 70220 67482 70220 4 DVDD
port 1 nsew
rlabel metal5 s 70444 44321 70444 44321 4 DVDD
port 1 nsew
rlabel metal5 s 70444 53176 70444 53176 4 DVDD
port 1 nsew
rlabel metal5 s 70444 54611 70444 54611 4 DVDD
port 1 nsew
rlabel metal5 s 70444 56376 70444 56376 4 DVDD
port 1 nsew
rlabel metal5 s 70444 59576 70444 59576 4 DVDD
port 1 nsew
rlabel metal5 s 70444 67411 70444 67411 4 DVDD
port 1 nsew
rlabel metal5 s 44292 70220 44292 70220 4 DVDD
port 1 nsew
rlabel metal5 s 53064 70220 53064 70220 4 DVDD
port 1 nsew
rlabel metal5 s 54690 70220 54690 70220 4 DVDD
port 1 nsew
rlabel metal5 s 56327 70220 56327 70220 4 DVDD
port 1 nsew
rlabel metal5 s 59509 70220 59509 70220 4 DVDD
port 1 nsew
rlabel metal5 s 67482 70220 67482 70220 4 DVDD
port 1 nsew
rlabel metal5 s 70444 44321 70444 44321 4 DVDD
port 1 nsew
rlabel metal5 s 70444 53176 70444 53176 4 DVDD
port 1 nsew
rlabel metal5 s 70444 54611 70444 54611 4 DVDD
port 1 nsew
rlabel metal5 s 70444 56376 70444 56376 4 DVDD
port 1 nsew
rlabel metal5 s 70444 59576 70444 59576 4 DVDD
port 1 nsew
rlabel metal5 s 70444 67411 70444 67411 4 DVDD
port 1 nsew
rlabel metal5 s 44292 70220 44292 70220 4 DVDD
port 1 nsew
rlabel metal5 s 53064 70220 53064 70220 4 DVDD
port 1 nsew
rlabel metal5 s 54690 70220 54690 70220 4 DVDD
port 1 nsew
rlabel metal5 s 56327 70220 56327 70220 4 DVDD
port 1 nsew
rlabel metal5 s 59509 70220 59509 70220 4 DVDD
port 1 nsew
rlabel metal5 s 67482 70220 67482 70220 4 DVDD
port 1 nsew
rlabel metal5 s 70444 44321 70444 44321 4 DVDD
port 1 nsew
rlabel metal5 s 70444 53176 70444 53176 4 DVDD
port 1 nsew
rlabel metal5 s 70444 54611 70444 54611 4 DVDD
port 1 nsew
rlabel metal5 s 70444 56376 70444 56376 4 DVDD
port 1 nsew
rlabel metal5 s 70444 59576 70444 59576 4 DVDD
port 1 nsew
rlabel metal5 s 70444 67411 70444 67411 4 DVDD
port 1 nsew
rlabel metal5 s 44292 70220 44292 70220 4 DVDD
port 1 nsew
rlabel metal5 s 53064 70220 53064 70220 4 DVDD
port 1 nsew
rlabel metal5 s 54690 70220 54690 70220 4 DVDD
port 1 nsew
rlabel metal5 s 56327 70220 56327 70220 4 DVDD
port 1 nsew
rlabel metal5 s 59509 70220 59509 70220 4 DVDD
port 1 nsew
rlabel metal5 s 41877 70220 41877 70220 4 DVDD
port 1 nsew
rlabel metal5 s 37671 70220 37671 70220 4 DVDD
port 1 nsew
rlabel metal5 s 41877 70220 41877 70220 4 DVDD
port 1 nsew
rlabel metal5 s 23985 70220 23985 70220 4 DVDD
port 1 nsew
rlabel metal5 s 23985 70220 23985 70220 4 DVDD
port 1 nsew
rlabel metal5 s 28097 70220 28097 70220 4 DVDD
port 1 nsew
rlabel metal5 s 31313 70220 31313 70220 4 DVDD
port 1 nsew
rlabel metal5 s 34449 70220 34449 70220 4 DVDD
port 1 nsew
rlabel metal5 s 37671 70220 37671 70220 4 DVDD
port 1 nsew
rlabel metal5 s 41877 70220 41877 70220 4 DVDD
port 1 nsew
rlabel metal5 s 28097 70220 28097 70220 4 DVDD
port 1 nsew
rlabel metal5 s 31313 70220 31313 70220 4 DVDD
port 1 nsew
rlabel metal5 s 34449 70220 34449 70220 4 DVDD
port 1 nsew
rlabel metal5 s 23985 70220 23985 70220 4 DVDD
port 1 nsew
rlabel metal5 s 28097 70220 28097 70220 4 DVDD
port 1 nsew
rlabel metal5 s 31313 70220 31313 70220 4 DVDD
port 1 nsew
rlabel metal5 s 34449 70220 34449 70220 4 DVDD
port 1 nsew
rlabel metal5 s 37671 70220 37671 70220 4 DVDD
port 1 nsew
rlabel metal5 s 70444 37912 70444 37912 4 DVDD
port 1 nsew
rlabel metal5 s 70444 41930 70444 41930 4 DVDD
port 1 nsew
rlabel metal5 s 70444 31562 70444 31562 4 DVDD
port 1 nsew
rlabel metal5 s 70444 34676 70444 34676 4 DVDD
port 1 nsew
rlabel metal5 s 70444 37912 70444 37912 4 DVDD
port 1 nsew
rlabel metal5 s 70444 41930 70444 41930 4 DVDD
port 1 nsew
rlabel metal5 s 70444 34676 70444 34676 4 DVDD
port 1 nsew
rlabel metal5 s 70444 37912 70444 37912 4 DVDD
port 1 nsew
rlabel metal5 s 70444 41930 70444 41930 4 DVDD
port 1 nsew
rlabel metal5 s 70444 24237 70444 24237 4 DVDD
port 1 nsew
rlabel metal5 s 70444 28347 70444 28347 4 DVDD
port 1 nsew
rlabel metal5 s 70444 31562 70444 31562 4 DVDD
port 1 nsew
rlabel metal5 s 70444 24237 70444 24237 4 DVDD
port 1 nsew
rlabel metal5 s 70444 28347 70444 28347 4 DVDD
port 1 nsew
rlabel metal5 s 70444 24237 70444 24237 4 DVDD
port 1 nsew
rlabel metal5 s 70444 28347 70444 28347 4 DVDD
port 1 nsew
rlabel metal5 s 70444 31562 70444 31562 4 DVDD
port 1 nsew
rlabel metal5 s 70444 34676 70444 34676 4 DVDD
port 1 nsew
rlabel metal4 s 59509 70220 59509 70220 4 DVDD
port 1 nsew
rlabel metal4 s 56327 70220 56327 70220 4 DVDD
port 1 nsew
rlabel metal4 s 53064 70220 53064 70220 4 DVDD
port 1 nsew
rlabel metal4 s 44292 70220 44292 70220 4 DVDD
port 1 nsew
rlabel metal4 s 34449 70220 34449 70220 4 DVDD
port 1 nsew
rlabel metal4 s 28097 70220 28097 70220 4 DVDD
port 1 nsew
rlabel metal4 s 23985 70220 23985 70220 4 DVDD
port 1 nsew
rlabel metal4 s 70444 67411 70444 67411 4 DVDD
port 1 nsew
rlabel metal4 s 70444 59576 70444 59576 4 DVDD
port 1 nsew
rlabel metal4 s 70444 54611 70444 54611 4 DVDD
port 1 nsew
rlabel metal4 s 70444 44321 70444 44321 4 DVDD
port 1 nsew
rlabel metal4 s 70444 37912 70444 37912 4 DVDD
port 1 nsew
rlabel metal4 s 70444 31562 70444 31562 4 DVDD
port 1 nsew
rlabel metal4 s 70444 24237 70444 24237 4 DVDD
port 1 nsew
rlabel metal4 s 67482 70220 67482 70220 4 DVDD
port 1 nsew
rlabel metal4 s 54690 70220 54690 70220 4 DVDD
port 1 nsew
rlabel metal4 s 41877 70220 41877 70220 4 DVDD
port 1 nsew
rlabel metal4 s 37671 70220 37671 70220 4 DVDD
port 1 nsew
rlabel metal4 s 31313 70220 31313 70220 4 DVDD
port 1 nsew
rlabel metal4 s 70444 56376 70444 56376 4 DVDD
port 1 nsew
rlabel metal4 s 70444 53176 70444 53176 4 DVDD
port 1 nsew
rlabel metal4 s 70444 41930 70444 41930 4 DVDD
port 1 nsew
rlabel metal4 s 70444 34676 70444 34676 4 DVDD
port 1 nsew
rlabel metal4 s 70444 28347 70444 28347 4 DVDD
port 1 nsew
rlabel metal3 s 53064 70220 53064 70220 4 DVDD
port 1 nsew
rlabel metal3 s 44292 70220 44292 70220 4 DVDD
port 1 nsew
rlabel metal3 s 41877 70220 41877 70220 4 DVDD
port 1 nsew
rlabel metal3 s 37671 70220 37671 70220 4 DVDD
port 1 nsew
rlabel metal3 s 34449 70220 34449 70220 4 DVDD
port 1 nsew
rlabel metal3 s 31313 70220 31313 70220 4 DVDD
port 1 nsew
rlabel metal3 s 28097 70220 28097 70220 4 DVDD
port 1 nsew
rlabel metal3 s 70444 59576 70444 59576 4 DVDD
port 1 nsew
rlabel metal3 s 70444 56376 70444 56376 4 DVDD
port 1 nsew
rlabel metal3 s 70444 54611 70444 54611 4 DVDD
port 1 nsew
rlabel metal3 s 70444 53176 70444 53176 4 DVDD
port 1 nsew
rlabel metal3 s 70444 44321 70444 44321 4 DVDD
port 1 nsew
rlabel metal3 s 70444 41930 70444 41930 4 DVDD
port 1 nsew
rlabel metal3 s 70444 37912 70444 37912 4 DVDD
port 1 nsew
rlabel metal3 s 70444 34676 70444 34676 4 DVDD
port 1 nsew
rlabel metal3 s 70444 31562 70444 31562 4 DVDD
port 1 nsew
rlabel metal3 s 70444 28347 70444 28347 4 DVDD
port 1 nsew
rlabel metal3 s 70444 24237 70444 24237 4 DVDD
port 1 nsew
rlabel metal3 s 56327 70220 56327 70220 4 DVDD
port 1 nsew
rlabel metal3 s 70444 67411 70444 67411 4 DVDD
port 1 nsew
rlabel metal3 s 23985 70220 23985 70220 4 DVDD
port 1 nsew
rlabel metal3 s 59509 70220 59509 70220 4 DVDD
port 1 nsew
rlabel metal3 s 67482 70220 67482 70220 4 DVDD
port 1 nsew
rlabel metal3 s 54690 70220 54690 70220 4 DVDD
port 1 nsew
rlabel metal5 s 69026 70220 69026 70220 4 DVSS
port 2 nsew
rlabel metal5 s 70444 47548 70444 47548 4 DVSS
port 2 nsew
rlabel metal5 s 70444 57811 70444 57811 4 DVSS
port 2 nsew
rlabel metal5 s 70444 61011 70444 61011 4 DVSS
port 2 nsew
rlabel metal5 s 70444 65976 70444 65976 4 DVSS
port 2 nsew
rlabel metal5 s 70444 69002 70444 69002 4 DVSS
port 2 nsew
rlabel metal5 s 47523 70220 47523 70220 4 DVSS
port 2 nsew
rlabel metal5 s 57931 70220 57931 70220 4 DVSS
port 2 nsew
rlabel metal5 s 61124 70220 61124 70220 4 DVSS
port 2 nsew
rlabel metal5 s 65891 70220 65891 70220 4 DVSS
port 2 nsew
rlabel metal5 s 69026 70220 69026 70220 4 DVSS
port 2 nsew
rlabel metal5 s 70444 47548 70444 47548 4 DVSS
port 2 nsew
rlabel metal5 s 70444 57811 70444 57811 4 DVSS
port 2 nsew
rlabel metal5 s 70444 61011 70444 61011 4 DVSS
port 2 nsew
rlabel metal5 s 70444 65976 70444 65976 4 DVSS
port 2 nsew
rlabel metal5 s 70444 69002 70444 69002 4 DVSS
port 2 nsew
rlabel metal5 s 47523 70220 47523 70220 4 DVSS
port 2 nsew
rlabel metal5 s 57931 70220 57931 70220 4 DVSS
port 2 nsew
rlabel metal5 s 61124 70220 61124 70220 4 DVSS
port 2 nsew
rlabel metal5 s 65891 70220 65891 70220 4 DVSS
port 2 nsew
rlabel metal5 s 69026 70220 69026 70220 4 DVSS
port 2 nsew
rlabel metal5 s 70444 47548 70444 47548 4 DVSS
port 2 nsew
rlabel metal5 s 70444 57811 70444 57811 4 DVSS
port 2 nsew
rlabel metal5 s 70444 61011 70444 61011 4 DVSS
port 2 nsew
rlabel metal5 s 70444 65976 70444 65976 4 DVSS
port 2 nsew
rlabel metal5 s 70444 69002 70444 69002 4 DVSS
port 2 nsew
rlabel metal5 s 47523 70220 47523 70220 4 DVSS
port 2 nsew
rlabel metal5 s 57931 70220 57931 70220 4 DVSS
port 2 nsew
rlabel metal5 s 61124 70220 61124 70220 4 DVSS
port 2 nsew
rlabel metal5 s 65891 70220 65891 70220 4 DVSS
port 2 nsew
rlabel metal5 s 40319 70220 40319 70220 4 DVSS
port 2 nsew
rlabel metal5 s 40319 70220 40319 70220 4 DVSS
port 2 nsew
rlabel metal5 s 15448 70196 15448 70196 4 DVSS
port 2 nsew
rlabel metal5 s 18634 70150 18634 70150 4 DVSS
port 2 nsew
rlabel metal5 s 21613 70220 21613 70220 4 DVSS
port 2 nsew
rlabel metal5 s 15448 70196 15448 70196 4 DVSS
port 2 nsew
rlabel metal5 s 18634 70150 18634 70150 4 DVSS
port 2 nsew
rlabel metal5 s 21613 70220 21613 70220 4 DVSS
port 2 nsew
rlabel metal5 s 25800 70220 25800 70220 4 DVSS
port 2 nsew
rlabel metal5 s 40319 70220 40319 70220 4 DVSS
port 2 nsew
rlabel metal5 s 25800 70220 25800 70220 4 DVSS
port 2 nsew
rlabel metal5 s 15448 70196 15448 70196 4 DVSS
port 2 nsew
rlabel metal5 s 18634 70150 18634 70150 4 DVSS
port 2 nsew
rlabel metal5 s 21613 70220 21613 70220 4 DVSS
port 2 nsew
rlabel metal5 s 25800 70220 25800 70220 4 DVSS
port 2 nsew
rlabel metal5 s 70375 18874 70375 18874 4 DVSS
port 2 nsew
rlabel metal5 s 70422 15703 70422 15703 4 DVSS
port 2 nsew
rlabel metal5 s 70444 21860 70444 21860 4 DVSS
port 2 nsew
rlabel metal5 s 70444 21860 70444 21860 4 DVSS
port 2 nsew
rlabel metal5 s 70444 26053 70444 26053 4 DVSS
port 2 nsew
rlabel metal5 s 70444 40295 70444 40295 4 DVSS
port 2 nsew
rlabel metal5 s 70444 26053 70444 26053 4 DVSS
port 2 nsew
rlabel metal5 s 70444 40295 70444 40295 4 DVSS
port 2 nsew
rlabel metal5 s 70422 15703 70422 15703 4 DVSS
port 2 nsew
rlabel metal5 s 70375 18874 70375 18874 4 DVSS
port 2 nsew
rlabel metal5 s 70375 18874 70375 18874 4 DVSS
port 2 nsew
rlabel metal5 s 70422 15703 70422 15703 4 DVSS
port 2 nsew
rlabel metal5 s 70444 21860 70444 21860 4 DVSS
port 2 nsew
rlabel metal5 s 70444 26053 70444 26053 4 DVSS
port 2 nsew
rlabel metal5 s 70444 40295 70444 40295 4 DVSS
port 2 nsew
rlabel metal4 s 69026 70220 69026 70220 4 DVSS
port 2 nsew
rlabel metal4 s 65891 70220 65891 70220 4 DVSS
port 2 nsew
rlabel metal4 s 40319 70220 40319 70220 4 DVSS
port 2 nsew
rlabel metal4 s 18634 70150 18634 70150 4 DVSS
port 2 nsew
rlabel metal4 s 70444 69002 70444 69002 4 DVSS
port 2 nsew
rlabel metal4 s 70444 61011 70444 61011 4 DVSS
port 2 nsew
rlabel metal4 s 70444 47548 70444 47548 4 DVSS
port 2 nsew
rlabel metal4 s 70444 26053 70444 26053 4 DVSS
port 2 nsew
rlabel metal4 s 70422 15703 70422 15703 4 DVSS
port 2 nsew
rlabel metal4 s 61124 70220 61124 70220 4 DVSS
port 2 nsew
rlabel metal4 s 57931 70220 57931 70220 4 DVSS
port 2 nsew
rlabel metal4 s 47523 70220 47523 70220 4 DVSS
port 2 nsew
rlabel metal4 s 25800 70220 25800 70220 4 DVSS
port 2 nsew
rlabel metal4 s 21613 70220 21613 70220 4 DVSS
port 2 nsew
rlabel metal4 s 15448 70196 15448 70196 4 DVSS
port 2 nsew
rlabel metal4 s 70444 65976 70444 65976 4 DVSS
port 2 nsew
rlabel metal4 s 70444 57811 70444 57811 4 DVSS
port 2 nsew
rlabel metal4 s 70444 40295 70444 40295 4 DVSS
port 2 nsew
rlabel metal4 s 70444 21860 70444 21860 4 DVSS
port 2 nsew
rlabel metal4 s 70375 18874 70375 18874 4 DVSS
port 2 nsew
rlabel metal3 s 40319 70220 40319 70220 4 DVSS
port 2 nsew
rlabel metal3 s 57931 70220 57931 70220 4 DVSS
port 2 nsew
rlabel metal3 s 70444 69002 70444 69002 4 DVSS
port 2 nsew
rlabel metal3 s 47523 70220 47523 70220 4 DVSS
port 2 nsew
rlabel metal3 s 15448 70196 15448 70196 4 DVSS
port 2 nsew
rlabel metal3 s 18634 70150 18634 70150 4 DVSS
port 2 nsew
rlabel metal3 s 21613 70220 21613 70220 4 DVSS
port 2 nsew
rlabel metal3 s 25800 70220 25800 70220 4 DVSS
port 2 nsew
rlabel metal3 s 61124 70220 61124 70220 4 DVSS
port 2 nsew
rlabel metal3 s 65891 70220 65891 70220 4 DVSS
port 2 nsew
rlabel metal3 s 69026 70220 69026 70220 4 DVSS
port 2 nsew
rlabel metal3 s 70375 18874 70375 18874 4 DVSS
port 2 nsew
rlabel metal3 s 70422 15703 70422 15703 4 DVSS
port 2 nsew
rlabel metal3 s 70444 21860 70444 21860 4 DVSS
port 2 nsew
rlabel metal3 s 70444 26053 70444 26053 4 DVSS
port 2 nsew
rlabel metal3 s 70444 40295 70444 40295 4 DVSS
port 2 nsew
rlabel metal3 s 70444 47548 70444 47548 4 DVSS
port 2 nsew
rlabel metal3 s 70444 57811 70444 57811 4 DVSS
port 2 nsew
rlabel metal3 s 70444 61011 70444 61011 4 DVSS
port 2 nsew
rlabel metal3 s 70444 65976 70444 65976 4 DVSS
port 2 nsew
rlabel metal5 s 70548 51411 70548 51411 4 VDD
port 3 nsew
rlabel metal5 s 70444 62776 70444 62776 4 VDD
port 3 nsew
rlabel metal5 s 51498 70220 51498 70220 4 VDD
port 3 nsew
rlabel metal5 s 62716 70220 62716 70220 4 VDD
port 3 nsew
rlabel metal5 s 70548 51411 70548 51411 4 VDD
port 3 nsew
rlabel metal5 s 70444 62776 70444 62776 4 VDD
port 3 nsew
rlabel metal5 s 51498 70220 51498 70220 4 VDD
port 3 nsew
rlabel metal5 s 62716 70220 62716 70220 4 VDD
port 3 nsew
rlabel metal5 s 70548 51411 70548 51411 4 VDD
port 3 nsew
rlabel metal5 s 70444 62776 70444 62776 4 VDD
port 3 nsew
rlabel metal5 s 51498 70220 51498 70220 4 VDD
port 3 nsew
rlabel metal5 s 62716 70220 62716 70220 4 VDD
port 3 nsew
rlabel metal4 s 70548 51411 70548 51411 4 VDD
port 3 nsew
rlabel metal4 s 62716 70220 62716 70220 4 VDD
port 3 nsew
rlabel metal4 s 51498 70220 51498 70220 4 VDD
port 3 nsew
rlabel metal4 s 70444 62776 70444 62776 4 VDD
port 3 nsew
rlabel metal3 s 62716 70220 62716 70220 4 VDD
port 3 nsew
rlabel metal3 s 51498 70220 51498 70220 4 VDD
port 3 nsew
rlabel metal3 s 70443 62776 70443 62776 4 VDD
port 3 nsew
rlabel metal3 s 70548 51411 70548 51411 4 VDD
port 3 nsew
rlabel metal5 s 70547 49976 70547 49976 4 VSS
port 4 nsew
rlabel metal5 s 70444 64211 70444 64211 4 VSS
port 4 nsew
rlabel metal5 s 49849 70219 49849 70219 4 VSS
port 4 nsew
rlabel metal5 s 64328 70220 64328 70220 4 VSS
port 4 nsew
rlabel metal5 s 70547 49976 70547 49976 4 VSS
port 4 nsew
rlabel metal5 s 70444 64211 70444 64211 4 VSS
port 4 nsew
rlabel metal5 s 49849 70219 49849 70219 4 VSS
port 4 nsew
rlabel metal5 s 64328 70220 64328 70220 4 VSS
port 4 nsew
rlabel metal5 s 70547 49976 70547 49976 4 VSS
port 4 nsew
rlabel metal5 s 49849 70219 49849 70219 4 VSS
port 4 nsew
rlabel metal5 s 64328 70220 64328 70220 4 VSS
port 4 nsew
rlabel metal4 s 49849 70219 49849 70219 4 VSS
port 4 nsew
rlabel metal4 s 70547 49976 70547 49976 4 VSS
port 4 nsew
rlabel metal4 s 64328 70220 64328 70220 4 VSS
port 4 nsew
rlabel metal4 s 70444 64211 70444 64211 4 VSS
port 4 nsew
rlabel metal3 s 49849 70219 49849 70219 4 VSS
port 4 nsew
rlabel metal3 s 64328 70220 64328 70220 4 VSS
port 4 nsew
rlabel metal3 s 70444 64211 70444 64211 4 VSS
port 4 nsew
rlabel metal3 s 70547 49976 70547 49976 4 VSS
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 71000 71000
<< end >>
