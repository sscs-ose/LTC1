magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1703 -1133 1703 1133
<< metal2 >>
rect -703 128 703 133
rect -703 100 -698 128
rect -670 100 -622 128
rect -594 100 -546 128
rect -518 100 -470 128
rect -442 100 -394 128
rect -366 100 -318 128
rect -290 100 -242 128
rect -214 100 -166 128
rect -138 100 -90 128
rect -62 100 -14 128
rect 14 100 62 128
rect 90 100 138 128
rect 166 100 214 128
rect 242 100 290 128
rect 318 100 366 128
rect 394 100 442 128
rect 470 100 518 128
rect 546 100 594 128
rect 622 100 670 128
rect 698 100 703 128
rect -703 52 703 100
rect -703 24 -698 52
rect -670 24 -622 52
rect -594 24 -546 52
rect -518 24 -470 52
rect -442 24 -394 52
rect -366 24 -318 52
rect -290 24 -242 52
rect -214 24 -166 52
rect -138 24 -90 52
rect -62 24 -14 52
rect 14 24 62 52
rect 90 24 138 52
rect 166 24 214 52
rect 242 24 290 52
rect 318 24 366 52
rect 394 24 442 52
rect 470 24 518 52
rect 546 24 594 52
rect 622 24 670 52
rect 698 24 703 52
rect -703 -24 703 24
rect -703 -52 -698 -24
rect -670 -52 -622 -24
rect -594 -52 -546 -24
rect -518 -52 -470 -24
rect -442 -52 -394 -24
rect -366 -52 -318 -24
rect -290 -52 -242 -24
rect -214 -52 -166 -24
rect -138 -52 -90 -24
rect -62 -52 -14 -24
rect 14 -52 62 -24
rect 90 -52 138 -24
rect 166 -52 214 -24
rect 242 -52 290 -24
rect 318 -52 366 -24
rect 394 -52 442 -24
rect 470 -52 518 -24
rect 546 -52 594 -24
rect 622 -52 670 -24
rect 698 -52 703 -24
rect -703 -100 703 -52
rect -703 -128 -698 -100
rect -670 -128 -622 -100
rect -594 -128 -546 -100
rect -518 -128 -470 -100
rect -442 -128 -394 -100
rect -366 -128 -318 -100
rect -290 -128 -242 -100
rect -214 -128 -166 -100
rect -138 -128 -90 -100
rect -62 -128 -14 -100
rect 14 -128 62 -100
rect 90 -128 138 -100
rect 166 -128 214 -100
rect 242 -128 290 -100
rect 318 -128 366 -100
rect 394 -128 442 -100
rect 470 -128 518 -100
rect 546 -128 594 -100
rect 622 -128 670 -100
rect 698 -128 703 -100
rect -703 -133 703 -128
<< via2 >>
rect -698 100 -670 128
rect -622 100 -594 128
rect -546 100 -518 128
rect -470 100 -442 128
rect -394 100 -366 128
rect -318 100 -290 128
rect -242 100 -214 128
rect -166 100 -138 128
rect -90 100 -62 128
rect -14 100 14 128
rect 62 100 90 128
rect 138 100 166 128
rect 214 100 242 128
rect 290 100 318 128
rect 366 100 394 128
rect 442 100 470 128
rect 518 100 546 128
rect 594 100 622 128
rect 670 100 698 128
rect -698 24 -670 52
rect -622 24 -594 52
rect -546 24 -518 52
rect -470 24 -442 52
rect -394 24 -366 52
rect -318 24 -290 52
rect -242 24 -214 52
rect -166 24 -138 52
rect -90 24 -62 52
rect -14 24 14 52
rect 62 24 90 52
rect 138 24 166 52
rect 214 24 242 52
rect 290 24 318 52
rect 366 24 394 52
rect 442 24 470 52
rect 518 24 546 52
rect 594 24 622 52
rect 670 24 698 52
rect -698 -52 -670 -24
rect -622 -52 -594 -24
rect -546 -52 -518 -24
rect -470 -52 -442 -24
rect -394 -52 -366 -24
rect -318 -52 -290 -24
rect -242 -52 -214 -24
rect -166 -52 -138 -24
rect -90 -52 -62 -24
rect -14 -52 14 -24
rect 62 -52 90 -24
rect 138 -52 166 -24
rect 214 -52 242 -24
rect 290 -52 318 -24
rect 366 -52 394 -24
rect 442 -52 470 -24
rect 518 -52 546 -24
rect 594 -52 622 -24
rect 670 -52 698 -24
rect -698 -128 -670 -100
rect -622 -128 -594 -100
rect -546 -128 -518 -100
rect -470 -128 -442 -100
rect -394 -128 -366 -100
rect -318 -128 -290 -100
rect -242 -128 -214 -100
rect -166 -128 -138 -100
rect -90 -128 -62 -100
rect -14 -128 14 -100
rect 62 -128 90 -100
rect 138 -128 166 -100
rect 214 -128 242 -100
rect 290 -128 318 -100
rect 366 -128 394 -100
rect 442 -128 470 -100
rect 518 -128 546 -100
rect 594 -128 622 -100
rect 670 -128 698 -100
<< metal3 >>
rect -703 128 703 133
rect -703 100 -698 128
rect -670 100 -622 128
rect -594 100 -546 128
rect -518 100 -470 128
rect -442 100 -394 128
rect -366 100 -318 128
rect -290 100 -242 128
rect -214 100 -166 128
rect -138 100 -90 128
rect -62 100 -14 128
rect 14 100 62 128
rect 90 100 138 128
rect 166 100 214 128
rect 242 100 290 128
rect 318 100 366 128
rect 394 100 442 128
rect 470 100 518 128
rect 546 100 594 128
rect 622 100 670 128
rect 698 100 703 128
rect -703 52 703 100
rect -703 24 -698 52
rect -670 24 -622 52
rect -594 24 -546 52
rect -518 24 -470 52
rect -442 24 -394 52
rect -366 24 -318 52
rect -290 24 -242 52
rect -214 24 -166 52
rect -138 24 -90 52
rect -62 24 -14 52
rect 14 24 62 52
rect 90 24 138 52
rect 166 24 214 52
rect 242 24 290 52
rect 318 24 366 52
rect 394 24 442 52
rect 470 24 518 52
rect 546 24 594 52
rect 622 24 670 52
rect 698 24 703 52
rect -703 -24 703 24
rect -703 -52 -698 -24
rect -670 -52 -622 -24
rect -594 -52 -546 -24
rect -518 -52 -470 -24
rect -442 -52 -394 -24
rect -366 -52 -318 -24
rect -290 -52 -242 -24
rect -214 -52 -166 -24
rect -138 -52 -90 -24
rect -62 -52 -14 -24
rect 14 -52 62 -24
rect 90 -52 138 -24
rect 166 -52 214 -24
rect 242 -52 290 -24
rect 318 -52 366 -24
rect 394 -52 442 -24
rect 470 -52 518 -24
rect 546 -52 594 -24
rect 622 -52 670 -24
rect 698 -52 703 -24
rect -703 -100 703 -52
rect -703 -128 -698 -100
rect -670 -128 -622 -100
rect -594 -128 -546 -100
rect -518 -128 -470 -100
rect -442 -128 -394 -100
rect -366 -128 -318 -100
rect -290 -128 -242 -100
rect -214 -128 -166 -100
rect -138 -128 -90 -100
rect -62 -128 -14 -100
rect 14 -128 62 -100
rect 90 -128 138 -100
rect 166 -128 214 -100
rect 242 -128 290 -100
rect 318 -128 366 -100
rect 394 -128 442 -100
rect 470 -128 518 -100
rect 546 -128 594 -100
rect 622 -128 670 -100
rect 698 -128 703 -100
rect -703 -133 703 -128
<< end >>
