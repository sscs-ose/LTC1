** sch_path: /home/shahid/GF180Projects/GF_INV/DAC_low_curr/untitled-18.sch
**.subckt untitled-18 VDD VSS B7 B11 B8 B12 B9 B10
*.iopin VDD
*.iopin VSS
*.ipin B7
*.ipin B11
*.ipin B8
*.ipin B12
*.ipin B9
*.ipin B10
x2 OUT+ OUT- VDD R4 R5 C1 net5 net6 VSS MSB_UNIT_CELL
x3 OUT+ OUT- VDD R3 R4 C4 net5 net6 VSS MSB_UNIT_CELL
x4 OUT+ OUT- VDD R2 R3 C4 net1 net2 VSS MSB_UNIT_CELL
x5 OUT+ OUT- VDD R3 R4 C3 net7 net8 VSS MSB_UNIT_CELL
x6 OUT+ OUT- VDD R2 R3 C3 net3 net4 VSS MSB_UNIT_CELL
x7 OUT+ OUT- VDD R1 R2 C6 net3 net4 VSS MSB_UNIT_CELL
x8 VDD C32_U net5 C32_D net6 VSS CM_32_s
x9 VDD C32_U net7 C32_D net8 VSS CM_32_s
x10 VDD C32_U net1 C32_D net2 VSS CM_32_s
x11 VDD C32_U net3 C32_D net4 VSS CM_32_s
x12 OUT+ OUT- VDD R5 R6 C3 net25 net26 VSS MSB_UNIT_CELL
x13 OUT+ OUT- VDD R5 R6 C4 net23 net24 VSS MSB_UNIT_CELL
x14 OUT+ OUT- VDD R5 R6 C5 net23 net24 VSS MSB_UNIT_CELL
x15 OUT+ OUT- VDD R5 R6 C2 net25 net26 VSS MSB_UNIT_CELL
x16 OUT+ OUT- VDD R5 R6 C6 net21 net22 VSS MSB_UNIT_CELL
x17 OUT+ OUT- VDD R4 R5 C0 net7 net8 VSS MSB_UNIT_CELL
x18 OUT+ OUT- VDD R3 R4 C2 net9 net10 VSS MSB_UNIT_CELL
x19 OUT+ OUT- VDD R2 R3 C2 net11 net12 VSS MSB_UNIT_CELL
x20 OUT+ OUT- VDD R1 R2 C3 net11 net12 VSS MSB_UNIT_CELL
x21 OUT+ OUT- VDD R1 R2 C2 net15 net16 VSS MSB_UNIT_CELL
x22 OUT+ OUT- VDD R1 R2 C4 net15 net16 VSS MSB_UNIT_CELL
x23 OUT+ OUT- VDD R1 R2 C5 net15 net16 VSS MSB_UNIT_CELL
x24 OUT+ OUT- VDD R0 R1 C4 net17 net18 VSS MSB_UNIT_CELL
x25 OUT+ OUT- VDD R0 R1 C5 net17 net18 VSS MSB_UNIT_CELL
x26 OUT+ OUT- VDD R1 R2 VSS net1 net2 VSS MSB_UNIT_CELL
x27 OUT+ OUT- VDD R2 R3 C5 net19 net20 VSS MSB_UNIT_CELL
x28 OUT+ OUT- VDD R3 R4 C5 net21 net22 VSS MSB_UNIT_CELL
x29 OUT+ OUT- VDD R4 R5 C2 net21 net22 VSS MSB_UNIT_CELL
x30 OUT+ OUT- VDD R5 R6 C1 net9 net10 VSS MSB_UNIT_CELL
x31 VDD net7 net9 net8 net10 VSS CM_32_s
x32 OUT+ OUT- VDD R3 R4 C1 net9 net10 VSS MSB_UNIT_CELL
x35 OUT+ OUT- VDD R2 R3 C1 net11 net12 VSS MSB_UNIT_CELL
x33 VDD net11 net13 net12 net14 VSS CM_32_s
x34 VDD net3 net11 net4 net12 VSS CM_32_s
x36 OUT+ OUT- VDD R5 R6 C0 net27 net28 VSS MSB_UNIT_CELL
x37 VDD net9 net27 net10 net28 VSS CM_32_s
x38 OUT+ OUT- VDD R3 R4 C0 net27 net28 VSS MSB_UNIT_CELL
x39 OUT+ OUT- VDD R1 R2 C0 net13 net14 VSS MSB_UNIT_CELL
x40 OUT+ OUT- VDD R2 R3 C0 net27 net28 VSS MSB_UNIT_CELL
x41 OUT+ OUT- VDD R1 R2 C1 net13 net14 VSS MSB_UNIT_CELL
x42 OUT+ OUT- VDD R4 R5 C4 net35 net36 VSS MSB_UNIT_CELL
x43 VDD net21 net35 net22 net36 VSS CM_32_s
x44 OUT+ OUT- VDD R3 R4 VSS net33 net34 VSS MSB_UNIT_CELL
x45 OUT+ OUT- VDD R0 R1 VSS net33 net34 VSS MSB_UNIT_CELL
x47 VDD net19 net33 net20 net34 VSS CM_32_s
x48 OUT+ OUT- VDD R4 R5 C3 net35 net36 VSS MSB_UNIT_CELL
x49 VDD net5 net21 net6 net22 VSS CM_32_s
x50 OUT+ OUT- VDD R3 R4 C6 net35 net36 VSS MSB_UNIT_CELL
x51 OUT+ OUT- VDD R0 R1 C6 net19 net20 VSS MSB_UNIT_CELL
x52 OUT+ OUT- VDD R2 R3 C6 net19 net20 VSS MSB_UNIT_CELL
x46 OUT+ OUT- VDD R2 R3 VSS net33 net34 VSS MSB_UNIT_CELL
x53 VDD net1 net19 net2 net20 VSS CM_32_s
x54 OUT+ OUT- VDD R0 R1 C2 net29 net30 VSS MSB_UNIT_CELL
x55 OUT+ OUT- VDD R0 R1 C1 net13 net14 VSS MSB_UNIT_CELL
x56 OUT+ OUT- VDD R0 R1 C0 net13 net14 VSS MSB_UNIT_CELL
x57 VDD net3 net15 net4 net16 VSS CM_32_s
x58 OUT+ OUT- VDD R0 R1 C3 net17 net18 VSS MSB_UNIT_CELL
x59 VDD net1 net17 net2 net18 VSS CM_32_s
x60 OUT+ OUT- VDD VDD R0 C4 net31 net32 VSS MSB_UNIT_CELL
x61 OUT+ OUT- VDD VDD R0 VSS net33 net34 VSS MSB_UNIT_CELL
x62 OUT+ OUT- VDD VDD R0 C5 net31 net32 VSS MSB_UNIT_CELL
x63 OUT+ OUT- VDD VDD R0 C1 net29 net30 VSS MSB_UNIT_CELL
x64 OUT+ OUT- VDD VDD R0 C0 net29 net30 VSS MSB_UNIT_CELL
x65 VDD net15 net29 net16 net30 VSS CM_32_s
x66 OUT+ OUT- VDD VDD R0 C2 net29 net30 VSS MSB_UNIT_CELL
x67 OUT+ OUT- VDD VDD R0 C3 net31 net32 VSS MSB_UNIT_CELL
x68 VDD net17 net31 net18 net32 VSS CM_32_s
x69 OUT+ OUT- VDD VDD R0 C6 net31 net32 VSS MSB_UNIT_CELL
x70 OUT+ OUT- VDD R6 VSS C2 net25 net26 VSS MSB_UNIT_CELL
x71 OUT+ OUT- VDD R6 VSS C1 net27 net28 VSS MSB_UNIT_CELL
x73 VDD net7 net25 net8 net26 VSS CM_32_s
x74 OUT+ OUT- VDD R6 VSS C4 net23 net24 VSS MSB_UNIT_CELL
x75 VDD net5 net23 net6 net24 VSS CM_32_s
x76 OUT+ OUT- VDD R5 R6 VSS net37 net38 VSS MSB_UNIT_CELL
x77 OUT+ OUT- VDD R4 R5 C5 net35 net36 VSS MSB_UNIT_CELL
x78 OUT+ OUT- VDD R4 R5 C6 net37 net38 VSS MSB_UNIT_CELL
x72 OUT+ OUT- VDD R6 VSS C3 net39 net40 VSS MSB_UNIT_CELL
x79 OUT+ OUT- VDD R6 VSS C0 net39 net40 VSS MSB_UNIT_CELL
x80 VDD net25 net39 net26 net40 VSS CM_32_s
x81 OUT+ OUT- VDD R6 VSS C5 net39 net40 VSS MSB_UNIT_CELL
x82 VDD net23 net37 net24 net38 VSS CM_32_s
x83 OUT+ OUT- VDD R6 VSS C6 net37 net38 VSS MSB_UNIT_CELL
x85 OUT+ OUT- VDD R4 R5 VSS net37 net38 VSS MSB_UNIT_CELL
x84 R6 VDD R5 VSS R4 B12 R3 R2 B11 R1 B10 R0 Thermo_Decoder
x86 C6 VDD C5 VSS C4 B9 C3 C2 B8 C1 B7 C0 Thermo_Decoder
XM11 C32_U C32_U C32_D VSS nfet_03v3 L=0.5u W=19.2u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM12 C32_D C32_D VSS VSS nfet_03v3 L=0.5u W=19.2u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
V1 VSS GND 0
.save i(v1)
V2 VDD VSS 3.3
.save i(v2)
I1 VDD C32_U 80u
V13 B8 VSS pulse(0 3.3 0 10p 10p 6.4u 12.8u)
.save i(v13)
V14 B7 VSS pulse(0 3.3 0 10p 10p 3.2u 6.4u)
.save i(v14)
V9 B9 VSS pulse(0 3.3 0 10p 10p 12.8u 25.6u)
.save i(v9)
V3 B10 VSS pulse(0 3.3 0 10p 10p 25.6u 51.2u)
.save i(v3)
V4 B11 VSS pulse(0 3.3 0 10p 10p 51.2u 102.4u)
.save i(v4)
V5 B12 VSS pulse(0 3.3 0 10p 10p 102.4u 204.8u)
.save i(v5)
R1 OUT+ VDD 200 m=1
R2 OUT- VDD 200 m=1
**** begin user architecture code

.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical



.options savecurrents
.control
*save all
op

tran tmax 205u
plot v(OUT+) v(OUT-)

*write DAC_12Bit_TB.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  MSB_UNIT_CELL.sym # of pins=9
** sym_path: /home/shahid/GF180Projects/GF_INV/DAC_low_curr/MSB_UNIT_CELL.sym
** sch_path: /home/shahid/GF180Projects/GF_INV/DAC_low_curr/MSB_UNIT_CELL.sch
.subckt MSB_UNIT_CELL IOUT+ IOUT- VDD Ri-1 Ri Ci IM_T IM VSS
*.iopin VDD
*.iopin VSS
*.ipin Ri-1
*.ipin Ri
*.ipin Ci
*.ipin IM_T
*.ipin IM
*.opin IOUT+
*.opin IOUT-
x1 VDD VSS Ri-1 Ri Ci net2 net3 Local_Enc
XM1 IOUT+ net2 net1 VSS nfet_03v3 L=0.5u W=38.4u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 IOUT- net3 net1 VSS nfet_03v3 L=0.5u W=38.4u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 net1 IM_T net4 VSS nfet_03v3 L=0.5u W=38.4u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 net4 IM VSS VSS nfet_03v3 L=0.5u W=38.4u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  CM_32_s.sym # of pins=6
** sym_path: /home/shahid/GF180Projects/GF_INV/DAC_low_curr/CM_32_s.sym
** sch_path: /home/shahid/GF180Projects/GF_INV/DAC_low_curr/CM_32_s.sch
.subckt CM_32_s VDD G0_2 G3_2 G0_1 G3_1 VSS
*.ipin G0_2
*.iopin VDD
*.iopin VSS
*.opin G3_2
*.ipin G0_1
*.opin G3_1
XM1 net2 G0_2 net1 VSS nfet_03v3 L=0.5u W=19.2u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 net1 G0_1 VSS VSS nfet_03v3 L=0.5u W=19.2u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM7 net2 net2 net3 VDD pfet_03v3 L=0.5u W=19.2u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM8 net3 net3 VDD VDD pfet_03v3 L=0.5u W=19.2u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM9 G3_2 net2 net4 VDD pfet_03v3 L=0.5u W=19.2u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM10 net4 net3 VDD VDD pfet_03v3 L=0.5u W=19.2u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM11 G3_2 G3_2 G3_1 VSS nfet_03v3 L=0.5u W=19.2u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM12 G3_1 G3_1 VSS VSS nfet_03v3 L=0.5u W=19.2u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  Thermo_Decoder.sym # of pins=12
** sym_path: /home/shahid/GF180Projects/GF_INV/DAC_low_curr/Thermo_Decoder.sym
** sch_path: /home/shahid/GF180Projects/GF_INV/DAC_low_curr/Thermo_Decoder.sch
.subckt Thermo_Decoder D1 VDD D2 VSS D3 B1 D4 D5 B2 D6 B3 D7
*.iopin VDD
*.iopin VSS
*.ipin B1
*.ipin B2
*.ipin B3
*.opin D3
*.opin D4
*.opin D1
*.opin D2
*.opin D6
*.opin D7
*.opin D5
x1 VDD VSS B1 B2 net8 AND
x2 VDD VSS net1 D1 inv
x3 VDD VSS B1 B2 net4 OR
x4 VDD VSS B2 B3 net9 OR
x5 VDD VSS B1 B2 net2 AND
x6 VDD VSS B3 net8 net1 AND
x7 VDD VSS net2 D2 inv
x8 VDD VSS B1 net9 net3 AND
x9 VDD VSS net3 D3 inv
x10 VDD VSS B1 D4 inv
x11 VDD VSS net4 D6 inv
x12 VDD VSS B2 B3 net6 AND
x13 VDD VSS B1 net6 net7 OR
x14 VDD VSS net7 D5 inv
x15 VDD VSS B1 B2 net10 OR
x16 VDD VSS B3 net10 net5 OR
x17 VDD VSS net5 D7 inv
.ends


* expanding   symbol:  Local_Enc.sym # of pins=7
** sym_path: /home/shahid/GF180Projects/GF_INV/DAC_low_curr/Local_Enc.sym
** sch_path: /home/shahid/GF180Projects/GF_INV/DAC_low_curr/Local_Enc.sch
.subckt Local_Enc VDD VSS Ri-1 Ri Ci Q QB
*.iopin VDD
*.iopin VSS
*.ipin Ri-1
*.ipin Ri
*.ipin Ci
*.opin Q
*.opin QB
x1 VDD VSS Ri-1 Ri-1 net5 NAND
x2 VDD VSS Ri Ri net6 NAND
x3 VDD VSS Ci Ci net7 NAND
x4 VDD VSS net5 net5 net3 NAND
x5 VDD VSS net6 net7 net4 NAND
x6 VDD VSS net4 net3 net2 NAND
x7 VDD VSS net2 net2 net1 NAND
x8 VDD VSS Q net1 QB NAND
x9 VDD VSS net2 QB Q NAND
.ends


* expanding   symbol:  AND.sym # of pins=5
** sym_path: /home/shahid/GF180Projects/GF_INV/DAC_low_curr/AND.sym
** sch_path: /home/shahid/GF180Projects/GF_INV/DAC_low_curr/AND.sch
.subckt AND VDD VSS A B OUT
*.iopin VDD
*.iopin VSS
*.ipin A
*.ipin B
*.opin OUT
XM1 net2 A VSS VSS nfet_03v3 L=0.28u W=0.5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 net1 B VDD VDD pfet_03v3 L=0.28u W=0.5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 net1 A VDD VDD pfet_03v3 L=0.28u W=0.5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 net1 B net2 VSS nfet_03v3 L=0.28u W=0.5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
x1 VSS VDD OUT net1 GF_INV
.ends


* expanding   symbol:  inv.sym # of pins=4
** sym_path: /home/shahid/GF180Projects/GF_INV/DAC_low_curr/inv.sym
** sch_path: /home/shahid/GF180Projects/GF_INV/DAC_low_curr/inv.sch
.subckt inv VDD VSS IN OUT
*.opin OUT
*.iopin VDD
*.iopin VSS
*.ipin IN
x1 VSS VDD net1 IN GF_INV
x2 VSS VDD OUT net1 GF_INV
.ends


* expanding   symbol:  OR.sym # of pins=5
** sym_path: /home/shahid/GF180Projects/GF_INV/DAC_low_curr/OR.sym
** sch_path: /home/shahid/GF180Projects/GF_INV/DAC_low_curr/OR.sch
.subckt OR VDD VSS A B OUT
*.iopin VDD
*.iopin VSS
*.ipin A
*.ipin B
*.opin OUT
x1 VSS VDD OUT net1 GF_INV
XM1 net1 A VSS VSS nfet_03v3 L=0.28u W=0.25u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 net2 B VDD VDD pfet_03v3 L=0.28u W=1u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM5 net1 A net2 VDD pfet_03v3 L=0.28u W=1u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM6 net1 B VSS VSS nfet_03v3 L=0.28u W=0.25u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  NAND.sym # of pins=5
** sym_path: /home/shahid/GF180Projects/GF_INV/DAC_low_curr/NAND.sym
** sch_path: /home/shahid/GF180Projects/GF_INV/DAC_low_curr/NAND.sch
.subckt NAND VDD VSS A B OUT
*.iopin VDD
*.iopin VSS
*.ipin A
*.ipin B
*.opin OUT
XM2 OUT A VDD VDD pfet_03v3 L=0.28u W=0.5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 OUT B VDD VDD pfet_03v3 L=0.28u W=0.5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM1 OUT A net1 VSS nfet_03v3 L=0.28u W=0.5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 net1 B VSS VSS nfet_03v3 L=0.28u W=0.5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  GF_INV.sym # of pins=4
** sym_path: /home/shahid/GF180Projects/GF_INV/DAC_low_curr/GF_INV.sym
** sch_path: /home/shahid/GF180Projects/GF_INV/DAC_low_curr/GF_INV.sch
.subckt GF_INV VSS VDD OUT IN
*.iopin VDD
*.iopin VSS
*.ipin IN
*.opin OUT
XM1 OUT IN VSS VSS nfet_03v3 L=0.28u W=0.25u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 OUT IN VDD VDD pfet_03v3 L=0.28u W=0.5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends

.GLOBAL GND
.end
