magic
tech gf180mcuC
magscale 1 10
timestamp 1714126980
<< error_p >>
rect -343 -48 -297 48
rect -183 -48 -137 48
rect -23 -48 23 48
rect 137 -48 183 48
rect 297 -48 343 48
<< pwell >>
rect -380 -118 380 118
<< nmos >>
rect -268 -50 -212 50
rect -108 -50 -52 50
rect 52 -50 108 50
rect 212 -50 268 50
<< ndiff >>
rect -356 37 -268 50
rect -356 -37 -343 37
rect -297 -37 -268 37
rect -356 -50 -268 -37
rect -212 37 -108 50
rect -212 -37 -183 37
rect -137 -37 -108 37
rect -212 -50 -108 -37
rect -52 37 52 50
rect -52 -37 -23 37
rect 23 -37 52 37
rect -52 -50 52 -37
rect 108 37 212 50
rect 108 -37 137 37
rect 183 -37 212 37
rect 108 -50 212 -37
rect 268 37 356 50
rect 268 -37 297 37
rect 343 -37 356 37
rect 268 -50 356 -37
<< ndiffc >>
rect -343 -37 -297 37
rect -183 -37 -137 37
rect -23 -37 23 37
rect 137 -37 183 37
rect 297 -37 343 37
<< polysilicon >>
rect -268 50 -212 94
rect -108 50 -52 94
rect 52 50 108 94
rect 212 50 268 94
rect -268 -94 -212 -50
rect -108 -94 -52 -50
rect 52 -94 108 -50
rect 212 -94 268 -50
<< metal1 >>
rect -343 37 -297 48
rect -343 -48 -297 -37
rect -183 37 -137 48
rect -183 -48 -137 -37
rect -23 37 23 48
rect -23 -48 23 -37
rect 137 37 183 48
rect 137 -48 183 -37
rect 297 37 343 48
rect 297 -48 343 -37
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 0.5 l 0.280 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
