* NGSPICE file created from nand2_flat.ext - technology: gf180mcuC

.subckt NAND_PEX IN1 VSS VDD OUT IN2
X0 OUT IN1.t0 a_168_68# VSS.t0 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1 OUT IN2.t0 VDD.t4 VDD.t3 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2 a_168_68# IN2.t1 VSS.t2 VSS.t1 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X3 VDD IN1.t1 OUT.t1 VDD.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
R0 IN1.n0 IN1.t0 31.528
R1 IN1.n0 IN1.t1 15.3826
R2 IN1 IN1.n0 8.85806
R3 OUT OUT.n2 7.15141
R4 OUT OUT.n1 3.22776
R5 OUT.n1 OUT.t1 2.2755
R6 OUT.n1 OUT.n0 2.2755
R7 VSS.n0 VSS.t0 596.558
R8 VSS.n0 VSS.t1 397.707
R9 VSS VSS.t2 7.30963
R10 VSS VSS.n1 5.2005
R11 VSS VSS.n1 5.2005
R12 VSS.n1 VSS.n0 2.6005
R13 IN2.n0 IN2.t0 30.9379
R14 IN2.n0 IN2.t1 21.6422
R15 IN2 IN2.n0 4.005
R16 VDD.n2 VDD.t0 193.183
R17 VDD.n2 VDD.t3 109.849
R18 VDD VDD.n0 5.23855
R19 VDD.n4 VDD.t4 5.21701
R20 VDD.n4 VDD.n3 3.1505
R21 VDD.n3 VDD.n2 3.1505
R22 VDD.n3 VDD.n1 0.109121
R23 VDD VDD.n4 0.00166129
C0 a_168_68# OUT 0.069f
C1 OUT IN1 0.191f
C2 VDD IN2 0.146f
C3 VDD a_168_68# 3.14e-19
C4 a_168_68# IN2 0.00347f
C5 VDD IN1 0.225f
C6 IN1 IN2 0.0466f
C7 a_168_68# IN1 0.00348f
C8 VDD OUT 0.206f
C9 OUT IN2 0.0956f
.ends

