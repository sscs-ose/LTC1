magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2045 -2609 2045 2609
<< psubdiff >>
rect -45 587 45 609
rect -45 -587 -23 587
rect 23 -587 45 587
rect -45 -609 45 -587
<< psubdiffcont >>
rect -23 -587 23 587
<< metal1 >>
rect -34 587 34 598
rect -34 -587 -23 587
rect 23 -587 34 587
rect -34 -598 34 -587
<< end >>
