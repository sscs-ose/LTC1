magic
tech gf180mcuC
magscale 1 10
timestamp 1699203423
<< nwell >>
rect -1824 -516 1824 516
<< nsubdiff >>
rect -1800 420 1800 492
rect -1800 -420 -1728 420
rect 1728 -420 1800 420
rect -1800 -492 1800 -420
<< polysilicon >>
rect -1640 319 -1440 332
rect -1640 273 -1627 319
rect -1453 273 -1440 319
rect -1640 230 -1440 273
rect -1640 -273 -1440 -230
rect -1640 -319 -1627 -273
rect -1453 -319 -1440 -273
rect -1640 -332 -1440 -319
rect -1360 319 -1160 332
rect -1360 273 -1347 319
rect -1173 273 -1160 319
rect -1360 230 -1160 273
rect -1360 -273 -1160 -230
rect -1360 -319 -1347 -273
rect -1173 -319 -1160 -273
rect -1360 -332 -1160 -319
rect -1080 319 -880 332
rect -1080 273 -1067 319
rect -893 273 -880 319
rect -1080 230 -880 273
rect -1080 -273 -880 -230
rect -1080 -319 -1067 -273
rect -893 -319 -880 -273
rect -1080 -332 -880 -319
rect -800 319 -600 332
rect -800 273 -787 319
rect -613 273 -600 319
rect -800 230 -600 273
rect -800 -273 -600 -230
rect -800 -319 -787 -273
rect -613 -319 -600 -273
rect -800 -332 -600 -319
rect -520 319 -320 332
rect -520 273 -507 319
rect -333 273 -320 319
rect -520 230 -320 273
rect -520 -273 -320 -230
rect -520 -319 -507 -273
rect -333 -319 -320 -273
rect -520 -332 -320 -319
rect -240 319 -40 332
rect -240 273 -227 319
rect -53 273 -40 319
rect -240 230 -40 273
rect -240 -273 -40 -230
rect -240 -319 -227 -273
rect -53 -319 -40 -273
rect -240 -332 -40 -319
rect 40 319 240 332
rect 40 273 53 319
rect 227 273 240 319
rect 40 230 240 273
rect 40 -273 240 -230
rect 40 -319 53 -273
rect 227 -319 240 -273
rect 40 -332 240 -319
rect 320 319 520 332
rect 320 273 333 319
rect 507 273 520 319
rect 320 230 520 273
rect 320 -273 520 -230
rect 320 -319 333 -273
rect 507 -319 520 -273
rect 320 -332 520 -319
rect 600 319 800 332
rect 600 273 613 319
rect 787 273 800 319
rect 600 230 800 273
rect 600 -273 800 -230
rect 600 -319 613 -273
rect 787 -319 800 -273
rect 600 -332 800 -319
rect 880 319 1080 332
rect 880 273 893 319
rect 1067 273 1080 319
rect 880 230 1080 273
rect 880 -273 1080 -230
rect 880 -319 893 -273
rect 1067 -319 1080 -273
rect 880 -332 1080 -319
rect 1160 319 1360 332
rect 1160 273 1173 319
rect 1347 273 1360 319
rect 1160 230 1360 273
rect 1160 -273 1360 -230
rect 1160 -319 1173 -273
rect 1347 -319 1360 -273
rect 1160 -332 1360 -319
rect 1440 319 1640 332
rect 1440 273 1453 319
rect 1627 273 1640 319
rect 1440 230 1640 273
rect 1440 -273 1640 -230
rect 1440 -319 1453 -273
rect 1627 -319 1640 -273
rect 1440 -332 1640 -319
<< polycontact >>
rect -1627 273 -1453 319
rect -1627 -319 -1453 -273
rect -1347 273 -1173 319
rect -1347 -319 -1173 -273
rect -1067 273 -893 319
rect -1067 -319 -893 -273
rect -787 273 -613 319
rect -787 -319 -613 -273
rect -507 273 -333 319
rect -507 -319 -333 -273
rect -227 273 -53 319
rect -227 -319 -53 -273
rect 53 273 227 319
rect 53 -319 227 -273
rect 333 273 507 319
rect 333 -319 507 -273
rect 613 273 787 319
rect 613 -319 787 -273
rect 893 273 1067 319
rect 893 -319 1067 -273
rect 1173 273 1347 319
rect 1173 -319 1347 -273
rect 1453 273 1627 319
rect 1453 -319 1627 -273
<< ppolyres >>
rect -1640 -230 -1440 230
rect -1360 -230 -1160 230
rect -1080 -230 -880 230
rect -800 -230 -600 230
rect -520 -230 -320 230
rect -240 -230 -40 230
rect 40 -230 240 230
rect 320 -230 520 230
rect 600 -230 800 230
rect 880 -230 1080 230
rect 1160 -230 1360 230
rect 1440 -230 1640 230
<< metal1 >>
rect -1638 273 -1627 319
rect -1453 273 -1442 319
rect -1358 273 -1347 319
rect -1173 273 -1162 319
rect -1078 273 -1067 319
rect -893 273 -882 319
rect -798 273 -787 319
rect -613 273 -602 319
rect -518 273 -507 319
rect -333 273 -322 319
rect -238 273 -227 319
rect -53 273 -42 319
rect 42 273 53 319
rect 227 273 238 319
rect 322 273 333 319
rect 507 273 518 319
rect 602 273 613 319
rect 787 273 798 319
rect 882 273 893 319
rect 1067 273 1078 319
rect 1162 273 1173 319
rect 1347 273 1358 319
rect 1442 273 1453 319
rect 1627 273 1638 319
rect -1638 -319 -1627 -273
rect -1453 -319 -1442 -273
rect -1358 -319 -1347 -273
rect -1173 -319 -1162 -273
rect -1078 -319 -1067 -273
rect -893 -319 -882 -273
rect -798 -319 -787 -273
rect -613 -319 -602 -273
rect -518 -319 -507 -273
rect -333 -319 -322 -273
rect -238 -319 -227 -273
rect -53 -319 -42 -273
rect 42 -319 53 -273
rect 227 -319 238 -273
rect 322 -319 333 -273
rect 507 -319 518 -273
rect 602 -319 613 -273
rect 787 -319 798 -273
rect 882 -319 893 -273
rect 1067 -319 1078 -273
rect 1162 -319 1173 -273
rect 1347 -319 1358 -273
rect 1442 -319 1453 -273
rect 1627 -319 1638 -273
<< properties >>
string FIXED_BBOX -1764 -456 1764 456
string gencell ppolyf_u
string library gf180mcu
string parameters w 1.0 l 2.3 m 1 nx 12 wmin 0.80 lmin 1.00 rho 315 val 779.032 dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 0 grc 0 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 0
<< end >>
