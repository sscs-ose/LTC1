magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -2446 -2242 2446 2242
<< nwell >>
rect -446 -242 446 242
<< pmos >>
rect -272 -112 -160 112
rect -56 -112 56 112
rect 160 -112 272 112
<< pdiff >>
rect -360 70 -272 112
rect -360 -70 -347 70
rect -301 -70 -272 70
rect -360 -112 -272 -70
rect -160 70 -56 112
rect -160 -70 -131 70
rect -85 -70 -56 70
rect -160 -112 -56 -70
rect 56 70 160 112
rect 56 -70 85 70
rect 131 -70 160 70
rect 56 -112 160 -70
rect 272 70 360 112
rect 272 -70 301 70
rect 347 -70 360 70
rect 272 -112 360 -70
<< pdiffc >>
rect -347 -70 -301 70
rect -131 -70 -85 70
rect 85 -70 131 70
rect 301 -70 347 70
<< polysilicon >>
rect -272 112 -160 156
rect -56 112 56 156
rect 160 112 272 156
rect -272 -156 -160 -112
rect -56 -156 56 -112
rect 160 -156 272 -112
<< metal1 >>
rect -347 70 -301 110
rect -347 -110 -301 -70
rect -131 70 -85 110
rect -131 -110 -85 -70
rect 85 70 131 110
rect 85 -110 131 -70
rect 301 70 347 110
rect 301 -110 347 -70
<< end >>
