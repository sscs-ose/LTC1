magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -4916 -2348 4916 2348
<< pwell >>
rect -2916 -348 2916 348
<< nmos >>
rect -2804 -280 -2704 280
rect -2600 -280 -2500 280
rect -2396 -280 -2296 280
rect -2192 -280 -2092 280
rect -1988 -280 -1888 280
rect -1784 -280 -1684 280
rect -1580 -280 -1480 280
rect -1376 -280 -1276 280
rect -1172 -280 -1072 280
rect -968 -280 -868 280
rect -764 -280 -664 280
rect -560 -280 -460 280
rect -356 -280 -256 280
rect -152 -280 -52 280
rect 52 -280 152 280
rect 256 -280 356 280
rect 460 -280 560 280
rect 664 -280 764 280
rect 868 -280 968 280
rect 1072 -280 1172 280
rect 1276 -280 1376 280
rect 1480 -280 1580 280
rect 1684 -280 1784 280
rect 1888 -280 1988 280
rect 2092 -280 2192 280
rect 2296 -280 2396 280
rect 2500 -280 2600 280
rect 2704 -280 2804 280
<< ndiff >>
rect -2892 258 -2804 280
rect -2892 -258 -2879 258
rect -2833 -258 -2804 258
rect -2892 -280 -2804 -258
rect -2704 258 -2600 280
rect -2704 -258 -2675 258
rect -2629 -258 -2600 258
rect -2704 -280 -2600 -258
rect -2500 258 -2396 280
rect -2500 -258 -2471 258
rect -2425 -258 -2396 258
rect -2500 -280 -2396 -258
rect -2296 258 -2192 280
rect -2296 -258 -2267 258
rect -2221 -258 -2192 258
rect -2296 -280 -2192 -258
rect -2092 258 -1988 280
rect -2092 -258 -2063 258
rect -2017 -258 -1988 258
rect -2092 -280 -1988 -258
rect -1888 258 -1784 280
rect -1888 -258 -1859 258
rect -1813 -258 -1784 258
rect -1888 -280 -1784 -258
rect -1684 258 -1580 280
rect -1684 -258 -1655 258
rect -1609 -258 -1580 258
rect -1684 -280 -1580 -258
rect -1480 258 -1376 280
rect -1480 -258 -1451 258
rect -1405 -258 -1376 258
rect -1480 -280 -1376 -258
rect -1276 258 -1172 280
rect -1276 -258 -1247 258
rect -1201 -258 -1172 258
rect -1276 -280 -1172 -258
rect -1072 258 -968 280
rect -1072 -258 -1043 258
rect -997 -258 -968 258
rect -1072 -280 -968 -258
rect -868 258 -764 280
rect -868 -258 -839 258
rect -793 -258 -764 258
rect -868 -280 -764 -258
rect -664 258 -560 280
rect -664 -258 -635 258
rect -589 -258 -560 258
rect -664 -280 -560 -258
rect -460 258 -356 280
rect -460 -258 -431 258
rect -385 -258 -356 258
rect -460 -280 -356 -258
rect -256 258 -152 280
rect -256 -258 -227 258
rect -181 -258 -152 258
rect -256 -280 -152 -258
rect -52 258 52 280
rect -52 -258 -23 258
rect 23 -258 52 258
rect -52 -280 52 -258
rect 152 258 256 280
rect 152 -258 181 258
rect 227 -258 256 258
rect 152 -280 256 -258
rect 356 258 460 280
rect 356 -258 385 258
rect 431 -258 460 258
rect 356 -280 460 -258
rect 560 258 664 280
rect 560 -258 589 258
rect 635 -258 664 258
rect 560 -280 664 -258
rect 764 258 868 280
rect 764 -258 793 258
rect 839 -258 868 258
rect 764 -280 868 -258
rect 968 258 1072 280
rect 968 -258 997 258
rect 1043 -258 1072 258
rect 968 -280 1072 -258
rect 1172 258 1276 280
rect 1172 -258 1201 258
rect 1247 -258 1276 258
rect 1172 -280 1276 -258
rect 1376 258 1480 280
rect 1376 -258 1405 258
rect 1451 -258 1480 258
rect 1376 -280 1480 -258
rect 1580 258 1684 280
rect 1580 -258 1609 258
rect 1655 -258 1684 258
rect 1580 -280 1684 -258
rect 1784 258 1888 280
rect 1784 -258 1813 258
rect 1859 -258 1888 258
rect 1784 -280 1888 -258
rect 1988 258 2092 280
rect 1988 -258 2017 258
rect 2063 -258 2092 258
rect 1988 -280 2092 -258
rect 2192 258 2296 280
rect 2192 -258 2221 258
rect 2267 -258 2296 258
rect 2192 -280 2296 -258
rect 2396 258 2500 280
rect 2396 -258 2425 258
rect 2471 -258 2500 258
rect 2396 -280 2500 -258
rect 2600 258 2704 280
rect 2600 -258 2629 258
rect 2675 -258 2704 258
rect 2600 -280 2704 -258
rect 2804 258 2892 280
rect 2804 -258 2833 258
rect 2879 -258 2892 258
rect 2804 -280 2892 -258
<< ndiffc >>
rect -2879 -258 -2833 258
rect -2675 -258 -2629 258
rect -2471 -258 -2425 258
rect -2267 -258 -2221 258
rect -2063 -258 -2017 258
rect -1859 -258 -1813 258
rect -1655 -258 -1609 258
rect -1451 -258 -1405 258
rect -1247 -258 -1201 258
rect -1043 -258 -997 258
rect -839 -258 -793 258
rect -635 -258 -589 258
rect -431 -258 -385 258
rect -227 -258 -181 258
rect -23 -258 23 258
rect 181 -258 227 258
rect 385 -258 431 258
rect 589 -258 635 258
rect 793 -258 839 258
rect 997 -258 1043 258
rect 1201 -258 1247 258
rect 1405 -258 1451 258
rect 1609 -258 1655 258
rect 1813 -258 1859 258
rect 2017 -258 2063 258
rect 2221 -258 2267 258
rect 2425 -258 2471 258
rect 2629 -258 2675 258
rect 2833 -258 2879 258
<< polysilicon >>
rect -2804 280 -2704 324
rect -2600 280 -2500 324
rect -2396 280 -2296 324
rect -2192 280 -2092 324
rect -1988 280 -1888 324
rect -1784 280 -1684 324
rect -1580 280 -1480 324
rect -1376 280 -1276 324
rect -1172 280 -1072 324
rect -968 280 -868 324
rect -764 280 -664 324
rect -560 280 -460 324
rect -356 280 -256 324
rect -152 280 -52 324
rect 52 280 152 324
rect 256 280 356 324
rect 460 280 560 324
rect 664 280 764 324
rect 868 280 968 324
rect 1072 280 1172 324
rect 1276 280 1376 324
rect 1480 280 1580 324
rect 1684 280 1784 324
rect 1888 280 1988 324
rect 2092 280 2192 324
rect 2296 280 2396 324
rect 2500 280 2600 324
rect 2704 280 2804 324
rect -2804 -324 -2704 -280
rect -2600 -324 -2500 -280
rect -2396 -324 -2296 -280
rect -2192 -324 -2092 -280
rect -1988 -324 -1888 -280
rect -1784 -324 -1684 -280
rect -1580 -324 -1480 -280
rect -1376 -324 -1276 -280
rect -1172 -324 -1072 -280
rect -968 -324 -868 -280
rect -764 -324 -664 -280
rect -560 -324 -460 -280
rect -356 -324 -256 -280
rect -152 -324 -52 -280
rect 52 -324 152 -280
rect 256 -324 356 -280
rect 460 -324 560 -280
rect 664 -324 764 -280
rect 868 -324 968 -280
rect 1072 -324 1172 -280
rect 1276 -324 1376 -280
rect 1480 -324 1580 -280
rect 1684 -324 1784 -280
rect 1888 -324 1988 -280
rect 2092 -324 2192 -280
rect 2296 -324 2396 -280
rect 2500 -324 2600 -280
rect 2704 -324 2804 -280
<< metal1 >>
rect -2879 258 -2833 278
rect -2879 -278 -2833 -258
rect -2675 258 -2629 278
rect -2675 -278 -2629 -258
rect -2471 258 -2425 278
rect -2471 -278 -2425 -258
rect -2267 258 -2221 278
rect -2267 -278 -2221 -258
rect -2063 258 -2017 278
rect -2063 -278 -2017 -258
rect -1859 258 -1813 278
rect -1859 -278 -1813 -258
rect -1655 258 -1609 278
rect -1655 -278 -1609 -258
rect -1451 258 -1405 278
rect -1451 -278 -1405 -258
rect -1247 258 -1201 278
rect -1247 -278 -1201 -258
rect -1043 258 -997 278
rect -1043 -278 -997 -258
rect -839 258 -793 278
rect -839 -278 -793 -258
rect -635 258 -589 278
rect -635 -278 -589 -258
rect -431 258 -385 278
rect -431 -278 -385 -258
rect -227 258 -181 278
rect -227 -278 -181 -258
rect -23 258 23 278
rect -23 -278 23 -258
rect 181 258 227 278
rect 181 -278 227 -258
rect 385 258 431 278
rect 385 -278 431 -258
rect 589 258 635 278
rect 589 -278 635 -258
rect 793 258 839 278
rect 793 -278 839 -258
rect 997 258 1043 278
rect 997 -278 1043 -258
rect 1201 258 1247 278
rect 1201 -278 1247 -258
rect 1405 258 1451 278
rect 1405 -278 1451 -258
rect 1609 258 1655 278
rect 1609 -278 1655 -258
rect 1813 258 1859 278
rect 1813 -278 1859 -258
rect 2017 258 2063 278
rect 2017 -278 2063 -258
rect 2221 258 2267 278
rect 2221 -278 2267 -258
rect 2425 258 2471 278
rect 2425 -278 2471 -258
rect 2629 258 2675 278
rect 2629 -278 2675 -258
rect 2833 258 2879 278
rect 2833 -278 2879 -258
<< end >>
