magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2457 -2128 2457 2128
<< nwell >>
rect -457 -128 457 128
<< nsubdiff >>
rect -374 23 374 45
rect -374 -23 -352 23
rect 352 -23 374 23
rect -374 -45 374 -23
<< nsubdiffcont >>
rect -352 -23 352 23
<< metal1 >>
rect -363 23 363 34
rect -363 -23 -352 23
rect 352 -23 363 23
rect -363 -34 363 -23
<< end >>
