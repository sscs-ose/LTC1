* NGSPICE file created from res_48k_mag_flat.ext - technology: gf180mcuC

.subckt res_48k_mag_flat A B VDD
X0 a_364_2267# a_124_124# VDD.t6 ppolyf_u r_width=0.8u r_length=10.2u
X1 a_844_2267# a_604_124# VDD.t8 ppolyf_u r_width=0.8u r_length=10.2u
X2 a_1324_2267# a_1084_124# VDD.t9 ppolyf_u r_width=0.8u r_length=10.2u
X3 a_1804_2267# a_1564_124# VDD.t10 ppolyf_u r_width=0.8u r_length=10.2u
X4 a_1804_2267# a_2044_124# VDD.t5 ppolyf_u r_width=0.8u r_length=10.2u
X5 a_2284_2267# B.t0 VDD.t3 ppolyf_u r_width=0.8u r_length=10.2u
X6 a_844_2267# a_1084_124# VDD.t2 ppolyf_u r_width=0.8u r_length=10.2u
X7 a_1324_2267# a_1564_124# VDD.t0 ppolyf_u r_width=0.8u r_length=10.2u
X8 A.t0 a_124_124# VDD.t4 ppolyf_u r_width=0.8u r_length=10.2u
X9 a_364_2267# a_604_124# VDD.t7 ppolyf_u r_width=0.8u r_length=10.2u
X10 a_2284_2267# a_2044_124# VDD.t1 ppolyf_u r_width=0.8u r_length=10.2u
R0 VDD.t1 VDD.t3 85.9604
R1 VDD.t5 VDD.t1 85.9604
R2 VDD.t10 VDD.t5 85.9604
R3 VDD.t0 VDD.t10 85.9604
R4 VDD.t9 VDD.t0 85.9604
R5 VDD.t2 VDD.t9 85.9604
R6 VDD.t8 VDD.t7 85.9604
R7 VDD.t7 VDD.t6 85.9604
R8 VDD.t6 VDD.t4 85.9604
R9 VDD.n0 VDD.t2 58.3816
R10 VDD.n0 VDD.t8 27.5793
R11 VDD VDD.n2 3.15512
R12 VDD.n2 VDD.n0 3.1505
R13 VDD.n2 VDD.n1 0.320839
R14 B B.t0 7.17944
R15 A A.t0 7.18956
C0 a_1804_2267# a_364_2267# 6.05e-21
C1 a_844_2267# a_1804_2267# 1.62e-20
C2 A VDD 0.178f
C3 a_2044_124# B 0.0759f
C4 VDD a_1324_2267# 0.249f
C5 B VDD 0.252f
C6 A a_364_2267# 0.0615f
C7 B a_1084_124# 3.93e-20
C8 a_604_124# a_1564_124# 7.37e-20
C9 A a_1804_2267# 9.36e-22
C10 a_844_2267# a_1324_2267# 0.0759f
C11 a_604_124# a_124_124# 0.0759f
C12 a_604_124# VDD 0.304f
C13 a_1804_2267# a_1324_2267# 0.0755f
C14 a_2044_124# a_1564_124# 0.0759f
C15 a_1564_124# VDD 0.276f
C16 a_604_124# a_1084_124# 0.0755f
C17 a_124_124# VDD 0.286f
C18 a_2044_124# VDD 0.276f
C19 a_1084_124# a_1564_124# 0.0755f
C20 a_2284_2267# VDD 0.259f
C21 a_1084_124# VDD 0.289f
C22 VDD a_364_2267# 0.25f
C23 a_844_2267# VDD 0.249f
C24 a_1804_2267# VDD 0.249f
C25 a_2284_2267# a_1804_2267# 0.0759f
C26 a_844_2267# a_364_2267# 0.0759f
C27 B VSUBS 0.198f
C28 A VSUBS 0.186f
C29 VDD VSUBS 24.6f
C30 a_2284_2267# VSUBS 0.245f
C31 a_2044_124# VSUBS 0.197f
C32 a_1804_2267# VSUBS 0.224f
C33 a_1564_124# VSUBS 0.197f
C34 a_1324_2267# VSUBS 0.224f
C35 a_1084_124# VSUBS 0.19f
C36 a_844_2267# VSUBS 0.224f
C37 a_604_124# VSUBS 0.182f
C38 a_364_2267# VSUBS 0.227f
C39 a_124_124# VSUBS 0.218f
.ends

