magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1217 -1811 1217 1811
<< metal1 >>
rect -217 805 217 811
rect -217 779 -211 805
rect -185 779 -145 805
rect -119 779 -79 805
rect -53 779 -13 805
rect 13 779 53 805
rect 79 779 119 805
rect 145 779 185 805
rect 211 779 217 805
rect -217 739 217 779
rect -217 713 -211 739
rect -185 713 -145 739
rect -119 713 -79 739
rect -53 713 -13 739
rect 13 713 53 739
rect 79 713 119 739
rect 145 713 185 739
rect 211 713 217 739
rect -217 673 217 713
rect -217 647 -211 673
rect -185 647 -145 673
rect -119 647 -79 673
rect -53 647 -13 673
rect 13 647 53 673
rect 79 647 119 673
rect 145 647 185 673
rect 211 647 217 673
rect -217 607 217 647
rect -217 581 -211 607
rect -185 581 -145 607
rect -119 581 -79 607
rect -53 581 -13 607
rect 13 581 53 607
rect 79 581 119 607
rect 145 581 185 607
rect 211 581 217 607
rect -217 541 217 581
rect -217 515 -211 541
rect -185 515 -145 541
rect -119 515 -79 541
rect -53 515 -13 541
rect 13 515 53 541
rect 79 515 119 541
rect 145 515 185 541
rect 211 515 217 541
rect -217 475 217 515
rect -217 449 -211 475
rect -185 449 -145 475
rect -119 449 -79 475
rect -53 449 -13 475
rect 13 449 53 475
rect 79 449 119 475
rect 145 449 185 475
rect 211 449 217 475
rect -217 409 217 449
rect -217 383 -211 409
rect -185 383 -145 409
rect -119 383 -79 409
rect -53 383 -13 409
rect 13 383 53 409
rect 79 383 119 409
rect 145 383 185 409
rect 211 383 217 409
rect -217 343 217 383
rect -217 317 -211 343
rect -185 317 -145 343
rect -119 317 -79 343
rect -53 317 -13 343
rect 13 317 53 343
rect 79 317 119 343
rect 145 317 185 343
rect 211 317 217 343
rect -217 277 217 317
rect -217 251 -211 277
rect -185 251 -145 277
rect -119 251 -79 277
rect -53 251 -13 277
rect 13 251 53 277
rect 79 251 119 277
rect 145 251 185 277
rect 211 251 217 277
rect -217 211 217 251
rect -217 185 -211 211
rect -185 185 -145 211
rect -119 185 -79 211
rect -53 185 -13 211
rect 13 185 53 211
rect 79 185 119 211
rect 145 185 185 211
rect 211 185 217 211
rect -217 145 217 185
rect -217 119 -211 145
rect -185 119 -145 145
rect -119 119 -79 145
rect -53 119 -13 145
rect 13 119 53 145
rect 79 119 119 145
rect 145 119 185 145
rect 211 119 217 145
rect -217 79 217 119
rect -217 53 -211 79
rect -185 53 -145 79
rect -119 53 -79 79
rect -53 53 -13 79
rect 13 53 53 79
rect 79 53 119 79
rect 145 53 185 79
rect 211 53 217 79
rect -217 13 217 53
rect -217 -13 -211 13
rect -185 -13 -145 13
rect -119 -13 -79 13
rect -53 -13 -13 13
rect 13 -13 53 13
rect 79 -13 119 13
rect 145 -13 185 13
rect 211 -13 217 13
rect -217 -53 217 -13
rect -217 -79 -211 -53
rect -185 -79 -145 -53
rect -119 -79 -79 -53
rect -53 -79 -13 -53
rect 13 -79 53 -53
rect 79 -79 119 -53
rect 145 -79 185 -53
rect 211 -79 217 -53
rect -217 -119 217 -79
rect -217 -145 -211 -119
rect -185 -145 -145 -119
rect -119 -145 -79 -119
rect -53 -145 -13 -119
rect 13 -145 53 -119
rect 79 -145 119 -119
rect 145 -145 185 -119
rect 211 -145 217 -119
rect -217 -185 217 -145
rect -217 -211 -211 -185
rect -185 -211 -145 -185
rect -119 -211 -79 -185
rect -53 -211 -13 -185
rect 13 -211 53 -185
rect 79 -211 119 -185
rect 145 -211 185 -185
rect 211 -211 217 -185
rect -217 -251 217 -211
rect -217 -277 -211 -251
rect -185 -277 -145 -251
rect -119 -277 -79 -251
rect -53 -277 -13 -251
rect 13 -277 53 -251
rect 79 -277 119 -251
rect 145 -277 185 -251
rect 211 -277 217 -251
rect -217 -317 217 -277
rect -217 -343 -211 -317
rect -185 -343 -145 -317
rect -119 -343 -79 -317
rect -53 -343 -13 -317
rect 13 -343 53 -317
rect 79 -343 119 -317
rect 145 -343 185 -317
rect 211 -343 217 -317
rect -217 -383 217 -343
rect -217 -409 -211 -383
rect -185 -409 -145 -383
rect -119 -409 -79 -383
rect -53 -409 -13 -383
rect 13 -409 53 -383
rect 79 -409 119 -383
rect 145 -409 185 -383
rect 211 -409 217 -383
rect -217 -449 217 -409
rect -217 -475 -211 -449
rect -185 -475 -145 -449
rect -119 -475 -79 -449
rect -53 -475 -13 -449
rect 13 -475 53 -449
rect 79 -475 119 -449
rect 145 -475 185 -449
rect 211 -475 217 -449
rect -217 -515 217 -475
rect -217 -541 -211 -515
rect -185 -541 -145 -515
rect -119 -541 -79 -515
rect -53 -541 -13 -515
rect 13 -541 53 -515
rect 79 -541 119 -515
rect 145 -541 185 -515
rect 211 -541 217 -515
rect -217 -581 217 -541
rect -217 -607 -211 -581
rect -185 -607 -145 -581
rect -119 -607 -79 -581
rect -53 -607 -13 -581
rect 13 -607 53 -581
rect 79 -607 119 -581
rect 145 -607 185 -581
rect 211 -607 217 -581
rect -217 -647 217 -607
rect -217 -673 -211 -647
rect -185 -673 -145 -647
rect -119 -673 -79 -647
rect -53 -673 -13 -647
rect 13 -673 53 -647
rect 79 -673 119 -647
rect 145 -673 185 -647
rect 211 -673 217 -647
rect -217 -713 217 -673
rect -217 -739 -211 -713
rect -185 -739 -145 -713
rect -119 -739 -79 -713
rect -53 -739 -13 -713
rect 13 -739 53 -713
rect 79 -739 119 -713
rect 145 -739 185 -713
rect 211 -739 217 -713
rect -217 -779 217 -739
rect -217 -805 -211 -779
rect -185 -805 -145 -779
rect -119 -805 -79 -779
rect -53 -805 -13 -779
rect 13 -805 53 -779
rect 79 -805 119 -779
rect 145 -805 185 -779
rect 211 -805 217 -779
rect -217 -811 217 -805
<< via1 >>
rect -211 779 -185 805
rect -145 779 -119 805
rect -79 779 -53 805
rect -13 779 13 805
rect 53 779 79 805
rect 119 779 145 805
rect 185 779 211 805
rect -211 713 -185 739
rect -145 713 -119 739
rect -79 713 -53 739
rect -13 713 13 739
rect 53 713 79 739
rect 119 713 145 739
rect 185 713 211 739
rect -211 647 -185 673
rect -145 647 -119 673
rect -79 647 -53 673
rect -13 647 13 673
rect 53 647 79 673
rect 119 647 145 673
rect 185 647 211 673
rect -211 581 -185 607
rect -145 581 -119 607
rect -79 581 -53 607
rect -13 581 13 607
rect 53 581 79 607
rect 119 581 145 607
rect 185 581 211 607
rect -211 515 -185 541
rect -145 515 -119 541
rect -79 515 -53 541
rect -13 515 13 541
rect 53 515 79 541
rect 119 515 145 541
rect 185 515 211 541
rect -211 449 -185 475
rect -145 449 -119 475
rect -79 449 -53 475
rect -13 449 13 475
rect 53 449 79 475
rect 119 449 145 475
rect 185 449 211 475
rect -211 383 -185 409
rect -145 383 -119 409
rect -79 383 -53 409
rect -13 383 13 409
rect 53 383 79 409
rect 119 383 145 409
rect 185 383 211 409
rect -211 317 -185 343
rect -145 317 -119 343
rect -79 317 -53 343
rect -13 317 13 343
rect 53 317 79 343
rect 119 317 145 343
rect 185 317 211 343
rect -211 251 -185 277
rect -145 251 -119 277
rect -79 251 -53 277
rect -13 251 13 277
rect 53 251 79 277
rect 119 251 145 277
rect 185 251 211 277
rect -211 185 -185 211
rect -145 185 -119 211
rect -79 185 -53 211
rect -13 185 13 211
rect 53 185 79 211
rect 119 185 145 211
rect 185 185 211 211
rect -211 119 -185 145
rect -145 119 -119 145
rect -79 119 -53 145
rect -13 119 13 145
rect 53 119 79 145
rect 119 119 145 145
rect 185 119 211 145
rect -211 53 -185 79
rect -145 53 -119 79
rect -79 53 -53 79
rect -13 53 13 79
rect 53 53 79 79
rect 119 53 145 79
rect 185 53 211 79
rect -211 -13 -185 13
rect -145 -13 -119 13
rect -79 -13 -53 13
rect -13 -13 13 13
rect 53 -13 79 13
rect 119 -13 145 13
rect 185 -13 211 13
rect -211 -79 -185 -53
rect -145 -79 -119 -53
rect -79 -79 -53 -53
rect -13 -79 13 -53
rect 53 -79 79 -53
rect 119 -79 145 -53
rect 185 -79 211 -53
rect -211 -145 -185 -119
rect -145 -145 -119 -119
rect -79 -145 -53 -119
rect -13 -145 13 -119
rect 53 -145 79 -119
rect 119 -145 145 -119
rect 185 -145 211 -119
rect -211 -211 -185 -185
rect -145 -211 -119 -185
rect -79 -211 -53 -185
rect -13 -211 13 -185
rect 53 -211 79 -185
rect 119 -211 145 -185
rect 185 -211 211 -185
rect -211 -277 -185 -251
rect -145 -277 -119 -251
rect -79 -277 -53 -251
rect -13 -277 13 -251
rect 53 -277 79 -251
rect 119 -277 145 -251
rect 185 -277 211 -251
rect -211 -343 -185 -317
rect -145 -343 -119 -317
rect -79 -343 -53 -317
rect -13 -343 13 -317
rect 53 -343 79 -317
rect 119 -343 145 -317
rect 185 -343 211 -317
rect -211 -409 -185 -383
rect -145 -409 -119 -383
rect -79 -409 -53 -383
rect -13 -409 13 -383
rect 53 -409 79 -383
rect 119 -409 145 -383
rect 185 -409 211 -383
rect -211 -475 -185 -449
rect -145 -475 -119 -449
rect -79 -475 -53 -449
rect -13 -475 13 -449
rect 53 -475 79 -449
rect 119 -475 145 -449
rect 185 -475 211 -449
rect -211 -541 -185 -515
rect -145 -541 -119 -515
rect -79 -541 -53 -515
rect -13 -541 13 -515
rect 53 -541 79 -515
rect 119 -541 145 -515
rect 185 -541 211 -515
rect -211 -607 -185 -581
rect -145 -607 -119 -581
rect -79 -607 -53 -581
rect -13 -607 13 -581
rect 53 -607 79 -581
rect 119 -607 145 -581
rect 185 -607 211 -581
rect -211 -673 -185 -647
rect -145 -673 -119 -647
rect -79 -673 -53 -647
rect -13 -673 13 -647
rect 53 -673 79 -647
rect 119 -673 145 -647
rect 185 -673 211 -647
rect -211 -739 -185 -713
rect -145 -739 -119 -713
rect -79 -739 -53 -713
rect -13 -739 13 -713
rect 53 -739 79 -713
rect 119 -739 145 -713
rect 185 -739 211 -713
rect -211 -805 -185 -779
rect -145 -805 -119 -779
rect -79 -805 -53 -779
rect -13 -805 13 -779
rect 53 -805 79 -779
rect 119 -805 145 -779
rect 185 -805 211 -779
<< metal2 >>
rect -217 805 217 811
rect -217 779 -211 805
rect -185 779 -145 805
rect -119 779 -79 805
rect -53 779 -13 805
rect 13 779 53 805
rect 79 779 119 805
rect 145 779 185 805
rect 211 779 217 805
rect -217 739 217 779
rect -217 713 -211 739
rect -185 713 -145 739
rect -119 713 -79 739
rect -53 713 -13 739
rect 13 713 53 739
rect 79 713 119 739
rect 145 713 185 739
rect 211 713 217 739
rect -217 673 217 713
rect -217 647 -211 673
rect -185 647 -145 673
rect -119 647 -79 673
rect -53 647 -13 673
rect 13 647 53 673
rect 79 647 119 673
rect 145 647 185 673
rect 211 647 217 673
rect -217 607 217 647
rect -217 581 -211 607
rect -185 581 -145 607
rect -119 581 -79 607
rect -53 581 -13 607
rect 13 581 53 607
rect 79 581 119 607
rect 145 581 185 607
rect 211 581 217 607
rect -217 541 217 581
rect -217 515 -211 541
rect -185 515 -145 541
rect -119 515 -79 541
rect -53 515 -13 541
rect 13 515 53 541
rect 79 515 119 541
rect 145 515 185 541
rect 211 515 217 541
rect -217 475 217 515
rect -217 449 -211 475
rect -185 449 -145 475
rect -119 449 -79 475
rect -53 449 -13 475
rect 13 449 53 475
rect 79 449 119 475
rect 145 449 185 475
rect 211 449 217 475
rect -217 409 217 449
rect -217 383 -211 409
rect -185 383 -145 409
rect -119 383 -79 409
rect -53 383 -13 409
rect 13 383 53 409
rect 79 383 119 409
rect 145 383 185 409
rect 211 383 217 409
rect -217 343 217 383
rect -217 317 -211 343
rect -185 317 -145 343
rect -119 317 -79 343
rect -53 317 -13 343
rect 13 317 53 343
rect 79 317 119 343
rect 145 317 185 343
rect 211 317 217 343
rect -217 277 217 317
rect -217 251 -211 277
rect -185 251 -145 277
rect -119 251 -79 277
rect -53 251 -13 277
rect 13 251 53 277
rect 79 251 119 277
rect 145 251 185 277
rect 211 251 217 277
rect -217 211 217 251
rect -217 185 -211 211
rect -185 185 -145 211
rect -119 185 -79 211
rect -53 185 -13 211
rect 13 185 53 211
rect 79 185 119 211
rect 145 185 185 211
rect 211 185 217 211
rect -217 145 217 185
rect -217 119 -211 145
rect -185 119 -145 145
rect -119 119 -79 145
rect -53 119 -13 145
rect 13 119 53 145
rect 79 119 119 145
rect 145 119 185 145
rect 211 119 217 145
rect -217 79 217 119
rect -217 53 -211 79
rect -185 53 -145 79
rect -119 53 -79 79
rect -53 53 -13 79
rect 13 53 53 79
rect 79 53 119 79
rect 145 53 185 79
rect 211 53 217 79
rect -217 13 217 53
rect -217 -13 -211 13
rect -185 -13 -145 13
rect -119 -13 -79 13
rect -53 -13 -13 13
rect 13 -13 53 13
rect 79 -13 119 13
rect 145 -13 185 13
rect 211 -13 217 13
rect -217 -53 217 -13
rect -217 -79 -211 -53
rect -185 -79 -145 -53
rect -119 -79 -79 -53
rect -53 -79 -13 -53
rect 13 -79 53 -53
rect 79 -79 119 -53
rect 145 -79 185 -53
rect 211 -79 217 -53
rect -217 -119 217 -79
rect -217 -145 -211 -119
rect -185 -145 -145 -119
rect -119 -145 -79 -119
rect -53 -145 -13 -119
rect 13 -145 53 -119
rect 79 -145 119 -119
rect 145 -145 185 -119
rect 211 -145 217 -119
rect -217 -185 217 -145
rect -217 -211 -211 -185
rect -185 -211 -145 -185
rect -119 -211 -79 -185
rect -53 -211 -13 -185
rect 13 -211 53 -185
rect 79 -211 119 -185
rect 145 -211 185 -185
rect 211 -211 217 -185
rect -217 -251 217 -211
rect -217 -277 -211 -251
rect -185 -277 -145 -251
rect -119 -277 -79 -251
rect -53 -277 -13 -251
rect 13 -277 53 -251
rect 79 -277 119 -251
rect 145 -277 185 -251
rect 211 -277 217 -251
rect -217 -317 217 -277
rect -217 -343 -211 -317
rect -185 -343 -145 -317
rect -119 -343 -79 -317
rect -53 -343 -13 -317
rect 13 -343 53 -317
rect 79 -343 119 -317
rect 145 -343 185 -317
rect 211 -343 217 -317
rect -217 -383 217 -343
rect -217 -409 -211 -383
rect -185 -409 -145 -383
rect -119 -409 -79 -383
rect -53 -409 -13 -383
rect 13 -409 53 -383
rect 79 -409 119 -383
rect 145 -409 185 -383
rect 211 -409 217 -383
rect -217 -449 217 -409
rect -217 -475 -211 -449
rect -185 -475 -145 -449
rect -119 -475 -79 -449
rect -53 -475 -13 -449
rect 13 -475 53 -449
rect 79 -475 119 -449
rect 145 -475 185 -449
rect 211 -475 217 -449
rect -217 -515 217 -475
rect -217 -541 -211 -515
rect -185 -541 -145 -515
rect -119 -541 -79 -515
rect -53 -541 -13 -515
rect 13 -541 53 -515
rect 79 -541 119 -515
rect 145 -541 185 -515
rect 211 -541 217 -515
rect -217 -581 217 -541
rect -217 -607 -211 -581
rect -185 -607 -145 -581
rect -119 -607 -79 -581
rect -53 -607 -13 -581
rect 13 -607 53 -581
rect 79 -607 119 -581
rect 145 -607 185 -581
rect 211 -607 217 -581
rect -217 -647 217 -607
rect -217 -673 -211 -647
rect -185 -673 -145 -647
rect -119 -673 -79 -647
rect -53 -673 -13 -647
rect 13 -673 53 -647
rect 79 -673 119 -647
rect 145 -673 185 -647
rect 211 -673 217 -647
rect -217 -713 217 -673
rect -217 -739 -211 -713
rect -185 -739 -145 -713
rect -119 -739 -79 -713
rect -53 -739 -13 -713
rect 13 -739 53 -713
rect 79 -739 119 -713
rect 145 -739 185 -713
rect 211 -739 217 -713
rect -217 -779 217 -739
rect -217 -805 -211 -779
rect -185 -805 -145 -779
rect -119 -805 -79 -779
rect -53 -805 -13 -779
rect 13 -805 53 -779
rect 79 -805 119 -779
rect 145 -805 185 -779
rect 211 -805 217 -779
rect -217 -811 217 -805
<< end >>
