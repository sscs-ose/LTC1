magic
tech gf180mcuC
magscale 1 10
timestamp 1694584912
<< nwell >>
rect -62 668 502 818
rect 243 394 306 398
rect 38 393 127 394
rect 38 332 125 393
rect 243 392 403 394
rect 310 379 476 380
rect 310 352 502 379
rect 272 348 502 352
rect 272 346 328 348
rect 357 346 502 348
rect 112 322 122 332
rect 310 328 502 346
<< pwell >>
rect 229 280 289 281
rect 229 221 292 280
rect 87 211 218 212
rect 303 211 416 212
<< psubdiff >>
rect -50 -26 504 -10
rect -50 -74 -19 -26
rect 450 -74 504 -26
rect -50 -92 504 -74
<< nsubdiff >>
rect 16 772 422 792
rect 16 716 53 772
rect 365 716 422 772
rect 16 695 422 716
<< psubdiffcont >>
rect -19 -74 450 -26
<< nsubdiffcont >>
rect 53 716 365 772
<< polysilicon >>
rect 38 380 168 394
rect 38 321 52 380
rect 115 321 168 380
rect 38 306 168 321
rect 112 212 168 306
rect 272 293 328 394
rect 216 280 328 293
rect 216 221 229 280
rect 292 221 328 280
rect 216 212 328 221
rect 216 208 303 212
<< polycontact >>
rect 52 321 115 380
rect 229 221 292 280
<< metal1 >>
rect -62 772 502 818
rect -62 716 53 772
rect 365 716 502 772
rect -62 668 502 716
rect 34 449 85 668
rect 209 447 230 454
rect 197 440 242 447
rect 357 440 403 668
rect 197 398 243 440
rect 197 394 306 398
rect 38 380 127 394
rect 38 352 52 380
rect -63 321 52 352
rect 115 321 127 380
rect 197 352 502 394
rect 273 348 502 352
rect -63 306 127 321
rect 218 280 303 291
rect 218 258 229 280
rect -61 221 229 258
rect 292 221 303 280
rect -61 212 303 221
rect 37 1 83 166
rect 184 67 251 165
rect 357 70 403 348
rect -86 -26 530 1
rect -86 -74 -19 -26
rect 450 -74 530 -26
rect -86 -97 530 -74
use nmos_3p3_HZS5UA  nmos_3p3_HZS5UA_0
timestamp 1690264421
transform 1 0 300 0 1 118
box -140 -118 140 118
use nmos_3p3_HZS5UA  nmos_3p3_HZS5UA_1
timestamp 1690264421
transform 1 0 140 0 1 118
box -140 -118 140 118
use pmos_3p3_M8RWPS  pmos_3p3_M8RWPS_0
timestamp 1692705520
transform -1 0 300 0 1 488
box -202 -180 202 180
use pmos_3p3_M8RWPS  pmos_3p3_M8RWPS_1
timestamp 1692705520
transform 1 0 140 0 1 488
box -202 -180 202 180
<< labels >>
flabel nsubdiffcont 207 744 207 744 0 FreeSans 320 0 0 0 VDD
port 0 nsew
flabel psubdiffcont 216 -48 216 -48 0 FreeSans 320 0 0 0 VSS
port 1 nsew
flabel metal1 -33 330 -33 330 0 FreeSans 480 0 0 0 B
port 2 nsew
flabel metal1 -30 232 -30 232 0 FreeSans 480 0 0 0 A
port 3 nsew
flabel metal1 469 376 469 376 0 FreeSans 480 0 0 0 OUT
port 4 nsew
flabel metal1 218 109 218 109 0 FreeSans 480 0 0 0 SD
port 5 nsew
<< end >>
