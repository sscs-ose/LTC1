magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2045 -3972 2045 3972
<< psubdiff >>
rect -45 1950 45 1972
rect -45 -1950 -23 1950
rect 23 -1950 45 1950
rect -45 -1972 45 -1950
<< psubdiffcont >>
rect -23 -1950 23 1950
<< metal1 >>
rect -34 1950 34 1961
rect -34 -1950 -23 1950
rect 23 -1950 34 1950
rect -34 -1961 34 -1950
<< end >>
