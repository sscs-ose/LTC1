magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2461 -2097 2461 2097
<< psubdiff >>
rect -461 75 461 97
rect -461 29 -439 75
rect -393 29 -335 75
rect -289 29 -231 75
rect -185 29 -127 75
rect -81 29 -23 75
rect 23 29 81 75
rect 127 29 185 75
rect 231 29 289 75
rect 335 29 393 75
rect 439 29 461 75
rect -461 -29 461 29
rect -461 -75 -439 -29
rect -393 -75 -335 -29
rect -289 -75 -231 -29
rect -185 -75 -127 -29
rect -81 -75 -23 -29
rect 23 -75 81 -29
rect 127 -75 185 -29
rect 231 -75 289 -29
rect 335 -75 393 -29
rect 439 -75 461 -29
rect -461 -97 461 -75
<< psubdiffcont >>
rect -439 29 -393 75
rect -335 29 -289 75
rect -231 29 -185 75
rect -127 29 -81 75
rect -23 29 23 75
rect 81 29 127 75
rect 185 29 231 75
rect 289 29 335 75
rect 393 29 439 75
rect -439 -75 -393 -29
rect -335 -75 -289 -29
rect -231 -75 -185 -29
rect -127 -75 -81 -29
rect -23 -75 23 -29
rect 81 -75 127 -29
rect 185 -75 231 -29
rect 289 -75 335 -29
rect 393 -75 439 -29
<< metal1 >>
rect -450 75 450 86
rect -450 29 -439 75
rect -393 29 -335 75
rect -289 29 -231 75
rect -185 29 -127 75
rect -81 29 -23 75
rect 23 29 81 75
rect 127 29 185 75
rect 231 29 289 75
rect 335 29 393 75
rect 439 29 450 75
rect -450 -29 450 29
rect -450 -75 -439 -29
rect -393 -75 -335 -29
rect -289 -75 -231 -29
rect -185 -75 -127 -29
rect -81 -75 -23 -29
rect 23 -75 81 -29
rect 127 -75 185 -29
rect 231 -75 289 -29
rect 335 -75 393 -29
rect 439 -75 450 -29
rect -450 -86 450 -75
<< end >>
