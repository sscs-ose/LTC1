magic
tech gf180mcuC
magscale 1 10
timestamp 1692057126
<< nwell >>
rect -224 -410 224 410
<< pmos >>
rect -50 -280 50 280
<< pdiff >>
rect -138 267 -50 280
rect -138 -267 -125 267
rect -79 -267 -50 267
rect -138 -280 -50 -267
rect 50 267 138 280
rect 50 -267 79 267
rect 125 -267 138 267
rect 50 -280 138 -267
<< pdiffc >>
rect -125 -267 -79 267
rect 79 -267 125 267
<< polysilicon >>
rect -50 280 50 324
rect -50 -324 50 -280
<< metal1 >>
rect -125 267 -79 278
rect -125 -278 -79 -267
rect 79 267 125 278
rect 79 -278 125 -267
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 2.8 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
