magic
tech gf180mcuC
magscale 1 10
timestamp 1698511765
<< pwell >>
rect 7871 -745 7937 -717
<< polysilicon >>
rect 7863 -679 7935 -671
rect 7861 -684 7937 -679
rect 7861 -730 7876 -684
rect 7922 -730 7937 -684
rect 7861 -735 7937 -730
rect 7863 -743 7935 -735
<< polycontact >>
rect 7876 -730 7922 -684
<< metal1 >>
rect -1039 2772 10 2884
rect -16 2440 60 2452
rect -16 2437 -4 2440
rect -749 2391 -4 2437
rect -16 2388 -4 2391
rect 48 2388 60 2440
rect -16 2376 60 2388
rect -138 1558 -62 1570
rect -138 1555 -126 1558
rect -866 1509 -126 1555
rect -138 1506 -126 1509
rect -74 1506 -62 1558
rect -138 1494 -62 1506
rect 254 1389 330 1401
rect 254 1337 266 1389
rect 318 1337 330 1389
rect 10886 1389 10962 1401
rect 5391 1340 5825 1386
rect 254 1325 330 1337
rect 10886 1337 10898 1389
rect 10950 1337 10962 1389
rect 11373 1389 11449 1401
rect 11373 1386 11385 1389
rect 10987 1340 11385 1386
rect 10886 1325 10962 1337
rect 11373 1337 11385 1340
rect 11437 1337 11449 1389
rect 11373 1325 11449 1337
rect -261 730 -185 742
rect -261 727 -249 730
rect -843 681 -249 727
rect -261 678 -249 681
rect -197 678 -185 730
rect -261 666 -185 678
rect 7871 530 7927 532
rect 7861 477 7873 530
rect 7925 477 7937 530
rect 7871 475 7927 477
rect -261 -152 -185 -140
rect -261 -155 -249 -152
rect -743 -201 -249 -155
rect -261 -204 -249 -201
rect -197 -204 -185 -152
rect -261 -216 -185 -204
rect 7865 -680 7933 -673
rect 7861 -733 7873 -680
rect 7925 -733 7937 -680
rect 7865 -741 7933 -733
rect -393 -980 -317 -968
rect -393 -983 -381 -980
rect -764 -1029 -381 -983
rect -393 -1032 -381 -1029
rect -329 -1032 -317 -980
rect -393 -1044 -317 -1032
rect 254 -1541 330 -1529
rect 254 -1593 266 -1541
rect 318 -1593 330 -1541
rect 10886 -1541 10962 -1529
rect 5391 -1590 5834 -1544
rect 254 -1605 330 -1593
rect 10886 -1593 10898 -1541
rect 10950 -1593 10962 -1541
rect 10886 -1605 10962 -1593
rect -526 -1862 -450 -1850
rect -526 -1865 -514 -1862
rect -843 -1911 -514 -1865
rect -526 -1914 -514 -1911
rect -462 -1914 -450 -1862
rect -526 -1926 -450 -1914
rect -1440 -3088 136 -2976
rect 254 -4471 330 -4459
rect 254 -4523 266 -4471
rect 318 -4523 330 -4471
rect 10886 -4471 10962 -4459
rect 5393 -4520 5824 -4474
rect 254 -4535 330 -4523
rect 10886 -4523 10898 -4471
rect 10950 -4523 10962 -4471
rect 10886 -4535 10962 -4523
rect 11373 -4578 11449 -4566
rect 11373 -4581 11385 -4578
rect 10572 -4627 11385 -4581
rect 11373 -4630 11385 -4627
rect 11437 -4630 11449 -4578
rect 11373 -4642 11449 -4630
rect -393 -5329 -317 -5317
rect -393 -5332 -381 -5329
rect -1489 -5378 -381 -5332
rect -393 -5381 -381 -5378
rect -329 -5381 -317 -5329
rect -393 -5393 -317 -5381
rect -1440 -6018 10 -5906
<< via1 >>
rect -4 2388 48 2440
rect -126 1506 -74 1558
rect 266 1337 318 1389
rect 10898 1337 10950 1389
rect 11385 1337 11437 1389
rect -249 678 -197 730
rect 2275 477 2327 529
rect 7873 477 7925 530
rect -249 -204 -197 -152
rect 2275 -733 2327 -681
rect 7873 -684 7925 -680
rect 7873 -730 7876 -684
rect 7876 -730 7922 -684
rect 7922 -730 7925 -684
rect 7873 -733 7925 -730
rect -381 -1032 -329 -980
rect 266 -1593 318 -1541
rect 10898 -1593 10950 -1541
rect -514 -1914 -462 -1862
rect 266 -4523 318 -4471
rect 10898 -4523 10950 -4471
rect 11385 -4630 11437 -4578
rect -6545 -5383 -6493 -5331
rect -381 -5381 -329 -5329
rect 2275 -5383 2327 -5331
rect 8889 -5383 8941 -5331
<< metal2 >>
rect -16 2440 60 2452
rect -16 2388 -4 2440
rect 48 2388 60 2440
rect -16 2376 60 2388
rect -138 1558 -62 1570
rect -138 1506 -126 1558
rect -74 1506 -62 1558
rect -138 1494 -62 1506
rect -261 732 -185 742
rect -261 676 -251 732
rect -195 676 -185 732
rect -261 666 -185 676
rect -261 -152 -185 -140
rect -261 -204 -249 -152
rect -197 -204 -185 -152
rect -261 -216 -185 -204
rect -393 -980 -317 -968
rect -393 -1032 -381 -980
rect -329 -1032 -317 -980
rect -393 -1044 -317 -1032
rect -526 -1862 -450 -1850
rect -526 -1914 -514 -1862
rect -462 -1914 -450 -1862
rect -526 -1926 -450 -1914
rect -516 -5319 -460 -1926
rect -383 -5317 -327 -1044
rect -6557 -5329 -6481 -5319
rect -6557 -5385 -6547 -5329
rect -6491 -5385 -6481 -5329
rect -6557 -5395 -6481 -5385
rect -526 -5329 -450 -5319
rect -526 -5385 -516 -5329
rect -460 -5385 -450 -5329
rect -526 -5395 -450 -5385
rect -393 -5329 -317 -5317
rect -251 -5319 -195 -216
rect -128 -669 -72 1494
rect -6 541 50 2376
rect 254 1391 330 1401
rect 254 1335 264 1391
rect 320 1335 330 1391
rect 254 1325 330 1335
rect 10886 1391 10962 1401
rect 10886 1335 10896 1391
rect 10952 1335 10962 1391
rect 10886 1325 10962 1335
rect 11373 1389 11449 1401
rect 11373 1337 11385 1389
rect 11437 1337 11449 1389
rect 11373 1325 11449 1337
rect 8877 732 8953 742
rect 8877 676 8887 732
rect 8943 676 8953 732
rect 8877 666 8953 676
rect -16 531 60 541
rect -16 475 -6 531
rect 50 475 60 531
rect -16 465 60 475
rect 2263 531 2339 541
rect 2263 475 2273 531
rect 2329 475 2339 531
rect 2263 465 2339 475
rect 7861 530 7937 542
rect 7861 477 7873 530
rect 7925 477 7937 530
rect 7861 465 7937 477
rect 2273 -669 2329 465
rect 7871 -668 7927 465
rect -138 -679 -62 -669
rect -138 -735 -128 -679
rect -72 -735 -62 -679
rect -138 -745 -62 -735
rect 2263 -681 2339 -669
rect 2263 -733 2275 -681
rect 2327 -733 2339 -681
rect 2263 -745 2339 -733
rect 7861 -678 7937 -668
rect 7861 -735 7871 -678
rect 7927 -735 7937 -678
rect 7861 -745 7937 -735
rect 254 -1539 330 -1529
rect 254 -1595 264 -1539
rect 320 -1595 330 -1539
rect 254 -1605 330 -1595
rect 254 -4469 330 -4459
rect 254 -4525 264 -4469
rect 320 -4525 330 -4469
rect 254 -4535 330 -4525
rect 8887 -5319 8943 666
rect 10886 -1539 10962 -1529
rect 10886 -1595 10896 -1539
rect 10952 -1595 10962 -1539
rect 10886 -1605 10962 -1595
rect 10886 -4469 10962 -4459
rect 10886 -4525 10896 -4469
rect 10952 -4525 10962 -4469
rect 10886 -4535 10962 -4525
rect 11383 -4566 11439 1325
rect 11373 -4578 11449 -4566
rect 11373 -4630 11385 -4578
rect 11437 -4630 11449 -4578
rect 11373 -4642 11449 -4630
rect -393 -5381 -381 -5329
rect -329 -5381 -317 -5329
rect -393 -5393 -317 -5381
rect -261 -5329 -185 -5319
rect -261 -5385 -251 -5329
rect -195 -5385 -185 -5329
rect -261 -5395 -185 -5385
rect 2263 -5329 2339 -5319
rect 2263 -5385 2273 -5329
rect 2329 -5385 2339 -5329
rect 2263 -5395 2339 -5385
rect 8877 -5331 8953 -5319
rect 8877 -5383 8889 -5331
rect 8941 -5383 8953 -5331
rect 8877 -5395 8953 -5383
<< via2 >>
rect -251 730 -195 732
rect -251 678 -249 730
rect -249 678 -197 730
rect -197 678 -195 730
rect -251 676 -195 678
rect -6547 -5331 -6491 -5329
rect -6547 -5383 -6545 -5331
rect -6545 -5383 -6493 -5331
rect -6493 -5383 -6491 -5331
rect -6547 -5385 -6491 -5383
rect -516 -5385 -460 -5329
rect 264 1389 320 1391
rect 264 1337 266 1389
rect 266 1337 318 1389
rect 318 1337 320 1389
rect 264 1335 320 1337
rect 10896 1389 10952 1391
rect 10896 1337 10898 1389
rect 10898 1337 10950 1389
rect 10950 1337 10952 1389
rect 10896 1335 10952 1337
rect 8887 676 8943 732
rect -6 475 50 531
rect 2273 529 2329 531
rect 2273 477 2275 529
rect 2275 477 2327 529
rect 2327 477 2329 529
rect 2273 475 2329 477
rect -128 -735 -72 -679
rect 7871 -680 7927 -678
rect 7871 -733 7873 -680
rect 7873 -733 7925 -680
rect 7925 -733 7927 -680
rect 7871 -735 7927 -733
rect 264 -1541 320 -1539
rect 264 -1593 266 -1541
rect 266 -1593 318 -1541
rect 318 -1593 320 -1541
rect 264 -1595 320 -1593
rect 264 -4471 320 -4469
rect 264 -4523 266 -4471
rect 266 -4523 318 -4471
rect 318 -4523 320 -4471
rect 264 -4525 320 -4523
rect 10896 -1541 10952 -1539
rect 10896 -1593 10898 -1541
rect 10898 -1593 10950 -1541
rect 10950 -1593 10952 -1541
rect 10896 -1595 10952 -1593
rect 10896 -4471 10952 -4469
rect 10896 -4523 10898 -4471
rect 10898 -4523 10950 -4471
rect 10950 -4523 10952 -4471
rect 10896 -4525 10952 -4523
rect -251 -5385 -195 -5329
rect 2273 -5331 2329 -5329
rect 2273 -5383 2275 -5331
rect 2275 -5383 2327 -5331
rect 2327 -5383 2329 -5331
rect 2273 -5385 2329 -5383
<< metal3 >>
rect 254 1391 330 1401
rect 10886 1391 10962 1401
rect 254 1335 264 1391
rect 320 1335 10896 1391
rect 10952 1335 10962 1391
rect 254 1325 330 1335
rect 10886 1325 10962 1335
rect -261 732 -185 742
rect 8877 732 8953 742
rect -261 676 -251 732
rect -195 676 8887 732
rect 8943 676 8953 732
rect -261 666 -185 676
rect 8877 666 8953 676
rect -16 531 60 541
rect 2263 531 2339 541
rect -16 475 -6 531
rect 50 475 2273 531
rect 2329 475 2339 531
rect -16 465 60 475
rect 2263 465 2339 475
rect -138 -679 -62 -669
rect 7861 -678 7937 -668
rect 7861 -679 7871 -678
rect -138 -735 -128 -679
rect -72 -735 7871 -679
rect 7927 -735 7937 -678
rect -138 -745 -62 -735
rect 7861 -745 7937 -735
rect 254 -1539 330 -1529
rect 10886 -1539 10962 -1529
rect 254 -1595 264 -1539
rect 320 -1595 10896 -1539
rect 10952 -1595 10962 -1539
rect 254 -1605 330 -1595
rect 10886 -1605 10962 -1595
rect 254 -4469 330 -4459
rect 10886 -4469 10962 -4459
rect 254 -4525 264 -4469
rect 320 -4525 10896 -4469
rect 10952 -4525 10962 -4469
rect 254 -4535 330 -4525
rect 10886 -4535 10962 -4525
rect -6557 -5329 -6481 -5319
rect -526 -5329 -450 -5319
rect -6557 -5385 -6547 -5329
rect -6491 -5385 -516 -5329
rect -460 -5385 -450 -5329
rect -6557 -5395 -6481 -5385
rect -526 -5395 -450 -5385
rect -261 -5329 -185 -5319
rect 2263 -5329 2339 -5319
rect -261 -5385 -251 -5329
rect -195 -5385 2273 -5329
rect 2329 -5385 2339 -5329
rect -261 -5395 -185 -5385
rect 2263 -5395 2339 -5385
use Non_Ovl_CLK_Gen_Layout  Non_Ovl_CLK_Gen_Layout_0 ~/GF180Projects/Tapeout/Magic/Non_Ovl_CLK_Gen
timestamp 1698511765
transform 1 0 -3813 0 1 -1503
box -1478 -868 3162 980
use Non_Ovl_CLK_Gen_Layout  Non_Ovl_CLK_Gen_Layout_1
timestamp 1698511765
transform 1 0 -3813 0 1 1917
box -1478 -868 3162 980
use Non_Ovl_CLK_Gen_Layout  Non_Ovl_CLK_Gen_Layout_2
timestamp 1698511765
transform 1 0 -3813 0 -1 319
box -1478 -868 3162 980
use TG_Layout  TG_Layout_0 ~/GF180Projects/Tapeout/Magic/Logic_Gates/Transmission_Gate
timestamp 1698511765
transform 1 0 8341 0 1 -6
box 45 -152 2865 2894
use TG_Layout  TG_Layout_1
timestamp 1698511765
transform 1 0 8341 0 -1 -198
box 45 -152 2865 2894
use TG_Layout  TG_Layout_2
timestamp 1698511765
transform -1 0 8473 0 1 -6
box 45 -152 2865 2894
use TG_Layout  TG_Layout_3
timestamp 1698511765
transform -1 0 8473 0 -1 -198
box 45 -152 2865 2894
use TG_Layout  TG_Layout_4
timestamp 1698511765
transform 1 0 8341 0 1 -5866
box 45 -152 2865 2894
use TG_Layout  TG_Layout_5
timestamp 1698511765
transform -1 0 2875 0 1 -6
box 45 -152 2865 2894
use TG_Layout  TG_Layout_6
timestamp 1698511765
transform 1 0 2743 0 -1 -198
box 45 -152 2865 2894
use TG_Layout  TG_Layout_7
timestamp 1698511765
transform 1 0 2743 0 1 -6
box 45 -152 2865 2894
use TG_Layout  TG_Layout_8
timestamp 1698511765
transform -1 0 2875 0 -1 -198
box 45 -152 2865 2894
use TG_Layout  TG_Layout_9
timestamp 1698511765
transform -1 0 2875 0 1 -5866
box 45 -152 2865 2894
use TG_Layout  TG_Layout_10
timestamp 1698511765
transform 1 0 2743 0 1 -5866
box 45 -152 2865 2894
use TG_Layout  TG_Layout_11
timestamp 1698511765
transform -1 0 8473 0 1 -5866
box 45 -152 2865 2894
use TG_Layout  TG_Layout_12
timestamp 1698511765
transform -1 0 -1379 0 1 -5866
box 45 -152 2865 2894
use TG_Layout  TG_Layout_13
timestamp 1698511765
transform 1 0 -7093 0 1 -5866
box 45 -152 2865 2894
<< end >>
