magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect 11097 11097 73000 73000
<< psubdiff >>
rect 69813 70674 69968 71000
rect 70671 69774 71000 69968
rect 70802 69642 71000 69774
rect 13097 44921 13291 45178
tri 13291 44921 13295 44925 sw
rect 13097 44913 13295 44921
tri 13295 44913 13303 44921 sw
rect 13097 44905 13303 44913
tri 13303 44905 13311 44913 sw
rect 13097 44897 13311 44905
tri 13311 44897 13319 44905 sw
rect 13097 44889 13319 44897
tri 13319 44889 13327 44897 sw
rect 13097 44881 13327 44889
tri 13327 44881 13335 44889 sw
rect 13097 44873 13335 44881
tri 13335 44873 13343 44881 sw
rect 13097 44865 13343 44873
tri 13343 44865 13351 44873 sw
rect 13097 44857 13351 44865
tri 13351 44857 13359 44865 sw
rect 13097 44849 13359 44857
tri 13359 44849 13367 44857 sw
rect 13097 44843 13367 44849
tri 13097 44839 13101 44843 ne
rect 13101 44841 13367 44843
tri 13367 44841 13375 44849 sw
rect 13101 44839 13375 44841
tri 13101 44831 13109 44839 ne
rect 13109 44833 13375 44839
tri 13375 44833 13383 44841 sw
rect 13109 44831 13383 44833
tri 13109 44823 13117 44831 ne
rect 13117 44825 13383 44831
tri 13383 44825 13391 44833 sw
rect 13117 44823 13391 44825
tri 13117 44815 13125 44823 ne
rect 13125 44817 13391 44823
tri 13391 44817 13399 44825 sw
rect 13125 44815 13399 44817
tri 13125 44807 13133 44815 ne
rect 13133 44809 13399 44815
tri 13399 44809 13407 44817 sw
rect 13133 44807 13407 44809
tri 13133 44799 13141 44807 ne
rect 13141 44801 13407 44807
tri 13407 44801 13415 44809 sw
rect 13141 44799 13415 44801
tri 13141 44791 13149 44799 ne
rect 13149 44793 13415 44799
tri 13415 44793 13423 44801 sw
rect 13149 44791 13423 44793
tri 13149 44783 13157 44791 ne
rect 13157 44787 13423 44791
tri 13423 44787 13429 44793 sw
rect 13157 44783 13429 44787
tri 13157 44775 13165 44783 ne
rect 13165 44779 13429 44783
tri 13429 44779 13437 44787 sw
rect 13165 44775 13437 44779
tri 13165 44767 13173 44775 ne
rect 13173 44771 13437 44775
tri 13437 44771 13445 44779 sw
rect 13173 44767 13445 44771
tri 13173 44759 13181 44767 ne
rect 13181 44763 13445 44767
tri 13445 44763 13453 44771 sw
rect 13181 44759 13453 44763
tri 13181 44751 13189 44759 ne
rect 13189 44755 13453 44759
tri 13453 44755 13461 44763 sw
rect 13189 44751 13461 44755
tri 13189 44743 13197 44751 ne
rect 13197 44747 13461 44751
tri 13461 44747 13469 44755 sw
rect 13197 44743 13469 44747
tri 13197 44735 13205 44743 ne
rect 13205 44739 13469 44743
tri 13469 44739 13477 44747 sw
rect 13205 44735 13477 44739
tri 13205 44727 13213 44735 ne
rect 13213 44731 13477 44735
tri 13477 44731 13485 44739 sw
rect 13213 44727 13485 44731
tri 13213 44719 13221 44727 ne
rect 13221 44723 13485 44727
tri 13485 44723 13493 44731 sw
rect 13221 44719 13493 44723
tri 13221 44711 13229 44719 ne
rect 13229 44715 13493 44719
tri 13493 44715 13501 44723 sw
rect 13229 44711 13501 44715
tri 13229 44703 13237 44711 ne
rect 13237 44707 13501 44711
tri 13501 44707 13509 44715 sw
rect 13237 44703 13509 44707
tri 13237 44695 13245 44703 ne
rect 13245 44699 13509 44703
tri 13509 44699 13517 44707 sw
rect 13245 44695 13517 44699
tri 13245 44687 13253 44695 ne
rect 13253 44691 13517 44695
tri 13517 44691 13525 44699 sw
rect 13253 44687 13525 44691
tri 13253 44679 13261 44687 ne
rect 13261 44683 13525 44687
tri 13525 44683 13533 44691 sw
rect 13261 44679 13533 44683
tri 13261 44671 13269 44679 ne
rect 13269 44675 13533 44679
tri 13533 44675 13541 44683 sw
rect 13269 44671 13541 44675
tri 13269 44663 13277 44671 ne
rect 13277 44667 13541 44671
tri 13541 44667 13549 44675 sw
rect 13277 44663 13549 44667
tri 13277 44655 13285 44663 ne
rect 13285 44659 13549 44663
tri 13549 44659 13557 44667 sw
rect 13285 44655 13557 44659
tri 13285 44651 13289 44655 ne
rect 13289 44651 13557 44655
tri 13557 44651 13565 44659 sw
tri 13289 44647 13293 44651 ne
rect 13293 44647 13565 44651
tri 13565 44647 13569 44651 sw
tri 13293 44639 13301 44647 ne
rect 13301 44639 13569 44647
tri 13569 44639 13577 44647 sw
tri 13301 44631 13309 44639 ne
rect 13309 44631 13577 44639
tri 13577 44631 13585 44639 sw
tri 13309 44623 13317 44631 ne
rect 13317 44623 13585 44631
tri 13585 44623 13593 44631 sw
tri 13317 44615 13325 44623 ne
rect 13325 44615 13593 44623
tri 13593 44615 13601 44623 sw
tri 13325 44607 13333 44615 ne
rect 13333 44607 13601 44615
tri 13601 44607 13609 44615 sw
tri 13333 44599 13341 44607 ne
rect 13341 44599 13609 44607
tri 13609 44599 13617 44607 sw
tri 13341 44591 13349 44599 ne
rect 13349 44591 13617 44599
tri 13617 44591 13625 44599 sw
tri 13349 44583 13357 44591 ne
rect 13357 44583 13625 44591
tri 13625 44583 13633 44591 sw
tri 13357 44575 13365 44583 ne
rect 13365 44575 13633 44583
tri 13633 44575 13641 44583 sw
tri 13365 44567 13373 44575 ne
rect 13373 44567 13641 44575
tri 13641 44567 13649 44575 sw
tri 13373 44559 13381 44567 ne
rect 13381 44559 13649 44567
tri 13649 44559 13657 44567 sw
tri 13381 44551 13389 44559 ne
rect 13389 44551 13657 44559
tri 13657 44551 13665 44559 sw
tri 13389 44543 13397 44551 ne
rect 13397 44543 13665 44551
tri 13665 44543 13673 44551 sw
tri 13397 44535 13405 44543 ne
rect 13405 44535 13673 44543
tri 13673 44535 13681 44543 sw
tri 13405 44527 13413 44535 ne
rect 13413 44527 13681 44535
tri 13681 44527 13689 44535 sw
tri 13413 44519 13421 44527 ne
rect 13421 44519 13689 44527
tri 13689 44519 13697 44527 sw
tri 13421 44511 13429 44519 ne
rect 13429 44511 13697 44519
tri 13697 44511 13705 44519 sw
tri 13429 44507 13433 44511 ne
rect 13433 44507 13705 44511
tri 13433 44499 13441 44507 ne
rect 13441 44503 13705 44507
tri 13705 44503 13713 44511 sw
rect 13441 44499 13713 44503
tri 13441 44491 13449 44499 ne
rect 13449 44495 13713 44499
tri 13713 44495 13721 44503 sw
rect 13449 44491 13721 44495
tri 13449 44483 13457 44491 ne
rect 13457 44487 13721 44491
tri 13721 44487 13729 44495 sw
rect 13457 44483 13729 44487
tri 13457 44475 13465 44483 ne
rect 13465 44479 13729 44483
tri 13729 44479 13737 44487 sw
rect 13465 44475 13737 44479
tri 13465 44467 13473 44475 ne
rect 13473 44471 13737 44475
tri 13737 44471 13745 44479 sw
rect 13473 44467 13745 44471
tri 13473 44459 13481 44467 ne
rect 13481 44463 13745 44467
tri 13745 44463 13753 44471 sw
rect 13481 44459 13753 44463
tri 13481 44451 13489 44459 ne
rect 13489 44455 13753 44459
tri 13753 44455 13761 44463 sw
rect 13489 44451 13761 44455
tri 13489 44443 13497 44451 ne
rect 13497 44447 13761 44451
tri 13761 44447 13769 44455 sw
rect 13497 44443 13769 44447
tri 13497 44435 13505 44443 ne
rect 13505 44439 13769 44443
tri 13769 44439 13777 44447 sw
rect 13505 44435 13777 44439
tri 13505 44427 13513 44435 ne
rect 13513 44431 13777 44435
tri 13777 44431 13785 44439 sw
rect 13513 44427 13785 44431
tri 13513 44419 13521 44427 ne
rect 13521 44423 13785 44427
tri 13785 44423 13793 44431 sw
rect 13521 44419 13793 44423
tri 13521 44411 13529 44419 ne
rect 13529 44415 13793 44419
tri 13793 44415 13801 44423 sw
rect 13529 44411 13801 44415
tri 13529 44403 13537 44411 ne
rect 13537 44407 13801 44411
tri 13801 44407 13809 44415 sw
rect 13537 44403 13809 44407
tri 13537 44395 13545 44403 ne
rect 13545 44399 13809 44403
tri 13809 44399 13817 44407 sw
rect 13545 44395 13817 44399
tri 13545 44387 13553 44395 ne
rect 13553 44391 13817 44395
tri 13817 44391 13825 44399 sw
rect 13553 44387 13825 44391
tri 13553 44379 13561 44387 ne
rect 13561 44383 13825 44387
tri 13825 44383 13833 44391 sw
rect 13561 44379 13833 44383
tri 13561 44375 13565 44379 ne
rect 13565 44375 13833 44379
tri 13833 44375 13841 44383 sw
tri 13565 44371 13569 44375 ne
rect 13569 44371 13841 44375
tri 13841 44371 13845 44375 sw
tri 13569 44363 13577 44371 ne
rect 13577 44363 13845 44371
tri 13845 44363 13853 44371 sw
tri 13577 44355 13585 44363 ne
rect 13585 44355 13853 44363
tri 13853 44355 13861 44363 sw
tri 13585 44347 13593 44355 ne
rect 13593 44347 13861 44355
tri 13861 44347 13869 44355 sw
tri 13593 44339 13601 44347 ne
rect 13601 44339 13869 44347
tri 13869 44339 13877 44347 sw
tri 13601 44331 13609 44339 ne
rect 13609 44331 13877 44339
tri 13877 44331 13885 44339 sw
tri 13609 44323 13617 44331 ne
rect 13617 44323 13885 44331
tri 13885 44323 13893 44331 sw
tri 13617 44315 13625 44323 ne
rect 13625 44315 13893 44323
tri 13893 44315 13901 44323 sw
tri 13625 44307 13633 44315 ne
rect 13633 44307 13901 44315
tri 13901 44307 13909 44315 sw
tri 13633 44299 13641 44307 ne
rect 13641 44299 13909 44307
tri 13909 44299 13917 44307 sw
tri 13641 44291 13649 44299 ne
rect 13649 44291 13917 44299
tri 13917 44291 13925 44299 sw
tri 13649 44283 13657 44291 ne
rect 13657 44283 13925 44291
tri 13925 44283 13933 44291 sw
tri 13657 44275 13665 44283 ne
rect 13665 44275 13933 44283
tri 13933 44275 13941 44283 sw
tri 13665 44267 13673 44275 ne
rect 13673 44267 13941 44275
tri 13941 44267 13949 44275 sw
tri 13673 44259 13681 44267 ne
rect 13681 44259 13949 44267
tri 13949 44259 13957 44267 sw
tri 13681 44251 13689 44259 ne
rect 13689 44251 13957 44259
tri 13957 44251 13965 44259 sw
tri 13689 44246 13694 44251 ne
rect 13694 44250 13965 44251
tri 13965 44250 13966 44251 sw
rect 13694 44246 13966 44250
tri 13694 44238 13702 44246 ne
rect 13702 44242 13966 44246
tri 13966 44242 13974 44250 sw
rect 13702 44238 13974 44242
tri 13702 44230 13710 44238 ne
rect 13710 44234 13974 44238
tri 13974 44234 13982 44242 sw
rect 13710 44230 13982 44234
tri 13710 44222 13718 44230 ne
rect 13718 44226 13982 44230
tri 13982 44226 13990 44234 sw
rect 13718 44222 13990 44226
tri 13718 44214 13726 44222 ne
rect 13726 44218 13990 44222
tri 13990 44218 13998 44226 sw
rect 13726 44214 13998 44218
tri 13726 44206 13734 44214 ne
rect 13734 44210 13998 44214
tri 13998 44210 14006 44218 sw
rect 13734 44206 14006 44210
tri 13734 44198 13742 44206 ne
rect 13742 44202 14006 44206
tri 14006 44202 14014 44210 sw
rect 13742 44198 14014 44202
tri 13742 44190 13750 44198 ne
rect 13750 44194 14014 44198
tri 14014 44194 14022 44202 sw
rect 13750 44190 14022 44194
tri 13750 44182 13758 44190 ne
rect 13758 44186 14022 44190
tri 14022 44186 14030 44194 sw
rect 13758 44182 14030 44186
tri 13758 44174 13766 44182 ne
rect 13766 44178 14030 44182
tri 14030 44178 14038 44186 sw
rect 13766 44174 14038 44178
tri 13766 44166 13774 44174 ne
rect 13774 44170 14038 44174
tri 14038 44170 14046 44178 sw
rect 13774 44166 14046 44170
tri 13774 44158 13782 44166 ne
rect 13782 44162 14046 44166
tri 14046 44162 14054 44170 sw
rect 13782 44158 14054 44162
tri 13782 44150 13790 44158 ne
rect 13790 44154 14054 44158
tri 14054 44154 14062 44162 sw
rect 13790 44150 14062 44154
tri 13790 44142 13798 44150 ne
rect 13798 44146 14062 44150
tri 14062 44146 14070 44154 sw
rect 13798 44142 14070 44146
tri 13798 44134 13806 44142 ne
rect 13806 44138 14070 44142
tri 14070 44138 14078 44146 sw
rect 13806 44134 14078 44138
tri 13806 44130 13810 44134 ne
rect 13810 44130 14078 44134
tri 14078 44130 14086 44138 sw
tri 13810 44126 13814 44130 ne
rect 13814 44126 14086 44130
tri 14086 44126 14090 44130 sw
tri 13814 44118 13822 44126 ne
rect 13822 44118 14090 44126
tri 14090 44118 14098 44126 sw
tri 13822 44110 13830 44118 ne
rect 13830 44110 14098 44118
tri 14098 44110 14106 44118 sw
tri 13830 44102 13838 44110 ne
rect 13838 44102 14106 44110
tri 14106 44102 14114 44110 sw
tri 13838 44094 13846 44102 ne
rect 13846 44094 14114 44102
tri 14114 44094 14122 44102 sw
tri 13846 44086 13854 44094 ne
rect 13854 44086 14122 44094
tri 14122 44086 14130 44094 sw
tri 13854 44078 13862 44086 ne
rect 13862 44078 14130 44086
tri 14130 44078 14138 44086 sw
tri 13862 44070 13870 44078 ne
rect 13870 44070 14138 44078
tri 14138 44070 14146 44078 sw
tri 13870 44062 13878 44070 ne
rect 13878 44062 14146 44070
tri 14146 44062 14154 44070 sw
tri 13878 44054 13886 44062 ne
rect 13886 44054 14154 44062
tri 14154 44054 14162 44062 sw
tri 13886 44046 13894 44054 ne
rect 13894 44046 14162 44054
tri 14162 44046 14170 44054 sw
tri 13894 44038 13902 44046 ne
rect 13902 44038 14170 44046
tri 14170 44038 14178 44046 sw
tri 13902 44030 13910 44038 ne
rect 13910 44030 14178 44038
tri 14178 44030 14186 44038 sw
tri 13910 44022 13918 44030 ne
rect 13918 44022 14186 44030
tri 14186 44022 14194 44030 sw
tri 13918 44014 13926 44022 ne
rect 13926 44014 14194 44022
tri 14194 44014 14202 44022 sw
tri 13926 44006 13934 44014 ne
rect 13934 44006 14202 44014
tri 14202 44006 14210 44014 sw
tri 13934 43998 13942 44006 ne
rect 13942 43998 14210 44006
tri 14210 43998 14218 44006 sw
tri 13942 43990 13950 43998 ne
rect 13950 43990 14218 43998
tri 14218 43990 14226 43998 sw
tri 13950 43986 13954 43990 ne
rect 13954 43986 14226 43990
tri 13954 43978 13962 43986 ne
rect 13962 43982 14226 43986
tri 14226 43982 14234 43990 sw
rect 13962 43978 14234 43982
tri 13962 43970 13970 43978 ne
rect 13970 43974 14234 43978
tri 14234 43974 14242 43982 sw
rect 13970 43970 14242 43974
tri 13970 43962 13978 43970 ne
rect 13978 43966 14242 43970
tri 14242 43966 14250 43974 sw
rect 13978 43962 14250 43966
tri 13978 43954 13986 43962 ne
rect 13986 43958 14250 43962
tri 14250 43958 14258 43966 sw
rect 13986 43954 14258 43958
tri 13986 43946 13994 43954 ne
rect 13994 43950 14258 43954
tri 14258 43950 14266 43958 sw
rect 13994 43946 14266 43950
tri 13994 43938 14002 43946 ne
rect 14002 43942 14266 43946
tri 14266 43942 14274 43950 sw
rect 14002 43938 14274 43942
tri 14002 43930 14010 43938 ne
rect 14010 43934 14274 43938
tri 14274 43934 14282 43942 sw
rect 14010 43930 14282 43934
tri 14010 43922 14018 43930 ne
rect 14018 43926 14282 43930
tri 14282 43926 14290 43934 sw
rect 14018 43922 14290 43926
tri 14018 43914 14026 43922 ne
rect 14026 43918 14290 43922
tri 14290 43918 14298 43926 sw
rect 14026 43914 14298 43918
tri 14026 43906 14034 43914 ne
rect 14034 43910 14298 43914
tri 14298 43910 14306 43918 sw
rect 14034 43906 14306 43910
tri 14034 43898 14042 43906 ne
rect 14042 43902 14306 43906
tri 14306 43902 14314 43910 sw
rect 14042 43898 14314 43902
tri 14042 43890 14050 43898 ne
rect 14050 43894 14314 43898
tri 14314 43894 14322 43902 sw
rect 14050 43890 14322 43894
tri 14050 43882 14058 43890 ne
rect 14058 43886 14322 43890
tri 14322 43886 14330 43894 sw
rect 14058 43882 14330 43886
tri 14058 43874 14066 43882 ne
rect 14066 43878 14330 43882
tri 14330 43878 14338 43886 sw
rect 14066 43874 14338 43878
tri 14066 43866 14074 43874 ne
rect 14074 43870 14338 43874
tri 14338 43870 14346 43878 sw
rect 14074 43866 14346 43870
tri 14074 43858 14082 43866 ne
rect 14082 43862 14346 43866
tri 14346 43862 14354 43870 sw
rect 14082 43858 14354 43862
tri 14082 43854 14086 43858 ne
rect 14086 43854 14354 43858
tri 14354 43854 14362 43862 sw
tri 14086 43850 14090 43854 ne
rect 14090 43850 14362 43854
tri 14362 43850 14366 43854 sw
tri 14090 43842 14098 43850 ne
rect 14098 43842 14366 43850
tri 14366 43842 14374 43850 sw
tri 14098 43834 14106 43842 ne
rect 14106 43834 14374 43842
tri 14374 43834 14382 43842 sw
tri 14106 43826 14114 43834 ne
rect 14114 43826 14382 43834
tri 14382 43826 14390 43834 sw
tri 14114 43818 14122 43826 ne
rect 14122 43818 14390 43826
tri 14390 43818 14398 43826 sw
tri 14122 43810 14130 43818 ne
rect 14130 43810 14398 43818
tri 14398 43810 14406 43818 sw
tri 14130 43802 14138 43810 ne
rect 14138 43802 14406 43810
tri 14406 43802 14414 43810 sw
tri 14138 43794 14146 43802 ne
rect 14146 43794 14414 43802
tri 14414 43794 14422 43802 sw
tri 14146 43786 14154 43794 ne
rect 14154 43786 14422 43794
tri 14422 43786 14430 43794 sw
tri 14154 43778 14162 43786 ne
rect 14162 43778 14430 43786
tri 14430 43778 14438 43786 sw
tri 14162 43770 14170 43778 ne
rect 14170 43770 14438 43778
tri 14438 43770 14446 43778 sw
tri 14170 43762 14178 43770 ne
rect 14178 43762 14446 43770
tri 14446 43762 14454 43770 sw
tri 14178 43754 14186 43762 ne
rect 14186 43754 14454 43762
tri 14454 43754 14462 43762 sw
tri 14186 43746 14194 43754 ne
rect 14194 43746 14462 43754
tri 14462 43746 14470 43754 sw
tri 14194 43738 14202 43746 ne
rect 14202 43738 14470 43746
tri 14470 43738 14478 43746 sw
tri 14202 43730 14210 43738 ne
rect 14210 43730 14478 43738
tri 14478 43730 14486 43738 sw
tri 14210 43722 14218 43730 ne
rect 14218 43722 14486 43730
tri 14486 43722 14494 43730 sw
tri 14218 43714 14226 43722 ne
rect 14226 43720 14494 43722
tri 14494 43720 14496 43722 sw
rect 14226 43714 14496 43720
tri 14226 43710 14230 43714 ne
rect 14230 43712 14496 43714
tri 14496 43712 14504 43720 sw
rect 14230 43710 14504 43712
tri 14230 43702 14238 43710 ne
rect 14238 43704 14504 43710
tri 14504 43704 14512 43712 sw
rect 14238 43702 14512 43704
tri 14238 43694 14246 43702 ne
rect 14246 43696 14512 43702
tri 14512 43696 14520 43704 sw
rect 14246 43694 14520 43696
tri 14246 43686 14254 43694 ne
rect 14254 43688 14520 43694
tri 14520 43688 14528 43696 sw
rect 14254 43686 14528 43688
tri 14254 43678 14262 43686 ne
rect 14262 43680 14528 43686
tri 14528 43680 14536 43688 sw
rect 14262 43678 14536 43680
tri 14262 43670 14270 43678 ne
rect 14270 43672 14536 43678
tri 14536 43672 14544 43680 sw
rect 14270 43670 14544 43672
tri 14270 43662 14278 43670 ne
rect 14278 43664 14544 43670
tri 14544 43664 14552 43672 sw
rect 14278 43662 14552 43664
tri 14278 43654 14286 43662 ne
rect 14286 43656 14552 43662
tri 14552 43656 14560 43664 sw
rect 14286 43654 14560 43656
tri 14286 43646 14294 43654 ne
rect 14294 43648 14560 43654
tri 14560 43648 14568 43656 sw
rect 14294 43646 14568 43648
tri 14294 43638 14302 43646 ne
rect 14302 43640 14568 43646
tri 14568 43640 14576 43648 sw
rect 14302 43638 14576 43640
tri 14302 43630 14310 43638 ne
rect 14310 43632 14576 43638
tri 14576 43632 14584 43640 sw
rect 14310 43630 14584 43632
tri 14310 43622 14318 43630 ne
rect 14318 43624 14584 43630
tri 14584 43624 14592 43632 sw
rect 14318 43622 14592 43624
tri 14318 43614 14326 43622 ne
rect 14326 43616 14592 43622
tri 14592 43616 14600 43624 sw
rect 14326 43614 14600 43616
tri 14326 43606 14334 43614 ne
rect 14334 43608 14600 43614
tri 14600 43608 14608 43616 sw
rect 14334 43606 14608 43608
tri 14334 43598 14342 43606 ne
rect 14342 43600 14608 43606
tri 14608 43600 14616 43608 sw
rect 14342 43598 14616 43600
tri 14342 43590 14350 43598 ne
rect 14350 43592 14616 43598
tri 14616 43592 14624 43600 sw
rect 14350 43590 14624 43592
tri 14350 43582 14358 43590 ne
rect 14358 43584 14624 43590
tri 14624 43584 14632 43592 sw
rect 14358 43582 14632 43584
tri 14632 43582 14634 43584 sw
tri 14358 43578 14362 43582 ne
rect 14362 43578 14634 43582
tri 14362 43574 14366 43578 ne
rect 14366 43574 14634 43578
tri 14634 43574 14642 43582 sw
tri 14366 43566 14374 43574 ne
rect 14374 43566 14642 43574
tri 14642 43566 14650 43574 sw
tri 14374 43558 14382 43566 ne
rect 14382 43558 14650 43566
tri 14650 43558 14658 43566 sw
tri 14382 43550 14390 43558 ne
rect 14390 43550 14658 43558
tri 14658 43550 14666 43558 sw
tri 14390 43542 14398 43550 ne
rect 14398 43542 14666 43550
tri 14666 43542 14674 43550 sw
tri 14398 43534 14406 43542 ne
rect 14406 43534 14674 43542
tri 14674 43534 14682 43542 sw
tri 14406 43526 14414 43534 ne
rect 14414 43526 14682 43534
tri 14682 43526 14690 43534 sw
tri 14414 43518 14422 43526 ne
rect 14422 43518 14690 43526
tri 14690 43518 14698 43526 sw
tri 14422 43510 14430 43518 ne
rect 14430 43510 14698 43518
tri 14698 43510 14706 43518 sw
tri 14430 43502 14438 43510 ne
rect 14438 43502 14706 43510
tri 14706 43502 14714 43510 sw
tri 14438 43494 14446 43502 ne
rect 14446 43494 14714 43502
tri 14714 43494 14722 43502 sw
tri 14446 43486 14454 43494 ne
rect 14454 43486 14722 43494
tri 14722 43486 14730 43494 sw
tri 14454 43478 14462 43486 ne
rect 14462 43478 14730 43486
tri 14730 43478 14738 43486 sw
tri 14462 43470 14470 43478 ne
rect 14470 43470 14738 43478
tri 14738 43470 14746 43478 sw
tri 14470 43462 14478 43470 ne
rect 14478 43462 14746 43470
tri 14746 43462 14754 43470 sw
tri 14478 43461 14479 43462 ne
rect 14479 43461 14754 43462
tri 14479 43453 14487 43461 ne
rect 14487 43457 14754 43461
tri 14754 43457 14759 43462 sw
rect 14487 43453 14759 43457
tri 14487 43445 14495 43453 ne
rect 14495 43449 14759 43453
tri 14759 43449 14767 43457 sw
rect 14495 43445 14767 43449
tri 14495 43437 14503 43445 ne
rect 14503 43441 14767 43445
tri 14767 43441 14775 43449 sw
rect 14503 43437 14775 43441
tri 14503 43429 14511 43437 ne
rect 14511 43433 14775 43437
tri 14775 43433 14783 43441 sw
rect 14511 43429 14783 43433
tri 14511 43421 14519 43429 ne
rect 14519 43425 14783 43429
tri 14783 43425 14791 43433 sw
rect 14519 43421 14791 43425
tri 14519 43413 14527 43421 ne
rect 14527 43417 14791 43421
tri 14791 43417 14799 43425 sw
rect 14527 43413 14799 43417
tri 14527 43405 14535 43413 ne
rect 14535 43409 14799 43413
tri 14799 43409 14807 43417 sw
rect 14535 43405 14807 43409
tri 14535 43397 14543 43405 ne
rect 14543 43401 14807 43405
tri 14807 43401 14815 43409 sw
rect 14543 43397 14815 43401
tri 14543 43389 14551 43397 ne
rect 14551 43393 14815 43397
tri 14815 43393 14823 43401 sw
rect 14551 43389 14823 43393
tri 14551 43381 14559 43389 ne
rect 14559 43385 14823 43389
tri 14823 43385 14831 43393 sw
rect 14559 43381 14831 43385
tri 14559 43373 14567 43381 ne
rect 14567 43377 14831 43381
tri 14831 43377 14839 43385 sw
rect 14567 43373 14839 43377
tri 14567 43365 14575 43373 ne
rect 14575 43369 14839 43373
tri 14839 43369 14847 43377 sw
rect 14575 43365 14847 43369
tri 14575 43357 14583 43365 ne
rect 14583 43361 14847 43365
tri 14847 43361 14855 43369 sw
rect 14583 43357 14855 43361
tri 14583 43353 14587 43357 ne
rect 14587 43353 14855 43357
tri 14855 43353 14863 43361 sw
tri 14587 43349 14591 43353 ne
rect 14591 43349 14863 43353
tri 14863 43349 14867 43353 sw
tri 14591 43341 14599 43349 ne
rect 14599 43341 14867 43349
tri 14867 43341 14875 43349 sw
tri 14599 43333 14607 43341 ne
rect 14607 43333 14875 43341
tri 14875 43333 14883 43341 sw
tri 14607 43325 14615 43333 ne
rect 14615 43325 14883 43333
tri 14883 43325 14891 43333 sw
tri 14615 43317 14623 43325 ne
rect 14623 43317 14891 43325
tri 14891 43317 14899 43325 sw
tri 14623 43309 14631 43317 ne
rect 14631 43309 14899 43317
tri 14899 43309 14907 43317 sw
tri 14631 43301 14639 43309 ne
rect 14639 43301 14907 43309
tri 14907 43301 14915 43309 sw
tri 14639 43293 14647 43301 ne
rect 14647 43293 14915 43301
tri 14915 43293 14923 43301 sw
tri 14647 43285 14655 43293 ne
rect 14655 43285 14923 43293
tri 14923 43285 14931 43293 sw
tri 14655 43277 14663 43285 ne
rect 14663 43277 14931 43285
tri 14931 43277 14939 43285 sw
tri 14663 43269 14671 43277 ne
rect 14671 43269 14939 43277
tri 14939 43269 14947 43277 sw
tri 14671 43261 14679 43269 ne
rect 14679 43261 14947 43269
tri 14947 43261 14955 43269 sw
tri 14679 43253 14687 43261 ne
rect 14687 43253 14955 43261
tri 14955 43253 14963 43261 sw
tri 14687 43245 14695 43253 ne
rect 14695 43245 14963 43253
tri 14963 43245 14971 43253 sw
tri 14695 43237 14703 43245 ne
rect 14703 43237 14971 43245
tri 14971 43237 14979 43245 sw
tri 14703 43229 14711 43237 ne
rect 14711 43229 14979 43237
tri 14979 43229 14987 43237 sw
tri 14711 43221 14719 43229 ne
rect 14719 43221 14987 43229
tri 14987 43221 14995 43229 sw
tri 14719 43213 14727 43221 ne
rect 14727 43213 14995 43221
tri 14995 43213 15003 43221 sw
tri 14727 43209 14731 43213 ne
rect 14731 43209 15003 43213
tri 14731 43201 14739 43209 ne
rect 14739 43205 15003 43209
tri 15003 43205 15011 43213 sw
rect 14739 43201 15011 43205
tri 14739 43193 14747 43201 ne
rect 14747 43197 15011 43201
tri 15011 43197 15019 43205 sw
rect 14747 43193 15019 43197
tri 14747 43185 14755 43193 ne
rect 14755 43189 15019 43193
tri 15019 43189 15027 43197 sw
rect 14755 43185 15027 43189
tri 14755 43177 14763 43185 ne
rect 14763 43181 15027 43185
tri 15027 43181 15035 43189 sw
rect 14763 43177 15035 43181
tri 14763 43169 14771 43177 ne
rect 14771 43173 15035 43177
tri 15035 43173 15043 43181 sw
rect 14771 43169 15043 43173
tri 14771 43161 14779 43169 ne
rect 14779 43165 15043 43169
tri 15043 43165 15051 43173 sw
rect 14779 43161 15051 43165
tri 14779 43153 14787 43161 ne
rect 14787 43157 15051 43161
tri 15051 43157 15059 43165 sw
rect 14787 43153 15059 43157
tri 14787 43145 14795 43153 ne
rect 14795 43149 15059 43153
tri 15059 43149 15067 43157 sw
rect 14795 43145 15067 43149
tri 14795 43137 14803 43145 ne
rect 14803 43141 15067 43145
tri 15067 43141 15075 43149 sw
rect 14803 43137 15075 43141
tri 14803 43129 14811 43137 ne
rect 14811 43133 15075 43137
tri 15075 43133 15083 43141 sw
rect 14811 43129 15083 43133
tri 14811 43121 14819 43129 ne
rect 14819 43125 15083 43129
tri 15083 43125 15091 43133 sw
rect 14819 43121 15091 43125
tri 14819 43113 14827 43121 ne
rect 14827 43117 15091 43121
tri 15091 43117 15099 43125 sw
rect 14827 43113 15099 43117
tri 14827 43105 14835 43113 ne
rect 14835 43109 15099 43113
tri 15099 43109 15107 43117 sw
rect 14835 43105 15107 43109
tri 14835 43097 14843 43105 ne
rect 14843 43101 15107 43105
tri 15107 43101 15115 43109 sw
rect 14843 43097 15115 43101
tri 14843 43089 14851 43097 ne
rect 14851 43093 15115 43097
tri 15115 43093 15123 43101 sw
rect 14851 43089 15123 43093
tri 14851 43081 14859 43089 ne
rect 14859 43085 15123 43089
tri 15123 43085 15131 43093 sw
rect 14859 43081 15131 43085
tri 14859 43077 14863 43081 ne
rect 14863 43077 15131 43081
tri 15131 43077 15139 43085 sw
tri 14863 43073 14867 43077 ne
rect 14867 43073 15139 43077
tri 15139 43073 15143 43077 sw
tri 14867 43065 14875 43073 ne
rect 14875 43065 15143 43073
tri 15143 43065 15151 43073 sw
tri 14875 43057 14883 43065 ne
rect 14883 43057 15151 43065
tri 15151 43057 15159 43065 sw
tri 14883 43049 14891 43057 ne
rect 14891 43049 15159 43057
tri 15159 43049 15167 43057 sw
tri 14891 43041 14899 43049 ne
rect 14899 43041 15167 43049
tri 15167 43041 15175 43049 sw
tri 14899 43033 14907 43041 ne
rect 14907 43033 15175 43041
tri 15175 43033 15183 43041 sw
tri 14907 43025 14915 43033 ne
rect 14915 43025 15183 43033
tri 15183 43025 15191 43033 sw
tri 14915 43017 14923 43025 ne
rect 14923 43017 15191 43025
tri 15191 43017 15199 43025 sw
tri 14923 43009 14931 43017 ne
rect 14931 43009 15199 43017
tri 15199 43009 15207 43017 sw
tri 14931 43001 14939 43009 ne
rect 14939 43001 15207 43009
tri 15207 43001 15215 43009 sw
tri 14939 42993 14947 43001 ne
rect 14947 42993 15215 43001
tri 15215 42993 15223 43001 sw
tri 14947 42985 14955 42993 ne
rect 14955 42985 15223 42993
tri 15223 42985 15231 42993 sw
tri 14955 42977 14963 42985 ne
rect 14963 42977 15231 42985
tri 15231 42977 15239 42985 sw
tri 14963 42969 14971 42977 ne
rect 14971 42969 15239 42977
tri 15239 42969 15247 42977 sw
tri 14971 42961 14979 42969 ne
rect 14979 42961 15247 42969
tri 15247 42961 15255 42969 sw
tri 14979 42953 14987 42961 ne
rect 14987 42953 15255 42961
tri 15255 42953 15263 42961 sw
tri 14987 42945 14995 42953 ne
rect 14995 42945 15263 42953
tri 15263 42945 15271 42953 sw
tri 14995 42937 15003 42945 ne
rect 15003 42937 15271 42945
tri 15271 42937 15279 42945 sw
tri 15003 42933 15007 42937 ne
rect 15007 42933 15279 42937
tri 15007 42925 15015 42933 ne
rect 15015 42929 15279 42933
tri 15279 42929 15287 42937 sw
rect 15015 42925 15287 42929
tri 15015 42917 15023 42925 ne
rect 15023 42921 15287 42925
tri 15287 42921 15295 42929 sw
rect 15023 42917 15295 42921
tri 15023 42909 15031 42917 ne
rect 15031 42913 15295 42917
tri 15295 42913 15303 42921 sw
rect 15031 42909 15303 42913
tri 15031 42901 15039 42909 ne
rect 15039 42905 15303 42909
tri 15303 42905 15311 42913 sw
rect 15039 42901 15311 42905
tri 15039 42893 15047 42901 ne
rect 15047 42897 15311 42901
tri 15311 42897 15319 42905 sw
rect 15047 42893 15319 42897
tri 15047 42885 15055 42893 ne
rect 15055 42889 15319 42893
tri 15319 42889 15327 42897 sw
rect 15055 42885 15327 42889
tri 15055 42877 15063 42885 ne
rect 15063 42881 15327 42885
tri 15327 42881 15335 42889 sw
rect 15063 42877 15335 42881
tri 15063 42869 15071 42877 ne
rect 15071 42873 15335 42877
tri 15335 42873 15343 42881 sw
rect 15071 42869 15343 42873
tri 15071 42861 15079 42869 ne
rect 15079 42865 15343 42869
tri 15343 42865 15351 42873 sw
rect 15079 42861 15351 42865
tri 15079 42853 15087 42861 ne
rect 15087 42857 15351 42861
tri 15351 42857 15359 42865 sw
rect 15087 42853 15359 42857
tri 15087 42845 15095 42853 ne
rect 15095 42849 15359 42853
tri 15359 42849 15367 42857 sw
rect 15095 42845 15367 42849
tri 15095 42837 15103 42845 ne
rect 15103 42841 15367 42845
tri 15367 42841 15375 42849 sw
rect 15103 42837 15375 42841
tri 15103 42829 15111 42837 ne
rect 15111 42833 15375 42837
tri 15375 42833 15383 42841 sw
rect 15111 42829 15383 42833
tri 15111 42821 15119 42829 ne
rect 15119 42825 15383 42829
tri 15383 42825 15391 42833 sw
rect 15119 42821 15391 42825
tri 15119 42813 15127 42821 ne
rect 15127 42817 15391 42821
tri 15391 42817 15399 42825 sw
rect 15127 42813 15399 42817
tri 15127 42805 15135 42813 ne
rect 15135 42809 15399 42813
tri 15399 42809 15407 42817 sw
rect 15135 42805 15407 42809
tri 15135 42801 15139 42805 ne
rect 15139 42801 15407 42805
tri 15407 42801 15415 42809 sw
tri 15139 42797 15143 42801 ne
rect 15143 42797 15415 42801
tri 15415 42797 15419 42801 sw
tri 15143 42789 15151 42797 ne
rect 15151 42789 15419 42797
tri 15419 42789 15427 42797 sw
tri 15151 42781 15159 42789 ne
rect 15159 42781 15427 42789
tri 15427 42781 15435 42789 sw
tri 15159 42773 15167 42781 ne
rect 15167 42773 15435 42781
tri 15435 42773 15443 42781 sw
tri 15167 42765 15175 42773 ne
rect 15175 42765 15443 42773
tri 15443 42765 15451 42773 sw
tri 15175 42757 15183 42765 ne
rect 15183 42757 15451 42765
tri 15451 42757 15459 42765 sw
tri 15183 42749 15191 42757 ne
rect 15191 42749 15459 42757
tri 15459 42749 15467 42757 sw
tri 15191 42741 15199 42749 ne
rect 15199 42741 15467 42749
tri 15467 42741 15475 42749 sw
tri 15199 42733 15207 42741 ne
rect 15207 42733 15475 42741
tri 15475 42733 15483 42741 sw
tri 15207 42725 15215 42733 ne
rect 15215 42725 15483 42733
tri 15483 42725 15491 42733 sw
tri 15215 42717 15223 42725 ne
rect 15223 42717 15491 42725
tri 15491 42717 15499 42725 sw
tri 15223 42709 15231 42717 ne
rect 15231 42709 15499 42717
tri 15499 42709 15507 42717 sw
tri 15231 42701 15239 42709 ne
rect 15239 42701 15507 42709
tri 15507 42701 15515 42709 sw
tri 15239 42693 15247 42701 ne
rect 15247 42693 15515 42701
tri 15515 42693 15523 42701 sw
tri 15247 42685 15255 42693 ne
rect 15255 42685 15523 42693
tri 15523 42685 15531 42693 sw
tri 15255 42677 15263 42685 ne
rect 15263 42677 15531 42685
tri 15531 42677 15539 42685 sw
tri 15263 42669 15271 42677 ne
rect 15271 42669 15539 42677
tri 15539 42669 15547 42677 sw
tri 15271 42663 15277 42669 ne
rect 15277 42667 15547 42669
tri 15547 42667 15549 42669 sw
rect 15277 42663 15549 42667
tri 15277 42655 15285 42663 ne
rect 15285 42659 15549 42663
tri 15549 42659 15557 42667 sw
rect 15285 42655 15557 42659
tri 15285 42647 15293 42655 ne
rect 15293 42651 15557 42655
tri 15557 42651 15565 42659 sw
rect 15293 42647 15565 42651
tri 15293 42639 15301 42647 ne
rect 15301 42643 15565 42647
tri 15565 42643 15573 42651 sw
rect 15301 42639 15573 42643
tri 15301 42631 15309 42639 ne
rect 15309 42635 15573 42639
tri 15573 42635 15581 42643 sw
rect 15309 42631 15581 42635
tri 15309 42623 15317 42631 ne
rect 15317 42627 15581 42631
tri 15581 42627 15589 42635 sw
rect 15317 42623 15589 42627
tri 15317 42615 15325 42623 ne
rect 15325 42619 15589 42623
tri 15589 42619 15597 42627 sw
rect 15325 42615 15597 42619
tri 15325 42607 15333 42615 ne
rect 15333 42611 15597 42615
tri 15597 42611 15605 42619 sw
rect 15333 42607 15605 42611
tri 15333 42599 15341 42607 ne
rect 15341 42603 15605 42607
tri 15605 42603 15613 42611 sw
rect 15341 42599 15613 42603
tri 15341 42591 15349 42599 ne
rect 15349 42595 15613 42599
tri 15613 42595 15621 42603 sw
rect 15349 42591 15621 42595
tri 15349 42583 15357 42591 ne
rect 15357 42587 15621 42591
tri 15621 42587 15629 42595 sw
rect 15357 42583 15629 42587
tri 15357 42575 15365 42583 ne
rect 15365 42579 15629 42583
tri 15629 42579 15637 42587 sw
rect 15365 42575 15637 42579
tri 15365 42567 15373 42575 ne
rect 15373 42571 15637 42575
tri 15637 42571 15645 42579 sw
rect 15373 42567 15645 42571
tri 15373 42559 15381 42567 ne
rect 15381 42563 15645 42567
tri 15645 42563 15653 42571 sw
rect 15381 42559 15653 42563
tri 15381 42551 15389 42559 ne
rect 15389 42555 15653 42559
tri 15653 42555 15661 42563 sw
rect 15389 42551 15661 42555
tri 15389 42543 15397 42551 ne
rect 15397 42547 15661 42551
tri 15661 42547 15669 42555 sw
rect 15397 42543 15669 42547
tri 15397 42539 15401 42543 ne
rect 15401 42539 15669 42543
tri 15669 42539 15677 42547 sw
tri 15401 42535 15405 42539 ne
rect 15405 42535 15677 42539
tri 15677 42535 15681 42539 sw
tri 15405 42527 15413 42535 ne
rect 15413 42527 15681 42535
tri 15681 42527 15689 42535 sw
tri 15413 42519 15421 42527 ne
rect 15421 42519 15689 42527
tri 15689 42519 15697 42527 sw
tri 15421 42511 15429 42519 ne
rect 15429 42511 15697 42519
tri 15697 42511 15705 42519 sw
tri 15429 42503 15437 42511 ne
rect 15437 42503 15705 42511
tri 15705 42503 15713 42511 sw
tri 15437 42495 15445 42503 ne
rect 15445 42495 15713 42503
tri 15713 42495 15721 42503 sw
tri 15445 42487 15453 42495 ne
rect 15453 42487 15721 42495
tri 15721 42487 15729 42495 sw
tri 15453 42479 15461 42487 ne
rect 15461 42479 15729 42487
tri 15729 42479 15737 42487 sw
tri 15461 42471 15469 42479 ne
rect 15469 42471 15737 42479
tri 15737 42471 15745 42479 sw
tri 15469 42463 15477 42471 ne
rect 15477 42463 15745 42471
tri 15745 42463 15753 42471 sw
tri 15477 42455 15485 42463 ne
rect 15485 42455 15753 42463
tri 15753 42455 15761 42463 sw
tri 15485 42447 15493 42455 ne
rect 15493 42447 15761 42455
tri 15761 42447 15769 42455 sw
tri 15493 42439 15501 42447 ne
rect 15501 42439 15769 42447
tri 15769 42439 15777 42447 sw
tri 15501 42431 15509 42439 ne
rect 15509 42431 15777 42439
tri 15777 42431 15785 42439 sw
tri 15509 42423 15517 42431 ne
rect 15517 42423 15785 42431
tri 15785 42423 15793 42431 sw
tri 15517 42416 15524 42423 ne
rect 15524 42416 15793 42423
tri 15524 42408 15532 42416 ne
rect 15532 42415 15793 42416
tri 15793 42415 15801 42423 sw
rect 15532 42412 15801 42415
tri 15801 42412 15804 42415 sw
rect 15532 42408 15804 42412
tri 15532 42400 15540 42408 ne
rect 15540 42404 15804 42408
tri 15804 42404 15812 42412 sw
rect 15540 42400 15812 42404
tri 15540 42392 15548 42400 ne
rect 15548 42396 15812 42400
tri 15812 42396 15820 42404 sw
rect 15548 42392 15820 42396
tri 15548 42384 15556 42392 ne
rect 15556 42388 15820 42392
tri 15820 42388 15828 42396 sw
rect 15556 42384 15828 42388
tri 15556 42376 15564 42384 ne
rect 15564 42380 15828 42384
tri 15828 42380 15836 42388 sw
rect 15564 42376 15836 42380
tri 15564 42368 15572 42376 ne
rect 15572 42372 15836 42376
tri 15836 42372 15844 42380 sw
rect 15572 42368 15844 42372
tri 15572 42360 15580 42368 ne
rect 15580 42364 15844 42368
tri 15844 42364 15852 42372 sw
rect 15580 42360 15852 42364
tri 15580 42352 15588 42360 ne
rect 15588 42356 15852 42360
tri 15852 42356 15860 42364 sw
rect 15588 42352 15860 42356
tri 15588 42344 15596 42352 ne
rect 15596 42348 15860 42352
tri 15860 42348 15868 42356 sw
rect 15596 42344 15868 42348
tri 15596 42336 15604 42344 ne
rect 15604 42340 15868 42344
tri 15868 42340 15876 42348 sw
rect 15604 42336 15876 42340
tri 15604 42328 15612 42336 ne
rect 15612 42332 15876 42336
tri 15876 42332 15884 42340 sw
rect 15612 42328 15884 42332
tri 15612 42320 15620 42328 ne
rect 15620 42324 15884 42328
tri 15884 42324 15892 42332 sw
rect 15620 42320 15892 42324
tri 15620 42312 15628 42320 ne
rect 15628 42316 15892 42320
tri 15892 42316 15900 42324 sw
rect 15628 42312 15900 42316
tri 15628 42304 15636 42312 ne
rect 15636 42308 15900 42312
tri 15900 42308 15908 42316 sw
rect 15636 42304 15908 42308
tri 15636 42300 15640 42304 ne
rect 15640 42300 15908 42304
tri 15908 42300 15916 42308 sw
tri 15640 42296 15644 42300 ne
rect 15644 42296 15916 42300
tri 15916 42296 15920 42300 sw
tri 15644 42288 15652 42296 ne
rect 15652 42288 15920 42296
tri 15920 42288 15928 42296 sw
tri 15652 42280 15660 42288 ne
rect 15660 42280 15928 42288
tri 15928 42280 15936 42288 sw
tri 15660 42272 15668 42280 ne
rect 15668 42272 15936 42280
tri 15936 42272 15944 42280 sw
tri 15668 42264 15676 42272 ne
rect 15676 42264 15944 42272
tri 15944 42264 15952 42272 sw
tri 15676 42256 15684 42264 ne
rect 15684 42256 15952 42264
tri 15952 42256 15960 42264 sw
tri 15684 42248 15692 42256 ne
rect 15692 42248 15960 42256
tri 15960 42248 15968 42256 sw
tri 15692 42240 15700 42248 ne
rect 15700 42240 15968 42248
tri 15968 42240 15976 42248 sw
tri 15700 42232 15708 42240 ne
rect 15708 42232 15976 42240
tri 15976 42232 15984 42240 sw
tri 15708 42224 15716 42232 ne
rect 15716 42224 15984 42232
tri 15984 42224 15992 42232 sw
tri 15716 42216 15724 42224 ne
rect 15724 42216 15992 42224
tri 15992 42216 16000 42224 sw
tri 15724 42208 15732 42216 ne
rect 15732 42208 16000 42216
tri 16000 42208 16008 42216 sw
tri 15732 42200 15740 42208 ne
rect 15740 42200 16008 42208
tri 16008 42200 16016 42208 sw
tri 15740 42192 15748 42200 ne
rect 15748 42192 16016 42200
tri 16016 42192 16024 42200 sw
tri 15748 42184 15756 42192 ne
rect 15756 42184 16024 42192
tri 16024 42184 16032 42192 sw
tri 15756 42176 15764 42184 ne
rect 15764 42176 16032 42184
tri 16032 42176 16040 42184 sw
tri 15764 42168 15772 42176 ne
rect 15772 42168 16040 42176
tri 16040 42168 16048 42176 sw
tri 15772 42160 15780 42168 ne
rect 15780 42160 16048 42168
tri 16048 42160 16056 42168 sw
tri 15780 42156 15784 42160 ne
rect 15784 42156 16056 42160
tri 15784 42148 15792 42156 ne
rect 15792 42152 16056 42156
tri 16056 42152 16064 42160 sw
rect 15792 42148 16064 42152
tri 15792 42140 15800 42148 ne
rect 15800 42144 16064 42148
tri 16064 42144 16072 42152 sw
rect 15800 42140 16072 42144
tri 15800 42132 15808 42140 ne
rect 15808 42136 16072 42140
tri 16072 42136 16080 42144 sw
rect 15808 42132 16080 42136
tri 15808 42124 15816 42132 ne
rect 15816 42128 16080 42132
tri 16080 42128 16088 42136 sw
rect 15816 42124 16088 42128
tri 15816 42116 15824 42124 ne
rect 15824 42120 16088 42124
tri 16088 42120 16096 42128 sw
rect 15824 42116 16096 42120
tri 15824 42108 15832 42116 ne
rect 15832 42112 16096 42116
tri 16096 42112 16104 42120 sw
rect 15832 42108 16104 42112
tri 15832 42100 15840 42108 ne
rect 15840 42104 16104 42108
tri 16104 42104 16112 42112 sw
rect 15840 42100 16112 42104
tri 15840 42092 15848 42100 ne
rect 15848 42096 16112 42100
tri 16112 42096 16120 42104 sw
rect 15848 42092 16120 42096
tri 15848 42084 15856 42092 ne
rect 15856 42088 16120 42092
tri 16120 42088 16128 42096 sw
rect 15856 42084 16128 42088
tri 15856 42076 15864 42084 ne
rect 15864 42080 16128 42084
tri 16128 42080 16136 42088 sw
rect 15864 42076 16136 42080
tri 15864 42068 15872 42076 ne
rect 15872 42072 16136 42076
tri 16136 42072 16144 42080 sw
rect 15872 42068 16144 42072
tri 15872 42060 15880 42068 ne
rect 15880 42064 16144 42068
tri 16144 42064 16152 42072 sw
rect 15880 42060 16152 42064
tri 15880 42052 15888 42060 ne
rect 15888 42056 16152 42060
tri 16152 42056 16160 42064 sw
rect 15888 42052 16160 42056
tri 15888 42044 15896 42052 ne
rect 15896 42048 16160 42052
tri 16160 42048 16168 42056 sw
rect 15896 42044 16168 42048
tri 15896 42036 15904 42044 ne
rect 15904 42040 16168 42044
tri 16168 42040 16176 42048 sw
rect 15904 42036 16176 42040
tri 15904 42028 15912 42036 ne
rect 15912 42032 16176 42036
tri 16176 42032 16184 42040 sw
rect 15912 42028 16184 42032
tri 15912 42024 15916 42028 ne
rect 15916 42024 16184 42028
tri 16184 42024 16192 42032 sw
tri 15916 42020 15920 42024 ne
rect 15920 42020 16192 42024
tri 16192 42020 16196 42024 sw
tri 15920 42012 15928 42020 ne
rect 15928 42012 16196 42020
tri 16196 42012 16204 42020 sw
tri 15928 42004 15936 42012 ne
rect 15936 42004 16204 42012
tri 16204 42004 16212 42012 sw
tri 15936 41996 15944 42004 ne
rect 15944 41996 16212 42004
tri 16212 41996 16220 42004 sw
tri 15944 41988 15952 41996 ne
rect 15952 41988 16220 41996
tri 16220 41988 16228 41996 sw
tri 15952 41980 15960 41988 ne
rect 15960 41980 16228 41988
tri 16228 41980 16236 41988 sw
tri 15960 41972 15968 41980 ne
rect 15968 41972 16236 41980
tri 16236 41972 16244 41980 sw
tri 15968 41964 15976 41972 ne
rect 15976 41964 16244 41972
tri 16244 41964 16252 41972 sw
tri 15976 41956 15984 41964 ne
rect 15984 41956 16252 41964
tri 16252 41956 16260 41964 sw
tri 15984 41948 15992 41956 ne
rect 15992 41948 16260 41956
tri 16260 41948 16268 41956 sw
tri 15992 41940 16000 41948 ne
rect 16000 41940 16268 41948
tri 16268 41940 16276 41948 sw
tri 16000 41932 16008 41940 ne
rect 16008 41932 16276 41940
tri 16276 41932 16284 41940 sw
tri 16008 41924 16016 41932 ne
rect 16016 41924 16284 41932
tri 16284 41924 16292 41932 sw
tri 16016 41916 16024 41924 ne
rect 16024 41916 16292 41924
tri 16292 41916 16300 41924 sw
tri 16024 41908 16032 41916 ne
rect 16032 41908 16300 41916
tri 16300 41908 16308 41916 sw
tri 16032 41900 16040 41908 ne
rect 16040 41900 16308 41908
tri 16308 41900 16316 41908 sw
tri 16040 41892 16048 41900 ne
rect 16048 41892 16316 41900
tri 16316 41892 16324 41900 sw
tri 16048 41888 16052 41892 ne
rect 16052 41888 16324 41892
tri 16052 41880 16060 41888 ne
rect 16060 41884 16324 41888
tri 16324 41884 16332 41892 sw
rect 16060 41880 16332 41884
tri 16060 41872 16068 41880 ne
rect 16068 41876 16332 41880
tri 16332 41876 16340 41884 sw
rect 16068 41872 16340 41876
tri 16068 41864 16076 41872 ne
rect 16076 41868 16340 41872
tri 16340 41868 16348 41876 sw
rect 16076 41864 16348 41868
tri 16076 41856 16084 41864 ne
rect 16084 41860 16348 41864
tri 16348 41860 16356 41868 sw
rect 16084 41856 16356 41860
tri 16084 41848 16092 41856 ne
rect 16092 41852 16356 41856
tri 16356 41852 16364 41860 sw
rect 16092 41848 16364 41852
tri 16092 41840 16100 41848 ne
rect 16100 41844 16364 41848
tri 16364 41844 16372 41852 sw
rect 16100 41840 16372 41844
tri 16100 41832 16108 41840 ne
rect 16108 41836 16372 41840
tri 16372 41836 16380 41844 sw
rect 16108 41832 16380 41836
tri 16108 41824 16116 41832 ne
rect 16116 41828 16380 41832
tri 16380 41828 16388 41836 sw
rect 16116 41824 16388 41828
tri 16116 41816 16124 41824 ne
rect 16124 41820 16388 41824
tri 16388 41820 16396 41828 sw
rect 16124 41816 16396 41820
tri 16124 41808 16132 41816 ne
rect 16132 41812 16396 41816
tri 16396 41812 16404 41820 sw
rect 16132 41808 16404 41812
tri 16132 41800 16140 41808 ne
rect 16140 41804 16404 41808
tri 16404 41804 16412 41812 sw
rect 16140 41800 16412 41804
tri 16140 41792 16148 41800 ne
rect 16148 41796 16412 41800
tri 16412 41796 16420 41804 sw
rect 16148 41792 16420 41796
tri 16148 41784 16156 41792 ne
rect 16156 41788 16420 41792
tri 16420 41788 16428 41796 sw
rect 16156 41784 16428 41788
tri 16156 41776 16164 41784 ne
rect 16164 41780 16428 41784
tri 16428 41780 16436 41788 sw
rect 16164 41776 16436 41780
tri 16164 41768 16172 41776 ne
rect 16172 41772 16436 41776
tri 16436 41772 16444 41780 sw
rect 16172 41768 16444 41772
tri 16172 41760 16180 41768 ne
rect 16180 41764 16444 41768
tri 16444 41764 16452 41772 sw
rect 16180 41760 16452 41764
tri 16180 41756 16184 41760 ne
rect 16184 41756 16452 41760
tri 16452 41756 16460 41764 sw
tri 16184 41752 16188 41756 ne
rect 16188 41752 16460 41756
tri 16460 41752 16464 41756 sw
tri 16188 41744 16196 41752 ne
rect 16196 41744 16464 41752
tri 16464 41744 16472 41752 sw
tri 16196 41736 16204 41744 ne
rect 16204 41736 16472 41744
tri 16472 41736 16480 41744 sw
tri 16204 41728 16212 41736 ne
rect 16212 41728 16480 41736
tri 16480 41728 16488 41736 sw
tri 16212 41720 16220 41728 ne
rect 16220 41720 16488 41728
tri 16488 41720 16496 41728 sw
tri 16220 41712 16228 41720 ne
rect 16228 41712 16496 41720
tri 16496 41712 16504 41720 sw
tri 16228 41704 16236 41712 ne
rect 16236 41704 16504 41712
tri 16504 41704 16512 41712 sw
tri 16236 41696 16244 41704 ne
rect 16244 41696 16512 41704
tri 16512 41696 16520 41704 sw
tri 16244 41688 16252 41696 ne
rect 16252 41688 16520 41696
tri 16520 41688 16528 41696 sw
tri 16252 41680 16260 41688 ne
rect 16260 41680 16528 41688
tri 16528 41680 16536 41688 sw
tri 16260 41672 16268 41680 ne
rect 16268 41672 16536 41680
tri 16536 41672 16544 41680 sw
tri 16268 41664 16276 41672 ne
rect 16276 41664 16544 41672
tri 16544 41664 16552 41672 sw
tri 16276 41656 16284 41664 ne
rect 16284 41656 16552 41664
tri 16552 41656 16560 41664 sw
tri 16284 41648 16292 41656 ne
rect 16292 41648 16560 41656
tri 16560 41648 16568 41656 sw
tri 16292 41640 16300 41648 ne
rect 16300 41640 16568 41648
tri 16568 41640 16576 41648 sw
tri 16300 41632 16308 41640 ne
rect 16308 41632 16576 41640
tri 16576 41632 16584 41640 sw
tri 16308 41624 16316 41632 ne
rect 16316 41624 16584 41632
tri 16584 41624 16592 41632 sw
tri 16316 41616 16324 41624 ne
rect 16324 41616 16592 41624
tri 16592 41616 16600 41624 sw
tri 16324 41612 16328 41616 ne
rect 16328 41612 16600 41616
tri 16328 41604 16336 41612 ne
rect 16336 41608 16600 41612
tri 16600 41608 16608 41616 sw
rect 16336 41604 16608 41608
tri 16336 41596 16344 41604 ne
rect 16344 41600 16608 41604
tri 16608 41600 16616 41608 sw
rect 16344 41596 16616 41600
tri 16344 41588 16352 41596 ne
rect 16352 41592 16616 41596
tri 16616 41592 16624 41600 sw
rect 16352 41588 16624 41592
tri 16352 41580 16360 41588 ne
rect 16360 41584 16624 41588
tri 16624 41584 16632 41592 sw
rect 16360 41580 16632 41584
tri 16360 41572 16368 41580 ne
rect 16368 41576 16632 41580
tri 16632 41576 16640 41584 sw
rect 16368 41572 16640 41576
tri 16368 41564 16376 41572 ne
rect 16376 41568 16640 41572
tri 16640 41568 16648 41576 sw
rect 16376 41564 16648 41568
tri 16376 41556 16384 41564 ne
rect 16384 41560 16648 41564
tri 16648 41560 16656 41568 sw
rect 16384 41556 16656 41560
tri 16384 41548 16392 41556 ne
rect 16392 41552 16656 41556
tri 16656 41552 16664 41560 sw
rect 16392 41548 16664 41552
tri 16392 41540 16400 41548 ne
rect 16400 41544 16664 41548
tri 16664 41544 16672 41552 sw
rect 16400 41540 16672 41544
tri 16400 41532 16408 41540 ne
rect 16408 41536 16672 41540
tri 16672 41536 16680 41544 sw
rect 16408 41532 16680 41536
tri 16408 41524 16416 41532 ne
rect 16416 41528 16680 41532
tri 16680 41528 16688 41536 sw
rect 16416 41524 16688 41528
tri 16416 41516 16424 41524 ne
rect 16424 41520 16688 41524
tri 16688 41520 16696 41528 sw
rect 16424 41516 16696 41520
tri 16424 41508 16432 41516 ne
rect 16432 41512 16696 41516
tri 16696 41512 16704 41520 sw
rect 16432 41508 16704 41512
tri 16432 41500 16440 41508 ne
rect 16440 41504 16704 41508
tri 16704 41504 16712 41512 sw
rect 16440 41500 16712 41504
tri 16440 41492 16448 41500 ne
rect 16448 41496 16712 41500
tri 16712 41496 16720 41504 sw
rect 16448 41492 16720 41496
tri 16448 41484 16456 41492 ne
rect 16456 41488 16720 41492
tri 16720 41488 16728 41496 sw
rect 16456 41484 16728 41488
tri 16456 41480 16460 41484 ne
rect 16460 41480 16728 41484
tri 16728 41480 16736 41488 sw
tri 16460 41476 16464 41480 ne
rect 16464 41476 16736 41480
tri 16736 41476 16740 41480 sw
tri 16464 41468 16472 41476 ne
rect 16472 41468 16740 41476
tri 16740 41468 16748 41476 sw
tri 16472 41460 16480 41468 ne
rect 16480 41460 16748 41468
tri 16748 41460 16756 41468 sw
tri 16480 41452 16488 41460 ne
rect 16488 41452 16756 41460
tri 16756 41452 16764 41460 sw
tri 16488 41444 16496 41452 ne
rect 16496 41444 16764 41452
tri 16764 41444 16772 41452 sw
tri 16496 41436 16504 41444 ne
rect 16504 41436 16772 41444
tri 16772 41436 16780 41444 sw
tri 16504 41428 16512 41436 ne
rect 16512 41428 16780 41436
tri 16780 41428 16788 41436 sw
tri 16512 41420 16520 41428 ne
rect 16520 41420 16788 41428
tri 16788 41420 16796 41428 sw
tri 16520 41412 16528 41420 ne
rect 16528 41412 16796 41420
tri 16796 41412 16804 41420 sw
tri 16528 41404 16536 41412 ne
rect 16536 41404 16804 41412
tri 16804 41404 16812 41412 sw
tri 16536 41396 16544 41404 ne
rect 16544 41396 16812 41404
tri 16812 41396 16820 41404 sw
tri 16544 41388 16552 41396 ne
rect 16552 41388 16820 41396
tri 16820 41388 16828 41396 sw
tri 16552 41380 16560 41388 ne
rect 16560 41380 16828 41388
tri 16828 41380 16836 41388 sw
tri 16560 41372 16568 41380 ne
rect 16568 41372 16836 41380
tri 16836 41372 16844 41380 sw
tri 16568 41364 16576 41372 ne
rect 16576 41364 16844 41372
tri 16844 41364 16852 41372 sw
tri 16576 41363 16577 41364 ne
rect 16577 41363 16852 41364
tri 16577 41355 16585 41363 ne
rect 16585 41359 16852 41363
tri 16852 41359 16857 41364 sw
rect 16585 41355 16857 41359
tri 16585 41347 16593 41355 ne
rect 16593 41351 16857 41355
tri 16857 41351 16865 41359 sw
rect 16593 41347 16865 41351
tri 16593 41339 16601 41347 ne
rect 16601 41343 16865 41347
tri 16865 41343 16873 41351 sw
rect 16601 41339 16873 41343
tri 16601 41331 16609 41339 ne
rect 16609 41335 16873 41339
tri 16873 41335 16881 41343 sw
rect 16609 41331 16881 41335
tri 16609 41323 16617 41331 ne
rect 16617 41327 16881 41331
tri 16881 41327 16889 41335 sw
rect 16617 41323 16889 41327
tri 16617 41315 16625 41323 ne
rect 16625 41319 16889 41323
tri 16889 41319 16897 41327 sw
rect 16625 41315 16897 41319
tri 16625 41307 16633 41315 ne
rect 16633 41311 16897 41315
tri 16897 41311 16905 41319 sw
rect 16633 41307 16905 41311
tri 16633 41299 16641 41307 ne
rect 16641 41303 16905 41307
tri 16905 41303 16913 41311 sw
rect 16641 41299 16913 41303
tri 16641 41291 16649 41299 ne
rect 16649 41295 16913 41299
tri 16913 41295 16921 41303 sw
rect 16649 41291 16921 41295
tri 16649 41283 16657 41291 ne
rect 16657 41287 16921 41291
tri 16921 41287 16929 41295 sw
rect 16657 41283 16929 41287
tri 16657 41275 16665 41283 ne
rect 16665 41279 16929 41283
tri 16929 41279 16937 41287 sw
rect 16665 41275 16937 41279
tri 16665 41267 16673 41275 ne
rect 16673 41271 16937 41275
tri 16937 41271 16945 41279 sw
rect 16673 41267 16945 41271
tri 16673 41259 16681 41267 ne
rect 16681 41263 16945 41267
tri 16945 41263 16953 41271 sw
rect 16681 41259 16953 41263
tri 16681 41251 16689 41259 ne
rect 16689 41255 16953 41259
tri 16953 41255 16961 41263 sw
rect 16689 41251 16961 41255
tri 16689 41247 16693 41251 ne
rect 16693 41247 16961 41251
tri 16961 41247 16969 41255 sw
tri 16693 41243 16697 41247 ne
rect 16697 41243 16969 41247
tri 16969 41243 16973 41247 sw
tri 16697 41235 16705 41243 ne
rect 16705 41235 16973 41243
tri 16973 41235 16981 41243 sw
tri 16705 41227 16713 41235 ne
rect 16713 41227 16981 41235
tri 16981 41227 16989 41235 sw
tri 16713 41219 16721 41227 ne
rect 16721 41219 16989 41227
tri 16989 41219 16997 41227 sw
tri 16721 41211 16729 41219 ne
rect 16729 41211 16997 41219
tri 16997 41211 17005 41219 sw
tri 16729 41203 16737 41211 ne
rect 16737 41203 17005 41211
tri 17005 41203 17013 41211 sw
tri 16737 41195 16745 41203 ne
rect 16745 41195 17013 41203
tri 17013 41195 17021 41203 sw
tri 16745 41187 16753 41195 ne
rect 16753 41187 17021 41195
tri 17021 41187 17029 41195 sw
tri 16753 41179 16761 41187 ne
rect 16761 41179 17029 41187
tri 17029 41179 17037 41187 sw
tri 16761 41171 16769 41179 ne
rect 16769 41171 17037 41179
tri 17037 41171 17045 41179 sw
tri 16769 41163 16777 41171 ne
rect 16777 41163 17045 41171
tri 17045 41163 17053 41171 sw
tri 16777 41155 16785 41163 ne
rect 16785 41155 17053 41163
tri 17053 41155 17061 41163 sw
tri 16785 41147 16793 41155 ne
rect 16793 41147 17061 41155
tri 17061 41147 17069 41155 sw
tri 16793 41139 16801 41147 ne
rect 16801 41139 17069 41147
tri 17069 41139 17077 41147 sw
tri 16801 41131 16809 41139 ne
rect 16809 41131 17077 41139
tri 17077 41131 17085 41139 sw
tri 16809 41123 16817 41131 ne
rect 16817 41123 17085 41131
tri 17085 41123 17093 41131 sw
tri 16817 41115 16825 41123 ne
rect 16825 41115 17093 41123
tri 17093 41115 17101 41123 sw
tri 16825 41107 16833 41115 ne
rect 16833 41107 17101 41115
tri 17101 41107 17109 41115 sw
tri 16833 41105 16835 41107 ne
rect 16835 41105 17109 41107
tri 16835 41097 16843 41105 ne
rect 16843 41101 17109 41105
tri 17109 41101 17115 41107 sw
rect 16843 41097 17115 41101
tri 16843 41089 16851 41097 ne
rect 16851 41093 17115 41097
tri 17115 41093 17123 41101 sw
rect 16851 41089 17123 41093
tri 16851 41081 16859 41089 ne
rect 16859 41085 17123 41089
tri 17123 41085 17131 41093 sw
rect 16859 41081 17131 41085
tri 16859 41073 16867 41081 ne
rect 16867 41077 17131 41081
tri 17131 41077 17139 41085 sw
rect 16867 41073 17139 41077
tri 16867 41065 16875 41073 ne
rect 16875 41069 17139 41073
tri 17139 41069 17147 41077 sw
rect 16875 41065 17147 41069
tri 16875 41057 16883 41065 ne
rect 16883 41061 17147 41065
tri 17147 41061 17155 41069 sw
rect 16883 41057 17155 41061
tri 16883 41049 16891 41057 ne
rect 16891 41053 17155 41057
tri 17155 41053 17163 41061 sw
rect 16891 41049 17163 41053
tri 16891 41041 16899 41049 ne
rect 16899 41045 17163 41049
tri 17163 41045 17171 41053 sw
rect 16899 41041 17171 41045
tri 16899 41033 16907 41041 ne
rect 16907 41037 17171 41041
tri 17171 41037 17179 41045 sw
rect 16907 41033 17179 41037
tri 16907 41025 16915 41033 ne
rect 16915 41029 17179 41033
tri 17179 41029 17187 41037 sw
rect 16915 41025 17187 41029
tri 16915 41017 16923 41025 ne
rect 16923 41021 17187 41025
tri 17187 41021 17195 41029 sw
rect 16923 41017 17195 41021
tri 16923 41009 16931 41017 ne
rect 16931 41013 17195 41017
tri 17195 41013 17203 41021 sw
rect 16931 41009 17203 41013
tri 16931 41001 16939 41009 ne
rect 16939 41005 17203 41009
tri 17203 41005 17211 41013 sw
rect 16939 41001 17211 41005
tri 16939 40993 16947 41001 ne
rect 16947 40997 17211 41001
tri 17211 40997 17219 41005 sw
rect 16947 40993 17219 40997
tri 16947 40985 16955 40993 ne
rect 16955 40989 17219 40993
tri 17219 40989 17227 40997 sw
rect 16955 40985 17227 40989
tri 16955 40977 16963 40985 ne
rect 16963 40981 17227 40985
tri 17227 40981 17235 40989 sw
rect 16963 40977 17235 40981
tri 16963 40973 16967 40977 ne
rect 16967 40973 17235 40977
tri 17235 40973 17243 40981 sw
tri 16967 40969 16971 40973 ne
rect 16971 40969 17243 40973
tri 17243 40969 17247 40973 sw
tri 16971 40961 16979 40969 ne
rect 16979 40961 17247 40969
tri 17247 40961 17255 40969 sw
tri 16979 40953 16987 40961 ne
rect 16987 40953 17255 40961
tri 17255 40953 17263 40961 sw
tri 16987 40945 16995 40953 ne
rect 16995 40945 17263 40953
tri 17263 40945 17271 40953 sw
tri 16995 40937 17003 40945 ne
rect 17003 40937 17271 40945
tri 17271 40937 17279 40945 sw
tri 17003 40929 17011 40937 ne
rect 17011 40929 17279 40937
tri 17279 40929 17287 40937 sw
tri 17011 40921 17019 40929 ne
rect 17019 40921 17287 40929
tri 17287 40921 17295 40929 sw
tri 17019 40913 17027 40921 ne
rect 17027 40913 17295 40921
tri 17295 40913 17303 40921 sw
tri 17027 40905 17035 40913 ne
rect 17035 40905 17303 40913
tri 17303 40905 17311 40913 sw
tri 17035 40897 17043 40905 ne
rect 17043 40897 17311 40905
tri 17311 40897 17319 40905 sw
tri 17043 40889 17051 40897 ne
rect 17051 40889 17319 40897
tri 17319 40889 17327 40897 sw
tri 17051 40881 17059 40889 ne
rect 17059 40881 17327 40889
tri 17327 40881 17335 40889 sw
tri 17059 40873 17067 40881 ne
rect 17067 40873 17335 40881
tri 17335 40873 17343 40881 sw
tri 17067 40865 17075 40873 ne
rect 17075 40865 17343 40873
tri 17343 40865 17351 40873 sw
tri 17075 40857 17083 40865 ne
rect 17083 40857 17351 40865
tri 17351 40857 17359 40865 sw
tri 17083 40849 17091 40857 ne
rect 17091 40849 17359 40857
tri 17359 40849 17367 40857 sw
tri 17091 40841 17099 40849 ne
rect 17099 40841 17367 40849
tri 17367 40841 17375 40849 sw
tri 17099 40833 17107 40841 ne
rect 17107 40833 17375 40841
tri 17375 40833 17383 40841 sw
tri 17107 40829 17111 40833 ne
rect 17111 40829 17383 40833
tri 17111 40821 17119 40829 ne
rect 17119 40825 17383 40829
tri 17383 40825 17391 40833 sw
rect 17119 40821 17391 40825
tri 17119 40813 17127 40821 ne
rect 17127 40817 17391 40821
tri 17391 40817 17399 40825 sw
rect 17127 40813 17399 40817
tri 17127 40805 17135 40813 ne
rect 17135 40809 17399 40813
tri 17399 40809 17407 40817 sw
rect 17135 40805 17407 40809
tri 17135 40797 17143 40805 ne
rect 17143 40801 17407 40805
tri 17407 40801 17415 40809 sw
rect 17143 40797 17415 40801
tri 17143 40789 17151 40797 ne
rect 17151 40793 17415 40797
tri 17415 40793 17423 40801 sw
rect 17151 40789 17423 40793
tri 17151 40781 17159 40789 ne
rect 17159 40785 17423 40789
tri 17423 40785 17431 40793 sw
rect 17159 40781 17431 40785
tri 17159 40773 17167 40781 ne
rect 17167 40777 17431 40781
tri 17431 40777 17439 40785 sw
rect 17167 40773 17439 40777
tri 17167 40765 17175 40773 ne
rect 17175 40769 17439 40773
tri 17439 40769 17447 40777 sw
rect 17175 40765 17447 40769
tri 17175 40757 17183 40765 ne
rect 17183 40761 17447 40765
tri 17447 40761 17455 40769 sw
rect 17183 40757 17455 40761
tri 17183 40749 17191 40757 ne
rect 17191 40753 17455 40757
tri 17455 40753 17463 40761 sw
rect 17191 40749 17463 40753
tri 17191 40741 17199 40749 ne
rect 17199 40745 17463 40749
tri 17463 40745 17471 40753 sw
rect 17199 40741 17471 40745
tri 17199 40733 17207 40741 ne
rect 17207 40737 17471 40741
tri 17471 40737 17479 40745 sw
rect 17207 40733 17479 40737
tri 17207 40725 17215 40733 ne
rect 17215 40729 17479 40733
tri 17479 40729 17487 40737 sw
rect 17215 40725 17487 40729
tri 17215 40717 17223 40725 ne
rect 17223 40721 17487 40725
tri 17487 40721 17495 40729 sw
rect 17223 40717 17495 40721
tri 17223 40709 17231 40717 ne
rect 17231 40713 17495 40717
tri 17495 40713 17503 40721 sw
rect 17231 40709 17503 40713
tri 17231 40701 17239 40709 ne
rect 17239 40705 17503 40709
tri 17503 40705 17511 40713 sw
rect 17239 40701 17511 40705
tri 17239 40697 17243 40701 ne
rect 17243 40697 17511 40701
tri 17511 40697 17519 40705 sw
tri 17243 40693 17247 40697 ne
rect 17247 40693 17519 40697
tri 17519 40693 17523 40697 sw
tri 17247 40685 17255 40693 ne
rect 17255 40685 17523 40693
tri 17523 40685 17531 40693 sw
tri 17255 40677 17263 40685 ne
rect 17263 40677 17531 40685
tri 17531 40677 17539 40685 sw
tri 17263 40669 17271 40677 ne
rect 17271 40669 17539 40677
tri 17539 40669 17547 40677 sw
tri 17271 40661 17279 40669 ne
rect 17279 40661 17547 40669
tri 17547 40661 17555 40669 sw
tri 17279 40653 17287 40661 ne
rect 17287 40653 17555 40661
tri 17555 40653 17563 40661 sw
tri 17287 40645 17295 40653 ne
rect 17295 40645 17563 40653
tri 17563 40645 17571 40653 sw
tri 17295 40637 17303 40645 ne
rect 17303 40637 17571 40645
tri 17571 40637 17579 40645 sw
tri 17303 40629 17311 40637 ne
rect 17311 40629 17579 40637
tri 17579 40629 17587 40637 sw
tri 17311 40621 17319 40629 ne
rect 17319 40621 17587 40629
tri 17587 40621 17595 40629 sw
tri 17319 40613 17327 40621 ne
rect 17327 40613 17595 40621
tri 17595 40613 17603 40621 sw
tri 17327 40605 17335 40613 ne
rect 17335 40605 17603 40613
tri 17603 40605 17611 40613 sw
tri 17335 40597 17343 40605 ne
rect 17343 40597 17611 40605
tri 17611 40597 17619 40605 sw
tri 17343 40589 17351 40597 ne
rect 17351 40589 17619 40597
tri 17619 40589 17627 40597 sw
tri 17351 40581 17359 40589 ne
rect 17359 40581 17627 40589
tri 17627 40581 17635 40589 sw
tri 17359 40573 17367 40581 ne
rect 17367 40573 17635 40581
tri 17635 40573 17643 40581 sw
tri 17367 40565 17375 40573 ne
rect 17375 40565 17643 40573
tri 17643 40565 17651 40573 sw
tri 17375 40557 17383 40565 ne
rect 17383 40557 17651 40565
tri 17651 40557 17659 40565 sw
tri 17383 40553 17387 40557 ne
rect 17387 40553 17659 40557
tri 17387 40545 17395 40553 ne
rect 17395 40549 17659 40553
tri 17659 40549 17667 40557 sw
rect 17395 40545 17667 40549
tri 17395 40537 17403 40545 ne
rect 17403 40541 17667 40545
tri 17667 40541 17675 40549 sw
rect 17403 40537 17675 40541
tri 17403 40529 17411 40537 ne
rect 17411 40533 17675 40537
tri 17675 40533 17683 40541 sw
rect 17411 40529 17683 40533
tri 17411 40521 17419 40529 ne
rect 17419 40525 17683 40529
tri 17683 40525 17691 40533 sw
rect 17419 40521 17691 40525
tri 17419 40513 17427 40521 ne
rect 17427 40517 17691 40521
tri 17691 40517 17699 40525 sw
rect 17427 40513 17699 40517
tri 17427 40505 17435 40513 ne
rect 17435 40509 17699 40513
tri 17699 40509 17707 40517 sw
rect 17435 40505 17707 40509
tri 17435 40497 17443 40505 ne
rect 17443 40501 17707 40505
tri 17707 40501 17715 40509 sw
rect 17443 40497 17715 40501
tri 17443 40489 17451 40497 ne
rect 17451 40493 17715 40497
tri 17715 40493 17723 40501 sw
rect 17451 40489 17723 40493
tri 17451 40481 17459 40489 ne
rect 17459 40485 17723 40489
tri 17723 40485 17731 40493 sw
rect 17459 40481 17731 40485
tri 17459 40473 17467 40481 ne
rect 17467 40477 17731 40481
tri 17731 40477 17739 40485 sw
rect 17467 40473 17739 40477
tri 17467 40465 17475 40473 ne
rect 17475 40469 17739 40473
tri 17739 40469 17747 40477 sw
rect 17475 40465 17747 40469
tri 17475 40457 17483 40465 ne
rect 17483 40461 17747 40465
tri 17747 40461 17755 40469 sw
rect 17483 40457 17755 40461
tri 17483 40449 17491 40457 ne
rect 17491 40453 17755 40457
tri 17755 40453 17763 40461 sw
rect 17491 40449 17763 40453
tri 17491 40441 17499 40449 ne
rect 17499 40445 17763 40449
tri 17763 40445 17771 40453 sw
rect 17499 40441 17771 40445
tri 17499 40433 17507 40441 ne
rect 17507 40437 17771 40441
tri 17771 40437 17779 40445 sw
rect 17507 40433 17779 40437
tri 17507 40425 17515 40433 ne
rect 17515 40429 17779 40433
tri 17779 40429 17787 40437 sw
rect 17515 40425 17787 40429
tri 17515 40421 17519 40425 ne
rect 17519 40421 17787 40425
tri 17787 40421 17795 40429 sw
tri 17519 40417 17523 40421 ne
rect 17523 40417 17795 40421
tri 17795 40417 17799 40421 sw
tri 17523 40409 17531 40417 ne
rect 17531 40409 17799 40417
tri 17799 40409 17807 40417 sw
tri 17531 40401 17539 40409 ne
rect 17539 40401 17807 40409
tri 17807 40401 17815 40409 sw
tri 17539 40393 17547 40401 ne
rect 17547 40393 17815 40401
tri 17815 40393 17823 40401 sw
tri 17547 40385 17555 40393 ne
rect 17555 40385 17823 40393
tri 17823 40385 17831 40393 sw
tri 17555 40377 17563 40385 ne
rect 17563 40377 17831 40385
tri 17831 40377 17839 40385 sw
tri 17563 40369 17571 40377 ne
rect 17571 40369 17839 40377
tri 17839 40369 17847 40377 sw
tri 17571 40361 17579 40369 ne
rect 17579 40361 17847 40369
tri 17847 40361 17855 40369 sw
tri 17579 40353 17587 40361 ne
rect 17587 40353 17855 40361
tri 17855 40353 17863 40361 sw
tri 17587 40345 17595 40353 ne
rect 17595 40345 17863 40353
tri 17863 40345 17871 40353 sw
tri 17595 40337 17603 40345 ne
rect 17603 40337 17871 40345
tri 17871 40337 17879 40345 sw
tri 17603 40329 17611 40337 ne
rect 17611 40329 17879 40337
tri 17879 40329 17887 40337 sw
tri 17611 40321 17619 40329 ne
rect 17619 40321 17887 40329
tri 17887 40321 17895 40329 sw
tri 17619 40313 17627 40321 ne
rect 17627 40313 17895 40321
tri 17895 40313 17903 40321 sw
tri 17627 40305 17635 40313 ne
rect 17635 40305 17903 40313
tri 17903 40305 17911 40313 sw
tri 17635 40297 17643 40305 ne
rect 17643 40297 17911 40305
tri 17911 40297 17919 40305 sw
tri 17643 40289 17651 40297 ne
rect 17651 40289 17919 40297
tri 17919 40289 17927 40297 sw
tri 17651 40281 17659 40289 ne
rect 17659 40281 17927 40289
tri 17927 40281 17935 40289 sw
tri 17659 40277 17663 40281 ne
rect 17663 40277 17935 40281
tri 17663 40269 17671 40277 ne
rect 17671 40273 17935 40277
tri 17935 40273 17943 40281 sw
rect 17671 40269 17943 40273
tri 17671 40261 17679 40269 ne
rect 17679 40265 17943 40269
tri 17943 40265 17951 40273 sw
rect 17679 40261 17951 40265
tri 17679 40253 17687 40261 ne
rect 17687 40257 17951 40261
tri 17951 40257 17959 40265 sw
rect 17687 40253 17959 40257
tri 17687 40245 17695 40253 ne
rect 17695 40249 17959 40253
tri 17959 40249 17967 40257 sw
rect 17695 40245 17967 40249
tri 17695 40237 17703 40245 ne
rect 17703 40241 17967 40245
tri 17967 40241 17975 40249 sw
rect 17703 40237 17975 40241
tri 17703 40229 17711 40237 ne
rect 17711 40233 17975 40237
tri 17975 40233 17983 40241 sw
rect 17711 40229 17983 40233
tri 17711 40221 17719 40229 ne
rect 17719 40225 17983 40229
tri 17983 40225 17991 40233 sw
rect 17719 40221 17991 40225
tri 17719 40213 17727 40221 ne
rect 17727 40217 17991 40221
tri 17991 40217 17999 40225 sw
rect 17727 40213 17999 40217
tri 17727 40205 17735 40213 ne
rect 17735 40209 17999 40213
tri 17999 40209 18007 40217 sw
rect 17735 40205 18007 40209
tri 17735 40197 17743 40205 ne
rect 17743 40201 18007 40205
tri 18007 40201 18015 40209 sw
rect 17743 40197 18015 40201
tri 17743 40189 17751 40197 ne
rect 17751 40193 18015 40197
tri 18015 40193 18023 40201 sw
rect 17751 40189 18023 40193
tri 17751 40181 17759 40189 ne
rect 17759 40185 18023 40189
tri 18023 40185 18031 40193 sw
rect 17759 40181 18031 40185
tri 17759 40173 17767 40181 ne
rect 17767 40177 18031 40181
tri 18031 40177 18039 40185 sw
rect 17767 40173 18039 40177
tri 17767 40165 17775 40173 ne
rect 17775 40169 18039 40173
tri 18039 40169 18047 40177 sw
rect 17775 40165 18047 40169
tri 17775 40157 17783 40165 ne
rect 17783 40161 18047 40165
tri 18047 40161 18055 40169 sw
rect 17783 40157 18055 40161
tri 17783 40149 17791 40157 ne
rect 17791 40153 18055 40157
tri 18055 40153 18063 40161 sw
rect 17791 40149 18063 40153
tri 17791 40145 17795 40149 ne
rect 17795 40145 18063 40149
tri 18063 40145 18071 40153 sw
tri 17795 40141 17799 40145 ne
rect 17799 40141 18071 40145
tri 18071 40141 18075 40145 sw
tri 17799 40133 17807 40141 ne
rect 17807 40133 18075 40141
tri 18075 40133 18083 40141 sw
tri 17807 40125 17815 40133 ne
rect 17815 40125 18083 40133
tri 18083 40125 18091 40133 sw
tri 17815 40117 17823 40125 ne
rect 17823 40117 18091 40125
tri 18091 40117 18099 40125 sw
tri 17823 40109 17831 40117 ne
rect 17831 40109 18099 40117
tri 18099 40109 18107 40117 sw
tri 17831 40101 17839 40109 ne
rect 17839 40101 18107 40109
tri 18107 40101 18115 40109 sw
tri 17839 40093 17847 40101 ne
rect 17847 40093 18115 40101
tri 18115 40093 18123 40101 sw
tri 17847 40085 17855 40093 ne
rect 17855 40085 18123 40093
tri 18123 40085 18131 40093 sw
tri 17855 40077 17863 40085 ne
rect 17863 40077 18131 40085
tri 18131 40077 18139 40085 sw
tri 17863 40069 17871 40077 ne
rect 17871 40069 18139 40077
tri 18139 40069 18147 40077 sw
tri 17871 40061 17879 40069 ne
rect 17879 40061 18147 40069
tri 18147 40061 18155 40069 sw
tri 17879 40053 17887 40061 ne
rect 17887 40053 18155 40061
tri 18155 40053 18163 40061 sw
tri 17887 40045 17895 40053 ne
rect 17895 40045 18163 40053
tri 18163 40045 18171 40053 sw
tri 17895 40037 17903 40045 ne
rect 17903 40037 18171 40045
tri 18171 40037 18179 40045 sw
tri 17903 40029 17911 40037 ne
rect 17911 40029 18179 40037
tri 18179 40029 18187 40037 sw
tri 17911 40021 17919 40029 ne
rect 17919 40021 18187 40029
tri 18187 40021 18195 40029 sw
tri 17919 40013 17927 40021 ne
rect 17927 40013 18195 40021
tri 18195 40013 18203 40021 sw
tri 17927 40005 17935 40013 ne
rect 17935 40005 18203 40013
tri 18203 40005 18211 40013 sw
tri 17935 40001 17939 40005 ne
rect 17939 40001 18211 40005
tri 17939 39993 17947 40001 ne
rect 17947 39997 18211 40001
tri 18211 39997 18219 40005 sw
rect 17947 39993 18219 39997
tri 17947 39985 17955 39993 ne
rect 17955 39989 18219 39993
tri 18219 39989 18227 39997 sw
rect 17955 39985 18227 39989
tri 17955 39977 17963 39985 ne
rect 17963 39981 18227 39985
tri 18227 39981 18235 39989 sw
rect 17963 39977 18235 39981
tri 17963 39969 17971 39977 ne
rect 17971 39973 18235 39977
tri 18235 39973 18243 39981 sw
rect 17971 39969 18243 39973
tri 17971 39961 17979 39969 ne
rect 17979 39965 18243 39969
tri 18243 39965 18251 39973 sw
rect 17979 39961 18251 39965
tri 17979 39953 17987 39961 ne
rect 17987 39957 18251 39961
tri 18251 39957 18259 39965 sw
rect 17987 39953 18259 39957
tri 17987 39945 17995 39953 ne
rect 17995 39949 18259 39953
tri 18259 39949 18267 39957 sw
rect 17995 39945 18267 39949
tri 17995 39937 18003 39945 ne
rect 18003 39941 18267 39945
tri 18267 39941 18275 39949 sw
rect 18003 39937 18275 39941
tri 18003 39929 18011 39937 ne
rect 18011 39933 18275 39937
tri 18275 39933 18283 39941 sw
rect 18011 39929 18283 39933
tri 18011 39921 18019 39929 ne
rect 18019 39925 18283 39929
tri 18283 39925 18291 39933 sw
rect 18019 39921 18291 39925
tri 18019 39913 18027 39921 ne
rect 18027 39917 18291 39921
tri 18291 39917 18299 39925 sw
rect 18027 39913 18299 39917
tri 18027 39905 18035 39913 ne
rect 18035 39909 18299 39913
tri 18299 39909 18307 39917 sw
rect 18035 39905 18307 39909
tri 18035 39897 18043 39905 ne
rect 18043 39901 18307 39905
tri 18307 39901 18315 39909 sw
rect 18043 39897 18315 39901
tri 18043 39889 18051 39897 ne
rect 18051 39893 18315 39897
tri 18315 39893 18323 39901 sw
rect 18051 39889 18323 39893
tri 18051 39881 18059 39889 ne
rect 18059 39885 18323 39889
tri 18323 39885 18331 39893 sw
rect 18059 39881 18331 39885
tri 18059 39873 18067 39881 ne
rect 18067 39877 18331 39881
tri 18331 39877 18339 39885 sw
rect 18067 39873 18339 39877
tri 18067 39869 18071 39873 ne
rect 18071 39869 18339 39873
tri 18339 39869 18347 39877 sw
tri 18071 39865 18075 39869 ne
rect 18075 39865 18347 39869
tri 18347 39865 18351 39869 sw
tri 18075 39857 18083 39865 ne
rect 18083 39857 18351 39865
tri 18351 39857 18359 39865 sw
tri 18083 39849 18091 39857 ne
rect 18091 39849 18359 39857
tri 18359 39849 18367 39857 sw
tri 18091 39841 18099 39849 ne
rect 18099 39841 18367 39849
tri 18367 39841 18375 39849 sw
tri 18099 39833 18107 39841 ne
rect 18107 39833 18375 39841
tri 18375 39833 18383 39841 sw
tri 18107 39825 18115 39833 ne
rect 18115 39825 18383 39833
tri 18383 39825 18391 39833 sw
tri 18115 39817 18123 39825 ne
rect 18123 39817 18391 39825
tri 18391 39817 18399 39825 sw
tri 18123 39809 18131 39817 ne
rect 18131 39809 18399 39817
tri 18399 39809 18407 39817 sw
tri 18131 39801 18139 39809 ne
rect 18139 39801 18407 39809
tri 18407 39801 18415 39809 sw
tri 18139 39793 18147 39801 ne
rect 18147 39793 18415 39801
tri 18415 39793 18423 39801 sw
tri 18147 39785 18155 39793 ne
rect 18155 39785 18423 39793
tri 18423 39785 18431 39793 sw
tri 18155 39777 18163 39785 ne
rect 18163 39777 18431 39785
tri 18431 39777 18439 39785 sw
tri 18163 39769 18171 39777 ne
rect 18171 39769 18439 39777
tri 18439 39769 18447 39777 sw
tri 18171 39761 18179 39769 ne
rect 18179 39761 18447 39769
tri 18447 39761 18455 39769 sw
tri 18179 39753 18187 39761 ne
rect 18187 39753 18455 39761
tri 18455 39753 18463 39761 sw
tri 18187 39745 18195 39753 ne
rect 18195 39745 18463 39753
tri 18463 39745 18471 39753 sw
tri 18195 39737 18203 39745 ne
rect 18203 39737 18471 39745
tri 18471 39737 18479 39745 sw
tri 18203 39729 18211 39737 ne
rect 18211 39729 18479 39737
tri 18479 39729 18487 39737 sw
tri 18211 39725 18215 39729 ne
rect 18215 39725 18487 39729
tri 18215 39717 18223 39725 ne
rect 18223 39721 18487 39725
tri 18487 39721 18495 39729 sw
rect 18223 39717 18495 39721
tri 18223 39709 18231 39717 ne
rect 18231 39713 18495 39717
tri 18495 39713 18503 39721 sw
rect 18231 39709 18503 39713
tri 18231 39701 18239 39709 ne
rect 18239 39705 18503 39709
tri 18503 39705 18511 39713 sw
rect 18239 39701 18511 39705
tri 18239 39693 18247 39701 ne
rect 18247 39697 18511 39701
tri 18511 39697 18519 39705 sw
rect 18247 39693 18519 39697
tri 18247 39685 18255 39693 ne
rect 18255 39689 18519 39693
tri 18519 39689 18527 39697 sw
rect 18255 39685 18527 39689
tri 18255 39677 18263 39685 ne
rect 18263 39681 18527 39685
tri 18527 39681 18535 39689 sw
rect 18263 39677 18535 39681
tri 18263 39669 18271 39677 ne
rect 18271 39673 18535 39677
tri 18535 39673 18543 39681 sw
rect 18271 39669 18543 39673
tri 18271 39661 18279 39669 ne
rect 18279 39665 18543 39669
tri 18543 39665 18551 39673 sw
rect 18279 39661 18551 39665
tri 18279 39653 18287 39661 ne
rect 18287 39657 18551 39661
tri 18551 39657 18559 39665 sw
rect 18287 39653 18559 39657
tri 18287 39645 18295 39653 ne
rect 18295 39649 18559 39653
tri 18559 39649 18567 39657 sw
rect 18295 39645 18567 39649
tri 18295 39637 18303 39645 ne
rect 18303 39641 18567 39645
tri 18567 39641 18575 39649 sw
rect 18303 39637 18575 39641
tri 18303 39629 18311 39637 ne
rect 18311 39633 18575 39637
tri 18575 39633 18583 39641 sw
rect 18311 39629 18583 39633
tri 18311 39621 18319 39629 ne
rect 18319 39625 18583 39629
tri 18583 39625 18591 39633 sw
rect 18319 39621 18591 39625
tri 18319 39613 18327 39621 ne
rect 18327 39617 18591 39621
tri 18591 39617 18599 39625 sw
rect 18327 39613 18599 39617
tri 18327 39605 18335 39613 ne
rect 18335 39609 18599 39613
tri 18599 39609 18607 39617 sw
rect 18335 39605 18607 39609
tri 18335 39597 18343 39605 ne
rect 18343 39601 18607 39605
tri 18607 39601 18615 39609 sw
rect 18343 39597 18615 39601
tri 18343 39593 18347 39597 ne
rect 18347 39593 18615 39597
tri 18615 39593 18623 39601 sw
tri 18347 39589 18351 39593 ne
rect 18351 39589 18623 39593
tri 18623 39589 18627 39593 sw
tri 18351 39581 18359 39589 ne
rect 18359 39581 18627 39589
tri 18627 39581 18635 39589 sw
tri 18359 39573 18367 39581 ne
rect 18367 39573 18635 39581
tri 18635 39573 18643 39581 sw
tri 18367 39565 18375 39573 ne
rect 18375 39565 18643 39573
tri 18643 39565 18651 39573 sw
tri 18375 39557 18383 39565 ne
rect 18383 39557 18651 39565
tri 18651 39557 18659 39565 sw
tri 18383 39549 18391 39557 ne
rect 18391 39549 18659 39557
tri 18659 39549 18667 39557 sw
tri 18391 39541 18399 39549 ne
rect 18399 39541 18667 39549
tri 18667 39541 18675 39549 sw
tri 18399 39533 18407 39541 ne
rect 18407 39533 18675 39541
tri 18675 39533 18683 39541 sw
tri 18407 39525 18415 39533 ne
rect 18415 39525 18683 39533
tri 18683 39525 18691 39533 sw
tri 18415 39517 18423 39525 ne
rect 18423 39517 18691 39525
tri 18691 39517 18699 39525 sw
tri 18423 39509 18431 39517 ne
rect 18431 39509 18699 39517
tri 18699 39509 18707 39517 sw
tri 18431 39501 18439 39509 ne
rect 18439 39501 18707 39509
tri 18707 39501 18715 39509 sw
tri 18439 39493 18447 39501 ne
rect 18447 39493 18715 39501
tri 18715 39493 18723 39501 sw
tri 18447 39485 18455 39493 ne
rect 18455 39485 18723 39493
tri 18723 39485 18731 39493 sw
tri 18455 39477 18463 39485 ne
rect 18463 39477 18731 39485
tri 18731 39477 18739 39485 sw
tri 18463 39469 18471 39477 ne
rect 18471 39469 18739 39477
tri 18739 39469 18747 39477 sw
tri 18471 39461 18479 39469 ne
rect 18479 39461 18747 39469
tri 18747 39461 18755 39469 sw
tri 18479 39453 18487 39461 ne
rect 18487 39453 18755 39461
tri 18755 39453 18763 39461 sw
tri 18487 39449 18491 39453 ne
rect 18491 39449 18763 39453
tri 18491 39441 18499 39449 ne
rect 18499 39445 18763 39449
tri 18763 39445 18771 39453 sw
rect 18499 39441 18771 39445
tri 18499 39433 18507 39441 ne
rect 18507 39437 18771 39441
tri 18771 39437 18779 39445 sw
rect 18507 39433 18779 39437
tri 18507 39425 18515 39433 ne
rect 18515 39429 18779 39433
tri 18779 39429 18787 39437 sw
rect 18515 39425 18787 39429
tri 18515 39417 18523 39425 ne
rect 18523 39421 18787 39425
tri 18787 39421 18795 39429 sw
rect 18523 39417 18795 39421
tri 18523 39409 18531 39417 ne
rect 18531 39413 18795 39417
tri 18795 39413 18803 39421 sw
rect 18531 39409 18803 39413
tri 18531 39401 18539 39409 ne
rect 18539 39405 18803 39409
tri 18803 39405 18811 39413 sw
rect 18539 39401 18811 39405
tri 18539 39393 18547 39401 ne
rect 18547 39397 18811 39401
tri 18811 39397 18819 39405 sw
rect 18547 39393 18819 39397
tri 18547 39385 18555 39393 ne
rect 18555 39389 18819 39393
tri 18819 39389 18827 39397 sw
rect 18555 39385 18827 39389
tri 18555 39377 18563 39385 ne
rect 18563 39381 18827 39385
tri 18827 39381 18835 39389 sw
rect 18563 39377 18835 39381
tri 18563 39369 18571 39377 ne
rect 18571 39373 18835 39377
tri 18835 39373 18843 39381 sw
rect 18571 39369 18843 39373
tri 18571 39361 18579 39369 ne
rect 18579 39365 18843 39369
tri 18843 39365 18851 39373 sw
rect 18579 39361 18851 39365
tri 18579 39353 18587 39361 ne
rect 18587 39357 18851 39361
tri 18851 39357 18859 39365 sw
rect 18587 39353 18859 39357
tri 18587 39345 18595 39353 ne
rect 18595 39349 18859 39353
tri 18859 39349 18867 39357 sw
rect 18595 39345 18867 39349
tri 18595 39337 18603 39345 ne
rect 18603 39341 18867 39345
tri 18867 39341 18875 39349 sw
rect 18603 39337 18875 39341
tri 18603 39329 18611 39337 ne
rect 18611 39333 18875 39337
tri 18875 39333 18883 39341 sw
rect 18611 39329 18883 39333
tri 18611 39321 18619 39329 ne
rect 18619 39325 18883 39329
tri 18883 39325 18891 39333 sw
rect 18619 39321 18891 39325
tri 18619 39317 18623 39321 ne
rect 18623 39317 18891 39321
tri 18891 39317 18899 39325 sw
tri 18623 39313 18627 39317 ne
rect 18627 39313 18899 39317
tri 18899 39313 18903 39317 sw
tri 18627 39305 18635 39313 ne
rect 18635 39305 18903 39313
tri 18903 39305 18911 39313 sw
tri 18635 39297 18643 39305 ne
rect 18643 39297 18911 39305
tri 18911 39297 18919 39305 sw
tri 18643 39289 18651 39297 ne
rect 18651 39289 18919 39297
tri 18919 39289 18927 39297 sw
tri 18651 39281 18659 39289 ne
rect 18659 39281 18927 39289
tri 18927 39281 18935 39289 sw
tri 18659 39273 18667 39281 ne
rect 18667 39273 18935 39281
tri 18935 39273 18943 39281 sw
tri 18667 39265 18675 39273 ne
rect 18675 39265 18943 39273
tri 18943 39265 18951 39273 sw
tri 18675 39257 18683 39265 ne
rect 18683 39257 18951 39265
tri 18951 39257 18959 39265 sw
tri 18683 39249 18691 39257 ne
rect 18691 39249 18959 39257
tri 18959 39249 18967 39257 sw
tri 18691 39241 18699 39249 ne
rect 18699 39241 18967 39249
tri 18967 39241 18975 39249 sw
tri 18699 39233 18707 39241 ne
rect 18707 39233 18975 39241
tri 18975 39233 18983 39241 sw
tri 18707 39225 18715 39233 ne
rect 18715 39225 18983 39233
tri 18983 39225 18991 39233 sw
tri 18715 39217 18723 39225 ne
rect 18723 39217 18991 39225
tri 18991 39217 18999 39225 sw
tri 18723 39209 18731 39217 ne
rect 18731 39209 18999 39217
tri 18999 39209 19007 39217 sw
tri 18731 39201 18739 39209 ne
rect 18739 39201 19007 39209
tri 19007 39201 19015 39209 sw
tri 18739 39193 18747 39201 ne
rect 18747 39193 19015 39201
tri 19015 39193 19023 39201 sw
tri 18747 39185 18755 39193 ne
rect 18755 39185 19023 39193
tri 19023 39185 19031 39193 sw
tri 18755 39177 18763 39185 ne
rect 18763 39177 19031 39185
tri 19031 39177 19039 39185 sw
tri 18763 39173 18767 39177 ne
rect 18767 39173 19039 39177
tri 18767 39165 18775 39173 ne
rect 18775 39169 19039 39173
tri 19039 39169 19047 39177 sw
rect 18775 39165 19047 39169
tri 18775 39157 18783 39165 ne
rect 18783 39161 19047 39165
tri 19047 39161 19055 39169 sw
rect 18783 39157 19055 39161
tri 18783 39149 18791 39157 ne
rect 18791 39153 19055 39157
tri 19055 39153 19063 39161 sw
rect 18791 39149 19063 39153
tri 18791 39141 18799 39149 ne
rect 18799 39145 19063 39149
tri 19063 39145 19071 39153 sw
rect 18799 39141 19071 39145
tri 18799 39133 18807 39141 ne
rect 18807 39137 19071 39141
tri 19071 39137 19079 39145 sw
rect 18807 39133 19079 39137
tri 18807 39125 18815 39133 ne
rect 18815 39129 19079 39133
tri 19079 39129 19087 39137 sw
rect 18815 39125 19087 39129
tri 18815 39117 18823 39125 ne
rect 18823 39121 19087 39125
tri 19087 39121 19095 39129 sw
rect 18823 39117 19095 39121
tri 18823 39109 18831 39117 ne
rect 18831 39113 19095 39117
tri 19095 39113 19103 39121 sw
rect 18831 39109 19103 39113
tri 18831 39101 18839 39109 ne
rect 18839 39105 19103 39109
tri 19103 39105 19111 39113 sw
rect 18839 39101 19111 39105
tri 18839 39093 18847 39101 ne
rect 18847 39097 19111 39101
tri 19111 39097 19119 39105 sw
rect 18847 39093 19119 39097
tri 18847 39085 18855 39093 ne
rect 18855 39089 19119 39093
tri 19119 39089 19127 39097 sw
rect 18855 39085 19127 39089
tri 18855 39077 18863 39085 ne
rect 18863 39081 19127 39085
tri 19127 39081 19135 39089 sw
rect 18863 39077 19135 39081
tri 18863 39069 18871 39077 ne
rect 18871 39073 19135 39077
tri 19135 39073 19143 39081 sw
rect 18871 39069 19143 39073
tri 18871 39061 18879 39069 ne
rect 18879 39065 19143 39069
tri 19143 39065 19151 39073 sw
rect 18879 39061 19151 39065
tri 18879 39053 18887 39061 ne
rect 18887 39057 19151 39061
tri 19151 39057 19159 39065 sw
rect 18887 39053 19159 39057
tri 18887 39045 18895 39053 ne
rect 18895 39049 19159 39053
tri 19159 39049 19167 39057 sw
rect 18895 39045 19167 39049
tri 18895 39041 18899 39045 ne
rect 18899 39041 19167 39045
tri 19167 39041 19175 39049 sw
tri 18899 39037 18903 39041 ne
rect 18903 39037 19175 39041
tri 19175 39037 19179 39041 sw
tri 18903 39029 18911 39037 ne
rect 18911 39029 19179 39037
tri 19179 39029 19187 39037 sw
tri 18911 39021 18919 39029 ne
rect 18919 39021 19187 39029
tri 19187 39021 19195 39029 sw
tri 18919 39013 18927 39021 ne
rect 18927 39013 19195 39021
tri 19195 39013 19203 39021 sw
tri 18927 39005 18935 39013 ne
rect 18935 39005 19203 39013
tri 19203 39005 19211 39013 sw
tri 18935 38997 18943 39005 ne
rect 18943 38997 19211 39005
tri 19211 38997 19219 39005 sw
tri 18943 38989 18951 38997 ne
rect 18951 38989 19219 38997
tri 19219 38989 19227 38997 sw
tri 18951 38981 18959 38989 ne
rect 18959 38981 19227 38989
tri 19227 38981 19235 38989 sw
tri 18959 38973 18967 38981 ne
rect 18967 38973 19235 38981
tri 19235 38973 19243 38981 sw
tri 18967 38965 18975 38973 ne
rect 18975 38965 19243 38973
tri 19243 38965 19251 38973 sw
tri 18975 38957 18983 38965 ne
rect 18983 38957 19251 38965
tri 19251 38957 19259 38965 sw
tri 18983 38949 18991 38957 ne
rect 18991 38949 19259 38957
tri 19259 38949 19267 38957 sw
tri 18991 38941 18999 38949 ne
rect 18999 38941 19267 38949
tri 19267 38941 19275 38949 sw
tri 18999 38933 19007 38941 ne
rect 19007 38933 19275 38941
tri 19275 38933 19283 38941 sw
tri 19007 38925 19015 38933 ne
rect 19015 38925 19283 38933
tri 19283 38925 19291 38933 sw
tri 19015 38917 19023 38925 ne
rect 19023 38917 19291 38925
tri 19291 38917 19299 38925 sw
tri 19023 38909 19031 38917 ne
rect 19031 38909 19299 38917
tri 19299 38909 19307 38917 sw
tri 19031 38901 19039 38909 ne
rect 19039 38901 19307 38909
tri 19307 38901 19315 38909 sw
tri 19039 38897 19043 38901 ne
rect 19043 38897 19315 38901
tri 19043 38889 19051 38897 ne
rect 19051 38893 19315 38897
tri 19315 38893 19323 38901 sw
rect 19051 38889 19323 38893
tri 19051 38881 19059 38889 ne
rect 19059 38885 19323 38889
tri 19323 38885 19331 38893 sw
rect 19059 38881 19331 38885
tri 19059 38873 19067 38881 ne
rect 19067 38877 19331 38881
tri 19331 38877 19339 38885 sw
rect 19067 38873 19339 38877
tri 19067 38865 19075 38873 ne
rect 19075 38869 19339 38873
tri 19339 38869 19347 38877 sw
rect 19075 38865 19347 38869
tri 19075 38857 19083 38865 ne
rect 19083 38861 19347 38865
tri 19347 38861 19355 38869 sw
rect 19083 38857 19355 38861
tri 19083 38849 19091 38857 ne
rect 19091 38853 19355 38857
tri 19355 38853 19363 38861 sw
rect 19091 38849 19363 38853
tri 19091 38841 19099 38849 ne
rect 19099 38845 19363 38849
tri 19363 38845 19371 38853 sw
rect 19099 38841 19371 38845
tri 19099 38833 19107 38841 ne
rect 19107 38837 19371 38841
tri 19371 38837 19379 38845 sw
rect 19107 38833 19379 38837
tri 19107 38825 19115 38833 ne
rect 19115 38829 19379 38833
tri 19379 38829 19387 38837 sw
rect 19115 38825 19387 38829
tri 19115 38817 19123 38825 ne
rect 19123 38821 19387 38825
tri 19387 38821 19395 38829 sw
rect 19123 38817 19395 38821
tri 19123 38809 19131 38817 ne
rect 19131 38813 19395 38817
tri 19395 38813 19403 38821 sw
rect 19131 38809 19403 38813
tri 19131 38801 19139 38809 ne
rect 19139 38805 19403 38809
tri 19403 38805 19411 38813 sw
rect 19139 38801 19411 38805
tri 19139 38793 19147 38801 ne
rect 19147 38797 19411 38801
tri 19411 38797 19419 38805 sw
rect 19147 38793 19419 38797
tri 19147 38785 19155 38793 ne
rect 19155 38789 19419 38793
tri 19419 38789 19427 38797 sw
rect 19155 38785 19427 38789
tri 19155 38777 19163 38785 ne
rect 19163 38781 19427 38785
tri 19427 38781 19435 38789 sw
rect 19163 38777 19435 38781
tri 19163 38769 19171 38777 ne
rect 19171 38773 19435 38777
tri 19435 38773 19443 38781 sw
rect 19171 38769 19443 38773
tri 19171 38765 19175 38769 ne
rect 19175 38765 19443 38769
tri 19443 38765 19451 38773 sw
tri 19175 38761 19179 38765 ne
rect 19179 38761 19451 38765
tri 19451 38761 19455 38765 sw
tri 19179 38753 19187 38761 ne
rect 19187 38753 19455 38761
tri 19455 38753 19463 38761 sw
tri 19187 38745 19195 38753 ne
rect 19195 38745 19463 38753
tri 19463 38745 19471 38753 sw
tri 19195 38737 19203 38745 ne
rect 19203 38737 19471 38745
tri 19471 38737 19479 38745 sw
tri 19203 38729 19211 38737 ne
rect 19211 38729 19479 38737
tri 19479 38729 19487 38737 sw
tri 19211 38721 19219 38729 ne
rect 19219 38721 19487 38729
tri 19487 38721 19495 38729 sw
tri 19219 38713 19227 38721 ne
rect 19227 38713 19495 38721
tri 19495 38713 19503 38721 sw
tri 19227 38705 19235 38713 ne
rect 19235 38705 19503 38713
tri 19503 38705 19511 38713 sw
tri 19235 38697 19243 38705 ne
rect 19243 38697 19511 38705
tri 19511 38697 19519 38705 sw
tri 19243 38689 19251 38697 ne
rect 19251 38689 19519 38697
tri 19519 38689 19527 38697 sw
tri 19251 38681 19259 38689 ne
rect 19259 38681 19527 38689
tri 19527 38681 19535 38689 sw
tri 19259 38673 19267 38681 ne
rect 19267 38673 19535 38681
tri 19535 38673 19543 38681 sw
tri 19267 38665 19275 38673 ne
rect 19275 38665 19543 38673
tri 19543 38665 19551 38673 sw
tri 19275 38657 19283 38665 ne
rect 19283 38657 19551 38665
tri 19551 38657 19559 38665 sw
tri 19283 38649 19291 38657 ne
rect 19291 38649 19559 38657
tri 19559 38649 19567 38657 sw
tri 19291 38641 19299 38649 ne
rect 19299 38641 19567 38649
tri 19567 38641 19575 38649 sw
tri 19299 38633 19307 38641 ne
rect 19307 38633 19575 38641
tri 19575 38633 19583 38641 sw
tri 19307 38625 19315 38633 ne
rect 19315 38625 19583 38633
tri 19583 38625 19591 38633 sw
tri 19315 38621 19319 38625 ne
rect 19319 38621 19591 38625
tri 19319 38613 19327 38621 ne
rect 19327 38617 19591 38621
tri 19591 38617 19599 38625 sw
rect 19327 38613 19599 38617
tri 19327 38605 19335 38613 ne
rect 19335 38609 19599 38613
tri 19599 38609 19607 38617 sw
rect 19335 38605 19607 38609
tri 19335 38597 19343 38605 ne
rect 19343 38601 19607 38605
tri 19607 38601 19615 38609 sw
rect 19343 38597 19615 38601
tri 19343 38589 19351 38597 ne
rect 19351 38593 19615 38597
tri 19615 38593 19623 38601 sw
rect 19351 38589 19623 38593
tri 19351 38581 19359 38589 ne
rect 19359 38585 19623 38589
tri 19623 38585 19631 38593 sw
rect 19359 38581 19631 38585
tri 19359 38573 19367 38581 ne
rect 19367 38577 19631 38581
tri 19631 38577 19639 38585 sw
rect 19367 38573 19639 38577
tri 19367 38565 19375 38573 ne
rect 19375 38569 19639 38573
tri 19639 38569 19647 38577 sw
rect 19375 38565 19647 38569
tri 19375 38557 19383 38565 ne
rect 19383 38561 19647 38565
tri 19647 38561 19655 38569 sw
rect 19383 38557 19655 38561
tri 19383 38549 19391 38557 ne
rect 19391 38553 19655 38557
tri 19655 38553 19663 38561 sw
rect 19391 38549 19663 38553
tri 19391 38541 19399 38549 ne
rect 19399 38545 19663 38549
tri 19663 38545 19671 38553 sw
rect 19399 38541 19671 38545
tri 19399 38533 19407 38541 ne
rect 19407 38537 19671 38541
tri 19671 38537 19679 38545 sw
rect 19407 38533 19679 38537
tri 19407 38525 19415 38533 ne
rect 19415 38529 19679 38533
tri 19679 38529 19687 38537 sw
rect 19415 38525 19687 38529
tri 19415 38517 19423 38525 ne
rect 19423 38521 19687 38525
tri 19687 38521 19695 38529 sw
rect 19423 38517 19695 38521
tri 19423 38509 19431 38517 ne
rect 19431 38513 19695 38517
tri 19695 38513 19703 38521 sw
rect 19431 38509 19703 38513
tri 19431 38501 19439 38509 ne
rect 19439 38505 19703 38509
tri 19703 38505 19711 38513 sw
rect 19439 38501 19711 38505
tri 19439 38493 19447 38501 ne
rect 19447 38497 19711 38501
tri 19711 38497 19719 38505 sw
rect 19447 38493 19719 38497
tri 19447 38489 19451 38493 ne
rect 19451 38489 19719 38493
tri 19719 38489 19727 38497 sw
tri 19451 38485 19455 38489 ne
rect 19455 38485 19727 38489
tri 19727 38485 19731 38489 sw
tri 19455 38477 19463 38485 ne
rect 19463 38477 19731 38485
tri 19731 38477 19739 38485 sw
tri 19463 38469 19471 38477 ne
rect 19471 38469 19739 38477
tri 19739 38469 19747 38477 sw
tri 19471 38461 19479 38469 ne
rect 19479 38461 19747 38469
tri 19747 38461 19755 38469 sw
tri 19479 38453 19487 38461 ne
rect 19487 38453 19755 38461
tri 19755 38453 19763 38461 sw
tri 19487 38445 19495 38453 ne
rect 19495 38445 19763 38453
tri 19763 38445 19771 38453 sw
tri 19495 38437 19503 38445 ne
rect 19503 38437 19771 38445
tri 19771 38437 19779 38445 sw
tri 19503 38429 19511 38437 ne
rect 19511 38429 19779 38437
tri 19779 38429 19787 38437 sw
tri 19511 38421 19519 38429 ne
rect 19519 38421 19787 38429
tri 19787 38421 19795 38429 sw
tri 19519 38413 19527 38421 ne
rect 19527 38413 19795 38421
tri 19795 38413 19803 38421 sw
tri 19527 38405 19535 38413 ne
rect 19535 38405 19803 38413
tri 19803 38405 19811 38413 sw
tri 19535 38397 19543 38405 ne
rect 19543 38397 19811 38405
tri 19811 38397 19819 38405 sw
tri 19543 38389 19551 38397 ne
rect 19551 38389 19819 38397
tri 19819 38389 19827 38397 sw
tri 19551 38381 19559 38389 ne
rect 19559 38381 19827 38389
tri 19827 38381 19835 38389 sw
tri 19559 38373 19567 38381 ne
rect 19567 38373 19835 38381
tri 19835 38373 19843 38381 sw
tri 19567 38365 19575 38373 ne
rect 19575 38365 19843 38373
tri 19843 38365 19851 38373 sw
tri 19575 38357 19583 38365 ne
rect 19583 38357 19851 38365
tri 19851 38357 19859 38365 sw
tri 19583 38349 19591 38357 ne
rect 19591 38349 19859 38357
tri 19859 38349 19867 38357 sw
tri 19591 38345 19595 38349 ne
rect 19595 38345 19867 38349
tri 19595 38337 19603 38345 ne
rect 19603 38341 19867 38345
tri 19867 38341 19875 38349 sw
rect 19603 38337 19875 38341
tri 19603 38329 19611 38337 ne
rect 19611 38333 19875 38337
tri 19875 38333 19883 38341 sw
rect 19611 38329 19883 38333
tri 19611 38321 19619 38329 ne
rect 19619 38325 19883 38329
tri 19883 38325 19891 38333 sw
rect 19619 38321 19891 38325
tri 19619 38313 19627 38321 ne
rect 19627 38317 19891 38321
tri 19891 38317 19899 38325 sw
rect 19627 38313 19899 38317
tri 19627 38305 19635 38313 ne
rect 19635 38309 19899 38313
tri 19899 38309 19907 38317 sw
rect 19635 38305 19907 38309
tri 19635 38297 19643 38305 ne
rect 19643 38301 19907 38305
tri 19907 38301 19915 38309 sw
rect 19643 38297 19915 38301
tri 19643 38289 19651 38297 ne
rect 19651 38293 19915 38297
tri 19915 38293 19923 38301 sw
rect 19651 38289 19923 38293
tri 19651 38281 19659 38289 ne
rect 19659 38285 19923 38289
tri 19923 38285 19931 38293 sw
rect 19659 38281 19931 38285
tri 19659 38273 19667 38281 ne
rect 19667 38277 19931 38281
tri 19931 38277 19939 38285 sw
rect 19667 38273 19939 38277
tri 19667 38265 19675 38273 ne
rect 19675 38269 19939 38273
tri 19939 38269 19947 38277 sw
rect 19675 38265 19947 38269
tri 19675 38257 19683 38265 ne
rect 19683 38261 19947 38265
tri 19947 38261 19955 38269 sw
rect 19683 38257 19955 38261
tri 19683 38249 19691 38257 ne
rect 19691 38253 19955 38257
tri 19955 38253 19963 38261 sw
rect 19691 38249 19963 38253
tri 19691 38241 19699 38249 ne
rect 19699 38245 19963 38249
tri 19963 38245 19971 38253 sw
rect 19699 38241 19971 38245
tri 19699 38233 19707 38241 ne
rect 19707 38237 19971 38241
tri 19971 38237 19979 38245 sw
rect 19707 38233 19979 38237
tri 19707 38225 19715 38233 ne
rect 19715 38229 19979 38233
tri 19979 38229 19987 38237 sw
rect 19715 38225 19987 38229
tri 19715 38217 19723 38225 ne
rect 19723 38221 19987 38225
tri 19987 38221 19995 38229 sw
rect 19723 38217 19995 38221
tri 19723 38213 19727 38217 ne
rect 19727 38213 19995 38217
tri 19995 38213 20003 38221 sw
tri 19727 38209 19731 38213 ne
rect 19731 38209 20003 38213
tri 20003 38209 20007 38213 sw
tri 19731 38201 19739 38209 ne
rect 19739 38201 20007 38209
tri 20007 38201 20015 38209 sw
tri 19739 38193 19747 38201 ne
rect 19747 38193 20015 38201
tri 20015 38193 20023 38201 sw
tri 19747 38185 19755 38193 ne
rect 19755 38185 20023 38193
tri 20023 38185 20031 38193 sw
tri 19755 38177 19763 38185 ne
rect 19763 38177 20031 38185
tri 20031 38177 20039 38185 sw
tri 19763 38169 19771 38177 ne
rect 19771 38169 20039 38177
tri 20039 38169 20047 38177 sw
tri 19771 38161 19779 38169 ne
rect 19779 38161 20047 38169
tri 20047 38161 20055 38169 sw
tri 19779 38153 19787 38161 ne
rect 19787 38153 20055 38161
tri 20055 38153 20063 38161 sw
tri 19787 38145 19795 38153 ne
rect 19795 38145 20063 38153
tri 20063 38145 20071 38153 sw
tri 19795 38137 19803 38145 ne
rect 19803 38137 20071 38145
tri 20071 38137 20079 38145 sw
tri 19803 38129 19811 38137 ne
rect 19811 38129 20079 38137
tri 20079 38129 20087 38137 sw
tri 19811 38121 19819 38129 ne
rect 19819 38121 20087 38129
tri 20087 38121 20095 38129 sw
tri 19819 38113 19827 38121 ne
rect 19827 38113 20095 38121
tri 20095 38113 20103 38121 sw
tri 19827 38105 19835 38113 ne
rect 19835 38105 20103 38113
tri 20103 38105 20111 38113 sw
tri 19835 38097 19843 38105 ne
rect 19843 38097 20111 38105
tri 20111 38097 20119 38105 sw
tri 19843 38089 19851 38097 ne
rect 19851 38089 20119 38097
tri 20119 38089 20127 38097 sw
tri 19851 38081 19859 38089 ne
rect 19859 38081 20127 38089
tri 20127 38081 20135 38089 sw
tri 19859 38073 19867 38081 ne
rect 19867 38073 20135 38081
tri 20135 38073 20143 38081 sw
tri 19867 38069 19871 38073 ne
rect 19871 38069 20143 38073
tri 19871 38061 19879 38069 ne
rect 19879 38065 20143 38069
tri 20143 38065 20151 38073 sw
rect 19879 38061 20151 38065
tri 19879 38053 19887 38061 ne
rect 19887 38057 20151 38061
tri 20151 38057 20159 38065 sw
rect 19887 38053 20159 38057
tri 19887 38045 19895 38053 ne
rect 19895 38049 20159 38053
tri 20159 38049 20167 38057 sw
rect 19895 38045 20167 38049
tri 19895 38037 19903 38045 ne
rect 19903 38041 20167 38045
tri 20167 38041 20175 38049 sw
rect 19903 38037 20175 38041
tri 19903 38029 19911 38037 ne
rect 19911 38033 20175 38037
tri 20175 38033 20183 38041 sw
rect 19911 38029 20183 38033
tri 19911 38021 19919 38029 ne
rect 19919 38025 20183 38029
tri 20183 38025 20191 38033 sw
rect 19919 38021 20191 38025
tri 19919 38013 19927 38021 ne
rect 19927 38017 20191 38021
tri 20191 38017 20199 38025 sw
rect 19927 38013 20199 38017
tri 19927 38005 19935 38013 ne
rect 19935 38009 20199 38013
tri 20199 38009 20207 38017 sw
rect 19935 38005 20207 38009
tri 19935 37997 19943 38005 ne
rect 19943 38001 20207 38005
tri 20207 38001 20215 38009 sw
rect 19943 37997 20215 38001
tri 19943 37989 19951 37997 ne
rect 19951 37993 20215 37997
tri 20215 37993 20223 38001 sw
rect 19951 37989 20223 37993
tri 19951 37981 19959 37989 ne
rect 19959 37985 20223 37989
tri 20223 37985 20231 37993 sw
rect 19959 37981 20231 37985
tri 19959 37973 19967 37981 ne
rect 19967 37977 20231 37981
tri 20231 37977 20239 37985 sw
rect 19967 37973 20239 37977
tri 19967 37965 19975 37973 ne
rect 19975 37969 20239 37973
tri 20239 37969 20247 37977 sw
rect 19975 37965 20247 37969
tri 19975 37957 19983 37965 ne
rect 19983 37961 20247 37965
tri 20247 37961 20255 37969 sw
rect 19983 37957 20255 37961
tri 19983 37949 19991 37957 ne
rect 19991 37953 20255 37957
tri 20255 37953 20263 37961 sw
rect 19991 37949 20263 37953
tri 19991 37941 19999 37949 ne
rect 19999 37945 20263 37949
tri 20263 37945 20271 37953 sw
rect 19999 37941 20271 37945
tri 19999 37937 20003 37941 ne
rect 20003 37937 20271 37941
tri 20271 37937 20279 37945 sw
tri 20003 37933 20007 37937 ne
rect 20007 37933 20279 37937
tri 20279 37933 20283 37937 sw
tri 20007 37925 20015 37933 ne
rect 20015 37925 20283 37933
tri 20283 37925 20291 37933 sw
tri 20015 37917 20023 37925 ne
rect 20023 37917 20291 37925
tri 20291 37917 20299 37925 sw
tri 20023 37909 20031 37917 ne
rect 20031 37909 20299 37917
tri 20299 37909 20307 37917 sw
tri 20031 37901 20039 37909 ne
rect 20039 37901 20307 37909
tri 20307 37901 20315 37909 sw
tri 20039 37893 20047 37901 ne
rect 20047 37893 20315 37901
tri 20315 37893 20323 37901 sw
tri 20047 37885 20055 37893 ne
rect 20055 37885 20323 37893
tri 20323 37885 20331 37893 sw
tri 20055 37877 20063 37885 ne
rect 20063 37877 20331 37885
tri 20331 37877 20339 37885 sw
tri 20063 37869 20071 37877 ne
rect 20071 37869 20339 37877
tri 20339 37869 20347 37877 sw
tri 20071 37861 20079 37869 ne
rect 20079 37861 20347 37869
tri 20347 37861 20355 37869 sw
tri 20079 37853 20087 37861 ne
rect 20087 37853 20355 37861
tri 20355 37853 20363 37861 sw
tri 20087 37845 20095 37853 ne
rect 20095 37845 20363 37853
tri 20363 37845 20371 37853 sw
tri 20095 37837 20103 37845 ne
rect 20103 37837 20371 37845
tri 20371 37837 20379 37845 sw
tri 20103 37829 20111 37837 ne
rect 20111 37829 20379 37837
tri 20379 37829 20387 37837 sw
tri 20111 37821 20119 37829 ne
rect 20119 37821 20387 37829
tri 20387 37821 20395 37829 sw
tri 20119 37813 20127 37821 ne
rect 20127 37813 20395 37821
tri 20395 37813 20403 37821 sw
tri 20127 37805 20135 37813 ne
rect 20135 37805 20403 37813
tri 20403 37805 20411 37813 sw
tri 20135 37797 20143 37805 ne
rect 20143 37797 20411 37805
tri 20411 37797 20419 37805 sw
tri 20143 37793 20147 37797 ne
rect 20147 37793 20419 37797
tri 20147 37785 20155 37793 ne
rect 20155 37789 20419 37793
tri 20419 37789 20427 37797 sw
rect 20155 37785 20427 37789
tri 20155 37777 20163 37785 ne
rect 20163 37781 20427 37785
tri 20427 37781 20435 37789 sw
rect 20163 37777 20435 37781
tri 20163 37769 20171 37777 ne
rect 20171 37773 20435 37777
tri 20435 37773 20443 37781 sw
rect 20171 37769 20443 37773
tri 20171 37761 20179 37769 ne
rect 20179 37765 20443 37769
tri 20443 37765 20451 37773 sw
rect 20179 37761 20451 37765
tri 20179 37753 20187 37761 ne
rect 20187 37757 20451 37761
tri 20451 37757 20459 37765 sw
rect 20187 37753 20459 37757
tri 20187 37745 20195 37753 ne
rect 20195 37749 20459 37753
tri 20459 37749 20467 37757 sw
rect 20195 37745 20467 37749
tri 20195 37737 20203 37745 ne
rect 20203 37741 20467 37745
tri 20467 37741 20475 37749 sw
rect 20203 37737 20475 37741
tri 20203 37729 20211 37737 ne
rect 20211 37733 20475 37737
tri 20475 37733 20483 37741 sw
rect 20211 37729 20483 37733
tri 20211 37721 20219 37729 ne
rect 20219 37725 20483 37729
tri 20483 37725 20491 37733 sw
rect 20219 37721 20491 37725
tri 20219 37713 20227 37721 ne
rect 20227 37717 20491 37721
tri 20491 37717 20499 37725 sw
rect 20227 37713 20499 37717
tri 20227 37705 20235 37713 ne
rect 20235 37709 20499 37713
tri 20499 37709 20507 37717 sw
rect 20235 37705 20507 37709
tri 20235 37697 20243 37705 ne
rect 20243 37701 20507 37705
tri 20507 37701 20515 37709 sw
rect 20243 37697 20515 37701
tri 20243 37689 20251 37697 ne
rect 20251 37693 20515 37697
tri 20515 37693 20523 37701 sw
rect 20251 37689 20523 37693
tri 20251 37681 20259 37689 ne
rect 20259 37685 20523 37689
tri 20523 37685 20531 37693 sw
rect 20259 37681 20531 37685
tri 20259 37673 20267 37681 ne
rect 20267 37677 20531 37681
tri 20531 37677 20539 37685 sw
rect 20267 37673 20539 37677
tri 20267 37665 20275 37673 ne
rect 20275 37669 20539 37673
tri 20539 37669 20547 37677 sw
rect 20275 37665 20547 37669
tri 20275 37661 20279 37665 ne
rect 20279 37661 20547 37665
tri 20547 37661 20555 37669 sw
tri 20279 37657 20283 37661 ne
rect 20283 37657 20555 37661
tri 20555 37657 20559 37661 sw
tri 20283 37649 20291 37657 ne
rect 20291 37649 20559 37657
tri 20559 37649 20567 37657 sw
tri 20291 37641 20299 37649 ne
rect 20299 37641 20567 37649
tri 20567 37641 20575 37649 sw
tri 20299 37633 20307 37641 ne
rect 20307 37633 20575 37641
tri 20575 37633 20583 37641 sw
tri 20307 37625 20315 37633 ne
rect 20315 37625 20583 37633
tri 20583 37625 20591 37633 sw
tri 20315 37617 20323 37625 ne
rect 20323 37617 20591 37625
tri 20591 37617 20599 37625 sw
tri 20323 37609 20331 37617 ne
rect 20331 37609 20599 37617
tri 20599 37609 20607 37617 sw
tri 20331 37601 20339 37609 ne
rect 20339 37601 20607 37609
tri 20607 37601 20615 37609 sw
tri 20339 37593 20347 37601 ne
rect 20347 37593 20615 37601
tri 20615 37593 20623 37601 sw
tri 20347 37585 20355 37593 ne
rect 20355 37585 20623 37593
tri 20623 37585 20631 37593 sw
tri 20355 37577 20363 37585 ne
rect 20363 37577 20631 37585
tri 20631 37577 20639 37585 sw
tri 20363 37569 20371 37577 ne
rect 20371 37569 20639 37577
tri 20639 37569 20647 37577 sw
tri 20371 37561 20379 37569 ne
rect 20379 37561 20647 37569
tri 20647 37561 20655 37569 sw
tri 20379 37553 20387 37561 ne
rect 20387 37553 20655 37561
tri 20655 37553 20663 37561 sw
tri 20387 37545 20395 37553 ne
rect 20395 37545 20663 37553
tri 20663 37545 20671 37553 sw
tri 20395 37537 20403 37545 ne
rect 20403 37537 20671 37545
tri 20671 37537 20679 37545 sw
tri 20403 37529 20411 37537 ne
rect 20411 37529 20679 37537
tri 20679 37529 20687 37537 sw
tri 20411 37521 20419 37529 ne
rect 20419 37521 20687 37529
tri 20687 37521 20695 37529 sw
tri 20419 37517 20423 37521 ne
rect 20423 37517 20695 37521
tri 20423 37509 20431 37517 ne
rect 20431 37513 20695 37517
tri 20695 37513 20703 37521 sw
rect 20431 37509 20703 37513
tri 20431 37501 20439 37509 ne
rect 20439 37505 20703 37509
tri 20703 37505 20711 37513 sw
rect 20439 37501 20711 37505
tri 20439 37493 20447 37501 ne
rect 20447 37497 20711 37501
tri 20711 37497 20719 37505 sw
rect 20447 37493 20719 37497
tri 20447 37485 20455 37493 ne
rect 20455 37489 20719 37493
tri 20719 37489 20727 37497 sw
rect 20455 37485 20727 37489
tri 20455 37477 20463 37485 ne
rect 20463 37481 20727 37485
tri 20727 37481 20735 37489 sw
rect 20463 37477 20735 37481
tri 20463 37469 20471 37477 ne
rect 20471 37473 20735 37477
tri 20735 37473 20743 37481 sw
rect 20471 37469 20743 37473
tri 20471 37461 20479 37469 ne
rect 20479 37465 20743 37469
tri 20743 37465 20751 37473 sw
rect 20479 37461 20751 37465
tri 20479 37453 20487 37461 ne
rect 20487 37457 20751 37461
tri 20751 37457 20759 37465 sw
rect 20487 37453 20759 37457
tri 20487 37445 20495 37453 ne
rect 20495 37449 20759 37453
tri 20759 37449 20767 37457 sw
rect 20495 37445 20767 37449
tri 20495 37437 20503 37445 ne
rect 20503 37441 20767 37445
tri 20767 37441 20775 37449 sw
rect 20503 37437 20775 37441
tri 20503 37429 20511 37437 ne
rect 20511 37433 20775 37437
tri 20775 37433 20783 37441 sw
rect 20511 37429 20783 37433
tri 20511 37421 20519 37429 ne
rect 20519 37425 20783 37429
tri 20783 37425 20791 37433 sw
rect 20519 37421 20791 37425
tri 20519 37413 20527 37421 ne
rect 20527 37417 20791 37421
tri 20791 37417 20799 37425 sw
rect 20527 37413 20799 37417
tri 20527 37405 20535 37413 ne
rect 20535 37409 20799 37413
tri 20799 37409 20807 37417 sw
rect 20535 37405 20807 37409
tri 20535 37397 20543 37405 ne
rect 20543 37401 20807 37405
tri 20807 37401 20815 37409 sw
rect 20543 37397 20815 37401
tri 20543 37389 20551 37397 ne
rect 20551 37393 20815 37397
tri 20815 37393 20823 37401 sw
rect 20551 37389 20823 37393
tri 20551 37385 20555 37389 ne
rect 20555 37385 20823 37389
tri 20823 37385 20831 37393 sw
tri 20555 37381 20559 37385 ne
rect 20559 37381 20831 37385
tri 20831 37381 20835 37385 sw
tri 20559 37373 20567 37381 ne
rect 20567 37373 20835 37381
tri 20835 37373 20843 37381 sw
tri 20567 37365 20575 37373 ne
rect 20575 37365 20843 37373
tri 20843 37365 20851 37373 sw
tri 20575 37357 20583 37365 ne
rect 20583 37357 20851 37365
tri 20851 37357 20859 37365 sw
tri 20583 37349 20591 37357 ne
rect 20591 37349 20859 37357
tri 20859 37349 20867 37357 sw
tri 20591 37341 20599 37349 ne
rect 20599 37341 20867 37349
tri 20867 37341 20875 37349 sw
tri 20599 37333 20607 37341 ne
rect 20607 37333 20875 37341
tri 20875 37333 20883 37341 sw
tri 20607 37325 20615 37333 ne
rect 20615 37325 20883 37333
tri 20883 37325 20891 37333 sw
tri 20615 37317 20623 37325 ne
rect 20623 37317 20891 37325
tri 20891 37317 20899 37325 sw
tri 20623 37309 20631 37317 ne
rect 20631 37309 20899 37317
tri 20899 37309 20907 37317 sw
tri 20631 37301 20639 37309 ne
rect 20639 37301 20907 37309
tri 20907 37301 20915 37309 sw
tri 20639 37293 20647 37301 ne
rect 20647 37293 20915 37301
tri 20915 37293 20923 37301 sw
tri 20647 37285 20655 37293 ne
rect 20655 37285 20923 37293
tri 20923 37285 20931 37293 sw
tri 20655 37277 20663 37285 ne
rect 20663 37277 20931 37285
tri 20931 37277 20939 37285 sw
tri 20663 37269 20671 37277 ne
rect 20671 37269 20939 37277
tri 20939 37269 20947 37277 sw
tri 20671 37261 20679 37269 ne
rect 20679 37261 20947 37269
tri 20947 37261 20955 37269 sw
tri 20679 37253 20687 37261 ne
rect 20687 37253 20955 37261
tri 20955 37253 20963 37261 sw
tri 20687 37245 20695 37253 ne
rect 20695 37245 20963 37253
tri 20963 37245 20971 37253 sw
tri 20695 37241 20699 37245 ne
rect 20699 37241 20971 37245
tri 20699 37233 20707 37241 ne
rect 20707 37237 20971 37241
tri 20971 37237 20979 37245 sw
rect 20707 37233 20979 37237
tri 20707 37225 20715 37233 ne
rect 20715 37229 20979 37233
tri 20979 37229 20987 37237 sw
rect 20715 37225 20987 37229
tri 20715 37217 20723 37225 ne
rect 20723 37221 20987 37225
tri 20987 37221 20995 37229 sw
rect 20723 37217 20995 37221
tri 20723 37209 20731 37217 ne
rect 20731 37213 20995 37217
tri 20995 37213 21003 37221 sw
rect 20731 37209 21003 37213
tri 20731 37201 20739 37209 ne
rect 20739 37205 21003 37209
tri 21003 37205 21011 37213 sw
rect 20739 37201 21011 37205
tri 20739 37193 20747 37201 ne
rect 20747 37197 21011 37201
tri 21011 37197 21019 37205 sw
rect 20747 37193 21019 37197
tri 20747 37185 20755 37193 ne
rect 20755 37189 21019 37193
tri 21019 37189 21027 37197 sw
rect 20755 37185 21027 37189
tri 20755 37177 20763 37185 ne
rect 20763 37181 21027 37185
tri 21027 37181 21035 37189 sw
rect 20763 37177 21035 37181
tri 20763 37169 20771 37177 ne
rect 20771 37173 21035 37177
tri 21035 37173 21043 37181 sw
rect 20771 37169 21043 37173
tri 20771 37161 20779 37169 ne
rect 20779 37165 21043 37169
tri 21043 37165 21051 37173 sw
rect 20779 37161 21051 37165
tri 20779 37153 20787 37161 ne
rect 20787 37157 21051 37161
tri 21051 37157 21059 37165 sw
rect 20787 37153 21059 37157
tri 20787 37145 20795 37153 ne
rect 20795 37149 21059 37153
tri 21059 37149 21067 37157 sw
rect 20795 37145 21067 37149
tri 20795 37137 20803 37145 ne
rect 20803 37141 21067 37145
tri 21067 37141 21075 37149 sw
rect 20803 37137 21075 37141
tri 20803 37129 20811 37137 ne
rect 20811 37133 21075 37137
tri 21075 37133 21083 37141 sw
rect 20811 37129 21083 37133
tri 20811 37121 20819 37129 ne
rect 20819 37125 21083 37129
tri 21083 37125 21091 37133 sw
rect 20819 37121 21091 37125
tri 20819 37113 20827 37121 ne
rect 20827 37117 21091 37121
tri 21091 37117 21099 37125 sw
rect 20827 37113 21099 37117
tri 20827 37109 20831 37113 ne
rect 20831 37109 21099 37113
tri 21099 37109 21107 37117 sw
tri 20831 37105 20835 37109 ne
rect 20835 37105 21107 37109
tri 21107 37105 21111 37109 sw
tri 20835 37097 20843 37105 ne
rect 20843 37097 21111 37105
tri 21111 37097 21119 37105 sw
tri 20843 37089 20851 37097 ne
rect 20851 37089 21119 37097
tri 21119 37089 21127 37097 sw
tri 20851 37081 20859 37089 ne
rect 20859 37081 21127 37089
tri 21127 37081 21135 37089 sw
tri 20859 37073 20867 37081 ne
rect 20867 37073 21135 37081
tri 21135 37073 21143 37081 sw
tri 20867 37065 20875 37073 ne
rect 20875 37065 21143 37073
tri 21143 37065 21151 37073 sw
tri 20875 37057 20883 37065 ne
rect 20883 37057 21151 37065
tri 21151 37057 21159 37065 sw
tri 20883 37049 20891 37057 ne
rect 20891 37049 21159 37057
tri 21159 37049 21167 37057 sw
tri 20891 37041 20899 37049 ne
rect 20899 37041 21167 37049
tri 21167 37041 21175 37049 sw
tri 20899 37033 20907 37041 ne
rect 20907 37033 21175 37041
tri 21175 37033 21183 37041 sw
tri 20907 37025 20915 37033 ne
rect 20915 37025 21183 37033
tri 21183 37025 21191 37033 sw
tri 20915 37017 20923 37025 ne
rect 20923 37017 21191 37025
tri 21191 37017 21199 37025 sw
tri 20923 37009 20931 37017 ne
rect 20931 37009 21199 37017
tri 21199 37009 21207 37017 sw
tri 20931 37001 20939 37009 ne
rect 20939 37001 21207 37009
tri 21207 37001 21215 37009 sw
tri 20939 36993 20947 37001 ne
rect 20947 36993 21215 37001
tri 21215 36993 21223 37001 sw
tri 20947 36985 20955 36993 ne
rect 20955 36985 21223 36993
tri 21223 36985 21231 36993 sw
tri 20955 36977 20963 36985 ne
rect 20963 36977 21231 36985
tri 21231 36977 21239 36985 sw
tri 20963 36969 20971 36977 ne
rect 20971 36969 21239 36977
tri 21239 36969 21247 36977 sw
tri 20971 36965 20975 36969 ne
rect 20975 36965 21247 36969
tri 20975 36957 20983 36965 ne
rect 20983 36961 21247 36965
tri 21247 36961 21255 36969 sw
rect 20983 36957 21255 36961
tri 20983 36949 20991 36957 ne
rect 20991 36953 21255 36957
tri 21255 36953 21263 36961 sw
rect 20991 36949 21263 36953
tri 20991 36941 20999 36949 ne
rect 20999 36945 21263 36949
tri 21263 36945 21271 36953 sw
rect 20999 36941 21271 36945
tri 20999 36933 21007 36941 ne
rect 21007 36937 21271 36941
tri 21271 36937 21279 36945 sw
rect 21007 36933 21279 36937
tri 21007 36925 21015 36933 ne
rect 21015 36929 21279 36933
tri 21279 36929 21287 36937 sw
rect 21015 36925 21287 36929
tri 21015 36917 21023 36925 ne
rect 21023 36921 21287 36925
tri 21287 36921 21295 36929 sw
rect 21023 36917 21295 36921
tri 21023 36909 21031 36917 ne
rect 21031 36913 21295 36917
tri 21295 36913 21303 36921 sw
rect 21031 36909 21303 36913
tri 21031 36901 21039 36909 ne
rect 21039 36905 21303 36909
tri 21303 36905 21311 36913 sw
rect 21039 36901 21311 36905
tri 21039 36893 21047 36901 ne
rect 21047 36897 21311 36901
tri 21311 36897 21319 36905 sw
rect 21047 36893 21319 36897
tri 21047 36885 21055 36893 ne
rect 21055 36889 21319 36893
tri 21319 36889 21327 36897 sw
rect 21055 36885 21327 36889
tri 21055 36877 21063 36885 ne
rect 21063 36881 21327 36885
tri 21327 36881 21335 36889 sw
rect 21063 36877 21335 36881
tri 21063 36869 21071 36877 ne
rect 21071 36873 21335 36877
tri 21335 36873 21343 36881 sw
rect 21071 36869 21343 36873
tri 21071 36861 21079 36869 ne
rect 21079 36865 21343 36869
tri 21343 36865 21351 36873 sw
rect 21079 36861 21351 36865
tri 21079 36853 21087 36861 ne
rect 21087 36857 21351 36861
tri 21351 36857 21359 36865 sw
rect 21087 36853 21359 36857
tri 21087 36845 21095 36853 ne
rect 21095 36849 21359 36853
tri 21359 36849 21367 36857 sw
rect 21095 36845 21367 36849
tri 21095 36837 21103 36845 ne
rect 21103 36841 21367 36845
tri 21367 36841 21375 36849 sw
rect 21103 36837 21375 36841
tri 21103 36833 21107 36837 ne
rect 21107 36833 21375 36837
tri 21375 36833 21383 36841 sw
tri 21107 36829 21111 36833 ne
rect 21111 36829 21383 36833
tri 21383 36829 21387 36833 sw
tri 21111 36821 21119 36829 ne
rect 21119 36821 21387 36829
tri 21387 36821 21395 36829 sw
tri 21119 36813 21127 36821 ne
rect 21127 36813 21395 36821
tri 21395 36813 21403 36821 sw
tri 21127 36805 21135 36813 ne
rect 21135 36805 21403 36813
tri 21403 36805 21411 36813 sw
tri 21135 36797 21143 36805 ne
rect 21143 36797 21411 36805
tri 21411 36797 21419 36805 sw
tri 21143 36789 21151 36797 ne
rect 21151 36789 21419 36797
tri 21419 36789 21427 36797 sw
tri 21151 36781 21159 36789 ne
rect 21159 36781 21427 36789
tri 21427 36781 21435 36789 sw
tri 21159 36773 21167 36781 ne
rect 21167 36773 21435 36781
tri 21435 36773 21443 36781 sw
tri 21167 36765 21175 36773 ne
rect 21175 36765 21443 36773
tri 21443 36765 21451 36773 sw
tri 21175 36757 21183 36765 ne
rect 21183 36757 21451 36765
tri 21451 36757 21459 36765 sw
tri 21183 36749 21191 36757 ne
rect 21191 36749 21459 36757
tri 21459 36749 21467 36757 sw
tri 21191 36741 21199 36749 ne
rect 21199 36741 21467 36749
tri 21467 36741 21475 36749 sw
tri 21199 36733 21207 36741 ne
rect 21207 36733 21475 36741
tri 21475 36733 21483 36741 sw
tri 21207 36725 21215 36733 ne
rect 21215 36725 21483 36733
tri 21483 36725 21491 36733 sw
tri 21215 36717 21223 36725 ne
rect 21223 36717 21491 36725
tri 21491 36717 21499 36725 sw
tri 21223 36709 21231 36717 ne
rect 21231 36709 21499 36717
tri 21499 36709 21507 36717 sw
tri 21231 36701 21239 36709 ne
rect 21239 36701 21507 36709
tri 21507 36701 21515 36709 sw
tri 21239 36693 21247 36701 ne
rect 21247 36693 21515 36701
tri 21515 36693 21523 36701 sw
tri 21247 36689 21251 36693 ne
rect 21251 36689 21523 36693
tri 21251 36681 21259 36689 ne
rect 21259 36685 21523 36689
tri 21523 36685 21531 36693 sw
rect 21259 36681 21531 36685
tri 21259 36673 21267 36681 ne
rect 21267 36677 21531 36681
tri 21531 36677 21539 36685 sw
rect 21267 36673 21539 36677
tri 21267 36665 21275 36673 ne
rect 21275 36669 21539 36673
tri 21539 36669 21547 36677 sw
rect 21275 36665 21547 36669
tri 21275 36657 21283 36665 ne
rect 21283 36661 21547 36665
tri 21547 36661 21555 36669 sw
rect 21283 36657 21555 36661
tri 21283 36649 21291 36657 ne
rect 21291 36653 21555 36657
tri 21555 36653 21563 36661 sw
rect 21291 36649 21563 36653
tri 21291 36641 21299 36649 ne
rect 21299 36645 21563 36649
tri 21563 36645 21571 36653 sw
rect 21299 36641 21571 36645
tri 21299 36633 21307 36641 ne
rect 21307 36637 21571 36641
tri 21571 36637 21579 36645 sw
rect 21307 36633 21579 36637
tri 21307 36625 21315 36633 ne
rect 21315 36629 21579 36633
tri 21579 36629 21587 36637 sw
rect 21315 36625 21587 36629
tri 21315 36617 21323 36625 ne
rect 21323 36621 21587 36625
tri 21587 36621 21595 36629 sw
rect 21323 36617 21595 36621
tri 21323 36609 21331 36617 ne
rect 21331 36613 21595 36617
tri 21595 36613 21603 36621 sw
rect 21331 36609 21603 36613
tri 21331 36601 21339 36609 ne
rect 21339 36605 21603 36609
tri 21603 36605 21611 36613 sw
rect 21339 36601 21611 36605
tri 21339 36593 21347 36601 ne
rect 21347 36597 21611 36601
tri 21611 36597 21619 36605 sw
rect 21347 36593 21619 36597
tri 21347 36585 21355 36593 ne
rect 21355 36589 21619 36593
tri 21619 36589 21627 36597 sw
rect 21355 36585 21627 36589
tri 21355 36577 21363 36585 ne
rect 21363 36581 21627 36585
tri 21627 36581 21635 36589 sw
rect 21363 36577 21635 36581
tri 21363 36569 21371 36577 ne
rect 21371 36573 21635 36577
tri 21635 36573 21643 36581 sw
rect 21371 36569 21643 36573
tri 21371 36561 21379 36569 ne
rect 21379 36565 21643 36569
tri 21643 36565 21651 36573 sw
rect 21379 36561 21651 36565
tri 21379 36557 21383 36561 ne
rect 21383 36557 21651 36561
tri 21651 36557 21659 36565 sw
tri 21383 36553 21387 36557 ne
rect 21387 36553 21659 36557
tri 21659 36553 21663 36557 sw
tri 21387 36545 21395 36553 ne
rect 21395 36545 21663 36553
tri 21663 36545 21671 36553 sw
tri 21395 36537 21403 36545 ne
rect 21403 36537 21671 36545
tri 21671 36537 21679 36545 sw
tri 21403 36529 21411 36537 ne
rect 21411 36529 21679 36537
tri 21679 36529 21687 36537 sw
tri 21411 36521 21419 36529 ne
rect 21419 36521 21687 36529
tri 21687 36521 21695 36529 sw
tri 21419 36513 21427 36521 ne
rect 21427 36513 21695 36521
tri 21695 36513 21703 36521 sw
tri 21427 36505 21435 36513 ne
rect 21435 36505 21703 36513
tri 21703 36505 21711 36513 sw
tri 21435 36497 21443 36505 ne
rect 21443 36497 21711 36505
tri 21711 36497 21719 36505 sw
tri 21443 36489 21451 36497 ne
rect 21451 36489 21719 36497
tri 21719 36489 21727 36497 sw
tri 21451 36481 21459 36489 ne
rect 21459 36481 21727 36489
tri 21727 36481 21735 36489 sw
tri 21459 36473 21467 36481 ne
rect 21467 36473 21735 36481
tri 21735 36473 21743 36481 sw
tri 21467 36465 21475 36473 ne
rect 21475 36465 21743 36473
tri 21743 36465 21751 36473 sw
tri 21475 36457 21483 36465 ne
rect 21483 36457 21751 36465
tri 21751 36457 21759 36465 sw
tri 21483 36449 21491 36457 ne
rect 21491 36449 21759 36457
tri 21759 36449 21767 36457 sw
tri 21491 36441 21499 36449 ne
rect 21499 36441 21767 36449
tri 21767 36441 21775 36449 sw
tri 21499 36433 21507 36441 ne
rect 21507 36433 21775 36441
tri 21775 36433 21783 36441 sw
tri 21507 36425 21515 36433 ne
rect 21515 36425 21783 36433
tri 21783 36425 21791 36433 sw
tri 21515 36417 21523 36425 ne
rect 21523 36417 21791 36425
tri 21791 36417 21799 36425 sw
tri 21523 36413 21527 36417 ne
rect 21527 36413 21799 36417
tri 21527 36405 21535 36413 ne
rect 21535 36409 21799 36413
tri 21799 36409 21807 36417 sw
rect 21535 36405 21807 36409
tri 21535 36397 21543 36405 ne
rect 21543 36401 21807 36405
tri 21807 36401 21815 36409 sw
rect 21543 36397 21815 36401
tri 21543 36389 21551 36397 ne
rect 21551 36393 21815 36397
tri 21815 36393 21823 36401 sw
rect 21551 36389 21823 36393
tri 21551 36381 21559 36389 ne
rect 21559 36385 21823 36389
tri 21823 36385 21831 36393 sw
rect 21559 36381 21831 36385
tri 21559 36373 21567 36381 ne
rect 21567 36377 21831 36381
tri 21831 36377 21839 36385 sw
rect 21567 36373 21839 36377
tri 21567 36365 21575 36373 ne
rect 21575 36369 21839 36373
tri 21839 36369 21847 36377 sw
rect 21575 36365 21847 36369
tri 21575 36357 21583 36365 ne
rect 21583 36361 21847 36365
tri 21847 36361 21855 36369 sw
rect 21583 36357 21855 36361
tri 21583 36349 21591 36357 ne
rect 21591 36353 21855 36357
tri 21855 36353 21863 36361 sw
rect 21591 36349 21863 36353
tri 21591 36341 21599 36349 ne
rect 21599 36345 21863 36349
tri 21863 36345 21871 36353 sw
rect 21599 36341 21871 36345
tri 21599 36333 21607 36341 ne
rect 21607 36337 21871 36341
tri 21871 36337 21879 36345 sw
rect 21607 36333 21879 36337
tri 21607 36325 21615 36333 ne
rect 21615 36329 21879 36333
tri 21879 36329 21887 36337 sw
rect 21615 36325 21887 36329
tri 21615 36317 21623 36325 ne
rect 21623 36321 21887 36325
tri 21887 36321 21895 36329 sw
rect 21623 36317 21895 36321
tri 21623 36309 21631 36317 ne
rect 21631 36313 21895 36317
tri 21895 36313 21903 36321 sw
rect 21631 36309 21903 36313
tri 21631 36301 21639 36309 ne
rect 21639 36305 21903 36309
tri 21903 36305 21911 36313 sw
rect 21639 36301 21911 36305
tri 21639 36293 21647 36301 ne
rect 21647 36297 21911 36301
tri 21911 36297 21919 36305 sw
rect 21647 36293 21919 36297
tri 21647 36285 21655 36293 ne
rect 21655 36289 21919 36293
tri 21919 36289 21927 36297 sw
rect 21655 36285 21927 36289
tri 21655 36281 21659 36285 ne
rect 21659 36281 21927 36285
tri 21927 36281 21935 36289 sw
tri 21659 36277 21663 36281 ne
rect 21663 36277 21935 36281
tri 21935 36277 21939 36281 sw
tri 21663 36269 21671 36277 ne
rect 21671 36269 21939 36277
tri 21939 36269 21947 36277 sw
tri 21671 36261 21679 36269 ne
rect 21679 36261 21947 36269
tri 21947 36261 21955 36269 sw
tri 21679 36253 21687 36261 ne
rect 21687 36253 21955 36261
tri 21955 36253 21963 36261 sw
tri 21687 36245 21695 36253 ne
rect 21695 36245 21963 36253
tri 21963 36245 21971 36253 sw
tri 21695 36237 21703 36245 ne
rect 21703 36237 21971 36245
tri 21971 36237 21979 36245 sw
tri 21703 36229 21711 36237 ne
rect 21711 36229 21979 36237
tri 21979 36229 21987 36237 sw
tri 21711 36221 21719 36229 ne
rect 21719 36221 21987 36229
tri 21987 36221 21995 36229 sw
tri 21719 36213 21727 36221 ne
rect 21727 36213 21995 36221
tri 21995 36213 22003 36221 sw
tri 21727 36205 21735 36213 ne
rect 21735 36205 22003 36213
tri 22003 36205 22011 36213 sw
tri 21735 36197 21743 36205 ne
rect 21743 36197 22011 36205
tri 22011 36197 22019 36205 sw
tri 21743 36189 21751 36197 ne
rect 21751 36189 22019 36197
tri 22019 36189 22027 36197 sw
tri 21751 36181 21759 36189 ne
rect 21759 36181 22027 36189
tri 22027 36181 22035 36189 sw
tri 21759 36173 21767 36181 ne
rect 21767 36173 22035 36181
tri 22035 36173 22043 36181 sw
tri 21767 36165 21775 36173 ne
rect 21775 36165 22043 36173
tri 22043 36165 22051 36173 sw
tri 21775 36157 21783 36165 ne
rect 21783 36157 22051 36165
tri 22051 36157 22059 36165 sw
tri 21783 36149 21791 36157 ne
rect 21791 36149 22059 36157
tri 22059 36149 22067 36157 sw
tri 21791 36141 21799 36149 ne
rect 21799 36141 22067 36149
tri 22067 36141 22075 36149 sw
tri 21799 36137 21803 36141 ne
rect 21803 36137 22075 36141
tri 21803 36129 21811 36137 ne
rect 21811 36133 22075 36137
tri 22075 36133 22083 36141 sw
rect 21811 36129 22083 36133
tri 21811 36121 21819 36129 ne
rect 21819 36125 22083 36129
tri 22083 36125 22091 36133 sw
rect 21819 36121 22091 36125
tri 21819 36113 21827 36121 ne
rect 21827 36117 22091 36121
tri 22091 36117 22099 36125 sw
rect 21827 36113 22099 36117
tri 21827 36105 21835 36113 ne
rect 21835 36109 22099 36113
tri 22099 36109 22107 36117 sw
rect 21835 36105 22107 36109
tri 21835 36097 21843 36105 ne
rect 21843 36101 22107 36105
tri 22107 36101 22115 36109 sw
rect 21843 36097 22115 36101
tri 21843 36089 21851 36097 ne
rect 21851 36093 22115 36097
tri 22115 36093 22123 36101 sw
rect 21851 36089 22123 36093
tri 21851 36081 21859 36089 ne
rect 21859 36085 22123 36089
tri 22123 36085 22131 36093 sw
rect 21859 36081 22131 36085
tri 21859 36073 21867 36081 ne
rect 21867 36077 22131 36081
tri 22131 36077 22139 36085 sw
rect 21867 36073 22139 36077
tri 21867 36065 21875 36073 ne
rect 21875 36069 22139 36073
tri 22139 36069 22147 36077 sw
rect 21875 36065 22147 36069
tri 21875 36057 21883 36065 ne
rect 21883 36061 22147 36065
tri 22147 36061 22155 36069 sw
rect 21883 36057 22155 36061
tri 21883 36049 21891 36057 ne
rect 21891 36053 22155 36057
tri 22155 36053 22163 36061 sw
rect 21891 36049 22163 36053
tri 21891 36041 21899 36049 ne
rect 21899 36045 22163 36049
tri 22163 36045 22171 36053 sw
rect 21899 36041 22171 36045
tri 21899 36033 21907 36041 ne
rect 21907 36037 22171 36041
tri 22171 36037 22179 36045 sw
rect 21907 36033 22179 36037
tri 21907 36025 21915 36033 ne
rect 21915 36029 22179 36033
tri 22179 36029 22187 36037 sw
rect 21915 36025 22187 36029
tri 21915 36017 21923 36025 ne
rect 21923 36021 22187 36025
tri 22187 36021 22195 36029 sw
rect 21923 36017 22195 36021
tri 21923 36009 21931 36017 ne
rect 21931 36013 22195 36017
tri 22195 36013 22203 36021 sw
rect 21931 36009 22203 36013
tri 21931 36005 21935 36009 ne
rect 21935 36005 22203 36009
tri 22203 36005 22211 36013 sw
tri 21935 36001 21939 36005 ne
rect 21939 36001 22211 36005
tri 22211 36001 22215 36005 sw
tri 21939 35993 21947 36001 ne
rect 21947 35993 22215 36001
tri 22215 35993 22223 36001 sw
tri 21947 35985 21955 35993 ne
rect 21955 35985 22223 35993
tri 22223 35985 22231 35993 sw
tri 21955 35977 21963 35985 ne
rect 21963 35977 22231 35985
tri 22231 35977 22239 35985 sw
tri 21963 35969 21971 35977 ne
rect 21971 35969 22239 35977
tri 22239 35969 22247 35977 sw
tri 21971 35961 21979 35969 ne
rect 21979 35961 22247 35969
tri 22247 35961 22255 35969 sw
tri 21979 35953 21987 35961 ne
rect 21987 35953 22255 35961
tri 22255 35953 22263 35961 sw
tri 21987 35945 21995 35953 ne
rect 21995 35945 22263 35953
tri 22263 35945 22271 35953 sw
tri 21995 35937 22003 35945 ne
rect 22003 35937 22271 35945
tri 22271 35937 22279 35945 sw
tri 22003 35929 22011 35937 ne
rect 22011 35929 22279 35937
tri 22279 35929 22287 35937 sw
tri 22011 35921 22019 35929 ne
rect 22019 35921 22287 35929
tri 22287 35921 22295 35929 sw
tri 22019 35913 22027 35921 ne
rect 22027 35913 22295 35921
tri 22295 35913 22303 35921 sw
tri 22027 35905 22035 35913 ne
rect 22035 35905 22303 35913
tri 22303 35905 22311 35913 sw
tri 22035 35897 22043 35905 ne
rect 22043 35897 22311 35905
tri 22311 35897 22319 35905 sw
tri 22043 35889 22051 35897 ne
rect 22051 35889 22319 35897
tri 22319 35889 22327 35897 sw
tri 22051 35881 22059 35889 ne
rect 22059 35881 22327 35889
tri 22327 35881 22335 35889 sw
tri 22059 35873 22067 35881 ne
rect 22067 35873 22335 35881
tri 22335 35873 22343 35881 sw
tri 22067 35865 22075 35873 ne
rect 22075 35865 22343 35873
tri 22343 35865 22351 35873 sw
tri 22075 35861 22079 35865 ne
rect 22079 35861 22351 35865
tri 22079 35853 22087 35861 ne
rect 22087 35857 22351 35861
tri 22351 35857 22359 35865 sw
rect 22087 35853 22359 35857
tri 22087 35845 22095 35853 ne
rect 22095 35849 22359 35853
tri 22359 35849 22367 35857 sw
rect 22095 35845 22367 35849
tri 22095 35837 22103 35845 ne
rect 22103 35841 22367 35845
tri 22367 35841 22375 35849 sw
rect 22103 35837 22375 35841
tri 22103 35829 22111 35837 ne
rect 22111 35833 22375 35837
tri 22375 35833 22383 35841 sw
rect 22111 35829 22383 35833
tri 22111 35821 22119 35829 ne
rect 22119 35825 22383 35829
tri 22383 35825 22391 35833 sw
rect 22119 35821 22391 35825
tri 22119 35813 22127 35821 ne
rect 22127 35817 22391 35821
tri 22391 35817 22399 35825 sw
rect 22127 35813 22399 35817
tri 22127 35805 22135 35813 ne
rect 22135 35809 22399 35813
tri 22399 35809 22407 35817 sw
rect 22135 35805 22407 35809
tri 22135 35797 22143 35805 ne
rect 22143 35801 22407 35805
tri 22407 35801 22415 35809 sw
rect 22143 35797 22415 35801
tri 22143 35789 22151 35797 ne
rect 22151 35793 22415 35797
tri 22415 35793 22423 35801 sw
rect 22151 35789 22423 35793
tri 22151 35781 22159 35789 ne
rect 22159 35785 22423 35789
tri 22423 35785 22431 35793 sw
rect 22159 35781 22431 35785
tri 22159 35773 22167 35781 ne
rect 22167 35777 22431 35781
tri 22431 35777 22439 35785 sw
rect 22167 35773 22439 35777
tri 22167 35765 22175 35773 ne
rect 22175 35769 22439 35773
tri 22439 35769 22447 35777 sw
rect 22175 35765 22447 35769
tri 22175 35757 22183 35765 ne
rect 22183 35761 22447 35765
tri 22447 35761 22455 35769 sw
rect 22183 35757 22455 35761
tri 22183 35749 22191 35757 ne
rect 22191 35753 22455 35757
tri 22455 35753 22463 35761 sw
rect 22191 35749 22463 35753
tri 22191 35741 22199 35749 ne
rect 22199 35745 22463 35749
tri 22463 35745 22471 35753 sw
rect 22199 35741 22471 35745
tri 22199 35733 22207 35741 ne
rect 22207 35737 22471 35741
tri 22471 35737 22479 35745 sw
rect 22207 35733 22479 35737
tri 22207 35729 22211 35733 ne
rect 22211 35729 22479 35733
tri 22479 35729 22487 35737 sw
tri 22211 35725 22215 35729 ne
rect 22215 35725 22487 35729
tri 22487 35725 22491 35729 sw
tri 22215 35717 22223 35725 ne
rect 22223 35717 22491 35725
tri 22491 35717 22499 35725 sw
tri 22223 35709 22231 35717 ne
rect 22231 35709 22499 35717
tri 22499 35709 22507 35717 sw
tri 22231 35701 22239 35709 ne
rect 22239 35701 22507 35709
tri 22507 35701 22515 35709 sw
tri 22239 35693 22247 35701 ne
rect 22247 35693 22515 35701
tri 22515 35693 22523 35701 sw
tri 22247 35685 22255 35693 ne
rect 22255 35685 22523 35693
tri 22523 35685 22531 35693 sw
tri 22255 35677 22263 35685 ne
rect 22263 35677 22531 35685
tri 22531 35677 22539 35685 sw
tri 22263 35669 22271 35677 ne
rect 22271 35669 22539 35677
tri 22539 35669 22547 35677 sw
tri 22271 35661 22279 35669 ne
rect 22279 35661 22547 35669
tri 22547 35661 22555 35669 sw
tri 22279 35653 22287 35661 ne
rect 22287 35653 22555 35661
tri 22555 35653 22563 35661 sw
tri 22287 35645 22295 35653 ne
rect 22295 35645 22563 35653
tri 22563 35645 22571 35653 sw
tri 22295 35637 22303 35645 ne
rect 22303 35637 22571 35645
tri 22571 35637 22579 35645 sw
tri 22303 35629 22311 35637 ne
rect 22311 35629 22579 35637
tri 22579 35629 22587 35637 sw
tri 22311 35621 22319 35629 ne
rect 22319 35621 22587 35629
tri 22587 35621 22595 35629 sw
tri 22319 35613 22327 35621 ne
rect 22327 35613 22595 35621
tri 22595 35613 22603 35621 sw
tri 22327 35605 22335 35613 ne
rect 22335 35605 22603 35613
tri 22603 35605 22611 35613 sw
tri 22335 35597 22343 35605 ne
rect 22343 35597 22611 35605
tri 22611 35597 22619 35605 sw
tri 22343 35589 22351 35597 ne
rect 22351 35589 22619 35597
tri 22619 35589 22627 35597 sw
tri 22351 35585 22355 35589 ne
rect 22355 35585 22627 35589
tri 22355 35577 22363 35585 ne
rect 22363 35581 22627 35585
tri 22627 35581 22635 35589 sw
rect 22363 35577 22635 35581
tri 22363 35569 22371 35577 ne
rect 22371 35573 22635 35577
tri 22635 35573 22643 35581 sw
rect 22371 35569 22643 35573
tri 22371 35561 22379 35569 ne
rect 22379 35565 22643 35569
tri 22643 35565 22651 35573 sw
rect 22379 35561 22651 35565
tri 22379 35553 22387 35561 ne
rect 22387 35557 22651 35561
tri 22651 35557 22659 35565 sw
rect 22387 35553 22659 35557
tri 22387 35545 22395 35553 ne
rect 22395 35549 22659 35553
tri 22659 35549 22667 35557 sw
rect 22395 35545 22667 35549
tri 22395 35537 22403 35545 ne
rect 22403 35541 22667 35545
tri 22667 35541 22675 35549 sw
rect 22403 35537 22675 35541
tri 22403 35529 22411 35537 ne
rect 22411 35533 22675 35537
tri 22675 35533 22683 35541 sw
rect 22411 35529 22683 35533
tri 22411 35521 22419 35529 ne
rect 22419 35525 22683 35529
tri 22683 35525 22691 35533 sw
rect 22419 35521 22691 35525
tri 22419 35513 22427 35521 ne
rect 22427 35517 22691 35521
tri 22691 35517 22699 35525 sw
rect 22427 35513 22699 35517
tri 22427 35505 22435 35513 ne
rect 22435 35509 22699 35513
tri 22699 35509 22707 35517 sw
rect 22435 35505 22707 35509
tri 22435 35497 22443 35505 ne
rect 22443 35501 22707 35505
tri 22707 35501 22715 35509 sw
rect 22443 35497 22715 35501
tri 22443 35489 22451 35497 ne
rect 22451 35493 22715 35497
tri 22715 35493 22723 35501 sw
rect 22451 35489 22723 35493
tri 22451 35481 22459 35489 ne
rect 22459 35485 22723 35489
tri 22723 35485 22731 35493 sw
rect 22459 35481 22731 35485
tri 22459 35473 22467 35481 ne
rect 22467 35477 22731 35481
tri 22731 35477 22739 35485 sw
rect 22467 35473 22739 35477
tri 22467 35465 22475 35473 ne
rect 22475 35469 22739 35473
tri 22739 35469 22747 35477 sw
rect 22475 35465 22747 35469
tri 22475 35457 22483 35465 ne
rect 22483 35461 22747 35465
tri 22747 35461 22755 35469 sw
rect 22483 35457 22755 35461
tri 22483 35453 22487 35457 ne
rect 22487 35453 22755 35457
tri 22755 35453 22763 35461 sw
tri 22487 35449 22491 35453 ne
rect 22491 35449 22763 35453
tri 22763 35449 22767 35453 sw
tri 22491 35441 22499 35449 ne
rect 22499 35441 22767 35449
tri 22767 35441 22775 35449 sw
tri 22499 35433 22507 35441 ne
rect 22507 35433 22775 35441
tri 22775 35433 22783 35441 sw
tri 22507 35425 22515 35433 ne
rect 22515 35425 22783 35433
tri 22783 35425 22791 35433 sw
tri 22515 35417 22523 35425 ne
rect 22523 35417 22791 35425
tri 22791 35417 22799 35425 sw
tri 22523 35409 22531 35417 ne
rect 22531 35409 22799 35417
tri 22799 35409 22807 35417 sw
tri 22531 35401 22539 35409 ne
rect 22539 35401 22807 35409
tri 22807 35401 22815 35409 sw
tri 22539 35393 22547 35401 ne
rect 22547 35393 22815 35401
tri 22815 35393 22823 35401 sw
tri 22547 35385 22555 35393 ne
rect 22555 35385 22823 35393
tri 22823 35385 22831 35393 sw
tri 22555 35377 22563 35385 ne
rect 22563 35377 22831 35385
tri 22831 35377 22839 35385 sw
tri 22563 35369 22571 35377 ne
rect 22571 35369 22839 35377
tri 22839 35369 22847 35377 sw
tri 22571 35361 22579 35369 ne
rect 22579 35361 22847 35369
tri 22847 35361 22855 35369 sw
tri 22579 35353 22587 35361 ne
rect 22587 35353 22855 35361
tri 22855 35353 22863 35361 sw
tri 22587 35345 22595 35353 ne
rect 22595 35345 22863 35353
tri 22863 35345 22871 35353 sw
tri 22595 35337 22603 35345 ne
rect 22603 35337 22871 35345
tri 22871 35337 22879 35345 sw
tri 22603 35329 22611 35337 ne
rect 22611 35329 22879 35337
tri 22879 35329 22887 35337 sw
tri 22611 35321 22619 35329 ne
rect 22619 35321 22887 35329
tri 22887 35321 22895 35329 sw
tri 22619 35313 22627 35321 ne
rect 22627 35313 22895 35321
tri 22895 35313 22903 35321 sw
tri 22627 35309 22631 35313 ne
rect 22631 35309 22903 35313
tri 22631 35301 22639 35309 ne
rect 22639 35305 22903 35309
tri 22903 35305 22911 35313 sw
rect 22639 35301 22911 35305
tri 22639 35293 22647 35301 ne
rect 22647 35297 22911 35301
tri 22911 35297 22919 35305 sw
rect 22647 35293 22919 35297
tri 22647 35285 22655 35293 ne
rect 22655 35289 22919 35293
tri 22919 35289 22927 35297 sw
rect 22655 35285 22927 35289
tri 22655 35277 22663 35285 ne
rect 22663 35281 22927 35285
tri 22927 35281 22935 35289 sw
rect 22663 35277 22935 35281
tri 22663 35269 22671 35277 ne
rect 22671 35273 22935 35277
tri 22935 35273 22943 35281 sw
rect 22671 35269 22943 35273
tri 22671 35261 22679 35269 ne
rect 22679 35265 22943 35269
tri 22943 35265 22951 35273 sw
rect 22679 35261 22951 35265
tri 22679 35253 22687 35261 ne
rect 22687 35257 22951 35261
tri 22951 35257 22959 35265 sw
rect 22687 35253 22959 35257
tri 22687 35245 22695 35253 ne
rect 22695 35249 22959 35253
tri 22959 35249 22967 35257 sw
rect 22695 35245 22967 35249
tri 22695 35237 22703 35245 ne
rect 22703 35241 22967 35245
tri 22967 35241 22975 35249 sw
rect 22703 35237 22975 35241
tri 22703 35229 22711 35237 ne
rect 22711 35233 22975 35237
tri 22975 35233 22983 35241 sw
rect 22711 35229 22983 35233
tri 22711 35221 22719 35229 ne
rect 22719 35225 22983 35229
tri 22983 35225 22991 35233 sw
rect 22719 35221 22991 35225
tri 22719 35213 22727 35221 ne
rect 22727 35217 22991 35221
tri 22991 35217 22999 35225 sw
rect 22727 35213 22999 35217
tri 22727 35205 22735 35213 ne
rect 22735 35209 22999 35213
tri 22999 35209 23007 35217 sw
rect 22735 35205 23007 35209
tri 22735 35197 22743 35205 ne
rect 22743 35201 23007 35205
tri 23007 35201 23015 35209 sw
rect 22743 35197 23015 35201
tri 22743 35189 22751 35197 ne
rect 22751 35193 23015 35197
tri 23015 35193 23023 35201 sw
rect 22751 35189 23023 35193
tri 22751 35181 22759 35189 ne
rect 22759 35185 23023 35189
tri 23023 35185 23031 35193 sw
rect 22759 35181 23031 35185
tri 22759 35177 22763 35181 ne
rect 22763 35177 23031 35181
tri 23031 35177 23039 35185 sw
tri 22763 35173 22767 35177 ne
rect 22767 35173 23039 35177
tri 23039 35173 23043 35177 sw
tri 22767 35165 22775 35173 ne
rect 22775 35165 23043 35173
tri 23043 35165 23051 35173 sw
tri 22775 35157 22783 35165 ne
rect 22783 35157 23051 35165
tri 23051 35157 23059 35165 sw
tri 22783 35149 22791 35157 ne
rect 22791 35149 23059 35157
tri 23059 35149 23067 35157 sw
tri 22791 35141 22799 35149 ne
rect 22799 35141 23067 35149
tri 23067 35141 23075 35149 sw
tri 22799 35133 22807 35141 ne
rect 22807 35133 23075 35141
tri 23075 35133 23083 35141 sw
tri 22807 35125 22815 35133 ne
rect 22815 35125 23083 35133
tri 23083 35125 23091 35133 sw
tri 22815 35117 22823 35125 ne
rect 22823 35117 23091 35125
tri 23091 35117 23099 35125 sw
tri 22823 35109 22831 35117 ne
rect 22831 35109 23099 35117
tri 23099 35109 23107 35117 sw
tri 22831 35101 22839 35109 ne
rect 22839 35101 23107 35109
tri 23107 35101 23115 35109 sw
tri 22839 35093 22847 35101 ne
rect 22847 35093 23115 35101
tri 23115 35093 23123 35101 sw
tri 22847 35085 22855 35093 ne
rect 22855 35085 23123 35093
tri 23123 35085 23131 35093 sw
tri 22855 35077 22863 35085 ne
rect 22863 35077 23131 35085
tri 23131 35077 23139 35085 sw
tri 22863 35069 22871 35077 ne
rect 22871 35069 23139 35077
tri 23139 35069 23147 35077 sw
tri 22871 35061 22879 35069 ne
rect 22879 35061 23147 35069
tri 23147 35061 23155 35069 sw
tri 22879 35053 22887 35061 ne
rect 22887 35053 23155 35061
tri 23155 35053 23163 35061 sw
tri 22887 35045 22895 35053 ne
rect 22895 35045 23163 35053
tri 23163 35045 23171 35053 sw
tri 22895 35037 22903 35045 ne
rect 22903 35037 23171 35045
tri 23171 35037 23179 35045 sw
tri 22903 35033 22907 35037 ne
rect 22907 35033 23179 35037
tri 22907 35025 22915 35033 ne
rect 22915 35029 23179 35033
tri 23179 35029 23187 35037 sw
rect 22915 35025 23187 35029
tri 22915 35017 22923 35025 ne
rect 22923 35021 23187 35025
tri 23187 35021 23195 35029 sw
rect 22923 35017 23195 35021
tri 22923 35009 22931 35017 ne
rect 22931 35013 23195 35017
tri 23195 35013 23203 35021 sw
rect 22931 35009 23203 35013
tri 22931 35001 22939 35009 ne
rect 22939 35005 23203 35009
tri 23203 35005 23211 35013 sw
rect 22939 35001 23211 35005
tri 22939 34993 22947 35001 ne
rect 22947 34997 23211 35001
tri 23211 34997 23219 35005 sw
rect 22947 34993 23219 34997
tri 22947 34985 22955 34993 ne
rect 22955 34989 23219 34993
tri 23219 34989 23227 34997 sw
rect 22955 34985 23227 34989
tri 22955 34977 22963 34985 ne
rect 22963 34981 23227 34985
tri 23227 34981 23235 34989 sw
rect 22963 34977 23235 34981
tri 22963 34969 22971 34977 ne
rect 22971 34973 23235 34977
tri 23235 34973 23243 34981 sw
rect 22971 34969 23243 34973
tri 22971 34961 22979 34969 ne
rect 22979 34965 23243 34969
tri 23243 34965 23251 34973 sw
rect 22979 34961 23251 34965
tri 22979 34953 22987 34961 ne
rect 22987 34957 23251 34961
tri 23251 34957 23259 34965 sw
rect 22987 34953 23259 34957
tri 22987 34945 22995 34953 ne
rect 22995 34949 23259 34953
tri 23259 34949 23267 34957 sw
rect 22995 34945 23267 34949
tri 22995 34937 23003 34945 ne
rect 23003 34941 23267 34945
tri 23267 34941 23275 34949 sw
rect 23003 34937 23275 34941
tri 23003 34929 23011 34937 ne
rect 23011 34933 23275 34937
tri 23275 34933 23283 34941 sw
rect 23011 34929 23283 34933
tri 23011 34921 23019 34929 ne
rect 23019 34925 23283 34929
tri 23283 34925 23291 34933 sw
rect 23019 34921 23291 34925
tri 23019 34913 23027 34921 ne
rect 23027 34917 23291 34921
tri 23291 34917 23299 34925 sw
rect 23027 34913 23299 34917
tri 23027 34905 23035 34913 ne
rect 23035 34909 23299 34913
tri 23299 34909 23307 34917 sw
rect 23035 34905 23307 34909
tri 23035 34901 23039 34905 ne
rect 23039 34901 23307 34905
tri 23307 34901 23315 34909 sw
tri 23039 34897 23043 34901 ne
rect 23043 34897 23315 34901
tri 23315 34897 23319 34901 sw
tri 23043 34889 23051 34897 ne
rect 23051 34889 23319 34897
tri 23319 34889 23327 34897 sw
tri 23051 34881 23059 34889 ne
rect 23059 34881 23327 34889
tri 23327 34881 23335 34889 sw
tri 23059 34873 23067 34881 ne
rect 23067 34873 23335 34881
tri 23335 34873 23343 34881 sw
tri 23067 34865 23075 34873 ne
rect 23075 34865 23343 34873
tri 23343 34865 23351 34873 sw
tri 23075 34857 23083 34865 ne
rect 23083 34857 23351 34865
tri 23351 34857 23359 34865 sw
tri 23083 34849 23091 34857 ne
rect 23091 34849 23359 34857
tri 23359 34849 23367 34857 sw
tri 23091 34841 23099 34849 ne
rect 23099 34841 23367 34849
tri 23367 34841 23375 34849 sw
tri 23099 34833 23107 34841 ne
rect 23107 34833 23375 34841
tri 23375 34833 23383 34841 sw
tri 23107 34825 23115 34833 ne
rect 23115 34825 23383 34833
tri 23383 34825 23391 34833 sw
tri 23115 34817 23123 34825 ne
rect 23123 34817 23391 34825
tri 23391 34817 23399 34825 sw
tri 23123 34809 23131 34817 ne
rect 23131 34809 23399 34817
tri 23399 34809 23407 34817 sw
tri 23131 34801 23139 34809 ne
rect 23139 34801 23407 34809
tri 23407 34801 23415 34809 sw
tri 23139 34793 23147 34801 ne
rect 23147 34793 23415 34801
tri 23415 34793 23423 34801 sw
tri 23147 34785 23155 34793 ne
rect 23155 34785 23423 34793
tri 23423 34785 23431 34793 sw
tri 23155 34777 23163 34785 ne
rect 23163 34777 23431 34785
tri 23431 34777 23439 34785 sw
tri 23163 34769 23171 34777 ne
rect 23171 34769 23439 34777
tri 23439 34769 23447 34777 sw
tri 23171 34761 23179 34769 ne
rect 23179 34761 23447 34769
tri 23447 34761 23455 34769 sw
tri 23179 34757 23183 34761 ne
rect 23183 34757 23455 34761
tri 23183 34749 23191 34757 ne
rect 23191 34753 23455 34757
tri 23455 34753 23463 34761 sw
rect 23191 34749 23463 34753
tri 23191 34741 23199 34749 ne
rect 23199 34745 23463 34749
tri 23463 34745 23471 34753 sw
rect 23199 34741 23471 34745
tri 23199 34733 23207 34741 ne
rect 23207 34737 23471 34741
tri 23471 34737 23479 34745 sw
rect 23207 34733 23479 34737
tri 23207 34725 23215 34733 ne
rect 23215 34729 23479 34733
tri 23479 34729 23487 34737 sw
rect 23215 34725 23487 34729
tri 23215 34717 23223 34725 ne
rect 23223 34721 23487 34725
tri 23487 34721 23495 34729 sw
rect 23223 34717 23495 34721
tri 23223 34709 23231 34717 ne
rect 23231 34713 23495 34717
tri 23495 34713 23503 34721 sw
rect 23231 34709 23503 34713
tri 23231 34701 23239 34709 ne
rect 23239 34705 23503 34709
tri 23503 34705 23511 34713 sw
rect 23239 34701 23511 34705
tri 23239 34693 23247 34701 ne
rect 23247 34697 23511 34701
tri 23511 34697 23519 34705 sw
rect 23247 34693 23519 34697
tri 23247 34685 23255 34693 ne
rect 23255 34689 23519 34693
tri 23519 34689 23527 34697 sw
rect 23255 34685 23527 34689
tri 23255 34677 23263 34685 ne
rect 23263 34681 23527 34685
tri 23527 34681 23535 34689 sw
rect 23263 34677 23535 34681
tri 23263 34669 23271 34677 ne
rect 23271 34673 23535 34677
tri 23535 34673 23543 34681 sw
rect 23271 34669 23543 34673
tri 23271 34661 23279 34669 ne
rect 23279 34665 23543 34669
tri 23543 34665 23551 34673 sw
rect 23279 34661 23551 34665
tri 23279 34653 23287 34661 ne
rect 23287 34657 23551 34661
tri 23551 34657 23559 34665 sw
rect 23287 34653 23559 34657
tri 23287 34645 23295 34653 ne
rect 23295 34649 23559 34653
tri 23559 34649 23567 34657 sw
rect 23295 34645 23567 34649
tri 23295 34637 23303 34645 ne
rect 23303 34641 23567 34645
tri 23567 34641 23575 34649 sw
rect 23303 34637 23575 34641
tri 23303 34629 23311 34637 ne
rect 23311 34633 23575 34637
tri 23575 34633 23583 34641 sw
rect 23311 34629 23583 34633
tri 23311 34625 23315 34629 ne
rect 23315 34625 23583 34629
tri 23583 34625 23591 34633 sw
tri 23315 34621 23319 34625 ne
rect 23319 34621 23591 34625
tri 23591 34621 23595 34625 sw
tri 23319 34613 23327 34621 ne
rect 23327 34613 23595 34621
tri 23595 34613 23603 34621 sw
tri 23327 34605 23335 34613 ne
rect 23335 34605 23603 34613
tri 23603 34605 23611 34613 sw
tri 23335 34597 23343 34605 ne
rect 23343 34597 23611 34605
tri 23611 34597 23619 34605 sw
tri 23343 34589 23351 34597 ne
rect 23351 34589 23619 34597
tri 23619 34589 23627 34597 sw
tri 23351 34581 23359 34589 ne
rect 23359 34581 23627 34589
tri 23627 34581 23635 34589 sw
tri 23359 34573 23367 34581 ne
rect 23367 34573 23635 34581
tri 23635 34573 23643 34581 sw
tri 23367 34565 23375 34573 ne
rect 23375 34565 23643 34573
tri 23643 34565 23651 34573 sw
tri 23375 34557 23383 34565 ne
rect 23383 34557 23651 34565
tri 23651 34557 23659 34565 sw
tri 23383 34549 23391 34557 ne
rect 23391 34549 23659 34557
tri 23659 34549 23667 34557 sw
tri 23391 34541 23399 34549 ne
rect 23399 34541 23667 34549
tri 23667 34541 23675 34549 sw
tri 23399 34533 23407 34541 ne
rect 23407 34533 23675 34541
tri 23675 34533 23683 34541 sw
tri 23407 34525 23415 34533 ne
rect 23415 34525 23683 34533
tri 23683 34525 23691 34533 sw
tri 23415 34517 23423 34525 ne
rect 23423 34517 23691 34525
tri 23691 34517 23699 34525 sw
tri 23423 34509 23431 34517 ne
rect 23431 34509 23699 34517
tri 23699 34509 23707 34517 sw
tri 23431 34501 23439 34509 ne
rect 23439 34501 23707 34509
tri 23707 34501 23715 34509 sw
tri 23439 34493 23447 34501 ne
rect 23447 34493 23715 34501
tri 23715 34493 23723 34501 sw
tri 23447 34485 23455 34493 ne
rect 23455 34485 23723 34493
tri 23723 34485 23731 34493 sw
tri 23455 34481 23459 34485 ne
rect 23459 34481 23731 34485
tri 23459 34473 23467 34481 ne
rect 23467 34477 23731 34481
tri 23731 34477 23739 34485 sw
rect 23467 34473 23739 34477
tri 23467 34465 23475 34473 ne
rect 23475 34469 23739 34473
tri 23739 34469 23747 34477 sw
rect 23475 34465 23747 34469
tri 23475 34457 23483 34465 ne
rect 23483 34461 23747 34465
tri 23747 34461 23755 34469 sw
rect 23483 34457 23755 34461
tri 23483 34449 23491 34457 ne
rect 23491 34453 23755 34457
tri 23755 34453 23763 34461 sw
rect 23491 34449 23763 34453
tri 23491 34441 23499 34449 ne
rect 23499 34445 23763 34449
tri 23763 34445 23771 34453 sw
rect 23499 34441 23771 34445
tri 23499 34433 23507 34441 ne
rect 23507 34437 23771 34441
tri 23771 34437 23779 34445 sw
rect 23507 34433 23779 34437
tri 23507 34425 23515 34433 ne
rect 23515 34429 23779 34433
tri 23779 34429 23787 34437 sw
rect 23515 34425 23787 34429
tri 23515 34417 23523 34425 ne
rect 23523 34421 23787 34425
tri 23787 34421 23795 34429 sw
rect 23523 34417 23795 34421
tri 23523 34409 23531 34417 ne
rect 23531 34413 23795 34417
tri 23795 34413 23803 34421 sw
rect 23531 34409 23803 34413
tri 23531 34401 23539 34409 ne
rect 23539 34405 23803 34409
tri 23803 34405 23811 34413 sw
rect 23539 34401 23811 34405
tri 23539 34393 23547 34401 ne
rect 23547 34397 23811 34401
tri 23811 34397 23819 34405 sw
rect 23547 34393 23819 34397
tri 23547 34385 23555 34393 ne
rect 23555 34389 23819 34393
tri 23819 34389 23827 34397 sw
rect 23555 34385 23827 34389
tri 23555 34377 23563 34385 ne
rect 23563 34381 23827 34385
tri 23827 34381 23835 34389 sw
rect 23563 34377 23835 34381
tri 23563 34369 23571 34377 ne
rect 23571 34373 23835 34377
tri 23835 34373 23843 34381 sw
rect 23571 34369 23843 34373
tri 23571 34361 23579 34369 ne
rect 23579 34365 23843 34369
tri 23843 34365 23851 34373 sw
rect 23579 34361 23851 34365
tri 23579 34353 23587 34361 ne
rect 23587 34357 23851 34361
tri 23851 34357 23859 34365 sw
rect 23587 34353 23859 34357
tri 23587 34349 23591 34353 ne
rect 23591 34349 23859 34353
tri 23859 34349 23867 34357 sw
tri 23591 34345 23595 34349 ne
rect 23595 34345 23867 34349
tri 23867 34345 23871 34349 sw
tri 23595 34337 23603 34345 ne
rect 23603 34337 23871 34345
tri 23871 34337 23879 34345 sw
tri 23603 34329 23611 34337 ne
rect 23611 34329 23879 34337
tri 23879 34329 23887 34337 sw
tri 23611 34321 23619 34329 ne
rect 23619 34321 23887 34329
tri 23887 34321 23895 34329 sw
tri 23619 34313 23627 34321 ne
rect 23627 34313 23895 34321
tri 23895 34313 23903 34321 sw
tri 23627 34305 23635 34313 ne
rect 23635 34305 23903 34313
tri 23903 34305 23911 34313 sw
tri 23635 34297 23643 34305 ne
rect 23643 34297 23911 34305
tri 23911 34297 23919 34305 sw
tri 23643 34289 23651 34297 ne
rect 23651 34289 23919 34297
tri 23919 34289 23927 34297 sw
tri 23651 34281 23659 34289 ne
rect 23659 34281 23927 34289
tri 23927 34281 23935 34289 sw
tri 23659 34273 23667 34281 ne
rect 23667 34273 23935 34281
tri 23935 34273 23943 34281 sw
tri 23667 34265 23675 34273 ne
rect 23675 34265 23943 34273
tri 23943 34265 23951 34273 sw
tri 23675 34257 23683 34265 ne
rect 23683 34257 23951 34265
tri 23951 34257 23959 34265 sw
tri 23683 34249 23691 34257 ne
rect 23691 34249 23959 34257
tri 23959 34249 23967 34257 sw
tri 23691 34241 23699 34249 ne
rect 23699 34241 23967 34249
tri 23967 34241 23975 34249 sw
tri 23699 34233 23707 34241 ne
rect 23707 34233 23975 34241
tri 23975 34233 23983 34241 sw
tri 23707 34225 23715 34233 ne
rect 23715 34225 23983 34233
tri 23983 34225 23991 34233 sw
tri 23715 34217 23723 34225 ne
rect 23723 34217 23991 34225
tri 23991 34217 23999 34225 sw
tri 23723 34209 23731 34217 ne
rect 23731 34209 23999 34217
tri 23999 34209 24007 34217 sw
tri 23731 34205 23735 34209 ne
rect 23735 34205 24007 34209
tri 23735 34197 23743 34205 ne
rect 23743 34201 24007 34205
tri 24007 34201 24015 34209 sw
rect 23743 34197 24015 34201
tri 23743 34189 23751 34197 ne
rect 23751 34193 24015 34197
tri 24015 34193 24023 34201 sw
rect 23751 34189 24023 34193
tri 23751 34181 23759 34189 ne
rect 23759 34185 24023 34189
tri 24023 34185 24031 34193 sw
rect 23759 34181 24031 34185
tri 23759 34173 23767 34181 ne
rect 23767 34177 24031 34181
tri 24031 34177 24039 34185 sw
rect 23767 34173 24039 34177
tri 23767 34165 23775 34173 ne
rect 23775 34169 24039 34173
tri 24039 34169 24047 34177 sw
rect 23775 34165 24047 34169
tri 23775 34157 23783 34165 ne
rect 23783 34161 24047 34165
tri 24047 34161 24055 34169 sw
rect 23783 34157 24055 34161
tri 23783 34149 23791 34157 ne
rect 23791 34153 24055 34157
tri 24055 34153 24063 34161 sw
rect 23791 34149 24063 34153
tri 23791 34141 23799 34149 ne
rect 23799 34145 24063 34149
tri 24063 34145 24071 34153 sw
rect 23799 34141 24071 34145
tri 23799 34133 23807 34141 ne
rect 23807 34137 24071 34141
tri 24071 34137 24079 34145 sw
rect 23807 34133 24079 34137
tri 23807 34125 23815 34133 ne
rect 23815 34129 24079 34133
tri 24079 34129 24087 34137 sw
rect 23815 34125 24087 34129
tri 23815 34117 23823 34125 ne
rect 23823 34121 24087 34125
tri 24087 34121 24095 34129 sw
rect 23823 34117 24095 34121
tri 23823 34109 23831 34117 ne
rect 23831 34113 24095 34117
tri 24095 34113 24103 34121 sw
rect 23831 34109 24103 34113
tri 23831 34101 23839 34109 ne
rect 23839 34105 24103 34109
tri 24103 34105 24111 34113 sw
rect 23839 34101 24111 34105
tri 23839 34093 23847 34101 ne
rect 23847 34097 24111 34101
tri 24111 34097 24119 34105 sw
rect 23847 34093 24119 34097
tri 23847 34085 23855 34093 ne
rect 23855 34089 24119 34093
tri 24119 34089 24127 34097 sw
rect 23855 34085 24127 34089
tri 23855 34077 23863 34085 ne
rect 23863 34081 24127 34085
tri 24127 34081 24135 34089 sw
rect 23863 34077 24135 34081
tri 23863 34073 23867 34077 ne
rect 23867 34073 24135 34077
tri 24135 34073 24143 34081 sw
tri 23867 34069 23871 34073 ne
rect 23871 34069 24143 34073
tri 24143 34069 24147 34073 sw
tri 23871 34061 23879 34069 ne
rect 23879 34061 24147 34069
tri 24147 34061 24155 34069 sw
tri 23879 34053 23887 34061 ne
rect 23887 34053 24155 34061
tri 24155 34053 24163 34061 sw
tri 23887 34045 23895 34053 ne
rect 23895 34045 24163 34053
tri 24163 34045 24171 34053 sw
tri 23895 34037 23903 34045 ne
rect 23903 34037 24171 34045
tri 24171 34037 24179 34045 sw
tri 23903 34029 23911 34037 ne
rect 23911 34029 24179 34037
tri 24179 34029 24187 34037 sw
tri 23911 34021 23919 34029 ne
rect 23919 34021 24187 34029
tri 24187 34021 24195 34029 sw
tri 23919 34013 23927 34021 ne
rect 23927 34013 24195 34021
tri 24195 34013 24203 34021 sw
tri 23927 34005 23935 34013 ne
rect 23935 34005 24203 34013
tri 24203 34005 24211 34013 sw
tri 23935 33997 23943 34005 ne
rect 23943 33997 24211 34005
tri 24211 33997 24219 34005 sw
tri 23943 33989 23951 33997 ne
rect 23951 33989 24219 33997
tri 24219 33989 24227 33997 sw
tri 23951 33981 23959 33989 ne
rect 23959 33981 24227 33989
tri 24227 33981 24235 33989 sw
tri 23959 33973 23967 33981 ne
rect 23967 33973 24235 33981
tri 24235 33973 24243 33981 sw
tri 23967 33965 23975 33973 ne
rect 23975 33965 24243 33973
tri 24243 33965 24251 33973 sw
tri 23975 33957 23983 33965 ne
rect 23983 33957 24251 33965
tri 24251 33957 24259 33965 sw
tri 23983 33949 23991 33957 ne
rect 23991 33949 24259 33957
tri 24259 33949 24267 33957 sw
tri 23991 33941 23999 33949 ne
rect 23999 33941 24267 33949
tri 24267 33941 24275 33949 sw
tri 23999 33933 24007 33941 ne
rect 24007 33933 24275 33941
tri 24275 33933 24283 33941 sw
tri 24007 33929 24011 33933 ne
rect 24011 33929 24283 33933
tri 24011 33921 24019 33929 ne
rect 24019 33925 24283 33929
tri 24283 33925 24291 33933 sw
rect 24019 33921 24291 33925
tri 24019 33913 24027 33921 ne
rect 24027 33917 24291 33921
tri 24291 33917 24299 33925 sw
rect 24027 33913 24299 33917
tri 24027 33905 24035 33913 ne
rect 24035 33909 24299 33913
tri 24299 33909 24307 33917 sw
rect 24035 33905 24307 33909
tri 24035 33897 24043 33905 ne
rect 24043 33901 24307 33905
tri 24307 33901 24315 33909 sw
rect 24043 33897 24315 33901
tri 24043 33889 24051 33897 ne
rect 24051 33893 24315 33897
tri 24315 33893 24323 33901 sw
rect 24051 33889 24323 33893
tri 24051 33881 24059 33889 ne
rect 24059 33885 24323 33889
tri 24323 33885 24331 33893 sw
rect 24059 33881 24331 33885
tri 24059 33873 24067 33881 ne
rect 24067 33877 24331 33881
tri 24331 33877 24339 33885 sw
rect 24067 33873 24339 33877
tri 24067 33865 24075 33873 ne
rect 24075 33869 24339 33873
tri 24339 33869 24347 33877 sw
rect 24075 33865 24347 33869
tri 24075 33857 24083 33865 ne
rect 24083 33861 24347 33865
tri 24347 33861 24355 33869 sw
rect 24083 33857 24355 33861
tri 24083 33849 24091 33857 ne
rect 24091 33853 24355 33857
tri 24355 33853 24363 33861 sw
rect 24091 33849 24363 33853
tri 24091 33841 24099 33849 ne
rect 24099 33845 24363 33849
tri 24363 33845 24371 33853 sw
rect 24099 33841 24371 33845
tri 24099 33833 24107 33841 ne
rect 24107 33837 24371 33841
tri 24371 33837 24379 33845 sw
rect 24107 33833 24379 33837
tri 24107 33825 24115 33833 ne
rect 24115 33829 24379 33833
tri 24379 33829 24387 33837 sw
rect 24115 33825 24387 33829
tri 24115 33817 24123 33825 ne
rect 24123 33821 24387 33825
tri 24387 33821 24395 33829 sw
rect 24123 33817 24395 33821
tri 24123 33809 24131 33817 ne
rect 24131 33813 24395 33817
tri 24395 33813 24403 33821 sw
rect 24131 33809 24403 33813
tri 24131 33801 24139 33809 ne
rect 24139 33805 24403 33809
tri 24403 33805 24411 33813 sw
rect 24139 33801 24411 33805
tri 24139 33797 24143 33801 ne
rect 24143 33797 24411 33801
tri 24411 33797 24419 33805 sw
tri 24143 33793 24147 33797 ne
rect 24147 33793 24419 33797
tri 24419 33793 24423 33797 sw
tri 24147 33785 24155 33793 ne
rect 24155 33785 24423 33793
tri 24423 33785 24431 33793 sw
tri 24155 33777 24163 33785 ne
rect 24163 33777 24431 33785
tri 24431 33777 24439 33785 sw
tri 24163 33769 24171 33777 ne
rect 24171 33769 24439 33777
tri 24439 33769 24447 33777 sw
tri 24171 33761 24179 33769 ne
rect 24179 33761 24447 33769
tri 24447 33761 24455 33769 sw
tri 24179 33753 24187 33761 ne
rect 24187 33753 24455 33761
tri 24455 33753 24463 33761 sw
tri 24187 33745 24195 33753 ne
rect 24195 33745 24463 33753
tri 24463 33745 24471 33753 sw
tri 24195 33737 24203 33745 ne
rect 24203 33737 24471 33745
tri 24471 33737 24479 33745 sw
tri 24203 33729 24211 33737 ne
rect 24211 33729 24479 33737
tri 24479 33729 24487 33737 sw
tri 24211 33721 24219 33729 ne
rect 24219 33721 24487 33729
tri 24487 33721 24495 33729 sw
tri 24219 33713 24227 33721 ne
rect 24227 33713 24495 33721
tri 24495 33713 24503 33721 sw
tri 24227 33705 24235 33713 ne
rect 24235 33705 24503 33713
tri 24503 33705 24511 33713 sw
tri 24235 33697 24243 33705 ne
rect 24243 33697 24511 33705
tri 24511 33697 24519 33705 sw
tri 24243 33689 24251 33697 ne
rect 24251 33689 24519 33697
tri 24519 33689 24527 33697 sw
tri 24251 33681 24259 33689 ne
rect 24259 33681 24527 33689
tri 24527 33681 24535 33689 sw
tri 24259 33673 24267 33681 ne
rect 24267 33673 24535 33681
tri 24535 33673 24543 33681 sw
tri 24267 33665 24275 33673 ne
rect 24275 33665 24543 33673
tri 24543 33665 24551 33673 sw
tri 24275 33657 24283 33665 ne
rect 24283 33657 24551 33665
tri 24551 33657 24559 33665 sw
tri 24283 33653 24287 33657 ne
rect 24287 33653 24559 33657
tri 24287 33645 24295 33653 ne
rect 24295 33649 24559 33653
tri 24559 33649 24567 33657 sw
rect 24295 33645 24567 33649
tri 24295 33637 24303 33645 ne
rect 24303 33641 24567 33645
tri 24567 33641 24575 33649 sw
rect 24303 33637 24575 33641
tri 24303 33629 24311 33637 ne
rect 24311 33633 24575 33637
tri 24575 33633 24583 33641 sw
rect 24311 33629 24583 33633
tri 24311 33621 24319 33629 ne
rect 24319 33625 24583 33629
tri 24583 33625 24591 33633 sw
rect 24319 33621 24591 33625
tri 24319 33613 24327 33621 ne
rect 24327 33617 24591 33621
tri 24591 33617 24599 33625 sw
rect 24327 33613 24599 33617
tri 24327 33605 24335 33613 ne
rect 24335 33609 24599 33613
tri 24599 33609 24607 33617 sw
rect 24335 33605 24607 33609
tri 24335 33597 24343 33605 ne
rect 24343 33601 24607 33605
tri 24607 33601 24615 33609 sw
rect 24343 33597 24615 33601
tri 24343 33589 24351 33597 ne
rect 24351 33593 24615 33597
tri 24615 33593 24623 33601 sw
rect 24351 33589 24623 33593
tri 24351 33581 24359 33589 ne
rect 24359 33585 24623 33589
tri 24623 33585 24631 33593 sw
rect 24359 33581 24631 33585
tri 24359 33573 24367 33581 ne
rect 24367 33577 24631 33581
tri 24631 33577 24639 33585 sw
rect 24367 33573 24639 33577
tri 24367 33565 24375 33573 ne
rect 24375 33569 24639 33573
tri 24639 33569 24647 33577 sw
rect 24375 33565 24647 33569
tri 24375 33557 24383 33565 ne
rect 24383 33561 24647 33565
tri 24647 33561 24655 33569 sw
rect 24383 33557 24655 33561
tri 24383 33549 24391 33557 ne
rect 24391 33553 24655 33557
tri 24655 33553 24663 33561 sw
rect 24391 33549 24663 33553
tri 24391 33541 24399 33549 ne
rect 24399 33545 24663 33549
tri 24663 33545 24671 33553 sw
rect 24399 33541 24671 33545
tri 24399 33533 24407 33541 ne
rect 24407 33537 24671 33541
tri 24671 33537 24679 33545 sw
rect 24407 33533 24679 33537
tri 24407 33525 24415 33533 ne
rect 24415 33529 24679 33533
tri 24679 33529 24687 33537 sw
rect 24415 33525 24687 33529
tri 24415 33521 24419 33525 ne
rect 24419 33521 24687 33525
tri 24687 33521 24695 33529 sw
tri 24419 33517 24423 33521 ne
rect 24423 33517 24695 33521
tri 24695 33517 24699 33521 sw
tri 24423 33509 24431 33517 ne
rect 24431 33509 24699 33517
tri 24699 33509 24707 33517 sw
tri 24431 33501 24439 33509 ne
rect 24439 33501 24707 33509
tri 24707 33501 24715 33509 sw
tri 24439 33493 24447 33501 ne
rect 24447 33493 24715 33501
tri 24715 33493 24723 33501 sw
tri 24447 33485 24455 33493 ne
rect 24455 33485 24723 33493
tri 24723 33485 24731 33493 sw
tri 24455 33477 24463 33485 ne
rect 24463 33477 24731 33485
tri 24731 33477 24739 33485 sw
tri 24463 33469 24471 33477 ne
rect 24471 33469 24739 33477
tri 24739 33469 24747 33477 sw
tri 24471 33461 24479 33469 ne
rect 24479 33461 24747 33469
tri 24747 33461 24755 33469 sw
tri 24479 33453 24487 33461 ne
rect 24487 33453 24755 33461
tri 24755 33453 24763 33461 sw
tri 24487 33445 24495 33453 ne
rect 24495 33445 24763 33453
tri 24763 33445 24771 33453 sw
tri 24495 33437 24503 33445 ne
rect 24503 33437 24771 33445
tri 24771 33437 24779 33445 sw
tri 24503 33429 24511 33437 ne
rect 24511 33429 24779 33437
tri 24779 33429 24787 33437 sw
tri 24511 33421 24519 33429 ne
rect 24519 33421 24787 33429
tri 24787 33421 24795 33429 sw
tri 24519 33413 24527 33421 ne
rect 24527 33413 24795 33421
tri 24795 33413 24803 33421 sw
tri 24527 33405 24535 33413 ne
rect 24535 33405 24803 33413
tri 24803 33405 24811 33413 sw
tri 24535 33397 24543 33405 ne
rect 24543 33397 24811 33405
tri 24811 33397 24819 33405 sw
tri 24543 33389 24551 33397 ne
rect 24551 33389 24819 33397
tri 24819 33389 24827 33397 sw
tri 24551 33381 24559 33389 ne
rect 24559 33381 24827 33389
tri 24827 33381 24835 33389 sw
tri 24559 33377 24563 33381 ne
rect 24563 33377 24835 33381
tri 24563 33369 24571 33377 ne
rect 24571 33373 24835 33377
tri 24835 33373 24843 33381 sw
rect 24571 33369 24843 33373
tri 24571 33361 24579 33369 ne
rect 24579 33365 24843 33369
tri 24843 33365 24851 33373 sw
rect 24579 33361 24851 33365
tri 24579 33353 24587 33361 ne
rect 24587 33357 24851 33361
tri 24851 33357 24859 33365 sw
rect 24587 33353 24859 33357
tri 24587 33345 24595 33353 ne
rect 24595 33349 24859 33353
tri 24859 33349 24867 33357 sw
rect 24595 33345 24867 33349
tri 24595 33337 24603 33345 ne
rect 24603 33341 24867 33345
tri 24867 33341 24875 33349 sw
rect 24603 33337 24875 33341
tri 24603 33329 24611 33337 ne
rect 24611 33333 24875 33337
tri 24875 33333 24883 33341 sw
rect 24611 33329 24883 33333
tri 24611 33321 24619 33329 ne
rect 24619 33325 24883 33329
tri 24883 33325 24891 33333 sw
rect 24619 33321 24891 33325
tri 24619 33313 24627 33321 ne
rect 24627 33317 24891 33321
tri 24891 33317 24899 33325 sw
rect 24627 33313 24899 33317
tri 24627 33305 24635 33313 ne
rect 24635 33309 24899 33313
tri 24899 33309 24907 33317 sw
rect 24635 33305 24907 33309
tri 24635 33297 24643 33305 ne
rect 24643 33301 24907 33305
tri 24907 33301 24915 33309 sw
rect 24643 33297 24915 33301
tri 24643 33289 24651 33297 ne
rect 24651 33293 24915 33297
tri 24915 33293 24923 33301 sw
rect 24651 33289 24923 33293
tri 24651 33281 24659 33289 ne
rect 24659 33285 24923 33289
tri 24923 33285 24931 33293 sw
rect 24659 33281 24931 33285
tri 24659 33273 24667 33281 ne
rect 24667 33277 24931 33281
tri 24931 33277 24939 33285 sw
rect 24667 33273 24939 33277
tri 24667 33265 24675 33273 ne
rect 24675 33269 24939 33273
tri 24939 33269 24947 33277 sw
rect 24675 33265 24947 33269
tri 24675 33257 24683 33265 ne
rect 24683 33261 24947 33265
tri 24947 33261 24955 33269 sw
rect 24683 33257 24955 33261
tri 24683 33249 24691 33257 ne
rect 24691 33253 24955 33257
tri 24955 33253 24963 33261 sw
rect 24691 33249 24963 33253
tri 24691 33245 24695 33249 ne
rect 24695 33245 24963 33249
tri 24963 33245 24971 33253 sw
tri 24695 33241 24699 33245 ne
rect 24699 33241 24971 33245
tri 24971 33241 24975 33245 sw
tri 24699 33233 24707 33241 ne
rect 24707 33233 24975 33241
tri 24975 33233 24983 33241 sw
tri 24707 33225 24715 33233 ne
rect 24715 33225 24983 33233
tri 24983 33225 24991 33233 sw
tri 24715 33217 24723 33225 ne
rect 24723 33217 24991 33225
tri 24991 33217 24999 33225 sw
tri 24723 33209 24731 33217 ne
rect 24731 33209 24999 33217
tri 24999 33209 25007 33217 sw
tri 24731 33201 24739 33209 ne
rect 24739 33201 25007 33209
tri 25007 33201 25015 33209 sw
tri 24739 33193 24747 33201 ne
rect 24747 33193 25015 33201
tri 25015 33193 25023 33201 sw
tri 24747 33185 24755 33193 ne
rect 24755 33185 25023 33193
tri 25023 33185 25031 33193 sw
tri 24755 33177 24763 33185 ne
rect 24763 33177 25031 33185
tri 25031 33177 25039 33185 sw
tri 24763 33169 24771 33177 ne
rect 24771 33169 25039 33177
tri 25039 33169 25047 33177 sw
tri 24771 33161 24779 33169 ne
rect 24779 33161 25047 33169
tri 25047 33161 25055 33169 sw
tri 24779 33153 24787 33161 ne
rect 24787 33153 25055 33161
tri 25055 33153 25063 33161 sw
tri 24787 33145 24795 33153 ne
rect 24795 33145 25063 33153
tri 25063 33145 25071 33153 sw
tri 24795 33137 24803 33145 ne
rect 24803 33137 25071 33145
tri 25071 33137 25079 33145 sw
tri 24803 33129 24811 33137 ne
rect 24811 33129 25079 33137
tri 25079 33129 25087 33137 sw
tri 24811 33121 24819 33129 ne
rect 24819 33121 25087 33129
tri 25087 33121 25095 33129 sw
tri 24819 33113 24827 33121 ne
rect 24827 33113 25095 33121
tri 25095 33113 25103 33121 sw
tri 24827 33105 24835 33113 ne
rect 24835 33105 25103 33113
tri 25103 33105 25111 33113 sw
tri 24835 33101 24839 33105 ne
rect 24839 33101 25111 33105
tri 24839 33093 24847 33101 ne
rect 24847 33097 25111 33101
tri 25111 33097 25119 33105 sw
rect 24847 33093 25119 33097
tri 24847 33085 24855 33093 ne
rect 24855 33089 25119 33093
tri 25119 33089 25127 33097 sw
rect 24855 33085 25127 33089
tri 24855 33077 24863 33085 ne
rect 24863 33081 25127 33085
tri 25127 33081 25135 33089 sw
rect 24863 33077 25135 33081
tri 24863 33069 24871 33077 ne
rect 24871 33073 25135 33077
tri 25135 33073 25143 33081 sw
rect 24871 33069 25143 33073
tri 24871 33061 24879 33069 ne
rect 24879 33065 25143 33069
tri 25143 33065 25151 33073 sw
rect 24879 33061 25151 33065
tri 24879 33053 24887 33061 ne
rect 24887 33057 25151 33061
tri 25151 33057 25159 33065 sw
rect 24887 33053 25159 33057
tri 24887 33045 24895 33053 ne
rect 24895 33049 25159 33053
tri 25159 33049 25167 33057 sw
rect 24895 33045 25167 33049
tri 24895 33037 24903 33045 ne
rect 24903 33041 25167 33045
tri 25167 33041 25175 33049 sw
rect 24903 33037 25175 33041
tri 24903 33029 24911 33037 ne
rect 24911 33033 25175 33037
tri 25175 33033 25183 33041 sw
rect 24911 33029 25183 33033
tri 24911 33021 24919 33029 ne
rect 24919 33025 25183 33029
tri 25183 33025 25191 33033 sw
rect 24919 33021 25191 33025
tri 24919 33013 24927 33021 ne
rect 24927 33017 25191 33021
tri 25191 33017 25199 33025 sw
rect 24927 33013 25199 33017
tri 24927 33005 24935 33013 ne
rect 24935 33009 25199 33013
tri 25199 33009 25207 33017 sw
rect 24935 33005 25207 33009
tri 24935 32997 24943 33005 ne
rect 24943 33001 25207 33005
tri 25207 33001 25215 33009 sw
rect 24943 32997 25215 33001
tri 24943 32989 24951 32997 ne
rect 24951 32993 25215 32997
tri 25215 32993 25223 33001 sw
rect 24951 32989 25223 32993
tri 24951 32981 24959 32989 ne
rect 24959 32985 25223 32989
tri 25223 32985 25231 32993 sw
rect 24959 32981 25231 32985
tri 24959 32973 24967 32981 ne
rect 24967 32977 25231 32981
tri 25231 32977 25239 32985 sw
rect 24967 32973 25239 32977
tri 24967 32969 24971 32973 ne
rect 24971 32969 25239 32973
tri 25239 32969 25247 32977 sw
tri 24971 32965 24975 32969 ne
rect 24975 32965 25247 32969
tri 25247 32965 25251 32969 sw
tri 24975 32957 24983 32965 ne
rect 24983 32957 25251 32965
tri 25251 32957 25259 32965 sw
tri 24983 32949 24991 32957 ne
rect 24991 32949 25259 32957
tri 25259 32949 25267 32957 sw
tri 24991 32941 24999 32949 ne
rect 24999 32941 25267 32949
tri 25267 32941 25275 32949 sw
tri 24999 32933 25007 32941 ne
rect 25007 32933 25275 32941
tri 25275 32933 25283 32941 sw
tri 25007 32925 25015 32933 ne
rect 25015 32925 25283 32933
tri 25283 32925 25291 32933 sw
tri 25015 32917 25023 32925 ne
rect 25023 32917 25291 32925
tri 25291 32917 25299 32925 sw
tri 25023 32909 25031 32917 ne
rect 25031 32909 25299 32917
tri 25299 32909 25307 32917 sw
tri 25031 32901 25039 32909 ne
rect 25039 32901 25307 32909
tri 25307 32901 25315 32909 sw
tri 25039 32893 25047 32901 ne
rect 25047 32893 25315 32901
tri 25315 32893 25323 32901 sw
tri 25047 32885 25055 32893 ne
rect 25055 32885 25323 32893
tri 25323 32885 25331 32893 sw
tri 25055 32877 25063 32885 ne
rect 25063 32877 25331 32885
tri 25331 32877 25339 32885 sw
tri 25063 32869 25071 32877 ne
rect 25071 32869 25339 32877
tri 25339 32869 25347 32877 sw
tri 25071 32861 25079 32869 ne
rect 25079 32861 25347 32869
tri 25347 32861 25355 32869 sw
tri 25079 32853 25087 32861 ne
rect 25087 32853 25355 32861
tri 25355 32853 25363 32861 sw
tri 25087 32845 25095 32853 ne
rect 25095 32845 25363 32853
tri 25363 32845 25371 32853 sw
tri 25095 32837 25103 32845 ne
rect 25103 32837 25371 32845
tri 25371 32837 25379 32845 sw
tri 25103 32829 25111 32837 ne
rect 25111 32829 25379 32837
tri 25379 32829 25387 32837 sw
tri 25111 32825 25115 32829 ne
rect 25115 32825 25387 32829
tri 25115 32817 25123 32825 ne
rect 25123 32821 25387 32825
tri 25387 32821 25395 32829 sw
rect 25123 32817 25395 32821
tri 25123 32809 25131 32817 ne
rect 25131 32813 25395 32817
tri 25395 32813 25403 32821 sw
rect 25131 32809 25403 32813
tri 25131 32801 25139 32809 ne
rect 25139 32805 25403 32809
tri 25403 32805 25411 32813 sw
rect 25139 32801 25411 32805
tri 25139 32793 25147 32801 ne
rect 25147 32797 25411 32801
tri 25411 32797 25419 32805 sw
rect 25147 32793 25419 32797
tri 25147 32785 25155 32793 ne
rect 25155 32789 25419 32793
tri 25419 32789 25427 32797 sw
rect 25155 32785 25427 32789
tri 25155 32777 25163 32785 ne
rect 25163 32781 25427 32785
tri 25427 32781 25435 32789 sw
rect 25163 32777 25435 32781
tri 25163 32769 25171 32777 ne
rect 25171 32773 25435 32777
tri 25435 32773 25443 32781 sw
rect 25171 32769 25443 32773
tri 25171 32761 25179 32769 ne
rect 25179 32765 25443 32769
tri 25443 32765 25451 32773 sw
rect 25179 32761 25451 32765
tri 25179 32753 25187 32761 ne
rect 25187 32757 25451 32761
tri 25451 32757 25459 32765 sw
rect 25187 32753 25459 32757
tri 25187 32745 25195 32753 ne
rect 25195 32749 25459 32753
tri 25459 32749 25467 32757 sw
rect 25195 32745 25467 32749
tri 25195 32737 25203 32745 ne
rect 25203 32741 25467 32745
tri 25467 32741 25475 32749 sw
rect 25203 32737 25475 32741
tri 25203 32729 25211 32737 ne
rect 25211 32733 25475 32737
tri 25475 32733 25483 32741 sw
rect 25211 32729 25483 32733
tri 25211 32721 25219 32729 ne
rect 25219 32725 25483 32729
tri 25483 32725 25491 32733 sw
rect 25219 32721 25491 32725
tri 25219 32713 25227 32721 ne
rect 25227 32717 25491 32721
tri 25491 32717 25499 32725 sw
rect 25227 32713 25499 32717
tri 25227 32705 25235 32713 ne
rect 25235 32709 25499 32713
tri 25499 32709 25507 32717 sw
rect 25235 32705 25507 32709
tri 25235 32697 25243 32705 ne
rect 25243 32701 25507 32705
tri 25507 32701 25515 32709 sw
rect 25243 32697 25515 32701
tri 25243 32693 25247 32697 ne
rect 25247 32693 25515 32697
tri 25515 32693 25523 32701 sw
tri 25247 32689 25251 32693 ne
rect 25251 32689 25523 32693
tri 25523 32689 25527 32693 sw
tri 25251 32681 25259 32689 ne
rect 25259 32681 25527 32689
tri 25527 32681 25535 32689 sw
tri 25259 32673 25267 32681 ne
rect 25267 32673 25535 32681
tri 25535 32673 25543 32681 sw
tri 25267 32665 25275 32673 ne
rect 25275 32665 25543 32673
tri 25543 32665 25551 32673 sw
tri 25275 32657 25283 32665 ne
rect 25283 32657 25551 32665
tri 25551 32657 25559 32665 sw
tri 25283 32649 25291 32657 ne
rect 25291 32649 25559 32657
tri 25559 32649 25567 32657 sw
tri 25291 32641 25299 32649 ne
rect 25299 32641 25567 32649
tri 25567 32641 25575 32649 sw
tri 25299 32633 25307 32641 ne
rect 25307 32633 25575 32641
tri 25575 32633 25583 32641 sw
tri 25307 32625 25315 32633 ne
rect 25315 32625 25583 32633
tri 25583 32625 25591 32633 sw
tri 25315 32617 25323 32625 ne
rect 25323 32617 25591 32625
tri 25591 32617 25599 32625 sw
tri 25323 32609 25331 32617 ne
rect 25331 32609 25599 32617
tri 25599 32609 25607 32617 sw
tri 25331 32601 25339 32609 ne
rect 25339 32601 25607 32609
tri 25607 32601 25615 32609 sw
tri 25339 32593 25347 32601 ne
rect 25347 32593 25615 32601
tri 25615 32593 25623 32601 sw
tri 25347 32585 25355 32593 ne
rect 25355 32585 25623 32593
tri 25623 32585 25631 32593 sw
tri 25355 32577 25363 32585 ne
rect 25363 32577 25631 32585
tri 25631 32577 25639 32585 sw
tri 25363 32569 25371 32577 ne
rect 25371 32569 25639 32577
tri 25639 32569 25647 32577 sw
tri 25371 32561 25379 32569 ne
rect 25379 32561 25647 32569
tri 25647 32561 25655 32569 sw
tri 25379 32553 25387 32561 ne
rect 25387 32553 25655 32561
tri 25655 32553 25663 32561 sw
tri 25387 32549 25391 32553 ne
rect 25391 32549 25663 32553
tri 25391 32541 25399 32549 ne
rect 25399 32545 25663 32549
tri 25663 32545 25671 32553 sw
rect 25399 32541 25671 32545
tri 25399 32533 25407 32541 ne
rect 25407 32537 25671 32541
tri 25671 32537 25679 32545 sw
rect 25407 32533 25679 32537
tri 25407 32525 25415 32533 ne
rect 25415 32529 25679 32533
tri 25679 32529 25687 32537 sw
rect 25415 32525 25687 32529
tri 25415 32517 25423 32525 ne
rect 25423 32521 25687 32525
tri 25687 32521 25695 32529 sw
rect 25423 32517 25695 32521
tri 25423 32509 25431 32517 ne
rect 25431 32513 25695 32517
tri 25695 32513 25703 32521 sw
rect 25431 32509 25703 32513
tri 25431 32501 25439 32509 ne
rect 25439 32505 25703 32509
tri 25703 32505 25711 32513 sw
rect 25439 32501 25711 32505
tri 25439 32493 25447 32501 ne
rect 25447 32497 25711 32501
tri 25711 32497 25719 32505 sw
rect 25447 32493 25719 32497
tri 25447 32485 25455 32493 ne
rect 25455 32489 25719 32493
tri 25719 32489 25727 32497 sw
rect 25455 32485 25727 32489
tri 25455 32477 25463 32485 ne
rect 25463 32481 25727 32485
tri 25727 32481 25735 32489 sw
rect 25463 32477 25735 32481
tri 25463 32469 25471 32477 ne
rect 25471 32473 25735 32477
tri 25735 32473 25743 32481 sw
rect 25471 32469 25743 32473
tri 25471 32461 25479 32469 ne
rect 25479 32465 25743 32469
tri 25743 32465 25751 32473 sw
rect 25479 32461 25751 32465
tri 25479 32453 25487 32461 ne
rect 25487 32457 25751 32461
tri 25751 32457 25759 32465 sw
rect 25487 32453 25759 32457
tri 25487 32445 25495 32453 ne
rect 25495 32449 25759 32453
tri 25759 32449 25767 32457 sw
rect 25495 32445 25767 32449
tri 25495 32437 25503 32445 ne
rect 25503 32441 25767 32445
tri 25767 32441 25775 32449 sw
rect 25503 32437 25775 32441
tri 25503 32429 25511 32437 ne
rect 25511 32433 25775 32437
tri 25775 32433 25783 32441 sw
rect 25511 32429 25783 32433
tri 25511 32421 25519 32429 ne
rect 25519 32425 25783 32429
tri 25783 32425 25791 32433 sw
rect 25519 32421 25791 32425
tri 25519 32417 25523 32421 ne
rect 25523 32417 25791 32421
tri 25791 32417 25799 32425 sw
tri 25523 32413 25527 32417 ne
rect 25527 32413 25799 32417
tri 25799 32413 25803 32417 sw
tri 25527 32405 25535 32413 ne
rect 25535 32405 25803 32413
tri 25803 32405 25811 32413 sw
tri 25535 32397 25543 32405 ne
rect 25543 32397 25811 32405
tri 25811 32397 25819 32405 sw
tri 25543 32389 25551 32397 ne
rect 25551 32389 25819 32397
tri 25819 32389 25827 32397 sw
tri 25551 32381 25559 32389 ne
rect 25559 32381 25827 32389
tri 25827 32381 25835 32389 sw
tri 25559 32373 25567 32381 ne
rect 25567 32373 25835 32381
tri 25835 32373 25843 32381 sw
tri 25567 32365 25575 32373 ne
rect 25575 32365 25843 32373
tri 25843 32365 25851 32373 sw
tri 25575 32357 25583 32365 ne
rect 25583 32357 25851 32365
tri 25851 32357 25859 32365 sw
tri 25583 32349 25591 32357 ne
rect 25591 32349 25859 32357
tri 25859 32349 25867 32357 sw
tri 25591 32341 25599 32349 ne
rect 25599 32341 25867 32349
tri 25867 32341 25875 32349 sw
tri 25599 32333 25607 32341 ne
rect 25607 32333 25875 32341
tri 25875 32333 25883 32341 sw
tri 25607 32325 25615 32333 ne
rect 25615 32325 25883 32333
tri 25883 32325 25891 32333 sw
tri 25615 32317 25623 32325 ne
rect 25623 32317 25891 32325
tri 25891 32317 25899 32325 sw
tri 25623 32309 25631 32317 ne
rect 25631 32309 25899 32317
tri 25899 32309 25907 32317 sw
tri 25631 32301 25639 32309 ne
rect 25639 32301 25907 32309
tri 25907 32301 25915 32309 sw
tri 25639 32293 25647 32301 ne
rect 25647 32293 25915 32301
tri 25915 32293 25923 32301 sw
tri 25647 32285 25655 32293 ne
rect 25655 32285 25923 32293
tri 25923 32285 25931 32293 sw
tri 25655 32277 25663 32285 ne
rect 25663 32277 25931 32285
tri 25931 32277 25939 32285 sw
tri 25663 32273 25667 32277 ne
rect 25667 32273 25939 32277
tri 25667 32265 25675 32273 ne
rect 25675 32269 25939 32273
tri 25939 32269 25947 32277 sw
rect 25675 32265 25947 32269
tri 25675 32257 25683 32265 ne
rect 25683 32261 25947 32265
tri 25947 32261 25955 32269 sw
rect 25683 32257 25955 32261
tri 25683 32249 25691 32257 ne
rect 25691 32253 25955 32257
tri 25955 32253 25963 32261 sw
rect 25691 32249 25963 32253
tri 25691 32241 25699 32249 ne
rect 25699 32245 25963 32249
tri 25963 32245 25971 32253 sw
rect 25699 32241 25971 32245
tri 25699 32233 25707 32241 ne
rect 25707 32237 25971 32241
tri 25971 32237 25979 32245 sw
rect 25707 32233 25979 32237
tri 25707 32225 25715 32233 ne
rect 25715 32229 25979 32233
tri 25979 32229 25987 32237 sw
rect 25715 32225 25987 32229
tri 25715 32217 25723 32225 ne
rect 25723 32221 25987 32225
tri 25987 32221 25995 32229 sw
rect 25723 32217 25995 32221
tri 25723 32209 25731 32217 ne
rect 25731 32213 25995 32217
tri 25995 32213 26003 32221 sw
rect 25731 32209 26003 32213
tri 25731 32201 25739 32209 ne
rect 25739 32205 26003 32209
tri 26003 32205 26011 32213 sw
rect 25739 32201 26011 32205
tri 25739 32193 25747 32201 ne
rect 25747 32197 26011 32201
tri 26011 32197 26019 32205 sw
rect 25747 32193 26019 32197
tri 25747 32185 25755 32193 ne
rect 25755 32189 26019 32193
tri 26019 32189 26027 32197 sw
rect 25755 32185 26027 32189
tri 25755 32177 25763 32185 ne
rect 25763 32181 26027 32185
tri 26027 32181 26035 32189 sw
rect 25763 32177 26035 32181
tri 25763 32169 25771 32177 ne
rect 25771 32173 26035 32177
tri 26035 32173 26043 32181 sw
rect 25771 32169 26043 32173
tri 25771 32161 25779 32169 ne
rect 25779 32165 26043 32169
tri 26043 32165 26051 32173 sw
rect 25779 32161 26051 32165
tri 25779 32153 25787 32161 ne
rect 25787 32157 26051 32161
tri 26051 32157 26059 32165 sw
rect 25787 32153 26059 32157
tri 25787 32145 25795 32153 ne
rect 25795 32149 26059 32153
tri 26059 32149 26067 32157 sw
rect 25795 32145 26067 32149
tri 25795 32141 25799 32145 ne
rect 25799 32141 26067 32145
tri 26067 32141 26075 32149 sw
tri 25799 32137 25803 32141 ne
rect 25803 32137 26075 32141
tri 26075 32137 26079 32141 sw
tri 25803 32129 25811 32137 ne
rect 25811 32129 26079 32137
tri 26079 32129 26087 32137 sw
tri 25811 32121 25819 32129 ne
rect 25819 32121 26087 32129
tri 26087 32121 26095 32129 sw
tri 25819 32113 25827 32121 ne
rect 25827 32113 26095 32121
tri 26095 32113 26103 32121 sw
tri 25827 32105 25835 32113 ne
rect 25835 32105 26103 32113
tri 26103 32105 26111 32113 sw
tri 25835 32097 25843 32105 ne
rect 25843 32097 26111 32105
tri 26111 32097 26119 32105 sw
tri 25843 32089 25851 32097 ne
rect 25851 32089 26119 32097
tri 26119 32089 26127 32097 sw
tri 25851 32081 25859 32089 ne
rect 25859 32081 26127 32089
tri 26127 32081 26135 32089 sw
tri 25859 32073 25867 32081 ne
rect 25867 32073 26135 32081
tri 26135 32073 26143 32081 sw
tri 25867 32065 25875 32073 ne
rect 25875 32065 26143 32073
tri 26143 32065 26151 32073 sw
tri 25875 32057 25883 32065 ne
rect 25883 32057 26151 32065
tri 26151 32057 26159 32065 sw
tri 25883 32049 25891 32057 ne
rect 25891 32049 26159 32057
tri 26159 32049 26167 32057 sw
tri 25891 32041 25899 32049 ne
rect 25899 32041 26167 32049
tri 26167 32041 26175 32049 sw
tri 25899 32033 25907 32041 ne
rect 25907 32033 26175 32041
tri 26175 32033 26183 32041 sw
tri 25907 32025 25915 32033 ne
rect 25915 32025 26183 32033
tri 26183 32025 26191 32033 sw
tri 25915 32017 25923 32025 ne
rect 25923 32017 26191 32025
tri 26191 32017 26199 32025 sw
tri 25923 32009 25931 32017 ne
rect 25931 32009 26199 32017
tri 26199 32009 26207 32017 sw
tri 25931 32001 25939 32009 ne
rect 25939 32001 26207 32009
tri 26207 32001 26215 32009 sw
tri 25939 31997 25943 32001 ne
rect 25943 31997 26215 32001
tri 25943 31989 25951 31997 ne
rect 25951 31993 26215 31997
tri 26215 31993 26223 32001 sw
rect 25951 31989 26223 31993
tri 25951 31981 25959 31989 ne
rect 25959 31985 26223 31989
tri 26223 31985 26231 31993 sw
rect 25959 31981 26231 31985
tri 25959 31973 25967 31981 ne
rect 25967 31977 26231 31981
tri 26231 31977 26239 31985 sw
rect 25967 31973 26239 31977
tri 25967 31965 25975 31973 ne
rect 25975 31969 26239 31973
tri 26239 31969 26247 31977 sw
rect 25975 31965 26247 31969
tri 25975 31957 25983 31965 ne
rect 25983 31961 26247 31965
tri 26247 31961 26255 31969 sw
rect 25983 31957 26255 31961
tri 25983 31949 25991 31957 ne
rect 25991 31953 26255 31957
tri 26255 31953 26263 31961 sw
rect 25991 31949 26263 31953
tri 25991 31941 25999 31949 ne
rect 25999 31945 26263 31949
tri 26263 31945 26271 31953 sw
rect 25999 31941 26271 31945
tri 25999 31933 26007 31941 ne
rect 26007 31937 26271 31941
tri 26271 31937 26279 31945 sw
rect 26007 31933 26279 31937
tri 26007 31925 26015 31933 ne
rect 26015 31929 26279 31933
tri 26279 31929 26287 31937 sw
rect 26015 31925 26287 31929
tri 26015 31917 26023 31925 ne
rect 26023 31921 26287 31925
tri 26287 31921 26295 31929 sw
rect 26023 31917 26295 31921
tri 26023 31909 26031 31917 ne
rect 26031 31913 26295 31917
tri 26295 31913 26303 31921 sw
rect 26031 31909 26303 31913
tri 26031 31901 26039 31909 ne
rect 26039 31905 26303 31909
tri 26303 31905 26311 31913 sw
rect 26039 31901 26311 31905
tri 26039 31893 26047 31901 ne
rect 26047 31897 26311 31901
tri 26311 31897 26319 31905 sw
rect 26047 31893 26319 31897
tri 26047 31885 26055 31893 ne
rect 26055 31889 26319 31893
tri 26319 31889 26327 31897 sw
rect 26055 31885 26327 31889
tri 26055 31877 26063 31885 ne
rect 26063 31881 26327 31885
tri 26327 31881 26335 31889 sw
rect 26063 31877 26335 31881
tri 26063 31869 26071 31877 ne
rect 26071 31873 26335 31877
tri 26335 31873 26343 31881 sw
rect 26071 31869 26343 31873
tri 26071 31865 26075 31869 ne
rect 26075 31865 26343 31869
tri 26343 31865 26351 31873 sw
tri 26075 31861 26079 31865 ne
rect 26079 31861 26351 31865
tri 26351 31861 26355 31865 sw
tri 26079 31853 26087 31861 ne
rect 26087 31853 26355 31861
tri 26355 31853 26363 31861 sw
tri 26087 31845 26095 31853 ne
rect 26095 31845 26363 31853
tri 26363 31845 26371 31853 sw
tri 26095 31837 26103 31845 ne
rect 26103 31837 26371 31845
tri 26371 31837 26379 31845 sw
tri 26103 31829 26111 31837 ne
rect 26111 31829 26379 31837
tri 26379 31829 26387 31837 sw
tri 26111 31821 26119 31829 ne
rect 26119 31821 26387 31829
tri 26387 31821 26395 31829 sw
tri 26119 31813 26127 31821 ne
rect 26127 31813 26395 31821
tri 26395 31813 26403 31821 sw
tri 26127 31805 26135 31813 ne
rect 26135 31805 26403 31813
tri 26403 31805 26411 31813 sw
tri 26135 31797 26143 31805 ne
rect 26143 31797 26411 31805
tri 26411 31797 26419 31805 sw
tri 26143 31789 26151 31797 ne
rect 26151 31789 26419 31797
tri 26419 31789 26427 31797 sw
tri 26151 31781 26159 31789 ne
rect 26159 31781 26427 31789
tri 26427 31781 26435 31789 sw
tri 26159 31773 26167 31781 ne
rect 26167 31773 26435 31781
tri 26435 31773 26443 31781 sw
tri 26167 31765 26175 31773 ne
rect 26175 31765 26443 31773
tri 26443 31765 26451 31773 sw
tri 26175 31757 26183 31765 ne
rect 26183 31757 26451 31765
tri 26451 31757 26459 31765 sw
tri 26183 31749 26191 31757 ne
rect 26191 31749 26459 31757
tri 26459 31749 26467 31757 sw
tri 26191 31741 26199 31749 ne
rect 26199 31741 26467 31749
tri 26467 31741 26475 31749 sw
tri 26199 31733 26207 31741 ne
rect 26207 31733 26475 31741
tri 26475 31733 26483 31741 sw
tri 26207 31725 26215 31733 ne
rect 26215 31725 26483 31733
tri 26483 31725 26491 31733 sw
tri 26215 31721 26219 31725 ne
rect 26219 31721 26491 31725
tri 26219 31713 26227 31721 ne
rect 26227 31717 26491 31721
tri 26491 31717 26499 31725 sw
rect 26227 31713 26499 31717
tri 26227 31705 26235 31713 ne
rect 26235 31709 26499 31713
tri 26499 31709 26507 31717 sw
rect 26235 31705 26507 31709
tri 26235 31697 26243 31705 ne
rect 26243 31701 26507 31705
tri 26507 31701 26515 31709 sw
rect 26243 31697 26515 31701
tri 26243 31689 26251 31697 ne
rect 26251 31693 26515 31697
tri 26515 31693 26523 31701 sw
rect 26251 31689 26523 31693
tri 26251 31681 26259 31689 ne
rect 26259 31685 26523 31689
tri 26523 31685 26531 31693 sw
rect 26259 31681 26531 31685
tri 26259 31673 26267 31681 ne
rect 26267 31677 26531 31681
tri 26531 31677 26539 31685 sw
rect 26267 31673 26539 31677
tri 26267 31665 26275 31673 ne
rect 26275 31669 26539 31673
tri 26539 31669 26547 31677 sw
rect 26275 31665 26547 31669
tri 26275 31657 26283 31665 ne
rect 26283 31661 26547 31665
tri 26547 31661 26555 31669 sw
rect 26283 31657 26555 31661
tri 26283 31649 26291 31657 ne
rect 26291 31653 26555 31657
tri 26555 31653 26563 31661 sw
rect 26291 31649 26563 31653
tri 26291 31641 26299 31649 ne
rect 26299 31645 26563 31649
tri 26563 31645 26571 31653 sw
rect 26299 31641 26571 31645
tri 26299 31633 26307 31641 ne
rect 26307 31637 26571 31641
tri 26571 31637 26579 31645 sw
rect 26307 31633 26579 31637
tri 26307 31625 26315 31633 ne
rect 26315 31629 26579 31633
tri 26579 31629 26587 31637 sw
rect 26315 31625 26587 31629
tri 26315 31617 26323 31625 ne
rect 26323 31621 26587 31625
tri 26587 31621 26595 31629 sw
rect 26323 31617 26595 31621
tri 26323 31609 26331 31617 ne
rect 26331 31613 26595 31617
tri 26595 31613 26603 31621 sw
rect 26331 31609 26603 31613
tri 26331 31601 26339 31609 ne
rect 26339 31605 26603 31609
tri 26603 31605 26611 31613 sw
rect 26339 31601 26611 31605
tri 26339 31593 26347 31601 ne
rect 26347 31597 26611 31601
tri 26611 31597 26619 31605 sw
rect 26347 31593 26619 31597
tri 26347 31589 26351 31593 ne
rect 26351 31589 26619 31593
tri 26619 31589 26627 31597 sw
tri 26351 31585 26355 31589 ne
rect 26355 31585 26627 31589
tri 26627 31585 26631 31589 sw
tri 26355 31577 26363 31585 ne
rect 26363 31577 26631 31585
tri 26631 31577 26639 31585 sw
tri 26363 31569 26371 31577 ne
rect 26371 31569 26639 31577
tri 26639 31569 26647 31577 sw
tri 26371 31561 26379 31569 ne
rect 26379 31561 26647 31569
tri 26647 31561 26655 31569 sw
tri 26379 31553 26387 31561 ne
rect 26387 31553 26655 31561
tri 26655 31553 26663 31561 sw
tri 26387 31545 26395 31553 ne
rect 26395 31545 26663 31553
tri 26663 31545 26671 31553 sw
tri 26395 31537 26403 31545 ne
rect 26403 31537 26671 31545
tri 26671 31537 26679 31545 sw
tri 26403 31529 26411 31537 ne
rect 26411 31529 26679 31537
tri 26679 31529 26687 31537 sw
tri 26411 31521 26419 31529 ne
rect 26419 31521 26687 31529
tri 26687 31521 26695 31529 sw
tri 26419 31513 26427 31521 ne
rect 26427 31513 26695 31521
tri 26695 31513 26703 31521 sw
tri 26427 31505 26435 31513 ne
rect 26435 31505 26703 31513
tri 26703 31505 26711 31513 sw
tri 26435 31497 26443 31505 ne
rect 26443 31497 26711 31505
tri 26711 31497 26719 31505 sw
tri 26443 31489 26451 31497 ne
rect 26451 31489 26719 31497
tri 26719 31489 26727 31497 sw
tri 26451 31481 26459 31489 ne
rect 26459 31481 26727 31489
tri 26727 31481 26735 31489 sw
tri 26459 31473 26467 31481 ne
rect 26467 31473 26735 31481
tri 26735 31473 26743 31481 sw
tri 26467 31465 26475 31473 ne
rect 26475 31465 26743 31473
tri 26743 31465 26751 31473 sw
tri 26475 31457 26483 31465 ne
rect 26483 31457 26751 31465
tri 26751 31457 26759 31465 sw
tri 26483 31449 26491 31457 ne
rect 26491 31449 26759 31457
tri 26759 31449 26767 31457 sw
tri 26491 31445 26495 31449 ne
rect 26495 31445 26767 31449
tri 26495 31437 26503 31445 ne
rect 26503 31441 26767 31445
tri 26767 31441 26775 31449 sw
rect 26503 31437 26775 31441
tri 26503 31429 26511 31437 ne
rect 26511 31433 26775 31437
tri 26775 31433 26783 31441 sw
rect 26511 31429 26783 31433
tri 26511 31421 26519 31429 ne
rect 26519 31425 26783 31429
tri 26783 31425 26791 31433 sw
rect 26519 31421 26791 31425
tri 26519 31413 26527 31421 ne
rect 26527 31417 26791 31421
tri 26791 31417 26799 31425 sw
rect 26527 31413 26799 31417
tri 26527 31405 26535 31413 ne
rect 26535 31409 26799 31413
tri 26799 31409 26807 31417 sw
rect 26535 31405 26807 31409
tri 26535 31397 26543 31405 ne
rect 26543 31401 26807 31405
tri 26807 31401 26815 31409 sw
rect 26543 31397 26815 31401
tri 26543 31389 26551 31397 ne
rect 26551 31393 26815 31397
tri 26815 31393 26823 31401 sw
rect 26551 31389 26823 31393
tri 26551 31381 26559 31389 ne
rect 26559 31385 26823 31389
tri 26823 31385 26831 31393 sw
rect 26559 31381 26831 31385
tri 26559 31373 26567 31381 ne
rect 26567 31377 26831 31381
tri 26831 31377 26839 31385 sw
rect 26567 31373 26839 31377
tri 26567 31365 26575 31373 ne
rect 26575 31369 26839 31373
tri 26839 31369 26847 31377 sw
rect 26575 31365 26847 31369
tri 26575 31357 26583 31365 ne
rect 26583 31361 26847 31365
tri 26847 31361 26855 31369 sw
rect 26583 31357 26855 31361
tri 26583 31349 26591 31357 ne
rect 26591 31353 26855 31357
tri 26855 31353 26863 31361 sw
rect 26591 31349 26863 31353
tri 26591 31341 26599 31349 ne
rect 26599 31345 26863 31349
tri 26863 31345 26871 31353 sw
rect 26599 31341 26871 31345
tri 26599 31333 26607 31341 ne
rect 26607 31337 26871 31341
tri 26871 31337 26879 31345 sw
rect 26607 31333 26879 31337
tri 26607 31325 26615 31333 ne
rect 26615 31329 26879 31333
tri 26879 31329 26887 31337 sw
rect 26615 31325 26887 31329
tri 26615 31317 26623 31325 ne
rect 26623 31321 26887 31325
tri 26887 31321 26895 31329 sw
rect 26623 31317 26895 31321
tri 26623 31313 26627 31317 ne
rect 26627 31313 26895 31317
tri 26895 31313 26903 31321 sw
tri 26627 31309 26631 31313 ne
rect 26631 31309 26903 31313
tri 26903 31309 26907 31313 sw
tri 26631 31301 26639 31309 ne
rect 26639 31301 26907 31309
tri 26907 31301 26915 31309 sw
tri 26639 31293 26647 31301 ne
rect 26647 31293 26915 31301
tri 26915 31293 26923 31301 sw
tri 26647 31285 26655 31293 ne
rect 26655 31285 26923 31293
tri 26923 31285 26931 31293 sw
tri 26655 31277 26663 31285 ne
rect 26663 31277 26931 31285
tri 26931 31277 26939 31285 sw
tri 26663 31269 26671 31277 ne
rect 26671 31269 26939 31277
tri 26939 31269 26947 31277 sw
tri 26671 31261 26679 31269 ne
rect 26679 31261 26947 31269
tri 26947 31261 26955 31269 sw
tri 26679 31253 26687 31261 ne
rect 26687 31253 26955 31261
tri 26955 31253 26963 31261 sw
tri 26687 31245 26695 31253 ne
rect 26695 31245 26963 31253
tri 26963 31245 26971 31253 sw
tri 26695 31237 26703 31245 ne
rect 26703 31237 26971 31245
tri 26971 31237 26979 31245 sw
tri 26703 31229 26711 31237 ne
rect 26711 31229 26979 31237
tri 26979 31229 26987 31237 sw
tri 26711 31221 26719 31229 ne
rect 26719 31221 26987 31229
tri 26987 31221 26995 31229 sw
tri 26719 31213 26727 31221 ne
rect 26727 31213 26995 31221
tri 26995 31213 27003 31221 sw
tri 26727 31205 26735 31213 ne
rect 26735 31205 27003 31213
tri 27003 31205 27011 31213 sw
tri 26735 31197 26743 31205 ne
rect 26743 31197 27011 31205
tri 27011 31197 27019 31205 sw
tri 26743 31189 26751 31197 ne
rect 26751 31189 27019 31197
tri 27019 31189 27027 31197 sw
tri 26751 31181 26759 31189 ne
rect 26759 31181 27027 31189
tri 27027 31181 27035 31189 sw
tri 26759 31173 26767 31181 ne
rect 26767 31173 27035 31181
tri 27035 31173 27043 31181 sw
tri 26767 31169 26771 31173 ne
rect 26771 31169 27043 31173
tri 26771 31161 26779 31169 ne
rect 26779 31165 27043 31169
tri 27043 31165 27051 31173 sw
rect 26779 31161 27051 31165
tri 26779 31153 26787 31161 ne
rect 26787 31157 27051 31161
tri 27051 31157 27059 31165 sw
rect 26787 31153 27059 31157
tri 26787 31145 26795 31153 ne
rect 26795 31149 27059 31153
tri 27059 31149 27067 31157 sw
rect 26795 31145 27067 31149
tri 26795 31137 26803 31145 ne
rect 26803 31141 27067 31145
tri 27067 31141 27075 31149 sw
rect 26803 31137 27075 31141
tri 26803 31129 26811 31137 ne
rect 26811 31133 27075 31137
tri 27075 31133 27083 31141 sw
rect 26811 31129 27083 31133
tri 26811 31121 26819 31129 ne
rect 26819 31125 27083 31129
tri 27083 31125 27091 31133 sw
rect 26819 31121 27091 31125
tri 26819 31113 26827 31121 ne
rect 26827 31117 27091 31121
tri 27091 31117 27099 31125 sw
rect 26827 31113 27099 31117
tri 26827 31105 26835 31113 ne
rect 26835 31109 27099 31113
tri 27099 31109 27107 31117 sw
rect 26835 31105 27107 31109
tri 26835 31097 26843 31105 ne
rect 26843 31101 27107 31105
tri 27107 31101 27115 31109 sw
rect 26843 31097 27115 31101
tri 26843 31089 26851 31097 ne
rect 26851 31093 27115 31097
tri 27115 31093 27123 31101 sw
rect 26851 31089 27123 31093
tri 26851 31081 26859 31089 ne
rect 26859 31085 27123 31089
tri 27123 31085 27131 31093 sw
rect 26859 31081 27131 31085
tri 26859 31073 26867 31081 ne
rect 26867 31077 27131 31081
tri 27131 31077 27139 31085 sw
rect 26867 31073 27139 31077
tri 26867 31065 26875 31073 ne
rect 26875 31069 27139 31073
tri 27139 31069 27147 31077 sw
rect 26875 31065 27147 31069
tri 26875 31057 26883 31065 ne
rect 26883 31061 27147 31065
tri 27147 31061 27155 31069 sw
rect 26883 31057 27155 31061
tri 26883 31049 26891 31057 ne
rect 26891 31053 27155 31057
tri 27155 31053 27163 31061 sw
rect 26891 31049 27163 31053
tri 26891 31041 26899 31049 ne
rect 26899 31045 27163 31049
tri 27163 31045 27171 31053 sw
rect 26899 31041 27171 31045
tri 26899 31037 26903 31041 ne
rect 26903 31037 27171 31041
tri 27171 31037 27179 31045 sw
tri 26903 31033 26907 31037 ne
rect 26907 31033 27179 31037
tri 27179 31033 27183 31037 sw
tri 26907 31025 26915 31033 ne
rect 26915 31025 27183 31033
tri 27183 31025 27191 31033 sw
tri 26915 31017 26923 31025 ne
rect 26923 31017 27191 31025
tri 27191 31017 27199 31025 sw
tri 26923 31009 26931 31017 ne
rect 26931 31009 27199 31017
tri 27199 31009 27207 31017 sw
tri 26931 31001 26939 31009 ne
rect 26939 31001 27207 31009
tri 27207 31001 27215 31009 sw
tri 26939 30993 26947 31001 ne
rect 26947 30993 27215 31001
tri 27215 30993 27223 31001 sw
tri 26947 30985 26955 30993 ne
rect 26955 30985 27223 30993
tri 27223 30985 27231 30993 sw
tri 26955 30977 26963 30985 ne
rect 26963 30977 27231 30985
tri 27231 30977 27239 30985 sw
tri 26963 30969 26971 30977 ne
rect 26971 30969 27239 30977
tri 27239 30969 27247 30977 sw
tri 26971 30961 26979 30969 ne
rect 26979 30961 27247 30969
tri 27247 30961 27255 30969 sw
tri 26979 30953 26987 30961 ne
rect 26987 30953 27255 30961
tri 27255 30953 27263 30961 sw
tri 26987 30945 26995 30953 ne
rect 26995 30945 27263 30953
tri 27263 30945 27271 30953 sw
tri 26995 30937 27003 30945 ne
rect 27003 30937 27271 30945
tri 27271 30937 27279 30945 sw
tri 27003 30929 27011 30937 ne
rect 27011 30929 27279 30937
tri 27279 30929 27287 30937 sw
tri 27011 30921 27019 30929 ne
rect 27019 30921 27287 30929
tri 27287 30921 27295 30929 sw
tri 27019 30913 27027 30921 ne
rect 27027 30913 27295 30921
tri 27295 30913 27303 30921 sw
tri 27027 30905 27035 30913 ne
rect 27035 30905 27303 30913
tri 27303 30905 27311 30913 sw
tri 27035 30897 27043 30905 ne
rect 27043 30897 27311 30905
tri 27311 30897 27319 30905 sw
tri 27043 30893 27047 30897 ne
rect 27047 30893 27319 30897
tri 27047 30885 27055 30893 ne
rect 27055 30889 27319 30893
tri 27319 30889 27327 30897 sw
rect 27055 30885 27327 30889
tri 27055 30877 27063 30885 ne
rect 27063 30881 27327 30885
tri 27327 30881 27335 30889 sw
rect 27063 30877 27335 30881
tri 27063 30869 27071 30877 ne
rect 27071 30873 27335 30877
tri 27335 30873 27343 30881 sw
rect 27071 30869 27343 30873
tri 27071 30861 27079 30869 ne
rect 27079 30865 27343 30869
tri 27343 30865 27351 30873 sw
rect 27079 30861 27351 30865
tri 27079 30853 27087 30861 ne
rect 27087 30857 27351 30861
tri 27351 30857 27359 30865 sw
rect 27087 30853 27359 30857
tri 27087 30845 27095 30853 ne
rect 27095 30849 27359 30853
tri 27359 30849 27367 30857 sw
rect 27095 30845 27367 30849
tri 27095 30837 27103 30845 ne
rect 27103 30841 27367 30845
tri 27367 30841 27375 30849 sw
rect 27103 30837 27375 30841
tri 27103 30829 27111 30837 ne
rect 27111 30833 27375 30837
tri 27375 30833 27383 30841 sw
rect 27111 30829 27383 30833
tri 27111 30821 27119 30829 ne
rect 27119 30825 27383 30829
tri 27383 30825 27391 30833 sw
rect 27119 30821 27391 30825
tri 27119 30813 27127 30821 ne
rect 27127 30817 27391 30821
tri 27391 30817 27399 30825 sw
rect 27127 30813 27399 30817
tri 27127 30805 27135 30813 ne
rect 27135 30809 27399 30813
tri 27399 30809 27407 30817 sw
rect 27135 30805 27407 30809
tri 27135 30797 27143 30805 ne
rect 27143 30801 27407 30805
tri 27407 30801 27415 30809 sw
rect 27143 30797 27415 30801
tri 27143 30789 27151 30797 ne
rect 27151 30793 27415 30797
tri 27415 30793 27423 30801 sw
rect 27151 30789 27423 30793
tri 27151 30781 27159 30789 ne
rect 27159 30785 27423 30789
tri 27423 30785 27431 30793 sw
rect 27159 30781 27431 30785
tri 27159 30773 27167 30781 ne
rect 27167 30777 27431 30781
tri 27431 30777 27439 30785 sw
rect 27167 30773 27439 30777
tri 27167 30765 27175 30773 ne
rect 27175 30769 27439 30773
tri 27439 30769 27447 30777 sw
rect 27175 30765 27447 30769
tri 27175 30761 27179 30765 ne
rect 27179 30761 27447 30765
tri 27447 30761 27455 30769 sw
tri 27179 30757 27183 30761 ne
rect 27183 30757 27455 30761
tri 27455 30757 27459 30761 sw
tri 27183 30749 27191 30757 ne
rect 27191 30749 27459 30757
tri 27459 30749 27467 30757 sw
tri 27191 30741 27199 30749 ne
rect 27199 30741 27467 30749
tri 27467 30741 27475 30749 sw
tri 27199 30733 27207 30741 ne
rect 27207 30733 27475 30741
tri 27475 30733 27483 30741 sw
tri 27207 30725 27215 30733 ne
rect 27215 30725 27483 30733
tri 27483 30725 27491 30733 sw
tri 27215 30717 27223 30725 ne
rect 27223 30717 27491 30725
tri 27491 30717 27499 30725 sw
tri 27223 30709 27231 30717 ne
rect 27231 30709 27499 30717
tri 27499 30709 27507 30717 sw
tri 27231 30701 27239 30709 ne
rect 27239 30701 27507 30709
tri 27507 30701 27515 30709 sw
tri 27239 30693 27247 30701 ne
rect 27247 30693 27515 30701
tri 27515 30693 27523 30701 sw
tri 27247 30685 27255 30693 ne
rect 27255 30685 27523 30693
tri 27523 30685 27531 30693 sw
tri 27255 30677 27263 30685 ne
rect 27263 30677 27531 30685
tri 27531 30677 27539 30685 sw
tri 27263 30669 27271 30677 ne
rect 27271 30669 27539 30677
tri 27539 30669 27547 30677 sw
tri 27271 30661 27279 30669 ne
rect 27279 30661 27547 30669
tri 27547 30661 27555 30669 sw
tri 27279 30653 27287 30661 ne
rect 27287 30653 27555 30661
tri 27555 30653 27563 30661 sw
tri 27287 30645 27295 30653 ne
rect 27295 30645 27563 30653
tri 27563 30645 27571 30653 sw
tri 27295 30637 27303 30645 ne
rect 27303 30637 27571 30645
tri 27571 30637 27579 30645 sw
tri 27303 30629 27311 30637 ne
rect 27311 30629 27579 30637
tri 27579 30629 27587 30637 sw
tri 27311 30621 27319 30629 ne
rect 27319 30621 27587 30629
tri 27587 30621 27595 30629 sw
tri 27319 30617 27323 30621 ne
rect 27323 30617 27595 30621
tri 27323 30609 27331 30617 ne
rect 27331 30613 27595 30617
tri 27595 30613 27603 30621 sw
rect 27331 30609 27603 30613
tri 27331 30601 27339 30609 ne
rect 27339 30605 27603 30609
tri 27603 30605 27611 30613 sw
rect 27339 30601 27611 30605
tri 27339 30593 27347 30601 ne
rect 27347 30597 27611 30601
tri 27611 30597 27619 30605 sw
rect 27347 30593 27619 30597
tri 27347 30585 27355 30593 ne
rect 27355 30589 27619 30593
tri 27619 30589 27627 30597 sw
rect 27355 30585 27627 30589
tri 27355 30577 27363 30585 ne
rect 27363 30581 27627 30585
tri 27627 30581 27635 30589 sw
rect 27363 30577 27635 30581
tri 27363 30569 27371 30577 ne
rect 27371 30573 27635 30577
tri 27635 30573 27643 30581 sw
rect 27371 30569 27643 30573
tri 27371 30561 27379 30569 ne
rect 27379 30565 27643 30569
tri 27643 30565 27651 30573 sw
rect 27379 30561 27651 30565
tri 27379 30553 27387 30561 ne
rect 27387 30557 27651 30561
tri 27651 30557 27659 30565 sw
rect 27387 30553 27659 30557
tri 27387 30545 27395 30553 ne
rect 27395 30549 27659 30553
tri 27659 30549 27667 30557 sw
rect 27395 30545 27667 30549
tri 27395 30537 27403 30545 ne
rect 27403 30541 27667 30545
tri 27667 30541 27675 30549 sw
rect 27403 30537 27675 30541
tri 27403 30529 27411 30537 ne
rect 27411 30533 27675 30537
tri 27675 30533 27683 30541 sw
rect 27411 30529 27683 30533
tri 27411 30521 27419 30529 ne
rect 27419 30525 27683 30529
tri 27683 30525 27691 30533 sw
rect 27419 30521 27691 30525
tri 27419 30513 27427 30521 ne
rect 27427 30517 27691 30521
tri 27691 30517 27699 30525 sw
rect 27427 30513 27699 30517
tri 27427 30505 27435 30513 ne
rect 27435 30509 27699 30513
tri 27699 30509 27707 30517 sw
rect 27435 30505 27707 30509
tri 27435 30497 27443 30505 ne
rect 27443 30501 27707 30505
tri 27707 30501 27715 30509 sw
rect 27443 30497 27715 30501
tri 27443 30489 27451 30497 ne
rect 27451 30493 27715 30497
tri 27715 30493 27723 30501 sw
rect 27451 30489 27723 30493
tri 27451 30485 27455 30489 ne
rect 27455 30485 27723 30489
tri 27723 30485 27731 30493 sw
tri 27455 30481 27459 30485 ne
rect 27459 30481 27731 30485
tri 27731 30481 27735 30485 sw
tri 27459 30473 27467 30481 ne
rect 27467 30473 27735 30481
tri 27735 30473 27743 30481 sw
tri 27467 30465 27475 30473 ne
rect 27475 30465 27743 30473
tri 27743 30465 27751 30473 sw
tri 27475 30457 27483 30465 ne
rect 27483 30457 27751 30465
tri 27751 30457 27759 30465 sw
tri 27483 30449 27491 30457 ne
rect 27491 30449 27759 30457
tri 27759 30449 27767 30457 sw
tri 27491 30441 27499 30449 ne
rect 27499 30441 27767 30449
tri 27767 30441 27775 30449 sw
tri 27499 30433 27507 30441 ne
rect 27507 30433 27775 30441
tri 27775 30433 27783 30441 sw
tri 27507 30425 27515 30433 ne
rect 27515 30425 27783 30433
tri 27783 30425 27791 30433 sw
tri 27515 30417 27523 30425 ne
rect 27523 30417 27791 30425
tri 27791 30417 27799 30425 sw
tri 27523 30409 27531 30417 ne
rect 27531 30409 27799 30417
tri 27799 30409 27807 30417 sw
tri 27531 30401 27539 30409 ne
rect 27539 30401 27807 30409
tri 27807 30401 27815 30409 sw
tri 27539 30393 27547 30401 ne
rect 27547 30393 27815 30401
tri 27815 30393 27823 30401 sw
tri 27547 30385 27555 30393 ne
rect 27555 30385 27823 30393
tri 27823 30385 27831 30393 sw
tri 27555 30377 27563 30385 ne
rect 27563 30377 27831 30385
tri 27831 30377 27839 30385 sw
tri 27563 30369 27571 30377 ne
rect 27571 30369 27839 30377
tri 27839 30369 27847 30377 sw
tri 27571 30361 27579 30369 ne
rect 27579 30361 27847 30369
tri 27847 30361 27855 30369 sw
tri 27579 30353 27587 30361 ne
rect 27587 30353 27855 30361
tri 27855 30353 27863 30361 sw
tri 27587 30345 27595 30353 ne
rect 27595 30345 27863 30353
tri 27863 30345 27871 30353 sw
tri 27595 30341 27599 30345 ne
rect 27599 30341 27871 30345
tri 27599 30333 27607 30341 ne
rect 27607 30337 27871 30341
tri 27871 30337 27879 30345 sw
rect 27607 30333 27879 30337
tri 27607 30325 27615 30333 ne
rect 27615 30329 27879 30333
tri 27879 30329 27887 30337 sw
rect 27615 30325 27887 30329
tri 27615 30317 27623 30325 ne
rect 27623 30321 27887 30325
tri 27887 30321 27895 30329 sw
rect 27623 30317 27895 30321
tri 27623 30309 27631 30317 ne
rect 27631 30313 27895 30317
tri 27895 30313 27903 30321 sw
rect 27631 30309 27903 30313
tri 27631 30301 27639 30309 ne
rect 27639 30305 27903 30309
tri 27903 30305 27911 30313 sw
rect 27639 30301 27911 30305
tri 27639 30293 27647 30301 ne
rect 27647 30297 27911 30301
tri 27911 30297 27919 30305 sw
rect 27647 30293 27919 30297
tri 27647 30285 27655 30293 ne
rect 27655 30289 27919 30293
tri 27919 30289 27927 30297 sw
rect 27655 30285 27927 30289
tri 27655 30277 27663 30285 ne
rect 27663 30281 27927 30285
tri 27927 30281 27935 30289 sw
rect 27663 30277 27935 30281
tri 27663 30269 27671 30277 ne
rect 27671 30273 27935 30277
tri 27935 30273 27943 30281 sw
rect 27671 30269 27943 30273
tri 27671 30261 27679 30269 ne
rect 27679 30265 27943 30269
tri 27943 30265 27951 30273 sw
rect 27679 30261 27951 30265
tri 27679 30253 27687 30261 ne
rect 27687 30257 27951 30261
tri 27951 30257 27959 30265 sw
rect 27687 30253 27959 30257
tri 27687 30245 27695 30253 ne
rect 27695 30249 27959 30253
tri 27959 30249 27967 30257 sw
rect 27695 30245 27967 30249
tri 27695 30237 27703 30245 ne
rect 27703 30241 27967 30245
tri 27967 30241 27975 30249 sw
rect 27703 30237 27975 30241
tri 27703 30229 27711 30237 ne
rect 27711 30233 27975 30237
tri 27975 30233 27983 30241 sw
rect 27711 30229 27983 30233
tri 27711 30221 27719 30229 ne
rect 27719 30225 27983 30229
tri 27983 30225 27991 30233 sw
rect 27719 30221 27991 30225
tri 27719 30213 27727 30221 ne
rect 27727 30217 27991 30221
tri 27991 30217 27999 30225 sw
rect 27727 30213 27999 30217
tri 27727 30209 27731 30213 ne
rect 27731 30209 27999 30213
tri 27999 30209 28007 30217 sw
tri 27731 30205 27735 30209 ne
rect 27735 30205 28007 30209
tri 28007 30205 28011 30209 sw
tri 27735 30197 27743 30205 ne
rect 27743 30197 28011 30205
tri 28011 30197 28019 30205 sw
tri 27743 30189 27751 30197 ne
rect 27751 30189 28019 30197
tri 28019 30189 28027 30197 sw
tri 27751 30181 27759 30189 ne
rect 27759 30181 28027 30189
tri 28027 30181 28035 30189 sw
tri 27759 30173 27767 30181 ne
rect 27767 30173 28035 30181
tri 28035 30173 28043 30181 sw
tri 27767 30165 27775 30173 ne
rect 27775 30165 28043 30173
tri 28043 30165 28051 30173 sw
tri 27775 30157 27783 30165 ne
rect 27783 30157 28051 30165
tri 28051 30157 28059 30165 sw
tri 27783 30149 27791 30157 ne
rect 27791 30149 28059 30157
tri 28059 30149 28067 30157 sw
tri 27791 30141 27799 30149 ne
rect 27799 30141 28067 30149
tri 28067 30141 28075 30149 sw
tri 27799 30133 27807 30141 ne
rect 27807 30133 28075 30141
tri 28075 30133 28083 30141 sw
tri 27807 30125 27815 30133 ne
rect 27815 30125 28083 30133
tri 28083 30125 28091 30133 sw
tri 27815 30117 27823 30125 ne
rect 27823 30117 28091 30125
tri 28091 30117 28099 30125 sw
tri 27823 30109 27831 30117 ne
rect 27831 30109 28099 30117
tri 28099 30109 28107 30117 sw
tri 27831 30101 27839 30109 ne
rect 27839 30101 28107 30109
tri 28107 30101 28115 30109 sw
tri 27839 30093 27847 30101 ne
rect 27847 30093 28115 30101
tri 28115 30093 28123 30101 sw
tri 27847 30085 27855 30093 ne
rect 27855 30085 28123 30093
tri 28123 30085 28131 30093 sw
tri 27855 30077 27863 30085 ne
rect 27863 30077 28131 30085
tri 28131 30077 28139 30085 sw
tri 27863 30069 27871 30077 ne
rect 27871 30069 28139 30077
tri 28139 30069 28147 30077 sw
tri 27871 30065 27875 30069 ne
rect 27875 30065 28147 30069
tri 27875 30057 27883 30065 ne
rect 27883 30061 28147 30065
tri 28147 30061 28155 30069 sw
rect 27883 30057 28155 30061
tri 27883 30049 27891 30057 ne
rect 27891 30053 28155 30057
tri 28155 30053 28163 30061 sw
rect 27891 30049 28163 30053
tri 27891 30041 27899 30049 ne
rect 27899 30045 28163 30049
tri 28163 30045 28171 30053 sw
rect 27899 30041 28171 30045
tri 27899 30033 27907 30041 ne
rect 27907 30037 28171 30041
tri 28171 30037 28179 30045 sw
rect 27907 30033 28179 30037
tri 27907 30025 27915 30033 ne
rect 27915 30029 28179 30033
tri 28179 30029 28187 30037 sw
rect 27915 30025 28187 30029
tri 27915 30017 27923 30025 ne
rect 27923 30021 28187 30025
tri 28187 30021 28195 30029 sw
rect 27923 30017 28195 30021
tri 27923 30009 27931 30017 ne
rect 27931 30013 28195 30017
tri 28195 30013 28203 30021 sw
rect 27931 30009 28203 30013
tri 27931 30001 27939 30009 ne
rect 27939 30005 28203 30009
tri 28203 30005 28211 30013 sw
rect 27939 30001 28211 30005
tri 27939 29993 27947 30001 ne
rect 27947 29997 28211 30001
tri 28211 29997 28219 30005 sw
rect 27947 29993 28219 29997
tri 27947 29985 27955 29993 ne
rect 27955 29989 28219 29993
tri 28219 29989 28227 29997 sw
rect 27955 29985 28227 29989
tri 27955 29977 27963 29985 ne
rect 27963 29981 28227 29985
tri 28227 29981 28235 29989 sw
rect 27963 29977 28235 29981
tri 27963 29969 27971 29977 ne
rect 27971 29973 28235 29977
tri 28235 29973 28243 29981 sw
rect 27971 29969 28243 29973
tri 27971 29961 27979 29969 ne
rect 27979 29965 28243 29969
tri 28243 29965 28251 29973 sw
rect 27979 29961 28251 29965
tri 27979 29953 27987 29961 ne
rect 27987 29957 28251 29961
tri 28251 29957 28259 29965 sw
rect 27987 29953 28259 29957
tri 27987 29945 27995 29953 ne
rect 27995 29949 28259 29953
tri 28259 29949 28267 29957 sw
rect 27995 29945 28267 29949
tri 27995 29937 28003 29945 ne
rect 28003 29941 28267 29945
tri 28267 29941 28275 29949 sw
rect 28003 29937 28275 29941
tri 28003 29933 28007 29937 ne
rect 28007 29933 28275 29937
tri 28275 29933 28283 29941 sw
tri 28007 29929 28011 29933 ne
rect 28011 29929 28283 29933
tri 28283 29929 28287 29933 sw
tri 28011 29921 28019 29929 ne
rect 28019 29921 28287 29929
tri 28287 29921 28295 29929 sw
tri 28019 29913 28027 29921 ne
rect 28027 29913 28295 29921
tri 28295 29913 28303 29921 sw
tri 28027 29905 28035 29913 ne
rect 28035 29905 28303 29913
tri 28303 29905 28311 29913 sw
tri 28035 29897 28043 29905 ne
rect 28043 29897 28311 29905
tri 28311 29897 28319 29905 sw
tri 28043 29889 28051 29897 ne
rect 28051 29889 28319 29897
tri 28319 29889 28327 29897 sw
tri 28051 29881 28059 29889 ne
rect 28059 29881 28327 29889
tri 28327 29881 28335 29889 sw
tri 28059 29873 28067 29881 ne
rect 28067 29873 28335 29881
tri 28335 29873 28343 29881 sw
tri 28067 29865 28075 29873 ne
rect 28075 29865 28343 29873
tri 28343 29865 28351 29873 sw
tri 28075 29857 28083 29865 ne
rect 28083 29857 28351 29865
tri 28351 29857 28359 29865 sw
tri 28083 29849 28091 29857 ne
rect 28091 29849 28359 29857
tri 28359 29849 28367 29857 sw
tri 28091 29841 28099 29849 ne
rect 28099 29841 28367 29849
tri 28367 29841 28375 29849 sw
tri 28099 29833 28107 29841 ne
rect 28107 29833 28375 29841
tri 28375 29833 28383 29841 sw
tri 28107 29825 28115 29833 ne
rect 28115 29825 28383 29833
tri 28383 29825 28391 29833 sw
tri 28115 29817 28123 29825 ne
rect 28123 29817 28391 29825
tri 28391 29817 28399 29825 sw
tri 28123 29809 28131 29817 ne
rect 28131 29809 28399 29817
tri 28399 29809 28407 29817 sw
tri 28131 29801 28139 29809 ne
rect 28139 29801 28407 29809
tri 28407 29801 28415 29809 sw
tri 28139 29793 28147 29801 ne
rect 28147 29793 28415 29801
tri 28415 29793 28423 29801 sw
tri 28147 29789 28151 29793 ne
rect 28151 29789 28423 29793
tri 28151 29781 28159 29789 ne
rect 28159 29785 28423 29789
tri 28423 29785 28431 29793 sw
rect 28159 29781 28431 29785
tri 28159 29773 28167 29781 ne
rect 28167 29777 28431 29781
tri 28431 29777 28439 29785 sw
rect 28167 29773 28439 29777
tri 28167 29765 28175 29773 ne
rect 28175 29769 28439 29773
tri 28439 29769 28447 29777 sw
rect 28175 29765 28447 29769
tri 28175 29757 28183 29765 ne
rect 28183 29761 28447 29765
tri 28447 29761 28455 29769 sw
rect 28183 29757 28455 29761
tri 28183 29749 28191 29757 ne
rect 28191 29753 28455 29757
tri 28455 29753 28463 29761 sw
rect 28191 29749 28463 29753
tri 28191 29741 28199 29749 ne
rect 28199 29745 28463 29749
tri 28463 29745 28471 29753 sw
rect 28199 29741 28471 29745
tri 28199 29733 28207 29741 ne
rect 28207 29737 28471 29741
tri 28471 29737 28479 29745 sw
rect 28207 29733 28479 29737
tri 28207 29725 28215 29733 ne
rect 28215 29729 28479 29733
tri 28479 29729 28487 29737 sw
rect 28215 29725 28487 29729
tri 28215 29717 28223 29725 ne
rect 28223 29721 28487 29725
tri 28487 29721 28495 29729 sw
rect 28223 29717 28495 29721
tri 28223 29709 28231 29717 ne
rect 28231 29713 28495 29717
tri 28495 29713 28503 29721 sw
rect 28231 29709 28503 29713
tri 28231 29701 28239 29709 ne
rect 28239 29705 28503 29709
tri 28503 29705 28511 29713 sw
rect 28239 29701 28511 29705
tri 28239 29693 28247 29701 ne
rect 28247 29697 28511 29701
tri 28511 29697 28519 29705 sw
rect 28247 29693 28519 29697
tri 28247 29685 28255 29693 ne
rect 28255 29689 28519 29693
tri 28519 29689 28527 29697 sw
rect 28255 29685 28527 29689
tri 28255 29677 28263 29685 ne
rect 28263 29681 28527 29685
tri 28527 29681 28535 29689 sw
rect 28263 29677 28535 29681
tri 28263 29669 28271 29677 ne
rect 28271 29673 28535 29677
tri 28535 29673 28543 29681 sw
rect 28271 29669 28543 29673
tri 28271 29661 28279 29669 ne
rect 28279 29665 28543 29669
tri 28543 29665 28551 29673 sw
rect 28279 29661 28551 29665
tri 28279 29657 28283 29661 ne
rect 28283 29657 28551 29661
tri 28551 29657 28559 29665 sw
tri 28283 29653 28287 29657 ne
rect 28287 29653 28559 29657
tri 28559 29653 28563 29657 sw
tri 28287 29645 28295 29653 ne
rect 28295 29645 28563 29653
tri 28563 29645 28571 29653 sw
tri 28295 29637 28303 29645 ne
rect 28303 29637 28571 29645
tri 28571 29637 28579 29645 sw
tri 28303 29629 28311 29637 ne
rect 28311 29629 28579 29637
tri 28579 29629 28587 29637 sw
tri 28311 29621 28319 29629 ne
rect 28319 29621 28587 29629
tri 28587 29621 28595 29629 sw
tri 28319 29613 28327 29621 ne
rect 28327 29613 28595 29621
tri 28595 29613 28603 29621 sw
tri 28327 29605 28335 29613 ne
rect 28335 29605 28603 29613
tri 28603 29605 28611 29613 sw
tri 28335 29597 28343 29605 ne
rect 28343 29597 28611 29605
tri 28611 29597 28619 29605 sw
tri 28343 29589 28351 29597 ne
rect 28351 29589 28619 29597
tri 28619 29589 28627 29597 sw
tri 28351 29581 28359 29589 ne
rect 28359 29581 28627 29589
tri 28627 29581 28635 29589 sw
tri 28359 29573 28367 29581 ne
rect 28367 29573 28635 29581
tri 28635 29573 28643 29581 sw
tri 28367 29565 28375 29573 ne
rect 28375 29565 28643 29573
tri 28643 29565 28651 29573 sw
tri 28375 29557 28383 29565 ne
rect 28383 29557 28651 29565
tri 28651 29557 28659 29565 sw
tri 28383 29549 28391 29557 ne
rect 28391 29549 28659 29557
tri 28659 29549 28667 29557 sw
tri 28391 29541 28399 29549 ne
rect 28399 29541 28667 29549
tri 28667 29541 28675 29549 sw
tri 28399 29533 28407 29541 ne
rect 28407 29533 28675 29541
tri 28675 29533 28683 29541 sw
tri 28407 29525 28415 29533 ne
rect 28415 29525 28683 29533
tri 28683 29525 28691 29533 sw
tri 28415 29517 28423 29525 ne
rect 28423 29517 28691 29525
tri 28691 29517 28699 29525 sw
tri 28423 29513 28427 29517 ne
rect 28427 29513 28699 29517
tri 28427 29505 28435 29513 ne
rect 28435 29509 28699 29513
tri 28699 29509 28707 29517 sw
rect 28435 29505 28707 29509
tri 28435 29497 28443 29505 ne
rect 28443 29501 28707 29505
tri 28707 29501 28715 29509 sw
rect 28443 29497 28715 29501
tri 28443 29489 28451 29497 ne
rect 28451 29493 28715 29497
tri 28715 29493 28723 29501 sw
rect 28451 29489 28723 29493
tri 28451 29481 28459 29489 ne
rect 28459 29485 28723 29489
tri 28723 29485 28731 29493 sw
rect 28459 29481 28731 29485
tri 28459 29473 28467 29481 ne
rect 28467 29477 28731 29481
tri 28731 29477 28739 29485 sw
rect 28467 29473 28739 29477
tri 28467 29465 28475 29473 ne
rect 28475 29469 28739 29473
tri 28739 29469 28747 29477 sw
rect 28475 29465 28747 29469
tri 28475 29457 28483 29465 ne
rect 28483 29461 28747 29465
tri 28747 29461 28755 29469 sw
rect 28483 29457 28755 29461
tri 28483 29449 28491 29457 ne
rect 28491 29453 28755 29457
tri 28755 29453 28763 29461 sw
rect 28491 29449 28763 29453
tri 28491 29441 28499 29449 ne
rect 28499 29445 28763 29449
tri 28763 29445 28771 29453 sw
rect 28499 29441 28771 29445
tri 28499 29433 28507 29441 ne
rect 28507 29437 28771 29441
tri 28771 29437 28779 29445 sw
rect 28507 29433 28779 29437
tri 28507 29425 28515 29433 ne
rect 28515 29429 28779 29433
tri 28779 29429 28787 29437 sw
rect 28515 29425 28787 29429
tri 28515 29417 28523 29425 ne
rect 28523 29421 28787 29425
tri 28787 29421 28795 29429 sw
rect 28523 29417 28795 29421
tri 28523 29409 28531 29417 ne
rect 28531 29413 28795 29417
tri 28795 29413 28803 29421 sw
rect 28531 29409 28803 29413
tri 28531 29401 28539 29409 ne
rect 28539 29405 28803 29409
tri 28803 29405 28811 29413 sw
rect 28539 29401 28811 29405
tri 28539 29393 28547 29401 ne
rect 28547 29397 28811 29401
tri 28811 29397 28819 29405 sw
rect 28547 29393 28819 29397
tri 28547 29385 28555 29393 ne
rect 28555 29389 28819 29393
tri 28819 29389 28827 29397 sw
rect 28555 29385 28827 29389
tri 28555 29381 28559 29385 ne
rect 28559 29381 28827 29385
tri 28827 29381 28835 29389 sw
tri 28559 29377 28563 29381 ne
rect 28563 29377 28835 29381
tri 28835 29377 28839 29381 sw
tri 28563 29369 28571 29377 ne
rect 28571 29369 28839 29377
tri 28839 29369 28847 29377 sw
tri 28571 29361 28579 29369 ne
rect 28579 29361 28847 29369
tri 28847 29361 28855 29369 sw
tri 28579 29353 28587 29361 ne
rect 28587 29353 28855 29361
tri 28855 29353 28863 29361 sw
tri 28587 29345 28595 29353 ne
rect 28595 29345 28863 29353
tri 28863 29345 28871 29353 sw
tri 28595 29337 28603 29345 ne
rect 28603 29337 28871 29345
tri 28871 29337 28879 29345 sw
tri 28603 29329 28611 29337 ne
rect 28611 29329 28879 29337
tri 28879 29329 28887 29337 sw
tri 28611 29321 28619 29329 ne
rect 28619 29321 28887 29329
tri 28887 29321 28895 29329 sw
tri 28619 29313 28627 29321 ne
rect 28627 29313 28895 29321
tri 28895 29313 28903 29321 sw
tri 28627 29305 28635 29313 ne
rect 28635 29305 28903 29313
tri 28903 29305 28911 29313 sw
tri 28635 29297 28643 29305 ne
rect 28643 29297 28911 29305
tri 28911 29297 28919 29305 sw
tri 28643 29289 28651 29297 ne
rect 28651 29289 28919 29297
tri 28919 29289 28927 29297 sw
tri 28651 29281 28659 29289 ne
rect 28659 29281 28927 29289
tri 28927 29281 28935 29289 sw
tri 28659 29273 28667 29281 ne
rect 28667 29273 28935 29281
tri 28935 29273 28943 29281 sw
tri 28667 29265 28675 29273 ne
rect 28675 29265 28943 29273
tri 28943 29265 28951 29273 sw
tri 28675 29257 28683 29265 ne
rect 28683 29257 28951 29265
tri 28951 29257 28959 29265 sw
tri 28683 29249 28691 29257 ne
rect 28691 29249 28959 29257
tri 28959 29249 28967 29257 sw
tri 28691 29241 28699 29249 ne
rect 28699 29241 28967 29249
tri 28967 29241 28975 29249 sw
tri 28699 29237 28703 29241 ne
rect 28703 29237 28975 29241
tri 28703 29229 28711 29237 ne
rect 28711 29233 28975 29237
tri 28975 29233 28983 29241 sw
rect 28711 29229 28983 29233
tri 28711 29221 28719 29229 ne
rect 28719 29225 28983 29229
tri 28983 29225 28991 29233 sw
rect 28719 29221 28991 29225
tri 28719 29213 28727 29221 ne
rect 28727 29217 28991 29221
tri 28991 29217 28999 29225 sw
rect 28727 29213 28999 29217
tri 28727 29205 28735 29213 ne
rect 28735 29209 28999 29213
tri 28999 29209 29007 29217 sw
rect 28735 29205 29007 29209
tri 28735 29197 28743 29205 ne
rect 28743 29201 29007 29205
tri 29007 29201 29015 29209 sw
rect 28743 29197 29015 29201
tri 28743 29189 28751 29197 ne
rect 28751 29193 29015 29197
tri 29015 29193 29023 29201 sw
rect 28751 29189 29023 29193
tri 28751 29181 28759 29189 ne
rect 28759 29185 29023 29189
tri 29023 29185 29031 29193 sw
rect 28759 29181 29031 29185
tri 28759 29173 28767 29181 ne
rect 28767 29177 29031 29181
tri 29031 29177 29039 29185 sw
rect 28767 29173 29039 29177
tri 28767 29165 28775 29173 ne
rect 28775 29169 29039 29173
tri 29039 29169 29047 29177 sw
rect 28775 29165 29047 29169
tri 28775 29157 28783 29165 ne
rect 28783 29161 29047 29165
tri 29047 29161 29055 29169 sw
rect 28783 29157 29055 29161
tri 28783 29149 28791 29157 ne
rect 28791 29153 29055 29157
tri 29055 29153 29063 29161 sw
rect 28791 29149 29063 29153
tri 28791 29141 28799 29149 ne
rect 28799 29145 29063 29149
tri 29063 29145 29071 29153 sw
rect 28799 29141 29071 29145
tri 28799 29133 28807 29141 ne
rect 28807 29137 29071 29141
tri 29071 29137 29079 29145 sw
rect 28807 29133 29079 29137
tri 28807 29125 28815 29133 ne
rect 28815 29129 29079 29133
tri 29079 29129 29087 29137 sw
rect 28815 29125 29087 29129
tri 28815 29117 28823 29125 ne
rect 28823 29121 29087 29125
tri 29087 29121 29095 29129 sw
rect 28823 29117 29095 29121
tri 28823 29109 28831 29117 ne
rect 28831 29113 29095 29117
tri 29095 29113 29103 29121 sw
rect 28831 29109 29103 29113
tri 28831 29105 28835 29109 ne
rect 28835 29105 29103 29109
tri 29103 29105 29111 29113 sw
tri 28835 29101 28839 29105 ne
rect 28839 29101 29111 29105
tri 29111 29101 29115 29105 sw
tri 28839 29093 28847 29101 ne
rect 28847 29093 29115 29101
tri 29115 29093 29123 29101 sw
tri 28847 29085 28855 29093 ne
rect 28855 29085 29123 29093
tri 29123 29085 29131 29093 sw
tri 28855 29077 28863 29085 ne
rect 28863 29077 29131 29085
tri 29131 29077 29139 29085 sw
tri 28863 29069 28871 29077 ne
rect 28871 29069 29139 29077
tri 29139 29069 29147 29077 sw
tri 28871 29061 28879 29069 ne
rect 28879 29061 29147 29069
tri 29147 29061 29155 29069 sw
tri 28879 29053 28887 29061 ne
rect 28887 29053 29155 29061
tri 29155 29053 29163 29061 sw
tri 28887 29045 28895 29053 ne
rect 28895 29045 29163 29053
tri 29163 29045 29171 29053 sw
tri 28895 29037 28903 29045 ne
rect 28903 29037 29171 29045
tri 29171 29037 29179 29045 sw
tri 28903 29029 28911 29037 ne
rect 28911 29029 29179 29037
tri 29179 29029 29187 29037 sw
tri 28911 29021 28919 29029 ne
rect 28919 29021 29187 29029
tri 29187 29021 29195 29029 sw
tri 28919 29013 28927 29021 ne
rect 28927 29013 29195 29021
tri 29195 29013 29203 29021 sw
tri 28927 29005 28935 29013 ne
rect 28935 29005 29203 29013
tri 29203 29005 29211 29013 sw
tri 28935 28997 28943 29005 ne
rect 28943 28997 29211 29005
tri 29211 28997 29219 29005 sw
tri 28943 28989 28951 28997 ne
rect 28951 28989 29219 28997
tri 29219 28989 29227 28997 sw
tri 28951 28981 28959 28989 ne
rect 28959 28981 29227 28989
tri 29227 28981 29235 28989 sw
tri 28959 28973 28967 28981 ne
rect 28967 28973 29235 28981
tri 29235 28973 29243 28981 sw
tri 28967 28965 28975 28973 ne
rect 28975 28965 29243 28973
tri 29243 28965 29251 28973 sw
tri 28975 28961 28979 28965 ne
rect 28979 28961 29251 28965
tri 28979 28953 28987 28961 ne
rect 28987 28957 29251 28961
tri 29251 28957 29259 28965 sw
rect 28987 28953 29259 28957
tri 28987 28945 28995 28953 ne
rect 28995 28949 29259 28953
tri 29259 28949 29267 28957 sw
rect 28995 28945 29267 28949
tri 28995 28937 29003 28945 ne
rect 29003 28941 29267 28945
tri 29267 28941 29275 28949 sw
rect 29003 28937 29275 28941
tri 29003 28929 29011 28937 ne
rect 29011 28933 29275 28937
tri 29275 28933 29283 28941 sw
rect 29011 28929 29283 28933
tri 29011 28921 29019 28929 ne
rect 29019 28925 29283 28929
tri 29283 28925 29291 28933 sw
rect 29019 28921 29291 28925
tri 29019 28913 29027 28921 ne
rect 29027 28917 29291 28921
tri 29291 28917 29299 28925 sw
rect 29027 28913 29299 28917
tri 29027 28905 29035 28913 ne
rect 29035 28909 29299 28913
tri 29299 28909 29307 28917 sw
rect 29035 28905 29307 28909
tri 29035 28897 29043 28905 ne
rect 29043 28901 29307 28905
tri 29307 28901 29315 28909 sw
rect 29043 28897 29315 28901
tri 29043 28889 29051 28897 ne
rect 29051 28893 29315 28897
tri 29315 28893 29323 28901 sw
rect 29051 28889 29323 28893
tri 29051 28881 29059 28889 ne
rect 29059 28885 29323 28889
tri 29323 28885 29331 28893 sw
rect 29059 28881 29331 28885
tri 29059 28873 29067 28881 ne
rect 29067 28877 29331 28881
tri 29331 28877 29339 28885 sw
rect 29067 28873 29339 28877
tri 29067 28865 29075 28873 ne
rect 29075 28869 29339 28873
tri 29339 28869 29347 28877 sw
rect 29075 28865 29347 28869
tri 29075 28857 29083 28865 ne
rect 29083 28861 29347 28865
tri 29347 28861 29355 28869 sw
rect 29083 28857 29355 28861
tri 29083 28849 29091 28857 ne
rect 29091 28853 29355 28857
tri 29355 28853 29363 28861 sw
rect 29091 28849 29363 28853
tri 29091 28841 29099 28849 ne
rect 29099 28845 29363 28849
tri 29363 28845 29371 28853 sw
rect 29099 28841 29371 28845
tri 29099 28833 29107 28841 ne
rect 29107 28837 29371 28841
tri 29371 28837 29379 28845 sw
rect 29107 28833 29379 28837
tri 29107 28829 29111 28833 ne
rect 29111 28829 29379 28833
tri 29379 28829 29387 28837 sw
tri 29111 28825 29115 28829 ne
rect 29115 28825 29387 28829
tri 29387 28825 29391 28829 sw
tri 29115 28817 29123 28825 ne
rect 29123 28817 29391 28825
tri 29391 28817 29399 28825 sw
tri 29123 28809 29131 28817 ne
rect 29131 28809 29399 28817
tri 29399 28809 29407 28817 sw
tri 29131 28801 29139 28809 ne
rect 29139 28801 29407 28809
tri 29407 28801 29415 28809 sw
tri 29139 28793 29147 28801 ne
rect 29147 28793 29415 28801
tri 29415 28793 29423 28801 sw
tri 29147 28785 29155 28793 ne
rect 29155 28785 29423 28793
tri 29423 28785 29431 28793 sw
tri 29155 28777 29163 28785 ne
rect 29163 28777 29431 28785
tri 29431 28777 29439 28785 sw
tri 29163 28769 29171 28777 ne
rect 29171 28769 29439 28777
tri 29439 28769 29447 28777 sw
tri 29171 28761 29179 28769 ne
rect 29179 28761 29447 28769
tri 29447 28761 29455 28769 sw
tri 29179 28753 29187 28761 ne
rect 29187 28753 29455 28761
tri 29455 28753 29463 28761 sw
tri 29187 28745 29195 28753 ne
rect 29195 28745 29463 28753
tri 29463 28745 29471 28753 sw
tri 29195 28737 29203 28745 ne
rect 29203 28737 29471 28745
tri 29471 28737 29479 28745 sw
tri 29203 28729 29211 28737 ne
rect 29211 28729 29479 28737
tri 29479 28729 29487 28737 sw
tri 29211 28721 29219 28729 ne
rect 29219 28721 29487 28729
tri 29487 28721 29495 28729 sw
tri 29219 28713 29227 28721 ne
rect 29227 28713 29495 28721
tri 29495 28713 29503 28721 sw
tri 29227 28705 29235 28713 ne
rect 29235 28705 29503 28713
tri 29503 28705 29511 28713 sw
tri 29235 28697 29243 28705 ne
rect 29243 28697 29511 28705
tri 29511 28697 29519 28705 sw
tri 29243 28689 29251 28697 ne
rect 29251 28689 29519 28697
tri 29519 28689 29527 28697 sw
tri 29251 28685 29255 28689 ne
rect 29255 28685 29527 28689
tri 29255 28677 29263 28685 ne
rect 29263 28681 29527 28685
tri 29527 28681 29535 28689 sw
rect 29263 28677 29535 28681
tri 29263 28669 29271 28677 ne
rect 29271 28673 29535 28677
tri 29535 28673 29543 28681 sw
rect 29271 28669 29543 28673
tri 29271 28661 29279 28669 ne
rect 29279 28665 29543 28669
tri 29543 28665 29551 28673 sw
rect 29279 28661 29551 28665
tri 29279 28653 29287 28661 ne
rect 29287 28657 29551 28661
tri 29551 28657 29559 28665 sw
rect 29287 28653 29559 28657
tri 29287 28645 29295 28653 ne
rect 29295 28649 29559 28653
tri 29559 28649 29567 28657 sw
rect 29295 28645 29567 28649
tri 29295 28637 29303 28645 ne
rect 29303 28641 29567 28645
tri 29567 28641 29575 28649 sw
rect 29303 28637 29575 28641
tri 29303 28629 29311 28637 ne
rect 29311 28633 29575 28637
tri 29575 28633 29583 28641 sw
rect 29311 28629 29583 28633
tri 29311 28621 29319 28629 ne
rect 29319 28625 29583 28629
tri 29583 28625 29591 28633 sw
rect 29319 28621 29591 28625
tri 29319 28613 29327 28621 ne
rect 29327 28617 29591 28621
tri 29591 28617 29599 28625 sw
rect 29327 28613 29599 28617
tri 29327 28605 29335 28613 ne
rect 29335 28609 29599 28613
tri 29599 28609 29607 28617 sw
rect 29335 28605 29607 28609
tri 29335 28597 29343 28605 ne
rect 29343 28601 29607 28605
tri 29607 28601 29615 28609 sw
rect 29343 28597 29615 28601
tri 29343 28589 29351 28597 ne
rect 29351 28593 29615 28597
tri 29615 28593 29623 28601 sw
rect 29351 28589 29623 28593
tri 29351 28581 29359 28589 ne
rect 29359 28585 29623 28589
tri 29623 28585 29631 28593 sw
rect 29359 28581 29631 28585
tri 29359 28573 29367 28581 ne
rect 29367 28577 29631 28581
tri 29631 28577 29639 28585 sw
rect 29367 28573 29639 28577
tri 29367 28565 29375 28573 ne
rect 29375 28569 29639 28573
tri 29639 28569 29647 28577 sw
rect 29375 28565 29647 28569
tri 29375 28557 29383 28565 ne
rect 29383 28561 29647 28565
tri 29647 28561 29655 28569 sw
rect 29383 28557 29655 28561
tri 29383 28553 29387 28557 ne
rect 29387 28553 29655 28557
tri 29655 28553 29663 28561 sw
tri 29387 28549 29391 28553 ne
rect 29391 28549 29663 28553
tri 29663 28549 29667 28553 sw
tri 29391 28541 29399 28549 ne
rect 29399 28541 29667 28549
tri 29667 28541 29675 28549 sw
tri 29399 28533 29407 28541 ne
rect 29407 28533 29675 28541
tri 29675 28533 29683 28541 sw
tri 29407 28525 29415 28533 ne
rect 29415 28525 29683 28533
tri 29683 28525 29691 28533 sw
tri 29415 28517 29423 28525 ne
rect 29423 28517 29691 28525
tri 29691 28517 29699 28525 sw
tri 29423 28509 29431 28517 ne
rect 29431 28509 29699 28517
tri 29699 28509 29707 28517 sw
tri 29431 28501 29439 28509 ne
rect 29439 28501 29707 28509
tri 29707 28501 29715 28509 sw
tri 29439 28493 29447 28501 ne
rect 29447 28493 29715 28501
tri 29715 28493 29723 28501 sw
tri 29447 28485 29455 28493 ne
rect 29455 28485 29723 28493
tri 29723 28485 29731 28493 sw
tri 29455 28477 29463 28485 ne
rect 29463 28477 29731 28485
tri 29731 28477 29739 28485 sw
tri 29463 28469 29471 28477 ne
rect 29471 28469 29739 28477
tri 29739 28469 29747 28477 sw
tri 29471 28461 29479 28469 ne
rect 29479 28461 29747 28469
tri 29747 28461 29755 28469 sw
tri 29479 28453 29487 28461 ne
rect 29487 28453 29755 28461
tri 29755 28453 29763 28461 sw
tri 29487 28445 29495 28453 ne
rect 29495 28445 29763 28453
tri 29763 28445 29771 28453 sw
tri 29495 28437 29503 28445 ne
rect 29503 28437 29771 28445
tri 29771 28437 29779 28445 sw
tri 29503 28429 29511 28437 ne
rect 29511 28429 29779 28437
tri 29779 28429 29787 28437 sw
tri 29511 28421 29519 28429 ne
rect 29519 28421 29787 28429
tri 29787 28421 29795 28429 sw
tri 29519 28413 29527 28421 ne
rect 29527 28413 29795 28421
tri 29795 28413 29803 28421 sw
tri 29527 28409 29531 28413 ne
rect 29531 28409 29803 28413
tri 29531 28401 29539 28409 ne
rect 29539 28405 29803 28409
tri 29803 28405 29811 28413 sw
rect 29539 28401 29811 28405
tri 29539 28393 29547 28401 ne
rect 29547 28397 29811 28401
tri 29811 28397 29819 28405 sw
rect 29547 28393 29819 28397
tri 29547 28385 29555 28393 ne
rect 29555 28389 29819 28393
tri 29819 28389 29827 28397 sw
rect 29555 28385 29827 28389
tri 29555 28377 29563 28385 ne
rect 29563 28381 29827 28385
tri 29827 28381 29835 28389 sw
rect 29563 28377 29835 28381
tri 29563 28369 29571 28377 ne
rect 29571 28373 29835 28377
tri 29835 28373 29843 28381 sw
rect 29571 28369 29843 28373
tri 29571 28361 29579 28369 ne
rect 29579 28365 29843 28369
tri 29843 28365 29851 28373 sw
rect 29579 28361 29851 28365
tri 29579 28353 29587 28361 ne
rect 29587 28357 29851 28361
tri 29851 28357 29859 28365 sw
rect 29587 28353 29859 28357
tri 29587 28345 29595 28353 ne
rect 29595 28349 29859 28353
tri 29859 28349 29867 28357 sw
rect 29595 28345 29867 28349
tri 29595 28337 29603 28345 ne
rect 29603 28341 29867 28345
tri 29867 28341 29875 28349 sw
rect 29603 28337 29875 28341
tri 29603 28329 29611 28337 ne
rect 29611 28333 29875 28337
tri 29875 28333 29883 28341 sw
rect 29611 28329 29883 28333
tri 29611 28321 29619 28329 ne
rect 29619 28325 29883 28329
tri 29883 28325 29891 28333 sw
rect 29619 28321 29891 28325
tri 29619 28313 29627 28321 ne
rect 29627 28317 29891 28321
tri 29891 28317 29899 28325 sw
rect 29627 28313 29899 28317
tri 29627 28305 29635 28313 ne
rect 29635 28309 29899 28313
tri 29899 28309 29907 28317 sw
rect 29635 28305 29907 28309
tri 29635 28297 29643 28305 ne
rect 29643 28301 29907 28305
tri 29907 28301 29915 28309 sw
rect 29643 28297 29915 28301
tri 29643 28289 29651 28297 ne
rect 29651 28293 29915 28297
tri 29915 28293 29923 28301 sw
rect 29651 28289 29923 28293
tri 29651 28281 29659 28289 ne
rect 29659 28285 29923 28289
tri 29923 28285 29931 28293 sw
rect 29659 28281 29931 28285
tri 29659 28277 29663 28281 ne
rect 29663 28277 29931 28281
tri 29931 28277 29939 28285 sw
tri 29663 28273 29667 28277 ne
rect 29667 28273 29939 28277
tri 29939 28273 29943 28277 sw
tri 29667 28265 29675 28273 ne
rect 29675 28265 29943 28273
tri 29943 28265 29951 28273 sw
tri 29675 28257 29683 28265 ne
rect 29683 28257 29951 28265
tri 29951 28257 29959 28265 sw
tri 29683 28249 29691 28257 ne
rect 29691 28249 29959 28257
tri 29959 28249 29967 28257 sw
tri 29691 28241 29699 28249 ne
rect 29699 28241 29967 28249
tri 29967 28241 29975 28249 sw
tri 29699 28233 29707 28241 ne
rect 29707 28233 29975 28241
tri 29975 28233 29983 28241 sw
tri 29707 28225 29715 28233 ne
rect 29715 28225 29983 28233
tri 29983 28225 29991 28233 sw
tri 29715 28217 29723 28225 ne
rect 29723 28217 29991 28225
tri 29991 28217 29999 28225 sw
tri 29723 28209 29731 28217 ne
rect 29731 28209 29999 28217
tri 29999 28209 30007 28217 sw
tri 29731 28201 29739 28209 ne
rect 29739 28201 30007 28209
tri 30007 28201 30015 28209 sw
tri 29739 28193 29747 28201 ne
rect 29747 28193 30015 28201
tri 30015 28193 30023 28201 sw
tri 29747 28185 29755 28193 ne
rect 29755 28185 30023 28193
tri 30023 28185 30031 28193 sw
tri 29755 28177 29763 28185 ne
rect 29763 28177 30031 28185
tri 30031 28177 30039 28185 sw
tri 29763 28169 29771 28177 ne
rect 29771 28169 30039 28177
tri 30039 28169 30047 28177 sw
tri 29771 28161 29779 28169 ne
rect 29779 28161 30047 28169
tri 30047 28161 30055 28169 sw
tri 29779 28153 29787 28161 ne
rect 29787 28153 30055 28161
tri 30055 28153 30063 28161 sw
tri 29787 28145 29795 28153 ne
rect 29795 28145 30063 28153
tri 30063 28145 30071 28153 sw
tri 29795 28137 29803 28145 ne
rect 29803 28137 30071 28145
tri 30071 28137 30079 28145 sw
tri 29803 28133 29807 28137 ne
rect 29807 28133 30079 28137
tri 29807 28125 29815 28133 ne
rect 29815 28129 30079 28133
tri 30079 28129 30087 28137 sw
rect 29815 28125 30087 28129
tri 29815 28117 29823 28125 ne
rect 29823 28121 30087 28125
tri 30087 28121 30095 28129 sw
rect 29823 28117 30095 28121
tri 29823 28109 29831 28117 ne
rect 29831 28113 30095 28117
tri 30095 28113 30103 28121 sw
rect 29831 28109 30103 28113
tri 29831 28101 29839 28109 ne
rect 29839 28105 30103 28109
tri 30103 28105 30111 28113 sw
rect 29839 28101 30111 28105
tri 29839 28093 29847 28101 ne
rect 29847 28097 30111 28101
tri 30111 28097 30119 28105 sw
rect 29847 28093 30119 28097
tri 29847 28085 29855 28093 ne
rect 29855 28089 30119 28093
tri 30119 28089 30127 28097 sw
rect 29855 28085 30127 28089
tri 29855 28077 29863 28085 ne
rect 29863 28081 30127 28085
tri 30127 28081 30135 28089 sw
rect 29863 28077 30135 28081
tri 29863 28069 29871 28077 ne
rect 29871 28073 30135 28077
tri 30135 28073 30143 28081 sw
rect 29871 28069 30143 28073
tri 29871 28061 29879 28069 ne
rect 29879 28065 30143 28069
tri 30143 28065 30151 28073 sw
rect 29879 28061 30151 28065
tri 29879 28053 29887 28061 ne
rect 29887 28057 30151 28061
tri 30151 28057 30159 28065 sw
rect 29887 28053 30159 28057
tri 29887 28045 29895 28053 ne
rect 29895 28049 30159 28053
tri 30159 28049 30167 28057 sw
rect 29895 28045 30167 28049
tri 29895 28037 29903 28045 ne
rect 29903 28041 30167 28045
tri 30167 28041 30175 28049 sw
rect 29903 28037 30175 28041
tri 29903 28029 29911 28037 ne
rect 29911 28033 30175 28037
tri 30175 28033 30183 28041 sw
rect 29911 28029 30183 28033
tri 29911 28021 29919 28029 ne
rect 29919 28025 30183 28029
tri 30183 28025 30191 28033 sw
rect 29919 28021 30191 28025
tri 29919 28013 29927 28021 ne
rect 29927 28017 30191 28021
tri 30191 28017 30199 28025 sw
rect 29927 28013 30199 28017
tri 29927 28005 29935 28013 ne
rect 29935 28009 30199 28013
tri 30199 28009 30207 28017 sw
rect 29935 28005 30207 28009
tri 29935 28001 29939 28005 ne
rect 29939 28001 30207 28005
tri 30207 28001 30215 28009 sw
tri 29939 27997 29943 28001 ne
rect 29943 27997 30215 28001
tri 30215 27997 30219 28001 sw
tri 29943 27989 29951 27997 ne
rect 29951 27989 30219 27997
tri 30219 27989 30227 27997 sw
tri 29951 27981 29959 27989 ne
rect 29959 27981 30227 27989
tri 30227 27981 30235 27989 sw
tri 29959 27973 29967 27981 ne
rect 29967 27973 30235 27981
tri 30235 27973 30243 27981 sw
tri 29967 27965 29975 27973 ne
rect 29975 27965 30243 27973
tri 30243 27965 30251 27973 sw
tri 29975 27957 29983 27965 ne
rect 29983 27957 30251 27965
tri 30251 27957 30259 27965 sw
tri 29983 27949 29991 27957 ne
rect 29991 27949 30259 27957
tri 30259 27949 30267 27957 sw
tri 29991 27941 29999 27949 ne
rect 29999 27941 30267 27949
tri 30267 27941 30275 27949 sw
tri 29999 27933 30007 27941 ne
rect 30007 27933 30275 27941
tri 30275 27933 30283 27941 sw
tri 30007 27925 30015 27933 ne
rect 30015 27925 30283 27933
tri 30283 27925 30291 27933 sw
tri 30015 27917 30023 27925 ne
rect 30023 27917 30291 27925
tri 30291 27917 30299 27925 sw
tri 30023 27909 30031 27917 ne
rect 30031 27909 30299 27917
tri 30299 27909 30307 27917 sw
tri 30031 27901 30039 27909 ne
rect 30039 27901 30307 27909
tri 30307 27901 30315 27909 sw
tri 30039 27893 30047 27901 ne
rect 30047 27893 30315 27901
tri 30315 27893 30323 27901 sw
tri 30047 27885 30055 27893 ne
rect 30055 27885 30323 27893
tri 30323 27885 30331 27893 sw
tri 30055 27877 30063 27885 ne
rect 30063 27877 30331 27885
tri 30331 27877 30339 27885 sw
tri 30063 27869 30071 27877 ne
rect 30071 27869 30339 27877
tri 30339 27869 30347 27877 sw
tri 30071 27861 30079 27869 ne
rect 30079 27861 30347 27869
tri 30347 27861 30355 27869 sw
tri 30079 27857 30083 27861 ne
rect 30083 27857 30355 27861
tri 30083 27849 30091 27857 ne
rect 30091 27853 30355 27857
tri 30355 27853 30363 27861 sw
rect 30091 27849 30363 27853
tri 30091 27841 30099 27849 ne
rect 30099 27845 30363 27849
tri 30363 27845 30371 27853 sw
rect 30099 27841 30371 27845
tri 30099 27833 30107 27841 ne
rect 30107 27837 30371 27841
tri 30371 27837 30379 27845 sw
rect 30107 27833 30379 27837
tri 30107 27825 30115 27833 ne
rect 30115 27829 30379 27833
tri 30379 27829 30387 27837 sw
rect 30115 27825 30387 27829
tri 30115 27817 30123 27825 ne
rect 30123 27821 30387 27825
tri 30387 27821 30395 27829 sw
rect 30123 27817 30395 27821
tri 30123 27809 30131 27817 ne
rect 30131 27813 30395 27817
tri 30395 27813 30403 27821 sw
rect 30131 27809 30403 27813
tri 30131 27801 30139 27809 ne
rect 30139 27805 30403 27809
tri 30403 27805 30411 27813 sw
rect 30139 27801 30411 27805
tri 30139 27793 30147 27801 ne
rect 30147 27797 30411 27801
tri 30411 27797 30419 27805 sw
rect 30147 27793 30419 27797
tri 30147 27785 30155 27793 ne
rect 30155 27789 30419 27793
tri 30419 27789 30427 27797 sw
rect 30155 27785 30427 27789
tri 30155 27777 30163 27785 ne
rect 30163 27781 30427 27785
tri 30427 27781 30435 27789 sw
rect 30163 27777 30435 27781
tri 30163 27769 30171 27777 ne
rect 30171 27773 30435 27777
tri 30435 27773 30443 27781 sw
rect 30171 27769 30443 27773
tri 30171 27761 30179 27769 ne
rect 30179 27765 30443 27769
tri 30443 27765 30451 27773 sw
rect 30179 27761 30451 27765
tri 30179 27753 30187 27761 ne
rect 30187 27757 30451 27761
tri 30451 27757 30459 27765 sw
rect 30187 27753 30459 27757
tri 30187 27745 30195 27753 ne
rect 30195 27749 30459 27753
tri 30459 27749 30467 27757 sw
rect 30195 27745 30467 27749
tri 30195 27737 30203 27745 ne
rect 30203 27741 30467 27745
tri 30467 27741 30475 27749 sw
rect 30203 27737 30475 27741
tri 30203 27729 30211 27737 ne
rect 30211 27733 30475 27737
tri 30475 27733 30483 27741 sw
rect 30211 27729 30483 27733
tri 30211 27725 30215 27729 ne
rect 30215 27725 30483 27729
tri 30483 27725 30491 27733 sw
tri 30215 27721 30219 27725 ne
rect 30219 27721 30491 27725
tri 30491 27721 30495 27725 sw
tri 30219 27713 30227 27721 ne
rect 30227 27713 30495 27721
tri 30495 27713 30503 27721 sw
tri 30227 27705 30235 27713 ne
rect 30235 27705 30503 27713
tri 30503 27705 30511 27713 sw
tri 30235 27697 30243 27705 ne
rect 30243 27697 30511 27705
tri 30511 27697 30519 27705 sw
tri 30243 27689 30251 27697 ne
rect 30251 27689 30519 27697
tri 30519 27689 30527 27697 sw
tri 30251 27681 30259 27689 ne
rect 30259 27681 30527 27689
tri 30527 27681 30535 27689 sw
tri 30259 27673 30267 27681 ne
rect 30267 27673 30535 27681
tri 30535 27673 30543 27681 sw
tri 30267 27665 30275 27673 ne
rect 30275 27665 30543 27673
tri 30543 27665 30551 27673 sw
tri 30275 27657 30283 27665 ne
rect 30283 27657 30551 27665
tri 30551 27657 30559 27665 sw
tri 30283 27649 30291 27657 ne
rect 30291 27649 30559 27657
tri 30559 27649 30567 27657 sw
tri 30291 27641 30299 27649 ne
rect 30299 27641 30567 27649
tri 30567 27641 30575 27649 sw
tri 30299 27633 30307 27641 ne
rect 30307 27633 30575 27641
tri 30575 27633 30583 27641 sw
tri 30307 27625 30315 27633 ne
rect 30315 27625 30583 27633
tri 30583 27625 30591 27633 sw
tri 30315 27617 30323 27625 ne
rect 30323 27617 30591 27625
tri 30591 27617 30599 27625 sw
tri 30323 27609 30331 27617 ne
rect 30331 27609 30599 27617
tri 30599 27609 30607 27617 sw
tri 30331 27601 30339 27609 ne
rect 30339 27601 30607 27609
tri 30607 27601 30615 27609 sw
tri 30339 27593 30347 27601 ne
rect 30347 27593 30615 27601
tri 30615 27593 30623 27601 sw
tri 30347 27585 30355 27593 ne
rect 30355 27585 30623 27593
tri 30623 27585 30631 27593 sw
tri 30355 27581 30359 27585 ne
rect 30359 27581 30631 27585
tri 30359 27573 30367 27581 ne
rect 30367 27577 30631 27581
tri 30631 27577 30639 27585 sw
rect 30367 27573 30639 27577
tri 30367 27565 30375 27573 ne
rect 30375 27569 30639 27573
tri 30639 27569 30647 27577 sw
rect 30375 27565 30647 27569
tri 30375 27557 30383 27565 ne
rect 30383 27561 30647 27565
tri 30647 27561 30655 27569 sw
rect 30383 27557 30655 27561
tri 30383 27549 30391 27557 ne
rect 30391 27553 30655 27557
tri 30655 27553 30663 27561 sw
rect 30391 27549 30663 27553
tri 30391 27541 30399 27549 ne
rect 30399 27545 30663 27549
tri 30663 27545 30671 27553 sw
rect 30399 27541 30671 27545
tri 30399 27533 30407 27541 ne
rect 30407 27537 30671 27541
tri 30671 27537 30679 27545 sw
rect 30407 27533 30679 27537
tri 30407 27525 30415 27533 ne
rect 30415 27529 30679 27533
tri 30679 27529 30687 27537 sw
rect 30415 27525 30687 27529
tri 30415 27517 30423 27525 ne
rect 30423 27521 30687 27525
tri 30687 27521 30695 27529 sw
rect 30423 27517 30695 27521
tri 30423 27509 30431 27517 ne
rect 30431 27513 30695 27517
tri 30695 27513 30703 27521 sw
rect 30431 27509 30703 27513
tri 30431 27501 30439 27509 ne
rect 30439 27505 30703 27509
tri 30703 27505 30711 27513 sw
rect 30439 27501 30711 27505
tri 30439 27493 30447 27501 ne
rect 30447 27497 30711 27501
tri 30711 27497 30719 27505 sw
rect 30447 27493 30719 27497
tri 30447 27485 30455 27493 ne
rect 30455 27489 30719 27493
tri 30719 27489 30727 27497 sw
rect 30455 27485 30727 27489
tri 30455 27477 30463 27485 ne
rect 30463 27481 30727 27485
tri 30727 27481 30735 27489 sw
rect 30463 27477 30735 27481
tri 30463 27469 30471 27477 ne
rect 30471 27473 30735 27477
tri 30735 27473 30743 27481 sw
rect 30471 27469 30743 27473
tri 30471 27461 30479 27469 ne
rect 30479 27465 30743 27469
tri 30743 27465 30751 27473 sw
rect 30479 27461 30751 27465
tri 30479 27453 30487 27461 ne
rect 30487 27457 30751 27461
tri 30751 27457 30759 27465 sw
rect 30487 27453 30759 27457
tri 30487 27449 30491 27453 ne
rect 30491 27449 30759 27453
tri 30759 27449 30767 27457 sw
tri 30491 27445 30495 27449 ne
rect 30495 27445 30767 27449
tri 30767 27445 30771 27449 sw
tri 30495 27437 30503 27445 ne
rect 30503 27437 30771 27445
tri 30771 27437 30779 27445 sw
tri 30503 27429 30511 27437 ne
rect 30511 27429 30779 27437
tri 30779 27429 30787 27437 sw
tri 30511 27421 30519 27429 ne
rect 30519 27421 30787 27429
tri 30787 27421 30795 27429 sw
tri 30519 27413 30527 27421 ne
rect 30527 27413 30795 27421
tri 30795 27413 30803 27421 sw
tri 30527 27405 30535 27413 ne
rect 30535 27405 30803 27413
tri 30803 27405 30811 27413 sw
tri 30535 27397 30543 27405 ne
rect 30543 27397 30811 27405
tri 30811 27397 30819 27405 sw
tri 30543 27389 30551 27397 ne
rect 30551 27389 30819 27397
tri 30819 27389 30827 27397 sw
tri 30551 27381 30559 27389 ne
rect 30559 27381 30827 27389
tri 30827 27381 30835 27389 sw
tri 30559 27373 30567 27381 ne
rect 30567 27373 30835 27381
tri 30835 27373 30843 27381 sw
tri 30567 27365 30575 27373 ne
rect 30575 27365 30843 27373
tri 30843 27365 30851 27373 sw
tri 30575 27357 30583 27365 ne
rect 30583 27357 30851 27365
tri 30851 27357 30859 27365 sw
tri 30583 27349 30591 27357 ne
rect 30591 27349 30859 27357
tri 30859 27349 30867 27357 sw
tri 30591 27341 30599 27349 ne
rect 30599 27341 30867 27349
tri 30867 27341 30875 27349 sw
tri 30599 27333 30607 27341 ne
rect 30607 27333 30875 27341
tri 30875 27333 30883 27341 sw
tri 30607 27325 30615 27333 ne
rect 30615 27325 30883 27333
tri 30883 27325 30891 27333 sw
tri 30615 27317 30623 27325 ne
rect 30623 27317 30891 27325
tri 30891 27317 30899 27325 sw
tri 30623 27309 30631 27317 ne
rect 30631 27309 30899 27317
tri 30899 27309 30907 27317 sw
tri 30631 27305 30635 27309 ne
rect 30635 27305 30907 27309
tri 30635 27297 30643 27305 ne
rect 30643 27301 30907 27305
tri 30907 27301 30915 27309 sw
rect 30643 27297 30915 27301
tri 30643 27289 30651 27297 ne
rect 30651 27293 30915 27297
tri 30915 27293 30923 27301 sw
rect 30651 27289 30923 27293
tri 30651 27281 30659 27289 ne
rect 30659 27285 30923 27289
tri 30923 27285 30931 27293 sw
rect 30659 27281 30931 27285
tri 30659 27273 30667 27281 ne
rect 30667 27277 30931 27281
tri 30931 27277 30939 27285 sw
rect 30667 27273 30939 27277
tri 30667 27265 30675 27273 ne
rect 30675 27269 30939 27273
tri 30939 27269 30947 27277 sw
rect 30675 27265 30947 27269
tri 30675 27257 30683 27265 ne
rect 30683 27261 30947 27265
tri 30947 27261 30955 27269 sw
rect 30683 27257 30955 27261
tri 30683 27249 30691 27257 ne
rect 30691 27253 30955 27257
tri 30955 27253 30963 27261 sw
rect 30691 27249 30963 27253
tri 30691 27241 30699 27249 ne
rect 30699 27245 30963 27249
tri 30963 27245 30971 27253 sw
rect 30699 27241 30971 27245
tri 30699 27233 30707 27241 ne
rect 30707 27237 30971 27241
tri 30971 27237 30979 27245 sw
rect 30707 27233 30979 27237
tri 30707 27225 30715 27233 ne
rect 30715 27229 30979 27233
tri 30979 27229 30987 27237 sw
rect 30715 27225 30987 27229
tri 30715 27217 30723 27225 ne
rect 30723 27221 30987 27225
tri 30987 27221 30995 27229 sw
rect 30723 27217 30995 27221
tri 30723 27209 30731 27217 ne
rect 30731 27213 30995 27217
tri 30995 27213 31003 27221 sw
rect 30731 27209 31003 27213
tri 30731 27201 30739 27209 ne
rect 30739 27205 31003 27209
tri 31003 27205 31011 27213 sw
rect 30739 27201 31011 27205
tri 30739 27193 30747 27201 ne
rect 30747 27197 31011 27201
tri 31011 27197 31019 27205 sw
rect 30747 27193 31019 27197
tri 30747 27185 30755 27193 ne
rect 30755 27189 31019 27193
tri 31019 27189 31027 27197 sw
rect 30755 27185 31027 27189
tri 30755 27177 30763 27185 ne
rect 30763 27181 31027 27185
tri 31027 27181 31035 27189 sw
rect 30763 27177 31035 27181
tri 30763 27173 30767 27177 ne
rect 30767 27173 31035 27177
tri 31035 27173 31043 27181 sw
tri 30767 27169 30771 27173 ne
rect 30771 27169 31043 27173
tri 31043 27169 31047 27173 sw
tri 30771 27161 30779 27169 ne
rect 30779 27161 31047 27169
tri 31047 27161 31055 27169 sw
tri 30779 27153 30787 27161 ne
rect 30787 27153 31055 27161
tri 31055 27153 31063 27161 sw
tri 30787 27145 30795 27153 ne
rect 30795 27145 31063 27153
tri 31063 27145 31071 27153 sw
tri 30795 27137 30803 27145 ne
rect 30803 27137 31071 27145
tri 31071 27137 31079 27145 sw
tri 30803 27129 30811 27137 ne
rect 30811 27129 31079 27137
tri 31079 27129 31087 27137 sw
tri 30811 27121 30819 27129 ne
rect 30819 27121 31087 27129
tri 31087 27121 31095 27129 sw
tri 30819 27113 30827 27121 ne
rect 30827 27113 31095 27121
tri 31095 27113 31103 27121 sw
tri 30827 27105 30835 27113 ne
rect 30835 27105 31103 27113
tri 31103 27105 31111 27113 sw
tri 30835 27097 30843 27105 ne
rect 30843 27097 31111 27105
tri 31111 27097 31119 27105 sw
tri 30843 27089 30851 27097 ne
rect 30851 27089 31119 27097
tri 31119 27089 31127 27097 sw
tri 30851 27081 30859 27089 ne
rect 30859 27081 31127 27089
tri 31127 27081 31135 27089 sw
tri 30859 27073 30867 27081 ne
rect 30867 27073 31135 27081
tri 31135 27073 31143 27081 sw
tri 30867 27065 30875 27073 ne
rect 30875 27065 31143 27073
tri 31143 27065 31151 27073 sw
tri 30875 27057 30883 27065 ne
rect 30883 27057 31151 27065
tri 31151 27057 31159 27065 sw
tri 30883 27049 30891 27057 ne
rect 30891 27049 31159 27057
tri 31159 27049 31167 27057 sw
tri 30891 27041 30899 27049 ne
rect 30899 27041 31167 27049
tri 31167 27041 31175 27049 sw
tri 30899 27033 30907 27041 ne
rect 30907 27033 31175 27041
tri 31175 27033 31183 27041 sw
tri 30907 27029 30911 27033 ne
rect 30911 27029 31183 27033
tri 30911 27021 30919 27029 ne
rect 30919 27025 31183 27029
tri 31183 27025 31191 27033 sw
rect 30919 27021 31191 27025
tri 30919 27013 30927 27021 ne
rect 30927 27017 31191 27021
tri 31191 27017 31199 27025 sw
rect 30927 27013 31199 27017
tri 30927 27005 30935 27013 ne
rect 30935 27009 31199 27013
tri 31199 27009 31207 27017 sw
rect 30935 27005 31207 27009
tri 30935 26997 30943 27005 ne
rect 30943 27001 31207 27005
tri 31207 27001 31215 27009 sw
rect 30943 26997 31215 27001
tri 30943 26989 30951 26997 ne
rect 30951 26993 31215 26997
tri 31215 26993 31223 27001 sw
rect 30951 26989 31223 26993
tri 30951 26981 30959 26989 ne
rect 30959 26985 31223 26989
tri 31223 26985 31231 26993 sw
rect 30959 26981 31231 26985
tri 30959 26973 30967 26981 ne
rect 30967 26977 31231 26981
tri 31231 26977 31239 26985 sw
rect 30967 26973 31239 26977
tri 30967 26965 30975 26973 ne
rect 30975 26969 31239 26973
tri 31239 26969 31247 26977 sw
rect 30975 26965 31247 26969
tri 30975 26957 30983 26965 ne
rect 30983 26961 31247 26965
tri 31247 26961 31255 26969 sw
rect 30983 26957 31255 26961
tri 30983 26949 30991 26957 ne
rect 30991 26953 31255 26957
tri 31255 26953 31263 26961 sw
rect 30991 26949 31263 26953
tri 30991 26941 30999 26949 ne
rect 30999 26945 31263 26949
tri 31263 26945 31271 26953 sw
rect 30999 26941 31271 26945
tri 30999 26933 31007 26941 ne
rect 31007 26937 31271 26941
tri 31271 26937 31279 26945 sw
rect 31007 26933 31279 26937
tri 31007 26925 31015 26933 ne
rect 31015 26929 31279 26933
tri 31279 26929 31287 26937 sw
rect 31015 26925 31287 26929
tri 31015 26917 31023 26925 ne
rect 31023 26921 31287 26925
tri 31287 26921 31295 26929 sw
rect 31023 26917 31295 26921
tri 31023 26909 31031 26917 ne
rect 31031 26913 31295 26917
tri 31295 26913 31303 26921 sw
rect 31031 26909 31303 26913
tri 31031 26901 31039 26909 ne
rect 31039 26905 31303 26909
tri 31303 26905 31311 26913 sw
rect 31039 26901 31311 26905
tri 31039 26897 31043 26901 ne
rect 31043 26897 31311 26901
tri 31311 26897 31319 26905 sw
tri 31043 26893 31047 26897 ne
rect 31047 26893 31319 26897
tri 31319 26893 31323 26897 sw
tri 31047 26885 31055 26893 ne
rect 31055 26885 31323 26893
tri 31323 26885 31331 26893 sw
tri 31055 26877 31063 26885 ne
rect 31063 26877 31331 26885
tri 31331 26877 31339 26885 sw
tri 31063 26869 31071 26877 ne
rect 31071 26869 31339 26877
tri 31339 26869 31347 26877 sw
tri 31071 26861 31079 26869 ne
rect 31079 26861 31347 26869
tri 31347 26861 31355 26869 sw
tri 31079 26853 31087 26861 ne
rect 31087 26853 31355 26861
tri 31355 26853 31363 26861 sw
tri 31087 26845 31095 26853 ne
rect 31095 26845 31363 26853
tri 31363 26845 31371 26853 sw
tri 31095 26837 31103 26845 ne
rect 31103 26837 31371 26845
tri 31371 26837 31379 26845 sw
tri 31103 26829 31111 26837 ne
rect 31111 26829 31379 26837
tri 31379 26829 31387 26837 sw
tri 31111 26821 31119 26829 ne
rect 31119 26821 31387 26829
tri 31387 26821 31395 26829 sw
tri 31119 26813 31127 26821 ne
rect 31127 26813 31395 26821
tri 31395 26813 31403 26821 sw
tri 31127 26805 31135 26813 ne
rect 31135 26805 31403 26813
tri 31403 26805 31411 26813 sw
tri 31135 26797 31143 26805 ne
rect 31143 26797 31411 26805
tri 31411 26797 31419 26805 sw
tri 31143 26789 31151 26797 ne
rect 31151 26789 31419 26797
tri 31419 26789 31427 26797 sw
tri 31151 26781 31159 26789 ne
rect 31159 26781 31427 26789
tri 31427 26781 31435 26789 sw
tri 31159 26773 31167 26781 ne
rect 31167 26773 31435 26781
tri 31435 26773 31443 26781 sw
tri 31167 26765 31175 26773 ne
rect 31175 26765 31443 26773
tri 31443 26765 31451 26773 sw
tri 31175 26757 31183 26765 ne
rect 31183 26757 31451 26765
tri 31451 26757 31459 26765 sw
tri 31183 26753 31187 26757 ne
rect 31187 26753 31459 26757
tri 31187 26745 31195 26753 ne
rect 31195 26749 31459 26753
tri 31459 26749 31467 26757 sw
rect 31195 26745 31467 26749
tri 31195 26737 31203 26745 ne
rect 31203 26741 31467 26745
tri 31467 26741 31475 26749 sw
rect 31203 26737 31475 26741
tri 31203 26729 31211 26737 ne
rect 31211 26733 31475 26737
tri 31475 26733 31483 26741 sw
rect 31211 26729 31483 26733
tri 31211 26721 31219 26729 ne
rect 31219 26725 31483 26729
tri 31483 26725 31491 26733 sw
rect 31219 26721 31491 26725
tri 31219 26713 31227 26721 ne
rect 31227 26717 31491 26721
tri 31491 26717 31499 26725 sw
rect 31227 26713 31499 26717
tri 31227 26705 31235 26713 ne
rect 31235 26709 31499 26713
tri 31499 26709 31507 26717 sw
rect 31235 26705 31507 26709
tri 31235 26697 31243 26705 ne
rect 31243 26701 31507 26705
tri 31507 26701 31515 26709 sw
rect 31243 26697 31515 26701
tri 31243 26689 31251 26697 ne
rect 31251 26693 31515 26697
tri 31515 26693 31523 26701 sw
rect 31251 26689 31523 26693
tri 31251 26681 31259 26689 ne
rect 31259 26685 31523 26689
tri 31523 26685 31531 26693 sw
rect 31259 26681 31531 26685
tri 31259 26673 31267 26681 ne
rect 31267 26677 31531 26681
tri 31531 26677 31539 26685 sw
rect 31267 26673 31539 26677
tri 31267 26665 31275 26673 ne
rect 31275 26669 31539 26673
tri 31539 26669 31547 26677 sw
rect 31275 26665 31547 26669
tri 31275 26657 31283 26665 ne
rect 31283 26661 31547 26665
tri 31547 26661 31555 26669 sw
rect 31283 26657 31555 26661
tri 31283 26649 31291 26657 ne
rect 31291 26653 31555 26657
tri 31555 26653 31563 26661 sw
rect 31291 26649 31563 26653
tri 31291 26641 31299 26649 ne
rect 31299 26645 31563 26649
tri 31563 26645 31571 26653 sw
rect 31299 26641 31571 26645
tri 31299 26633 31307 26641 ne
rect 31307 26637 31571 26641
tri 31571 26637 31579 26645 sw
rect 31307 26633 31579 26637
tri 31307 26625 31315 26633 ne
rect 31315 26629 31579 26633
tri 31579 26629 31587 26637 sw
rect 31315 26625 31587 26629
tri 31315 26621 31319 26625 ne
rect 31319 26621 31587 26625
tri 31587 26621 31595 26629 sw
tri 31319 26617 31323 26621 ne
rect 31323 26617 31595 26621
tri 31595 26617 31599 26621 sw
tri 31323 26609 31331 26617 ne
rect 31331 26609 31599 26617
tri 31599 26609 31607 26617 sw
tri 31331 26601 31339 26609 ne
rect 31339 26601 31607 26609
tri 31607 26601 31615 26609 sw
tri 31339 26593 31347 26601 ne
rect 31347 26593 31615 26601
tri 31615 26593 31623 26601 sw
tri 31347 26585 31355 26593 ne
rect 31355 26585 31623 26593
tri 31623 26585 31631 26593 sw
tri 31355 26577 31363 26585 ne
rect 31363 26577 31631 26585
tri 31631 26577 31639 26585 sw
tri 31363 26569 31371 26577 ne
rect 31371 26569 31639 26577
tri 31639 26569 31647 26577 sw
tri 31371 26561 31379 26569 ne
rect 31379 26561 31647 26569
tri 31647 26561 31655 26569 sw
tri 31379 26553 31387 26561 ne
rect 31387 26553 31655 26561
tri 31655 26553 31663 26561 sw
tri 31387 26545 31395 26553 ne
rect 31395 26545 31663 26553
tri 31663 26545 31671 26553 sw
tri 31395 26537 31403 26545 ne
rect 31403 26537 31671 26545
tri 31671 26537 31679 26545 sw
tri 31403 26529 31411 26537 ne
rect 31411 26529 31679 26537
tri 31679 26529 31687 26537 sw
tri 31411 26521 31419 26529 ne
rect 31419 26521 31687 26529
tri 31687 26521 31695 26529 sw
tri 31419 26513 31427 26521 ne
rect 31427 26513 31695 26521
tri 31695 26513 31703 26521 sw
tri 31427 26505 31435 26513 ne
rect 31435 26505 31703 26513
tri 31703 26505 31711 26513 sw
tri 31435 26497 31443 26505 ne
rect 31443 26497 31711 26505
tri 31711 26497 31719 26505 sw
tri 31443 26489 31451 26497 ne
rect 31451 26489 31719 26497
tri 31719 26489 31727 26497 sw
tri 31451 26481 31459 26489 ne
rect 31459 26481 31727 26489
tri 31727 26481 31735 26489 sw
tri 31459 26477 31463 26481 ne
rect 31463 26477 31735 26481
tri 31463 26469 31471 26477 ne
rect 31471 26473 31735 26477
tri 31735 26473 31743 26481 sw
rect 31471 26469 31743 26473
tri 31471 26461 31479 26469 ne
rect 31479 26465 31743 26469
tri 31743 26465 31751 26473 sw
rect 31479 26461 31751 26465
tri 31479 26453 31487 26461 ne
rect 31487 26457 31751 26461
tri 31751 26457 31759 26465 sw
rect 31487 26453 31759 26457
tri 31487 26445 31495 26453 ne
rect 31495 26449 31759 26453
tri 31759 26449 31767 26457 sw
rect 31495 26445 31767 26449
tri 31495 26437 31503 26445 ne
rect 31503 26441 31767 26445
tri 31767 26441 31775 26449 sw
rect 31503 26437 31775 26441
tri 31503 26429 31511 26437 ne
rect 31511 26433 31775 26437
tri 31775 26433 31783 26441 sw
rect 31511 26429 31783 26433
tri 31511 26421 31519 26429 ne
rect 31519 26425 31783 26429
tri 31783 26425 31791 26433 sw
rect 31519 26421 31791 26425
tri 31519 26413 31527 26421 ne
rect 31527 26417 31791 26421
tri 31791 26417 31799 26425 sw
rect 31527 26413 31799 26417
tri 31527 26405 31535 26413 ne
rect 31535 26409 31799 26413
tri 31799 26409 31807 26417 sw
rect 31535 26405 31807 26409
tri 31535 26397 31543 26405 ne
rect 31543 26401 31807 26405
tri 31807 26401 31815 26409 sw
rect 31543 26397 31815 26401
tri 31543 26389 31551 26397 ne
rect 31551 26393 31815 26397
tri 31815 26393 31823 26401 sw
rect 31551 26389 31823 26393
tri 31551 26381 31559 26389 ne
rect 31559 26385 31823 26389
tri 31823 26385 31831 26393 sw
rect 31559 26381 31831 26385
tri 31559 26373 31567 26381 ne
rect 31567 26377 31831 26381
tri 31831 26377 31839 26385 sw
rect 31567 26373 31839 26377
tri 31567 26365 31575 26373 ne
rect 31575 26369 31839 26373
tri 31839 26369 31847 26377 sw
rect 31575 26365 31847 26369
tri 31575 26357 31583 26365 ne
rect 31583 26361 31847 26365
tri 31847 26361 31855 26369 sw
rect 31583 26357 31855 26361
tri 31583 26349 31591 26357 ne
rect 31591 26353 31855 26357
tri 31855 26353 31863 26361 sw
rect 31591 26349 31863 26353
tri 31591 26345 31595 26349 ne
rect 31595 26345 31863 26349
tri 31863 26345 31871 26353 sw
tri 31595 26341 31599 26345 ne
rect 31599 26341 31871 26345
tri 31871 26341 31875 26345 sw
tri 31599 26333 31607 26341 ne
rect 31607 26333 31875 26341
tri 31875 26333 31883 26341 sw
tri 31607 26325 31615 26333 ne
rect 31615 26325 31883 26333
tri 31883 26325 31891 26333 sw
tri 31615 26317 31623 26325 ne
rect 31623 26317 31891 26325
tri 31891 26317 31899 26325 sw
tri 31623 26309 31631 26317 ne
rect 31631 26309 31899 26317
tri 31899 26309 31907 26317 sw
tri 31631 26301 31639 26309 ne
rect 31639 26301 31907 26309
tri 31907 26301 31915 26309 sw
tri 31639 26293 31647 26301 ne
rect 31647 26293 31915 26301
tri 31915 26293 31923 26301 sw
tri 31647 26285 31655 26293 ne
rect 31655 26285 31923 26293
tri 31923 26285 31931 26293 sw
tri 31655 26277 31663 26285 ne
rect 31663 26277 31931 26285
tri 31931 26277 31939 26285 sw
tri 31663 26269 31671 26277 ne
rect 31671 26269 31939 26277
tri 31939 26269 31947 26277 sw
tri 31671 26261 31679 26269 ne
rect 31679 26261 31947 26269
tri 31947 26261 31955 26269 sw
tri 31679 26253 31687 26261 ne
rect 31687 26253 31955 26261
tri 31955 26253 31963 26261 sw
tri 31687 26245 31695 26253 ne
rect 31695 26245 31963 26253
tri 31963 26245 31971 26253 sw
tri 31695 26237 31703 26245 ne
rect 31703 26237 31971 26245
tri 31971 26237 31979 26245 sw
tri 31703 26229 31711 26237 ne
rect 31711 26229 31979 26237
tri 31979 26229 31987 26237 sw
tri 31711 26221 31719 26229 ne
rect 31719 26221 31987 26229
tri 31987 26221 31995 26229 sw
tri 31719 26213 31727 26221 ne
rect 31727 26213 31995 26221
tri 31995 26213 32003 26221 sw
tri 31727 26205 31735 26213 ne
rect 31735 26205 32003 26213
tri 32003 26205 32011 26213 sw
tri 31735 26201 31739 26205 ne
rect 31739 26201 32011 26205
tri 31739 26193 31747 26201 ne
rect 31747 26197 32011 26201
tri 32011 26197 32019 26205 sw
rect 31747 26193 32019 26197
tri 31747 26185 31755 26193 ne
rect 31755 26189 32019 26193
tri 32019 26189 32027 26197 sw
rect 31755 26185 32027 26189
tri 31755 26177 31763 26185 ne
rect 31763 26181 32027 26185
tri 32027 26181 32035 26189 sw
rect 31763 26177 32035 26181
tri 31763 26169 31771 26177 ne
rect 31771 26173 32035 26177
tri 32035 26173 32043 26181 sw
rect 31771 26169 32043 26173
tri 31771 26161 31779 26169 ne
rect 31779 26165 32043 26169
tri 32043 26165 32051 26173 sw
rect 31779 26161 32051 26165
tri 31779 26153 31787 26161 ne
rect 31787 26157 32051 26161
tri 32051 26157 32059 26165 sw
rect 31787 26153 32059 26157
tri 31787 26145 31795 26153 ne
rect 31795 26149 32059 26153
tri 32059 26149 32067 26157 sw
rect 31795 26145 32067 26149
tri 31795 26137 31803 26145 ne
rect 31803 26141 32067 26145
tri 32067 26141 32075 26149 sw
rect 31803 26137 32075 26141
tri 31803 26129 31811 26137 ne
rect 31811 26133 32075 26137
tri 32075 26133 32083 26141 sw
rect 31811 26129 32083 26133
tri 31811 26121 31819 26129 ne
rect 31819 26125 32083 26129
tri 32083 26125 32091 26133 sw
rect 31819 26121 32091 26125
tri 31819 26113 31827 26121 ne
rect 31827 26117 32091 26121
tri 32091 26117 32099 26125 sw
rect 31827 26113 32099 26117
tri 31827 26105 31835 26113 ne
rect 31835 26109 32099 26113
tri 32099 26109 32107 26117 sw
rect 31835 26105 32107 26109
tri 31835 26097 31843 26105 ne
rect 31843 26101 32107 26105
tri 32107 26101 32115 26109 sw
rect 31843 26097 32115 26101
tri 31843 26089 31851 26097 ne
rect 31851 26093 32115 26097
tri 32115 26093 32123 26101 sw
rect 31851 26089 32123 26093
tri 31851 26081 31859 26089 ne
rect 31859 26085 32123 26089
tri 32123 26085 32131 26093 sw
rect 31859 26081 32131 26085
tri 31859 26073 31867 26081 ne
rect 31867 26077 32131 26081
tri 32131 26077 32139 26085 sw
rect 31867 26073 32139 26077
tri 31867 26069 31871 26073 ne
rect 31871 26069 32139 26073
tri 32139 26069 32147 26077 sw
tri 31871 26065 31875 26069 ne
rect 31875 26065 32147 26069
tri 32147 26065 32151 26069 sw
tri 31875 26057 31883 26065 ne
rect 31883 26057 32151 26065
tri 32151 26057 32159 26065 sw
tri 31883 26049 31891 26057 ne
rect 31891 26049 32159 26057
tri 32159 26049 32167 26057 sw
tri 31891 26041 31899 26049 ne
rect 31899 26041 32167 26049
tri 32167 26041 32175 26049 sw
tri 31899 26033 31907 26041 ne
rect 31907 26033 32175 26041
tri 32175 26033 32183 26041 sw
tri 31907 26025 31915 26033 ne
rect 31915 26025 32183 26033
tri 32183 26025 32191 26033 sw
tri 31915 26017 31923 26025 ne
rect 31923 26017 32191 26025
tri 32191 26017 32199 26025 sw
tri 31923 26009 31931 26017 ne
rect 31931 26009 32199 26017
tri 32199 26009 32207 26017 sw
tri 31931 26001 31939 26009 ne
rect 31939 26001 32207 26009
tri 32207 26001 32215 26009 sw
tri 31939 25993 31947 26001 ne
rect 31947 25993 32215 26001
tri 32215 25993 32223 26001 sw
tri 31947 25985 31955 25993 ne
rect 31955 25985 32223 25993
tri 32223 25985 32231 25993 sw
tri 31955 25977 31963 25985 ne
rect 31963 25977 32231 25985
tri 32231 25977 32239 25985 sw
tri 31963 25969 31971 25977 ne
rect 31971 25969 32239 25977
tri 32239 25969 32247 25977 sw
tri 31971 25961 31979 25969 ne
rect 31979 25961 32247 25969
tri 32247 25961 32255 25969 sw
tri 31979 25953 31987 25961 ne
rect 31987 25953 32255 25961
tri 32255 25953 32263 25961 sw
tri 31987 25945 31995 25953 ne
rect 31995 25945 32263 25953
tri 32263 25945 32271 25953 sw
tri 31995 25937 32003 25945 ne
rect 32003 25937 32271 25945
tri 32271 25937 32279 25945 sw
tri 32003 25929 32011 25937 ne
rect 32011 25929 32279 25937
tri 32279 25929 32287 25937 sw
tri 32011 25925 32015 25929 ne
rect 32015 25925 32287 25929
tri 32015 25917 32023 25925 ne
rect 32023 25921 32287 25925
tri 32287 25921 32295 25929 sw
rect 32023 25917 32295 25921
tri 32023 25909 32031 25917 ne
rect 32031 25913 32295 25917
tri 32295 25913 32303 25921 sw
rect 32031 25909 32303 25913
tri 32031 25901 32039 25909 ne
rect 32039 25905 32303 25909
tri 32303 25905 32311 25913 sw
rect 32039 25901 32311 25905
tri 32039 25893 32047 25901 ne
rect 32047 25897 32311 25901
tri 32311 25897 32319 25905 sw
rect 32047 25893 32319 25897
tri 32047 25885 32055 25893 ne
rect 32055 25889 32319 25893
tri 32319 25889 32327 25897 sw
rect 32055 25885 32327 25889
tri 32055 25877 32063 25885 ne
rect 32063 25881 32327 25885
tri 32327 25881 32335 25889 sw
rect 32063 25877 32335 25881
tri 32063 25869 32071 25877 ne
rect 32071 25873 32335 25877
tri 32335 25873 32343 25881 sw
rect 32071 25869 32343 25873
tri 32071 25861 32079 25869 ne
rect 32079 25865 32343 25869
tri 32343 25865 32351 25873 sw
rect 32079 25861 32351 25865
tri 32079 25853 32087 25861 ne
rect 32087 25857 32351 25861
tri 32351 25857 32359 25865 sw
rect 32087 25853 32359 25857
tri 32087 25845 32095 25853 ne
rect 32095 25849 32359 25853
tri 32359 25849 32367 25857 sw
rect 32095 25845 32367 25849
tri 32095 25837 32103 25845 ne
rect 32103 25841 32367 25845
tri 32367 25841 32375 25849 sw
rect 32103 25837 32375 25841
tri 32103 25829 32111 25837 ne
rect 32111 25833 32375 25837
tri 32375 25833 32383 25841 sw
rect 32111 25829 32383 25833
tri 32111 25821 32119 25829 ne
rect 32119 25825 32383 25829
tri 32383 25825 32391 25833 sw
rect 32119 25821 32391 25825
tri 32119 25813 32127 25821 ne
rect 32127 25817 32391 25821
tri 32391 25817 32399 25825 sw
rect 32127 25813 32399 25817
tri 32127 25805 32135 25813 ne
rect 32135 25809 32399 25813
tri 32399 25809 32407 25817 sw
rect 32135 25805 32407 25809
tri 32135 25797 32143 25805 ne
rect 32143 25801 32407 25805
tri 32407 25801 32415 25809 sw
rect 32143 25797 32415 25801
tri 32143 25793 32147 25797 ne
rect 32147 25793 32415 25797
tri 32415 25793 32423 25801 sw
tri 32147 25789 32151 25793 ne
rect 32151 25789 32423 25793
tri 32423 25789 32427 25793 sw
tri 32151 25781 32159 25789 ne
rect 32159 25781 32427 25789
tri 32427 25781 32435 25789 sw
tri 32159 25773 32167 25781 ne
rect 32167 25773 32435 25781
tri 32435 25773 32443 25781 sw
tri 32167 25765 32175 25773 ne
rect 32175 25765 32443 25773
tri 32443 25765 32451 25773 sw
tri 32175 25757 32183 25765 ne
rect 32183 25757 32451 25765
tri 32451 25757 32459 25765 sw
tri 32183 25749 32191 25757 ne
rect 32191 25749 32459 25757
tri 32459 25749 32467 25757 sw
tri 32191 25741 32199 25749 ne
rect 32199 25741 32467 25749
tri 32467 25741 32475 25749 sw
tri 32199 25733 32207 25741 ne
rect 32207 25733 32475 25741
tri 32475 25733 32483 25741 sw
tri 32207 25725 32215 25733 ne
rect 32215 25725 32483 25733
tri 32483 25725 32491 25733 sw
tri 32215 25717 32223 25725 ne
rect 32223 25717 32491 25725
tri 32491 25717 32499 25725 sw
tri 32223 25709 32231 25717 ne
rect 32231 25709 32499 25717
tri 32499 25709 32507 25717 sw
tri 32231 25701 32239 25709 ne
rect 32239 25701 32507 25709
tri 32507 25701 32515 25709 sw
tri 32239 25693 32247 25701 ne
rect 32247 25693 32515 25701
tri 32515 25693 32523 25701 sw
tri 32247 25685 32255 25693 ne
rect 32255 25685 32523 25693
tri 32523 25685 32531 25693 sw
tri 32255 25677 32263 25685 ne
rect 32263 25677 32531 25685
tri 32531 25677 32539 25685 sw
tri 32263 25669 32271 25677 ne
rect 32271 25669 32539 25677
tri 32539 25669 32547 25677 sw
tri 32271 25661 32279 25669 ne
rect 32279 25661 32547 25669
tri 32547 25661 32555 25669 sw
tri 32279 25653 32287 25661 ne
rect 32287 25653 32555 25661
tri 32555 25653 32563 25661 sw
tri 32287 25649 32291 25653 ne
rect 32291 25649 32563 25653
tri 32291 25641 32299 25649 ne
rect 32299 25645 32563 25649
tri 32563 25645 32571 25653 sw
rect 32299 25641 32571 25645
tri 32299 25633 32307 25641 ne
rect 32307 25637 32571 25641
tri 32571 25637 32579 25645 sw
rect 32307 25633 32579 25637
tri 32307 25625 32315 25633 ne
rect 32315 25629 32579 25633
tri 32579 25629 32587 25637 sw
rect 32315 25625 32587 25629
tri 32315 25617 32323 25625 ne
rect 32323 25621 32587 25625
tri 32587 25621 32595 25629 sw
rect 32323 25617 32595 25621
tri 32323 25609 32331 25617 ne
rect 32331 25613 32595 25617
tri 32595 25613 32603 25621 sw
rect 32331 25609 32603 25613
tri 32331 25601 32339 25609 ne
rect 32339 25605 32603 25609
tri 32603 25605 32611 25613 sw
rect 32339 25601 32611 25605
tri 32339 25593 32347 25601 ne
rect 32347 25597 32611 25601
tri 32611 25597 32619 25605 sw
rect 32347 25593 32619 25597
tri 32347 25585 32355 25593 ne
rect 32355 25589 32619 25593
tri 32619 25589 32627 25597 sw
rect 32355 25585 32627 25589
tri 32355 25577 32363 25585 ne
rect 32363 25581 32627 25585
tri 32627 25581 32635 25589 sw
rect 32363 25577 32635 25581
tri 32363 25569 32371 25577 ne
rect 32371 25573 32635 25577
tri 32635 25573 32643 25581 sw
rect 32371 25569 32643 25573
tri 32371 25561 32379 25569 ne
rect 32379 25565 32643 25569
tri 32643 25565 32651 25573 sw
rect 32379 25561 32651 25565
tri 32379 25553 32387 25561 ne
rect 32387 25557 32651 25561
tri 32651 25557 32659 25565 sw
rect 32387 25553 32659 25557
tri 32387 25545 32395 25553 ne
rect 32395 25549 32659 25553
tri 32659 25549 32667 25557 sw
rect 32395 25545 32667 25549
tri 32395 25537 32403 25545 ne
rect 32403 25541 32667 25545
tri 32667 25541 32675 25549 sw
rect 32403 25537 32675 25541
tri 32403 25529 32411 25537 ne
rect 32411 25533 32675 25537
tri 32675 25533 32683 25541 sw
rect 32411 25529 32683 25533
tri 32411 25521 32419 25529 ne
rect 32419 25525 32683 25529
tri 32683 25525 32691 25533 sw
rect 32419 25521 32691 25525
tri 32419 25517 32423 25521 ne
rect 32423 25517 32691 25521
tri 32691 25517 32699 25525 sw
tri 32423 25513 32427 25517 ne
rect 32427 25513 32699 25517
tri 32699 25513 32703 25517 sw
tri 32427 25505 32435 25513 ne
rect 32435 25505 32703 25513
tri 32703 25505 32711 25513 sw
tri 32435 25497 32443 25505 ne
rect 32443 25497 32711 25505
tri 32711 25497 32719 25505 sw
tri 32443 25489 32451 25497 ne
rect 32451 25489 32719 25497
tri 32719 25489 32727 25497 sw
tri 32451 25481 32459 25489 ne
rect 32459 25481 32727 25489
tri 32727 25481 32735 25489 sw
tri 32459 25473 32467 25481 ne
rect 32467 25473 32735 25481
tri 32735 25473 32743 25481 sw
tri 32467 25465 32475 25473 ne
rect 32475 25465 32743 25473
tri 32743 25465 32751 25473 sw
tri 32475 25457 32483 25465 ne
rect 32483 25457 32751 25465
tri 32751 25457 32759 25465 sw
tri 32483 25449 32491 25457 ne
rect 32491 25449 32759 25457
tri 32759 25449 32767 25457 sw
tri 32491 25441 32499 25449 ne
rect 32499 25441 32767 25449
tri 32767 25441 32775 25449 sw
tri 32499 25433 32507 25441 ne
rect 32507 25433 32775 25441
tri 32775 25433 32783 25441 sw
tri 32507 25425 32515 25433 ne
rect 32515 25425 32783 25433
tri 32783 25425 32791 25433 sw
tri 32515 25417 32523 25425 ne
rect 32523 25417 32791 25425
tri 32791 25417 32799 25425 sw
tri 32523 25409 32531 25417 ne
rect 32531 25409 32799 25417
tri 32799 25409 32807 25417 sw
tri 32531 25401 32539 25409 ne
rect 32539 25401 32807 25409
tri 32807 25401 32815 25409 sw
tri 32539 25393 32547 25401 ne
rect 32547 25393 32815 25401
tri 32815 25393 32823 25401 sw
tri 32547 25385 32555 25393 ne
rect 32555 25385 32823 25393
tri 32823 25385 32831 25393 sw
tri 32555 25377 32563 25385 ne
rect 32563 25377 32831 25385
tri 32831 25377 32839 25385 sw
tri 32563 25373 32567 25377 ne
rect 32567 25373 32839 25377
tri 32567 25365 32575 25373 ne
rect 32575 25369 32839 25373
tri 32839 25369 32847 25377 sw
rect 32575 25365 32847 25369
tri 32575 25357 32583 25365 ne
rect 32583 25361 32847 25365
tri 32847 25361 32855 25369 sw
rect 32583 25357 32855 25361
tri 32583 25349 32591 25357 ne
rect 32591 25353 32855 25357
tri 32855 25353 32863 25361 sw
rect 32591 25349 32863 25353
tri 32591 25341 32599 25349 ne
rect 32599 25345 32863 25349
tri 32863 25345 32871 25353 sw
rect 32599 25341 32871 25345
tri 32599 25333 32607 25341 ne
rect 32607 25337 32871 25341
tri 32871 25337 32879 25345 sw
rect 32607 25333 32879 25337
tri 32607 25325 32615 25333 ne
rect 32615 25329 32879 25333
tri 32879 25329 32887 25337 sw
rect 32615 25325 32887 25329
tri 32615 25317 32623 25325 ne
rect 32623 25321 32887 25325
tri 32887 25321 32895 25329 sw
rect 32623 25317 32895 25321
tri 32623 25309 32631 25317 ne
rect 32631 25313 32895 25317
tri 32895 25313 32903 25321 sw
rect 32631 25309 32903 25313
tri 32631 25301 32639 25309 ne
rect 32639 25305 32903 25309
tri 32903 25305 32911 25313 sw
rect 32639 25301 32911 25305
tri 32639 25293 32647 25301 ne
rect 32647 25297 32911 25301
tri 32911 25297 32919 25305 sw
rect 32647 25293 32919 25297
tri 32647 25285 32655 25293 ne
rect 32655 25289 32919 25293
tri 32919 25289 32927 25297 sw
rect 32655 25285 32927 25289
tri 32655 25277 32663 25285 ne
rect 32663 25281 32927 25285
tri 32927 25281 32935 25289 sw
rect 32663 25277 32935 25281
tri 32663 25269 32671 25277 ne
rect 32671 25273 32935 25277
tri 32935 25273 32943 25281 sw
rect 32671 25269 32943 25273
tri 32671 25261 32679 25269 ne
rect 32679 25265 32943 25269
tri 32943 25265 32951 25273 sw
rect 32679 25261 32951 25265
tri 32679 25253 32687 25261 ne
rect 32687 25257 32951 25261
tri 32951 25257 32959 25265 sw
rect 32687 25253 32959 25257
tri 32687 25245 32695 25253 ne
rect 32695 25249 32959 25253
tri 32959 25249 32967 25257 sw
rect 32695 25245 32967 25249
tri 32695 25241 32699 25245 ne
rect 32699 25241 32967 25245
tri 32967 25241 32975 25249 sw
tri 32699 25237 32703 25241 ne
rect 32703 25237 32975 25241
tri 32975 25237 32979 25241 sw
tri 32703 25229 32711 25237 ne
rect 32711 25229 32979 25237
tri 32979 25229 32987 25237 sw
tri 32711 25221 32719 25229 ne
rect 32719 25221 32987 25229
tri 32987 25221 32995 25229 sw
tri 32719 25213 32727 25221 ne
rect 32727 25213 32995 25221
tri 32995 25213 33003 25221 sw
tri 32727 25205 32735 25213 ne
rect 32735 25205 33003 25213
tri 33003 25205 33011 25213 sw
tri 32735 25197 32743 25205 ne
rect 32743 25197 33011 25205
tri 33011 25197 33019 25205 sw
tri 32743 25189 32751 25197 ne
rect 32751 25189 33019 25197
tri 33019 25189 33027 25197 sw
tri 32751 25181 32759 25189 ne
rect 32759 25181 33027 25189
tri 33027 25181 33035 25189 sw
tri 32759 25173 32767 25181 ne
rect 32767 25173 33035 25181
tri 33035 25173 33043 25181 sw
tri 32767 25165 32775 25173 ne
rect 32775 25165 33043 25173
tri 33043 25165 33051 25173 sw
tri 32775 25157 32783 25165 ne
rect 32783 25157 33051 25165
tri 33051 25157 33059 25165 sw
tri 32783 25149 32791 25157 ne
rect 32791 25149 33059 25157
tri 33059 25149 33067 25157 sw
tri 32791 25141 32799 25149 ne
rect 32799 25141 33067 25149
tri 33067 25141 33075 25149 sw
tri 32799 25133 32807 25141 ne
rect 32807 25133 33075 25141
tri 33075 25133 33083 25141 sw
tri 32807 25125 32815 25133 ne
rect 32815 25125 33083 25133
tri 33083 25125 33091 25133 sw
tri 32815 25117 32823 25125 ne
rect 32823 25117 33091 25125
tri 33091 25117 33099 25125 sw
tri 32823 25109 32831 25117 ne
rect 32831 25109 33099 25117
tri 33099 25109 33107 25117 sw
tri 32831 25101 32839 25109 ne
rect 32839 25101 33107 25109
tri 33107 25101 33115 25109 sw
tri 32839 25097 32843 25101 ne
rect 32843 25097 33115 25101
tri 32843 25089 32851 25097 ne
rect 32851 25093 33115 25097
tri 33115 25093 33123 25101 sw
rect 32851 25089 33123 25093
tri 32851 25081 32859 25089 ne
rect 32859 25085 33123 25089
tri 33123 25085 33131 25093 sw
rect 32859 25081 33131 25085
tri 32859 25073 32867 25081 ne
rect 32867 25077 33131 25081
tri 33131 25077 33139 25085 sw
rect 32867 25073 33139 25077
tri 32867 25065 32875 25073 ne
rect 32875 25069 33139 25073
tri 33139 25069 33147 25077 sw
rect 32875 25065 33147 25069
tri 32875 25057 32883 25065 ne
rect 32883 25061 33147 25065
tri 33147 25061 33155 25069 sw
rect 32883 25057 33155 25061
tri 32883 25049 32891 25057 ne
rect 32891 25053 33155 25057
tri 33155 25053 33163 25061 sw
rect 32891 25049 33163 25053
tri 32891 25041 32899 25049 ne
rect 32899 25045 33163 25049
tri 33163 25045 33171 25053 sw
rect 32899 25041 33171 25045
tri 32899 25033 32907 25041 ne
rect 32907 25037 33171 25041
tri 33171 25037 33179 25045 sw
rect 32907 25033 33179 25037
tri 32907 25025 32915 25033 ne
rect 32915 25029 33179 25033
tri 33179 25029 33187 25037 sw
rect 32915 25025 33187 25029
tri 32915 25017 32923 25025 ne
rect 32923 25021 33187 25025
tri 33187 25021 33195 25029 sw
rect 32923 25017 33195 25021
tri 32923 25009 32931 25017 ne
rect 32931 25013 33195 25017
tri 33195 25013 33203 25021 sw
rect 32931 25009 33203 25013
tri 32931 25001 32939 25009 ne
rect 32939 25005 33203 25009
tri 33203 25005 33211 25013 sw
rect 32939 25001 33211 25005
tri 32939 24993 32947 25001 ne
rect 32947 24997 33211 25001
tri 33211 24997 33219 25005 sw
rect 32947 24993 33219 24997
tri 32947 24985 32955 24993 ne
rect 32955 24989 33219 24993
tri 33219 24989 33227 24997 sw
rect 32955 24985 33227 24989
tri 32955 24977 32963 24985 ne
rect 32963 24981 33227 24985
tri 33227 24981 33235 24989 sw
rect 32963 24977 33235 24981
tri 32963 24969 32971 24977 ne
rect 32971 24973 33235 24977
tri 33235 24973 33243 24981 sw
rect 32971 24969 33243 24973
tri 32971 24965 32975 24969 ne
rect 32975 24965 33243 24969
tri 33243 24965 33251 24973 sw
tri 32975 24961 32979 24965 ne
rect 32979 24961 33251 24965
tri 33251 24961 33255 24965 sw
tri 32979 24953 32987 24961 ne
rect 32987 24953 33255 24961
tri 33255 24953 33263 24961 sw
tri 32987 24945 32995 24953 ne
rect 32995 24945 33263 24953
tri 33263 24945 33271 24953 sw
tri 32995 24937 33003 24945 ne
rect 33003 24937 33271 24945
tri 33271 24937 33279 24945 sw
tri 33003 24929 33011 24937 ne
rect 33011 24929 33279 24937
tri 33279 24929 33287 24937 sw
tri 33011 24921 33019 24929 ne
rect 33019 24921 33287 24929
tri 33287 24921 33295 24929 sw
tri 33019 24913 33027 24921 ne
rect 33027 24913 33295 24921
tri 33295 24913 33303 24921 sw
tri 33027 24905 33035 24913 ne
rect 33035 24905 33303 24913
tri 33303 24905 33311 24913 sw
tri 33035 24897 33043 24905 ne
rect 33043 24897 33311 24905
tri 33311 24897 33319 24905 sw
tri 33043 24889 33051 24897 ne
rect 33051 24889 33319 24897
tri 33319 24889 33327 24897 sw
tri 33051 24881 33059 24889 ne
rect 33059 24881 33327 24889
tri 33327 24881 33335 24889 sw
tri 33059 24873 33067 24881 ne
rect 33067 24873 33335 24881
tri 33335 24873 33343 24881 sw
tri 33067 24865 33075 24873 ne
rect 33075 24865 33343 24873
tri 33343 24865 33351 24873 sw
tri 33075 24857 33083 24865 ne
rect 33083 24857 33351 24865
tri 33351 24857 33359 24865 sw
tri 33083 24849 33091 24857 ne
rect 33091 24849 33359 24857
tri 33359 24849 33367 24857 sw
tri 33091 24841 33099 24849 ne
rect 33099 24841 33367 24849
tri 33367 24841 33375 24849 sw
tri 33099 24833 33107 24841 ne
rect 33107 24833 33375 24841
tri 33375 24833 33383 24841 sw
tri 33107 24825 33115 24833 ne
rect 33115 24825 33383 24833
tri 33383 24825 33391 24833 sw
tri 33115 24821 33119 24825 ne
rect 33119 24821 33391 24825
tri 33119 24813 33127 24821 ne
rect 33127 24817 33391 24821
tri 33391 24817 33399 24825 sw
rect 33127 24813 33399 24817
tri 33127 24805 33135 24813 ne
rect 33135 24809 33399 24813
tri 33399 24809 33407 24817 sw
rect 33135 24805 33407 24809
tri 33135 24797 33143 24805 ne
rect 33143 24801 33407 24805
tri 33407 24801 33415 24809 sw
rect 33143 24797 33415 24801
tri 33143 24789 33151 24797 ne
rect 33151 24793 33415 24797
tri 33415 24793 33423 24801 sw
rect 33151 24789 33423 24793
tri 33151 24781 33159 24789 ne
rect 33159 24785 33423 24789
tri 33423 24785 33431 24793 sw
rect 33159 24781 33431 24785
tri 33159 24773 33167 24781 ne
rect 33167 24777 33431 24781
tri 33431 24777 33439 24785 sw
rect 33167 24773 33439 24777
tri 33167 24765 33175 24773 ne
rect 33175 24769 33439 24773
tri 33439 24769 33447 24777 sw
rect 33175 24765 33447 24769
tri 33175 24757 33183 24765 ne
rect 33183 24761 33447 24765
tri 33447 24761 33455 24769 sw
rect 33183 24757 33455 24761
tri 33183 24749 33191 24757 ne
rect 33191 24753 33455 24757
tri 33455 24753 33463 24761 sw
rect 33191 24749 33463 24753
tri 33191 24741 33199 24749 ne
rect 33199 24745 33463 24749
tri 33463 24745 33471 24753 sw
rect 33199 24741 33471 24745
tri 33199 24733 33207 24741 ne
rect 33207 24737 33471 24741
tri 33471 24737 33479 24745 sw
rect 33207 24733 33479 24737
tri 33207 24725 33215 24733 ne
rect 33215 24729 33479 24733
tri 33479 24729 33487 24737 sw
rect 33215 24725 33487 24729
tri 33215 24717 33223 24725 ne
rect 33223 24721 33487 24725
tri 33487 24721 33495 24729 sw
rect 33223 24717 33495 24721
tri 33223 24709 33231 24717 ne
rect 33231 24713 33495 24717
tri 33495 24713 33503 24721 sw
rect 33231 24709 33503 24713
tri 33231 24701 33239 24709 ne
rect 33239 24705 33503 24709
tri 33503 24705 33511 24713 sw
rect 33239 24701 33511 24705
tri 33239 24693 33247 24701 ne
rect 33247 24697 33511 24701
tri 33511 24697 33519 24705 sw
rect 33247 24693 33519 24697
tri 33247 24689 33251 24693 ne
rect 33251 24689 33519 24693
tri 33519 24689 33527 24697 sw
tri 33251 24685 33255 24689 ne
rect 33255 24685 33527 24689
tri 33527 24685 33531 24689 sw
tri 33255 24677 33263 24685 ne
rect 33263 24677 33531 24685
tri 33531 24677 33539 24685 sw
tri 33263 24669 33271 24677 ne
rect 33271 24669 33539 24677
tri 33539 24669 33547 24677 sw
tri 33271 24661 33279 24669 ne
rect 33279 24661 33547 24669
tri 33547 24661 33555 24669 sw
tri 33279 24653 33287 24661 ne
rect 33287 24653 33555 24661
tri 33555 24653 33563 24661 sw
tri 33287 24645 33295 24653 ne
rect 33295 24645 33563 24653
tri 33563 24645 33571 24653 sw
tri 33295 24637 33303 24645 ne
rect 33303 24637 33571 24645
tri 33571 24637 33579 24645 sw
tri 33303 24629 33311 24637 ne
rect 33311 24629 33579 24637
tri 33579 24629 33587 24637 sw
tri 33311 24621 33319 24629 ne
rect 33319 24621 33587 24629
tri 33587 24621 33595 24629 sw
tri 33319 24613 33327 24621 ne
rect 33327 24613 33595 24621
tri 33595 24613 33603 24621 sw
tri 33327 24605 33335 24613 ne
rect 33335 24605 33603 24613
tri 33603 24605 33611 24613 sw
tri 33335 24597 33343 24605 ne
rect 33343 24597 33611 24605
tri 33611 24597 33619 24605 sw
tri 33343 24589 33351 24597 ne
rect 33351 24589 33619 24597
tri 33619 24589 33627 24597 sw
tri 33351 24581 33359 24589 ne
rect 33359 24581 33627 24589
tri 33627 24581 33635 24589 sw
tri 33359 24573 33367 24581 ne
rect 33367 24573 33635 24581
tri 33635 24573 33643 24581 sw
tri 33367 24565 33375 24573 ne
rect 33375 24565 33643 24573
tri 33643 24565 33651 24573 sw
tri 33375 24557 33383 24565 ne
rect 33383 24557 33651 24565
tri 33651 24557 33659 24565 sw
tri 33383 24549 33391 24557 ne
rect 33391 24549 33659 24557
tri 33659 24549 33667 24557 sw
tri 33391 24545 33395 24549 ne
rect 33395 24545 33667 24549
tri 33395 24537 33403 24545 ne
rect 33403 24541 33667 24545
tri 33667 24541 33675 24549 sw
rect 33403 24537 33675 24541
tri 33403 24529 33411 24537 ne
rect 33411 24533 33675 24537
tri 33675 24533 33683 24541 sw
rect 33411 24529 33683 24533
tri 33411 24521 33419 24529 ne
rect 33419 24525 33683 24529
tri 33683 24525 33691 24533 sw
rect 33419 24521 33691 24525
tri 33419 24513 33427 24521 ne
rect 33427 24517 33691 24521
tri 33691 24517 33699 24525 sw
rect 33427 24513 33699 24517
tri 33427 24505 33435 24513 ne
rect 33435 24509 33699 24513
tri 33699 24509 33707 24517 sw
rect 33435 24505 33707 24509
tri 33435 24497 33443 24505 ne
rect 33443 24501 33707 24505
tri 33707 24501 33715 24509 sw
rect 33443 24497 33715 24501
tri 33443 24489 33451 24497 ne
rect 33451 24493 33715 24497
tri 33715 24493 33723 24501 sw
rect 33451 24489 33723 24493
tri 33451 24481 33459 24489 ne
rect 33459 24485 33723 24489
tri 33723 24485 33731 24493 sw
rect 33459 24481 33731 24485
tri 33459 24473 33467 24481 ne
rect 33467 24477 33731 24481
tri 33731 24477 33739 24485 sw
rect 33467 24473 33739 24477
tri 33467 24465 33475 24473 ne
rect 33475 24469 33739 24473
tri 33739 24469 33747 24477 sw
rect 33475 24465 33747 24469
tri 33475 24457 33483 24465 ne
rect 33483 24461 33747 24465
tri 33747 24461 33755 24469 sw
rect 33483 24457 33755 24461
tri 33483 24449 33491 24457 ne
rect 33491 24453 33755 24457
tri 33755 24453 33763 24461 sw
rect 33491 24449 33763 24453
tri 33491 24441 33499 24449 ne
rect 33499 24445 33763 24449
tri 33763 24445 33771 24453 sw
rect 33499 24441 33771 24445
tri 33499 24433 33507 24441 ne
rect 33507 24437 33771 24441
tri 33771 24437 33779 24445 sw
rect 33507 24433 33779 24437
tri 33507 24425 33515 24433 ne
rect 33515 24429 33779 24433
tri 33779 24429 33787 24437 sw
rect 33515 24425 33787 24429
tri 33515 24417 33523 24425 ne
rect 33523 24421 33787 24425
tri 33787 24421 33795 24429 sw
rect 33523 24417 33795 24421
tri 33523 24413 33527 24417 ne
rect 33527 24413 33795 24417
tri 33795 24413 33803 24421 sw
tri 33527 24409 33531 24413 ne
rect 33531 24409 33803 24413
tri 33803 24409 33807 24413 sw
tri 33531 24401 33539 24409 ne
rect 33539 24401 33807 24409
tri 33807 24401 33815 24409 sw
tri 33539 24393 33547 24401 ne
rect 33547 24393 33815 24401
tri 33815 24393 33823 24401 sw
tri 33547 24385 33555 24393 ne
rect 33555 24385 33823 24393
tri 33823 24385 33831 24393 sw
tri 33555 24377 33563 24385 ne
rect 33563 24377 33831 24385
tri 33831 24377 33839 24385 sw
tri 33563 24369 33571 24377 ne
rect 33571 24369 33839 24377
tri 33839 24369 33847 24377 sw
tri 33571 24361 33579 24369 ne
rect 33579 24361 33847 24369
tri 33847 24361 33855 24369 sw
tri 33579 24353 33587 24361 ne
rect 33587 24353 33855 24361
tri 33855 24353 33863 24361 sw
tri 33587 24345 33595 24353 ne
rect 33595 24345 33863 24353
tri 33863 24345 33871 24353 sw
tri 33595 24337 33603 24345 ne
rect 33603 24337 33871 24345
tri 33871 24337 33879 24345 sw
tri 33603 24329 33611 24337 ne
rect 33611 24329 33879 24337
tri 33879 24329 33887 24337 sw
tri 33611 24321 33619 24329 ne
rect 33619 24321 33887 24329
tri 33887 24321 33895 24329 sw
tri 33619 24313 33627 24321 ne
rect 33627 24313 33895 24321
tri 33895 24313 33903 24321 sw
tri 33627 24305 33635 24313 ne
rect 33635 24305 33903 24313
tri 33903 24305 33911 24313 sw
tri 33635 24297 33643 24305 ne
rect 33643 24297 33911 24305
tri 33911 24297 33919 24305 sw
tri 33643 24289 33651 24297 ne
rect 33651 24289 33919 24297
tri 33919 24289 33927 24297 sw
tri 33651 24281 33659 24289 ne
rect 33659 24281 33927 24289
tri 33927 24281 33935 24289 sw
tri 33659 24273 33667 24281 ne
rect 33667 24273 33935 24281
tri 33935 24273 33943 24281 sw
tri 33667 24269 33671 24273 ne
rect 33671 24269 33943 24273
tri 33671 24261 33679 24269 ne
rect 33679 24265 33943 24269
tri 33943 24265 33951 24273 sw
rect 33679 24261 33951 24265
tri 33679 24253 33687 24261 ne
rect 33687 24257 33951 24261
tri 33951 24257 33959 24265 sw
rect 33687 24253 33959 24257
tri 33687 24245 33695 24253 ne
rect 33695 24249 33959 24253
tri 33959 24249 33967 24257 sw
rect 33695 24245 33967 24249
tri 33695 24237 33703 24245 ne
rect 33703 24241 33967 24245
tri 33967 24241 33975 24249 sw
rect 33703 24237 33975 24241
tri 33703 24229 33711 24237 ne
rect 33711 24233 33975 24237
tri 33975 24233 33983 24241 sw
rect 33711 24229 33983 24233
tri 33711 24221 33719 24229 ne
rect 33719 24225 33983 24229
tri 33983 24225 33991 24233 sw
rect 33719 24221 33991 24225
tri 33719 24213 33727 24221 ne
rect 33727 24217 33991 24221
tri 33991 24217 33999 24225 sw
rect 33727 24213 33999 24217
tri 33727 24205 33735 24213 ne
rect 33735 24209 33999 24213
tri 33999 24209 34007 24217 sw
rect 33735 24205 34007 24209
tri 33735 24197 33743 24205 ne
rect 33743 24201 34007 24205
tri 34007 24201 34015 24209 sw
rect 33743 24197 34015 24201
tri 33743 24189 33751 24197 ne
rect 33751 24193 34015 24197
tri 34015 24193 34023 24201 sw
rect 33751 24189 34023 24193
tri 33751 24181 33759 24189 ne
rect 33759 24185 34023 24189
tri 34023 24185 34031 24193 sw
rect 33759 24181 34031 24185
tri 33759 24173 33767 24181 ne
rect 33767 24177 34031 24181
tri 34031 24177 34039 24185 sw
rect 33767 24173 34039 24177
tri 33767 24165 33775 24173 ne
rect 33775 24169 34039 24173
tri 34039 24169 34047 24177 sw
rect 33775 24165 34047 24169
tri 33775 24157 33783 24165 ne
rect 33783 24161 34047 24165
tri 34047 24161 34055 24169 sw
rect 33783 24157 34055 24161
tri 33783 24149 33791 24157 ne
rect 33791 24153 34055 24157
tri 34055 24153 34063 24161 sw
rect 33791 24149 34063 24153
tri 33791 24141 33799 24149 ne
rect 33799 24145 34063 24149
tri 34063 24145 34071 24153 sw
rect 33799 24141 34071 24145
tri 33799 24137 33803 24141 ne
rect 33803 24137 34071 24141
tri 34071 24137 34079 24145 sw
tri 33803 24133 33807 24137 ne
rect 33807 24133 34079 24137
tri 34079 24133 34083 24137 sw
tri 33807 24125 33815 24133 ne
rect 33815 24125 34083 24133
tri 34083 24125 34091 24133 sw
tri 33815 24117 33823 24125 ne
rect 33823 24117 34091 24125
tri 34091 24117 34099 24125 sw
tri 33823 24109 33831 24117 ne
rect 33831 24109 34099 24117
tri 34099 24109 34107 24117 sw
tri 33831 24101 33839 24109 ne
rect 33839 24101 34107 24109
tri 34107 24101 34115 24109 sw
tri 33839 24093 33847 24101 ne
rect 33847 24093 34115 24101
tri 34115 24093 34123 24101 sw
tri 33847 24085 33855 24093 ne
rect 33855 24085 34123 24093
tri 34123 24085 34131 24093 sw
tri 33855 24077 33863 24085 ne
rect 33863 24077 34131 24085
tri 34131 24077 34139 24085 sw
tri 33863 24069 33871 24077 ne
rect 33871 24069 34139 24077
tri 34139 24069 34147 24077 sw
tri 33871 24061 33879 24069 ne
rect 33879 24061 34147 24069
tri 34147 24061 34155 24069 sw
tri 33879 24053 33887 24061 ne
rect 33887 24053 34155 24061
tri 34155 24053 34163 24061 sw
tri 33887 24045 33895 24053 ne
rect 33895 24045 34163 24053
tri 34163 24045 34171 24053 sw
tri 33895 24037 33903 24045 ne
rect 33903 24037 34171 24045
tri 34171 24037 34179 24045 sw
tri 33903 24029 33911 24037 ne
rect 33911 24029 34179 24037
tri 34179 24029 34187 24037 sw
tri 33911 24021 33919 24029 ne
rect 33919 24021 34187 24029
tri 34187 24021 34195 24029 sw
tri 33919 24013 33927 24021 ne
rect 33927 24013 34195 24021
tri 34195 24013 34203 24021 sw
tri 33927 24005 33935 24013 ne
rect 33935 24005 34203 24013
tri 34203 24005 34211 24013 sw
tri 33935 23997 33943 24005 ne
rect 33943 23997 34211 24005
tri 34211 23997 34219 24005 sw
tri 33943 23993 33947 23997 ne
rect 33947 23993 34219 23997
tri 33947 23985 33955 23993 ne
rect 33955 23989 34219 23993
tri 34219 23989 34227 23997 sw
rect 33955 23985 34227 23989
tri 33955 23977 33963 23985 ne
rect 33963 23981 34227 23985
tri 34227 23981 34235 23989 sw
rect 33963 23977 34235 23981
tri 33963 23969 33971 23977 ne
rect 33971 23973 34235 23977
tri 34235 23973 34243 23981 sw
rect 33971 23969 34243 23973
tri 33971 23961 33979 23969 ne
rect 33979 23965 34243 23969
tri 34243 23965 34251 23973 sw
rect 33979 23961 34251 23965
tri 33979 23953 33987 23961 ne
rect 33987 23957 34251 23961
tri 34251 23957 34259 23965 sw
rect 33987 23953 34259 23957
tri 33987 23945 33995 23953 ne
rect 33995 23949 34259 23953
tri 34259 23949 34267 23957 sw
rect 33995 23945 34267 23949
tri 33995 23937 34003 23945 ne
rect 34003 23941 34267 23945
tri 34267 23941 34275 23949 sw
rect 34003 23937 34275 23941
tri 34003 23929 34011 23937 ne
rect 34011 23933 34275 23937
tri 34275 23933 34283 23941 sw
rect 34011 23929 34283 23933
tri 34011 23921 34019 23929 ne
rect 34019 23925 34283 23929
tri 34283 23925 34291 23933 sw
rect 34019 23921 34291 23925
tri 34019 23913 34027 23921 ne
rect 34027 23917 34291 23921
tri 34291 23917 34299 23925 sw
rect 34027 23913 34299 23917
tri 34027 23905 34035 23913 ne
rect 34035 23909 34299 23913
tri 34299 23909 34307 23917 sw
rect 34035 23905 34307 23909
tri 34035 23897 34043 23905 ne
rect 34043 23901 34307 23905
tri 34307 23901 34315 23909 sw
rect 34043 23897 34315 23901
tri 34043 23889 34051 23897 ne
rect 34051 23893 34315 23897
tri 34315 23893 34323 23901 sw
rect 34051 23889 34323 23893
tri 34051 23881 34059 23889 ne
rect 34059 23885 34323 23889
tri 34323 23885 34331 23893 sw
rect 34059 23881 34331 23885
tri 34059 23873 34067 23881 ne
rect 34067 23877 34331 23881
tri 34331 23877 34339 23885 sw
rect 34067 23873 34339 23877
tri 34067 23865 34075 23873 ne
rect 34075 23869 34339 23873
tri 34339 23869 34347 23877 sw
rect 34075 23865 34347 23869
tri 34075 23861 34079 23865 ne
rect 34079 23861 34347 23865
tri 34347 23861 34355 23869 sw
tri 34079 23857 34083 23861 ne
rect 34083 23857 34355 23861
tri 34355 23857 34359 23861 sw
tri 34083 23849 34091 23857 ne
rect 34091 23849 34359 23857
tri 34359 23849 34367 23857 sw
tri 34091 23841 34099 23849 ne
rect 34099 23841 34367 23849
tri 34367 23841 34375 23849 sw
tri 34099 23833 34107 23841 ne
rect 34107 23833 34375 23841
tri 34375 23833 34383 23841 sw
tri 34107 23825 34115 23833 ne
rect 34115 23825 34383 23833
tri 34383 23825 34391 23833 sw
tri 34115 23817 34123 23825 ne
rect 34123 23817 34391 23825
tri 34391 23817 34399 23825 sw
tri 34123 23809 34131 23817 ne
rect 34131 23809 34399 23817
tri 34399 23809 34407 23817 sw
tri 34131 23801 34139 23809 ne
rect 34139 23801 34407 23809
tri 34407 23801 34415 23809 sw
tri 34139 23793 34147 23801 ne
rect 34147 23793 34415 23801
tri 34415 23793 34423 23801 sw
tri 34147 23785 34155 23793 ne
rect 34155 23785 34423 23793
tri 34423 23785 34431 23793 sw
tri 34155 23777 34163 23785 ne
rect 34163 23777 34431 23785
tri 34431 23777 34439 23785 sw
tri 34163 23769 34171 23777 ne
rect 34171 23769 34439 23777
tri 34439 23769 34447 23777 sw
tri 34171 23761 34179 23769 ne
rect 34179 23761 34447 23769
tri 34447 23761 34455 23769 sw
tri 34179 23753 34187 23761 ne
rect 34187 23753 34455 23761
tri 34455 23753 34463 23761 sw
tri 34187 23745 34195 23753 ne
rect 34195 23745 34463 23753
tri 34463 23745 34471 23753 sw
tri 34195 23737 34203 23745 ne
rect 34203 23737 34471 23745
tri 34471 23737 34479 23745 sw
tri 34203 23729 34211 23737 ne
rect 34211 23729 34479 23737
tri 34479 23729 34487 23737 sw
tri 34211 23721 34219 23729 ne
rect 34219 23721 34487 23729
tri 34487 23721 34495 23729 sw
tri 34219 23717 34223 23721 ne
rect 34223 23717 34495 23721
tri 34223 23709 34231 23717 ne
rect 34231 23713 34495 23717
tri 34495 23713 34503 23721 sw
rect 34231 23709 34503 23713
tri 34231 23701 34239 23709 ne
rect 34239 23705 34503 23709
tri 34503 23705 34511 23713 sw
rect 34239 23701 34511 23705
tri 34239 23693 34247 23701 ne
rect 34247 23697 34511 23701
tri 34511 23697 34519 23705 sw
rect 34247 23693 34519 23697
tri 34247 23685 34255 23693 ne
rect 34255 23689 34519 23693
tri 34519 23689 34527 23697 sw
rect 34255 23685 34527 23689
tri 34255 23677 34263 23685 ne
rect 34263 23681 34527 23685
tri 34527 23681 34535 23689 sw
rect 34263 23677 34535 23681
tri 34263 23669 34271 23677 ne
rect 34271 23673 34535 23677
tri 34535 23673 34543 23681 sw
rect 34271 23669 34543 23673
tri 34271 23661 34279 23669 ne
rect 34279 23665 34543 23669
tri 34543 23665 34551 23673 sw
rect 34279 23661 34551 23665
tri 34279 23653 34287 23661 ne
rect 34287 23657 34551 23661
tri 34551 23657 34559 23665 sw
rect 34287 23653 34559 23657
tri 34287 23645 34295 23653 ne
rect 34295 23649 34559 23653
tri 34559 23649 34567 23657 sw
rect 34295 23645 34567 23649
tri 34295 23637 34303 23645 ne
rect 34303 23641 34567 23645
tri 34567 23641 34575 23649 sw
rect 34303 23637 34575 23641
tri 34303 23629 34311 23637 ne
rect 34311 23633 34575 23637
tri 34575 23633 34583 23641 sw
rect 34311 23629 34583 23633
tri 34311 23621 34319 23629 ne
rect 34319 23625 34583 23629
tri 34583 23625 34591 23633 sw
rect 34319 23621 34591 23625
tri 34319 23613 34327 23621 ne
rect 34327 23617 34591 23621
tri 34591 23617 34599 23625 sw
rect 34327 23613 34599 23617
tri 34327 23605 34335 23613 ne
rect 34335 23609 34599 23613
tri 34599 23609 34607 23617 sw
rect 34335 23605 34607 23609
tri 34335 23597 34343 23605 ne
rect 34343 23601 34607 23605
tri 34607 23601 34615 23609 sw
rect 34343 23597 34615 23601
tri 34343 23589 34351 23597 ne
rect 34351 23593 34615 23597
tri 34615 23593 34623 23601 sw
rect 34351 23589 34623 23593
tri 34351 23585 34355 23589 ne
rect 34355 23585 34623 23589
tri 34623 23585 34631 23593 sw
tri 34355 23581 34359 23585 ne
rect 34359 23581 34631 23585
tri 34631 23581 34635 23585 sw
tri 34359 23573 34367 23581 ne
rect 34367 23573 34635 23581
tri 34635 23573 34643 23581 sw
tri 34367 23565 34375 23573 ne
rect 34375 23565 34643 23573
tri 34643 23565 34651 23573 sw
tri 34375 23557 34383 23565 ne
rect 34383 23557 34651 23565
tri 34651 23557 34659 23565 sw
tri 34383 23549 34391 23557 ne
rect 34391 23549 34659 23557
tri 34659 23549 34667 23557 sw
tri 34391 23541 34399 23549 ne
rect 34399 23541 34667 23549
tri 34667 23541 34675 23549 sw
tri 34399 23533 34407 23541 ne
rect 34407 23533 34675 23541
tri 34675 23533 34683 23541 sw
tri 34407 23525 34415 23533 ne
rect 34415 23525 34683 23533
tri 34683 23525 34691 23533 sw
tri 34415 23517 34423 23525 ne
rect 34423 23517 34691 23525
tri 34691 23517 34699 23525 sw
tri 34423 23509 34431 23517 ne
rect 34431 23509 34699 23517
tri 34699 23509 34707 23517 sw
tri 34431 23501 34439 23509 ne
rect 34439 23501 34707 23509
tri 34707 23501 34715 23509 sw
tri 34439 23493 34447 23501 ne
rect 34447 23493 34715 23501
tri 34715 23493 34723 23501 sw
tri 34447 23485 34455 23493 ne
rect 34455 23485 34723 23493
tri 34723 23485 34731 23493 sw
tri 34455 23477 34463 23485 ne
rect 34463 23477 34731 23485
tri 34731 23477 34739 23485 sw
tri 34463 23469 34471 23477 ne
rect 34471 23469 34739 23477
tri 34739 23469 34747 23477 sw
tri 34471 23461 34479 23469 ne
rect 34479 23461 34747 23469
tri 34747 23461 34755 23469 sw
tri 34479 23453 34487 23461 ne
rect 34487 23453 34755 23461
tri 34755 23453 34763 23461 sw
tri 34487 23445 34495 23453 ne
rect 34495 23445 34763 23453
tri 34763 23445 34771 23453 sw
tri 34495 23441 34499 23445 ne
rect 34499 23441 34771 23445
tri 34499 23433 34507 23441 ne
rect 34507 23437 34771 23441
tri 34771 23437 34779 23445 sw
rect 34507 23433 34779 23437
tri 34507 23425 34515 23433 ne
rect 34515 23429 34779 23433
tri 34779 23429 34787 23437 sw
rect 34515 23425 34787 23429
tri 34515 23417 34523 23425 ne
rect 34523 23421 34787 23425
tri 34787 23421 34795 23429 sw
rect 34523 23417 34795 23421
tri 34523 23409 34531 23417 ne
rect 34531 23413 34795 23417
tri 34795 23413 34803 23421 sw
rect 34531 23409 34803 23413
tri 34531 23401 34539 23409 ne
rect 34539 23405 34803 23409
tri 34803 23405 34811 23413 sw
rect 34539 23401 34811 23405
tri 34539 23393 34547 23401 ne
rect 34547 23397 34811 23401
tri 34811 23397 34819 23405 sw
rect 34547 23393 34819 23397
tri 34547 23385 34555 23393 ne
rect 34555 23389 34819 23393
tri 34819 23389 34827 23397 sw
rect 34555 23385 34827 23389
tri 34555 23377 34563 23385 ne
rect 34563 23381 34827 23385
tri 34827 23381 34835 23389 sw
rect 34563 23377 34835 23381
tri 34563 23369 34571 23377 ne
rect 34571 23373 34835 23377
tri 34835 23373 34843 23381 sw
rect 34571 23369 34843 23373
tri 34571 23361 34579 23369 ne
rect 34579 23365 34843 23369
tri 34843 23365 34851 23373 sw
rect 34579 23361 34851 23365
tri 34579 23353 34587 23361 ne
rect 34587 23357 34851 23361
tri 34851 23357 34859 23365 sw
rect 34587 23353 34859 23357
tri 34587 23345 34595 23353 ne
rect 34595 23349 34859 23353
tri 34859 23349 34867 23357 sw
rect 34595 23345 34867 23349
tri 34595 23337 34603 23345 ne
rect 34603 23341 34867 23345
tri 34867 23341 34875 23349 sw
rect 34603 23337 34875 23341
tri 34603 23329 34611 23337 ne
rect 34611 23333 34875 23337
tri 34875 23333 34883 23341 sw
rect 34611 23329 34883 23333
tri 34611 23321 34619 23329 ne
rect 34619 23325 34883 23329
tri 34883 23325 34891 23333 sw
rect 34619 23321 34891 23325
tri 34619 23313 34627 23321 ne
rect 34627 23317 34891 23321
tri 34891 23317 34899 23325 sw
rect 34627 23313 34899 23317
tri 34627 23309 34631 23313 ne
rect 34631 23309 34899 23313
tri 34899 23309 34907 23317 sw
tri 34631 23305 34635 23309 ne
rect 34635 23305 34907 23309
tri 34907 23305 34911 23309 sw
tri 34635 23297 34643 23305 ne
rect 34643 23297 34911 23305
tri 34911 23297 34919 23305 sw
tri 34643 23289 34651 23297 ne
rect 34651 23289 34919 23297
tri 34919 23289 34927 23297 sw
tri 34651 23281 34659 23289 ne
rect 34659 23281 34927 23289
tri 34927 23281 34935 23289 sw
tri 34659 23273 34667 23281 ne
rect 34667 23273 34935 23281
tri 34935 23273 34943 23281 sw
tri 34667 23265 34675 23273 ne
rect 34675 23265 34943 23273
tri 34943 23265 34951 23273 sw
tri 34675 23257 34683 23265 ne
rect 34683 23257 34951 23265
tri 34951 23257 34959 23265 sw
tri 34683 23249 34691 23257 ne
rect 34691 23249 34959 23257
tri 34959 23249 34967 23257 sw
tri 34691 23241 34699 23249 ne
rect 34699 23241 34967 23249
tri 34967 23241 34975 23249 sw
tri 34699 23233 34707 23241 ne
rect 34707 23233 34975 23241
tri 34975 23233 34983 23241 sw
tri 34707 23225 34715 23233 ne
rect 34715 23225 34983 23233
tri 34983 23225 34991 23233 sw
tri 34715 23217 34723 23225 ne
rect 34723 23217 34991 23225
tri 34991 23217 34999 23225 sw
tri 34723 23209 34731 23217 ne
rect 34731 23209 34999 23217
tri 34999 23209 35007 23217 sw
tri 34731 23201 34739 23209 ne
rect 34739 23201 35007 23209
tri 35007 23201 35015 23209 sw
tri 34739 23193 34747 23201 ne
rect 34747 23193 35015 23201
tri 35015 23193 35023 23201 sw
tri 34747 23185 34755 23193 ne
rect 34755 23185 35023 23193
tri 35023 23185 35031 23193 sw
tri 34755 23177 34763 23185 ne
rect 34763 23177 35031 23185
tri 35031 23177 35039 23185 sw
tri 34763 23169 34771 23177 ne
rect 34771 23169 35039 23177
tri 35039 23169 35047 23177 sw
tri 34771 23165 34775 23169 ne
rect 34775 23165 35047 23169
tri 34775 23157 34783 23165 ne
rect 34783 23161 35047 23165
tri 35047 23161 35055 23169 sw
rect 34783 23157 35055 23161
tri 34783 23149 34791 23157 ne
rect 34791 23153 35055 23157
tri 35055 23153 35063 23161 sw
rect 34791 23149 35063 23153
tri 34791 23141 34799 23149 ne
rect 34799 23145 35063 23149
tri 35063 23145 35071 23153 sw
rect 34799 23141 35071 23145
tri 34799 23133 34807 23141 ne
rect 34807 23137 35071 23141
tri 35071 23137 35079 23145 sw
rect 34807 23133 35079 23137
tri 34807 23125 34815 23133 ne
rect 34815 23129 35079 23133
tri 35079 23129 35087 23137 sw
rect 34815 23125 35087 23129
tri 34815 23117 34823 23125 ne
rect 34823 23121 35087 23125
tri 35087 23121 35095 23129 sw
rect 34823 23117 35095 23121
tri 34823 23109 34831 23117 ne
rect 34831 23113 35095 23117
tri 35095 23113 35103 23121 sw
rect 34831 23109 35103 23113
tri 34831 23101 34839 23109 ne
rect 34839 23105 35103 23109
tri 35103 23105 35111 23113 sw
rect 34839 23101 35111 23105
tri 34839 23093 34847 23101 ne
rect 34847 23097 35111 23101
tri 35111 23097 35119 23105 sw
rect 34847 23093 35119 23097
tri 34847 23085 34855 23093 ne
rect 34855 23089 35119 23093
tri 35119 23089 35127 23097 sw
rect 34855 23085 35127 23089
tri 34855 23077 34863 23085 ne
rect 34863 23081 35127 23085
tri 35127 23081 35135 23089 sw
rect 34863 23077 35135 23081
tri 34863 23069 34871 23077 ne
rect 34871 23073 35135 23077
tri 35135 23073 35143 23081 sw
rect 34871 23069 35143 23073
tri 34871 23061 34879 23069 ne
rect 34879 23065 35143 23069
tri 35143 23065 35151 23073 sw
rect 34879 23061 35151 23065
tri 34879 23053 34887 23061 ne
rect 34887 23057 35151 23061
tri 35151 23057 35159 23065 sw
rect 34887 23053 35159 23057
tri 34887 23045 34895 23053 ne
rect 34895 23049 35159 23053
tri 35159 23049 35167 23057 sw
rect 34895 23045 35167 23049
tri 34895 23037 34903 23045 ne
rect 34903 23041 35167 23045
tri 35167 23041 35175 23049 sw
rect 34903 23037 35175 23041
tri 34903 23033 34907 23037 ne
rect 34907 23033 35175 23037
tri 35175 23033 35183 23041 sw
tri 34907 23029 34911 23033 ne
rect 34911 23029 35183 23033
tri 35183 23029 35187 23033 sw
tri 34911 23021 34919 23029 ne
rect 34919 23021 35187 23029
tri 35187 23021 35195 23029 sw
tri 34919 23013 34927 23021 ne
rect 34927 23013 35195 23021
tri 35195 23013 35203 23021 sw
tri 34927 23005 34935 23013 ne
rect 34935 23005 35203 23013
tri 35203 23005 35211 23013 sw
tri 34935 22997 34943 23005 ne
rect 34943 22997 35211 23005
tri 35211 22997 35219 23005 sw
tri 34943 22989 34951 22997 ne
rect 34951 22989 35219 22997
tri 35219 22989 35227 22997 sw
tri 34951 22981 34959 22989 ne
rect 34959 22981 35227 22989
tri 35227 22981 35235 22989 sw
tri 34959 22973 34967 22981 ne
rect 34967 22973 35235 22981
tri 35235 22973 35243 22981 sw
tri 34967 22965 34975 22973 ne
rect 34975 22965 35243 22973
tri 35243 22965 35251 22973 sw
tri 34975 22957 34983 22965 ne
rect 34983 22957 35251 22965
tri 35251 22957 35259 22965 sw
tri 34983 22949 34991 22957 ne
rect 34991 22949 35259 22957
tri 35259 22949 35267 22957 sw
tri 34991 22941 34999 22949 ne
rect 34999 22941 35267 22949
tri 35267 22941 35275 22949 sw
tri 34999 22933 35007 22941 ne
rect 35007 22933 35275 22941
tri 35275 22933 35283 22941 sw
tri 35007 22925 35015 22933 ne
rect 35015 22925 35283 22933
tri 35283 22925 35291 22933 sw
tri 35015 22917 35023 22925 ne
rect 35023 22917 35291 22925
tri 35291 22917 35299 22925 sw
tri 35023 22909 35031 22917 ne
rect 35031 22909 35299 22917
tri 35299 22909 35307 22917 sw
tri 35031 22901 35039 22909 ne
rect 35039 22901 35307 22909
tri 35307 22901 35315 22909 sw
tri 35039 22893 35047 22901 ne
rect 35047 22893 35315 22901
tri 35315 22893 35323 22901 sw
tri 35047 22889 35051 22893 ne
rect 35051 22889 35323 22893
tri 35051 22881 35059 22889 ne
rect 35059 22885 35323 22889
tri 35323 22885 35331 22893 sw
rect 35059 22881 35331 22885
tri 35059 22873 35067 22881 ne
rect 35067 22877 35331 22881
tri 35331 22877 35339 22885 sw
rect 35067 22873 35339 22877
tri 35067 22865 35075 22873 ne
rect 35075 22869 35339 22873
tri 35339 22869 35347 22877 sw
rect 35075 22865 35347 22869
tri 35075 22857 35083 22865 ne
rect 35083 22861 35347 22865
tri 35347 22861 35355 22869 sw
rect 35083 22857 35355 22861
tri 35083 22849 35091 22857 ne
rect 35091 22853 35355 22857
tri 35355 22853 35363 22861 sw
rect 35091 22849 35363 22853
tri 35091 22841 35099 22849 ne
rect 35099 22845 35363 22849
tri 35363 22845 35371 22853 sw
rect 35099 22841 35371 22845
tri 35099 22833 35107 22841 ne
rect 35107 22837 35371 22841
tri 35371 22837 35379 22845 sw
rect 35107 22833 35379 22837
tri 35107 22825 35115 22833 ne
rect 35115 22829 35379 22833
tri 35379 22829 35387 22837 sw
rect 35115 22825 35387 22829
tri 35115 22817 35123 22825 ne
rect 35123 22821 35387 22825
tri 35387 22821 35395 22829 sw
rect 35123 22817 35395 22821
tri 35123 22809 35131 22817 ne
rect 35131 22813 35395 22817
tri 35395 22813 35403 22821 sw
rect 35131 22809 35403 22813
tri 35131 22801 35139 22809 ne
rect 35139 22805 35403 22809
tri 35403 22805 35411 22813 sw
rect 35139 22801 35411 22805
tri 35139 22793 35147 22801 ne
rect 35147 22797 35411 22801
tri 35411 22797 35419 22805 sw
rect 35147 22793 35419 22797
tri 35147 22785 35155 22793 ne
rect 35155 22789 35419 22793
tri 35419 22789 35427 22797 sw
rect 35155 22785 35427 22789
tri 35155 22777 35163 22785 ne
rect 35163 22781 35427 22785
tri 35427 22781 35435 22789 sw
rect 35163 22777 35435 22781
tri 35163 22769 35171 22777 ne
rect 35171 22773 35435 22777
tri 35435 22773 35443 22781 sw
rect 35171 22769 35443 22773
tri 35171 22761 35179 22769 ne
rect 35179 22765 35443 22769
tri 35443 22765 35451 22773 sw
rect 35179 22761 35451 22765
tri 35179 22757 35183 22761 ne
rect 35183 22757 35451 22761
tri 35451 22757 35459 22765 sw
tri 35183 22753 35187 22757 ne
rect 35187 22753 35459 22757
tri 35459 22753 35463 22757 sw
tri 35187 22745 35195 22753 ne
rect 35195 22745 35463 22753
tri 35463 22745 35471 22753 sw
tri 35195 22737 35203 22745 ne
rect 35203 22737 35471 22745
tri 35471 22737 35479 22745 sw
tri 35203 22729 35211 22737 ne
rect 35211 22729 35479 22737
tri 35479 22729 35487 22737 sw
tri 35211 22721 35219 22729 ne
rect 35219 22721 35487 22729
tri 35487 22721 35495 22729 sw
tri 35219 22713 35227 22721 ne
rect 35227 22713 35495 22721
tri 35495 22713 35503 22721 sw
tri 35227 22705 35235 22713 ne
rect 35235 22705 35503 22713
tri 35503 22705 35511 22713 sw
tri 35235 22697 35243 22705 ne
rect 35243 22697 35511 22705
tri 35511 22697 35519 22705 sw
tri 35243 22689 35251 22697 ne
rect 35251 22689 35519 22697
tri 35519 22689 35527 22697 sw
tri 35251 22681 35259 22689 ne
rect 35259 22681 35527 22689
tri 35527 22681 35535 22689 sw
tri 35259 22673 35267 22681 ne
rect 35267 22673 35535 22681
tri 35535 22673 35543 22681 sw
tri 35267 22665 35275 22673 ne
rect 35275 22665 35543 22673
tri 35543 22665 35551 22673 sw
tri 35275 22657 35283 22665 ne
rect 35283 22657 35551 22665
tri 35551 22657 35559 22665 sw
tri 35283 22649 35291 22657 ne
rect 35291 22649 35559 22657
tri 35559 22649 35567 22657 sw
tri 35291 22641 35299 22649 ne
rect 35299 22641 35567 22649
tri 35567 22641 35575 22649 sw
tri 35299 22633 35307 22641 ne
rect 35307 22633 35575 22641
tri 35575 22633 35583 22641 sw
tri 35307 22625 35315 22633 ne
rect 35315 22625 35583 22633
tri 35583 22625 35591 22633 sw
tri 35315 22617 35323 22625 ne
rect 35323 22617 35591 22625
tri 35591 22617 35599 22625 sw
tri 35323 22613 35327 22617 ne
rect 35327 22613 35599 22617
tri 35327 22605 35335 22613 ne
rect 35335 22609 35599 22613
tri 35599 22609 35607 22617 sw
rect 35335 22605 35607 22609
tri 35335 22597 35343 22605 ne
rect 35343 22601 35607 22605
tri 35607 22601 35615 22609 sw
rect 35343 22597 35615 22601
tri 35343 22589 35351 22597 ne
rect 35351 22593 35615 22597
tri 35615 22593 35623 22601 sw
rect 35351 22589 35623 22593
tri 35351 22581 35359 22589 ne
rect 35359 22585 35623 22589
tri 35623 22585 35631 22593 sw
rect 35359 22581 35631 22585
tri 35359 22573 35367 22581 ne
rect 35367 22577 35631 22581
tri 35631 22577 35639 22585 sw
rect 35367 22573 35639 22577
tri 35367 22565 35375 22573 ne
rect 35375 22569 35639 22573
tri 35639 22569 35647 22577 sw
rect 35375 22565 35647 22569
tri 35375 22557 35383 22565 ne
rect 35383 22561 35647 22565
tri 35647 22561 35655 22569 sw
rect 35383 22557 35655 22561
tri 35383 22549 35391 22557 ne
rect 35391 22553 35655 22557
tri 35655 22553 35663 22561 sw
rect 35391 22549 35663 22553
tri 35391 22541 35399 22549 ne
rect 35399 22545 35663 22549
tri 35663 22545 35671 22553 sw
rect 35399 22541 35671 22545
tri 35399 22533 35407 22541 ne
rect 35407 22537 35671 22541
tri 35671 22537 35679 22545 sw
rect 35407 22533 35679 22537
tri 35407 22525 35415 22533 ne
rect 35415 22529 35679 22533
tri 35679 22529 35687 22537 sw
rect 35415 22525 35687 22529
tri 35415 22517 35423 22525 ne
rect 35423 22521 35687 22525
tri 35687 22521 35695 22529 sw
rect 35423 22517 35695 22521
tri 35423 22509 35431 22517 ne
rect 35431 22513 35695 22517
tri 35695 22513 35703 22521 sw
rect 35431 22509 35703 22513
tri 35431 22501 35439 22509 ne
rect 35439 22505 35703 22509
tri 35703 22505 35711 22513 sw
rect 35439 22501 35711 22505
tri 35439 22493 35447 22501 ne
rect 35447 22497 35711 22501
tri 35711 22497 35719 22505 sw
rect 35447 22493 35719 22497
tri 35447 22485 35455 22493 ne
rect 35455 22489 35719 22493
tri 35719 22489 35727 22497 sw
rect 35455 22485 35727 22489
tri 35455 22481 35459 22485 ne
rect 35459 22481 35727 22485
tri 35727 22481 35735 22489 sw
tri 35459 22477 35463 22481 ne
rect 35463 22477 35735 22481
tri 35735 22477 35739 22481 sw
tri 35463 22469 35471 22477 ne
rect 35471 22469 35739 22477
tri 35739 22469 35747 22477 sw
tri 35471 22461 35479 22469 ne
rect 35479 22461 35747 22469
tri 35747 22461 35755 22469 sw
tri 35479 22453 35487 22461 ne
rect 35487 22453 35755 22461
tri 35755 22453 35763 22461 sw
tri 35487 22445 35495 22453 ne
rect 35495 22445 35763 22453
tri 35763 22445 35771 22453 sw
tri 35495 22437 35503 22445 ne
rect 35503 22437 35771 22445
tri 35771 22437 35779 22445 sw
tri 35503 22429 35511 22437 ne
rect 35511 22429 35779 22437
tri 35779 22429 35787 22437 sw
tri 35511 22421 35519 22429 ne
rect 35519 22421 35787 22429
tri 35787 22421 35795 22429 sw
tri 35519 22413 35527 22421 ne
rect 35527 22413 35795 22421
tri 35795 22413 35803 22421 sw
tri 35527 22405 35535 22413 ne
rect 35535 22405 35803 22413
tri 35803 22405 35811 22413 sw
tri 35535 22397 35543 22405 ne
rect 35543 22397 35811 22405
tri 35811 22397 35819 22405 sw
tri 35543 22389 35551 22397 ne
rect 35551 22389 35819 22397
tri 35819 22389 35827 22397 sw
tri 35551 22381 35559 22389 ne
rect 35559 22381 35827 22389
tri 35827 22381 35835 22389 sw
tri 35559 22373 35567 22381 ne
rect 35567 22373 35835 22381
tri 35835 22373 35843 22381 sw
tri 35567 22365 35575 22373 ne
rect 35575 22365 35843 22373
tri 35843 22365 35851 22373 sw
tri 35575 22357 35583 22365 ne
rect 35583 22357 35851 22365
tri 35851 22357 35859 22365 sw
tri 35583 22349 35591 22357 ne
rect 35591 22349 35859 22357
tri 35859 22349 35867 22357 sw
tri 35591 22341 35599 22349 ne
rect 35599 22341 35867 22349
tri 35867 22341 35875 22349 sw
tri 35599 22337 35603 22341 ne
rect 35603 22337 35875 22341
tri 35603 22329 35611 22337 ne
rect 35611 22333 35875 22337
tri 35875 22333 35883 22341 sw
rect 35611 22329 35883 22333
tri 35611 22321 35619 22329 ne
rect 35619 22325 35883 22329
tri 35883 22325 35891 22333 sw
rect 35619 22321 35891 22325
tri 35619 22313 35627 22321 ne
rect 35627 22317 35891 22321
tri 35891 22317 35899 22325 sw
rect 35627 22313 35899 22317
tri 35627 22305 35635 22313 ne
rect 35635 22309 35899 22313
tri 35899 22309 35907 22317 sw
rect 35635 22305 35907 22309
tri 35635 22297 35643 22305 ne
rect 35643 22301 35907 22305
tri 35907 22301 35915 22309 sw
rect 35643 22297 35915 22301
tri 35643 22289 35651 22297 ne
rect 35651 22293 35915 22297
tri 35915 22293 35923 22301 sw
rect 35651 22289 35923 22293
tri 35651 22281 35659 22289 ne
rect 35659 22285 35923 22289
tri 35923 22285 35931 22293 sw
rect 35659 22281 35931 22285
tri 35659 22273 35667 22281 ne
rect 35667 22277 35931 22281
tri 35931 22277 35939 22285 sw
rect 35667 22273 35939 22277
tri 35667 22265 35675 22273 ne
rect 35675 22269 35939 22273
tri 35939 22269 35947 22277 sw
rect 35675 22265 35947 22269
tri 35675 22257 35683 22265 ne
rect 35683 22261 35947 22265
tri 35947 22261 35955 22269 sw
rect 35683 22257 35955 22261
tri 35683 22249 35691 22257 ne
rect 35691 22253 35955 22257
tri 35955 22253 35963 22261 sw
rect 35691 22249 35963 22253
tri 35691 22241 35699 22249 ne
rect 35699 22245 35963 22249
tri 35963 22245 35971 22253 sw
rect 35699 22241 35971 22245
tri 35699 22233 35707 22241 ne
rect 35707 22237 35971 22241
tri 35971 22237 35979 22245 sw
rect 35707 22233 35979 22237
tri 35707 22225 35715 22233 ne
rect 35715 22229 35979 22233
tri 35979 22229 35987 22237 sw
rect 35715 22225 35987 22229
tri 35715 22217 35723 22225 ne
rect 35723 22221 35987 22225
tri 35987 22221 35995 22229 sw
rect 35723 22217 35995 22221
tri 35723 22209 35731 22217 ne
rect 35731 22213 35995 22217
tri 35995 22213 36003 22221 sw
rect 35731 22209 36003 22213
tri 35731 22205 35735 22209 ne
rect 35735 22205 36003 22209
tri 36003 22205 36011 22213 sw
tri 35735 22201 35739 22205 ne
rect 35739 22201 36011 22205
tri 36011 22201 36015 22205 sw
tri 35739 22193 35747 22201 ne
rect 35747 22193 36015 22201
tri 36015 22193 36023 22201 sw
tri 35747 22185 35755 22193 ne
rect 35755 22185 36023 22193
tri 36023 22185 36031 22193 sw
tri 35755 22177 35763 22185 ne
rect 35763 22177 36031 22185
tri 36031 22177 36039 22185 sw
tri 35763 22169 35771 22177 ne
rect 35771 22169 36039 22177
tri 36039 22169 36047 22177 sw
tri 35771 22161 35779 22169 ne
rect 35779 22161 36047 22169
tri 36047 22161 36055 22169 sw
tri 35779 22153 35787 22161 ne
rect 35787 22153 36055 22161
tri 36055 22153 36063 22161 sw
tri 35787 22145 35795 22153 ne
rect 35795 22145 36063 22153
tri 36063 22145 36071 22153 sw
tri 35795 22137 35803 22145 ne
rect 35803 22137 36071 22145
tri 36071 22137 36079 22145 sw
tri 35803 22129 35811 22137 ne
rect 35811 22129 36079 22137
tri 36079 22129 36087 22137 sw
tri 35811 22121 35819 22129 ne
rect 35819 22121 36087 22129
tri 36087 22121 36095 22129 sw
tri 35819 22113 35827 22121 ne
rect 35827 22113 36095 22121
tri 36095 22113 36103 22121 sw
tri 35827 22105 35835 22113 ne
rect 35835 22105 36103 22113
tri 36103 22105 36111 22113 sw
tri 35835 22097 35843 22105 ne
rect 35843 22097 36111 22105
tri 36111 22097 36119 22105 sw
tri 35843 22089 35851 22097 ne
rect 35851 22089 36119 22097
tri 36119 22089 36127 22097 sw
tri 35851 22081 35859 22089 ne
rect 35859 22081 36127 22089
tri 36127 22081 36135 22089 sw
tri 35859 22073 35867 22081 ne
rect 35867 22073 36135 22081
tri 36135 22073 36143 22081 sw
tri 35867 22065 35875 22073 ne
rect 35875 22065 36143 22073
tri 36143 22065 36151 22073 sw
tri 35875 22061 35879 22065 ne
rect 35879 22061 36151 22065
tri 35879 22053 35887 22061 ne
rect 35887 22057 36151 22061
tri 36151 22057 36159 22065 sw
rect 35887 22053 36159 22057
tri 35887 22045 35895 22053 ne
rect 35895 22049 36159 22053
tri 36159 22049 36167 22057 sw
rect 35895 22045 36167 22049
tri 35895 22037 35903 22045 ne
rect 35903 22041 36167 22045
tri 36167 22041 36175 22049 sw
rect 35903 22037 36175 22041
tri 35903 22029 35911 22037 ne
rect 35911 22033 36175 22037
tri 36175 22033 36183 22041 sw
rect 35911 22029 36183 22033
tri 35911 22021 35919 22029 ne
rect 35919 22025 36183 22029
tri 36183 22025 36191 22033 sw
rect 35919 22021 36191 22025
tri 35919 22013 35927 22021 ne
rect 35927 22017 36191 22021
tri 36191 22017 36199 22025 sw
rect 35927 22013 36199 22017
tri 35927 22005 35935 22013 ne
rect 35935 22009 36199 22013
tri 36199 22009 36207 22017 sw
rect 35935 22005 36207 22009
tri 35935 21997 35943 22005 ne
rect 35943 22001 36207 22005
tri 36207 22001 36215 22009 sw
rect 35943 21997 36215 22001
tri 35943 21989 35951 21997 ne
rect 35951 21993 36215 21997
tri 36215 21993 36223 22001 sw
rect 35951 21989 36223 21993
tri 35951 21981 35959 21989 ne
rect 35959 21985 36223 21989
tri 36223 21985 36231 21993 sw
rect 35959 21981 36231 21985
tri 35959 21973 35967 21981 ne
rect 35967 21977 36231 21981
tri 36231 21977 36239 21985 sw
rect 35967 21973 36239 21977
tri 35967 21965 35975 21973 ne
rect 35975 21969 36239 21973
tri 36239 21969 36247 21977 sw
rect 35975 21965 36247 21969
tri 35975 21957 35983 21965 ne
rect 35983 21961 36247 21965
tri 36247 21961 36255 21969 sw
rect 35983 21957 36255 21961
tri 35983 21949 35991 21957 ne
rect 35991 21953 36255 21957
tri 36255 21953 36263 21961 sw
rect 35991 21949 36263 21953
tri 35991 21941 35999 21949 ne
rect 35999 21945 36263 21949
tri 36263 21945 36271 21953 sw
rect 35999 21941 36271 21945
tri 35999 21933 36007 21941 ne
rect 36007 21937 36271 21941
tri 36271 21937 36279 21945 sw
rect 36007 21933 36279 21937
tri 36007 21929 36011 21933 ne
rect 36011 21929 36279 21933
tri 36279 21929 36287 21937 sw
tri 36011 21925 36015 21929 ne
rect 36015 21925 36287 21929
tri 36287 21925 36291 21929 sw
tri 36015 21917 36023 21925 ne
rect 36023 21917 36291 21925
tri 36291 21917 36299 21925 sw
tri 36023 21909 36031 21917 ne
rect 36031 21909 36299 21917
tri 36299 21909 36307 21917 sw
tri 36031 21901 36039 21909 ne
rect 36039 21901 36307 21909
tri 36307 21901 36315 21909 sw
tri 36039 21893 36047 21901 ne
rect 36047 21893 36315 21901
tri 36315 21893 36323 21901 sw
tri 36047 21885 36055 21893 ne
rect 36055 21885 36323 21893
tri 36323 21885 36331 21893 sw
tri 36055 21877 36063 21885 ne
rect 36063 21877 36331 21885
tri 36331 21877 36339 21885 sw
tri 36063 21869 36071 21877 ne
rect 36071 21869 36339 21877
tri 36339 21869 36347 21877 sw
tri 36071 21861 36079 21869 ne
rect 36079 21861 36347 21869
tri 36347 21861 36355 21869 sw
tri 36079 21853 36087 21861 ne
rect 36087 21853 36355 21861
tri 36355 21853 36363 21861 sw
tri 36087 21845 36095 21853 ne
rect 36095 21845 36363 21853
tri 36363 21845 36371 21853 sw
tri 36095 21837 36103 21845 ne
rect 36103 21837 36371 21845
tri 36371 21837 36379 21845 sw
tri 36103 21829 36111 21837 ne
rect 36111 21829 36379 21837
tri 36379 21829 36387 21837 sw
tri 36111 21821 36119 21829 ne
rect 36119 21821 36387 21829
tri 36387 21821 36395 21829 sw
tri 36119 21813 36127 21821 ne
rect 36127 21813 36395 21821
tri 36395 21813 36403 21821 sw
tri 36127 21805 36135 21813 ne
rect 36135 21805 36403 21813
tri 36403 21805 36411 21813 sw
tri 36135 21797 36143 21805 ne
rect 36143 21797 36411 21805
tri 36411 21797 36419 21805 sw
tri 36143 21789 36151 21797 ne
rect 36151 21789 36419 21797
tri 36419 21789 36427 21797 sw
tri 36151 21785 36155 21789 ne
rect 36155 21785 36427 21789
tri 36155 21777 36163 21785 ne
rect 36163 21781 36427 21785
tri 36427 21781 36435 21789 sw
rect 36163 21777 36435 21781
tri 36163 21769 36171 21777 ne
rect 36171 21773 36435 21777
tri 36435 21773 36443 21781 sw
rect 36171 21769 36443 21773
tri 36171 21761 36179 21769 ne
rect 36179 21765 36443 21769
tri 36443 21765 36451 21773 sw
rect 36179 21761 36451 21765
tri 36179 21753 36187 21761 ne
rect 36187 21757 36451 21761
tri 36451 21757 36459 21765 sw
rect 36187 21753 36459 21757
tri 36187 21745 36195 21753 ne
rect 36195 21749 36459 21753
tri 36459 21749 36467 21757 sw
rect 36195 21745 36467 21749
tri 36195 21737 36203 21745 ne
rect 36203 21741 36467 21745
tri 36467 21741 36475 21749 sw
rect 36203 21737 36475 21741
tri 36203 21729 36211 21737 ne
rect 36211 21733 36475 21737
tri 36475 21733 36483 21741 sw
rect 36211 21729 36483 21733
tri 36211 21721 36219 21729 ne
rect 36219 21725 36483 21729
tri 36483 21725 36491 21733 sw
rect 36219 21721 36491 21725
tri 36219 21713 36227 21721 ne
rect 36227 21717 36491 21721
tri 36491 21717 36499 21725 sw
rect 36227 21713 36499 21717
tri 36227 21705 36235 21713 ne
rect 36235 21709 36499 21713
tri 36499 21709 36507 21717 sw
rect 36235 21705 36507 21709
tri 36235 21697 36243 21705 ne
rect 36243 21701 36507 21705
tri 36507 21701 36515 21709 sw
rect 36243 21697 36515 21701
tri 36243 21689 36251 21697 ne
rect 36251 21693 36515 21697
tri 36515 21693 36523 21701 sw
rect 36251 21689 36523 21693
tri 36251 21681 36259 21689 ne
rect 36259 21685 36523 21689
tri 36523 21685 36531 21693 sw
rect 36259 21681 36531 21685
tri 36259 21673 36267 21681 ne
rect 36267 21677 36531 21681
tri 36531 21677 36539 21685 sw
rect 36267 21673 36539 21677
tri 36267 21665 36275 21673 ne
rect 36275 21669 36539 21673
tri 36539 21669 36547 21677 sw
rect 36275 21665 36547 21669
tri 36275 21657 36283 21665 ne
rect 36283 21661 36547 21665
tri 36547 21661 36555 21669 sw
rect 36283 21657 36555 21661
tri 36283 21653 36287 21657 ne
rect 36287 21653 36555 21657
tri 36555 21653 36563 21661 sw
tri 36287 21649 36291 21653 ne
rect 36291 21649 36563 21653
tri 36563 21649 36567 21653 sw
tri 36291 21641 36299 21649 ne
rect 36299 21641 36567 21649
tri 36567 21641 36575 21649 sw
tri 36299 21633 36307 21641 ne
rect 36307 21633 36575 21641
tri 36575 21633 36583 21641 sw
tri 36307 21625 36315 21633 ne
rect 36315 21625 36583 21633
tri 36583 21625 36591 21633 sw
tri 36315 21617 36323 21625 ne
rect 36323 21617 36591 21625
tri 36591 21617 36599 21625 sw
tri 36323 21609 36331 21617 ne
rect 36331 21609 36599 21617
tri 36599 21609 36607 21617 sw
tri 36331 21601 36339 21609 ne
rect 36339 21601 36607 21609
tri 36607 21601 36615 21609 sw
tri 36339 21593 36347 21601 ne
rect 36347 21593 36615 21601
tri 36615 21593 36623 21601 sw
tri 36347 21585 36355 21593 ne
rect 36355 21585 36623 21593
tri 36623 21585 36631 21593 sw
tri 36355 21577 36363 21585 ne
rect 36363 21577 36631 21585
tri 36631 21577 36639 21585 sw
tri 36363 21569 36371 21577 ne
rect 36371 21569 36639 21577
tri 36639 21569 36647 21577 sw
tri 36371 21561 36379 21569 ne
rect 36379 21561 36647 21569
tri 36647 21561 36655 21569 sw
tri 36379 21553 36387 21561 ne
rect 36387 21553 36655 21561
tri 36655 21553 36663 21561 sw
tri 36387 21545 36395 21553 ne
rect 36395 21545 36663 21553
tri 36663 21545 36671 21553 sw
tri 36395 21537 36403 21545 ne
rect 36403 21537 36671 21545
tri 36671 21537 36679 21545 sw
tri 36403 21529 36411 21537 ne
rect 36411 21529 36679 21537
tri 36679 21529 36687 21537 sw
tri 36411 21521 36419 21529 ne
rect 36419 21521 36687 21529
tri 36687 21521 36695 21529 sw
tri 36419 21513 36427 21521 ne
rect 36427 21513 36695 21521
tri 36695 21513 36703 21521 sw
tri 36427 21509 36431 21513 ne
rect 36431 21509 36703 21513
tri 36431 21501 36439 21509 ne
rect 36439 21505 36703 21509
tri 36703 21505 36711 21513 sw
rect 36439 21501 36711 21505
tri 36439 21493 36447 21501 ne
rect 36447 21497 36711 21501
tri 36711 21497 36719 21505 sw
rect 36447 21493 36719 21497
tri 36447 21485 36455 21493 ne
rect 36455 21489 36719 21493
tri 36719 21489 36727 21497 sw
rect 36455 21485 36727 21489
tri 36455 21477 36463 21485 ne
rect 36463 21481 36727 21485
tri 36727 21481 36735 21489 sw
rect 36463 21477 36735 21481
tri 36463 21469 36471 21477 ne
rect 36471 21473 36735 21477
tri 36735 21473 36743 21481 sw
rect 36471 21469 36743 21473
tri 36471 21461 36479 21469 ne
rect 36479 21465 36743 21469
tri 36743 21465 36751 21473 sw
rect 36479 21461 36751 21465
tri 36479 21453 36487 21461 ne
rect 36487 21457 36751 21461
tri 36751 21457 36759 21465 sw
rect 36487 21453 36759 21457
tri 36487 21445 36495 21453 ne
rect 36495 21449 36759 21453
tri 36759 21449 36767 21457 sw
rect 36495 21445 36767 21449
tri 36495 21437 36503 21445 ne
rect 36503 21441 36767 21445
tri 36767 21441 36775 21449 sw
rect 36503 21437 36775 21441
tri 36503 21429 36511 21437 ne
rect 36511 21433 36775 21437
tri 36775 21433 36783 21441 sw
rect 36511 21429 36783 21433
tri 36511 21421 36519 21429 ne
rect 36519 21425 36783 21429
tri 36783 21425 36791 21433 sw
rect 36519 21421 36791 21425
tri 36519 21413 36527 21421 ne
rect 36527 21417 36791 21421
tri 36791 21417 36799 21425 sw
rect 36527 21413 36799 21417
tri 36527 21405 36535 21413 ne
rect 36535 21409 36799 21413
tri 36799 21409 36807 21417 sw
rect 36535 21405 36807 21409
tri 36535 21397 36543 21405 ne
rect 36543 21401 36807 21405
tri 36807 21401 36815 21409 sw
rect 36543 21397 36815 21401
tri 36543 21389 36551 21397 ne
rect 36551 21393 36815 21397
tri 36815 21393 36823 21401 sw
rect 36551 21389 36823 21393
tri 36551 21381 36559 21389 ne
rect 36559 21385 36823 21389
tri 36823 21385 36831 21393 sw
rect 36559 21381 36831 21385
tri 36559 21377 36563 21381 ne
rect 36563 21377 36831 21381
tri 36831 21377 36839 21385 sw
tri 36563 21373 36567 21377 ne
rect 36567 21373 36839 21377
tri 36839 21373 36843 21377 sw
tri 36567 21365 36575 21373 ne
rect 36575 21365 36843 21373
tri 36843 21365 36851 21373 sw
tri 36575 21357 36583 21365 ne
rect 36583 21357 36851 21365
tri 36851 21357 36859 21365 sw
tri 36583 21349 36591 21357 ne
rect 36591 21349 36859 21357
tri 36859 21349 36867 21357 sw
tri 36591 21341 36599 21349 ne
rect 36599 21341 36867 21349
tri 36867 21341 36875 21349 sw
tri 36599 21333 36607 21341 ne
rect 36607 21333 36875 21341
tri 36875 21333 36883 21341 sw
tri 36607 21325 36615 21333 ne
rect 36615 21325 36883 21333
tri 36883 21325 36891 21333 sw
tri 36615 21317 36623 21325 ne
rect 36623 21317 36891 21325
tri 36891 21317 36899 21325 sw
tri 36623 21309 36631 21317 ne
rect 36631 21309 36899 21317
tri 36899 21309 36907 21317 sw
tri 36631 21301 36639 21309 ne
rect 36639 21301 36907 21309
tri 36907 21301 36915 21309 sw
tri 36639 21293 36647 21301 ne
rect 36647 21293 36915 21301
tri 36915 21293 36923 21301 sw
tri 36647 21285 36655 21293 ne
rect 36655 21285 36923 21293
tri 36923 21285 36931 21293 sw
tri 36655 21277 36663 21285 ne
rect 36663 21277 36931 21285
tri 36931 21277 36939 21285 sw
tri 36663 21269 36671 21277 ne
rect 36671 21269 36939 21277
tri 36939 21269 36947 21277 sw
tri 36671 21261 36679 21269 ne
rect 36679 21261 36947 21269
tri 36947 21261 36955 21269 sw
tri 36679 21253 36687 21261 ne
rect 36687 21253 36955 21261
tri 36955 21253 36963 21261 sw
tri 36687 21245 36695 21253 ne
rect 36695 21245 36963 21253
tri 36963 21245 36971 21253 sw
tri 36695 21237 36703 21245 ne
rect 36703 21237 36971 21245
tri 36971 21237 36979 21245 sw
tri 36703 21233 36707 21237 ne
rect 36707 21233 36979 21237
tri 36707 21225 36715 21233 ne
rect 36715 21229 36979 21233
tri 36979 21229 36987 21237 sw
rect 36715 21225 36987 21229
tri 36715 21217 36723 21225 ne
rect 36723 21221 36987 21225
tri 36987 21221 36995 21229 sw
rect 36723 21217 36995 21221
tri 36723 21209 36731 21217 ne
rect 36731 21213 36995 21217
tri 36995 21213 37003 21221 sw
rect 36731 21209 37003 21213
tri 36731 21201 36739 21209 ne
rect 36739 21205 37003 21209
tri 37003 21205 37011 21213 sw
rect 36739 21201 37011 21205
tri 36739 21193 36747 21201 ne
rect 36747 21197 37011 21201
tri 37011 21197 37019 21205 sw
rect 36747 21193 37019 21197
tri 36747 21185 36755 21193 ne
rect 36755 21189 37019 21193
tri 37019 21189 37027 21197 sw
rect 36755 21185 37027 21189
tri 36755 21177 36763 21185 ne
rect 36763 21181 37027 21185
tri 37027 21181 37035 21189 sw
rect 36763 21177 37035 21181
tri 36763 21169 36771 21177 ne
rect 36771 21173 37035 21177
tri 37035 21173 37043 21181 sw
rect 36771 21169 37043 21173
tri 36771 21161 36779 21169 ne
rect 36779 21165 37043 21169
tri 37043 21165 37051 21173 sw
rect 36779 21161 37051 21165
tri 36779 21153 36787 21161 ne
rect 36787 21157 37051 21161
tri 37051 21157 37059 21165 sw
rect 36787 21153 37059 21157
tri 36787 21145 36795 21153 ne
rect 36795 21149 37059 21153
tri 37059 21149 37067 21157 sw
rect 36795 21145 37067 21149
tri 36795 21137 36803 21145 ne
rect 36803 21141 37067 21145
tri 37067 21141 37075 21149 sw
rect 36803 21137 37075 21141
tri 36803 21129 36811 21137 ne
rect 36811 21133 37075 21137
tri 37075 21133 37083 21141 sw
rect 36811 21129 37083 21133
tri 36811 21121 36819 21129 ne
rect 36819 21125 37083 21129
tri 37083 21125 37091 21133 sw
rect 36819 21121 37091 21125
tri 36819 21113 36827 21121 ne
rect 36827 21117 37091 21121
tri 37091 21117 37099 21125 sw
rect 36827 21113 37099 21117
tri 36827 21105 36835 21113 ne
rect 36835 21109 37099 21113
tri 37099 21109 37107 21117 sw
rect 36835 21105 37107 21109
tri 36835 21101 36839 21105 ne
rect 36839 21101 37107 21105
tri 37107 21101 37115 21109 sw
tri 36839 21097 36843 21101 ne
rect 36843 21097 37115 21101
tri 37115 21097 37119 21101 sw
tri 36843 21089 36851 21097 ne
rect 36851 21089 37119 21097
tri 37119 21089 37127 21097 sw
tri 36851 21081 36859 21089 ne
rect 36859 21081 37127 21089
tri 37127 21081 37135 21089 sw
tri 36859 21073 36867 21081 ne
rect 36867 21073 37135 21081
tri 37135 21073 37143 21081 sw
tri 36867 21065 36875 21073 ne
rect 36875 21065 37143 21073
tri 37143 21065 37151 21073 sw
tri 36875 21057 36883 21065 ne
rect 36883 21057 37151 21065
tri 37151 21057 37159 21065 sw
tri 36883 21049 36891 21057 ne
rect 36891 21049 37159 21057
tri 37159 21049 37167 21057 sw
tri 36891 21041 36899 21049 ne
rect 36899 21041 37167 21049
tri 37167 21041 37175 21049 sw
tri 36899 21033 36907 21041 ne
rect 36907 21033 37175 21041
tri 37175 21033 37183 21041 sw
tri 36907 21025 36915 21033 ne
rect 36915 21025 37183 21033
tri 37183 21025 37191 21033 sw
tri 36915 21017 36923 21025 ne
rect 36923 21017 37191 21025
tri 37191 21017 37199 21025 sw
tri 36923 21009 36931 21017 ne
rect 36931 21009 37199 21017
tri 37199 21009 37207 21017 sw
tri 36931 21001 36939 21009 ne
rect 36939 21001 37207 21009
tri 37207 21001 37215 21009 sw
tri 36939 20993 36947 21001 ne
rect 36947 20993 37215 21001
tri 37215 20993 37223 21001 sw
tri 36947 20985 36955 20993 ne
rect 36955 20985 37223 20993
tri 37223 20985 37231 20993 sw
tri 36955 20977 36963 20985 ne
rect 36963 20977 37231 20985
tri 37231 20977 37239 20985 sw
tri 36963 20969 36971 20977 ne
rect 36971 20969 37239 20977
tri 37239 20969 37247 20977 sw
tri 36971 20961 36979 20969 ne
rect 36979 20961 37247 20969
tri 37247 20961 37255 20969 sw
tri 36979 20957 36983 20961 ne
rect 36983 20957 37255 20961
tri 36983 20949 36991 20957 ne
rect 36991 20953 37255 20957
tri 37255 20953 37263 20961 sw
rect 36991 20949 37263 20953
tri 36991 20941 36999 20949 ne
rect 36999 20945 37263 20949
tri 37263 20945 37271 20953 sw
rect 36999 20941 37271 20945
tri 36999 20933 37007 20941 ne
rect 37007 20937 37271 20941
tri 37271 20937 37279 20945 sw
rect 37007 20933 37279 20937
tri 37007 20925 37015 20933 ne
rect 37015 20929 37279 20933
tri 37279 20929 37287 20937 sw
rect 37015 20925 37287 20929
tri 37015 20917 37023 20925 ne
rect 37023 20921 37287 20925
tri 37287 20921 37295 20929 sw
rect 37023 20917 37295 20921
tri 37023 20909 37031 20917 ne
rect 37031 20913 37295 20917
tri 37295 20913 37303 20921 sw
rect 37031 20909 37303 20913
tri 37031 20901 37039 20909 ne
rect 37039 20905 37303 20909
tri 37303 20905 37311 20913 sw
rect 37039 20901 37311 20905
tri 37039 20893 37047 20901 ne
rect 37047 20897 37311 20901
tri 37311 20897 37319 20905 sw
rect 37047 20893 37319 20897
tri 37047 20885 37055 20893 ne
rect 37055 20889 37319 20893
tri 37319 20889 37327 20897 sw
rect 37055 20885 37327 20889
tri 37055 20877 37063 20885 ne
rect 37063 20881 37327 20885
tri 37327 20881 37335 20889 sw
rect 37063 20877 37335 20881
tri 37063 20869 37071 20877 ne
rect 37071 20873 37335 20877
tri 37335 20873 37343 20881 sw
rect 37071 20869 37343 20873
tri 37071 20861 37079 20869 ne
rect 37079 20865 37343 20869
tri 37343 20865 37351 20873 sw
rect 37079 20861 37351 20865
tri 37079 20853 37087 20861 ne
rect 37087 20857 37351 20861
tri 37351 20857 37359 20865 sw
rect 37087 20853 37359 20857
tri 37087 20845 37095 20853 ne
rect 37095 20849 37359 20853
tri 37359 20849 37367 20857 sw
rect 37095 20845 37367 20849
tri 37095 20837 37103 20845 ne
rect 37103 20841 37367 20845
tri 37367 20841 37375 20849 sw
rect 37103 20837 37375 20841
tri 37103 20829 37111 20837 ne
rect 37111 20833 37375 20837
tri 37375 20833 37383 20841 sw
rect 37111 20829 37383 20833
tri 37111 20825 37115 20829 ne
rect 37115 20825 37383 20829
tri 37383 20825 37391 20833 sw
tri 37115 20821 37119 20825 ne
rect 37119 20821 37391 20825
tri 37391 20821 37395 20825 sw
tri 37119 20813 37127 20821 ne
rect 37127 20813 37395 20821
tri 37395 20813 37403 20821 sw
tri 37127 20805 37135 20813 ne
rect 37135 20805 37403 20813
tri 37403 20805 37411 20813 sw
tri 37135 20797 37143 20805 ne
rect 37143 20797 37411 20805
tri 37411 20797 37419 20805 sw
tri 37143 20789 37151 20797 ne
rect 37151 20789 37419 20797
tri 37419 20789 37427 20797 sw
tri 37151 20781 37159 20789 ne
rect 37159 20781 37427 20789
tri 37427 20781 37435 20789 sw
tri 37159 20773 37167 20781 ne
rect 37167 20773 37435 20781
tri 37435 20773 37443 20781 sw
tri 37167 20765 37175 20773 ne
rect 37175 20765 37443 20773
tri 37443 20765 37451 20773 sw
tri 37175 20757 37183 20765 ne
rect 37183 20757 37451 20765
tri 37451 20757 37459 20765 sw
tri 37183 20749 37191 20757 ne
rect 37191 20749 37459 20757
tri 37459 20749 37467 20757 sw
tri 37191 20741 37199 20749 ne
rect 37199 20741 37467 20749
tri 37467 20741 37475 20749 sw
tri 37199 20733 37207 20741 ne
rect 37207 20733 37475 20741
tri 37475 20733 37483 20741 sw
tri 37207 20725 37215 20733 ne
rect 37215 20725 37483 20733
tri 37483 20725 37491 20733 sw
tri 37215 20717 37223 20725 ne
rect 37223 20717 37491 20725
tri 37491 20717 37499 20725 sw
tri 37223 20709 37231 20717 ne
rect 37231 20709 37499 20717
tri 37499 20709 37507 20717 sw
tri 37231 20701 37239 20709 ne
rect 37239 20701 37507 20709
tri 37507 20701 37515 20709 sw
tri 37239 20693 37247 20701 ne
rect 37247 20693 37515 20701
tri 37515 20693 37523 20701 sw
tri 37247 20685 37255 20693 ne
rect 37255 20685 37523 20693
tri 37523 20685 37531 20693 sw
tri 37255 20681 37259 20685 ne
rect 37259 20681 37531 20685
tri 37259 20673 37267 20681 ne
rect 37267 20677 37531 20681
tri 37531 20677 37539 20685 sw
rect 37267 20673 37539 20677
tri 37267 20665 37275 20673 ne
rect 37275 20669 37539 20673
tri 37539 20669 37547 20677 sw
rect 37275 20665 37547 20669
tri 37275 20657 37283 20665 ne
rect 37283 20661 37547 20665
tri 37547 20661 37555 20669 sw
rect 37283 20657 37555 20661
tri 37283 20649 37291 20657 ne
rect 37291 20653 37555 20657
tri 37555 20653 37563 20661 sw
rect 37291 20649 37563 20653
tri 37291 20641 37299 20649 ne
rect 37299 20645 37563 20649
tri 37563 20645 37571 20653 sw
rect 37299 20641 37571 20645
tri 37299 20633 37307 20641 ne
rect 37307 20637 37571 20641
tri 37571 20637 37579 20645 sw
rect 37307 20633 37579 20637
tri 37307 20625 37315 20633 ne
rect 37315 20629 37579 20633
tri 37579 20629 37587 20637 sw
rect 37315 20625 37587 20629
tri 37315 20617 37323 20625 ne
rect 37323 20621 37587 20625
tri 37587 20621 37595 20629 sw
rect 37323 20617 37595 20621
tri 37323 20609 37331 20617 ne
rect 37331 20613 37595 20617
tri 37595 20613 37603 20621 sw
rect 37331 20609 37603 20613
tri 37331 20601 37339 20609 ne
rect 37339 20605 37603 20609
tri 37603 20605 37611 20613 sw
rect 37339 20601 37611 20605
tri 37339 20593 37347 20601 ne
rect 37347 20597 37611 20601
tri 37611 20597 37619 20605 sw
rect 37347 20593 37619 20597
tri 37347 20585 37355 20593 ne
rect 37355 20589 37619 20593
tri 37619 20589 37627 20597 sw
rect 37355 20585 37627 20589
tri 37355 20577 37363 20585 ne
rect 37363 20581 37627 20585
tri 37627 20581 37635 20589 sw
rect 37363 20577 37635 20581
tri 37363 20569 37371 20577 ne
rect 37371 20573 37635 20577
tri 37635 20573 37643 20581 sw
rect 37371 20569 37643 20573
tri 37371 20561 37379 20569 ne
rect 37379 20565 37643 20569
tri 37643 20565 37651 20573 sw
rect 37379 20561 37651 20565
tri 37379 20553 37387 20561 ne
rect 37387 20557 37651 20561
tri 37651 20557 37659 20565 sw
rect 37387 20553 37659 20557
tri 37387 20549 37391 20553 ne
rect 37391 20549 37659 20553
tri 37659 20549 37667 20557 sw
tri 37391 20545 37395 20549 ne
rect 37395 20545 37667 20549
tri 37667 20545 37671 20549 sw
tri 37395 20537 37403 20545 ne
rect 37403 20537 37671 20545
tri 37671 20537 37679 20545 sw
tri 37403 20529 37411 20537 ne
rect 37411 20529 37679 20537
tri 37679 20529 37687 20537 sw
tri 37411 20521 37419 20529 ne
rect 37419 20521 37687 20529
tri 37687 20521 37695 20529 sw
tri 37419 20513 37427 20521 ne
rect 37427 20513 37695 20521
tri 37695 20513 37703 20521 sw
tri 37427 20505 37435 20513 ne
rect 37435 20505 37703 20513
tri 37703 20505 37711 20513 sw
tri 37435 20497 37443 20505 ne
rect 37443 20497 37711 20505
tri 37711 20497 37719 20505 sw
tri 37443 20489 37451 20497 ne
rect 37451 20489 37719 20497
tri 37719 20489 37727 20497 sw
tri 37451 20481 37459 20489 ne
rect 37459 20481 37727 20489
tri 37727 20481 37735 20489 sw
tri 37459 20473 37467 20481 ne
rect 37467 20473 37735 20481
tri 37735 20473 37743 20481 sw
tri 37467 20465 37475 20473 ne
rect 37475 20465 37743 20473
tri 37743 20465 37751 20473 sw
tri 37475 20457 37483 20465 ne
rect 37483 20457 37751 20465
tri 37751 20457 37759 20465 sw
tri 37483 20449 37491 20457 ne
rect 37491 20449 37759 20457
tri 37759 20449 37767 20457 sw
tri 37491 20441 37499 20449 ne
rect 37499 20441 37767 20449
tri 37767 20441 37775 20449 sw
tri 37499 20433 37507 20441 ne
rect 37507 20433 37775 20441
tri 37775 20433 37783 20441 sw
tri 37507 20425 37515 20433 ne
rect 37515 20425 37783 20433
tri 37783 20425 37791 20433 sw
tri 37515 20417 37523 20425 ne
rect 37523 20417 37791 20425
tri 37791 20417 37799 20425 sw
tri 37523 20409 37531 20417 ne
rect 37531 20409 37799 20417
tri 37799 20409 37807 20417 sw
tri 37531 20405 37535 20409 ne
rect 37535 20405 37807 20409
tri 37535 20397 37543 20405 ne
rect 37543 20401 37807 20405
tri 37807 20401 37815 20409 sw
rect 37543 20397 37815 20401
tri 37543 20389 37551 20397 ne
rect 37551 20393 37815 20397
tri 37815 20393 37823 20401 sw
rect 37551 20389 37823 20393
tri 37551 20381 37559 20389 ne
rect 37559 20385 37823 20389
tri 37823 20385 37831 20393 sw
rect 37559 20381 37831 20385
tri 37559 20373 37567 20381 ne
rect 37567 20377 37831 20381
tri 37831 20377 37839 20385 sw
rect 37567 20373 37839 20377
tri 37567 20365 37575 20373 ne
rect 37575 20369 37839 20373
tri 37839 20369 37847 20377 sw
rect 37575 20365 37847 20369
tri 37575 20357 37583 20365 ne
rect 37583 20361 37847 20365
tri 37847 20361 37855 20369 sw
rect 37583 20357 37855 20361
tri 37583 20349 37591 20357 ne
rect 37591 20353 37855 20357
tri 37855 20353 37863 20361 sw
rect 37591 20349 37863 20353
tri 37591 20341 37599 20349 ne
rect 37599 20345 37863 20349
tri 37863 20345 37871 20353 sw
rect 37599 20341 37871 20345
tri 37599 20333 37607 20341 ne
rect 37607 20337 37871 20341
tri 37871 20337 37879 20345 sw
rect 37607 20333 37879 20337
tri 37607 20325 37615 20333 ne
rect 37615 20329 37879 20333
tri 37879 20329 37887 20337 sw
rect 37615 20325 37887 20329
tri 37615 20317 37623 20325 ne
rect 37623 20321 37887 20325
tri 37887 20321 37895 20329 sw
rect 37623 20317 37895 20321
tri 37623 20309 37631 20317 ne
rect 37631 20313 37895 20317
tri 37895 20313 37903 20321 sw
rect 37631 20309 37903 20313
tri 37631 20301 37639 20309 ne
rect 37639 20305 37903 20309
tri 37903 20305 37911 20313 sw
rect 37639 20301 37911 20305
tri 37639 20293 37647 20301 ne
rect 37647 20297 37911 20301
tri 37911 20297 37919 20305 sw
rect 37647 20293 37919 20297
tri 37647 20285 37655 20293 ne
rect 37655 20289 37919 20293
tri 37919 20289 37927 20297 sw
rect 37655 20285 37927 20289
tri 37655 20277 37663 20285 ne
rect 37663 20281 37927 20285
tri 37927 20281 37935 20289 sw
rect 37663 20277 37935 20281
tri 37663 20273 37667 20277 ne
rect 37667 20273 37935 20277
tri 37935 20273 37943 20281 sw
tri 37667 20269 37671 20273 ne
rect 37671 20269 37943 20273
tri 37943 20269 37947 20273 sw
tri 37671 20261 37679 20269 ne
rect 37679 20261 37947 20269
tri 37947 20261 37955 20269 sw
tri 37679 20253 37687 20261 ne
rect 37687 20253 37955 20261
tri 37955 20253 37963 20261 sw
tri 37687 20245 37695 20253 ne
rect 37695 20245 37963 20253
tri 37963 20245 37971 20253 sw
tri 37695 20237 37703 20245 ne
rect 37703 20237 37971 20245
tri 37971 20237 37979 20245 sw
tri 37703 20229 37711 20237 ne
rect 37711 20229 37979 20237
tri 37979 20229 37987 20237 sw
tri 37711 20221 37719 20229 ne
rect 37719 20221 37987 20229
tri 37987 20221 37995 20229 sw
tri 37719 20213 37727 20221 ne
rect 37727 20213 37995 20221
tri 37995 20213 38003 20221 sw
tri 37727 20205 37735 20213 ne
rect 37735 20205 38003 20213
tri 38003 20205 38011 20213 sw
tri 37735 20197 37743 20205 ne
rect 37743 20197 38011 20205
tri 38011 20197 38019 20205 sw
tri 37743 20189 37751 20197 ne
rect 37751 20189 38019 20197
tri 38019 20189 38027 20197 sw
tri 37751 20181 37759 20189 ne
rect 37759 20181 38027 20189
tri 38027 20181 38035 20189 sw
tri 37759 20173 37767 20181 ne
rect 37767 20173 38035 20181
tri 38035 20173 38043 20181 sw
tri 37767 20165 37775 20173 ne
rect 37775 20165 38043 20173
tri 38043 20165 38051 20173 sw
tri 37775 20157 37783 20165 ne
rect 37783 20157 38051 20165
tri 38051 20157 38059 20165 sw
tri 37783 20149 37791 20157 ne
rect 37791 20149 38059 20157
tri 38059 20149 38067 20157 sw
tri 37791 20141 37799 20149 ne
rect 37799 20141 38067 20149
tri 38067 20141 38075 20149 sw
tri 37799 20133 37807 20141 ne
rect 37807 20133 38075 20141
tri 38075 20133 38083 20141 sw
tri 37807 20129 37811 20133 ne
rect 37811 20129 38083 20133
tri 37811 20121 37819 20129 ne
rect 37819 20125 38083 20129
tri 38083 20125 38091 20133 sw
rect 37819 20121 38091 20125
tri 37819 20113 37827 20121 ne
rect 37827 20117 38091 20121
tri 38091 20117 38099 20125 sw
rect 37827 20113 38099 20117
tri 37827 20105 37835 20113 ne
rect 37835 20109 38099 20113
tri 38099 20109 38107 20117 sw
rect 37835 20105 38107 20109
tri 37835 20097 37843 20105 ne
rect 37843 20101 38107 20105
tri 38107 20101 38115 20109 sw
rect 37843 20097 38115 20101
tri 37843 20089 37851 20097 ne
rect 37851 20093 38115 20097
tri 38115 20093 38123 20101 sw
rect 37851 20089 38123 20093
tri 37851 20081 37859 20089 ne
rect 37859 20085 38123 20089
tri 38123 20085 38131 20093 sw
rect 37859 20081 38131 20085
tri 37859 20073 37867 20081 ne
rect 37867 20077 38131 20081
tri 38131 20077 38139 20085 sw
rect 37867 20073 38139 20077
tri 37867 20065 37875 20073 ne
rect 37875 20069 38139 20073
tri 38139 20069 38147 20077 sw
rect 37875 20065 38147 20069
tri 37875 20057 37883 20065 ne
rect 37883 20061 38147 20065
tri 38147 20061 38155 20069 sw
rect 37883 20057 38155 20061
tri 37883 20049 37891 20057 ne
rect 37891 20053 38155 20057
tri 38155 20053 38163 20061 sw
rect 37891 20049 38163 20053
tri 37891 20041 37899 20049 ne
rect 37899 20045 38163 20049
tri 38163 20045 38171 20053 sw
rect 37899 20041 38171 20045
tri 37899 20033 37907 20041 ne
rect 37907 20037 38171 20041
tri 38171 20037 38179 20045 sw
rect 37907 20033 38179 20037
tri 37907 20025 37915 20033 ne
rect 37915 20029 38179 20033
tri 38179 20029 38187 20037 sw
rect 37915 20025 38187 20029
tri 37915 20017 37923 20025 ne
rect 37923 20021 38187 20025
tri 38187 20021 38195 20029 sw
rect 37923 20017 38195 20021
tri 37923 20009 37931 20017 ne
rect 37931 20013 38195 20017
tri 38195 20013 38203 20021 sw
rect 37931 20009 38203 20013
tri 37931 20001 37939 20009 ne
rect 37939 20005 38203 20009
tri 38203 20005 38211 20013 sw
rect 37939 20001 38211 20005
tri 37939 19997 37943 20001 ne
rect 37943 19997 38211 20001
tri 38211 19997 38219 20005 sw
tri 37943 19993 37947 19997 ne
rect 37947 19993 38219 19997
tri 38219 19993 38223 19997 sw
tri 37947 19985 37955 19993 ne
rect 37955 19985 38223 19993
tri 38223 19985 38231 19993 sw
tri 37955 19977 37963 19985 ne
rect 37963 19977 38231 19985
tri 38231 19977 38239 19985 sw
tri 37963 19969 37971 19977 ne
rect 37971 19969 38239 19977
tri 38239 19969 38247 19977 sw
tri 37971 19961 37979 19969 ne
rect 37979 19961 38247 19969
tri 38247 19961 38255 19969 sw
tri 37979 19953 37987 19961 ne
rect 37987 19953 38255 19961
tri 38255 19953 38263 19961 sw
tri 37987 19945 37995 19953 ne
rect 37995 19945 38263 19953
tri 38263 19945 38271 19953 sw
tri 37995 19937 38003 19945 ne
rect 38003 19937 38271 19945
tri 38271 19937 38279 19945 sw
tri 38003 19929 38011 19937 ne
rect 38011 19929 38279 19937
tri 38279 19929 38287 19937 sw
tri 38011 19921 38019 19929 ne
rect 38019 19921 38287 19929
tri 38287 19921 38295 19929 sw
tri 38019 19913 38027 19921 ne
rect 38027 19913 38295 19921
tri 38295 19913 38303 19921 sw
tri 38027 19905 38035 19913 ne
rect 38035 19905 38303 19913
tri 38303 19905 38311 19913 sw
tri 38035 19897 38043 19905 ne
rect 38043 19897 38311 19905
tri 38311 19897 38319 19905 sw
tri 38043 19889 38051 19897 ne
rect 38051 19889 38319 19897
tri 38319 19889 38327 19897 sw
tri 38051 19881 38059 19889 ne
rect 38059 19881 38327 19889
tri 38327 19881 38335 19889 sw
tri 38059 19873 38067 19881 ne
rect 38067 19873 38335 19881
tri 38335 19873 38343 19881 sw
tri 38067 19865 38075 19873 ne
rect 38075 19865 38343 19873
tri 38343 19865 38351 19873 sw
tri 38075 19857 38083 19865 ne
rect 38083 19857 38351 19865
tri 38351 19857 38359 19865 sw
tri 38083 19853 38087 19857 ne
rect 38087 19853 38359 19857
tri 38087 19845 38095 19853 ne
rect 38095 19849 38359 19853
tri 38359 19849 38367 19857 sw
rect 38095 19845 38367 19849
tri 38095 19837 38103 19845 ne
rect 38103 19841 38367 19845
tri 38367 19841 38375 19849 sw
rect 38103 19837 38375 19841
tri 38103 19829 38111 19837 ne
rect 38111 19833 38375 19837
tri 38375 19833 38383 19841 sw
rect 38111 19829 38383 19833
tri 38111 19821 38119 19829 ne
rect 38119 19825 38383 19829
tri 38383 19825 38391 19833 sw
rect 38119 19821 38391 19825
tri 38119 19813 38127 19821 ne
rect 38127 19817 38391 19821
tri 38391 19817 38399 19825 sw
rect 38127 19813 38399 19817
tri 38127 19805 38135 19813 ne
rect 38135 19809 38399 19813
tri 38399 19809 38407 19817 sw
rect 38135 19805 38407 19809
tri 38135 19797 38143 19805 ne
rect 38143 19801 38407 19805
tri 38407 19801 38415 19809 sw
rect 38143 19797 38415 19801
tri 38143 19789 38151 19797 ne
rect 38151 19793 38415 19797
tri 38415 19793 38423 19801 sw
rect 38151 19789 38423 19793
tri 38151 19781 38159 19789 ne
rect 38159 19785 38423 19789
tri 38423 19785 38431 19793 sw
rect 38159 19781 38431 19785
tri 38159 19773 38167 19781 ne
rect 38167 19777 38431 19781
tri 38431 19777 38439 19785 sw
rect 38167 19773 38439 19777
tri 38167 19765 38175 19773 ne
rect 38175 19769 38439 19773
tri 38439 19769 38447 19777 sw
rect 38175 19765 38447 19769
tri 38175 19757 38183 19765 ne
rect 38183 19761 38447 19765
tri 38447 19761 38455 19769 sw
rect 38183 19757 38455 19761
tri 38183 19749 38191 19757 ne
rect 38191 19753 38455 19757
tri 38455 19753 38463 19761 sw
rect 38191 19749 38463 19753
tri 38191 19741 38199 19749 ne
rect 38199 19745 38463 19749
tri 38463 19745 38471 19753 sw
rect 38199 19741 38471 19745
tri 38199 19733 38207 19741 ne
rect 38207 19737 38471 19741
tri 38471 19737 38479 19745 sw
rect 38207 19733 38479 19737
tri 38207 19725 38215 19733 ne
rect 38215 19729 38479 19733
tri 38479 19729 38487 19737 sw
rect 38215 19725 38487 19729
tri 38215 19721 38219 19725 ne
rect 38219 19721 38487 19725
tri 38487 19721 38495 19729 sw
tri 38219 19717 38223 19721 ne
rect 38223 19717 38495 19721
tri 38495 19717 38499 19721 sw
tri 38223 19709 38231 19717 ne
rect 38231 19709 38499 19717
tri 38499 19709 38507 19717 sw
tri 38231 19701 38239 19709 ne
rect 38239 19701 38507 19709
tri 38507 19701 38515 19709 sw
tri 38239 19693 38247 19701 ne
rect 38247 19693 38515 19701
tri 38515 19693 38523 19701 sw
tri 38247 19685 38255 19693 ne
rect 38255 19685 38523 19693
tri 38523 19685 38531 19693 sw
tri 38255 19677 38263 19685 ne
rect 38263 19677 38531 19685
tri 38531 19677 38539 19685 sw
tri 38263 19669 38271 19677 ne
rect 38271 19669 38539 19677
tri 38539 19669 38547 19677 sw
tri 38271 19661 38279 19669 ne
rect 38279 19661 38547 19669
tri 38547 19661 38555 19669 sw
tri 38279 19653 38287 19661 ne
rect 38287 19653 38555 19661
tri 38555 19653 38563 19661 sw
tri 38287 19645 38295 19653 ne
rect 38295 19645 38563 19653
tri 38563 19645 38571 19653 sw
tri 38295 19637 38303 19645 ne
rect 38303 19637 38571 19645
tri 38571 19637 38579 19645 sw
tri 38303 19629 38311 19637 ne
rect 38311 19629 38579 19637
tri 38579 19629 38587 19637 sw
tri 38311 19621 38319 19629 ne
rect 38319 19621 38587 19629
tri 38587 19621 38595 19629 sw
tri 38319 19613 38327 19621 ne
rect 38327 19613 38595 19621
tri 38595 19613 38603 19621 sw
tri 38327 19605 38335 19613 ne
rect 38335 19605 38603 19613
tri 38603 19605 38611 19613 sw
tri 38335 19597 38343 19605 ne
rect 38343 19597 38611 19605
tri 38611 19597 38619 19605 sw
tri 38343 19589 38351 19597 ne
rect 38351 19589 38619 19597
tri 38619 19589 38627 19597 sw
tri 38351 19581 38359 19589 ne
rect 38359 19581 38627 19589
tri 38627 19581 38635 19589 sw
tri 38359 19577 38363 19581 ne
rect 38363 19577 38635 19581
tri 38363 19569 38371 19577 ne
rect 38371 19573 38635 19577
tri 38635 19573 38643 19581 sw
rect 38371 19569 38643 19573
tri 38371 19561 38379 19569 ne
rect 38379 19565 38643 19569
tri 38643 19565 38651 19573 sw
rect 38379 19561 38651 19565
tri 38379 19553 38387 19561 ne
rect 38387 19557 38651 19561
tri 38651 19557 38659 19565 sw
rect 38387 19553 38659 19557
tri 38387 19545 38395 19553 ne
rect 38395 19549 38659 19553
tri 38659 19549 38667 19557 sw
rect 38395 19545 38667 19549
tri 38395 19537 38403 19545 ne
rect 38403 19541 38667 19545
tri 38667 19541 38675 19549 sw
rect 38403 19537 38675 19541
tri 38403 19529 38411 19537 ne
rect 38411 19533 38675 19537
tri 38675 19533 38683 19541 sw
rect 38411 19529 38683 19533
tri 38411 19521 38419 19529 ne
rect 38419 19525 38683 19529
tri 38683 19525 38691 19533 sw
rect 38419 19521 38691 19525
tri 38419 19513 38427 19521 ne
rect 38427 19517 38691 19521
tri 38691 19517 38699 19525 sw
rect 38427 19513 38699 19517
tri 38427 19505 38435 19513 ne
rect 38435 19509 38699 19513
tri 38699 19509 38707 19517 sw
rect 38435 19505 38707 19509
tri 38435 19497 38443 19505 ne
rect 38443 19501 38707 19505
tri 38707 19501 38715 19509 sw
rect 38443 19497 38715 19501
tri 38443 19489 38451 19497 ne
rect 38451 19493 38715 19497
tri 38715 19493 38723 19501 sw
rect 38451 19489 38723 19493
tri 38451 19481 38459 19489 ne
rect 38459 19485 38723 19489
tri 38723 19485 38731 19493 sw
rect 38459 19481 38731 19485
tri 38459 19473 38467 19481 ne
rect 38467 19477 38731 19481
tri 38731 19477 38739 19485 sw
rect 38467 19473 38739 19477
tri 38467 19465 38475 19473 ne
rect 38475 19469 38739 19473
tri 38739 19469 38747 19477 sw
rect 38475 19465 38747 19469
tri 38475 19457 38483 19465 ne
rect 38483 19461 38747 19465
tri 38747 19461 38755 19469 sw
rect 38483 19457 38755 19461
tri 38483 19449 38491 19457 ne
rect 38491 19453 38755 19457
tri 38755 19453 38763 19461 sw
rect 38491 19449 38763 19453
tri 38491 19445 38495 19449 ne
rect 38495 19445 38763 19449
tri 38763 19445 38771 19453 sw
tri 38495 19441 38499 19445 ne
rect 38499 19441 38771 19445
tri 38771 19441 38775 19445 sw
tri 38499 19433 38507 19441 ne
rect 38507 19433 38775 19441
tri 38775 19433 38783 19441 sw
tri 38507 19425 38515 19433 ne
rect 38515 19425 38783 19433
tri 38783 19425 38791 19433 sw
tri 38515 19417 38523 19425 ne
rect 38523 19417 38791 19425
tri 38791 19417 38799 19425 sw
tri 38523 19409 38531 19417 ne
rect 38531 19409 38799 19417
tri 38799 19409 38807 19417 sw
tri 38531 19401 38539 19409 ne
rect 38539 19401 38807 19409
tri 38807 19401 38815 19409 sw
tri 38539 19393 38547 19401 ne
rect 38547 19393 38815 19401
tri 38815 19393 38823 19401 sw
tri 38547 19385 38555 19393 ne
rect 38555 19385 38823 19393
tri 38823 19385 38831 19393 sw
tri 38555 19377 38563 19385 ne
rect 38563 19377 38831 19385
tri 38831 19377 38839 19385 sw
tri 38563 19369 38571 19377 ne
rect 38571 19369 38839 19377
tri 38839 19369 38847 19377 sw
tri 38571 19361 38579 19369 ne
rect 38579 19361 38847 19369
tri 38847 19361 38855 19369 sw
tri 38579 19353 38587 19361 ne
rect 38587 19353 38855 19361
tri 38855 19353 38863 19361 sw
tri 38587 19345 38595 19353 ne
rect 38595 19345 38863 19353
tri 38863 19345 38871 19353 sw
tri 38595 19337 38603 19345 ne
rect 38603 19337 38871 19345
tri 38871 19337 38879 19345 sw
tri 38603 19329 38611 19337 ne
rect 38611 19329 38879 19337
tri 38879 19329 38887 19337 sw
tri 38611 19321 38619 19329 ne
rect 38619 19321 38887 19329
tri 38887 19321 38895 19329 sw
tri 38619 19313 38627 19321 ne
rect 38627 19313 38895 19321
tri 38895 19313 38903 19321 sw
tri 38627 19305 38635 19313 ne
rect 38635 19305 38903 19313
tri 38903 19305 38911 19313 sw
tri 38635 19301 38639 19305 ne
rect 38639 19301 38911 19305
tri 38639 19293 38647 19301 ne
rect 38647 19297 38911 19301
tri 38911 19297 38919 19305 sw
rect 38647 19293 38919 19297
tri 38647 19285 38655 19293 ne
rect 38655 19289 38919 19293
tri 38919 19289 38927 19297 sw
rect 38655 19285 38927 19289
tri 38655 19277 38663 19285 ne
rect 38663 19281 38927 19285
tri 38927 19281 38935 19289 sw
rect 38663 19277 38935 19281
tri 38663 19269 38671 19277 ne
rect 38671 19273 38935 19277
tri 38935 19273 38943 19281 sw
rect 38671 19269 38943 19273
tri 38671 19261 38679 19269 ne
rect 38679 19265 38943 19269
tri 38943 19265 38951 19273 sw
rect 38679 19261 38951 19265
tri 38679 19253 38687 19261 ne
rect 38687 19257 38951 19261
tri 38951 19257 38959 19265 sw
rect 38687 19253 38959 19257
tri 38687 19245 38695 19253 ne
rect 38695 19249 38959 19253
tri 38959 19249 38967 19257 sw
rect 38695 19245 38967 19249
tri 38695 19237 38703 19245 ne
rect 38703 19241 38967 19245
tri 38967 19241 38975 19249 sw
rect 38703 19237 38975 19241
tri 38703 19229 38711 19237 ne
rect 38711 19233 38975 19237
tri 38975 19233 38983 19241 sw
rect 38711 19229 38983 19233
tri 38711 19221 38719 19229 ne
rect 38719 19225 38983 19229
tri 38983 19225 38991 19233 sw
rect 38719 19221 38991 19225
tri 38719 19213 38727 19221 ne
rect 38727 19217 38991 19221
tri 38991 19217 38999 19225 sw
rect 38727 19213 38999 19217
tri 38727 19205 38735 19213 ne
rect 38735 19209 38999 19213
tri 38999 19209 39007 19217 sw
rect 38735 19205 39007 19209
tri 38735 19197 38743 19205 ne
rect 38743 19201 39007 19205
tri 39007 19201 39015 19209 sw
rect 38743 19197 39015 19201
tri 38743 19189 38751 19197 ne
rect 38751 19193 39015 19197
tri 39015 19193 39023 19201 sw
rect 38751 19189 39023 19193
tri 38751 19181 38759 19189 ne
rect 38759 19185 39023 19189
tri 39023 19185 39031 19193 sw
rect 38759 19181 39031 19185
tri 38759 19173 38767 19181 ne
rect 38767 19177 39031 19181
tri 39031 19177 39039 19185 sw
rect 38767 19173 39039 19177
tri 38767 19169 38771 19173 ne
rect 38771 19169 39039 19173
tri 39039 19169 39047 19177 sw
tri 38771 19165 38775 19169 ne
rect 38775 19165 39047 19169
tri 39047 19165 39051 19169 sw
tri 38775 19157 38783 19165 ne
rect 38783 19157 39051 19165
tri 39051 19157 39059 19165 sw
tri 38783 19149 38791 19157 ne
rect 38791 19149 39059 19157
tri 39059 19149 39067 19157 sw
tri 38791 19141 38799 19149 ne
rect 38799 19141 39067 19149
tri 39067 19141 39075 19149 sw
tri 38799 19133 38807 19141 ne
rect 38807 19133 39075 19141
tri 39075 19133 39083 19141 sw
tri 38807 19125 38815 19133 ne
rect 38815 19125 39083 19133
tri 39083 19125 39091 19133 sw
tri 38815 19117 38823 19125 ne
rect 38823 19117 39091 19125
tri 39091 19117 39099 19125 sw
tri 38823 19109 38831 19117 ne
rect 38831 19109 39099 19117
tri 39099 19109 39107 19117 sw
tri 38831 19101 38839 19109 ne
rect 38839 19101 39107 19109
tri 39107 19101 39115 19109 sw
tri 38839 19093 38847 19101 ne
rect 38847 19093 39115 19101
tri 39115 19093 39123 19101 sw
tri 38847 19085 38855 19093 ne
rect 38855 19085 39123 19093
tri 39123 19085 39131 19093 sw
tri 38855 19077 38863 19085 ne
rect 38863 19077 39131 19085
tri 39131 19077 39139 19085 sw
tri 38863 19069 38871 19077 ne
rect 38871 19069 39139 19077
tri 39139 19069 39147 19077 sw
tri 38871 19061 38879 19069 ne
rect 38879 19061 39147 19069
tri 39147 19061 39155 19069 sw
tri 38879 19053 38887 19061 ne
rect 38887 19053 39155 19061
tri 39155 19053 39163 19061 sw
tri 38887 19045 38895 19053 ne
rect 38895 19045 39163 19053
tri 39163 19045 39171 19053 sw
tri 38895 19037 38903 19045 ne
rect 38903 19037 39171 19045
tri 39171 19037 39179 19045 sw
tri 38903 19029 38911 19037 ne
rect 38911 19029 39179 19037
tri 39179 19029 39187 19037 sw
tri 38911 19025 38915 19029 ne
rect 38915 19025 39187 19029
tri 38915 19017 38923 19025 ne
rect 38923 19021 39187 19025
tri 39187 19021 39195 19029 sw
rect 38923 19017 39195 19021
tri 38923 19009 38931 19017 ne
rect 38931 19013 39195 19017
tri 39195 19013 39203 19021 sw
rect 38931 19009 39203 19013
tri 38931 19001 38939 19009 ne
rect 38939 19005 39203 19009
tri 39203 19005 39211 19013 sw
rect 38939 19001 39211 19005
tri 38939 18993 38947 19001 ne
rect 38947 18997 39211 19001
tri 39211 18997 39219 19005 sw
rect 38947 18993 39219 18997
tri 38947 18985 38955 18993 ne
rect 38955 18989 39219 18993
tri 39219 18989 39227 18997 sw
rect 38955 18985 39227 18989
tri 38955 18977 38963 18985 ne
rect 38963 18981 39227 18985
tri 39227 18981 39235 18989 sw
rect 38963 18977 39235 18981
tri 38963 18969 38971 18977 ne
rect 38971 18973 39235 18977
tri 39235 18973 39243 18981 sw
rect 38971 18969 39243 18973
tri 38971 18961 38979 18969 ne
rect 38979 18965 39243 18969
tri 39243 18965 39251 18973 sw
rect 38979 18961 39251 18965
tri 38979 18953 38987 18961 ne
rect 38987 18957 39251 18961
tri 39251 18957 39259 18965 sw
rect 38987 18953 39259 18957
tri 38987 18945 38995 18953 ne
rect 38995 18949 39259 18953
tri 39259 18949 39267 18957 sw
rect 38995 18945 39267 18949
tri 38995 18937 39003 18945 ne
rect 39003 18941 39267 18945
tri 39267 18941 39275 18949 sw
rect 39003 18937 39275 18941
tri 39003 18929 39011 18937 ne
rect 39011 18933 39275 18937
tri 39275 18933 39283 18941 sw
rect 39011 18929 39283 18933
tri 39011 18921 39019 18929 ne
rect 39019 18925 39283 18929
tri 39283 18925 39291 18933 sw
rect 39019 18921 39291 18925
tri 39019 18913 39027 18921 ne
rect 39027 18917 39291 18921
tri 39291 18917 39299 18925 sw
rect 39027 18913 39299 18917
tri 39027 18905 39035 18913 ne
rect 39035 18909 39299 18913
tri 39299 18909 39307 18917 sw
rect 39035 18905 39307 18909
tri 39035 18897 39043 18905 ne
rect 39043 18901 39307 18905
tri 39307 18901 39315 18909 sw
rect 39043 18897 39315 18901
tri 39043 18893 39047 18897 ne
rect 39047 18893 39315 18897
tri 39315 18893 39323 18901 sw
tri 39047 18889 39051 18893 ne
rect 39051 18889 39323 18893
tri 39323 18889 39327 18893 sw
tri 39051 18881 39059 18889 ne
rect 39059 18881 39327 18889
tri 39327 18881 39335 18889 sw
tri 39059 18873 39067 18881 ne
rect 39067 18873 39335 18881
tri 39335 18873 39343 18881 sw
tri 39067 18865 39075 18873 ne
rect 39075 18865 39343 18873
tri 39343 18865 39351 18873 sw
tri 39075 18857 39083 18865 ne
rect 39083 18857 39351 18865
tri 39351 18857 39359 18865 sw
tri 39083 18849 39091 18857 ne
rect 39091 18849 39359 18857
tri 39359 18849 39367 18857 sw
tri 39091 18841 39099 18849 ne
rect 39099 18841 39367 18849
tri 39367 18841 39375 18849 sw
tri 39099 18833 39107 18841 ne
rect 39107 18833 39375 18841
tri 39375 18833 39383 18841 sw
tri 39107 18825 39115 18833 ne
rect 39115 18825 39383 18833
tri 39383 18825 39391 18833 sw
tri 39115 18817 39123 18825 ne
rect 39123 18817 39391 18825
tri 39391 18817 39399 18825 sw
tri 39123 18809 39131 18817 ne
rect 39131 18809 39399 18817
tri 39399 18809 39407 18817 sw
tri 39131 18801 39139 18809 ne
rect 39139 18801 39407 18809
tri 39407 18801 39415 18809 sw
tri 39139 18793 39147 18801 ne
rect 39147 18793 39415 18801
tri 39415 18793 39423 18801 sw
tri 39147 18785 39155 18793 ne
rect 39155 18785 39423 18793
tri 39423 18785 39431 18793 sw
tri 39155 18777 39163 18785 ne
rect 39163 18777 39431 18785
tri 39431 18777 39439 18785 sw
tri 39163 18769 39171 18777 ne
rect 39171 18769 39439 18777
tri 39439 18769 39447 18777 sw
tri 39171 18761 39179 18769 ne
rect 39179 18761 39447 18769
tri 39447 18761 39455 18769 sw
tri 39179 18753 39187 18761 ne
rect 39187 18753 39455 18761
tri 39455 18753 39463 18761 sw
tri 39187 18749 39191 18753 ne
rect 39191 18749 39463 18753
tri 39191 18741 39199 18749 ne
rect 39199 18745 39463 18749
tri 39463 18745 39471 18753 sw
rect 39199 18741 39471 18745
tri 39199 18733 39207 18741 ne
rect 39207 18737 39471 18741
tri 39471 18737 39479 18745 sw
rect 39207 18733 39479 18737
tri 39207 18725 39215 18733 ne
rect 39215 18729 39479 18733
tri 39479 18729 39487 18737 sw
rect 39215 18725 39487 18729
tri 39215 18717 39223 18725 ne
rect 39223 18721 39487 18725
tri 39487 18721 39495 18729 sw
rect 39223 18717 39495 18721
tri 39223 18709 39231 18717 ne
rect 39231 18713 39495 18717
tri 39495 18713 39503 18721 sw
rect 39231 18709 39503 18713
tri 39231 18701 39239 18709 ne
rect 39239 18705 39503 18709
tri 39503 18705 39511 18713 sw
rect 39239 18701 39511 18705
tri 39239 18693 39247 18701 ne
rect 39247 18697 39511 18701
tri 39511 18697 39519 18705 sw
rect 39247 18693 39519 18697
tri 39247 18685 39255 18693 ne
rect 39255 18689 39519 18693
tri 39519 18689 39527 18697 sw
rect 39255 18685 39527 18689
tri 39255 18677 39263 18685 ne
rect 39263 18681 39527 18685
tri 39527 18681 39535 18689 sw
rect 39263 18677 39535 18681
tri 39263 18669 39271 18677 ne
rect 39271 18673 39535 18677
tri 39535 18673 39543 18681 sw
rect 39271 18669 39543 18673
tri 39271 18661 39279 18669 ne
rect 39279 18665 39543 18669
tri 39543 18665 39551 18673 sw
rect 39279 18661 39551 18665
tri 39279 18653 39287 18661 ne
rect 39287 18657 39551 18661
tri 39551 18657 39559 18665 sw
rect 39287 18653 39559 18657
tri 39287 18645 39295 18653 ne
rect 39295 18649 39559 18653
tri 39559 18649 39567 18657 sw
rect 39295 18645 39567 18649
tri 39295 18637 39303 18645 ne
rect 39303 18641 39567 18645
tri 39567 18641 39575 18649 sw
rect 39303 18637 39575 18641
tri 39303 18629 39311 18637 ne
rect 39311 18633 39575 18637
tri 39575 18633 39583 18641 sw
rect 39311 18629 39583 18633
tri 39311 18621 39319 18629 ne
rect 39319 18625 39583 18629
tri 39583 18625 39591 18633 sw
rect 39319 18621 39591 18625
tri 39319 18617 39323 18621 ne
rect 39323 18617 39591 18621
tri 39591 18617 39599 18625 sw
tri 39323 18613 39327 18617 ne
rect 39327 18613 39599 18617
tri 39599 18613 39603 18617 sw
tri 39327 18605 39335 18613 ne
rect 39335 18605 39603 18613
tri 39603 18605 39611 18613 sw
tri 39335 18597 39343 18605 ne
rect 39343 18597 39611 18605
tri 39611 18597 39619 18605 sw
tri 39343 18589 39351 18597 ne
rect 39351 18589 39619 18597
tri 39619 18589 39627 18597 sw
tri 39351 18581 39359 18589 ne
rect 39359 18581 39627 18589
tri 39627 18581 39635 18589 sw
tri 39359 18573 39367 18581 ne
rect 39367 18573 39635 18581
tri 39635 18573 39643 18581 sw
tri 39367 18565 39375 18573 ne
rect 39375 18565 39643 18573
tri 39643 18565 39651 18573 sw
tri 39375 18557 39383 18565 ne
rect 39383 18557 39651 18565
tri 39651 18557 39659 18565 sw
tri 39383 18549 39391 18557 ne
rect 39391 18549 39659 18557
tri 39659 18549 39667 18557 sw
tri 39391 18541 39399 18549 ne
rect 39399 18541 39667 18549
tri 39667 18541 39675 18549 sw
tri 39399 18533 39407 18541 ne
rect 39407 18533 39675 18541
tri 39675 18533 39683 18541 sw
tri 39407 18525 39415 18533 ne
rect 39415 18525 39683 18533
tri 39683 18525 39691 18533 sw
tri 39415 18517 39423 18525 ne
rect 39423 18517 39691 18525
tri 39691 18517 39699 18525 sw
tri 39423 18509 39431 18517 ne
rect 39431 18509 39699 18517
tri 39699 18509 39707 18517 sw
tri 39431 18501 39439 18509 ne
rect 39439 18501 39707 18509
tri 39707 18501 39715 18509 sw
tri 39439 18493 39447 18501 ne
rect 39447 18493 39715 18501
tri 39715 18493 39723 18501 sw
tri 39447 18485 39455 18493 ne
rect 39455 18485 39723 18493
tri 39723 18485 39731 18493 sw
tri 39455 18477 39463 18485 ne
rect 39463 18477 39731 18485
tri 39731 18477 39739 18485 sw
tri 39463 18473 39467 18477 ne
rect 39467 18473 39739 18477
tri 39467 18465 39475 18473 ne
rect 39475 18469 39739 18473
tri 39739 18469 39747 18477 sw
rect 39475 18465 39747 18469
tri 39475 18457 39483 18465 ne
rect 39483 18461 39747 18465
tri 39747 18461 39755 18469 sw
rect 39483 18457 39755 18461
tri 39483 18449 39491 18457 ne
rect 39491 18453 39755 18457
tri 39755 18453 39763 18461 sw
rect 39491 18449 39763 18453
tri 39491 18441 39499 18449 ne
rect 39499 18445 39763 18449
tri 39763 18445 39771 18453 sw
rect 39499 18441 39771 18445
tri 39499 18433 39507 18441 ne
rect 39507 18437 39771 18441
tri 39771 18437 39779 18445 sw
rect 39507 18433 39779 18437
tri 39507 18425 39515 18433 ne
rect 39515 18429 39779 18433
tri 39779 18429 39787 18437 sw
rect 39515 18425 39787 18429
tri 39515 18417 39523 18425 ne
rect 39523 18421 39787 18425
tri 39787 18421 39795 18429 sw
rect 39523 18417 39795 18421
tri 39523 18409 39531 18417 ne
rect 39531 18413 39795 18417
tri 39795 18413 39803 18421 sw
rect 39531 18409 39803 18413
tri 39531 18401 39539 18409 ne
rect 39539 18405 39803 18409
tri 39803 18405 39811 18413 sw
rect 39539 18401 39811 18405
tri 39539 18393 39547 18401 ne
rect 39547 18397 39811 18401
tri 39811 18397 39819 18405 sw
rect 39547 18393 39819 18397
tri 39547 18385 39555 18393 ne
rect 39555 18389 39819 18393
tri 39819 18389 39827 18397 sw
rect 39555 18385 39827 18389
tri 39555 18377 39563 18385 ne
rect 39563 18381 39827 18385
tri 39827 18381 39835 18389 sw
rect 39563 18377 39835 18381
tri 39563 18369 39571 18377 ne
rect 39571 18373 39835 18377
tri 39835 18373 39843 18381 sw
rect 39571 18369 39843 18373
tri 39571 18361 39579 18369 ne
rect 39579 18365 39843 18369
tri 39843 18365 39851 18373 sw
rect 39579 18361 39851 18365
tri 39579 18353 39587 18361 ne
rect 39587 18357 39851 18361
tri 39851 18357 39859 18365 sw
rect 39587 18353 39859 18357
tri 39587 18345 39595 18353 ne
rect 39595 18349 39859 18353
tri 39859 18349 39867 18357 sw
rect 39595 18345 39867 18349
tri 39595 18341 39599 18345 ne
rect 39599 18341 39867 18345
tri 39867 18341 39875 18349 sw
tri 39599 18337 39603 18341 ne
rect 39603 18337 39875 18341
tri 39875 18337 39879 18341 sw
tri 39603 18329 39611 18337 ne
rect 39611 18329 39879 18337
tri 39879 18329 39887 18337 sw
tri 39611 18321 39619 18329 ne
rect 39619 18321 39887 18329
tri 39887 18321 39895 18329 sw
tri 39619 18313 39627 18321 ne
rect 39627 18313 39895 18321
tri 39895 18313 39903 18321 sw
tri 39627 18305 39635 18313 ne
rect 39635 18305 39903 18313
tri 39903 18305 39911 18313 sw
tri 39635 18297 39643 18305 ne
rect 39643 18297 39911 18305
tri 39911 18297 39919 18305 sw
tri 39643 18289 39651 18297 ne
rect 39651 18289 39919 18297
tri 39919 18289 39927 18297 sw
tri 39651 18281 39659 18289 ne
rect 39659 18281 39927 18289
tri 39927 18281 39935 18289 sw
tri 39659 18273 39667 18281 ne
rect 39667 18273 39935 18281
tri 39935 18273 39943 18281 sw
tri 39667 18265 39675 18273 ne
rect 39675 18265 39943 18273
tri 39943 18265 39951 18273 sw
tri 39675 18257 39683 18265 ne
rect 39683 18257 39951 18265
tri 39951 18257 39959 18265 sw
tri 39683 18249 39691 18257 ne
rect 39691 18249 39959 18257
tri 39959 18249 39967 18257 sw
tri 39691 18241 39699 18249 ne
rect 39699 18241 39967 18249
tri 39967 18241 39975 18249 sw
tri 39699 18233 39707 18241 ne
rect 39707 18233 39975 18241
tri 39975 18233 39983 18241 sw
tri 39707 18225 39715 18233 ne
rect 39715 18225 39983 18233
tri 39983 18225 39991 18233 sw
tri 39715 18217 39723 18225 ne
rect 39723 18217 39991 18225
tri 39991 18217 39999 18225 sw
tri 39723 18209 39731 18217 ne
rect 39731 18209 39999 18217
tri 39999 18209 40007 18217 sw
tri 39731 18201 39739 18209 ne
rect 39739 18201 40007 18209
tri 40007 18201 40015 18209 sw
tri 39739 18197 39743 18201 ne
rect 39743 18197 40015 18201
tri 39743 18189 39751 18197 ne
rect 39751 18193 40015 18197
tri 40015 18193 40023 18201 sw
rect 39751 18189 40023 18193
tri 39751 18181 39759 18189 ne
rect 39759 18185 40023 18189
tri 40023 18185 40031 18193 sw
rect 39759 18181 40031 18185
tri 39759 18173 39767 18181 ne
rect 39767 18177 40031 18181
tri 40031 18177 40039 18185 sw
rect 39767 18173 40039 18177
tri 39767 18165 39775 18173 ne
rect 39775 18169 40039 18173
tri 40039 18169 40047 18177 sw
rect 39775 18165 40047 18169
tri 39775 18157 39783 18165 ne
rect 39783 18161 40047 18165
tri 40047 18161 40055 18169 sw
rect 39783 18157 40055 18161
tri 39783 18149 39791 18157 ne
rect 39791 18153 40055 18157
tri 40055 18153 40063 18161 sw
rect 39791 18149 40063 18153
tri 39791 18141 39799 18149 ne
rect 39799 18145 40063 18149
tri 40063 18145 40071 18153 sw
rect 39799 18141 40071 18145
tri 39799 18133 39807 18141 ne
rect 39807 18137 40071 18141
tri 40071 18137 40079 18145 sw
rect 39807 18133 40079 18137
tri 39807 18125 39815 18133 ne
rect 39815 18129 40079 18133
tri 40079 18129 40087 18137 sw
rect 39815 18125 40087 18129
tri 39815 18117 39823 18125 ne
rect 39823 18121 40087 18125
tri 40087 18121 40095 18129 sw
rect 39823 18117 40095 18121
tri 39823 18109 39831 18117 ne
rect 39831 18113 40095 18117
tri 40095 18113 40103 18121 sw
rect 39831 18109 40103 18113
tri 39831 18101 39839 18109 ne
rect 39839 18105 40103 18109
tri 40103 18105 40111 18113 sw
rect 39839 18101 40111 18105
tri 39839 18093 39847 18101 ne
rect 39847 18097 40111 18101
tri 40111 18097 40119 18105 sw
rect 39847 18093 40119 18097
tri 39847 18085 39855 18093 ne
rect 39855 18089 40119 18093
tri 40119 18089 40127 18097 sw
rect 39855 18085 40127 18089
tri 39855 18077 39863 18085 ne
rect 39863 18081 40127 18085
tri 40127 18081 40135 18089 sw
rect 39863 18077 40135 18081
tri 39863 18069 39871 18077 ne
rect 39871 18073 40135 18077
tri 40135 18073 40143 18081 sw
rect 39871 18069 40143 18073
tri 39871 18065 39875 18069 ne
rect 39875 18065 40143 18069
tri 40143 18065 40151 18073 sw
tri 39875 18061 39879 18065 ne
rect 39879 18061 40151 18065
tri 40151 18061 40155 18065 sw
tri 39879 18053 39887 18061 ne
rect 39887 18053 40155 18061
tri 40155 18053 40163 18061 sw
tri 39887 18045 39895 18053 ne
rect 39895 18045 40163 18053
tri 40163 18045 40171 18053 sw
tri 39895 18037 39903 18045 ne
rect 39903 18037 40171 18045
tri 40171 18037 40179 18045 sw
tri 39903 18029 39911 18037 ne
rect 39911 18029 40179 18037
tri 40179 18029 40187 18037 sw
tri 39911 18021 39919 18029 ne
rect 39919 18021 40187 18029
tri 40187 18021 40195 18029 sw
tri 39919 18013 39927 18021 ne
rect 39927 18013 40195 18021
tri 40195 18013 40203 18021 sw
tri 39927 18005 39935 18013 ne
rect 39935 18005 40203 18013
tri 40203 18005 40211 18013 sw
tri 39935 17997 39943 18005 ne
rect 39943 17997 40211 18005
tri 40211 17997 40219 18005 sw
tri 39943 17989 39951 17997 ne
rect 39951 17989 40219 17997
tri 40219 17989 40227 17997 sw
tri 39951 17981 39959 17989 ne
rect 39959 17981 40227 17989
tri 40227 17981 40235 17989 sw
tri 39959 17973 39967 17981 ne
rect 39967 17973 40235 17981
tri 40235 17973 40243 17981 sw
tri 39967 17965 39975 17973 ne
rect 39975 17965 40243 17973
tri 40243 17965 40251 17973 sw
tri 39975 17957 39983 17965 ne
rect 39983 17957 40251 17965
tri 40251 17957 40259 17965 sw
tri 39983 17949 39991 17957 ne
rect 39991 17949 40259 17957
tri 40259 17949 40267 17957 sw
tri 39991 17941 39999 17949 ne
rect 39999 17941 40267 17949
tri 40267 17941 40275 17949 sw
tri 39999 17933 40007 17941 ne
rect 40007 17933 40275 17941
tri 40275 17933 40283 17941 sw
tri 40007 17925 40015 17933 ne
rect 40015 17925 40283 17933
tri 40283 17925 40291 17933 sw
tri 40015 17921 40019 17925 ne
rect 40019 17921 40291 17925
tri 40019 17913 40027 17921 ne
rect 40027 17917 40291 17921
tri 40291 17917 40299 17925 sw
rect 40027 17913 40299 17917
tri 40027 17905 40035 17913 ne
rect 40035 17909 40299 17913
tri 40299 17909 40307 17917 sw
rect 40035 17905 40307 17909
tri 40035 17897 40043 17905 ne
rect 40043 17901 40307 17905
tri 40307 17901 40315 17909 sw
rect 40043 17897 40315 17901
tri 40043 17889 40051 17897 ne
rect 40051 17893 40315 17897
tri 40315 17893 40323 17901 sw
rect 40051 17889 40323 17893
tri 40051 17881 40059 17889 ne
rect 40059 17885 40323 17889
tri 40323 17885 40331 17893 sw
rect 40059 17881 40331 17885
tri 40059 17873 40067 17881 ne
rect 40067 17877 40331 17881
tri 40331 17877 40339 17885 sw
rect 40067 17873 40339 17877
tri 40067 17865 40075 17873 ne
rect 40075 17869 40339 17873
tri 40339 17869 40347 17877 sw
rect 40075 17865 40347 17869
tri 40075 17857 40083 17865 ne
rect 40083 17861 40347 17865
tri 40347 17861 40355 17869 sw
rect 40083 17857 40355 17861
tri 40083 17849 40091 17857 ne
rect 40091 17853 40355 17857
tri 40355 17853 40363 17861 sw
rect 40091 17849 40363 17853
tri 40091 17841 40099 17849 ne
rect 40099 17845 40363 17849
tri 40363 17845 40371 17853 sw
rect 40099 17841 40371 17845
tri 40099 17833 40107 17841 ne
rect 40107 17837 40371 17841
tri 40371 17837 40379 17845 sw
rect 40107 17833 40379 17837
tri 40107 17825 40115 17833 ne
rect 40115 17829 40379 17833
tri 40379 17829 40387 17837 sw
rect 40115 17825 40387 17829
tri 40115 17817 40123 17825 ne
rect 40123 17821 40387 17825
tri 40387 17821 40395 17829 sw
rect 40123 17817 40395 17821
tri 40123 17809 40131 17817 ne
rect 40131 17813 40395 17817
tri 40395 17813 40403 17821 sw
rect 40131 17809 40403 17813
tri 40131 17801 40139 17809 ne
rect 40139 17805 40403 17809
tri 40403 17805 40411 17813 sw
rect 40139 17801 40411 17805
tri 40139 17793 40147 17801 ne
rect 40147 17797 40411 17801
tri 40411 17797 40419 17805 sw
rect 40147 17793 40419 17797
tri 40147 17789 40151 17793 ne
rect 40151 17789 40419 17793
tri 40419 17789 40427 17797 sw
tri 40151 17785 40155 17789 ne
rect 40155 17785 40427 17789
tri 40427 17785 40431 17789 sw
tri 40155 17777 40163 17785 ne
rect 40163 17777 40431 17785
tri 40431 17777 40439 17785 sw
tri 40163 17769 40171 17777 ne
rect 40171 17769 40439 17777
tri 40439 17769 40447 17777 sw
tri 40171 17761 40179 17769 ne
rect 40179 17761 40447 17769
tri 40447 17761 40455 17769 sw
tri 40179 17753 40187 17761 ne
rect 40187 17753 40455 17761
tri 40455 17753 40463 17761 sw
tri 40187 17745 40195 17753 ne
rect 40195 17745 40463 17753
tri 40463 17745 40471 17753 sw
tri 40195 17737 40203 17745 ne
rect 40203 17737 40471 17745
tri 40471 17737 40479 17745 sw
tri 40203 17729 40211 17737 ne
rect 40211 17729 40479 17737
tri 40479 17729 40487 17737 sw
tri 40211 17721 40219 17729 ne
rect 40219 17721 40487 17729
tri 40487 17721 40495 17729 sw
tri 40219 17713 40227 17721 ne
rect 40227 17713 40495 17721
tri 40495 17713 40503 17721 sw
tri 40227 17705 40235 17713 ne
rect 40235 17705 40503 17713
tri 40503 17705 40511 17713 sw
tri 40235 17697 40243 17705 ne
rect 40243 17697 40511 17705
tri 40511 17697 40519 17705 sw
tri 40243 17689 40251 17697 ne
rect 40251 17689 40519 17697
tri 40519 17689 40527 17697 sw
tri 40251 17681 40259 17689 ne
rect 40259 17681 40527 17689
tri 40527 17681 40535 17689 sw
tri 40259 17673 40267 17681 ne
rect 40267 17673 40535 17681
tri 40535 17673 40543 17681 sw
tri 40267 17665 40275 17673 ne
rect 40275 17665 40543 17673
tri 40543 17665 40551 17673 sw
tri 40275 17657 40283 17665 ne
rect 40283 17657 40551 17665
tri 40551 17657 40559 17665 sw
tri 40283 17649 40291 17657 ne
rect 40291 17649 40559 17657
tri 40559 17649 40567 17657 sw
tri 40291 17645 40295 17649 ne
rect 40295 17645 40567 17649
tri 40295 17637 40303 17645 ne
rect 40303 17641 40567 17645
tri 40567 17641 40575 17649 sw
rect 40303 17637 40575 17641
tri 40303 17629 40311 17637 ne
rect 40311 17633 40575 17637
tri 40575 17633 40583 17641 sw
rect 40311 17629 40583 17633
tri 40311 17621 40319 17629 ne
rect 40319 17625 40583 17629
tri 40583 17625 40591 17633 sw
rect 40319 17621 40591 17625
tri 40319 17613 40327 17621 ne
rect 40327 17617 40591 17621
tri 40591 17617 40599 17625 sw
rect 40327 17613 40599 17617
tri 40327 17605 40335 17613 ne
rect 40335 17609 40599 17613
tri 40599 17609 40607 17617 sw
rect 40335 17605 40607 17609
tri 40335 17597 40343 17605 ne
rect 40343 17601 40607 17605
tri 40607 17601 40615 17609 sw
rect 40343 17597 40615 17601
tri 40343 17589 40351 17597 ne
rect 40351 17593 40615 17597
tri 40615 17593 40623 17601 sw
rect 40351 17589 40623 17593
tri 40351 17581 40359 17589 ne
rect 40359 17585 40623 17589
tri 40623 17585 40631 17593 sw
rect 40359 17581 40631 17585
tri 40359 17573 40367 17581 ne
rect 40367 17577 40631 17581
tri 40631 17577 40639 17585 sw
rect 40367 17573 40639 17577
tri 40367 17565 40375 17573 ne
rect 40375 17569 40639 17573
tri 40639 17569 40647 17577 sw
rect 40375 17565 40647 17569
tri 40375 17557 40383 17565 ne
rect 40383 17561 40647 17565
tri 40647 17561 40655 17569 sw
rect 40383 17557 40655 17561
tri 40383 17549 40391 17557 ne
rect 40391 17553 40655 17557
tri 40655 17553 40663 17561 sw
rect 40391 17549 40663 17553
tri 40391 17541 40399 17549 ne
rect 40399 17545 40663 17549
tri 40663 17545 40671 17553 sw
rect 40399 17541 40671 17545
tri 40399 17533 40407 17541 ne
rect 40407 17537 40671 17541
tri 40671 17537 40679 17545 sw
rect 40407 17533 40679 17537
tri 40407 17525 40415 17533 ne
rect 40415 17529 40679 17533
tri 40679 17529 40687 17537 sw
rect 40415 17525 40687 17529
tri 40415 17517 40423 17525 ne
rect 40423 17521 40687 17525
tri 40687 17521 40695 17529 sw
rect 40423 17517 40695 17521
tri 40423 17513 40427 17517 ne
rect 40427 17513 40695 17517
tri 40695 17513 40703 17521 sw
tri 40427 17509 40431 17513 ne
rect 40431 17509 40703 17513
tri 40703 17509 40707 17513 sw
tri 40431 17501 40439 17509 ne
rect 40439 17501 40707 17509
tri 40707 17501 40715 17509 sw
tri 40439 17493 40447 17501 ne
rect 40447 17493 40715 17501
tri 40715 17493 40723 17501 sw
tri 40447 17485 40455 17493 ne
rect 40455 17485 40723 17493
tri 40723 17485 40731 17493 sw
tri 40455 17477 40463 17485 ne
rect 40463 17477 40731 17485
tri 40731 17477 40739 17485 sw
tri 40463 17469 40471 17477 ne
rect 40471 17469 40739 17477
tri 40739 17469 40747 17477 sw
tri 40471 17461 40479 17469 ne
rect 40479 17461 40747 17469
tri 40747 17461 40755 17469 sw
tri 40479 17453 40487 17461 ne
rect 40487 17453 40755 17461
tri 40755 17453 40763 17461 sw
tri 40487 17445 40495 17453 ne
rect 40495 17445 40763 17453
tri 40763 17445 40771 17453 sw
tri 40495 17437 40503 17445 ne
rect 40503 17437 40771 17445
tri 40771 17437 40779 17445 sw
tri 40503 17429 40511 17437 ne
rect 40511 17429 40779 17437
tri 40779 17429 40787 17437 sw
tri 40511 17421 40519 17429 ne
rect 40519 17421 40787 17429
tri 40787 17421 40795 17429 sw
tri 40519 17413 40527 17421 ne
rect 40527 17413 40795 17421
tri 40795 17413 40803 17421 sw
tri 40527 17405 40535 17413 ne
rect 40535 17405 40803 17413
tri 40803 17405 40811 17413 sw
tri 40535 17397 40543 17405 ne
rect 40543 17397 40811 17405
tri 40811 17397 40819 17405 sw
tri 40543 17389 40551 17397 ne
rect 40551 17389 40819 17397
tri 40819 17389 40827 17397 sw
tri 40551 17381 40559 17389 ne
rect 40559 17381 40827 17389
tri 40827 17381 40835 17389 sw
tri 40559 17373 40567 17381 ne
rect 40567 17373 40835 17381
tri 40835 17373 40843 17381 sw
tri 40567 17369 40571 17373 ne
rect 40571 17369 40843 17373
tri 40571 17361 40579 17369 ne
rect 40579 17365 40843 17369
tri 40843 17365 40851 17373 sw
rect 40579 17361 40851 17365
tri 40579 17353 40587 17361 ne
rect 40587 17357 40851 17361
tri 40851 17357 40859 17365 sw
rect 40587 17353 40859 17357
tri 40587 17345 40595 17353 ne
rect 40595 17349 40859 17353
tri 40859 17349 40867 17357 sw
rect 40595 17345 40867 17349
tri 40595 17337 40603 17345 ne
rect 40603 17341 40867 17345
tri 40867 17341 40875 17349 sw
rect 40603 17337 40875 17341
tri 40603 17329 40611 17337 ne
rect 40611 17333 40875 17337
tri 40875 17333 40883 17341 sw
rect 40611 17329 40883 17333
tri 40611 17321 40619 17329 ne
rect 40619 17325 40883 17329
tri 40883 17325 40891 17333 sw
rect 40619 17321 40891 17325
tri 40619 17313 40627 17321 ne
rect 40627 17317 40891 17321
tri 40891 17317 40899 17325 sw
rect 40627 17313 40899 17317
tri 40627 17305 40635 17313 ne
rect 40635 17309 40899 17313
tri 40899 17309 40907 17317 sw
rect 40635 17305 40907 17309
tri 40635 17297 40643 17305 ne
rect 40643 17301 40907 17305
tri 40907 17301 40915 17309 sw
rect 40643 17297 40915 17301
tri 40643 17289 40651 17297 ne
rect 40651 17293 40915 17297
tri 40915 17293 40923 17301 sw
rect 40651 17289 40923 17293
tri 40651 17281 40659 17289 ne
rect 40659 17285 40923 17289
tri 40923 17285 40931 17293 sw
rect 40659 17281 40931 17285
tri 40659 17273 40667 17281 ne
rect 40667 17277 40931 17281
tri 40931 17277 40939 17285 sw
rect 40667 17273 40939 17277
tri 40667 17265 40675 17273 ne
rect 40675 17269 40939 17273
tri 40939 17269 40947 17277 sw
rect 40675 17265 40947 17269
tri 40675 17257 40683 17265 ne
rect 40683 17261 40947 17265
tri 40947 17261 40955 17269 sw
rect 40683 17257 40955 17261
tri 40683 17249 40691 17257 ne
rect 40691 17253 40955 17257
tri 40955 17253 40963 17261 sw
rect 40691 17249 40963 17253
tri 40691 17241 40699 17249 ne
rect 40699 17245 40963 17249
tri 40963 17245 40971 17253 sw
rect 40699 17241 40971 17245
tri 40699 17237 40703 17241 ne
rect 40703 17237 40971 17241
tri 40971 17237 40979 17245 sw
tri 40703 17233 40707 17237 ne
rect 40707 17233 40979 17237
tri 40979 17233 40983 17237 sw
tri 40707 17225 40715 17233 ne
rect 40715 17225 40983 17233
tri 40983 17225 40991 17233 sw
tri 40715 17217 40723 17225 ne
rect 40723 17217 40991 17225
tri 40991 17217 40999 17225 sw
tri 40723 17209 40731 17217 ne
rect 40731 17209 40999 17217
tri 40999 17209 41007 17217 sw
tri 40731 17201 40739 17209 ne
rect 40739 17201 41007 17209
tri 41007 17201 41015 17209 sw
tri 40739 17193 40747 17201 ne
rect 40747 17193 41015 17201
tri 41015 17193 41023 17201 sw
tri 40747 17185 40755 17193 ne
rect 40755 17185 41023 17193
tri 41023 17185 41031 17193 sw
tri 40755 17177 40763 17185 ne
rect 40763 17177 41031 17185
tri 41031 17177 41039 17185 sw
tri 40763 17169 40771 17177 ne
rect 40771 17169 41039 17177
tri 41039 17169 41047 17177 sw
tri 40771 17161 40779 17169 ne
rect 40779 17161 41047 17169
tri 41047 17161 41055 17169 sw
tri 40779 17153 40787 17161 ne
rect 40787 17153 41055 17161
tri 41055 17153 41063 17161 sw
tri 40787 17145 40795 17153 ne
rect 40795 17145 41063 17153
tri 41063 17145 41071 17153 sw
tri 40795 17137 40803 17145 ne
rect 40803 17137 41071 17145
tri 41071 17137 41079 17145 sw
tri 40803 17129 40811 17137 ne
rect 40811 17129 41079 17137
tri 41079 17129 41087 17137 sw
tri 40811 17121 40819 17129 ne
rect 40819 17121 41087 17129
tri 41087 17121 41095 17129 sw
tri 40819 17113 40827 17121 ne
rect 40827 17113 41095 17121
tri 41095 17113 41103 17121 sw
tri 40827 17105 40835 17113 ne
rect 40835 17105 41103 17113
tri 41103 17105 41111 17113 sw
tri 40835 17097 40843 17105 ne
rect 40843 17097 41111 17105
tri 41111 17097 41119 17105 sw
tri 40843 17093 40847 17097 ne
rect 40847 17093 41119 17097
tri 40847 17085 40855 17093 ne
rect 40855 17089 41119 17093
tri 41119 17089 41127 17097 sw
rect 40855 17085 41127 17089
tri 40855 17077 40863 17085 ne
rect 40863 17081 41127 17085
tri 41127 17081 41135 17089 sw
rect 40863 17077 41135 17081
tri 40863 17069 40871 17077 ne
rect 40871 17073 41135 17077
tri 41135 17073 41143 17081 sw
rect 40871 17069 41143 17073
tri 40871 17061 40879 17069 ne
rect 40879 17065 41143 17069
tri 41143 17065 41151 17073 sw
rect 40879 17061 41151 17065
tri 40879 17053 40887 17061 ne
rect 40887 17057 41151 17061
tri 41151 17057 41159 17065 sw
rect 40887 17053 41159 17057
tri 40887 17045 40895 17053 ne
rect 40895 17049 41159 17053
tri 41159 17049 41167 17057 sw
rect 40895 17045 41167 17049
tri 40895 17037 40903 17045 ne
rect 40903 17041 41167 17045
tri 41167 17041 41175 17049 sw
rect 40903 17037 41175 17041
tri 40903 17029 40911 17037 ne
rect 40911 17033 41175 17037
tri 41175 17033 41183 17041 sw
rect 40911 17029 41183 17033
tri 40911 17021 40919 17029 ne
rect 40919 17025 41183 17029
tri 41183 17025 41191 17033 sw
rect 40919 17021 41191 17025
tri 40919 17013 40927 17021 ne
rect 40927 17017 41191 17021
tri 41191 17017 41199 17025 sw
rect 40927 17013 41199 17017
tri 40927 17005 40935 17013 ne
rect 40935 17009 41199 17013
tri 41199 17009 41207 17017 sw
rect 40935 17005 41207 17009
tri 40935 16997 40943 17005 ne
rect 40943 17001 41207 17005
tri 41207 17001 41215 17009 sw
rect 40943 16997 41215 17001
tri 40943 16989 40951 16997 ne
rect 40951 16993 41215 16997
tri 41215 16993 41223 17001 sw
rect 40951 16989 41223 16993
tri 40951 16981 40959 16989 ne
rect 40959 16985 41223 16989
tri 41223 16985 41231 16993 sw
rect 40959 16981 41231 16985
tri 40959 16973 40967 16981 ne
rect 40967 16977 41231 16981
tri 41231 16977 41239 16985 sw
rect 40967 16973 41239 16977
tri 40967 16965 40975 16973 ne
rect 40975 16969 41239 16973
tri 41239 16969 41247 16977 sw
rect 40975 16965 41247 16969
tri 40975 16961 40979 16965 ne
rect 40979 16961 41247 16965
tri 41247 16961 41255 16969 sw
tri 40979 16957 40983 16961 ne
rect 40983 16957 41255 16961
tri 41255 16957 41259 16961 sw
tri 40983 16949 40991 16957 ne
rect 40991 16949 41259 16957
tri 41259 16949 41267 16957 sw
tri 40991 16941 40999 16949 ne
rect 40999 16941 41267 16949
tri 41267 16941 41275 16949 sw
tri 40999 16933 41007 16941 ne
rect 41007 16933 41275 16941
tri 41275 16933 41283 16941 sw
tri 41007 16925 41015 16933 ne
rect 41015 16925 41283 16933
tri 41283 16925 41291 16933 sw
tri 41015 16917 41023 16925 ne
rect 41023 16917 41291 16925
tri 41291 16917 41299 16925 sw
tri 41023 16909 41031 16917 ne
rect 41031 16909 41299 16917
tri 41299 16909 41307 16917 sw
tri 41031 16901 41039 16909 ne
rect 41039 16901 41307 16909
tri 41307 16901 41315 16909 sw
tri 41039 16893 41047 16901 ne
rect 41047 16893 41315 16901
tri 41315 16893 41323 16901 sw
tri 41047 16885 41055 16893 ne
rect 41055 16885 41323 16893
tri 41323 16885 41331 16893 sw
tri 41055 16877 41063 16885 ne
rect 41063 16877 41331 16885
tri 41331 16877 41339 16885 sw
tri 41063 16869 41071 16877 ne
rect 41071 16869 41339 16877
tri 41339 16869 41347 16877 sw
tri 41071 16861 41079 16869 ne
rect 41079 16861 41347 16869
tri 41347 16861 41355 16869 sw
tri 41079 16853 41087 16861 ne
rect 41087 16853 41355 16861
tri 41355 16853 41363 16861 sw
tri 41087 16845 41095 16853 ne
rect 41095 16845 41363 16853
tri 41363 16845 41371 16853 sw
tri 41095 16837 41103 16845 ne
rect 41103 16837 41371 16845
tri 41371 16837 41379 16845 sw
tri 41103 16829 41111 16837 ne
rect 41111 16829 41379 16837
tri 41379 16829 41387 16837 sw
tri 41111 16821 41119 16829 ne
rect 41119 16821 41387 16829
tri 41387 16821 41395 16829 sw
tri 41119 16817 41123 16821 ne
rect 41123 16817 41395 16821
tri 41123 16809 41131 16817 ne
rect 41131 16813 41395 16817
tri 41395 16813 41403 16821 sw
rect 41131 16809 41403 16813
tri 41131 16801 41139 16809 ne
rect 41139 16805 41403 16809
tri 41403 16805 41411 16813 sw
rect 41139 16801 41411 16805
tri 41139 16793 41147 16801 ne
rect 41147 16797 41411 16801
tri 41411 16797 41419 16805 sw
rect 41147 16793 41419 16797
tri 41147 16785 41155 16793 ne
rect 41155 16789 41419 16793
tri 41419 16789 41427 16797 sw
rect 41155 16785 41427 16789
tri 41155 16777 41163 16785 ne
rect 41163 16781 41427 16785
tri 41427 16781 41435 16789 sw
rect 41163 16777 41435 16781
tri 41163 16769 41171 16777 ne
rect 41171 16773 41435 16777
tri 41435 16773 41443 16781 sw
rect 41171 16769 41443 16773
tri 41171 16761 41179 16769 ne
rect 41179 16765 41443 16769
tri 41443 16765 41451 16773 sw
rect 41179 16761 41451 16765
tri 41179 16753 41187 16761 ne
rect 41187 16757 41451 16761
tri 41451 16757 41459 16765 sw
rect 41187 16753 41459 16757
tri 41187 16745 41195 16753 ne
rect 41195 16749 41459 16753
tri 41459 16749 41467 16757 sw
rect 41195 16745 41467 16749
tri 41195 16737 41203 16745 ne
rect 41203 16741 41467 16745
tri 41467 16741 41475 16749 sw
rect 41203 16737 41475 16741
tri 41203 16729 41211 16737 ne
rect 41211 16733 41475 16737
tri 41475 16733 41483 16741 sw
rect 41211 16729 41483 16733
tri 41211 16721 41219 16729 ne
rect 41219 16725 41483 16729
tri 41483 16725 41491 16733 sw
rect 41219 16721 41491 16725
tri 41219 16713 41227 16721 ne
rect 41227 16717 41491 16721
tri 41491 16717 41499 16725 sw
rect 41227 16713 41499 16717
tri 41227 16705 41235 16713 ne
rect 41235 16709 41499 16713
tri 41499 16709 41507 16717 sw
rect 41235 16705 41507 16709
tri 41235 16697 41243 16705 ne
rect 41243 16701 41507 16705
tri 41507 16701 41515 16709 sw
rect 41243 16697 41515 16701
tri 41243 16689 41251 16697 ne
rect 41251 16693 41515 16697
tri 41515 16693 41523 16701 sw
rect 41251 16689 41523 16693
tri 41251 16685 41255 16689 ne
rect 41255 16685 41523 16689
tri 41523 16685 41531 16693 sw
tri 41255 16681 41259 16685 ne
rect 41259 16681 41531 16685
tri 41531 16681 41535 16685 sw
tri 41259 16673 41267 16681 ne
rect 41267 16673 41535 16681
tri 41535 16673 41543 16681 sw
tri 41267 16665 41275 16673 ne
rect 41275 16665 41543 16673
tri 41543 16665 41551 16673 sw
tri 41275 16657 41283 16665 ne
rect 41283 16657 41551 16665
tri 41551 16657 41559 16665 sw
tri 41283 16649 41291 16657 ne
rect 41291 16649 41559 16657
tri 41559 16649 41567 16657 sw
tri 41291 16641 41299 16649 ne
rect 41299 16641 41567 16649
tri 41567 16641 41575 16649 sw
tri 41299 16633 41307 16641 ne
rect 41307 16633 41575 16641
tri 41575 16633 41583 16641 sw
tri 41307 16625 41315 16633 ne
rect 41315 16625 41583 16633
tri 41583 16625 41591 16633 sw
tri 41315 16617 41323 16625 ne
rect 41323 16617 41591 16625
tri 41591 16617 41599 16625 sw
tri 41323 16609 41331 16617 ne
rect 41331 16609 41599 16617
tri 41599 16609 41607 16617 sw
tri 41331 16601 41339 16609 ne
rect 41339 16601 41607 16609
tri 41607 16601 41615 16609 sw
tri 41339 16593 41347 16601 ne
rect 41347 16593 41615 16601
tri 41615 16593 41623 16601 sw
tri 41347 16585 41355 16593 ne
rect 41355 16585 41623 16593
tri 41623 16585 41631 16593 sw
tri 41355 16577 41363 16585 ne
rect 41363 16577 41631 16585
tri 41631 16577 41639 16585 sw
tri 41363 16569 41371 16577 ne
rect 41371 16569 41639 16577
tri 41639 16569 41647 16577 sw
tri 41371 16561 41379 16569 ne
rect 41379 16561 41647 16569
tri 41647 16561 41655 16569 sw
tri 41379 16553 41387 16561 ne
rect 41387 16553 41655 16561
tri 41655 16553 41663 16561 sw
tri 41387 16545 41395 16553 ne
rect 41395 16545 41663 16553
tri 41663 16545 41671 16553 sw
tri 41395 16541 41399 16545 ne
rect 41399 16541 41671 16545
tri 41399 16533 41407 16541 ne
rect 41407 16537 41671 16541
tri 41671 16537 41679 16545 sw
rect 41407 16533 41679 16537
tri 41407 16525 41415 16533 ne
rect 41415 16529 41679 16533
tri 41679 16529 41687 16537 sw
rect 41415 16525 41687 16529
tri 41415 16517 41423 16525 ne
rect 41423 16521 41687 16525
tri 41687 16521 41695 16529 sw
rect 41423 16517 41695 16521
tri 41423 16509 41431 16517 ne
rect 41431 16513 41695 16517
tri 41695 16513 41703 16521 sw
rect 41431 16509 41703 16513
tri 41431 16501 41439 16509 ne
rect 41439 16505 41703 16509
tri 41703 16505 41711 16513 sw
rect 41439 16501 41711 16505
tri 41439 16493 41447 16501 ne
rect 41447 16497 41711 16501
tri 41711 16497 41719 16505 sw
rect 41447 16493 41719 16497
tri 41447 16485 41455 16493 ne
rect 41455 16489 41719 16493
tri 41719 16489 41727 16497 sw
rect 41455 16485 41727 16489
tri 41455 16477 41463 16485 ne
rect 41463 16481 41727 16485
tri 41727 16481 41735 16489 sw
rect 41463 16477 41735 16481
tri 41463 16469 41471 16477 ne
rect 41471 16473 41735 16477
tri 41735 16473 41743 16481 sw
rect 41471 16469 41743 16473
tri 41471 16461 41479 16469 ne
rect 41479 16465 41743 16469
tri 41743 16465 41751 16473 sw
rect 41479 16461 41751 16465
tri 41479 16453 41487 16461 ne
rect 41487 16457 41751 16461
tri 41751 16457 41759 16465 sw
rect 41487 16453 41759 16457
tri 41487 16445 41495 16453 ne
rect 41495 16449 41759 16453
tri 41759 16449 41767 16457 sw
rect 41495 16445 41767 16449
tri 41495 16437 41503 16445 ne
rect 41503 16441 41767 16445
tri 41767 16441 41775 16449 sw
rect 41503 16437 41775 16441
tri 41503 16429 41511 16437 ne
rect 41511 16433 41775 16437
tri 41775 16433 41783 16441 sw
rect 41511 16429 41783 16433
tri 41511 16421 41519 16429 ne
rect 41519 16425 41783 16429
tri 41783 16425 41791 16433 sw
rect 41519 16421 41791 16425
tri 41519 16413 41527 16421 ne
rect 41527 16417 41791 16421
tri 41791 16417 41799 16425 sw
rect 41527 16413 41799 16417
tri 41527 16409 41531 16413 ne
rect 41531 16409 41799 16413
tri 41799 16409 41807 16417 sw
tri 41531 16405 41535 16409 ne
rect 41535 16405 41807 16409
tri 41807 16405 41811 16409 sw
tri 41535 16397 41543 16405 ne
rect 41543 16397 41811 16405
tri 41811 16397 41819 16405 sw
tri 41543 16389 41551 16397 ne
rect 41551 16389 41819 16397
tri 41819 16389 41827 16397 sw
tri 41551 16381 41559 16389 ne
rect 41559 16381 41827 16389
tri 41827 16381 41835 16389 sw
tri 41559 16373 41567 16381 ne
rect 41567 16373 41835 16381
tri 41835 16373 41843 16381 sw
tri 41567 16365 41575 16373 ne
rect 41575 16365 41843 16373
tri 41843 16365 41851 16373 sw
tri 41575 16357 41583 16365 ne
rect 41583 16357 41851 16365
tri 41851 16357 41859 16365 sw
tri 41583 16349 41591 16357 ne
rect 41591 16349 41859 16357
tri 41859 16349 41867 16357 sw
tri 41591 16341 41599 16349 ne
rect 41599 16341 41867 16349
tri 41867 16341 41875 16349 sw
tri 41599 16333 41607 16341 ne
rect 41607 16333 41875 16341
tri 41875 16333 41883 16341 sw
tri 41607 16325 41615 16333 ne
rect 41615 16325 41883 16333
tri 41883 16325 41891 16333 sw
tri 41615 16317 41623 16325 ne
rect 41623 16317 41891 16325
tri 41891 16317 41899 16325 sw
tri 41623 16309 41631 16317 ne
rect 41631 16309 41899 16317
tri 41899 16309 41907 16317 sw
tri 41631 16301 41639 16309 ne
rect 41639 16301 41907 16309
tri 41907 16301 41915 16309 sw
tri 41639 16293 41647 16301 ne
rect 41647 16293 41915 16301
tri 41915 16293 41923 16301 sw
tri 41647 16285 41655 16293 ne
rect 41655 16285 41923 16293
tri 41923 16285 41931 16293 sw
tri 41655 16277 41663 16285 ne
rect 41663 16277 41931 16285
tri 41931 16277 41939 16285 sw
tri 41663 16269 41671 16277 ne
rect 41671 16269 41939 16277
tri 41939 16269 41947 16277 sw
tri 41671 16265 41675 16269 ne
rect 41675 16265 41947 16269
tri 41675 16257 41683 16265 ne
rect 41683 16261 41947 16265
tri 41947 16261 41955 16269 sw
rect 41683 16257 41955 16261
tri 41683 16249 41691 16257 ne
rect 41691 16253 41955 16257
tri 41955 16253 41963 16261 sw
rect 41691 16249 41963 16253
tri 41691 16241 41699 16249 ne
rect 41699 16245 41963 16249
tri 41963 16245 41971 16253 sw
rect 41699 16241 41971 16245
tri 41699 16233 41707 16241 ne
rect 41707 16237 41971 16241
tri 41971 16237 41979 16245 sw
rect 41707 16233 41979 16237
tri 41707 16225 41715 16233 ne
rect 41715 16229 41979 16233
tri 41979 16229 41987 16237 sw
rect 41715 16225 41987 16229
tri 41715 16217 41723 16225 ne
rect 41723 16221 41987 16225
tri 41987 16221 41995 16229 sw
rect 41723 16217 41995 16221
tri 41723 16209 41731 16217 ne
rect 41731 16213 41995 16217
tri 41995 16213 42003 16221 sw
rect 41731 16209 42003 16213
tri 41731 16201 41739 16209 ne
rect 41739 16205 42003 16209
tri 42003 16205 42011 16213 sw
rect 41739 16201 42011 16205
tri 41739 16193 41747 16201 ne
rect 41747 16197 42011 16201
tri 42011 16197 42019 16205 sw
rect 41747 16193 42019 16197
tri 41747 16185 41755 16193 ne
rect 41755 16189 42019 16193
tri 42019 16189 42027 16197 sw
rect 41755 16185 42027 16189
tri 41755 16177 41763 16185 ne
rect 41763 16181 42027 16185
tri 42027 16181 42035 16189 sw
rect 41763 16177 42035 16181
tri 41763 16169 41771 16177 ne
rect 41771 16173 42035 16177
tri 42035 16173 42043 16181 sw
rect 41771 16169 42043 16173
tri 41771 16161 41779 16169 ne
rect 41779 16165 42043 16169
tri 42043 16165 42051 16173 sw
rect 41779 16161 42051 16165
tri 41779 16153 41787 16161 ne
rect 41787 16157 42051 16161
tri 42051 16157 42059 16165 sw
rect 41787 16153 42059 16157
tri 41787 16145 41795 16153 ne
rect 41795 16149 42059 16153
tri 42059 16149 42067 16157 sw
rect 41795 16145 42067 16149
tri 41795 16137 41803 16145 ne
rect 41803 16141 42067 16145
tri 42067 16141 42075 16149 sw
rect 41803 16137 42075 16141
tri 41803 16133 41807 16137 ne
rect 41807 16133 42075 16137
tri 42075 16133 42083 16141 sw
tri 41807 16129 41811 16133 ne
rect 41811 16129 42083 16133
tri 42083 16129 42087 16133 sw
tri 41811 16121 41819 16129 ne
rect 41819 16121 42087 16129
tri 42087 16121 42095 16129 sw
tri 41819 16113 41827 16121 ne
rect 41827 16113 42095 16121
tri 42095 16113 42103 16121 sw
tri 41827 16105 41835 16113 ne
rect 41835 16105 42103 16113
tri 42103 16105 42111 16113 sw
tri 41835 16097 41843 16105 ne
rect 41843 16097 42111 16105
tri 42111 16097 42119 16105 sw
tri 41843 16089 41851 16097 ne
rect 41851 16089 42119 16097
tri 42119 16089 42127 16097 sw
tri 41851 16081 41859 16089 ne
rect 41859 16081 42127 16089
tri 42127 16081 42135 16089 sw
tri 41859 16073 41867 16081 ne
rect 41867 16073 42135 16081
tri 42135 16073 42143 16081 sw
tri 41867 16065 41875 16073 ne
rect 41875 16065 42143 16073
tri 42143 16065 42151 16073 sw
tri 41875 16057 41883 16065 ne
rect 41883 16057 42151 16065
tri 42151 16057 42159 16065 sw
tri 41883 16049 41891 16057 ne
rect 41891 16049 42159 16057
tri 42159 16049 42167 16057 sw
tri 41891 16041 41899 16049 ne
rect 41899 16041 42167 16049
tri 42167 16041 42175 16049 sw
tri 41899 16033 41907 16041 ne
rect 41907 16033 42175 16041
tri 42175 16033 42183 16041 sw
tri 41907 16025 41915 16033 ne
rect 41915 16025 42183 16033
tri 42183 16025 42191 16033 sw
tri 41915 16017 41923 16025 ne
rect 41923 16017 42191 16025
tri 42191 16017 42199 16025 sw
tri 41923 16009 41931 16017 ne
rect 41931 16009 42199 16017
tri 42199 16009 42207 16017 sw
tri 41931 16001 41939 16009 ne
rect 41939 16001 42207 16009
tri 42207 16001 42215 16009 sw
tri 41939 15993 41947 16001 ne
rect 41947 15993 42215 16001
tri 42215 15993 42223 16001 sw
tri 41947 15989 41951 15993 ne
rect 41951 15989 42223 15993
tri 41951 15981 41959 15989 ne
rect 41959 15985 42223 15989
tri 42223 15985 42231 15993 sw
rect 41959 15981 42231 15985
tri 41959 15973 41967 15981 ne
rect 41967 15977 42231 15981
tri 42231 15977 42239 15985 sw
rect 41967 15973 42239 15977
tri 41967 15965 41975 15973 ne
rect 41975 15969 42239 15973
tri 42239 15969 42247 15977 sw
rect 41975 15965 42247 15969
tri 41975 15957 41983 15965 ne
rect 41983 15961 42247 15965
tri 42247 15961 42255 15969 sw
rect 41983 15957 42255 15961
tri 41983 15949 41991 15957 ne
rect 41991 15953 42255 15957
tri 42255 15953 42263 15961 sw
rect 41991 15949 42263 15953
tri 41991 15941 41999 15949 ne
rect 41999 15945 42263 15949
tri 42263 15945 42271 15953 sw
rect 41999 15941 42271 15945
tri 41999 15933 42007 15941 ne
rect 42007 15937 42271 15941
tri 42271 15937 42279 15945 sw
rect 42007 15933 42279 15937
tri 42007 15925 42015 15933 ne
rect 42015 15929 42279 15933
tri 42279 15929 42287 15937 sw
rect 42015 15925 42287 15929
tri 42015 15917 42023 15925 ne
rect 42023 15921 42287 15925
tri 42287 15921 42295 15929 sw
rect 42023 15917 42295 15921
tri 42023 15909 42031 15917 ne
rect 42031 15913 42295 15917
tri 42295 15913 42303 15921 sw
rect 42031 15909 42303 15913
tri 42031 15901 42039 15909 ne
rect 42039 15905 42303 15909
tri 42303 15905 42311 15913 sw
rect 42039 15901 42311 15905
tri 42039 15893 42047 15901 ne
rect 42047 15897 42311 15901
tri 42311 15897 42319 15905 sw
rect 42047 15893 42319 15897
tri 42047 15885 42055 15893 ne
rect 42055 15889 42319 15893
tri 42319 15889 42327 15897 sw
rect 42055 15885 42327 15889
tri 42055 15877 42063 15885 ne
rect 42063 15881 42327 15885
tri 42327 15881 42335 15889 sw
rect 42063 15877 42335 15881
tri 42063 15869 42071 15877 ne
rect 42071 15873 42335 15877
tri 42335 15873 42343 15881 sw
rect 42071 15869 42343 15873
tri 42071 15861 42079 15869 ne
rect 42079 15865 42343 15869
tri 42343 15865 42351 15873 sw
rect 42079 15861 42351 15865
tri 42079 15857 42083 15861 ne
rect 42083 15857 42351 15861
tri 42351 15857 42359 15865 sw
tri 42083 15853 42087 15857 ne
rect 42087 15853 42359 15857
tri 42359 15853 42363 15857 sw
tri 42087 15845 42095 15853 ne
rect 42095 15845 42363 15853
tri 42363 15845 42371 15853 sw
tri 42095 15837 42103 15845 ne
rect 42103 15837 42371 15845
tri 42371 15837 42379 15845 sw
tri 42103 15829 42111 15837 ne
rect 42111 15829 42379 15837
tri 42379 15829 42387 15837 sw
tri 42111 15821 42119 15829 ne
rect 42119 15821 42387 15829
tri 42387 15821 42395 15829 sw
tri 42119 15813 42127 15821 ne
rect 42127 15813 42395 15821
tri 42395 15813 42403 15821 sw
tri 42127 15805 42135 15813 ne
rect 42135 15805 42403 15813
tri 42403 15805 42411 15813 sw
tri 42135 15797 42143 15805 ne
rect 42143 15797 42411 15805
tri 42411 15797 42419 15805 sw
tri 42143 15789 42151 15797 ne
rect 42151 15789 42419 15797
tri 42419 15789 42427 15797 sw
tri 42151 15781 42159 15789 ne
rect 42159 15781 42427 15789
tri 42427 15781 42435 15789 sw
tri 42159 15773 42167 15781 ne
rect 42167 15773 42435 15781
tri 42435 15773 42443 15781 sw
tri 42167 15765 42175 15773 ne
rect 42175 15765 42443 15773
tri 42443 15765 42451 15773 sw
tri 42175 15757 42183 15765 ne
rect 42183 15757 42451 15765
tri 42451 15757 42459 15765 sw
tri 42183 15749 42191 15757 ne
rect 42191 15749 42459 15757
tri 42459 15749 42467 15757 sw
tri 42191 15741 42199 15749 ne
rect 42199 15741 42467 15749
tri 42467 15741 42475 15749 sw
tri 42199 15733 42207 15741 ne
rect 42207 15733 42475 15741
tri 42475 15733 42483 15741 sw
tri 42207 15725 42215 15733 ne
rect 42215 15725 42483 15733
tri 42483 15725 42491 15733 sw
tri 42215 15717 42223 15725 ne
rect 42223 15717 42491 15725
tri 42491 15717 42499 15725 sw
tri 42223 15713 42227 15717 ne
rect 42227 15713 42499 15717
tri 42227 15705 42235 15713 ne
rect 42235 15709 42499 15713
tri 42499 15709 42507 15717 sw
rect 42235 15705 42507 15709
tri 42235 15697 42243 15705 ne
rect 42243 15701 42507 15705
tri 42507 15701 42515 15709 sw
rect 42243 15697 42515 15701
tri 42243 15689 42251 15697 ne
rect 42251 15693 42515 15697
tri 42515 15693 42523 15701 sw
rect 42251 15689 42523 15693
tri 42251 15681 42259 15689 ne
rect 42259 15685 42523 15689
tri 42523 15685 42531 15693 sw
rect 42259 15681 42531 15685
tri 42259 15673 42267 15681 ne
rect 42267 15677 42531 15681
tri 42531 15677 42539 15685 sw
rect 42267 15673 42539 15677
tri 42267 15665 42275 15673 ne
rect 42275 15669 42539 15673
tri 42539 15669 42547 15677 sw
rect 42275 15665 42547 15669
tri 42275 15657 42283 15665 ne
rect 42283 15661 42547 15665
tri 42547 15661 42555 15669 sw
rect 42283 15657 42555 15661
tri 42283 15649 42291 15657 ne
rect 42291 15653 42555 15657
tri 42555 15653 42563 15661 sw
rect 42291 15649 42563 15653
tri 42291 15641 42299 15649 ne
rect 42299 15645 42563 15649
tri 42563 15645 42571 15653 sw
rect 42299 15641 42571 15645
tri 42299 15633 42307 15641 ne
rect 42307 15637 42571 15641
tri 42571 15637 42579 15645 sw
rect 42307 15633 42579 15637
tri 42307 15625 42315 15633 ne
rect 42315 15629 42579 15633
tri 42579 15629 42587 15637 sw
rect 42315 15625 42587 15629
tri 42315 15617 42323 15625 ne
rect 42323 15621 42587 15625
tri 42587 15621 42595 15629 sw
rect 42323 15617 42595 15621
tri 42323 15609 42331 15617 ne
rect 42331 15613 42595 15617
tri 42595 15613 42603 15621 sw
rect 42331 15609 42603 15613
tri 42331 15601 42339 15609 ne
rect 42339 15605 42603 15609
tri 42603 15605 42611 15613 sw
rect 42339 15601 42611 15605
tri 42339 15593 42347 15601 ne
rect 42347 15597 42611 15601
tri 42611 15597 42619 15605 sw
rect 42347 15593 42619 15597
tri 42347 15585 42355 15593 ne
rect 42355 15589 42619 15593
tri 42619 15589 42627 15597 sw
rect 42355 15585 42627 15589
tri 42355 15581 42359 15585 ne
rect 42359 15581 42627 15585
tri 42627 15581 42635 15589 sw
tri 42359 15577 42363 15581 ne
rect 42363 15577 42635 15581
tri 42635 15577 42639 15581 sw
tri 42363 15569 42371 15577 ne
rect 42371 15569 42639 15577
tri 42639 15569 42647 15577 sw
tri 42371 15561 42379 15569 ne
rect 42379 15561 42647 15569
tri 42647 15561 42655 15569 sw
tri 42379 15553 42387 15561 ne
rect 42387 15553 42655 15561
tri 42655 15553 42663 15561 sw
tri 42387 15545 42395 15553 ne
rect 42395 15545 42663 15553
tri 42663 15545 42671 15553 sw
tri 42395 15537 42403 15545 ne
rect 42403 15537 42671 15545
tri 42671 15537 42679 15545 sw
tri 42403 15529 42411 15537 ne
rect 42411 15529 42679 15537
tri 42679 15529 42687 15537 sw
tri 42411 15521 42419 15529 ne
rect 42419 15521 42687 15529
tri 42687 15521 42695 15529 sw
tri 42419 15513 42427 15521 ne
rect 42427 15513 42695 15521
tri 42695 15513 42703 15521 sw
tri 42427 15505 42435 15513 ne
rect 42435 15505 42703 15513
tri 42703 15505 42711 15513 sw
tri 42435 15497 42443 15505 ne
rect 42443 15497 42711 15505
tri 42711 15497 42719 15505 sw
tri 42443 15489 42451 15497 ne
rect 42451 15489 42719 15497
tri 42719 15489 42727 15497 sw
tri 42451 15481 42459 15489 ne
rect 42459 15481 42727 15489
tri 42727 15481 42735 15489 sw
tri 42459 15473 42467 15481 ne
rect 42467 15473 42735 15481
tri 42735 15473 42743 15481 sw
tri 42467 15465 42475 15473 ne
rect 42475 15465 42743 15473
tri 42743 15465 42751 15473 sw
tri 42475 15457 42483 15465 ne
rect 42483 15457 42751 15465
tri 42751 15457 42759 15465 sw
tri 42483 15449 42491 15457 ne
rect 42491 15449 42759 15457
tri 42759 15449 42767 15457 sw
tri 42491 15441 42499 15449 ne
rect 42499 15441 42767 15449
tri 42767 15441 42775 15449 sw
tri 42499 15437 42503 15441 ne
rect 42503 15437 42775 15441
tri 42503 15429 42511 15437 ne
rect 42511 15433 42775 15437
tri 42775 15433 42783 15441 sw
rect 42511 15429 42783 15433
tri 42511 15421 42519 15429 ne
rect 42519 15425 42783 15429
tri 42783 15425 42791 15433 sw
rect 42519 15421 42791 15425
tri 42519 15413 42527 15421 ne
rect 42527 15417 42791 15421
tri 42791 15417 42799 15425 sw
rect 42527 15413 42799 15417
tri 42527 15405 42535 15413 ne
rect 42535 15409 42799 15413
tri 42799 15409 42807 15417 sw
rect 42535 15405 42807 15409
tri 42535 15397 42543 15405 ne
rect 42543 15401 42807 15405
tri 42807 15401 42815 15409 sw
rect 42543 15397 42815 15401
tri 42543 15389 42551 15397 ne
rect 42551 15393 42815 15397
tri 42815 15393 42823 15401 sw
rect 42551 15389 42823 15393
tri 42551 15381 42559 15389 ne
rect 42559 15385 42823 15389
tri 42823 15385 42831 15393 sw
rect 42559 15381 42831 15385
tri 42559 15373 42567 15381 ne
rect 42567 15377 42831 15381
tri 42831 15377 42839 15385 sw
rect 42567 15373 42839 15377
tri 42567 15365 42575 15373 ne
rect 42575 15369 42839 15373
tri 42839 15369 42847 15377 sw
rect 42575 15365 42847 15369
tri 42575 15357 42583 15365 ne
rect 42583 15361 42847 15365
tri 42847 15361 42855 15369 sw
rect 42583 15357 42855 15361
tri 42583 15349 42591 15357 ne
rect 42591 15353 42855 15357
tri 42855 15353 42863 15361 sw
rect 42591 15349 42863 15353
tri 42591 15341 42599 15349 ne
rect 42599 15345 42863 15349
tri 42863 15345 42871 15353 sw
rect 42599 15341 42871 15345
tri 42599 15333 42607 15341 ne
rect 42607 15337 42871 15341
tri 42871 15337 42879 15345 sw
rect 42607 15333 42879 15337
tri 42607 15325 42615 15333 ne
rect 42615 15329 42879 15333
tri 42879 15329 42887 15337 sw
rect 42615 15325 42887 15329
tri 42615 15317 42623 15325 ne
rect 42623 15321 42887 15325
tri 42887 15321 42895 15329 sw
rect 42623 15317 42895 15321
tri 42623 15309 42631 15317 ne
rect 42631 15313 42895 15317
tri 42895 15313 42903 15321 sw
rect 42631 15309 42903 15313
tri 42631 15305 42635 15309 ne
rect 42635 15305 42903 15309
tri 42903 15305 42911 15313 sw
tri 42635 15301 42639 15305 ne
rect 42639 15301 42911 15305
tri 42911 15301 42915 15305 sw
tri 42639 15293 42647 15301 ne
rect 42647 15293 42915 15301
tri 42915 15293 42923 15301 sw
tri 42647 15285 42655 15293 ne
rect 42655 15285 42923 15293
tri 42923 15285 42931 15293 sw
tri 42655 15277 42663 15285 ne
rect 42663 15277 42931 15285
tri 42931 15277 42939 15285 sw
tri 42663 15269 42671 15277 ne
rect 42671 15269 42939 15277
tri 42939 15269 42947 15277 sw
tri 42671 15261 42679 15269 ne
rect 42679 15261 42947 15269
tri 42947 15261 42955 15269 sw
tri 42679 15253 42687 15261 ne
rect 42687 15253 42955 15261
tri 42955 15253 42963 15261 sw
tri 42687 15245 42695 15253 ne
rect 42695 15245 42963 15253
tri 42963 15245 42971 15253 sw
tri 42695 15237 42703 15245 ne
rect 42703 15237 42971 15245
tri 42971 15237 42979 15245 sw
tri 42703 15229 42711 15237 ne
rect 42711 15229 42979 15237
tri 42979 15229 42987 15237 sw
tri 42711 15221 42719 15229 ne
rect 42719 15221 42987 15229
tri 42987 15221 42995 15229 sw
tri 42719 15213 42727 15221 ne
rect 42727 15213 42995 15221
tri 42995 15213 43003 15221 sw
tri 42727 15205 42735 15213 ne
rect 42735 15205 43003 15213
tri 43003 15205 43011 15213 sw
tri 42735 15197 42743 15205 ne
rect 42743 15197 43011 15205
tri 43011 15197 43019 15205 sw
tri 42743 15189 42751 15197 ne
rect 42751 15189 43019 15197
tri 43019 15189 43027 15197 sw
tri 42751 15181 42759 15189 ne
rect 42759 15181 43027 15189
tri 43027 15181 43035 15189 sw
tri 42759 15173 42767 15181 ne
rect 42767 15173 43035 15181
tri 43035 15173 43043 15181 sw
tri 42767 15165 42775 15173 ne
rect 42775 15165 43043 15173
tri 43043 15165 43051 15173 sw
tri 42775 15161 42779 15165 ne
rect 42779 15161 43051 15165
tri 42779 15153 42787 15161 ne
rect 42787 15157 43051 15161
tri 43051 15157 43059 15165 sw
rect 42787 15153 43059 15157
tri 42787 15145 42795 15153 ne
rect 42795 15149 43059 15153
tri 43059 15149 43067 15157 sw
rect 42795 15145 43067 15149
tri 42795 15137 42803 15145 ne
rect 42803 15141 43067 15145
tri 43067 15141 43075 15149 sw
rect 42803 15137 43075 15141
tri 42803 15129 42811 15137 ne
rect 42811 15133 43075 15137
tri 43075 15133 43083 15141 sw
rect 42811 15129 43083 15133
tri 42811 15121 42819 15129 ne
rect 42819 15125 43083 15129
tri 43083 15125 43091 15133 sw
rect 42819 15121 43091 15125
tri 42819 15113 42827 15121 ne
rect 42827 15117 43091 15121
tri 43091 15117 43099 15125 sw
rect 42827 15113 43099 15117
tri 42827 15105 42835 15113 ne
rect 42835 15109 43099 15113
tri 43099 15109 43107 15117 sw
rect 42835 15105 43107 15109
tri 42835 15097 42843 15105 ne
rect 42843 15101 43107 15105
tri 43107 15101 43115 15109 sw
rect 42843 15097 43115 15101
tri 42843 15089 42851 15097 ne
rect 42851 15093 43115 15097
tri 43115 15093 43123 15101 sw
rect 42851 15089 43123 15093
tri 42851 15081 42859 15089 ne
rect 42859 15085 43123 15089
tri 43123 15085 43131 15093 sw
rect 42859 15081 43131 15085
tri 42859 15073 42867 15081 ne
rect 42867 15077 43131 15081
tri 43131 15077 43139 15085 sw
rect 42867 15073 43139 15077
tri 42867 15065 42875 15073 ne
rect 42875 15069 43139 15073
tri 43139 15069 43147 15077 sw
rect 42875 15065 43147 15069
tri 42875 15057 42883 15065 ne
rect 42883 15061 43147 15065
tri 43147 15061 43155 15069 sw
rect 42883 15057 43155 15061
tri 42883 15049 42891 15057 ne
rect 42891 15053 43155 15057
tri 43155 15053 43163 15061 sw
rect 42891 15049 43163 15053
tri 42891 15041 42899 15049 ne
rect 42899 15045 43163 15049
tri 43163 15045 43171 15053 sw
rect 42899 15041 43171 15045
tri 42899 15033 42907 15041 ne
rect 42907 15037 43171 15041
tri 43171 15037 43179 15045 sw
rect 42907 15033 43179 15037
tri 42907 15029 42911 15033 ne
rect 42911 15029 43179 15033
tri 43179 15029 43187 15037 sw
tri 42911 15025 42915 15029 ne
rect 42915 15025 43187 15029
tri 43187 15025 43191 15029 sw
tri 42915 15017 42923 15025 ne
rect 42923 15017 43191 15025
tri 43191 15017 43199 15025 sw
tri 42923 15009 42931 15017 ne
rect 42931 15009 43199 15017
tri 43199 15009 43207 15017 sw
tri 42931 15001 42939 15009 ne
rect 42939 15001 43207 15009
tri 43207 15001 43215 15009 sw
tri 42939 14993 42947 15001 ne
rect 42947 14993 43215 15001
tri 43215 14993 43223 15001 sw
tri 42947 14985 42955 14993 ne
rect 42955 14985 43223 14993
tri 43223 14985 43231 14993 sw
tri 42955 14977 42963 14985 ne
rect 42963 14977 43231 14985
tri 43231 14977 43239 14985 sw
tri 42963 14969 42971 14977 ne
rect 42971 14969 43239 14977
tri 43239 14969 43247 14977 sw
tri 42971 14961 42979 14969 ne
rect 42979 14961 43247 14969
tri 43247 14961 43255 14969 sw
tri 42979 14953 42987 14961 ne
rect 42987 14953 43255 14961
tri 43255 14953 43263 14961 sw
tri 42987 14945 42995 14953 ne
rect 42995 14945 43263 14953
tri 43263 14945 43271 14953 sw
tri 42995 14937 43003 14945 ne
rect 43003 14937 43271 14945
tri 43271 14937 43279 14945 sw
tri 43003 14929 43011 14937 ne
rect 43011 14929 43279 14937
tri 43279 14929 43287 14937 sw
tri 43011 14921 43019 14929 ne
rect 43019 14921 43287 14929
tri 43287 14921 43295 14929 sw
tri 43019 14913 43027 14921 ne
rect 43027 14913 43295 14921
tri 43295 14913 43303 14921 sw
tri 43027 14905 43035 14913 ne
rect 43035 14905 43303 14913
tri 43303 14905 43311 14913 sw
tri 43035 14897 43043 14905 ne
rect 43043 14897 43311 14905
tri 43311 14897 43319 14905 sw
tri 43043 14889 43051 14897 ne
rect 43051 14889 43319 14897
tri 43319 14889 43327 14897 sw
tri 43051 14885 43055 14889 ne
rect 43055 14885 43327 14889
tri 43055 14877 43063 14885 ne
rect 43063 14881 43327 14885
tri 43327 14881 43335 14889 sw
rect 43063 14877 43335 14881
tri 43063 14869 43071 14877 ne
rect 43071 14873 43335 14877
tri 43335 14873 43343 14881 sw
rect 43071 14869 43343 14873
tri 43071 14861 43079 14869 ne
rect 43079 14865 43343 14869
tri 43343 14865 43351 14873 sw
rect 43079 14861 43351 14865
tri 43079 14853 43087 14861 ne
rect 43087 14857 43351 14861
tri 43351 14857 43359 14865 sw
rect 43087 14853 43359 14857
tri 43087 14845 43095 14853 ne
rect 43095 14849 43359 14853
tri 43359 14849 43367 14857 sw
rect 43095 14845 43367 14849
tri 43095 14837 43103 14845 ne
rect 43103 14841 43367 14845
tri 43367 14841 43375 14849 sw
rect 43103 14837 43375 14841
tri 43103 14829 43111 14837 ne
rect 43111 14833 43375 14837
tri 43375 14833 43383 14841 sw
rect 43111 14829 43383 14833
tri 43111 14821 43119 14829 ne
rect 43119 14825 43383 14829
tri 43383 14825 43391 14833 sw
rect 43119 14821 43391 14825
tri 43119 14813 43127 14821 ne
rect 43127 14817 43391 14821
tri 43391 14817 43399 14825 sw
rect 43127 14813 43399 14817
tri 43127 14805 43135 14813 ne
rect 43135 14809 43399 14813
tri 43399 14809 43407 14817 sw
rect 43135 14805 43407 14809
tri 43135 14797 43143 14805 ne
rect 43143 14801 43407 14805
tri 43407 14801 43415 14809 sw
rect 43143 14797 43415 14801
tri 43143 14789 43151 14797 ne
rect 43151 14793 43415 14797
tri 43415 14793 43423 14801 sw
rect 43151 14789 43423 14793
tri 43151 14781 43159 14789 ne
rect 43159 14785 43423 14789
tri 43423 14785 43431 14793 sw
rect 43159 14781 43431 14785
tri 43159 14773 43167 14781 ne
rect 43167 14777 43431 14781
tri 43431 14777 43439 14785 sw
rect 43167 14773 43439 14777
tri 43167 14765 43175 14773 ne
rect 43175 14769 43439 14773
tri 43439 14769 43447 14777 sw
rect 43175 14765 43447 14769
tri 43175 14757 43183 14765 ne
rect 43183 14761 43447 14765
tri 43447 14761 43455 14769 sw
rect 43183 14757 43455 14761
tri 43183 14753 43187 14757 ne
rect 43187 14753 43455 14757
tri 43455 14753 43463 14761 sw
tri 43187 14749 43191 14753 ne
rect 43191 14749 43463 14753
tri 43463 14749 43467 14753 sw
tri 43191 14741 43199 14749 ne
rect 43199 14741 43467 14749
tri 43467 14741 43475 14749 sw
tri 43199 14733 43207 14741 ne
rect 43207 14733 43475 14741
tri 43475 14733 43483 14741 sw
tri 43207 14725 43215 14733 ne
rect 43215 14725 43483 14733
tri 43483 14725 43491 14733 sw
tri 43215 14717 43223 14725 ne
rect 43223 14717 43491 14725
tri 43491 14717 43499 14725 sw
tri 43223 14709 43231 14717 ne
rect 43231 14709 43499 14717
tri 43499 14709 43507 14717 sw
tri 43231 14701 43239 14709 ne
rect 43239 14701 43507 14709
tri 43507 14701 43515 14709 sw
tri 43239 14693 43247 14701 ne
rect 43247 14693 43515 14701
tri 43515 14693 43523 14701 sw
tri 43247 14685 43255 14693 ne
rect 43255 14685 43523 14693
tri 43523 14685 43531 14693 sw
tri 43255 14677 43263 14685 ne
rect 43263 14677 43531 14685
tri 43531 14677 43539 14685 sw
tri 43263 14669 43271 14677 ne
rect 43271 14669 43539 14677
tri 43539 14669 43547 14677 sw
tri 43271 14661 43279 14669 ne
rect 43279 14661 43547 14669
tri 43547 14661 43555 14669 sw
tri 43279 14653 43287 14661 ne
rect 43287 14653 43555 14661
tri 43555 14653 43563 14661 sw
tri 43287 14645 43295 14653 ne
rect 43295 14645 43563 14653
tri 43563 14645 43571 14653 sw
tri 43295 14637 43303 14645 ne
rect 43303 14637 43571 14645
tri 43571 14637 43579 14645 sw
tri 43303 14629 43311 14637 ne
rect 43311 14629 43579 14637
tri 43579 14629 43587 14637 sw
tri 43311 14621 43319 14629 ne
rect 43319 14621 43587 14629
tri 43587 14621 43595 14629 sw
tri 43319 14613 43327 14621 ne
rect 43327 14613 43595 14621
tri 43595 14613 43603 14621 sw
tri 43327 14609 43331 14613 ne
rect 43331 14609 43603 14613
tri 43331 14601 43339 14609 ne
rect 43339 14605 43603 14609
tri 43603 14605 43611 14613 sw
rect 43339 14601 43611 14605
tri 43339 14593 43347 14601 ne
rect 43347 14597 43611 14601
tri 43611 14597 43619 14605 sw
rect 43347 14593 43619 14597
tri 43347 14585 43355 14593 ne
rect 43355 14589 43619 14593
tri 43619 14589 43627 14597 sw
rect 43355 14585 43627 14589
tri 43355 14577 43363 14585 ne
rect 43363 14581 43627 14585
tri 43627 14581 43635 14589 sw
rect 43363 14577 43635 14581
tri 43363 14569 43371 14577 ne
rect 43371 14573 43635 14577
tri 43635 14573 43643 14581 sw
rect 43371 14569 43643 14573
tri 43371 14561 43379 14569 ne
rect 43379 14565 43643 14569
tri 43643 14565 43651 14573 sw
rect 43379 14561 43651 14565
tri 43379 14553 43387 14561 ne
rect 43387 14557 43651 14561
tri 43651 14557 43659 14565 sw
rect 43387 14553 43659 14557
tri 43387 14545 43395 14553 ne
rect 43395 14549 43659 14553
tri 43659 14549 43667 14557 sw
rect 43395 14545 43667 14549
tri 43395 14537 43403 14545 ne
rect 43403 14541 43667 14545
tri 43667 14541 43675 14549 sw
rect 43403 14537 43675 14541
tri 43403 14529 43411 14537 ne
rect 43411 14533 43675 14537
tri 43675 14533 43683 14541 sw
rect 43411 14529 43683 14533
tri 43411 14521 43419 14529 ne
rect 43419 14525 43683 14529
tri 43683 14525 43691 14533 sw
rect 43419 14521 43691 14525
tri 43419 14513 43427 14521 ne
rect 43427 14517 43691 14521
tri 43691 14517 43699 14525 sw
rect 43427 14513 43699 14517
tri 43427 14505 43435 14513 ne
rect 43435 14509 43699 14513
tri 43699 14509 43707 14517 sw
rect 43435 14505 43707 14509
tri 43435 14497 43443 14505 ne
rect 43443 14501 43707 14505
tri 43707 14501 43715 14509 sw
rect 43443 14497 43715 14501
tri 43443 14489 43451 14497 ne
rect 43451 14493 43715 14497
tri 43715 14493 43723 14501 sw
rect 43451 14489 43723 14493
tri 43451 14481 43459 14489 ne
rect 43459 14485 43723 14489
tri 43723 14485 43731 14493 sw
rect 43459 14481 43731 14485
tri 43459 14477 43463 14481 ne
rect 43463 14477 43731 14481
tri 43731 14477 43739 14485 sw
tri 43463 14473 43467 14477 ne
rect 43467 14473 43739 14477
tri 43739 14473 43743 14477 sw
tri 43467 14465 43475 14473 ne
rect 43475 14465 43743 14473
tri 43743 14465 43751 14473 sw
tri 43475 14457 43483 14465 ne
rect 43483 14457 43751 14465
tri 43751 14457 43759 14465 sw
tri 43483 14449 43491 14457 ne
rect 43491 14449 43759 14457
tri 43759 14449 43767 14457 sw
tri 43491 14441 43499 14449 ne
rect 43499 14441 43767 14449
tri 43767 14441 43775 14449 sw
tri 43499 14433 43507 14441 ne
rect 43507 14433 43775 14441
tri 43775 14433 43783 14441 sw
tri 43507 14425 43515 14433 ne
rect 43515 14425 43783 14433
tri 43783 14425 43791 14433 sw
tri 43515 14417 43523 14425 ne
rect 43523 14417 43791 14425
tri 43791 14417 43799 14425 sw
tri 43523 14409 43531 14417 ne
rect 43531 14409 43799 14417
tri 43799 14409 43807 14417 sw
tri 43531 14401 43539 14409 ne
rect 43539 14401 43807 14409
tri 43807 14401 43815 14409 sw
tri 43539 14393 43547 14401 ne
rect 43547 14393 43815 14401
tri 43815 14393 43823 14401 sw
tri 43547 14385 43555 14393 ne
rect 43555 14385 43823 14393
tri 43823 14385 43831 14393 sw
tri 43555 14377 43563 14385 ne
rect 43563 14377 43831 14385
tri 43831 14377 43839 14385 sw
tri 43563 14369 43571 14377 ne
rect 43571 14369 43839 14377
tri 43839 14369 43847 14377 sw
tri 43571 14361 43579 14369 ne
rect 43579 14361 43847 14369
tri 43847 14361 43855 14369 sw
tri 43579 14353 43587 14361 ne
rect 43587 14353 43855 14361
tri 43855 14353 43863 14361 sw
tri 43587 14345 43595 14353 ne
rect 43595 14345 43863 14353
tri 43863 14345 43871 14353 sw
tri 43595 14337 43603 14345 ne
rect 43603 14337 43871 14345
tri 43871 14337 43879 14345 sw
tri 43603 14333 43607 14337 ne
rect 43607 14333 43879 14337
tri 43607 14325 43615 14333 ne
rect 43615 14329 43879 14333
tri 43879 14329 43887 14337 sw
rect 43615 14325 43887 14329
tri 43615 14317 43623 14325 ne
rect 43623 14321 43887 14325
tri 43887 14321 43895 14329 sw
rect 43623 14317 43895 14321
tri 43623 14309 43631 14317 ne
rect 43631 14313 43895 14317
tri 43895 14313 43903 14321 sw
rect 43631 14309 43903 14313
tri 43631 14301 43639 14309 ne
rect 43639 14305 43903 14309
tri 43903 14305 43911 14313 sw
rect 43639 14301 43911 14305
tri 43639 14293 43647 14301 ne
rect 43647 14297 43911 14301
tri 43911 14297 43919 14305 sw
rect 43647 14293 43919 14297
tri 43647 14285 43655 14293 ne
rect 43655 14289 43919 14293
tri 43919 14289 43927 14297 sw
rect 43655 14285 43927 14289
tri 43655 14277 43663 14285 ne
rect 43663 14281 43927 14285
tri 43927 14281 43935 14289 sw
rect 43663 14277 43935 14281
tri 43663 14269 43671 14277 ne
rect 43671 14273 43935 14277
tri 43935 14273 43943 14281 sw
rect 43671 14269 43943 14273
tri 43671 14261 43679 14269 ne
rect 43679 14265 43943 14269
tri 43943 14265 43951 14273 sw
rect 43679 14261 43951 14265
tri 43679 14253 43687 14261 ne
rect 43687 14257 43951 14261
tri 43951 14257 43959 14265 sw
rect 43687 14253 43959 14257
tri 43687 14245 43695 14253 ne
rect 43695 14249 43959 14253
tri 43959 14249 43967 14257 sw
rect 43695 14245 43967 14249
tri 43695 14237 43703 14245 ne
rect 43703 14241 43967 14245
tri 43967 14241 43975 14249 sw
rect 43703 14237 43975 14241
tri 43703 14229 43711 14237 ne
rect 43711 14233 43975 14237
tri 43975 14233 43983 14241 sw
rect 43711 14229 43983 14233
tri 43711 14221 43719 14229 ne
rect 43719 14225 43983 14229
tri 43983 14225 43991 14233 sw
rect 43719 14221 43991 14225
tri 43719 14213 43727 14221 ne
rect 43727 14217 43991 14221
tri 43991 14217 43999 14225 sw
rect 43727 14213 43999 14217
tri 43727 14205 43735 14213 ne
rect 43735 14209 43999 14213
tri 43999 14209 44007 14217 sw
rect 43735 14205 44007 14209
tri 43735 14201 43739 14205 ne
rect 43739 14201 44007 14205
tri 44007 14201 44015 14209 sw
tri 43739 14197 43743 14201 ne
rect 43743 14197 44015 14201
tri 44015 14197 44019 14201 sw
tri 43743 14189 43751 14197 ne
rect 43751 14189 44019 14197
tri 44019 14189 44027 14197 sw
tri 43751 14181 43759 14189 ne
rect 43759 14181 44027 14189
tri 44027 14181 44035 14189 sw
tri 43759 14173 43767 14181 ne
rect 43767 14173 44035 14181
tri 44035 14173 44043 14181 sw
tri 43767 14165 43775 14173 ne
rect 43775 14165 44043 14173
tri 44043 14165 44051 14173 sw
tri 43775 14157 43783 14165 ne
rect 43783 14157 44051 14165
tri 44051 14157 44059 14165 sw
tri 43783 14149 43791 14157 ne
rect 43791 14149 44059 14157
tri 44059 14149 44067 14157 sw
tri 43791 14141 43799 14149 ne
rect 43799 14141 44067 14149
tri 44067 14141 44075 14149 sw
tri 43799 14133 43807 14141 ne
rect 43807 14133 44075 14141
tri 44075 14133 44083 14141 sw
tri 43807 14125 43815 14133 ne
rect 43815 14125 44083 14133
tri 44083 14125 44091 14133 sw
tri 43815 14117 43823 14125 ne
rect 43823 14117 44091 14125
tri 44091 14117 44099 14125 sw
tri 43823 14109 43831 14117 ne
rect 43831 14109 44099 14117
tri 44099 14109 44107 14117 sw
tri 43831 14101 43839 14109 ne
rect 43839 14101 44107 14109
tri 44107 14101 44115 14109 sw
tri 43839 14093 43847 14101 ne
rect 43847 14093 44115 14101
tri 44115 14093 44123 14101 sw
tri 43847 14085 43855 14093 ne
rect 43855 14085 44123 14093
tri 44123 14085 44131 14093 sw
tri 43855 14077 43863 14085 ne
rect 43863 14077 44131 14085
tri 44131 14077 44139 14085 sw
tri 43863 14069 43871 14077 ne
rect 43871 14069 44139 14077
tri 44139 14069 44147 14077 sw
tri 43871 14061 43879 14069 ne
rect 43879 14061 44147 14069
tri 44147 14061 44155 14069 sw
tri 43879 14057 43883 14061 ne
rect 43883 14057 44155 14061
tri 43883 14049 43891 14057 ne
rect 43891 14053 44155 14057
tri 44155 14053 44163 14061 sw
rect 43891 14049 44163 14053
tri 43891 14041 43899 14049 ne
rect 43899 14045 44163 14049
tri 44163 14045 44171 14053 sw
rect 43899 14041 44171 14045
tri 43899 14033 43907 14041 ne
rect 43907 14037 44171 14041
tri 44171 14037 44179 14045 sw
rect 43907 14033 44179 14037
tri 43907 14025 43915 14033 ne
rect 43915 14029 44179 14033
tri 44179 14029 44187 14037 sw
rect 43915 14025 44187 14029
tri 43915 14017 43923 14025 ne
rect 43923 14021 44187 14025
tri 44187 14021 44195 14029 sw
rect 43923 14017 44195 14021
tri 43923 14009 43931 14017 ne
rect 43931 14013 44195 14017
tri 44195 14013 44203 14021 sw
rect 43931 14009 44203 14013
tri 43931 14001 43939 14009 ne
rect 43939 14005 44203 14009
tri 44203 14005 44211 14013 sw
rect 43939 14001 44211 14005
tri 43939 13993 43947 14001 ne
rect 43947 13997 44211 14001
tri 44211 13997 44219 14005 sw
rect 43947 13993 44219 13997
tri 43947 13985 43955 13993 ne
rect 43955 13989 44219 13993
tri 44219 13989 44227 13997 sw
rect 43955 13985 44227 13989
tri 43955 13977 43963 13985 ne
rect 43963 13981 44227 13985
tri 44227 13981 44235 13989 sw
rect 43963 13977 44235 13981
tri 43963 13969 43971 13977 ne
rect 43971 13973 44235 13977
tri 44235 13973 44243 13981 sw
rect 43971 13969 44243 13973
tri 43971 13961 43979 13969 ne
rect 43979 13965 44243 13969
tri 44243 13965 44251 13973 sw
rect 43979 13961 44251 13965
tri 43979 13953 43987 13961 ne
rect 43987 13957 44251 13961
tri 44251 13957 44259 13965 sw
rect 43987 13953 44259 13957
tri 43987 13945 43995 13953 ne
rect 43995 13949 44259 13953
tri 44259 13949 44267 13957 sw
rect 43995 13945 44267 13949
tri 43995 13937 44003 13945 ne
rect 44003 13941 44267 13945
tri 44267 13941 44275 13949 sw
rect 44003 13937 44275 13941
tri 44003 13929 44011 13937 ne
rect 44011 13933 44275 13937
tri 44275 13933 44283 13941 sw
rect 44011 13929 44283 13933
tri 44011 13925 44015 13929 ne
rect 44015 13925 44283 13929
tri 44283 13925 44291 13933 sw
tri 44015 13921 44019 13925 ne
rect 44019 13921 44291 13925
tri 44291 13921 44295 13925 sw
tri 44019 13913 44027 13921 ne
rect 44027 13913 44295 13921
tri 44295 13913 44303 13921 sw
tri 44027 13905 44035 13913 ne
rect 44035 13905 44303 13913
tri 44303 13905 44311 13913 sw
tri 44035 13897 44043 13905 ne
rect 44043 13897 44311 13905
tri 44311 13897 44319 13905 sw
tri 44043 13889 44051 13897 ne
rect 44051 13889 44319 13897
tri 44319 13889 44327 13897 sw
tri 44051 13881 44059 13889 ne
rect 44059 13881 44327 13889
tri 44327 13881 44335 13889 sw
tri 44059 13873 44067 13881 ne
rect 44067 13873 44335 13881
tri 44335 13873 44343 13881 sw
tri 44067 13865 44075 13873 ne
rect 44075 13865 44343 13873
tri 44343 13865 44351 13873 sw
tri 44075 13857 44083 13865 ne
rect 44083 13857 44351 13865
tri 44351 13857 44359 13865 sw
tri 44083 13849 44091 13857 ne
rect 44091 13849 44359 13857
tri 44359 13849 44367 13857 sw
tri 44091 13841 44099 13849 ne
rect 44099 13841 44367 13849
tri 44367 13841 44375 13849 sw
tri 44099 13833 44107 13841 ne
rect 44107 13833 44375 13841
tri 44375 13833 44383 13841 sw
tri 44107 13825 44115 13833 ne
rect 44115 13825 44383 13833
tri 44383 13825 44391 13833 sw
tri 44115 13817 44123 13825 ne
rect 44123 13817 44391 13825
tri 44391 13817 44399 13825 sw
tri 44123 13809 44131 13817 ne
rect 44131 13809 44399 13817
tri 44399 13809 44407 13817 sw
tri 44131 13801 44139 13809 ne
rect 44139 13801 44407 13809
tri 44407 13801 44415 13809 sw
tri 44139 13793 44147 13801 ne
rect 44147 13793 44415 13801
tri 44415 13793 44423 13801 sw
tri 44147 13785 44155 13793 ne
rect 44155 13785 44423 13793
tri 44423 13785 44431 13793 sw
tri 44155 13781 44159 13785 ne
rect 44159 13781 44431 13785
tri 44159 13773 44167 13781 ne
rect 44167 13777 44431 13781
tri 44431 13777 44439 13785 sw
rect 44167 13773 44439 13777
tri 44167 13765 44175 13773 ne
rect 44175 13769 44439 13773
tri 44439 13769 44447 13777 sw
rect 44175 13765 44447 13769
tri 44175 13757 44183 13765 ne
rect 44183 13761 44447 13765
tri 44447 13761 44455 13769 sw
rect 44183 13757 44455 13761
tri 44183 13749 44191 13757 ne
rect 44191 13753 44455 13757
tri 44455 13753 44463 13761 sw
rect 44191 13749 44463 13753
tri 44191 13741 44199 13749 ne
rect 44199 13745 44463 13749
tri 44463 13745 44471 13753 sw
rect 44199 13741 44471 13745
tri 44199 13733 44207 13741 ne
rect 44207 13737 44471 13741
tri 44471 13737 44479 13745 sw
rect 44207 13733 44479 13737
tri 44207 13725 44215 13733 ne
rect 44215 13729 44479 13733
tri 44479 13729 44487 13737 sw
rect 44215 13725 44487 13729
tri 44215 13717 44223 13725 ne
rect 44223 13721 44487 13725
tri 44487 13721 44495 13729 sw
rect 44223 13717 44495 13721
tri 44223 13709 44231 13717 ne
rect 44231 13713 44495 13717
tri 44495 13713 44503 13721 sw
rect 44231 13709 44503 13713
tri 44231 13701 44239 13709 ne
rect 44239 13705 44503 13709
tri 44503 13705 44511 13713 sw
rect 44239 13701 44511 13705
tri 44239 13693 44247 13701 ne
rect 44247 13697 44511 13701
tri 44511 13697 44519 13705 sw
rect 44247 13693 44519 13697
tri 44247 13685 44255 13693 ne
rect 44255 13689 44519 13693
tri 44519 13689 44527 13697 sw
rect 44255 13685 44527 13689
tri 44255 13677 44263 13685 ne
rect 44263 13681 44527 13685
tri 44527 13681 44535 13689 sw
rect 44263 13677 44535 13681
tri 44263 13669 44271 13677 ne
rect 44271 13673 44535 13677
tri 44535 13673 44543 13681 sw
rect 44271 13669 44543 13673
tri 44271 13661 44279 13669 ne
rect 44279 13665 44543 13669
tri 44543 13665 44551 13673 sw
rect 44279 13661 44551 13665
tri 44279 13653 44287 13661 ne
rect 44287 13657 44551 13661
tri 44551 13657 44559 13665 sw
rect 44287 13653 44559 13657
tri 44287 13649 44291 13653 ne
rect 44291 13649 44559 13653
tri 44559 13649 44567 13657 sw
tri 44291 13645 44295 13649 ne
rect 44295 13645 44567 13649
tri 44567 13645 44571 13649 sw
tri 44295 13637 44303 13645 ne
rect 44303 13637 44571 13645
tri 44571 13637 44579 13645 sw
tri 44303 13629 44311 13637 ne
rect 44311 13629 44579 13637
tri 44579 13629 44587 13637 sw
tri 44311 13621 44319 13629 ne
rect 44319 13621 44587 13629
tri 44587 13621 44595 13629 sw
tri 44319 13613 44327 13621 ne
rect 44327 13613 44595 13621
tri 44595 13613 44603 13621 sw
tri 44327 13605 44335 13613 ne
rect 44335 13605 44603 13613
tri 44603 13605 44611 13613 sw
tri 44335 13597 44343 13605 ne
rect 44343 13597 44611 13605
tri 44611 13597 44619 13605 sw
tri 44343 13589 44351 13597 ne
rect 44351 13589 44619 13597
tri 44619 13589 44627 13597 sw
tri 44351 13581 44359 13589 ne
rect 44359 13581 44627 13589
tri 44627 13581 44635 13589 sw
tri 44359 13573 44367 13581 ne
rect 44367 13573 44635 13581
tri 44635 13573 44643 13581 sw
tri 44367 13565 44375 13573 ne
rect 44375 13565 44643 13573
tri 44643 13565 44651 13573 sw
tri 44375 13557 44383 13565 ne
rect 44383 13557 44651 13565
tri 44651 13557 44659 13565 sw
tri 44383 13549 44391 13557 ne
rect 44391 13549 44659 13557
tri 44659 13549 44667 13557 sw
tri 44391 13541 44399 13549 ne
rect 44399 13541 44667 13549
tri 44667 13541 44675 13549 sw
tri 44399 13533 44407 13541 ne
rect 44407 13533 44675 13541
tri 44675 13533 44683 13541 sw
tri 44407 13525 44415 13533 ne
rect 44415 13525 44683 13533
tri 44683 13525 44691 13533 sw
tri 44415 13517 44423 13525 ne
rect 44423 13517 44691 13525
tri 44691 13517 44699 13525 sw
tri 44423 13509 44431 13517 ne
rect 44431 13509 44699 13517
tri 44699 13509 44707 13517 sw
tri 44431 13505 44435 13509 ne
rect 44435 13505 44707 13509
tri 44707 13505 44711 13509 sw
tri 44435 13497 44443 13505 ne
rect 44443 13497 44711 13505
tri 44711 13497 44719 13505 sw
tri 44443 13489 44451 13497 ne
rect 44451 13489 44719 13497
tri 44719 13489 44727 13497 sw
tri 44451 13481 44459 13489 ne
rect 44459 13481 44727 13489
tri 44727 13481 44735 13489 sw
tri 44459 13473 44467 13481 ne
rect 44467 13473 44735 13481
tri 44735 13473 44743 13481 sw
tri 44467 13465 44475 13473 ne
rect 44475 13465 44743 13473
tri 44743 13465 44751 13473 sw
tri 44475 13457 44483 13465 ne
rect 44483 13457 44751 13465
tri 44751 13457 44759 13465 sw
tri 44483 13449 44491 13457 ne
rect 44491 13449 44759 13457
tri 44759 13449 44767 13457 sw
tri 44491 13441 44499 13449 ne
rect 44499 13441 44767 13449
tri 44767 13441 44775 13449 sw
tri 44499 13433 44507 13441 ne
rect 44507 13433 44775 13441
tri 44775 13433 44783 13441 sw
tri 44507 13425 44515 13433 ne
rect 44515 13425 44783 13433
tri 44783 13425 44791 13433 sw
tri 44515 13417 44523 13425 ne
rect 44523 13417 44791 13425
tri 44791 13417 44799 13425 sw
tri 44523 13409 44531 13417 ne
rect 44531 13409 44799 13417
tri 44799 13409 44807 13417 sw
tri 44531 13401 44539 13409 ne
rect 44539 13401 44807 13409
tri 44807 13401 44815 13409 sw
tri 44539 13393 44547 13401 ne
rect 44547 13393 44815 13401
tri 44815 13393 44823 13401 sw
tri 44547 13385 44555 13393 ne
rect 44555 13385 44823 13393
tri 44823 13385 44831 13393 sw
tri 44555 13377 44563 13385 ne
rect 44563 13377 44831 13385
tri 44831 13377 44839 13385 sw
tri 44563 13373 44567 13377 ne
rect 44567 13373 44839 13377
tri 44839 13373 44843 13377 sw
tri 44567 13369 44571 13373 ne
rect 44571 13369 44843 13373
tri 44843 13369 44847 13373 sw
tri 44571 13361 44579 13369 ne
rect 44579 13361 44847 13369
tri 44847 13361 44855 13369 sw
tri 44579 13353 44587 13361 ne
rect 44587 13353 44855 13361
tri 44855 13353 44863 13361 sw
tri 44587 13345 44595 13353 ne
rect 44595 13345 44863 13353
tri 44863 13345 44871 13353 sw
tri 44595 13337 44603 13345 ne
rect 44603 13337 44871 13345
tri 44871 13337 44879 13345 sw
tri 44603 13329 44611 13337 ne
rect 44611 13335 44879 13337
tri 44879 13335 44881 13337 sw
rect 44611 13329 44881 13335
tri 44611 13321 44619 13329 ne
rect 44619 13327 44881 13329
tri 44881 13327 44889 13335 sw
rect 44619 13321 44889 13327
tri 44619 13313 44627 13321 ne
rect 44627 13319 44889 13321
tri 44889 13319 44897 13327 sw
rect 44627 13313 44897 13319
tri 44627 13305 44635 13313 ne
rect 44635 13311 44897 13313
tri 44897 13311 44905 13319 sw
rect 44635 13305 44905 13311
tri 44635 13297 44643 13305 ne
rect 44643 13303 44905 13305
tri 44905 13303 44913 13311 sw
rect 44643 13297 44913 13303
tri 44643 13289 44651 13297 ne
rect 44651 13295 44913 13297
tri 44913 13295 44921 13303 sw
rect 44651 13291 44921 13295
tri 44921 13291 44925 13295 sw
rect 44651 13289 46172 13291
tri 44651 13281 44659 13289 ne
rect 44659 13281 46172 13289
tri 44659 13273 44667 13281 ne
rect 44667 13273 46172 13281
tri 44667 13265 44675 13273 ne
rect 44675 13265 46172 13273
tri 44675 13257 44683 13265 ne
rect 44683 13257 46172 13265
tri 44683 13249 44691 13257 ne
rect 44691 13249 46172 13257
tri 44691 13241 44699 13249 ne
rect 44699 13241 46172 13249
tri 44699 13233 44707 13241 ne
rect 44707 13233 46172 13241
tri 44707 13229 44711 13233 ne
rect 44711 13229 46172 13233
tri 44711 13221 44719 13229 ne
rect 44719 13221 46172 13229
tri 44719 13213 44727 13221 ne
rect 44727 13213 46172 13221
tri 44727 13205 44735 13213 ne
rect 44735 13205 46172 13213
tri 44735 13197 44743 13205 ne
rect 44743 13197 46172 13205
tri 44743 13189 44751 13197 ne
rect 44751 13189 46172 13197
tri 44751 13181 44759 13189 ne
rect 44759 13181 46172 13189
tri 44759 13173 44767 13181 ne
rect 44767 13173 46172 13181
tri 44767 13165 44775 13173 ne
rect 44775 13165 46172 13173
tri 44775 13157 44783 13165 ne
rect 44783 13157 46172 13165
tri 44783 13149 44791 13157 ne
rect 44791 13149 46172 13157
tri 44791 13141 44799 13149 ne
rect 44799 13141 46172 13149
tri 44799 13133 44807 13141 ne
rect 44807 13133 46172 13141
tri 44807 13125 44815 13133 ne
rect 44815 13125 46172 13133
tri 44815 13117 44823 13125 ne
rect 44823 13117 46172 13125
tri 44823 13109 44831 13117 ne
rect 44831 13109 46172 13117
tri 44831 13101 44839 13109 ne
rect 44839 13101 46172 13109
tri 44839 13097 44843 13101 ne
rect 44843 13097 46172 13101
rect 70802 13097 71000 13436
<< metal1 >>
rect 13108 70814 69957 71000
rect 69785 69930 69957 70814
rect 70656 69785 71000 69957
rect 13108 44848 13280 45051
tri 13108 44828 13128 44848 ne
rect 13128 44828 13280 44848
tri 13280 44828 13372 44920 sw
tri 13128 44584 13372 44828 ne
tri 13372 44584 13616 44828 sw
tri 13372 44340 13616 44584 ne
tri 13616 44340 13860 44584 sw
tri 13616 44096 13860 44340 ne
tri 13860 44096 14104 44340 sw
tri 13860 43852 14104 44096 ne
tri 14104 43852 14348 44096 sw
tri 14104 43608 14348 43852 ne
tri 14348 43608 14592 43852 sw
tri 14348 43364 14592 43608 ne
tri 14592 43364 14836 43608 sw
tri 14592 43120 14836 43364 ne
tri 14836 43120 15080 43364 sw
tri 14836 42876 15080 43120 ne
tri 15080 42876 15324 43120 sw
tri 15080 42632 15324 42876 ne
tri 15324 42632 15568 42876 sw
tri 15324 42388 15568 42632 ne
tri 15568 42388 15812 42632 sw
tri 15568 42144 15812 42388 ne
tri 15812 42144 16056 42388 sw
tri 15812 41900 16056 42144 ne
tri 16056 41900 16300 42144 sw
tri 16056 41656 16300 41900 ne
tri 16300 41656 16544 41900 sw
tri 16300 41412 16544 41656 ne
tri 16544 41412 16788 41656 sw
tri 16544 41168 16788 41412 ne
tri 16788 41168 17032 41412 sw
tri 16788 40924 17032 41168 ne
tri 17032 40924 17276 41168 sw
tri 17032 40680 17276 40924 ne
tri 17276 40680 17520 40924 sw
tri 17276 40436 17520 40680 ne
tri 17520 40436 17764 40680 sw
tri 17520 40192 17764 40436 ne
tri 17764 40192 18008 40436 sw
tri 17764 39948 18008 40192 ne
tri 18008 39948 18252 40192 sw
tri 18008 39704 18252 39948 ne
tri 18252 39704 18496 39948 sw
tri 18252 39460 18496 39704 ne
tri 18496 39460 18740 39704 sw
tri 18496 39216 18740 39460 ne
tri 18740 39216 18984 39460 sw
tri 18740 38972 18984 39216 ne
tri 18984 38972 19228 39216 sw
tri 18984 38728 19228 38972 ne
tri 19228 38728 19472 38972 sw
tri 19228 38484 19472 38728 ne
tri 19472 38484 19716 38728 sw
tri 19472 38240 19716 38484 ne
tri 19716 38240 19960 38484 sw
tri 19716 37996 19960 38240 ne
tri 19960 37996 20204 38240 sw
tri 19960 37752 20204 37996 ne
tri 20204 37752 20448 37996 sw
tri 20204 37508 20448 37752 ne
tri 20448 37508 20692 37752 sw
tri 20448 37264 20692 37508 ne
tri 20692 37264 20936 37508 sw
tri 20692 37020 20936 37264 ne
tri 20936 37020 21180 37264 sw
tri 20936 36776 21180 37020 ne
tri 21180 36776 21424 37020 sw
tri 21180 36532 21424 36776 ne
tri 21424 36532 21668 36776 sw
tri 21424 36288 21668 36532 ne
tri 21668 36288 21912 36532 sw
tri 21668 36044 21912 36288 ne
tri 21912 36044 22156 36288 sw
tri 21912 35800 22156 36044 ne
tri 22156 35800 22400 36044 sw
tri 22156 35556 22400 35800 ne
tri 22400 35556 22644 35800 sw
tri 22400 35312 22644 35556 ne
tri 22644 35312 22888 35556 sw
tri 22644 35068 22888 35312 ne
tri 22888 35068 23132 35312 sw
tri 22888 34824 23132 35068 ne
tri 23132 34824 23376 35068 sw
tri 23132 34580 23376 34824 ne
tri 23376 34580 23620 34824 sw
tri 23376 34336 23620 34580 ne
tri 23620 34336 23864 34580 sw
tri 23620 34092 23864 34336 ne
tri 23864 34092 24108 34336 sw
tri 23864 33848 24108 34092 ne
tri 24108 33848 24352 34092 sw
tri 24108 33604 24352 33848 ne
tri 24352 33604 24596 33848 sw
tri 24352 33360 24596 33604 ne
tri 24596 33360 24840 33604 sw
tri 24596 33116 24840 33360 ne
tri 24840 33116 25084 33360 sw
tri 24840 32872 25084 33116 ne
tri 25084 32872 25328 33116 sw
tri 25084 32628 25328 32872 ne
tri 25328 32628 25572 32872 sw
tri 25328 32384 25572 32628 ne
tri 25572 32384 25816 32628 sw
tri 25572 32140 25816 32384 ne
tri 25816 32140 26060 32384 sw
tri 25816 31896 26060 32140 ne
tri 26060 31896 26304 32140 sw
tri 26060 31652 26304 31896 ne
tri 26304 31652 26548 31896 sw
tri 26304 31408 26548 31652 ne
tri 26548 31408 26792 31652 sw
tri 26548 31164 26792 31408 ne
tri 26792 31164 27036 31408 sw
tri 26792 30920 27036 31164 ne
tri 27036 30920 27280 31164 sw
tri 27036 30676 27280 30920 ne
tri 27280 30676 27524 30920 sw
tri 27280 30432 27524 30676 ne
tri 27524 30432 27768 30676 sw
tri 27524 30188 27768 30432 ne
tri 27768 30188 28012 30432 sw
tri 27768 29944 28012 30188 ne
tri 28012 29944 28256 30188 sw
tri 28012 29700 28256 29944 ne
tri 28256 29700 28500 29944 sw
tri 28256 29456 28500 29700 ne
tri 28500 29456 28744 29700 sw
tri 28500 29212 28744 29456 ne
tri 28744 29212 28988 29456 sw
tri 28744 28968 28988 29212 ne
tri 28988 28968 29232 29212 sw
tri 28988 28724 29232 28968 ne
tri 29232 28724 29476 28968 sw
tri 29232 28480 29476 28724 ne
tri 29476 28480 29720 28724 sw
tri 29476 28236 29720 28480 ne
tri 29720 28236 29964 28480 sw
tri 29720 27992 29964 28236 ne
tri 29964 27992 30208 28236 sw
tri 29964 27748 30208 27992 ne
tri 30208 27748 30452 27992 sw
tri 30208 27504 30452 27748 ne
tri 30452 27504 30696 27748 sw
tri 30452 27260 30696 27504 ne
tri 30696 27260 30940 27504 sw
tri 30696 27016 30940 27260 ne
tri 30940 27016 31184 27260 sw
tri 30940 26772 31184 27016 ne
tri 31184 26772 31428 27016 sw
tri 31184 26528 31428 26772 ne
tri 31428 26528 31672 26772 sw
tri 31428 26284 31672 26528 ne
tri 31672 26284 31916 26528 sw
tri 31672 26040 31916 26284 ne
tri 31916 26040 32160 26284 sw
tri 31916 25796 32160 26040 ne
tri 32160 25796 32404 26040 sw
tri 32160 25552 32404 25796 ne
tri 32404 25552 32648 25796 sw
tri 32404 25308 32648 25552 ne
tri 32648 25308 32892 25552 sw
tri 32648 25064 32892 25308 ne
tri 32892 25064 33136 25308 sw
tri 32892 24820 33136 25064 ne
tri 33136 24820 33380 25064 sw
tri 33136 24576 33380 24820 ne
tri 33380 24576 33624 24820 sw
tri 33380 24332 33624 24576 ne
tri 33624 24332 33868 24576 sw
tri 33624 24088 33868 24332 ne
tri 33868 24088 34112 24332 sw
tri 33868 23844 34112 24088 ne
tri 34112 23844 34356 24088 sw
tri 34112 23600 34356 23844 ne
tri 34356 23600 34600 23844 sw
tri 34356 23356 34600 23600 ne
tri 34600 23356 34844 23600 sw
tri 34600 23112 34844 23356 ne
tri 34844 23112 35088 23356 sw
tri 34844 22868 35088 23112 ne
tri 35088 22868 35332 23112 sw
tri 35088 22624 35332 22868 ne
tri 35332 22624 35576 22868 sw
tri 35332 22380 35576 22624 ne
tri 35576 22380 35820 22624 sw
tri 35576 22136 35820 22380 ne
tri 35820 22136 36064 22380 sw
tri 35820 21892 36064 22136 ne
tri 36064 21892 36308 22136 sw
tri 36064 21648 36308 21892 ne
tri 36308 21648 36552 21892 sw
tri 36308 21404 36552 21648 ne
tri 36552 21404 36796 21648 sw
tri 36552 21160 36796 21404 ne
tri 36796 21160 37040 21404 sw
tri 36796 20916 37040 21160 ne
tri 37040 20916 37284 21160 sw
tri 37040 20672 37284 20916 ne
tri 37284 20672 37528 20916 sw
tri 37284 20428 37528 20672 ne
tri 37528 20428 37772 20672 sw
tri 37528 20184 37772 20428 ne
tri 37772 20184 38016 20428 sw
tri 37772 19940 38016 20184 ne
tri 38016 19940 38260 20184 sw
tri 38016 19696 38260 19940 ne
tri 38260 19696 38504 19940 sw
tri 38260 19452 38504 19696 ne
tri 38504 19452 38748 19696 sw
tri 38504 19208 38748 19452 ne
tri 38748 19208 38992 19452 sw
tri 38748 18964 38992 19208 ne
tri 38992 18964 39236 19208 sw
tri 38992 18720 39236 18964 ne
tri 39236 18720 39480 18964 sw
tri 39236 18476 39480 18720 ne
tri 39480 18476 39724 18720 sw
tri 39480 18232 39724 18476 ne
tri 39724 18232 39968 18476 sw
tri 39724 17988 39968 18232 ne
tri 39968 17988 40212 18232 sw
tri 39968 17744 40212 17988 ne
tri 40212 17744 40456 17988 sw
tri 40212 17500 40456 17744 ne
tri 40456 17500 40700 17744 sw
tri 40456 17256 40700 17500 ne
tri 40700 17256 40944 17500 sw
tri 40700 17012 40944 17256 ne
tri 40944 17012 41188 17256 sw
tri 40944 16768 41188 17012 ne
tri 41188 16768 41432 17012 sw
tri 41188 16524 41432 16768 ne
tri 41432 16524 41676 16768 sw
tri 41432 16280 41676 16524 ne
tri 41676 16280 41920 16524 sw
tri 41676 16036 41920 16280 ne
tri 41920 16036 42164 16280 sw
tri 41920 15792 42164 16036 ne
tri 42164 15792 42408 16036 sw
tri 42164 15548 42408 15792 ne
tri 42408 15548 42652 15792 sw
tri 42408 15304 42652 15548 ne
tri 42652 15304 42896 15548 sw
tri 42652 15060 42896 15304 ne
tri 42896 15060 43140 15304 sw
tri 42896 14816 43140 15060 ne
tri 43140 14816 43384 15060 sw
tri 43140 14572 43384 14816 ne
tri 43384 14572 43628 14816 sw
tri 43384 14328 43628 14572 ne
tri 43628 14328 43872 14572 sw
tri 43628 14084 43872 14328 ne
tri 43872 14084 44116 14328 sw
tri 43872 13840 44116 14084 ne
tri 44116 13840 44360 14084 sw
tri 44116 13596 44360 13840 ne
tri 44360 13596 44604 13840 sw
tri 44360 13352 44604 13596 ne
tri 44604 13352 44848 13596 sw
tri 44604 13108 44848 13352 ne
tri 44848 13280 44920 13352 sw
rect 44848 13108 46414 13280
rect 70813 13108 71000 69785
<< metal2 >>
rect 70584 23599 70702 68200
<< metal3 >>
rect 14000 47020 17000 71000
rect 17200 48366 20200 71000
rect 20400 49774 23400 71000
rect 23600 50362 25000 71000
rect 25200 51120 26600 71000
rect 26800 52360 29800 71000
rect 30000 53704 33000 71000
rect 33200 55027 36200 71000
rect 36400 56465 39400 71000
rect 39600 57132 41000 71000
rect 41200 57810 42600 71000
rect 42800 59044 45800 71000
rect 46000 60708 49000 71000
rect 49200 61091 50600 71000
rect 50800 61751 52200 71000
rect 52400 62421 53800 71000
rect 54000 63320 55400 71000
rect 55600 63753 57000 71000
rect 57200 64540 58600 71000
rect 58800 65081 60200 71000
rect 60400 65760 61800 71000
rect 62000 66402 63400 71000
rect 63600 67263 65000 71000
rect 65200 67745 66600 71000
rect 66800 68493 68200 71000
rect 68400 69678 69678 71000
rect 68400 68769 71000 69678
tri 68400 68693 68476 68769 ne
rect 68476 68693 71000 68769
tri 68200 68493 68400 68693 sw
tri 68476 68493 68676 68693 ne
rect 68676 68493 71000 68693
rect 66800 68400 68400 68493
tri 68400 68400 68493 68493 sw
tri 68676 68400 68769 68493 ne
rect 68769 68400 71000 68493
rect 66800 68200 68493 68400
tri 68493 68200 68693 68400 sw
rect 66800 68113 71000 68200
tri 66800 68029 66884 68113 ne
rect 66884 68029 71000 68113
tri 66600 67745 66884 68029 sw
tri 66884 67745 67168 68029 ne
rect 67168 67745 71000 68029
rect 65200 67461 66884 67745
tri 66884 67461 67168 67745 sw
tri 67168 67461 67452 67745 ne
rect 67452 67461 71000 67745
rect 65200 67452 67168 67461
tri 67168 67452 67177 67461 sw
tri 67452 67452 67461 67461 ne
rect 67461 67452 71000 67461
rect 65200 67449 67177 67452
tri 65200 67366 65283 67449 ne
rect 65283 67366 67177 67449
tri 65000 67263 65103 67366 sw
tri 65283 67263 65386 67366 ne
rect 65386 67263 67177 67366
rect 63600 66980 65103 67263
tri 65103 66980 65386 67263 sw
tri 65386 66980 65669 67263 ne
rect 65669 67168 67177 67263
tri 67177 67168 67461 67452 sw
tri 67461 67168 67745 67452 ne
rect 67745 67168 71000 67452
rect 65669 66980 67461 67168
rect 63600 66786 65386 66980
tri 63600 66694 63692 66786 ne
rect 63692 66697 65386 66786
tri 65386 66697 65669 66980 sw
tri 65669 66697 65952 66980 ne
rect 65952 66884 67461 66980
tri 67461 66884 67745 67168 sw
tri 67745 66884 68029 67168 ne
rect 68029 66884 71000 67168
rect 65952 66697 67745 66884
rect 63692 66694 65669 66697
tri 63400 66402 63692 66694 sw
tri 63692 66402 63984 66694 ne
rect 63984 66414 65669 66694
tri 65669 66414 65952 66697 sw
tri 65952 66414 66235 66697 ne
rect 66235 66600 67745 66697
tri 67745 66600 68029 66884 sw
tri 68029 66800 68113 66884 ne
rect 68113 66800 71000 66884
rect 66235 66414 71000 66600
rect 63984 66402 65952 66414
rect 62000 66114 63692 66402
tri 62000 66031 62083 66114 ne
rect 62083 66110 63692 66114
tri 63692 66110 63984 66402 sw
tri 63984 66110 64276 66402 ne
rect 64276 66332 65952 66402
tri 65952 66332 66034 66414 sw
tri 66235 66332 66317 66414 ne
rect 66317 66332 71000 66414
rect 64276 66110 66034 66332
rect 62083 66031 63984 66110
tri 61800 65760 62071 66031 sw
tri 62083 65760 62354 66031 ne
rect 62354 65964 63984 66031
tri 63984 65964 64130 66110 sw
tri 64276 65964 64422 66110 ne
rect 64422 66049 66034 66110
tri 66034 66049 66317 66332 sw
tri 66317 66049 66600 66332 ne
rect 66600 66049 71000 66332
rect 64422 65964 66317 66049
rect 62354 65760 64130 65964
rect 60400 65477 62071 65760
tri 62071 65477 62354 65760 sw
tri 62354 65477 62637 65760 ne
rect 62637 65672 64130 65760
tri 64130 65672 64422 65964 sw
tri 64422 65672 64714 65964 ne
rect 64714 65766 66317 65964
tri 66317 65766 66600 66049 sw
tri 66600 65766 66883 66049 ne
rect 66883 65766 71000 66049
rect 64714 65672 66600 65766
rect 62637 65477 64422 65672
rect 60400 65451 62354 65477
tri 60400 65366 60485 65451 ne
rect 60485 65366 62354 65451
tri 60200 65081 60485 65366 sw
tri 60485 65081 60770 65366 ne
rect 60770 65194 62354 65366
tri 62354 65194 62637 65477 sw
tri 62637 65194 62920 65477 ne
rect 62920 65380 64422 65477
tri 64422 65380 64714 65672 sw
tri 64714 65380 65006 65672 ne
rect 65006 65566 66600 65672
tri 66600 65566 66800 65766 sw
tri 66883 65566 67083 65766 ne
rect 67083 65566 71000 65766
rect 65006 65380 66800 65566
rect 62920 65194 64714 65380
rect 60770 65081 62637 65194
rect 58800 64796 60485 65081
tri 60485 64796 60770 65081 sw
tri 60770 64796 61055 65081 ne
rect 61055 64997 62637 65081
tri 62637 64997 62834 65194 sw
tri 62920 64997 63117 65194 ne
rect 63117 65088 64714 65194
tri 64714 65088 65006 65380 sw
tri 65006 65088 65298 65380 ne
rect 65298 65283 66800 65380
tri 66800 65283 67083 65566 sw
tri 67083 65283 67366 65566 ne
rect 67366 65283 71000 65566
rect 65298 65088 67083 65283
rect 63117 65000 65006 65088
tri 65006 65000 65094 65088 sw
tri 65298 65000 65386 65088 ne
rect 65386 65000 67083 65088
tri 67083 65000 67366 65283 sw
tri 67366 65200 67449 65283 ne
rect 67449 65200 71000 65283
rect 63117 64997 65094 65000
rect 61055 64796 62834 64997
rect 58800 64786 60770 64796
tri 58800 64699 58887 64786 ne
rect 58887 64730 60770 64786
tri 60770 64730 60836 64796 sw
tri 61055 64730 61121 64796 ne
rect 61121 64730 62834 64796
rect 58887 64699 60836 64730
tri 58600 64540 58759 64699 sw
tri 58887 64540 59046 64699 ne
rect 59046 64540 60836 64699
rect 57200 64253 58759 64540
tri 58759 64253 59046 64540 sw
tri 59046 64253 59333 64540 ne
rect 59333 64445 60836 64540
tri 60836 64445 61121 64730 sw
tri 61121 64445 61406 64730 ne
rect 61406 64714 62834 64730
tri 62834 64714 63117 64997 sw
tri 63117 64714 63400 64997 ne
rect 63400 64714 65094 64997
rect 61406 64445 63117 64714
rect 59333 64253 61121 64445
rect 57200 64119 59046 64253
tri 57200 64036 57283 64119 ne
rect 57283 64036 59046 64119
tri 57000 63753 57283 64036 sw
tri 57283 63753 57566 64036 ne
rect 57566 63966 59046 64036
tri 59046 63966 59333 64253 sw
tri 59333 63966 59620 64253 ne
rect 59620 64160 61121 64253
tri 61121 64160 61406 64445 sw
tri 61406 64160 61691 64445 ne
rect 61691 64431 63117 64445
tri 63117 64431 63400 64714 sw
tri 63400 64431 63683 64714 ne
rect 63683 64708 65094 64714
tri 65094 64708 65386 65000 sw
tri 65386 64708 65678 65000 ne
rect 65678 64708 71000 65000
rect 63683 64431 65386 64708
rect 61691 64346 63400 64431
tri 63400 64346 63485 64431 sw
tri 63683 64346 63768 64431 ne
rect 63768 64416 65386 64431
tri 65386 64416 65678 64708 sw
tri 65678 64416 65970 64708 ne
rect 65970 64416 71000 64708
rect 63768 64346 65678 64416
rect 61691 64160 63485 64346
rect 59620 63966 61406 64160
rect 57566 63960 59333 63966
tri 59333 63960 59339 63966 sw
tri 59620 63960 59626 63966 ne
rect 59626 63960 61406 63966
rect 57566 63753 59339 63960
rect 55600 63506 57283 63753
tri 57283 63506 57530 63753 sw
tri 57566 63506 57813 63753 ne
rect 57813 63673 59339 63753
tri 59339 63673 59626 63960 sw
tri 59626 63673 59913 63960 ne
rect 59913 63875 61406 63960
tri 61406 63875 61691 64160 sw
tri 61691 63875 61976 64160 ne
rect 61976 64063 63485 64160
tri 63485 64063 63768 64346 sw
tri 63768 64063 64051 64346 ne
rect 64051 64276 65678 64346
tri 65678 64276 65818 64416 sw
tri 65970 64276 66110 64416 ne
rect 66110 64276 71000 64416
rect 64051 64063 65818 64276
rect 61976 63875 63768 64063
rect 59913 63780 61691 63875
tri 61691 63780 61786 63875 sw
tri 61976 63780 62071 63875 ne
rect 62071 63780 63768 63875
tri 63768 63780 64051 64063 sw
tri 64051 63780 64334 64063 ne
rect 64334 63984 65818 64063
tri 65818 63984 66110 64276 sw
tri 66110 63984 66402 64276 ne
rect 66402 63984 71000 64276
rect 64334 63780 66110 63984
rect 59913 63673 61786 63780
rect 57813 63506 59626 63673
rect 55600 63456 57530 63506
tri 55600 63373 55683 63456 ne
rect 55683 63373 57530 63456
tri 55400 63320 55453 63373 sw
tri 55683 63320 55736 63373 ne
rect 55736 63320 57530 63373
rect 54000 63037 55453 63320
tri 55453 63037 55736 63320 sw
tri 55736 63037 56019 63320 ne
rect 56019 63223 57530 63320
tri 57530 63223 57813 63506 sw
tri 57813 63223 58096 63506 ne
rect 58096 63386 59626 63506
tri 59626 63386 59913 63673 sw
tri 59913 63386 60200 63673 ne
rect 60200 63495 61786 63673
tri 61786 63495 62071 63780 sw
tri 62071 63495 62356 63780 ne
rect 62356 63497 64051 63780
tri 64051 63497 64334 63780 sw
tri 64334 63497 64617 63780 ne
rect 64617 63692 66110 63780
tri 66110 63692 66402 63984 sw
tri 66402 63692 66694 63984 ne
rect 66694 63692 71000 63984
rect 64617 63497 66402 63692
rect 62356 63495 64334 63497
rect 60200 63386 62071 63495
rect 58096 63223 59913 63386
rect 56019 63037 57813 63223
rect 54000 62793 55736 63037
tri 54000 62707 54086 62793 ne
rect 54086 62754 55736 62793
tri 55736 62754 56019 63037 sw
tri 56019 62754 56302 63037 ne
rect 56302 62940 57813 63037
tri 57813 62940 58096 63223 sw
tri 58096 62940 58379 63223 ne
rect 58379 63099 59913 63223
tri 59913 63099 60200 63386 sw
tri 60200 63099 60487 63386 ne
rect 60487 63210 62071 63386
tri 62071 63210 62356 63495 sw
tri 62356 63210 62641 63495 ne
rect 62641 63400 64334 63495
tri 64334 63400 64431 63497 sw
tri 64617 63400 64714 63497 ne
rect 64714 63400 66402 63497
tri 66402 63400 66694 63692 sw
tri 66694 63600 66786 63692 ne
rect 66786 63600 71000 63692
rect 62641 63210 64431 63400
rect 60487 63099 62356 63210
rect 58379 62940 60200 63099
rect 56302 62754 58096 62940
rect 54086 62707 56019 62754
tri 53800 62421 54086 62707 sw
tri 54086 62421 54372 62707 ne
rect 54372 62622 56019 62707
tri 56019 62622 56151 62754 sw
tri 56302 62622 56434 62754 ne
rect 56434 62657 58096 62754
tri 58096 62657 58379 62940 sw
tri 58379 62657 58662 62940 ne
rect 58662 62847 60200 62940
tri 60200 62847 60452 63099 sw
tri 60487 62847 60739 63099 ne
rect 60739 63035 62356 63099
tri 62356 63035 62531 63210 sw
tri 62641 63035 62816 63210 ne
rect 62816 63117 64431 63210
tri 64431 63117 64714 63400 sw
tri 64714 63117 64997 63400 ne
rect 64997 63117 71000 63400
rect 62816 63035 64714 63117
rect 60739 62847 62531 63035
rect 58662 62657 60452 62847
rect 56434 62622 58379 62657
rect 54372 62421 56151 62622
rect 52400 62292 54086 62421
tri 54086 62292 54215 62421 sw
tri 54372 62292 54501 62421 ne
rect 54501 62339 56151 62421
tri 56151 62339 56434 62622 sw
tri 56434 62339 56717 62622 ne
rect 56717 62560 58379 62622
tri 58379 62560 58476 62657 sw
tri 58662 62560 58759 62657 ne
rect 58759 62560 60452 62657
tri 60452 62560 60739 62847 sw
tri 60739 62560 61026 62847 ne
rect 61026 62750 62531 62847
tri 62531 62750 62816 63035 sw
tri 62816 62750 63101 63035 ne
rect 63101 62834 64714 63035
tri 64714 62834 64997 63117 sw
tri 64997 62834 65280 63117 ne
rect 65280 62834 71000 63117
rect 63101 62750 64997 62834
rect 61026 62560 62816 62750
rect 56717 62339 58476 62560
rect 54501 62292 56434 62339
rect 52400 62127 54215 62292
tri 52400 62039 52488 62127 ne
rect 52488 62039 54215 62127
tri 52200 61751 52488 62039 sw
tri 52488 61751 52776 62039 ne
rect 52776 62006 54215 62039
tri 54215 62006 54501 62292 sw
tri 54501 62006 54787 62292 ne
rect 54787 62056 56434 62292
tri 56434 62056 56717 62339 sw
tri 56717 62056 57000 62339 ne
rect 57000 62277 58476 62339
tri 58476 62277 58759 62560 sw
tri 58759 62277 59042 62560 ne
rect 59042 62277 60739 62560
rect 57000 62056 58759 62277
rect 54787 62006 56717 62056
rect 52776 61751 54501 62006
rect 50800 61463 52488 61751
tri 52488 61463 52776 61751 sw
tri 52776 61463 53064 61751 ne
rect 53064 61720 54501 61751
tri 54501 61720 54787 62006 sw
tri 54787 61720 55073 62006 ne
rect 55073 61773 56717 62006
tri 56717 61773 57000 62056 sw
tri 57000 61773 57283 62056 ne
rect 57283 61994 58759 62056
tri 58759 61994 59042 62277 sw
tri 59042 61994 59325 62277 ne
rect 59325 62273 60739 62277
tri 60739 62273 61026 62560 sw
tri 61026 62273 61313 62560 ne
rect 61313 62465 62816 62560
tri 62816 62465 63101 62750 sw
tri 63101 62465 63386 62750 ne
rect 63386 62649 64997 62750
tri 64997 62649 65182 62834 sw
tri 65280 62649 65465 62834 ne
rect 65465 62649 71000 62834
rect 63386 62465 65182 62649
rect 61313 62273 63101 62465
rect 59325 62180 61026 62273
tri 61026 62180 61119 62273 sw
tri 61313 62180 61406 62273 ne
rect 61406 62180 63101 62273
tri 63101 62180 63386 62465 sw
tri 63386 62180 63671 62465 ne
rect 63671 62366 65182 62465
tri 65182 62366 65465 62649 sw
tri 65465 62366 65748 62649 ne
rect 65748 62366 71000 62649
rect 63671 62180 65465 62366
rect 59325 61994 61119 62180
rect 57283 61809 59042 61994
tri 59042 61809 59227 61994 sw
tri 59325 61809 59510 61994 ne
rect 59510 61893 61119 61994
tri 61119 61893 61406 62180 sw
tri 61406 61893 61693 62180 ne
rect 61693 61895 63386 62180
tri 63386 61895 63671 62180 sw
tri 63671 61895 63956 62180 ne
rect 63956 62083 65465 62180
tri 65465 62083 65748 62366 sw
tri 65748 62083 66031 62366 ne
rect 66031 62083 71000 62366
rect 63956 61895 65748 62083
rect 61693 61893 63671 61895
rect 59510 61809 61406 61893
rect 57283 61773 59227 61809
rect 55073 61720 57000 61773
rect 53064 61463 54787 61720
rect 50800 61459 52776 61463
tri 50800 61375 50884 61459 ne
rect 50884 61375 52776 61459
tri 50600 61091 50884 61375 sw
tri 50884 61091 51168 61375 ne
rect 51168 61303 52776 61375
tri 52776 61303 52936 61463 sw
tri 53064 61303 53224 61463 ne
rect 53224 61434 54787 61463
tri 54787 61434 55073 61720 sw
tri 55073 61434 55359 61720 ne
rect 55359 61623 57000 61720
tri 57000 61623 57150 61773 sw
tri 57283 61623 57433 61773 ne
rect 57433 61623 59227 61773
rect 55359 61434 57150 61623
rect 53224 61340 55073 61434
tri 55073 61340 55167 61434 sw
tri 55359 61340 55453 61434 ne
rect 55453 61340 57150 61434
tri 57150 61340 57433 61623 sw
tri 57433 61340 57716 61623 ne
rect 57716 61526 59227 61623
tri 59227 61526 59510 61809 sw
tri 59510 61526 59793 61809 ne
rect 59793 61606 61406 61809
tri 61406 61606 61693 61893 sw
tri 61693 61606 61980 61893 ne
rect 61980 61800 63671 61893
tri 63671 61800 63766 61895 sw
tri 63956 61800 64051 61895 ne
rect 64051 61800 65748 61895
tri 65748 61800 66031 62083 sw
tri 66031 62000 66114 62083 ne
rect 66114 62000 71000 62083
rect 61980 61606 63766 61800
rect 59793 61526 61693 61606
rect 57716 61340 59510 61526
rect 53224 61303 55167 61340
rect 51168 61091 52936 61303
rect 49200 61068 50884 61091
tri 50884 61068 50907 61091 sw
tri 51168 61068 51191 61091 ne
rect 51191 61068 52936 61091
rect 49200 60795 50907 61068
tri 49200 60710 49285 60795 ne
rect 49285 60784 50907 60795
tri 50907 60784 51191 61068 sw
tri 51191 60784 51475 61068 ne
rect 51475 61015 52936 61068
tri 52936 61015 53224 61303 sw
tri 53224 61015 53512 61303 ne
rect 53512 61054 55167 61303
tri 55167 61054 55453 61340 sw
tri 55453 61054 55739 61340 ne
rect 55739 61057 57433 61340
tri 57433 61057 57716 61340 sw
tri 57716 61057 57999 61340 ne
rect 57999 61243 59510 61340
tri 59510 61243 59793 61526 sw
tri 59793 61243 60076 61526 ne
rect 60076 61441 61693 61526
tri 61693 61441 61858 61606 sw
tri 61980 61441 62145 61606 ne
rect 62145 61515 63766 61606
tri 63766 61515 64051 61800 sw
tri 64051 61515 64336 61800 ne
rect 64336 61515 71000 61800
rect 62145 61441 64051 61515
rect 60076 61243 61858 61441
rect 57999 61057 59793 61243
rect 55739 61054 57716 61057
rect 53512 61015 55453 61054
rect 51475 60784 53224 61015
rect 49285 60710 51191 60784
tri 49000 60708 49002 60710 sw
tri 49285 60708 49287 60710 ne
rect 49287 60708 51191 60710
rect 46000 60423 49002 60708
tri 49002 60423 49287 60708 sw
tri 49287 60423 49572 60708 ne
rect 49572 60500 51191 60708
tri 51191 60500 51475 60784 sw
tri 51475 60500 51759 60784 ne
rect 51759 60727 53224 60784
tri 53224 60727 53512 61015 sw
tri 53512 60727 53800 61015 ne
rect 53800 60768 55453 61015
tri 55453 60768 55739 61054 sw
tri 55739 60768 56025 61054 ne
rect 56025 60960 57716 61054
tri 57716 60960 57813 61057 sw
tri 57999 60960 58096 61057 ne
rect 58096 60960 59793 61057
tri 59793 60960 60076 61243 sw
tri 60076 60960 60359 61243 ne
rect 60359 61154 61858 61243
tri 61858 61154 62145 61441 sw
tri 62145 61154 62432 61441 ne
rect 62432 61230 64051 61441
tri 64051 61230 64336 61515 sw
tri 64336 61230 64621 61515 ne
rect 64621 61230 71000 61515
rect 62432 61154 64336 61230
rect 60359 60960 62145 61154
rect 56025 60768 57813 60960
rect 53800 60727 55739 60768
rect 51759 60500 53512 60727
rect 49572 60423 51475 60500
rect 46000 60138 49287 60423
tri 49287 60138 49572 60423 sw
tri 49572 60138 49857 60423 ne
rect 49857 60216 51475 60423
tri 51475 60216 51759 60500 sw
tri 51759 60216 52043 60500 ne
rect 52043 60439 53512 60500
tri 53512 60439 53800 60727 sw
tri 53800 60439 54088 60727 ne
rect 54088 60598 55739 60727
tri 55739 60598 55909 60768 sw
tri 56025 60598 56195 60768 ne
rect 56195 60677 57813 60768
tri 57813 60677 58096 60960 sw
tri 58096 60677 58379 60960 ne
rect 58379 60677 60076 60960
tri 60076 60677 60359 60960 sw
tri 60359 60677 60642 60960 ne
rect 60642 60867 62145 60960
tri 62145 60867 62432 61154 sw
tri 62432 60867 62719 61154 ne
rect 62719 61055 64336 61154
tri 64336 61055 64511 61230 sw
tri 64621 61055 64796 61230 ne
rect 64796 61055 71000 61230
rect 62719 60867 64511 61055
rect 60642 60677 62432 60867
rect 56195 60598 58096 60677
rect 54088 60439 55909 60598
rect 52043 60408 53800 60439
tri 53800 60408 53831 60439 sw
tri 54088 60408 54119 60439 ne
rect 54119 60408 55909 60439
rect 52043 60216 53831 60408
rect 49857 60138 51759 60216
rect 46000 59853 49572 60138
tri 49572 59853 49857 60138 sw
tri 49857 59853 50142 60138 ne
rect 50142 60059 51759 60138
tri 51759 60059 51916 60216 sw
tri 52043 60059 52200 60216 ne
rect 52200 60120 53831 60216
tri 53831 60120 54119 60408 sw
tri 54119 60120 54407 60408 ne
rect 54407 60312 55909 60408
tri 55909 60312 56195 60598 sw
tri 56195 60312 56481 60598 ne
rect 56481 60394 58096 60598
tri 58096 60394 58379 60677 sw
tri 58379 60394 58662 60677 ne
rect 58662 60580 60359 60677
tri 60359 60580 60456 60677 sw
tri 60642 60580 60739 60677 ne
rect 60739 60580 62432 60677
tri 62432 60580 62719 60867 sw
tri 62719 60580 63006 60867 ne
rect 63006 60770 64511 60867
tri 64511 60770 64796 61055 sw
tri 64796 60770 65081 61055 ne
rect 65081 60770 71000 61055
rect 63006 60580 64796 60770
rect 58662 60394 60456 60580
rect 56481 60312 58379 60394
rect 54407 60120 56195 60312
rect 52200 60059 54119 60120
rect 50142 59853 51916 60059
rect 46000 59683 49857 59853
tri 49857 59683 50027 59853 sw
tri 50142 59683 50312 59853 ne
rect 50312 59775 51916 59853
tri 51916 59775 52200 60059 sw
tri 52200 59775 52484 60059 ne
rect 52484 59832 54119 60059
tri 54119 59832 54407 60120 sw
tri 54407 59832 54695 60120 ne
rect 54695 60026 56195 60120
tri 56195 60026 56481 60312 sw
tri 56481 60026 56767 60312 ne
rect 56767 60209 58379 60312
tri 58379 60209 58564 60394 sw
tri 58662 60209 58847 60394 ne
rect 58847 60297 60456 60394
tri 60456 60297 60739 60580 sw
tri 60739 60297 61022 60580 ne
rect 61022 60297 62719 60580
rect 58847 60209 60739 60297
rect 56767 60026 58564 60209
rect 54695 59832 56481 60026
rect 52484 59775 54407 59832
rect 50312 59683 52200 59775
rect 46000 59461 50027 59683
tri 46000 59350 46111 59461 ne
rect 46111 59398 50027 59461
tri 50027 59398 50312 59683 sw
tri 50312 59398 50597 59683 ne
rect 50597 59491 52200 59683
tri 52200 59491 52484 59775 sw
tri 52484 59491 52768 59775 ne
rect 52768 59740 54407 59775
tri 54407 59740 54499 59832 sw
tri 54695 59740 54787 59832 ne
rect 54787 59740 56481 59832
tri 56481 59740 56767 60026 sw
tri 56767 59740 57053 60026 ne
rect 57053 59926 58564 60026
tri 58564 59926 58847 60209 sw
tri 58847 59926 59130 60209 ne
rect 59130 60014 60739 60209
tri 60739 60014 61022 60297 sw
tri 61022 60014 61305 60297 ne
rect 61305 60293 62719 60297
tri 62719 60293 63006 60580 sw
tri 63006 60293 63293 60580 ne
rect 63293 60485 64796 60580
tri 64796 60485 65081 60770 sw
tri 65081 60485 65366 60770 ne
rect 65366 60485 71000 60770
rect 63293 60293 65081 60485
rect 61305 60200 63006 60293
tri 63006 60200 63099 60293 sw
tri 63293 60200 63386 60293 ne
rect 63386 60200 65081 60293
tri 65081 60200 65366 60485 sw
tri 65366 60400 65451 60485 ne
rect 65451 60400 71000 60485
rect 61305 60014 63099 60200
rect 59130 59926 61022 60014
rect 57053 59740 58847 59926
rect 52768 59491 54499 59740
rect 50597 59398 52484 59491
rect 46111 59397 50312 59398
tri 50312 59397 50313 59398 sw
tri 50597 59397 50598 59398 ne
rect 50598 59397 52484 59398
rect 46111 59350 50313 59397
tri 45800 59044 46106 59350 sw
tri 46111 59044 46417 59350 ne
rect 46417 59112 50313 59350
tri 50313 59112 50598 59397 sw
tri 50598 59112 50883 59397 ne
rect 50883 59372 52484 59397
tri 52484 59372 52603 59491 sw
tri 52768 59372 52887 59491 ne
rect 52887 59452 54499 59491
tri 54499 59452 54787 59740 sw
tri 54787 59452 55075 59740 ne
rect 55075 59454 56767 59740
tri 56767 59454 57053 59740 sw
tri 57053 59454 57339 59740 ne
rect 57339 59643 58847 59740
tri 58847 59643 59130 59926 sw
tri 59130 59643 59413 59926 ne
rect 59413 59829 61022 59926
tri 61022 59829 61207 60014 sw
tri 61305 59829 61490 60014 ne
rect 61490 59913 63099 60014
tri 63099 59913 63386 60200 sw
tri 63386 59913 63673 60200 ne
rect 63673 59913 71000 60200
rect 61490 59829 63386 59913
rect 59413 59643 61207 59829
rect 57339 59454 59130 59643
rect 55075 59452 57053 59454
rect 52887 59372 54787 59452
rect 50883 59112 52603 59372
rect 46417 59110 50598 59112
tri 50598 59110 50600 59112 sw
tri 50883 59110 50885 59112 ne
rect 50885 59110 52603 59112
rect 46417 59044 50600 59110
rect 42800 58834 46106 59044
tri 46106 58834 46316 59044 sw
tri 46417 58834 46627 59044 ne
rect 46627 58834 50600 59044
rect 42800 58551 46316 58834
tri 46316 58551 46599 58834 sw
tri 46627 58551 46910 58834 ne
rect 46910 58825 50600 58834
tri 50600 58825 50885 59110 sw
tri 50885 58825 51170 59110 ne
rect 51170 59088 52603 59110
tri 52603 59088 52887 59372 sw
tri 52887 59088 53171 59372 ne
rect 53171 59164 54787 59372
tri 54787 59164 55075 59452 sw
tri 55075 59164 55363 59452 ne
rect 55363 59360 57053 59452
tri 57053 59360 57147 59454 sw
tri 57339 59360 57433 59454 ne
rect 57433 59360 59130 59454
tri 59130 59360 59413 59643 sw
tri 59413 59360 59696 59643 ne
rect 59696 59546 61207 59643
tri 61207 59546 61490 59829 sw
tri 61490 59546 61773 59829 ne
rect 61773 59626 63386 59829
tri 63386 59626 63673 59913 sw
tri 63673 59626 63960 59913 ne
rect 63960 59626 71000 59913
rect 61773 59546 63673 59626
rect 59696 59360 61490 59546
rect 55363 59164 57147 59360
rect 53171 59088 55075 59164
rect 51170 58825 52887 59088
rect 46910 58551 50885 58825
rect 42800 58436 46599 58551
tri 46599 58436 46714 58551 sw
tri 46910 58436 47025 58551 ne
rect 47025 58541 50885 58551
tri 50885 58541 51169 58825 sw
tri 51170 58541 51454 58825 ne
rect 51454 58804 52887 58825
tri 52887 58804 53171 59088 sw
tri 53171 58804 53455 59088 ne
rect 53455 59004 55075 59088
tri 55075 59004 55235 59164 sw
tri 55363 59004 55523 59164 ne
rect 55523 59074 57147 59164
tri 57147 59074 57433 59360 sw
tri 57433 59074 57719 59360 ne
rect 57719 59077 59413 59360
tri 59413 59077 59696 59360 sw
tri 59696 59077 59979 59360 ne
rect 59979 59263 61490 59360
tri 61490 59263 61773 59546 sw
tri 61773 59263 62056 59546 ne
rect 62056 59461 63673 59546
tri 63673 59461 63838 59626 sw
tri 63960 59461 64125 59626 ne
rect 64125 59461 71000 59626
rect 62056 59263 63838 59461
rect 59979 59077 61773 59263
rect 57719 59074 59696 59077
rect 55523 59004 57433 59074
rect 53455 58804 55235 59004
rect 51454 58541 53171 58804
rect 47025 58520 51169 58541
tri 51169 58520 51190 58541 sw
tri 51454 58520 51475 58541 ne
rect 51475 58520 53171 58541
tri 53171 58520 53455 58804 sw
tri 53455 58520 53739 58804 ne
rect 53739 58716 55235 58804
tri 55235 58716 55523 59004 sw
tri 55523 58716 55811 59004 ne
rect 55811 58788 57433 59004
tri 57433 58788 57719 59074 sw
tri 57719 58788 58005 59074 ne
rect 58005 58980 59696 59074
tri 59696 58980 59793 59077 sw
tri 59979 58980 60076 59077 ne
rect 60076 58980 61773 59077
tri 61773 58980 62056 59263 sw
tri 62056 58980 62339 59263 ne
rect 62339 59174 63838 59263
tri 63838 59174 64125 59461 sw
tri 64125 59174 64412 59461 ne
rect 64412 59174 71000 59461
rect 62339 58980 64125 59174
rect 58005 58788 59793 58980
rect 55811 58716 57719 58788
rect 53739 58520 55523 58716
rect 47025 58436 51190 58520
rect 42800 58131 46714 58436
tri 46714 58131 47019 58436 sw
tri 47025 58131 47330 58436 ne
rect 47330 58235 51190 58436
tri 51190 58235 51475 58520 sw
tri 51475 58235 51760 58520 ne
rect 51760 58236 53455 58520
tri 53455 58236 53739 58520 sw
tri 53739 58236 54023 58520 ne
rect 54023 58428 55523 58520
tri 55523 58428 55811 58716 sw
tri 55811 58428 56099 58716 ne
rect 56099 58618 57719 58716
tri 57719 58618 57889 58788 sw
tri 58005 58618 58175 58788 ne
rect 58175 58697 59793 58788
tri 59793 58697 60076 58980 sw
tri 60076 58697 60359 58980 ne
rect 60359 58697 62056 58980
tri 62056 58697 62339 58980 sw
tri 62339 58697 62622 58980 ne
rect 62622 58887 64125 58980
tri 64125 58887 64412 59174 sw
tri 64412 58887 64699 59174 ne
rect 64699 58887 71000 59174
rect 62622 58697 64412 58887
rect 58175 58618 60076 58697
rect 56099 58428 57889 58618
rect 54023 58236 55811 58428
rect 51760 58235 53739 58236
rect 47330 58131 51475 58235
rect 42800 58097 47019 58131
tri 42800 58010 42887 58097 ne
rect 42887 58010 47019 58097
tri 42600 57810 42800 58010 sw
tri 42887 57810 43087 58010 ne
rect 43087 57888 47019 58010
tri 47019 57888 47262 58131 sw
tri 47330 57888 47573 58131 ne
rect 47573 57950 51475 58131
tri 51475 57950 51760 58235 sw
tri 51760 57950 52045 58235 ne
rect 52045 58140 53739 58235
tri 53739 58140 53835 58236 sw
tri 54023 58140 54119 58236 ne
rect 54119 58140 55811 58236
tri 55811 58140 56099 58428 sw
tri 56099 58140 56387 58428 ne
rect 56387 58332 57889 58428
tri 57889 58332 58175 58618 sw
tri 58175 58332 58461 58618 ne
rect 58461 58414 60076 58618
tri 60076 58414 60359 58697 sw
tri 60359 58414 60642 58697 ne
rect 60642 58600 62339 58697
tri 62339 58600 62436 58697 sw
tri 62622 58600 62719 58697 ne
rect 62719 58600 64412 58697
tri 64412 58600 64699 58887 sw
tri 64699 58800 64786 58887 ne
rect 64786 58800 71000 58887
rect 60642 58414 62436 58600
rect 58461 58332 60359 58414
rect 56387 58140 58175 58332
rect 52045 57950 53835 58140
rect 47573 57888 51760 57950
rect 43087 57810 47262 57888
rect 41200 57722 42800 57810
tri 42800 57722 42888 57810 sw
tri 43087 57722 43175 57810 ne
rect 43175 57722 47262 57810
rect 41200 57435 42888 57722
tri 42888 57435 43175 57722 sw
tri 43175 57435 43462 57722 ne
rect 43462 57582 47262 57722
tri 47262 57582 47568 57888 sw
tri 47573 57582 47879 57888 ne
rect 47879 57774 51760 57888
tri 51760 57774 51936 57950 sw
tri 52045 57774 52221 57950 ne
rect 52221 57856 53835 57950
tri 53835 57856 54119 58140 sw
tri 54119 57856 54403 58140 ne
rect 54403 57856 56099 58140
rect 52221 57774 54119 57856
rect 47879 57582 51936 57774
rect 43462 57562 47568 57582
tri 47568 57562 47588 57582 sw
tri 47879 57562 47899 57582 ne
rect 47899 57562 51936 57582
rect 43462 57435 47588 57562
rect 41200 57430 43175 57435
tri 41200 57338 41292 57430 ne
rect 41292 57338 43175 57430
tri 41000 57132 41206 57338 sw
tri 41292 57132 41498 57338 ne
rect 41498 57322 43175 57338
tri 43175 57322 43288 57435 sw
tri 43462 57322 43575 57435 ne
rect 43575 57322 47588 57435
rect 41498 57132 43288 57322
rect 39600 56840 41206 57132
tri 41206 56840 41498 57132 sw
tri 41498 56840 41790 57132 ne
rect 41790 57035 43288 57132
tri 43288 57035 43575 57322 sw
tri 43575 57035 43862 57322 ne
rect 43862 57260 47588 57322
tri 47588 57260 47890 57562 sw
tri 47899 57260 48201 57562 ne
rect 48201 57489 51936 57562
tri 51936 57489 52221 57774 sw
tri 52221 57489 52506 57774 ne
rect 52506 57572 54119 57774
tri 54119 57572 54403 57856 sw
tri 54403 57572 54687 57856 ne
rect 54687 57852 56099 57856
tri 56099 57852 56387 58140 sw
tri 56387 57852 56675 58140 ne
rect 56675 58046 58175 58140
tri 58175 58046 58461 58332 sw
tri 58461 58046 58747 58332 ne
rect 58747 58229 60359 58332
tri 60359 58229 60544 58414 sw
tri 60642 58229 60827 58414 ne
rect 60827 58317 62436 58414
tri 62436 58317 62719 58600 sw
tri 62719 58317 63002 58600 ne
rect 63002 58317 71000 58600
rect 60827 58229 62719 58317
rect 58747 58046 60544 58229
rect 56675 57852 58461 58046
rect 54687 57760 56387 57852
tri 56387 57760 56479 57852 sw
tri 56675 57760 56767 57852 ne
rect 56767 57760 58461 57852
tri 58461 57760 58747 58046 sw
tri 58747 57760 59033 58046 ne
rect 59033 57946 60544 58046
tri 60544 57946 60827 58229 sw
tri 60827 57946 61110 58229 ne
rect 61110 58034 62719 58229
tri 62719 58034 63002 58317 sw
tri 63002 58034 63285 58317 ne
rect 63285 58034 71000 58317
rect 61110 57946 63002 58034
rect 59033 57760 60827 57946
rect 54687 57572 56479 57760
rect 52506 57489 54403 57572
rect 48201 57487 52221 57489
tri 52221 57487 52223 57489 sw
tri 52506 57487 52508 57489 ne
rect 52508 57487 54403 57489
rect 48201 57260 52223 57487
rect 43862 57126 47890 57260
tri 47890 57126 48024 57260 sw
tri 48201 57126 48335 57260 ne
rect 48335 57202 52223 57260
tri 52223 57202 52508 57487 sw
tri 52508 57202 52793 57487 ne
rect 52793 57392 54403 57487
tri 54403 57392 54583 57572 sw
tri 54687 57392 54867 57572 ne
rect 54867 57472 56479 57572
tri 56479 57472 56767 57760 sw
tri 56767 57472 57055 57760 ne
rect 57055 57474 58747 57760
tri 58747 57474 59033 57760 sw
tri 59033 57474 59319 57760 ne
rect 59319 57663 60827 57760
tri 60827 57663 61110 57946 sw
tri 61110 57663 61393 57946 ne
rect 61393 57849 63002 57946
tri 63002 57849 63187 58034 sw
tri 63285 57849 63470 58034 ne
rect 63470 57849 71000 58034
rect 61393 57663 63187 57849
rect 59319 57474 61110 57663
rect 57055 57472 59033 57474
rect 54867 57392 56767 57472
rect 52793 57202 54583 57392
rect 48335 57201 52508 57202
tri 52508 57201 52509 57202 sw
tri 52793 57201 52794 57202 ne
rect 52794 57201 54583 57202
rect 48335 57126 52509 57201
rect 43862 57035 48024 57126
rect 41790 56840 43575 57035
rect 39600 56758 41498 56840
tri 39600 56665 39693 56758 ne
rect 39693 56665 41498 56758
tri 39400 56465 39600 56665 sw
tri 39693 56465 39893 56665 ne
rect 39893 56548 41498 56665
tri 41498 56548 41790 56840 sw
tri 41790 56548 42082 56840 ne
rect 42082 56748 43575 56840
tri 43575 56748 43862 57035 sw
tri 43862 56748 44149 57035 ne
rect 44149 56820 48024 57035
tri 48024 56820 48330 57126 sw
tri 48335 56820 48641 57126 ne
rect 48641 56916 52509 57126
tri 52509 56916 52794 57201 sw
tri 52794 56916 53079 57201 ne
rect 53079 57108 54583 57201
tri 54583 57108 54867 57392 sw
tri 54867 57108 55151 57392 ne
rect 55151 57184 56767 57392
tri 56767 57184 57055 57472 sw
tri 57055 57184 57343 57472 ne
rect 57343 57380 59033 57472
tri 59033 57380 59127 57474 sw
tri 59319 57380 59413 57474 ne
rect 59413 57380 61110 57474
tri 61110 57380 61393 57663 sw
tri 61393 57380 61676 57663 ne
rect 61676 57566 63187 57663
tri 63187 57566 63470 57849 sw
tri 63470 57566 63753 57849 ne
rect 63753 57566 71000 57849
rect 61676 57380 63470 57566
rect 57343 57184 59127 57380
rect 55151 57108 57055 57184
rect 53079 56916 54867 57108
rect 48641 56914 52794 56916
tri 52794 56914 52796 56916 sw
tri 53079 56914 53081 56916 ne
rect 53081 56914 54867 56916
rect 48641 56820 52796 56914
rect 44149 56800 48330 56820
tri 48330 56800 48350 56820 sw
tri 48641 56800 48661 56820 ne
rect 48661 56800 52796 56820
rect 44149 56748 48350 56800
rect 42082 56747 43862 56748
tri 43862 56747 43863 56748 sw
tri 44149 56747 44150 56748 ne
rect 44150 56747 48350 56748
rect 42082 56548 43863 56747
rect 39893 56465 41790 56548
rect 36400 56371 39600 56465
tri 39600 56371 39694 56465 sw
tri 39893 56371 39987 56465 ne
rect 39987 56371 41790 56465
rect 36400 56078 39694 56371
tri 39694 56078 39987 56371 sw
tri 39987 56078 40280 56371 ne
rect 40280 56322 41790 56371
tri 41790 56322 42016 56548 sw
tri 42082 56322 42308 56548 ne
rect 42308 56460 43863 56548
tri 43863 56460 44150 56747 sw
tri 44150 56460 44437 56747 ne
rect 44437 56494 48350 56747
tri 48350 56494 48656 56800 sw
tri 48661 56494 48967 56800 ne
rect 48967 56630 52796 56800
tri 52796 56630 53080 56914 sw
tri 53081 56630 53365 56914 ne
rect 53365 56824 54867 56914
tri 54867 56824 55151 57108 sw
tri 55151 56824 55435 57108 ne
rect 55435 57024 57055 57108
tri 57055 57024 57215 57184 sw
tri 57343 57024 57503 57184 ne
rect 57503 57094 59127 57184
tri 59127 57094 59413 57380 sw
tri 59413 57094 59699 57380 ne
rect 59699 57097 61393 57380
tri 61393 57097 61676 57380 sw
tri 61676 57097 61959 57380 ne
rect 61959 57283 63470 57380
tri 63470 57283 63753 57566 sw
tri 63753 57283 64036 57566 ne
rect 64036 57283 71000 57566
rect 61959 57097 63753 57283
rect 59699 57094 61676 57097
rect 57503 57024 59413 57094
rect 55435 56824 57215 57024
rect 53365 56630 55151 56824
rect 48967 56540 53080 56630
tri 53080 56540 53170 56630 sw
tri 53365 56540 53455 56630 ne
rect 53455 56540 55151 56630
tri 55151 56540 55435 56824 sw
tri 55435 56540 55719 56824 ne
rect 55719 56736 57215 56824
tri 57215 56736 57503 57024 sw
tri 57503 56736 57791 57024 ne
rect 57791 56808 59413 57024
tri 59413 56808 59699 57094 sw
tri 59699 56808 59985 57094 ne
rect 59985 57000 61676 57094
tri 61676 57000 61773 57097 sw
tri 61959 57000 62056 57097 ne
rect 62056 57000 63753 57097
tri 63753 57000 64036 57283 sw
tri 64036 57200 64119 57283 ne
rect 64119 57200 71000 57283
rect 59985 56808 61773 57000
rect 57791 56736 59699 56808
rect 55719 56540 57503 56736
rect 48967 56494 53170 56540
rect 44437 56475 48656 56494
tri 48656 56475 48675 56494 sw
tri 48967 56475 48986 56494 ne
rect 48986 56475 53170 56494
rect 44437 56460 48675 56475
rect 42308 56459 44150 56460
tri 44150 56459 44151 56460 sw
tri 44437 56459 44438 56460 ne
rect 44438 56459 48675 56460
rect 42308 56322 44151 56459
rect 40280 56078 42016 56322
rect 36400 55785 39987 56078
tri 39987 55785 40280 56078 sw
tri 40280 55785 40573 56078 ne
rect 40573 56030 42016 56078
tri 42016 56030 42308 56322 sw
tri 42308 56030 42600 56322 ne
rect 42600 56172 44151 56322
tri 44151 56172 44438 56459 sw
tri 44438 56172 44725 56459 ne
rect 44725 56172 48675 56459
rect 42600 56030 44438 56172
rect 40573 55785 42308 56030
rect 36400 55492 40280 55785
tri 40280 55492 40573 55785 sw
tri 40573 55492 40866 55785 ne
rect 40866 55738 42308 55785
tri 42308 55738 42600 56030 sw
tri 42600 55738 42892 56030 ne
rect 42892 55885 44438 56030
tri 44438 55885 44725 56172 sw
tri 44725 55885 45012 56172 ne
rect 45012 56169 48675 56172
tri 48675 56169 48981 56475 sw
tri 48986 56169 49292 56475 ne
rect 49292 56255 53170 56475
tri 53170 56255 53455 56540 sw
tri 53455 56255 53740 56540 ne
rect 53740 56256 55435 56540
tri 55435 56256 55719 56540 sw
tri 55719 56256 56003 56540 ne
rect 56003 56448 57503 56540
tri 57503 56448 57791 56736 sw
tri 57791 56448 58079 56736 ne
rect 58079 56638 59699 56736
tri 59699 56638 59869 56808 sw
tri 59985 56638 60155 56808 ne
rect 60155 56717 61773 56808
tri 61773 56717 62056 57000 sw
tri 62056 56717 62339 57000 ne
rect 62339 56717 71000 57000
rect 60155 56638 62056 56717
rect 58079 56448 59869 56638
rect 56003 56256 57791 56448
rect 53740 56255 55719 56256
rect 49292 56169 53455 56255
rect 45012 56150 48981 56169
tri 48981 56150 49000 56169 sw
tri 49292 56150 49311 56169 ne
rect 49311 56150 53455 56169
rect 45012 55885 49000 56150
rect 42892 55884 44725 55885
tri 44725 55884 44726 55885 sw
tri 45012 55884 45013 55885 ne
rect 45013 55884 49000 55885
rect 42892 55738 44726 55884
rect 40866 55492 42600 55738
rect 36400 55421 40573 55492
tri 36400 55324 36497 55421 ne
rect 36497 55324 40573 55421
tri 36200 55027 36497 55324 sw
tri 36497 55027 36794 55324 ne
rect 36794 55199 40573 55324
tri 40573 55199 40866 55492 sw
tri 40866 55199 41159 55492 ne
rect 41159 55446 42600 55492
tri 42600 55446 42892 55738 sw
tri 42892 55446 43184 55738 ne
rect 43184 55597 44726 55738
tri 44726 55597 45013 55884 sw
tri 45013 55597 45300 55884 ne
rect 45300 55844 49000 55884
tri 49000 55844 49306 56150 sw
tri 49311 55844 49617 56150 ne
rect 49617 55970 53455 56150
tri 53455 55970 53740 56255 sw
tri 53740 55970 54025 56255 ne
rect 54025 56160 55719 56255
tri 55719 56160 55815 56256 sw
tri 56003 56160 56099 56256 ne
rect 56099 56160 57791 56256
tri 57791 56160 58079 56448 sw
tri 58079 56160 58367 56448 ne
rect 58367 56352 59869 56448
tri 59869 56352 60155 56638 sw
tri 60155 56352 60441 56638 ne
rect 60441 56434 62056 56638
tri 62056 56434 62339 56717 sw
tri 62339 56434 62622 56717 ne
rect 62622 56434 71000 56717
rect 60441 56352 62339 56434
rect 58367 56160 60155 56352
rect 54025 55970 55815 56160
rect 49617 55968 53740 55970
tri 53740 55968 53742 55970 sw
tri 54025 55968 54027 55970 ne
rect 54027 55968 55815 55970
rect 49617 55844 53742 55968
rect 45300 55597 49306 55844
rect 43184 55446 45013 55597
rect 41159 55444 42892 55446
tri 42892 55444 42894 55446 sw
tri 43184 55444 43186 55446 ne
rect 43186 55444 45013 55446
rect 41159 55199 42894 55444
rect 36794 55154 40866 55199
tri 40866 55154 40911 55199 sw
tri 41159 55154 41204 55199 ne
rect 41204 55154 42894 55199
rect 36794 55027 40911 55154
rect 33200 54827 36497 55027
tri 36497 54827 36697 55027 sw
tri 36794 54827 36994 55027 ne
rect 36994 54861 40911 55027
tri 40911 54861 41204 55154 sw
tri 41204 54861 41497 55154 ne
rect 41497 55152 42894 55154
tri 42894 55152 43186 55444 sw
tri 43186 55152 43478 55444 ne
rect 43478 55343 45013 55444
tri 45013 55343 45267 55597 sw
tri 45300 55343 45554 55597 ne
rect 45554 55559 49306 55597
tri 49306 55559 49591 55844 sw
tri 49617 55559 49902 55844 ne
rect 49902 55683 53742 55844
tri 53742 55683 54027 55968 sw
tri 54027 55683 54312 55968 ne
rect 54312 55876 55815 55968
tri 55815 55876 56099 56160 sw
tri 56099 55876 56383 56160 ne
rect 56383 55876 58079 56160
rect 54312 55683 56099 55876
rect 49902 55682 54027 55683
tri 54027 55682 54028 55683 sw
tri 54312 55682 54313 55683 ne
rect 54313 55682 56099 55683
rect 49902 55559 54028 55682
rect 45554 55343 49591 55559
rect 43478 55272 45267 55343
tri 45267 55272 45338 55343 sw
tri 45554 55272 45625 55343 ne
rect 45625 55272 49591 55343
rect 43478 55152 45338 55272
rect 41497 54861 43186 55152
rect 36994 54827 41204 54861
rect 33200 54728 36697 54827
tri 36697 54728 36796 54827 sw
tri 36994 54728 37093 54827 ne
rect 37093 54728 41204 54827
rect 33200 54431 36796 54728
tri 36796 54431 37093 54728 sw
tri 37093 54431 37390 54728 ne
rect 37390 54568 41204 54728
tri 41204 54568 41497 54861 sw
tri 41497 54568 41790 54861 ne
rect 41790 54860 43186 54861
tri 43186 54860 43478 55152 sw
tri 43478 54860 43770 55152 ne
rect 43770 55055 45338 55152
tri 45338 55055 45555 55272 sw
tri 45625 55055 45842 55272 ne
rect 45842 55257 49591 55272
tri 49591 55257 49893 55559 sw
tri 49902 55257 50204 55559 ne
rect 50204 55397 54028 55559
tri 54028 55397 54313 55682 sw
tri 54313 55397 54598 55682 ne
rect 54598 55592 56099 55682
tri 56099 55592 56383 55876 sw
tri 56383 55592 56667 55876 ne
rect 56667 55872 58079 55876
tri 58079 55872 58367 56160 sw
tri 58367 55872 58655 56160 ne
rect 58655 56066 60155 56160
tri 60155 56066 60441 56352 sw
tri 60441 56066 60727 56352 ne
rect 60727 56249 62339 56352
tri 62339 56249 62524 56434 sw
tri 62622 56249 62807 56434 ne
rect 62807 56249 71000 56434
rect 60727 56066 62524 56249
rect 58655 55872 60441 56066
rect 56667 55780 58367 55872
tri 58367 55780 58459 55872 sw
tri 58655 55780 58747 55872 ne
rect 58747 55780 60441 55872
tri 60441 55780 60727 56066 sw
tri 60727 55780 61013 56066 ne
rect 61013 55966 62524 56066
tri 62524 55966 62807 56249 sw
tri 62807 55966 63090 56249 ne
rect 63090 55966 71000 56249
rect 61013 55780 62807 55966
rect 56667 55592 58459 55780
rect 54598 55412 56383 55592
tri 56383 55412 56563 55592 sw
tri 56667 55412 56847 55592 ne
rect 56847 55492 58459 55592
tri 58459 55492 58747 55780 sw
tri 58747 55492 59035 55780 ne
rect 59035 55494 60727 55780
tri 60727 55494 61013 55780 sw
tri 61013 55494 61299 55780 ne
rect 61299 55683 62807 55780
tri 62807 55683 63090 55966 sw
tri 63090 55683 63373 55966 ne
rect 63373 55683 71000 55966
rect 61299 55494 63090 55683
rect 59035 55492 61013 55494
rect 56847 55412 58747 55492
rect 54598 55397 56563 55412
rect 50204 55257 54313 55397
rect 45842 55055 49893 55257
rect 43770 54860 45555 55055
rect 41790 54568 43478 54860
tri 43478 54568 43770 54860 sw
tri 43770 54568 44062 54860 ne
rect 44062 54768 45555 54860
tri 45555 54768 45842 55055 sw
tri 45842 54768 46129 55055 ne
rect 46129 54946 49893 55055
tri 49893 54946 50204 55257 sw
tri 50204 54946 50515 55257 ne
rect 50515 55135 54313 55257
tri 54313 55135 54575 55397 sw
tri 54598 55135 54860 55397 ne
rect 54860 55135 56563 55397
rect 50515 54946 54575 55135
rect 46129 54768 50204 54946
rect 44062 54767 45842 54768
tri 45842 54767 45843 54768 sw
tri 46129 54767 46130 54768 ne
rect 46130 54767 50204 54768
rect 44062 54568 45843 54767
rect 37390 54567 41497 54568
tri 41497 54567 41498 54568 sw
tri 41790 54567 41791 54568 ne
rect 41791 54567 43770 54568
rect 37390 54431 41498 54567
rect 33200 54429 37093 54431
tri 37093 54429 37095 54431 sw
tri 37390 54429 37392 54431 ne
rect 37392 54429 41498 54431
rect 33200 54133 37095 54429
tri 37095 54133 37391 54429 sw
tri 37392 54133 37688 54429 ne
rect 37688 54274 41498 54429
tri 41498 54274 41791 54567 sw
tri 41791 54274 42084 54567 ne
rect 42084 54402 43770 54567
tri 43770 54402 43936 54568 sw
tri 44062 54402 44228 54568 ne
rect 44228 54480 45843 54568
tri 45843 54480 46130 54767 sw
tri 46130 54480 46417 54767 ne
rect 46417 54640 50204 54767
tri 50204 54640 50510 54946 sw
tri 50515 54640 50821 54946 ne
rect 50821 54850 54575 54946
tri 54575 54850 54860 55135 sw
tri 54860 54850 55145 55135 ne
rect 55145 55128 56563 55135
tri 56563 55128 56847 55412 sw
tri 56847 55128 57131 55412 ne
rect 57131 55204 58747 55412
tri 58747 55204 59035 55492 sw
tri 59035 55204 59323 55492 ne
rect 59323 55400 61013 55492
tri 61013 55400 61107 55494 sw
tri 61299 55400 61393 55494 ne
rect 61393 55400 63090 55494
tri 63090 55400 63373 55683 sw
tri 63373 55600 63456 55683 ne
rect 63456 55600 71000 55683
rect 59323 55204 61107 55400
rect 57131 55128 59035 55204
rect 55145 54850 56847 55128
rect 50821 54848 54860 54850
tri 54860 54848 54862 54850 sw
tri 55145 54848 55147 54850 ne
rect 55147 54848 56847 54850
rect 50821 54640 54862 54848
rect 46417 54620 50510 54640
tri 50510 54620 50530 54640 sw
tri 50821 54620 50841 54640 ne
rect 50841 54620 54862 54640
rect 46417 54480 50530 54620
rect 44228 54402 46130 54480
rect 42084 54274 43936 54402
rect 37688 54273 41791 54274
tri 41791 54273 41792 54274 sw
tri 42084 54273 42085 54274 ne
rect 42085 54273 43936 54274
rect 37688 54133 41792 54273
rect 33200 54080 37391 54133
tri 37391 54080 37444 54133 sw
tri 37688 54080 37741 54133 ne
rect 37741 54080 41792 54133
tri 33200 53992 33288 54080 ne
rect 33288 53992 37444 54080
tri 33000 53704 33288 53992 sw
tri 33288 53704 33576 53992 ne
rect 33576 53783 37444 53992
tri 37444 53783 37741 54080 sw
tri 37741 53783 38038 54080 ne
rect 38038 53980 41792 54080
tri 41792 53980 42085 54273 sw
tri 42085 53980 42378 54273 ne
rect 42378 54188 43936 54273
tri 43936 54188 44150 54402 sw
tri 44228 54188 44442 54402 ne
rect 44442 54285 46130 54402
tri 46130 54285 46325 54480 sw
tri 46417 54285 46612 54480 ne
rect 46612 54312 50530 54480
tri 50530 54312 50838 54620 sw
tri 50841 54312 51149 54620 ne
rect 51149 54563 54862 54620
tri 54862 54563 55147 54848 sw
tri 55147 54563 55432 54848 ne
rect 55432 54844 56847 54848
tri 56847 54844 57131 55128 sw
tri 57131 54844 57415 55128 ne
rect 57415 55044 59035 55128
tri 59035 55044 59195 55204 sw
tri 59323 55044 59483 55204 ne
rect 59483 55114 61107 55204
tri 61107 55114 61393 55400 sw
tri 61393 55114 61679 55400 ne
rect 61679 55114 71000 55400
rect 59483 55044 61393 55114
rect 57415 54844 59195 55044
rect 55432 54563 57131 54844
rect 51149 54312 55147 54563
rect 46612 54285 50838 54312
rect 44442 54188 46325 54285
rect 42378 53980 44150 54188
rect 38038 53783 42085 53980
rect 33576 53768 37741 53783
tri 37741 53768 37756 53783 sw
tri 38038 53768 38053 53783 ne
rect 38053 53768 42085 53783
rect 33576 53704 37756 53768
rect 30000 53504 33288 53704
tri 33288 53504 33488 53704 sw
tri 33576 53504 33776 53704 ne
rect 33776 53504 37756 53704
rect 30000 53414 33488 53504
tri 33488 53414 33578 53504 sw
tri 33776 53414 33866 53504 ne
rect 33866 53471 37756 53504
tri 37756 53471 38053 53768 sw
tri 38053 53471 38350 53768 ne
rect 38350 53687 42085 53768
tri 42085 53687 42378 53980 sw
tri 42378 53687 42671 53980 ne
rect 42671 53896 44150 53980
tri 44150 53896 44442 54188 sw
tri 44442 53896 44734 54188 ne
rect 44734 53998 46325 54188
tri 46325 53998 46612 54285 sw
tri 46612 53998 46899 54285 ne
rect 46899 54187 50838 54285
tri 50838 54187 50963 54312 sw
tri 51149 54187 51274 54312 ne
rect 51274 54278 55147 54312
tri 55147 54278 55432 54563 sw
tri 55432 54278 55717 54563 ne
rect 55717 54560 57131 54563
tri 57131 54560 57415 54844 sw
tri 57415 54560 57699 54844 ne
rect 57699 54756 59195 54844
tri 59195 54756 59483 55044 sw
tri 59483 54756 59771 55044 ne
rect 59771 54828 61393 55044
tri 61393 54828 61679 55114 sw
tri 61679 54828 61965 55114 ne
rect 61965 54828 71000 55114
rect 59771 54756 61679 54828
rect 57699 54560 59483 54756
rect 55717 54278 57415 54560
rect 51274 54273 55432 54278
tri 55432 54273 55437 54278 sw
tri 55717 54273 55722 54278 ne
rect 55722 54276 57415 54278
tri 57415 54276 57699 54560 sw
tri 57699 54276 57983 54560 ne
rect 57983 54468 59483 54560
tri 59483 54468 59771 54756 sw
tri 59771 54468 60059 54756 ne
rect 60059 54658 61679 54756
tri 61679 54658 61849 54828 sw
tri 61965 54658 62135 54828 ne
rect 62135 54658 71000 54828
rect 60059 54468 61849 54658
rect 57983 54276 59771 54468
rect 55722 54273 57699 54276
rect 51274 54187 55437 54273
rect 46899 53998 50963 54187
rect 44734 53997 46612 53998
tri 46612 53997 46613 53998 sw
tri 46899 53997 46900 53998 ne
rect 46900 53997 50963 53998
rect 44734 53896 46613 53997
rect 42671 53756 44442 53896
tri 44442 53756 44582 53896 sw
tri 44734 53756 44874 53896 ne
rect 44874 53756 46613 53896
rect 42671 53687 44582 53756
rect 38350 53471 42378 53687
rect 33866 53470 38053 53471
tri 38053 53470 38054 53471 sw
tri 38350 53470 38351 53471 ne
rect 38351 53470 42378 53471
rect 33866 53414 38054 53470
rect 30000 53126 33578 53414
tri 33578 53126 33866 53414 sw
tri 33866 53126 34154 53414 ne
rect 34154 53173 38054 53414
tri 38054 53173 38351 53470 sw
tri 38351 53173 38648 53470 ne
rect 38648 53468 42378 53470
tri 42378 53468 42597 53687 sw
tri 42671 53468 42890 53687 ne
rect 42890 53468 44582 53687
rect 38648 53175 42597 53468
tri 42597 53175 42890 53468 sw
tri 42890 53175 43183 53468 ne
rect 43183 53464 44582 53468
tri 44582 53464 44874 53756 sw
tri 44874 53464 45166 53756 ne
rect 45166 53710 46613 53756
tri 46613 53710 46900 53997 sw
tri 46900 53710 47187 53997 ne
rect 47187 53879 50963 53997
tri 50963 53879 51271 54187 sw
tri 51274 53879 51582 54187 ne
rect 51582 53988 55437 54187
tri 55437 53988 55722 54273 sw
tri 55722 53988 56007 54273 ne
rect 56007 54180 57699 54273
tri 57699 54180 57795 54276 sw
tri 57983 54180 58079 54276 ne
rect 58079 54180 59771 54276
tri 59771 54180 60059 54468 sw
tri 60059 54180 60347 54468 ne
rect 60347 54372 61849 54468
tri 61849 54372 62135 54658 sw
tri 62135 54372 62421 54658 ne
rect 62421 54372 71000 54658
rect 60347 54180 62135 54372
rect 56007 53988 57795 54180
rect 51582 53879 55722 53988
rect 47187 53710 51271 53879
rect 45166 53464 46900 53710
rect 43183 53175 44874 53464
rect 38648 53173 42890 53175
rect 34154 53126 38351 53173
rect 30000 53124 33866 53126
tri 33866 53124 33868 53126 sw
tri 34154 53124 34156 53126 ne
rect 34156 53124 38351 53126
rect 30000 52836 33868 53124
tri 33868 52836 34156 53124 sw
tri 34156 52836 34444 53124 ne
rect 34444 53079 38351 53124
tri 38351 53079 38445 53173 sw
tri 38648 53079 38742 53173 ne
rect 38742 53079 42890 53173
rect 34444 52836 38445 53079
rect 30000 52835 34156 52836
tri 34156 52835 34157 52836 sw
tri 34444 52835 34445 52836 ne
rect 34445 52835 38445 52836
rect 30000 52748 34157 52835
tri 30000 52654 30094 52748 ne
rect 30094 52654 34157 52748
tri 29800 52360 30094 52654 sw
tri 30094 52360 30388 52654 ne
rect 30388 52547 34157 52654
tri 34157 52547 34445 52835 sw
tri 34445 52547 34733 52835 ne
rect 34733 52782 38445 52835
tri 38445 52782 38742 53079 sw
tri 38742 52782 39039 53079 ne
rect 39039 52882 42890 53079
tri 42890 52882 43183 53175 sw
tri 43183 52882 43476 53175 ne
rect 43476 53172 44874 53175
tri 44874 53172 45166 53464 sw
tri 45166 53172 45458 53464 ne
rect 45458 53423 46900 53464
tri 46900 53423 47187 53710 sw
tri 47187 53423 47474 53710 ne
rect 47474 53645 51271 53710
tri 51271 53645 51505 53879 sw
tri 51582 53645 51816 53879 ne
rect 51816 53704 55722 53879
tri 55722 53704 56006 53988 sw
tri 56007 53704 56291 53988 ne
rect 56291 53896 57795 53988
tri 57795 53896 58079 54180 sw
tri 58079 53896 58363 54180 ne
rect 58363 53896 60059 54180
rect 56291 53704 58079 53896
rect 51816 53645 56006 53704
rect 47474 53423 51505 53645
rect 45458 53362 47187 53423
tri 47187 53362 47248 53423 sw
tri 47474 53362 47535 53423 ne
rect 47535 53362 51505 53423
rect 45458 53172 47248 53362
rect 43476 52882 45166 53172
rect 39039 52881 43183 52882
tri 43183 52881 43184 52882 sw
tri 43476 52881 43477 52882 ne
rect 43477 52881 45166 52882
rect 39039 52782 43184 52881
rect 34733 52575 38742 52782
tri 38742 52575 38949 52782 sw
tri 39039 52575 39246 52782 ne
rect 39246 52588 43184 52782
tri 43184 52588 43477 52881 sw
tri 43477 52588 43770 52881 ne
rect 43770 52880 45166 52881
tri 45166 52880 45458 53172 sw
tri 45458 52880 45750 53172 ne
rect 45750 53075 47248 53172
tri 47248 53075 47535 53362 sw
tri 47535 53075 47822 53362 ne
rect 47822 53339 51505 53362
tri 51505 53339 51811 53645 sw
tri 51816 53339 52122 53645 ne
rect 52122 53531 56006 53645
tri 56006 53531 56179 53704 sw
tri 56291 53531 56464 53704 ne
rect 56464 53612 58079 53704
tri 58079 53612 58363 53896 sw
tri 58363 53612 58647 53896 ne
rect 58647 53892 60059 53896
tri 60059 53892 60347 54180 sw
tri 60347 53892 60635 54180 ne
rect 60635 54086 62135 54180
tri 62135 54086 62421 54372 sw
tri 62421 54086 62707 54372 ne
rect 62707 54086 71000 54372
rect 60635 53892 62421 54086
rect 58647 53800 60347 53892
tri 60347 53800 60439 53892 sw
tri 60635 53800 60727 53892 ne
rect 60727 53800 62421 53892
tri 62421 53800 62707 54086 sw
tri 62707 54000 62793 54086 ne
rect 62793 54000 71000 54086
rect 58647 53612 60439 53800
rect 56464 53531 58363 53612
rect 52122 53339 56179 53531
rect 47822 53252 51811 53339
tri 51811 53252 51898 53339 sw
tri 52122 53252 52209 53339 ne
rect 52209 53252 56179 53339
rect 47822 53075 51898 53252
rect 45750 52880 47535 53075
rect 43770 52588 45458 52880
tri 45458 52588 45750 52880 sw
tri 45750 52588 46042 52880 ne
rect 46042 52788 47535 52880
tri 47535 52788 47822 53075 sw
tri 47822 52788 48109 53075 ne
rect 48109 52946 51898 53075
tri 51898 52946 52204 53252 sw
tri 52209 52946 52515 53252 ne
rect 52515 53246 56179 53252
tri 56179 53246 56464 53531 sw
tri 56464 53246 56749 53531 ne
rect 56749 53432 58363 53531
tri 58363 53432 58543 53612 sw
tri 58647 53432 58827 53612 ne
rect 58827 53512 60439 53612
tri 60439 53512 60727 53800 sw
tri 60727 53512 61015 53800 ne
rect 61015 53512 71000 53800
rect 58827 53432 60727 53512
rect 56749 53246 58543 53432
rect 52515 53244 56464 53246
tri 56464 53244 56466 53246 sw
tri 56749 53244 56751 53246 ne
rect 56751 53244 58543 53246
rect 52515 52959 56466 53244
tri 56466 52959 56751 53244 sw
tri 56751 52959 57036 53244 ne
rect 57036 53148 58543 53244
tri 58543 53148 58827 53432 sw
tri 58827 53148 59111 53432 ne
rect 59111 53224 60727 53432
tri 60727 53224 61015 53512 sw
tri 61015 53224 61303 53512 ne
rect 61303 53224 71000 53512
rect 59111 53148 61015 53224
rect 57036 52959 58827 53148
rect 52515 52958 56751 52959
tri 56751 52958 56752 52959 sw
tri 57036 52958 57037 52959 ne
rect 57037 52958 58827 52959
rect 52515 52946 56752 52958
rect 48109 52927 52204 52946
tri 52204 52927 52223 52946 sw
tri 52515 52927 52534 52946 ne
rect 52534 52927 56752 52946
rect 48109 52788 52223 52927
rect 46042 52787 47822 52788
tri 47822 52787 47823 52788 sw
tri 48109 52787 48110 52788 ne
rect 48110 52787 52223 52788
rect 46042 52588 47823 52787
rect 39246 52587 43477 52588
tri 43477 52587 43478 52588 sw
tri 43770 52587 43771 52588 ne
rect 43771 52587 45750 52588
rect 39246 52575 43478 52587
rect 34733 52547 38949 52575
rect 30388 52546 34445 52547
tri 34445 52546 34446 52547 sw
tri 34733 52546 34734 52547 ne
rect 34734 52546 38949 52547
rect 30388 52360 34446 52546
rect 26800 52160 30094 52360
tri 30094 52160 30294 52360 sw
tri 30388 52160 30588 52360 ne
rect 30588 52258 34446 52360
tri 34446 52258 34734 52546 sw
tri 34734 52258 35022 52546 ne
rect 35022 52278 38949 52546
tri 38949 52278 39246 52575 sw
tri 39246 52278 39543 52575 ne
rect 39543 52294 43478 52575
tri 43478 52294 43771 52587 sw
tri 43771 52294 44064 52587 ne
rect 44064 52500 45750 52587
tri 45750 52500 45838 52588 sw
tri 46042 52500 46130 52588 ne
rect 46130 52500 47823 52588
tri 47823 52500 48110 52787 sw
tri 48110 52500 48397 52787 ne
rect 48397 52621 52223 52787
tri 52223 52621 52529 52927 sw
tri 52534 52621 52840 52927 ne
rect 52840 52673 56752 52927
tri 56752 52673 57037 52958 sw
tri 57037 52673 57322 52958 ne
rect 57322 52864 58827 52958
tri 58827 52864 59111 53148 sw
tri 59111 52864 59395 53148 ne
rect 59395 53064 61015 53148
tri 61015 53064 61175 53224 sw
tri 61303 53064 61463 53224 ne
rect 61463 53064 71000 53224
rect 59395 52864 61175 53064
rect 57322 52673 59111 52864
rect 52840 52621 57037 52673
rect 48397 52602 52529 52621
tri 52529 52602 52548 52621 sw
tri 52840 52602 52859 52621 ne
rect 52859 52602 57037 52621
rect 48397 52500 52548 52602
rect 44064 52294 45838 52500
rect 39543 52278 43771 52294
rect 35022 52258 39246 52278
rect 30588 52238 34734 52258
tri 34734 52238 34754 52258 sw
tri 35022 52238 35042 52258 ne
rect 35042 52238 39246 52258
rect 30588 52160 34754 52238
rect 26800 52064 30294 52160
tri 30294 52064 30390 52160 sw
tri 30588 52064 30684 52160 ne
rect 30684 52064 34754 52160
rect 26800 51770 30390 52064
tri 30390 51770 30684 52064 sw
tri 30684 51770 30978 52064 ne
rect 30978 51950 34754 52064
tri 34754 51950 35042 52238 sw
tri 35042 51950 35330 52238 ne
rect 35330 52129 39246 52238
tri 39246 52129 39395 52278 sw
tri 39543 52129 39692 52278 ne
rect 39692 52129 43771 52278
tri 43771 52129 43936 52294 sw
tri 44064 52129 44229 52294 ne
rect 44229 52208 45838 52294
tri 45838 52208 46130 52500 sw
tri 46130 52208 46422 52500 ne
rect 46422 52499 48110 52500
tri 48110 52499 48111 52500 sw
tri 48397 52499 48398 52500 ne
rect 48398 52499 52548 52500
rect 46422 52212 48111 52499
tri 48111 52212 48398 52499 sw
tri 48398 52212 48685 52499 ne
rect 48685 52296 52548 52499
tri 52548 52296 52854 52602 sw
tri 52859 52296 53165 52602 ne
rect 53165 52582 57037 52602
tri 57037 52582 57128 52673 sw
tri 57322 52582 57413 52673 ne
rect 57413 52582 59111 52673
rect 53165 52297 57128 52582
tri 57128 52297 57413 52582 sw
tri 57413 52297 57698 52582 ne
rect 57698 52580 59111 52582
tri 59111 52580 59395 52864 sw
tri 59395 52580 59679 52864 ne
rect 59679 52776 61175 52864
tri 61175 52776 61463 53064 sw
tri 61463 52776 61751 53064 ne
rect 61751 52776 71000 53064
rect 59679 52580 61463 52776
rect 57698 52297 59395 52580
rect 53165 52296 57413 52297
rect 48685 52277 52854 52296
tri 52854 52277 52873 52296 sw
tri 53165 52277 53184 52296 ne
rect 53184 52295 57413 52296
tri 57413 52295 57415 52297 sw
tri 57698 52295 57700 52297 ne
rect 57700 52296 59395 52297
tri 59395 52296 59679 52580 sw
tri 59679 52296 59963 52580 ne
rect 59963 52488 61463 52580
tri 61463 52488 61751 52776 sw
tri 61751 52488 62039 52776 ne
rect 62039 52488 71000 52776
rect 59963 52296 61751 52488
rect 57700 52295 59679 52296
rect 53184 52277 57415 52295
rect 48685 52212 52873 52277
rect 46422 52208 48398 52212
rect 44229 52129 46130 52208
rect 35330 51950 39395 52129
rect 30978 51949 35042 51950
tri 35042 51949 35043 51950 sw
tri 35330 51949 35331 51950 ne
rect 35331 51949 39395 51950
rect 30978 51770 35043 51949
rect 26800 51605 30684 51770
tri 30684 51605 30849 51770 sw
tri 30978 51605 31143 51770 ne
rect 31143 51661 35043 51770
tri 35043 51661 35331 51949 sw
tri 35331 51661 35619 51949 ne
rect 35619 51832 39395 51949
tri 39395 51832 39692 52129 sw
tri 39692 51832 39989 52129 ne
rect 39989 51836 43936 52129
tri 43936 51836 44229 52129 sw
tri 44229 51836 44522 52129 ne
rect 44522 51916 46130 52129
tri 46130 51916 46422 52208 sw
tri 46422 51916 46714 52208 ne
rect 46714 51925 48398 52208
tri 48398 51925 48685 52212 sw
tri 48685 51925 48972 52212 ne
rect 48972 51971 52873 52212
tri 52873 51971 53179 52277 sw
tri 53184 51971 53490 52277 ne
rect 53490 52010 57415 52277
tri 57415 52010 57700 52295 sw
tri 57700 52010 57985 52295 ne
rect 57985 52200 59679 52295
tri 59679 52200 59775 52296 sw
tri 59963 52200 60059 52296 ne
rect 60059 52200 61751 52296
tri 61751 52200 62039 52488 sw
tri 62039 52400 62127 52488 ne
rect 62127 52400 71000 52488
rect 57985 52010 59775 52200
rect 53490 52008 57700 52010
tri 57700 52008 57702 52010 sw
tri 57985 52008 57987 52010 ne
rect 57987 52008 59775 52010
rect 53490 51971 57702 52008
rect 48972 51952 53179 51971
tri 53179 51952 53198 51971 sw
tri 53490 51952 53509 51971 ne
rect 53509 51952 57702 51971
rect 48972 51925 53198 51952
rect 46714 51924 48685 51925
tri 48685 51924 48686 51925 sw
tri 48972 51924 48973 51925 ne
rect 48973 51924 53198 51925
rect 46714 51916 48686 51924
rect 44522 51836 46422 51916
rect 39989 51835 44229 51836
tri 44229 51835 44230 51836 sw
tri 44522 51835 44523 51836 ne
rect 44523 51835 46422 51836
rect 39989 51832 44230 51835
rect 35619 51831 39692 51832
tri 39692 51831 39693 51832 sw
tri 39989 51831 39990 51832 ne
rect 39990 51831 44230 51832
rect 35619 51661 39693 51831
rect 31143 51660 35331 51661
tri 35331 51660 35332 51661 sw
tri 35619 51660 35620 51661 ne
rect 35620 51660 39693 51661
rect 31143 51605 35332 51660
rect 26800 51410 30849 51605
tri 30849 51410 31044 51605 sw
tri 31143 51410 31338 51605 ne
rect 31338 51410 35332 51605
tri 26800 51320 26890 51410 ne
rect 26890 51320 31044 51410
tri 26600 51120 26800 51320 sw
tri 26890 51120 27090 51320 ne
rect 27090 51120 31044 51320
rect 25200 50941 26800 51120
tri 26800 50941 26979 51120 sw
tri 27090 50941 27269 51120 ne
rect 27269 51116 31044 51120
tri 31044 51116 31338 51410 sw
tri 31338 51116 31632 51410 ne
rect 31632 51372 35332 51410
tri 35332 51372 35620 51660 sw
tri 35620 51372 35908 51660 ne
rect 35908 51534 39693 51660
tri 39693 51534 39990 51831 sw
tri 39990 51534 40287 51831 ne
rect 40287 51542 44230 51831
tri 44230 51542 44523 51835 sw
tri 44523 51542 44816 51835 ne
rect 44816 51776 46422 51835
tri 46422 51776 46562 51916 sw
tri 46714 51776 46854 51916 ne
rect 46854 51776 48686 51916
rect 44816 51542 46562 51776
rect 40287 51534 44523 51542
rect 35908 51533 39990 51534
tri 39990 51533 39991 51534 sw
tri 40287 51533 40288 51534 ne
rect 40288 51533 44523 51534
rect 35908 51372 39991 51533
rect 31632 51220 35620 51372
tri 35620 51220 35772 51372 sw
tri 35908 51220 36060 51372 ne
rect 36060 51236 39991 51372
tri 39991 51236 40288 51533 sw
tri 40288 51236 40585 51533 ne
rect 40585 51249 44523 51533
tri 44523 51249 44816 51542 sw
tri 44816 51249 45109 51542 ne
rect 45109 51484 46562 51542
tri 46562 51484 46854 51776 sw
tri 46854 51484 47146 51776 ne
rect 47146 51637 48686 51776
tri 48686 51637 48973 51924 sw
tri 48973 51637 49260 51924 ne
rect 49260 51645 53198 51924
tri 53198 51645 53505 51952 sw
tri 53509 51645 53816 51952 ne
rect 53816 51723 57702 51952
tri 57702 51723 57987 52008 sw
tri 57987 51723 58272 52008 ne
rect 58272 51916 59775 52008
tri 59775 51916 60059 52200 sw
tri 60059 51916 60343 52200 ne
rect 60343 51916 71000 52200
rect 58272 51723 60059 51916
rect 53816 51722 57987 51723
tri 57987 51722 57988 51723 sw
tri 58272 51722 58273 51723 ne
rect 58273 51722 60059 51723
rect 53816 51645 57988 51722
rect 49260 51637 53505 51645
rect 47146 51484 48973 51637
rect 45109 51249 46854 51484
rect 40585 51236 44816 51249
rect 36060 51234 40288 51236
tri 40288 51234 40290 51236 sw
tri 40585 51234 40587 51236 ne
rect 40587 51234 44816 51236
rect 36060 51220 40290 51234
rect 31632 51116 35772 51220
rect 27269 50941 31338 51116
rect 25200 50740 26979 50941
tri 25200 50651 25289 50740 ne
rect 25289 50651 26979 50740
tri 26979 50651 27269 50941 sw
tri 27269 50651 27559 50941 ne
rect 27559 50926 31338 50941
tri 31338 50926 31528 51116 sw
tri 31632 50926 31822 51116 ne
rect 31822 50932 35772 51116
tri 35772 50932 36060 51220 sw
tri 36060 50932 36348 51220 ne
rect 36348 50937 40290 51220
tri 40290 50937 40587 51234 sw
tri 40587 50937 40884 51234 ne
rect 40884 50956 44816 51234
tri 44816 50956 45109 51249 sw
tri 45109 50956 45402 51249 ne
rect 45402 51192 46854 51249
tri 46854 51192 47146 51484 sw
tri 47146 51192 47438 51484 ne
rect 47438 51383 48973 51484
tri 48973 51383 49227 51637 sw
tri 49260 51383 49514 51637 ne
rect 49514 51383 53505 51637
rect 47438 51306 49227 51383
tri 49227 51306 49304 51383 sw
tri 49514 51306 49591 51383 ne
rect 49591 51353 53505 51383
tri 53505 51353 53797 51645 sw
tri 53816 51353 54108 51645 ne
rect 54108 51437 57988 51645
tri 57988 51437 58273 51722 sw
tri 58273 51437 58558 51722 ne
rect 58558 51632 60059 51722
tri 60059 51632 60343 51916 sw
tri 60343 51632 60627 51916 ne
rect 60627 51632 71000 51916
rect 58558 51452 60343 51632
tri 60343 51452 60523 51632 sw
tri 60627 51452 60807 51632 ne
rect 60807 51452 71000 51632
rect 58558 51437 60523 51452
rect 54108 51353 58273 51437
rect 49591 51306 53797 51353
tri 53797 51306 53844 51353 sw
tri 54108 51306 54155 51353 ne
rect 54155 51306 58273 51353
rect 47438 51192 49304 51306
rect 45402 50956 47146 51192
rect 40884 50937 45109 50956
rect 36348 50936 40587 50937
tri 40587 50936 40588 50937 sw
tri 40884 50936 40885 50937 ne
rect 40885 50936 45109 50937
rect 36348 50932 40588 50936
rect 31822 50926 36060 50932
rect 27559 50651 31528 50926
tri 25000 50362 25289 50651 sw
tri 25289 50362 25578 50651 ne
rect 25578 50650 27269 50651
tri 27269 50650 27270 50651 sw
tri 27559 50650 27560 50651 ne
rect 27560 50650 31528 50651
rect 25578 50362 27270 50650
rect 23600 50073 25289 50362
tri 25289 50073 25578 50362 sw
tri 25578 50073 25867 50362 ne
rect 25867 50360 27270 50362
tri 27270 50360 27560 50650 sw
tri 27560 50360 27850 50650 ne
rect 27850 50632 31528 50650
tri 31528 50632 31822 50926 sw
tri 31822 50632 32116 50926 ne
rect 32116 50792 36060 50926
tri 36060 50792 36200 50932 sw
tri 36348 50792 36488 50932 ne
rect 36488 50792 40588 50932
rect 32116 50632 36200 50792
rect 27850 50424 31822 50632
tri 31822 50424 32030 50632 sw
tri 32116 50424 32324 50632 ne
rect 32324 50504 36200 50632
tri 36200 50504 36488 50792 sw
tri 36488 50504 36776 50792 ne
rect 36776 50639 40588 50792
tri 40588 50639 40885 50936 sw
tri 40885 50639 41182 50936 ne
rect 41182 50901 45109 50936
tri 45109 50901 45164 50956 sw
tri 45402 50901 45457 50956 ne
rect 45457 50901 47146 50956
rect 41182 50639 45164 50901
rect 36776 50638 40885 50639
tri 40885 50638 40886 50639 sw
tri 41182 50638 41183 50639 ne
rect 41183 50638 45164 50639
rect 36776 50504 40886 50638
rect 32324 50424 36488 50504
rect 27850 50360 32030 50424
rect 25867 50359 27560 50360
tri 27560 50359 27561 50360 sw
tri 27850 50359 27851 50360 ne
rect 27851 50359 32030 50360
rect 25867 50073 27561 50359
rect 23600 50071 25578 50073
tri 23600 49974 23697 50071 ne
rect 23697 49974 25578 50071
tri 23400 49774 23600 49974 sw
tri 23697 49774 23897 49974 ne
rect 23897 49918 25578 49974
tri 25578 49918 25733 50073 sw
tri 25867 49918 26022 50073 ne
rect 26022 50069 27561 50073
tri 27561 50069 27851 50359 sw
tri 27851 50069 28141 50359 ne
rect 28141 50130 32030 50359
tri 32030 50130 32324 50424 sw
tri 32324 50130 32618 50424 ne
rect 32618 50261 36488 50424
tri 36488 50261 36731 50504 sw
tri 36776 50261 37019 50504 ne
rect 37019 50341 40886 50504
tri 40886 50341 41183 50638 sw
tri 41183 50341 41480 50638 ne
rect 41480 50608 45164 50638
tri 45164 50608 45457 50901 sw
tri 45457 50608 45750 50901 ne
rect 45750 50900 47146 50901
tri 47146 50900 47438 51192 sw
tri 47438 50900 47730 51192 ne
rect 47730 51019 49304 51192
tri 49304 51019 49591 51306 sw
tri 49591 51019 49878 51306 ne
rect 49878 51019 53844 51306
rect 47730 50900 49591 51019
rect 45750 50608 47438 50900
tri 47438 50608 47730 50900 sw
tri 47730 50608 48022 50900 ne
rect 48022 50807 49591 50900
tri 49591 50807 49803 51019 sw
tri 49878 50807 50090 51019 ne
rect 50090 51004 53844 51019
tri 53844 51004 54146 51306 sw
tri 54155 51004 54457 51306 ne
rect 54457 51175 58273 51306
tri 58273 51175 58535 51437 sw
tri 58558 51175 58820 51437 ne
rect 58820 51175 60523 51437
rect 54457 51004 58535 51175
rect 50090 50807 54146 51004
rect 48022 50608 49803 50807
rect 41480 50607 45457 50608
tri 45457 50607 45458 50608 sw
tri 45750 50607 45751 50608 ne
rect 45751 50607 47730 50608
rect 41480 50341 45458 50607
rect 37019 50261 41183 50341
rect 32618 50130 36731 50261
rect 28141 50069 32324 50130
rect 26022 49918 27851 50069
rect 23897 49774 25733 49918
rect 20400 49676 23600 49774
tri 23600 49676 23698 49774 sw
tri 23897 49676 23995 49774 ne
rect 23995 49676 25733 49774
rect 20400 49379 23698 49676
tri 23698 49379 23995 49676 sw
tri 23995 49379 24292 49676 ne
rect 24292 49629 25733 49676
tri 25733 49629 26022 49918 sw
tri 26022 49629 26311 49918 ne
rect 26311 49779 27851 49918
tri 27851 49779 28141 50069 sw
tri 28141 49779 28431 50069 ne
rect 28431 50044 32324 50069
tri 32324 50044 32410 50130 sw
tri 32618 50044 32704 50130 ne
rect 32704 50044 36731 50130
rect 28431 49779 32410 50044
rect 26311 49778 28141 49779
tri 28141 49778 28142 49779 sw
tri 28431 49778 28432 49779 ne
rect 28432 49778 32410 49779
rect 26311 49629 28142 49778
rect 24292 49379 26022 49629
rect 20400 49155 23995 49379
tri 23995 49155 24219 49379 sw
tri 24292 49155 24516 49379 ne
rect 24516 49340 26022 49379
tri 26022 49340 26311 49629 sw
tri 26311 49340 26600 49629 ne
rect 26600 49488 28142 49629
tri 28142 49488 28432 49778 sw
tri 28432 49488 28722 49778 ne
rect 28722 49750 32410 49778
tri 32410 49750 32704 50044 sw
tri 32704 49750 32998 50044 ne
rect 32998 49973 36731 50044
tri 36731 49973 37019 50261 sw
tri 37019 49973 37307 50261 ne
rect 37307 50122 41183 50261
tri 41183 50122 41402 50341 sw
tri 41480 50122 41699 50341 ne
rect 41699 50314 45458 50341
tri 45458 50314 45751 50607 sw
tri 45751 50314 46044 50607 ne
rect 46044 50520 47730 50607
tri 47730 50520 47818 50608 sw
tri 48022 50520 48110 50608 ne
rect 48110 50520 49803 50608
tri 49803 50520 50090 50807 sw
tri 50090 50520 50377 50807 ne
rect 50377 50703 54146 50807
tri 54146 50703 54447 51004 sw
tri 54457 50703 54758 51004 ne
rect 54758 50890 58535 51004
tri 58535 50890 58820 51175 sw
tri 58820 50890 59105 51175 ne
rect 59105 51168 60523 51175
tri 60523 51168 60807 51452 sw
tri 60807 51168 61091 51452 ne
rect 61091 51168 71000 51452
rect 59105 50890 60807 51168
rect 54758 50888 58820 50890
tri 58820 50888 58822 50890 sw
tri 59105 50888 59107 50890 ne
rect 59107 50888 60807 50890
rect 54758 50703 58822 50888
rect 50377 50520 54447 50703
rect 46044 50314 47818 50520
rect 41699 50313 45751 50314
tri 45751 50313 45752 50314 sw
tri 46044 50313 46045 50314 ne
rect 46045 50313 47818 50314
rect 41699 50122 45752 50313
rect 37307 49973 41402 50122
rect 32998 49888 37019 49973
tri 37019 49888 37104 49973 sw
tri 37307 49888 37392 49973 ne
rect 37392 49888 41402 49973
rect 32998 49750 37104 49888
rect 28722 49749 32704 49750
tri 32704 49749 32705 49750 sw
tri 32998 49749 32999 49750 ne
rect 32999 49749 37104 49750
rect 28722 49488 32705 49749
rect 26600 49340 28432 49488
rect 24516 49155 26311 49340
rect 20400 48858 24219 49155
tri 24219 48858 24516 49155 sw
tri 24516 48858 24813 49155 ne
rect 24813 49051 26311 49155
tri 26311 49051 26600 49340 sw
tri 26600 49051 26889 49340 ne
rect 26889 49251 28432 49340
tri 28432 49251 28669 49488 sw
tri 28722 49251 28959 49488 ne
rect 28959 49455 32705 49488
tri 32705 49455 32999 49749 sw
tri 32999 49455 33293 49749 ne
rect 33293 49600 37104 49749
tri 37104 49600 37392 49888 sw
tri 37392 49600 37680 49888 ne
rect 37680 49879 41402 49888
tri 41402 49879 41645 50122 sw
tri 41699 49879 41942 50122 ne
rect 41942 50020 45752 50122
tri 45752 50020 46045 50313 sw
tri 46045 50020 46338 50313 ne
rect 46338 50228 47818 50313
tri 47818 50228 48110 50520 sw
tri 48110 50228 48402 50520 ne
rect 48402 50519 50090 50520
tri 50090 50519 50091 50520 sw
tri 50377 50519 50378 50520 ne
rect 50378 50519 54447 50520
rect 48402 50232 50091 50519
tri 50091 50232 50378 50519 sw
tri 50378 50232 50665 50519 ne
rect 50665 50397 54447 50519
tri 54447 50397 54753 50703 sw
tri 54758 50397 55064 50703 ne
rect 55064 50603 58822 50703
tri 58822 50603 59107 50888 sw
tri 59107 50603 59392 50888 ne
rect 59392 50884 60807 50888
tri 60807 50884 61091 51168 sw
tri 61091 50884 61375 51168 ne
rect 61375 50884 71000 51168
rect 59392 50603 61091 50884
rect 55064 50602 59107 50603
tri 59107 50602 59108 50603 sw
tri 59392 50602 59393 50603 ne
rect 59393 50602 61091 50603
rect 55064 50397 59108 50602
rect 50665 50378 54753 50397
tri 54753 50378 54772 50397 sw
tri 55064 50378 55083 50397 ne
rect 55083 50378 59108 50397
rect 50665 50232 54772 50378
rect 48402 50228 50378 50232
rect 46338 50020 48110 50228
rect 41942 49879 46045 50020
rect 37680 49824 41645 49879
tri 41645 49824 41700 49879 sw
tri 41942 49824 41997 49879 ne
rect 41997 49824 46045 49879
rect 37680 49600 41700 49824
rect 33293 49455 37392 49600
rect 28959 49454 32999 49455
tri 32999 49454 33000 49455 sw
tri 33293 49454 33294 49455 ne
rect 33294 49454 37392 49455
rect 28959 49251 33000 49454
rect 26889 49051 28669 49251
rect 24813 49049 26600 49051
tri 26600 49049 26602 49051 sw
tri 26889 49049 26891 49051 ne
rect 26891 49049 28669 49051
rect 24813 48858 26602 49049
rect 20400 48730 24516 48858
tri 20400 48648 20482 48730 ne
rect 20482 48648 24516 48730
tri 20200 48366 20482 48648 sw
tri 20482 48366 20764 48648 ne
rect 20764 48561 24516 48648
tri 24516 48561 24813 48858 sw
tri 24813 48561 25110 48858 ne
rect 25110 48760 26602 48858
tri 26602 48760 26891 49049 sw
tri 26891 48760 27180 49049 ne
rect 27180 48961 28669 49049
tri 28669 48961 28959 49251 sw
tri 28959 48961 29249 49251 ne
rect 29249 49160 33000 49251
tri 33000 49160 33294 49454 sw
tri 33294 49160 33588 49454 ne
rect 33588 49393 37392 49454
tri 37392 49393 37599 49600 sw
tri 37680 49393 37887 49600 ne
rect 37887 49527 41700 49600
tri 41700 49527 41997 49824 sw
tri 41997 49527 42294 49824 ne
rect 42294 49727 46045 49824
tri 46045 49727 46338 50020 sw
tri 46338 49727 46631 50020 ne
rect 46631 49936 48110 50020
tri 48110 49936 48402 50228 sw
tri 48402 49936 48694 50228 ne
rect 48694 50042 50378 50228
tri 50378 50042 50568 50232 sw
tri 50665 50042 50855 50232 ne
rect 50855 50072 54772 50232
tri 54772 50072 55078 50378 sw
tri 55083 50072 55389 50378 ne
rect 55389 50317 59108 50378
tri 59108 50317 59393 50602 sw
tri 59393 50317 59678 50602 ne
rect 59678 50600 61091 50602
tri 61091 50600 61375 50884 sw
tri 61375 50800 61459 50884 ne
rect 61459 50800 71000 50884
rect 59678 50317 71000 50600
rect 55389 50249 59393 50317
tri 59393 50249 59461 50317 sw
tri 59678 50249 59746 50317 ne
rect 59746 50249 71000 50317
rect 55389 50072 59461 50249
rect 50855 50042 55078 50072
rect 48694 49936 50568 50042
rect 46631 49796 48402 49936
tri 48402 49796 48542 49936 sw
tri 48694 49796 48834 49936 ne
rect 48834 49796 50568 49936
rect 46631 49727 48542 49796
rect 42294 49527 46338 49727
rect 37887 49525 41997 49527
tri 41997 49525 41999 49527 sw
tri 42294 49525 42296 49527 ne
rect 42296 49525 46338 49527
rect 37887 49393 41999 49525
rect 33588 49160 37599 49393
rect 29249 49159 33294 49160
tri 33294 49159 33295 49160 sw
tri 33588 49159 33589 49160 ne
rect 33589 49159 37599 49160
rect 29249 48961 33295 49159
rect 27180 48760 28959 48961
rect 25110 48561 26891 48760
rect 20764 48374 24813 48561
tri 24813 48374 25000 48561 sw
tri 25110 48374 25297 48561 ne
rect 25297 48471 26891 48561
tri 26891 48471 27180 48760 sw
tri 27180 48471 27469 48760 ne
rect 27469 48671 28959 48760
tri 28959 48671 29249 48961 sw
tri 29249 48671 29539 48961 ne
rect 29539 48865 33295 48961
tri 33295 48865 33589 49159 sw
tri 33589 48865 33883 49159 ne
rect 33883 49105 37599 49159
tri 37599 49105 37887 49393 sw
tri 37887 49105 38175 49393 ne
rect 38175 49228 41999 49393
tri 41999 49228 42296 49525 sw
tri 42296 49228 42593 49525 ne
rect 42593 49508 46338 49525
tri 46338 49508 46557 49727 sw
tri 46631 49508 46850 49727 ne
rect 46850 49508 48542 49727
rect 42593 49228 46557 49508
rect 38175 49227 42296 49228
tri 42296 49227 42297 49228 sw
tri 42593 49227 42594 49228 ne
rect 42594 49227 46557 49228
rect 38175 49105 42297 49227
rect 33883 48929 37887 49105
tri 37887 48929 38063 49105 sw
tri 38175 48929 38351 49105 ne
rect 38351 48930 42297 49105
tri 42297 48930 42594 49227 sw
tri 42594 48930 42891 49227 ne
rect 42891 49215 46557 49227
tri 46557 49215 46850 49508 sw
tri 46850 49215 47143 49508 ne
rect 47143 49504 48542 49508
tri 48542 49504 48834 49796 sw
tri 48834 49504 49126 49796 ne
rect 49126 49755 50568 49796
tri 50568 49755 50855 50042 sw
tri 50855 49755 51142 50042 ne
rect 51142 49938 55078 50042
tri 55078 49938 55212 50072 sw
tri 55389 49938 55523 50072 ne
rect 55523 49964 59461 50072
tri 59461 49964 59746 50249 sw
tri 59746 49964 60031 50249 ne
rect 60031 49964 71000 50249
rect 55523 49938 59746 49964
rect 51142 49755 55212 49938
rect 49126 49504 50855 49755
rect 47143 49215 48834 49504
rect 42891 48930 46850 49215
rect 38351 48929 42594 48930
rect 33883 48865 38063 48929
rect 29539 48864 33589 48865
tri 33589 48864 33590 48865 sw
tri 33883 48864 33884 48865 ne
rect 33884 48864 38063 48865
rect 29539 48671 33590 48864
rect 27469 48670 29249 48671
tri 29249 48670 29250 48671 sw
tri 29539 48670 29540 48671 ne
rect 29540 48670 33590 48671
rect 27469 48471 29250 48670
rect 25297 48380 27180 48471
tri 27180 48380 27271 48471 sw
tri 27469 48380 27560 48471 ne
rect 27560 48380 29250 48471
tri 29250 48380 29540 48670 sw
tri 29540 48380 29830 48670 ne
rect 29830 48570 33590 48670
tri 33590 48570 33884 48864 sw
tri 33884 48570 34178 48864 ne
rect 34178 48641 38063 48864
tri 38063 48641 38351 48929 sw
tri 38351 48641 38639 48929 ne
rect 38639 48835 42594 48929
tri 42594 48835 42689 48930 sw
tri 42891 48835 42986 48930 ne
rect 42986 48922 46850 48930
tri 46850 48922 47143 49215 sw
tri 47143 48922 47436 49215 ne
rect 47436 49212 48834 49215
tri 48834 49212 49126 49504 sw
tri 49126 49212 49418 49504 ne
rect 49418 49468 50855 49504
tri 50855 49468 51142 49755 sw
tri 51142 49468 51429 49755 ne
rect 51429 49636 55212 49755
tri 55212 49636 55514 49938 sw
tri 55523 49636 55825 49938 ne
rect 55825 49743 59746 49938
tri 59746 49743 59967 49964 sw
tri 60031 49743 60252 49964 ne
rect 60252 49743 71000 49964
rect 55825 49636 59967 49743
rect 51429 49468 55514 49636
rect 49418 49402 51142 49468
tri 51142 49402 51208 49468 sw
tri 51429 49402 51495 49468 ne
rect 51495 49402 55514 49468
tri 55514 49402 55748 49636 sw
tri 55825 49402 56059 49636 ne
rect 56059 49575 59967 49636
tri 59967 49575 60135 49743 sw
tri 60252 49575 60420 49743 ne
rect 60420 49575 71000 49743
rect 56059 49402 60135 49575
rect 49418 49212 51208 49402
rect 47436 48922 49126 49212
rect 42986 48920 47143 48922
tri 47143 48920 47145 48922 sw
tri 47436 48920 47438 48922 ne
rect 47438 48920 49126 48922
tri 49126 48920 49418 49212 sw
tri 49418 48920 49710 49212 ne
rect 49710 49115 51208 49212
tri 51208 49115 51495 49402 sw
tri 51495 49115 51782 49402 ne
rect 51782 49115 55748 49402
rect 49710 48920 51495 49115
rect 42986 48835 47145 48920
rect 38639 48641 42689 48835
rect 34178 48640 38351 48641
tri 38351 48640 38352 48641 sw
tri 38639 48640 38640 48641 ne
rect 38640 48640 42689 48641
rect 34178 48570 38352 48640
rect 29830 48568 33884 48570
tri 33884 48568 33886 48570 sw
tri 34178 48568 34180 48570 ne
rect 34180 48568 38352 48570
rect 29830 48380 33886 48568
rect 25297 48374 27271 48380
rect 20764 48366 25000 48374
rect 17200 48166 20482 48366
tri 20482 48166 20682 48366 sw
tri 20764 48166 20964 48366 ne
rect 20964 48166 25000 48366
rect 17200 48082 20682 48166
tri 20682 48082 20766 48166 sw
tri 20964 48082 21048 48166 ne
rect 21048 48082 25000 48166
rect 17200 47800 20766 48082
tri 20766 47800 21048 48082 sw
tri 21048 47800 21330 48082 ne
rect 21330 48077 25000 48082
tri 25000 48077 25297 48374 sw
tri 25297 48077 25594 48374 ne
rect 25594 48091 27271 48374
tri 27271 48091 27560 48380 sw
tri 27560 48091 27849 48380 ne
rect 27849 48379 29540 48380
tri 29540 48379 29541 48380 sw
tri 29830 48379 29831 48380 ne
rect 29831 48379 33886 48380
rect 27849 48091 29541 48379
rect 25594 48077 27560 48091
rect 21330 48076 25297 48077
tri 25297 48076 25298 48077 sw
tri 25594 48076 25595 48077 ne
rect 25595 48076 27560 48077
rect 21330 47800 25298 48076
rect 17200 47798 21048 47800
tri 21048 47798 21050 47800 sw
tri 21330 47798 21332 47800 ne
rect 21332 47798 25298 47800
rect 17200 47516 21050 47798
tri 21050 47516 21332 47798 sw
tri 21332 47516 21614 47798 ne
rect 21614 47779 25298 47798
tri 25298 47779 25595 48076 sw
tri 25595 47779 25892 48076 ne
rect 25892 47802 27560 48076
tri 27560 47802 27849 48091 sw
tri 27849 47802 28138 48091 ne
rect 28138 48089 29541 48091
tri 29541 48089 29831 48379 sw
tri 29831 48089 30121 48379 ne
rect 30121 48274 33886 48379
tri 33886 48274 34180 48568 sw
tri 34180 48274 34474 48568 ne
rect 34474 48352 38352 48568
tri 38352 48352 38640 48640 sw
tri 38640 48352 38928 48640 ne
rect 38928 48538 42689 48640
tri 42689 48538 42986 48835 sw
tri 42986 48538 43283 48835 ne
rect 43283 48627 47145 48835
tri 47145 48627 47438 48920 sw
tri 47438 48627 47731 48920 ne
rect 47731 48628 49418 48920
tri 49418 48628 49710 48920 sw
tri 49710 48628 50002 48920 ne
rect 50002 48828 51495 48920
tri 51495 48828 51782 49115 sw
tri 51782 48828 52069 49115 ne
rect 52069 49096 55748 49115
tri 55748 49096 56054 49402 sw
tri 56059 49096 56365 49402 ne
rect 56365 49290 60135 49402
tri 60135 49290 60420 49575 sw
tri 60420 49290 60705 49575 ne
rect 60705 49290 71000 49575
rect 56365 49288 60420 49290
tri 60420 49288 60422 49290 sw
tri 60705 49288 60707 49290 ne
rect 60707 49288 71000 49290
rect 56365 49096 60422 49288
rect 52069 49010 56054 49096
tri 56054 49010 56140 49096 sw
tri 56365 49010 56451 49096 ne
rect 56451 49010 60422 49096
rect 52069 48828 56140 49010
rect 50002 48827 51782 48828
tri 51782 48827 51783 48828 sw
tri 52069 48827 52070 48828 ne
rect 52070 48827 56140 48828
rect 50002 48628 51783 48827
rect 47731 48627 49710 48628
rect 43283 48538 47438 48627
rect 38928 48352 42986 48538
rect 34474 48351 38640 48352
tri 38640 48351 38641 48352 sw
tri 38928 48351 38929 48352 ne
rect 38929 48351 42986 48352
rect 34474 48274 38641 48351
rect 30121 48089 34180 48274
rect 28138 48020 29831 48089
tri 29831 48020 29900 48089 sw
tri 30121 48020 30190 48089 ne
rect 30190 48020 34180 48089
tri 34180 48020 34434 48274 sw
tri 34474 48020 34728 48274 ne
rect 34728 48063 38641 48274
tri 38641 48063 38929 48351 sw
tri 38929 48063 39217 48351 ne
rect 39217 48333 42986 48351
tri 42986 48333 43191 48538 sw
tri 43283 48333 43488 48538 ne
rect 43488 48334 47438 48538
tri 47438 48334 47731 48627 sw
tri 47731 48334 48024 48627 ne
rect 48024 48540 49710 48627
tri 49710 48540 49798 48628 sw
tri 50002 48540 50090 48628 ne
rect 50090 48540 51783 48628
tri 51783 48540 52070 48827 sw
tri 52070 48540 52357 48827 ne
rect 52357 48704 56140 48827
tri 56140 48704 56446 49010 sw
tri 56451 48704 56757 49010 ne
rect 56757 49003 60422 49010
tri 60422 49003 60707 49288 sw
tri 60707 49200 60795 49288 ne
rect 60795 49200 71000 49288
rect 56757 49000 60707 49003
tri 60707 49000 60710 49003 sw
rect 56757 48704 71000 49000
rect 52357 48684 56446 48704
tri 56446 48684 56466 48704 sw
tri 56757 48684 56777 48704 ne
rect 56777 48684 71000 48704
rect 52357 48540 56466 48684
rect 48024 48334 49798 48540
rect 43488 48333 47731 48334
rect 39217 48063 43191 48333
rect 34728 48061 38929 48063
tri 38929 48061 38931 48063 sw
tri 39217 48061 39219 48063 ne
rect 39219 48061 43191 48063
rect 34728 48020 38931 48061
rect 28138 47802 29900 48020
rect 25892 47779 27849 47802
rect 21614 47516 25595 47779
rect 17200 47515 21332 47516
tri 21332 47515 21333 47516 sw
tri 21614 47515 21615 47516 ne
rect 21615 47515 25595 47516
rect 17200 47404 21333 47515
tri 17200 47312 17292 47404 ne
rect 17292 47312 21333 47404
tri 17000 47020 17292 47312 sw
tri 17292 47020 17584 47312 ne
rect 17584 47233 21333 47312
tri 21333 47233 21615 47515 sw
tri 21615 47233 21897 47515 ne
rect 21897 47482 25595 47515
tri 25595 47482 25892 47779 sw
tri 25892 47482 26189 47779 ne
rect 26189 47647 27849 47779
tri 27849 47647 28004 47802 sw
tri 28138 47647 28293 47802 ne
rect 28293 47730 29900 47802
tri 29900 47730 30190 48020 sw
tri 30190 47730 30480 48020 ne
rect 30480 47730 34434 48020
rect 28293 47647 30190 47730
rect 26189 47482 28004 47647
rect 21897 47376 25892 47482
tri 25892 47376 25998 47482 sw
tri 26189 47376 26295 47482 ne
rect 26295 47376 28004 47482
rect 21897 47233 25998 47376
rect 17584 47232 21615 47233
tri 21615 47232 21616 47233 sw
tri 21897 47232 21898 47233 ne
rect 21898 47232 25998 47233
rect 17584 47020 21616 47232
rect 14000 46820 17292 47020
tri 17292 46820 17492 47020 sw
tri 17584 46820 17784 47020 ne
rect 17784 46950 21616 47020
tri 21616 46950 21898 47232 sw
tri 21898 46950 22180 47232 ne
rect 22180 47079 25998 47232
tri 25998 47079 26295 47376 sw
tri 26295 47079 26592 47376 ne
rect 26592 47358 28004 47376
tri 28004 47358 28293 47647 sw
tri 28293 47358 28582 47647 ne
rect 28582 47508 30190 47647
tri 30190 47508 30412 47730 sw
tri 30480 47508 30702 47730 ne
rect 30702 47726 34434 47730
tri 34434 47726 34728 48020 sw
tri 34728 47726 35022 48020 ne
rect 35022 47773 38931 48020
tri 38931 47773 39219 48061 sw
tri 39219 47773 39507 48061 ne
rect 39507 48036 43191 48061
tri 43191 48036 43488 48333 sw
tri 43488 48036 43785 48333 ne
rect 43785 48180 47731 48333
tri 47731 48180 47885 48334 sw
tri 48024 48180 48178 48334 ne
rect 48178 48248 49798 48334
tri 49798 48248 50090 48540 sw
tri 50090 48248 50382 48540 ne
rect 50382 48539 52070 48540
tri 52070 48539 52071 48540 sw
tri 52357 48539 52358 48540 ne
rect 52358 48539 56466 48540
rect 50382 48252 52071 48539
tri 52071 48252 52358 48539 sw
tri 52358 48252 52645 48539 ne
rect 52645 48378 56466 48539
tri 56466 48378 56772 48684 sw
tri 56777 48378 57083 48684 ne
rect 57083 48378 71000 48684
rect 52645 48359 56772 48378
tri 56772 48359 56791 48378 sw
tri 57083 48359 57102 48378 ne
rect 57102 48359 71000 48378
rect 52645 48252 56791 48359
rect 50382 48248 52358 48252
rect 48178 48180 50090 48248
rect 43785 48036 47885 48180
rect 39507 47886 43488 48036
tri 43488 47886 43638 48036 sw
tri 43785 47886 43935 48036 ne
rect 43935 47887 47885 48036
tri 47885 47887 48178 48180 sw
tri 48178 47887 48471 48180 ne
rect 48471 47956 50090 48180
tri 50090 47956 50382 48248 sw
tri 50382 47956 50674 48248 ne
rect 50674 47965 52358 48248
tri 52358 47965 52645 48252 sw
tri 52645 47965 52932 48252 ne
rect 52932 48053 56791 48252
tri 56791 48053 57097 48359 sw
tri 57102 48053 57408 48359 ne
rect 57408 48053 71000 48359
rect 52932 48034 57097 48053
tri 57097 48034 57116 48053 sw
tri 57408 48034 57427 48053 ne
rect 57427 48034 71000 48053
rect 52932 47965 57116 48034
rect 50674 47964 52645 47965
tri 52645 47964 52646 47965 sw
tri 52932 47964 52933 47965 ne
rect 52933 47964 57116 47965
rect 50674 47956 52646 47964
rect 48471 47887 50382 47956
rect 43935 47886 48178 47887
tri 48178 47886 48179 47887 sw
tri 48471 47886 48472 47887 ne
rect 48472 47886 50382 47887
rect 39507 47773 43638 47886
rect 35022 47772 39219 47773
tri 39219 47772 39220 47773 sw
tri 39507 47772 39508 47773 ne
rect 39508 47772 43638 47773
rect 35022 47726 39220 47772
rect 30702 47657 34728 47726
tri 34728 47657 34797 47726 sw
tri 35022 47657 35091 47726 ne
rect 35091 47657 39220 47726
rect 30702 47508 34797 47657
rect 28582 47358 30412 47508
rect 26592 47079 28293 47358
rect 22180 47078 26295 47079
tri 26295 47078 26296 47079 sw
tri 26592 47078 26593 47079 ne
rect 26593 47078 28293 47079
rect 22180 46950 26296 47078
rect 17784 46820 21898 46950
rect 14000 46616 17492 46820
tri 17492 46616 17696 46820 sw
tri 17784 46616 17988 46820 ne
rect 17988 46790 21898 46820
tri 21898 46790 22058 46950 sw
tri 22180 46790 22340 46950 ne
rect 22340 46790 26296 46950
rect 17988 46626 22058 46790
tri 22058 46626 22222 46790 sw
tri 22340 46626 22504 46790 ne
rect 22504 46781 26296 46790
tri 26296 46781 26593 47078 sw
tri 26593 46781 26890 47078 ne
rect 26890 47069 28293 47078
tri 28293 47069 28582 47358 sw
tri 28582 47069 28871 47358 ne
rect 28871 47352 30412 47358
tri 30412 47352 30568 47508 sw
tri 30702 47352 30858 47508 ne
rect 30858 47363 34797 47508
tri 34797 47363 35091 47657 sw
tri 35091 47363 35385 47657 ne
rect 35385 47484 39220 47657
tri 39220 47484 39508 47772 sw
tri 39508 47484 39796 47772 ne
rect 39796 47589 43638 47772
tri 43638 47589 43935 47886 sw
tri 43935 47589 44232 47886 ne
rect 44232 47593 48179 47886
tri 48179 47593 48472 47886 sw
tri 48472 47593 48765 47886 ne
rect 48765 47816 50382 47886
tri 50382 47816 50522 47956 sw
tri 50674 47816 50814 47956 ne
rect 50814 47816 52646 47956
rect 48765 47593 50522 47816
rect 44232 47589 48472 47593
rect 39796 47588 43935 47589
tri 43935 47588 43936 47589 sw
tri 44232 47588 44233 47589 ne
rect 44233 47588 48472 47589
rect 39796 47484 43936 47588
rect 35385 47483 39508 47484
tri 39508 47483 39509 47484 sw
tri 39796 47483 39797 47484 ne
rect 39797 47483 43936 47484
rect 35385 47363 39509 47483
rect 30858 47362 35091 47363
tri 35091 47362 35092 47363 sw
tri 35385 47362 35386 47363 ne
rect 35386 47362 39509 47363
rect 30858 47352 35092 47362
rect 28871 47069 30568 47352
rect 26890 46781 28582 47069
rect 22504 46626 26593 46781
rect 17988 46616 22222 46626
rect 14000 46324 17696 46616
tri 17696 46324 17988 46616 sw
tri 17988 46324 18280 46616 ne
rect 18280 46507 22222 46616
tri 22222 46507 22341 46626 sw
tri 22504 46507 22623 46626 ne
rect 22623 46507 26593 46626
rect 18280 46324 22341 46507
rect 14000 46114 17988 46324
tri 17988 46114 18198 46324 sw
tri 18280 46114 18490 46324 ne
rect 18490 46225 22341 46324
tri 22341 46225 22623 46507 sw
tri 22623 46225 22905 46507 ne
rect 22905 46484 26593 46507
tri 26593 46484 26890 46781 sw
tri 26890 46484 27187 46781 ne
rect 27187 46780 28582 46781
tri 28582 46780 28871 47069 sw
tri 28871 46780 29160 47069 ne
rect 29160 47062 30568 47069
tri 30568 47062 30858 47352 sw
tri 30858 47062 31148 47352 ne
rect 31148 47068 35092 47352
tri 35092 47068 35386 47362 sw
tri 35386 47068 35680 47362 ne
rect 35680 47195 39509 47362
tri 39509 47195 39797 47483 sw
tri 39797 47195 40085 47483 ne
rect 40085 47291 43936 47483
tri 43936 47291 44233 47588 sw
tri 44233 47291 44530 47588 ne
rect 44530 47300 48472 47588
tri 48472 47300 48765 47593 sw
tri 48765 47300 49058 47593 ne
rect 49058 47524 50522 47593
tri 50522 47524 50814 47816 sw
tri 50814 47524 51106 47816 ne
rect 51106 47677 52646 47816
tri 52646 47677 52933 47964 sw
tri 52933 47677 53220 47964 ne
rect 53220 47728 57116 47964
tri 57116 47728 57422 48034 sw
tri 57427 47728 57733 48034 ne
rect 57733 47728 71000 48034
rect 53220 47709 57422 47728
tri 57422 47709 57441 47728 sw
tri 57733 47709 57752 47728 ne
rect 57752 47709 71000 47728
rect 53220 47677 57441 47709
rect 51106 47524 52933 47677
rect 49058 47300 50814 47524
rect 44530 47299 48765 47300
tri 48765 47299 48766 47300 sw
tri 49058 47299 49059 47300 ne
rect 49059 47299 50814 47300
rect 44530 47291 48766 47299
rect 40085 47290 44233 47291
tri 44233 47290 44234 47291 sw
tri 44530 47290 44531 47291 ne
rect 44531 47290 48766 47291
rect 40085 47195 44234 47290
rect 35680 47068 39797 47195
rect 31148 47067 35386 47068
tri 35386 47067 35387 47068 sw
tri 35680 47067 35681 47068 ne
rect 35681 47067 39797 47068
rect 31148 47062 35387 47067
rect 29160 47061 30858 47062
tri 30858 47061 30859 47062 sw
tri 31148 47061 31149 47062 ne
rect 31149 47061 35387 47062
rect 29160 46780 30859 47061
rect 27187 46491 28871 46780
tri 28871 46491 29160 46780 sw
tri 29160 46491 29449 46780 ne
rect 29449 46771 30859 46780
tri 30859 46771 31149 47061 sw
tri 31149 46771 31439 47061 ne
rect 31439 46773 35387 47061
tri 35387 46773 35681 47067 sw
tri 35681 46773 35975 47067 ne
rect 35975 46976 39797 47067
tri 39797 46976 40016 47195 sw
tri 40085 46976 40304 47195 ne
rect 40304 46993 44234 47195
tri 44234 46993 44531 47290 sw
tri 44531 46993 44828 47290 ne
rect 44828 47006 48766 47290
tri 48766 47006 49059 47299 sw
tri 49059 47006 49352 47299 ne
rect 49352 47232 50814 47299
tri 50814 47232 51106 47524 sw
tri 51106 47232 51398 47524 ne
rect 51398 47422 52933 47524
tri 52933 47422 53188 47677 sw
tri 53220 47422 53475 47677 ne
rect 53475 47422 57441 47677
rect 51398 47232 53188 47422
rect 49352 47006 51106 47232
rect 44828 46993 49059 47006
rect 40304 46992 44531 46993
tri 44531 46992 44532 46993 sw
tri 44828 46992 44829 46993 ne
rect 44829 46992 49059 46993
rect 40304 46976 44532 46992
rect 35975 46773 40016 46976
rect 31439 46771 35681 46773
rect 29449 46690 31149 46771
tri 31149 46690 31230 46771 sw
tri 31439 46690 31520 46771 ne
rect 31520 46690 35681 46771
rect 29449 46491 31230 46690
rect 27187 46484 29160 46491
rect 22905 46483 26890 46484
tri 26890 46483 26891 46484 sw
tri 27187 46483 27188 46484 ne
rect 27188 46483 29160 46484
rect 22905 46225 26891 46483
rect 18490 46224 22623 46225
tri 22623 46224 22624 46225 sw
tri 22905 46224 22906 46225 ne
rect 22906 46224 26891 46225
rect 18490 46114 22624 46224
rect 14000 46068 18198 46114
tri 14000 43708 16360 46068 ne
rect 16360 45822 18198 46068
tri 18198 45822 18490 46114 sw
tri 18490 45822 18782 46114 ne
rect 18782 45942 22624 46114
tri 22624 45942 22906 46224 sw
tri 22906 45942 23188 46224 ne
rect 23188 46186 26891 46224
tri 26891 46186 27188 46483 sw
tri 27188 46186 27485 46483 ne
rect 27485 46400 29160 46483
tri 29160 46400 29251 46491 sw
tri 29449 46400 29540 46491 ne
rect 29540 46400 31230 46491
tri 31230 46400 31520 46690 sw
tri 31520 46400 31810 46690 ne
rect 31810 46682 35681 46690
tri 35681 46682 35772 46773 sw
tri 35975 46682 36066 46773 ne
rect 36066 46688 40016 46773
tri 40016 46688 40304 46976 sw
tri 40304 46688 40592 46976 ne
rect 40592 46695 44532 46976
tri 44532 46695 44829 46992 sw
tri 44829 46695 45126 46992 ne
rect 45126 46940 49059 46992
tri 49059 46940 49125 47006 sw
tri 49352 46940 49418 47006 ne
rect 49418 46940 51106 47006
tri 51106 46940 51398 47232 sw
tri 51398 46940 51690 47232 ne
rect 51690 47135 53188 47232
tri 53188 47135 53475 47422 sw
tri 53475 47135 53762 47422 ne
rect 53762 47402 57441 47422
tri 57441 47402 57748 47709 sw
tri 57752 47402 58059 47709 ne
rect 58059 47402 71000 47709
rect 53762 47135 57748 47402
rect 51690 47053 53475 47135
tri 53475 47053 53557 47135 sw
tri 53762 47053 53844 47135 ne
rect 53844 47110 57748 47135
tri 57748 47110 58040 47402 sw
tri 58059 47110 58351 47402 ne
rect 58351 47110 71000 47402
rect 53844 47053 58040 47110
tri 58040 47053 58097 47110 sw
tri 58351 47053 58408 47110 ne
rect 58408 47053 71000 47110
rect 51690 46940 53557 47053
rect 45126 46695 49125 46940
rect 40592 46693 44829 46695
tri 44829 46693 44831 46695 sw
tri 45126 46693 45128 46695 ne
rect 45128 46693 49125 46695
rect 40592 46688 44831 46693
rect 36066 46682 40304 46688
rect 31810 46400 35772 46682
rect 27485 46186 29251 46400
rect 23188 46185 27188 46186
tri 27188 46185 27189 46186 sw
tri 27485 46185 27486 46186 ne
rect 27486 46185 29251 46186
rect 23188 45942 27189 46185
rect 18782 45941 22906 45942
tri 22906 45941 22907 45942 sw
tri 23188 45941 23189 45942 ne
rect 23189 45941 27189 45942
rect 18782 45822 22907 45941
rect 16360 45821 18490 45822
tri 18490 45821 18491 45822 sw
tri 18782 45821 18783 45822 ne
rect 18783 45821 22907 45822
rect 16360 45529 18491 45821
tri 18491 45529 18783 45821 sw
tri 18783 45529 19075 45821 ne
rect 19075 45659 22907 45821
tri 22907 45659 23189 45941 sw
tri 23189 45659 23471 45941 ne
rect 23471 45888 27189 45941
tri 27189 45888 27486 46185 sw
tri 27486 45888 27783 46185 ne
rect 27783 46111 29251 46185
tri 29251 46111 29540 46400 sw
tri 29540 46111 29829 46400 ne
rect 29829 46399 31520 46400
tri 31520 46399 31521 46400 sw
tri 31810 46399 31811 46400 ne
rect 31811 46399 35772 46400
rect 29829 46111 31521 46399
rect 27783 45888 29540 46111
rect 23471 45804 27486 45888
tri 27486 45804 27570 45888 sw
tri 27783 45804 27867 45888 ne
rect 27867 45822 29540 45888
tri 29540 45822 29829 46111 sw
tri 29829 45822 30118 46111 ne
rect 30118 46109 31521 46111
tri 31521 46109 31811 46399 sw
tri 31811 46109 32101 46399 ne
rect 32101 46388 35772 46399
tri 35772 46388 36066 46682 sw
tri 36066 46388 36360 46682 ne
rect 36360 46597 40304 46682
tri 40304 46597 40395 46688 sw
tri 40592 46597 40683 46688 ne
rect 40683 46597 44831 46688
rect 36360 46388 40395 46597
rect 32101 46181 36066 46388
tri 36066 46181 36273 46388 sw
tri 36360 46181 36567 46388 ne
rect 36567 46309 40395 46388
tri 40395 46309 40683 46597 sw
tri 40683 46309 40971 46597 ne
rect 40971 46396 44831 46597
tri 44831 46396 45128 46693 sw
tri 45128 46396 45425 46693 ne
rect 45425 46647 49125 46693
tri 49125 46647 49418 46940 sw
tri 49418 46647 49711 46940 ne
rect 49711 46648 51398 46940
tri 51398 46648 51690 46940 sw
tri 51690 46648 51982 46940 ne
rect 51982 46766 53557 46940
tri 53557 46766 53844 47053 sw
tri 53844 46766 54131 47053 ne
rect 54131 46766 58097 47053
rect 51982 46648 53844 46766
rect 49711 46647 51690 46648
rect 45425 46396 49418 46647
rect 40971 46309 45128 46396
rect 36567 46307 40683 46309
tri 40683 46307 40685 46309 sw
tri 40971 46307 40973 46309 ne
rect 40973 46307 45128 46309
rect 36567 46181 40685 46307
rect 32101 46109 36273 46181
rect 30118 45822 31811 46109
rect 27867 45804 29829 45822
rect 23471 45659 27570 45804
rect 19075 45582 23189 45659
tri 23189 45582 23266 45659 sw
tri 23471 45582 23548 45659 ne
rect 23548 45582 27570 45659
rect 19075 45529 23266 45582
rect 16360 45527 18783 45529
tri 18783 45527 18785 45529 sw
tri 19075 45527 19077 45529 ne
rect 19077 45527 23266 45529
rect 16360 45236 18785 45527
tri 18785 45236 19076 45527 sw
tri 19077 45236 19368 45527 ne
rect 19368 45300 23266 45527
tri 23266 45300 23548 45582 sw
tri 23548 45300 23830 45582 ne
rect 23830 45507 27570 45582
tri 27570 45507 27867 45804 sw
tri 27867 45507 28164 45804 ne
rect 28164 45667 29829 45804
tri 29829 45667 29984 45822 sw
tri 30118 45667 30273 45822 ne
rect 30273 45819 31811 45822
tri 31811 45819 32101 46109 sw
tri 32101 45819 32391 46109 ne
rect 32391 45887 36273 46109
tri 36273 45887 36567 46181 sw
tri 36567 45887 36861 46181 ne
rect 36861 46019 40685 46181
tri 40685 46019 40973 46307 sw
tri 40973 46019 41261 46307 ne
rect 41261 46099 45128 46307
tri 45128 46099 45425 46396 sw
tri 45425 46099 45722 46396 ne
rect 45722 46354 49418 46396
tri 49418 46354 49711 46647 sw
tri 49711 46354 50004 46647 ne
rect 50004 46560 51690 46647
tri 51690 46560 51778 46648 sw
tri 51982 46560 52070 46648 ne
rect 52070 46560 53844 46648
rect 50004 46354 51778 46560
rect 45722 46353 49711 46354
tri 49711 46353 49712 46354 sw
tri 50004 46353 50005 46354 ne
rect 50005 46353 51778 46354
rect 45722 46099 49712 46353
rect 41261 46019 45425 46099
rect 36861 46018 40973 46019
tri 40973 46018 40974 46019 sw
tri 41261 46018 41262 46019 ne
rect 41262 46018 45425 46019
rect 36861 45887 40974 46018
rect 32391 45819 36567 45887
rect 30273 45818 32101 45819
tri 32101 45818 32102 45819 sw
tri 32391 45818 32392 45819 ne
rect 32392 45818 36567 45819
rect 30273 45667 32102 45818
rect 28164 45507 29984 45667
rect 23830 45300 27867 45507
rect 19368 45236 23548 45300
rect 16360 44992 19076 45236
tri 19076 44992 19320 45236 sw
tri 19368 44992 19612 45236 ne
rect 19612 45091 23548 45236
tri 23548 45091 23757 45300 sw
tri 23830 45091 24039 45300 ne
rect 24039 45210 27867 45300
tri 27867 45210 28164 45507 sw
tri 28164 45210 28461 45507 ne
rect 28461 45378 29984 45507
tri 29984 45378 30273 45667 sw
tri 30273 45378 30562 45667 ne
rect 30562 45528 32102 45667
tri 32102 45528 32392 45818 sw
tri 32392 45528 32682 45818 ne
rect 32682 45729 36567 45818
tri 36567 45729 36725 45887 sw
tri 36861 45729 37019 45887 ne
rect 37019 45730 40974 45887
tri 40974 45730 41262 46018 sw
tri 41262 45730 41550 46018 ne
rect 41550 45879 45425 46018
tri 45425 45879 45645 46099 sw
tri 45722 45879 45942 46099 ne
rect 45942 46060 49712 46099
tri 49712 46060 50005 46353 sw
tri 50005 46060 50298 46353 ne
rect 50298 46268 51778 46353
tri 51778 46268 52070 46560 sw
tri 52070 46268 52362 46560 ne
rect 52362 46559 53844 46560
tri 53844 46559 54051 46766 sw
tri 54131 46559 54338 46766 ne
rect 54338 46742 58097 46766
tri 58097 46742 58408 47053 sw
tri 58408 46742 58719 47053 ne
rect 58719 46742 71000 47053
rect 54338 46559 58408 46742
rect 52362 46272 54051 46559
tri 54051 46272 54338 46559 sw
tri 54338 46272 54625 46559 ne
rect 54625 46460 58408 46559
tri 58408 46460 58690 46742 sw
tri 58719 46460 59001 46742 ne
rect 59001 46460 71000 46742
rect 54625 46272 58690 46460
rect 52362 46268 54338 46272
rect 50298 46060 52070 46268
rect 45942 45879 50005 46060
rect 41550 45730 45645 45879
rect 37019 45729 41262 45730
rect 32682 45528 36725 45729
rect 30562 45378 32392 45528
rect 28461 45210 30273 45378
rect 24039 45091 28164 45210
rect 19612 44992 23757 45091
rect 16360 44700 19320 44992
tri 19320 44700 19612 44992 sw
tri 19612 44700 19904 44992 ne
rect 19904 44809 23757 44992
tri 23757 44809 24039 45091 sw
tri 24039 44809 24321 45091 ne
rect 24321 44913 28164 45091
tri 28164 44913 28461 45210 sw
tri 28461 44913 28758 45210 ne
rect 28758 45089 30273 45210
tri 30273 45089 30562 45378 sw
tri 30562 45089 30851 45378 ne
rect 30851 45291 32392 45378
tri 32392 45291 32629 45528 sw
tri 32682 45291 32919 45528 ne
rect 32919 45435 36725 45528
tri 36725 45435 37019 45729 sw
tri 37019 45435 37313 45729 ne
rect 37313 45644 41262 45729
tri 41262 45644 41348 45730 sw
tri 41550 45644 41636 45730 ne
rect 41636 45644 45645 45730
rect 37313 45435 41348 45644
rect 32919 45434 37019 45435
tri 37019 45434 37020 45435 sw
tri 37313 45434 37314 45435 ne
rect 37314 45434 41348 45435
rect 32919 45291 37020 45434
rect 30851 45089 32629 45291
rect 28758 44913 30562 45089
rect 24321 44912 28461 44913
tri 28461 44912 28462 44913 sw
tri 28758 44912 28759 44913 ne
rect 28759 44912 30562 44913
rect 24321 44809 28462 44912
rect 19904 44700 24039 44809
rect 16360 44698 19612 44700
tri 19612 44698 19614 44700 sw
tri 19904 44698 19906 44700 ne
rect 19906 44698 24039 44700
rect 16360 44406 19614 44698
tri 19614 44406 19906 44698 sw
tri 19906 44406 20198 44698 ne
rect 20198 44615 24039 44698
tri 24039 44615 24233 44809 sw
tri 24321 44615 24515 44809 ne
rect 24515 44615 28462 44809
tri 28462 44615 28759 44912 sw
tri 28759 44615 29056 44912 ne
rect 29056 44800 30562 44912
tri 30562 44800 30851 45089 sw
tri 30851 44800 31140 45089 ne
rect 31140 45001 32629 45089
tri 32629 45001 32919 45291 sw
tri 32919 45001 33209 45291 ne
rect 33209 45140 37020 45291
tri 37020 45140 37314 45434 sw
tri 37314 45140 37608 45434 ne
rect 37608 45356 41348 45434
tri 41348 45356 41636 45644 sw
tri 41636 45356 41924 45644 ne
rect 41924 45635 45645 45644
tri 45645 45635 45889 45879 sw
tri 45942 45635 46186 45879 ne
rect 46186 45767 50005 45879
tri 50005 45767 50298 46060 sw
tri 50298 45767 50591 46060 ne
rect 50591 45976 52070 46060
tri 52070 45976 52362 46268 sw
tri 52362 45976 52654 46268 ne
rect 52654 46087 54338 46268
tri 54338 46087 54523 46272 sw
tri 54625 46087 54810 46272 ne
rect 54810 46154 58690 46272
tri 58690 46154 58996 46460 sw
tri 59001 46154 59307 46460 ne
rect 59307 46154 71000 46460
rect 54810 46135 58996 46154
tri 58996 46135 59015 46154 sw
tri 59307 46135 59326 46154 ne
rect 59326 46135 71000 46154
rect 54810 46087 59015 46135
rect 52654 45976 54523 46087
rect 50591 45836 52362 45976
tri 52362 45836 52502 45976 sw
tri 52654 45836 52794 45976 ne
rect 52794 45836 54523 45976
rect 50591 45767 52502 45836
rect 46186 45635 50298 45767
rect 41924 45581 45889 45635
tri 45889 45581 45943 45635 sw
tri 46186 45581 46240 45635 ne
rect 46240 45581 50298 45635
rect 41924 45356 45943 45581
rect 37608 45151 41636 45356
tri 41636 45151 41841 45356 sw
tri 41924 45151 42129 45356 ne
rect 42129 45284 45943 45356
tri 45943 45284 46240 45581 sw
tri 46240 45284 46537 45581 ne
rect 46537 45548 50298 45581
tri 50298 45548 50517 45767 sw
tri 50591 45548 50810 45767 ne
rect 50810 45548 52502 45767
rect 46537 45284 50517 45548
rect 42129 45283 46240 45284
tri 46240 45283 46241 45284 sw
tri 46537 45283 46538 45284 ne
rect 46538 45283 50517 45284
rect 42129 45151 46241 45283
rect 37608 45140 41841 45151
rect 33209 45139 37314 45140
tri 37314 45139 37315 45140 sw
tri 37608 45139 37609 45140 ne
rect 37609 45139 41841 45140
rect 33209 45001 37315 45139
rect 31140 44800 32919 45001
rect 29056 44615 30851 44800
rect 20198 44406 24233 44615
rect 16360 44405 19906 44406
tri 19906 44405 19907 44406 sw
tri 20198 44405 20199 44406 ne
rect 20199 44405 24233 44406
rect 16360 44113 19907 44405
tri 19907 44113 20199 44405 sw
tri 20199 44113 20491 44405 ne
rect 20491 44333 24233 44405
tri 24233 44333 24515 44615 sw
tri 24515 44333 24797 44615 ne
rect 24797 44333 28759 44615
rect 20491 44331 24515 44333
tri 24515 44331 24517 44333 sw
tri 24797 44331 24799 44333 ne
rect 24799 44331 28759 44333
rect 20491 44113 24517 44331
rect 16360 44112 20199 44113
tri 20199 44112 20200 44113 sw
tri 20491 44112 20492 44113 ne
rect 20492 44112 24517 44113
rect 16360 43820 20200 44112
tri 20200 43820 20492 44112 sw
tri 20492 43820 20784 44112 ne
rect 20784 44049 24517 44112
tri 24517 44049 24799 44331 sw
tri 24799 44049 25081 44331 ne
rect 25081 44318 28759 44331
tri 28759 44318 29056 44615 sw
tri 29056 44318 29353 44615 ne
rect 29353 44511 30851 44615
tri 30851 44511 31140 44800 sw
tri 31140 44511 31429 44800 ne
rect 31429 44711 32919 44800
tri 32919 44711 33209 45001 sw
tri 33209 44711 33499 45001 ne
rect 33499 44845 37315 45001
tri 37315 44845 37609 45139 sw
tri 37609 44845 37903 45139 ne
rect 37903 44863 41841 45139
tri 41841 44863 42129 45151 sw
tri 42129 44863 42417 45151 ne
rect 42417 44986 46241 45151
tri 46241 44986 46538 45283 sw
tri 46538 44986 46835 45283 ne
rect 46835 45255 50517 45283
tri 50517 45255 50810 45548 sw
tri 50810 45255 51103 45548 ne
rect 51103 45544 52502 45548
tri 52502 45544 52794 45836 sw
tri 52794 45544 53086 45836 ne
rect 53086 45800 54523 45836
tri 54523 45800 54810 46087 sw
tri 54810 45800 55097 46087 ne
rect 55097 45829 59015 46087
tri 59015 45829 59321 46135 sw
tri 59326 46000 59461 46135 ne
rect 59461 46000 71000 46135
rect 55097 45800 59321 45829
tri 59321 45800 59350 45829 sw
rect 53086 45799 54810 45800
tri 54810 45799 54811 45800 sw
tri 55097 45799 55098 45800 ne
rect 55098 45799 71000 45800
rect 53086 45544 54811 45799
rect 51103 45255 52794 45544
rect 46835 45254 50810 45255
tri 50810 45254 50811 45255 sw
tri 51103 45254 51104 45255 ne
rect 51104 45254 52794 45255
rect 46835 44986 50811 45254
rect 42417 44984 46538 44986
tri 46538 44984 46540 44986 sw
tri 46835 44984 46837 44986 ne
rect 46837 44984 50811 44986
rect 42417 44863 46540 44984
rect 37903 44845 42129 44863
rect 33499 44843 37609 44845
tri 37609 44843 37611 44845 sw
tri 37903 44843 37905 44845 ne
rect 37905 44843 42129 44845
rect 33499 44711 37611 44843
rect 31429 44710 33209 44711
tri 33209 44710 33210 44711 sw
tri 33499 44710 33500 44711 ne
rect 33500 44710 37611 44711
rect 31429 44511 33210 44710
rect 29353 44420 31140 44511
tri 31140 44420 31231 44511 sw
tri 31429 44420 31520 44511 ne
rect 31520 44420 33210 44511
tri 33210 44420 33500 44710 sw
tri 33500 44420 33790 44710 ne
rect 33790 44549 37611 44710
tri 37611 44549 37905 44843 sw
tri 37905 44549 38199 44843 ne
rect 38199 44686 42129 44843
tri 42129 44686 42306 44863 sw
tri 42417 44686 42594 44863 ne
rect 42594 44688 46540 44863
tri 46540 44688 46836 44984 sw
tri 46837 44688 47133 44984 ne
rect 47133 44961 50811 44984
tri 50811 44961 51104 45254 sw
tri 51104 44961 51397 45254 ne
rect 51397 45252 52794 45254
tri 52794 45252 53086 45544 sw
tri 53086 45252 53378 45544 ne
rect 53378 45512 54811 45544
tri 54811 45512 55098 45799 sw
tri 55098 45512 55385 45799 ne
rect 55385 45512 71000 45799
rect 53378 45252 55098 45512
rect 51397 44961 53086 45252
rect 47133 44688 51104 44961
rect 42594 44686 46836 44688
rect 38199 44549 42306 44686
rect 33790 44548 37905 44549
tri 37905 44548 37906 44549 sw
tri 38199 44548 38200 44549 ne
rect 38200 44548 42306 44549
rect 33790 44420 37906 44548
rect 29353 44318 31231 44420
rect 25081 44317 29056 44318
tri 29056 44317 29057 44318 sw
tri 29353 44317 29354 44318 ne
rect 29354 44317 31231 44318
rect 25081 44049 29057 44317
rect 20784 44048 24799 44049
tri 24799 44048 24800 44049 sw
tri 25081 44048 25082 44049 ne
rect 25082 44048 29057 44049
rect 20784 43820 24800 44048
rect 16360 43708 20492 43820
tri 20492 43708 20604 43820 sw
tri 20784 43708 20896 43820 ne
rect 20896 43766 24800 43820
tri 24800 43766 25082 44048 sw
tri 25082 43766 25364 44048 ne
rect 25364 44020 29057 44048
tri 29057 44020 29354 44317 sw
tri 29354 44020 29651 44317 ne
rect 29651 44131 31231 44317
tri 31231 44131 31520 44420 sw
tri 31520 44131 31809 44420 ne
rect 31809 44419 33500 44420
tri 33500 44419 33501 44420 sw
tri 33790 44419 33791 44420 ne
rect 33791 44419 37906 44420
rect 31809 44131 33501 44419
rect 29651 44020 31520 44131
rect 25364 44019 29354 44020
tri 29354 44019 29355 44020 sw
tri 29651 44019 29652 44020 ne
rect 29652 44019 31520 44020
rect 25364 43766 29355 44019
rect 20896 43765 25082 43766
tri 25082 43765 25083 43766 sw
tri 25364 43765 25365 43766 ne
rect 25365 43765 29355 43766
rect 20896 43708 25083 43765
tri 16360 39464 20604 43708 ne
tri 20604 43416 20896 43708 sw
tri 20896 43416 21188 43708 ne
rect 21188 43483 25083 43708
tri 25083 43483 25365 43765 sw
tri 25365 43483 25647 43765 ne
rect 25647 43722 29355 43765
tri 29355 43722 29652 44019 sw
tri 29652 43722 29949 44019 ne
rect 29949 43842 31520 44019
tri 31520 43842 31809 44131 sw
tri 31809 43842 32098 44131 ne
rect 32098 44129 33501 44131
tri 33501 44129 33791 44419 sw
tri 33791 44129 34081 44419 ne
rect 34081 44254 37906 44419
tri 37906 44254 38200 44548 sw
tri 38200 44254 38494 44548 ne
rect 38494 44398 42306 44548
tri 42306 44398 42594 44686 sw
tri 42594 44398 42882 44686 ne
rect 42882 44591 46836 44686
tri 46836 44591 46933 44688 sw
tri 47133 44591 47230 44688 ne
rect 47230 44668 51104 44688
tri 51104 44668 51397 44961 sw
tri 51397 44668 51690 44961 ne
rect 51690 44960 53086 44961
tri 53086 44960 53378 45252 sw
tri 53378 44960 53670 45252 ne
rect 53670 45225 55098 45252
tri 55098 45225 55385 45512 sw
tri 55385 45225 55672 45512 ne
rect 55672 45225 71000 45512
rect 53670 45155 55385 45225
tri 55385 45155 55455 45225 sw
tri 55672 45155 55742 45225 ne
rect 55742 45155 71000 45225
rect 53670 44960 55455 45155
rect 51690 44668 53378 44960
tri 53378 44668 53670 44960 sw
tri 53670 44668 53962 44960 ne
rect 53962 44868 55455 44960
tri 55455 44868 55742 45155 sw
tri 55742 44868 56029 45155 ne
rect 56029 44868 71000 45155
rect 53962 44867 55742 44868
tri 55742 44867 55743 44868 sw
tri 56029 44867 56030 44868 ne
rect 56030 44867 71000 44868
rect 53962 44668 55743 44867
rect 47230 44666 51397 44668
tri 51397 44666 51399 44668 sw
tri 51690 44666 51692 44668 ne
rect 51692 44666 53670 44668
rect 47230 44591 51399 44666
rect 42882 44398 46933 44591
rect 38494 44397 42594 44398
tri 42594 44397 42595 44398 sw
tri 42882 44397 42883 44398 ne
rect 42883 44397 46933 44398
rect 38494 44254 42595 44397
rect 34081 44253 38200 44254
tri 38200 44253 38201 44254 sw
tri 38494 44253 38495 44254 ne
rect 38495 44253 42595 44254
rect 34081 44129 38201 44253
rect 32098 43842 33791 44129
rect 29949 43722 31809 43842
rect 25647 43483 29652 43722
rect 21188 43482 25365 43483
tri 25365 43482 25366 43483 sw
tri 25647 43482 25648 43483 ne
rect 25648 43482 29652 43483
rect 21188 43416 25366 43482
rect 20604 43233 20896 43416
tri 20896 43233 21079 43416 sw
tri 21188 43233 21371 43416 ne
rect 21371 43233 25366 43416
rect 20604 43044 21079 43233
tri 21079 43044 21268 43233 sw
tri 21371 43044 21560 43233 ne
rect 21560 43200 25366 43233
tri 25366 43200 25648 43482 sw
tri 25648 43200 25930 43482 ne
rect 25930 43425 29652 43482
tri 29652 43425 29949 43722 sw
tri 29949 43425 30246 43722 ne
rect 30246 43687 31809 43722
tri 31809 43687 31964 43842 sw
tri 32098 43687 32253 43842 ne
rect 32253 43839 33791 43842
tri 33791 43839 34081 44129 sw
tri 34081 43839 34371 44129 ne
rect 34371 43959 38201 44129
tri 38201 43959 38495 44253 sw
tri 38495 43959 38789 44253 ne
rect 38789 44109 42595 44253
tri 42595 44109 42883 44397 sw
tri 42883 44109 43171 44397 ne
rect 43171 44294 46933 44397
tri 46933 44294 47230 44591 sw
tri 47230 44294 47527 44591 ne
rect 47527 44373 51399 44591
tri 51399 44373 51692 44666 sw
tri 51692 44373 51985 44666 ne
rect 51985 44580 53670 44666
tri 53670 44580 53758 44668 sw
tri 53962 44580 54050 44668 ne
rect 54050 44580 55743 44668
tri 55743 44580 56030 44867 sw
tri 56030 44580 56317 44867 ne
rect 56317 44580 71000 44867
rect 51985 44373 53758 44580
rect 47527 44294 51692 44373
rect 43171 44109 47230 44294
rect 38789 44108 42883 44109
tri 42883 44108 42884 44109 sw
tri 43171 44108 43172 44109 ne
rect 43172 44108 47230 44109
rect 38789 43959 42884 44108
rect 34371 43839 38495 43959
rect 32253 43776 34081 43839
tri 34081 43776 34144 43839 sw
tri 34371 43776 34434 43839 ne
rect 34434 43776 38495 43839
rect 32253 43687 34144 43776
rect 30246 43425 31964 43687
rect 25930 43416 29949 43425
tri 29949 43416 29958 43425 sw
tri 30246 43416 30255 43425 ne
rect 30255 43416 31964 43425
rect 25930 43200 29958 43416
rect 21560 43199 25648 43200
tri 25648 43199 25649 43200 sw
tri 25930 43199 25931 43200 ne
rect 25931 43199 29958 43200
rect 21560 43044 25649 43199
rect 20604 42752 21268 43044
tri 21268 42752 21560 43044 sw
tri 21560 42752 21852 43044 ne
rect 21852 42917 25649 43044
tri 25649 42917 25931 43199 sw
tri 25931 42917 26213 43199 ne
rect 26213 43119 29958 43199
tri 29958 43119 30255 43416 sw
tri 30255 43119 30552 43416 ne
rect 30552 43398 31964 43416
tri 31964 43398 32253 43687 sw
tri 32253 43398 32542 43687 ne
rect 32542 43486 34144 43687
tri 34144 43486 34434 43776 sw
tri 34434 43486 34724 43776 ne
rect 34724 43710 38495 43776
tri 38495 43710 38744 43959 sw
tri 38789 43710 39038 43959 ne
rect 39038 43820 42884 43959
tri 42884 43820 43172 44108 sw
tri 43172 43820 43460 44108 ne
rect 43460 44090 47230 44108
tri 47230 44090 47434 44294 sw
tri 47527 44090 47731 44294 ne
rect 47731 44090 51692 44294
rect 43460 43820 47434 44090
rect 39038 43819 43172 43820
tri 43172 43819 43173 43820 sw
tri 43460 43819 43461 43820 ne
rect 43461 43819 47434 43820
rect 39038 43710 43173 43819
rect 34724 43486 38744 43710
rect 32542 43398 34434 43486
rect 30552 43119 32253 43398
rect 26213 43118 30255 43119
tri 30255 43118 30256 43119 sw
tri 30552 43118 30553 43119 ne
rect 30553 43118 32253 43119
rect 26213 42917 30256 43118
rect 21852 42752 25931 42917
rect 20604 42751 21560 42752
tri 21560 42751 21561 42752 sw
tri 21852 42751 21853 42752 ne
rect 21853 42751 25931 42752
rect 20604 42459 21561 42751
tri 21561 42459 21853 42751 sw
tri 21853 42459 22145 42751 ne
rect 22145 42664 25931 42751
tri 25931 42664 26184 42917 sw
tri 26213 42664 26466 42917 ne
rect 26466 42821 30256 42917
tri 30256 42821 30553 43118 sw
tri 30553 42821 30850 43118 ne
rect 30850 43109 32253 43118
tri 32253 43109 32542 43398 sw
tri 32542 43109 32831 43398 ne
rect 32831 43311 34434 43398
tri 34434 43311 34609 43486 sw
tri 34724 43311 34899 43486 ne
rect 34899 43482 38744 43486
tri 38744 43482 38972 43710 sw
tri 39038 43482 39266 43710 ne
rect 39266 43531 43173 43710
tri 43173 43531 43461 43819 sw
tri 43461 43531 43749 43819 ne
rect 43749 43793 47434 43819
tri 47434 43793 47731 44090 sw
tri 47731 43793 48028 44090 ne
rect 48028 44080 51692 44090
tri 51692 44080 51985 44373 sw
tri 51985 44080 52278 44373 ne
rect 52278 44288 53758 44373
tri 53758 44288 54050 44580 sw
tri 54050 44288 54342 44580 ne
rect 54342 44579 56030 44580
tri 56030 44579 56031 44580 sw
tri 56317 44579 56318 44580 ne
rect 56318 44579 71000 44580
rect 54342 44292 56031 44579
tri 56031 44292 56318 44579 sw
tri 56318 44292 56605 44579 ne
rect 56605 44292 71000 44579
rect 54342 44288 56318 44292
rect 52278 44080 54050 44288
rect 48028 43937 51985 44080
tri 51985 43937 52128 44080 sw
tri 52278 43937 52421 44080 ne
rect 52421 43996 54050 44080
tri 54050 43996 54342 44288 sw
tri 54342 43996 54634 44288 ne
rect 54634 44005 56318 44288
tri 56318 44005 56605 44292 sw
tri 56605 44005 56892 44292 ne
rect 56892 44005 71000 44292
rect 54634 44004 56605 44005
tri 56605 44004 56606 44005 sw
tri 56892 44004 56893 44005 ne
rect 56893 44004 71000 44005
rect 54634 43996 56606 44004
rect 52421 43937 54342 43996
rect 48028 43793 52128 43937
rect 43749 43643 47731 43793
tri 47731 43643 47881 43793 sw
tri 48028 43643 48178 43793 ne
rect 48178 43644 52128 43793
tri 52128 43644 52421 43937 sw
tri 52421 43644 52714 43937 ne
rect 52714 43856 54342 43937
tri 54342 43856 54482 43996 sw
tri 54634 43856 54774 43996 ne
rect 54774 43856 56606 43996
rect 52714 43644 54482 43856
rect 48178 43643 52421 43644
tri 52421 43643 52422 43644 sw
tri 52714 43643 52715 43644 ne
rect 52715 43643 54482 43644
rect 43749 43531 47881 43643
rect 39266 43529 43461 43531
tri 43461 43529 43463 43531 sw
tri 43749 43529 43751 43531 ne
rect 43751 43529 47881 43531
rect 39266 43482 43463 43529
rect 34899 43415 38972 43482
tri 38972 43415 39039 43482 sw
tri 39266 43415 39333 43482 ne
rect 39333 43415 43463 43482
rect 34899 43311 39039 43415
rect 32831 43109 34609 43311
rect 30850 42821 32542 43109
rect 26466 42664 30553 42821
rect 22145 42459 26184 42664
rect 20604 42372 21853 42459
tri 21853 42372 21940 42459 sw
tri 22145 42372 22232 42459 ne
rect 22232 42382 26184 42459
tri 26184 42382 26466 42664 sw
tri 26466 42382 26748 42664 ne
rect 26748 42524 30553 42664
tri 30553 42524 30850 42821 sw
tri 30850 42524 31147 42821 ne
rect 31147 42820 32542 42821
tri 32542 42820 32831 43109 sw
tri 32831 42820 33120 43109 ne
rect 33120 43021 34609 43109
tri 34609 43021 34899 43311 sw
tri 34899 43021 35189 43311 ne
rect 35189 43121 39039 43311
tri 39039 43121 39333 43415 sw
tri 39333 43121 39627 43415 ne
rect 39627 43241 43463 43415
tri 43463 43241 43751 43529 sw
tri 43751 43241 44039 43529 ne
rect 44039 43346 47881 43529
tri 47881 43346 48178 43643 sw
tri 48178 43346 48475 43643 ne
rect 48475 43350 52422 43643
tri 52422 43350 52715 43643 sw
tri 52715 43350 53008 43643 ne
rect 53008 43564 54482 43643
tri 54482 43564 54774 43856 sw
tri 54774 43564 55066 43856 ne
rect 55066 43717 56606 43856
tri 56606 43717 56893 44004 sw
tri 56893 43717 57180 44004 ne
rect 57180 43717 71000 44004
rect 55066 43564 56893 43717
rect 53008 43350 54774 43564
rect 48475 43346 52715 43350
rect 44039 43345 48178 43346
tri 48178 43345 48179 43346 sw
tri 48475 43345 48476 43346 ne
rect 48476 43345 52715 43346
rect 44039 43241 48179 43345
rect 39627 43121 43751 43241
rect 35189 43119 39333 43121
tri 39333 43119 39335 43121 sw
tri 39627 43119 39629 43121 ne
rect 39629 43119 43751 43121
rect 35189 43021 39335 43119
rect 33120 42820 34899 43021
rect 31147 42531 32831 42820
tri 32831 42531 33120 42820 sw
tri 33120 42531 33409 42820 ne
rect 33409 42731 34899 42820
tri 34899 42731 35189 43021 sw
tri 35189 42731 35479 43021 ne
rect 35479 42825 39335 43021
tri 39335 42825 39629 43119 sw
tri 39629 42825 39923 43119 ne
rect 39923 42953 43751 43119
tri 43751 42953 44039 43241 sw
tri 44039 42953 44327 43241 ne
rect 44327 43048 48179 43241
tri 48179 43048 48476 43345 sw
tri 48476 43048 48773 43345 ne
rect 48773 43057 52715 43345
tri 52715 43057 53008 43350 sw
tri 53008 43057 53301 43350 ne
rect 53301 43272 54774 43350
tri 54774 43272 55066 43564 sw
tri 55066 43272 55358 43564 ne
rect 55358 43462 56893 43564
tri 56893 43462 57148 43717 sw
tri 57180 43462 57435 43717 ne
rect 57435 43462 71000 43717
rect 55358 43272 57148 43462
rect 53301 43057 55066 43272
rect 48773 43048 53008 43057
rect 44327 43047 48476 43048
tri 48476 43047 48477 43048 sw
tri 48773 43047 48774 43048 ne
rect 48774 43047 53008 43048
rect 44327 42953 48477 43047
rect 39923 42825 44039 42953
rect 35479 42824 39629 42825
tri 39629 42824 39630 42825 sw
tri 39923 42824 39924 42825 ne
rect 39924 42824 44039 42825
rect 35479 42731 39630 42824
rect 33409 42730 35189 42731
tri 35189 42730 35190 42731 sw
tri 35479 42730 35480 42731 ne
rect 35480 42730 39630 42731
rect 33409 42531 35190 42730
rect 31147 42524 33120 42531
rect 26748 42523 30850 42524
tri 30850 42523 30851 42524 sw
tri 31147 42523 31148 42524 ne
rect 31148 42523 33120 42524
rect 26748 42382 30851 42523
rect 22232 42372 26466 42382
rect 20604 42080 21940 42372
tri 21940 42080 22232 42372 sw
tri 22232 42080 22524 42372 ne
rect 22524 42264 26466 42372
tri 26466 42264 26584 42382 sw
tri 26748 42264 26866 42382 ne
rect 26866 42264 30851 42382
rect 22524 42080 26584 42264
rect 20604 41871 22232 42080
tri 22232 41871 22441 42080 sw
tri 22524 41871 22733 42080 ne
rect 22733 41982 26584 42080
tri 26584 41982 26866 42264 sw
tri 26866 41982 27148 42264 ne
rect 27148 42226 30851 42264
tri 30851 42226 31148 42523 sw
tri 31148 42226 31445 42523 ne
rect 31445 42440 33120 42523
tri 33120 42440 33211 42531 sw
tri 33409 42440 33500 42531 ne
rect 33500 42440 35190 42531
tri 35190 42440 35480 42730 sw
tri 35480 42440 35770 42730 ne
rect 35770 42530 39630 42730
tri 39630 42530 39924 42824 sw
tri 39924 42530 40218 42824 ne
rect 40218 42732 44039 42824
tri 44039 42732 44260 42953 sw
tri 44327 42732 44548 42953 ne
rect 44548 42750 48477 42953
tri 48477 42750 48774 43047 sw
tri 48774 42750 49071 43047 ne
rect 49071 42981 53008 43047
tri 53008 42981 53084 43057 sw
tri 53301 42981 53377 43057 ne
rect 53377 42981 55066 43057
rect 49071 42750 53084 42981
rect 44548 42749 48774 42750
tri 48774 42749 48775 42750 sw
tri 49071 42749 49072 42750 ne
rect 49072 42749 53084 42750
rect 44548 42732 48775 42749
rect 40218 42530 44260 42732
rect 35770 42440 39924 42530
rect 31445 42226 33211 42440
rect 27148 42225 31148 42226
tri 31148 42225 31149 42226 sw
tri 31445 42225 31446 42226 ne
rect 31446 42225 33211 42226
rect 27148 41982 31149 42225
rect 22733 41981 26866 41982
tri 26866 41981 26867 41982 sw
tri 27148 41981 27149 41982 ne
rect 27149 41981 31149 41982
rect 22733 41871 26867 41981
rect 20604 41579 22441 41871
tri 22441 41579 22733 41871 sw
tri 22733 41579 23025 41871 ne
rect 23025 41699 26867 41871
tri 26867 41699 27149 41981 sw
tri 27149 41699 27431 41981 ne
rect 27431 41928 31149 41981
tri 31149 41928 31446 42225 sw
tri 31446 41928 31743 42225 ne
rect 31743 42151 33211 42225
tri 33211 42151 33500 42440 sw
tri 33500 42151 33789 42440 ne
rect 33789 42439 35480 42440
tri 35480 42439 35481 42440 sw
tri 35770 42439 35771 42440 ne
rect 35771 42439 39924 42440
rect 33789 42151 35481 42439
rect 31743 41928 33500 42151
rect 27431 41699 31446 41928
rect 23025 41698 27149 41699
tri 27149 41698 27150 41699 sw
tri 27431 41698 27432 41699 ne
rect 27432 41698 31446 41699
rect 23025 41579 27150 41698
rect 20604 41415 22733 41579
tri 22733 41415 22897 41579 sw
tri 23025 41415 23189 41579 ne
rect 23189 41416 27150 41579
tri 27150 41416 27432 41698 sw
tri 27432 41416 27714 41698 ne
rect 27714 41631 31446 41698
tri 31446 41631 31743 41928 sw
tri 31743 41631 32040 41928 ne
rect 32040 41862 33500 41928
tri 33500 41862 33789 42151 sw
tri 33789 41862 34078 42151 ne
rect 34078 42149 35481 42151
tri 35481 42149 35771 42439 sw
tri 35771 42149 36061 42439 ne
rect 36061 42438 39924 42439
tri 39924 42438 40016 42530 sw
tri 40218 42438 40310 42530 ne
rect 40310 42444 44260 42530
tri 44260 42444 44548 42732 sw
tri 44548 42444 44836 42732 ne
rect 44836 42452 48775 42732
tri 48775 42452 49072 42749 sw
tri 49072 42452 49369 42749 ne
rect 49369 42688 53084 42749
tri 53084 42688 53377 42981 sw
tri 53377 42688 53670 42981 ne
rect 53670 42980 55066 42981
tri 55066 42980 55358 43272 sw
tri 55358 42980 55650 43272 ne
rect 55650 43175 57148 43272
tri 57148 43175 57435 43462 sw
tri 57435 43175 57722 43462 ne
rect 57722 43175 71000 43462
rect 55650 42980 57435 43175
rect 53670 42688 55358 42980
tri 55358 42688 55650 42980 sw
tri 55650 42688 55942 42980 ne
rect 55942 42888 57435 42980
tri 57435 42888 57722 43175 sw
tri 57722 42888 58009 43175 ne
rect 58009 42888 71000 43175
rect 55942 42800 57722 42888
tri 57722 42800 57810 42888 sw
tri 58009 42800 58097 42888 ne
rect 58097 42800 71000 42888
rect 55942 42688 57810 42800
rect 49369 42687 53377 42688
tri 53377 42687 53378 42688 sw
tri 53670 42687 53671 42688 ne
rect 53671 42687 55650 42688
rect 49369 42452 53378 42687
rect 44836 42451 49072 42452
tri 49072 42451 49073 42452 sw
tri 49369 42451 49370 42452 ne
rect 49370 42451 53378 42452
rect 44836 42444 49073 42451
rect 40310 42438 44548 42444
rect 36061 42149 40016 42438
rect 34078 41862 35771 42149
rect 32040 41707 33789 41862
tri 33789 41707 33944 41862 sw
tri 34078 41707 34233 41862 ne
rect 34233 41859 35771 41862
tri 35771 41859 36061 42149 sw
tri 36061 41859 36351 42149 ne
rect 36351 42144 40016 42149
tri 40016 42144 40310 42438 sw
tri 40310 42144 40604 42438 ne
rect 40604 42354 44548 42438
tri 44548 42354 44638 42444 sw
tri 44836 42354 44926 42444 ne
rect 44926 42354 49073 42444
rect 40604 42144 44638 42354
rect 36351 41939 40310 42144
tri 40310 41939 40515 42144 sw
tri 40604 41939 40809 42144 ne
rect 40809 42066 44638 42144
tri 44638 42066 44926 42354 sw
tri 44926 42066 45214 42354 ne
rect 45214 42154 49073 42354
tri 49073 42154 49370 42451 sw
tri 49370 42154 49667 42451 ne
rect 49667 42394 53378 42451
tri 53378 42394 53671 42687 sw
tri 53671 42394 53964 42687 ne
rect 53964 42600 55650 42687
tri 55650 42600 55738 42688 sw
tri 55942 42600 56030 42688 ne
rect 56030 42600 57810 42688
tri 57810 42600 58010 42800 sw
rect 53964 42394 55738 42600
rect 49667 42393 53671 42394
tri 53671 42393 53672 42394 sw
tri 53964 42393 53965 42394 ne
rect 53965 42393 55738 42394
rect 49667 42154 53672 42393
rect 45214 42152 49370 42154
tri 49370 42152 49372 42154 sw
tri 49667 42152 49669 42154 ne
rect 49669 42152 53672 42154
rect 45214 42066 49372 42152
rect 40809 42065 44926 42066
tri 44926 42065 44927 42066 sw
tri 45214 42065 45215 42066 ne
rect 45215 42065 49372 42066
rect 40809 41939 44927 42065
rect 36351 41859 40515 41939
rect 34233 41858 36061 41859
tri 36061 41858 36062 41859 sw
tri 36351 41858 36352 41859 ne
rect 36352 41858 40515 41859
rect 34233 41707 36062 41858
rect 32040 41631 33944 41707
rect 27714 41416 31743 41631
rect 23189 41415 27432 41416
rect 20604 41123 22897 41415
tri 22897 41123 23189 41415 sw
tri 23189 41123 23481 41415 ne
rect 23481 41338 27432 41415
tri 27432 41338 27510 41416 sw
tri 27714 41338 27792 41416 ne
rect 27792 41338 31743 41416
rect 23481 41123 27510 41338
rect 20604 41121 23189 41123
tri 23189 41121 23191 41123 sw
tri 23481 41121 23483 41123 ne
rect 23483 41121 27510 41123
rect 20604 40829 23191 41121
tri 23191 40829 23483 41121 sw
tri 23483 40829 23775 41121 ne
rect 23775 41056 27510 41121
tri 27510 41056 27792 41338 sw
tri 27792 41056 28074 41338 ne
rect 28074 41334 31743 41338
tri 31743 41334 32040 41631 sw
tri 32040 41334 32337 41631 ne
rect 32337 41418 33944 41631
tri 33944 41418 34233 41707 sw
tri 34233 41418 34522 41707 ne
rect 34522 41568 36062 41707
tri 36062 41568 36352 41858 sw
tri 36352 41568 36642 41858 ne
rect 36642 41645 40515 41858
tri 40515 41645 40809 41939 sw
tri 40809 41645 41103 41939 ne
rect 41103 41777 44927 41939
tri 44927 41777 45215 42065 sw
tri 45215 41777 45503 42065 ne
rect 45503 41856 49372 42065
tri 49372 41856 49668 42152 sw
tri 49669 41856 49965 42152 ne
rect 49965 42100 53672 42152
tri 53672 42100 53965 42393 sw
tri 53965 42100 54258 42393 ne
rect 54258 42308 55738 42393
tri 55738 42308 56030 42600 sw
tri 56030 42308 56322 42600 ne
rect 56322 42308 71000 42600
rect 54258 42100 56030 42308
rect 49965 41856 53965 42100
rect 45503 41777 49668 41856
rect 41103 41775 45215 41777
tri 45215 41775 45217 41777 sw
tri 45503 41775 45505 41777 ne
rect 45505 41775 49668 41777
rect 41103 41645 45217 41775
rect 36642 41568 40809 41645
rect 34522 41418 36352 41568
rect 32337 41334 34233 41418
rect 28074 41138 32040 41334
tri 32040 41138 32236 41334 sw
tri 32337 41138 32533 41334 ne
rect 32533 41138 34233 41334
rect 28074 41056 32236 41138
rect 23775 40848 27792 41056
tri 27792 40848 28000 41056 sw
tri 28074 40848 28282 41056 ne
rect 28282 40848 32236 41056
rect 23775 40829 28000 40848
rect 20604 40828 23483 40829
tri 23483 40828 23484 40829 sw
tri 23775 40828 23776 40829 ne
rect 23776 40828 28000 40829
rect 20604 40536 23484 40828
tri 23484 40536 23776 40828 sw
tri 23776 40536 24068 40828 ne
rect 24068 40566 28000 40828
tri 28000 40566 28282 40848 sw
tri 28282 40566 28564 40848 ne
rect 28564 40841 32236 40848
tri 32236 40841 32533 41138 sw
tri 32533 40841 32830 41138 ne
rect 32830 41129 34233 41138
tri 34233 41129 34522 41418 sw
tri 34522 41129 34811 41418 ne
rect 34811 41331 36352 41418
tri 36352 41331 36589 41568 sw
tri 36642 41331 36879 41568 ne
rect 36879 41486 40809 41568
tri 40809 41486 40968 41645 sw
tri 41103 41486 41262 41645 ne
rect 41262 41488 45217 41645
tri 45217 41488 45504 41775 sw
tri 45505 41488 45792 41775 ne
rect 45792 41636 49668 41775
tri 49668 41636 49888 41856 sw
tri 49965 41636 50185 41856 ne
rect 50185 41807 53965 41856
tri 53965 41807 54258 42100 sw
tri 54258 41807 54551 42100 ne
rect 54551 42016 56030 42100
tri 56030 42016 56322 42308 sw
tri 56322 42016 56614 42308 ne
rect 56614 42016 71000 42308
rect 54551 41876 56322 42016
tri 56322 41876 56462 42016 sw
tri 56614 41876 56754 42016 ne
rect 56754 41876 71000 42016
rect 54551 41807 56462 41876
rect 50185 41636 54258 41807
rect 45792 41488 49888 41636
rect 41262 41486 45504 41488
rect 36879 41331 40968 41486
rect 34811 41129 36589 41331
rect 32830 40841 34522 41129
rect 28564 40566 32533 40841
rect 24068 40536 28282 40566
rect 20604 40535 23776 40536
tri 23776 40535 23777 40536 sw
tri 24068 40535 24069 40536 ne
rect 24069 40535 28282 40536
rect 20604 40243 23777 40535
tri 23777 40243 24069 40535 sw
tri 24069 40243 24361 40535 ne
rect 24361 40372 28282 40535
tri 28282 40372 28476 40566 sw
tri 28564 40372 28758 40566 ne
rect 28758 40544 32533 40566
tri 32533 40544 32830 40841 sw
tri 32830 40544 33127 40841 ne
rect 33127 40840 34522 40841
tri 34522 40840 34811 41129 sw
tri 34811 40840 35100 41129 ne
rect 35100 41041 36589 41129
tri 36589 41041 36879 41331 sw
tri 36879 41041 37169 41331 ne
rect 37169 41192 40968 41331
tri 40968 41192 41262 41486 sw
tri 41262 41192 41556 41486 ne
rect 41556 41400 45504 41486
tri 45504 41400 45592 41488 sw
tri 45792 41400 45880 41488 ne
rect 45880 41400 49888 41488
rect 41556 41192 45592 41400
rect 37169 41191 41262 41192
tri 41262 41191 41263 41192 sw
tri 41556 41191 41557 41192 ne
rect 41557 41191 45592 41192
rect 37169 41041 41263 41191
rect 35100 40840 36879 41041
rect 33127 40551 34811 40840
tri 34811 40551 35100 40840 sw
tri 35100 40551 35389 40840 ne
rect 35389 40751 36879 40840
tri 36879 40751 37169 41041 sw
tri 37169 40751 37459 41041 ne
rect 37459 40897 41263 41041
tri 41263 40897 41557 41191 sw
tri 41557 40897 41851 41191 ne
rect 41851 41112 45592 41191
tri 45592 41112 45880 41400 sw
tri 45880 41112 46168 41400 ne
rect 46168 41391 49888 41400
tri 49888 41391 50133 41636 sw
tri 50185 41391 50430 41636 ne
rect 50430 41588 54258 41636
tri 54258 41588 54477 41807 sw
tri 54551 41588 54770 41807 ne
rect 54770 41588 56462 41807
rect 50430 41391 54477 41588
rect 46168 41338 50133 41391
tri 50133 41338 50186 41391 sw
tri 50430 41338 50483 41391 ne
rect 50483 41338 54477 41391
rect 46168 41112 50186 41338
rect 41851 40908 45880 41112
tri 45880 40908 46084 41112 sw
tri 46168 40908 46372 41112 ne
rect 46372 41041 50186 41112
tri 50186 41041 50483 41338 sw
tri 50483 41041 50780 41338 ne
rect 50780 41295 54477 41338
tri 54477 41295 54770 41588 sw
tri 54770 41295 55063 41588 ne
rect 55063 41584 56462 41588
tri 56462 41584 56754 41876 sw
tri 56754 41584 57046 41876 ne
rect 57046 41584 71000 41876
rect 55063 41295 56754 41584
rect 50780 41294 54770 41295
tri 54770 41294 54771 41295 sw
tri 55063 41294 55064 41295 ne
rect 55064 41294 56754 41295
rect 50780 41041 54771 41294
rect 46372 41040 50483 41041
tri 50483 41040 50484 41041 sw
tri 50780 41040 50781 41041 ne
rect 50781 41040 54771 41041
rect 46372 40908 50484 41040
rect 41851 40897 46084 40908
rect 37459 40896 41557 40897
tri 41557 40896 41558 40897 sw
tri 41851 40896 41852 40897 ne
rect 41852 40896 46084 40897
rect 37459 40751 41558 40896
rect 35389 40750 37169 40751
tri 37169 40750 37170 40751 sw
tri 37459 40750 37460 40751 ne
rect 37460 40750 41558 40751
rect 35389 40551 37170 40750
rect 33127 40544 35100 40551
rect 28758 40372 32830 40544
tri 32830 40372 33002 40544 sw
tri 33127 40372 33299 40544 ne
rect 33299 40460 35100 40544
tri 35100 40460 35191 40551 sw
tri 35389 40460 35480 40551 ne
rect 35480 40460 37170 40551
tri 37170 40460 37460 40750 sw
tri 37460 40460 37750 40750 ne
rect 37750 40602 41558 40750
tri 41558 40602 41852 40896 sw
tri 41852 40602 42146 40896 ne
rect 42146 40620 46084 40896
tri 46084 40620 46372 40908 sw
tri 46372 40620 46660 40908 ne
rect 46660 40743 50484 40908
tri 50484 40743 50781 41040 sw
tri 50781 40743 51078 41040 ne
rect 51078 41001 54771 41040
tri 54771 41001 55064 41294 sw
tri 55064 41001 55357 41294 ne
rect 55357 41292 56754 41294
tri 56754 41292 57046 41584 sw
tri 57046 41292 57338 41584 ne
rect 57338 41292 71000 41584
rect 55357 41001 57046 41292
rect 51078 40743 55064 41001
rect 46660 40742 50781 40743
tri 50781 40742 50782 40743 sw
tri 51078 40742 51079 40743 ne
rect 51079 40742 55064 40743
rect 46660 40620 50782 40742
rect 42146 40602 46372 40620
rect 37750 40601 41852 40602
tri 41852 40601 41853 40602 sw
tri 42146 40601 42147 40602 ne
rect 42147 40601 46372 40602
rect 37750 40460 41853 40601
rect 33299 40372 35191 40460
rect 24361 40243 28476 40372
rect 20604 40242 24069 40243
tri 24069 40242 24070 40243 sw
tri 24361 40242 24362 40243 ne
rect 24362 40242 28476 40243
rect 20604 39950 24070 40242
tri 24070 39950 24362 40242 sw
tri 24362 39950 24654 40242 ne
rect 24654 40090 28476 40242
tri 28476 40090 28758 40372 sw
tri 28758 40090 29040 40372 ne
rect 29040 40090 33002 40372
rect 24654 40089 28758 40090
tri 28758 40089 28759 40090 sw
tri 29040 40089 29041 40090 ne
rect 29041 40089 33002 40090
rect 24654 39950 28759 40089
rect 20604 39949 24362 39950
tri 24362 39949 24363 39950 sw
tri 24654 39949 24655 39950 ne
rect 24655 39949 28759 39950
rect 20604 39657 24363 39949
tri 24363 39657 24655 39949 sw
tri 24655 39657 24947 39949 ne
rect 24947 39807 28759 39949
tri 28759 39807 29041 40089 sw
tri 29041 39807 29323 40089 ne
rect 29323 40075 33002 40089
tri 33002 40075 33299 40372 sw
tri 33299 40075 33596 40372 ne
rect 33596 40171 35191 40372
tri 35191 40171 35480 40460 sw
tri 35480 40171 35769 40460 ne
rect 35769 40459 37460 40460
tri 37460 40459 37461 40460 sw
tri 37750 40459 37751 40460 ne
rect 37751 40459 41853 40460
rect 35769 40171 37461 40459
rect 33596 40075 35480 40171
rect 29323 40074 33299 40075
tri 33299 40074 33300 40075 sw
tri 33596 40074 33597 40075 ne
rect 33597 40074 35480 40075
rect 29323 39807 33300 40074
rect 24947 39805 29041 39807
tri 29041 39805 29043 39807 sw
tri 29323 39805 29325 39807 ne
rect 29325 39805 33300 39807
rect 24947 39657 29043 39805
rect 20604 39464 24655 39657
tri 24655 39464 24848 39657 sw
tri 24947 39464 25140 39657 ne
rect 25140 39523 29043 39657
tri 29043 39523 29325 39805 sw
tri 29325 39523 29607 39805 ne
rect 29607 39777 33300 39805
tri 33300 39777 33597 40074 sw
tri 33597 39777 33894 40074 ne
rect 33894 39882 35480 40074
tri 35480 39882 35769 40171 sw
tri 35769 39882 36058 40171 ne
rect 36058 40169 37461 40171
tri 37461 40169 37751 40459 sw
tri 37751 40169 38041 40459 ne
rect 38041 40307 41853 40459
tri 41853 40307 42147 40601 sw
tri 42147 40307 42441 40601 ne
rect 42441 40443 46372 40601
tri 46372 40443 46549 40620 sw
tri 46660 40443 46837 40620 ne
rect 46837 40445 50782 40620
tri 50782 40445 51079 40742 sw
tri 51079 40445 51376 40742 ne
rect 51376 40708 55064 40742
tri 55064 40708 55357 41001 sw
tri 55357 40708 55650 41001 ne
rect 55650 41000 57046 41001
tri 57046 41000 57338 41292 sw
tri 57338 41200 57430 41292 ne
rect 57430 41200 71000 41292
rect 55650 40708 71000 41000
rect 51376 40644 55357 40708
tri 55357 40644 55421 40708 sw
tri 55650 40644 55714 40708 ne
rect 55714 40644 71000 40708
rect 51376 40445 55421 40644
rect 46837 40443 51079 40445
rect 42441 40307 46549 40443
rect 38041 40305 42147 40307
tri 42147 40305 42149 40307 sw
tri 42441 40305 42443 40307 ne
rect 42443 40305 46549 40307
rect 38041 40169 42149 40305
rect 36058 39882 37751 40169
rect 33894 39777 35769 39882
rect 29607 39523 33597 39777
rect 25140 39522 29325 39523
tri 29325 39522 29326 39523 sw
tri 29607 39522 29608 39523 ne
rect 29608 39522 33597 39523
rect 25140 39464 29326 39522
tri 20604 35220 24848 39464 ne
tri 24848 39172 25140 39464 sw
tri 25140 39172 25432 39464 ne
rect 25432 39240 29326 39464
tri 29326 39240 29608 39522 sw
tri 29608 39240 29890 39522 ne
rect 29890 39480 33597 39522
tri 33597 39480 33894 39777 sw
tri 33894 39480 34191 39777 ne
rect 34191 39653 35769 39777
tri 35769 39653 35998 39882 sw
tri 36058 39653 36287 39882 ne
rect 36287 39879 37751 39882
tri 37751 39879 38041 40169 sw
tri 38041 39879 38331 40169 ne
rect 38331 40011 42149 40169
tri 42149 40011 42443 40305 sw
tri 42443 40011 42737 40305 ne
rect 42737 40155 46549 40305
tri 46549 40155 46837 40443 sw
tri 46837 40155 47125 40443 ne
rect 47125 40347 51079 40443
tri 51079 40347 51177 40445 sw
tri 51376 40347 51474 40445 ne
rect 51474 40351 55421 40445
tri 55421 40351 55714 40644 sw
tri 55714 40351 56007 40644 ne
rect 56007 40351 71000 40644
rect 51474 40347 55714 40351
rect 47125 40155 51177 40347
rect 42737 40154 46837 40155
tri 46837 40154 46838 40155 sw
tri 47125 40154 47126 40155 ne
rect 47126 40154 51177 40155
rect 42737 40011 46838 40154
rect 38331 39879 42443 40011
rect 36287 39878 38041 39879
tri 38041 39878 38042 39879 sw
tri 38331 39878 38332 39879 ne
rect 38332 39878 42443 39879
rect 36287 39653 38042 39878
rect 34191 39480 35998 39653
rect 29890 39479 33894 39480
tri 33894 39479 33895 39480 sw
tri 34191 39479 34192 39480 ne
rect 34192 39479 35998 39480
rect 29890 39240 33895 39479
rect 25432 39239 29608 39240
tri 29608 39239 29609 39240 sw
tri 29890 39239 29891 39240 ne
rect 29891 39239 33895 39240
rect 25432 39172 29609 39239
rect 24848 39094 25140 39172
tri 25140 39094 25218 39172 sw
tri 25432 39094 25510 39172 ne
rect 25510 39094 29609 39172
rect 24848 38802 25218 39094
tri 25218 38802 25510 39094 sw
tri 25510 38802 25802 39094 ne
rect 25802 38957 29609 39094
tri 29609 38957 29891 39239 sw
tri 29891 38957 30173 39239 ne
rect 30173 39182 33895 39239
tri 33895 39182 34192 39479 sw
tri 34192 39182 34489 39479 ne
rect 34489 39438 35998 39479
tri 35998 39438 36213 39653 sw
tri 36287 39438 36502 39653 ne
rect 36502 39588 38042 39653
tri 38042 39588 38332 39878 sw
tri 38332 39588 38622 39878 ne
rect 38622 39717 42443 39878
tri 42443 39717 42737 40011 sw
tri 42737 39717 43031 40011 ne
rect 43031 39866 46838 40011
tri 46838 39866 47126 40154 sw
tri 47126 39866 47414 40154 ne
rect 47414 40050 51177 40154
tri 51177 40050 51474 40347 sw
tri 51474 40050 51771 40347 ne
rect 51771 40120 55714 40347
tri 55714 40120 55945 40351 sw
tri 56007 40120 56238 40351 ne
rect 56238 40120 71000 40351
rect 51771 40050 55945 40120
rect 47414 39866 51474 40050
rect 43031 39865 47126 39866
tri 47126 39865 47127 39866 sw
tri 47414 39865 47415 39866 ne
rect 47415 39865 51474 39866
rect 43031 39717 47127 39865
rect 38622 39588 42737 39717
rect 36502 39438 38332 39588
rect 34489 39182 36213 39438
rect 30173 39158 34192 39182
tri 34192 39158 34216 39182 sw
tri 34489 39158 34513 39182 ne
rect 34513 39158 36213 39182
rect 30173 38957 34216 39158
rect 25802 38956 29891 38957
tri 29891 38956 29892 38957 sw
tri 30173 38956 30174 38957 ne
rect 30174 38956 34216 38957
rect 25802 38802 29892 38956
rect 24848 38801 25510 38802
tri 25510 38801 25511 38802 sw
tri 25802 38801 25803 38802 ne
rect 25803 38801 29892 38802
rect 24848 38509 25511 38801
tri 25511 38509 25803 38801 sw
tri 25803 38509 26095 38801 ne
rect 26095 38674 29892 38801
tri 29892 38674 30174 38956 sw
tri 30174 38674 30456 38956 ne
rect 30456 38861 34216 38956
tri 34216 38861 34513 39158 sw
tri 34513 38861 34810 39158 ne
rect 34810 39149 36213 39158
tri 36213 39149 36502 39438 sw
tri 36502 39149 36791 39438 ne
rect 36791 39352 38332 39438
tri 38332 39352 38568 39588 sw
tri 38622 39352 38858 39588 ne
rect 38858 39467 42737 39588
tri 42737 39467 42987 39717 sw
tri 43031 39467 43281 39717 ne
rect 43281 39577 47127 39717
tri 47127 39577 47415 39865 sw
tri 47415 39577 47703 39865 ne
rect 47703 39847 51474 39865
tri 51474 39847 51677 40050 sw
tri 51771 39847 51974 40050 ne
rect 51974 39988 55945 40050
tri 55945 39988 56077 40120 sw
tri 56238 39988 56370 40120 ne
rect 56370 39988 71000 40120
rect 51974 39847 56077 39988
rect 47703 39577 51677 39847
rect 43281 39576 47415 39577
tri 47415 39576 47416 39577 sw
tri 47703 39576 47704 39577 ne
rect 47704 39576 51677 39577
rect 43281 39467 47416 39576
rect 38858 39352 42987 39467
rect 36791 39242 38568 39352
tri 38568 39242 38678 39352 sw
tri 38858 39242 38968 39352 ne
rect 38968 39242 42987 39352
rect 36791 39149 38678 39242
rect 34810 38861 36502 39149
rect 30456 38674 34513 38861
rect 26095 38509 30174 38674
rect 24848 38508 25803 38509
tri 25803 38508 25804 38509 sw
tri 26095 38508 26096 38509 ne
rect 26096 38508 30174 38509
rect 24848 38216 25804 38508
tri 25804 38216 26096 38508 sw
tri 26096 38216 26388 38508 ne
rect 26388 38420 30174 38508
tri 30174 38420 30428 38674 sw
tri 30456 38420 30710 38674 ne
rect 30710 38564 34513 38674
tri 34513 38564 34810 38861 sw
tri 34810 38564 35107 38861 ne
rect 35107 38860 36502 38861
tri 36502 38860 36791 39149 sw
tri 36791 38860 37080 39149 ne
rect 37080 39061 38678 39149
tri 38678 39061 38859 39242 sw
tri 38968 39061 39149 39242 ne
rect 39149 39238 42987 39242
tri 42987 39238 43216 39467 sw
tri 43281 39238 43510 39467 ne
rect 43510 39288 47416 39467
tri 47416 39288 47704 39576 sw
tri 47704 39288 47992 39576 ne
rect 47992 39550 51677 39576
tri 51677 39550 51974 39847 sw
tri 51974 39550 52271 39847 ne
rect 52271 39695 56077 39847
tri 56077 39695 56370 39988 sw
tri 56370 39695 56663 39988 ne
rect 56663 39695 71000 39988
rect 52271 39694 56370 39695
tri 56370 39694 56371 39695 sw
tri 56663 39694 56664 39695 ne
rect 56664 39694 71000 39695
rect 52271 39550 56371 39694
rect 47992 39401 51974 39550
tri 51974 39401 52123 39550 sw
tri 52271 39401 52420 39550 ne
rect 52420 39401 56371 39550
tri 56371 39401 56664 39694 sw
tri 56664 39600 56758 39694 ne
rect 56758 39600 71000 39694
rect 47992 39288 52123 39401
rect 43510 39287 47704 39288
tri 47704 39287 47705 39288 sw
tri 47992 39287 47993 39288 ne
rect 47993 39287 52123 39288
rect 43510 39238 47705 39287
rect 39149 39172 43216 39238
tri 43216 39172 43282 39238 sw
tri 43510 39172 43576 39238 ne
rect 43576 39172 47705 39238
rect 39149 39061 43282 39172
rect 37080 38860 38859 39061
rect 35107 38571 36791 38860
tri 36791 38571 37080 38860 sw
tri 37080 38571 37369 38860 ne
rect 37369 38771 38859 38860
tri 38859 38771 39149 39061 sw
tri 39149 38771 39439 39061 ne
rect 39439 38878 43282 39061
tri 43282 38878 43576 39172 sw
tri 43576 38878 43870 39172 ne
rect 43870 38999 47705 39172
tri 47705 38999 47993 39287 sw
tri 47993 38999 48281 39287 ne
rect 48281 39104 52123 39287
tri 52123 39104 52420 39401 sw
tri 52420 39104 52717 39401 ne
rect 52717 39400 56664 39401
tri 56664 39400 56665 39401 sw
rect 52717 39104 71000 39400
rect 48281 39102 52420 39104
tri 52420 39102 52422 39104 sw
tri 52717 39102 52719 39104 ne
rect 52719 39102 71000 39104
rect 48281 38999 52422 39102
rect 43870 38997 47993 38999
tri 47993 38997 47995 38999 sw
tri 48281 38997 48283 38999 ne
rect 48283 38997 52422 38999
rect 43870 38878 47995 38997
rect 39439 38877 43576 38878
tri 43576 38877 43577 38878 sw
tri 43870 38877 43871 38878 ne
rect 43871 38877 47995 38878
rect 39439 38771 43577 38877
rect 37369 38770 39149 38771
tri 39149 38770 39150 38771 sw
tri 39439 38770 39440 38771 ne
rect 39440 38770 43577 38771
rect 37369 38571 39150 38770
rect 35107 38564 37080 38571
rect 30710 38563 34810 38564
tri 34810 38563 34811 38564 sw
tri 35107 38563 35108 38564 ne
rect 35108 38563 37080 38564
rect 30710 38420 34811 38563
rect 26388 38216 30428 38420
rect 24848 38128 26096 38216
tri 26096 38128 26184 38216 sw
tri 26388 38128 26476 38216 ne
rect 26476 38138 30428 38216
tri 30428 38138 30710 38420 sw
tri 30710 38138 30992 38420 ne
rect 30992 38266 34811 38420
tri 34811 38266 35108 38563 sw
tri 35108 38266 35405 38563 ne
rect 35405 38406 37080 38563
tri 37080 38406 37245 38571 sw
tri 37369 38406 37534 38571 ne
rect 37534 38480 39150 38571
tri 39150 38480 39440 38770 sw
tri 39440 38480 39730 38770 ne
rect 39730 38583 43577 38770
tri 43577 38583 43871 38877 sw
tri 43871 38583 44165 38877 ne
rect 44165 38710 47995 38877
tri 47995 38710 48282 38997 sw
tri 48283 38710 48570 38997 ne
rect 48570 38805 52422 38997
tri 52422 38805 52719 39102 sw
tri 52719 38805 53016 39102 ne
rect 53016 38805 71000 39102
rect 48570 38804 52719 38805
tri 52719 38804 52720 38805 sw
tri 53016 38804 53017 38805 ne
rect 53017 38804 71000 38805
rect 48570 38710 52720 38804
rect 44165 38583 48282 38710
rect 39730 38581 43871 38583
tri 43871 38581 43873 38583 sw
tri 44165 38581 44167 38583 ne
rect 44167 38581 48282 38583
rect 39730 38480 43873 38581
rect 37534 38406 39440 38480
rect 35405 38266 37245 38406
rect 30992 38265 35108 38266
tri 35108 38265 35109 38266 sw
tri 35405 38265 35406 38266 ne
rect 35406 38265 37245 38266
rect 30992 38138 35109 38265
rect 26476 38128 30710 38138
rect 24848 37836 26184 38128
tri 26184 37836 26476 38128 sw
tri 26476 37836 26768 38128 ne
rect 26768 38021 30710 38128
tri 30710 38021 30827 38138 sw
tri 30992 38021 31109 38138 ne
rect 31109 38021 35109 38138
rect 26768 37836 30827 38021
rect 24848 37628 26476 37836
tri 26476 37628 26684 37836 sw
tri 26768 37628 26976 37836 ne
rect 26976 37739 30827 37836
tri 30827 37739 31109 38021 sw
tri 31109 37739 31391 38021 ne
rect 31391 37968 35109 38021
tri 35109 37968 35406 38265 sw
tri 35406 37968 35703 38265 ne
rect 35703 38191 37245 38265
tri 37245 38191 37460 38406 sw
tri 37534 38191 37749 38406 ne
rect 37749 38285 39440 38406
tri 39440 38285 39635 38480 sw
tri 39730 38285 39925 38480 ne
rect 39925 38288 43873 38480
tri 43873 38288 44166 38581 sw
tri 44167 38288 44460 38581 ne
rect 44460 38488 48282 38581
tri 48282 38488 48504 38710 sw
tri 48570 38488 48792 38710 ne
rect 48792 38507 52720 38710
tri 52720 38507 53017 38804 sw
tri 53017 38507 53314 38804 ne
rect 53314 38507 71000 38804
rect 48792 38506 53017 38507
tri 53017 38506 53018 38507 sw
tri 53314 38506 53315 38507 ne
rect 53315 38506 71000 38507
rect 48792 38488 53018 38506
rect 44460 38288 48504 38488
rect 39925 38285 44166 38288
rect 37749 38191 39635 38285
rect 35703 37968 37460 38191
rect 31391 37739 35406 37968
rect 26976 37738 31109 37739
tri 31109 37738 31110 37739 sw
tri 31391 37738 31392 37739 ne
rect 31392 37738 35406 37739
rect 26976 37628 31110 37738
rect 24848 37337 26684 37628
tri 26684 37337 26975 37628 sw
tri 26976 37337 27267 37628 ne
rect 27267 37456 31110 37628
tri 31110 37456 31392 37738 sw
tri 31392 37456 31674 37738 ne
rect 31674 37671 35406 37738
tri 35406 37671 35703 37968 sw
tri 35703 37671 36000 37968 ne
rect 36000 37902 37460 37968
tri 37460 37902 37749 38191 sw
tri 37749 37902 38038 38191 ne
rect 38038 37995 39635 38191
tri 39635 37995 39925 38285 sw
tri 39925 37995 40215 38285 ne
rect 40215 38194 44166 38285
tri 44166 38194 44260 38288 sw
tri 44460 38194 44554 38288 ne
rect 44554 38200 48504 38288
tri 48504 38200 48792 38488 sw
tri 48792 38200 49080 38488 ne
rect 49080 38209 53018 38488
tri 53018 38209 53315 38506 sw
tri 53315 38209 53612 38506 ne
rect 53612 38209 71000 38506
rect 49080 38208 53315 38209
tri 53315 38208 53316 38209 sw
tri 53612 38208 53613 38209 ne
rect 53613 38208 71000 38209
rect 49080 38200 53316 38208
rect 44554 38194 48792 38200
rect 40215 37995 44260 38194
rect 38038 37994 39925 37995
tri 39925 37994 39926 37995 sw
tri 40215 37994 40216 37995 ne
rect 40216 37994 44260 37995
rect 38038 37902 39926 37994
rect 36000 37747 37749 37902
tri 37749 37747 37904 37902 sw
tri 38038 37747 38193 37902 ne
rect 38193 37747 39926 37902
rect 36000 37671 37904 37747
rect 31674 37456 35703 37671
rect 27267 37455 31392 37456
tri 31392 37455 31393 37456 sw
tri 31674 37455 31675 37456 ne
rect 31675 37455 35703 37456
rect 27267 37337 31393 37455
rect 24848 37172 26975 37337
tri 26975 37172 27140 37337 sw
tri 27267 37172 27432 37337 ne
rect 27432 37173 31393 37337
tri 31393 37173 31675 37455 sw
tri 31675 37173 31957 37455 ne
rect 31957 37374 35703 37455
tri 35703 37374 36000 37671 sw
tri 36000 37374 36297 37671 ne
rect 36297 37458 37904 37671
tri 37904 37458 38193 37747 sw
tri 38193 37458 38482 37747 ne
rect 38482 37704 39926 37747
tri 39926 37704 40216 37994 sw
tri 40216 37704 40506 37994 ne
rect 40506 37900 44260 37994
tri 44260 37900 44554 38194 sw
tri 44554 37900 44848 38194 ne
rect 44848 38111 48792 38194
tri 48792 38111 48881 38200 sw
tri 49080 38111 49169 38200 ne
rect 49169 38111 53316 38200
rect 44848 37900 48881 38111
rect 40506 37704 44554 37900
rect 38482 37458 40216 37704
rect 36297 37374 38193 37458
rect 31957 37173 36000 37374
rect 27432 37172 31675 37173
rect 24848 36880 27140 37172
tri 27140 36880 27432 37172 sw
tri 27432 36880 27724 37172 ne
rect 27724 37094 31675 37172
tri 31675 37094 31754 37173 sw
tri 31957 37094 32036 37173 ne
rect 32036 37094 36000 37173
rect 27724 36880 31754 37094
rect 24848 36879 27432 36880
tri 27432 36879 27433 36880 sw
tri 27724 36879 27725 36880 ne
rect 27725 36879 31754 36880
rect 24848 36587 27433 36879
tri 27433 36587 27725 36879 sw
tri 27725 36587 28017 36879 ne
rect 28017 36812 31754 36879
tri 31754 36812 32036 37094 sw
tri 32036 36812 32318 37094 ne
rect 32318 37077 36000 37094
tri 36000 37077 36297 37374 sw
tri 36297 37077 36594 37374 ne
rect 36594 37169 38193 37374
tri 38193 37169 38482 37458 sw
tri 38482 37169 38771 37458 ne
rect 38771 37414 40216 37458
tri 40216 37414 40506 37704 sw
tri 40506 37414 40796 37704 ne
rect 40796 37696 44554 37704
tri 44554 37696 44758 37900 sw
tri 44848 37696 45052 37900 ne
rect 45052 37823 48881 37900
tri 48881 37823 49169 38111 sw
tri 49169 37823 49457 38111 ne
rect 49457 37911 53316 38111
tri 53316 37911 53613 38208 sw
tri 53613 37911 53910 38208 ne
rect 53910 37911 71000 38208
rect 49457 37910 53613 37911
tri 53613 37910 53614 37911 sw
tri 53910 37910 53911 37911 ne
rect 53911 37910 71000 37911
rect 49457 37823 53614 37910
rect 45052 37822 49169 37823
tri 49169 37822 49170 37823 sw
tri 49457 37822 49458 37823 ne
rect 49458 37822 53614 37823
rect 45052 37696 49170 37822
rect 40796 37414 44758 37696
rect 38771 37371 40506 37414
tri 40506 37371 40549 37414 sw
tri 40796 37371 40839 37414 ne
rect 40839 37402 44758 37414
tri 44758 37402 45052 37696 sw
tri 45052 37402 45346 37696 ne
rect 45346 37534 49170 37696
tri 49170 37534 49458 37822 sw
tri 49458 37534 49746 37822 ne
rect 49746 37613 53614 37822
tri 53614 37613 53911 37910 sw
tri 53911 37613 54208 37910 ne
rect 54208 37613 71000 37910
rect 49746 37534 53911 37613
rect 45346 37533 49458 37534
tri 49458 37533 49459 37534 sw
tri 49746 37533 49747 37534 ne
rect 49747 37533 53911 37534
rect 45346 37402 49459 37533
rect 40839 37371 45052 37402
rect 38771 37169 40549 37371
rect 36594 37077 38482 37169
rect 32318 36881 36297 37077
tri 36297 36881 36493 37077 sw
tri 36594 36881 36790 37077 ne
rect 36790 36881 38482 37077
rect 32318 36812 36493 36881
rect 28017 36605 32036 36812
tri 32036 36605 32243 36812 sw
tri 32318 36605 32525 36812 ne
rect 32525 36605 36493 36812
rect 28017 36587 32243 36605
rect 24848 36585 27725 36587
tri 27725 36585 27727 36587 sw
tri 28017 36585 28019 36587 ne
rect 28019 36585 32243 36587
rect 24848 36293 27727 36585
tri 27727 36293 28019 36585 sw
tri 28019 36293 28311 36585 ne
rect 28311 36323 32243 36585
tri 32243 36323 32525 36605 sw
tri 32525 36323 32807 36605 ne
rect 32807 36584 36493 36605
tri 36493 36584 36790 36881 sw
tri 36790 36584 37087 36881 ne
rect 37087 36880 38482 36881
tri 38482 36880 38771 37169 sw
tri 38771 36880 39060 37169 ne
rect 39060 37081 40549 37169
tri 40549 37081 40839 37371 sw
tri 40839 37081 41129 37371 ne
rect 41129 37243 45052 37371
tri 45052 37243 45211 37402 sw
tri 45346 37243 45505 37402 ne
rect 45505 37245 49459 37402
tri 49459 37245 49747 37533 sw
tri 49747 37245 50035 37533 ne
rect 50035 37393 53911 37533
tri 53911 37393 54131 37613 sw
tri 54208 37393 54428 37613 ne
rect 54428 37393 71000 37613
rect 50035 37245 54131 37393
rect 45505 37243 49747 37245
rect 41129 37081 45211 37243
rect 39060 36880 40839 37081
rect 37087 36591 38771 36880
tri 38771 36591 39060 36880 sw
tri 39060 36591 39349 36880 ne
rect 39349 36791 40839 36880
tri 40839 36791 41129 37081 sw
tri 41129 36791 41419 37081 ne
rect 41419 36949 45211 37081
tri 45211 36949 45505 37243 sw
tri 45505 36949 45799 37243 ne
rect 45799 37156 49747 37243
tri 49747 37156 49836 37245 sw
tri 50035 37156 50124 37245 ne
rect 50124 37156 54131 37245
rect 45799 36949 49836 37156
rect 41419 36948 45505 36949
tri 45505 36948 45506 36949 sw
tri 45799 36948 45800 36949 ne
rect 45800 36948 49836 36949
rect 41419 36791 45506 36948
rect 39349 36790 41129 36791
tri 41129 36790 41130 36791 sw
tri 41419 36790 41420 36791 ne
rect 41420 36790 45506 36791
rect 39349 36591 41130 36790
rect 37087 36584 39060 36591
rect 32807 36583 36790 36584
tri 36790 36583 36791 36584 sw
tri 37087 36583 37088 36584 ne
rect 37088 36583 39060 36584
rect 32807 36323 36791 36583
rect 28311 36293 32525 36323
rect 24848 36292 28019 36293
tri 28019 36292 28020 36293 sw
tri 28311 36292 28312 36293 ne
rect 28312 36292 32525 36293
rect 24848 36000 28020 36292
tri 28020 36000 28312 36292 sw
tri 28312 36000 28604 36292 ne
rect 28604 36129 32525 36292
tri 32525 36129 32719 36323 sw
tri 32807 36129 33001 36323 ne
rect 33001 36286 36791 36323
tri 36791 36286 37088 36583 sw
tri 37088 36286 37385 36583 ne
rect 37385 36500 39060 36583
tri 39060 36500 39151 36591 sw
tri 39349 36500 39440 36591 ne
rect 39440 36500 41130 36591
tri 41130 36500 41420 36790 sw
tri 41420 36500 41710 36790 ne
rect 41710 36654 45506 36790
tri 45506 36654 45800 36948 sw
tri 45800 36654 46094 36948 ne
rect 46094 36868 49836 36948
tri 49836 36868 50124 37156 sw
tri 50124 36868 50412 37156 ne
rect 50412 37147 54131 37156
tri 54131 37147 54377 37393 sw
tri 54428 37147 54674 37393 ne
rect 54674 37147 71000 37393
rect 50412 37095 54377 37147
tri 54377 37095 54429 37147 sw
tri 54674 37095 54726 37147 ne
rect 54726 37095 71000 37147
rect 50412 36868 54429 37095
rect 46094 36665 50124 36868
tri 50124 36665 50327 36868 sw
tri 50412 36665 50615 36868 ne
rect 50615 36798 54429 36868
tri 54429 36798 54726 37095 sw
tri 54726 36798 55023 37095 ne
rect 55023 36798 71000 37095
rect 50615 36797 54726 36798
tri 54726 36797 54727 36798 sw
tri 55023 36797 55024 36798 ne
rect 55024 36797 71000 36798
rect 50615 36665 54727 36797
rect 46094 36654 50327 36665
rect 41710 36653 45800 36654
tri 45800 36653 45801 36654 sw
tri 46094 36653 46095 36654 ne
rect 46095 36653 50327 36654
rect 41710 36500 45801 36653
rect 37385 36286 39151 36500
rect 33001 36129 37088 36286
tri 37088 36129 37245 36286 sw
tri 37385 36129 37542 36286 ne
rect 37542 36211 39151 36286
tri 39151 36211 39440 36500 sw
tri 39440 36211 39729 36500 ne
rect 39729 36499 41420 36500
tri 41420 36499 41421 36500 sw
tri 41710 36499 41711 36500 ne
rect 41711 36499 45801 36500
rect 39729 36211 41421 36499
rect 37542 36129 39440 36211
rect 28604 36000 32719 36129
rect 24848 35999 28312 36000
tri 28312 35999 28313 36000 sw
tri 28604 35999 28605 36000 ne
rect 28605 35999 32719 36000
rect 24848 35707 28313 35999
tri 28313 35707 28605 35999 sw
tri 28605 35707 28897 35999 ne
rect 28897 35847 32719 35999
tri 32719 35847 33001 36129 sw
tri 33001 35847 33283 36129 ne
rect 33283 35847 37245 36129
rect 28897 35846 33001 35847
tri 33001 35846 33002 35847 sw
tri 33283 35846 33284 35847 ne
rect 33284 35846 37245 35847
rect 28897 35707 33002 35846
rect 24848 35706 28605 35707
tri 28605 35706 28606 35707 sw
tri 28897 35706 28898 35707 ne
rect 28898 35706 33002 35707
rect 24848 35414 28606 35706
tri 28606 35414 28898 35706 sw
tri 28898 35414 29190 35706 ne
rect 29190 35564 33002 35706
tri 33002 35564 33284 35846 sw
tri 33284 35564 33566 35846 ne
rect 33566 35832 37245 35846
tri 37245 35832 37542 36129 sw
tri 37542 35832 37839 36129 ne
rect 37839 35922 39440 36129
tri 39440 35922 39729 36211 sw
tri 39729 35922 40018 36211 ne
rect 40018 36209 41421 36211
tri 41421 36209 41711 36499 sw
tri 41711 36209 42001 36499 ne
rect 42001 36359 45801 36499
tri 45801 36359 46095 36653 sw
tri 46095 36359 46389 36653 ne
rect 46389 36377 50327 36653
tri 50327 36377 50615 36665 sw
tri 50615 36377 50903 36665 ne
rect 50903 36500 54727 36665
tri 54727 36500 55024 36797 sw
tri 55024 36500 55321 36797 ne
rect 55321 36500 71000 36797
rect 50903 36499 55024 36500
tri 55024 36499 55025 36500 sw
tri 55321 36499 55322 36500 ne
rect 55322 36499 71000 36500
rect 50903 36377 55025 36499
rect 46389 36359 50615 36377
rect 42001 36358 46095 36359
tri 46095 36358 46096 36359 sw
tri 46389 36358 46390 36359 ne
rect 46390 36358 50615 36359
rect 42001 36209 46096 36358
rect 40018 35922 41711 36209
rect 37839 35832 39729 35922
rect 33566 35831 37542 35832
tri 37542 35831 37543 35832 sw
tri 37839 35831 37840 35832 ne
rect 37840 35831 39729 35832
rect 33566 35564 37543 35831
rect 29190 35563 33284 35564
tri 33284 35563 33285 35564 sw
tri 33566 35563 33567 35564 ne
rect 33567 35563 37543 35564
rect 29190 35414 33285 35563
rect 24848 35220 28898 35414
tri 28898 35220 29092 35414 sw
tri 29190 35220 29384 35414 ne
rect 29384 35281 33285 35414
tri 33285 35281 33567 35563 sw
tri 33567 35281 33849 35563 ne
rect 33849 35534 37543 35563
tri 37543 35534 37840 35831 sw
tri 37840 35534 38137 35831 ne
rect 38137 35767 39729 35831
tri 39729 35767 39884 35922 sw
tri 40018 35767 40173 35922 ne
rect 40173 35919 41711 35922
tri 41711 35919 42001 36209 sw
tri 42001 35919 42291 36209 ne
rect 42291 36064 46096 36209
tri 46096 36064 46390 36358 sw
tri 46390 36064 46684 36358 ne
rect 46684 36201 50615 36358
tri 50615 36201 50791 36377 sw
tri 50903 36201 51079 36377 ne
rect 51079 36202 55025 36377
tri 55025 36202 55322 36499 sw
tri 55322 36400 55421 36499 ne
rect 55421 36400 71000 36499
rect 51079 36201 55322 36202
rect 46684 36064 50791 36201
rect 42291 36063 46390 36064
tri 46390 36063 46391 36064 sw
tri 46684 36063 46685 36064 ne
rect 46685 36063 50791 36064
rect 42291 35919 46391 36063
rect 40173 35918 42001 35919
tri 42001 35918 42002 35919 sw
tri 42291 35918 42292 35919 ne
rect 42292 35918 46391 35919
rect 40173 35767 42002 35918
rect 38137 35534 39884 35767
rect 33849 35281 37840 35534
rect 29384 35279 33567 35281
tri 33567 35279 33569 35281 sw
tri 33849 35279 33851 35281 ne
rect 33851 35279 37840 35281
rect 29384 35220 33569 35279
tri 24848 30976 29092 35220 ne
tri 29092 34928 29384 35220 sw
tri 29384 34928 29676 35220 ne
rect 29676 34997 33569 35220
tri 33569 34997 33851 35279 sw
tri 33851 34997 34133 35279 ne
rect 34133 35237 37840 35279
tri 37840 35237 38137 35534 sw
tri 38137 35237 38434 35534 ne
rect 38434 35478 39884 35534
tri 39884 35478 40173 35767 sw
tri 40173 35478 40462 35767 ne
rect 40462 35628 42002 35767
tri 42002 35628 42292 35918 sw
tri 42292 35628 42582 35918 ne
rect 42582 35769 46391 35918
tri 46391 35769 46685 36063 sw
tri 46685 35769 46979 36063 ne
rect 46979 35913 50791 36063
tri 50791 35913 51079 36201 sw
tri 51079 35913 51367 36201 ne
rect 51367 36200 55322 36201
tri 55322 36200 55324 36202 sw
rect 51367 35913 71000 36200
rect 46979 35911 51079 35913
tri 51079 35911 51081 35913 sw
tri 51367 35911 51369 35913 ne
rect 51369 35911 71000 35913
rect 46979 35769 51081 35911
rect 42582 35767 46685 35769
tri 46685 35767 46687 35769 sw
tri 46979 35767 46981 35769 ne
rect 46981 35767 51081 35769
rect 42582 35628 46687 35767
rect 40462 35478 42292 35628
rect 38434 35237 40173 35478
rect 34133 34997 38137 35237
rect 29676 34996 33851 34997
tri 33851 34996 33852 34997 sw
tri 34133 34996 34134 34997 ne
rect 34134 34996 38137 34997
rect 29676 34928 33852 34996
rect 29092 34851 29384 34928
tri 29384 34851 29461 34928 sw
tri 29676 34851 29753 34928 ne
rect 29753 34851 33852 34928
rect 29092 34559 29461 34851
tri 29461 34559 29753 34851 sw
tri 29753 34559 30045 34851 ne
rect 30045 34714 33852 34851
tri 33852 34714 34134 34996 sw
tri 34134 34714 34416 34996 ne
rect 34416 34940 38137 34996
tri 38137 34940 38434 35237 sw
tri 38434 34940 38731 35237 ne
rect 38731 35189 40173 35237
tri 40173 35189 40462 35478 sw
tri 40462 35189 40751 35478 ne
rect 40751 35392 42292 35478
tri 42292 35392 42528 35628 sw
tri 42582 35392 42818 35628 ne
rect 42818 35474 46687 35628
tri 46687 35474 46980 35767 sw
tri 46981 35474 47274 35767 ne
rect 47274 35623 51081 35767
tri 51081 35623 51369 35911 sw
tri 51369 35623 51657 35911 ne
rect 51657 35623 71000 35911
rect 47274 35622 51369 35623
tri 51369 35622 51370 35623 sw
tri 51657 35622 51658 35623 ne
rect 51658 35622 71000 35623
rect 47274 35474 51370 35622
rect 42818 35392 46980 35474
rect 40751 35288 42528 35392
tri 42528 35288 42632 35392 sw
tri 42818 35288 42922 35392 ne
rect 42922 35288 46980 35392
rect 40751 35189 42632 35288
rect 38731 34940 40462 35189
rect 34416 34901 38434 34940
tri 38434 34901 38473 34940 sw
tri 38731 34901 38770 34940 ne
rect 38770 34901 40462 34940
rect 34416 34714 38473 34901
rect 30045 34713 34134 34714
tri 34134 34713 34135 34714 sw
tri 34416 34713 34417 34714 ne
rect 34417 34713 38473 34714
rect 30045 34559 34135 34713
rect 29092 34558 29753 34559
tri 29753 34558 29754 34559 sw
tri 30045 34558 30046 34559 ne
rect 30046 34558 34135 34559
rect 29092 34266 29754 34558
tri 29754 34266 30046 34558 sw
tri 30046 34266 30338 34558 ne
rect 30338 34431 34135 34558
tri 34135 34431 34417 34713 sw
tri 34417 34431 34699 34713 ne
rect 34699 34604 38473 34713
tri 38473 34604 38770 34901 sw
tri 38770 34604 39067 34901 ne
rect 39067 34900 40462 34901
tri 40462 34900 40751 35189 sw
tri 40751 34900 41040 35189 ne
rect 41040 34998 42632 35189
tri 42632 34998 42922 35288 sw
tri 42922 34998 43212 35288 ne
rect 43212 35224 46980 35288
tri 46980 35224 47230 35474 sw
tri 47274 35224 47524 35474 ne
rect 47524 35334 51370 35474
tri 51370 35334 51658 35622 sw
tri 51658 35334 51946 35622 ne
rect 51946 35334 71000 35622
rect 47524 35333 51658 35334
tri 51658 35333 51659 35334 sw
tri 51946 35333 51947 35334 ne
rect 51947 35333 71000 35334
rect 47524 35224 51659 35333
rect 43212 34998 47230 35224
rect 41040 34900 42922 34998
rect 39067 34611 40751 34900
tri 40751 34611 41040 34900 sw
tri 41040 34611 41329 34900 ne
rect 41329 34810 42922 34900
tri 42922 34810 43110 34998 sw
tri 43212 34810 43400 34998 ne
rect 43400 34994 47230 34998
tri 47230 34994 47460 35224 sw
tri 47524 34994 47754 35224 ne
rect 47754 35045 51659 35224
tri 51659 35045 51947 35333 sw
tri 51947 35045 52235 35333 ne
rect 52235 35045 71000 35333
rect 47754 35044 51947 35045
tri 51947 35044 51948 35045 sw
tri 52235 35044 52236 35045 ne
rect 52236 35044 71000 35045
rect 47754 34994 51948 35044
rect 43400 34929 47460 34994
tri 47460 34929 47525 34994 sw
tri 47754 34929 47819 34994 ne
rect 47819 34929 51948 34994
rect 43400 34810 47525 34929
rect 41329 34611 43110 34810
rect 39067 34604 41040 34611
rect 34699 34603 38770 34604
tri 38770 34603 38771 34604 sw
tri 39067 34603 39068 34604 ne
rect 39068 34603 41040 34604
rect 34699 34431 38771 34603
rect 30338 34266 34417 34431
rect 29092 34265 30046 34266
tri 30046 34265 30047 34266 sw
tri 30338 34265 30339 34266 ne
rect 30339 34265 34417 34266
rect 29092 33973 30047 34265
tri 30047 33973 30339 34265 sw
tri 30339 33973 30631 34265 ne
rect 30631 34176 34417 34265
tri 34417 34176 34672 34431 sw
tri 34699 34176 34954 34431 ne
rect 34954 34306 38771 34431
tri 38771 34306 39068 34603 sw
tri 39068 34306 39365 34603 ne
rect 39365 34520 41040 34603
tri 41040 34520 41131 34611 sw
tri 41329 34520 41420 34611 ne
rect 41420 34520 43110 34611
tri 43110 34520 43400 34810 sw
tri 43400 34520 43690 34810 ne
rect 43690 34635 47525 34810
tri 47525 34635 47819 34929 sw
tri 47819 34635 48113 34929 ne
rect 48113 34756 51948 34929
tri 51948 34756 52236 35044 sw
tri 52236 34756 52524 35044 ne
rect 52524 34756 71000 35044
rect 48113 34755 52236 34756
tri 52236 34755 52237 34756 sw
tri 52524 34755 52525 34756 ne
rect 52525 34755 71000 34756
rect 48113 34635 52237 34755
rect 43690 34634 47819 34635
tri 47819 34634 47820 34635 sw
tri 48113 34634 48114 34635 ne
rect 48114 34634 52237 34635
rect 43690 34520 47820 34634
rect 39365 34306 41131 34520
rect 34954 34305 39068 34306
tri 39068 34305 39069 34306 sw
tri 39365 34305 39366 34306 ne
rect 39366 34305 41131 34306
rect 34954 34176 39069 34305
rect 30631 33973 34672 34176
rect 29092 33884 30339 33973
tri 30339 33884 30428 33973 sw
tri 30631 33884 30720 33973 ne
rect 30720 33894 34672 33973
tri 34672 33894 34954 34176 sw
tri 34954 33894 35236 34176 ne
rect 35236 34008 39069 34176
tri 39069 34008 39366 34305 sw
tri 39366 34008 39663 34305 ne
rect 39663 34231 41131 34305
tri 41131 34231 41420 34520 sw
tri 41420 34231 41709 34520 ne
rect 41709 34519 43400 34520
tri 43400 34519 43401 34520 sw
tri 43690 34519 43691 34520 ne
rect 43691 34519 47820 34520
rect 41709 34231 43401 34519
rect 39663 34008 41420 34231
rect 35236 33894 39366 34008
rect 30720 33884 34954 33894
rect 29092 33592 30428 33884
tri 30428 33592 30720 33884 sw
tri 30720 33592 31012 33884 ne
rect 31012 33779 34954 33884
tri 34954 33779 35069 33894 sw
tri 35236 33779 35351 33894 ne
rect 35351 33779 39366 33894
rect 31012 33592 35069 33779
rect 29092 33385 30720 33592
tri 30720 33385 30927 33592 sw
tri 31012 33385 31219 33592 ne
rect 31219 33497 35069 33592
tri 35069 33497 35351 33779 sw
tri 35351 33497 35633 33779 ne
rect 35633 33711 39366 33779
tri 39366 33711 39663 34008 sw
tri 39663 33711 39960 34008 ne
rect 39960 33942 41420 34008
tri 41420 33942 41709 34231 sw
tri 41709 33942 41998 34231 ne
rect 41998 34229 43401 34231
tri 43401 34229 43691 34519 sw
tri 43691 34229 43981 34519 ne
rect 43981 34340 47820 34519
tri 47820 34340 48114 34634 sw
tri 48114 34340 48408 34634 ne
rect 48408 34467 52237 34634
tri 52237 34467 52525 34755 sw
tri 52525 34467 52813 34755 ne
rect 52813 34467 71000 34755
rect 48408 34340 52525 34467
rect 43981 34339 48114 34340
tri 48114 34339 48115 34340 sw
tri 48408 34339 48409 34340 ne
rect 48409 34339 52525 34340
rect 43981 34229 48115 34339
rect 41998 34042 43691 34229
tri 43691 34042 43878 34229 sw
tri 43981 34042 44168 34229 ne
rect 44168 34045 48115 34229
tri 48115 34045 48409 34339 sw
tri 48409 34045 48703 34339 ne
rect 48703 34244 52525 34339
tri 52525 34244 52748 34467 sw
tri 52813 34244 53036 34467 ne
rect 53036 34244 71000 34467
rect 48703 34045 52748 34244
rect 44168 34042 48409 34045
rect 41998 33942 43878 34042
rect 39960 33787 41709 33942
tri 41709 33787 41864 33942 sw
tri 41998 33787 42153 33942 ne
rect 42153 33787 43878 33942
rect 39960 33711 41864 33787
rect 35633 33516 39663 33711
tri 39663 33516 39858 33711 sw
tri 39960 33516 40155 33711 ne
rect 40155 33516 41864 33711
rect 35633 33497 39858 33516
rect 31219 33495 35351 33497
tri 35351 33495 35353 33497 sw
tri 35633 33495 35635 33497 ne
rect 35635 33495 39858 33497
rect 31219 33385 35353 33495
rect 29092 33094 30927 33385
tri 30927 33094 31218 33385 sw
tri 31219 33094 31510 33385 ne
rect 31510 33213 35353 33385
tri 35353 33213 35635 33495 sw
tri 35635 33213 35917 33495 ne
rect 35917 33219 39858 33495
tri 39858 33219 40155 33516 sw
tri 40155 33219 40452 33516 ne
rect 40452 33498 41864 33516
tri 41864 33498 42153 33787 sw
tri 42153 33498 42442 33787 ne
rect 42442 33752 43878 33787
tri 43878 33752 44168 34042 sw
tri 44168 33752 44458 34042 ne
rect 44458 33950 48409 34042
tri 48409 33950 48504 34045 sw
tri 48703 33950 48798 34045 ne
rect 48798 33956 52748 34045
tri 52748 33956 53036 34244 sw
tri 53036 33956 53324 34244 ne
rect 53324 33956 71000 34244
rect 48798 33950 53036 33956
rect 44458 33752 48504 33950
rect 42442 33498 44168 33752
rect 40452 33219 42153 33498
rect 35917 33213 40155 33219
rect 31510 33212 35635 33213
tri 35635 33212 35636 33213 sw
tri 35917 33212 35918 33213 ne
rect 35918 33212 40155 33213
rect 31510 33094 35636 33212
rect 29092 32929 31218 33094
tri 31218 32929 31383 33094 sw
tri 31510 32929 31675 33094 ne
rect 31675 32930 35636 33094
tri 35636 32930 35918 33212 sw
tri 35918 32930 36200 33212 ne
rect 36200 32930 40155 33212
rect 31675 32929 35918 32930
rect 29092 32637 31383 32929
tri 31383 32637 31675 32929 sw
tri 31675 32637 31967 32929 ne
rect 31967 32850 35918 32929
tri 35918 32850 35998 32930 sw
tri 36200 32850 36280 32930 ne
rect 36280 32922 40155 32930
tri 40155 32922 40452 33219 sw
tri 40452 32922 40749 33219 ne
rect 40749 33209 42153 33219
tri 42153 33209 42442 33498 sw
tri 42442 33209 42731 33498 ne
rect 42731 33462 44168 33498
tri 44168 33462 44458 33752 sw
tri 44458 33462 44748 33752 ne
rect 44748 33656 48504 33752
tri 48504 33656 48798 33950 sw
tri 48798 33656 49092 33950 ne
rect 49092 33868 53036 33950
tri 53036 33868 53124 33956 sw
tri 53324 33868 53412 33956 ne
rect 53412 33868 71000 33956
rect 49092 33656 53124 33868
rect 44748 33462 48798 33656
rect 42731 33411 44458 33462
tri 44458 33411 44509 33462 sw
tri 44748 33411 44799 33462 ne
rect 44799 33453 48798 33462
tri 48798 33453 49001 33656 sw
tri 49092 33453 49295 33656 ne
rect 49295 33580 53124 33656
tri 53124 33580 53412 33868 sw
tri 53412 33580 53700 33868 ne
rect 53700 33580 71000 33868
rect 49295 33579 53412 33580
tri 53412 33579 53413 33580 sw
tri 53700 33579 53701 33580 ne
rect 53701 33579 71000 33580
rect 49295 33453 53413 33579
rect 44799 33411 49001 33453
rect 42731 33209 44509 33411
rect 40749 32922 42442 33209
rect 36280 32920 40452 32922
tri 40452 32920 40454 32922 sw
tri 40749 32920 40751 32922 ne
rect 40751 32920 42442 32922
tri 42442 32920 42731 33209 sw
tri 42731 32920 43020 33209 ne
rect 43020 33121 44509 33209
tri 44509 33121 44799 33411 sw
tri 44799 33121 45089 33411 ne
rect 45089 33159 49001 33411
tri 49001 33159 49295 33453 sw
tri 49295 33159 49589 33453 ne
rect 49589 33291 53413 33453
tri 53413 33291 53701 33579 sw
tri 53701 33291 53989 33579 ne
rect 53989 33291 71000 33579
rect 49589 33290 53701 33291
tri 53701 33290 53702 33291 sw
tri 53989 33290 53990 33291 ne
rect 53990 33290 71000 33291
rect 49589 33159 53702 33290
rect 45089 33121 49295 33159
rect 43020 32920 44799 33121
rect 36280 32850 40454 32920
rect 31967 32637 35998 32850
rect 29092 32636 31675 32637
tri 31675 32636 31676 32637 sw
tri 31967 32636 31968 32637 ne
rect 31968 32636 35998 32637
rect 29092 32344 31676 32636
tri 31676 32344 31968 32636 sw
tri 31968 32344 32260 32636 ne
rect 32260 32568 35998 32636
tri 35998 32568 36280 32850 sw
tri 36280 32568 36562 32850 ne
rect 36562 32623 40454 32850
tri 40454 32623 40751 32920 sw
tri 40751 32623 41048 32920 ne
rect 41048 32631 42731 32920
tri 42731 32631 43020 32920 sw
tri 43020 32631 43309 32920 ne
rect 43309 32831 44799 32920
tri 44799 32831 45089 33121 sw
tri 45089 32831 45379 33121 ne
rect 45379 33001 49295 33121
tri 49295 33001 49453 33159 sw
tri 49589 33001 49747 33159 ne
rect 49747 33002 53702 33159
tri 53702 33002 53990 33290 sw
tri 53990 33200 54080 33290 ne
rect 54080 33200 71000 33290
rect 49747 33001 53990 33002
rect 45379 32831 49453 33001
rect 43309 32830 45089 32831
tri 45089 32830 45090 32831 sw
tri 45379 32830 45380 32831 ne
rect 45380 32830 49453 32831
rect 43309 32631 45090 32830
rect 41048 32623 43020 32631
rect 36562 32568 40751 32623
rect 32260 32363 36280 32568
tri 36280 32363 36485 32568 sw
tri 36562 32363 36767 32568 ne
rect 36767 32363 40751 32568
rect 32260 32344 36485 32363
rect 29092 32343 31968 32344
tri 31968 32343 31969 32344 sw
tri 32260 32343 32261 32344 ne
rect 32261 32343 36485 32344
rect 29092 32051 31969 32343
tri 31969 32051 32261 32343 sw
tri 32261 32051 32553 32343 ne
rect 32553 32081 36485 32343
tri 36485 32081 36767 32363 sw
tri 36767 32081 37049 32363 ne
rect 37049 32326 40751 32363
tri 40751 32326 41048 32623 sw
tri 41048 32326 41345 32623 ne
rect 41345 32540 43020 32623
tri 43020 32540 43111 32631 sw
tri 43309 32540 43400 32631 ne
rect 43400 32540 45090 32631
tri 45090 32540 45380 32830 sw
tri 45380 32540 45670 32830 ne
rect 45670 32707 49453 32830
tri 49453 32707 49747 33001 sw
tri 49747 32707 50041 33001 ne
rect 50041 33000 53990 33001
tri 53990 33000 53992 33002 sw
rect 50041 32707 71000 33000
rect 45670 32705 49747 32707
tri 49747 32705 49749 32707 sw
tri 50041 32705 50043 32707 ne
rect 50043 32705 71000 32707
rect 45670 32540 49749 32705
rect 41345 32326 43111 32540
rect 37049 32184 41048 32326
tri 41048 32184 41190 32326 sw
tri 41345 32184 41487 32326 ne
rect 41487 32251 43111 32326
tri 43111 32251 43400 32540 sw
tri 43400 32251 43689 32540 ne
rect 43689 32539 45380 32540
tri 45380 32539 45381 32540 sw
tri 45670 32539 45671 32540 ne
rect 45671 32539 49749 32540
rect 43689 32251 45381 32539
rect 41487 32184 43400 32251
rect 37049 32081 41190 32184
rect 32553 32051 36767 32081
rect 29092 32049 32261 32051
tri 32261 32049 32263 32051 sw
tri 32553 32049 32555 32051 ne
rect 32555 32049 36767 32051
rect 29092 31757 32263 32049
tri 32263 31757 32555 32049 sw
tri 32555 31757 32847 32049 ne
rect 32847 31886 36767 32049
tri 36767 31886 36962 32081 sw
tri 37049 31886 37244 32081 ne
rect 37244 31887 41190 32081
tri 41190 31887 41487 32184 sw
tri 41487 31887 41784 32184 ne
rect 41784 31962 43400 32184
tri 43400 31962 43689 32251 sw
tri 43689 31962 43978 32251 ne
rect 43978 32249 45381 32251
tri 45381 32249 45671 32539 sw
tri 45671 32249 45961 32539 ne
rect 45961 32411 49749 32539
tri 49749 32411 50043 32705 sw
tri 50043 32411 50337 32705 ne
rect 50337 32411 71000 32705
rect 45961 32410 50043 32411
tri 50043 32410 50044 32411 sw
tri 50337 32410 50338 32411 ne
rect 50338 32410 71000 32411
rect 45961 32249 50044 32410
rect 43978 31962 45671 32249
rect 41784 31887 43689 31962
rect 37244 31886 41487 31887
tri 41487 31886 41488 31887 sw
tri 41784 31886 41785 31887 ne
rect 41785 31886 43689 31887
rect 32847 31757 36962 31886
rect 29092 31756 32555 31757
tri 32555 31756 32556 31757 sw
tri 32847 31756 32848 31757 ne
rect 32848 31756 36962 31757
rect 29092 31464 32556 31756
tri 32556 31464 32848 31756 sw
tri 32848 31464 33140 31756 ne
rect 33140 31604 36962 31756
tri 36962 31604 37244 31886 sw
tri 37244 31604 37526 31886 ne
rect 37526 31604 41488 31886
rect 33140 31603 37244 31604
tri 37244 31603 37245 31604 sw
tri 37526 31603 37527 31604 ne
rect 37527 31603 41488 31604
rect 33140 31464 37245 31603
rect 29092 31463 32848 31464
tri 32848 31463 32849 31464 sw
tri 33140 31463 33141 31464 ne
rect 33141 31463 37245 31464
rect 29092 31171 32849 31463
tri 32849 31171 33141 31463 sw
tri 33141 31171 33433 31463 ne
rect 33433 31321 37245 31463
tri 37245 31321 37527 31603 sw
tri 37527 31321 37809 31603 ne
rect 37809 31589 41488 31603
tri 41488 31589 41785 31886 sw
tri 41785 31589 42082 31886 ne
rect 42082 31807 43689 31886
tri 43689 31807 43844 31962 sw
tri 43978 31807 44133 31962 ne
rect 44133 31959 45671 31962
tri 45671 31959 45961 32249 sw
tri 45961 31959 46251 32249 ne
rect 46251 32116 50044 32249
tri 50044 32116 50338 32410 sw
tri 50338 32116 50632 32410 ne
rect 50632 32116 71000 32410
rect 46251 32115 50338 32116
tri 50338 32115 50339 32116 sw
tri 50632 32115 50633 32116 ne
rect 50633 32115 71000 32116
rect 46251 31959 50339 32115
rect 44133 31958 45961 31959
tri 45961 31958 45962 31959 sw
tri 46251 31958 46252 31959 ne
rect 46252 31958 50339 31959
rect 44133 31807 45962 31958
rect 42082 31589 43844 31807
rect 37809 31321 41785 31589
rect 33433 31320 37527 31321
tri 37527 31320 37528 31321 sw
tri 37809 31320 37810 31321 ne
rect 37810 31320 41785 31321
rect 33433 31171 37528 31320
rect 29092 30976 33141 31171
tri 33141 30976 33336 31171 sw
tri 33433 30976 33628 31171 ne
rect 33628 31038 37528 31171
tri 37528 31038 37810 31320 sw
tri 37810 31038 38092 31320 ne
rect 38092 31292 41785 31320
tri 41785 31292 42082 31589 sw
tri 42082 31292 42379 31589 ne
rect 42379 31518 43844 31589
tri 43844 31518 44133 31807 sw
tri 44133 31518 44422 31807 ne
rect 44422 31668 45962 31807
tri 45962 31668 46252 31958 sw
tri 46252 31668 46542 31958 ne
rect 46542 31821 50339 31958
tri 50339 31821 50633 32115 sw
tri 50633 31821 50927 32115 ne
rect 50927 31821 71000 32115
rect 46542 31820 50633 31821
tri 50633 31820 50634 31821 sw
tri 50927 31820 50928 31821 ne
rect 50928 31820 71000 31821
rect 46542 31668 50634 31820
rect 44422 31518 46252 31668
rect 42379 31292 44133 31518
rect 38092 31291 42082 31292
tri 42082 31291 42083 31292 sw
tri 42379 31291 42380 31292 ne
rect 42380 31291 44133 31292
rect 38092 31038 42083 31291
rect 33628 31037 37810 31038
tri 37810 31037 37811 31038 sw
tri 38092 31037 38093 31038 ne
rect 38093 31037 42083 31038
rect 33628 30976 37811 31037
tri 29092 26732 33336 30976 ne
tri 33336 30684 33628 30976 sw
tri 33628 30684 33920 30976 ne
rect 33920 30755 37811 30976
tri 37811 30755 38093 31037 sw
tri 38093 30755 38375 31037 ne
rect 38375 30994 42083 31037
tri 42083 30994 42380 31291 sw
tri 42380 30994 42677 31291 ne
rect 42677 31229 44133 31291
tri 44133 31229 44422 31518 sw
tri 44422 31229 44711 31518 ne
rect 44711 31431 46252 31518
tri 46252 31431 46489 31668 sw
tri 46542 31431 46779 31668 ne
rect 46779 31526 50634 31668
tri 50634 31526 50928 31820 sw
tri 50928 31526 51222 31820 ne
rect 51222 31526 71000 31820
rect 46779 31525 50928 31526
tri 50928 31525 50929 31526 sw
tri 51222 31525 51223 31526 ne
rect 51223 31525 71000 31526
rect 46779 31431 50929 31525
rect 44711 31229 46489 31431
rect 42677 30994 44422 31229
rect 38375 30940 42380 30994
tri 42380 30940 42434 30994 sw
tri 42677 30940 42731 30994 ne
rect 42731 30940 44422 30994
tri 44422 30940 44711 31229 sw
tri 44711 30940 45000 31229 ne
rect 45000 31141 46489 31229
tri 46489 31141 46779 31431 sw
tri 46779 31141 47069 31431 ne
rect 47069 31231 50929 31431
tri 50929 31231 51223 31525 sw
tri 51223 31231 51517 31525 ne
rect 51517 31231 71000 31525
rect 47069 31141 51223 31231
rect 45000 31044 46779 31141
tri 46779 31044 46876 31141 sw
tri 47069 31044 47166 31141 ne
rect 47166 31044 51223 31141
rect 45000 30940 46876 31044
rect 38375 30755 42434 30940
rect 33920 30753 38093 30755
tri 38093 30753 38095 30755 sw
tri 38375 30753 38377 30755 ne
rect 38377 30753 42434 30755
rect 33920 30684 38095 30753
rect 33336 30609 33628 30684
tri 33628 30609 33703 30684 sw
tri 33920 30609 33995 30684 ne
rect 33995 30609 38095 30684
rect 33336 30317 33703 30609
tri 33703 30317 33995 30609 sw
tri 33995 30317 34287 30609 ne
rect 34287 30471 38095 30609
tri 38095 30471 38377 30753 sw
tri 38377 30471 38659 30753 ne
rect 38659 30643 42434 30753
tri 42434 30643 42731 30940 sw
tri 42731 30643 43028 30940 ne
rect 43028 30651 44711 30940
tri 44711 30651 45000 30940 sw
tri 45000 30651 45289 30940 ne
rect 45289 30754 46876 30940
tri 46876 30754 47166 31044 sw
tri 47166 30754 47456 31044 ne
rect 47456 30981 51223 31044
tri 51223 30981 51473 31231 sw
tri 51517 30981 51767 31231 ne
rect 51767 30981 71000 31231
rect 47456 30754 51473 30981
rect 45289 30651 47166 30754
rect 43028 30643 45000 30651
rect 38659 30471 42731 30643
rect 34287 30317 38377 30471
rect 33336 30315 33995 30317
tri 33995 30315 33997 30317 sw
tri 34287 30315 34289 30317 ne
rect 34289 30315 38377 30317
rect 33336 30023 33997 30315
tri 33997 30023 34289 30315 sw
tri 34289 30023 34581 30315 ne
rect 34581 30189 38377 30315
tri 38377 30189 38659 30471 sw
tri 38659 30189 38941 30471 ne
rect 38941 30346 42731 30471
tri 42731 30346 43028 30643 sw
tri 43028 30346 43325 30643 ne
rect 43325 30560 45000 30643
tri 45000 30560 45091 30651 sw
tri 45289 30560 45380 30651 ne
rect 45380 30560 47166 30651
rect 43325 30346 45091 30560
rect 38941 30345 43028 30346
tri 43028 30345 43029 30346 sw
tri 43325 30345 43326 30346 ne
rect 43326 30345 45091 30346
rect 38941 30189 43029 30345
rect 34581 30023 38659 30189
rect 33336 30022 34289 30023
tri 34289 30022 34290 30023 sw
tri 34581 30022 34582 30023 ne
rect 34582 30022 38659 30023
rect 33336 29730 34290 30022
tri 34290 29730 34582 30022 sw
tri 34582 29730 34874 30022 ne
rect 34874 29932 38659 30022
tri 38659 29932 38916 30189 sw
tri 38941 29932 39198 30189 ne
rect 39198 30048 43029 30189
tri 43029 30048 43326 30345 sw
tri 43326 30048 43623 30345 ne
rect 43623 30271 45091 30345
tri 45091 30271 45380 30560 sw
tri 45380 30271 45669 30560 ne
rect 45669 30559 47166 30560
tri 47166 30559 47361 30754 sw
tri 47456 30559 47651 30754 ne
rect 47651 30750 51473 30754
tri 51473 30750 51704 30981 sw
tri 51767 30750 51998 30981 ne
rect 51998 30750 71000 30981
rect 47651 30686 51704 30750
tri 51704 30686 51768 30750 sw
tri 51998 30686 52062 30750 ne
rect 52062 30686 71000 30750
rect 47651 30559 51768 30686
rect 45669 30271 47361 30559
rect 43623 30048 45380 30271
rect 39198 29932 43326 30048
rect 34874 29730 38916 29932
rect 33336 29640 34582 29730
tri 34582 29640 34672 29730 sw
tri 34874 29640 34964 29730 ne
rect 34964 29650 38916 29730
tri 38916 29650 39198 29932 sw
tri 39198 29650 39480 29932 ne
rect 39480 29751 43326 29932
tri 43326 29751 43623 30048 sw
tri 43623 29751 43920 30048 ne
rect 43920 29982 45380 30048
tri 45380 29982 45669 30271 sw
tri 45669 29982 45958 30271 ne
rect 45958 30269 47361 30271
tri 47361 30269 47651 30559 sw
tri 47651 30269 47941 30559 ne
rect 47941 30392 51768 30559
tri 51768 30392 52062 30686 sw
tri 52062 30392 52356 30686 ne
rect 52356 30392 71000 30686
rect 47941 30391 52062 30392
tri 52062 30391 52063 30392 sw
tri 52356 30391 52357 30392 ne
rect 52357 30391 71000 30392
rect 47941 30269 52063 30391
rect 45958 30090 47651 30269
tri 47651 30090 47830 30269 sw
tri 47941 30090 48120 30269 ne
rect 48120 30097 52063 30269
tri 52063 30097 52357 30391 sw
tri 52357 30097 52651 30391 ne
rect 52651 30097 71000 30391
rect 48120 30096 52357 30097
tri 52357 30096 52358 30097 sw
tri 52651 30096 52652 30097 ne
rect 52652 30096 71000 30097
rect 48120 30090 52358 30096
rect 45958 29982 47830 30090
rect 43920 29827 45669 29982
tri 45669 29827 45824 29982 sw
tri 45958 29827 46113 29982 ne
rect 46113 29827 47830 29982
rect 43920 29751 45824 29827
rect 39480 29650 43623 29751
rect 34964 29640 39198 29650
rect 33336 29348 34672 29640
tri 34672 29348 34964 29640 sw
tri 34964 29348 35256 29640 ne
rect 35256 29536 39198 29640
tri 39198 29536 39312 29650 sw
tri 39480 29536 39594 29650 ne
rect 39594 29556 43623 29650
tri 43623 29556 43818 29751 sw
tri 43920 29556 44115 29751 ne
rect 44115 29556 45824 29751
rect 39594 29536 43818 29556
rect 35256 29348 39312 29536
rect 33336 29143 34964 29348
tri 34964 29143 35169 29348 sw
tri 35256 29143 35461 29348 ne
rect 35461 29254 39312 29348
tri 39312 29254 39594 29536 sw
tri 39594 29254 39876 29536 ne
rect 39876 29259 43818 29536
tri 43818 29259 44115 29556 sw
tri 44115 29259 44412 29556 ne
rect 44412 29538 45824 29556
tri 45824 29538 46113 29827 sw
tri 46113 29538 46402 29827 ne
rect 46402 29800 47830 29827
tri 47830 29800 48120 30090 sw
tri 48120 29800 48410 30090 ne
rect 48410 29802 52358 30090
tri 52358 29802 52652 30096 sw
tri 52652 30000 52748 30096 ne
rect 52748 30000 71000 30096
rect 48410 29800 52652 29802
tri 52652 29800 52654 29802 sw
rect 46402 29799 48120 29800
tri 48120 29799 48121 29800 sw
tri 48410 29799 48411 29800 ne
rect 48411 29799 71000 29800
rect 46402 29538 48121 29799
rect 44412 29259 46113 29538
rect 39876 29258 44115 29259
tri 44115 29258 44116 29259 sw
tri 44412 29258 44413 29259 ne
rect 44413 29258 46113 29259
rect 39876 29254 44116 29258
rect 35461 29253 39594 29254
tri 39594 29253 39595 29254 sw
tri 39876 29253 39877 29254 ne
rect 39877 29253 44116 29254
rect 35461 29143 39595 29253
rect 33336 28851 35169 29143
tri 35169 28851 35461 29143 sw
tri 35461 28851 35753 29143 ne
rect 35753 28971 39595 29143
tri 39595 28971 39877 29253 sw
tri 39877 28971 40159 29253 ne
rect 40159 28971 44116 29253
rect 35753 28969 39877 28971
tri 39877 28969 39879 28971 sw
tri 40159 28969 40161 28971 ne
rect 40161 28969 44116 28971
rect 35753 28851 39879 28969
rect 33336 28686 35461 28851
tri 35461 28686 35626 28851 sw
tri 35753 28686 35918 28851 ne
rect 35918 28688 39879 28851
tri 39879 28688 40160 28969 sw
tri 40161 28688 40442 28969 ne
rect 40442 28961 44116 28969
tri 44116 28961 44413 29258 sw
tri 44413 28961 44710 29258 ne
rect 44710 29249 46113 29258
tri 46113 29249 46402 29538 sw
tri 46402 29249 46691 29538 ne
rect 46691 29509 48121 29538
tri 48121 29509 48411 29799 sw
tri 48411 29509 48701 29799 ne
rect 48701 29509 71000 29799
rect 46691 29249 48411 29509
rect 44710 28961 46402 29249
rect 40442 28688 44413 28961
rect 35918 28686 40160 28688
rect 33336 28394 35626 28686
tri 35626 28394 35918 28686 sw
tri 35918 28394 36210 28686 ne
rect 36210 28606 40160 28686
tri 40160 28606 40242 28688 sw
tri 40442 28606 40524 28688 ne
rect 40524 28664 44413 28688
tri 44413 28664 44710 28961 sw
tri 44710 28664 45007 28961 ne
rect 45007 28960 46402 28961
tri 46402 28960 46691 29249 sw
tri 46691 28960 46980 29249 ne
rect 46980 29219 48411 29249
tri 48411 29219 48701 29509 sw
tri 48701 29219 48991 29509 ne
rect 48991 29219 71000 29509
rect 46980 29161 48701 29219
tri 48701 29161 48759 29219 sw
tri 48991 29161 49049 29219 ne
rect 49049 29161 71000 29219
rect 46980 28960 48759 29161
rect 45007 28671 46691 28960
tri 46691 28671 46980 28960 sw
tri 46980 28671 47269 28960 ne
rect 47269 28871 48759 28960
tri 48759 28871 49049 29161 sw
tri 49049 28871 49339 29161 ne
rect 49339 28871 71000 29161
rect 47269 28870 49049 28871
tri 49049 28870 49050 28871 sw
tri 49339 28870 49340 28871 ne
rect 49340 28870 71000 28871
rect 47269 28671 49050 28870
rect 45007 28664 46980 28671
rect 40524 28662 44710 28664
tri 44710 28662 44712 28664 sw
tri 45007 28662 45009 28664 ne
rect 45009 28662 46980 28664
rect 40524 28606 44712 28662
rect 36210 28394 40242 28606
rect 33336 28393 35918 28394
tri 35918 28393 35919 28394 sw
tri 36210 28393 36211 28394 ne
rect 36211 28393 40242 28394
rect 33336 28101 35919 28393
tri 35919 28101 36211 28393 sw
tri 36211 28101 36503 28393 ne
rect 36503 28324 40242 28393
tri 40242 28324 40524 28606 sw
tri 40524 28324 40806 28606 ne
rect 40806 28365 44712 28606
tri 44712 28365 45009 28662 sw
tri 45009 28365 45306 28662 ne
rect 45306 28580 46980 28662
tri 46980 28580 47071 28671 sw
tri 47269 28580 47360 28671 ne
rect 47360 28580 49050 28671
tri 49050 28580 49340 28870 sw
tri 49340 28580 49630 28870 ne
rect 49630 28580 71000 28870
rect 45306 28365 47071 28580
rect 40806 28324 45009 28365
rect 36503 28120 40524 28324
tri 40524 28120 40728 28324 sw
tri 40806 28120 41010 28324 ne
rect 41010 28120 45009 28324
rect 36503 28101 40728 28120
rect 33336 28100 36211 28101
tri 36211 28100 36212 28101 sw
tri 36503 28100 36504 28101 ne
rect 36504 28100 40728 28101
rect 33336 27808 36212 28100
tri 36212 27808 36504 28100 sw
tri 36504 27808 36796 28100 ne
rect 36796 27838 40728 28100
tri 40728 27838 41010 28120 sw
tri 41010 27838 41292 28120 ne
rect 41292 28069 45009 28120
tri 45009 28069 45305 28365 sw
tri 45306 28069 45602 28365 ne
rect 45602 28291 47071 28365
tri 47071 28291 47360 28580 sw
tri 47360 28291 47649 28580 ne
rect 47649 28579 49340 28580
tri 49340 28579 49341 28580 sw
tri 49630 28579 49631 28580 ne
rect 49631 28579 71000 28580
rect 47649 28291 49341 28579
rect 45602 28069 47360 28291
rect 41292 27941 45305 28069
tri 45305 27941 45433 28069 sw
tri 45602 27941 45730 28069 ne
rect 45730 28002 47360 28069
tri 47360 28002 47649 28291 sw
tri 47649 28002 47938 28291 ne
rect 47938 28289 49341 28291
tri 49341 28289 49631 28579 sw
tri 49631 28289 49921 28579 ne
rect 49921 28289 71000 28579
rect 47938 28002 49631 28289
rect 45730 27941 47649 28002
rect 41292 27838 45433 27941
rect 36796 27808 41010 27838
rect 33336 27807 36504 27808
tri 36504 27807 36505 27808 sw
tri 36796 27807 36797 27808 ne
rect 36797 27807 41010 27808
rect 33336 27515 36505 27807
tri 36505 27515 36797 27807 sw
tri 36797 27515 37089 27807 ne
rect 37089 27643 41010 27807
tri 41010 27643 41205 27838 sw
tri 41292 27643 41487 27838 ne
rect 41487 27644 45433 27838
tri 45433 27644 45730 27941 sw
tri 45730 27644 46027 27941 ne
rect 46027 27847 47649 27941
tri 47649 27847 47804 28002 sw
tri 47938 27847 48093 28002 ne
rect 48093 27999 49631 28002
tri 49631 27999 49921 28289 sw
tri 49921 27999 50211 28289 ne
rect 50211 27999 71000 28289
rect 48093 27998 49921 27999
tri 49921 27998 49922 27999 sw
tri 50211 27998 50212 27999 ne
rect 50212 27998 71000 27999
rect 48093 27847 49922 27998
rect 46027 27644 47804 27847
rect 41487 27643 45730 27644
tri 45730 27643 45731 27644 sw
tri 46027 27643 46028 27644 ne
rect 46028 27643 47804 27644
rect 37089 27515 41205 27643
rect 33336 27513 36797 27515
tri 36797 27513 36799 27515 sw
tri 37089 27513 37091 27515 ne
rect 37091 27513 41205 27515
rect 33336 27221 36799 27513
tri 36799 27221 37091 27513 sw
tri 37091 27221 37383 27513 ne
rect 37383 27361 41205 27513
tri 41205 27361 41487 27643 sw
tri 41487 27361 41769 27643 ne
rect 41769 27361 45731 27643
rect 37383 27360 41487 27361
tri 41487 27360 41488 27361 sw
tri 41769 27360 41770 27361 ne
rect 41770 27360 45731 27361
rect 37383 27221 41488 27360
rect 33336 27220 37091 27221
tri 37091 27220 37092 27221 sw
tri 37383 27220 37384 27221 ne
rect 37384 27220 41488 27221
rect 33336 26928 37092 27220
tri 37092 26928 37384 27220 sw
tri 37384 26928 37676 27220 ne
rect 37676 27078 41488 27220
tri 41488 27078 41770 27360 sw
tri 41770 27078 42052 27360 ne
rect 42052 27346 45731 27360
tri 45731 27346 46028 27643 sw
tri 46028 27346 46325 27643 ne
rect 46325 27558 47804 27643
tri 47804 27558 48093 27847 sw
tri 48093 27558 48382 27847 ne
rect 48382 27708 49922 27847
tri 49922 27708 50212 27998 sw
tri 50212 27708 50502 27998 ne
rect 50502 27708 71000 27998
rect 48382 27558 50212 27708
rect 46325 27346 48093 27558
rect 42052 27078 46028 27346
rect 37676 27077 41770 27078
tri 41770 27077 41771 27078 sw
tri 42052 27077 42053 27078 ne
rect 42053 27077 46028 27078
rect 37676 26928 41771 27077
rect 33336 26732 37384 26928
tri 37384 26732 37580 26928 sw
tri 37676 26732 37872 26928 ne
rect 37872 26795 41771 26928
tri 41771 26795 42053 27077 sw
tri 42053 26795 42335 27077 ne
rect 42335 27049 46028 27077
tri 46028 27049 46325 27346 sw
tri 46325 27049 46622 27346 ne
rect 46622 27269 48093 27346
tri 48093 27269 48382 27558 sw
tri 48382 27269 48671 27558 ne
rect 48671 27471 50212 27558
tri 50212 27471 50449 27708 sw
tri 50502 27471 50739 27708 ne
rect 50739 27471 71000 27708
rect 48671 27269 50449 27471
rect 46622 27049 48382 27269
rect 42335 26981 46325 27049
tri 46325 26981 46393 27049 sw
tri 46622 26981 46690 27049 ne
rect 46690 26981 48382 27049
rect 42335 26795 46393 26981
rect 37872 26794 42053 26795
tri 42053 26794 42054 26795 sw
tri 42335 26794 42336 26795 ne
rect 42336 26794 46393 26795
rect 37872 26732 42054 26794
tri 33336 22488 37580 26732 ne
tri 37580 26440 37872 26732 sw
tri 37872 26440 38164 26732 ne
rect 38164 26512 42054 26732
tri 42054 26512 42336 26794 sw
tri 42336 26512 42618 26794 ne
rect 42618 26684 46393 26794
tri 46393 26684 46690 26981 sw
tri 46690 26684 46987 26981 ne
rect 46987 26980 48382 26981
tri 48382 26980 48671 27269 sw
tri 48671 26980 48960 27269 ne
rect 48960 27181 50449 27269
tri 50449 27181 50739 27471 sw
tri 50739 27181 51029 27471 ne
rect 51029 27181 71000 27471
rect 48960 26980 50739 27181
rect 46987 26691 48671 26980
tri 48671 26691 48960 26980 sw
tri 48960 26691 49249 26980 ne
rect 49249 26891 50739 26980
tri 50739 26891 51029 27181 sw
tri 51029 26891 51319 27181 ne
rect 51319 26891 71000 27181
rect 49249 26800 51029 26891
tri 51029 26800 51120 26891 sw
tri 51319 26800 51410 26891 ne
rect 51410 26800 71000 26891
rect 49249 26691 51120 26800
rect 46987 26684 48960 26691
rect 42618 26683 46690 26684
tri 46690 26683 46691 26684 sw
tri 46987 26683 46988 26684 ne
rect 46988 26683 48960 26684
rect 42618 26512 46691 26683
rect 38164 26511 42336 26512
tri 42336 26511 42337 26512 sw
tri 42618 26511 42619 26512 ne
rect 42619 26511 46691 26512
rect 38164 26440 42337 26511
rect 37580 26366 37872 26440
tri 37872 26366 37946 26440 sw
tri 38164 26366 38238 26440 ne
rect 38238 26366 42337 26440
rect 37580 26074 37946 26366
tri 37946 26074 38238 26366 sw
tri 38238 26074 38530 26366 ne
rect 38530 26229 42337 26366
tri 42337 26229 42619 26511 sw
tri 42619 26229 42901 26511 ne
rect 42901 26386 46691 26511
tri 46691 26386 46988 26683 sw
tri 46988 26386 47285 26683 ne
rect 47285 26600 48960 26683
tri 48960 26600 49051 26691 sw
tri 49249 26600 49340 26691 ne
rect 49340 26600 51120 26691
tri 51120 26600 51320 26800 sw
rect 47285 26386 49051 26600
rect 42901 26385 46988 26386
tri 46988 26385 46989 26386 sw
tri 47285 26385 47286 26386 ne
rect 47286 26385 49051 26386
rect 42901 26229 46989 26385
rect 38530 26227 42619 26229
tri 42619 26227 42621 26229 sw
tri 42901 26227 42903 26229 ne
rect 42903 26227 46989 26229
rect 38530 26074 42621 26227
rect 37580 26073 38238 26074
tri 38238 26073 38239 26074 sw
tri 38530 26073 38531 26074 ne
rect 38531 26073 42621 26074
rect 37580 25781 38239 26073
tri 38239 25781 38531 26073 sw
tri 38531 25781 38823 26073 ne
rect 38823 25946 42621 26073
tri 42621 25946 42902 26227 sw
tri 42903 25946 43184 26227 ne
rect 43184 26088 46989 26227
tri 46989 26088 47286 26385 sw
tri 47286 26088 47583 26385 ne
rect 47583 26311 49051 26385
tri 49051 26311 49340 26600 sw
tri 49340 26311 49629 26600 ne
rect 49629 26311 71000 26600
rect 47583 26088 49340 26311
rect 43184 25946 47286 26088
rect 38823 25781 42902 25946
rect 37580 25779 38531 25781
tri 38531 25779 38533 25781 sw
tri 38823 25779 38825 25781 ne
rect 38825 25779 42902 25781
rect 37580 25487 38533 25779
tri 38533 25487 38825 25779 sw
tri 38825 25487 39117 25779 ne
rect 39117 25688 42902 25779
tri 42902 25688 43160 25946 sw
tri 43184 25688 43442 25946 ne
rect 43442 25791 47286 25946
tri 47286 25791 47583 26088 sw
tri 47583 25791 47880 26088 ne
rect 47880 26022 49340 26088
tri 49340 26022 49629 26311 sw
tri 49629 26022 49918 26311 ne
rect 49918 26022 71000 26311
rect 47880 25867 49629 26022
tri 49629 25867 49784 26022 sw
tri 49918 25867 50073 26022 ne
rect 50073 25867 71000 26022
rect 47880 25791 49784 25867
rect 43442 25688 47583 25791
rect 39117 25487 43160 25688
rect 37580 25396 38825 25487
tri 38825 25396 38916 25487 sw
tri 39117 25396 39208 25487 ne
rect 39208 25406 43160 25487
tri 43160 25406 43442 25688 sw
tri 43442 25406 43724 25688 ne
rect 43724 25596 47583 25688
tri 47583 25596 47778 25791 sw
tri 47880 25596 48075 25791 ne
rect 48075 25596 49784 25791
rect 43724 25406 47778 25596
rect 39208 25396 43442 25406
rect 37580 25104 38916 25396
tri 38916 25104 39208 25396 sw
tri 39208 25104 39500 25396 ne
rect 39500 25293 43442 25396
tri 43442 25293 43555 25406 sw
tri 43724 25293 43837 25406 ne
rect 43837 25299 47778 25406
tri 47778 25299 48075 25596 sw
tri 48075 25299 48372 25596 ne
rect 48372 25578 49784 25596
tri 49784 25578 50073 25867 sw
tri 50073 25578 50362 25867 ne
rect 50362 25578 71000 25867
rect 48372 25299 50073 25578
rect 43837 25298 48075 25299
tri 48075 25298 48076 25299 sw
tri 48372 25298 48373 25299 ne
rect 48373 25298 50073 25299
rect 43837 25293 48076 25298
rect 39500 25104 43555 25293
rect 37580 24900 39208 25104
tri 39208 24900 39412 25104 sw
tri 39500 24900 39704 25104 ne
rect 39704 25011 43555 25104
tri 43555 25011 43837 25293 sw
tri 43837 25011 44119 25293 ne
rect 44119 25011 48076 25293
rect 39704 25010 43837 25011
tri 43837 25010 43838 25011 sw
tri 44119 25010 44120 25011 ne
rect 44120 25010 48076 25011
rect 39704 24900 43838 25010
rect 37580 24608 39412 24900
tri 39412 24608 39704 24900 sw
tri 39704 24608 39996 24900 ne
rect 39996 24728 43838 24900
tri 43838 24728 44120 25010 sw
tri 44120 24728 44402 25010 ne
rect 44402 25001 48076 25010
tri 48076 25001 48373 25298 sw
tri 48373 25001 48670 25298 ne
rect 48670 25289 50073 25298
tri 50073 25289 50362 25578 sw
tri 50362 25289 50651 25578 ne
rect 50651 25289 71000 25578
rect 48670 25001 50362 25289
rect 44402 24728 48373 25001
rect 39996 24727 44120 24728
tri 44120 24727 44121 24728 sw
tri 44402 24727 44403 24728 ne
rect 44403 24727 48373 24728
rect 39996 24608 44121 24727
rect 37580 24443 39704 24608
tri 39704 24443 39869 24608 sw
tri 39996 24443 40161 24608 ne
rect 40161 24445 44121 24608
tri 44121 24445 44403 24727 sw
tri 44403 24445 44685 24727 ne
rect 44685 24704 48373 24727
tri 48373 24704 48670 25001 sw
tri 48670 24704 48967 25001 ne
rect 48967 25000 50362 25001
tri 50362 25000 50651 25289 sw
tri 50651 25200 50740 25289 ne
rect 50740 25200 71000 25289
rect 48967 24704 71000 25000
rect 44685 24644 48670 24704
tri 48670 24644 48730 24704 sw
tri 48967 24644 49027 24704 ne
rect 49027 24644 71000 24704
rect 44685 24445 48730 24644
rect 40161 24443 44403 24445
rect 37580 24151 39869 24443
tri 39869 24151 40161 24443 sw
tri 40161 24151 40453 24443 ne
rect 40453 24362 44403 24443
tri 44403 24362 44486 24445 sw
tri 44685 24362 44768 24445 ne
rect 44768 24362 48730 24445
rect 40453 24151 44486 24362
rect 37580 24150 40161 24151
tri 40161 24150 40162 24151 sw
tri 40453 24150 40454 24151 ne
rect 40454 24150 44486 24151
rect 37580 23858 40162 24150
tri 40162 23858 40454 24150 sw
tri 40454 23858 40746 24150 ne
rect 40746 24080 44486 24150
tri 44486 24080 44768 24362 sw
tri 44768 24080 45050 24362 ne
rect 45050 24347 48730 24362
tri 48730 24347 49027 24644 sw
tri 49027 24347 49324 24644 ne
rect 49324 24347 71000 24644
rect 45050 24108 49027 24347
tri 49027 24108 49266 24347 sw
tri 49324 24108 49563 24347 ne
rect 49563 24108 71000 24347
rect 45050 24080 49266 24108
rect 40746 23877 44768 24080
tri 44768 23877 44971 24080 sw
tri 45050 23877 45253 24080 ne
rect 45253 23996 49266 24080
tri 49266 23996 49378 24108 sw
tri 49563 23996 49675 24108 ne
rect 49675 23996 71000 24108
rect 45253 23877 49378 23996
rect 40746 23858 44971 23877
rect 37580 23857 40454 23858
tri 40454 23857 40455 23858 sw
tri 40746 23857 40747 23858 ne
rect 40747 23857 44971 23858
rect 37580 23565 40455 23857
tri 40455 23565 40747 23857 sw
tri 40747 23565 41039 23857 ne
rect 41039 23595 44971 23857
tri 44971 23595 45253 23877 sw
tri 45253 23595 45535 23877 ne
rect 45535 23699 49378 23877
tri 49378 23699 49675 23996 sw
tri 49675 23699 49972 23996 ne
rect 49972 23699 71000 23996
rect 45535 23698 49675 23699
tri 49675 23698 49676 23699 sw
tri 49972 23698 49973 23699 ne
rect 49973 23698 71000 23699
rect 45535 23595 49676 23698
rect 41039 23565 45253 23595
rect 37580 23564 40747 23565
tri 40747 23564 40748 23565 sw
tri 41039 23564 41040 23565 ne
rect 41040 23564 45253 23565
rect 37580 23272 40748 23564
tri 40748 23272 41040 23564 sw
tri 41040 23272 41332 23564 ne
rect 41332 23401 45253 23564
tri 45253 23401 45447 23595 sw
tri 45535 23401 45729 23595 ne
rect 45729 23401 49676 23595
tri 49676 23401 49973 23698 sw
tri 49973 23600 50071 23698 ne
rect 50071 23600 71000 23698
rect 41332 23272 45447 23401
rect 37580 23271 41040 23272
tri 41040 23271 41041 23272 sw
tri 41332 23271 41333 23272 ne
rect 41333 23271 45447 23272
rect 37580 22979 41041 23271
tri 41041 22979 41333 23271 sw
tri 41333 22979 41625 23271 ne
rect 41625 23119 45447 23271
tri 45447 23119 45729 23401 sw
tri 45729 23119 46011 23401 ne
rect 46011 23400 49973 23401
tri 49973 23400 49974 23401 sw
rect 46011 23119 71000 23400
rect 41625 23117 45729 23119
tri 45729 23117 45731 23119 sw
tri 46011 23117 46013 23119 ne
rect 46013 23117 71000 23119
rect 41625 22979 45731 23117
rect 37580 22977 41333 22979
tri 41333 22977 41335 22979 sw
tri 41625 22977 41627 22979 ne
rect 41627 22977 45731 22979
rect 37580 22685 41335 22977
tri 41335 22685 41627 22977 sw
tri 41627 22685 41919 22977 ne
rect 41919 22835 45731 22977
tri 45731 22835 46013 23117 sw
tri 46013 22835 46295 23117 ne
rect 46295 22835 71000 23117
rect 41919 22834 46013 22835
tri 46013 22834 46014 22835 sw
tri 46295 22834 46296 22835 ne
rect 46296 22834 71000 22835
rect 41919 22685 46014 22834
rect 37580 22488 41627 22685
tri 41627 22488 41824 22685 sw
tri 41919 22488 42116 22685 ne
rect 42116 22552 46014 22685
tri 46014 22552 46296 22834 sw
tri 46296 22552 46578 22834 ne
rect 46578 22552 71000 22834
rect 42116 22551 46296 22552
tri 46296 22551 46297 22552 sw
tri 46578 22551 46579 22552 ne
rect 46579 22551 71000 22552
rect 42116 22488 46297 22551
tri 37580 18244 41824 22488 ne
tri 41824 22196 42116 22488 sw
tri 42116 22196 42408 22488 ne
rect 42408 22269 46297 22488
tri 46297 22269 46579 22551 sw
tri 46579 22269 46861 22551 ne
rect 46861 22269 71000 22551
rect 42408 22268 46579 22269
tri 46579 22268 46580 22269 sw
tri 46861 22268 46862 22269 ne
rect 46862 22268 71000 22269
rect 42408 22196 46580 22268
rect 41824 22123 42116 22196
tri 42116 22123 42189 22196 sw
tri 42408 22123 42481 22196 ne
rect 42481 22123 46580 22196
rect 41824 21831 42189 22123
tri 42189 21831 42481 22123 sw
tri 42481 21831 42773 22123 ne
rect 42773 21986 46580 22123
tri 46580 21986 46862 22268 sw
tri 46862 21986 47144 22268 ne
rect 47144 21986 71000 22268
rect 42773 21985 46862 21986
tri 46862 21985 46863 21986 sw
tri 47144 21985 47145 21986 ne
rect 47145 21985 71000 21986
rect 42773 21831 46863 21985
rect 41824 21830 42481 21831
tri 42481 21830 42482 21831 sw
tri 42773 21830 42774 21831 ne
rect 42774 21830 46863 21831
rect 41824 21538 42482 21830
tri 42482 21538 42774 21830 sw
tri 42774 21538 43066 21830 ne
rect 43066 21703 46863 21830
tri 46863 21703 47145 21985 sw
tri 47145 21703 47427 21985 ne
rect 47427 21703 71000 21985
rect 43066 21538 47145 21703
rect 41824 21537 42774 21538
tri 42774 21537 42775 21538 sw
tri 43066 21537 43067 21538 ne
rect 43067 21537 47145 21538
rect 41824 21245 42775 21537
tri 42775 21245 43067 21537 sw
tri 43067 21245 43359 21537 ne
rect 43359 21444 47145 21537
tri 47145 21444 47404 21703 sw
tri 47427 21444 47686 21703 ne
rect 47686 21444 71000 21703
rect 43359 21245 47404 21444
rect 41824 21152 43067 21245
tri 43067 21152 43160 21245 sw
tri 43359 21152 43452 21245 ne
rect 43452 21162 47404 21245
tri 47404 21162 47686 21444 sw
tri 47686 21162 47968 21444 ne
rect 47968 21162 71000 21444
rect 43452 21152 47686 21162
rect 41824 20860 43160 21152
tri 43160 20860 43452 21152 sw
tri 43452 20860 43744 21152 ne
rect 43744 21050 47686 21152
tri 47686 21050 47798 21162 sw
tri 47968 21050 48080 21162 ne
rect 48080 21050 71000 21162
rect 43744 20860 47798 21050
rect 41824 20657 43452 20860
tri 43452 20657 43655 20860 sw
tri 43744 20657 43947 20860 ne
rect 43947 20768 47798 20860
tri 47798 20768 48080 21050 sw
tri 48080 20768 48362 21050 ne
rect 48362 20768 71000 21050
rect 43947 20767 48080 20768
tri 48080 20767 48081 20768 sw
tri 48362 20767 48363 20768 ne
rect 48363 20767 71000 20768
rect 43947 20657 48081 20767
rect 41824 20365 43655 20657
tri 43655 20365 43947 20657 sw
tri 43947 20365 44239 20657 ne
rect 44239 20485 48081 20657
tri 48081 20485 48363 20767 sw
tri 48363 20485 48645 20767 ne
rect 48645 20485 71000 20767
rect 44239 20484 48363 20485
tri 48363 20484 48364 20485 sw
tri 48645 20484 48646 20485 ne
rect 48646 20484 71000 20485
rect 44239 20365 48364 20484
rect 41824 20201 43947 20365
tri 43947 20201 44111 20365 sw
tri 44239 20201 44403 20365 ne
rect 44403 20202 48364 20365
tri 48364 20202 48646 20484 sw
tri 48646 20400 48730 20484 ne
rect 48730 20400 71000 20484
rect 44403 20201 48646 20202
rect 41824 19909 44111 20201
tri 44111 19909 44403 20201 sw
tri 44403 19909 44695 20201 ne
rect 44695 20200 48646 20201
tri 48646 20200 48648 20202 sw
rect 44695 19909 71000 20200
rect 41824 19907 44403 19909
tri 44403 19907 44405 19909 sw
tri 44695 19907 44697 19909 ne
rect 44697 19907 71000 19909
rect 41824 19615 44405 19907
tri 44405 19615 44697 19907 sw
tri 44697 19615 44989 19907 ne
rect 44989 19615 71000 19907
rect 41824 19614 44697 19615
tri 44697 19614 44698 19615 sw
tri 44989 19614 44990 19615 ne
rect 44990 19614 71000 19615
rect 41824 19322 44698 19614
tri 44698 19322 44990 19614 sw
tri 44990 19322 45282 19614 ne
rect 45282 19322 71000 19614
rect 41824 19321 44990 19322
tri 44990 19321 44991 19322 sw
tri 45282 19321 45283 19322 ne
rect 45283 19321 71000 19322
rect 41824 19029 44991 19321
tri 44991 19029 45283 19321 sw
tri 45283 19029 45575 19321 ne
rect 45575 19029 71000 19321
rect 41824 19028 45283 19029
tri 45283 19028 45284 19029 sw
tri 45575 19028 45576 19029 ne
rect 45576 19028 71000 19029
rect 41824 18736 45284 19028
tri 45284 18736 45576 19028 sw
tri 45576 18736 45868 19028 ne
rect 45868 18736 71000 19028
rect 41824 18735 45576 18736
tri 45576 18735 45577 18736 sw
tri 45868 18735 45869 18736 ne
rect 45869 18735 71000 18736
rect 41824 18443 45577 18735
tri 45577 18443 45869 18735 sw
tri 45869 18443 46161 18735 ne
rect 46161 18443 71000 18735
rect 41824 18244 45869 18443
tri 45869 18244 46068 18443 sw
tri 46161 18244 46360 18443 ne
rect 46360 18244 71000 18443
tri 41824 14000 46068 18244 ne
tri 46068 17952 46360 18244 sw
tri 46360 17952 46652 18244 ne
rect 46652 17952 71000 18244
rect 46068 17880 46360 17952
tri 46360 17880 46432 17952 sw
tri 46652 17880 46724 17952 ne
rect 46724 17880 71000 17952
rect 46068 17588 46432 17880
tri 46432 17588 46724 17880 sw
tri 46724 17588 47016 17880 ne
rect 47016 17588 71000 17880
rect 46068 17587 46724 17588
tri 46724 17587 46725 17588 sw
tri 47016 17587 47017 17588 ne
rect 47017 17587 71000 17588
rect 46068 17295 46725 17587
tri 46725 17295 47017 17587 sw
tri 47017 17295 47309 17587 ne
rect 47309 17295 71000 17587
rect 46068 17294 47017 17295
tri 47017 17294 47018 17295 sw
tri 47309 17294 47310 17295 ne
rect 47310 17294 71000 17295
rect 46068 17002 47018 17294
tri 47018 17002 47310 17294 sw
tri 47310 17200 47404 17294 ne
rect 47404 17200 71000 17294
rect 46068 17000 47310 17002
tri 47310 17000 47312 17002 sw
rect 46068 14000 71000 17000
use M1_PSUB_CDNS_69033583165334  M1_PSUB_CDNS_69033583165334_0
timestamp 1713338890
transform 1 0 41636 0 1 70900
box -28281 -97 28281 97
use M1_PSUB_CDNS_69033583165334  M1_PSUB_CDNS_69033583165334_1
timestamp 1713338890
transform 0 -1 70899 1 0 41649
box -28281 -97 28281 97
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_0
timestamp 1713338890
transform 1 0 44873 0 1 13233
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_1
timestamp 1713338890
transform 1 0 44561 0 1 13517
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_2
timestamp 1713338890
transform 1 0 44693 0 1 13385
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_3
timestamp 1713338890
transform 1 0 44429 0 1 13649
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_4
timestamp 1713338890
transform 1 0 44165 0 1 13913
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_5
timestamp 1713338890
transform 1 0 44297 0 1 13781
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_6
timestamp 1713338890
transform 1 0 44033 0 1 14045
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_7
timestamp 1713338890
transform 1 0 43769 0 1 14309
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_8
timestamp 1713338890
transform 1 0 43901 0 1 14177
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_9
timestamp 1713338890
transform 1 0 43637 0 1 14441
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_10
timestamp 1713338890
transform 1 0 43505 0 1 14573
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_11
timestamp 1713338890
transform 1 0 43241 0 1 14837
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_12
timestamp 1713338890
transform 1 0 43373 0 1 14705
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_13
timestamp 1713338890
transform 1 0 43109 0 1 14969
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_14
timestamp 1713338890
transform 1 0 42845 0 1 15233
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_15
timestamp 1713338890
transform 1 0 42977 0 1 15101
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_16
timestamp 1713338890
transform 1 0 42713 0 1 15365
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_17
timestamp 1713338890
transform 1 0 42449 0 1 15629
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_18
timestamp 1713338890
transform 1 0 42581 0 1 15497
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_19
timestamp 1713338890
transform 1 0 42317 0 1 15761
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_20
timestamp 1713338890
transform 1 0 42053 0 1 16025
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_21
timestamp 1713338890
transform 1 0 42185 0 1 15893
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_22
timestamp 1713338890
transform 1 0 39545 0 1 18533
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_23
timestamp 1713338890
transform 1 0 39677 0 1 18401
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_24
timestamp 1713338890
transform 1 0 39809 0 1 18269
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_25
timestamp 1713338890
transform 1 0 39941 0 1 18137
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_26
timestamp 1713338890
transform 1 0 40073 0 1 18005
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_27
timestamp 1713338890
transform 1 0 40205 0 1 17873
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_28
timestamp 1713338890
transform 1 0 39281 0 1 18797
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_29
timestamp 1713338890
transform 1 0 39413 0 1 18665
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_30
timestamp 1713338890
transform 1 0 40337 0 1 17741
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_31
timestamp 1713338890
transform 1 0 40469 0 1 17609
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_32
timestamp 1713338890
transform 1 0 40601 0 1 17477
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_33
timestamp 1713338890
transform 1 0 40733 0 1 17345
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_34
timestamp 1713338890
transform 1 0 40865 0 1 17213
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_35
timestamp 1713338890
transform 1 0 40997 0 1 17081
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_36
timestamp 1713338890
transform 1 0 41129 0 1 16949
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_37
timestamp 1713338890
transform 1 0 41393 0 1 16685
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_38
timestamp 1713338890
transform 1 0 41261 0 1 16817
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_39
timestamp 1713338890
transform 1 0 41525 0 1 16553
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_40
timestamp 1713338890
transform 1 0 41657 0 1 16421
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_41
timestamp 1713338890
transform 1 0 41789 0 1 16289
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_42
timestamp 1713338890
transform 1 0 41921 0 1 16157
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_43
timestamp 1713338890
transform 1 0 36377 0 1 21701
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_44
timestamp 1713338890
transform 1 0 36509 0 1 21569
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_45
timestamp 1713338890
transform 1 0 37433 0 1 20645
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_46
timestamp 1713338890
transform 1 0 37565 0 1 20513
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_47
timestamp 1713338890
transform 1 0 37697 0 1 20381
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_48
timestamp 1713338890
transform 1 0 36641 0 1 21437
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_49
timestamp 1713338890
transform 1 0 36773 0 1 21305
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_50
timestamp 1713338890
transform 1 0 36905 0 1 21173
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_51
timestamp 1713338890
transform 1 0 37037 0 1 21041
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_52
timestamp 1713338890
transform 1 0 37169 0 1 20909
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_53
timestamp 1713338890
transform 1 0 37301 0 1 20777
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_54
timestamp 1713338890
transform 1 0 37829 0 1 20249
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_55
timestamp 1713338890
transform 1 0 37961 0 1 20117
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_56
timestamp 1713338890
transform 1 0 38093 0 1 19985
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_57
timestamp 1713338890
transform 1 0 38225 0 1 19853
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_58
timestamp 1713338890
transform 1 0 38357 0 1 19721
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_59
timestamp 1713338890
transform 1 0 38489 0 1 19589
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_60
timestamp 1713338890
transform 1 0 38621 0 1 19457
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_61
timestamp 1713338890
transform 1 0 38753 0 1 19325
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_62
timestamp 1713338890
transform 1 0 38885 0 1 19193
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_63
timestamp 1713338890
transform 1 0 39017 0 1 19061
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_64
timestamp 1713338890
transform 1 0 39149 0 1 18929
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_65
timestamp 1713338890
transform 1 0 33473 0 1 24605
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_66
timestamp 1713338890
transform 1 0 34265 0 1 23813
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_67
timestamp 1713338890
transform 1 0 34133 0 1 23945
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_68
timestamp 1713338890
transform 1 0 34001 0 1 24077
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_69
timestamp 1713338890
transform 1 0 33869 0 1 24209
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_70
timestamp 1713338890
transform 1 0 33737 0 1 24341
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_71
timestamp 1713338890
transform 1 0 33605 0 1 24473
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_72
timestamp 1713338890
transform 1 0 35057 0 1 23021
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_73
timestamp 1713338890
transform 1 0 34925 0 1 23153
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_74
timestamp 1713338890
transform 1 0 35189 0 1 22889
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_75
timestamp 1713338890
transform 1 0 35321 0 1 22757
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_76
timestamp 1713338890
transform 1 0 35453 0 1 22625
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_77
timestamp 1713338890
transform 1 0 34793 0 1 23285
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_78
timestamp 1713338890
transform 1 0 34661 0 1 23417
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_79
timestamp 1713338890
transform 1 0 34529 0 1 23549
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_80
timestamp 1713338890
transform 1 0 34397 0 1 23681
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_81
timestamp 1713338890
transform 1 0 35585 0 1 22493
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_82
timestamp 1713338890
transform 1 0 35717 0 1 22361
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_83
timestamp 1713338890
transform 1 0 35849 0 1 22229
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_84
timestamp 1713338890
transform 1 0 35981 0 1 22097
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_85
timestamp 1713338890
transform 1 0 36113 0 1 21965
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_86
timestamp 1713338890
transform 1 0 36245 0 1 21833
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_87
timestamp 1713338890
transform 1 0 30569 0 1 27509
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_88
timestamp 1713338890
transform 1 0 30701 0 1 27377
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_89
timestamp 1713338890
transform 1 0 31097 0 1 26981
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_90
timestamp 1713338890
transform 1 0 30833 0 1 27245
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_91
timestamp 1713338890
transform 1 0 30965 0 1 27113
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_92
timestamp 1713338890
transform 1 0 31229 0 1 26849
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_93
timestamp 1713338890
transform 1 0 31361 0 1 26717
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_94
timestamp 1713338890
transform 1 0 31493 0 1 26585
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_95
timestamp 1713338890
transform 1 0 31625 0 1 26453
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_96
timestamp 1713338890
transform 1 0 31757 0 1 26321
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_97
timestamp 1713338890
transform 1 0 31889 0 1 26189
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_98
timestamp 1713338890
transform 1 0 33077 0 1 25001
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_99
timestamp 1713338890
transform 1 0 32021 0 1 26057
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_100
timestamp 1713338890
transform 1 0 32153 0 1 25925
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_101
timestamp 1713338890
transform 1 0 32285 0 1 25793
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_102
timestamp 1713338890
transform 1 0 32417 0 1 25661
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_103
timestamp 1713338890
transform 1 0 32549 0 1 25529
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_104
timestamp 1713338890
transform 1 0 32681 0 1 25397
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_105
timestamp 1713338890
transform 1 0 32813 0 1 25265
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_106
timestamp 1713338890
transform 1 0 32945 0 1 25133
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_107
timestamp 1713338890
transform 1 0 33341 0 1 24737
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_108
timestamp 1713338890
transform 1 0 33209 0 1 24869
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_109
timestamp 1713338890
transform 1 0 27665 0 1 30413
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_110
timestamp 1713338890
transform 1 0 27797 0 1 30281
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_111
timestamp 1713338890
transform 1 0 27929 0 1 30149
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_112
timestamp 1713338890
transform 1 0 28061 0 1 30017
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_113
timestamp 1713338890
transform 1 0 28193 0 1 29885
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_114
timestamp 1713338890
transform 1 0 28325 0 1 29753
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_115
timestamp 1713338890
transform 1 0 29381 0 1 28697
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_116
timestamp 1713338890
transform 1 0 29513 0 1 28565
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_117
timestamp 1713338890
transform 1 0 28853 0 1 29225
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_118
timestamp 1713338890
transform 1 0 29249 0 1 28829
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_119
timestamp 1713338890
transform 1 0 28457 0 1 29621
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_120
timestamp 1713338890
transform 1 0 28589 0 1 29489
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_121
timestamp 1713338890
transform 1 0 28721 0 1 29357
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_122
timestamp 1713338890
transform 1 0 28985 0 1 29093
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_123
timestamp 1713338890
transform 1 0 29117 0 1 28961
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_124
timestamp 1713338890
transform 1 0 29645 0 1 28433
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_125
timestamp 1713338890
transform 1 0 29777 0 1 28301
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_126
timestamp 1713338890
transform 1 0 29909 0 1 28169
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_127
timestamp 1713338890
transform 1 0 30041 0 1 28037
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_128
timestamp 1713338890
transform 1 0 30173 0 1 27905
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_129
timestamp 1713338890
transform 1 0 30305 0 1 27773
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_130
timestamp 1713338890
transform 1 0 30437 0 1 27641
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_131
timestamp 1713338890
transform 1 0 24893 0 1 33185
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_132
timestamp 1713338890
transform 1 0 24761 0 1 33317
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_133
timestamp 1713338890
transform 1 0 25157 0 1 32921
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_134
timestamp 1713338890
transform 1 0 25289 0 1 32789
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_135
timestamp 1713338890
transform 1 0 25421 0 1 32657
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_136
timestamp 1713338890
transform 1 0 25553 0 1 32525
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_137
timestamp 1713338890
transform 1 0 25685 0 1 32393
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_138
timestamp 1713338890
transform 1 0 25817 0 1 32261
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_139
timestamp 1713338890
transform 1 0 25949 0 1 32129
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_140
timestamp 1713338890
transform 1 0 25025 0 1 33053
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_141
timestamp 1713338890
transform 1 0 27005 0 1 31073
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_142
timestamp 1713338890
transform 1 0 26081 0 1 31997
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_143
timestamp 1713338890
transform 1 0 26213 0 1 31865
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_144
timestamp 1713338890
transform 1 0 26345 0 1 31733
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_145
timestamp 1713338890
transform 1 0 26477 0 1 31601
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_146
timestamp 1713338890
transform 1 0 26609 0 1 31469
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_147
timestamp 1713338890
transform 1 0 26741 0 1 31337
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_148
timestamp 1713338890
transform 1 0 26873 0 1 31205
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_149
timestamp 1713338890
transform 1 0 27137 0 1 30941
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_150
timestamp 1713338890
transform 1 0 27533 0 1 30545
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_151
timestamp 1713338890
transform 1 0 27269 0 1 30809
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_152
timestamp 1713338890
transform 1 0 27401 0 1 30677
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_153
timestamp 1713338890
transform 1 0 21857 0 1 36221
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_154
timestamp 1713338890
transform 1 0 21989 0 1 36089
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_155
timestamp 1713338890
transform 1 0 22121 0 1 35957
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_156
timestamp 1713338890
transform 1 0 22253 0 1 35825
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_157
timestamp 1713338890
transform 1 0 22385 0 1 35693
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_158
timestamp 1713338890
transform 1 0 22517 0 1 35561
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_159
timestamp 1713338890
transform 1 0 22649 0 1 35429
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_160
timestamp 1713338890
transform 1 0 22781 0 1 35297
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_161
timestamp 1713338890
transform 1 0 22913 0 1 35165
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_162
timestamp 1713338890
transform 1 0 23177 0 1 34901
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_163
timestamp 1713338890
transform 1 0 23705 0 1 34373
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_164
timestamp 1713338890
transform 1 0 23573 0 1 34505
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_165
timestamp 1713338890
transform 1 0 23441 0 1 34637
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_166
timestamp 1713338890
transform 1 0 23309 0 1 34769
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_167
timestamp 1713338890
transform 1 0 23045 0 1 35033
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_168
timestamp 1713338890
transform 1 0 24629 0 1 33449
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_169
timestamp 1713338890
transform 1 0 24497 0 1 33581
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_170
timestamp 1713338890
transform 1 0 24365 0 1 33713
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_171
timestamp 1713338890
transform 1 0 24233 0 1 33845
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_172
timestamp 1713338890
transform 1 0 24101 0 1 33977
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_173
timestamp 1713338890
transform 1 0 23837 0 1 34241
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_174
timestamp 1713338890
transform 1 0 23969 0 1 34109
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_175
timestamp 1713338890
transform 1 0 19217 0 1 38861
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_176
timestamp 1713338890
transform 1 0 19085 0 1 38993
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_177
timestamp 1713338890
transform 1 0 19349 0 1 38729
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_178
timestamp 1713338890
transform 1 0 19481 0 1 38597
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_179
timestamp 1713338890
transform 1 0 19613 0 1 38465
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_180
timestamp 1713338890
transform 1 0 19745 0 1 38333
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_181
timestamp 1713338890
transform 1 0 19877 0 1 38201
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_182
timestamp 1713338890
transform 1 0 20009 0 1 38069
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_183
timestamp 1713338890
transform 1 0 20141 0 1 37937
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_184
timestamp 1713338890
transform 1 0 20273 0 1 37805
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_185
timestamp 1713338890
transform 1 0 20405 0 1 37673
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_186
timestamp 1713338890
transform 1 0 21329 0 1 36749
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_187
timestamp 1713338890
transform 1 0 21461 0 1 36617
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_188
timestamp 1713338890
transform 1 0 21593 0 1 36485
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_189
timestamp 1713338890
transform 1 0 21725 0 1 36353
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_190
timestamp 1713338890
transform 1 0 20669 0 1 37409
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_191
timestamp 1713338890
transform 1 0 20801 0 1 37277
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_192
timestamp 1713338890
transform 1 0 20933 0 1 37145
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_193
timestamp 1713338890
transform 1 0 21065 0 1 37013
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_194
timestamp 1713338890
transform 1 0 21197 0 1 36881
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_195
timestamp 1713338890
transform 1 0 20537 0 1 37541
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_196
timestamp 1713338890
transform 1 0 16181 0 1 41897
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_197
timestamp 1713338890
transform 1 0 16313 0 1 41765
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_198
timestamp 1713338890
transform 1 0 16445 0 1 41633
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_199
timestamp 1713338890
transform 1 0 16577 0 1 41501
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_200
timestamp 1713338890
transform 1 0 17237 0 1 40841
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_201
timestamp 1713338890
transform 1 0 16709 0 1 41369
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_202
timestamp 1713338890
transform 1 0 16841 0 1 41237
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_203
timestamp 1713338890
transform 1 0 17105 0 1 40973
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_204
timestamp 1713338890
transform 1 0 17369 0 1 40709
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_205
timestamp 1713338890
transform 1 0 17501 0 1 40577
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_206
timestamp 1713338890
transform 1 0 17633 0 1 40445
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_207
timestamp 1713338890
transform 1 0 17765 0 1 40313
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_208
timestamp 1713338890
transform 1 0 16973 0 1 41105
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_209
timestamp 1713338890
transform 1 0 18821 0 1 39257
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_210
timestamp 1713338890
transform 1 0 18953 0 1 39125
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_211
timestamp 1713338890
transform 1 0 17897 0 1 40181
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_212
timestamp 1713338890
transform 1 0 18029 0 1 40049
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_213
timestamp 1713338890
transform 1 0 18161 0 1 39917
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_214
timestamp 1713338890
transform 1 0 18293 0 1 39785
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_215
timestamp 1713338890
transform 1 0 18425 0 1 39653
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_216
timestamp 1713338890
transform 1 0 18557 0 1 39521
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_217
timestamp 1713338890
transform 1 0 18689 0 1 39389
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_218
timestamp 1713338890
transform 1 0 16049 0 1 42029
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_219
timestamp 1713338890
transform 1 0 14729 0 1 43349
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_220
timestamp 1713338890
transform 1 0 14861 0 1 43217
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_221
timestamp 1713338890
transform 1 0 14993 0 1 43085
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_222
timestamp 1713338890
transform 1 0 15257 0 1 42821
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_223
timestamp 1713338890
transform 1 0 15389 0 1 42689
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_224
timestamp 1713338890
transform 1 0 15521 0 1 42557
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_225
timestamp 1713338890
transform 1 0 15653 0 1 42425
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_226
timestamp 1713338890
transform 1 0 15125 0 1 42953
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_227
timestamp 1713338890
transform 1 0 15785 0 1 42293
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_228
timestamp 1713338890
transform 1 0 15917 0 1 42161
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_229
timestamp 1713338890
transform 1 0 14069 0 1 44009
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_230
timestamp 1713338890
transform 1 0 14201 0 1 43877
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_231
timestamp 1713338890
transform 1 0 14333 0 1 43745
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_232
timestamp 1713338890
transform 1 0 13541 0 1 44537
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_233
timestamp 1713338890
transform 1 0 13673 0 1 44405
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_234
timestamp 1713338890
transform 1 0 13805 0 1 44273
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_235
timestamp 1713338890
transform 1 0 13937 0 1 44141
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_236
timestamp 1713338890
transform 1 0 14465 0 1 43613
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_237
timestamp 1713338890
transform 1 0 14597 0 1 43481
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_238
timestamp 1713338890
transform 1 0 13277 0 1 44801
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165335  M1_PSUB_CDNS_69033583165335_239
timestamp 1713338890
transform 1 0 13409 0 1 44669
box -45 -45 45 45
use M1_PSUB_CDNS_69033583165337  M1_PSUB_CDNS_69033583165337_0
timestamp 1713338890
transform 1 0 70235 0 1 69871
box -461 -97 461 97
use M1_PSUB_CDNS_69033583165338  M1_PSUB_CDNS_69033583165338_0
timestamp 1713338890
transform 0 -1 69871 1 0 70385
box -357 -97 357 97
use M1_PSUB_CDNS_69033583165340  M1_PSUB_CDNS_69033583165340_0
timestamp 1713338890
transform 0 -1 13194 1 0 58004
box -12993 -97 12993 97
use M1_PSUB_CDNS_69033583165341  M1_PSUB_CDNS_69033583165341_0
timestamp 1713338890
transform -1 0 58007 0 -1 13194
box -12941 -97 12941 97
use M3_M2_CDNS_69033583165336  M3_M2_CDNS_69033583165336_0
timestamp 1713338890
transform 1 0 70641 0 1 24306
box -38 -610 38 610
use M3_M2_CDNS_69033583165336  M3_M2_CDNS_69033583165336_1
timestamp 1713338890
transform 1 0 70641 0 1 41897
box -38 -610 38 610
use M3_M2_CDNS_69033583165336  M3_M2_CDNS_69033583165336_2
timestamp 1713338890
transform 1 0 70641 0 1 53122
box -38 -610 38 610
use M3_M2_CDNS_69033583165336  M3_M2_CDNS_69033583165336_3
timestamp 1713338890
transform 1 0 70641 0 1 56310
box -38 -610 38 610
use M3_M2_CDNS_69033583165336  M3_M2_CDNS_69033583165336_4
timestamp 1713338890
transform 1 0 70641 0 1 54702
box -38 -610 38 610
use M3_M2_CDNS_69033583165336  M3_M2_CDNS_69033583165336_5
timestamp 1713338890
transform 1 0 70641 0 1 59520
box -38 -610 38 610
use M3_M2_CDNS_69033583165336  M3_M2_CDNS_69033583165336_6
timestamp 1713338890
transform 1 0 70641 0 1 67516
box -38 -610 38 610
use M3_M2_CDNS_69033583165339  M3_M2_CDNS_69033583165339_0
timestamp 1713338890
transform 1 0 70641 0 1 28320
box -38 -1442 38 1442
use M3_M2_CDNS_69033583165339  M3_M2_CDNS_69033583165339_1
timestamp 1713338890
transform 1 0 70641 0 1 31488
box -38 -1442 38 1442
use M3_M2_CDNS_69033583165339  M3_M2_CDNS_69033583165339_2
timestamp 1713338890
transform 1 0 70641 0 1 34700
box -38 -1442 38 1442
use M3_M2_CDNS_69033583165339  M3_M2_CDNS_69033583165339_3
timestamp 1713338890
transform 1 0 70641 0 1 37900
box -38 -1442 38 1442
use M3_M2_CDNS_69033583165339  M3_M2_CDNS_69033583165339_4
timestamp 1713338890
transform 1 0 70641 0 1 44307
box -38 -1442 38 1442
<< labels >>
rlabel metal3 s 70454 61011 70454 61011 4 DVSS
port 1 nsew
rlabel metal3 s 70454 65976 70454 65976 4 DVSS
port 1 nsew
rlabel metal3 s 70454 69002 70454 69002 4 DVSS
port 1 nsew
rlabel metal3 s 70454 57811 70454 57811 4 DVSS
port 1 nsew
rlabel metal3 s 70454 47548 70454 47548 4 DVSS
port 1 nsew
rlabel metal3 s 70454 40295 70454 40295 4 DVSS
port 1 nsew
rlabel metal3 s 70454 26053 70454 26053 4 DVSS
port 1 nsew
rlabel metal3 s 70454 21860 70454 21860 4 DVSS
port 1 nsew
rlabel metal3 s 70385 18874 70385 18874 4 DVSS
port 1 nsew
rlabel metal3 s 70432 15703 70432 15703 4 DVSS
port 1 nsew
rlabel metal3 s 70454 67411 70454 67411 4 DVDD
port 2 nsew
rlabel metal3 s 70454 59576 70454 59576 4 DVDD
port 2 nsew
rlabel metal3 s 70454 56376 70454 56376 4 DVDD
port 2 nsew
rlabel metal3 s 70454 54611 70454 54611 4 DVDD
port 2 nsew
rlabel metal3 s 70454 53176 70454 53176 4 DVDD
port 2 nsew
rlabel metal3 s 70454 44321 70454 44321 4 DVDD
port 2 nsew
rlabel metal3 s 70454 41930 70454 41930 4 DVDD
port 2 nsew
rlabel metal3 s 70454 37912 70454 37912 4 DVDD
port 2 nsew
rlabel metal3 s 70454 34676 70454 34676 4 DVDD
port 2 nsew
rlabel metal3 s 70454 31562 70454 31562 4 DVDD
port 2 nsew
rlabel metal3 s 70454 28347 70454 28347 4 DVDD
port 2 nsew
rlabel metal3 s 70454 24237 70454 24237 4 DVDD
port 2 nsew
rlabel metal3 s 70454 64211 70454 64211 4 VSS
port 3 nsew
rlabel metal3 s 70559 49976 70559 49976 4 VSS
port 3 nsew
rlabel metal3 s 70454 62776 70454 62776 4 VDD
port 4 nsew
rlabel metal3 s 70559 51411 70559 51411 4 VDD
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 71000 71000
<< end >>
