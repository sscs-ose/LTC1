magic
tech gf180mcuC
magscale 1 10
timestamp 1691402935
<< nwell >>
rect -1082 -834 1082 834
<< pmos >>
rect -908 454 -852 704
rect -748 454 -692 704
rect -588 454 -532 704
rect -428 454 -372 704
rect -268 454 -212 704
rect -108 454 -52 704
rect 52 454 108 704
rect 212 454 268 704
rect 372 454 428 704
rect 532 454 588 704
rect 692 454 748 704
rect 852 454 908 704
rect -908 68 -852 318
rect -748 68 -692 318
rect -588 68 -532 318
rect -428 68 -372 318
rect -268 68 -212 318
rect -108 68 -52 318
rect 52 68 108 318
rect 212 68 268 318
rect 372 68 428 318
rect 532 68 588 318
rect 692 68 748 318
rect 852 68 908 318
rect -908 -318 -852 -68
rect -748 -318 -692 -68
rect -588 -318 -532 -68
rect -428 -318 -372 -68
rect -268 -318 -212 -68
rect -108 -318 -52 -68
rect 52 -318 108 -68
rect 212 -318 268 -68
rect 372 -318 428 -68
rect 532 -318 588 -68
rect 692 -318 748 -68
rect 852 -318 908 -68
rect -908 -704 -852 -454
rect -748 -704 -692 -454
rect -588 -704 -532 -454
rect -428 -704 -372 -454
rect -268 -704 -212 -454
rect -108 -704 -52 -454
rect 52 -704 108 -454
rect 212 -704 268 -454
rect 372 -704 428 -454
rect 532 -704 588 -454
rect 692 -704 748 -454
rect 852 -704 908 -454
<< pdiff >>
rect -996 691 -908 704
rect -996 467 -983 691
rect -937 467 -908 691
rect -996 454 -908 467
rect -852 691 -748 704
rect -852 467 -823 691
rect -777 467 -748 691
rect -852 454 -748 467
rect -692 691 -588 704
rect -692 467 -663 691
rect -617 467 -588 691
rect -692 454 -588 467
rect -532 691 -428 704
rect -532 467 -503 691
rect -457 467 -428 691
rect -532 454 -428 467
rect -372 691 -268 704
rect -372 467 -343 691
rect -297 467 -268 691
rect -372 454 -268 467
rect -212 691 -108 704
rect -212 467 -183 691
rect -137 467 -108 691
rect -212 454 -108 467
rect -52 691 52 704
rect -52 467 -23 691
rect 23 467 52 691
rect -52 454 52 467
rect 108 691 212 704
rect 108 467 137 691
rect 183 467 212 691
rect 108 454 212 467
rect 268 691 372 704
rect 268 467 297 691
rect 343 467 372 691
rect 268 454 372 467
rect 428 691 532 704
rect 428 467 457 691
rect 503 467 532 691
rect 428 454 532 467
rect 588 691 692 704
rect 588 467 617 691
rect 663 467 692 691
rect 588 454 692 467
rect 748 691 852 704
rect 748 467 777 691
rect 823 467 852 691
rect 748 454 852 467
rect 908 691 996 704
rect 908 467 937 691
rect 983 467 996 691
rect 908 454 996 467
rect -996 305 -908 318
rect -996 81 -983 305
rect -937 81 -908 305
rect -996 68 -908 81
rect -852 305 -748 318
rect -852 81 -823 305
rect -777 81 -748 305
rect -852 68 -748 81
rect -692 305 -588 318
rect -692 81 -663 305
rect -617 81 -588 305
rect -692 68 -588 81
rect -532 305 -428 318
rect -532 81 -503 305
rect -457 81 -428 305
rect -532 68 -428 81
rect -372 305 -268 318
rect -372 81 -343 305
rect -297 81 -268 305
rect -372 68 -268 81
rect -212 305 -108 318
rect -212 81 -183 305
rect -137 81 -108 305
rect -212 68 -108 81
rect -52 305 52 318
rect -52 81 -23 305
rect 23 81 52 305
rect -52 68 52 81
rect 108 305 212 318
rect 108 81 137 305
rect 183 81 212 305
rect 108 68 212 81
rect 268 305 372 318
rect 268 81 297 305
rect 343 81 372 305
rect 268 68 372 81
rect 428 305 532 318
rect 428 81 457 305
rect 503 81 532 305
rect 428 68 532 81
rect 588 305 692 318
rect 588 81 617 305
rect 663 81 692 305
rect 588 68 692 81
rect 748 305 852 318
rect 748 81 777 305
rect 823 81 852 305
rect 748 68 852 81
rect 908 305 996 318
rect 908 81 937 305
rect 983 81 996 305
rect 908 68 996 81
rect -996 -81 -908 -68
rect -996 -305 -983 -81
rect -937 -305 -908 -81
rect -996 -318 -908 -305
rect -852 -81 -748 -68
rect -852 -305 -823 -81
rect -777 -305 -748 -81
rect -852 -318 -748 -305
rect -692 -81 -588 -68
rect -692 -305 -663 -81
rect -617 -305 -588 -81
rect -692 -318 -588 -305
rect -532 -81 -428 -68
rect -532 -305 -503 -81
rect -457 -305 -428 -81
rect -532 -318 -428 -305
rect -372 -81 -268 -68
rect -372 -305 -343 -81
rect -297 -305 -268 -81
rect -372 -318 -268 -305
rect -212 -81 -108 -68
rect -212 -305 -183 -81
rect -137 -305 -108 -81
rect -212 -318 -108 -305
rect -52 -81 52 -68
rect -52 -305 -23 -81
rect 23 -305 52 -81
rect -52 -318 52 -305
rect 108 -81 212 -68
rect 108 -305 137 -81
rect 183 -305 212 -81
rect 108 -318 212 -305
rect 268 -81 372 -68
rect 268 -305 297 -81
rect 343 -305 372 -81
rect 268 -318 372 -305
rect 428 -81 532 -68
rect 428 -305 457 -81
rect 503 -305 532 -81
rect 428 -318 532 -305
rect 588 -81 692 -68
rect 588 -305 617 -81
rect 663 -305 692 -81
rect 588 -318 692 -305
rect 748 -81 852 -68
rect 748 -305 777 -81
rect 823 -305 852 -81
rect 748 -318 852 -305
rect 908 -81 996 -68
rect 908 -305 937 -81
rect 983 -305 996 -81
rect 908 -318 996 -305
rect -996 -467 -908 -454
rect -996 -691 -983 -467
rect -937 -691 -908 -467
rect -996 -704 -908 -691
rect -852 -467 -748 -454
rect -852 -691 -823 -467
rect -777 -691 -748 -467
rect -852 -704 -748 -691
rect -692 -467 -588 -454
rect -692 -691 -663 -467
rect -617 -691 -588 -467
rect -692 -704 -588 -691
rect -532 -467 -428 -454
rect -532 -691 -503 -467
rect -457 -691 -428 -467
rect -532 -704 -428 -691
rect -372 -467 -268 -454
rect -372 -691 -343 -467
rect -297 -691 -268 -467
rect -372 -704 -268 -691
rect -212 -467 -108 -454
rect -212 -691 -183 -467
rect -137 -691 -108 -467
rect -212 -704 -108 -691
rect -52 -467 52 -454
rect -52 -691 -23 -467
rect 23 -691 52 -467
rect -52 -704 52 -691
rect 108 -467 212 -454
rect 108 -691 137 -467
rect 183 -691 212 -467
rect 108 -704 212 -691
rect 268 -467 372 -454
rect 268 -691 297 -467
rect 343 -691 372 -467
rect 268 -704 372 -691
rect 428 -467 532 -454
rect 428 -691 457 -467
rect 503 -691 532 -467
rect 428 -704 532 -691
rect 588 -467 692 -454
rect 588 -691 617 -467
rect 663 -691 692 -467
rect 588 -704 692 -691
rect 748 -467 852 -454
rect 748 -691 777 -467
rect 823 -691 852 -467
rect 748 -704 852 -691
rect 908 -467 996 -454
rect 908 -691 937 -467
rect 983 -691 996 -467
rect 908 -704 996 -691
<< pdiffc >>
rect -983 467 -937 691
rect -823 467 -777 691
rect -663 467 -617 691
rect -503 467 -457 691
rect -343 467 -297 691
rect -183 467 -137 691
rect -23 467 23 691
rect 137 467 183 691
rect 297 467 343 691
rect 457 467 503 691
rect 617 467 663 691
rect 777 467 823 691
rect 937 467 983 691
rect -983 81 -937 305
rect -823 81 -777 305
rect -663 81 -617 305
rect -503 81 -457 305
rect -343 81 -297 305
rect -183 81 -137 305
rect -23 81 23 305
rect 137 81 183 305
rect 297 81 343 305
rect 457 81 503 305
rect 617 81 663 305
rect 777 81 823 305
rect 937 81 983 305
rect -983 -305 -937 -81
rect -823 -305 -777 -81
rect -663 -305 -617 -81
rect -503 -305 -457 -81
rect -343 -305 -297 -81
rect -183 -305 -137 -81
rect -23 -305 23 -81
rect 137 -305 183 -81
rect 297 -305 343 -81
rect 457 -305 503 -81
rect 617 -305 663 -81
rect 777 -305 823 -81
rect 937 -305 983 -81
rect -983 -691 -937 -467
rect -823 -691 -777 -467
rect -663 -691 -617 -467
rect -503 -691 -457 -467
rect -343 -691 -297 -467
rect -183 -691 -137 -467
rect -23 -691 23 -467
rect 137 -691 183 -467
rect 297 -691 343 -467
rect 457 -691 503 -467
rect 617 -691 663 -467
rect 777 -691 823 -467
rect 937 -691 983 -467
<< polysilicon >>
rect -908 704 -852 748
rect -748 704 -692 748
rect -588 704 -532 748
rect -428 704 -372 748
rect -268 704 -212 748
rect -108 704 -52 748
rect 52 704 108 748
rect 212 704 268 748
rect 372 704 428 748
rect 532 704 588 748
rect 692 704 748 748
rect 852 704 908 748
rect -908 410 -852 454
rect -748 410 -692 454
rect -588 410 -532 454
rect -428 410 -372 454
rect -268 410 -212 454
rect -108 410 -52 454
rect 52 410 108 454
rect 212 410 268 454
rect 372 410 428 454
rect 532 410 588 454
rect 692 410 748 454
rect 852 410 908 454
rect -908 318 -852 362
rect -748 318 -692 362
rect -588 318 -532 362
rect -428 318 -372 362
rect -268 318 -212 362
rect -108 318 -52 362
rect 52 318 108 362
rect 212 318 268 362
rect 372 318 428 362
rect 532 318 588 362
rect 692 318 748 362
rect 852 318 908 362
rect -908 24 -852 68
rect -748 24 -692 68
rect -588 24 -532 68
rect -428 24 -372 68
rect -268 24 -212 68
rect -108 24 -52 68
rect 52 24 108 68
rect 212 24 268 68
rect 372 24 428 68
rect 532 24 588 68
rect 692 24 748 68
rect 852 24 908 68
rect -908 -68 -852 -24
rect -748 -68 -692 -24
rect -588 -68 -532 -24
rect -428 -68 -372 -24
rect -268 -68 -212 -24
rect -108 -68 -52 -24
rect 52 -68 108 -24
rect 212 -68 268 -24
rect 372 -68 428 -24
rect 532 -68 588 -24
rect 692 -68 748 -24
rect 852 -68 908 -24
rect -908 -362 -852 -318
rect -748 -362 -692 -318
rect -588 -362 -532 -318
rect -428 -362 -372 -318
rect -268 -362 -212 -318
rect -108 -362 -52 -318
rect 52 -362 108 -318
rect 212 -362 268 -318
rect 372 -362 428 -318
rect 532 -362 588 -318
rect 692 -362 748 -318
rect 852 -362 908 -318
rect -908 -454 -852 -410
rect -748 -454 -692 -410
rect -588 -454 -532 -410
rect -428 -454 -372 -410
rect -268 -454 -212 -410
rect -108 -454 -52 -410
rect 52 -454 108 -410
rect 212 -454 268 -410
rect 372 -454 428 -410
rect 532 -454 588 -410
rect 692 -454 748 -410
rect 852 -454 908 -410
rect -908 -748 -852 -704
rect -748 -748 -692 -704
rect -588 -748 -532 -704
rect -428 -748 -372 -704
rect -268 -748 -212 -704
rect -108 -748 -52 -704
rect 52 -748 108 -704
rect 212 -748 268 -704
rect 372 -748 428 -704
rect 532 -748 588 -704
rect 692 -748 748 -704
rect 852 -748 908 -704
<< metal1 >>
rect -983 691 -937 702
rect -983 456 -937 467
rect -823 691 -777 702
rect -823 456 -777 467
rect -663 691 -617 702
rect -663 456 -617 467
rect -503 691 -457 702
rect -503 456 -457 467
rect -343 691 -297 702
rect -343 456 -297 467
rect -183 691 -137 702
rect -183 456 -137 467
rect -23 691 23 702
rect -23 456 23 467
rect 137 691 183 702
rect 137 456 183 467
rect 297 691 343 702
rect 297 456 343 467
rect 457 691 503 702
rect 457 456 503 467
rect 617 691 663 702
rect 617 456 663 467
rect 777 691 823 702
rect 777 456 823 467
rect 937 691 983 702
rect 937 456 983 467
rect -983 305 -937 316
rect -983 70 -937 81
rect -823 305 -777 316
rect -823 70 -777 81
rect -663 305 -617 316
rect -663 70 -617 81
rect -503 305 -457 316
rect -503 70 -457 81
rect -343 305 -297 316
rect -343 70 -297 81
rect -183 305 -137 316
rect -183 70 -137 81
rect -23 305 23 316
rect -23 70 23 81
rect 137 305 183 316
rect 137 70 183 81
rect 297 305 343 316
rect 297 70 343 81
rect 457 305 503 316
rect 457 70 503 81
rect 617 305 663 316
rect 617 70 663 81
rect 777 305 823 316
rect 777 70 823 81
rect 937 305 983 316
rect 937 70 983 81
rect -983 -81 -937 -70
rect -983 -316 -937 -305
rect -823 -81 -777 -70
rect -823 -316 -777 -305
rect -663 -81 -617 -70
rect -663 -316 -617 -305
rect -503 -81 -457 -70
rect -503 -316 -457 -305
rect -343 -81 -297 -70
rect -343 -316 -297 -305
rect -183 -81 -137 -70
rect -183 -316 -137 -305
rect -23 -81 23 -70
rect -23 -316 23 -305
rect 137 -81 183 -70
rect 137 -316 183 -305
rect 297 -81 343 -70
rect 297 -316 343 -305
rect 457 -81 503 -70
rect 457 -316 503 -305
rect 617 -81 663 -70
rect 617 -316 663 -305
rect 777 -81 823 -70
rect 777 -316 823 -305
rect 937 -81 983 -70
rect 937 -316 983 -305
rect -983 -467 -937 -456
rect -983 -702 -937 -691
rect -823 -467 -777 -456
rect -823 -702 -777 -691
rect -663 -467 -617 -456
rect -663 -702 -617 -691
rect -503 -467 -457 -456
rect -503 -702 -457 -691
rect -343 -467 -297 -456
rect -343 -702 -297 -691
rect -183 -467 -137 -456
rect -183 -702 -137 -691
rect -23 -467 23 -456
rect -23 -702 23 -691
rect 137 -467 183 -456
rect 137 -702 183 -691
rect 297 -467 343 -456
rect 297 -702 343 -691
rect 457 -467 503 -456
rect 457 -702 503 -691
rect 617 -467 663 -456
rect 617 -702 663 -691
rect 777 -467 823 -456
rect 777 -702 823 -691
rect 937 -467 983 -456
rect 937 -702 983 -691
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 1.25 l 0.280 m 4 nf 12 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
