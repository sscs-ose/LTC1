magic
tech gf180mcuC
magscale 1 10
timestamp 1699925801
<< pwell >>
rect -264 -308 264 308
<< nmos >>
rect -152 -240 -52 240
rect 52 -240 152 240
<< ndiff >>
rect -240 227 -152 240
rect -240 -227 -227 227
rect -181 -227 -152 227
rect -240 -240 -152 -227
rect -52 227 52 240
rect -52 -227 -23 227
rect 23 -227 52 227
rect -52 -240 52 -227
rect 152 227 240 240
rect 152 -227 181 227
rect 227 -227 240 227
rect 152 -240 240 -227
<< ndiffc >>
rect -227 -227 -181 227
rect -23 -227 23 227
rect 181 -227 227 227
<< polysilicon >>
rect -152 240 -52 284
rect 52 240 152 284
rect -152 -284 -52 -240
rect 52 -284 152 -240
<< metal1 >>
rect -227 227 -181 238
rect -227 -238 -181 -227
rect -23 227 23 238
rect -23 -238 23 -227
rect 181 227 227 238
rect 181 -238 227 -227
<< properties >>
string gencell nfet_03v3
string library gf180mcu
string parameters w 2.4 l 0.5 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt}
<< end >>
