magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1513 -3641 1513 3641
<< metal2 >>
rect -513 2636 513 2641
rect -513 2608 -508 2636
rect -480 2608 -432 2636
rect -404 2608 -356 2636
rect -328 2608 -280 2636
rect -252 2608 -204 2636
rect -176 2608 -128 2636
rect -100 2608 -52 2636
rect -24 2608 24 2636
rect 52 2608 100 2636
rect 128 2608 176 2636
rect 204 2608 252 2636
rect 280 2608 328 2636
rect 356 2608 404 2636
rect 432 2608 480 2636
rect 508 2608 513 2636
rect -513 2560 513 2608
rect -513 2532 -508 2560
rect -480 2532 -432 2560
rect -404 2532 -356 2560
rect -328 2532 -280 2560
rect -252 2532 -204 2560
rect -176 2532 -128 2560
rect -100 2532 -52 2560
rect -24 2532 24 2560
rect 52 2532 100 2560
rect 128 2532 176 2560
rect 204 2532 252 2560
rect 280 2532 328 2560
rect 356 2532 404 2560
rect 432 2532 480 2560
rect 508 2532 513 2560
rect -513 2484 513 2532
rect -513 2456 -508 2484
rect -480 2456 -432 2484
rect -404 2456 -356 2484
rect -328 2456 -280 2484
rect -252 2456 -204 2484
rect -176 2456 -128 2484
rect -100 2456 -52 2484
rect -24 2456 24 2484
rect 52 2456 100 2484
rect 128 2456 176 2484
rect 204 2456 252 2484
rect 280 2456 328 2484
rect 356 2456 404 2484
rect 432 2456 480 2484
rect 508 2456 513 2484
rect -513 2408 513 2456
rect -513 2380 -508 2408
rect -480 2380 -432 2408
rect -404 2380 -356 2408
rect -328 2380 -280 2408
rect -252 2380 -204 2408
rect -176 2380 -128 2408
rect -100 2380 -52 2408
rect -24 2380 24 2408
rect 52 2380 100 2408
rect 128 2380 176 2408
rect 204 2380 252 2408
rect 280 2380 328 2408
rect 356 2380 404 2408
rect 432 2380 480 2408
rect 508 2380 513 2408
rect -513 2332 513 2380
rect -513 2304 -508 2332
rect -480 2304 -432 2332
rect -404 2304 -356 2332
rect -328 2304 -280 2332
rect -252 2304 -204 2332
rect -176 2304 -128 2332
rect -100 2304 -52 2332
rect -24 2304 24 2332
rect 52 2304 100 2332
rect 128 2304 176 2332
rect 204 2304 252 2332
rect 280 2304 328 2332
rect 356 2304 404 2332
rect 432 2304 480 2332
rect 508 2304 513 2332
rect -513 2256 513 2304
rect -513 2228 -508 2256
rect -480 2228 -432 2256
rect -404 2228 -356 2256
rect -328 2228 -280 2256
rect -252 2228 -204 2256
rect -176 2228 -128 2256
rect -100 2228 -52 2256
rect -24 2228 24 2256
rect 52 2228 100 2256
rect 128 2228 176 2256
rect 204 2228 252 2256
rect 280 2228 328 2256
rect 356 2228 404 2256
rect 432 2228 480 2256
rect 508 2228 513 2256
rect -513 2180 513 2228
rect -513 2152 -508 2180
rect -480 2152 -432 2180
rect -404 2152 -356 2180
rect -328 2152 -280 2180
rect -252 2152 -204 2180
rect -176 2152 -128 2180
rect -100 2152 -52 2180
rect -24 2152 24 2180
rect 52 2152 100 2180
rect 128 2152 176 2180
rect 204 2152 252 2180
rect 280 2152 328 2180
rect 356 2152 404 2180
rect 432 2152 480 2180
rect 508 2152 513 2180
rect -513 2104 513 2152
rect -513 2076 -508 2104
rect -480 2076 -432 2104
rect -404 2076 -356 2104
rect -328 2076 -280 2104
rect -252 2076 -204 2104
rect -176 2076 -128 2104
rect -100 2076 -52 2104
rect -24 2076 24 2104
rect 52 2076 100 2104
rect 128 2076 176 2104
rect 204 2076 252 2104
rect 280 2076 328 2104
rect 356 2076 404 2104
rect 432 2076 480 2104
rect 508 2076 513 2104
rect -513 2028 513 2076
rect -513 2000 -508 2028
rect -480 2000 -432 2028
rect -404 2000 -356 2028
rect -328 2000 -280 2028
rect -252 2000 -204 2028
rect -176 2000 -128 2028
rect -100 2000 -52 2028
rect -24 2000 24 2028
rect 52 2000 100 2028
rect 128 2000 176 2028
rect 204 2000 252 2028
rect 280 2000 328 2028
rect 356 2000 404 2028
rect 432 2000 480 2028
rect 508 2000 513 2028
rect -513 1952 513 2000
rect -513 1924 -508 1952
rect -480 1924 -432 1952
rect -404 1924 -356 1952
rect -328 1924 -280 1952
rect -252 1924 -204 1952
rect -176 1924 -128 1952
rect -100 1924 -52 1952
rect -24 1924 24 1952
rect 52 1924 100 1952
rect 128 1924 176 1952
rect 204 1924 252 1952
rect 280 1924 328 1952
rect 356 1924 404 1952
rect 432 1924 480 1952
rect 508 1924 513 1952
rect -513 1876 513 1924
rect -513 1848 -508 1876
rect -480 1848 -432 1876
rect -404 1848 -356 1876
rect -328 1848 -280 1876
rect -252 1848 -204 1876
rect -176 1848 -128 1876
rect -100 1848 -52 1876
rect -24 1848 24 1876
rect 52 1848 100 1876
rect 128 1848 176 1876
rect 204 1848 252 1876
rect 280 1848 328 1876
rect 356 1848 404 1876
rect 432 1848 480 1876
rect 508 1848 513 1876
rect -513 1800 513 1848
rect -513 1772 -508 1800
rect -480 1772 -432 1800
rect -404 1772 -356 1800
rect -328 1772 -280 1800
rect -252 1772 -204 1800
rect -176 1772 -128 1800
rect -100 1772 -52 1800
rect -24 1772 24 1800
rect 52 1772 100 1800
rect 128 1772 176 1800
rect 204 1772 252 1800
rect 280 1772 328 1800
rect 356 1772 404 1800
rect 432 1772 480 1800
rect 508 1772 513 1800
rect -513 1724 513 1772
rect -513 1696 -508 1724
rect -480 1696 -432 1724
rect -404 1696 -356 1724
rect -328 1696 -280 1724
rect -252 1696 -204 1724
rect -176 1696 -128 1724
rect -100 1696 -52 1724
rect -24 1696 24 1724
rect 52 1696 100 1724
rect 128 1696 176 1724
rect 204 1696 252 1724
rect 280 1696 328 1724
rect 356 1696 404 1724
rect 432 1696 480 1724
rect 508 1696 513 1724
rect -513 1648 513 1696
rect -513 1620 -508 1648
rect -480 1620 -432 1648
rect -404 1620 -356 1648
rect -328 1620 -280 1648
rect -252 1620 -204 1648
rect -176 1620 -128 1648
rect -100 1620 -52 1648
rect -24 1620 24 1648
rect 52 1620 100 1648
rect 128 1620 176 1648
rect 204 1620 252 1648
rect 280 1620 328 1648
rect 356 1620 404 1648
rect 432 1620 480 1648
rect 508 1620 513 1648
rect -513 1572 513 1620
rect -513 1544 -508 1572
rect -480 1544 -432 1572
rect -404 1544 -356 1572
rect -328 1544 -280 1572
rect -252 1544 -204 1572
rect -176 1544 -128 1572
rect -100 1544 -52 1572
rect -24 1544 24 1572
rect 52 1544 100 1572
rect 128 1544 176 1572
rect 204 1544 252 1572
rect 280 1544 328 1572
rect 356 1544 404 1572
rect 432 1544 480 1572
rect 508 1544 513 1572
rect -513 1496 513 1544
rect -513 1468 -508 1496
rect -480 1468 -432 1496
rect -404 1468 -356 1496
rect -328 1468 -280 1496
rect -252 1468 -204 1496
rect -176 1468 -128 1496
rect -100 1468 -52 1496
rect -24 1468 24 1496
rect 52 1468 100 1496
rect 128 1468 176 1496
rect 204 1468 252 1496
rect 280 1468 328 1496
rect 356 1468 404 1496
rect 432 1468 480 1496
rect 508 1468 513 1496
rect -513 1420 513 1468
rect -513 1392 -508 1420
rect -480 1392 -432 1420
rect -404 1392 -356 1420
rect -328 1392 -280 1420
rect -252 1392 -204 1420
rect -176 1392 -128 1420
rect -100 1392 -52 1420
rect -24 1392 24 1420
rect 52 1392 100 1420
rect 128 1392 176 1420
rect 204 1392 252 1420
rect 280 1392 328 1420
rect 356 1392 404 1420
rect 432 1392 480 1420
rect 508 1392 513 1420
rect -513 1344 513 1392
rect -513 1316 -508 1344
rect -480 1316 -432 1344
rect -404 1316 -356 1344
rect -328 1316 -280 1344
rect -252 1316 -204 1344
rect -176 1316 -128 1344
rect -100 1316 -52 1344
rect -24 1316 24 1344
rect 52 1316 100 1344
rect 128 1316 176 1344
rect 204 1316 252 1344
rect 280 1316 328 1344
rect 356 1316 404 1344
rect 432 1316 480 1344
rect 508 1316 513 1344
rect -513 1268 513 1316
rect -513 1240 -508 1268
rect -480 1240 -432 1268
rect -404 1240 -356 1268
rect -328 1240 -280 1268
rect -252 1240 -204 1268
rect -176 1240 -128 1268
rect -100 1240 -52 1268
rect -24 1240 24 1268
rect 52 1240 100 1268
rect 128 1240 176 1268
rect 204 1240 252 1268
rect 280 1240 328 1268
rect 356 1240 404 1268
rect 432 1240 480 1268
rect 508 1240 513 1268
rect -513 1192 513 1240
rect -513 1164 -508 1192
rect -480 1164 -432 1192
rect -404 1164 -356 1192
rect -328 1164 -280 1192
rect -252 1164 -204 1192
rect -176 1164 -128 1192
rect -100 1164 -52 1192
rect -24 1164 24 1192
rect 52 1164 100 1192
rect 128 1164 176 1192
rect 204 1164 252 1192
rect 280 1164 328 1192
rect 356 1164 404 1192
rect 432 1164 480 1192
rect 508 1164 513 1192
rect -513 1116 513 1164
rect -513 1088 -508 1116
rect -480 1088 -432 1116
rect -404 1088 -356 1116
rect -328 1088 -280 1116
rect -252 1088 -204 1116
rect -176 1088 -128 1116
rect -100 1088 -52 1116
rect -24 1088 24 1116
rect 52 1088 100 1116
rect 128 1088 176 1116
rect 204 1088 252 1116
rect 280 1088 328 1116
rect 356 1088 404 1116
rect 432 1088 480 1116
rect 508 1088 513 1116
rect -513 1040 513 1088
rect -513 1012 -508 1040
rect -480 1012 -432 1040
rect -404 1012 -356 1040
rect -328 1012 -280 1040
rect -252 1012 -204 1040
rect -176 1012 -128 1040
rect -100 1012 -52 1040
rect -24 1012 24 1040
rect 52 1012 100 1040
rect 128 1012 176 1040
rect 204 1012 252 1040
rect 280 1012 328 1040
rect 356 1012 404 1040
rect 432 1012 480 1040
rect 508 1012 513 1040
rect -513 964 513 1012
rect -513 936 -508 964
rect -480 936 -432 964
rect -404 936 -356 964
rect -328 936 -280 964
rect -252 936 -204 964
rect -176 936 -128 964
rect -100 936 -52 964
rect -24 936 24 964
rect 52 936 100 964
rect 128 936 176 964
rect 204 936 252 964
rect 280 936 328 964
rect 356 936 404 964
rect 432 936 480 964
rect 508 936 513 964
rect -513 888 513 936
rect -513 860 -508 888
rect -480 860 -432 888
rect -404 860 -356 888
rect -328 860 -280 888
rect -252 860 -204 888
rect -176 860 -128 888
rect -100 860 -52 888
rect -24 860 24 888
rect 52 860 100 888
rect 128 860 176 888
rect 204 860 252 888
rect 280 860 328 888
rect 356 860 404 888
rect 432 860 480 888
rect 508 860 513 888
rect -513 812 513 860
rect -513 784 -508 812
rect -480 784 -432 812
rect -404 784 -356 812
rect -328 784 -280 812
rect -252 784 -204 812
rect -176 784 -128 812
rect -100 784 -52 812
rect -24 784 24 812
rect 52 784 100 812
rect 128 784 176 812
rect 204 784 252 812
rect 280 784 328 812
rect 356 784 404 812
rect 432 784 480 812
rect 508 784 513 812
rect -513 736 513 784
rect -513 708 -508 736
rect -480 708 -432 736
rect -404 708 -356 736
rect -328 708 -280 736
rect -252 708 -204 736
rect -176 708 -128 736
rect -100 708 -52 736
rect -24 708 24 736
rect 52 708 100 736
rect 128 708 176 736
rect 204 708 252 736
rect 280 708 328 736
rect 356 708 404 736
rect 432 708 480 736
rect 508 708 513 736
rect -513 660 513 708
rect -513 632 -508 660
rect -480 632 -432 660
rect -404 632 -356 660
rect -328 632 -280 660
rect -252 632 -204 660
rect -176 632 -128 660
rect -100 632 -52 660
rect -24 632 24 660
rect 52 632 100 660
rect 128 632 176 660
rect 204 632 252 660
rect 280 632 328 660
rect 356 632 404 660
rect 432 632 480 660
rect 508 632 513 660
rect -513 584 513 632
rect -513 556 -508 584
rect -480 556 -432 584
rect -404 556 -356 584
rect -328 556 -280 584
rect -252 556 -204 584
rect -176 556 -128 584
rect -100 556 -52 584
rect -24 556 24 584
rect 52 556 100 584
rect 128 556 176 584
rect 204 556 252 584
rect 280 556 328 584
rect 356 556 404 584
rect 432 556 480 584
rect 508 556 513 584
rect -513 508 513 556
rect -513 480 -508 508
rect -480 480 -432 508
rect -404 480 -356 508
rect -328 480 -280 508
rect -252 480 -204 508
rect -176 480 -128 508
rect -100 480 -52 508
rect -24 480 24 508
rect 52 480 100 508
rect 128 480 176 508
rect 204 480 252 508
rect 280 480 328 508
rect 356 480 404 508
rect 432 480 480 508
rect 508 480 513 508
rect -513 432 513 480
rect -513 404 -508 432
rect -480 404 -432 432
rect -404 404 -356 432
rect -328 404 -280 432
rect -252 404 -204 432
rect -176 404 -128 432
rect -100 404 -52 432
rect -24 404 24 432
rect 52 404 100 432
rect 128 404 176 432
rect 204 404 252 432
rect 280 404 328 432
rect 356 404 404 432
rect 432 404 480 432
rect 508 404 513 432
rect -513 356 513 404
rect -513 328 -508 356
rect -480 328 -432 356
rect -404 328 -356 356
rect -328 328 -280 356
rect -252 328 -204 356
rect -176 328 -128 356
rect -100 328 -52 356
rect -24 328 24 356
rect 52 328 100 356
rect 128 328 176 356
rect 204 328 252 356
rect 280 328 328 356
rect 356 328 404 356
rect 432 328 480 356
rect 508 328 513 356
rect -513 280 513 328
rect -513 252 -508 280
rect -480 252 -432 280
rect -404 252 -356 280
rect -328 252 -280 280
rect -252 252 -204 280
rect -176 252 -128 280
rect -100 252 -52 280
rect -24 252 24 280
rect 52 252 100 280
rect 128 252 176 280
rect 204 252 252 280
rect 280 252 328 280
rect 356 252 404 280
rect 432 252 480 280
rect 508 252 513 280
rect -513 204 513 252
rect -513 176 -508 204
rect -480 176 -432 204
rect -404 176 -356 204
rect -328 176 -280 204
rect -252 176 -204 204
rect -176 176 -128 204
rect -100 176 -52 204
rect -24 176 24 204
rect 52 176 100 204
rect 128 176 176 204
rect 204 176 252 204
rect 280 176 328 204
rect 356 176 404 204
rect 432 176 480 204
rect 508 176 513 204
rect -513 128 513 176
rect -513 100 -508 128
rect -480 100 -432 128
rect -404 100 -356 128
rect -328 100 -280 128
rect -252 100 -204 128
rect -176 100 -128 128
rect -100 100 -52 128
rect -24 100 24 128
rect 52 100 100 128
rect 128 100 176 128
rect 204 100 252 128
rect 280 100 328 128
rect 356 100 404 128
rect 432 100 480 128
rect 508 100 513 128
rect -513 52 513 100
rect -513 24 -508 52
rect -480 24 -432 52
rect -404 24 -356 52
rect -328 24 -280 52
rect -252 24 -204 52
rect -176 24 -128 52
rect -100 24 -52 52
rect -24 24 24 52
rect 52 24 100 52
rect 128 24 176 52
rect 204 24 252 52
rect 280 24 328 52
rect 356 24 404 52
rect 432 24 480 52
rect 508 24 513 52
rect -513 -24 513 24
rect -513 -52 -508 -24
rect -480 -52 -432 -24
rect -404 -52 -356 -24
rect -328 -52 -280 -24
rect -252 -52 -204 -24
rect -176 -52 -128 -24
rect -100 -52 -52 -24
rect -24 -52 24 -24
rect 52 -52 100 -24
rect 128 -52 176 -24
rect 204 -52 252 -24
rect 280 -52 328 -24
rect 356 -52 404 -24
rect 432 -52 480 -24
rect 508 -52 513 -24
rect -513 -100 513 -52
rect -513 -128 -508 -100
rect -480 -128 -432 -100
rect -404 -128 -356 -100
rect -328 -128 -280 -100
rect -252 -128 -204 -100
rect -176 -128 -128 -100
rect -100 -128 -52 -100
rect -24 -128 24 -100
rect 52 -128 100 -100
rect 128 -128 176 -100
rect 204 -128 252 -100
rect 280 -128 328 -100
rect 356 -128 404 -100
rect 432 -128 480 -100
rect 508 -128 513 -100
rect -513 -176 513 -128
rect -513 -204 -508 -176
rect -480 -204 -432 -176
rect -404 -204 -356 -176
rect -328 -204 -280 -176
rect -252 -204 -204 -176
rect -176 -204 -128 -176
rect -100 -204 -52 -176
rect -24 -204 24 -176
rect 52 -204 100 -176
rect 128 -204 176 -176
rect 204 -204 252 -176
rect 280 -204 328 -176
rect 356 -204 404 -176
rect 432 -204 480 -176
rect 508 -204 513 -176
rect -513 -252 513 -204
rect -513 -280 -508 -252
rect -480 -280 -432 -252
rect -404 -280 -356 -252
rect -328 -280 -280 -252
rect -252 -280 -204 -252
rect -176 -280 -128 -252
rect -100 -280 -52 -252
rect -24 -280 24 -252
rect 52 -280 100 -252
rect 128 -280 176 -252
rect 204 -280 252 -252
rect 280 -280 328 -252
rect 356 -280 404 -252
rect 432 -280 480 -252
rect 508 -280 513 -252
rect -513 -328 513 -280
rect -513 -356 -508 -328
rect -480 -356 -432 -328
rect -404 -356 -356 -328
rect -328 -356 -280 -328
rect -252 -356 -204 -328
rect -176 -356 -128 -328
rect -100 -356 -52 -328
rect -24 -356 24 -328
rect 52 -356 100 -328
rect 128 -356 176 -328
rect 204 -356 252 -328
rect 280 -356 328 -328
rect 356 -356 404 -328
rect 432 -356 480 -328
rect 508 -356 513 -328
rect -513 -404 513 -356
rect -513 -432 -508 -404
rect -480 -432 -432 -404
rect -404 -432 -356 -404
rect -328 -432 -280 -404
rect -252 -432 -204 -404
rect -176 -432 -128 -404
rect -100 -432 -52 -404
rect -24 -432 24 -404
rect 52 -432 100 -404
rect 128 -432 176 -404
rect 204 -432 252 -404
rect 280 -432 328 -404
rect 356 -432 404 -404
rect 432 -432 480 -404
rect 508 -432 513 -404
rect -513 -480 513 -432
rect -513 -508 -508 -480
rect -480 -508 -432 -480
rect -404 -508 -356 -480
rect -328 -508 -280 -480
rect -252 -508 -204 -480
rect -176 -508 -128 -480
rect -100 -508 -52 -480
rect -24 -508 24 -480
rect 52 -508 100 -480
rect 128 -508 176 -480
rect 204 -508 252 -480
rect 280 -508 328 -480
rect 356 -508 404 -480
rect 432 -508 480 -480
rect 508 -508 513 -480
rect -513 -556 513 -508
rect -513 -584 -508 -556
rect -480 -584 -432 -556
rect -404 -584 -356 -556
rect -328 -584 -280 -556
rect -252 -584 -204 -556
rect -176 -584 -128 -556
rect -100 -584 -52 -556
rect -24 -584 24 -556
rect 52 -584 100 -556
rect 128 -584 176 -556
rect 204 -584 252 -556
rect 280 -584 328 -556
rect 356 -584 404 -556
rect 432 -584 480 -556
rect 508 -584 513 -556
rect -513 -632 513 -584
rect -513 -660 -508 -632
rect -480 -660 -432 -632
rect -404 -660 -356 -632
rect -328 -660 -280 -632
rect -252 -660 -204 -632
rect -176 -660 -128 -632
rect -100 -660 -52 -632
rect -24 -660 24 -632
rect 52 -660 100 -632
rect 128 -660 176 -632
rect 204 -660 252 -632
rect 280 -660 328 -632
rect 356 -660 404 -632
rect 432 -660 480 -632
rect 508 -660 513 -632
rect -513 -708 513 -660
rect -513 -736 -508 -708
rect -480 -736 -432 -708
rect -404 -736 -356 -708
rect -328 -736 -280 -708
rect -252 -736 -204 -708
rect -176 -736 -128 -708
rect -100 -736 -52 -708
rect -24 -736 24 -708
rect 52 -736 100 -708
rect 128 -736 176 -708
rect 204 -736 252 -708
rect 280 -736 328 -708
rect 356 -736 404 -708
rect 432 -736 480 -708
rect 508 -736 513 -708
rect -513 -784 513 -736
rect -513 -812 -508 -784
rect -480 -812 -432 -784
rect -404 -812 -356 -784
rect -328 -812 -280 -784
rect -252 -812 -204 -784
rect -176 -812 -128 -784
rect -100 -812 -52 -784
rect -24 -812 24 -784
rect 52 -812 100 -784
rect 128 -812 176 -784
rect 204 -812 252 -784
rect 280 -812 328 -784
rect 356 -812 404 -784
rect 432 -812 480 -784
rect 508 -812 513 -784
rect -513 -860 513 -812
rect -513 -888 -508 -860
rect -480 -888 -432 -860
rect -404 -888 -356 -860
rect -328 -888 -280 -860
rect -252 -888 -204 -860
rect -176 -888 -128 -860
rect -100 -888 -52 -860
rect -24 -888 24 -860
rect 52 -888 100 -860
rect 128 -888 176 -860
rect 204 -888 252 -860
rect 280 -888 328 -860
rect 356 -888 404 -860
rect 432 -888 480 -860
rect 508 -888 513 -860
rect -513 -936 513 -888
rect -513 -964 -508 -936
rect -480 -964 -432 -936
rect -404 -964 -356 -936
rect -328 -964 -280 -936
rect -252 -964 -204 -936
rect -176 -964 -128 -936
rect -100 -964 -52 -936
rect -24 -964 24 -936
rect 52 -964 100 -936
rect 128 -964 176 -936
rect 204 -964 252 -936
rect 280 -964 328 -936
rect 356 -964 404 -936
rect 432 -964 480 -936
rect 508 -964 513 -936
rect -513 -1012 513 -964
rect -513 -1040 -508 -1012
rect -480 -1040 -432 -1012
rect -404 -1040 -356 -1012
rect -328 -1040 -280 -1012
rect -252 -1040 -204 -1012
rect -176 -1040 -128 -1012
rect -100 -1040 -52 -1012
rect -24 -1040 24 -1012
rect 52 -1040 100 -1012
rect 128 -1040 176 -1012
rect 204 -1040 252 -1012
rect 280 -1040 328 -1012
rect 356 -1040 404 -1012
rect 432 -1040 480 -1012
rect 508 -1040 513 -1012
rect -513 -1088 513 -1040
rect -513 -1116 -508 -1088
rect -480 -1116 -432 -1088
rect -404 -1116 -356 -1088
rect -328 -1116 -280 -1088
rect -252 -1116 -204 -1088
rect -176 -1116 -128 -1088
rect -100 -1116 -52 -1088
rect -24 -1116 24 -1088
rect 52 -1116 100 -1088
rect 128 -1116 176 -1088
rect 204 -1116 252 -1088
rect 280 -1116 328 -1088
rect 356 -1116 404 -1088
rect 432 -1116 480 -1088
rect 508 -1116 513 -1088
rect -513 -1164 513 -1116
rect -513 -1192 -508 -1164
rect -480 -1192 -432 -1164
rect -404 -1192 -356 -1164
rect -328 -1192 -280 -1164
rect -252 -1192 -204 -1164
rect -176 -1192 -128 -1164
rect -100 -1192 -52 -1164
rect -24 -1192 24 -1164
rect 52 -1192 100 -1164
rect 128 -1192 176 -1164
rect 204 -1192 252 -1164
rect 280 -1192 328 -1164
rect 356 -1192 404 -1164
rect 432 -1192 480 -1164
rect 508 -1192 513 -1164
rect -513 -1240 513 -1192
rect -513 -1268 -508 -1240
rect -480 -1268 -432 -1240
rect -404 -1268 -356 -1240
rect -328 -1268 -280 -1240
rect -252 -1268 -204 -1240
rect -176 -1268 -128 -1240
rect -100 -1268 -52 -1240
rect -24 -1268 24 -1240
rect 52 -1268 100 -1240
rect 128 -1268 176 -1240
rect 204 -1268 252 -1240
rect 280 -1268 328 -1240
rect 356 -1268 404 -1240
rect 432 -1268 480 -1240
rect 508 -1268 513 -1240
rect -513 -1316 513 -1268
rect -513 -1344 -508 -1316
rect -480 -1344 -432 -1316
rect -404 -1344 -356 -1316
rect -328 -1344 -280 -1316
rect -252 -1344 -204 -1316
rect -176 -1344 -128 -1316
rect -100 -1344 -52 -1316
rect -24 -1344 24 -1316
rect 52 -1344 100 -1316
rect 128 -1344 176 -1316
rect 204 -1344 252 -1316
rect 280 -1344 328 -1316
rect 356 -1344 404 -1316
rect 432 -1344 480 -1316
rect 508 -1344 513 -1316
rect -513 -1392 513 -1344
rect -513 -1420 -508 -1392
rect -480 -1420 -432 -1392
rect -404 -1420 -356 -1392
rect -328 -1420 -280 -1392
rect -252 -1420 -204 -1392
rect -176 -1420 -128 -1392
rect -100 -1420 -52 -1392
rect -24 -1420 24 -1392
rect 52 -1420 100 -1392
rect 128 -1420 176 -1392
rect 204 -1420 252 -1392
rect 280 -1420 328 -1392
rect 356 -1420 404 -1392
rect 432 -1420 480 -1392
rect 508 -1420 513 -1392
rect -513 -1468 513 -1420
rect -513 -1496 -508 -1468
rect -480 -1496 -432 -1468
rect -404 -1496 -356 -1468
rect -328 -1496 -280 -1468
rect -252 -1496 -204 -1468
rect -176 -1496 -128 -1468
rect -100 -1496 -52 -1468
rect -24 -1496 24 -1468
rect 52 -1496 100 -1468
rect 128 -1496 176 -1468
rect 204 -1496 252 -1468
rect 280 -1496 328 -1468
rect 356 -1496 404 -1468
rect 432 -1496 480 -1468
rect 508 -1496 513 -1468
rect -513 -1544 513 -1496
rect -513 -1572 -508 -1544
rect -480 -1572 -432 -1544
rect -404 -1572 -356 -1544
rect -328 -1572 -280 -1544
rect -252 -1572 -204 -1544
rect -176 -1572 -128 -1544
rect -100 -1572 -52 -1544
rect -24 -1572 24 -1544
rect 52 -1572 100 -1544
rect 128 -1572 176 -1544
rect 204 -1572 252 -1544
rect 280 -1572 328 -1544
rect 356 -1572 404 -1544
rect 432 -1572 480 -1544
rect 508 -1572 513 -1544
rect -513 -1620 513 -1572
rect -513 -1648 -508 -1620
rect -480 -1648 -432 -1620
rect -404 -1648 -356 -1620
rect -328 -1648 -280 -1620
rect -252 -1648 -204 -1620
rect -176 -1648 -128 -1620
rect -100 -1648 -52 -1620
rect -24 -1648 24 -1620
rect 52 -1648 100 -1620
rect 128 -1648 176 -1620
rect 204 -1648 252 -1620
rect 280 -1648 328 -1620
rect 356 -1648 404 -1620
rect 432 -1648 480 -1620
rect 508 -1648 513 -1620
rect -513 -1696 513 -1648
rect -513 -1724 -508 -1696
rect -480 -1724 -432 -1696
rect -404 -1724 -356 -1696
rect -328 -1724 -280 -1696
rect -252 -1724 -204 -1696
rect -176 -1724 -128 -1696
rect -100 -1724 -52 -1696
rect -24 -1724 24 -1696
rect 52 -1724 100 -1696
rect 128 -1724 176 -1696
rect 204 -1724 252 -1696
rect 280 -1724 328 -1696
rect 356 -1724 404 -1696
rect 432 -1724 480 -1696
rect 508 -1724 513 -1696
rect -513 -1772 513 -1724
rect -513 -1800 -508 -1772
rect -480 -1800 -432 -1772
rect -404 -1800 -356 -1772
rect -328 -1800 -280 -1772
rect -252 -1800 -204 -1772
rect -176 -1800 -128 -1772
rect -100 -1800 -52 -1772
rect -24 -1800 24 -1772
rect 52 -1800 100 -1772
rect 128 -1800 176 -1772
rect 204 -1800 252 -1772
rect 280 -1800 328 -1772
rect 356 -1800 404 -1772
rect 432 -1800 480 -1772
rect 508 -1800 513 -1772
rect -513 -1848 513 -1800
rect -513 -1876 -508 -1848
rect -480 -1876 -432 -1848
rect -404 -1876 -356 -1848
rect -328 -1876 -280 -1848
rect -252 -1876 -204 -1848
rect -176 -1876 -128 -1848
rect -100 -1876 -52 -1848
rect -24 -1876 24 -1848
rect 52 -1876 100 -1848
rect 128 -1876 176 -1848
rect 204 -1876 252 -1848
rect 280 -1876 328 -1848
rect 356 -1876 404 -1848
rect 432 -1876 480 -1848
rect 508 -1876 513 -1848
rect -513 -1924 513 -1876
rect -513 -1952 -508 -1924
rect -480 -1952 -432 -1924
rect -404 -1952 -356 -1924
rect -328 -1952 -280 -1924
rect -252 -1952 -204 -1924
rect -176 -1952 -128 -1924
rect -100 -1952 -52 -1924
rect -24 -1952 24 -1924
rect 52 -1952 100 -1924
rect 128 -1952 176 -1924
rect 204 -1952 252 -1924
rect 280 -1952 328 -1924
rect 356 -1952 404 -1924
rect 432 -1952 480 -1924
rect 508 -1952 513 -1924
rect -513 -2000 513 -1952
rect -513 -2028 -508 -2000
rect -480 -2028 -432 -2000
rect -404 -2028 -356 -2000
rect -328 -2028 -280 -2000
rect -252 -2028 -204 -2000
rect -176 -2028 -128 -2000
rect -100 -2028 -52 -2000
rect -24 -2028 24 -2000
rect 52 -2028 100 -2000
rect 128 -2028 176 -2000
rect 204 -2028 252 -2000
rect 280 -2028 328 -2000
rect 356 -2028 404 -2000
rect 432 -2028 480 -2000
rect 508 -2028 513 -2000
rect -513 -2076 513 -2028
rect -513 -2104 -508 -2076
rect -480 -2104 -432 -2076
rect -404 -2104 -356 -2076
rect -328 -2104 -280 -2076
rect -252 -2104 -204 -2076
rect -176 -2104 -128 -2076
rect -100 -2104 -52 -2076
rect -24 -2104 24 -2076
rect 52 -2104 100 -2076
rect 128 -2104 176 -2076
rect 204 -2104 252 -2076
rect 280 -2104 328 -2076
rect 356 -2104 404 -2076
rect 432 -2104 480 -2076
rect 508 -2104 513 -2076
rect -513 -2152 513 -2104
rect -513 -2180 -508 -2152
rect -480 -2180 -432 -2152
rect -404 -2180 -356 -2152
rect -328 -2180 -280 -2152
rect -252 -2180 -204 -2152
rect -176 -2180 -128 -2152
rect -100 -2180 -52 -2152
rect -24 -2180 24 -2152
rect 52 -2180 100 -2152
rect 128 -2180 176 -2152
rect 204 -2180 252 -2152
rect 280 -2180 328 -2152
rect 356 -2180 404 -2152
rect 432 -2180 480 -2152
rect 508 -2180 513 -2152
rect -513 -2228 513 -2180
rect -513 -2256 -508 -2228
rect -480 -2256 -432 -2228
rect -404 -2256 -356 -2228
rect -328 -2256 -280 -2228
rect -252 -2256 -204 -2228
rect -176 -2256 -128 -2228
rect -100 -2256 -52 -2228
rect -24 -2256 24 -2228
rect 52 -2256 100 -2228
rect 128 -2256 176 -2228
rect 204 -2256 252 -2228
rect 280 -2256 328 -2228
rect 356 -2256 404 -2228
rect 432 -2256 480 -2228
rect 508 -2256 513 -2228
rect -513 -2304 513 -2256
rect -513 -2332 -508 -2304
rect -480 -2332 -432 -2304
rect -404 -2332 -356 -2304
rect -328 -2332 -280 -2304
rect -252 -2332 -204 -2304
rect -176 -2332 -128 -2304
rect -100 -2332 -52 -2304
rect -24 -2332 24 -2304
rect 52 -2332 100 -2304
rect 128 -2332 176 -2304
rect 204 -2332 252 -2304
rect 280 -2332 328 -2304
rect 356 -2332 404 -2304
rect 432 -2332 480 -2304
rect 508 -2332 513 -2304
rect -513 -2380 513 -2332
rect -513 -2408 -508 -2380
rect -480 -2408 -432 -2380
rect -404 -2408 -356 -2380
rect -328 -2408 -280 -2380
rect -252 -2408 -204 -2380
rect -176 -2408 -128 -2380
rect -100 -2408 -52 -2380
rect -24 -2408 24 -2380
rect 52 -2408 100 -2380
rect 128 -2408 176 -2380
rect 204 -2408 252 -2380
rect 280 -2408 328 -2380
rect 356 -2408 404 -2380
rect 432 -2408 480 -2380
rect 508 -2408 513 -2380
rect -513 -2456 513 -2408
rect -513 -2484 -508 -2456
rect -480 -2484 -432 -2456
rect -404 -2484 -356 -2456
rect -328 -2484 -280 -2456
rect -252 -2484 -204 -2456
rect -176 -2484 -128 -2456
rect -100 -2484 -52 -2456
rect -24 -2484 24 -2456
rect 52 -2484 100 -2456
rect 128 -2484 176 -2456
rect 204 -2484 252 -2456
rect 280 -2484 328 -2456
rect 356 -2484 404 -2456
rect 432 -2484 480 -2456
rect 508 -2484 513 -2456
rect -513 -2532 513 -2484
rect -513 -2560 -508 -2532
rect -480 -2560 -432 -2532
rect -404 -2560 -356 -2532
rect -328 -2560 -280 -2532
rect -252 -2560 -204 -2532
rect -176 -2560 -128 -2532
rect -100 -2560 -52 -2532
rect -24 -2560 24 -2532
rect 52 -2560 100 -2532
rect 128 -2560 176 -2532
rect 204 -2560 252 -2532
rect 280 -2560 328 -2532
rect 356 -2560 404 -2532
rect 432 -2560 480 -2532
rect 508 -2560 513 -2532
rect -513 -2608 513 -2560
rect -513 -2636 -508 -2608
rect -480 -2636 -432 -2608
rect -404 -2636 -356 -2608
rect -328 -2636 -280 -2608
rect -252 -2636 -204 -2608
rect -176 -2636 -128 -2608
rect -100 -2636 -52 -2608
rect -24 -2636 24 -2608
rect 52 -2636 100 -2608
rect 128 -2636 176 -2608
rect 204 -2636 252 -2608
rect 280 -2636 328 -2608
rect 356 -2636 404 -2608
rect 432 -2636 480 -2608
rect 508 -2636 513 -2608
rect -513 -2641 513 -2636
<< via2 >>
rect -508 2608 -480 2636
rect -432 2608 -404 2636
rect -356 2608 -328 2636
rect -280 2608 -252 2636
rect -204 2608 -176 2636
rect -128 2608 -100 2636
rect -52 2608 -24 2636
rect 24 2608 52 2636
rect 100 2608 128 2636
rect 176 2608 204 2636
rect 252 2608 280 2636
rect 328 2608 356 2636
rect 404 2608 432 2636
rect 480 2608 508 2636
rect -508 2532 -480 2560
rect -432 2532 -404 2560
rect -356 2532 -328 2560
rect -280 2532 -252 2560
rect -204 2532 -176 2560
rect -128 2532 -100 2560
rect -52 2532 -24 2560
rect 24 2532 52 2560
rect 100 2532 128 2560
rect 176 2532 204 2560
rect 252 2532 280 2560
rect 328 2532 356 2560
rect 404 2532 432 2560
rect 480 2532 508 2560
rect -508 2456 -480 2484
rect -432 2456 -404 2484
rect -356 2456 -328 2484
rect -280 2456 -252 2484
rect -204 2456 -176 2484
rect -128 2456 -100 2484
rect -52 2456 -24 2484
rect 24 2456 52 2484
rect 100 2456 128 2484
rect 176 2456 204 2484
rect 252 2456 280 2484
rect 328 2456 356 2484
rect 404 2456 432 2484
rect 480 2456 508 2484
rect -508 2380 -480 2408
rect -432 2380 -404 2408
rect -356 2380 -328 2408
rect -280 2380 -252 2408
rect -204 2380 -176 2408
rect -128 2380 -100 2408
rect -52 2380 -24 2408
rect 24 2380 52 2408
rect 100 2380 128 2408
rect 176 2380 204 2408
rect 252 2380 280 2408
rect 328 2380 356 2408
rect 404 2380 432 2408
rect 480 2380 508 2408
rect -508 2304 -480 2332
rect -432 2304 -404 2332
rect -356 2304 -328 2332
rect -280 2304 -252 2332
rect -204 2304 -176 2332
rect -128 2304 -100 2332
rect -52 2304 -24 2332
rect 24 2304 52 2332
rect 100 2304 128 2332
rect 176 2304 204 2332
rect 252 2304 280 2332
rect 328 2304 356 2332
rect 404 2304 432 2332
rect 480 2304 508 2332
rect -508 2228 -480 2256
rect -432 2228 -404 2256
rect -356 2228 -328 2256
rect -280 2228 -252 2256
rect -204 2228 -176 2256
rect -128 2228 -100 2256
rect -52 2228 -24 2256
rect 24 2228 52 2256
rect 100 2228 128 2256
rect 176 2228 204 2256
rect 252 2228 280 2256
rect 328 2228 356 2256
rect 404 2228 432 2256
rect 480 2228 508 2256
rect -508 2152 -480 2180
rect -432 2152 -404 2180
rect -356 2152 -328 2180
rect -280 2152 -252 2180
rect -204 2152 -176 2180
rect -128 2152 -100 2180
rect -52 2152 -24 2180
rect 24 2152 52 2180
rect 100 2152 128 2180
rect 176 2152 204 2180
rect 252 2152 280 2180
rect 328 2152 356 2180
rect 404 2152 432 2180
rect 480 2152 508 2180
rect -508 2076 -480 2104
rect -432 2076 -404 2104
rect -356 2076 -328 2104
rect -280 2076 -252 2104
rect -204 2076 -176 2104
rect -128 2076 -100 2104
rect -52 2076 -24 2104
rect 24 2076 52 2104
rect 100 2076 128 2104
rect 176 2076 204 2104
rect 252 2076 280 2104
rect 328 2076 356 2104
rect 404 2076 432 2104
rect 480 2076 508 2104
rect -508 2000 -480 2028
rect -432 2000 -404 2028
rect -356 2000 -328 2028
rect -280 2000 -252 2028
rect -204 2000 -176 2028
rect -128 2000 -100 2028
rect -52 2000 -24 2028
rect 24 2000 52 2028
rect 100 2000 128 2028
rect 176 2000 204 2028
rect 252 2000 280 2028
rect 328 2000 356 2028
rect 404 2000 432 2028
rect 480 2000 508 2028
rect -508 1924 -480 1952
rect -432 1924 -404 1952
rect -356 1924 -328 1952
rect -280 1924 -252 1952
rect -204 1924 -176 1952
rect -128 1924 -100 1952
rect -52 1924 -24 1952
rect 24 1924 52 1952
rect 100 1924 128 1952
rect 176 1924 204 1952
rect 252 1924 280 1952
rect 328 1924 356 1952
rect 404 1924 432 1952
rect 480 1924 508 1952
rect -508 1848 -480 1876
rect -432 1848 -404 1876
rect -356 1848 -328 1876
rect -280 1848 -252 1876
rect -204 1848 -176 1876
rect -128 1848 -100 1876
rect -52 1848 -24 1876
rect 24 1848 52 1876
rect 100 1848 128 1876
rect 176 1848 204 1876
rect 252 1848 280 1876
rect 328 1848 356 1876
rect 404 1848 432 1876
rect 480 1848 508 1876
rect -508 1772 -480 1800
rect -432 1772 -404 1800
rect -356 1772 -328 1800
rect -280 1772 -252 1800
rect -204 1772 -176 1800
rect -128 1772 -100 1800
rect -52 1772 -24 1800
rect 24 1772 52 1800
rect 100 1772 128 1800
rect 176 1772 204 1800
rect 252 1772 280 1800
rect 328 1772 356 1800
rect 404 1772 432 1800
rect 480 1772 508 1800
rect -508 1696 -480 1724
rect -432 1696 -404 1724
rect -356 1696 -328 1724
rect -280 1696 -252 1724
rect -204 1696 -176 1724
rect -128 1696 -100 1724
rect -52 1696 -24 1724
rect 24 1696 52 1724
rect 100 1696 128 1724
rect 176 1696 204 1724
rect 252 1696 280 1724
rect 328 1696 356 1724
rect 404 1696 432 1724
rect 480 1696 508 1724
rect -508 1620 -480 1648
rect -432 1620 -404 1648
rect -356 1620 -328 1648
rect -280 1620 -252 1648
rect -204 1620 -176 1648
rect -128 1620 -100 1648
rect -52 1620 -24 1648
rect 24 1620 52 1648
rect 100 1620 128 1648
rect 176 1620 204 1648
rect 252 1620 280 1648
rect 328 1620 356 1648
rect 404 1620 432 1648
rect 480 1620 508 1648
rect -508 1544 -480 1572
rect -432 1544 -404 1572
rect -356 1544 -328 1572
rect -280 1544 -252 1572
rect -204 1544 -176 1572
rect -128 1544 -100 1572
rect -52 1544 -24 1572
rect 24 1544 52 1572
rect 100 1544 128 1572
rect 176 1544 204 1572
rect 252 1544 280 1572
rect 328 1544 356 1572
rect 404 1544 432 1572
rect 480 1544 508 1572
rect -508 1468 -480 1496
rect -432 1468 -404 1496
rect -356 1468 -328 1496
rect -280 1468 -252 1496
rect -204 1468 -176 1496
rect -128 1468 -100 1496
rect -52 1468 -24 1496
rect 24 1468 52 1496
rect 100 1468 128 1496
rect 176 1468 204 1496
rect 252 1468 280 1496
rect 328 1468 356 1496
rect 404 1468 432 1496
rect 480 1468 508 1496
rect -508 1392 -480 1420
rect -432 1392 -404 1420
rect -356 1392 -328 1420
rect -280 1392 -252 1420
rect -204 1392 -176 1420
rect -128 1392 -100 1420
rect -52 1392 -24 1420
rect 24 1392 52 1420
rect 100 1392 128 1420
rect 176 1392 204 1420
rect 252 1392 280 1420
rect 328 1392 356 1420
rect 404 1392 432 1420
rect 480 1392 508 1420
rect -508 1316 -480 1344
rect -432 1316 -404 1344
rect -356 1316 -328 1344
rect -280 1316 -252 1344
rect -204 1316 -176 1344
rect -128 1316 -100 1344
rect -52 1316 -24 1344
rect 24 1316 52 1344
rect 100 1316 128 1344
rect 176 1316 204 1344
rect 252 1316 280 1344
rect 328 1316 356 1344
rect 404 1316 432 1344
rect 480 1316 508 1344
rect -508 1240 -480 1268
rect -432 1240 -404 1268
rect -356 1240 -328 1268
rect -280 1240 -252 1268
rect -204 1240 -176 1268
rect -128 1240 -100 1268
rect -52 1240 -24 1268
rect 24 1240 52 1268
rect 100 1240 128 1268
rect 176 1240 204 1268
rect 252 1240 280 1268
rect 328 1240 356 1268
rect 404 1240 432 1268
rect 480 1240 508 1268
rect -508 1164 -480 1192
rect -432 1164 -404 1192
rect -356 1164 -328 1192
rect -280 1164 -252 1192
rect -204 1164 -176 1192
rect -128 1164 -100 1192
rect -52 1164 -24 1192
rect 24 1164 52 1192
rect 100 1164 128 1192
rect 176 1164 204 1192
rect 252 1164 280 1192
rect 328 1164 356 1192
rect 404 1164 432 1192
rect 480 1164 508 1192
rect -508 1088 -480 1116
rect -432 1088 -404 1116
rect -356 1088 -328 1116
rect -280 1088 -252 1116
rect -204 1088 -176 1116
rect -128 1088 -100 1116
rect -52 1088 -24 1116
rect 24 1088 52 1116
rect 100 1088 128 1116
rect 176 1088 204 1116
rect 252 1088 280 1116
rect 328 1088 356 1116
rect 404 1088 432 1116
rect 480 1088 508 1116
rect -508 1012 -480 1040
rect -432 1012 -404 1040
rect -356 1012 -328 1040
rect -280 1012 -252 1040
rect -204 1012 -176 1040
rect -128 1012 -100 1040
rect -52 1012 -24 1040
rect 24 1012 52 1040
rect 100 1012 128 1040
rect 176 1012 204 1040
rect 252 1012 280 1040
rect 328 1012 356 1040
rect 404 1012 432 1040
rect 480 1012 508 1040
rect -508 936 -480 964
rect -432 936 -404 964
rect -356 936 -328 964
rect -280 936 -252 964
rect -204 936 -176 964
rect -128 936 -100 964
rect -52 936 -24 964
rect 24 936 52 964
rect 100 936 128 964
rect 176 936 204 964
rect 252 936 280 964
rect 328 936 356 964
rect 404 936 432 964
rect 480 936 508 964
rect -508 860 -480 888
rect -432 860 -404 888
rect -356 860 -328 888
rect -280 860 -252 888
rect -204 860 -176 888
rect -128 860 -100 888
rect -52 860 -24 888
rect 24 860 52 888
rect 100 860 128 888
rect 176 860 204 888
rect 252 860 280 888
rect 328 860 356 888
rect 404 860 432 888
rect 480 860 508 888
rect -508 784 -480 812
rect -432 784 -404 812
rect -356 784 -328 812
rect -280 784 -252 812
rect -204 784 -176 812
rect -128 784 -100 812
rect -52 784 -24 812
rect 24 784 52 812
rect 100 784 128 812
rect 176 784 204 812
rect 252 784 280 812
rect 328 784 356 812
rect 404 784 432 812
rect 480 784 508 812
rect -508 708 -480 736
rect -432 708 -404 736
rect -356 708 -328 736
rect -280 708 -252 736
rect -204 708 -176 736
rect -128 708 -100 736
rect -52 708 -24 736
rect 24 708 52 736
rect 100 708 128 736
rect 176 708 204 736
rect 252 708 280 736
rect 328 708 356 736
rect 404 708 432 736
rect 480 708 508 736
rect -508 632 -480 660
rect -432 632 -404 660
rect -356 632 -328 660
rect -280 632 -252 660
rect -204 632 -176 660
rect -128 632 -100 660
rect -52 632 -24 660
rect 24 632 52 660
rect 100 632 128 660
rect 176 632 204 660
rect 252 632 280 660
rect 328 632 356 660
rect 404 632 432 660
rect 480 632 508 660
rect -508 556 -480 584
rect -432 556 -404 584
rect -356 556 -328 584
rect -280 556 -252 584
rect -204 556 -176 584
rect -128 556 -100 584
rect -52 556 -24 584
rect 24 556 52 584
rect 100 556 128 584
rect 176 556 204 584
rect 252 556 280 584
rect 328 556 356 584
rect 404 556 432 584
rect 480 556 508 584
rect -508 480 -480 508
rect -432 480 -404 508
rect -356 480 -328 508
rect -280 480 -252 508
rect -204 480 -176 508
rect -128 480 -100 508
rect -52 480 -24 508
rect 24 480 52 508
rect 100 480 128 508
rect 176 480 204 508
rect 252 480 280 508
rect 328 480 356 508
rect 404 480 432 508
rect 480 480 508 508
rect -508 404 -480 432
rect -432 404 -404 432
rect -356 404 -328 432
rect -280 404 -252 432
rect -204 404 -176 432
rect -128 404 -100 432
rect -52 404 -24 432
rect 24 404 52 432
rect 100 404 128 432
rect 176 404 204 432
rect 252 404 280 432
rect 328 404 356 432
rect 404 404 432 432
rect 480 404 508 432
rect -508 328 -480 356
rect -432 328 -404 356
rect -356 328 -328 356
rect -280 328 -252 356
rect -204 328 -176 356
rect -128 328 -100 356
rect -52 328 -24 356
rect 24 328 52 356
rect 100 328 128 356
rect 176 328 204 356
rect 252 328 280 356
rect 328 328 356 356
rect 404 328 432 356
rect 480 328 508 356
rect -508 252 -480 280
rect -432 252 -404 280
rect -356 252 -328 280
rect -280 252 -252 280
rect -204 252 -176 280
rect -128 252 -100 280
rect -52 252 -24 280
rect 24 252 52 280
rect 100 252 128 280
rect 176 252 204 280
rect 252 252 280 280
rect 328 252 356 280
rect 404 252 432 280
rect 480 252 508 280
rect -508 176 -480 204
rect -432 176 -404 204
rect -356 176 -328 204
rect -280 176 -252 204
rect -204 176 -176 204
rect -128 176 -100 204
rect -52 176 -24 204
rect 24 176 52 204
rect 100 176 128 204
rect 176 176 204 204
rect 252 176 280 204
rect 328 176 356 204
rect 404 176 432 204
rect 480 176 508 204
rect -508 100 -480 128
rect -432 100 -404 128
rect -356 100 -328 128
rect -280 100 -252 128
rect -204 100 -176 128
rect -128 100 -100 128
rect -52 100 -24 128
rect 24 100 52 128
rect 100 100 128 128
rect 176 100 204 128
rect 252 100 280 128
rect 328 100 356 128
rect 404 100 432 128
rect 480 100 508 128
rect -508 24 -480 52
rect -432 24 -404 52
rect -356 24 -328 52
rect -280 24 -252 52
rect -204 24 -176 52
rect -128 24 -100 52
rect -52 24 -24 52
rect 24 24 52 52
rect 100 24 128 52
rect 176 24 204 52
rect 252 24 280 52
rect 328 24 356 52
rect 404 24 432 52
rect 480 24 508 52
rect -508 -52 -480 -24
rect -432 -52 -404 -24
rect -356 -52 -328 -24
rect -280 -52 -252 -24
rect -204 -52 -176 -24
rect -128 -52 -100 -24
rect -52 -52 -24 -24
rect 24 -52 52 -24
rect 100 -52 128 -24
rect 176 -52 204 -24
rect 252 -52 280 -24
rect 328 -52 356 -24
rect 404 -52 432 -24
rect 480 -52 508 -24
rect -508 -128 -480 -100
rect -432 -128 -404 -100
rect -356 -128 -328 -100
rect -280 -128 -252 -100
rect -204 -128 -176 -100
rect -128 -128 -100 -100
rect -52 -128 -24 -100
rect 24 -128 52 -100
rect 100 -128 128 -100
rect 176 -128 204 -100
rect 252 -128 280 -100
rect 328 -128 356 -100
rect 404 -128 432 -100
rect 480 -128 508 -100
rect -508 -204 -480 -176
rect -432 -204 -404 -176
rect -356 -204 -328 -176
rect -280 -204 -252 -176
rect -204 -204 -176 -176
rect -128 -204 -100 -176
rect -52 -204 -24 -176
rect 24 -204 52 -176
rect 100 -204 128 -176
rect 176 -204 204 -176
rect 252 -204 280 -176
rect 328 -204 356 -176
rect 404 -204 432 -176
rect 480 -204 508 -176
rect -508 -280 -480 -252
rect -432 -280 -404 -252
rect -356 -280 -328 -252
rect -280 -280 -252 -252
rect -204 -280 -176 -252
rect -128 -280 -100 -252
rect -52 -280 -24 -252
rect 24 -280 52 -252
rect 100 -280 128 -252
rect 176 -280 204 -252
rect 252 -280 280 -252
rect 328 -280 356 -252
rect 404 -280 432 -252
rect 480 -280 508 -252
rect -508 -356 -480 -328
rect -432 -356 -404 -328
rect -356 -356 -328 -328
rect -280 -356 -252 -328
rect -204 -356 -176 -328
rect -128 -356 -100 -328
rect -52 -356 -24 -328
rect 24 -356 52 -328
rect 100 -356 128 -328
rect 176 -356 204 -328
rect 252 -356 280 -328
rect 328 -356 356 -328
rect 404 -356 432 -328
rect 480 -356 508 -328
rect -508 -432 -480 -404
rect -432 -432 -404 -404
rect -356 -432 -328 -404
rect -280 -432 -252 -404
rect -204 -432 -176 -404
rect -128 -432 -100 -404
rect -52 -432 -24 -404
rect 24 -432 52 -404
rect 100 -432 128 -404
rect 176 -432 204 -404
rect 252 -432 280 -404
rect 328 -432 356 -404
rect 404 -432 432 -404
rect 480 -432 508 -404
rect -508 -508 -480 -480
rect -432 -508 -404 -480
rect -356 -508 -328 -480
rect -280 -508 -252 -480
rect -204 -508 -176 -480
rect -128 -508 -100 -480
rect -52 -508 -24 -480
rect 24 -508 52 -480
rect 100 -508 128 -480
rect 176 -508 204 -480
rect 252 -508 280 -480
rect 328 -508 356 -480
rect 404 -508 432 -480
rect 480 -508 508 -480
rect -508 -584 -480 -556
rect -432 -584 -404 -556
rect -356 -584 -328 -556
rect -280 -584 -252 -556
rect -204 -584 -176 -556
rect -128 -584 -100 -556
rect -52 -584 -24 -556
rect 24 -584 52 -556
rect 100 -584 128 -556
rect 176 -584 204 -556
rect 252 -584 280 -556
rect 328 -584 356 -556
rect 404 -584 432 -556
rect 480 -584 508 -556
rect -508 -660 -480 -632
rect -432 -660 -404 -632
rect -356 -660 -328 -632
rect -280 -660 -252 -632
rect -204 -660 -176 -632
rect -128 -660 -100 -632
rect -52 -660 -24 -632
rect 24 -660 52 -632
rect 100 -660 128 -632
rect 176 -660 204 -632
rect 252 -660 280 -632
rect 328 -660 356 -632
rect 404 -660 432 -632
rect 480 -660 508 -632
rect -508 -736 -480 -708
rect -432 -736 -404 -708
rect -356 -736 -328 -708
rect -280 -736 -252 -708
rect -204 -736 -176 -708
rect -128 -736 -100 -708
rect -52 -736 -24 -708
rect 24 -736 52 -708
rect 100 -736 128 -708
rect 176 -736 204 -708
rect 252 -736 280 -708
rect 328 -736 356 -708
rect 404 -736 432 -708
rect 480 -736 508 -708
rect -508 -812 -480 -784
rect -432 -812 -404 -784
rect -356 -812 -328 -784
rect -280 -812 -252 -784
rect -204 -812 -176 -784
rect -128 -812 -100 -784
rect -52 -812 -24 -784
rect 24 -812 52 -784
rect 100 -812 128 -784
rect 176 -812 204 -784
rect 252 -812 280 -784
rect 328 -812 356 -784
rect 404 -812 432 -784
rect 480 -812 508 -784
rect -508 -888 -480 -860
rect -432 -888 -404 -860
rect -356 -888 -328 -860
rect -280 -888 -252 -860
rect -204 -888 -176 -860
rect -128 -888 -100 -860
rect -52 -888 -24 -860
rect 24 -888 52 -860
rect 100 -888 128 -860
rect 176 -888 204 -860
rect 252 -888 280 -860
rect 328 -888 356 -860
rect 404 -888 432 -860
rect 480 -888 508 -860
rect -508 -964 -480 -936
rect -432 -964 -404 -936
rect -356 -964 -328 -936
rect -280 -964 -252 -936
rect -204 -964 -176 -936
rect -128 -964 -100 -936
rect -52 -964 -24 -936
rect 24 -964 52 -936
rect 100 -964 128 -936
rect 176 -964 204 -936
rect 252 -964 280 -936
rect 328 -964 356 -936
rect 404 -964 432 -936
rect 480 -964 508 -936
rect -508 -1040 -480 -1012
rect -432 -1040 -404 -1012
rect -356 -1040 -328 -1012
rect -280 -1040 -252 -1012
rect -204 -1040 -176 -1012
rect -128 -1040 -100 -1012
rect -52 -1040 -24 -1012
rect 24 -1040 52 -1012
rect 100 -1040 128 -1012
rect 176 -1040 204 -1012
rect 252 -1040 280 -1012
rect 328 -1040 356 -1012
rect 404 -1040 432 -1012
rect 480 -1040 508 -1012
rect -508 -1116 -480 -1088
rect -432 -1116 -404 -1088
rect -356 -1116 -328 -1088
rect -280 -1116 -252 -1088
rect -204 -1116 -176 -1088
rect -128 -1116 -100 -1088
rect -52 -1116 -24 -1088
rect 24 -1116 52 -1088
rect 100 -1116 128 -1088
rect 176 -1116 204 -1088
rect 252 -1116 280 -1088
rect 328 -1116 356 -1088
rect 404 -1116 432 -1088
rect 480 -1116 508 -1088
rect -508 -1192 -480 -1164
rect -432 -1192 -404 -1164
rect -356 -1192 -328 -1164
rect -280 -1192 -252 -1164
rect -204 -1192 -176 -1164
rect -128 -1192 -100 -1164
rect -52 -1192 -24 -1164
rect 24 -1192 52 -1164
rect 100 -1192 128 -1164
rect 176 -1192 204 -1164
rect 252 -1192 280 -1164
rect 328 -1192 356 -1164
rect 404 -1192 432 -1164
rect 480 -1192 508 -1164
rect -508 -1268 -480 -1240
rect -432 -1268 -404 -1240
rect -356 -1268 -328 -1240
rect -280 -1268 -252 -1240
rect -204 -1268 -176 -1240
rect -128 -1268 -100 -1240
rect -52 -1268 -24 -1240
rect 24 -1268 52 -1240
rect 100 -1268 128 -1240
rect 176 -1268 204 -1240
rect 252 -1268 280 -1240
rect 328 -1268 356 -1240
rect 404 -1268 432 -1240
rect 480 -1268 508 -1240
rect -508 -1344 -480 -1316
rect -432 -1344 -404 -1316
rect -356 -1344 -328 -1316
rect -280 -1344 -252 -1316
rect -204 -1344 -176 -1316
rect -128 -1344 -100 -1316
rect -52 -1344 -24 -1316
rect 24 -1344 52 -1316
rect 100 -1344 128 -1316
rect 176 -1344 204 -1316
rect 252 -1344 280 -1316
rect 328 -1344 356 -1316
rect 404 -1344 432 -1316
rect 480 -1344 508 -1316
rect -508 -1420 -480 -1392
rect -432 -1420 -404 -1392
rect -356 -1420 -328 -1392
rect -280 -1420 -252 -1392
rect -204 -1420 -176 -1392
rect -128 -1420 -100 -1392
rect -52 -1420 -24 -1392
rect 24 -1420 52 -1392
rect 100 -1420 128 -1392
rect 176 -1420 204 -1392
rect 252 -1420 280 -1392
rect 328 -1420 356 -1392
rect 404 -1420 432 -1392
rect 480 -1420 508 -1392
rect -508 -1496 -480 -1468
rect -432 -1496 -404 -1468
rect -356 -1496 -328 -1468
rect -280 -1496 -252 -1468
rect -204 -1496 -176 -1468
rect -128 -1496 -100 -1468
rect -52 -1496 -24 -1468
rect 24 -1496 52 -1468
rect 100 -1496 128 -1468
rect 176 -1496 204 -1468
rect 252 -1496 280 -1468
rect 328 -1496 356 -1468
rect 404 -1496 432 -1468
rect 480 -1496 508 -1468
rect -508 -1572 -480 -1544
rect -432 -1572 -404 -1544
rect -356 -1572 -328 -1544
rect -280 -1572 -252 -1544
rect -204 -1572 -176 -1544
rect -128 -1572 -100 -1544
rect -52 -1572 -24 -1544
rect 24 -1572 52 -1544
rect 100 -1572 128 -1544
rect 176 -1572 204 -1544
rect 252 -1572 280 -1544
rect 328 -1572 356 -1544
rect 404 -1572 432 -1544
rect 480 -1572 508 -1544
rect -508 -1648 -480 -1620
rect -432 -1648 -404 -1620
rect -356 -1648 -328 -1620
rect -280 -1648 -252 -1620
rect -204 -1648 -176 -1620
rect -128 -1648 -100 -1620
rect -52 -1648 -24 -1620
rect 24 -1648 52 -1620
rect 100 -1648 128 -1620
rect 176 -1648 204 -1620
rect 252 -1648 280 -1620
rect 328 -1648 356 -1620
rect 404 -1648 432 -1620
rect 480 -1648 508 -1620
rect -508 -1724 -480 -1696
rect -432 -1724 -404 -1696
rect -356 -1724 -328 -1696
rect -280 -1724 -252 -1696
rect -204 -1724 -176 -1696
rect -128 -1724 -100 -1696
rect -52 -1724 -24 -1696
rect 24 -1724 52 -1696
rect 100 -1724 128 -1696
rect 176 -1724 204 -1696
rect 252 -1724 280 -1696
rect 328 -1724 356 -1696
rect 404 -1724 432 -1696
rect 480 -1724 508 -1696
rect -508 -1800 -480 -1772
rect -432 -1800 -404 -1772
rect -356 -1800 -328 -1772
rect -280 -1800 -252 -1772
rect -204 -1800 -176 -1772
rect -128 -1800 -100 -1772
rect -52 -1800 -24 -1772
rect 24 -1800 52 -1772
rect 100 -1800 128 -1772
rect 176 -1800 204 -1772
rect 252 -1800 280 -1772
rect 328 -1800 356 -1772
rect 404 -1800 432 -1772
rect 480 -1800 508 -1772
rect -508 -1876 -480 -1848
rect -432 -1876 -404 -1848
rect -356 -1876 -328 -1848
rect -280 -1876 -252 -1848
rect -204 -1876 -176 -1848
rect -128 -1876 -100 -1848
rect -52 -1876 -24 -1848
rect 24 -1876 52 -1848
rect 100 -1876 128 -1848
rect 176 -1876 204 -1848
rect 252 -1876 280 -1848
rect 328 -1876 356 -1848
rect 404 -1876 432 -1848
rect 480 -1876 508 -1848
rect -508 -1952 -480 -1924
rect -432 -1952 -404 -1924
rect -356 -1952 -328 -1924
rect -280 -1952 -252 -1924
rect -204 -1952 -176 -1924
rect -128 -1952 -100 -1924
rect -52 -1952 -24 -1924
rect 24 -1952 52 -1924
rect 100 -1952 128 -1924
rect 176 -1952 204 -1924
rect 252 -1952 280 -1924
rect 328 -1952 356 -1924
rect 404 -1952 432 -1924
rect 480 -1952 508 -1924
rect -508 -2028 -480 -2000
rect -432 -2028 -404 -2000
rect -356 -2028 -328 -2000
rect -280 -2028 -252 -2000
rect -204 -2028 -176 -2000
rect -128 -2028 -100 -2000
rect -52 -2028 -24 -2000
rect 24 -2028 52 -2000
rect 100 -2028 128 -2000
rect 176 -2028 204 -2000
rect 252 -2028 280 -2000
rect 328 -2028 356 -2000
rect 404 -2028 432 -2000
rect 480 -2028 508 -2000
rect -508 -2104 -480 -2076
rect -432 -2104 -404 -2076
rect -356 -2104 -328 -2076
rect -280 -2104 -252 -2076
rect -204 -2104 -176 -2076
rect -128 -2104 -100 -2076
rect -52 -2104 -24 -2076
rect 24 -2104 52 -2076
rect 100 -2104 128 -2076
rect 176 -2104 204 -2076
rect 252 -2104 280 -2076
rect 328 -2104 356 -2076
rect 404 -2104 432 -2076
rect 480 -2104 508 -2076
rect -508 -2180 -480 -2152
rect -432 -2180 -404 -2152
rect -356 -2180 -328 -2152
rect -280 -2180 -252 -2152
rect -204 -2180 -176 -2152
rect -128 -2180 -100 -2152
rect -52 -2180 -24 -2152
rect 24 -2180 52 -2152
rect 100 -2180 128 -2152
rect 176 -2180 204 -2152
rect 252 -2180 280 -2152
rect 328 -2180 356 -2152
rect 404 -2180 432 -2152
rect 480 -2180 508 -2152
rect -508 -2256 -480 -2228
rect -432 -2256 -404 -2228
rect -356 -2256 -328 -2228
rect -280 -2256 -252 -2228
rect -204 -2256 -176 -2228
rect -128 -2256 -100 -2228
rect -52 -2256 -24 -2228
rect 24 -2256 52 -2228
rect 100 -2256 128 -2228
rect 176 -2256 204 -2228
rect 252 -2256 280 -2228
rect 328 -2256 356 -2228
rect 404 -2256 432 -2228
rect 480 -2256 508 -2228
rect -508 -2332 -480 -2304
rect -432 -2332 -404 -2304
rect -356 -2332 -328 -2304
rect -280 -2332 -252 -2304
rect -204 -2332 -176 -2304
rect -128 -2332 -100 -2304
rect -52 -2332 -24 -2304
rect 24 -2332 52 -2304
rect 100 -2332 128 -2304
rect 176 -2332 204 -2304
rect 252 -2332 280 -2304
rect 328 -2332 356 -2304
rect 404 -2332 432 -2304
rect 480 -2332 508 -2304
rect -508 -2408 -480 -2380
rect -432 -2408 -404 -2380
rect -356 -2408 -328 -2380
rect -280 -2408 -252 -2380
rect -204 -2408 -176 -2380
rect -128 -2408 -100 -2380
rect -52 -2408 -24 -2380
rect 24 -2408 52 -2380
rect 100 -2408 128 -2380
rect 176 -2408 204 -2380
rect 252 -2408 280 -2380
rect 328 -2408 356 -2380
rect 404 -2408 432 -2380
rect 480 -2408 508 -2380
rect -508 -2484 -480 -2456
rect -432 -2484 -404 -2456
rect -356 -2484 -328 -2456
rect -280 -2484 -252 -2456
rect -204 -2484 -176 -2456
rect -128 -2484 -100 -2456
rect -52 -2484 -24 -2456
rect 24 -2484 52 -2456
rect 100 -2484 128 -2456
rect 176 -2484 204 -2456
rect 252 -2484 280 -2456
rect 328 -2484 356 -2456
rect 404 -2484 432 -2456
rect 480 -2484 508 -2456
rect -508 -2560 -480 -2532
rect -432 -2560 -404 -2532
rect -356 -2560 -328 -2532
rect -280 -2560 -252 -2532
rect -204 -2560 -176 -2532
rect -128 -2560 -100 -2532
rect -52 -2560 -24 -2532
rect 24 -2560 52 -2532
rect 100 -2560 128 -2532
rect 176 -2560 204 -2532
rect 252 -2560 280 -2532
rect 328 -2560 356 -2532
rect 404 -2560 432 -2532
rect 480 -2560 508 -2532
rect -508 -2636 -480 -2608
rect -432 -2636 -404 -2608
rect -356 -2636 -328 -2608
rect -280 -2636 -252 -2608
rect -204 -2636 -176 -2608
rect -128 -2636 -100 -2608
rect -52 -2636 -24 -2608
rect 24 -2636 52 -2608
rect 100 -2636 128 -2608
rect 176 -2636 204 -2608
rect 252 -2636 280 -2608
rect 328 -2636 356 -2608
rect 404 -2636 432 -2608
rect 480 -2636 508 -2608
<< metal3 >>
rect -513 2636 513 2641
rect -513 2608 -508 2636
rect -480 2608 -432 2636
rect -404 2608 -356 2636
rect -328 2608 -280 2636
rect -252 2608 -204 2636
rect -176 2608 -128 2636
rect -100 2608 -52 2636
rect -24 2608 24 2636
rect 52 2608 100 2636
rect 128 2608 176 2636
rect 204 2608 252 2636
rect 280 2608 328 2636
rect 356 2608 404 2636
rect 432 2608 480 2636
rect 508 2608 513 2636
rect -513 2560 513 2608
rect -513 2532 -508 2560
rect -480 2532 -432 2560
rect -404 2532 -356 2560
rect -328 2532 -280 2560
rect -252 2532 -204 2560
rect -176 2532 -128 2560
rect -100 2532 -52 2560
rect -24 2532 24 2560
rect 52 2532 100 2560
rect 128 2532 176 2560
rect 204 2532 252 2560
rect 280 2532 328 2560
rect 356 2532 404 2560
rect 432 2532 480 2560
rect 508 2532 513 2560
rect -513 2484 513 2532
rect -513 2456 -508 2484
rect -480 2456 -432 2484
rect -404 2456 -356 2484
rect -328 2456 -280 2484
rect -252 2456 -204 2484
rect -176 2456 -128 2484
rect -100 2456 -52 2484
rect -24 2456 24 2484
rect 52 2456 100 2484
rect 128 2456 176 2484
rect 204 2456 252 2484
rect 280 2456 328 2484
rect 356 2456 404 2484
rect 432 2456 480 2484
rect 508 2456 513 2484
rect -513 2408 513 2456
rect -513 2380 -508 2408
rect -480 2380 -432 2408
rect -404 2380 -356 2408
rect -328 2380 -280 2408
rect -252 2380 -204 2408
rect -176 2380 -128 2408
rect -100 2380 -52 2408
rect -24 2380 24 2408
rect 52 2380 100 2408
rect 128 2380 176 2408
rect 204 2380 252 2408
rect 280 2380 328 2408
rect 356 2380 404 2408
rect 432 2380 480 2408
rect 508 2380 513 2408
rect -513 2332 513 2380
rect -513 2304 -508 2332
rect -480 2304 -432 2332
rect -404 2304 -356 2332
rect -328 2304 -280 2332
rect -252 2304 -204 2332
rect -176 2304 -128 2332
rect -100 2304 -52 2332
rect -24 2304 24 2332
rect 52 2304 100 2332
rect 128 2304 176 2332
rect 204 2304 252 2332
rect 280 2304 328 2332
rect 356 2304 404 2332
rect 432 2304 480 2332
rect 508 2304 513 2332
rect -513 2256 513 2304
rect -513 2228 -508 2256
rect -480 2228 -432 2256
rect -404 2228 -356 2256
rect -328 2228 -280 2256
rect -252 2228 -204 2256
rect -176 2228 -128 2256
rect -100 2228 -52 2256
rect -24 2228 24 2256
rect 52 2228 100 2256
rect 128 2228 176 2256
rect 204 2228 252 2256
rect 280 2228 328 2256
rect 356 2228 404 2256
rect 432 2228 480 2256
rect 508 2228 513 2256
rect -513 2180 513 2228
rect -513 2152 -508 2180
rect -480 2152 -432 2180
rect -404 2152 -356 2180
rect -328 2152 -280 2180
rect -252 2152 -204 2180
rect -176 2152 -128 2180
rect -100 2152 -52 2180
rect -24 2152 24 2180
rect 52 2152 100 2180
rect 128 2152 176 2180
rect 204 2152 252 2180
rect 280 2152 328 2180
rect 356 2152 404 2180
rect 432 2152 480 2180
rect 508 2152 513 2180
rect -513 2104 513 2152
rect -513 2076 -508 2104
rect -480 2076 -432 2104
rect -404 2076 -356 2104
rect -328 2076 -280 2104
rect -252 2076 -204 2104
rect -176 2076 -128 2104
rect -100 2076 -52 2104
rect -24 2076 24 2104
rect 52 2076 100 2104
rect 128 2076 176 2104
rect 204 2076 252 2104
rect 280 2076 328 2104
rect 356 2076 404 2104
rect 432 2076 480 2104
rect 508 2076 513 2104
rect -513 2028 513 2076
rect -513 2000 -508 2028
rect -480 2000 -432 2028
rect -404 2000 -356 2028
rect -328 2000 -280 2028
rect -252 2000 -204 2028
rect -176 2000 -128 2028
rect -100 2000 -52 2028
rect -24 2000 24 2028
rect 52 2000 100 2028
rect 128 2000 176 2028
rect 204 2000 252 2028
rect 280 2000 328 2028
rect 356 2000 404 2028
rect 432 2000 480 2028
rect 508 2000 513 2028
rect -513 1952 513 2000
rect -513 1924 -508 1952
rect -480 1924 -432 1952
rect -404 1924 -356 1952
rect -328 1924 -280 1952
rect -252 1924 -204 1952
rect -176 1924 -128 1952
rect -100 1924 -52 1952
rect -24 1924 24 1952
rect 52 1924 100 1952
rect 128 1924 176 1952
rect 204 1924 252 1952
rect 280 1924 328 1952
rect 356 1924 404 1952
rect 432 1924 480 1952
rect 508 1924 513 1952
rect -513 1876 513 1924
rect -513 1848 -508 1876
rect -480 1848 -432 1876
rect -404 1848 -356 1876
rect -328 1848 -280 1876
rect -252 1848 -204 1876
rect -176 1848 -128 1876
rect -100 1848 -52 1876
rect -24 1848 24 1876
rect 52 1848 100 1876
rect 128 1848 176 1876
rect 204 1848 252 1876
rect 280 1848 328 1876
rect 356 1848 404 1876
rect 432 1848 480 1876
rect 508 1848 513 1876
rect -513 1800 513 1848
rect -513 1772 -508 1800
rect -480 1772 -432 1800
rect -404 1772 -356 1800
rect -328 1772 -280 1800
rect -252 1772 -204 1800
rect -176 1772 -128 1800
rect -100 1772 -52 1800
rect -24 1772 24 1800
rect 52 1772 100 1800
rect 128 1772 176 1800
rect 204 1772 252 1800
rect 280 1772 328 1800
rect 356 1772 404 1800
rect 432 1772 480 1800
rect 508 1772 513 1800
rect -513 1724 513 1772
rect -513 1696 -508 1724
rect -480 1696 -432 1724
rect -404 1696 -356 1724
rect -328 1696 -280 1724
rect -252 1696 -204 1724
rect -176 1696 -128 1724
rect -100 1696 -52 1724
rect -24 1696 24 1724
rect 52 1696 100 1724
rect 128 1696 176 1724
rect 204 1696 252 1724
rect 280 1696 328 1724
rect 356 1696 404 1724
rect 432 1696 480 1724
rect 508 1696 513 1724
rect -513 1648 513 1696
rect -513 1620 -508 1648
rect -480 1620 -432 1648
rect -404 1620 -356 1648
rect -328 1620 -280 1648
rect -252 1620 -204 1648
rect -176 1620 -128 1648
rect -100 1620 -52 1648
rect -24 1620 24 1648
rect 52 1620 100 1648
rect 128 1620 176 1648
rect 204 1620 252 1648
rect 280 1620 328 1648
rect 356 1620 404 1648
rect 432 1620 480 1648
rect 508 1620 513 1648
rect -513 1572 513 1620
rect -513 1544 -508 1572
rect -480 1544 -432 1572
rect -404 1544 -356 1572
rect -328 1544 -280 1572
rect -252 1544 -204 1572
rect -176 1544 -128 1572
rect -100 1544 -52 1572
rect -24 1544 24 1572
rect 52 1544 100 1572
rect 128 1544 176 1572
rect 204 1544 252 1572
rect 280 1544 328 1572
rect 356 1544 404 1572
rect 432 1544 480 1572
rect 508 1544 513 1572
rect -513 1496 513 1544
rect -513 1468 -508 1496
rect -480 1468 -432 1496
rect -404 1468 -356 1496
rect -328 1468 -280 1496
rect -252 1468 -204 1496
rect -176 1468 -128 1496
rect -100 1468 -52 1496
rect -24 1468 24 1496
rect 52 1468 100 1496
rect 128 1468 176 1496
rect 204 1468 252 1496
rect 280 1468 328 1496
rect 356 1468 404 1496
rect 432 1468 480 1496
rect 508 1468 513 1496
rect -513 1420 513 1468
rect -513 1392 -508 1420
rect -480 1392 -432 1420
rect -404 1392 -356 1420
rect -328 1392 -280 1420
rect -252 1392 -204 1420
rect -176 1392 -128 1420
rect -100 1392 -52 1420
rect -24 1392 24 1420
rect 52 1392 100 1420
rect 128 1392 176 1420
rect 204 1392 252 1420
rect 280 1392 328 1420
rect 356 1392 404 1420
rect 432 1392 480 1420
rect 508 1392 513 1420
rect -513 1344 513 1392
rect -513 1316 -508 1344
rect -480 1316 -432 1344
rect -404 1316 -356 1344
rect -328 1316 -280 1344
rect -252 1316 -204 1344
rect -176 1316 -128 1344
rect -100 1316 -52 1344
rect -24 1316 24 1344
rect 52 1316 100 1344
rect 128 1316 176 1344
rect 204 1316 252 1344
rect 280 1316 328 1344
rect 356 1316 404 1344
rect 432 1316 480 1344
rect 508 1316 513 1344
rect -513 1268 513 1316
rect -513 1240 -508 1268
rect -480 1240 -432 1268
rect -404 1240 -356 1268
rect -328 1240 -280 1268
rect -252 1240 -204 1268
rect -176 1240 -128 1268
rect -100 1240 -52 1268
rect -24 1240 24 1268
rect 52 1240 100 1268
rect 128 1240 176 1268
rect 204 1240 252 1268
rect 280 1240 328 1268
rect 356 1240 404 1268
rect 432 1240 480 1268
rect 508 1240 513 1268
rect -513 1192 513 1240
rect -513 1164 -508 1192
rect -480 1164 -432 1192
rect -404 1164 -356 1192
rect -328 1164 -280 1192
rect -252 1164 -204 1192
rect -176 1164 -128 1192
rect -100 1164 -52 1192
rect -24 1164 24 1192
rect 52 1164 100 1192
rect 128 1164 176 1192
rect 204 1164 252 1192
rect 280 1164 328 1192
rect 356 1164 404 1192
rect 432 1164 480 1192
rect 508 1164 513 1192
rect -513 1116 513 1164
rect -513 1088 -508 1116
rect -480 1088 -432 1116
rect -404 1088 -356 1116
rect -328 1088 -280 1116
rect -252 1088 -204 1116
rect -176 1088 -128 1116
rect -100 1088 -52 1116
rect -24 1088 24 1116
rect 52 1088 100 1116
rect 128 1088 176 1116
rect 204 1088 252 1116
rect 280 1088 328 1116
rect 356 1088 404 1116
rect 432 1088 480 1116
rect 508 1088 513 1116
rect -513 1040 513 1088
rect -513 1012 -508 1040
rect -480 1012 -432 1040
rect -404 1012 -356 1040
rect -328 1012 -280 1040
rect -252 1012 -204 1040
rect -176 1012 -128 1040
rect -100 1012 -52 1040
rect -24 1012 24 1040
rect 52 1012 100 1040
rect 128 1012 176 1040
rect 204 1012 252 1040
rect 280 1012 328 1040
rect 356 1012 404 1040
rect 432 1012 480 1040
rect 508 1012 513 1040
rect -513 964 513 1012
rect -513 936 -508 964
rect -480 936 -432 964
rect -404 936 -356 964
rect -328 936 -280 964
rect -252 936 -204 964
rect -176 936 -128 964
rect -100 936 -52 964
rect -24 936 24 964
rect 52 936 100 964
rect 128 936 176 964
rect 204 936 252 964
rect 280 936 328 964
rect 356 936 404 964
rect 432 936 480 964
rect 508 936 513 964
rect -513 888 513 936
rect -513 860 -508 888
rect -480 860 -432 888
rect -404 860 -356 888
rect -328 860 -280 888
rect -252 860 -204 888
rect -176 860 -128 888
rect -100 860 -52 888
rect -24 860 24 888
rect 52 860 100 888
rect 128 860 176 888
rect 204 860 252 888
rect 280 860 328 888
rect 356 860 404 888
rect 432 860 480 888
rect 508 860 513 888
rect -513 812 513 860
rect -513 784 -508 812
rect -480 784 -432 812
rect -404 784 -356 812
rect -328 784 -280 812
rect -252 784 -204 812
rect -176 784 -128 812
rect -100 784 -52 812
rect -24 784 24 812
rect 52 784 100 812
rect 128 784 176 812
rect 204 784 252 812
rect 280 784 328 812
rect 356 784 404 812
rect 432 784 480 812
rect 508 784 513 812
rect -513 736 513 784
rect -513 708 -508 736
rect -480 708 -432 736
rect -404 708 -356 736
rect -328 708 -280 736
rect -252 708 -204 736
rect -176 708 -128 736
rect -100 708 -52 736
rect -24 708 24 736
rect 52 708 100 736
rect 128 708 176 736
rect 204 708 252 736
rect 280 708 328 736
rect 356 708 404 736
rect 432 708 480 736
rect 508 708 513 736
rect -513 660 513 708
rect -513 632 -508 660
rect -480 632 -432 660
rect -404 632 -356 660
rect -328 632 -280 660
rect -252 632 -204 660
rect -176 632 -128 660
rect -100 632 -52 660
rect -24 632 24 660
rect 52 632 100 660
rect 128 632 176 660
rect 204 632 252 660
rect 280 632 328 660
rect 356 632 404 660
rect 432 632 480 660
rect 508 632 513 660
rect -513 584 513 632
rect -513 556 -508 584
rect -480 556 -432 584
rect -404 556 -356 584
rect -328 556 -280 584
rect -252 556 -204 584
rect -176 556 -128 584
rect -100 556 -52 584
rect -24 556 24 584
rect 52 556 100 584
rect 128 556 176 584
rect 204 556 252 584
rect 280 556 328 584
rect 356 556 404 584
rect 432 556 480 584
rect 508 556 513 584
rect -513 508 513 556
rect -513 480 -508 508
rect -480 480 -432 508
rect -404 480 -356 508
rect -328 480 -280 508
rect -252 480 -204 508
rect -176 480 -128 508
rect -100 480 -52 508
rect -24 480 24 508
rect 52 480 100 508
rect 128 480 176 508
rect 204 480 252 508
rect 280 480 328 508
rect 356 480 404 508
rect 432 480 480 508
rect 508 480 513 508
rect -513 432 513 480
rect -513 404 -508 432
rect -480 404 -432 432
rect -404 404 -356 432
rect -328 404 -280 432
rect -252 404 -204 432
rect -176 404 -128 432
rect -100 404 -52 432
rect -24 404 24 432
rect 52 404 100 432
rect 128 404 176 432
rect 204 404 252 432
rect 280 404 328 432
rect 356 404 404 432
rect 432 404 480 432
rect 508 404 513 432
rect -513 356 513 404
rect -513 328 -508 356
rect -480 328 -432 356
rect -404 328 -356 356
rect -328 328 -280 356
rect -252 328 -204 356
rect -176 328 -128 356
rect -100 328 -52 356
rect -24 328 24 356
rect 52 328 100 356
rect 128 328 176 356
rect 204 328 252 356
rect 280 328 328 356
rect 356 328 404 356
rect 432 328 480 356
rect 508 328 513 356
rect -513 280 513 328
rect -513 252 -508 280
rect -480 252 -432 280
rect -404 252 -356 280
rect -328 252 -280 280
rect -252 252 -204 280
rect -176 252 -128 280
rect -100 252 -52 280
rect -24 252 24 280
rect 52 252 100 280
rect 128 252 176 280
rect 204 252 252 280
rect 280 252 328 280
rect 356 252 404 280
rect 432 252 480 280
rect 508 252 513 280
rect -513 204 513 252
rect -513 176 -508 204
rect -480 176 -432 204
rect -404 176 -356 204
rect -328 176 -280 204
rect -252 176 -204 204
rect -176 176 -128 204
rect -100 176 -52 204
rect -24 176 24 204
rect 52 176 100 204
rect 128 176 176 204
rect 204 176 252 204
rect 280 176 328 204
rect 356 176 404 204
rect 432 176 480 204
rect 508 176 513 204
rect -513 128 513 176
rect -513 100 -508 128
rect -480 100 -432 128
rect -404 100 -356 128
rect -328 100 -280 128
rect -252 100 -204 128
rect -176 100 -128 128
rect -100 100 -52 128
rect -24 100 24 128
rect 52 100 100 128
rect 128 100 176 128
rect 204 100 252 128
rect 280 100 328 128
rect 356 100 404 128
rect 432 100 480 128
rect 508 100 513 128
rect -513 52 513 100
rect -513 24 -508 52
rect -480 24 -432 52
rect -404 24 -356 52
rect -328 24 -280 52
rect -252 24 -204 52
rect -176 24 -128 52
rect -100 24 -52 52
rect -24 24 24 52
rect 52 24 100 52
rect 128 24 176 52
rect 204 24 252 52
rect 280 24 328 52
rect 356 24 404 52
rect 432 24 480 52
rect 508 24 513 52
rect -513 -24 513 24
rect -513 -52 -508 -24
rect -480 -52 -432 -24
rect -404 -52 -356 -24
rect -328 -52 -280 -24
rect -252 -52 -204 -24
rect -176 -52 -128 -24
rect -100 -52 -52 -24
rect -24 -52 24 -24
rect 52 -52 100 -24
rect 128 -52 176 -24
rect 204 -52 252 -24
rect 280 -52 328 -24
rect 356 -52 404 -24
rect 432 -52 480 -24
rect 508 -52 513 -24
rect -513 -100 513 -52
rect -513 -128 -508 -100
rect -480 -128 -432 -100
rect -404 -128 -356 -100
rect -328 -128 -280 -100
rect -252 -128 -204 -100
rect -176 -128 -128 -100
rect -100 -128 -52 -100
rect -24 -128 24 -100
rect 52 -128 100 -100
rect 128 -128 176 -100
rect 204 -128 252 -100
rect 280 -128 328 -100
rect 356 -128 404 -100
rect 432 -128 480 -100
rect 508 -128 513 -100
rect -513 -176 513 -128
rect -513 -204 -508 -176
rect -480 -204 -432 -176
rect -404 -204 -356 -176
rect -328 -204 -280 -176
rect -252 -204 -204 -176
rect -176 -204 -128 -176
rect -100 -204 -52 -176
rect -24 -204 24 -176
rect 52 -204 100 -176
rect 128 -204 176 -176
rect 204 -204 252 -176
rect 280 -204 328 -176
rect 356 -204 404 -176
rect 432 -204 480 -176
rect 508 -204 513 -176
rect -513 -252 513 -204
rect -513 -280 -508 -252
rect -480 -280 -432 -252
rect -404 -280 -356 -252
rect -328 -280 -280 -252
rect -252 -280 -204 -252
rect -176 -280 -128 -252
rect -100 -280 -52 -252
rect -24 -280 24 -252
rect 52 -280 100 -252
rect 128 -280 176 -252
rect 204 -280 252 -252
rect 280 -280 328 -252
rect 356 -280 404 -252
rect 432 -280 480 -252
rect 508 -280 513 -252
rect -513 -328 513 -280
rect -513 -356 -508 -328
rect -480 -356 -432 -328
rect -404 -356 -356 -328
rect -328 -356 -280 -328
rect -252 -356 -204 -328
rect -176 -356 -128 -328
rect -100 -356 -52 -328
rect -24 -356 24 -328
rect 52 -356 100 -328
rect 128 -356 176 -328
rect 204 -356 252 -328
rect 280 -356 328 -328
rect 356 -356 404 -328
rect 432 -356 480 -328
rect 508 -356 513 -328
rect -513 -404 513 -356
rect -513 -432 -508 -404
rect -480 -432 -432 -404
rect -404 -432 -356 -404
rect -328 -432 -280 -404
rect -252 -432 -204 -404
rect -176 -432 -128 -404
rect -100 -432 -52 -404
rect -24 -432 24 -404
rect 52 -432 100 -404
rect 128 -432 176 -404
rect 204 -432 252 -404
rect 280 -432 328 -404
rect 356 -432 404 -404
rect 432 -432 480 -404
rect 508 -432 513 -404
rect -513 -480 513 -432
rect -513 -508 -508 -480
rect -480 -508 -432 -480
rect -404 -508 -356 -480
rect -328 -508 -280 -480
rect -252 -508 -204 -480
rect -176 -508 -128 -480
rect -100 -508 -52 -480
rect -24 -508 24 -480
rect 52 -508 100 -480
rect 128 -508 176 -480
rect 204 -508 252 -480
rect 280 -508 328 -480
rect 356 -508 404 -480
rect 432 -508 480 -480
rect 508 -508 513 -480
rect -513 -556 513 -508
rect -513 -584 -508 -556
rect -480 -584 -432 -556
rect -404 -584 -356 -556
rect -328 -584 -280 -556
rect -252 -584 -204 -556
rect -176 -584 -128 -556
rect -100 -584 -52 -556
rect -24 -584 24 -556
rect 52 -584 100 -556
rect 128 -584 176 -556
rect 204 -584 252 -556
rect 280 -584 328 -556
rect 356 -584 404 -556
rect 432 -584 480 -556
rect 508 -584 513 -556
rect -513 -632 513 -584
rect -513 -660 -508 -632
rect -480 -660 -432 -632
rect -404 -660 -356 -632
rect -328 -660 -280 -632
rect -252 -660 -204 -632
rect -176 -660 -128 -632
rect -100 -660 -52 -632
rect -24 -660 24 -632
rect 52 -660 100 -632
rect 128 -660 176 -632
rect 204 -660 252 -632
rect 280 -660 328 -632
rect 356 -660 404 -632
rect 432 -660 480 -632
rect 508 -660 513 -632
rect -513 -708 513 -660
rect -513 -736 -508 -708
rect -480 -736 -432 -708
rect -404 -736 -356 -708
rect -328 -736 -280 -708
rect -252 -736 -204 -708
rect -176 -736 -128 -708
rect -100 -736 -52 -708
rect -24 -736 24 -708
rect 52 -736 100 -708
rect 128 -736 176 -708
rect 204 -736 252 -708
rect 280 -736 328 -708
rect 356 -736 404 -708
rect 432 -736 480 -708
rect 508 -736 513 -708
rect -513 -784 513 -736
rect -513 -812 -508 -784
rect -480 -812 -432 -784
rect -404 -812 -356 -784
rect -328 -812 -280 -784
rect -252 -812 -204 -784
rect -176 -812 -128 -784
rect -100 -812 -52 -784
rect -24 -812 24 -784
rect 52 -812 100 -784
rect 128 -812 176 -784
rect 204 -812 252 -784
rect 280 -812 328 -784
rect 356 -812 404 -784
rect 432 -812 480 -784
rect 508 -812 513 -784
rect -513 -860 513 -812
rect -513 -888 -508 -860
rect -480 -888 -432 -860
rect -404 -888 -356 -860
rect -328 -888 -280 -860
rect -252 -888 -204 -860
rect -176 -888 -128 -860
rect -100 -888 -52 -860
rect -24 -888 24 -860
rect 52 -888 100 -860
rect 128 -888 176 -860
rect 204 -888 252 -860
rect 280 -888 328 -860
rect 356 -888 404 -860
rect 432 -888 480 -860
rect 508 -888 513 -860
rect -513 -936 513 -888
rect -513 -964 -508 -936
rect -480 -964 -432 -936
rect -404 -964 -356 -936
rect -328 -964 -280 -936
rect -252 -964 -204 -936
rect -176 -964 -128 -936
rect -100 -964 -52 -936
rect -24 -964 24 -936
rect 52 -964 100 -936
rect 128 -964 176 -936
rect 204 -964 252 -936
rect 280 -964 328 -936
rect 356 -964 404 -936
rect 432 -964 480 -936
rect 508 -964 513 -936
rect -513 -1012 513 -964
rect -513 -1040 -508 -1012
rect -480 -1040 -432 -1012
rect -404 -1040 -356 -1012
rect -328 -1040 -280 -1012
rect -252 -1040 -204 -1012
rect -176 -1040 -128 -1012
rect -100 -1040 -52 -1012
rect -24 -1040 24 -1012
rect 52 -1040 100 -1012
rect 128 -1040 176 -1012
rect 204 -1040 252 -1012
rect 280 -1040 328 -1012
rect 356 -1040 404 -1012
rect 432 -1040 480 -1012
rect 508 -1040 513 -1012
rect -513 -1088 513 -1040
rect -513 -1116 -508 -1088
rect -480 -1116 -432 -1088
rect -404 -1116 -356 -1088
rect -328 -1116 -280 -1088
rect -252 -1116 -204 -1088
rect -176 -1116 -128 -1088
rect -100 -1116 -52 -1088
rect -24 -1116 24 -1088
rect 52 -1116 100 -1088
rect 128 -1116 176 -1088
rect 204 -1116 252 -1088
rect 280 -1116 328 -1088
rect 356 -1116 404 -1088
rect 432 -1116 480 -1088
rect 508 -1116 513 -1088
rect -513 -1164 513 -1116
rect -513 -1192 -508 -1164
rect -480 -1192 -432 -1164
rect -404 -1192 -356 -1164
rect -328 -1192 -280 -1164
rect -252 -1192 -204 -1164
rect -176 -1192 -128 -1164
rect -100 -1192 -52 -1164
rect -24 -1192 24 -1164
rect 52 -1192 100 -1164
rect 128 -1192 176 -1164
rect 204 -1192 252 -1164
rect 280 -1192 328 -1164
rect 356 -1192 404 -1164
rect 432 -1192 480 -1164
rect 508 -1192 513 -1164
rect -513 -1240 513 -1192
rect -513 -1268 -508 -1240
rect -480 -1268 -432 -1240
rect -404 -1268 -356 -1240
rect -328 -1268 -280 -1240
rect -252 -1268 -204 -1240
rect -176 -1268 -128 -1240
rect -100 -1268 -52 -1240
rect -24 -1268 24 -1240
rect 52 -1268 100 -1240
rect 128 -1268 176 -1240
rect 204 -1268 252 -1240
rect 280 -1268 328 -1240
rect 356 -1268 404 -1240
rect 432 -1268 480 -1240
rect 508 -1268 513 -1240
rect -513 -1316 513 -1268
rect -513 -1344 -508 -1316
rect -480 -1344 -432 -1316
rect -404 -1344 -356 -1316
rect -328 -1344 -280 -1316
rect -252 -1344 -204 -1316
rect -176 -1344 -128 -1316
rect -100 -1344 -52 -1316
rect -24 -1344 24 -1316
rect 52 -1344 100 -1316
rect 128 -1344 176 -1316
rect 204 -1344 252 -1316
rect 280 -1344 328 -1316
rect 356 -1344 404 -1316
rect 432 -1344 480 -1316
rect 508 -1344 513 -1316
rect -513 -1392 513 -1344
rect -513 -1420 -508 -1392
rect -480 -1420 -432 -1392
rect -404 -1420 -356 -1392
rect -328 -1420 -280 -1392
rect -252 -1420 -204 -1392
rect -176 -1420 -128 -1392
rect -100 -1420 -52 -1392
rect -24 -1420 24 -1392
rect 52 -1420 100 -1392
rect 128 -1420 176 -1392
rect 204 -1420 252 -1392
rect 280 -1420 328 -1392
rect 356 -1420 404 -1392
rect 432 -1420 480 -1392
rect 508 -1420 513 -1392
rect -513 -1468 513 -1420
rect -513 -1496 -508 -1468
rect -480 -1496 -432 -1468
rect -404 -1496 -356 -1468
rect -328 -1496 -280 -1468
rect -252 -1496 -204 -1468
rect -176 -1496 -128 -1468
rect -100 -1496 -52 -1468
rect -24 -1496 24 -1468
rect 52 -1496 100 -1468
rect 128 -1496 176 -1468
rect 204 -1496 252 -1468
rect 280 -1496 328 -1468
rect 356 -1496 404 -1468
rect 432 -1496 480 -1468
rect 508 -1496 513 -1468
rect -513 -1544 513 -1496
rect -513 -1572 -508 -1544
rect -480 -1572 -432 -1544
rect -404 -1572 -356 -1544
rect -328 -1572 -280 -1544
rect -252 -1572 -204 -1544
rect -176 -1572 -128 -1544
rect -100 -1572 -52 -1544
rect -24 -1572 24 -1544
rect 52 -1572 100 -1544
rect 128 -1572 176 -1544
rect 204 -1572 252 -1544
rect 280 -1572 328 -1544
rect 356 -1572 404 -1544
rect 432 -1572 480 -1544
rect 508 -1572 513 -1544
rect -513 -1620 513 -1572
rect -513 -1648 -508 -1620
rect -480 -1648 -432 -1620
rect -404 -1648 -356 -1620
rect -328 -1648 -280 -1620
rect -252 -1648 -204 -1620
rect -176 -1648 -128 -1620
rect -100 -1648 -52 -1620
rect -24 -1648 24 -1620
rect 52 -1648 100 -1620
rect 128 -1648 176 -1620
rect 204 -1648 252 -1620
rect 280 -1648 328 -1620
rect 356 -1648 404 -1620
rect 432 -1648 480 -1620
rect 508 -1648 513 -1620
rect -513 -1696 513 -1648
rect -513 -1724 -508 -1696
rect -480 -1724 -432 -1696
rect -404 -1724 -356 -1696
rect -328 -1724 -280 -1696
rect -252 -1724 -204 -1696
rect -176 -1724 -128 -1696
rect -100 -1724 -52 -1696
rect -24 -1724 24 -1696
rect 52 -1724 100 -1696
rect 128 -1724 176 -1696
rect 204 -1724 252 -1696
rect 280 -1724 328 -1696
rect 356 -1724 404 -1696
rect 432 -1724 480 -1696
rect 508 -1724 513 -1696
rect -513 -1772 513 -1724
rect -513 -1800 -508 -1772
rect -480 -1800 -432 -1772
rect -404 -1800 -356 -1772
rect -328 -1800 -280 -1772
rect -252 -1800 -204 -1772
rect -176 -1800 -128 -1772
rect -100 -1800 -52 -1772
rect -24 -1800 24 -1772
rect 52 -1800 100 -1772
rect 128 -1800 176 -1772
rect 204 -1800 252 -1772
rect 280 -1800 328 -1772
rect 356 -1800 404 -1772
rect 432 -1800 480 -1772
rect 508 -1800 513 -1772
rect -513 -1848 513 -1800
rect -513 -1876 -508 -1848
rect -480 -1876 -432 -1848
rect -404 -1876 -356 -1848
rect -328 -1876 -280 -1848
rect -252 -1876 -204 -1848
rect -176 -1876 -128 -1848
rect -100 -1876 -52 -1848
rect -24 -1876 24 -1848
rect 52 -1876 100 -1848
rect 128 -1876 176 -1848
rect 204 -1876 252 -1848
rect 280 -1876 328 -1848
rect 356 -1876 404 -1848
rect 432 -1876 480 -1848
rect 508 -1876 513 -1848
rect -513 -1924 513 -1876
rect -513 -1952 -508 -1924
rect -480 -1952 -432 -1924
rect -404 -1952 -356 -1924
rect -328 -1952 -280 -1924
rect -252 -1952 -204 -1924
rect -176 -1952 -128 -1924
rect -100 -1952 -52 -1924
rect -24 -1952 24 -1924
rect 52 -1952 100 -1924
rect 128 -1952 176 -1924
rect 204 -1952 252 -1924
rect 280 -1952 328 -1924
rect 356 -1952 404 -1924
rect 432 -1952 480 -1924
rect 508 -1952 513 -1924
rect -513 -2000 513 -1952
rect -513 -2028 -508 -2000
rect -480 -2028 -432 -2000
rect -404 -2028 -356 -2000
rect -328 -2028 -280 -2000
rect -252 -2028 -204 -2000
rect -176 -2028 -128 -2000
rect -100 -2028 -52 -2000
rect -24 -2028 24 -2000
rect 52 -2028 100 -2000
rect 128 -2028 176 -2000
rect 204 -2028 252 -2000
rect 280 -2028 328 -2000
rect 356 -2028 404 -2000
rect 432 -2028 480 -2000
rect 508 -2028 513 -2000
rect -513 -2076 513 -2028
rect -513 -2104 -508 -2076
rect -480 -2104 -432 -2076
rect -404 -2104 -356 -2076
rect -328 -2104 -280 -2076
rect -252 -2104 -204 -2076
rect -176 -2104 -128 -2076
rect -100 -2104 -52 -2076
rect -24 -2104 24 -2076
rect 52 -2104 100 -2076
rect 128 -2104 176 -2076
rect 204 -2104 252 -2076
rect 280 -2104 328 -2076
rect 356 -2104 404 -2076
rect 432 -2104 480 -2076
rect 508 -2104 513 -2076
rect -513 -2152 513 -2104
rect -513 -2180 -508 -2152
rect -480 -2180 -432 -2152
rect -404 -2180 -356 -2152
rect -328 -2180 -280 -2152
rect -252 -2180 -204 -2152
rect -176 -2180 -128 -2152
rect -100 -2180 -52 -2152
rect -24 -2180 24 -2152
rect 52 -2180 100 -2152
rect 128 -2180 176 -2152
rect 204 -2180 252 -2152
rect 280 -2180 328 -2152
rect 356 -2180 404 -2152
rect 432 -2180 480 -2152
rect 508 -2180 513 -2152
rect -513 -2228 513 -2180
rect -513 -2256 -508 -2228
rect -480 -2256 -432 -2228
rect -404 -2256 -356 -2228
rect -328 -2256 -280 -2228
rect -252 -2256 -204 -2228
rect -176 -2256 -128 -2228
rect -100 -2256 -52 -2228
rect -24 -2256 24 -2228
rect 52 -2256 100 -2228
rect 128 -2256 176 -2228
rect 204 -2256 252 -2228
rect 280 -2256 328 -2228
rect 356 -2256 404 -2228
rect 432 -2256 480 -2228
rect 508 -2256 513 -2228
rect -513 -2304 513 -2256
rect -513 -2332 -508 -2304
rect -480 -2332 -432 -2304
rect -404 -2332 -356 -2304
rect -328 -2332 -280 -2304
rect -252 -2332 -204 -2304
rect -176 -2332 -128 -2304
rect -100 -2332 -52 -2304
rect -24 -2332 24 -2304
rect 52 -2332 100 -2304
rect 128 -2332 176 -2304
rect 204 -2332 252 -2304
rect 280 -2332 328 -2304
rect 356 -2332 404 -2304
rect 432 -2332 480 -2304
rect 508 -2332 513 -2304
rect -513 -2380 513 -2332
rect -513 -2408 -508 -2380
rect -480 -2408 -432 -2380
rect -404 -2408 -356 -2380
rect -328 -2408 -280 -2380
rect -252 -2408 -204 -2380
rect -176 -2408 -128 -2380
rect -100 -2408 -52 -2380
rect -24 -2408 24 -2380
rect 52 -2408 100 -2380
rect 128 -2408 176 -2380
rect 204 -2408 252 -2380
rect 280 -2408 328 -2380
rect 356 -2408 404 -2380
rect 432 -2408 480 -2380
rect 508 -2408 513 -2380
rect -513 -2456 513 -2408
rect -513 -2484 -508 -2456
rect -480 -2484 -432 -2456
rect -404 -2484 -356 -2456
rect -328 -2484 -280 -2456
rect -252 -2484 -204 -2456
rect -176 -2484 -128 -2456
rect -100 -2484 -52 -2456
rect -24 -2484 24 -2456
rect 52 -2484 100 -2456
rect 128 -2484 176 -2456
rect 204 -2484 252 -2456
rect 280 -2484 328 -2456
rect 356 -2484 404 -2456
rect 432 -2484 480 -2456
rect 508 -2484 513 -2456
rect -513 -2532 513 -2484
rect -513 -2560 -508 -2532
rect -480 -2560 -432 -2532
rect -404 -2560 -356 -2532
rect -328 -2560 -280 -2532
rect -252 -2560 -204 -2532
rect -176 -2560 -128 -2532
rect -100 -2560 -52 -2532
rect -24 -2560 24 -2532
rect 52 -2560 100 -2532
rect 128 -2560 176 -2532
rect 204 -2560 252 -2532
rect 280 -2560 328 -2532
rect 356 -2560 404 -2532
rect 432 -2560 480 -2532
rect 508 -2560 513 -2532
rect -513 -2608 513 -2560
rect -513 -2636 -508 -2608
rect -480 -2636 -432 -2608
rect -404 -2636 -356 -2608
rect -328 -2636 -280 -2608
rect -252 -2636 -204 -2608
rect -176 -2636 -128 -2608
rect -100 -2636 -52 -2608
rect -24 -2636 24 -2608
rect 52 -2636 100 -2608
rect 128 -2636 176 -2608
rect 204 -2636 252 -2608
rect 280 -2636 328 -2608
rect 356 -2636 404 -2608
rect 432 -2636 480 -2608
rect 508 -2636 513 -2608
rect -513 -2641 513 -2636
<< end >>
