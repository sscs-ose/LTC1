* NGSPICE file created from buffer_loading_mag_flat.ext - technology: gf180mcuC

.subckt buffer_loading_mag_flat VDD VSS OUT IN
X0 OUT a_168_68# VDD.t14 VDD.t13 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 VSS IN.t0 a_168_68# VSS.t7 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X2 OUT a_168_68# VSS.t19 VSS.t18 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X3 a_168_68# IN.t1 VDD.t1 VDD.t0 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X4 a_168_68# IN.t2 VSS.t6 VSS.t5 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X5 VDD IN.t3 a_168_68# VDD.t15 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X6 VSS a_168_68# OUT.t1 VSS.t15 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X7 OUT a_168_68# VDD.t12 VDD.t11 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X8 VDD a_168_68# OUT.t4 VDD.t8 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X9 a_168_68# IN.t4 VDD.t19 VDD.t18 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X10 OUT a_168_68# VSS.t14 VSS.t13 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X11 VSS IN.t5 a_168_68# VSS.t2 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X12 VDD IN.t6 a_168_68# VDD.t2 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X13 VSS a_168_68# OUT.t0 VSS.t10 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X14 a_168_68# IN.t7 VSS.t1 VSS.t0 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X15 VDD a_168_68# OUT.t3 VDD.t5 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
R0 VDD.n11 VDD.t11 289.017
R1 VDD.n11 VDD.t15 265.897
R2 VDD.t13 VDD.t8 231.214
R3 VDD.t5 VDD.t13 231.214
R4 VDD.t11 VDD.t5 231.214
R5 VDD.t15 VDD.t0 231.214
R6 VDD.t0 VDD.t2 231.214
R7 VDD.t2 VDD.t18 231.214
R8 VDD.n8 VDD.t19 4.87751
R9 VDD.n3 VDD.n2 4.87713
R10 VDD.n9 VDD.n5 4.7565
R11 VDD.n4 VDD.t12 4.7565
R12 VDD.n13 VDD.n12 3.1505
R13 VDD.n12 VDD.n11 3.1505
R14 VDD.n8 VDD.n7 2.9365
R15 VDD.n3 VDD.n1 2.9365
R16 VDD.n7 VDD.t1 1.8205
R17 VDD.n7 VDD.n6 1.8205
R18 VDD.n1 VDD.t14 1.8205
R19 VDD.n1 VDD.n0 1.8205
R20 VDD.n12 VDD.n10 0.152307
R21 VDD.n4 VDD.n3 0.121508
R22 VDD.n9 VDD.n8 0.12113
R23 VDD VDD.n4 0.0436092
R24 VDD.n13 VDD.n9 0.0409622
R25 VDD VDD.n13 0.00201261
R26 OUT.n4 OUT.n3 3.416
R27 OUT.n9 OUT.n8 3.416
R28 OUT.n3 OUT.t0 3.2765
R29 OUT.n3 OUT.n2 3.2765
R30 OUT.n8 OUT.t1 3.2765
R31 OUT.n8 OUT.n7 3.2765
R32 OUT.n4 OUT.n1 3.013
R33 OUT.n9 OUT.n6 3.013
R34 OUT.n1 OUT.t3 1.8205
R35 OUT.n1 OUT.n0 1.8205
R36 OUT.n6 OUT.t4 1.8205
R37 OUT.n6 OUT.n5 1.8205
R38 OUT.n9 OUT.n4 0.445308
R39 OUT OUT.n9 0.310308
R40 IN.n1 IN.t1 34.8567
R41 IN.n2 IN.t6 34.85
R42 IN.n0 IN.t3 34.8414
R43 IN.n3 IN.t4 31.3659
R44 IN.n0 IN.t5 22.634
R45 IN.n2 IN.t0 22.6274
R46 IN.n1 IN.t7 22.6208
R47 IN.n4 IN.t2 16.7006
R48 IN.n2 IN.n1 14.3197
R49 IN.n3 IN.n2 14.3197
R50 IN.n1 IN.n0 13.8986
R51 IN IN.n4 4.12947
R52 IN.n4 IN.n3 0.604959
R53 VSS.n5 VSS.t18 1543.12
R54 VSS.t13 VSS.t15 1007.75
R55 VSS.t10 VSS.t13 1007.75
R56 VSS.t18 VSS.t10 1007.75
R57 VSS.t2 VSS.t0 1007.75
R58 VSS.t0 VSS.t7 1007.75
R59 VSS.t7 VSS.t5 1007.75
R60 VSS.n5 VSS.t2 875.485
R61 VSS.n12 VSS.t6 6.77222
R62 VSS.n3 VSS.n2 6.77171
R63 VSS.n4 VSS.t19 6.61132
R64 VSS.n13 VSS.n9 6.61132
R65 VSS.n3 VSS.n1 3.33532
R66 VSS.n12 VSS.n11 3.33532
R67 VSS.n1 VSS.t14 3.2765
R68 VSS.n1 VSS.n0 3.2765
R69 VSS.n11 VSS.t1 3.2765
R70 VSS.n11 VSS.n10 3.2765
R71 VSS.n8 VSS.n7 2.6005
R72 VSS.n7 VSS.n5 2.6005
R73 VSS.n7 VSS.n6 0.477773
R74 VSS.n4 VSS.n3 0.161394
R75 VSS.n13 VSS.n12 0.160891
R76 VSS.n8 VSS.n4 0.0824553
R77 VSS VSS.n13 0.027148
R78 VSS VSS.n8 0.00502514
C0 VDD OUT 0.579f
C1 IN OUT 0.00154f
C2 VDD a_168_68# 1.17f
C3 IN a_168_68# 0.329f
C4 IN VDD 0.59f
C5 OUT a_168_68# 0.33f
.ends

