magic
tech gf180mcuC
magscale 1 10
timestamp 1693394299
<< error_p >>
rect -3287 -58 -3241 58
rect -3083 -58 -3037 58
rect -2879 -58 -2833 58
rect -2675 -58 -2629 58
rect -2471 -58 -2425 58
rect -2267 -58 -2221 58
rect -2063 -58 -2017 58
rect -1859 -58 -1813 58
rect -1655 -58 -1609 58
rect -1451 -58 -1405 58
rect -1247 -58 -1201 58
rect -1043 -58 -997 58
rect -839 -58 -793 58
rect -635 -58 -589 58
rect -431 -58 -385 58
rect -227 -58 -181 58
rect -23 -58 23 58
rect 181 -58 227 58
rect 385 -58 431 58
rect 589 -58 635 58
rect 793 -58 839 58
rect 997 -58 1043 58
rect 1201 -58 1247 58
rect 1405 -58 1451 58
rect 1609 -58 1655 58
rect 1813 -58 1859 58
rect 2017 -58 2063 58
rect 2221 -58 2267 58
rect 2425 -58 2471 58
rect 2629 -58 2675 58
rect 2833 -58 2879 58
rect 3037 -58 3083 58
rect 3241 -58 3287 58
<< nwell >>
rect -3386 -190 3386 190
<< pmos >>
rect -3212 -60 -3112 60
rect -3008 -60 -2908 60
rect -2804 -60 -2704 60
rect -2600 -60 -2500 60
rect -2396 -60 -2296 60
rect -2192 -60 -2092 60
rect -1988 -60 -1888 60
rect -1784 -60 -1684 60
rect -1580 -60 -1480 60
rect -1376 -60 -1276 60
rect -1172 -60 -1072 60
rect -968 -60 -868 60
rect -764 -60 -664 60
rect -560 -60 -460 60
rect -356 -60 -256 60
rect -152 -60 -52 60
rect 52 -60 152 60
rect 256 -60 356 60
rect 460 -60 560 60
rect 664 -60 764 60
rect 868 -60 968 60
rect 1072 -60 1172 60
rect 1276 -60 1376 60
rect 1480 -60 1580 60
rect 1684 -60 1784 60
rect 1888 -60 1988 60
rect 2092 -60 2192 60
rect 2296 -60 2396 60
rect 2500 -60 2600 60
rect 2704 -60 2804 60
rect 2908 -60 3008 60
rect 3112 -60 3212 60
<< pdiff >>
rect -3300 47 -3212 60
rect -3300 -47 -3287 47
rect -3241 -47 -3212 47
rect -3300 -60 -3212 -47
rect -3112 47 -3008 60
rect -3112 -47 -3083 47
rect -3037 -47 -3008 47
rect -3112 -60 -3008 -47
rect -2908 47 -2804 60
rect -2908 -47 -2879 47
rect -2833 -47 -2804 47
rect -2908 -60 -2804 -47
rect -2704 47 -2600 60
rect -2704 -47 -2675 47
rect -2629 -47 -2600 47
rect -2704 -60 -2600 -47
rect -2500 47 -2396 60
rect -2500 -47 -2471 47
rect -2425 -47 -2396 47
rect -2500 -60 -2396 -47
rect -2296 47 -2192 60
rect -2296 -47 -2267 47
rect -2221 -47 -2192 47
rect -2296 -60 -2192 -47
rect -2092 47 -1988 60
rect -2092 -47 -2063 47
rect -2017 -47 -1988 47
rect -2092 -60 -1988 -47
rect -1888 47 -1784 60
rect -1888 -47 -1859 47
rect -1813 -47 -1784 47
rect -1888 -60 -1784 -47
rect -1684 47 -1580 60
rect -1684 -47 -1655 47
rect -1609 -47 -1580 47
rect -1684 -60 -1580 -47
rect -1480 47 -1376 60
rect -1480 -47 -1451 47
rect -1405 -47 -1376 47
rect -1480 -60 -1376 -47
rect -1276 47 -1172 60
rect -1276 -47 -1247 47
rect -1201 -47 -1172 47
rect -1276 -60 -1172 -47
rect -1072 47 -968 60
rect -1072 -47 -1043 47
rect -997 -47 -968 47
rect -1072 -60 -968 -47
rect -868 47 -764 60
rect -868 -47 -839 47
rect -793 -47 -764 47
rect -868 -60 -764 -47
rect -664 47 -560 60
rect -664 -47 -635 47
rect -589 -47 -560 47
rect -664 -60 -560 -47
rect -460 47 -356 60
rect -460 -47 -431 47
rect -385 -47 -356 47
rect -460 -60 -356 -47
rect -256 47 -152 60
rect -256 -47 -227 47
rect -181 -47 -152 47
rect -256 -60 -152 -47
rect -52 47 52 60
rect -52 -47 -23 47
rect 23 -47 52 47
rect -52 -60 52 -47
rect 152 47 256 60
rect 152 -47 181 47
rect 227 -47 256 47
rect 152 -60 256 -47
rect 356 47 460 60
rect 356 -47 385 47
rect 431 -47 460 47
rect 356 -60 460 -47
rect 560 47 664 60
rect 560 -47 589 47
rect 635 -47 664 47
rect 560 -60 664 -47
rect 764 47 868 60
rect 764 -47 793 47
rect 839 -47 868 47
rect 764 -60 868 -47
rect 968 47 1072 60
rect 968 -47 997 47
rect 1043 -47 1072 47
rect 968 -60 1072 -47
rect 1172 47 1276 60
rect 1172 -47 1201 47
rect 1247 -47 1276 47
rect 1172 -60 1276 -47
rect 1376 47 1480 60
rect 1376 -47 1405 47
rect 1451 -47 1480 47
rect 1376 -60 1480 -47
rect 1580 47 1684 60
rect 1580 -47 1609 47
rect 1655 -47 1684 47
rect 1580 -60 1684 -47
rect 1784 47 1888 60
rect 1784 -47 1813 47
rect 1859 -47 1888 47
rect 1784 -60 1888 -47
rect 1988 47 2092 60
rect 1988 -47 2017 47
rect 2063 -47 2092 47
rect 1988 -60 2092 -47
rect 2192 47 2296 60
rect 2192 -47 2221 47
rect 2267 -47 2296 47
rect 2192 -60 2296 -47
rect 2396 47 2500 60
rect 2396 -47 2425 47
rect 2471 -47 2500 47
rect 2396 -60 2500 -47
rect 2600 47 2704 60
rect 2600 -47 2629 47
rect 2675 -47 2704 47
rect 2600 -60 2704 -47
rect 2804 47 2908 60
rect 2804 -47 2833 47
rect 2879 -47 2908 47
rect 2804 -60 2908 -47
rect 3008 47 3112 60
rect 3008 -47 3037 47
rect 3083 -47 3112 47
rect 3008 -60 3112 -47
rect 3212 47 3300 60
rect 3212 -47 3241 47
rect 3287 -47 3300 47
rect 3212 -60 3300 -47
<< pdiffc >>
rect -3287 -47 -3241 47
rect -3083 -47 -3037 47
rect -2879 -47 -2833 47
rect -2675 -47 -2629 47
rect -2471 -47 -2425 47
rect -2267 -47 -2221 47
rect -2063 -47 -2017 47
rect -1859 -47 -1813 47
rect -1655 -47 -1609 47
rect -1451 -47 -1405 47
rect -1247 -47 -1201 47
rect -1043 -47 -997 47
rect -839 -47 -793 47
rect -635 -47 -589 47
rect -431 -47 -385 47
rect -227 -47 -181 47
rect -23 -47 23 47
rect 181 -47 227 47
rect 385 -47 431 47
rect 589 -47 635 47
rect 793 -47 839 47
rect 997 -47 1043 47
rect 1201 -47 1247 47
rect 1405 -47 1451 47
rect 1609 -47 1655 47
rect 1813 -47 1859 47
rect 2017 -47 2063 47
rect 2221 -47 2267 47
rect 2425 -47 2471 47
rect 2629 -47 2675 47
rect 2833 -47 2879 47
rect 3037 -47 3083 47
rect 3241 -47 3287 47
<< polysilicon >>
rect -3212 60 -3112 104
rect -3008 60 -2908 104
rect -2804 60 -2704 104
rect -2600 60 -2500 104
rect -2396 60 -2296 104
rect -2192 60 -2092 104
rect -1988 60 -1888 104
rect -1784 60 -1684 104
rect -1580 60 -1480 104
rect -1376 60 -1276 104
rect -1172 60 -1072 104
rect -968 60 -868 104
rect -764 60 -664 104
rect -560 60 -460 104
rect -356 60 -256 104
rect -152 60 -52 104
rect 52 60 152 104
rect 256 60 356 104
rect 460 60 560 104
rect 664 60 764 104
rect 868 60 968 104
rect 1072 60 1172 104
rect 1276 60 1376 104
rect 1480 60 1580 104
rect 1684 60 1784 104
rect 1888 60 1988 104
rect 2092 60 2192 104
rect 2296 60 2396 104
rect 2500 60 2600 104
rect 2704 60 2804 104
rect 2908 60 3008 104
rect 3112 60 3212 104
rect -3212 -104 -3112 -60
rect -3008 -104 -2908 -60
rect -2804 -104 -2704 -60
rect -2600 -104 -2500 -60
rect -2396 -104 -2296 -60
rect -2192 -104 -2092 -60
rect -1988 -104 -1888 -60
rect -1784 -104 -1684 -60
rect -1580 -104 -1480 -60
rect -1376 -104 -1276 -60
rect -1172 -104 -1072 -60
rect -968 -104 -868 -60
rect -764 -104 -664 -60
rect -560 -104 -460 -60
rect -356 -104 -256 -60
rect -152 -104 -52 -60
rect 52 -104 152 -60
rect 256 -104 356 -60
rect 460 -104 560 -60
rect 664 -104 764 -60
rect 868 -104 968 -60
rect 1072 -104 1172 -60
rect 1276 -104 1376 -60
rect 1480 -104 1580 -60
rect 1684 -104 1784 -60
rect 1888 -104 1988 -60
rect 2092 -104 2192 -60
rect 2296 -104 2396 -60
rect 2500 -104 2600 -60
rect 2704 -104 2804 -60
rect 2908 -104 3008 -60
rect 3112 -104 3212 -60
<< metal1 >>
rect -3287 47 -3241 58
rect -3287 -58 -3241 -47
rect -3083 47 -3037 58
rect -3083 -58 -3037 -47
rect -2879 47 -2833 58
rect -2879 -58 -2833 -47
rect -2675 47 -2629 58
rect -2675 -58 -2629 -47
rect -2471 47 -2425 58
rect -2471 -58 -2425 -47
rect -2267 47 -2221 58
rect -2267 -58 -2221 -47
rect -2063 47 -2017 58
rect -2063 -58 -2017 -47
rect -1859 47 -1813 58
rect -1859 -58 -1813 -47
rect -1655 47 -1609 58
rect -1655 -58 -1609 -47
rect -1451 47 -1405 58
rect -1451 -58 -1405 -47
rect -1247 47 -1201 58
rect -1247 -58 -1201 -47
rect -1043 47 -997 58
rect -1043 -58 -997 -47
rect -839 47 -793 58
rect -839 -58 -793 -47
rect -635 47 -589 58
rect -635 -58 -589 -47
rect -431 47 -385 58
rect -431 -58 -385 -47
rect -227 47 -181 58
rect -227 -58 -181 -47
rect -23 47 23 58
rect -23 -58 23 -47
rect 181 47 227 58
rect 181 -58 227 -47
rect 385 47 431 58
rect 385 -58 431 -47
rect 589 47 635 58
rect 589 -58 635 -47
rect 793 47 839 58
rect 793 -58 839 -47
rect 997 47 1043 58
rect 997 -58 1043 -47
rect 1201 47 1247 58
rect 1201 -58 1247 -47
rect 1405 47 1451 58
rect 1405 -58 1451 -47
rect 1609 47 1655 58
rect 1609 -58 1655 -47
rect 1813 47 1859 58
rect 1813 -58 1859 -47
rect 2017 47 2063 58
rect 2017 -58 2063 -47
rect 2221 47 2267 58
rect 2221 -58 2267 -47
rect 2425 47 2471 58
rect 2425 -58 2471 -47
rect 2629 47 2675 58
rect 2629 -58 2675 -47
rect 2833 47 2879 58
rect 2833 -58 2879 -47
rect 3037 47 3083 58
rect 3037 -58 3083 -47
rect 3241 47 3287 58
rect 3241 -58 3287 -47
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 0.6 l 0.5 m 1 nf 32 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
