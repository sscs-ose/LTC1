magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1112 -1143 1112 1143
<< metal1 >>
rect -112 137 112 143
rect -112 111 -106 137
rect -80 111 -44 137
rect -18 111 18 137
rect 44 111 80 137
rect 106 111 112 137
rect -112 75 112 111
rect -112 49 -106 75
rect -80 49 -44 75
rect -18 49 18 75
rect 44 49 80 75
rect 106 49 112 75
rect -112 13 112 49
rect -112 -13 -106 13
rect -80 -13 -44 13
rect -18 -13 18 13
rect 44 -13 80 13
rect 106 -13 112 13
rect -112 -49 112 -13
rect -112 -75 -106 -49
rect -80 -75 -44 -49
rect -18 -75 18 -49
rect 44 -75 80 -49
rect 106 -75 112 -49
rect -112 -111 112 -75
rect -112 -137 -106 -111
rect -80 -137 -44 -111
rect -18 -137 18 -111
rect 44 -137 80 -111
rect 106 -137 112 -111
rect -112 -143 112 -137
<< via1 >>
rect -106 111 -80 137
rect -44 111 -18 137
rect 18 111 44 137
rect 80 111 106 137
rect -106 49 -80 75
rect -44 49 -18 75
rect 18 49 44 75
rect 80 49 106 75
rect -106 -13 -80 13
rect -44 -13 -18 13
rect 18 -13 44 13
rect 80 -13 106 13
rect -106 -75 -80 -49
rect -44 -75 -18 -49
rect 18 -75 44 -49
rect 80 -75 106 -49
rect -106 -137 -80 -111
rect -44 -137 -18 -111
rect 18 -137 44 -111
rect 80 -137 106 -111
<< metal2 >>
rect -112 137 112 143
rect -112 111 -106 137
rect -80 111 -44 137
rect -18 111 18 137
rect 44 111 80 137
rect 106 111 112 137
rect -112 75 112 111
rect -112 49 -106 75
rect -80 49 -44 75
rect -18 49 18 75
rect 44 49 80 75
rect 106 49 112 75
rect -112 13 112 49
rect -112 -13 -106 13
rect -80 -13 -44 13
rect -18 -13 18 13
rect 44 -13 80 13
rect 106 -13 112 13
rect -112 -49 112 -13
rect -112 -75 -106 -49
rect -80 -75 -44 -49
rect -18 -75 18 -49
rect 44 -75 80 -49
rect 106 -75 112 -49
rect -112 -111 112 -75
rect -112 -137 -106 -111
rect -80 -137 -44 -111
rect -18 -137 18 -111
rect 44 -137 80 -111
rect 106 -137 112 -111
rect -112 -143 112 -137
<< end >>
