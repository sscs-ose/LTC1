* NGSPICE file created from MSB_Unit_Cell.ext - technology: gf180mcuC

.subckt nmos_3p3_AGPLV7 a_n138_n60# a_50_n60# a_n50_n104# VSUBS
X0 a_50_n60# a_n50_n104# a_n138_n60# VSUBS nfet_03v3 ad=0.264p pd=2.08u as=0.264p ps=2.08u w=0.6u l=0.5u
.ends

.subckt nmos_3p3_AQEADK a_n138_n60# a_50_n60# a_n50_n104# VSUBS
X0 a_50_n60# a_n50_n104# a_n138_n60# VSUBS nfet_03v3 ad=0.264p pd=2.08u as=0.264p ps=2.08u w=0.6u l=0.5u
.ends

.subckt MSB_Unit_Cell_p2 m1_34_n336# a_316_n480# a_51_258# a_316_26# m1_23_6# a_3095_69#
+ VSUBS
Xnmos_3p3_AGPLV7_5 m1_34_n336# a_3095_69# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_6 a_3095_69# m1_23_6# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_7 m1_23_6# a_3095_69# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_8 a_3095_69# m1_34_n336# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_9 m1_34_n336# a_3095_69# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AQEADK_0 a_3095_69# m1_34_n336# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_1 m1_23_6# a_3095_69# a_51_258# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_2 a_3095_69# m1_34_n336# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_4 a_3095_69# m1_23_6# a_51_258# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_3 m1_34_n336# a_3095_69# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_5 m1_23_6# a_3095_69# a_51_258# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_10 a_3095_69# m1_23_6# a_51_258# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_6 a_3095_69# m1_34_n336# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_11 m1_34_n336# a_3095_69# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_7 m1_34_n336# a_3095_69# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_12 a_3095_69# m1_23_6# a_51_258# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_8 a_3095_69# m1_23_6# a_51_258# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_13 m1_23_6# a_3095_69# a_51_258# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_9 m1_23_6# a_3095_69# a_51_258# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_15 m1_34_n336# a_3095_69# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_14 a_3095_69# m1_34_n336# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AGPLV7_10 a_3095_69# m1_23_6# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_12 a_3095_69# m1_23_6# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_11 m1_23_6# a_3095_69# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_13 m1_34_n336# a_3095_69# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_14 m1_23_6# a_3095_69# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_15 a_3095_69# m1_34_n336# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_0 a_3095_69# m1_34_n336# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_1 m1_34_n336# a_3095_69# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_2 a_3095_69# m1_23_6# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_3 m1_23_6# a_3095_69# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_4 a_3095_69# m1_34_n336# a_316_26# VSUBS nmos_3p3_AGPLV7
.ends

.subckt pmos_3p3_M8RWPS a_n28_n94# w_n202_n180# a_n116_n50# a_28_n50#
X0 a_28_n50# a_n28_n94# a_n116_n50# w_n202_n180# pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
.ends

.subckt nmos_3p3_HZS5UA a_n28_n94# a_n116_n50# a_28_n50# VSUBS
X0 a_28_n50# a_n28_n94# a_n116_n50# VSUBS nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
.ends

.subckt NAND VDD VSS B A OUT
Xpmos_3p3_M8RWPS_0 A VDD VDD OUT pmos_3p3_M8RWPS
Xpmos_3p3_M8RWPS_1 B VDD VDD OUT pmos_3p3_M8RWPS
Xnmos_3p3_HZS5UA_0 A m1_184_67# OUT VSS nmos_3p3_HZS5UA
Xnmos_3p3_HZS5UA_1 B VSS m1_184_67# VSS nmos_3p3_HZS5UA
.ends

.subckt Local_Enc Ri-1 VDD Q QB Ci Ri VSS
XNAND_0 VDD VSS Ri-1 Ri-1 NAND_1/B NAND
XNAND_1 VDD VSS NAND_1/B NAND_1/B NAND_5/B NAND
XNAND_2 VDD VSS Ci Ci NAND_6/B NAND
XNAND_3 VDD VSS Ri Ri NAND_6/A NAND
XNAND_4 VDD VSS NAND_4/B Q QB NAND
XNAND_5 VDD VSS NAND_5/B NAND_5/A NAND_8/A NAND
XNAND_6 VDD VSS NAND_6/B NAND_6/A NAND_5/A NAND
XNAND_7 VDD VSS NAND_8/A NAND_8/A NAND_4/B NAND
XNAND_8 VDD VSS QB NAND_8/A Q NAND
.ends

.subckt MSB_Unit_Cell_p1 a_3095_69# a_86_241# m1_37_n24# a_316_n480# m1_0_379# m1_0_n631#
+ a_316_26# VSUBS
Xnmos_3p3_AGPLV7_5 m1_0_n631# a_3095_69# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_6 a_3095_69# m1_37_n24# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_7 m1_37_n24# a_3095_69# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_8 a_3095_69# m1_0_n631# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_9 m1_0_n631# a_3095_69# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AQEADK_0 a_3095_69# m1_0_379# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_1 m1_37_n24# a_3095_69# a_86_241# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_2 a_3095_69# m1_0_379# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_30 a_3095_69# m1_37_n24# a_86_241# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_4 a_3095_69# m1_37_n24# a_86_241# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_3 m1_0_379# a_3095_69# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_31 m1_0_379# a_3095_69# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_20 a_3095_69# m1_37_n24# a_86_241# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_5 m1_37_n24# a_3095_69# a_86_241# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_21 m1_37_n24# a_3095_69# a_86_241# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_10 a_3095_69# m1_37_n24# a_86_241# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_6 a_3095_69# m1_0_379# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_22 a_3095_69# m1_0_379# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_11 m1_0_379# a_3095_69# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_7 m1_0_379# a_3095_69# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_23 m1_0_379# a_3095_69# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_12 a_3095_69# m1_37_n24# a_86_241# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_8 a_3095_69# m1_37_n24# a_86_241# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AGPLV7_30 a_3095_69# m1_0_n631# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AQEADK_24 a_3095_69# m1_37_n24# a_86_241# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_13 m1_37_n24# a_3095_69# a_86_241# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_9 m1_37_n24# a_3095_69# a_86_241# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AGPLV7_31 m1_37_n24# a_3095_69# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_20 a_3095_69# m1_0_n631# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AQEADK_26 a_3095_69# m1_0_379# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_25 m1_37_n24# a_3095_69# a_86_241# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_15 m1_0_379# a_3095_69# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_14 a_3095_69# m1_0_379# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AGPLV7_21 a_3095_69# m1_37_n24# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_10 a_3095_69# m1_37_n24# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AQEADK_27 a_3095_69# m1_0_379# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_16 m1_0_379# a_3095_69# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AGPLV7_23 m1_37_n24# a_3095_69# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_22 a_3095_69# m1_0_n631# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_12 a_3095_69# m1_37_n24# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_11 m1_37_n24# a_3095_69# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AQEADK_28 a_3095_69# m1_37_n24# a_86_241# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_17 m1_37_n24# a_3095_69# a_86_241# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AGPLV7_24 m1_0_n631# a_3095_69# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_13 m1_0_n631# a_3095_69# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AQEADK_29 m1_37_n24# a_3095_69# a_86_241# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_18 a_3095_69# m1_0_379# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AGPLV7_25 m1_37_n24# a_3095_69# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_14 m1_37_n24# a_3095_69# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AQEADK_19 m1_0_379# a_3095_69# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AGPLV7_26 a_3095_69# m1_37_n24# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_15 a_3095_69# m1_0_n631# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_27 a_3095_69# m1_37_n24# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_16 a_3095_69# m1_37_n24# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_28 a_3095_69# m1_0_n631# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_17 m1_0_n631# a_3095_69# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_29 m1_0_n631# a_3095_69# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_18 m1_37_n24# a_3095_69# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_19 m1_0_n631# a_3095_69# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_0 a_3095_69# m1_0_n631# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_1 m1_0_n631# a_3095_69# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_2 a_3095_69# m1_37_n24# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_3 m1_37_n24# a_3095_69# a_316_n480# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_4 a_3095_69# m1_0_n631# a_316_26# VSUBS nmos_3p3_AGPLV7
.ends

.subckt MSB_Unit_Cell Ri-1 Ci Ri VSS VDD IM_T IM IOUT+
XMSB_Unit_Cell_p2_3 m2_3332_6234# Local_Enc_0/Q Local_Enc_0/Q Local_Enc_0/QB IOUT+
+ m1_3106_3593# VSS MSB_Unit_Cell_p2
XLocal_Enc_0 Ri-1 VDD Local_Enc_0/Q Local_Enc_0/QB Ci Ri VSS Local_Enc
XMSB_Unit_Cell_p1_1 m2_643_2191# IM_T m1_3106_3593# IM_T VSS VSS IM VSS MSB_Unit_Cell_p1
XMSB_Unit_Cell_p1_0 m2_643_2191# IM_T m1_3106_3593# IM_T VSS VSS IM VSS MSB_Unit_Cell_p1
XMSB_Unit_Cell_p2_0 m2_3332_6234# Local_Enc_0/Q Local_Enc_0/Q Local_Enc_0/QB IOUT+
+ m1_3106_3593# VSS MSB_Unit_Cell_p2
XMSB_Unit_Cell_p2_1 m2_3332_6234# Local_Enc_0/Q Local_Enc_0/Q Local_Enc_0/QB IOUT+
+ m1_3106_3593# VSS MSB_Unit_Cell_p2
XMSB_Unit_Cell_p2_2 m2_3332_6234# Local_Enc_0/Q Local_Enc_0/Q Local_Enc_0/QB IOUT+
+ m1_3106_3593# VSS MSB_Unit_Cell_p2
.ends

