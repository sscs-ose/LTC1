magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1236 -1763 1236 1763
<< metal1 >>
rect -236 757 236 763
rect -236 731 -230 757
rect -204 731 -168 757
rect -142 731 -106 757
rect -80 731 -44 757
rect -18 731 18 757
rect 44 731 80 757
rect 106 731 142 757
rect 168 731 204 757
rect 230 731 236 757
rect -236 695 236 731
rect -236 669 -230 695
rect -204 669 -168 695
rect -142 669 -106 695
rect -80 669 -44 695
rect -18 669 18 695
rect 44 669 80 695
rect 106 669 142 695
rect 168 669 204 695
rect 230 669 236 695
rect -236 633 236 669
rect -236 607 -230 633
rect -204 607 -168 633
rect -142 607 -106 633
rect -80 607 -44 633
rect -18 607 18 633
rect 44 607 80 633
rect 106 607 142 633
rect 168 607 204 633
rect 230 607 236 633
rect -236 571 236 607
rect -236 545 -230 571
rect -204 545 -168 571
rect -142 545 -106 571
rect -80 545 -44 571
rect -18 545 18 571
rect 44 545 80 571
rect 106 545 142 571
rect 168 545 204 571
rect 230 545 236 571
rect -236 509 236 545
rect -236 483 -230 509
rect -204 483 -168 509
rect -142 483 -106 509
rect -80 483 -44 509
rect -18 483 18 509
rect 44 483 80 509
rect 106 483 142 509
rect 168 483 204 509
rect 230 483 236 509
rect -236 447 236 483
rect -236 421 -230 447
rect -204 421 -168 447
rect -142 421 -106 447
rect -80 421 -44 447
rect -18 421 18 447
rect 44 421 80 447
rect 106 421 142 447
rect 168 421 204 447
rect 230 421 236 447
rect -236 385 236 421
rect -236 359 -230 385
rect -204 359 -168 385
rect -142 359 -106 385
rect -80 359 -44 385
rect -18 359 18 385
rect 44 359 80 385
rect 106 359 142 385
rect 168 359 204 385
rect 230 359 236 385
rect -236 323 236 359
rect -236 297 -230 323
rect -204 297 -168 323
rect -142 297 -106 323
rect -80 297 -44 323
rect -18 297 18 323
rect 44 297 80 323
rect 106 297 142 323
rect 168 297 204 323
rect 230 297 236 323
rect -236 261 236 297
rect -236 235 -230 261
rect -204 235 -168 261
rect -142 235 -106 261
rect -80 235 -44 261
rect -18 235 18 261
rect 44 235 80 261
rect 106 235 142 261
rect 168 235 204 261
rect 230 235 236 261
rect -236 199 236 235
rect -236 173 -230 199
rect -204 173 -168 199
rect -142 173 -106 199
rect -80 173 -44 199
rect -18 173 18 199
rect 44 173 80 199
rect 106 173 142 199
rect 168 173 204 199
rect 230 173 236 199
rect -236 137 236 173
rect -236 111 -230 137
rect -204 111 -168 137
rect -142 111 -106 137
rect -80 111 -44 137
rect -18 111 18 137
rect 44 111 80 137
rect 106 111 142 137
rect 168 111 204 137
rect 230 111 236 137
rect -236 75 236 111
rect -236 49 -230 75
rect -204 49 -168 75
rect -142 49 -106 75
rect -80 49 -44 75
rect -18 49 18 75
rect 44 49 80 75
rect 106 49 142 75
rect 168 49 204 75
rect 230 49 236 75
rect -236 13 236 49
rect -236 -13 -230 13
rect -204 -13 -168 13
rect -142 -13 -106 13
rect -80 -13 -44 13
rect -18 -13 18 13
rect 44 -13 80 13
rect 106 -13 142 13
rect 168 -13 204 13
rect 230 -13 236 13
rect -236 -49 236 -13
rect -236 -75 -230 -49
rect -204 -75 -168 -49
rect -142 -75 -106 -49
rect -80 -75 -44 -49
rect -18 -75 18 -49
rect 44 -75 80 -49
rect 106 -75 142 -49
rect 168 -75 204 -49
rect 230 -75 236 -49
rect -236 -111 236 -75
rect -236 -137 -230 -111
rect -204 -137 -168 -111
rect -142 -137 -106 -111
rect -80 -137 -44 -111
rect -18 -137 18 -111
rect 44 -137 80 -111
rect 106 -137 142 -111
rect 168 -137 204 -111
rect 230 -137 236 -111
rect -236 -173 236 -137
rect -236 -199 -230 -173
rect -204 -199 -168 -173
rect -142 -199 -106 -173
rect -80 -199 -44 -173
rect -18 -199 18 -173
rect 44 -199 80 -173
rect 106 -199 142 -173
rect 168 -199 204 -173
rect 230 -199 236 -173
rect -236 -235 236 -199
rect -236 -261 -230 -235
rect -204 -261 -168 -235
rect -142 -261 -106 -235
rect -80 -261 -44 -235
rect -18 -261 18 -235
rect 44 -261 80 -235
rect 106 -261 142 -235
rect 168 -261 204 -235
rect 230 -261 236 -235
rect -236 -297 236 -261
rect -236 -323 -230 -297
rect -204 -323 -168 -297
rect -142 -323 -106 -297
rect -80 -323 -44 -297
rect -18 -323 18 -297
rect 44 -323 80 -297
rect 106 -323 142 -297
rect 168 -323 204 -297
rect 230 -323 236 -297
rect -236 -359 236 -323
rect -236 -385 -230 -359
rect -204 -385 -168 -359
rect -142 -385 -106 -359
rect -80 -385 -44 -359
rect -18 -385 18 -359
rect 44 -385 80 -359
rect 106 -385 142 -359
rect 168 -385 204 -359
rect 230 -385 236 -359
rect -236 -421 236 -385
rect -236 -447 -230 -421
rect -204 -447 -168 -421
rect -142 -447 -106 -421
rect -80 -447 -44 -421
rect -18 -447 18 -421
rect 44 -447 80 -421
rect 106 -447 142 -421
rect 168 -447 204 -421
rect 230 -447 236 -421
rect -236 -483 236 -447
rect -236 -509 -230 -483
rect -204 -509 -168 -483
rect -142 -509 -106 -483
rect -80 -509 -44 -483
rect -18 -509 18 -483
rect 44 -509 80 -483
rect 106 -509 142 -483
rect 168 -509 204 -483
rect 230 -509 236 -483
rect -236 -545 236 -509
rect -236 -571 -230 -545
rect -204 -571 -168 -545
rect -142 -571 -106 -545
rect -80 -571 -44 -545
rect -18 -571 18 -545
rect 44 -571 80 -545
rect 106 -571 142 -545
rect 168 -571 204 -545
rect 230 -571 236 -545
rect -236 -607 236 -571
rect -236 -633 -230 -607
rect -204 -633 -168 -607
rect -142 -633 -106 -607
rect -80 -633 -44 -607
rect -18 -633 18 -607
rect 44 -633 80 -607
rect 106 -633 142 -607
rect 168 -633 204 -607
rect 230 -633 236 -607
rect -236 -669 236 -633
rect -236 -695 -230 -669
rect -204 -695 -168 -669
rect -142 -695 -106 -669
rect -80 -695 -44 -669
rect -18 -695 18 -669
rect 44 -695 80 -669
rect 106 -695 142 -669
rect 168 -695 204 -669
rect 230 -695 236 -669
rect -236 -731 236 -695
rect -236 -757 -230 -731
rect -204 -757 -168 -731
rect -142 -757 -106 -731
rect -80 -757 -44 -731
rect -18 -757 18 -731
rect 44 -757 80 -731
rect 106 -757 142 -731
rect 168 -757 204 -731
rect 230 -757 236 -731
rect -236 -763 236 -757
<< via1 >>
rect -230 731 -204 757
rect -168 731 -142 757
rect -106 731 -80 757
rect -44 731 -18 757
rect 18 731 44 757
rect 80 731 106 757
rect 142 731 168 757
rect 204 731 230 757
rect -230 669 -204 695
rect -168 669 -142 695
rect -106 669 -80 695
rect -44 669 -18 695
rect 18 669 44 695
rect 80 669 106 695
rect 142 669 168 695
rect 204 669 230 695
rect -230 607 -204 633
rect -168 607 -142 633
rect -106 607 -80 633
rect -44 607 -18 633
rect 18 607 44 633
rect 80 607 106 633
rect 142 607 168 633
rect 204 607 230 633
rect -230 545 -204 571
rect -168 545 -142 571
rect -106 545 -80 571
rect -44 545 -18 571
rect 18 545 44 571
rect 80 545 106 571
rect 142 545 168 571
rect 204 545 230 571
rect -230 483 -204 509
rect -168 483 -142 509
rect -106 483 -80 509
rect -44 483 -18 509
rect 18 483 44 509
rect 80 483 106 509
rect 142 483 168 509
rect 204 483 230 509
rect -230 421 -204 447
rect -168 421 -142 447
rect -106 421 -80 447
rect -44 421 -18 447
rect 18 421 44 447
rect 80 421 106 447
rect 142 421 168 447
rect 204 421 230 447
rect -230 359 -204 385
rect -168 359 -142 385
rect -106 359 -80 385
rect -44 359 -18 385
rect 18 359 44 385
rect 80 359 106 385
rect 142 359 168 385
rect 204 359 230 385
rect -230 297 -204 323
rect -168 297 -142 323
rect -106 297 -80 323
rect -44 297 -18 323
rect 18 297 44 323
rect 80 297 106 323
rect 142 297 168 323
rect 204 297 230 323
rect -230 235 -204 261
rect -168 235 -142 261
rect -106 235 -80 261
rect -44 235 -18 261
rect 18 235 44 261
rect 80 235 106 261
rect 142 235 168 261
rect 204 235 230 261
rect -230 173 -204 199
rect -168 173 -142 199
rect -106 173 -80 199
rect -44 173 -18 199
rect 18 173 44 199
rect 80 173 106 199
rect 142 173 168 199
rect 204 173 230 199
rect -230 111 -204 137
rect -168 111 -142 137
rect -106 111 -80 137
rect -44 111 -18 137
rect 18 111 44 137
rect 80 111 106 137
rect 142 111 168 137
rect 204 111 230 137
rect -230 49 -204 75
rect -168 49 -142 75
rect -106 49 -80 75
rect -44 49 -18 75
rect 18 49 44 75
rect 80 49 106 75
rect 142 49 168 75
rect 204 49 230 75
rect -230 -13 -204 13
rect -168 -13 -142 13
rect -106 -13 -80 13
rect -44 -13 -18 13
rect 18 -13 44 13
rect 80 -13 106 13
rect 142 -13 168 13
rect 204 -13 230 13
rect -230 -75 -204 -49
rect -168 -75 -142 -49
rect -106 -75 -80 -49
rect -44 -75 -18 -49
rect 18 -75 44 -49
rect 80 -75 106 -49
rect 142 -75 168 -49
rect 204 -75 230 -49
rect -230 -137 -204 -111
rect -168 -137 -142 -111
rect -106 -137 -80 -111
rect -44 -137 -18 -111
rect 18 -137 44 -111
rect 80 -137 106 -111
rect 142 -137 168 -111
rect 204 -137 230 -111
rect -230 -199 -204 -173
rect -168 -199 -142 -173
rect -106 -199 -80 -173
rect -44 -199 -18 -173
rect 18 -199 44 -173
rect 80 -199 106 -173
rect 142 -199 168 -173
rect 204 -199 230 -173
rect -230 -261 -204 -235
rect -168 -261 -142 -235
rect -106 -261 -80 -235
rect -44 -261 -18 -235
rect 18 -261 44 -235
rect 80 -261 106 -235
rect 142 -261 168 -235
rect 204 -261 230 -235
rect -230 -323 -204 -297
rect -168 -323 -142 -297
rect -106 -323 -80 -297
rect -44 -323 -18 -297
rect 18 -323 44 -297
rect 80 -323 106 -297
rect 142 -323 168 -297
rect 204 -323 230 -297
rect -230 -385 -204 -359
rect -168 -385 -142 -359
rect -106 -385 -80 -359
rect -44 -385 -18 -359
rect 18 -385 44 -359
rect 80 -385 106 -359
rect 142 -385 168 -359
rect 204 -385 230 -359
rect -230 -447 -204 -421
rect -168 -447 -142 -421
rect -106 -447 -80 -421
rect -44 -447 -18 -421
rect 18 -447 44 -421
rect 80 -447 106 -421
rect 142 -447 168 -421
rect 204 -447 230 -421
rect -230 -509 -204 -483
rect -168 -509 -142 -483
rect -106 -509 -80 -483
rect -44 -509 -18 -483
rect 18 -509 44 -483
rect 80 -509 106 -483
rect 142 -509 168 -483
rect 204 -509 230 -483
rect -230 -571 -204 -545
rect -168 -571 -142 -545
rect -106 -571 -80 -545
rect -44 -571 -18 -545
rect 18 -571 44 -545
rect 80 -571 106 -545
rect 142 -571 168 -545
rect 204 -571 230 -545
rect -230 -633 -204 -607
rect -168 -633 -142 -607
rect -106 -633 -80 -607
rect -44 -633 -18 -607
rect 18 -633 44 -607
rect 80 -633 106 -607
rect 142 -633 168 -607
rect 204 -633 230 -607
rect -230 -695 -204 -669
rect -168 -695 -142 -669
rect -106 -695 -80 -669
rect -44 -695 -18 -669
rect 18 -695 44 -669
rect 80 -695 106 -669
rect 142 -695 168 -669
rect 204 -695 230 -669
rect -230 -757 -204 -731
rect -168 -757 -142 -731
rect -106 -757 -80 -731
rect -44 -757 -18 -731
rect 18 -757 44 -731
rect 80 -757 106 -731
rect 142 -757 168 -731
rect 204 -757 230 -731
<< metal2 >>
rect -236 757 236 763
rect -236 731 -230 757
rect -204 731 -168 757
rect -142 731 -106 757
rect -80 731 -44 757
rect -18 731 18 757
rect 44 731 80 757
rect 106 731 142 757
rect 168 731 204 757
rect 230 731 236 757
rect -236 695 236 731
rect -236 669 -230 695
rect -204 669 -168 695
rect -142 669 -106 695
rect -80 669 -44 695
rect -18 669 18 695
rect 44 669 80 695
rect 106 669 142 695
rect 168 669 204 695
rect 230 669 236 695
rect -236 633 236 669
rect -236 607 -230 633
rect -204 607 -168 633
rect -142 607 -106 633
rect -80 607 -44 633
rect -18 607 18 633
rect 44 607 80 633
rect 106 607 142 633
rect 168 607 204 633
rect 230 607 236 633
rect -236 571 236 607
rect -236 545 -230 571
rect -204 545 -168 571
rect -142 545 -106 571
rect -80 545 -44 571
rect -18 545 18 571
rect 44 545 80 571
rect 106 545 142 571
rect 168 545 204 571
rect 230 545 236 571
rect -236 509 236 545
rect -236 483 -230 509
rect -204 483 -168 509
rect -142 483 -106 509
rect -80 483 -44 509
rect -18 483 18 509
rect 44 483 80 509
rect 106 483 142 509
rect 168 483 204 509
rect 230 483 236 509
rect -236 447 236 483
rect -236 421 -230 447
rect -204 421 -168 447
rect -142 421 -106 447
rect -80 421 -44 447
rect -18 421 18 447
rect 44 421 80 447
rect 106 421 142 447
rect 168 421 204 447
rect 230 421 236 447
rect -236 385 236 421
rect -236 359 -230 385
rect -204 359 -168 385
rect -142 359 -106 385
rect -80 359 -44 385
rect -18 359 18 385
rect 44 359 80 385
rect 106 359 142 385
rect 168 359 204 385
rect 230 359 236 385
rect -236 323 236 359
rect -236 297 -230 323
rect -204 297 -168 323
rect -142 297 -106 323
rect -80 297 -44 323
rect -18 297 18 323
rect 44 297 80 323
rect 106 297 142 323
rect 168 297 204 323
rect 230 297 236 323
rect -236 261 236 297
rect -236 235 -230 261
rect -204 235 -168 261
rect -142 235 -106 261
rect -80 235 -44 261
rect -18 235 18 261
rect 44 235 80 261
rect 106 235 142 261
rect 168 235 204 261
rect 230 235 236 261
rect -236 199 236 235
rect -236 173 -230 199
rect -204 173 -168 199
rect -142 173 -106 199
rect -80 173 -44 199
rect -18 173 18 199
rect 44 173 80 199
rect 106 173 142 199
rect 168 173 204 199
rect 230 173 236 199
rect -236 137 236 173
rect -236 111 -230 137
rect -204 111 -168 137
rect -142 111 -106 137
rect -80 111 -44 137
rect -18 111 18 137
rect 44 111 80 137
rect 106 111 142 137
rect 168 111 204 137
rect 230 111 236 137
rect -236 75 236 111
rect -236 49 -230 75
rect -204 49 -168 75
rect -142 49 -106 75
rect -80 49 -44 75
rect -18 49 18 75
rect 44 49 80 75
rect 106 49 142 75
rect 168 49 204 75
rect 230 49 236 75
rect -236 13 236 49
rect -236 -13 -230 13
rect -204 -13 -168 13
rect -142 -13 -106 13
rect -80 -13 -44 13
rect -18 -13 18 13
rect 44 -13 80 13
rect 106 -13 142 13
rect 168 -13 204 13
rect 230 -13 236 13
rect -236 -49 236 -13
rect -236 -75 -230 -49
rect -204 -75 -168 -49
rect -142 -75 -106 -49
rect -80 -75 -44 -49
rect -18 -75 18 -49
rect 44 -75 80 -49
rect 106 -75 142 -49
rect 168 -75 204 -49
rect 230 -75 236 -49
rect -236 -111 236 -75
rect -236 -137 -230 -111
rect -204 -137 -168 -111
rect -142 -137 -106 -111
rect -80 -137 -44 -111
rect -18 -137 18 -111
rect 44 -137 80 -111
rect 106 -137 142 -111
rect 168 -137 204 -111
rect 230 -137 236 -111
rect -236 -173 236 -137
rect -236 -199 -230 -173
rect -204 -199 -168 -173
rect -142 -199 -106 -173
rect -80 -199 -44 -173
rect -18 -199 18 -173
rect 44 -199 80 -173
rect 106 -199 142 -173
rect 168 -199 204 -173
rect 230 -199 236 -173
rect -236 -235 236 -199
rect -236 -261 -230 -235
rect -204 -261 -168 -235
rect -142 -261 -106 -235
rect -80 -261 -44 -235
rect -18 -261 18 -235
rect 44 -261 80 -235
rect 106 -261 142 -235
rect 168 -261 204 -235
rect 230 -261 236 -235
rect -236 -297 236 -261
rect -236 -323 -230 -297
rect -204 -323 -168 -297
rect -142 -323 -106 -297
rect -80 -323 -44 -297
rect -18 -323 18 -297
rect 44 -323 80 -297
rect 106 -323 142 -297
rect 168 -323 204 -297
rect 230 -323 236 -297
rect -236 -359 236 -323
rect -236 -385 -230 -359
rect -204 -385 -168 -359
rect -142 -385 -106 -359
rect -80 -385 -44 -359
rect -18 -385 18 -359
rect 44 -385 80 -359
rect 106 -385 142 -359
rect 168 -385 204 -359
rect 230 -385 236 -359
rect -236 -421 236 -385
rect -236 -447 -230 -421
rect -204 -447 -168 -421
rect -142 -447 -106 -421
rect -80 -447 -44 -421
rect -18 -447 18 -421
rect 44 -447 80 -421
rect 106 -447 142 -421
rect 168 -447 204 -421
rect 230 -447 236 -421
rect -236 -483 236 -447
rect -236 -509 -230 -483
rect -204 -509 -168 -483
rect -142 -509 -106 -483
rect -80 -509 -44 -483
rect -18 -509 18 -483
rect 44 -509 80 -483
rect 106 -509 142 -483
rect 168 -509 204 -483
rect 230 -509 236 -483
rect -236 -545 236 -509
rect -236 -571 -230 -545
rect -204 -571 -168 -545
rect -142 -571 -106 -545
rect -80 -571 -44 -545
rect -18 -571 18 -545
rect 44 -571 80 -545
rect 106 -571 142 -545
rect 168 -571 204 -545
rect 230 -571 236 -545
rect -236 -607 236 -571
rect -236 -633 -230 -607
rect -204 -633 -168 -607
rect -142 -633 -106 -607
rect -80 -633 -44 -607
rect -18 -633 18 -607
rect 44 -633 80 -607
rect 106 -633 142 -607
rect 168 -633 204 -607
rect 230 -633 236 -607
rect -236 -669 236 -633
rect -236 -695 -230 -669
rect -204 -695 -168 -669
rect -142 -695 -106 -669
rect -80 -695 -44 -669
rect -18 -695 18 -669
rect 44 -695 80 -669
rect 106 -695 142 -669
rect 168 -695 204 -669
rect 230 -695 236 -669
rect -236 -731 236 -695
rect -236 -757 -230 -731
rect -204 -757 -168 -731
rect -142 -757 -106 -731
rect -80 -757 -44 -731
rect -18 -757 18 -731
rect 44 -757 80 -731
rect 106 -757 142 -731
rect 168 -757 204 -731
rect 230 -757 236 -731
rect -236 -763 236 -757
<< end >>
