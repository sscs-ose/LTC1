* NGSPICE file created from a2x1mux_mag_flat.ext - technology: gf180mcuC

.subckt a2x1mux_mag_flat IN2 SEL VOUT VDD VSS IN1
X0 IN1 Transmission_gate_mag_0.inv_my_mag_0.OUT VOUT.t36 VDD.t16 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 IN2 SEL.t0 VOUT.t14 VSS.t25 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X2 inv_my_mag_0.OUT SEL.t1 VDD.t3 VDD.t2 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X3 IN1 inv_my_mag_0.OUT VOUT.t7 VSS.t11 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X4 VOUT SEL.t2 IN2.t8 VSS.t24 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X5 IN2 SEL.t3 VOUT.t13 VSS.t23 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X6 IN1 Transmission_gate_mag_0.inv_my_mag_0.OUT VOUT.t35 VDD.t15 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X7 VOUT Transmission_gate_mag_1.inv_my_mag_0.OUT IN2.t19 VDD.t6 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X8 VOUT inv_my_mag_0.OUT IN1.t8 VSS.t10 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X9 IN2 Transmission_gate_mag_1.inv_my_mag_0.OUT VOUT.t22 VDD.t6 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X10 VOUT Transmission_gate_mag_0.inv_my_mag_0.OUT IN1.t17 VDD.t14 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X11 VOUT Transmission_gate_mag_1.inv_my_mag_0.OUT IN2.t17 VDD.t6 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X12 IN1 inv_my_mag_0.OUT VOUT.t6 VSS.t9 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X13 Transmission_gate_mag_0.inv_my_mag_0.OUT inv_my_mag_0.OUT VSS.t8 VSS.t7 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X14 VOUT inv_my_mag_0.OUT IN1.t6 VSS.t6 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X15 VOUT Transmission_gate_mag_0.inv_my_mag_0.OUT IN1.t16 VDD.t13 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X16 VOUT SEL.t4 IN2.t6 VSS.t22 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X17 inv_my_mag_0.OUT SEL.t5 VSS.t21 VSS.t20 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X18 Transmission_gate_mag_0.inv_my_mag_0.OUT inv_my_mag_0.OUT VDD.t1 VDD.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X19 Transmission_gate_mag_1.inv_my_mag_0.OUT SEL.t6 VSS.t19 VSS.t18 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X20 IN2 SEL.t7 VOUT.t11 VSS.t17 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X21 IN2 SEL.t8 VOUT.t29 VSS.t16 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X22 VOUT SEL.t9 IN2.t3 VSS.t15 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X23 IN1 Transmission_gate_mag_0.inv_my_mag_0.OUT VOUT.t34 VDD.t12 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X24 VOUT Transmission_gate_mag_0.inv_my_mag_0.OUT IN1.t14 VDD.t11 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X25 IN1 inv_my_mag_0.OUT VOUT.t5 VSS.t5 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X26 IN2 Transmission_gate_mag_1.inv_my_mag_0.OUT VOUT.t21 VDD.t6 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X27 IN1 Transmission_gate_mag_0.inv_my_mag_0.OUT VOUT.t33 VDD.t10 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X28 VOUT Transmission_gate_mag_1.inv_my_mag_0.OUT IN2.t15 VDD.t6 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X29 IN1 inv_my_mag_0.OUT VOUT.t4 VSS.t4 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X30 IN2 Transmission_gate_mag_1.inv_my_mag_0.OUT VOUT.t20 VDD.t6 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X31 VOUT SEL.t10 IN2.t2 VSS.t14 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X32 Transmission_gate_mag_1.inv_my_mag_0.OUT SEL.t11 VDD.t5 VDD.t4 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X33 IN2 SEL.t12 VOUT.t16 VSS.t13 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X34 VOUT SEL.t13 IN2.t0 VSS.t12 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X35 VOUT inv_my_mag_0.OUT IN1.t3 VSS.t3 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X36 VOUT Transmission_gate_mag_0.inv_my_mag_0.OUT IN1.t12 VDD.t9 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X37 VOUT inv_my_mag_0.OUT IN1.t2 VSS.t2 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X38 IN1 Transmission_gate_mag_0.inv_my_mag_0.OUT VOUT.t32 VDD.t8 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X39 VOUT Transmission_gate_mag_0.inv_my_mag_0.OUT IN1.t10 VDD.t7 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X40 VOUT Transmission_gate_mag_1.inv_my_mag_0.OUT IN2.t13 VDD.t6 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X41 IN1 inv_my_mag_0.OUT VOUT.t3 VSS.t1 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X42 IN2 Transmission_gate_mag_1.inv_my_mag_0.OUT VOUT.t19 VDD.t6 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X43 IN2 Transmission_gate_mag_1.inv_my_mag_0.OUT VOUT.t18 VDD.t6 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X44 VOUT inv_my_mag_0.OUT IN1.t0 VSS.t0 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X45 VOUT Transmission_gate_mag_1.inv_my_mag_0.OUT IN2.t10 VDD.t6 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
R0 VOUT.n54 VOUT.n53 3.16355
R1 VOUT.n19 VOUT.n18 3.16355
R2 VOUT.n39 VOUT.n36 3.15771
R3 VOUT.n44 VOUT.n41 3.15771
R4 VOUT.n49 VOUT.n46 3.15771
R5 VOUT.n14 VOUT.n13 3.15771
R6 VOUT.n9 VOUT.n8 3.15771
R7 VOUT.n4 VOUT.n3 3.15771
R8 VOUT.n54 VOUT.n51 3.15264
R9 VOUT.n19 VOUT.n16 3.15264
R10 VOUT.n39 VOUT.n38 3.1505
R11 VOUT.n44 VOUT.n43 3.1505
R12 VOUT.n49 VOUT.n48 3.1505
R13 VOUT.n58 VOUT.n34 3.1505
R14 VOUT.n14 VOUT.n11 3.1505
R15 VOUT.n9 VOUT.n6 3.1505
R16 VOUT.n4 VOUT.n1 3.1505
R17 VOUT.n25 VOUT.n24 3.1505
R18 VOUT.n59 VOUT.n32 2.93535
R19 VOUT.n28 VOUT.n27 2.93403
R20 VOUT.n60 VOUT.n59 2.54229
R21 VOUT.n29 VOUT.n28 2.54091
R22 VOUT.n30 VOUT 2.40445
R23 VOUT.n32 VOUT.t20 1.8205
R24 VOUT.n32 VOUT.n31 1.8205
R25 VOUT.n36 VOUT.t18 1.8205
R26 VOUT.n36 VOUT.n35 1.8205
R27 VOUT.n41 VOUT.t22 1.8205
R28 VOUT.n41 VOUT.n40 1.8205
R29 VOUT.n46 VOUT.t21 1.8205
R30 VOUT.n46 VOUT.n45 1.8205
R31 VOUT.n53 VOUT.t19 1.8205
R32 VOUT.n53 VOUT.n52 1.8205
R33 VOUT.n27 VOUT.t33 1.8205
R34 VOUT.n27 VOUT.n26 1.8205
R35 VOUT.n18 VOUT.t35 1.8205
R36 VOUT.n18 VOUT.n17 1.8205
R37 VOUT.n13 VOUT.t32 1.8205
R38 VOUT.n13 VOUT.n12 1.8205
R39 VOUT.n8 VOUT.t34 1.8205
R40 VOUT.n8 VOUT.n7 1.8205
R41 VOUT.n3 VOUT.t36 1.8205
R42 VOUT.n3 VOUT.n2 1.8205
R43 VOUT.n34 VOUT.t13 1.6385
R44 VOUT.n34 VOUT.n33 1.6385
R45 VOUT.n38 VOUT.t29 1.6385
R46 VOUT.n38 VOUT.n37 1.6385
R47 VOUT.n43 VOUT.t16 1.6385
R48 VOUT.n43 VOUT.n42 1.6385
R49 VOUT.n48 VOUT.t14 1.6385
R50 VOUT.n48 VOUT.n47 1.6385
R51 VOUT.n51 VOUT.t11 1.6385
R52 VOUT.n51 VOUT.n50 1.6385
R53 VOUT.n24 VOUT.t7 1.6385
R54 VOUT.n24 VOUT.n23 1.6385
R55 VOUT.n16 VOUT.t4 1.6385
R56 VOUT.n16 VOUT.n15 1.6385
R57 VOUT.n11 VOUT.t6 1.6385
R58 VOUT.n11 VOUT.n10 1.6385
R59 VOUT.n6 VOUT.t3 1.6385
R60 VOUT.n6 VOUT.n5 1.6385
R61 VOUT.n1 VOUT.t5 1.6385
R62 VOUT.n1 VOUT.n0 1.6385
R63 VOUT.n60 VOUT.n30 0.773
R64 VOUT.n30 VOUT.n29 0.74925
R65 VOUT.n58 VOUT.n57 0.690059
R66 VOUT.n25 VOUT.n22 0.690059
R67 VOUT.n55 VOUT.n54 0.686845
R68 VOUT.n20 VOUT.n19 0.686845
R69 VOUT.n56 VOUT.n55 0.424029
R70 VOUT.n21 VOUT.n20 0.424029
R71 VOUT.n57 VOUT.n56 0.422706
R72 VOUT.n22 VOUT.n21 0.422706
R73 VOUT.n57 VOUT.n39 0.263882
R74 VOUT.n56 VOUT.n44 0.263882
R75 VOUT.n55 VOUT.n49 0.263882
R76 VOUT.n20 VOUT.n14 0.263882
R77 VOUT.n21 VOUT.n9 0.263882
R78 VOUT.n22 VOUT.n4 0.263882
R79 VOUT.n28 VOUT.n25 0.224176
R80 VOUT.n59 VOUT.n58 0.222853
R81 VOUT.n29 VOUT 0.0946163
R82 VOUT VOUT.n60 0.093312
R83 IN1.n2 IN1.t8 5.34571
R84 IN1.n28 IN1.n0 5.13526
R85 IN1.n27 IN1.n1 4.4205
R86 IN1.n2 IN1.t12 4.4205
R87 IN1.n7 IN1.n4 3.70771
R88 IN1.n13 IN1.n10 3.70771
R89 IN1.n19 IN1.n16 3.70771
R90 IN1.n25 IN1.n22 3.70771
R91 IN1.n7 IN1.n6 2.6005
R92 IN1.n13 IN1.n12 2.6005
R93 IN1.n19 IN1.n18 2.6005
R94 IN1.n25 IN1.n24 2.6005
R95 IN1.n6 IN1.t16 1.8205
R96 IN1.n6 IN1.n5 1.8205
R97 IN1.n12 IN1.t17 1.8205
R98 IN1.n12 IN1.n11 1.8205
R99 IN1.n18 IN1.t10 1.8205
R100 IN1.n18 IN1.n17 1.8205
R101 IN1.n24 IN1.t14 1.8205
R102 IN1.n24 IN1.n23 1.8205
R103 IN1.n4 IN1.t2 1.6385
R104 IN1.n4 IN1.n3 1.6385
R105 IN1.n10 IN1.t3 1.6385
R106 IN1.n10 IN1.n9 1.6385
R107 IN1.n16 IN1.t6 1.6385
R108 IN1.n16 IN1.n15 1.6385
R109 IN1.n22 IN1.t0 1.6385
R110 IN1.n22 IN1.n21 1.6385
R111 IN1.n8 IN1.n2 0.600059
R112 IN1.n27 IN1.n26 0.600059
R113 IN1.n14 IN1.n8 0.361929
R114 IN1.n26 IN1.n20 0.361929
R115 IN1.n20 IN1.n14 0.359071
R116 IN1 IN1.n28 0.282412
R117 IN1.n8 IN1.n7 0.240059
R118 IN1.n14 IN1.n13 0.240059
R119 IN1.n20 IN1.n19 0.240059
R120 IN1.n26 IN1.n25 0.240059
R121 IN1.n28 IN1.n27 0.120941
R122 VDD.n1 VDD.n0 438.12
R123 VDD.n3 VDD.t9 436.957
R124 VDD.n5 VDD.n4 417.5
R125 VDD.n4 VDD.n0 413.366
R126 VDD.t11 VDD.t10 347.827
R127 VDD.t16 VDD.t11 347.827
R128 VDD.t7 VDD.t16 347.827
R129 VDD.t12 VDD.t7 347.827
R130 VDD.t14 VDD.t12 347.827
R131 VDD.t8 VDD.t14 347.827
R132 VDD.t13 VDD.t8 347.827
R133 VDD.t15 VDD.t13 347.827
R134 VDD.t9 VDD.t15 347.827
R135 VDD.n2 VDD.n1 242.417
R136 VDD.n4 VDD.t2 150
R137 VDD.n4 VDD.n3 99.0104
R138 VDD.n2 VDD.t6 91.7103
R139 VDD.n3 VDD.t0 49.5054
R140 VDD.t6 VDD.t4 8.90522
R141 VDD VDD.n2 6.30798
R142 VDD VDD.n5 6.3005
R143 VDD VDD.n0 6.3005
R144 VDD VDD.t3 5.2211
R145 VDD.n7 VDD.t1 5.17584
R146 VDD.n6 VDD.t5 5.17584
R147 VDD VDD.n7 0.0163291
R148 VDD.n6 VDD 0.00185678
R149 VDD.n7 VDD.n6 0.000726131
R150 SEL.n2 SEL.t3 45.8862
R151 SEL.n1 SEL.t11 25.4398
R152 SEL.n0 SEL.t1 25.4398
R153 SEL.n2 SEL.t2 25.0291
R154 SEL.n3 SEL.t8 25.0291
R155 SEL.n4 SEL.t9 25.0291
R156 SEL.n5 SEL.t12 25.0291
R157 SEL.n6 SEL.t13 25.0291
R158 SEL.n7 SEL.t0 25.0291
R159 SEL.n8 SEL.t4 25.0291
R160 SEL.n9 SEL.t7 25.0291
R161 SEL.n10 SEL.t10 21.9714
R162 SEL.n3 SEL.n2 20.8576
R163 SEL.n4 SEL.n3 20.8576
R164 SEL.n5 SEL.n4 20.8576
R165 SEL.n6 SEL.n5 20.8576
R166 SEL.n7 SEL.n6 20.8576
R167 SEL.n8 SEL.n7 20.8576
R168 SEL.n9 SEL.n8 20.8576
R169 SEL.n10 SEL.n9 19.8874
R170 SEL.n1 SEL.t6 17.6975
R171 SEL.n0 SEL.t5 17.6975
R172 SEL.n11 SEL.n10 9.15922
R173 SEL SEL.n1 4.23025
R174 SEL.n12 SEL.n0 4.20407
R175 SEL.n11 SEL 2.26321
R176 SEL.n12 SEL 2.2505
R177 SEL SEL.n13 0.00789726
R178 SEL.n13 SEL.n12 0.00666438
R179 SEL SEL.n11 0.0053
R180 IN2.n0 IN2.t2 5.34571
R181 IN2.n28 IN2.n27 5.13526
R182 IN2.n26 IN2.n25 4.4205
R183 IN2.n0 IN2.t19 4.4205
R184 IN2.n5 IN2.n4 3.70771
R185 IN2.n11 IN2.n10 3.70771
R186 IN2.n17 IN2.n16 3.70771
R187 IN2.n23 IN2.n22 3.70771
R188 IN2.n5 IN2.n2 2.6005
R189 IN2.n11 IN2.n8 2.6005
R190 IN2.n17 IN2.n14 2.6005
R191 IN2.n23 IN2.n20 2.6005
R192 IN2.n2 IN2.t13 1.8205
R193 IN2.n2 IN2.n1 1.8205
R194 IN2.n8 IN2.t17 1.8205
R195 IN2.n8 IN2.n7 1.8205
R196 IN2.n14 IN2.t10 1.8205
R197 IN2.n14 IN2.n13 1.8205
R198 IN2.n20 IN2.t15 1.8205
R199 IN2.n20 IN2.n19 1.8205
R200 IN2.n4 IN2.t6 1.6385
R201 IN2.n4 IN2.n3 1.6385
R202 IN2.n10 IN2.t0 1.6385
R203 IN2.n10 IN2.n9 1.6385
R204 IN2.n16 IN2.t3 1.6385
R205 IN2.n16 IN2.n15 1.6385
R206 IN2.n22 IN2.t8 1.6385
R207 IN2.n22 IN2.n21 1.6385
R208 IN2.n6 IN2.n0 0.598735
R209 IN2.n26 IN2.n24 0.598735
R210 IN2.n12 IN2.n6 0.361929
R211 IN2.n24 IN2.n18 0.361929
R212 IN2.n18 IN2.n12 0.359071
R213 IN2 IN2.n28 0.283735
R214 IN2.n6 IN2.n5 0.238735
R215 IN2.n12 IN2.n11 0.238735
R216 IN2.n18 IN2.n17 0.238735
R217 IN2.n24 IN2.n23 0.238735
R218 IN2.n28 IN2.n26 0.120941
R219 VSS.t11 VSS.t23 22404.1
R220 VSS.t14 VSS.t18 2859.72
R221 VSS.t7 VSS.t10 2859.72
R222 VSS.t20 VSS.n3 2781.66
R223 VSS.t23 VSS.t24 1135.37
R224 VSS.t24 VSS.t16 1135.37
R225 VSS.t16 VSS.t15 1135.37
R226 VSS.t15 VSS.t13 1135.37
R227 VSS.t13 VSS.t12 1135.37
R228 VSS.t12 VSS.t25 1135.37
R229 VSS.t25 VSS.t22 1135.37
R230 VSS.t22 VSS.t17 1135.37
R231 VSS.t17 VSS.t14 1135.37
R232 VSS.t0 VSS.t11 1135.37
R233 VSS.t5 VSS.t0 1135.37
R234 VSS.t6 VSS.t5 1135.37
R235 VSS.t1 VSS.t6 1135.37
R236 VSS.t3 VSS.t1 1135.37
R237 VSS.t9 VSS.t3 1135.37
R238 VSS.t2 VSS.t9 1135.37
R239 VSS.t4 VSS.t2 1135.37
R240 VSS.t10 VSS.t4 1135.37
R241 VSS.t18 VSS.n2 63.8651
R242 VSS.n3 VSS.t7 63.8651
R243 VSS.n4 VSS.t20 63.8651
R244 VSS VSS.t19 9.43421
R245 VSS.n5 VSS.t21 9.43089
R246 VSS.n6 VSS.t8 9.36804
R247 VSS.n2 VSS.n1 5.2005
R248 VSS.n3 VSS.n0 5.2005
R249 VSS.n5 VSS.n4 5.2005
R250 VSS.n6 VSS 0.0765345
R251 VSS VSS.n6 0.0555862
R252 VSS.n1 VSS 0.00839474
R253 VSS VSS.n0 0.00825862
R254 VSS.n1 VSS 0.00128947
R255 VSS.n0 VSS 0.00127586
R256 VSS VSS.n5 0.00127586
C0 SEL Transmission_gate_mag_0.inv_my_mag_0.OUT 0.00848f
C1 inv_my_mag_0.OUT IN1 0.223f
C2 inv_my_mag_0.OUT IN2 0.00111f
C3 SEL IN1 0.00419f
C4 SEL IN2 0.226f
C5 Transmission_gate_mag_1.inv_my_mag_0.OUT VDD 1.32f
C6 VDD VOUT 0.23f
C7 Transmission_gate_mag_1.inv_my_mag_0.OUT VOUT 0.165f
C8 Transmission_gate_mag_0.inv_my_mag_0.OUT VDD 1.33f
C9 Transmission_gate_mag_1.inv_my_mag_0.OUT Transmission_gate_mag_0.inv_my_mag_0.OUT 0.176f
C10 VDD IN1 0.291f
C11 VDD IN2 0.292f
C12 Transmission_gate_mag_1.inv_my_mag_0.OUT IN1 0.0331f
C13 Transmission_gate_mag_1.inv_my_mag_0.OUT IN2 0.591f
C14 Transmission_gate_mag_0.inv_my_mag_0.OUT VOUT 0.165f
C15 VOUT IN1 3.92f
C16 IN2 VOUT 3.92f
C17 Transmission_gate_mag_0.inv_my_mag_0.OUT IN1 0.591f
C18 Transmission_gate_mag_0.inv_my_mag_0.OUT IN2 0.0331f
C19 SEL inv_my_mag_0.OUT 0.177f
C20 IN2 IN1 0.249f
C21 inv_my_mag_0.OUT VDD 0.471f
C22 Transmission_gate_mag_1.inv_my_mag_0.OUT inv_my_mag_0.OUT 0.00208f
C23 SEL VDD 0.631f
C24 Transmission_gate_mag_1.inv_my_mag_0.OUT SEL 0.234f
C25 inv_my_mag_0.OUT VOUT 0.498f
C26 inv_my_mag_0.OUT Transmission_gate_mag_0.inv_my_mag_0.OUT 0.247f
C27 SEL VOUT 0.501f
C28 IN2 VSS 0.43f
C29 Transmission_gate_mag_1.inv_my_mag_0.OUT VSS 1.08f
C30 VOUT VSS 1.82f
C31 Transmission_gate_mag_0.inv_my_mag_0.OUT VSS 1.06f
C32 SEL VSS 3.25f
C33 IN1 VSS 0.429f
C34 inv_my_mag_0.OUT VSS 2.58f
C35 VDD VSS 7.42f
C36 IN2.t19 VSS 0.0774f
C37 IN2.t2 VSS 0.0992f
C38 IN2.n0 VSS 0.36f
C39 IN2.t13 VSS 0.0322f
C40 IN2.n1 VSS 0.0322f
C41 IN2.n2 VSS 0.0645f
C42 IN2.t6 VSS 0.0322f
C43 IN2.n3 VSS 0.0322f
C44 IN2.n4 VSS 0.0841f
C45 IN2.n5 VSS 0.238f
C46 IN2.n6 VSS 0.19f
C47 IN2.t17 VSS 0.0322f
C48 IN2.n7 VSS 0.0322f
C49 IN2.n8 VSS 0.0645f
C50 IN2.t0 VSS 0.0322f
C51 IN2.n9 VSS 0.0322f
C52 IN2.n10 VSS 0.0841f
C53 IN2.n11 VSS 0.238f
C54 IN2.n12 VSS 0.15f
C55 IN2.t10 VSS 0.0322f
C56 IN2.n13 VSS 0.0322f
C57 IN2.n14 VSS 0.0645f
C58 IN2.t3 VSS 0.0322f
C59 IN2.n15 VSS 0.0322f
C60 IN2.n16 VSS 0.0841f
C61 IN2.n17 VSS 0.238f
C62 IN2.n18 VSS 0.15f
C63 IN2.t15 VSS 0.0322f
C64 IN2.n19 VSS 0.0322f
C65 IN2.n20 VSS 0.0645f
C66 IN2.t8 VSS 0.0322f
C67 IN2.n21 VSS 0.0322f
C68 IN2.n22 VSS 0.0841f
C69 IN2.n23 VSS 0.237f
C70 IN2.n24 VSS 0.189f
C71 IN2.n25 VSS 0.0774f
C72 IN2.n26 VSS 0.147f
C73 IN2.n27 VSS 0.0911f
C74 IN2.n28 VSS 0.249f
C75 IN1.n0 VSS 0.0911f
C76 IN1.n1 VSS 0.0774f
C77 IN1.t8 VSS 0.0992f
C78 IN1.t12 VSS 0.0774f
C79 IN1.n2 VSS 0.36f
C80 IN1.t2 VSS 0.0322f
C81 IN1.n3 VSS 0.0322f
C82 IN1.n4 VSS 0.0841f
C83 IN1.t16 VSS 0.0322f
C84 IN1.n5 VSS 0.0322f
C85 IN1.n6 VSS 0.0645f
C86 IN1.n7 VSS 0.238f
C87 IN1.n8 VSS 0.19f
C88 IN1.t3 VSS 0.0322f
C89 IN1.n9 VSS 0.0322f
C90 IN1.n10 VSS 0.0841f
C91 IN1.t17 VSS 0.0322f
C92 IN1.n11 VSS 0.0322f
C93 IN1.n12 VSS 0.0645f
C94 IN1.n13 VSS 0.238f
C95 IN1.n14 VSS 0.15f
C96 IN1.t6 VSS 0.0322f
C97 IN1.n15 VSS 0.0322f
C98 IN1.n16 VSS 0.0841f
C99 IN1.t10 VSS 0.0322f
C100 IN1.n17 VSS 0.0322f
C101 IN1.n18 VSS 0.0645f
C102 IN1.n19 VSS 0.238f
C103 IN1.n20 VSS 0.15f
C104 IN1.t0 VSS 0.0322f
C105 IN1.n21 VSS 0.0322f
C106 IN1.n22 VSS 0.0841f
C107 IN1.t14 VSS 0.0322f
C108 IN1.n23 VSS 0.0322f
C109 IN1.n24 VSS 0.0645f
C110 IN1.n25 VSS 0.238f
C111 IN1.n26 VSS 0.188f
C112 IN1.n27 VSS 0.147f
C113 IN1.n28 VSS 0.249f
C114 VOUT.t5 VSS 0.032f
C115 VOUT.n0 VSS 0.032f
C116 VOUT.n1 VSS 0.0641f
C117 VOUT.t36 VSS 0.032f
C118 VOUT.n2 VSS 0.032f
C119 VOUT.n3 VSS 0.087f
C120 VOUT.n4 VSS 0.237f
C121 VOUT.t3 VSS 0.032f
C122 VOUT.n5 VSS 0.032f
C123 VOUT.n6 VSS 0.0641f
C124 VOUT.t34 VSS 0.032f
C125 VOUT.n7 VSS 0.032f
C126 VOUT.n8 VSS 0.087f
C127 VOUT.n9 VSS 0.237f
C128 VOUT.t6 VSS 0.032f
C129 VOUT.n10 VSS 0.032f
C130 VOUT.n11 VSS 0.0641f
C131 VOUT.t32 VSS 0.032f
C132 VOUT.n12 VSS 0.032f
C133 VOUT.n13 VSS 0.087f
C134 VOUT.n14 VSS 0.237f
C135 VOUT.t4 VSS 0.032f
C136 VOUT.n15 VSS 0.032f
C137 VOUT.n16 VSS 0.0641f
C138 VOUT.t35 VSS 0.032f
C139 VOUT.n17 VSS 0.032f
C140 VOUT.n18 VSS 0.0871f
C141 VOUT.n19 VSS 0.312f
C142 VOUT.n20 VSS 0.223f
C143 VOUT.n21 VSS 0.176f
C144 VOUT.n22 VSS 0.223f
C145 VOUT.t7 VSS 0.032f
C146 VOUT.n23 VSS 0.032f
C147 VOUT.n24 VSS 0.0641f
C148 VOUT.n25 VSS 0.153f
C149 VOUT.t33 VSS 0.032f
C150 VOUT.n26 VSS 0.032f
C151 VOUT.n27 VSS 0.0748f
C152 VOUT.n28 VSS 0.18f
C153 VOUT.n29 VSS 0.263f
C154 VOUT.n30 VSS 0.273f
C155 VOUT.t20 VSS 0.032f
C156 VOUT.n31 VSS 0.032f
C157 VOUT.n32 VSS 0.0749f
C158 VOUT.t13 VSS 0.032f
C159 VOUT.n33 VSS 0.032f
C160 VOUT.n34 VSS 0.0641f
C161 VOUT.t18 VSS 0.032f
C162 VOUT.n35 VSS 0.032f
C163 VOUT.n36 VSS 0.087f
C164 VOUT.t29 VSS 0.032f
C165 VOUT.n37 VSS 0.032f
C166 VOUT.n38 VSS 0.0641f
C167 VOUT.n39 VSS 0.237f
C168 VOUT.t22 VSS 0.032f
C169 VOUT.n40 VSS 0.032f
C170 VOUT.n41 VSS 0.087f
C171 VOUT.t16 VSS 0.032f
C172 VOUT.n42 VSS 0.032f
C173 VOUT.n43 VSS 0.0641f
C174 VOUT.n44 VSS 0.237f
C175 VOUT.t21 VSS 0.032f
C176 VOUT.n45 VSS 0.032f
C177 VOUT.n46 VSS 0.087f
C178 VOUT.t14 VSS 0.032f
C179 VOUT.n47 VSS 0.032f
C180 VOUT.n48 VSS 0.0641f
C181 VOUT.n49 VSS 0.237f
C182 VOUT.t11 VSS 0.032f
C183 VOUT.n50 VSS 0.032f
C184 VOUT.n51 VSS 0.0641f
C185 VOUT.t19 VSS 0.032f
C186 VOUT.n52 VSS 0.032f
C187 VOUT.n53 VSS 0.0871f
C188 VOUT.n54 VSS 0.312f
C189 VOUT.n55 VSS 0.223f
C190 VOUT.n56 VSS 0.176f
C191 VOUT.n57 VSS 0.223f
C192 VOUT.n58 VSS 0.153f
C193 VOUT.n59 VSS 0.18f
C194 VOUT.n60 VSS 0.267f
.ends

