magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -4162 -2230 4162 2230
<< nwell >>
rect -2162 -230 2162 230
<< pmos >>
rect -1988 -100 -1888 100
rect -1784 -100 -1684 100
rect -1580 -100 -1480 100
rect -1376 -100 -1276 100
rect -1172 -100 -1072 100
rect -968 -100 -868 100
rect -764 -100 -664 100
rect -560 -100 -460 100
rect -356 -100 -256 100
rect -152 -100 -52 100
rect 52 -100 152 100
rect 256 -100 356 100
rect 460 -100 560 100
rect 664 -100 764 100
rect 868 -100 968 100
rect 1072 -100 1172 100
rect 1276 -100 1376 100
rect 1480 -100 1580 100
rect 1684 -100 1784 100
rect 1888 -100 1988 100
<< pdiff >>
rect -2076 70 -1988 100
rect -2076 -70 -2063 70
rect -2017 -70 -1988 70
rect -2076 -100 -1988 -70
rect -1888 70 -1784 100
rect -1888 -70 -1859 70
rect -1813 -70 -1784 70
rect -1888 -100 -1784 -70
rect -1684 70 -1580 100
rect -1684 -70 -1655 70
rect -1609 -70 -1580 70
rect -1684 -100 -1580 -70
rect -1480 70 -1376 100
rect -1480 -70 -1451 70
rect -1405 -70 -1376 70
rect -1480 -100 -1376 -70
rect -1276 70 -1172 100
rect -1276 -70 -1247 70
rect -1201 -70 -1172 70
rect -1276 -100 -1172 -70
rect -1072 70 -968 100
rect -1072 -70 -1043 70
rect -997 -70 -968 70
rect -1072 -100 -968 -70
rect -868 70 -764 100
rect -868 -70 -839 70
rect -793 -70 -764 70
rect -868 -100 -764 -70
rect -664 70 -560 100
rect -664 -70 -635 70
rect -589 -70 -560 70
rect -664 -100 -560 -70
rect -460 70 -356 100
rect -460 -70 -431 70
rect -385 -70 -356 70
rect -460 -100 -356 -70
rect -256 70 -152 100
rect -256 -70 -227 70
rect -181 -70 -152 70
rect -256 -100 -152 -70
rect -52 70 52 100
rect -52 -70 -23 70
rect 23 -70 52 70
rect -52 -100 52 -70
rect 152 70 256 100
rect 152 -70 181 70
rect 227 -70 256 70
rect 152 -100 256 -70
rect 356 70 460 100
rect 356 -70 385 70
rect 431 -70 460 70
rect 356 -100 460 -70
rect 560 70 664 100
rect 560 -70 589 70
rect 635 -70 664 70
rect 560 -100 664 -70
rect 764 70 868 100
rect 764 -70 793 70
rect 839 -70 868 70
rect 764 -100 868 -70
rect 968 70 1072 100
rect 968 -70 997 70
rect 1043 -70 1072 70
rect 968 -100 1072 -70
rect 1172 70 1276 100
rect 1172 -70 1201 70
rect 1247 -70 1276 70
rect 1172 -100 1276 -70
rect 1376 70 1480 100
rect 1376 -70 1405 70
rect 1451 -70 1480 70
rect 1376 -100 1480 -70
rect 1580 70 1684 100
rect 1580 -70 1609 70
rect 1655 -70 1684 70
rect 1580 -100 1684 -70
rect 1784 70 1888 100
rect 1784 -70 1813 70
rect 1859 -70 1888 70
rect 1784 -100 1888 -70
rect 1988 70 2076 100
rect 1988 -70 2017 70
rect 2063 -70 2076 70
rect 1988 -100 2076 -70
<< pdiffc >>
rect -2063 -70 -2017 70
rect -1859 -70 -1813 70
rect -1655 -70 -1609 70
rect -1451 -70 -1405 70
rect -1247 -70 -1201 70
rect -1043 -70 -997 70
rect -839 -70 -793 70
rect -635 -70 -589 70
rect -431 -70 -385 70
rect -227 -70 -181 70
rect -23 -70 23 70
rect 181 -70 227 70
rect 385 -70 431 70
rect 589 -70 635 70
rect 793 -70 839 70
rect 997 -70 1043 70
rect 1201 -70 1247 70
rect 1405 -70 1451 70
rect 1609 -70 1655 70
rect 1813 -70 1859 70
rect 2017 -70 2063 70
<< polysilicon >>
rect -1988 100 -1888 144
rect -1784 100 -1684 144
rect -1580 100 -1480 144
rect -1376 100 -1276 144
rect -1172 100 -1072 144
rect -968 100 -868 144
rect -764 100 -664 144
rect -560 100 -460 144
rect -356 100 -256 144
rect -152 100 -52 144
rect 52 100 152 144
rect 256 100 356 144
rect 460 100 560 144
rect 664 100 764 144
rect 868 100 968 144
rect 1072 100 1172 144
rect 1276 100 1376 144
rect 1480 100 1580 144
rect 1684 100 1784 144
rect 1888 100 1988 144
rect -1988 -144 -1888 -100
rect -1784 -144 -1684 -100
rect -1580 -144 -1480 -100
rect -1376 -144 -1276 -100
rect -1172 -144 -1072 -100
rect -968 -144 -868 -100
rect -764 -144 -664 -100
rect -560 -144 -460 -100
rect -356 -144 -256 -100
rect -152 -144 -52 -100
rect 52 -144 152 -100
rect 256 -144 356 -100
rect 460 -144 560 -100
rect 664 -144 764 -100
rect 868 -144 968 -100
rect 1072 -144 1172 -100
rect 1276 -144 1376 -100
rect 1480 -144 1580 -100
rect 1684 -144 1784 -100
rect 1888 -144 1988 -100
<< metal1 >>
rect -2063 70 -2017 98
rect -2063 -98 -2017 -70
rect -1859 70 -1813 98
rect -1859 -98 -1813 -70
rect -1655 70 -1609 98
rect -1655 -98 -1609 -70
rect -1451 70 -1405 98
rect -1451 -98 -1405 -70
rect -1247 70 -1201 98
rect -1247 -98 -1201 -70
rect -1043 70 -997 98
rect -1043 -98 -997 -70
rect -839 70 -793 98
rect -839 -98 -793 -70
rect -635 70 -589 98
rect -635 -98 -589 -70
rect -431 70 -385 98
rect -431 -98 -385 -70
rect -227 70 -181 98
rect -227 -98 -181 -70
rect -23 70 23 98
rect -23 -98 23 -70
rect 181 70 227 98
rect 181 -98 227 -70
rect 385 70 431 98
rect 385 -98 431 -70
rect 589 70 635 98
rect 589 -98 635 -70
rect 793 70 839 98
rect 793 -98 839 -70
rect 997 70 1043 98
rect 997 -98 1043 -70
rect 1201 70 1247 98
rect 1201 -98 1247 -70
rect 1405 70 1451 98
rect 1405 -98 1451 -70
rect 1609 70 1655 98
rect 1609 -98 1655 -70
rect 1813 70 1859 98
rect 1813 -98 1859 -70
rect 2017 70 2063 98
rect 2017 -98 2063 -70
<< end >>
