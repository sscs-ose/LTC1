magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1205 -1763 1205 1763
<< metal1 >>
rect -205 757 205 763
rect -205 731 -199 757
rect -173 731 -137 757
rect -111 731 -75 757
rect -49 731 -13 757
rect 13 731 49 757
rect 75 731 111 757
rect 137 731 173 757
rect 199 731 205 757
rect -205 695 205 731
rect -205 669 -199 695
rect -173 669 -137 695
rect -111 669 -75 695
rect -49 669 -13 695
rect 13 669 49 695
rect 75 669 111 695
rect 137 669 173 695
rect 199 669 205 695
rect -205 633 205 669
rect -205 607 -199 633
rect -173 607 -137 633
rect -111 607 -75 633
rect -49 607 -13 633
rect 13 607 49 633
rect 75 607 111 633
rect 137 607 173 633
rect 199 607 205 633
rect -205 571 205 607
rect -205 545 -199 571
rect -173 545 -137 571
rect -111 545 -75 571
rect -49 545 -13 571
rect 13 545 49 571
rect 75 545 111 571
rect 137 545 173 571
rect 199 545 205 571
rect -205 509 205 545
rect -205 483 -199 509
rect -173 483 -137 509
rect -111 483 -75 509
rect -49 483 -13 509
rect 13 483 49 509
rect 75 483 111 509
rect 137 483 173 509
rect 199 483 205 509
rect -205 447 205 483
rect -205 421 -199 447
rect -173 421 -137 447
rect -111 421 -75 447
rect -49 421 -13 447
rect 13 421 49 447
rect 75 421 111 447
rect 137 421 173 447
rect 199 421 205 447
rect -205 385 205 421
rect -205 359 -199 385
rect -173 359 -137 385
rect -111 359 -75 385
rect -49 359 -13 385
rect 13 359 49 385
rect 75 359 111 385
rect 137 359 173 385
rect 199 359 205 385
rect -205 323 205 359
rect -205 297 -199 323
rect -173 297 -137 323
rect -111 297 -75 323
rect -49 297 -13 323
rect 13 297 49 323
rect 75 297 111 323
rect 137 297 173 323
rect 199 297 205 323
rect -205 261 205 297
rect -205 235 -199 261
rect -173 235 -137 261
rect -111 235 -75 261
rect -49 235 -13 261
rect 13 235 49 261
rect 75 235 111 261
rect 137 235 173 261
rect 199 235 205 261
rect -205 199 205 235
rect -205 173 -199 199
rect -173 173 -137 199
rect -111 173 -75 199
rect -49 173 -13 199
rect 13 173 49 199
rect 75 173 111 199
rect 137 173 173 199
rect 199 173 205 199
rect -205 137 205 173
rect -205 111 -199 137
rect -173 111 -137 137
rect -111 111 -75 137
rect -49 111 -13 137
rect 13 111 49 137
rect 75 111 111 137
rect 137 111 173 137
rect 199 111 205 137
rect -205 75 205 111
rect -205 49 -199 75
rect -173 49 -137 75
rect -111 49 -75 75
rect -49 49 -13 75
rect 13 49 49 75
rect 75 49 111 75
rect 137 49 173 75
rect 199 49 205 75
rect -205 13 205 49
rect -205 -13 -199 13
rect -173 -13 -137 13
rect -111 -13 -75 13
rect -49 -13 -13 13
rect 13 -13 49 13
rect 75 -13 111 13
rect 137 -13 173 13
rect 199 -13 205 13
rect -205 -49 205 -13
rect -205 -75 -199 -49
rect -173 -75 -137 -49
rect -111 -75 -75 -49
rect -49 -75 -13 -49
rect 13 -75 49 -49
rect 75 -75 111 -49
rect 137 -75 173 -49
rect 199 -75 205 -49
rect -205 -111 205 -75
rect -205 -137 -199 -111
rect -173 -137 -137 -111
rect -111 -137 -75 -111
rect -49 -137 -13 -111
rect 13 -137 49 -111
rect 75 -137 111 -111
rect 137 -137 173 -111
rect 199 -137 205 -111
rect -205 -173 205 -137
rect -205 -199 -199 -173
rect -173 -199 -137 -173
rect -111 -199 -75 -173
rect -49 -199 -13 -173
rect 13 -199 49 -173
rect 75 -199 111 -173
rect 137 -199 173 -173
rect 199 -199 205 -173
rect -205 -235 205 -199
rect -205 -261 -199 -235
rect -173 -261 -137 -235
rect -111 -261 -75 -235
rect -49 -261 -13 -235
rect 13 -261 49 -235
rect 75 -261 111 -235
rect 137 -261 173 -235
rect 199 -261 205 -235
rect -205 -297 205 -261
rect -205 -323 -199 -297
rect -173 -323 -137 -297
rect -111 -323 -75 -297
rect -49 -323 -13 -297
rect 13 -323 49 -297
rect 75 -323 111 -297
rect 137 -323 173 -297
rect 199 -323 205 -297
rect -205 -359 205 -323
rect -205 -385 -199 -359
rect -173 -385 -137 -359
rect -111 -385 -75 -359
rect -49 -385 -13 -359
rect 13 -385 49 -359
rect 75 -385 111 -359
rect 137 -385 173 -359
rect 199 -385 205 -359
rect -205 -421 205 -385
rect -205 -447 -199 -421
rect -173 -447 -137 -421
rect -111 -447 -75 -421
rect -49 -447 -13 -421
rect 13 -447 49 -421
rect 75 -447 111 -421
rect 137 -447 173 -421
rect 199 -447 205 -421
rect -205 -483 205 -447
rect -205 -509 -199 -483
rect -173 -509 -137 -483
rect -111 -509 -75 -483
rect -49 -509 -13 -483
rect 13 -509 49 -483
rect 75 -509 111 -483
rect 137 -509 173 -483
rect 199 -509 205 -483
rect -205 -545 205 -509
rect -205 -571 -199 -545
rect -173 -571 -137 -545
rect -111 -571 -75 -545
rect -49 -571 -13 -545
rect 13 -571 49 -545
rect 75 -571 111 -545
rect 137 -571 173 -545
rect 199 -571 205 -545
rect -205 -607 205 -571
rect -205 -633 -199 -607
rect -173 -633 -137 -607
rect -111 -633 -75 -607
rect -49 -633 -13 -607
rect 13 -633 49 -607
rect 75 -633 111 -607
rect 137 -633 173 -607
rect 199 -633 205 -607
rect -205 -669 205 -633
rect -205 -695 -199 -669
rect -173 -695 -137 -669
rect -111 -695 -75 -669
rect -49 -695 -13 -669
rect 13 -695 49 -669
rect 75 -695 111 -669
rect 137 -695 173 -669
rect 199 -695 205 -669
rect -205 -731 205 -695
rect -205 -757 -199 -731
rect -173 -757 -137 -731
rect -111 -757 -75 -731
rect -49 -757 -13 -731
rect 13 -757 49 -731
rect 75 -757 111 -731
rect 137 -757 173 -731
rect 199 -757 205 -731
rect -205 -763 205 -757
<< via1 >>
rect -199 731 -173 757
rect -137 731 -111 757
rect -75 731 -49 757
rect -13 731 13 757
rect 49 731 75 757
rect 111 731 137 757
rect 173 731 199 757
rect -199 669 -173 695
rect -137 669 -111 695
rect -75 669 -49 695
rect -13 669 13 695
rect 49 669 75 695
rect 111 669 137 695
rect 173 669 199 695
rect -199 607 -173 633
rect -137 607 -111 633
rect -75 607 -49 633
rect -13 607 13 633
rect 49 607 75 633
rect 111 607 137 633
rect 173 607 199 633
rect -199 545 -173 571
rect -137 545 -111 571
rect -75 545 -49 571
rect -13 545 13 571
rect 49 545 75 571
rect 111 545 137 571
rect 173 545 199 571
rect -199 483 -173 509
rect -137 483 -111 509
rect -75 483 -49 509
rect -13 483 13 509
rect 49 483 75 509
rect 111 483 137 509
rect 173 483 199 509
rect -199 421 -173 447
rect -137 421 -111 447
rect -75 421 -49 447
rect -13 421 13 447
rect 49 421 75 447
rect 111 421 137 447
rect 173 421 199 447
rect -199 359 -173 385
rect -137 359 -111 385
rect -75 359 -49 385
rect -13 359 13 385
rect 49 359 75 385
rect 111 359 137 385
rect 173 359 199 385
rect -199 297 -173 323
rect -137 297 -111 323
rect -75 297 -49 323
rect -13 297 13 323
rect 49 297 75 323
rect 111 297 137 323
rect 173 297 199 323
rect -199 235 -173 261
rect -137 235 -111 261
rect -75 235 -49 261
rect -13 235 13 261
rect 49 235 75 261
rect 111 235 137 261
rect 173 235 199 261
rect -199 173 -173 199
rect -137 173 -111 199
rect -75 173 -49 199
rect -13 173 13 199
rect 49 173 75 199
rect 111 173 137 199
rect 173 173 199 199
rect -199 111 -173 137
rect -137 111 -111 137
rect -75 111 -49 137
rect -13 111 13 137
rect 49 111 75 137
rect 111 111 137 137
rect 173 111 199 137
rect -199 49 -173 75
rect -137 49 -111 75
rect -75 49 -49 75
rect -13 49 13 75
rect 49 49 75 75
rect 111 49 137 75
rect 173 49 199 75
rect -199 -13 -173 13
rect -137 -13 -111 13
rect -75 -13 -49 13
rect -13 -13 13 13
rect 49 -13 75 13
rect 111 -13 137 13
rect 173 -13 199 13
rect -199 -75 -173 -49
rect -137 -75 -111 -49
rect -75 -75 -49 -49
rect -13 -75 13 -49
rect 49 -75 75 -49
rect 111 -75 137 -49
rect 173 -75 199 -49
rect -199 -137 -173 -111
rect -137 -137 -111 -111
rect -75 -137 -49 -111
rect -13 -137 13 -111
rect 49 -137 75 -111
rect 111 -137 137 -111
rect 173 -137 199 -111
rect -199 -199 -173 -173
rect -137 -199 -111 -173
rect -75 -199 -49 -173
rect -13 -199 13 -173
rect 49 -199 75 -173
rect 111 -199 137 -173
rect 173 -199 199 -173
rect -199 -261 -173 -235
rect -137 -261 -111 -235
rect -75 -261 -49 -235
rect -13 -261 13 -235
rect 49 -261 75 -235
rect 111 -261 137 -235
rect 173 -261 199 -235
rect -199 -323 -173 -297
rect -137 -323 -111 -297
rect -75 -323 -49 -297
rect -13 -323 13 -297
rect 49 -323 75 -297
rect 111 -323 137 -297
rect 173 -323 199 -297
rect -199 -385 -173 -359
rect -137 -385 -111 -359
rect -75 -385 -49 -359
rect -13 -385 13 -359
rect 49 -385 75 -359
rect 111 -385 137 -359
rect 173 -385 199 -359
rect -199 -447 -173 -421
rect -137 -447 -111 -421
rect -75 -447 -49 -421
rect -13 -447 13 -421
rect 49 -447 75 -421
rect 111 -447 137 -421
rect 173 -447 199 -421
rect -199 -509 -173 -483
rect -137 -509 -111 -483
rect -75 -509 -49 -483
rect -13 -509 13 -483
rect 49 -509 75 -483
rect 111 -509 137 -483
rect 173 -509 199 -483
rect -199 -571 -173 -545
rect -137 -571 -111 -545
rect -75 -571 -49 -545
rect -13 -571 13 -545
rect 49 -571 75 -545
rect 111 -571 137 -545
rect 173 -571 199 -545
rect -199 -633 -173 -607
rect -137 -633 -111 -607
rect -75 -633 -49 -607
rect -13 -633 13 -607
rect 49 -633 75 -607
rect 111 -633 137 -607
rect 173 -633 199 -607
rect -199 -695 -173 -669
rect -137 -695 -111 -669
rect -75 -695 -49 -669
rect -13 -695 13 -669
rect 49 -695 75 -669
rect 111 -695 137 -669
rect 173 -695 199 -669
rect -199 -757 -173 -731
rect -137 -757 -111 -731
rect -75 -757 -49 -731
rect -13 -757 13 -731
rect 49 -757 75 -731
rect 111 -757 137 -731
rect 173 -757 199 -731
<< metal2 >>
rect -205 757 205 763
rect -205 731 -199 757
rect -173 731 -137 757
rect -111 731 -75 757
rect -49 731 -13 757
rect 13 731 49 757
rect 75 731 111 757
rect 137 731 173 757
rect 199 731 205 757
rect -205 695 205 731
rect -205 669 -199 695
rect -173 669 -137 695
rect -111 669 -75 695
rect -49 669 -13 695
rect 13 669 49 695
rect 75 669 111 695
rect 137 669 173 695
rect 199 669 205 695
rect -205 633 205 669
rect -205 607 -199 633
rect -173 607 -137 633
rect -111 607 -75 633
rect -49 607 -13 633
rect 13 607 49 633
rect 75 607 111 633
rect 137 607 173 633
rect 199 607 205 633
rect -205 571 205 607
rect -205 545 -199 571
rect -173 545 -137 571
rect -111 545 -75 571
rect -49 545 -13 571
rect 13 545 49 571
rect 75 545 111 571
rect 137 545 173 571
rect 199 545 205 571
rect -205 509 205 545
rect -205 483 -199 509
rect -173 483 -137 509
rect -111 483 -75 509
rect -49 483 -13 509
rect 13 483 49 509
rect 75 483 111 509
rect 137 483 173 509
rect 199 483 205 509
rect -205 447 205 483
rect -205 421 -199 447
rect -173 421 -137 447
rect -111 421 -75 447
rect -49 421 -13 447
rect 13 421 49 447
rect 75 421 111 447
rect 137 421 173 447
rect 199 421 205 447
rect -205 385 205 421
rect -205 359 -199 385
rect -173 359 -137 385
rect -111 359 -75 385
rect -49 359 -13 385
rect 13 359 49 385
rect 75 359 111 385
rect 137 359 173 385
rect 199 359 205 385
rect -205 323 205 359
rect -205 297 -199 323
rect -173 297 -137 323
rect -111 297 -75 323
rect -49 297 -13 323
rect 13 297 49 323
rect 75 297 111 323
rect 137 297 173 323
rect 199 297 205 323
rect -205 261 205 297
rect -205 235 -199 261
rect -173 235 -137 261
rect -111 235 -75 261
rect -49 235 -13 261
rect 13 235 49 261
rect 75 235 111 261
rect 137 235 173 261
rect 199 235 205 261
rect -205 199 205 235
rect -205 173 -199 199
rect -173 173 -137 199
rect -111 173 -75 199
rect -49 173 -13 199
rect 13 173 49 199
rect 75 173 111 199
rect 137 173 173 199
rect 199 173 205 199
rect -205 137 205 173
rect -205 111 -199 137
rect -173 111 -137 137
rect -111 111 -75 137
rect -49 111 -13 137
rect 13 111 49 137
rect 75 111 111 137
rect 137 111 173 137
rect 199 111 205 137
rect -205 75 205 111
rect -205 49 -199 75
rect -173 49 -137 75
rect -111 49 -75 75
rect -49 49 -13 75
rect 13 49 49 75
rect 75 49 111 75
rect 137 49 173 75
rect 199 49 205 75
rect -205 13 205 49
rect -205 -13 -199 13
rect -173 -13 -137 13
rect -111 -13 -75 13
rect -49 -13 -13 13
rect 13 -13 49 13
rect 75 -13 111 13
rect 137 -13 173 13
rect 199 -13 205 13
rect -205 -49 205 -13
rect -205 -75 -199 -49
rect -173 -75 -137 -49
rect -111 -75 -75 -49
rect -49 -75 -13 -49
rect 13 -75 49 -49
rect 75 -75 111 -49
rect 137 -75 173 -49
rect 199 -75 205 -49
rect -205 -111 205 -75
rect -205 -137 -199 -111
rect -173 -137 -137 -111
rect -111 -137 -75 -111
rect -49 -137 -13 -111
rect 13 -137 49 -111
rect 75 -137 111 -111
rect 137 -137 173 -111
rect 199 -137 205 -111
rect -205 -173 205 -137
rect -205 -199 -199 -173
rect -173 -199 -137 -173
rect -111 -199 -75 -173
rect -49 -199 -13 -173
rect 13 -199 49 -173
rect 75 -199 111 -173
rect 137 -199 173 -173
rect 199 -199 205 -173
rect -205 -235 205 -199
rect -205 -261 -199 -235
rect -173 -261 -137 -235
rect -111 -261 -75 -235
rect -49 -261 -13 -235
rect 13 -261 49 -235
rect 75 -261 111 -235
rect 137 -261 173 -235
rect 199 -261 205 -235
rect -205 -297 205 -261
rect -205 -323 -199 -297
rect -173 -323 -137 -297
rect -111 -323 -75 -297
rect -49 -323 -13 -297
rect 13 -323 49 -297
rect 75 -323 111 -297
rect 137 -323 173 -297
rect 199 -323 205 -297
rect -205 -359 205 -323
rect -205 -385 -199 -359
rect -173 -385 -137 -359
rect -111 -385 -75 -359
rect -49 -385 -13 -359
rect 13 -385 49 -359
rect 75 -385 111 -359
rect 137 -385 173 -359
rect 199 -385 205 -359
rect -205 -421 205 -385
rect -205 -447 -199 -421
rect -173 -447 -137 -421
rect -111 -447 -75 -421
rect -49 -447 -13 -421
rect 13 -447 49 -421
rect 75 -447 111 -421
rect 137 -447 173 -421
rect 199 -447 205 -421
rect -205 -483 205 -447
rect -205 -509 -199 -483
rect -173 -509 -137 -483
rect -111 -509 -75 -483
rect -49 -509 -13 -483
rect 13 -509 49 -483
rect 75 -509 111 -483
rect 137 -509 173 -483
rect 199 -509 205 -483
rect -205 -545 205 -509
rect -205 -571 -199 -545
rect -173 -571 -137 -545
rect -111 -571 -75 -545
rect -49 -571 -13 -545
rect 13 -571 49 -545
rect 75 -571 111 -545
rect 137 -571 173 -545
rect 199 -571 205 -545
rect -205 -607 205 -571
rect -205 -633 -199 -607
rect -173 -633 -137 -607
rect -111 -633 -75 -607
rect -49 -633 -13 -607
rect 13 -633 49 -607
rect 75 -633 111 -607
rect 137 -633 173 -607
rect 199 -633 205 -607
rect -205 -669 205 -633
rect -205 -695 -199 -669
rect -173 -695 -137 -669
rect -111 -695 -75 -669
rect -49 -695 -13 -669
rect 13 -695 49 -669
rect 75 -695 111 -669
rect 137 -695 173 -669
rect 199 -695 205 -669
rect -205 -731 205 -695
rect -205 -757 -199 -731
rect -173 -757 -137 -731
rect -111 -757 -75 -731
rect -49 -757 -13 -731
rect 13 -757 49 -731
rect 75 -757 111 -731
rect 137 -757 173 -731
rect 199 -757 205 -731
rect -205 -763 205 -757
<< end >>
