magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1305 1019 1305
<< metal2 >>
rect -19 300 19 305
rect -19 -300 -14 300
rect 14 -300 19 300
rect -19 -305 19 -300
<< via2 >>
rect -14 -300 14 300
<< metal3 >>
rect -19 300 19 305
rect -19 -300 -14 300
rect 14 -300 19 300
rect -19 -305 19 -300
<< end >>
