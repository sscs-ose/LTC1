magic
tech gf180mcuC
magscale 1 10
timestamp 1690963719
<< error_p >>
rect -538 247 -527 293
rect -370 247 -359 293
rect -202 247 -191 293
rect -34 247 -23 293
rect 134 247 145 293
rect 302 247 313 293
rect 470 247 481 293
rect -538 67 -527 113
rect -370 67 -359 113
rect -202 67 -191 113
rect -34 67 -23 113
rect 134 67 145 113
rect 302 67 313 113
rect 470 67 481 113
rect -538 -113 -527 -67
rect -370 -113 -359 -67
rect -202 -113 -191 -67
rect -34 -113 -23 -67
rect 134 -113 145 -67
rect 302 -113 313 -67
rect 470 -113 481 -67
rect -538 -293 -527 -247
rect -370 -293 -359 -247
rect -202 -293 -191 -247
rect -34 -293 -23 -247
rect 134 -293 145 -247
rect 302 -293 313 -247
rect 470 -293 481 -247
<< nwell >>
rect -626 -429 626 429
<< pmos >>
rect -448 248 -392 292
rect -280 248 -224 292
rect -112 248 -56 292
rect 56 248 112 292
rect 224 248 280 292
rect 392 248 448 292
rect -448 68 -392 112
rect -280 68 -224 112
rect -112 68 -56 112
rect 56 68 112 112
rect 224 68 280 112
rect 392 68 448 112
rect -448 -112 -392 -68
rect -280 -112 -224 -68
rect -112 -112 -56 -68
rect 56 -112 112 -68
rect 224 -112 280 -68
rect 392 -112 448 -68
rect -448 -292 -392 -248
rect -280 -292 -224 -248
rect -112 -292 -56 -248
rect 56 -292 112 -248
rect 224 -292 280 -248
rect 392 -292 448 -248
<< pdiff >>
rect -540 293 -468 306
rect -540 247 -527 293
rect -481 292 -468 293
rect -372 293 -300 306
rect -372 292 -359 293
rect -481 248 -448 292
rect -392 248 -359 292
rect -481 247 -468 248
rect -540 234 -468 247
rect -372 247 -359 248
rect -313 292 -300 293
rect -204 293 -132 306
rect -204 292 -191 293
rect -313 248 -280 292
rect -224 248 -191 292
rect -313 247 -300 248
rect -372 234 -300 247
rect -204 247 -191 248
rect -145 292 -132 293
rect -36 293 36 306
rect -36 292 -23 293
rect -145 248 -112 292
rect -56 248 -23 292
rect -145 247 -132 248
rect -204 234 -132 247
rect -36 247 -23 248
rect 23 292 36 293
rect 132 293 204 306
rect 132 292 145 293
rect 23 248 56 292
rect 112 248 145 292
rect 23 247 36 248
rect -36 234 36 247
rect 132 247 145 248
rect 191 292 204 293
rect 300 293 372 306
rect 300 292 313 293
rect 191 248 224 292
rect 280 248 313 292
rect 191 247 204 248
rect 132 234 204 247
rect 300 247 313 248
rect 359 292 372 293
rect 468 293 540 306
rect 468 292 481 293
rect 359 248 392 292
rect 448 248 481 292
rect 359 247 372 248
rect 300 234 372 247
rect 468 247 481 248
rect 527 247 540 293
rect 468 234 540 247
rect -540 113 -468 126
rect -540 67 -527 113
rect -481 112 -468 113
rect -372 113 -300 126
rect -372 112 -359 113
rect -481 68 -448 112
rect -392 68 -359 112
rect -481 67 -468 68
rect -540 54 -468 67
rect -372 67 -359 68
rect -313 112 -300 113
rect -204 113 -132 126
rect -204 112 -191 113
rect -313 68 -280 112
rect -224 68 -191 112
rect -313 67 -300 68
rect -372 54 -300 67
rect -204 67 -191 68
rect -145 112 -132 113
rect -36 113 36 126
rect -36 112 -23 113
rect -145 68 -112 112
rect -56 68 -23 112
rect -145 67 -132 68
rect -204 54 -132 67
rect -36 67 -23 68
rect 23 112 36 113
rect 132 113 204 126
rect 132 112 145 113
rect 23 68 56 112
rect 112 68 145 112
rect 23 67 36 68
rect -36 54 36 67
rect 132 67 145 68
rect 191 112 204 113
rect 300 113 372 126
rect 300 112 313 113
rect 191 68 224 112
rect 280 68 313 112
rect 191 67 204 68
rect 132 54 204 67
rect 300 67 313 68
rect 359 112 372 113
rect 468 113 540 126
rect 468 112 481 113
rect 359 68 392 112
rect 448 68 481 112
rect 359 67 372 68
rect 300 54 372 67
rect 468 67 481 68
rect 527 67 540 113
rect 468 54 540 67
rect -540 -67 -468 -54
rect -540 -113 -527 -67
rect -481 -68 -468 -67
rect -372 -67 -300 -54
rect -372 -68 -359 -67
rect -481 -112 -448 -68
rect -392 -112 -359 -68
rect -481 -113 -468 -112
rect -540 -126 -468 -113
rect -372 -113 -359 -112
rect -313 -68 -300 -67
rect -204 -67 -132 -54
rect -204 -68 -191 -67
rect -313 -112 -280 -68
rect -224 -112 -191 -68
rect -313 -113 -300 -112
rect -372 -126 -300 -113
rect -204 -113 -191 -112
rect -145 -68 -132 -67
rect -36 -67 36 -54
rect -36 -68 -23 -67
rect -145 -112 -112 -68
rect -56 -112 -23 -68
rect -145 -113 -132 -112
rect -204 -126 -132 -113
rect -36 -113 -23 -112
rect 23 -68 36 -67
rect 132 -67 204 -54
rect 132 -68 145 -67
rect 23 -112 56 -68
rect 112 -112 145 -68
rect 23 -113 36 -112
rect -36 -126 36 -113
rect 132 -113 145 -112
rect 191 -68 204 -67
rect 300 -67 372 -54
rect 300 -68 313 -67
rect 191 -112 224 -68
rect 280 -112 313 -68
rect 191 -113 204 -112
rect 132 -126 204 -113
rect 300 -113 313 -112
rect 359 -68 372 -67
rect 468 -67 540 -54
rect 468 -68 481 -67
rect 359 -112 392 -68
rect 448 -112 481 -68
rect 359 -113 372 -112
rect 300 -126 372 -113
rect 468 -113 481 -112
rect 527 -113 540 -67
rect 468 -126 540 -113
rect -540 -247 -468 -234
rect -540 -293 -527 -247
rect -481 -248 -468 -247
rect -372 -247 -300 -234
rect -372 -248 -359 -247
rect -481 -292 -448 -248
rect -392 -292 -359 -248
rect -481 -293 -468 -292
rect -540 -306 -468 -293
rect -372 -293 -359 -292
rect -313 -248 -300 -247
rect -204 -247 -132 -234
rect -204 -248 -191 -247
rect -313 -292 -280 -248
rect -224 -292 -191 -248
rect -313 -293 -300 -292
rect -372 -306 -300 -293
rect -204 -293 -191 -292
rect -145 -248 -132 -247
rect -36 -247 36 -234
rect -36 -248 -23 -247
rect -145 -292 -112 -248
rect -56 -292 -23 -248
rect -145 -293 -132 -292
rect -204 -306 -132 -293
rect -36 -293 -23 -292
rect 23 -248 36 -247
rect 132 -247 204 -234
rect 132 -248 145 -247
rect 23 -292 56 -248
rect 112 -292 145 -248
rect 23 -293 36 -292
rect -36 -306 36 -293
rect 132 -293 145 -292
rect 191 -248 204 -247
rect 300 -247 372 -234
rect 300 -248 313 -247
rect 191 -292 224 -248
rect 280 -292 313 -248
rect 191 -293 204 -292
rect 132 -306 204 -293
rect 300 -293 313 -292
rect 359 -248 372 -247
rect 468 -247 540 -234
rect 468 -248 481 -247
rect 359 -292 392 -248
rect 448 -292 481 -248
rect 359 -293 372 -292
rect 300 -306 372 -293
rect 468 -293 481 -292
rect 527 -293 540 -247
rect 468 -306 540 -293
<< pdiffc >>
rect -527 247 -481 293
rect -359 247 -313 293
rect -191 247 -145 293
rect -23 247 23 293
rect 145 247 191 293
rect 313 247 359 293
rect 481 247 527 293
rect -527 67 -481 113
rect -359 67 -313 113
rect -191 67 -145 113
rect -23 67 23 113
rect 145 67 191 113
rect 313 67 359 113
rect 481 67 527 113
rect -527 -113 -481 -67
rect -359 -113 -313 -67
rect -191 -113 -145 -67
rect -23 -113 23 -67
rect 145 -113 191 -67
rect 313 -113 359 -67
rect 481 -113 527 -67
rect -527 -293 -481 -247
rect -359 -293 -313 -247
rect -191 -293 -145 -247
rect -23 -293 23 -247
rect 145 -293 191 -247
rect 313 -293 359 -247
rect 481 -293 527 -247
<< polysilicon >>
rect -448 292 -392 336
rect -448 204 -392 248
rect -280 292 -224 336
rect -280 204 -224 248
rect -112 292 -56 336
rect -112 204 -56 248
rect 56 292 112 336
rect 56 204 112 248
rect 224 292 280 336
rect 224 204 280 248
rect 392 292 448 336
rect 392 204 448 248
rect -448 112 -392 156
rect -448 24 -392 68
rect -280 112 -224 156
rect -280 24 -224 68
rect -112 112 -56 156
rect -112 24 -56 68
rect 56 112 112 156
rect 56 24 112 68
rect 224 112 280 156
rect 224 24 280 68
rect 392 112 448 156
rect 392 24 448 68
rect -448 -68 -392 -24
rect -448 -156 -392 -112
rect -280 -68 -224 -24
rect -280 -156 -224 -112
rect -112 -68 -56 -24
rect -112 -156 -56 -112
rect 56 -68 112 -24
rect 56 -156 112 -112
rect 224 -68 280 -24
rect 224 -156 280 -112
rect 392 -68 448 -24
rect 392 -156 448 -112
rect -448 -248 -392 -204
rect -448 -336 -392 -292
rect -280 -248 -224 -204
rect -280 -336 -224 -292
rect -112 -248 -56 -204
rect -112 -336 -56 -292
rect 56 -248 112 -204
rect 56 -336 112 -292
rect 224 -248 280 -204
rect 224 -336 280 -292
rect 392 -248 448 -204
rect 392 -336 448 -292
<< metal1 >>
rect -538 247 -527 293
rect -481 247 -470 293
rect -370 247 -359 293
rect -313 247 -302 293
rect -202 247 -191 293
rect -145 247 -134 293
rect -34 247 -23 293
rect 23 247 34 293
rect 134 247 145 293
rect 191 247 202 293
rect 302 247 313 293
rect 359 247 370 293
rect 470 247 481 293
rect 527 247 538 293
rect -538 67 -527 113
rect -481 67 -470 113
rect -370 67 -359 113
rect -313 67 -302 113
rect -202 67 -191 113
rect -145 67 -134 113
rect -34 67 -23 113
rect 23 67 34 113
rect 134 67 145 113
rect 191 67 202 113
rect 302 67 313 113
rect 359 67 370 113
rect 470 67 481 113
rect 527 67 538 113
rect -538 -113 -527 -67
rect -481 -113 -470 -67
rect -370 -113 -359 -67
rect -313 -113 -302 -67
rect -202 -113 -191 -67
rect -145 -113 -134 -67
rect -34 -113 -23 -67
rect 23 -113 34 -67
rect 134 -113 145 -67
rect 191 -113 202 -67
rect 302 -113 313 -67
rect 359 -113 370 -67
rect 470 -113 481 -67
rect 527 -113 538 -67
rect -538 -293 -527 -247
rect -481 -293 -470 -247
rect -370 -293 -359 -247
rect -313 -293 -302 -247
rect -202 -293 -191 -247
rect -145 -293 -134 -247
rect -34 -293 -23 -247
rect 23 -293 34 -247
rect 134 -293 145 -247
rect 191 -293 202 -247
rect 302 -293 313 -247
rect 359 -293 370 -247
rect 470 -293 481 -247
rect 527 -293 538 -247
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 0.22 l 0.280 m 4 nf 6 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
