magic
tech gf180mcuC
magscale 1 10
timestamp 1691396512
<< pwell >>
rect -460 -940 460 940
<< nmos >>
rect -348 632 -292 872
rect -188 632 -132 872
rect -28 632 28 872
rect 132 632 188 872
rect 292 632 348 872
rect -348 256 -292 496
rect -188 256 -132 496
rect -28 256 28 496
rect 132 256 188 496
rect 292 256 348 496
rect -348 -120 -292 120
rect -188 -120 -132 120
rect -28 -120 28 120
rect 132 -120 188 120
rect 292 -120 348 120
rect -348 -496 -292 -256
rect -188 -496 -132 -256
rect -28 -496 28 -256
rect 132 -496 188 -256
rect 292 -496 348 -256
rect -348 -872 -292 -632
rect -188 -872 -132 -632
rect -28 -872 28 -632
rect 132 -872 188 -632
rect 292 -872 348 -632
<< ndiff >>
rect -436 859 -348 872
rect -436 645 -423 859
rect -377 645 -348 859
rect -436 632 -348 645
rect -292 859 -188 872
rect -292 645 -263 859
rect -217 645 -188 859
rect -292 632 -188 645
rect -132 859 -28 872
rect -132 645 -103 859
rect -57 645 -28 859
rect -132 632 -28 645
rect 28 859 132 872
rect 28 645 57 859
rect 103 645 132 859
rect 28 632 132 645
rect 188 859 292 872
rect 188 645 217 859
rect 263 645 292 859
rect 188 632 292 645
rect 348 859 436 872
rect 348 645 377 859
rect 423 645 436 859
rect 348 632 436 645
rect -436 483 -348 496
rect -436 269 -423 483
rect -377 269 -348 483
rect -436 256 -348 269
rect -292 483 -188 496
rect -292 269 -263 483
rect -217 269 -188 483
rect -292 256 -188 269
rect -132 483 -28 496
rect -132 269 -103 483
rect -57 269 -28 483
rect -132 256 -28 269
rect 28 483 132 496
rect 28 269 57 483
rect 103 269 132 483
rect 28 256 132 269
rect 188 483 292 496
rect 188 269 217 483
rect 263 269 292 483
rect 188 256 292 269
rect 348 483 436 496
rect 348 269 377 483
rect 423 269 436 483
rect 348 256 436 269
rect -436 107 -348 120
rect -436 -107 -423 107
rect -377 -107 -348 107
rect -436 -120 -348 -107
rect -292 107 -188 120
rect -292 -107 -263 107
rect -217 -107 -188 107
rect -292 -120 -188 -107
rect -132 107 -28 120
rect -132 -107 -103 107
rect -57 -107 -28 107
rect -132 -120 -28 -107
rect 28 107 132 120
rect 28 -107 57 107
rect 103 -107 132 107
rect 28 -120 132 -107
rect 188 107 292 120
rect 188 -107 217 107
rect 263 -107 292 107
rect 188 -120 292 -107
rect 348 107 436 120
rect 348 -107 377 107
rect 423 -107 436 107
rect 348 -120 436 -107
rect -436 -269 -348 -256
rect -436 -483 -423 -269
rect -377 -483 -348 -269
rect -436 -496 -348 -483
rect -292 -269 -188 -256
rect -292 -483 -263 -269
rect -217 -483 -188 -269
rect -292 -496 -188 -483
rect -132 -269 -28 -256
rect -132 -483 -103 -269
rect -57 -483 -28 -269
rect -132 -496 -28 -483
rect 28 -269 132 -256
rect 28 -483 57 -269
rect 103 -483 132 -269
rect 28 -496 132 -483
rect 188 -269 292 -256
rect 188 -483 217 -269
rect 263 -483 292 -269
rect 188 -496 292 -483
rect 348 -269 436 -256
rect 348 -483 377 -269
rect 423 -483 436 -269
rect 348 -496 436 -483
rect -436 -645 -348 -632
rect -436 -859 -423 -645
rect -377 -859 -348 -645
rect -436 -872 -348 -859
rect -292 -645 -188 -632
rect -292 -859 -263 -645
rect -217 -859 -188 -645
rect -292 -872 -188 -859
rect -132 -645 -28 -632
rect -132 -859 -103 -645
rect -57 -859 -28 -645
rect -132 -872 -28 -859
rect 28 -645 132 -632
rect 28 -859 57 -645
rect 103 -859 132 -645
rect 28 -872 132 -859
rect 188 -645 292 -632
rect 188 -859 217 -645
rect 263 -859 292 -645
rect 188 -872 292 -859
rect 348 -645 436 -632
rect 348 -859 377 -645
rect 423 -859 436 -645
rect 348 -872 436 -859
<< ndiffc >>
rect -423 645 -377 859
rect -263 645 -217 859
rect -103 645 -57 859
rect 57 645 103 859
rect 217 645 263 859
rect 377 645 423 859
rect -423 269 -377 483
rect -263 269 -217 483
rect -103 269 -57 483
rect 57 269 103 483
rect 217 269 263 483
rect 377 269 423 483
rect -423 -107 -377 107
rect -263 -107 -217 107
rect -103 -107 -57 107
rect 57 -107 103 107
rect 217 -107 263 107
rect 377 -107 423 107
rect -423 -483 -377 -269
rect -263 -483 -217 -269
rect -103 -483 -57 -269
rect 57 -483 103 -269
rect 217 -483 263 -269
rect 377 -483 423 -269
rect -423 -859 -377 -645
rect -263 -859 -217 -645
rect -103 -859 -57 -645
rect 57 -859 103 -645
rect 217 -859 263 -645
rect 377 -859 423 -645
<< polysilicon >>
rect -348 872 -292 916
rect -188 872 -132 916
rect -28 872 28 916
rect 132 872 188 916
rect 292 872 348 916
rect -348 588 -292 632
rect -188 588 -132 632
rect -28 588 28 632
rect 132 588 188 632
rect 292 588 348 632
rect -348 496 -292 540
rect -188 496 -132 540
rect -28 496 28 540
rect 132 496 188 540
rect 292 496 348 540
rect -348 212 -292 256
rect -188 212 -132 256
rect -28 212 28 256
rect 132 212 188 256
rect 292 212 348 256
rect -348 120 -292 164
rect -188 120 -132 164
rect -28 120 28 164
rect 132 120 188 164
rect 292 120 348 164
rect -348 -164 -292 -120
rect -188 -164 -132 -120
rect -28 -164 28 -120
rect 132 -164 188 -120
rect 292 -164 348 -120
rect -348 -256 -292 -212
rect -188 -256 -132 -212
rect -28 -256 28 -212
rect 132 -256 188 -212
rect 292 -256 348 -212
rect -348 -540 -292 -496
rect -188 -540 -132 -496
rect -28 -540 28 -496
rect 132 -540 188 -496
rect 292 -540 348 -496
rect -348 -632 -292 -588
rect -188 -632 -132 -588
rect -28 -632 28 -588
rect 132 -632 188 -588
rect 292 -632 348 -588
rect -348 -916 -292 -872
rect -188 -916 -132 -872
rect -28 -916 28 -872
rect 132 -916 188 -872
rect 292 -916 348 -872
<< metal1 >>
rect -423 859 -377 870
rect -423 634 -377 645
rect -263 859 -217 870
rect -263 634 -217 645
rect -103 859 -57 870
rect -103 634 -57 645
rect 57 859 103 870
rect 57 634 103 645
rect 217 859 263 870
rect 217 634 263 645
rect 377 859 423 870
rect 377 634 423 645
rect -423 483 -377 494
rect -423 258 -377 269
rect -263 483 -217 494
rect -263 258 -217 269
rect -103 483 -57 494
rect -103 258 -57 269
rect 57 483 103 494
rect 57 258 103 269
rect 217 483 263 494
rect 217 258 263 269
rect 377 483 423 494
rect 377 258 423 269
rect -423 107 -377 118
rect -423 -118 -377 -107
rect -263 107 -217 118
rect -263 -118 -217 -107
rect -103 107 -57 118
rect -103 -118 -57 -107
rect 57 107 103 118
rect 57 -118 103 -107
rect 217 107 263 118
rect 217 -118 263 -107
rect 377 107 423 118
rect 377 -118 423 -107
rect -423 -269 -377 -258
rect -423 -494 -377 -483
rect -263 -269 -217 -258
rect -263 -494 -217 -483
rect -103 -269 -57 -258
rect -103 -494 -57 -483
rect 57 -269 103 -258
rect 57 -494 103 -483
rect 217 -269 263 -258
rect 217 -494 263 -483
rect 377 -269 423 -258
rect 377 -494 423 -483
rect -423 -645 -377 -634
rect -423 -870 -377 -859
rect -263 -645 -217 -634
rect -263 -870 -217 -859
rect -103 -645 -57 -634
rect -103 -870 -57 -859
rect 57 -645 103 -634
rect 57 -870 103 -859
rect 217 -645 263 -634
rect 217 -870 263 -859
rect 377 -645 423 -634
rect 377 -870 423 -859
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 1.2 l 0.280 m 5 nf 5 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
