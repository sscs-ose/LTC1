* NGSPICE file created from Tappered_Buffer_flat.ext - technology: gf180mcuC

.subckt Tappered_Buffer_flat VDD IN OUT VSS
X0 VDD a_138_n2984.t24 OUT.t76 VDD.t64 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1 OUT a_138_n2984.t25 VDD.t125 VDD.t27 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X2 VDD a_138_n2984.t26 OUT.t75 VDD.t2 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X3 VSS.t50 VSS.t48 VSS.t50 VSS.t49 nfet_03v3 ad=0 pd=0 as=0.728p ps=3.32u w=2.8u l=0.5u
X4 OUT a_138_n2984.t27 VSS.t112 VSS.t106 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X5 OUT a_138_n2984.t28 VDD.t122 VDD.t0 pfet_03v3 ad=0.728p pd=3.32u as=1.23p ps=6.48u w=2.8u l=0.5u
X6 OUT a_138_n2984.t29 VDD.t121 VDD.t50 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X7 VSS.t47 VSS.t45 VSS.t47 VSS.t46 nfet_03v3 ad=0 pd=0 as=0.728p ps=3.32u w=2.8u l=0.5u
X8 VDD a_138_n2984.t30 OUT.t74 VDD.t16 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X9 VSS a_138_n2984.t31 OUT.t33 VSS.t34 nfet_03v3 ad=1.23p pd=6.48u as=0.728p ps=3.32u w=2.8u l=0.5u
X10 VDD a_138_n2984.t32 OUT.t73 VDD.t88 pfet_03v3 ad=1.23p pd=6.48u as=0.728p ps=3.32u w=2.8u l=0.5u
X11 OUT a_138_n2984.t33 VDD.t116 VDD.t45 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X12 VDD a_138_n2984.t34 OUT.t72 VDD.t16 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X13 VSS a_138_n2984.t35 OUT.t32 VSS.t31 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X14 VDD a_138_n2984.t36 OUT.t71 VDD.t55 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X15 VDD a_138_n2984.t37 OUT.t70 VDD.t83 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X16 VDD a_138_n2984.t38 OUT.t69 VDD.t77 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X17 VDD a_138_n2984.t39 OUT.t68 VDD.t19 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X18 VSS.t44 VSS.t42 VSS.t44 VSS.t43 nfet_03v3 ad=0 pd=0 as=0.728p ps=3.32u w=2.8u l=0.5u
X19 VSS.t41 VSS.t39 VSS.t41 VSS.t40 nfet_03v3 ad=0 pd=0 as=0.728p ps=3.32u w=2.8u l=0.5u
X20 VDD a_138_n2984.t40 OUT.t67 VDD.t24 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X21 VSS.t38 VSS.t36 VSS.t38 VSS.t37 nfet_03v3 ad=0 pd=0 as=0.728p ps=3.32u w=2.8u l=0.5u
X22 OUT a_138_n2984.t41 VDD.t103 VDD.t47 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X23 VDD a_138_n2984.t42 OUT.t66 VDD.t10 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X24 VDD a_240_n2164.t8 a_138_n2984.t3 VDD.t2 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X25 OUT a_138_n2984.t43 VSS.t107 VSS.t106 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X26 VDD a_138_n2984.t44 OUT.t65 VDD.t77 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X27 VDD a_138_n2984.t45 OUT.t64 VDD.t88 pfet_03v3 ad=1.23p pd=6.48u as=0.728p ps=3.32u w=2.8u l=0.5u
X28 VDD a_138_n2984.t46 OUT.t63 VDD.t24 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X29 VDD a_138_n2984.t47 OUT.t62 VDD.t37 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X30 VDD a_138_n2984.t48 OUT.t61 VDD.t61 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X31 VDD a_138_n2984.t49 OUT.t60 VDD.t88 pfet_03v3 ad=1.23p pd=6.48u as=0.728p ps=3.32u w=2.8u l=0.5u
X32 VDD a_240_n2164.t9 a_138_n2984.t10 VDD.t19 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X33 OUT a_138_n2984.t50 VSS.t105 VSS.t28 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X34 VSS.t35 VSS.t33 VSS.t35 VSS.t34 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.5u
X35 OUT a_138_n2984.t51 VSS.t104 VSS.t96 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X36 OUT a_138_n2984.t52 VDD.t87 VDD.t5 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X37 OUT a_138_n2984.t53 VDD.t86 VDD.t52 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X38 VSS.t32 VSS.t30 VSS.t32 VSS.t31 nfet_03v3 ad=0 pd=0 as=0.728p ps=3.32u w=2.8u l=0.5u
X39 OUT a_138_n2984.t54 VSS.t103 VSS.t102 nfet_03v3 ad=0.728p pd=3.32u as=1.23p ps=6.48u w=2.8u l=0.5u
X40 OUT a_138_n2984.t55 VSS.t101 VSS.t100 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X41 OUT a_138_n2984.t56 VSS.t99 VSS.t7 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X42 VDD IN.t2 a_240_n2164.t4 VDD.t64 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X43 OUT a_138_n2984.t57 VSS.t98 VSS.t25 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X44 VDD a_138_n2984.t58 OUT.t59 VDD.t83 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X45 OUT a_138_n2984.t59 VDD.t82 VDD.t67 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X46 OUT a_138_n2984.t60 VDD.t81 VDD.t5 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X47 OUT a_138_n2984.t61 VDD.t80 VDD.t0 pfet_03v3 ad=0.728p pd=3.32u as=1.23p ps=6.48u w=2.8u l=0.5u
X48 VDD a_138_n2984.t62 OUT.t58 VDD.t77 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X49 OUT a_138_n2984.t63 VDD.t76 VDD.t72 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X50 VDD a_240_n2164.t14 a_138_n2984.t7 VDD.t61 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X51 VSS.t29 VSS.t27 VSS.t29 VSS.t28 nfet_03v3 ad=0 pd=0 as=0.728p ps=3.32u w=2.8u l=0.5u
X52 OUT a_138_n2984.t64 VSS.t97 VSS.t96 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X53 OUT a_138_n2984.t65 VDD.t75 VDD.t42 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X54 OUT a_138_n2984.t66 VSS.t95 VSS.t22 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X55 OUT a_138_n2984.t67 VDD.t74 VDD.t47 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X56 OUT a_138_n2984.t68 VDD.t73 VDD.t72 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X57 OUT a_138_n2984.t69 VSS.t94 VSS.t19 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X58 OUT a_138_n2984.t70 VSS.t93 VSS.t16 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X59 OUT a_138_n2984.t71 VDD.t71 VDD.t22 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X60 OUT a_138_n2984.t72 VSS.t92 VSS.t13 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X61 OUT a_138_n2984.t73 VDD.t70 VDD.t22 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X62 OUT a_138_n2984.t74 VDD.t69 VDD.t29 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X63 OUT a_138_n2984.t75 VDD.t68 VDD.t67 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X64 VDD a_138_n2984.t76 OUT.t57 VDD.t64 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X65 VDD IN.t4 a_240_n2164.t2 VDD.t7 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X66 VDD a_138_n2984.t77 OUT.t56 VDD.t61 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X67 VSS.t26 VSS.t24 VSS.t26 VSS.t25 nfet_03v3 ad=0 pd=0 as=0.728p ps=3.32u w=2.8u l=0.5u
X68 OUT a_138_n2984.t78 VSS.t91 VSS.t3 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X69 VSS a_240_n2164.t17 a_138_n2984.t18 VSS.t82 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X70 OUT a_138_n2984.t79 VSS.t90 VSS.t5 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X71 VDD a_138_n2984.t80 OUT.t55 VDD.t2 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X72 VDD a_240_n2164.t18 a_138_n2984.t19 VDD.t83 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X73 OUT a_138_n2984.t81 VSS.t89 VSS.t10 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X74 OUT a_138_n2984.t82 VDD.t58 VDD.t27 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X75 VDD a_138_n2984.t83 OUT.t54 VDD.t55 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X76 OUT a_138_n2984.t84 VDD.t54 VDD.t33 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X77 OUT a_138_n2984.t85 VDD.t53 VDD.t52 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X78 OUT a_138_n2984.t86 VDD.t51 VDD.t50 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X79 VDD a_240_n2164.t20 a_138_n2984.t17 VDD.t37 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X80 VSS a_138_n2984.t87 OUT.t31 VSS.t79 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X81 VSS.t23 VSS.t21 VSS.t23 VSS.t22 nfet_03v3 ad=0 pd=0 as=0.728p ps=3.32u w=2.8u l=0.5u
X82 VSS a_138_n2984.t88 OUT.t30 VSS.t76 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X83 VSS.t20 VSS.t18 VSS.t20 VSS.t19 nfet_03v3 ad=0 pd=0 as=0.728p ps=3.32u w=2.8u l=0.5u
X84 VSS.t17 VSS.t15 VSS.t17 VSS.t16 nfet_03v3 ad=0 pd=0 as=0.728p ps=3.32u w=2.8u l=0.5u
X85 VSS.t14 VSS.t12 VSS.t14 VSS.t13 nfet_03v3 ad=0 pd=0 as=0.728p ps=3.32u w=2.8u l=0.5u
X86 OUT a_138_n2984.t89 VDD.t49 VDD.t33 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X87 VDD a_240_n2164.t22 a_138_n2984.t13 VDD.t10 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X88 VSS a_138_n2984.t90 OUT.t29 VSS.t82 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X89 OUT a_138_n2984.t91 VDD.t48 VDD.t47 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X90 OUT a_138_n2984.t92 VDD.t46 VDD.t45 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X91 VSS a_240_n2164.t23 a_138_n2984.t8 VSS.t69 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X92 OUT a_138_n2984.t93 VDD.t44 VDD.t31 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X93 VSS IN.t5 a_240_n2164.t0 VSS.t0 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X94 OUT a_138_n2984.t94 VDD.t43 VDD.t42 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X95 VDD a_240_n2164.t24 a_138_n2984.t9 VDD.t55 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X96 VDD a_138_n2984.t95 OUT.t53 VDD.t7 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X97 VDD a_138_n2984.t96 OUT.t52 VDD.t37 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X98 VSS a_240_n2164.t25 a_138_n2984.t4 VSS.t51 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X99 VSS.t11 VSS.t9 VSS.t11 VSS.t10 nfet_03v3 ad=0 pd=0 as=0.728p ps=3.32u w=2.8u l=0.5u
X100 VSS a_240_n2164.t26 a_138_n2984.t5 VSS.t54 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X101 VDD a_138_n2984.t97 OUT.t51 VDD.t13 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X102 VDD a_240_n2164.t27 a_138_n2984.t22 VDD.t13 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X103 OUT a_138_n2984.t98 VDD.t34 VDD.t33 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X104 VSS a_138_n2984.t99 OUT.t28 VSS.t79 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X105 VSS a_138_n2984.t100 OUT.t27 VSS.t76 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X106 VSS a_138_n2984.t101 OUT.t26 VSS.t49 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X107 OUT a_138_n2984.t102 VDD.t32 VDD.t31 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X108 VSS a_138_n2984.t103 OUT.t25 VSS.t46 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X109 OUT a_138_n2984.t104 VDD.t30 VDD.t29 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X110 OUT a_138_n2984.t105 VDD.t28 VDD.t27 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X111 VDD a_138_n2984.t106 OUT.t50 VDD.t24 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X112 VSS a_138_n2984.t107 OUT.t24 VSS.t69 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X113 VSS a_138_n2984.t108 OUT.t23 VSS.t0 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X114 OUT a_138_n2984.t109 VDD.t23 VDD.t22 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X115 VSS a_138_n2984.t110 OUT.t22 VSS.t51 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X116 VSS a_138_n2984.t111 OUT.t21 VSS.t54 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X117 VSS a_138_n2984.t112 OUT.t20 VSS.t43 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X118 VDD a_138_n2984.t113 OUT.t49 VDD.t19 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X119 VSS a_138_n2984.t114 OUT.t19 VSS.t40 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X120 VDD a_138_n2984.t115 OUT.t48 VDD.t16 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X121 VDD a_138_n2984.t116 OUT.t47 VDD.t13 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X122 VSS a_138_n2984.t117 OUT.t18 VSS.t37 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X123 VDD a_138_n2984.t118 OUT.t46 VDD.t10 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X124 VDD a_138_n2984.t119 OUT.t45 VDD.t7 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
R0 a_138_n2984.n75 a_138_n2984.t31 40.255
R1 a_138_n2984.n34 a_138_n2984.t54 37.7641
R2 a_138_n2984.t85 a_138_n2984.n32 30.4352
R3 a_138_n2984.t47 a_138_n2984.n50 28.4705
R4 a_138_n2984.t93 a_138_n2984.n57 28.4705
R5 a_138_n2984.t118 a_138_n2984.n64 28.4705
R6 a_138_n2984.t82 a_138_n2984.n71 28.4705
R7 a_138_n2984.t34 a_138_n2984.n79 28.4705
R8 a_138_n2984.n83 a_138_n2984.t45 27.3249
R9 a_138_n2984.n50 a_138_n2984.t87 27.1982
R10 a_138_n2984.t45 a_138_n2984.n82 25.4384
R11 a_138_n2984.n82 a_138_n2984.t32 25.4384
R12 a_138_n2984.n80 a_138_n2984.t115 25.4045
R13 a_138_n2984.n74 a_138_n2984.t73 25.4045
R14 a_138_n2984.n74 a_138_n2984.t71 25.4045
R15 a_138_n2984.n73 a_138_n2984.t62 25.4045
R16 a_138_n2984.n73 a_138_n2984.t44 25.4045
R17 a_138_n2984.n65 a_138_n2984.t42 25.4045
R18 a_138_n2984.n60 a_138_n2984.t33 25.4045
R19 a_138_n2984.n60 a_138_n2984.t92 25.4045
R20 a_138_n2984.n59 a_138_n2984.t83 25.4045
R21 a_138_n2984.n59 a_138_n2984.t36 25.4045
R22 a_138_n2984.n10 a_138_n2984.t28 25.4045
R23 a_138_n2984.n10 a_138_n2984.t61 25.4045
R24 a_138_n2984.n11 a_138_n2984.t76 25.4045
R25 a_138_n2984.n11 a_138_n2984.t24 25.4045
R26 a_138_n2984.n12 a_138_n2984.t52 25.4045
R27 a_138_n2984.n12 a_138_n2984.t60 25.4045
R28 a_138_n2984.n13 a_138_n2984.t95 25.4045
R29 a_138_n2984.n13 a_138_n2984.t119 25.4045
R30 a_138_n2984.n14 a_138_n2984.t75 25.4045
R31 a_138_n2984.n14 a_138_n2984.t59 25.4045
R32 a_138_n2984.n15 a_138_n2984.t116 25.4045
R33 a_138_n2984.n15 a_138_n2984.t97 25.4045
R34 a_138_n2984.n16 a_138_n2984.t68 25.4045
R35 a_138_n2984.n16 a_138_n2984.t63 25.4045
R36 a_138_n2984.n17 a_138_n2984.t113 25.4045
R37 a_138_n2984.n17 a_138_n2984.t39 25.4045
R38 a_138_n2984.n18 a_138_n2984.t65 25.4045
R39 a_138_n2984.n18 a_138_n2984.t94 25.4045
R40 a_138_n2984.n19 a_138_n2984.t80 25.4045
R41 a_138_n2984.n19 a_138_n2984.t26 25.4045
R42 a_138_n2984.n20 a_138_n2984.t29 25.4045
R43 a_138_n2984.n20 a_138_n2984.t86 25.4045
R44 a_138_n2984.n21 a_138_n2984.t77 25.4045
R45 a_138_n2984.n21 a_138_n2984.t48 25.4045
R46 a_138_n2984.n33 a_138_n2984.t53 25.4045
R47 a_138_n2984.n33 a_138_n2984.t85 25.4045
R48 a_138_n2984.n51 a_138_n2984.t96 25.4045
R49 a_138_n2984.n46 a_138_n2984.t88 25.4045
R50 a_138_n2984.n44 a_138_n2984.t27 25.4045
R51 a_138_n2984.n44 a_138_n2984.t43 25.4045
R52 a_138_n2984.n46 a_138_n2984.t100 25.4045
R53 a_138_n2984.n48 a_138_n2984.t51 25.4045
R54 a_138_n2984.n48 a_138_n2984.t64 25.4045
R55 a_138_n2984.n49 a_138_n2984.t99 25.4045
R56 a_138_n2984.t87 a_138_n2984.n49 25.4045
R57 a_138_n2984.n51 a_138_n2984.t47 25.4045
R58 a_138_n2984.n52 a_138_n2984.t104 25.4045
R59 a_138_n2984.n52 a_138_n2984.t74 25.4045
R60 a_138_n2984.n53 a_138_n2984.t58 25.4045
R61 a_138_n2984.n53 a_138_n2984.t37 25.4045
R62 a_138_n2984.n58 a_138_n2984.t102 25.4045
R63 a_138_n2984.n58 a_138_n2984.t93 25.4045
R64 a_138_n2984.n65 a_138_n2984.t118 25.4045
R65 a_138_n2984.n66 a_138_n2984.t89 25.4045
R66 a_138_n2984.n66 a_138_n2984.t84 25.4045
R67 a_138_n2984.n67 a_138_n2984.t40 25.4045
R68 a_138_n2984.n67 a_138_n2984.t46 25.4045
R69 a_138_n2984.n72 a_138_n2984.t105 25.4045
R70 a_138_n2984.n72 a_138_n2984.t82 25.4045
R71 a_138_n2984.n80 a_138_n2984.t34 25.4045
R72 a_138_n2984.n81 a_138_n2984.t67 25.4045
R73 a_138_n2984.n81 a_138_n2984.t91 25.4045
R74 a_138_n2984.n56 a_138_n2984.t72 23.6525
R75 a_138_n2984.n63 a_138_n2984.t117 23.6525
R76 a_138_n2984.n70 a_138_n2984.t81 23.6525
R77 a_138_n2984.n78 a_138_n2984.t101 23.6525
R78 a_138_n2984.n83 a_138_n2984.t49 23.5689
R79 a_138_n2984.n84 a_138_n2984.t41 23.5065
R80 a_138_n2984.n85 a_138_n2984.t30 23.5065
R81 a_138_n2984.n86 a_138_n2984.t109 23.5065
R82 a_138_n2984.n87 a_138_n2984.t38 23.5065
R83 a_138_n2984.n88 a_138_n2984.t25 23.5065
R84 a_138_n2984.n89 a_138_n2984.t106 23.5065
R85 a_138_n2984.n90 a_138_n2984.t98 23.5065
R86 a_138_n2984.n35 a_138_n2984.t79 22.4115
R87 a_138_n2984.n34 a_138_n2984.t108 22.4115
R88 a_138_n2984.n55 a_138_n2984.t103 20.4405
R89 a_138_n2984.n54 a_138_n2984.t50 20.4405
R90 a_138_n2984.n36 a_138_n2984.t107 20.4405
R91 a_138_n2984.n37 a_138_n2984.t78 20.4405
R92 a_138_n2984.n38 a_138_n2984.t90 20.4405
R93 a_138_n2984.n39 a_138_n2984.t56 20.4405
R94 a_138_n2984.n40 a_138_n2984.t111 20.4405
R95 a_138_n2984.n41 a_138_n2984.t55 20.4405
R96 a_138_n2984.n42 a_138_n2984.t110 20.4405
R97 a_138_n2984.t43 a_138_n2984.n43 20.4405
R98 a_138_n2984.t100 a_138_n2984.n45 20.4405
R99 a_138_n2984.t64 a_138_n2984.n47 20.4405
R100 a_138_n2984.n61 a_138_n2984.t35 20.4405
R101 a_138_n2984.n62 a_138_n2984.t70 20.4405
R102 a_138_n2984.n69 a_138_n2984.t114 20.4405
R103 a_138_n2984.n68 a_138_n2984.t57 20.4405
R104 a_138_n2984.n76 a_138_n2984.t112 20.4405
R105 a_138_n2984.n77 a_138_n2984.t69 20.4405
R106 a_138_n2984.n75 a_138_n2984.t66 20.4405
R107 a_138_n2984.n56 a_138_n2984.n55 19.2623
R108 a_138_n2984.n63 a_138_n2984.n62 19.2623
R109 a_138_n2984.n70 a_138_n2984.n69 19.2623
R110 a_138_n2984.n78 a_138_n2984.n77 19.2623
R111 a_138_n2984.n55 a_138_n2984.n54 17.2497
R112 a_138_n2984.n62 a_138_n2984.n61 17.2497
R113 a_138_n2984.n69 a_138_n2984.n68 17.2497
R114 a_138_n2984.n77 a_138_n2984.n76 17.2497
R115 a_138_n2984.n80 a_138_n2984.n74 15.8172
R116 a_138_n2984.n74 a_138_n2984.n73 15.8172
R117 a_138_n2984.n65 a_138_n2984.n60 15.8172
R118 a_138_n2984.n60 a_138_n2984.n59 15.8172
R119 a_138_n2984.n12 a_138_n2984.n11 15.8172
R120 a_138_n2984.n13 a_138_n2984.n12 15.8172
R121 a_138_n2984.n14 a_138_n2984.n13 15.8172
R122 a_138_n2984.n15 a_138_n2984.n14 15.8172
R123 a_138_n2984.n16 a_138_n2984.n15 15.8172
R124 a_138_n2984.n17 a_138_n2984.n16 15.8172
R125 a_138_n2984.n18 a_138_n2984.n17 15.8172
R126 a_138_n2984.n19 a_138_n2984.n18 15.8172
R127 a_138_n2984.n20 a_138_n2984.n19 15.8172
R128 a_138_n2984.n21 a_138_n2984.n20 15.8172
R129 a_138_n2984.n33 a_138_n2984.n21 15.8172
R130 a_138_n2984.n51 a_138_n2984.n33 15.8172
R131 a_138_n2984.n52 a_138_n2984.n51 15.8172
R132 a_138_n2984.n53 a_138_n2984.n52 15.8172
R133 a_138_n2984.n58 a_138_n2984.n53 15.8172
R134 a_138_n2984.n59 a_138_n2984.n58 15.8172
R135 a_138_n2984.n66 a_138_n2984.n65 15.8172
R136 a_138_n2984.n67 a_138_n2984.n66 15.8172
R137 a_138_n2984.n72 a_138_n2984.n67 15.8172
R138 a_138_n2984.n73 a_138_n2984.n72 15.8172
R139 a_138_n2984.n81 a_138_n2984.n80 15.8172
R140 a_138_n2984.n82 a_138_n2984.n81 15.8172
R141 a_138_n2984.n79 a_138_n2984.n75 15.7165
R142 a_138_n2984.n11 a_138_n2984.n10 15.4944
R143 a_138_n2984.n35 a_138_n2984.n34 15.3531
R144 a_138_n2984.n36 a_138_n2984.n35 15.2373
R145 a_138_n2984.n37 a_138_n2984.n36 14.4179
R146 a_138_n2984.n38 a_138_n2984.n37 14.4179
R147 a_138_n2984.n39 a_138_n2984.n38 14.4179
R148 a_138_n2984.n40 a_138_n2984.n39 14.4179
R149 a_138_n2984.n41 a_138_n2984.n40 14.4179
R150 a_138_n2984.n42 a_138_n2984.n41 14.4179
R151 a_138_n2984.n43 a_138_n2984.n42 14.3002
R152 a_138_n2984.n46 a_138_n2984.n44 13.3198
R153 a_138_n2984.n48 a_138_n2984.n46 13.3198
R154 a_138_n2984.n49 a_138_n2984.n48 13.3198
R155 a_138_n2984.n85 a_138_n2984.n84 12.7287
R156 a_138_n2984.n86 a_138_n2984.n85 12.7287
R157 a_138_n2984.n87 a_138_n2984.n86 12.7287
R158 a_138_n2984.n88 a_138_n2984.n87 12.7287
R159 a_138_n2984.n89 a_138_n2984.n88 12.7287
R160 a_138_n2984.n90 a_138_n2984.n89 12.7287
R161 a_138_n2984.n84 a_138_n2984.n83 12.6663
R162 a_138_n2984.n91 a_138_n2984.n90 4.60781
R163 a_138_n2984.n100 a_138_n2984.n99 3.69699
R164 a_138_n2984.n57 a_138_n2984.n56 3.54621
R165 a_138_n2984.n64 a_138_n2984.n63 3.54621
R166 a_138_n2984.n71 a_138_n2984.n70 3.54621
R167 a_138_n2984.n79 a_138_n2984.n78 3.54621
R168 a_138_n2984.n92 a_138_n2984.n7 3.23924
R169 a_138_n2984.n93 a_138_n2984.n5 3.23924
R170 a_138_n2984.n94 a_138_n2984.n3 3.23924
R171 a_138_n2984.n91 a_138_n2984.n9 3.2392
R172 a_138_n2984.n100 a_138_n2984.n97 3.2392
R173 a_138_n2984.n95 a_138_n2984.n1 3.23916
R174 a_138_n2984.n103 a_138_n2984.n101 3.23916
R175 a_138_n2984.n26 a_138_n2984.n23 2.91928
R176 a_138_n2984.n32 a_138_n2984.n31 2.58908
R177 a_138_n2984.n29 a_138_n2984.n28 2.58711
R178 a_138_n2984.n26 a_138_n2984.n25 2.58292
R179 a_138_n2984.n9 a_138_n2984.t13 0.6505
R180 a_138_n2984.n9 a_138_n2984.n8 0.6505
R181 a_138_n2984.n7 a_138_n2984.t9 0.6505
R182 a_138_n2984.n7 a_138_n2984.n6 0.6505
R183 a_138_n2984.n5 a_138_n2984.t19 0.6505
R184 a_138_n2984.n5 a_138_n2984.n4 0.6505
R185 a_138_n2984.n3 a_138_n2984.t17 0.6505
R186 a_138_n2984.n3 a_138_n2984.n2 0.6505
R187 a_138_n2984.n1 a_138_n2984.t7 0.6505
R188 a_138_n2984.n1 a_138_n2984.n0 0.6505
R189 a_138_n2984.n97 a_138_n2984.t10 0.6505
R190 a_138_n2984.n97 a_138_n2984.n96 0.6505
R191 a_138_n2984.n99 a_138_n2984.t22 0.6505
R192 a_138_n2984.n99 a_138_n2984.n98 0.6505
R193 a_138_n2984.t3 a_138_n2984.n103 0.6505
R194 a_138_n2984.n103 a_138_n2984.n102 0.6505
R195 a_138_n2984.n31 a_138_n2984.t4 0.5855
R196 a_138_n2984.n31 a_138_n2984.n30 0.5855
R197 a_138_n2984.n23 a_138_n2984.t8 0.5855
R198 a_138_n2984.n23 a_138_n2984.n22 0.5855
R199 a_138_n2984.n25 a_138_n2984.t18 0.5855
R200 a_138_n2984.n25 a_138_n2984.n24 0.5855
R201 a_138_n2984.n28 a_138_n2984.t5 0.5855
R202 a_138_n2984.n28 a_138_n2984.n27 0.5855
R203 a_138_n2984.n101 a_138_n2984.n95 0.466449
R204 a_138_n2984.n92 a_138_n2984.n91 0.46531
R205 a_138_n2984.n93 a_138_n2984.n92 0.46531
R206 a_138_n2984.n94 a_138_n2984.n93 0.46531
R207 a_138_n2984.n101 a_138_n2984.n100 0.46531
R208 a_138_n2984.n95 a_138_n2984.n94 0.464171
R209 a_138_n2984.n29 a_138_n2984.n26 0.341015
R210 a_138_n2984.n32 a_138_n2984.n29 0.337297
R211 OUT.n8 OUT.n7 3.74358
R212 OUT.n10 OUT.n1 3.24303
R213 OUT.n9 OUT.n3 3.24286
R214 OUT.n8 OUT.n5 3.24211
R215 OUT.n84 OUT.n21 3.23441
R216 OUT.n81 OUT.n27 3.23441
R217 OUT.n76 OUT.n39 3.23441
R218 OUT.n69 OUT.n55 3.23441
R219 OUT.n68 OUT.n59 3.23441
R220 OUT.n81 OUT.n29 3.23391
R221 OUT.n83 OUT.n23 3.23391
R222 OUT.n76 OUT.n41 3.23387
R223 OUT.n73 OUT.n47 3.23387
R224 OUT.n75 OUT.n43 3.23387
R225 OUT.n78 OUT.n35 3.23387
R226 OUT.n80 OUT.n31 3.23387
R227 OUT.n69 OUT.n57 3.23383
R228 OUT.n67 OUT.n61 3.23383
R229 OUT.n71 OUT.n51 3.23383
R230 OUT.n82 OUT.n25 3.23358
R231 OUT.n66 OUT.n65 3.2335
R232 OUT.n85 OUT.n19 3.23343
R233 OUT.n87 OUT.n15 3.23343
R234 OUT.n86 OUT.n17 3.23337
R235 OUT.n79 OUT.n33 3.23316
R236 OUT.n77 OUT.n37 3.23312
R237 OUT.n74 OUT.n45 3.23312
R238 OUT.n72 OUT.n49 3.23312
R239 OUT.n70 OUT.n53 3.23312
R240 OUT.n66 OUT.n63 3.2315
R241 OUT.n100 OUT.n97 2.98385
R242 OUT.n113 OUT.n95 2.87549
R243 OUT.n116 OUT.n115 2.70972
R244 OUT.n119 OUT.n118 2.62238
R245 OUT.n122 OUT.n121 2.62091
R246 OUT.n125 OUT.n124 2.61945
R247 OUT.n131 OUT.n130 2.61636
R248 OUT.n137 OUT.n136 2.61619
R249 OUT.n128 OUT.n127 2.61619
R250 OUT.n134 OUT.n133 2.61554
R251 OUT.n13 OUT.n12 2.6005
R252 OUT.n91 OUT.n90 2.6005
R253 OUT.n100 OUT.n99 2.58236
R254 OUT.n106 OUT.n105 2.58184
R255 OUT.n109 OUT.n108 2.5817
R256 OUT.n103 OUT.n102 2.58166
R257 OUT.n112 OUT.n111 2.58122
R258 OUT.n138 OUT.n137 1.60202
R259 OUT.n138 OUT.n93 1.34978
R260 OUT.n139 OUT.n138 0.888141
R261 OUT.n13 OUT.n10 0.79069
R262 OUT.n84 OUT.n83 0.781777
R263 OUT.n81 OUT.n80 0.781777
R264 OUT.n76 OUT.n75 0.781777
R265 OUT.n69 OUT.n68 0.781777
R266 OUT.n67 OUT.n66 0.781777
R267 OUT.n82 OUT.n81 0.779862
R268 OUT.n79 OUT.n78 0.779862
R269 OUT.n77 OUT.n76 0.779862
R270 OUT.n74 OUT.n73 0.779862
R271 OUT.n72 OUT.n71 0.779862
R272 OUT.n70 OUT.n69 0.779862
R273 OUT.n88 OUT.n87 0.777947
R274 OUT.n86 OUT.n85 0.777947
R275 OUT.n139 OUT.n91 0.655477
R276 OUT.n90 OUT.t73 0.6505
R277 OUT.n90 OUT.n89 0.6505
R278 OUT.n12 OUT.t64 0.6505
R279 OUT.n12 OUT.n11 0.6505
R280 OUT.n1 OUT.t60 0.6505
R281 OUT.n1 OUT.n0 0.6505
R282 OUT.n3 OUT.t74 0.6505
R283 OUT.n3 OUT.n2 0.6505
R284 OUT.n5 OUT.t69 0.6505
R285 OUT.n5 OUT.n4 0.6505
R286 OUT.n7 OUT.t50 0.6505
R287 OUT.n7 OUT.n6 0.6505
R288 OUT.n17 OUT.t48 0.6505
R289 OUT.n17 OUT.n16 0.6505
R290 OUT.n21 OUT.t58 0.6505
R291 OUT.n21 OUT.n20 0.6505
R292 OUT.n25 OUT.t67 0.6505
R293 OUT.n25 OUT.n24 0.6505
R294 OUT.n29 OUT.t46 0.6505
R295 OUT.n29 OUT.n28 0.6505
R296 OUT.n27 OUT.t66 0.6505
R297 OUT.n27 OUT.n26 0.6505
R298 OUT.n33 OUT.t54 0.6505
R299 OUT.n33 OUT.n32 0.6505
R300 OUT.n37 OUT.t59 0.6505
R301 OUT.n37 OUT.n36 0.6505
R302 OUT.n41 OUT.t62 0.6505
R303 OUT.n41 OUT.n40 0.6505
R304 OUT.n39 OUT.t52 0.6505
R305 OUT.n39 OUT.n38 0.6505
R306 OUT.n45 OUT.t56 0.6505
R307 OUT.n45 OUT.n44 0.6505
R308 OUT.n49 OUT.t55 0.6505
R309 OUT.n49 OUT.n48 0.6505
R310 OUT.n53 OUT.t49 0.6505
R311 OUT.n53 OUT.n52 0.6505
R312 OUT.n57 OUT.t51 0.6505
R313 OUT.n57 OUT.n56 0.6505
R314 OUT.n55 OUT.t47 0.6505
R315 OUT.n55 OUT.n54 0.6505
R316 OUT.n59 OUT.t53 0.6505
R317 OUT.n59 OUT.n58 0.6505
R318 OUT.n65 OUT.t76 0.6505
R319 OUT.n65 OUT.n64 0.6505
R320 OUT.n63 OUT.t57 0.6505
R321 OUT.n63 OUT.n62 0.6505
R322 OUT.n61 OUT.t45 0.6505
R323 OUT.n61 OUT.n60 0.6505
R324 OUT.n51 OUT.t68 0.6505
R325 OUT.n51 OUT.n50 0.6505
R326 OUT.n47 OUT.t75 0.6505
R327 OUT.n47 OUT.n46 0.6505
R328 OUT.n43 OUT.t61 0.6505
R329 OUT.n43 OUT.n42 0.6505
R330 OUT.n35 OUT.t70 0.6505
R331 OUT.n35 OUT.n34 0.6505
R332 OUT.n31 OUT.t71 0.6505
R333 OUT.n31 OUT.n30 0.6505
R334 OUT.n23 OUT.t63 0.6505
R335 OUT.n23 OUT.n22 0.6505
R336 OUT.n19 OUT.t65 0.6505
R337 OUT.n19 OUT.n18 0.6505
R338 OUT.n15 OUT.t72 0.6505
R339 OUT.n15 OUT.n14 0.6505
R340 OUT.n91 OUT.n88 0.633955
R341 OUT.n88 OUT.n13 0.631666
R342 OUT.n127 OUT.t18 0.5855
R343 OUT.n127 OUT.n126 0.5855
R344 OUT.n133 OUT.t20 0.5855
R345 OUT.n133 OUT.n132 0.5855
R346 OUT.n136 OUT.t26 0.5855
R347 OUT.n136 OUT.n135 0.5855
R348 OUT.n115 OUT.t30 0.5855
R349 OUT.n115 OUT.n114 0.5855
R350 OUT.n118 OUT.t31 0.5855
R351 OUT.n118 OUT.n117 0.5855
R352 OUT.n121 OUT.t25 0.5855
R353 OUT.n121 OUT.n120 0.5855
R354 OUT.n124 OUT.t32 0.5855
R355 OUT.n124 OUT.n123 0.5855
R356 OUT.n130 OUT.t19 0.5855
R357 OUT.n130 OUT.n129 0.5855
R358 OUT.n97 OUT.t23 0.5855
R359 OUT.n97 OUT.n96 0.5855
R360 OUT.n99 OUT.t24 0.5855
R361 OUT.n99 OUT.n98 0.5855
R362 OUT.n102 OUT.t29 0.5855
R363 OUT.n102 OUT.n101 0.5855
R364 OUT.n105 OUT.t21 0.5855
R365 OUT.n105 OUT.n104 0.5855
R366 OUT.n108 OUT.t22 0.5855
R367 OUT.n108 OUT.n107 0.5855
R368 OUT.n111 OUT.t27 0.5855
R369 OUT.n111 OUT.n110 0.5855
R370 OUT.n95 OUT.t28 0.5855
R371 OUT.n95 OUT.n94 0.5855
R372 OUT.n93 OUT.t33 0.5855
R373 OUT.n93 OUT.n92 0.5855
R374 OUT.n116 OUT.n113 0.510866
R375 OUT.n10 OUT.n9 0.504747
R376 OUT.n9 OUT.n8 0.504747
R377 OUT.n106 OUT.n103 0.403414
R378 OUT.n109 OUT.n106 0.402304
R379 OUT.n112 OUT.n109 0.400958
R380 OUT.n103 OUT.n100 0.400949
R381 OUT OUT.n139 0.354162
R382 OUT.n128 OUT.n125 0.334681
R383 OUT.n131 OUT.n128 0.334473
R384 OUT.n122 OUT.n119 0.334465
R385 OUT.n134 OUT.n131 0.334064
R386 OUT.n137 OUT.n134 0.333663
R387 OUT.n125 OUT.n122 0.333454
R388 OUT.n119 OUT.n116 0.244714
R389 OUT.n113 OUT.n112 0.107492
R390 OUT.n87 OUT.n86 0.00432979
R391 OUT.n85 OUT.n84 0.00241489
R392 OUT.n83 OUT.n82 0.00241489
R393 OUT.n80 OUT.n79 0.00241489
R394 OUT.n78 OUT.n77 0.00241489
R395 OUT.n75 OUT.n74 0.00241489
R396 OUT.n73 OUT.n72 0.00241489
R397 OUT.n71 OUT.n70 0.00241489
R398 OUT.n68 OUT.n67 0.00241489
R399 VDD.t22 VDD.t77 85.5351
R400 VDD.t64 VDD.t0 85.5351
R401 VDD.n100 VDD.t16 75.0529
R402 VDD.n103 VDD.t24 67.925
R403 VDD.n106 VDD.t10 62.055
R404 VDD.n109 VDD.t55 56.185
R405 VDD.n113 VDD.t83 51.1535
R406 VDD.n97 VDD.t88 46.9607
R407 VDD.n131 VDD.t42 46.9607
R408 VDD.n142 VDD.t5 46.5414
R409 VDD.n120 VDD.t29 44.0257
R410 VDD.n120 VDD.t37 41.5099
R411 VDD.n142 VDD.t64 38.9942
R412 VDD.n97 VDD.t47 38.5749
R413 VDD.n131 VDD.t19 38.5749
R414 VDD.n113 VDD.t31 34.382
R415 VDD.n128 VDD.t2 30.1892
R416 VDD.n139 VDD.t7 29.7699
R417 VDD.n109 VDD.t45 29.3506
R418 VDD.n106 VDD.t33 23.4806
R419 VDD.n132 VDD.t72 21.3841
R420 VDD.n121 VDD.t52 20.9649
R421 VDD.n103 VDD.t27 17.6106
R422 VDD.n125 VDD.t50 12.9984
R423 VDD.n136 VDD.t67 12.5791
R424 VDD.n100 VDD.t22 10.4827
R425 VDD.n98 VDD.n97 6.3005
R426 VDD.n101 VDD.n100 6.3005
R427 VDD.n104 VDD.n103 6.3005
R428 VDD.n107 VDD.n106 6.3005
R429 VDD.n110 VDD.n109 6.3005
R430 VDD.n159 VDD.n120 6.3005
R431 VDD.n158 VDD.n121 6.3005
R432 VDD.n156 VDD.n124 6.3005
R433 VDD.n155 VDD.n125 6.3005
R434 VDD.n153 VDD.n128 6.3005
R435 VDD.n151 VDD.n131 6.3005
R436 VDD.n150 VDD.n132 6.3005
R437 VDD.n148 VDD.n135 6.3005
R438 VDD.n147 VDD.n136 6.3005
R439 VDD.n145 VDD.n139 6.3005
R440 VDD.n143 VDD.n142 6.3005
R441 VDD.n143 VDD.t1 4.21354
R442 VDD.n124 VDD.t61 4.19337
R443 VDD.n135 VDD.t13 4.19337
R444 VDD.n14 VDD.t80 3.28543
R445 VDD.n55 VDD.t122 3.27944
R446 VDD.n144 VDD.n141 3.27159
R447 VDD.n149 VDD.n134 3.27159
R448 VDD.n152 VDD.n130 3.27159
R449 VDD.n154 VDD.n127 3.27159
R450 VDD.n157 VDD.n123 3.27159
R451 VDD.n160 VDD.n119 3.27159
R452 VDD.n161 VDD.n117 3.27159
R453 VDD.n111 VDD.n1 3.27159
R454 VDD.n105 VDD.n5 3.27159
R455 VDD.n102 VDD.n7 3.27159
R456 VDD.n99 VDD.n9 3.27159
R457 VDD.n146 VDD.n138 3.26834
R458 VDD.n108 VDD.n3 3.26449
R459 VDD.n96 VDD.n10 3.2505
R460 VDD.n115 VDD.n114 3.1505
R461 VDD.n114 VDD.n113 3.1505
R462 VDD.n91 VDD.n90 2.42419
R463 VDD.n79 VDD.n78 2.42339
R464 VDD.n76 VDD.n75 2.42315
R465 VDD.n82 VDD.n81 2.42282
R466 VDD.n88 VDD.n87 2.42265
R467 VDD.n85 VDD.n84 2.42222
R468 VDD.n73 VDD.n72 2.42152
R469 VDD.n70 VDD.n69 2.41849
R470 VDD.n67 VDD.n66 2.41843
R471 VDD.n64 VDD.n63 2.41556
R472 VDD.n61 VDD.n60 2.41444
R473 VDD.n50 VDD.n49 2.41251
R474 VDD.n58 VDD.n57 2.41018
R475 VDD.n47 VDD.n46 2.41016
R476 VDD.n55 VDD.n54 2.40994
R477 VDD.n14 VDD.n13 2.40758
R478 VDD.n20 VDD.n19 2.40707
R479 VDD.n44 VDD.n43 2.40667
R480 VDD.n17 VDD.n16 2.40626
R481 VDD.n23 VDD.n22 2.40299
R482 VDD.n26 VDD.n25 2.40275
R483 VDD.n38 VDD.n37 2.4026
R484 VDD.n41 VDD.n40 2.40255
R485 VDD.n35 VDD.n34 2.40212
R486 VDD.n29 VDD.n28 2.40139
R487 VDD.n32 VDD.n31 2.40019
R488 VDD.n95 VDD.n94 2.38241
R489 VDD.n51 VDD.n11 1.91067
R490 VDD.n51 VDD.n50 1.38687
R491 VDD.n92 VDD.n91 1.34148
R492 VDD.n96 VDD.n95 1.25144
R493 VDD.n52 VDD.n51 0.996686
R494 VDD.n98 VDD.n96 0.828172
R495 VDD.n141 VDD.t6 0.6505
R496 VDD.n141 VDD.n140 0.6505
R497 VDD.n138 VDD.t144 0.6505
R498 VDD.n138 VDD.n137 0.6505
R499 VDD.n134 VDD.t143 0.6505
R500 VDD.n134 VDD.n133 0.6505
R501 VDD.n130 VDD.t130 0.6505
R502 VDD.n130 VDD.n129 0.6505
R503 VDD.n127 VDD.t137 0.6505
R504 VDD.n127 VDD.n126 0.6505
R505 VDD.n123 VDD.t150 0.6505
R506 VDD.n123 VDD.n122 0.6505
R507 VDD.n119 VDD.t149 0.6505
R508 VDD.n119 VDD.n118 0.6505
R509 VDD.n117 VDD.t140 0.6505
R510 VDD.n117 VDD.n116 0.6505
R511 VDD.n1 VDD.t153 0.6505
R512 VDD.n1 VDD.n0 0.6505
R513 VDD.n3 VDD.t34 0.6505
R514 VDD.n3 VDD.n2 0.6505
R515 VDD.n5 VDD.t125 0.6505
R516 VDD.n5 VDD.n4 0.6505
R517 VDD.n7 VDD.t23 0.6505
R518 VDD.n7 VDD.n6 0.6505
R519 VDD.n9 VDD.t103 0.6505
R520 VDD.n9 VDD.n8 0.6505
R521 VDD.n78 VDD.t116 0.6505
R522 VDD.n78 VDD.n77 0.6505
R523 VDD.n54 VDD.t87 0.6505
R524 VDD.n54 VDD.n53 0.6505
R525 VDD.n57 VDD.t68 0.6505
R526 VDD.n57 VDD.n56 0.6505
R527 VDD.n60 VDD.t73 0.6505
R528 VDD.n60 VDD.n59 0.6505
R529 VDD.n63 VDD.t75 0.6505
R530 VDD.n63 VDD.n62 0.6505
R531 VDD.n66 VDD.t121 0.6505
R532 VDD.n66 VDD.n65 0.6505
R533 VDD.n69 VDD.t86 0.6505
R534 VDD.n69 VDD.n68 0.6505
R535 VDD.n72 VDD.t30 0.6505
R536 VDD.n72 VDD.n71 0.6505
R537 VDD.n75 VDD.t32 0.6505
R538 VDD.n75 VDD.n74 0.6505
R539 VDD.n81 VDD.t49 0.6505
R540 VDD.n81 VDD.n80 0.6505
R541 VDD.n84 VDD.t28 0.6505
R542 VDD.n84 VDD.n83 0.6505
R543 VDD.n87 VDD.t70 0.6505
R544 VDD.n87 VDD.n86 0.6505
R545 VDD.n90 VDD.t74 0.6505
R546 VDD.n90 VDD.n89 0.6505
R547 VDD.n94 VDD.n93 0.6505
R548 VDD.n13 VDD.t81 0.6505
R549 VDD.n13 VDD.n12 0.6505
R550 VDD.n16 VDD.t82 0.6505
R551 VDD.n16 VDD.n15 0.6505
R552 VDD.n19 VDD.t76 0.6505
R553 VDD.n19 VDD.n18 0.6505
R554 VDD.n22 VDD.t43 0.6505
R555 VDD.n22 VDD.n21 0.6505
R556 VDD.n25 VDD.t51 0.6505
R557 VDD.n25 VDD.n24 0.6505
R558 VDD.n28 VDD.t53 0.6505
R559 VDD.n28 VDD.n27 0.6505
R560 VDD.n31 VDD.t69 0.6505
R561 VDD.n31 VDD.n30 0.6505
R562 VDD.n34 VDD.t44 0.6505
R563 VDD.n34 VDD.n33 0.6505
R564 VDD.n37 VDD.t46 0.6505
R565 VDD.n37 VDD.n36 0.6505
R566 VDD.n40 VDD.t54 0.6505
R567 VDD.n40 VDD.n39 0.6505
R568 VDD.n43 VDD.t58 0.6505
R569 VDD.n43 VDD.n42 0.6505
R570 VDD.n46 VDD.t71 0.6505
R571 VDD.n46 VDD.n45 0.6505
R572 VDD.n49 VDD.t48 0.6505
R573 VDD.n49 VDD.n48 0.6505
R574 VDD.n161 VDD.n160 0.299037
R575 VDD.n115 VDD.n111 0.284402
R576 VDD.n110 VDD.n108 0.275622
R577 VDD.n92 VDD.n52 0.265556
R578 VDD.n107 VDD.n105 0.265378
R579 VDD.n104 VDD.n102 0.255134
R580 VDD.n47 VDD.n44 0.235837
R581 VDD.n32 VDD.n29 0.23543
R582 VDD.n35 VDD.n32 0.235271
R583 VDD.n23 VDD.n20 0.234863
R584 VDD.n29 VDD.n26 0.234297
R585 VDD.n26 VDD.n23 0.234297
R586 VDD.n17 VDD.n14 0.234293
R587 VDD.n50 VDD.n47 0.234291
R588 VDD.n38 VDD.n35 0.233514
R589 VDD.n44 VDD.n41 0.233447
R590 VDD.n20 VDD.n17 0.233445
R591 VDD.n41 VDD.n38 0.233389
R592 VDD.n91 VDD.n88 0.226747
R593 VDD.n79 VDD.n76 0.225529
R594 VDD.n70 VDD.n67 0.225387
R595 VDD.n85 VDD.n82 0.225121
R596 VDD.n67 VDD.n64 0.225121
R597 VDD.n76 VDD.n73 0.22512
R598 VDD.n61 VDD.n58 0.22512
R599 VDD.n64 VDD.n61 0.224578
R600 VDD.n58 VDD.n55 0.223901
R601 VDD.n82 VDD.n79 0.22363
R602 VDD.n88 VDD.n85 0.222816
R603 VDD.n73 VDD.n70 0.22281
R604 VDD.n101 VDD.n99 0.20611
R605 VDD.n159 VDD.n158 0.185622
R606 VDD.n156 VDD.n155 0.179768
R607 VDD.n151 VDD.n150 0.179768
R608 VDD.n148 VDD.n147 0.179037
R609 VDD.n145 VDD.n144 0.172451
R610 VDD.n153 VDD.n152 0.17172
R611 VDD.n114 VDD.n112 0.159994
R612 VDD.n99 VDD.n98 0.142451
R613 VDD.n154 VDD.n153 0.127817
R614 VDD.n146 VDD.n145 0.126354
R615 VDD.n150 VDD.n149 0.112451
R616 VDD.n158 VDD.n157 0.11172
R617 VDD.n102 VDD.n101 0.0934268
R618 VDD.n157 VDD.n156 0.0678171
R619 VDD.n149 VDD.n148 0.0678171
R620 VDD.n95 VDD.n92 0.0587571
R621 VDD.n147 VDD.n146 0.0539146
R622 VDD.n155 VDD.n154 0.0524512
R623 VDD.n105 VDD.n104 0.0444024
R624 VDD.n108 VDD.n107 0.0341585
R625 VDD.n111 VDD.n110 0.0239146
R626 VDD VDD.n161 0.0136707
R627 VDD.n152 VDD.n151 0.00781707
R628 VDD.n144 VDD.n143 0.00708537
R629 VDD.n160 VDD.n159 0.00269512
R630 VDD VDD.n115 0.00196341
R631 VSS.t96 VSS.t79 405.01
R632 VSS.n112 VSS.t82 295.815
R633 VSS.n126 VSS.t5 275.962
R634 VSS.n99 VSS.t100 271.991
R635 VSS.n66 VSS.t19 252.138
R636 VSS.n83 VSS.t76 248.167
R637 VSS.n70 VSS.t40 228.315
R638 VSS.n79 VSS.t28 224.344
R639 VSS.n74 VSS.t16 204.49
R640 VSS.n74 VSS.t31 200.519
R641 VSS.n79 VSS.t46 180.667
R642 VSS.n70 VSS.t25 176.696
R643 VSS.n83 VSS.t96 156.843
R644 VSS.n66 VSS.t43 152.871
R645 VSS.n99 VSS.t51 133.018
R646 VSS.n62 VSS.t22 131.879
R647 VSS.n126 VSS.t0 129.048
R648 VSS.n62 VSS.t34 122.9
R649 VSS.n112 VSS.t7 109.195
R650 VSS.n113 VSS.t3 105.224
R651 VSS.n125 VSS.t69 85.3701
R652 VSS.n111 VSS.t54 81.3994
R653 VSS.n129 VSS.t102 66.746
R654 VSS.n63 VSS.t49 61.546
R655 VSS.n98 VSS.t106 57.5753
R656 VSS.n68 VSS.t10 37.7219
R657 VSS.n13 VSS.t33 36.0467
R658 VSS.n24 VSS.t27 36.0467
R659 VSS.t79 VSS.n82 33.7513
R660 VSS.n13 VSS.t21 22.6305
R661 VSS.n14 VSS.t48 22.6305
R662 VSS.n15 VSS.t18 22.6305
R663 VSS.n16 VSS.t42 22.6305
R664 VSS.n17 VSS.t9 22.6305
R665 VSS.n18 VSS.t39 22.6305
R666 VSS.n19 VSS.t24 22.6305
R667 VSS.n20 VSS.t36 22.6305
R668 VSS.n21 VSS.t15 22.6305
R669 VSS.n22 VSS.t30 22.6305
R670 VSS.n23 VSS.t12 22.6305
R671 VSS.n24 VSS.t45 22.6305
R672 VSS.n72 VSS.t37 13.8979
R673 VSS.n14 VSS.n13 13.4167
R674 VSS.n15 VSS.n14 13.4167
R675 VSS.n16 VSS.n15 13.4167
R676 VSS.n17 VSS.n16 13.4167
R677 VSS.n18 VSS.n17 13.4167
R678 VSS.n19 VSS.n18 13.4167
R679 VSS.n20 VSS.n19 13.4167
R680 VSS.n21 VSS.n20 13.4167
R681 VSS.n22 VSS.n21 13.4167
R682 VSS.n23 VSS.n22 13.4167
R683 VSS.n25 VSS.n23 13.2852
R684 VSS.n77 VSS.t13 9.92719
R685 VSS.n130 VSS.n126 5.2005
R686 VSS.n131 VSS.n125 5.2005
R687 VSS.n133 VSS.n113 5.2005
R688 VSS.n134 VSS.n112 5.2005
R689 VSS.n135 VSS.n111 5.2005
R690 VSS.n137 VSS.n99 5.2005
R691 VSS.n138 VSS.n98 5.2005
R692 VSS.n140 VSS.n83 5.2005
R693 VSS.n80 VSS.n79 5.2005
R694 VSS.n78 VSS.n77 5.2005
R695 VSS.n75 VSS.n74 5.2005
R696 VSS.n73 VSS.n72 5.2005
R697 VSS.n71 VSS.n70 5.2005
R698 VSS.n69 VSS.n68 5.2005
R699 VSS.n67 VSS.n66 5.2005
R700 VSS.n64 VSS.n63 5.2005
R701 VSS VSS.n81 5.2005
R702 VSS VSS.n81 5.2005
R703 VSS.n32 VSS.n29 5.11535
R704 VSS.n51 VSS.n25 4.42582
R705 VSS.n127 VSS.t115 4.411
R706 VSS.n106 VSS.n105 3.82995
R707 VSS.n93 VSS.n92 3.82991
R708 VSS.n120 VSS.n119 3.82991
R709 VSS.n41 VSS.n40 3.826
R710 VSS.n44 VSS.n43 3.826
R711 VSS.n47 VSS.n46 3.826
R712 VSS.n93 VSS.n90 3.826
R713 VSS.n121 VSS.n115 3.826
R714 VSS.n35 VSS.n34 3.82596
R715 VSS.n38 VSS.n37 3.82596
R716 VSS.n107 VSS.n101 3.82596
R717 VSS.n106 VSS.n103 3.82596
R718 VSS.n32 VSS.n31 3.82592
R719 VSS.n94 VSS.n88 3.82592
R720 VSS.n120 VSS.n117 3.82592
R721 VSS.n86 VSS.n85 3.78196
R722 VSS.n128 VSS.t103 3.7355
R723 VSS.n49 VSS.n28 3.16517
R724 VSS.n57 VSS.n56 3.1505
R725 VSS.n59 VSS.n58 3.1505
R726 VSS.n61 VSS.n60 3.1505
R727 VSS.n1 VSS.n0 3.1505
R728 VSS.n3 VSS.n2 3.1505
R729 VSS.n5 VSS.n4 3.1505
R730 VSS.n7 VSS.n6 3.1505
R731 VSS.n9 VSS.n8 3.1505
R732 VSS.n54 VSS.n10 3.1505
R733 VSS.n53 VSS.n11 3.1505
R734 VSS.n52 VSS.n12 3.1505
R735 VSS.n50 VSS.n26 3.1505
R736 VSS.n97 VSS.n96 3.1505
R737 VSS.n110 VSS.n109 3.1505
R738 VSS.n124 VSS.n123 3.1505
R739 VSS.n82 VSS.n81 2.6005
R740 VSS.n64 VSS.n62 2.53633
R741 VSS.n57 VSS.n55 1.81655
R742 VSS.n129 VSS.n128 0.921147
R743 VSS.n132 VSS.n124 0.869196
R744 VSS.n55 VSS.t23 0.826268
R745 VSS.n139 VSS.n97 0.782913
R746 VSS.n136 VSS.n110 0.781543
R747 VSS.n94 VSS.n86 0.749848
R748 VSS.n48 VSS.n47 0.722457
R749 VSS.n47 VSS.n44 0.708761
R750 VSS.n94 VSS.n93 0.708761
R751 VSS.n121 VSS.n120 0.708761
R752 VSS.n35 VSS.n32 0.706804
R753 VSS.n38 VSS.n35 0.706804
R754 VSS.n41 VSS.n38 0.706804
R755 VSS.n44 VSS.n41 0.706804
R756 VSS.n107 VSS.n106 0.704848
R757 VSS.n97 VSS.n94 0.679996
R758 VSS.n110 VSS.n107 0.679954
R759 VSS.n124 VSS.n121 0.679913
R760 VSS.n128 VSS.n127 0.679913
R761 VSS.n65 VSS.n61 0.659848
R762 VSS.n76 VSS.n54 0.654826
R763 VSS.n31 VSS.t95 0.5855
R764 VSS.n31 VSS.n30 0.5855
R765 VSS.n34 VSS.t94 0.5855
R766 VSS.n34 VSS.n33 0.5855
R767 VSS.n37 VSS.t89 0.5855
R768 VSS.n37 VSS.n36 0.5855
R769 VSS.n40 VSS.t98 0.5855
R770 VSS.n40 VSS.n39 0.5855
R771 VSS.n43 VSS.t93 0.5855
R772 VSS.n43 VSS.n42 0.5855
R773 VSS.n46 VSS.t92 0.5855
R774 VSS.n46 VSS.n45 0.5855
R775 VSS.n85 VSS.t105 0.5855
R776 VSS.n85 VSS.n84 0.5855
R777 VSS.n26 VSS.t29 0.5855
R778 VSS.n12 VSS.t47 0.5855
R779 VSS.n11 VSS.t14 0.5855
R780 VSS.n10 VSS.t17 0.5855
R781 VSS.n10 VSS.t32 0.5855
R782 VSS.n8 VSS.t38 0.5855
R783 VSS.n6 VSS.t26 0.5855
R784 VSS.n4 VSS.t41 0.5855
R785 VSS.n2 VSS.t11 0.5855
R786 VSS.n60 VSS.t20 0.5855
R787 VSS.n60 VSS.t44 0.5855
R788 VSS.n58 VSS.t50 0.5855
R789 VSS.n28 VSS.n27 0.5855
R790 VSS.n88 VSS.t104 0.5855
R791 VSS.n88 VSS.n87 0.5855
R792 VSS.n96 VSS.t97 0.5855
R793 VSS.n96 VSS.n95 0.5855
R794 VSS.n90 VSS.t112 0.5855
R795 VSS.n90 VSS.n89 0.5855
R796 VSS.n92 VSS.t107 0.5855
R797 VSS.n92 VSS.n91 0.5855
R798 VSS.n101 VSS.t116 0.5855
R799 VSS.n101 VSS.n100 0.5855
R800 VSS.n109 VSS.t101 0.5855
R801 VSS.n109 VSS.n108 0.5855
R802 VSS.n103 VSS.t8 0.5855
R803 VSS.n103 VSS.n102 0.5855
R804 VSS.n105 VSS.t99 0.5855
R805 VSS.n105 VSS.n104 0.5855
R806 VSS.n115 VSS.t4 0.5855
R807 VSS.n115 VSS.n114 0.5855
R808 VSS.n123 VSS.t91 0.5855
R809 VSS.n123 VSS.n122 0.5855
R810 VSS.n117 VSS.t6 0.5855
R811 VSS.n117 VSS.n116 0.5855
R812 VSS.n119 VSS.t90 0.5855
R813 VSS.n119 VSS.n118 0.5855
R814 VSS.n49 VSS.n48 0.354579
R815 VSS.n55 VSS.t35 0.301111
R816 VSS.n69 VSS.n67 0.220012
R817 VSS.n71 VSS.n69 0.220012
R818 VSS.n73 VSS.n71 0.220012
R819 VSS.n75 VSS.n73 0.220012
R820 VSS.n80 VSS.n78 0.220012
R821 VSS VSS.n80 0.220012
R822 VSS VSS.n140 0.220012
R823 VSS.n138 VSS.n137 0.220012
R824 VSS.n135 VSS.n134 0.220012
R825 VSS.n134 VSS.n133 0.220012
R826 VSS.n131 VSS.n130 0.220012
R827 VSS.n130 VSS.n129 0.220012
R828 VSS.n78 VSS.n76 0.216354
R829 VSS.n65 VSS.n64 0.20172
R830 VSS.n139 VSS.n138 0.200988
R831 VSS.n59 VSS.n57 0.200065
R832 VSS.n61 VSS.n59 0.200065
R833 VSS.n3 VSS.n1 0.200065
R834 VSS.n5 VSS.n3 0.200065
R835 VSS.n7 VSS.n5 0.200065
R836 VSS.n9 VSS.n7 0.200065
R837 VSS.n54 VSS.n9 0.200065
R838 VSS.n54 VSS.n53 0.200065
R839 VSS.n53 VSS.n52 0.200065
R840 VSS.n50 VSS.n49 0.185391
R841 VSS.n137 VSS.n136 0.174646
R842 VSS.n25 VSS.n24 0.132032
R843 VSS.n133 VSS.n132 0.113915
R844 VSS.n132 VSS.n131 0.106598
R845 VSS.n51 VSS.n50 0.101261
R846 VSS.n52 VSS.n51 0.0993043
R847 VSS.n136 VSS.n135 0.0458659
R848 VSS.n140 VSS.n139 0.0195244
R849 VSS.n67 VSS.n65 0.0187927
R850 VSS.n76 VSS.n75 0.00415854
R851 IN.n3 IN.t5 37.6513
R852 IN IN.n3 34.0473
R853 IN.n0 IN.t4 32.7094
R854 IN IN.n2 25.749
R855 IN.n0 IN.t3 23.2875
R856 IN.n1 IN.t2 23.2875
R857 IN.n3 IN.t0 20.4405
R858 IN.n2 IN.t1 20.4405
R859 IN.n1 IN.n0 12.5148
R860 IN.n2 IN.n1 12.2081
R861 a_240_n2164.n26 a_240_n2164.n25 72.9524
R862 a_240_n2164.n20 a_240_n2164.t25 44.8231
R863 a_240_n2164.n2 a_240_n2164.t22 36.4904
R864 a_240_n2164.n26 a_240_n2164.t12 23.7985
R865 a_240_n2164.n2 a_240_n2164.t28 23.6525
R866 a_240_n2164.n3 a_240_n2164.t24 23.6525
R867 a_240_n2164.n4 a_240_n2164.t21 23.6525
R868 a_240_n2164.n5 a_240_n2164.t18 23.6525
R869 a_240_n2164.n6 a_240_n2164.t15 23.6525
R870 a_240_n2164.n7 a_240_n2164.t20 23.6525
R871 a_240_n2164.n8 a_240_n2164.t16 23.6525
R872 a_240_n2164.n9 a_240_n2164.t14 23.6525
R873 a_240_n2164.n10 a_240_n2164.t10 23.6525
R874 a_240_n2164.n11 a_240_n2164.t8 23.6525
R875 a_240_n2164.n12 a_240_n2164.t13 23.6525
R876 a_240_n2164.n13 a_240_n2164.t9 23.6525
R877 a_240_n2164.n14 a_240_n2164.t29 23.6525
R878 a_240_n2164.n15 a_240_n2164.t27 23.6525
R879 a_240_n2164.n16 a_240_n2164.t19 23.6525
R880 a_240_n2164.n21 a_240_n2164.n20 23.3438
R881 a_240_n2164.n22 a_240_n2164.n21 23.3438
R882 a_240_n2164.n23 a_240_n2164.n22 23.3438
R883 a_240_n2164.n24 a_240_n2164.n23 23.3438
R884 a_240_n2164.n25 a_240_n2164.n24 23.3438
R885 a_240_n2164.n20 a_240_n2164.t6 20.4405
R886 a_240_n2164.n21 a_240_n2164.t26 20.4405
R887 a_240_n2164.n22 a_240_n2164.t7 20.4405
R888 a_240_n2164.n23 a_240_n2164.t17 20.4405
R889 a_240_n2164.n24 a_240_n2164.t11 20.4405
R890 a_240_n2164.n25 a_240_n2164.t23 20.4405
R891 a_240_n2164.n3 a_240_n2164.n2 12.8384
R892 a_240_n2164.n4 a_240_n2164.n3 12.8384
R893 a_240_n2164.n5 a_240_n2164.n4 12.8384
R894 a_240_n2164.n6 a_240_n2164.n5 12.8384
R895 a_240_n2164.n7 a_240_n2164.n6 12.8384
R896 a_240_n2164.n8 a_240_n2164.n7 12.8384
R897 a_240_n2164.n9 a_240_n2164.n8 12.8384
R898 a_240_n2164.n10 a_240_n2164.n9 12.8384
R899 a_240_n2164.n11 a_240_n2164.n10 12.8384
R900 a_240_n2164.n12 a_240_n2164.n11 12.8384
R901 a_240_n2164.n13 a_240_n2164.n12 12.8384
R902 a_240_n2164.n14 a_240_n2164.n13 12.8384
R903 a_240_n2164.n15 a_240_n2164.n14 12.8384
R904 a_240_n2164.n16 a_240_n2164.n15 12.8384
R905 a_240_n2164.n27 a_240_n2164.n26 6.95492
R906 a_240_n2164.n17 a_240_n2164.n16 4.78319
R907 a_240_n2164.n28 a_240_n2164.n27 4.13676
R908 a_240_n2164.n27 a_240_n2164.n19 3.79615
R909 a_240_n2164.n17 a_240_n2164.n1 3.22711
R910 a_240_n2164.n29 a_240_n2164.n28 3.22482
R911 a_240_n2164.n1 a_240_n2164.t2 0.6505
R912 a_240_n2164.n1 a_240_n2164.n0 0.6505
R913 a_240_n2164.n29 a_240_n2164.t4 0.6505
R914 a_240_n2164.n30 a_240_n2164.n29 0.6505
R915 a_240_n2164.n19 a_240_n2164.t0 0.5855
R916 a_240_n2164.n19 a_240_n2164.n18 0.5855
R917 a_240_n2164.n28 a_240_n2164.n17 0.471269
C0 VDD IN 1.11f
C1 IN OUT 0.0149f
C2 VDD OUT 14.6f
.ends

