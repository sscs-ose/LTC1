magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2102 -4553 2102 4553
<< psubdiff >>
rect -102 2531 102 2553
rect -102 2485 -80 2531
rect -34 2485 34 2531
rect 80 2485 102 2531
rect -102 2417 102 2485
rect -102 2371 -80 2417
rect -34 2371 34 2417
rect 80 2371 102 2417
rect -102 2303 102 2371
rect -102 2257 -80 2303
rect -34 2257 34 2303
rect 80 2257 102 2303
rect -102 2189 102 2257
rect -102 2143 -80 2189
rect -34 2143 34 2189
rect 80 2143 102 2189
rect -102 2075 102 2143
rect -102 2029 -80 2075
rect -34 2029 34 2075
rect 80 2029 102 2075
rect -102 1961 102 2029
rect -102 1915 -80 1961
rect -34 1915 34 1961
rect 80 1915 102 1961
rect -102 1847 102 1915
rect -102 1801 -80 1847
rect -34 1801 34 1847
rect 80 1801 102 1847
rect -102 1733 102 1801
rect -102 1687 -80 1733
rect -34 1687 34 1733
rect 80 1687 102 1733
rect -102 1619 102 1687
rect -102 1573 -80 1619
rect -34 1573 34 1619
rect 80 1573 102 1619
rect -102 1505 102 1573
rect -102 1459 -80 1505
rect -34 1459 34 1505
rect 80 1459 102 1505
rect -102 1391 102 1459
rect -102 1345 -80 1391
rect -34 1345 34 1391
rect 80 1345 102 1391
rect -102 1277 102 1345
rect -102 1231 -80 1277
rect -34 1231 34 1277
rect 80 1231 102 1277
rect -102 1163 102 1231
rect -102 1117 -80 1163
rect -34 1117 34 1163
rect 80 1117 102 1163
rect -102 1049 102 1117
rect -102 1003 -80 1049
rect -34 1003 34 1049
rect 80 1003 102 1049
rect -102 935 102 1003
rect -102 889 -80 935
rect -34 889 34 935
rect 80 889 102 935
rect -102 821 102 889
rect -102 775 -80 821
rect -34 775 34 821
rect 80 775 102 821
rect -102 707 102 775
rect -102 661 -80 707
rect -34 661 34 707
rect 80 661 102 707
rect -102 593 102 661
rect -102 547 -80 593
rect -34 547 34 593
rect 80 547 102 593
rect -102 479 102 547
rect -102 433 -80 479
rect -34 433 34 479
rect 80 433 102 479
rect -102 365 102 433
rect -102 319 -80 365
rect -34 319 34 365
rect 80 319 102 365
rect -102 251 102 319
rect -102 205 -80 251
rect -34 205 34 251
rect 80 205 102 251
rect -102 137 102 205
rect -102 91 -80 137
rect -34 91 34 137
rect 80 91 102 137
rect -102 23 102 91
rect -102 -23 -80 23
rect -34 -23 34 23
rect 80 -23 102 23
rect -102 -91 102 -23
rect -102 -137 -80 -91
rect -34 -137 34 -91
rect 80 -137 102 -91
rect -102 -205 102 -137
rect -102 -251 -80 -205
rect -34 -251 34 -205
rect 80 -251 102 -205
rect -102 -319 102 -251
rect -102 -365 -80 -319
rect -34 -365 34 -319
rect 80 -365 102 -319
rect -102 -433 102 -365
rect -102 -479 -80 -433
rect -34 -479 34 -433
rect 80 -479 102 -433
rect -102 -547 102 -479
rect -102 -593 -80 -547
rect -34 -593 34 -547
rect 80 -593 102 -547
rect -102 -661 102 -593
rect -102 -707 -80 -661
rect -34 -707 34 -661
rect 80 -707 102 -661
rect -102 -775 102 -707
rect -102 -821 -80 -775
rect -34 -821 34 -775
rect 80 -821 102 -775
rect -102 -889 102 -821
rect -102 -935 -80 -889
rect -34 -935 34 -889
rect 80 -935 102 -889
rect -102 -1003 102 -935
rect -102 -1049 -80 -1003
rect -34 -1049 34 -1003
rect 80 -1049 102 -1003
rect -102 -1117 102 -1049
rect -102 -1163 -80 -1117
rect -34 -1163 34 -1117
rect 80 -1163 102 -1117
rect -102 -1231 102 -1163
rect -102 -1277 -80 -1231
rect -34 -1277 34 -1231
rect 80 -1277 102 -1231
rect -102 -1345 102 -1277
rect -102 -1391 -80 -1345
rect -34 -1391 34 -1345
rect 80 -1391 102 -1345
rect -102 -1459 102 -1391
rect -102 -1505 -80 -1459
rect -34 -1505 34 -1459
rect 80 -1505 102 -1459
rect -102 -1573 102 -1505
rect -102 -1619 -80 -1573
rect -34 -1619 34 -1573
rect 80 -1619 102 -1573
rect -102 -1687 102 -1619
rect -102 -1733 -80 -1687
rect -34 -1733 34 -1687
rect 80 -1733 102 -1687
rect -102 -1801 102 -1733
rect -102 -1847 -80 -1801
rect -34 -1847 34 -1801
rect 80 -1847 102 -1801
rect -102 -1915 102 -1847
rect -102 -1961 -80 -1915
rect -34 -1961 34 -1915
rect 80 -1961 102 -1915
rect -102 -2029 102 -1961
rect -102 -2075 -80 -2029
rect -34 -2075 34 -2029
rect 80 -2075 102 -2029
rect -102 -2143 102 -2075
rect -102 -2189 -80 -2143
rect -34 -2189 34 -2143
rect 80 -2189 102 -2143
rect -102 -2257 102 -2189
rect -102 -2303 -80 -2257
rect -34 -2303 34 -2257
rect 80 -2303 102 -2257
rect -102 -2371 102 -2303
rect -102 -2417 -80 -2371
rect -34 -2417 34 -2371
rect 80 -2417 102 -2371
rect -102 -2485 102 -2417
rect -102 -2531 -80 -2485
rect -34 -2531 34 -2485
rect 80 -2531 102 -2485
rect -102 -2553 102 -2531
<< psubdiffcont >>
rect -80 2485 -34 2531
rect 34 2485 80 2531
rect -80 2371 -34 2417
rect 34 2371 80 2417
rect -80 2257 -34 2303
rect 34 2257 80 2303
rect -80 2143 -34 2189
rect 34 2143 80 2189
rect -80 2029 -34 2075
rect 34 2029 80 2075
rect -80 1915 -34 1961
rect 34 1915 80 1961
rect -80 1801 -34 1847
rect 34 1801 80 1847
rect -80 1687 -34 1733
rect 34 1687 80 1733
rect -80 1573 -34 1619
rect 34 1573 80 1619
rect -80 1459 -34 1505
rect 34 1459 80 1505
rect -80 1345 -34 1391
rect 34 1345 80 1391
rect -80 1231 -34 1277
rect 34 1231 80 1277
rect -80 1117 -34 1163
rect 34 1117 80 1163
rect -80 1003 -34 1049
rect 34 1003 80 1049
rect -80 889 -34 935
rect 34 889 80 935
rect -80 775 -34 821
rect 34 775 80 821
rect -80 661 -34 707
rect 34 661 80 707
rect -80 547 -34 593
rect 34 547 80 593
rect -80 433 -34 479
rect 34 433 80 479
rect -80 319 -34 365
rect 34 319 80 365
rect -80 205 -34 251
rect 34 205 80 251
rect -80 91 -34 137
rect 34 91 80 137
rect -80 -23 -34 23
rect 34 -23 80 23
rect -80 -137 -34 -91
rect 34 -137 80 -91
rect -80 -251 -34 -205
rect 34 -251 80 -205
rect -80 -365 -34 -319
rect 34 -365 80 -319
rect -80 -479 -34 -433
rect 34 -479 80 -433
rect -80 -593 -34 -547
rect 34 -593 80 -547
rect -80 -707 -34 -661
rect 34 -707 80 -661
rect -80 -821 -34 -775
rect 34 -821 80 -775
rect -80 -935 -34 -889
rect 34 -935 80 -889
rect -80 -1049 -34 -1003
rect 34 -1049 80 -1003
rect -80 -1163 -34 -1117
rect 34 -1163 80 -1117
rect -80 -1277 -34 -1231
rect 34 -1277 80 -1231
rect -80 -1391 -34 -1345
rect 34 -1391 80 -1345
rect -80 -1505 -34 -1459
rect 34 -1505 80 -1459
rect -80 -1619 -34 -1573
rect 34 -1619 80 -1573
rect -80 -1733 -34 -1687
rect 34 -1733 80 -1687
rect -80 -1847 -34 -1801
rect 34 -1847 80 -1801
rect -80 -1961 -34 -1915
rect 34 -1961 80 -1915
rect -80 -2075 -34 -2029
rect 34 -2075 80 -2029
rect -80 -2189 -34 -2143
rect 34 -2189 80 -2143
rect -80 -2303 -34 -2257
rect 34 -2303 80 -2257
rect -80 -2417 -34 -2371
rect 34 -2417 80 -2371
rect -80 -2531 -34 -2485
rect 34 -2531 80 -2485
<< metal1 >>
rect -91 2531 91 2542
rect -91 2485 -80 2531
rect -34 2485 34 2531
rect 80 2485 91 2531
rect -91 2417 91 2485
rect -91 2371 -80 2417
rect -34 2371 34 2417
rect 80 2371 91 2417
rect -91 2303 91 2371
rect -91 2257 -80 2303
rect -34 2257 34 2303
rect 80 2257 91 2303
rect -91 2189 91 2257
rect -91 2143 -80 2189
rect -34 2143 34 2189
rect 80 2143 91 2189
rect -91 2075 91 2143
rect -91 2029 -80 2075
rect -34 2029 34 2075
rect 80 2029 91 2075
rect -91 1961 91 2029
rect -91 1915 -80 1961
rect -34 1915 34 1961
rect 80 1915 91 1961
rect -91 1847 91 1915
rect -91 1801 -80 1847
rect -34 1801 34 1847
rect 80 1801 91 1847
rect -91 1733 91 1801
rect -91 1687 -80 1733
rect -34 1687 34 1733
rect 80 1687 91 1733
rect -91 1619 91 1687
rect -91 1573 -80 1619
rect -34 1573 34 1619
rect 80 1573 91 1619
rect -91 1505 91 1573
rect -91 1459 -80 1505
rect -34 1459 34 1505
rect 80 1459 91 1505
rect -91 1391 91 1459
rect -91 1345 -80 1391
rect -34 1345 34 1391
rect 80 1345 91 1391
rect -91 1277 91 1345
rect -91 1231 -80 1277
rect -34 1231 34 1277
rect 80 1231 91 1277
rect -91 1163 91 1231
rect -91 1117 -80 1163
rect -34 1117 34 1163
rect 80 1117 91 1163
rect -91 1049 91 1117
rect -91 1003 -80 1049
rect -34 1003 34 1049
rect 80 1003 91 1049
rect -91 935 91 1003
rect -91 889 -80 935
rect -34 889 34 935
rect 80 889 91 935
rect -91 821 91 889
rect -91 775 -80 821
rect -34 775 34 821
rect 80 775 91 821
rect -91 707 91 775
rect -91 661 -80 707
rect -34 661 34 707
rect 80 661 91 707
rect -91 593 91 661
rect -91 547 -80 593
rect -34 547 34 593
rect 80 547 91 593
rect -91 479 91 547
rect -91 433 -80 479
rect -34 433 34 479
rect 80 433 91 479
rect -91 365 91 433
rect -91 319 -80 365
rect -34 319 34 365
rect 80 319 91 365
rect -91 251 91 319
rect -91 205 -80 251
rect -34 205 34 251
rect 80 205 91 251
rect -91 137 91 205
rect -91 91 -80 137
rect -34 91 34 137
rect 80 91 91 137
rect -91 23 91 91
rect -91 -23 -80 23
rect -34 -23 34 23
rect 80 -23 91 23
rect -91 -91 91 -23
rect -91 -137 -80 -91
rect -34 -137 34 -91
rect 80 -137 91 -91
rect -91 -205 91 -137
rect -91 -251 -80 -205
rect -34 -251 34 -205
rect 80 -251 91 -205
rect -91 -319 91 -251
rect -91 -365 -80 -319
rect -34 -365 34 -319
rect 80 -365 91 -319
rect -91 -433 91 -365
rect -91 -479 -80 -433
rect -34 -479 34 -433
rect 80 -479 91 -433
rect -91 -547 91 -479
rect -91 -593 -80 -547
rect -34 -593 34 -547
rect 80 -593 91 -547
rect -91 -661 91 -593
rect -91 -707 -80 -661
rect -34 -707 34 -661
rect 80 -707 91 -661
rect -91 -775 91 -707
rect -91 -821 -80 -775
rect -34 -821 34 -775
rect 80 -821 91 -775
rect -91 -889 91 -821
rect -91 -935 -80 -889
rect -34 -935 34 -889
rect 80 -935 91 -889
rect -91 -1003 91 -935
rect -91 -1049 -80 -1003
rect -34 -1049 34 -1003
rect 80 -1049 91 -1003
rect -91 -1117 91 -1049
rect -91 -1163 -80 -1117
rect -34 -1163 34 -1117
rect 80 -1163 91 -1117
rect -91 -1231 91 -1163
rect -91 -1277 -80 -1231
rect -34 -1277 34 -1231
rect 80 -1277 91 -1231
rect -91 -1345 91 -1277
rect -91 -1391 -80 -1345
rect -34 -1391 34 -1345
rect 80 -1391 91 -1345
rect -91 -1459 91 -1391
rect -91 -1505 -80 -1459
rect -34 -1505 34 -1459
rect 80 -1505 91 -1459
rect -91 -1573 91 -1505
rect -91 -1619 -80 -1573
rect -34 -1619 34 -1573
rect 80 -1619 91 -1573
rect -91 -1687 91 -1619
rect -91 -1733 -80 -1687
rect -34 -1733 34 -1687
rect 80 -1733 91 -1687
rect -91 -1801 91 -1733
rect -91 -1847 -80 -1801
rect -34 -1847 34 -1801
rect 80 -1847 91 -1801
rect -91 -1915 91 -1847
rect -91 -1961 -80 -1915
rect -34 -1961 34 -1915
rect 80 -1961 91 -1915
rect -91 -2029 91 -1961
rect -91 -2075 -80 -2029
rect -34 -2075 34 -2029
rect 80 -2075 91 -2029
rect -91 -2143 91 -2075
rect -91 -2189 -80 -2143
rect -34 -2189 34 -2143
rect 80 -2189 91 -2143
rect -91 -2257 91 -2189
rect -91 -2303 -80 -2257
rect -34 -2303 34 -2257
rect 80 -2303 91 -2257
rect -91 -2371 91 -2303
rect -91 -2417 -80 -2371
rect -34 -2417 34 -2371
rect 80 -2417 91 -2371
rect -91 -2485 91 -2417
rect -91 -2531 -80 -2485
rect -34 -2531 34 -2485
rect 80 -2531 91 -2485
rect -91 -2542 91 -2531
<< end >>
