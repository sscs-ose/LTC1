magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect 2904 -1968 12576 14320
<< psubdiff >>
rect 4904 12298 5263 12320
rect 4904 12252 4926 12298
rect 4972 12252 5040 12298
rect 5086 12252 5263 12298
rect 4904 12184 5263 12252
rect 4904 12138 4926 12184
rect 4972 12138 5040 12184
rect 5086 12138 5263 12184
rect 4904 12116 5263 12138
rect 10233 12116 10423 12320
rect 4904 12070 5108 12116
rect 4904 12024 4926 12070
rect 4972 12024 5040 12070
rect 5086 12024 5108 12070
rect 4904 11500 5108 12024
rect 4904 11454 4926 11500
rect 4972 11454 5040 11500
rect 5086 11454 5108 11500
rect 4904 11386 5108 11454
rect 4904 11340 4926 11386
rect 4972 11340 5040 11386
rect 5086 11340 5108 11386
rect 4904 11272 5108 11340
rect 4904 11226 4926 11272
rect 4972 11226 5040 11272
rect 5086 11226 5108 11272
rect 4904 11158 5108 11226
rect 4904 11112 4926 11158
rect 4972 11112 5040 11158
rect 5086 11112 5108 11158
rect 4904 11044 5108 11112
rect 4904 10998 4926 11044
rect 4972 10998 5040 11044
rect 5086 10998 5108 11044
rect 4904 10930 5108 10998
rect 4904 10884 4926 10930
rect 4972 10884 5040 10930
rect 5086 10884 5108 10930
rect 4904 10816 5108 10884
rect 4904 10770 4926 10816
rect 4972 10770 5040 10816
rect 5086 10770 5108 10816
rect 4904 10702 5108 10770
rect 4904 10656 4926 10702
rect 4972 10656 5040 10702
rect 5086 10656 5108 10702
rect 4904 10588 5108 10656
rect 4904 10542 4926 10588
rect 4972 10542 5040 10588
rect 5086 10542 5108 10588
rect 4904 10474 5108 10542
rect 4904 10428 4926 10474
rect 4972 10428 5040 10474
rect 5086 10428 5108 10474
rect 4904 10360 5108 10428
rect 4904 10314 4926 10360
rect 4972 10314 5040 10360
rect 5086 10314 5108 10360
rect 4904 10246 5108 10314
rect 4904 10200 4926 10246
rect 4972 10200 5040 10246
rect 5086 10200 5108 10246
rect 4904 10132 5108 10200
rect 4904 10086 4926 10132
rect 4972 10086 5040 10132
rect 5086 10086 5108 10132
rect 4904 10018 5108 10086
rect 4904 9972 4926 10018
rect 4972 9972 5040 10018
rect 5086 9972 5108 10018
rect 4904 9904 5108 9972
rect 4904 9858 4926 9904
rect 4972 9858 5040 9904
rect 5086 9858 5108 9904
rect 4904 9790 5108 9858
rect 4904 9744 4926 9790
rect 4972 9744 5040 9790
rect 5086 9744 5108 9790
rect 4904 9676 5108 9744
rect 4904 9630 4926 9676
rect 4972 9630 5040 9676
rect 5086 9630 5108 9676
rect 4904 9562 5108 9630
rect 4904 9516 4926 9562
rect 4972 9516 5040 9562
rect 5086 9516 5108 9562
rect 4904 9448 5108 9516
rect 4904 9402 4926 9448
rect 4972 9402 5040 9448
rect 5086 9402 5108 9448
rect 4904 9334 5108 9402
rect 4904 9288 4926 9334
rect 4972 9288 5040 9334
rect 5086 9288 5108 9334
rect 4904 9220 5108 9288
rect 4904 9174 4926 9220
rect 4972 9174 5040 9220
rect 5086 9174 5108 9220
rect 4904 9106 5108 9174
rect 4904 9060 4926 9106
rect 4972 9060 5040 9106
rect 5086 9060 5108 9106
rect 4904 8992 5108 9060
rect 4904 8946 4926 8992
rect 4972 8946 5040 8992
rect 5086 8946 5108 8992
rect 4904 8878 5108 8946
rect 4904 8832 4926 8878
rect 4972 8832 5040 8878
rect 5086 8832 5108 8878
rect 4904 8764 5108 8832
rect 4904 8718 4926 8764
rect 4972 8718 5040 8764
rect 5086 8718 5108 8764
rect 4904 8650 5108 8718
rect 4904 8604 4926 8650
rect 4972 8604 5040 8650
rect 5086 8604 5108 8650
rect 4904 8536 5108 8604
rect 4904 8490 4926 8536
rect 4972 8490 5040 8536
rect 5086 8490 5108 8536
rect 4904 8422 5108 8490
rect 4904 8376 4926 8422
rect 4972 8376 5040 8422
rect 5086 8376 5108 8422
rect 4904 8308 5108 8376
rect 4904 8262 4926 8308
rect 4972 8262 5040 8308
rect 5086 8262 5108 8308
rect 4904 8194 5108 8262
rect 4904 8148 4926 8194
rect 4972 8148 5040 8194
rect 5086 8148 5108 8194
rect 4904 8080 5108 8148
rect 4904 8034 4926 8080
rect 4972 8034 5040 8080
rect 5086 8034 5108 8080
rect 4904 7966 5108 8034
rect 4904 7920 4926 7966
rect 4972 7920 5040 7966
rect 5086 7920 5108 7966
rect 4904 7852 5108 7920
rect 4904 7806 4926 7852
rect 4972 7806 5040 7852
rect 5086 7806 5108 7852
rect 4904 7738 5108 7806
rect 4904 7692 4926 7738
rect 4972 7692 5040 7738
rect 5086 7692 5108 7738
rect 4904 7624 5108 7692
rect 4904 7578 4926 7624
rect 4972 7578 5040 7624
rect 5086 7578 5108 7624
rect 4904 7510 5108 7578
rect 4904 7464 4926 7510
rect 4972 7464 5040 7510
rect 5086 7464 5108 7510
rect 4904 7396 5108 7464
rect 4904 7350 4926 7396
rect 4972 7350 5040 7396
rect 5086 7350 5108 7396
rect 4904 7282 5108 7350
rect 4904 7236 4926 7282
rect 4972 7236 5040 7282
rect 5086 7236 5108 7282
rect 4904 7168 5108 7236
rect 4904 7122 4926 7168
rect 4972 7122 5040 7168
rect 5086 7122 5108 7168
rect 4904 7054 5108 7122
rect 4904 7008 4926 7054
rect 4972 7008 5040 7054
rect 5086 7008 5108 7054
rect 4904 6940 5108 7008
rect 4904 6894 4926 6940
rect 4972 6894 5040 6940
rect 5086 6894 5108 6940
rect 4904 6826 5108 6894
rect 4904 6780 4926 6826
rect 4972 6780 5040 6826
rect 5086 6780 5108 6826
rect 4904 6712 5108 6780
rect 4904 6666 4926 6712
rect 4972 6666 5040 6712
rect 5086 6666 5108 6712
rect 4904 6598 5108 6666
rect 4904 6552 4926 6598
rect 4972 6552 5040 6598
rect 5086 6552 5108 6598
rect 4904 6484 5108 6552
rect 4904 6438 4926 6484
rect 4972 6438 5040 6484
rect 5086 6438 5108 6484
rect 4904 6370 5108 6438
rect 4904 6324 4926 6370
rect 4972 6324 5040 6370
rect 5086 6324 5108 6370
rect 4904 6256 5108 6324
rect 4904 6210 4926 6256
rect 4972 6210 5040 6256
rect 5086 6229 5108 6256
rect 5086 6210 5206 6229
rect 4904 6142 5206 6210
rect 4904 6096 4926 6142
rect 4972 6096 5040 6142
rect 5086 6096 5206 6142
rect 4904 6028 5206 6096
rect 4904 5982 4926 6028
rect 4972 5982 5040 6028
rect 5086 6025 5206 6028
rect 10294 6025 10372 6229
rect 5086 5982 5108 6025
rect 4904 5914 5108 5982
rect 4904 5868 4926 5914
rect 4972 5868 5040 5914
rect 5086 5868 5108 5914
rect 4904 5800 5108 5868
rect 4904 5754 4926 5800
rect 4972 5754 5040 5800
rect 5086 5754 5108 5800
rect 4904 5686 5108 5754
rect 4904 5640 4926 5686
rect 4972 5640 5040 5686
rect 5086 5640 5108 5686
rect 4904 5572 5108 5640
rect 4904 5526 4926 5572
rect 4972 5526 5040 5572
rect 5086 5526 5108 5572
rect 4904 5458 5108 5526
rect 4904 5412 4926 5458
rect 4972 5412 5040 5458
rect 5086 5412 5108 5458
rect 4904 5344 5108 5412
rect 4904 5298 4926 5344
rect 4972 5298 5040 5344
rect 5086 5298 5108 5344
rect 4904 5230 5108 5298
rect 4904 5184 4926 5230
rect 4972 5184 5040 5230
rect 5086 5184 5108 5230
rect 4904 5116 5108 5184
rect 4904 5070 4926 5116
rect 4972 5070 5040 5116
rect 5086 5070 5108 5116
rect 4904 5002 5108 5070
rect 4904 4956 4926 5002
rect 4972 4956 5040 5002
rect 5086 4956 5108 5002
rect 4904 4888 5108 4956
rect 4904 4842 4926 4888
rect 4972 4842 5040 4888
rect 5086 4842 5108 4888
rect 4904 4774 5108 4842
rect 4904 4728 4926 4774
rect 4972 4728 5040 4774
rect 5086 4728 5108 4774
rect 4904 4660 5108 4728
rect 4904 4614 4926 4660
rect 4972 4614 5040 4660
rect 5086 4614 5108 4660
rect 4904 4546 5108 4614
rect 4904 4500 4926 4546
rect 4972 4500 5040 4546
rect 5086 4500 5108 4546
rect 4904 4432 5108 4500
rect 4904 4386 4926 4432
rect 4972 4386 5040 4432
rect 5086 4386 5108 4432
rect 4904 4318 5108 4386
rect 4904 4272 4926 4318
rect 4972 4272 5040 4318
rect 5086 4272 5108 4318
rect 4904 4204 5108 4272
rect 4904 4158 4926 4204
rect 4972 4158 5040 4204
rect 5086 4158 5108 4204
rect 4904 4090 5108 4158
rect 4904 4044 4926 4090
rect 4972 4044 5040 4090
rect 5086 4044 5108 4090
rect 4904 3976 5108 4044
rect 4904 3930 4926 3976
rect 4972 3930 5040 3976
rect 5086 3930 5108 3976
rect 4904 3862 5108 3930
rect 4904 3816 4926 3862
rect 4972 3816 5040 3862
rect 5086 3816 5108 3862
rect 4904 3748 5108 3816
rect 4904 3702 4926 3748
rect 4972 3702 5040 3748
rect 5086 3702 5108 3748
rect 4904 3634 5108 3702
rect 4904 3588 4926 3634
rect 4972 3588 5040 3634
rect 5086 3588 5108 3634
rect 4904 3520 5108 3588
rect 4904 3474 4926 3520
rect 4972 3474 5040 3520
rect 5086 3474 5108 3520
rect 4904 3406 5108 3474
rect 4904 3360 4926 3406
rect 4972 3360 5040 3406
rect 5086 3360 5108 3406
rect 4904 3292 5108 3360
rect 4904 3246 4926 3292
rect 4972 3246 5040 3292
rect 5086 3246 5108 3292
rect 4904 3178 5108 3246
rect 4904 3132 4926 3178
rect 4972 3132 5040 3178
rect 5086 3132 5108 3178
rect 4904 3064 5108 3132
rect 4904 3018 4926 3064
rect 4972 3018 5040 3064
rect 5086 3018 5108 3064
rect 4904 2950 5108 3018
rect 4904 2904 4926 2950
rect 4972 2904 5040 2950
rect 5086 2904 5108 2950
rect 4904 2836 5108 2904
rect 4904 2790 4926 2836
rect 4972 2790 5040 2836
rect 5086 2790 5108 2836
rect 4904 2722 5108 2790
rect 4904 2676 4926 2722
rect 4972 2676 5040 2722
rect 5086 2676 5108 2722
rect 4904 2608 5108 2676
rect 4904 2562 4926 2608
rect 4972 2562 5040 2608
rect 5086 2562 5108 2608
rect 4904 2494 5108 2562
rect 4904 2448 4926 2494
rect 4972 2448 5040 2494
rect 5086 2448 5108 2494
rect 4904 2380 5108 2448
rect 4904 2334 4926 2380
rect 4972 2334 5040 2380
rect 5086 2334 5108 2380
rect 4904 2266 5108 2334
rect 4904 2220 4926 2266
rect 4972 2220 5040 2266
rect 5086 2220 5108 2266
rect 4904 2152 5108 2220
rect 4904 2106 4926 2152
rect 4972 2106 5040 2152
rect 5086 2106 5108 2152
rect 4904 2038 5108 2106
rect 4904 1992 4926 2038
rect 4972 1992 5040 2038
rect 5086 1992 5108 2038
rect 4904 1924 5108 1992
rect 4904 1878 4926 1924
rect 4972 1878 5040 1924
rect 5086 1878 5108 1924
rect 4904 1810 5108 1878
rect 4904 1764 4926 1810
rect 4972 1764 5040 1810
rect 5086 1764 5108 1810
rect 4904 1696 5108 1764
rect 4904 1650 4926 1696
rect 4972 1650 5040 1696
rect 5086 1650 5108 1696
rect 4904 1582 5108 1650
rect 4904 1536 4926 1582
rect 4972 1536 5040 1582
rect 5086 1536 5108 1582
rect 4904 1468 5108 1536
rect 4904 1422 4926 1468
rect 4972 1422 5040 1468
rect 5086 1422 5108 1468
rect 4904 1354 5108 1422
rect 4904 1308 4926 1354
rect 4972 1308 5040 1354
rect 5086 1308 5108 1354
rect 4904 1240 5108 1308
rect 4904 1194 4926 1240
rect 4972 1194 5040 1240
rect 5086 1194 5108 1240
rect 4904 1126 5108 1194
rect 4904 1080 4926 1126
rect 4972 1080 5040 1126
rect 5086 1080 5108 1126
rect 4904 1012 5108 1080
rect 4904 966 4926 1012
rect 4972 966 5040 1012
rect 5086 966 5108 1012
rect 4904 898 5108 966
rect 4904 852 4926 898
rect 4972 852 5040 898
rect 5086 852 5108 898
rect 4904 784 5108 852
rect 4904 738 4926 784
rect 4972 738 5040 784
rect 5086 738 5108 784
rect 4904 328 5108 738
rect 4904 282 4926 328
rect 4972 282 5040 328
rect 5086 282 5108 328
rect 4904 236 5108 282
rect 4904 214 10423 236
rect 4904 168 4926 214
rect 4972 168 5040 214
rect 5086 168 10423 214
rect 4904 100 10423 168
rect 4904 54 4926 100
rect 4972 54 5040 100
rect 5086 54 10423 100
rect 4904 32 10423 54
<< psubdiffcont >>
rect 4926 12252 4972 12298
rect 5040 12252 5086 12298
rect 4926 12138 4972 12184
rect 5040 12138 5086 12184
rect 4926 12024 4972 12070
rect 5040 12024 5086 12070
rect 4926 11454 4972 11500
rect 5040 11454 5086 11500
rect 4926 11340 4972 11386
rect 5040 11340 5086 11386
rect 4926 11226 4972 11272
rect 5040 11226 5086 11272
rect 4926 11112 4972 11158
rect 5040 11112 5086 11158
rect 4926 10998 4972 11044
rect 5040 10998 5086 11044
rect 4926 10884 4972 10930
rect 5040 10884 5086 10930
rect 4926 10770 4972 10816
rect 5040 10770 5086 10816
rect 4926 10656 4972 10702
rect 5040 10656 5086 10702
rect 4926 10542 4972 10588
rect 5040 10542 5086 10588
rect 4926 10428 4972 10474
rect 5040 10428 5086 10474
rect 4926 10314 4972 10360
rect 5040 10314 5086 10360
rect 4926 10200 4972 10246
rect 5040 10200 5086 10246
rect 4926 10086 4972 10132
rect 5040 10086 5086 10132
rect 4926 9972 4972 10018
rect 5040 9972 5086 10018
rect 4926 9858 4972 9904
rect 5040 9858 5086 9904
rect 4926 9744 4972 9790
rect 5040 9744 5086 9790
rect 4926 9630 4972 9676
rect 5040 9630 5086 9676
rect 4926 9516 4972 9562
rect 5040 9516 5086 9562
rect 4926 9402 4972 9448
rect 5040 9402 5086 9448
rect 4926 9288 4972 9334
rect 5040 9288 5086 9334
rect 4926 9174 4972 9220
rect 5040 9174 5086 9220
rect 4926 9060 4972 9106
rect 5040 9060 5086 9106
rect 4926 8946 4972 8992
rect 5040 8946 5086 8992
rect 4926 8832 4972 8878
rect 5040 8832 5086 8878
rect 4926 8718 4972 8764
rect 5040 8718 5086 8764
rect 4926 8604 4972 8650
rect 5040 8604 5086 8650
rect 4926 8490 4972 8536
rect 5040 8490 5086 8536
rect 4926 8376 4972 8422
rect 5040 8376 5086 8422
rect 4926 8262 4972 8308
rect 5040 8262 5086 8308
rect 4926 8148 4972 8194
rect 5040 8148 5086 8194
rect 4926 8034 4972 8080
rect 5040 8034 5086 8080
rect 4926 7920 4972 7966
rect 5040 7920 5086 7966
rect 4926 7806 4972 7852
rect 5040 7806 5086 7852
rect 4926 7692 4972 7738
rect 5040 7692 5086 7738
rect 4926 7578 4972 7624
rect 5040 7578 5086 7624
rect 4926 7464 4972 7510
rect 5040 7464 5086 7510
rect 4926 7350 4972 7396
rect 5040 7350 5086 7396
rect 4926 7236 4972 7282
rect 5040 7236 5086 7282
rect 4926 7122 4972 7168
rect 5040 7122 5086 7168
rect 4926 7008 4972 7054
rect 5040 7008 5086 7054
rect 4926 6894 4972 6940
rect 5040 6894 5086 6940
rect 4926 6780 4972 6826
rect 5040 6780 5086 6826
rect 4926 6666 4972 6712
rect 5040 6666 5086 6712
rect 4926 6552 4972 6598
rect 5040 6552 5086 6598
rect 4926 6438 4972 6484
rect 5040 6438 5086 6484
rect 4926 6324 4972 6370
rect 5040 6324 5086 6370
rect 4926 6210 4972 6256
rect 5040 6210 5086 6256
rect 4926 6096 4972 6142
rect 5040 6096 5086 6142
rect 4926 5982 4972 6028
rect 5040 5982 5086 6028
rect 4926 5868 4972 5914
rect 5040 5868 5086 5914
rect 4926 5754 4972 5800
rect 5040 5754 5086 5800
rect 4926 5640 4972 5686
rect 5040 5640 5086 5686
rect 4926 5526 4972 5572
rect 5040 5526 5086 5572
rect 4926 5412 4972 5458
rect 5040 5412 5086 5458
rect 4926 5298 4972 5344
rect 5040 5298 5086 5344
rect 4926 5184 4972 5230
rect 5040 5184 5086 5230
rect 4926 5070 4972 5116
rect 5040 5070 5086 5116
rect 4926 4956 4972 5002
rect 5040 4956 5086 5002
rect 4926 4842 4972 4888
rect 5040 4842 5086 4888
rect 4926 4728 4972 4774
rect 5040 4728 5086 4774
rect 4926 4614 4972 4660
rect 5040 4614 5086 4660
rect 4926 4500 4972 4546
rect 5040 4500 5086 4546
rect 4926 4386 4972 4432
rect 5040 4386 5086 4432
rect 4926 4272 4972 4318
rect 5040 4272 5086 4318
rect 4926 4158 4972 4204
rect 5040 4158 5086 4204
rect 4926 4044 4972 4090
rect 5040 4044 5086 4090
rect 4926 3930 4972 3976
rect 5040 3930 5086 3976
rect 4926 3816 4972 3862
rect 5040 3816 5086 3862
rect 4926 3702 4972 3748
rect 5040 3702 5086 3748
rect 4926 3588 4972 3634
rect 5040 3588 5086 3634
rect 4926 3474 4972 3520
rect 5040 3474 5086 3520
rect 4926 3360 4972 3406
rect 5040 3360 5086 3406
rect 4926 3246 4972 3292
rect 5040 3246 5086 3292
rect 4926 3132 4972 3178
rect 5040 3132 5086 3178
rect 4926 3018 4972 3064
rect 5040 3018 5086 3064
rect 4926 2904 4972 2950
rect 5040 2904 5086 2950
rect 4926 2790 4972 2836
rect 5040 2790 5086 2836
rect 4926 2676 4972 2722
rect 5040 2676 5086 2722
rect 4926 2562 4972 2608
rect 5040 2562 5086 2608
rect 4926 2448 4972 2494
rect 5040 2448 5086 2494
rect 4926 2334 4972 2380
rect 5040 2334 5086 2380
rect 4926 2220 4972 2266
rect 5040 2220 5086 2266
rect 4926 2106 4972 2152
rect 5040 2106 5086 2152
rect 4926 1992 4972 2038
rect 5040 1992 5086 2038
rect 4926 1878 4972 1924
rect 5040 1878 5086 1924
rect 4926 1764 4972 1810
rect 5040 1764 5086 1810
rect 4926 1650 4972 1696
rect 5040 1650 5086 1696
rect 4926 1536 4972 1582
rect 5040 1536 5086 1582
rect 4926 1422 4972 1468
rect 5040 1422 5086 1468
rect 4926 1308 4972 1354
rect 5040 1308 5086 1354
rect 4926 1194 4972 1240
rect 5040 1194 5086 1240
rect 4926 1080 4972 1126
rect 5040 1080 5086 1126
rect 4926 966 4972 1012
rect 5040 966 5086 1012
rect 4926 852 4972 898
rect 5040 852 5086 898
rect 4926 738 4972 784
rect 5040 738 5086 784
rect 4926 282 4972 328
rect 5040 282 5086 328
rect 4926 168 4972 214
rect 5040 168 5086 214
rect 4926 54 4972 100
rect 5040 54 5086 100
<< metal1 >>
rect 4915 12298 10565 12310
rect 4915 12252 4926 12298
rect 4972 12252 5040 12298
rect 5086 12252 10565 12298
rect 4915 12184 10565 12252
rect 4915 12138 4926 12184
rect 4972 12138 5040 12184
rect 5086 12138 10565 12184
rect 4915 12126 10565 12138
rect 4915 12070 5097 12126
rect 4915 12024 4926 12070
rect 4972 12024 5040 12070
rect 5086 12024 5097 12070
rect 4915 11633 5097 12024
rect 5561 11723 9913 11855
rect 5561 11655 7477 11723
rect 7997 11655 9913 11723
rect 4915 11500 5301 11633
rect 4915 11454 4926 11500
rect 4972 11454 5040 11500
rect 5086 11454 5301 11500
rect 4915 11386 5301 11454
rect 4915 11340 4926 11386
rect 4972 11340 5040 11386
rect 5086 11340 5301 11386
rect 4915 11272 5301 11340
rect 4915 11226 4926 11272
rect 4972 11226 5040 11272
rect 5086 11226 5301 11272
rect 4915 11158 5301 11226
rect 4915 11112 4926 11158
rect 4972 11112 5040 11158
rect 5086 11112 5301 11158
rect 4915 11044 5301 11112
rect 4915 10998 4926 11044
rect 4972 10998 5040 11044
rect 5086 10998 5301 11044
rect 4915 10930 5301 10998
rect 4915 10884 4926 10930
rect 4972 10884 5040 10930
rect 5086 10884 5301 10930
rect 4915 10816 5301 10884
rect 4915 10770 4926 10816
rect 4972 10770 5040 10816
rect 5086 10770 5301 10816
rect 4915 10702 5301 10770
rect 4915 10656 4926 10702
rect 4972 10656 5040 10702
rect 5086 10656 5301 10702
rect 4915 10588 5301 10656
rect 4915 10542 4926 10588
rect 4972 10542 5040 10588
rect 5086 10542 5301 10588
rect 4915 10474 5301 10542
rect 4915 10428 4926 10474
rect 4972 10428 5040 10474
rect 5086 10428 5301 10474
rect 4915 10360 5301 10428
rect 4915 10314 4926 10360
rect 4972 10314 5040 10360
rect 5086 10314 5301 10360
rect 4915 10246 5301 10314
rect 4915 10200 4926 10246
rect 4972 10200 5040 10246
rect 5086 10200 5301 10246
rect 4915 10132 5301 10200
rect 4915 10086 4926 10132
rect 4972 10086 5040 10132
rect 5086 10086 5301 10132
rect 4915 10018 5301 10086
rect 4915 9972 4926 10018
rect 4972 9972 5040 10018
rect 5086 9972 5301 10018
rect 4915 9904 5301 9972
rect 4915 9858 4926 9904
rect 4972 9858 5040 9904
rect 5086 9858 5301 9904
rect 4915 9790 5301 9858
rect 4915 9744 4926 9790
rect 4972 9744 5040 9790
rect 5086 9744 5301 9790
rect 4915 9676 5301 9744
rect 4915 9630 4926 9676
rect 4972 9630 5040 9676
rect 5086 9630 5301 9676
rect 4915 9562 5301 9630
rect 4915 9516 4926 9562
rect 4972 9516 5040 9562
rect 5086 9516 5301 9562
rect 4915 9448 5301 9516
rect 4915 9402 4926 9448
rect 4972 9402 5040 9448
rect 5086 9402 5301 9448
rect 4915 9334 5301 9402
rect 4915 9288 4926 9334
rect 4972 9288 5040 9334
rect 5086 9288 5301 9334
rect 4915 9220 5301 9288
rect 4915 9174 4926 9220
rect 4972 9174 5040 9220
rect 5086 9174 5301 9220
rect 4915 9106 5301 9174
rect 4915 9060 4926 9106
rect 4972 9060 5040 9106
rect 5086 9060 5301 9106
rect 4915 8992 5301 9060
rect 4915 8946 4926 8992
rect 4972 8946 5040 8992
rect 5086 8946 5301 8992
rect 4915 8878 5301 8946
rect 4915 8832 4926 8878
rect 4972 8832 5040 8878
rect 5086 8832 5301 8878
rect 4915 8764 5301 8832
rect 4915 8718 4926 8764
rect 4972 8718 5040 8764
rect 5086 8718 5301 8764
rect 4915 8650 5301 8718
rect 4915 8604 4926 8650
rect 4972 8604 5040 8650
rect 5086 8604 5301 8650
rect 4915 8536 5301 8604
rect 4915 8490 4926 8536
rect 4972 8490 5040 8536
rect 5086 8490 5301 8536
rect 4915 8422 5301 8490
rect 4915 8376 4926 8422
rect 4972 8376 5040 8422
rect 5086 8376 5301 8422
rect 4915 8308 5301 8376
rect 4915 8262 4926 8308
rect 4972 8262 5040 8308
rect 5086 8262 5301 8308
rect 4915 8194 5301 8262
rect 4915 8148 4926 8194
rect 4972 8148 5040 8194
rect 5086 8148 5301 8194
rect 4915 8080 5301 8148
rect 4915 8034 4926 8080
rect 4972 8034 5040 8080
rect 5086 8034 5301 8080
rect 4915 7966 5301 8034
rect 4915 7920 4926 7966
rect 4972 7920 5040 7966
rect 5086 7920 5301 7966
rect 4915 7852 5301 7920
rect 4915 7806 4926 7852
rect 4972 7806 5040 7852
rect 5086 7806 5301 7852
rect 4915 7738 5301 7806
rect 4915 7692 4926 7738
rect 4972 7692 5040 7738
rect 5086 7692 5301 7738
rect 4915 7624 5301 7692
rect 4915 7578 4926 7624
rect 4972 7578 5040 7624
rect 5086 7578 5301 7624
rect 4915 7510 5301 7578
rect 4915 7464 4926 7510
rect 4972 7464 5040 7510
rect 5086 7464 5301 7510
rect 4915 7396 5301 7464
rect 4915 7350 4926 7396
rect 4972 7350 5040 7396
rect 5086 7350 5301 7396
rect 4915 7282 5301 7350
rect 4915 7236 4926 7282
rect 4972 7236 5040 7282
rect 5086 7236 5301 7282
rect 4915 7168 5301 7236
rect 4915 7122 4926 7168
rect 4972 7122 5040 7168
rect 5086 7122 5301 7168
rect 4915 7054 5301 7122
rect 4915 7008 4926 7054
rect 4972 7008 5040 7054
rect 5086 7008 5301 7054
rect 4915 6940 5301 7008
rect 4915 6894 4926 6940
rect 4972 6894 5040 6940
rect 5086 6894 5301 6940
rect 4915 6826 5301 6894
rect 4915 6780 4926 6826
rect 4972 6780 5040 6826
rect 5086 6780 5301 6826
rect 4915 6712 5301 6780
rect 4915 6666 4926 6712
rect 4972 6666 5040 6712
rect 5086 6666 5301 6712
rect 4915 6598 5301 6666
rect 4915 6552 4926 6598
rect 4972 6552 5040 6598
rect 5086 6552 5301 6598
rect 4915 6484 5301 6552
rect 4915 6438 4926 6484
rect 4972 6438 5040 6484
rect 5086 6483 5301 6484
rect 10173 6483 10383 11633
rect 5086 6438 10383 6483
rect 4915 6370 10383 6438
rect 4915 6324 4926 6370
rect 4972 6324 5040 6370
rect 5086 6324 10383 6370
rect 4915 6256 10383 6324
rect 4915 6210 4926 6256
rect 4972 6210 5040 6256
rect 5086 6210 10383 6256
rect 4915 6142 10383 6210
rect 4915 6096 4926 6142
rect 4972 6096 5040 6142
rect 5086 6096 10383 6142
rect 4915 6028 10383 6096
rect 4915 5982 4926 6028
rect 4972 5982 5040 6028
rect 5086 5982 10383 6028
rect 4915 5914 10383 5982
rect 4915 5868 4926 5914
rect 4972 5868 5040 5914
rect 5086 5868 10383 5914
rect 4915 5800 10383 5868
rect 4915 5754 4926 5800
rect 4972 5754 5040 5800
rect 5086 5771 10383 5800
rect 5086 5754 5301 5771
rect 4915 5686 5301 5754
rect 4915 5640 4926 5686
rect 4972 5640 5040 5686
rect 5086 5640 5301 5686
rect 4915 5572 5301 5640
rect 4915 5526 4926 5572
rect 4972 5526 5040 5572
rect 5086 5526 5301 5572
rect 4915 5458 5301 5526
rect 4915 5412 4926 5458
rect 4972 5412 5040 5458
rect 5086 5412 5301 5458
rect 4915 5344 5301 5412
rect 4915 5298 4926 5344
rect 4972 5298 5040 5344
rect 5086 5298 5301 5344
rect 4915 5230 5301 5298
rect 4915 5184 4926 5230
rect 4972 5184 5040 5230
rect 5086 5184 5301 5230
rect 4915 5116 5301 5184
rect 4915 5070 4926 5116
rect 4972 5070 5040 5116
rect 5086 5070 5301 5116
rect 4915 5002 5301 5070
rect 4915 4956 4926 5002
rect 4972 4956 5040 5002
rect 5086 4956 5301 5002
rect 4915 4888 5301 4956
rect 4915 4842 4926 4888
rect 4972 4842 5040 4888
rect 5086 4842 5301 4888
rect 4915 4774 5301 4842
rect 4915 4728 4926 4774
rect 4972 4728 5040 4774
rect 5086 4728 5301 4774
rect 4915 4660 5301 4728
rect 4915 4614 4926 4660
rect 4972 4614 5040 4660
rect 5086 4614 5301 4660
rect 4915 4546 5301 4614
rect 4915 4500 4926 4546
rect 4972 4500 5040 4546
rect 5086 4500 5301 4546
rect 4915 4432 5301 4500
rect 4915 4386 4926 4432
rect 4972 4386 5040 4432
rect 5086 4386 5301 4432
rect 4915 4318 5301 4386
rect 4915 4272 4926 4318
rect 4972 4272 5040 4318
rect 5086 4272 5301 4318
rect 4915 4204 5301 4272
rect 4915 4158 4926 4204
rect 4972 4158 5040 4204
rect 5086 4158 5301 4204
rect 4915 4090 5301 4158
rect 4915 4044 4926 4090
rect 4972 4044 5040 4090
rect 5086 4044 5301 4090
rect 4915 3976 5301 4044
rect 4915 3930 4926 3976
rect 4972 3930 5040 3976
rect 5086 3930 5301 3976
rect 4915 3862 5301 3930
rect 4915 3816 4926 3862
rect 4972 3816 5040 3862
rect 5086 3816 5301 3862
rect 4915 3748 5301 3816
rect 4915 3702 4926 3748
rect 4972 3702 5040 3748
rect 5086 3702 5301 3748
rect 4915 3634 5301 3702
rect 4915 3588 4926 3634
rect 4972 3588 5040 3634
rect 5086 3588 5301 3634
rect 4915 3520 5301 3588
rect 4915 3474 4926 3520
rect 4972 3474 5040 3520
rect 5086 3474 5301 3520
rect 4915 3406 5301 3474
rect 4915 3360 4926 3406
rect 4972 3360 5040 3406
rect 5086 3360 5301 3406
rect 4915 3292 5301 3360
rect 4915 3246 4926 3292
rect 4972 3246 5040 3292
rect 5086 3246 5301 3292
rect 4915 3178 5301 3246
rect 4915 3132 4926 3178
rect 4972 3132 5040 3178
rect 5086 3132 5301 3178
rect 4915 3064 5301 3132
rect 4915 3018 4926 3064
rect 4972 3018 5040 3064
rect 5086 3018 5301 3064
rect 4915 2950 5301 3018
rect 4915 2904 4926 2950
rect 4972 2904 5040 2950
rect 5086 2904 5301 2950
rect 4915 2836 5301 2904
rect 4915 2790 4926 2836
rect 4972 2790 5040 2836
rect 5086 2790 5301 2836
rect 4915 2722 5301 2790
rect 4915 2676 4926 2722
rect 4972 2676 5040 2722
rect 5086 2676 5301 2722
rect 4915 2608 5301 2676
rect 4915 2562 4926 2608
rect 4972 2562 5040 2608
rect 5086 2562 5301 2608
rect 4915 2494 5301 2562
rect 4915 2448 4926 2494
rect 4972 2448 5040 2494
rect 5086 2448 5301 2494
rect 4915 2380 5301 2448
rect 4915 2334 4926 2380
rect 4972 2334 5040 2380
rect 5086 2334 5301 2380
rect 4915 2266 5301 2334
rect 4915 2220 4926 2266
rect 4972 2220 5040 2266
rect 5086 2220 5301 2266
rect 4915 2152 5301 2220
rect 4915 2106 4926 2152
rect 4972 2106 5040 2152
rect 5086 2106 5301 2152
rect 4915 2038 5301 2106
rect 4915 1992 4926 2038
rect 4972 1992 5040 2038
rect 5086 1992 5301 2038
rect 4915 1924 5301 1992
rect 4915 1878 4926 1924
rect 4972 1878 5040 1924
rect 5086 1878 5301 1924
rect 4915 1810 5301 1878
rect 4915 1764 4926 1810
rect 4972 1764 5040 1810
rect 5086 1764 5301 1810
rect 4915 1696 5301 1764
rect 4915 1650 4926 1696
rect 4972 1650 5040 1696
rect 5086 1650 5301 1696
rect 4915 1582 5301 1650
rect 4915 1536 4926 1582
rect 4972 1536 5040 1582
rect 5086 1536 5301 1582
rect 4915 1468 5301 1536
rect 4915 1422 4926 1468
rect 4972 1422 5040 1468
rect 5086 1422 5301 1468
rect 4915 1354 5301 1422
rect 4915 1308 4926 1354
rect 4972 1308 5040 1354
rect 5086 1308 5301 1354
rect 4915 1240 5301 1308
rect 4915 1194 4926 1240
rect 4972 1194 5040 1240
rect 5086 1194 5301 1240
rect 4915 1126 5301 1194
rect 4915 1080 4926 1126
rect 4972 1080 5040 1126
rect 5086 1080 5301 1126
rect 4915 1012 5301 1080
rect 4915 966 4926 1012
rect 4972 966 5040 1012
rect 5086 966 5301 1012
rect 4915 898 5301 966
rect 4915 852 4926 898
rect 4972 852 5040 898
rect 5086 852 5301 898
rect 4915 784 5301 852
rect 4915 738 4926 784
rect 4972 738 5040 784
rect 5086 738 5301 784
rect 4915 621 5301 738
rect 10173 621 10383 5771
rect 4915 328 5097 621
rect 5561 531 7477 599
rect 7997 531 9913 599
rect 5561 399 9913 531
rect 4915 282 4926 328
rect 4972 282 5040 328
rect 5086 282 5097 328
rect 4915 226 5097 282
rect 4915 214 10565 226
rect 4915 168 4926 214
rect 4972 168 5040 214
rect 5086 168 10565 214
rect 4915 100 10565 168
rect 4915 54 4926 100
rect 4972 54 5040 100
rect 5086 54 10565 100
rect 4915 42 10565 54
use M1_PSUB_CDNS_69033583165351  M1_PSUB_CDNS_69033583165351_0
timestamp 1713338890
transform 1 0 10474 0 1 6176
box -102 -6144 102 6144
use M1_PSUB_CDNS_69033583165486  M1_PSUB_CDNS_69033583165486_0
timestamp 1713338890
transform 0 -1 7753 1 0 134
box -102 -2553 102 2553
use M1_PSUB_CDNS_69033583165486  M1_PSUB_CDNS_69033583165486_1
timestamp 1713338890
transform 0 -1 7745 1 0 6127
box -102 -2553 102 2553
use M1_PSUB_CDNS_69033583165486  M1_PSUB_CDNS_69033583165486_2
timestamp 1713338890
transform 0 -1 7748 1 0 12218
box -102 -2553 102 2553
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_0
timestamp 1713338890
transform 1 0 5519 0 1 6633
box -218 -350 2218 5092
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_1
timestamp 1713338890
transform 1 0 7955 0 1 6633
box -218 -350 2218 5092
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_2
timestamp 1713338890
transform 1 0 5519 0 -1 5621
box -218 -350 2218 5092
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_3
timestamp 1713338890
transform 1 0 7955 0 -1 5621
box -218 -350 2218 5092
<< end >>
