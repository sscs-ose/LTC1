magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1748 1019 1748
<< metal2 >>
rect -19 742 19 748
rect -19 -742 -14 742
rect 14 -742 19 742
rect -19 -748 19 -742
<< via2 >>
rect -14 -742 14 742
<< metal3 >>
rect -19 742 19 748
rect -19 -742 -14 742
rect 14 -742 19 742
rect -19 -748 19 -742
<< end >>
