magic
tech gf180mcuC
magscale 1 10
timestamp 1714126980
<< error_p >>
rect -2063 -38 -2017 38
rect -1859 -38 -1813 38
rect -1655 -38 -1609 38
rect -1451 -38 -1405 38
rect -1247 -38 -1201 38
rect -1043 -38 -997 38
rect -839 -38 -793 38
rect -635 -38 -589 38
rect -431 -38 -385 38
rect -227 -38 -181 38
rect -23 -38 23 38
rect 181 -38 227 38
rect 385 -38 431 38
rect 589 -38 635 38
rect 793 -38 839 38
rect 997 -38 1043 38
rect 1201 -38 1247 38
rect 1405 -38 1451 38
rect 1609 -38 1655 38
rect 1813 -38 1859 38
rect 2017 -38 2063 38
<< nwell >>
rect -2162 -170 2162 170
<< pmos >>
rect -1988 -40 -1888 40
rect -1784 -40 -1684 40
rect -1580 -40 -1480 40
rect -1376 -40 -1276 40
rect -1172 -40 -1072 40
rect -968 -40 -868 40
rect -764 -40 -664 40
rect -560 -40 -460 40
rect -356 -40 -256 40
rect -152 -40 -52 40
rect 52 -40 152 40
rect 256 -40 356 40
rect 460 -40 560 40
rect 664 -40 764 40
rect 868 -40 968 40
rect 1072 -40 1172 40
rect 1276 -40 1376 40
rect 1480 -40 1580 40
rect 1684 -40 1784 40
rect 1888 -40 1988 40
<< pdiff >>
rect -2076 27 -1988 40
rect -2076 -27 -2063 27
rect -2017 -27 -1988 27
rect -2076 -40 -1988 -27
rect -1888 27 -1784 40
rect -1888 -27 -1859 27
rect -1813 -27 -1784 27
rect -1888 -40 -1784 -27
rect -1684 27 -1580 40
rect -1684 -27 -1655 27
rect -1609 -27 -1580 27
rect -1684 -40 -1580 -27
rect -1480 27 -1376 40
rect -1480 -27 -1451 27
rect -1405 -27 -1376 27
rect -1480 -40 -1376 -27
rect -1276 27 -1172 40
rect -1276 -27 -1247 27
rect -1201 -27 -1172 27
rect -1276 -40 -1172 -27
rect -1072 27 -968 40
rect -1072 -27 -1043 27
rect -997 -27 -968 27
rect -1072 -40 -968 -27
rect -868 27 -764 40
rect -868 -27 -839 27
rect -793 -27 -764 27
rect -868 -40 -764 -27
rect -664 27 -560 40
rect -664 -27 -635 27
rect -589 -27 -560 27
rect -664 -40 -560 -27
rect -460 27 -356 40
rect -460 -27 -431 27
rect -385 -27 -356 27
rect -460 -40 -356 -27
rect -256 27 -152 40
rect -256 -27 -227 27
rect -181 -27 -152 27
rect -256 -40 -152 -27
rect -52 27 52 40
rect -52 -27 -23 27
rect 23 -27 52 27
rect -52 -40 52 -27
rect 152 27 256 40
rect 152 -27 181 27
rect 227 -27 256 27
rect 152 -40 256 -27
rect 356 27 460 40
rect 356 -27 385 27
rect 431 -27 460 27
rect 356 -40 460 -27
rect 560 27 664 40
rect 560 -27 589 27
rect 635 -27 664 27
rect 560 -40 664 -27
rect 764 27 868 40
rect 764 -27 793 27
rect 839 -27 868 27
rect 764 -40 868 -27
rect 968 27 1072 40
rect 968 -27 997 27
rect 1043 -27 1072 27
rect 968 -40 1072 -27
rect 1172 27 1276 40
rect 1172 -27 1201 27
rect 1247 -27 1276 27
rect 1172 -40 1276 -27
rect 1376 27 1480 40
rect 1376 -27 1405 27
rect 1451 -27 1480 27
rect 1376 -40 1480 -27
rect 1580 27 1684 40
rect 1580 -27 1609 27
rect 1655 -27 1684 27
rect 1580 -40 1684 -27
rect 1784 27 1888 40
rect 1784 -27 1813 27
rect 1859 -27 1888 27
rect 1784 -40 1888 -27
rect 1988 27 2076 40
rect 1988 -27 2017 27
rect 2063 -27 2076 27
rect 1988 -40 2076 -27
<< pdiffc >>
rect -2063 -27 -2017 27
rect -1859 -27 -1813 27
rect -1655 -27 -1609 27
rect -1451 -27 -1405 27
rect -1247 -27 -1201 27
rect -1043 -27 -997 27
rect -839 -27 -793 27
rect -635 -27 -589 27
rect -431 -27 -385 27
rect -227 -27 -181 27
rect -23 -27 23 27
rect 181 -27 227 27
rect 385 -27 431 27
rect 589 -27 635 27
rect 793 -27 839 27
rect 997 -27 1043 27
rect 1201 -27 1247 27
rect 1405 -27 1451 27
rect 1609 -27 1655 27
rect 1813 -27 1859 27
rect 2017 -27 2063 27
<< polysilicon >>
rect -1988 40 -1888 84
rect -1784 40 -1684 84
rect -1580 40 -1480 84
rect -1376 40 -1276 84
rect -1172 40 -1072 84
rect -968 40 -868 84
rect -764 40 -664 84
rect -560 40 -460 84
rect -356 40 -256 84
rect -152 40 -52 84
rect 52 40 152 84
rect 256 40 356 84
rect 460 40 560 84
rect 664 40 764 84
rect 868 40 968 84
rect 1072 40 1172 84
rect 1276 40 1376 84
rect 1480 40 1580 84
rect 1684 40 1784 84
rect 1888 40 1988 84
rect -1988 -84 -1888 -40
rect -1784 -84 -1684 -40
rect -1580 -84 -1480 -40
rect -1376 -84 -1276 -40
rect -1172 -84 -1072 -40
rect -968 -84 -868 -40
rect -764 -84 -664 -40
rect -560 -84 -460 -40
rect -356 -84 -256 -40
rect -152 -84 -52 -40
rect 52 -84 152 -40
rect 256 -84 356 -40
rect 460 -84 560 -40
rect 664 -84 764 -40
rect 868 -84 968 -40
rect 1072 -84 1172 -40
rect 1276 -84 1376 -40
rect 1480 -84 1580 -40
rect 1684 -84 1784 -40
rect 1888 -84 1988 -40
<< metal1 >>
rect -2063 27 -2017 38
rect -2063 -38 -2017 -27
rect -1859 27 -1813 38
rect -1859 -38 -1813 -27
rect -1655 27 -1609 38
rect -1655 -38 -1609 -27
rect -1451 27 -1405 38
rect -1451 -38 -1405 -27
rect -1247 27 -1201 38
rect -1247 -38 -1201 -27
rect -1043 27 -997 38
rect -1043 -38 -997 -27
rect -839 27 -793 38
rect -839 -38 -793 -27
rect -635 27 -589 38
rect -635 -38 -589 -27
rect -431 27 -385 38
rect -431 -38 -385 -27
rect -227 27 -181 38
rect -227 -38 -181 -27
rect -23 27 23 38
rect -23 -38 23 -27
rect 181 27 227 38
rect 181 -38 227 -27
rect 385 27 431 38
rect 385 -38 431 -27
rect 589 27 635 38
rect 589 -38 635 -27
rect 793 27 839 38
rect 793 -38 839 -27
rect 997 27 1043 38
rect 997 -38 1043 -27
rect 1201 27 1247 38
rect 1201 -38 1247 -27
rect 1405 27 1451 38
rect 1405 -38 1451 -27
rect 1609 27 1655 38
rect 1609 -38 1655 -27
rect 1813 27 1859 38
rect 1813 -38 1859 -27
rect 2017 27 2063 38
rect 2017 -38 2063 -27
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 0.4 l 0.5 m 1 nf 20 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
