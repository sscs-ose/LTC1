magic
tech gf180mcuC
magscale 1 10
timestamp 1692567440
<< error_p >>
rect -118 -23 -107 23
rect 50 -23 61 23
<< nwell >>
rect -206 -161 206 161
<< pmos >>
rect -28 -25 28 25
<< pdiff >>
rect -120 25 -48 36
rect 48 25 120 36
rect -120 23 -28 25
rect -120 -23 -107 23
rect -61 -23 -28 23
rect -120 -25 -28 -23
rect 28 23 120 25
rect 28 -23 61 23
rect 107 -23 120 23
rect 28 -25 120 -23
rect -120 -36 -48 -25
rect 48 -36 120 -25
<< pdiffc >>
rect -107 -23 -61 23
rect 61 -23 107 23
<< polysilicon >>
rect -28 25 28 69
rect -28 -69 28 -25
<< metal1 >>
rect -118 -23 -107 23
rect -61 -23 -50 23
rect 50 -23 61 23
rect 107 -23 118 23
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 0.250 l 0.280 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
