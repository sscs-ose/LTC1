magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1319 -3233 1319 3233
<< metal4 >>
rect -316 2225 316 2230
rect -316 2197 -311 2225
rect -283 2197 -245 2225
rect -217 2197 -179 2225
rect -151 2197 -113 2225
rect -85 2197 -47 2225
rect -19 2197 19 2225
rect 47 2197 85 2225
rect 113 2197 151 2225
rect 179 2197 217 2225
rect 245 2197 283 2225
rect 311 2197 316 2225
rect -316 2159 316 2197
rect -316 2131 -311 2159
rect -283 2131 -245 2159
rect -217 2131 -179 2159
rect -151 2131 -113 2159
rect -85 2131 -47 2159
rect -19 2131 19 2159
rect 47 2131 85 2159
rect 113 2131 151 2159
rect 179 2131 217 2159
rect 245 2131 283 2159
rect 311 2131 316 2159
rect -316 2093 316 2131
rect -316 2065 -311 2093
rect -283 2065 -245 2093
rect -217 2065 -179 2093
rect -151 2065 -113 2093
rect -85 2065 -47 2093
rect -19 2065 19 2093
rect 47 2065 85 2093
rect 113 2065 151 2093
rect 179 2065 217 2093
rect 245 2065 283 2093
rect 311 2065 316 2093
rect -316 2027 316 2065
rect -316 1999 -311 2027
rect -283 1999 -245 2027
rect -217 1999 -179 2027
rect -151 1999 -113 2027
rect -85 1999 -47 2027
rect -19 1999 19 2027
rect 47 1999 85 2027
rect 113 1999 151 2027
rect 179 1999 217 2027
rect 245 1999 283 2027
rect 311 1999 316 2027
rect -316 1961 316 1999
rect -316 1933 -311 1961
rect -283 1933 -245 1961
rect -217 1933 -179 1961
rect -151 1933 -113 1961
rect -85 1933 -47 1961
rect -19 1933 19 1961
rect 47 1933 85 1961
rect 113 1933 151 1961
rect 179 1933 217 1961
rect 245 1933 283 1961
rect 311 1933 316 1961
rect -316 1895 316 1933
rect -316 1867 -311 1895
rect -283 1867 -245 1895
rect -217 1867 -179 1895
rect -151 1867 -113 1895
rect -85 1867 -47 1895
rect -19 1867 19 1895
rect 47 1867 85 1895
rect 113 1867 151 1895
rect 179 1867 217 1895
rect 245 1867 283 1895
rect 311 1867 316 1895
rect -316 1829 316 1867
rect -316 1801 -311 1829
rect -283 1801 -245 1829
rect -217 1801 -179 1829
rect -151 1801 -113 1829
rect -85 1801 -47 1829
rect -19 1801 19 1829
rect 47 1801 85 1829
rect 113 1801 151 1829
rect 179 1801 217 1829
rect 245 1801 283 1829
rect 311 1801 316 1829
rect -316 1763 316 1801
rect -316 1735 -311 1763
rect -283 1735 -245 1763
rect -217 1735 -179 1763
rect -151 1735 -113 1763
rect -85 1735 -47 1763
rect -19 1735 19 1763
rect 47 1735 85 1763
rect 113 1735 151 1763
rect 179 1735 217 1763
rect 245 1735 283 1763
rect 311 1735 316 1763
rect -316 1697 316 1735
rect -316 1669 -311 1697
rect -283 1669 -245 1697
rect -217 1669 -179 1697
rect -151 1669 -113 1697
rect -85 1669 -47 1697
rect -19 1669 19 1697
rect 47 1669 85 1697
rect 113 1669 151 1697
rect 179 1669 217 1697
rect 245 1669 283 1697
rect 311 1669 316 1697
rect -316 1631 316 1669
rect -316 1603 -311 1631
rect -283 1603 -245 1631
rect -217 1603 -179 1631
rect -151 1603 -113 1631
rect -85 1603 -47 1631
rect -19 1603 19 1631
rect 47 1603 85 1631
rect 113 1603 151 1631
rect 179 1603 217 1631
rect 245 1603 283 1631
rect 311 1603 316 1631
rect -316 1565 316 1603
rect -316 1537 -311 1565
rect -283 1537 -245 1565
rect -217 1537 -179 1565
rect -151 1537 -113 1565
rect -85 1537 -47 1565
rect -19 1537 19 1565
rect 47 1537 85 1565
rect 113 1537 151 1565
rect 179 1537 217 1565
rect 245 1537 283 1565
rect 311 1537 316 1565
rect -316 1499 316 1537
rect -316 1471 -311 1499
rect -283 1471 -245 1499
rect -217 1471 -179 1499
rect -151 1471 -113 1499
rect -85 1471 -47 1499
rect -19 1471 19 1499
rect 47 1471 85 1499
rect 113 1471 151 1499
rect 179 1471 217 1499
rect 245 1471 283 1499
rect 311 1471 316 1499
rect -316 1433 316 1471
rect -316 1405 -311 1433
rect -283 1405 -245 1433
rect -217 1405 -179 1433
rect -151 1405 -113 1433
rect -85 1405 -47 1433
rect -19 1405 19 1433
rect 47 1405 85 1433
rect 113 1405 151 1433
rect 179 1405 217 1433
rect 245 1405 283 1433
rect 311 1405 316 1433
rect -316 1367 316 1405
rect -316 1339 -311 1367
rect -283 1339 -245 1367
rect -217 1339 -179 1367
rect -151 1339 -113 1367
rect -85 1339 -47 1367
rect -19 1339 19 1367
rect 47 1339 85 1367
rect 113 1339 151 1367
rect 179 1339 217 1367
rect 245 1339 283 1367
rect 311 1339 316 1367
rect -316 1301 316 1339
rect -316 1273 -311 1301
rect -283 1273 -245 1301
rect -217 1273 -179 1301
rect -151 1273 -113 1301
rect -85 1273 -47 1301
rect -19 1273 19 1301
rect 47 1273 85 1301
rect 113 1273 151 1301
rect 179 1273 217 1301
rect 245 1273 283 1301
rect 311 1273 316 1301
rect -316 1235 316 1273
rect -316 1207 -311 1235
rect -283 1207 -245 1235
rect -217 1207 -179 1235
rect -151 1207 -113 1235
rect -85 1207 -47 1235
rect -19 1207 19 1235
rect 47 1207 85 1235
rect 113 1207 151 1235
rect 179 1207 217 1235
rect 245 1207 283 1235
rect 311 1207 316 1235
rect -316 1169 316 1207
rect -316 1141 -311 1169
rect -283 1141 -245 1169
rect -217 1141 -179 1169
rect -151 1141 -113 1169
rect -85 1141 -47 1169
rect -19 1141 19 1169
rect 47 1141 85 1169
rect 113 1141 151 1169
rect 179 1141 217 1169
rect 245 1141 283 1169
rect 311 1141 316 1169
rect -316 1103 316 1141
rect -316 1075 -311 1103
rect -283 1075 -245 1103
rect -217 1075 -179 1103
rect -151 1075 -113 1103
rect -85 1075 -47 1103
rect -19 1075 19 1103
rect 47 1075 85 1103
rect 113 1075 151 1103
rect 179 1075 217 1103
rect 245 1075 283 1103
rect 311 1075 316 1103
rect -316 1037 316 1075
rect -316 1009 -311 1037
rect -283 1009 -245 1037
rect -217 1009 -179 1037
rect -151 1009 -113 1037
rect -85 1009 -47 1037
rect -19 1009 19 1037
rect 47 1009 85 1037
rect 113 1009 151 1037
rect 179 1009 217 1037
rect 245 1009 283 1037
rect 311 1009 316 1037
rect -316 971 316 1009
rect -316 943 -311 971
rect -283 943 -245 971
rect -217 943 -179 971
rect -151 943 -113 971
rect -85 943 -47 971
rect -19 943 19 971
rect 47 943 85 971
rect 113 943 151 971
rect 179 943 217 971
rect 245 943 283 971
rect 311 943 316 971
rect -316 905 316 943
rect -316 877 -311 905
rect -283 877 -245 905
rect -217 877 -179 905
rect -151 877 -113 905
rect -85 877 -47 905
rect -19 877 19 905
rect 47 877 85 905
rect 113 877 151 905
rect 179 877 217 905
rect 245 877 283 905
rect 311 877 316 905
rect -316 839 316 877
rect -316 811 -311 839
rect -283 811 -245 839
rect -217 811 -179 839
rect -151 811 -113 839
rect -85 811 -47 839
rect -19 811 19 839
rect 47 811 85 839
rect 113 811 151 839
rect 179 811 217 839
rect 245 811 283 839
rect 311 811 316 839
rect -316 773 316 811
rect -316 745 -311 773
rect -283 745 -245 773
rect -217 745 -179 773
rect -151 745 -113 773
rect -85 745 -47 773
rect -19 745 19 773
rect 47 745 85 773
rect 113 745 151 773
rect 179 745 217 773
rect 245 745 283 773
rect 311 745 316 773
rect -316 707 316 745
rect -316 679 -311 707
rect -283 679 -245 707
rect -217 679 -179 707
rect -151 679 -113 707
rect -85 679 -47 707
rect -19 679 19 707
rect 47 679 85 707
rect 113 679 151 707
rect 179 679 217 707
rect 245 679 283 707
rect 311 679 316 707
rect -316 641 316 679
rect -316 613 -311 641
rect -283 613 -245 641
rect -217 613 -179 641
rect -151 613 -113 641
rect -85 613 -47 641
rect -19 613 19 641
rect 47 613 85 641
rect 113 613 151 641
rect 179 613 217 641
rect 245 613 283 641
rect 311 613 316 641
rect -316 575 316 613
rect -316 547 -311 575
rect -283 547 -245 575
rect -217 547 -179 575
rect -151 547 -113 575
rect -85 547 -47 575
rect -19 547 19 575
rect 47 547 85 575
rect 113 547 151 575
rect 179 547 217 575
rect 245 547 283 575
rect 311 547 316 575
rect -316 509 316 547
rect -316 481 -311 509
rect -283 481 -245 509
rect -217 481 -179 509
rect -151 481 -113 509
rect -85 481 -47 509
rect -19 481 19 509
rect 47 481 85 509
rect 113 481 151 509
rect 179 481 217 509
rect 245 481 283 509
rect 311 481 316 509
rect -316 443 316 481
rect -316 415 -311 443
rect -283 415 -245 443
rect -217 415 -179 443
rect -151 415 -113 443
rect -85 415 -47 443
rect -19 415 19 443
rect 47 415 85 443
rect 113 415 151 443
rect 179 415 217 443
rect 245 415 283 443
rect 311 415 316 443
rect -316 377 316 415
rect -316 349 -311 377
rect -283 349 -245 377
rect -217 349 -179 377
rect -151 349 -113 377
rect -85 349 -47 377
rect -19 349 19 377
rect 47 349 85 377
rect 113 349 151 377
rect 179 349 217 377
rect 245 349 283 377
rect 311 349 316 377
rect -316 311 316 349
rect -316 283 -311 311
rect -283 283 -245 311
rect -217 283 -179 311
rect -151 283 -113 311
rect -85 283 -47 311
rect -19 283 19 311
rect 47 283 85 311
rect 113 283 151 311
rect 179 283 217 311
rect 245 283 283 311
rect 311 283 316 311
rect -316 245 316 283
rect -316 217 -311 245
rect -283 217 -245 245
rect -217 217 -179 245
rect -151 217 -113 245
rect -85 217 -47 245
rect -19 217 19 245
rect 47 217 85 245
rect 113 217 151 245
rect 179 217 217 245
rect 245 217 283 245
rect 311 217 316 245
rect -316 179 316 217
rect -316 151 -311 179
rect -283 151 -245 179
rect -217 151 -179 179
rect -151 151 -113 179
rect -85 151 -47 179
rect -19 151 19 179
rect 47 151 85 179
rect 113 151 151 179
rect 179 151 217 179
rect 245 151 283 179
rect 311 151 316 179
rect -316 113 316 151
rect -316 85 -311 113
rect -283 85 -245 113
rect -217 85 -179 113
rect -151 85 -113 113
rect -85 85 -47 113
rect -19 85 19 113
rect 47 85 85 113
rect 113 85 151 113
rect 179 85 217 113
rect 245 85 283 113
rect 311 85 316 113
rect -316 47 316 85
rect -316 19 -311 47
rect -283 19 -245 47
rect -217 19 -179 47
rect -151 19 -113 47
rect -85 19 -47 47
rect -19 19 19 47
rect 47 19 85 47
rect 113 19 151 47
rect 179 19 217 47
rect 245 19 283 47
rect 311 19 316 47
rect -316 -19 316 19
rect -316 -47 -311 -19
rect -283 -47 -245 -19
rect -217 -47 -179 -19
rect -151 -47 -113 -19
rect -85 -47 -47 -19
rect -19 -47 19 -19
rect 47 -47 85 -19
rect 113 -47 151 -19
rect 179 -47 217 -19
rect 245 -47 283 -19
rect 311 -47 316 -19
rect -316 -85 316 -47
rect -316 -113 -311 -85
rect -283 -113 -245 -85
rect -217 -113 -179 -85
rect -151 -113 -113 -85
rect -85 -113 -47 -85
rect -19 -113 19 -85
rect 47 -113 85 -85
rect 113 -113 151 -85
rect 179 -113 217 -85
rect 245 -113 283 -85
rect 311 -113 316 -85
rect -316 -151 316 -113
rect -316 -179 -311 -151
rect -283 -179 -245 -151
rect -217 -179 -179 -151
rect -151 -179 -113 -151
rect -85 -179 -47 -151
rect -19 -179 19 -151
rect 47 -179 85 -151
rect 113 -179 151 -151
rect 179 -179 217 -151
rect 245 -179 283 -151
rect 311 -179 316 -151
rect -316 -217 316 -179
rect -316 -245 -311 -217
rect -283 -245 -245 -217
rect -217 -245 -179 -217
rect -151 -245 -113 -217
rect -85 -245 -47 -217
rect -19 -245 19 -217
rect 47 -245 85 -217
rect 113 -245 151 -217
rect 179 -245 217 -217
rect 245 -245 283 -217
rect 311 -245 316 -217
rect -316 -283 316 -245
rect -316 -311 -311 -283
rect -283 -311 -245 -283
rect -217 -311 -179 -283
rect -151 -311 -113 -283
rect -85 -311 -47 -283
rect -19 -311 19 -283
rect 47 -311 85 -283
rect 113 -311 151 -283
rect 179 -311 217 -283
rect 245 -311 283 -283
rect 311 -311 316 -283
rect -316 -349 316 -311
rect -316 -377 -311 -349
rect -283 -377 -245 -349
rect -217 -377 -179 -349
rect -151 -377 -113 -349
rect -85 -377 -47 -349
rect -19 -377 19 -349
rect 47 -377 85 -349
rect 113 -377 151 -349
rect 179 -377 217 -349
rect 245 -377 283 -349
rect 311 -377 316 -349
rect -316 -415 316 -377
rect -316 -443 -311 -415
rect -283 -443 -245 -415
rect -217 -443 -179 -415
rect -151 -443 -113 -415
rect -85 -443 -47 -415
rect -19 -443 19 -415
rect 47 -443 85 -415
rect 113 -443 151 -415
rect 179 -443 217 -415
rect 245 -443 283 -415
rect 311 -443 316 -415
rect -316 -481 316 -443
rect -316 -509 -311 -481
rect -283 -509 -245 -481
rect -217 -509 -179 -481
rect -151 -509 -113 -481
rect -85 -509 -47 -481
rect -19 -509 19 -481
rect 47 -509 85 -481
rect 113 -509 151 -481
rect 179 -509 217 -481
rect 245 -509 283 -481
rect 311 -509 316 -481
rect -316 -547 316 -509
rect -316 -575 -311 -547
rect -283 -575 -245 -547
rect -217 -575 -179 -547
rect -151 -575 -113 -547
rect -85 -575 -47 -547
rect -19 -575 19 -547
rect 47 -575 85 -547
rect 113 -575 151 -547
rect 179 -575 217 -547
rect 245 -575 283 -547
rect 311 -575 316 -547
rect -316 -613 316 -575
rect -316 -641 -311 -613
rect -283 -641 -245 -613
rect -217 -641 -179 -613
rect -151 -641 -113 -613
rect -85 -641 -47 -613
rect -19 -641 19 -613
rect 47 -641 85 -613
rect 113 -641 151 -613
rect 179 -641 217 -613
rect 245 -641 283 -613
rect 311 -641 316 -613
rect -316 -679 316 -641
rect -316 -707 -311 -679
rect -283 -707 -245 -679
rect -217 -707 -179 -679
rect -151 -707 -113 -679
rect -85 -707 -47 -679
rect -19 -707 19 -679
rect 47 -707 85 -679
rect 113 -707 151 -679
rect 179 -707 217 -679
rect 245 -707 283 -679
rect 311 -707 316 -679
rect -316 -745 316 -707
rect -316 -773 -311 -745
rect -283 -773 -245 -745
rect -217 -773 -179 -745
rect -151 -773 -113 -745
rect -85 -773 -47 -745
rect -19 -773 19 -745
rect 47 -773 85 -745
rect 113 -773 151 -745
rect 179 -773 217 -745
rect 245 -773 283 -745
rect 311 -773 316 -745
rect -316 -811 316 -773
rect -316 -839 -311 -811
rect -283 -839 -245 -811
rect -217 -839 -179 -811
rect -151 -839 -113 -811
rect -85 -839 -47 -811
rect -19 -839 19 -811
rect 47 -839 85 -811
rect 113 -839 151 -811
rect 179 -839 217 -811
rect 245 -839 283 -811
rect 311 -839 316 -811
rect -316 -877 316 -839
rect -316 -905 -311 -877
rect -283 -905 -245 -877
rect -217 -905 -179 -877
rect -151 -905 -113 -877
rect -85 -905 -47 -877
rect -19 -905 19 -877
rect 47 -905 85 -877
rect 113 -905 151 -877
rect 179 -905 217 -877
rect 245 -905 283 -877
rect 311 -905 316 -877
rect -316 -943 316 -905
rect -316 -971 -311 -943
rect -283 -971 -245 -943
rect -217 -971 -179 -943
rect -151 -971 -113 -943
rect -85 -971 -47 -943
rect -19 -971 19 -943
rect 47 -971 85 -943
rect 113 -971 151 -943
rect 179 -971 217 -943
rect 245 -971 283 -943
rect 311 -971 316 -943
rect -316 -1009 316 -971
rect -316 -1037 -311 -1009
rect -283 -1037 -245 -1009
rect -217 -1037 -179 -1009
rect -151 -1037 -113 -1009
rect -85 -1037 -47 -1009
rect -19 -1037 19 -1009
rect 47 -1037 85 -1009
rect 113 -1037 151 -1009
rect 179 -1037 217 -1009
rect 245 -1037 283 -1009
rect 311 -1037 316 -1009
rect -316 -1075 316 -1037
rect -316 -1103 -311 -1075
rect -283 -1103 -245 -1075
rect -217 -1103 -179 -1075
rect -151 -1103 -113 -1075
rect -85 -1103 -47 -1075
rect -19 -1103 19 -1075
rect 47 -1103 85 -1075
rect 113 -1103 151 -1075
rect 179 -1103 217 -1075
rect 245 -1103 283 -1075
rect 311 -1103 316 -1075
rect -316 -1141 316 -1103
rect -316 -1169 -311 -1141
rect -283 -1169 -245 -1141
rect -217 -1169 -179 -1141
rect -151 -1169 -113 -1141
rect -85 -1169 -47 -1141
rect -19 -1169 19 -1141
rect 47 -1169 85 -1141
rect 113 -1169 151 -1141
rect 179 -1169 217 -1141
rect 245 -1169 283 -1141
rect 311 -1169 316 -1141
rect -316 -1207 316 -1169
rect -316 -1235 -311 -1207
rect -283 -1235 -245 -1207
rect -217 -1235 -179 -1207
rect -151 -1235 -113 -1207
rect -85 -1235 -47 -1207
rect -19 -1235 19 -1207
rect 47 -1235 85 -1207
rect 113 -1235 151 -1207
rect 179 -1235 217 -1207
rect 245 -1235 283 -1207
rect 311 -1235 316 -1207
rect -316 -1273 316 -1235
rect -316 -1301 -311 -1273
rect -283 -1301 -245 -1273
rect -217 -1301 -179 -1273
rect -151 -1301 -113 -1273
rect -85 -1301 -47 -1273
rect -19 -1301 19 -1273
rect 47 -1301 85 -1273
rect 113 -1301 151 -1273
rect 179 -1301 217 -1273
rect 245 -1301 283 -1273
rect 311 -1301 316 -1273
rect -316 -1339 316 -1301
rect -316 -1367 -311 -1339
rect -283 -1367 -245 -1339
rect -217 -1367 -179 -1339
rect -151 -1367 -113 -1339
rect -85 -1367 -47 -1339
rect -19 -1367 19 -1339
rect 47 -1367 85 -1339
rect 113 -1367 151 -1339
rect 179 -1367 217 -1339
rect 245 -1367 283 -1339
rect 311 -1367 316 -1339
rect -316 -1405 316 -1367
rect -316 -1433 -311 -1405
rect -283 -1433 -245 -1405
rect -217 -1433 -179 -1405
rect -151 -1433 -113 -1405
rect -85 -1433 -47 -1405
rect -19 -1433 19 -1405
rect 47 -1433 85 -1405
rect 113 -1433 151 -1405
rect 179 -1433 217 -1405
rect 245 -1433 283 -1405
rect 311 -1433 316 -1405
rect -316 -1471 316 -1433
rect -316 -1499 -311 -1471
rect -283 -1499 -245 -1471
rect -217 -1499 -179 -1471
rect -151 -1499 -113 -1471
rect -85 -1499 -47 -1471
rect -19 -1499 19 -1471
rect 47 -1499 85 -1471
rect 113 -1499 151 -1471
rect 179 -1499 217 -1471
rect 245 -1499 283 -1471
rect 311 -1499 316 -1471
rect -316 -1537 316 -1499
rect -316 -1565 -311 -1537
rect -283 -1565 -245 -1537
rect -217 -1565 -179 -1537
rect -151 -1565 -113 -1537
rect -85 -1565 -47 -1537
rect -19 -1565 19 -1537
rect 47 -1565 85 -1537
rect 113 -1565 151 -1537
rect 179 -1565 217 -1537
rect 245 -1565 283 -1537
rect 311 -1565 316 -1537
rect -316 -1603 316 -1565
rect -316 -1631 -311 -1603
rect -283 -1631 -245 -1603
rect -217 -1631 -179 -1603
rect -151 -1631 -113 -1603
rect -85 -1631 -47 -1603
rect -19 -1631 19 -1603
rect 47 -1631 85 -1603
rect 113 -1631 151 -1603
rect 179 -1631 217 -1603
rect 245 -1631 283 -1603
rect 311 -1631 316 -1603
rect -316 -1669 316 -1631
rect -316 -1697 -311 -1669
rect -283 -1697 -245 -1669
rect -217 -1697 -179 -1669
rect -151 -1697 -113 -1669
rect -85 -1697 -47 -1669
rect -19 -1697 19 -1669
rect 47 -1697 85 -1669
rect 113 -1697 151 -1669
rect 179 -1697 217 -1669
rect 245 -1697 283 -1669
rect 311 -1697 316 -1669
rect -316 -1735 316 -1697
rect -316 -1763 -311 -1735
rect -283 -1763 -245 -1735
rect -217 -1763 -179 -1735
rect -151 -1763 -113 -1735
rect -85 -1763 -47 -1735
rect -19 -1763 19 -1735
rect 47 -1763 85 -1735
rect 113 -1763 151 -1735
rect 179 -1763 217 -1735
rect 245 -1763 283 -1735
rect 311 -1763 316 -1735
rect -316 -1801 316 -1763
rect -316 -1829 -311 -1801
rect -283 -1829 -245 -1801
rect -217 -1829 -179 -1801
rect -151 -1829 -113 -1801
rect -85 -1829 -47 -1801
rect -19 -1829 19 -1801
rect 47 -1829 85 -1801
rect 113 -1829 151 -1801
rect 179 -1829 217 -1801
rect 245 -1829 283 -1801
rect 311 -1829 316 -1801
rect -316 -1867 316 -1829
rect -316 -1895 -311 -1867
rect -283 -1895 -245 -1867
rect -217 -1895 -179 -1867
rect -151 -1895 -113 -1867
rect -85 -1895 -47 -1867
rect -19 -1895 19 -1867
rect 47 -1895 85 -1867
rect 113 -1895 151 -1867
rect 179 -1895 217 -1867
rect 245 -1895 283 -1867
rect 311 -1895 316 -1867
rect -316 -1933 316 -1895
rect -316 -1961 -311 -1933
rect -283 -1961 -245 -1933
rect -217 -1961 -179 -1933
rect -151 -1961 -113 -1933
rect -85 -1961 -47 -1933
rect -19 -1961 19 -1933
rect 47 -1961 85 -1933
rect 113 -1961 151 -1933
rect 179 -1961 217 -1933
rect 245 -1961 283 -1933
rect 311 -1961 316 -1933
rect -316 -1999 316 -1961
rect -316 -2027 -311 -1999
rect -283 -2027 -245 -1999
rect -217 -2027 -179 -1999
rect -151 -2027 -113 -1999
rect -85 -2027 -47 -1999
rect -19 -2027 19 -1999
rect 47 -2027 85 -1999
rect 113 -2027 151 -1999
rect 179 -2027 217 -1999
rect 245 -2027 283 -1999
rect 311 -2027 316 -1999
rect -316 -2065 316 -2027
rect -316 -2093 -311 -2065
rect -283 -2093 -245 -2065
rect -217 -2093 -179 -2065
rect -151 -2093 -113 -2065
rect -85 -2093 -47 -2065
rect -19 -2093 19 -2065
rect 47 -2093 85 -2065
rect 113 -2093 151 -2065
rect 179 -2093 217 -2065
rect 245 -2093 283 -2065
rect 311 -2093 316 -2065
rect -316 -2131 316 -2093
rect -316 -2159 -311 -2131
rect -283 -2159 -245 -2131
rect -217 -2159 -179 -2131
rect -151 -2159 -113 -2131
rect -85 -2159 -47 -2131
rect -19 -2159 19 -2131
rect 47 -2159 85 -2131
rect 113 -2159 151 -2131
rect 179 -2159 217 -2131
rect 245 -2159 283 -2131
rect 311 -2159 316 -2131
rect -316 -2197 316 -2159
rect -316 -2225 -311 -2197
rect -283 -2225 -245 -2197
rect -217 -2225 -179 -2197
rect -151 -2225 -113 -2197
rect -85 -2225 -47 -2197
rect -19 -2225 19 -2197
rect 47 -2225 85 -2197
rect 113 -2225 151 -2197
rect 179 -2225 217 -2197
rect 245 -2225 283 -2197
rect 311 -2225 316 -2197
rect -316 -2230 316 -2225
<< via4 >>
rect -311 2197 -283 2225
rect -245 2197 -217 2225
rect -179 2197 -151 2225
rect -113 2197 -85 2225
rect -47 2197 -19 2225
rect 19 2197 47 2225
rect 85 2197 113 2225
rect 151 2197 179 2225
rect 217 2197 245 2225
rect 283 2197 311 2225
rect -311 2131 -283 2159
rect -245 2131 -217 2159
rect -179 2131 -151 2159
rect -113 2131 -85 2159
rect -47 2131 -19 2159
rect 19 2131 47 2159
rect 85 2131 113 2159
rect 151 2131 179 2159
rect 217 2131 245 2159
rect 283 2131 311 2159
rect -311 2065 -283 2093
rect -245 2065 -217 2093
rect -179 2065 -151 2093
rect -113 2065 -85 2093
rect -47 2065 -19 2093
rect 19 2065 47 2093
rect 85 2065 113 2093
rect 151 2065 179 2093
rect 217 2065 245 2093
rect 283 2065 311 2093
rect -311 1999 -283 2027
rect -245 1999 -217 2027
rect -179 1999 -151 2027
rect -113 1999 -85 2027
rect -47 1999 -19 2027
rect 19 1999 47 2027
rect 85 1999 113 2027
rect 151 1999 179 2027
rect 217 1999 245 2027
rect 283 1999 311 2027
rect -311 1933 -283 1961
rect -245 1933 -217 1961
rect -179 1933 -151 1961
rect -113 1933 -85 1961
rect -47 1933 -19 1961
rect 19 1933 47 1961
rect 85 1933 113 1961
rect 151 1933 179 1961
rect 217 1933 245 1961
rect 283 1933 311 1961
rect -311 1867 -283 1895
rect -245 1867 -217 1895
rect -179 1867 -151 1895
rect -113 1867 -85 1895
rect -47 1867 -19 1895
rect 19 1867 47 1895
rect 85 1867 113 1895
rect 151 1867 179 1895
rect 217 1867 245 1895
rect 283 1867 311 1895
rect -311 1801 -283 1829
rect -245 1801 -217 1829
rect -179 1801 -151 1829
rect -113 1801 -85 1829
rect -47 1801 -19 1829
rect 19 1801 47 1829
rect 85 1801 113 1829
rect 151 1801 179 1829
rect 217 1801 245 1829
rect 283 1801 311 1829
rect -311 1735 -283 1763
rect -245 1735 -217 1763
rect -179 1735 -151 1763
rect -113 1735 -85 1763
rect -47 1735 -19 1763
rect 19 1735 47 1763
rect 85 1735 113 1763
rect 151 1735 179 1763
rect 217 1735 245 1763
rect 283 1735 311 1763
rect -311 1669 -283 1697
rect -245 1669 -217 1697
rect -179 1669 -151 1697
rect -113 1669 -85 1697
rect -47 1669 -19 1697
rect 19 1669 47 1697
rect 85 1669 113 1697
rect 151 1669 179 1697
rect 217 1669 245 1697
rect 283 1669 311 1697
rect -311 1603 -283 1631
rect -245 1603 -217 1631
rect -179 1603 -151 1631
rect -113 1603 -85 1631
rect -47 1603 -19 1631
rect 19 1603 47 1631
rect 85 1603 113 1631
rect 151 1603 179 1631
rect 217 1603 245 1631
rect 283 1603 311 1631
rect -311 1537 -283 1565
rect -245 1537 -217 1565
rect -179 1537 -151 1565
rect -113 1537 -85 1565
rect -47 1537 -19 1565
rect 19 1537 47 1565
rect 85 1537 113 1565
rect 151 1537 179 1565
rect 217 1537 245 1565
rect 283 1537 311 1565
rect -311 1471 -283 1499
rect -245 1471 -217 1499
rect -179 1471 -151 1499
rect -113 1471 -85 1499
rect -47 1471 -19 1499
rect 19 1471 47 1499
rect 85 1471 113 1499
rect 151 1471 179 1499
rect 217 1471 245 1499
rect 283 1471 311 1499
rect -311 1405 -283 1433
rect -245 1405 -217 1433
rect -179 1405 -151 1433
rect -113 1405 -85 1433
rect -47 1405 -19 1433
rect 19 1405 47 1433
rect 85 1405 113 1433
rect 151 1405 179 1433
rect 217 1405 245 1433
rect 283 1405 311 1433
rect -311 1339 -283 1367
rect -245 1339 -217 1367
rect -179 1339 -151 1367
rect -113 1339 -85 1367
rect -47 1339 -19 1367
rect 19 1339 47 1367
rect 85 1339 113 1367
rect 151 1339 179 1367
rect 217 1339 245 1367
rect 283 1339 311 1367
rect -311 1273 -283 1301
rect -245 1273 -217 1301
rect -179 1273 -151 1301
rect -113 1273 -85 1301
rect -47 1273 -19 1301
rect 19 1273 47 1301
rect 85 1273 113 1301
rect 151 1273 179 1301
rect 217 1273 245 1301
rect 283 1273 311 1301
rect -311 1207 -283 1235
rect -245 1207 -217 1235
rect -179 1207 -151 1235
rect -113 1207 -85 1235
rect -47 1207 -19 1235
rect 19 1207 47 1235
rect 85 1207 113 1235
rect 151 1207 179 1235
rect 217 1207 245 1235
rect 283 1207 311 1235
rect -311 1141 -283 1169
rect -245 1141 -217 1169
rect -179 1141 -151 1169
rect -113 1141 -85 1169
rect -47 1141 -19 1169
rect 19 1141 47 1169
rect 85 1141 113 1169
rect 151 1141 179 1169
rect 217 1141 245 1169
rect 283 1141 311 1169
rect -311 1075 -283 1103
rect -245 1075 -217 1103
rect -179 1075 -151 1103
rect -113 1075 -85 1103
rect -47 1075 -19 1103
rect 19 1075 47 1103
rect 85 1075 113 1103
rect 151 1075 179 1103
rect 217 1075 245 1103
rect 283 1075 311 1103
rect -311 1009 -283 1037
rect -245 1009 -217 1037
rect -179 1009 -151 1037
rect -113 1009 -85 1037
rect -47 1009 -19 1037
rect 19 1009 47 1037
rect 85 1009 113 1037
rect 151 1009 179 1037
rect 217 1009 245 1037
rect 283 1009 311 1037
rect -311 943 -283 971
rect -245 943 -217 971
rect -179 943 -151 971
rect -113 943 -85 971
rect -47 943 -19 971
rect 19 943 47 971
rect 85 943 113 971
rect 151 943 179 971
rect 217 943 245 971
rect 283 943 311 971
rect -311 877 -283 905
rect -245 877 -217 905
rect -179 877 -151 905
rect -113 877 -85 905
rect -47 877 -19 905
rect 19 877 47 905
rect 85 877 113 905
rect 151 877 179 905
rect 217 877 245 905
rect 283 877 311 905
rect -311 811 -283 839
rect -245 811 -217 839
rect -179 811 -151 839
rect -113 811 -85 839
rect -47 811 -19 839
rect 19 811 47 839
rect 85 811 113 839
rect 151 811 179 839
rect 217 811 245 839
rect 283 811 311 839
rect -311 745 -283 773
rect -245 745 -217 773
rect -179 745 -151 773
rect -113 745 -85 773
rect -47 745 -19 773
rect 19 745 47 773
rect 85 745 113 773
rect 151 745 179 773
rect 217 745 245 773
rect 283 745 311 773
rect -311 679 -283 707
rect -245 679 -217 707
rect -179 679 -151 707
rect -113 679 -85 707
rect -47 679 -19 707
rect 19 679 47 707
rect 85 679 113 707
rect 151 679 179 707
rect 217 679 245 707
rect 283 679 311 707
rect -311 613 -283 641
rect -245 613 -217 641
rect -179 613 -151 641
rect -113 613 -85 641
rect -47 613 -19 641
rect 19 613 47 641
rect 85 613 113 641
rect 151 613 179 641
rect 217 613 245 641
rect 283 613 311 641
rect -311 547 -283 575
rect -245 547 -217 575
rect -179 547 -151 575
rect -113 547 -85 575
rect -47 547 -19 575
rect 19 547 47 575
rect 85 547 113 575
rect 151 547 179 575
rect 217 547 245 575
rect 283 547 311 575
rect -311 481 -283 509
rect -245 481 -217 509
rect -179 481 -151 509
rect -113 481 -85 509
rect -47 481 -19 509
rect 19 481 47 509
rect 85 481 113 509
rect 151 481 179 509
rect 217 481 245 509
rect 283 481 311 509
rect -311 415 -283 443
rect -245 415 -217 443
rect -179 415 -151 443
rect -113 415 -85 443
rect -47 415 -19 443
rect 19 415 47 443
rect 85 415 113 443
rect 151 415 179 443
rect 217 415 245 443
rect 283 415 311 443
rect -311 349 -283 377
rect -245 349 -217 377
rect -179 349 -151 377
rect -113 349 -85 377
rect -47 349 -19 377
rect 19 349 47 377
rect 85 349 113 377
rect 151 349 179 377
rect 217 349 245 377
rect 283 349 311 377
rect -311 283 -283 311
rect -245 283 -217 311
rect -179 283 -151 311
rect -113 283 -85 311
rect -47 283 -19 311
rect 19 283 47 311
rect 85 283 113 311
rect 151 283 179 311
rect 217 283 245 311
rect 283 283 311 311
rect -311 217 -283 245
rect -245 217 -217 245
rect -179 217 -151 245
rect -113 217 -85 245
rect -47 217 -19 245
rect 19 217 47 245
rect 85 217 113 245
rect 151 217 179 245
rect 217 217 245 245
rect 283 217 311 245
rect -311 151 -283 179
rect -245 151 -217 179
rect -179 151 -151 179
rect -113 151 -85 179
rect -47 151 -19 179
rect 19 151 47 179
rect 85 151 113 179
rect 151 151 179 179
rect 217 151 245 179
rect 283 151 311 179
rect -311 85 -283 113
rect -245 85 -217 113
rect -179 85 -151 113
rect -113 85 -85 113
rect -47 85 -19 113
rect 19 85 47 113
rect 85 85 113 113
rect 151 85 179 113
rect 217 85 245 113
rect 283 85 311 113
rect -311 19 -283 47
rect -245 19 -217 47
rect -179 19 -151 47
rect -113 19 -85 47
rect -47 19 -19 47
rect 19 19 47 47
rect 85 19 113 47
rect 151 19 179 47
rect 217 19 245 47
rect 283 19 311 47
rect -311 -47 -283 -19
rect -245 -47 -217 -19
rect -179 -47 -151 -19
rect -113 -47 -85 -19
rect -47 -47 -19 -19
rect 19 -47 47 -19
rect 85 -47 113 -19
rect 151 -47 179 -19
rect 217 -47 245 -19
rect 283 -47 311 -19
rect -311 -113 -283 -85
rect -245 -113 -217 -85
rect -179 -113 -151 -85
rect -113 -113 -85 -85
rect -47 -113 -19 -85
rect 19 -113 47 -85
rect 85 -113 113 -85
rect 151 -113 179 -85
rect 217 -113 245 -85
rect 283 -113 311 -85
rect -311 -179 -283 -151
rect -245 -179 -217 -151
rect -179 -179 -151 -151
rect -113 -179 -85 -151
rect -47 -179 -19 -151
rect 19 -179 47 -151
rect 85 -179 113 -151
rect 151 -179 179 -151
rect 217 -179 245 -151
rect 283 -179 311 -151
rect -311 -245 -283 -217
rect -245 -245 -217 -217
rect -179 -245 -151 -217
rect -113 -245 -85 -217
rect -47 -245 -19 -217
rect 19 -245 47 -217
rect 85 -245 113 -217
rect 151 -245 179 -217
rect 217 -245 245 -217
rect 283 -245 311 -217
rect -311 -311 -283 -283
rect -245 -311 -217 -283
rect -179 -311 -151 -283
rect -113 -311 -85 -283
rect -47 -311 -19 -283
rect 19 -311 47 -283
rect 85 -311 113 -283
rect 151 -311 179 -283
rect 217 -311 245 -283
rect 283 -311 311 -283
rect -311 -377 -283 -349
rect -245 -377 -217 -349
rect -179 -377 -151 -349
rect -113 -377 -85 -349
rect -47 -377 -19 -349
rect 19 -377 47 -349
rect 85 -377 113 -349
rect 151 -377 179 -349
rect 217 -377 245 -349
rect 283 -377 311 -349
rect -311 -443 -283 -415
rect -245 -443 -217 -415
rect -179 -443 -151 -415
rect -113 -443 -85 -415
rect -47 -443 -19 -415
rect 19 -443 47 -415
rect 85 -443 113 -415
rect 151 -443 179 -415
rect 217 -443 245 -415
rect 283 -443 311 -415
rect -311 -509 -283 -481
rect -245 -509 -217 -481
rect -179 -509 -151 -481
rect -113 -509 -85 -481
rect -47 -509 -19 -481
rect 19 -509 47 -481
rect 85 -509 113 -481
rect 151 -509 179 -481
rect 217 -509 245 -481
rect 283 -509 311 -481
rect -311 -575 -283 -547
rect -245 -575 -217 -547
rect -179 -575 -151 -547
rect -113 -575 -85 -547
rect -47 -575 -19 -547
rect 19 -575 47 -547
rect 85 -575 113 -547
rect 151 -575 179 -547
rect 217 -575 245 -547
rect 283 -575 311 -547
rect -311 -641 -283 -613
rect -245 -641 -217 -613
rect -179 -641 -151 -613
rect -113 -641 -85 -613
rect -47 -641 -19 -613
rect 19 -641 47 -613
rect 85 -641 113 -613
rect 151 -641 179 -613
rect 217 -641 245 -613
rect 283 -641 311 -613
rect -311 -707 -283 -679
rect -245 -707 -217 -679
rect -179 -707 -151 -679
rect -113 -707 -85 -679
rect -47 -707 -19 -679
rect 19 -707 47 -679
rect 85 -707 113 -679
rect 151 -707 179 -679
rect 217 -707 245 -679
rect 283 -707 311 -679
rect -311 -773 -283 -745
rect -245 -773 -217 -745
rect -179 -773 -151 -745
rect -113 -773 -85 -745
rect -47 -773 -19 -745
rect 19 -773 47 -745
rect 85 -773 113 -745
rect 151 -773 179 -745
rect 217 -773 245 -745
rect 283 -773 311 -745
rect -311 -839 -283 -811
rect -245 -839 -217 -811
rect -179 -839 -151 -811
rect -113 -839 -85 -811
rect -47 -839 -19 -811
rect 19 -839 47 -811
rect 85 -839 113 -811
rect 151 -839 179 -811
rect 217 -839 245 -811
rect 283 -839 311 -811
rect -311 -905 -283 -877
rect -245 -905 -217 -877
rect -179 -905 -151 -877
rect -113 -905 -85 -877
rect -47 -905 -19 -877
rect 19 -905 47 -877
rect 85 -905 113 -877
rect 151 -905 179 -877
rect 217 -905 245 -877
rect 283 -905 311 -877
rect -311 -971 -283 -943
rect -245 -971 -217 -943
rect -179 -971 -151 -943
rect -113 -971 -85 -943
rect -47 -971 -19 -943
rect 19 -971 47 -943
rect 85 -971 113 -943
rect 151 -971 179 -943
rect 217 -971 245 -943
rect 283 -971 311 -943
rect -311 -1037 -283 -1009
rect -245 -1037 -217 -1009
rect -179 -1037 -151 -1009
rect -113 -1037 -85 -1009
rect -47 -1037 -19 -1009
rect 19 -1037 47 -1009
rect 85 -1037 113 -1009
rect 151 -1037 179 -1009
rect 217 -1037 245 -1009
rect 283 -1037 311 -1009
rect -311 -1103 -283 -1075
rect -245 -1103 -217 -1075
rect -179 -1103 -151 -1075
rect -113 -1103 -85 -1075
rect -47 -1103 -19 -1075
rect 19 -1103 47 -1075
rect 85 -1103 113 -1075
rect 151 -1103 179 -1075
rect 217 -1103 245 -1075
rect 283 -1103 311 -1075
rect -311 -1169 -283 -1141
rect -245 -1169 -217 -1141
rect -179 -1169 -151 -1141
rect -113 -1169 -85 -1141
rect -47 -1169 -19 -1141
rect 19 -1169 47 -1141
rect 85 -1169 113 -1141
rect 151 -1169 179 -1141
rect 217 -1169 245 -1141
rect 283 -1169 311 -1141
rect -311 -1235 -283 -1207
rect -245 -1235 -217 -1207
rect -179 -1235 -151 -1207
rect -113 -1235 -85 -1207
rect -47 -1235 -19 -1207
rect 19 -1235 47 -1207
rect 85 -1235 113 -1207
rect 151 -1235 179 -1207
rect 217 -1235 245 -1207
rect 283 -1235 311 -1207
rect -311 -1301 -283 -1273
rect -245 -1301 -217 -1273
rect -179 -1301 -151 -1273
rect -113 -1301 -85 -1273
rect -47 -1301 -19 -1273
rect 19 -1301 47 -1273
rect 85 -1301 113 -1273
rect 151 -1301 179 -1273
rect 217 -1301 245 -1273
rect 283 -1301 311 -1273
rect -311 -1367 -283 -1339
rect -245 -1367 -217 -1339
rect -179 -1367 -151 -1339
rect -113 -1367 -85 -1339
rect -47 -1367 -19 -1339
rect 19 -1367 47 -1339
rect 85 -1367 113 -1339
rect 151 -1367 179 -1339
rect 217 -1367 245 -1339
rect 283 -1367 311 -1339
rect -311 -1433 -283 -1405
rect -245 -1433 -217 -1405
rect -179 -1433 -151 -1405
rect -113 -1433 -85 -1405
rect -47 -1433 -19 -1405
rect 19 -1433 47 -1405
rect 85 -1433 113 -1405
rect 151 -1433 179 -1405
rect 217 -1433 245 -1405
rect 283 -1433 311 -1405
rect -311 -1499 -283 -1471
rect -245 -1499 -217 -1471
rect -179 -1499 -151 -1471
rect -113 -1499 -85 -1471
rect -47 -1499 -19 -1471
rect 19 -1499 47 -1471
rect 85 -1499 113 -1471
rect 151 -1499 179 -1471
rect 217 -1499 245 -1471
rect 283 -1499 311 -1471
rect -311 -1565 -283 -1537
rect -245 -1565 -217 -1537
rect -179 -1565 -151 -1537
rect -113 -1565 -85 -1537
rect -47 -1565 -19 -1537
rect 19 -1565 47 -1537
rect 85 -1565 113 -1537
rect 151 -1565 179 -1537
rect 217 -1565 245 -1537
rect 283 -1565 311 -1537
rect -311 -1631 -283 -1603
rect -245 -1631 -217 -1603
rect -179 -1631 -151 -1603
rect -113 -1631 -85 -1603
rect -47 -1631 -19 -1603
rect 19 -1631 47 -1603
rect 85 -1631 113 -1603
rect 151 -1631 179 -1603
rect 217 -1631 245 -1603
rect 283 -1631 311 -1603
rect -311 -1697 -283 -1669
rect -245 -1697 -217 -1669
rect -179 -1697 -151 -1669
rect -113 -1697 -85 -1669
rect -47 -1697 -19 -1669
rect 19 -1697 47 -1669
rect 85 -1697 113 -1669
rect 151 -1697 179 -1669
rect 217 -1697 245 -1669
rect 283 -1697 311 -1669
rect -311 -1763 -283 -1735
rect -245 -1763 -217 -1735
rect -179 -1763 -151 -1735
rect -113 -1763 -85 -1735
rect -47 -1763 -19 -1735
rect 19 -1763 47 -1735
rect 85 -1763 113 -1735
rect 151 -1763 179 -1735
rect 217 -1763 245 -1735
rect 283 -1763 311 -1735
rect -311 -1829 -283 -1801
rect -245 -1829 -217 -1801
rect -179 -1829 -151 -1801
rect -113 -1829 -85 -1801
rect -47 -1829 -19 -1801
rect 19 -1829 47 -1801
rect 85 -1829 113 -1801
rect 151 -1829 179 -1801
rect 217 -1829 245 -1801
rect 283 -1829 311 -1801
rect -311 -1895 -283 -1867
rect -245 -1895 -217 -1867
rect -179 -1895 -151 -1867
rect -113 -1895 -85 -1867
rect -47 -1895 -19 -1867
rect 19 -1895 47 -1867
rect 85 -1895 113 -1867
rect 151 -1895 179 -1867
rect 217 -1895 245 -1867
rect 283 -1895 311 -1867
rect -311 -1961 -283 -1933
rect -245 -1961 -217 -1933
rect -179 -1961 -151 -1933
rect -113 -1961 -85 -1933
rect -47 -1961 -19 -1933
rect 19 -1961 47 -1933
rect 85 -1961 113 -1933
rect 151 -1961 179 -1933
rect 217 -1961 245 -1933
rect 283 -1961 311 -1933
rect -311 -2027 -283 -1999
rect -245 -2027 -217 -1999
rect -179 -2027 -151 -1999
rect -113 -2027 -85 -1999
rect -47 -2027 -19 -1999
rect 19 -2027 47 -1999
rect 85 -2027 113 -1999
rect 151 -2027 179 -1999
rect 217 -2027 245 -1999
rect 283 -2027 311 -1999
rect -311 -2093 -283 -2065
rect -245 -2093 -217 -2065
rect -179 -2093 -151 -2065
rect -113 -2093 -85 -2065
rect -47 -2093 -19 -2065
rect 19 -2093 47 -2065
rect 85 -2093 113 -2065
rect 151 -2093 179 -2065
rect 217 -2093 245 -2065
rect 283 -2093 311 -2065
rect -311 -2159 -283 -2131
rect -245 -2159 -217 -2131
rect -179 -2159 -151 -2131
rect -113 -2159 -85 -2131
rect -47 -2159 -19 -2131
rect 19 -2159 47 -2131
rect 85 -2159 113 -2131
rect 151 -2159 179 -2131
rect 217 -2159 245 -2131
rect 283 -2159 311 -2131
rect -311 -2225 -283 -2197
rect -245 -2225 -217 -2197
rect -179 -2225 -151 -2197
rect -113 -2225 -85 -2197
rect -47 -2225 -19 -2197
rect 19 -2225 47 -2197
rect 85 -2225 113 -2197
rect 151 -2225 179 -2197
rect 217 -2225 245 -2197
rect 283 -2225 311 -2197
<< metal5 >>
rect -319 2225 319 2233
rect -319 2197 -311 2225
rect -283 2197 -245 2225
rect -217 2197 -179 2225
rect -151 2197 -113 2225
rect -85 2197 -47 2225
rect -19 2197 19 2225
rect 47 2197 85 2225
rect 113 2197 151 2225
rect 179 2197 217 2225
rect 245 2197 283 2225
rect 311 2197 319 2225
rect -319 2159 319 2197
rect -319 2131 -311 2159
rect -283 2131 -245 2159
rect -217 2131 -179 2159
rect -151 2131 -113 2159
rect -85 2131 -47 2159
rect -19 2131 19 2159
rect 47 2131 85 2159
rect 113 2131 151 2159
rect 179 2131 217 2159
rect 245 2131 283 2159
rect 311 2131 319 2159
rect -319 2093 319 2131
rect -319 2065 -311 2093
rect -283 2065 -245 2093
rect -217 2065 -179 2093
rect -151 2065 -113 2093
rect -85 2065 -47 2093
rect -19 2065 19 2093
rect 47 2065 85 2093
rect 113 2065 151 2093
rect 179 2065 217 2093
rect 245 2065 283 2093
rect 311 2065 319 2093
rect -319 2027 319 2065
rect -319 1999 -311 2027
rect -283 1999 -245 2027
rect -217 1999 -179 2027
rect -151 1999 -113 2027
rect -85 1999 -47 2027
rect -19 1999 19 2027
rect 47 1999 85 2027
rect 113 1999 151 2027
rect 179 1999 217 2027
rect 245 1999 283 2027
rect 311 1999 319 2027
rect -319 1961 319 1999
rect -319 1933 -311 1961
rect -283 1933 -245 1961
rect -217 1933 -179 1961
rect -151 1933 -113 1961
rect -85 1933 -47 1961
rect -19 1933 19 1961
rect 47 1933 85 1961
rect 113 1933 151 1961
rect 179 1933 217 1961
rect 245 1933 283 1961
rect 311 1933 319 1961
rect -319 1895 319 1933
rect -319 1867 -311 1895
rect -283 1867 -245 1895
rect -217 1867 -179 1895
rect -151 1867 -113 1895
rect -85 1867 -47 1895
rect -19 1867 19 1895
rect 47 1867 85 1895
rect 113 1867 151 1895
rect 179 1867 217 1895
rect 245 1867 283 1895
rect 311 1867 319 1895
rect -319 1829 319 1867
rect -319 1801 -311 1829
rect -283 1801 -245 1829
rect -217 1801 -179 1829
rect -151 1801 -113 1829
rect -85 1801 -47 1829
rect -19 1801 19 1829
rect 47 1801 85 1829
rect 113 1801 151 1829
rect 179 1801 217 1829
rect 245 1801 283 1829
rect 311 1801 319 1829
rect -319 1763 319 1801
rect -319 1735 -311 1763
rect -283 1735 -245 1763
rect -217 1735 -179 1763
rect -151 1735 -113 1763
rect -85 1735 -47 1763
rect -19 1735 19 1763
rect 47 1735 85 1763
rect 113 1735 151 1763
rect 179 1735 217 1763
rect 245 1735 283 1763
rect 311 1735 319 1763
rect -319 1697 319 1735
rect -319 1669 -311 1697
rect -283 1669 -245 1697
rect -217 1669 -179 1697
rect -151 1669 -113 1697
rect -85 1669 -47 1697
rect -19 1669 19 1697
rect 47 1669 85 1697
rect 113 1669 151 1697
rect 179 1669 217 1697
rect 245 1669 283 1697
rect 311 1669 319 1697
rect -319 1631 319 1669
rect -319 1603 -311 1631
rect -283 1603 -245 1631
rect -217 1603 -179 1631
rect -151 1603 -113 1631
rect -85 1603 -47 1631
rect -19 1603 19 1631
rect 47 1603 85 1631
rect 113 1603 151 1631
rect 179 1603 217 1631
rect 245 1603 283 1631
rect 311 1603 319 1631
rect -319 1565 319 1603
rect -319 1537 -311 1565
rect -283 1537 -245 1565
rect -217 1537 -179 1565
rect -151 1537 -113 1565
rect -85 1537 -47 1565
rect -19 1537 19 1565
rect 47 1537 85 1565
rect 113 1537 151 1565
rect 179 1537 217 1565
rect 245 1537 283 1565
rect 311 1537 319 1565
rect -319 1499 319 1537
rect -319 1471 -311 1499
rect -283 1471 -245 1499
rect -217 1471 -179 1499
rect -151 1471 -113 1499
rect -85 1471 -47 1499
rect -19 1471 19 1499
rect 47 1471 85 1499
rect 113 1471 151 1499
rect 179 1471 217 1499
rect 245 1471 283 1499
rect 311 1471 319 1499
rect -319 1433 319 1471
rect -319 1405 -311 1433
rect -283 1405 -245 1433
rect -217 1405 -179 1433
rect -151 1405 -113 1433
rect -85 1405 -47 1433
rect -19 1405 19 1433
rect 47 1405 85 1433
rect 113 1405 151 1433
rect 179 1405 217 1433
rect 245 1405 283 1433
rect 311 1405 319 1433
rect -319 1367 319 1405
rect -319 1339 -311 1367
rect -283 1339 -245 1367
rect -217 1339 -179 1367
rect -151 1339 -113 1367
rect -85 1339 -47 1367
rect -19 1339 19 1367
rect 47 1339 85 1367
rect 113 1339 151 1367
rect 179 1339 217 1367
rect 245 1339 283 1367
rect 311 1339 319 1367
rect -319 1301 319 1339
rect -319 1273 -311 1301
rect -283 1273 -245 1301
rect -217 1273 -179 1301
rect -151 1273 -113 1301
rect -85 1273 -47 1301
rect -19 1273 19 1301
rect 47 1273 85 1301
rect 113 1273 151 1301
rect 179 1273 217 1301
rect 245 1273 283 1301
rect 311 1273 319 1301
rect -319 1235 319 1273
rect -319 1207 -311 1235
rect -283 1207 -245 1235
rect -217 1207 -179 1235
rect -151 1207 -113 1235
rect -85 1207 -47 1235
rect -19 1207 19 1235
rect 47 1207 85 1235
rect 113 1207 151 1235
rect 179 1207 217 1235
rect 245 1207 283 1235
rect 311 1207 319 1235
rect -319 1169 319 1207
rect -319 1141 -311 1169
rect -283 1141 -245 1169
rect -217 1141 -179 1169
rect -151 1141 -113 1169
rect -85 1141 -47 1169
rect -19 1141 19 1169
rect 47 1141 85 1169
rect 113 1141 151 1169
rect 179 1141 217 1169
rect 245 1141 283 1169
rect 311 1141 319 1169
rect -319 1103 319 1141
rect -319 1075 -311 1103
rect -283 1075 -245 1103
rect -217 1075 -179 1103
rect -151 1075 -113 1103
rect -85 1075 -47 1103
rect -19 1075 19 1103
rect 47 1075 85 1103
rect 113 1075 151 1103
rect 179 1075 217 1103
rect 245 1075 283 1103
rect 311 1075 319 1103
rect -319 1037 319 1075
rect -319 1009 -311 1037
rect -283 1009 -245 1037
rect -217 1009 -179 1037
rect -151 1009 -113 1037
rect -85 1009 -47 1037
rect -19 1009 19 1037
rect 47 1009 85 1037
rect 113 1009 151 1037
rect 179 1009 217 1037
rect 245 1009 283 1037
rect 311 1009 319 1037
rect -319 971 319 1009
rect -319 943 -311 971
rect -283 943 -245 971
rect -217 943 -179 971
rect -151 943 -113 971
rect -85 943 -47 971
rect -19 943 19 971
rect 47 943 85 971
rect 113 943 151 971
rect 179 943 217 971
rect 245 943 283 971
rect 311 943 319 971
rect -319 905 319 943
rect -319 877 -311 905
rect -283 877 -245 905
rect -217 877 -179 905
rect -151 877 -113 905
rect -85 877 -47 905
rect -19 877 19 905
rect 47 877 85 905
rect 113 877 151 905
rect 179 877 217 905
rect 245 877 283 905
rect 311 877 319 905
rect -319 839 319 877
rect -319 811 -311 839
rect -283 811 -245 839
rect -217 811 -179 839
rect -151 811 -113 839
rect -85 811 -47 839
rect -19 811 19 839
rect 47 811 85 839
rect 113 811 151 839
rect 179 811 217 839
rect 245 811 283 839
rect 311 811 319 839
rect -319 773 319 811
rect -319 745 -311 773
rect -283 745 -245 773
rect -217 745 -179 773
rect -151 745 -113 773
rect -85 745 -47 773
rect -19 745 19 773
rect 47 745 85 773
rect 113 745 151 773
rect 179 745 217 773
rect 245 745 283 773
rect 311 745 319 773
rect -319 707 319 745
rect -319 679 -311 707
rect -283 679 -245 707
rect -217 679 -179 707
rect -151 679 -113 707
rect -85 679 -47 707
rect -19 679 19 707
rect 47 679 85 707
rect 113 679 151 707
rect 179 679 217 707
rect 245 679 283 707
rect 311 679 319 707
rect -319 641 319 679
rect -319 613 -311 641
rect -283 613 -245 641
rect -217 613 -179 641
rect -151 613 -113 641
rect -85 613 -47 641
rect -19 613 19 641
rect 47 613 85 641
rect 113 613 151 641
rect 179 613 217 641
rect 245 613 283 641
rect 311 613 319 641
rect -319 575 319 613
rect -319 547 -311 575
rect -283 547 -245 575
rect -217 547 -179 575
rect -151 547 -113 575
rect -85 547 -47 575
rect -19 547 19 575
rect 47 547 85 575
rect 113 547 151 575
rect 179 547 217 575
rect 245 547 283 575
rect 311 547 319 575
rect -319 509 319 547
rect -319 481 -311 509
rect -283 481 -245 509
rect -217 481 -179 509
rect -151 481 -113 509
rect -85 481 -47 509
rect -19 481 19 509
rect 47 481 85 509
rect 113 481 151 509
rect 179 481 217 509
rect 245 481 283 509
rect 311 481 319 509
rect -319 443 319 481
rect -319 415 -311 443
rect -283 415 -245 443
rect -217 415 -179 443
rect -151 415 -113 443
rect -85 415 -47 443
rect -19 415 19 443
rect 47 415 85 443
rect 113 415 151 443
rect 179 415 217 443
rect 245 415 283 443
rect 311 415 319 443
rect -319 377 319 415
rect -319 349 -311 377
rect -283 349 -245 377
rect -217 349 -179 377
rect -151 349 -113 377
rect -85 349 -47 377
rect -19 349 19 377
rect 47 349 85 377
rect 113 349 151 377
rect 179 349 217 377
rect 245 349 283 377
rect 311 349 319 377
rect -319 311 319 349
rect -319 283 -311 311
rect -283 283 -245 311
rect -217 283 -179 311
rect -151 283 -113 311
rect -85 283 -47 311
rect -19 283 19 311
rect 47 283 85 311
rect 113 283 151 311
rect 179 283 217 311
rect 245 283 283 311
rect 311 283 319 311
rect -319 245 319 283
rect -319 217 -311 245
rect -283 217 -245 245
rect -217 217 -179 245
rect -151 217 -113 245
rect -85 217 -47 245
rect -19 217 19 245
rect 47 217 85 245
rect 113 217 151 245
rect 179 217 217 245
rect 245 217 283 245
rect 311 217 319 245
rect -319 179 319 217
rect -319 151 -311 179
rect -283 151 -245 179
rect -217 151 -179 179
rect -151 151 -113 179
rect -85 151 -47 179
rect -19 151 19 179
rect 47 151 85 179
rect 113 151 151 179
rect 179 151 217 179
rect 245 151 283 179
rect 311 151 319 179
rect -319 113 319 151
rect -319 85 -311 113
rect -283 85 -245 113
rect -217 85 -179 113
rect -151 85 -113 113
rect -85 85 -47 113
rect -19 85 19 113
rect 47 85 85 113
rect 113 85 151 113
rect 179 85 217 113
rect 245 85 283 113
rect 311 85 319 113
rect -319 47 319 85
rect -319 19 -311 47
rect -283 19 -245 47
rect -217 19 -179 47
rect -151 19 -113 47
rect -85 19 -47 47
rect -19 19 19 47
rect 47 19 85 47
rect 113 19 151 47
rect 179 19 217 47
rect 245 19 283 47
rect 311 19 319 47
rect -319 -19 319 19
rect -319 -47 -311 -19
rect -283 -47 -245 -19
rect -217 -47 -179 -19
rect -151 -47 -113 -19
rect -85 -47 -47 -19
rect -19 -47 19 -19
rect 47 -47 85 -19
rect 113 -47 151 -19
rect 179 -47 217 -19
rect 245 -47 283 -19
rect 311 -47 319 -19
rect -319 -85 319 -47
rect -319 -113 -311 -85
rect -283 -113 -245 -85
rect -217 -113 -179 -85
rect -151 -113 -113 -85
rect -85 -113 -47 -85
rect -19 -113 19 -85
rect 47 -113 85 -85
rect 113 -113 151 -85
rect 179 -113 217 -85
rect 245 -113 283 -85
rect 311 -113 319 -85
rect -319 -151 319 -113
rect -319 -179 -311 -151
rect -283 -179 -245 -151
rect -217 -179 -179 -151
rect -151 -179 -113 -151
rect -85 -179 -47 -151
rect -19 -179 19 -151
rect 47 -179 85 -151
rect 113 -179 151 -151
rect 179 -179 217 -151
rect 245 -179 283 -151
rect 311 -179 319 -151
rect -319 -217 319 -179
rect -319 -245 -311 -217
rect -283 -245 -245 -217
rect -217 -245 -179 -217
rect -151 -245 -113 -217
rect -85 -245 -47 -217
rect -19 -245 19 -217
rect 47 -245 85 -217
rect 113 -245 151 -217
rect 179 -245 217 -217
rect 245 -245 283 -217
rect 311 -245 319 -217
rect -319 -283 319 -245
rect -319 -311 -311 -283
rect -283 -311 -245 -283
rect -217 -311 -179 -283
rect -151 -311 -113 -283
rect -85 -311 -47 -283
rect -19 -311 19 -283
rect 47 -311 85 -283
rect 113 -311 151 -283
rect 179 -311 217 -283
rect 245 -311 283 -283
rect 311 -311 319 -283
rect -319 -349 319 -311
rect -319 -377 -311 -349
rect -283 -377 -245 -349
rect -217 -377 -179 -349
rect -151 -377 -113 -349
rect -85 -377 -47 -349
rect -19 -377 19 -349
rect 47 -377 85 -349
rect 113 -377 151 -349
rect 179 -377 217 -349
rect 245 -377 283 -349
rect 311 -377 319 -349
rect -319 -415 319 -377
rect -319 -443 -311 -415
rect -283 -443 -245 -415
rect -217 -443 -179 -415
rect -151 -443 -113 -415
rect -85 -443 -47 -415
rect -19 -443 19 -415
rect 47 -443 85 -415
rect 113 -443 151 -415
rect 179 -443 217 -415
rect 245 -443 283 -415
rect 311 -443 319 -415
rect -319 -481 319 -443
rect -319 -509 -311 -481
rect -283 -509 -245 -481
rect -217 -509 -179 -481
rect -151 -509 -113 -481
rect -85 -509 -47 -481
rect -19 -509 19 -481
rect 47 -509 85 -481
rect 113 -509 151 -481
rect 179 -509 217 -481
rect 245 -509 283 -481
rect 311 -509 319 -481
rect -319 -547 319 -509
rect -319 -575 -311 -547
rect -283 -575 -245 -547
rect -217 -575 -179 -547
rect -151 -575 -113 -547
rect -85 -575 -47 -547
rect -19 -575 19 -547
rect 47 -575 85 -547
rect 113 -575 151 -547
rect 179 -575 217 -547
rect 245 -575 283 -547
rect 311 -575 319 -547
rect -319 -613 319 -575
rect -319 -641 -311 -613
rect -283 -641 -245 -613
rect -217 -641 -179 -613
rect -151 -641 -113 -613
rect -85 -641 -47 -613
rect -19 -641 19 -613
rect 47 -641 85 -613
rect 113 -641 151 -613
rect 179 -641 217 -613
rect 245 -641 283 -613
rect 311 -641 319 -613
rect -319 -679 319 -641
rect -319 -707 -311 -679
rect -283 -707 -245 -679
rect -217 -707 -179 -679
rect -151 -707 -113 -679
rect -85 -707 -47 -679
rect -19 -707 19 -679
rect 47 -707 85 -679
rect 113 -707 151 -679
rect 179 -707 217 -679
rect 245 -707 283 -679
rect 311 -707 319 -679
rect -319 -745 319 -707
rect -319 -773 -311 -745
rect -283 -773 -245 -745
rect -217 -773 -179 -745
rect -151 -773 -113 -745
rect -85 -773 -47 -745
rect -19 -773 19 -745
rect 47 -773 85 -745
rect 113 -773 151 -745
rect 179 -773 217 -745
rect 245 -773 283 -745
rect 311 -773 319 -745
rect -319 -811 319 -773
rect -319 -839 -311 -811
rect -283 -839 -245 -811
rect -217 -839 -179 -811
rect -151 -839 -113 -811
rect -85 -839 -47 -811
rect -19 -839 19 -811
rect 47 -839 85 -811
rect 113 -839 151 -811
rect 179 -839 217 -811
rect 245 -839 283 -811
rect 311 -839 319 -811
rect -319 -877 319 -839
rect -319 -905 -311 -877
rect -283 -905 -245 -877
rect -217 -905 -179 -877
rect -151 -905 -113 -877
rect -85 -905 -47 -877
rect -19 -905 19 -877
rect 47 -905 85 -877
rect 113 -905 151 -877
rect 179 -905 217 -877
rect 245 -905 283 -877
rect 311 -905 319 -877
rect -319 -943 319 -905
rect -319 -971 -311 -943
rect -283 -971 -245 -943
rect -217 -971 -179 -943
rect -151 -971 -113 -943
rect -85 -971 -47 -943
rect -19 -971 19 -943
rect 47 -971 85 -943
rect 113 -971 151 -943
rect 179 -971 217 -943
rect 245 -971 283 -943
rect 311 -971 319 -943
rect -319 -1009 319 -971
rect -319 -1037 -311 -1009
rect -283 -1037 -245 -1009
rect -217 -1037 -179 -1009
rect -151 -1037 -113 -1009
rect -85 -1037 -47 -1009
rect -19 -1037 19 -1009
rect 47 -1037 85 -1009
rect 113 -1037 151 -1009
rect 179 -1037 217 -1009
rect 245 -1037 283 -1009
rect 311 -1037 319 -1009
rect -319 -1075 319 -1037
rect -319 -1103 -311 -1075
rect -283 -1103 -245 -1075
rect -217 -1103 -179 -1075
rect -151 -1103 -113 -1075
rect -85 -1103 -47 -1075
rect -19 -1103 19 -1075
rect 47 -1103 85 -1075
rect 113 -1103 151 -1075
rect 179 -1103 217 -1075
rect 245 -1103 283 -1075
rect 311 -1103 319 -1075
rect -319 -1141 319 -1103
rect -319 -1169 -311 -1141
rect -283 -1169 -245 -1141
rect -217 -1169 -179 -1141
rect -151 -1169 -113 -1141
rect -85 -1169 -47 -1141
rect -19 -1169 19 -1141
rect 47 -1169 85 -1141
rect 113 -1169 151 -1141
rect 179 -1169 217 -1141
rect 245 -1169 283 -1141
rect 311 -1169 319 -1141
rect -319 -1207 319 -1169
rect -319 -1235 -311 -1207
rect -283 -1235 -245 -1207
rect -217 -1235 -179 -1207
rect -151 -1235 -113 -1207
rect -85 -1235 -47 -1207
rect -19 -1235 19 -1207
rect 47 -1235 85 -1207
rect 113 -1235 151 -1207
rect 179 -1235 217 -1207
rect 245 -1235 283 -1207
rect 311 -1235 319 -1207
rect -319 -1273 319 -1235
rect -319 -1301 -311 -1273
rect -283 -1301 -245 -1273
rect -217 -1301 -179 -1273
rect -151 -1301 -113 -1273
rect -85 -1301 -47 -1273
rect -19 -1301 19 -1273
rect 47 -1301 85 -1273
rect 113 -1301 151 -1273
rect 179 -1301 217 -1273
rect 245 -1301 283 -1273
rect 311 -1301 319 -1273
rect -319 -1339 319 -1301
rect -319 -1367 -311 -1339
rect -283 -1367 -245 -1339
rect -217 -1367 -179 -1339
rect -151 -1367 -113 -1339
rect -85 -1367 -47 -1339
rect -19 -1367 19 -1339
rect 47 -1367 85 -1339
rect 113 -1367 151 -1339
rect 179 -1367 217 -1339
rect 245 -1367 283 -1339
rect 311 -1367 319 -1339
rect -319 -1405 319 -1367
rect -319 -1433 -311 -1405
rect -283 -1433 -245 -1405
rect -217 -1433 -179 -1405
rect -151 -1433 -113 -1405
rect -85 -1433 -47 -1405
rect -19 -1433 19 -1405
rect 47 -1433 85 -1405
rect 113 -1433 151 -1405
rect 179 -1433 217 -1405
rect 245 -1433 283 -1405
rect 311 -1433 319 -1405
rect -319 -1471 319 -1433
rect -319 -1499 -311 -1471
rect -283 -1499 -245 -1471
rect -217 -1499 -179 -1471
rect -151 -1499 -113 -1471
rect -85 -1499 -47 -1471
rect -19 -1499 19 -1471
rect 47 -1499 85 -1471
rect 113 -1499 151 -1471
rect 179 -1499 217 -1471
rect 245 -1499 283 -1471
rect 311 -1499 319 -1471
rect -319 -1537 319 -1499
rect -319 -1565 -311 -1537
rect -283 -1565 -245 -1537
rect -217 -1565 -179 -1537
rect -151 -1565 -113 -1537
rect -85 -1565 -47 -1537
rect -19 -1565 19 -1537
rect 47 -1565 85 -1537
rect 113 -1565 151 -1537
rect 179 -1565 217 -1537
rect 245 -1565 283 -1537
rect 311 -1565 319 -1537
rect -319 -1603 319 -1565
rect -319 -1631 -311 -1603
rect -283 -1631 -245 -1603
rect -217 -1631 -179 -1603
rect -151 -1631 -113 -1603
rect -85 -1631 -47 -1603
rect -19 -1631 19 -1603
rect 47 -1631 85 -1603
rect 113 -1631 151 -1603
rect 179 -1631 217 -1603
rect 245 -1631 283 -1603
rect 311 -1631 319 -1603
rect -319 -1669 319 -1631
rect -319 -1697 -311 -1669
rect -283 -1697 -245 -1669
rect -217 -1697 -179 -1669
rect -151 -1697 -113 -1669
rect -85 -1697 -47 -1669
rect -19 -1697 19 -1669
rect 47 -1697 85 -1669
rect 113 -1697 151 -1669
rect 179 -1697 217 -1669
rect 245 -1697 283 -1669
rect 311 -1697 319 -1669
rect -319 -1735 319 -1697
rect -319 -1763 -311 -1735
rect -283 -1763 -245 -1735
rect -217 -1763 -179 -1735
rect -151 -1763 -113 -1735
rect -85 -1763 -47 -1735
rect -19 -1763 19 -1735
rect 47 -1763 85 -1735
rect 113 -1763 151 -1735
rect 179 -1763 217 -1735
rect 245 -1763 283 -1735
rect 311 -1763 319 -1735
rect -319 -1801 319 -1763
rect -319 -1829 -311 -1801
rect -283 -1829 -245 -1801
rect -217 -1829 -179 -1801
rect -151 -1829 -113 -1801
rect -85 -1829 -47 -1801
rect -19 -1829 19 -1801
rect 47 -1829 85 -1801
rect 113 -1829 151 -1801
rect 179 -1829 217 -1801
rect 245 -1829 283 -1801
rect 311 -1829 319 -1801
rect -319 -1867 319 -1829
rect -319 -1895 -311 -1867
rect -283 -1895 -245 -1867
rect -217 -1895 -179 -1867
rect -151 -1895 -113 -1867
rect -85 -1895 -47 -1867
rect -19 -1895 19 -1867
rect 47 -1895 85 -1867
rect 113 -1895 151 -1867
rect 179 -1895 217 -1867
rect 245 -1895 283 -1867
rect 311 -1895 319 -1867
rect -319 -1933 319 -1895
rect -319 -1961 -311 -1933
rect -283 -1961 -245 -1933
rect -217 -1961 -179 -1933
rect -151 -1961 -113 -1933
rect -85 -1961 -47 -1933
rect -19 -1961 19 -1933
rect 47 -1961 85 -1933
rect 113 -1961 151 -1933
rect 179 -1961 217 -1933
rect 245 -1961 283 -1933
rect 311 -1961 319 -1933
rect -319 -1999 319 -1961
rect -319 -2027 -311 -1999
rect -283 -2027 -245 -1999
rect -217 -2027 -179 -1999
rect -151 -2027 -113 -1999
rect -85 -2027 -47 -1999
rect -19 -2027 19 -1999
rect 47 -2027 85 -1999
rect 113 -2027 151 -1999
rect 179 -2027 217 -1999
rect 245 -2027 283 -1999
rect 311 -2027 319 -1999
rect -319 -2065 319 -2027
rect -319 -2093 -311 -2065
rect -283 -2093 -245 -2065
rect -217 -2093 -179 -2065
rect -151 -2093 -113 -2065
rect -85 -2093 -47 -2065
rect -19 -2093 19 -2065
rect 47 -2093 85 -2065
rect 113 -2093 151 -2065
rect 179 -2093 217 -2065
rect 245 -2093 283 -2065
rect 311 -2093 319 -2065
rect -319 -2131 319 -2093
rect -319 -2159 -311 -2131
rect -283 -2159 -245 -2131
rect -217 -2159 -179 -2131
rect -151 -2159 -113 -2131
rect -85 -2159 -47 -2131
rect -19 -2159 19 -2131
rect 47 -2159 85 -2131
rect 113 -2159 151 -2131
rect 179 -2159 217 -2131
rect 245 -2159 283 -2131
rect 311 -2159 319 -2131
rect -319 -2197 319 -2159
rect -319 -2225 -311 -2197
rect -283 -2225 -245 -2197
rect -217 -2225 -179 -2197
rect -151 -2225 -113 -2197
rect -85 -2225 -47 -2197
rect -19 -2225 19 -2197
rect 47 -2225 85 -2197
rect 113 -2225 151 -2197
rect 179 -2225 217 -2197
rect 245 -2225 283 -2197
rect 311 -2225 319 -2197
rect -319 -2233 319 -2225
<< end >>
