magic
tech gf180mcuC
magscale 1 10
timestamp 1690000208
<< nwell >>
rect 0 294 1532 762
rect 1128 241 1532 294
rect 1128 222 1332 241
<< pwell >>
rect 218 0 910 198
rect 1186 -2 1474 196
<< nmos >>
rect 334 74 390 124
rect 738 74 794 124
rect 1302 72 1358 122
<< pmos >>
rect 174 424 230 524
rect 334 424 390 524
rect 738 424 794 524
rect 898 424 954 524
rect 1302 371 1358 471
<< ndiff >>
rect 242 124 314 135
rect 410 124 482 135
rect 242 122 334 124
rect 242 76 255 122
rect 301 76 334 122
rect 242 74 334 76
rect 390 122 482 124
rect 390 76 423 122
rect 469 76 482 122
rect 390 74 482 76
rect 242 63 314 74
rect 410 63 482 74
rect 646 124 718 135
rect 814 124 886 135
rect 646 122 738 124
rect 646 76 659 122
rect 705 76 738 122
rect 646 74 738 76
rect 794 122 886 124
rect 794 76 827 122
rect 873 76 886 122
rect 794 74 886 76
rect 646 63 718 74
rect 814 63 886 74
rect 1210 122 1282 133
rect 1378 122 1450 133
rect 1210 120 1302 122
rect 1210 74 1223 120
rect 1269 74 1302 120
rect 1210 72 1302 74
rect 1358 120 1450 122
rect 1358 74 1391 120
rect 1437 74 1450 120
rect 1358 72 1450 74
rect 1210 61 1282 72
rect 1378 61 1450 72
<< pdiff >>
rect 86 511 174 524
rect 86 437 99 511
rect 145 437 174 511
rect 86 424 174 437
rect 230 511 334 524
rect 230 437 259 511
rect 305 437 334 511
rect 230 424 334 437
rect 390 511 478 524
rect 390 437 419 511
rect 465 437 478 511
rect 390 424 478 437
rect 650 511 738 524
rect 650 437 663 511
rect 709 437 738 511
rect 650 424 738 437
rect 794 511 898 524
rect 794 437 823 511
rect 869 437 898 511
rect 794 424 898 437
rect 954 511 1042 524
rect 954 437 983 511
rect 1029 437 1042 511
rect 954 424 1042 437
rect 1214 458 1302 471
rect 1214 384 1227 458
rect 1273 384 1302 458
rect 1214 371 1302 384
rect 1358 458 1446 471
rect 1358 384 1387 458
rect 1433 384 1446 458
rect 1358 371 1446 384
<< ndiffc >>
rect 255 76 301 122
rect 423 76 469 122
rect 659 76 705 122
rect 827 76 873 122
rect 1223 74 1269 120
rect 1391 74 1437 120
<< pdiffc >>
rect 99 437 145 511
rect 259 437 305 511
rect 419 437 465 511
rect 663 437 709 511
rect 823 437 869 511
rect 983 437 1029 511
rect 1227 384 1273 458
rect 1387 384 1433 458
<< psubdiff >>
rect 34 -72 1077 -57
rect 34 -118 64 -72
rect 1048 -118 1077 -72
rect 34 -133 1077 -118
rect 1154 -72 1502 -59
rect 1154 -121 1173 -72
rect 1482 -121 1502 -72
rect 1154 -136 1502 -121
<< nsubdiff >>
rect 24 725 1096 738
rect 24 678 45 725
rect 1067 678 1096 725
rect 24 663 1096 678
rect 1168 619 1460 636
rect 1168 568 1188 619
rect 1438 568 1460 619
rect 1168 551 1460 568
<< psubdiffcont >>
rect 64 -118 1048 -72
rect 1173 -121 1482 -72
<< nsubdiffcont >>
rect 45 678 1067 725
rect 1188 568 1438 619
<< polysilicon >>
rect 174 552 390 588
rect 174 524 230 552
rect 334 524 390 552
rect 738 551 954 590
rect 738 524 794 551
rect 898 524 954 551
rect 1302 471 1358 515
rect 174 380 230 424
rect 334 262 390 424
rect 738 377 794 424
rect 898 380 954 424
rect 659 363 794 377
rect 659 304 672 363
rect 735 304 794 363
rect 1302 309 1358 371
rect 659 290 794 304
rect 258 249 390 262
rect 258 190 272 249
rect 335 190 390 249
rect 258 175 390 190
rect 334 124 390 175
rect 334 30 390 74
rect 738 124 794 290
rect 1243 295 1358 309
rect 1243 236 1257 295
rect 1320 236 1358 295
rect 1243 222 1358 236
rect 738 30 794 74
rect 1302 122 1358 222
rect 1302 28 1358 72
<< polycontact >>
rect 672 304 735 363
rect 272 190 335 249
rect 1257 236 1320 295
<< metal1 >>
rect 0 725 1532 762
rect 0 678 45 725
rect 1067 678 1532 725
rect 0 663 1532 678
rect 99 511 145 663
rect 242 612 321 614
rect 242 558 255 612
rect 309 558 321 612
rect 242 550 321 558
rect 99 426 145 437
rect 259 511 305 550
rect 259 426 305 437
rect 419 511 465 663
rect 1128 619 1532 663
rect 649 614 723 616
rect 649 603 1029 614
rect 649 549 659 603
rect 713 568 1029 603
rect 713 549 723 568
rect 649 536 723 549
rect 419 426 465 437
rect 663 511 709 536
rect 663 426 709 437
rect 823 511 869 522
rect 659 376 748 377
rect 0 363 748 376
rect 0 330 672 363
rect 659 304 672 330
rect 735 304 748 363
rect 659 290 748 304
rect 258 249 347 262
rect 258 241 272 249
rect 0 195 272 241
rect 258 190 272 195
rect 335 190 347 249
rect 823 214 869 437
rect 983 511 1029 568
rect 1128 568 1188 619
rect 1438 568 1532 619
rect 1128 550 1532 568
rect 983 426 1029 437
rect 1204 458 1274 550
rect 1204 384 1227 458
rect 1273 384 1274 458
rect 1204 369 1274 384
rect 1386 458 1450 471
rect 1386 384 1387 458
rect 1433 384 1450 458
rect 258 175 347 190
rect 419 168 869 214
rect 419 122 465 168
rect 823 162 869 168
rect 1088 295 1332 303
rect 1088 236 1257 295
rect 1320 236 1332 295
rect 1088 222 1332 236
rect 1386 268 1450 384
rect 1088 162 1134 222
rect 823 122 1134 162
rect 1386 221 1566 268
rect 244 76 255 122
rect 301 76 312 122
rect 412 76 423 122
rect 469 76 480 122
rect 648 76 659 122
rect 705 76 716 122
rect 816 76 827 122
rect 873 116 1134 122
rect 1201 120 1282 125
rect 1386 120 1450 221
rect 873 76 884 116
rect 244 -37 312 76
rect 648 -37 716 76
rect 1201 74 1223 120
rect 1269 74 1282 120
rect 1380 74 1391 120
rect 1437 74 1450 120
rect 1201 -37 1282 74
rect 1386 73 1450 74
rect 0 -72 1532 -37
rect 0 -118 64 -72
rect 1048 -118 1173 -72
rect 0 -121 1173 -118
rect 1482 -121 1532 -72
rect 0 -150 1532 -121
<< via1 >>
rect 255 558 309 612
rect 659 549 713 603
<< metal2 >>
rect 239 614 323 624
rect 649 614 723 616
rect 239 612 723 614
rect 239 558 255 612
rect 309 603 723 612
rect 309 558 659 603
rect 239 541 323 558
rect 649 549 659 558
rect 713 549 723 603
rect 649 536 723 549
<< labels >>
flabel metal1 13 353 13 353 0 FreeSans 640 0 0 0 A
port 1 nsew
flabel metal1 21 217 21 217 0 FreeSans 640 0 0 0 B
port 2 nsew
flabel psubdiffcont 556 -94 556 -94 0 FreeSans 640 0 0 0 VSS
port 3 nsew
flabel nsubdiffcont 555 703 555 703 0 FreeSans 640 0 0 0 VDD
port 4 nsew
flabel metal1 1542 239 1542 239 0 FreeSans 640 0 0 0 OUT
port 5 nsew
flabel nsubdiffcont 1313 594 1313 594 0 FreeSans 640 0 0 0 Inverter_0.VDD
flabel psubdiffcont 1327 -98 1327 -98 0 FreeSans 640 0 0 0 Inverter_0.VSS
flabel metal1 1151 263 1151 263 0 FreeSans 640 0 0 0 Inverter_0.IN
flabel metal1 1518 236 1518 236 0 FreeSans 640 0 0 0 Inverter_0.OUT
<< end >>
