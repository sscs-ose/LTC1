magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -2264 -2348 2264 2348
<< pwell >>
rect -264 -348 264 348
<< nmos >>
rect -152 -280 -52 280
rect 52 -280 152 280
<< ndiff >>
rect -240 258 -152 280
rect -240 -258 -227 258
rect -181 -258 -152 258
rect -240 -280 -152 -258
rect -52 258 52 280
rect -52 -258 -23 258
rect 23 -258 52 258
rect -52 -280 52 -258
rect 152 258 240 280
rect 152 -258 181 258
rect 227 -258 240 258
rect 152 -280 240 -258
<< ndiffc >>
rect -227 -258 -181 258
rect -23 -258 23 258
rect 181 -258 227 258
<< polysilicon >>
rect -152 280 -52 324
rect 52 280 152 324
rect -152 -324 -52 -280
rect 52 -324 152 -280
<< metal1 >>
rect -227 258 -181 278
rect -227 -278 -181 -258
rect -23 258 23 278
rect -23 -278 23 -258
rect 181 258 227 278
rect 181 -278 227 -258
<< end >>
