magic
tech gf180mcuC
magscale 1 10
timestamp 1691669315
<< nwell >>
rect 98 310 822 833
<< pwell >>
rect 0 0 760 236
rect 778 0 1058 236
<< nmos >>
rect 112 68 168 168
rect 272 68 328 168
rect 432 68 488 168
rect 592 68 648 168
rect 890 68 946 168
<< pmos >>
rect 272 440 328 640
rect 432 440 488 640
rect 592 440 648 640
<< ndiff >>
rect 24 155 112 168
rect 24 81 37 155
rect 83 81 112 155
rect 24 68 112 81
rect 168 155 272 168
rect 168 81 197 155
rect 243 81 272 155
rect 168 68 272 81
rect 328 155 432 168
rect 328 81 357 155
rect 403 81 432 155
rect 328 68 432 81
rect 488 155 592 168
rect 488 81 517 155
rect 563 81 592 155
rect 488 68 592 81
rect 648 155 736 168
rect 648 81 677 155
rect 723 81 736 155
rect 648 68 736 81
rect 802 155 890 168
rect 802 81 815 155
rect 861 81 890 155
rect 802 68 890 81
rect 946 155 1034 168
rect 946 81 975 155
rect 1021 81 1034 155
rect 946 68 1034 81
<< pdiff >>
rect 184 627 272 640
rect 184 453 197 627
rect 243 453 272 627
rect 184 440 272 453
rect 328 627 432 640
rect 328 453 357 627
rect 403 453 432 627
rect 328 440 432 453
rect 488 627 592 640
rect 488 453 517 627
rect 563 453 592 627
rect 488 440 592 453
rect 648 627 736 640
rect 648 453 677 627
rect 723 453 736 627
rect 648 440 736 453
<< ndiffc >>
rect 37 81 83 155
rect 197 81 243 155
rect 357 81 403 155
rect 517 81 563 155
rect 677 81 723 155
rect 815 81 861 155
rect 975 81 1021 155
<< pdiffc >>
rect 197 453 243 627
rect 357 453 403 627
rect 517 453 563 627
rect 677 453 723 627
<< psubdiff >>
rect 28 -229 1041 -216
rect 28 -275 41 -229
rect 87 -275 135 -229
rect 181 -275 229 -229
rect 275 -275 323 -229
rect 369 -275 417 -229
rect 463 -275 511 -229
rect 557 -275 605 -229
rect 651 -275 699 -229
rect 745 -275 793 -229
rect 839 -275 887 -229
rect 933 -275 981 -229
rect 1027 -275 1041 -229
rect 28 -288 1041 -275
<< nsubdiff >>
rect 142 787 778 800
rect 142 741 155 787
rect 201 741 249 787
rect 295 741 343 787
rect 389 741 437 787
rect 483 741 531 787
rect 577 741 625 787
rect 671 741 719 787
rect 765 741 778 787
rect 142 728 778 741
<< psubdiffcont >>
rect 41 -275 87 -229
rect 135 -275 181 -229
rect 229 -275 275 -229
rect 323 -275 369 -229
rect 417 -275 463 -229
rect 511 -275 557 -229
rect 605 -275 651 -229
rect 699 -275 745 -229
rect 793 -275 839 -229
rect 887 -275 933 -229
rect 981 -275 1027 -229
<< nsubdiffcont >>
rect 155 741 201 787
rect 249 741 295 787
rect 343 741 389 787
rect 437 741 483 787
rect 531 741 577 787
rect 625 741 671 787
rect 719 741 765 787
<< polysilicon >>
rect 272 640 328 684
rect 432 640 488 684
rect 592 640 648 684
rect 79 281 151 289
rect 272 281 328 440
rect 79 276 328 281
rect 79 230 92 276
rect 138 230 328 276
rect 79 225 328 230
rect 79 217 168 225
rect 112 168 168 217
rect 272 168 328 225
rect 432 168 488 440
rect 592 401 648 440
rect 589 393 661 401
rect 589 388 946 393
rect 589 342 602 388
rect 648 342 946 388
rect 589 337 946 342
rect 589 329 661 337
rect 592 168 648 217
rect 890 168 946 337
rect 112 24 168 68
rect 272 24 328 68
rect 432 48 488 68
rect 592 48 648 68
rect 432 -8 648 48
rect 890 24 946 68
rect 81 -74 153 -66
rect 432 -74 488 -8
rect 81 -79 488 -74
rect 81 -125 94 -79
rect 140 -125 488 -79
rect 81 -130 488 -125
rect 81 -138 153 -130
<< polycontact >>
rect 92 230 138 276
rect 602 342 648 388
rect 94 -125 140 -79
<< metal1 >>
rect 98 787 822 820
rect 98 741 155 787
rect 201 741 249 787
rect 295 741 343 787
rect 389 741 437 787
rect 483 741 531 787
rect 577 741 625 787
rect 671 741 719 787
rect 765 741 822 787
rect 98 708 822 741
rect 197 627 243 708
rect 197 442 243 453
rect 357 627 403 638
rect 357 388 403 453
rect 517 627 563 708
rect 517 442 563 453
rect 677 627 723 638
rect 723 453 1085 488
rect 677 442 1085 453
rect 591 388 659 399
rect 197 342 602 388
rect 648 342 659 388
rect 81 276 149 287
rect 41 230 92 276
rect 138 230 149 276
rect 81 219 149 230
rect 37 155 83 166
rect 37 24 83 81
rect 197 155 243 342
rect 591 331 659 342
rect 197 70 243 81
rect 357 212 723 258
rect 357 155 403 212
rect 357 24 403 81
rect 37 -22 403 24
rect 517 155 563 166
rect 83 -79 151 -68
rect 34 -125 94 -79
rect 140 -125 151 -79
rect 83 -136 151 -125
rect 517 -196 563 81
rect 677 155 723 212
rect 677 70 723 81
rect 815 155 861 166
rect 815 -196 861 81
rect 975 155 1021 442
rect 975 70 1021 81
rect 8 -229 1061 -196
rect 8 -275 41 -229
rect 87 -275 135 -229
rect 181 -275 229 -229
rect 275 -275 323 -229
rect 369 -275 417 -229
rect 463 -275 511 -229
rect 557 -275 605 -229
rect 651 -275 699 -229
rect 745 -275 793 -229
rect 839 -275 887 -229
rect 933 -275 981 -229
rect 1027 -275 1061 -229
rect 8 -308 1061 -275
<< labels >>
flabel metal1 71 253 71 253 0 FreeSans 320 0 0 0 A
port 2 nsew
flabel metal1 1025 465 1025 465 0 FreeSans 320 0 0 0 OUT
port 4 nsew
flabel nsubdiffcont 460 764 460 764 0 FreeSans 320 0 0 0 VDD
port 5 nsew
flabel metal1 48 -102 48 -102 0 FreeSans 320 0 0 0 B
port 3 nsew
flabel psubdiffcont 534 -252 534 -252 0 FreeSans 320 0 0 0 VSS
port 6 nsew
<< end >>
