magic
tech gf180mcuC
magscale 1 10
timestamp 1690971400
<< pwell >>
rect -700 -168 700 168
<< nmos >>
rect -588 -100 -532 100
rect -428 -100 -372 100
rect -268 -100 -212 100
rect -108 -100 -52 100
rect 52 -100 108 100
rect 212 -100 268 100
rect 372 -100 428 100
rect 532 -100 588 100
<< ndiff >>
rect -676 87 -588 100
rect -676 -87 -663 87
rect -617 -87 -588 87
rect -676 -100 -588 -87
rect -532 87 -428 100
rect -532 -87 -503 87
rect -457 -87 -428 87
rect -532 -100 -428 -87
rect -372 87 -268 100
rect -372 -87 -343 87
rect -297 -87 -268 87
rect -372 -100 -268 -87
rect -212 87 -108 100
rect -212 -87 -183 87
rect -137 -87 -108 87
rect -212 -100 -108 -87
rect -52 87 52 100
rect -52 -87 -23 87
rect 23 -87 52 87
rect -52 -100 52 -87
rect 108 87 212 100
rect 108 -87 137 87
rect 183 -87 212 87
rect 108 -100 212 -87
rect 268 87 372 100
rect 268 -87 297 87
rect 343 -87 372 87
rect 268 -100 372 -87
rect 428 87 532 100
rect 428 -87 457 87
rect 503 -87 532 87
rect 428 -100 532 -87
rect 588 87 676 100
rect 588 -87 617 87
rect 663 -87 676 87
rect 588 -100 676 -87
<< ndiffc >>
rect -663 -87 -617 87
rect -503 -87 -457 87
rect -343 -87 -297 87
rect -183 -87 -137 87
rect -23 -87 23 87
rect 137 -87 183 87
rect 297 -87 343 87
rect 457 -87 503 87
rect 617 -87 663 87
<< polysilicon >>
rect -588 100 -532 144
rect -428 100 -372 144
rect -268 100 -212 144
rect -108 100 -52 144
rect 52 100 108 144
rect 212 100 268 144
rect 372 100 428 144
rect 532 100 588 144
rect -588 -144 -532 -100
rect -428 -144 -372 -100
rect -268 -144 -212 -100
rect -108 -144 -52 -100
rect 52 -144 108 -100
rect 212 -144 268 -100
rect 372 -144 428 -100
rect 532 -144 588 -100
<< metal1 >>
rect -663 87 -617 98
rect -663 -98 -617 -87
rect -503 87 -457 98
rect -503 -98 -457 -87
rect -343 87 -297 98
rect -343 -98 -297 -87
rect -183 87 -137 98
rect -183 -98 -137 -87
rect -23 87 23 98
rect -23 -98 23 -87
rect 137 87 183 98
rect 137 -98 183 -87
rect 297 87 343 98
rect 297 -98 343 -87
rect 457 87 503 98
rect 457 -98 503 -87
rect 617 87 663 98
rect 617 -98 663 -87
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 1 l 0.280 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
