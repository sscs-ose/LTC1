magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -2224 -2180 2224 2180
<< nwell >>
rect -224 -180 224 180
<< pmos >>
rect -50 -50 50 50
<< pdiff >>
rect -138 23 -50 50
rect -138 -23 -125 23
rect -79 -23 -50 23
rect -138 -50 -50 -23
rect 50 23 138 50
rect 50 -23 79 23
rect 125 -23 138 23
rect 50 -50 138 -23
<< pdiffc >>
rect -125 -23 -79 23
rect 79 -23 125 23
<< polysilicon >>
rect -50 50 50 94
rect -50 -94 50 -50
<< metal1 >>
rect -125 23 -79 48
rect -125 -48 -79 -23
rect 79 23 125 48
rect 79 -48 125 -23
<< end >>
