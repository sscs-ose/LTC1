* NGSPICE file created from nmos_3p3_GGGST2_flat.ext - technology: gf180mcuC

.subckt nmos_3p3_GGGST2_flat A B OUT VDD VSS
X0 OUT A.t1 VSS.t4 VSS.t3 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X1 OUT B.t0 a_86_407.t2 VDD.t5 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X2 VDD A.t2 a_86_407.t0 VDD.t0 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X3 VSS B.t2 OUT.t0 VSS.t0 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
R0 A.n1 A.t2 34.6599
R1 A.n0 A.t0 32.1987
R2 A.n1 A.n0 17.2076
R3 A.n0 A.t1 11.2112
R4 A A.n1 4.11202
R5 VDD.n6 VDD.t5 135.364
R6 VDD.n2 VDD.t6 75.6093
R7 VDD.n12 VDD.t0 75.608
R8 VDD.t5 VDD.n5 23.6892
R9 VDD.n14 VDD.t3 23.6892
R10 VDD.n7 VDD.n4 8.2255
R11 VDD.n15 VDD.n7 8.2255
R12 VDD VDD.n7 6.3005
R13 VDD VDD.n7 6.3005
R14 VDD.n1 VDD.n0 3.1505
R15 VDD.n4 VDD.n3 3.1505
R16 VDD.n5 VDD.n4 3.1505
R17 VDD.n7 VDD.n6 3.1505
R18 VDD.n16 VDD.n15 3.1505
R19 VDD.n15 VDD.n14 3.1505
R20 VDD.n11 VDD.n10 3.1505
R21 VDD.n13 VDD.n9 3.06224
R22 VDD.n2 VDD.n1 1.87215
R23 VDD.n12 VDD.n11 1.87197
R24 VDD.n9 VDD.t4 1.8205
R25 VDD.n9 VDD.n8 1.8205
R26 VDD.n3 VDD.n2 0.641733
R27 VDD.n13 VDD.n12 0.588896
R28 VDD VDD.n3 0.0760357
R29 VDD VDD.n16 0.0760357
R30 VDD.n16 VDD.n13 0.0535357
R31 a_86_407.n1 a_86_407.n0 5.61007
R32 a_86_407.n1 a_86_407.t0 5.61007
R33 a_86_407.n2 a_86_407.n1 2.6005
R34 a_86_407.n2 a_86_407.t2 1.8205
R35 a_86_407.n3 a_86_407.n2 1.8205
R36 VSS.n3 VSS.t0 275.707
R37 VSS.n8 VSS.t3 275.707
R38 VSS.n2 VSS.n0 6.67264
R39 VSS.n7 VSS.t4 6.67264
R40 VSS.n7 VSS.n6 2.6005
R41 VSS.n5 VSS.n4 2.6005
R42 VSS.n4 VSS.n3 2.6005
R43 VSS.n10 VSS.n9 2.6005
R44 VSS.n9 VSS.n8 2.6005
R45 VSS.n2 VSS.n1 2.6005
R46 VSS.n5 VSS.n2 0.0760357
R47 VSS.n10 VSS.n7 0.0760357
R48 VSS VSS.n5 0.0422857
R49 VSS VSS.n10 0.03425
R50 OUT.n4 OUT.n3 3.76289
R51 OUT.n3 OUT.t0 3.2765
R52 OUT.n3 OUT.n2 3.2765
R53 OUT.n4 OUT.n1 2.88224
R54 OUT.n1 OUT.t3 1.8205
R55 OUT.n1 OUT.n0 1.8205
R56 OUT OUT.n4 0.155065
R57 B B.n1 25.611
R58 B.n0 B.t2 22.0309
R59 B.n1 B.t1 21.3791
R60 B.n0 B.t0 21.3791
R61 B.n1 B.n0 20.8576
C0 VDD B 0.247f
C1 A B 0.0387f
C2 VDD OUT 0.02f
C3 OUT A 0.0248f
C4 OUT B 0.0857f
C5 VDD A 0.225f
.ends

