* NGSPICE file created from mux_4x1_flat.ext - technology: gf180mcuC

.subckt mux_4x1_flat I1 I2 I3 S1 S0 OUT VDD VSS I0
X0 VDD S1.t0 mux_2x1_1.nand2_1.IN2 VDD.t27 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1 mux_2x1_0.nand2_2.IN2 S0.t0 VSS.t22 VSS.t21 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2 mux_2x1_1.I1 mux_2x1_0.nand2_1.IN2 VDD.t48 VDD.t47 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X3 mux_2x1_0.nand2_2.OUT I2.t0 a_733_712# VSS.t6 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X4 VDD I2.t1 mux_2x1_0.nand2_2.OUT VDD.t11 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X5 mux_2x1_1.I0 mux_2x1_2.nand2_1.IN2 VDD.t33 VDD.t32 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X6 mux_2x1_1.nand2_2.IN2 S1.t1 VDD.t26 VDD.t25 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X7 mux_2x1_2.nand2_1.IN2 S0.t1 a_n956_1312# VSS.t20 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X8 VDD mux_2x1_1.nand2_2.OUT OUT.t1 VDD.t8 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X9 a_1859_712# mux_2x1_1.nand2_2.IN2 VSS.t26 VSS.t15 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X10 mux_2x1_1.nand2_2.OUT mux_2x1_1.nand2_2.IN2 VDD.t50 VDD.t49 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X11 OUT mux_2x1_1.nand2_1.IN2 VDD.t35 VDD.t34 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X12 a_n393_712# mux_2x1_2.nand2_2.IN2 VSS.t10 VSS.t9 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X13 mux_2x1_2.nand2_2.OUT mux_2x1_2.nand2_2.IN2 VDD.t24 VDD.t23 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X14 mux_2x1_1.nand2_1.IN2 mux_2x1_1.I1 VDD.t22 VDD.t21 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X15 mux_2x1_0.nand2_1.IN2 S0.t2 a_170_1312# VSS.t19 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X16 mux_2x1_1.I1 mux_2x1_0.nand2_2.OUT a_733_1312# VSS.t6 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X17 mux_2x1_2.nand2_2.IN2 S0.t3 VDD.t17 VDD.t16 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X18 mux_2x1_2.nand2_1.IN2 I1.t0 VDD.t1 VDD.t0 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X19 VDD mux_2x1_2.nand2_2.OUT mux_2x1_1.I0 VDD.t2 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X20 a_170_1312# I3.t0 VSS.t1 VSS.t0 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X21 mux_2x1_1.nand2_2.OUT mux_2x1_1.I0 a_1859_712# VSS.t3 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X22 VDD mux_2x1_1.I0 mux_2x1_1.nand2_2.OUT VDD.t38 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X23 mux_2x1_1.nand2_2.IN2 S1.t2 VSS.t13 VSS.t12 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X24 mux_2x1_1.nand2_1.IN2 S1.t3 a_1296_1312# VSS.t11 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X25 a_733_1312# mux_2x1_0.nand2_1.IN2 VSS.t25 VSS.t4 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X26 VDD S0.t4 mux_2x1_2.nand2_1.IN2 VDD.t44 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X27 a_n393_1312# mux_2x1_2.nand2_1.IN2 VSS.t14 VSS.t9 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X28 mux_2x1_2.nand2_2.IN2 S0.t5 VSS.t18 VSS.t17 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X29 a_733_712# mux_2x1_0.nand2_2.IN2 VSS.t5 VSS.t4 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X30 mux_2x1_0.nand2_2.OUT mux_2x1_0.nand2_2.IN2 VDD.t15 VDD.t14 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X31 OUT mux_2x1_1.nand2_2.OUT a_1859_1312# VSS.t3 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X32 a_1859_1312# mux_2x1_1.nand2_1.IN2 VSS.t16 VSS.t15 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X33 mux_2x1_0.nand2_2.IN2 S0.t6 VDD.t37 VDD.t36 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X34 VDD mux_2x1_0.nand2_2.OUT mux_2x1_1.I1 VDD.t18 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X35 a_1296_1312# mux_2x1_1.I1 VSS.t8 VSS.t7 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X36 VDD S0.t7 mux_2x1_0.nand2_1.IN2 VDD.t5 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X37 VDD I0.t0 mux_2x1_2.nand2_2.OUT VDD.t41 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X38 mux_2x1_0.nand2_1.IN2 I3.t1 VDD.t31 VDD.t30 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X39 mux_2x1_2.nand2_2.OUT I0.t1 a_n393_712# VSS.t2 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X40 a_n956_1312# I1.t1 VSS.t24 VSS.t23 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X41 mux_2x1_1.I0 mux_2x1_2.nand2_2.OUT a_n393_1312# VSS.t2 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
R0 S1.n3 S1.t3 31.528
R1 S1.n0 S1.t1 25.7638
R2 S1.n3 S1.t0 15.3826
R3 S1.n0 S1.t2 13.2969
R4 S1.n4 S1.n3 7.62076
R5 S1.n6 S1.n5 4.54699
R6 S1.n2 S1 4.52833
R7 S1.n1 S1.n0 2.11815
R8 S1.n5 S1.n2 1.33848
R9 S1.n1 S1 1.13555
R10 S1.n5 S1.n4 1.12145
R11 S1 S1.n6 0.0780197
R12 S1.n6 S1 0.0359098
R13 S1.n2 S1 0.0252959
R14 S1.n4 S1 0.00197541
R15 S1 S1.n1 0.00142783
R16 VDD.t34 VDD.t27 763.259
R17 VDD.t18 VDD.t21 763.259
R18 VDD.t2 VDD.t30 763.259
R19 VDD.t44 VDD.t32 763.259
R20 VDD.n10 VDD.t49 386.348
R21 VDD.n36 VDD.t14 386.348
R22 VDD.n42 VDD.t23 386.348
R23 VDD.n10 VDD.t25 362.409
R24 VDD.n36 VDD.t36 362.409
R25 VDD.n42 VDD.t16 362.409
R26 VDD.n43 VDD.n42 319.75
R27 VDD.n37 VDD.n36 319.75
R28 VDD.n14 VDD.n10 319.75
R29 VDD.n19 VDD.t8 193.183
R30 VDD.n27 VDD.t27 193.183
R31 VDD.n28 VDD.t18 193.183
R32 VDD.n2 VDD.t5 193.183
R33 VDD.n4 VDD.t2 193.183
R34 VDD.n48 VDD.t44 193.183
R35 VDD.n9 VDD.t38 193.183
R36 VDD.n35 VDD.t11 193.183
R37 VDD.n41 VDD.t41 193.183
R38 VDD.n19 VDD.t34 109.849
R39 VDD.t21 VDD.n27 109.849
R40 VDD.n28 VDD.t47 109.849
R41 VDD.t30 VDD.n2 109.849
R42 VDD.t32 VDD.n4 109.849
R43 VDD.n48 VDD.t0 109.849
R44 VDD.t49 VDD.n9 109.849
R45 VDD.t14 VDD.n35 109.849
R46 VDD.t23 VDD.n41 109.849
R47 VDD.n15 VDD 11.7877
R48 VDD.n41 VDD.n40 6.3005
R49 VDD.n35 VDD.n34 6.3005
R50 VDD.n9 VDD.n8 6.3005
R51 VDD.n20 VDD.n19 6.3005
R52 VDD.n27 VDD.n26 6.3005
R53 VDD.n29 VDD.n28 6.3005
R54 VDD.n55 VDD.n2 6.3005
R55 VDD.n52 VDD.n4 6.3005
R56 VDD.n49 VDD.n48 6.3005
R57 VDD VDD.n7 5.23855
R58 VDD VDD.n18 5.23855
R59 VDD.n49 VDD.t1 5.21701
R60 VDD.n43 VDD.t17 5.19258
R61 VDD.n38 VDD.t37 5.14703
R62 VDD.n13 VDD.t26 5.14703
R63 VDD.n54 VDD.t31 5.13746
R64 VDD.n25 VDD.t22 5.13746
R65 VDD.n50 VDD.n47 5.13287
R66 VDD.n53 VDD.n3 5.13287
R67 VDD.n1 VDD.n0 5.13287
R68 VDD.n24 VDD.n23 5.13287
R69 VDD.n22 VDD.n6 5.13287
R70 VDD.n39 VDD.n5 5.13287
R71 VDD.n12 VDD.n11 5.13287
R72 VDD.n46 VDD.t33 3.91303
R73 VDD.n31 VDD.t48 3.91303
R74 VDD.n17 VDD.t35 3.91303
R75 VDD.n46 VDD.n45 3.87623
R76 VDD.n32 VDD.n31 3.87623
R77 VDD.n17 VDD.n16 3.87523
R78 VDD.n16 VDD.t50 3.51093
R79 VDD.n45 VDD.t24 3.51093
R80 VDD.n32 VDD.t15 3.51093
R81 VDD.n13 VDD.n12 0.852084
R82 VDD.n44 VDD 0.31523
R83 VDD.n33 VDD 0.31523
R84 VDD.n45 VDD.n44 0.272927
R85 VDD.n33 VDD.n32 0.272927
R86 VDD.n16 VDD.n15 0.272927
R87 VDD.n51 VDD.n46 0.22389
R88 VDD.n31 VDD.n30 0.22389
R89 VDD.n21 VDD.n17 0.22389
R90 VDD.n39 VDD.n38 0.197419
R91 VDD.n22 VDD.n21 0.141016
R92 VDD.n25 VDD.n24 0.141016
R93 VDD.n30 VDD.n1 0.141016
R94 VDD.n54 VDD.n53 0.141016
R95 VDD.n51 VDD.n50 0.141016
R96 VDD VDD.n39 0.106177
R97 VDD.n12 VDD 0.106177
R98 VDD VDD.n22 0.106177
R99 VDD.n24 VDD 0.106177
R100 VDD VDD.n1 0.106177
R101 VDD.n53 VDD 0.106177
R102 VDD.n50 VDD 0.106177
R103 VDD.n21 VDD.n20 0.0800484
R104 VDD.n26 VDD.n25 0.0800484
R105 VDD.n30 VDD.n29 0.0800484
R106 VDD.n52 VDD.n51 0.0800484
R107 VDD VDD.n54 0.0788871
R108 VDD.n44 VDD 0.0783065
R109 VDD VDD.n33 0.0783065
R110 VDD.n15 VDD 0.0783065
R111 VDD.n38 VDD.n37 0.0460556
R112 VDD.n14 VDD.n13 0.0460556
R113 VDD.n40 VDD 0.00224194
R114 VDD.n34 VDD 0.00224194
R115 VDD.n8 VDD 0.00224194
R116 VDD.n40 VDD 0.00166129
R117 VDD.n34 VDD 0.00166129
R118 VDD.n8 VDD 0.00166129
R119 VDD.n20 VDD 0.00166129
R120 VDD.n26 VDD 0.00166129
R121 VDD.n29 VDD 0.00166129
R122 VDD VDD.n55 0.00166129
R123 VDD.n55 VDD 0.00166129
R124 VDD VDD.n52 0.00166129
R125 VDD VDD.n49 0.00166129
R126 VDD VDD.n43 0.00105556
R127 VDD.n37 VDD 0.00105556
R128 VDD VDD.n14 0.00105556
R129 S0.n3 S0.t1 31.528
R130 S0.n0 S0.t2 31.528
R131 S0.n6 S0.t3 25.7638
R132 S0.n13 S0.t6 25.7638
R133 S0.n3 S0.t4 15.3826
R134 S0.n0 S0.t7 15.3826
R135 S0.n6 S0.t5 13.2969
R136 S0.n13 S0.t0 13.2969
R137 S0.n1 S0.n0 7.6289
R138 S0.n4 S0.n3 7.62076
R139 S0.n2 S0 4.53443
R140 S0.n8 S0 4.52833
R141 S0 S0.n12 4.52833
R142 S0.n11 S0.n10 2.19776
R143 S0.n7 S0.n6 2.11815
R144 S0.n14 S0.n13 2.11815
R145 S0.n5 S0.n4 1.5005
R146 S0.n9 S0.n8 1.31042
R147 S0.n12 S0.n11 1.28387
R148 S0.n7 S0 1.13555
R149 S0 S0.n14 1.13555
R150 S0.n11 S0.n1 0.948428
R151 S0.n1 S0 0.108522
R152 S0.n2 S0 0.0780742
R153 S0.n4 S0.n2 0.0373852
R154 S0.n10 S0.n9 0.0359098
R155 S0.n8 S0 0.0252959
R156 S0 S0.n12 0.0252959
R157 S0.n5 S0 0.00345082
R158 S0.n10 S0.n5 0.00197541
R159 S0 S0.n7 0.00142783
R160 S0.n14 S0 0.00142783
R161 VSS.t11 VSS.t15 1483.3
R162 VSS.t7 VSS.t6 1483.3
R163 VSS.t19 VSS.t4 1483.3
R164 VSS.t2 VSS.t0 1483.3
R165 VSS.t20 VSS.t9 1483.3
R166 VSS.n5 VSS.t3 353.341
R167 VSS.n11 VSS.t6 353.341
R168 VSS.n15 VSS.t2 353.341
R169 VSS.t15 VSS.n5 235.561
R170 VSS.n7 VSS.t7 235.561
R171 VSS.t4 VSS.n11 235.561
R172 VSS.t0 VSS.n14 235.561
R173 VSS.t9 VSS.n15 235.561
R174 VSS.n17 VSS.t23 235.561
R175 VSS.n16 VSS.t18 9.34566
R176 VSS.n2 VSS.t13 9.34566
R177 VSS.n0 VSS.t22 9.34566
R178 VSS VSS.t24 7.24801
R179 VSS.n21 VSS.t14 7.19156
R180 VSS.n21 VSS.t10 7.19156
R181 VSS.n4 VSS.t16 7.19156
R182 VSS.n4 VSS.t26 7.19156
R183 VSS.n9 VSS.t8 7.19156
R184 VSS.n10 VSS.t25 7.19156
R185 VSS.n10 VSS.t5 7.19156
R186 VSS.n22 VSS.t1 7.19156
R187 VSS.t12 VSS.t11 3.68113
R188 VSS.t21 VSS.t19 3.68113
R189 VSS.t17 VSS.t20 3.68113
R190 VSS.n13 VSS.n12 3.37613
R191 VSS.n8 VSS.n6 3.37613
R192 VSS.n19 VSS.n18 3.37613
R193 VSS VSS.n15 2.6035
R194 VSS.n11 VSS 2.6035
R195 VSS.n5 VSS 2.60269
R196 VSS.n18 VSS 2.6005
R197 VSS.n18 VSS.n17 2.6005
R198 VSS.n20 VSS.n19 2.6005
R199 VSS.n19 VSS.t17 2.6005
R200 VSS VSS.n8 2.6005
R201 VSS.n8 VSS.n7 2.6005
R202 VSS.n6 VSS.n3 2.6005
R203 VSS.n6 VSS.t12 2.6005
R204 VSS VSS.n13 2.6005
R205 VSS.n14 VSS.n13 2.6005
R206 VSS.n12 VSS.n1 2.6005
R207 VSS.n12 VSS.t21 2.6005
R208 VSS.n22 VSS 0.171522
R209 VSS VSS.n9 0.171522
R210 VSS.n21 VSS 0.117596
R211 VSS.n4 VSS 0.117596
R212 VSS.n10 VSS 0.117596
R213 VSS VSS.n21 0.0595367
R214 VSS VSS.n4 0.0595367
R215 VSS VSS.n10 0.0595367
R216 VSS.n9 VSS 0.0569474
R217 VSS VSS.n22 0.0569474
R218 VSS.n16 VSS 0.0340526
R219 VSS VSS.n2 0.0340526
R220 VSS VSS.n0 0.0340526
R221 VSS VSS.n20 0.0139211
R222 VSS VSS.n3 0.0139211
R223 VSS VSS.n1 0.0139211
R224 VSS VSS.n16 0.00405263
R225 VSS VSS.n2 0.00405263
R226 VSS.n0 VSS 0.00247368
R227 VSS.n20 VSS 0.000894737
R228 VSS.n3 VSS 0.000894737
R229 VSS.n1 VSS 0.000894737
R230 I2.n0 I2.t0 31.528
R231 I2.n0 I2.t1 15.3826
R232 I2.n1 I2.n0 8.74076
R233 I2.n1 I2 0.116779
R234 I2 I2.n1 0.00202542
R235 OUT OUT.n2 7.15141
R236 OUT.n3 OUT.n1 3.2163
R237 OUT.n1 OUT.t1 2.2755
R238 OUT.n1 OUT.n0 2.2755
R239 OUT OUT.n3 0.0445816
R240 OUT.n3 OUT 0.0119545
R241 I1.n0 I1.t0 30.9379
R242 I1.n0 I1.t1 21.6422
R243 I1 I1.n0 4.00388
R244 I3.n0 I3.t1 30.9379
R245 I3.n0 I3.t0 21.6422
R246 I3 I3.n0 4.0005
R247 I0.n0 I0.t1 31.528
R248 I0.n0 I0.t0 15.3826
R249 I0 I0.n0 8.74076
C0 VDD mux_2x1_1.nand2_2.OUT 0.634f
C1 mux_2x1_2.nand2_1.IN2 a_n393_1312# 0.00372f
C2 mux_2x1_1.nand2_1.IN2 S0 4.45e-19
C3 mux_2x1_1.nand2_2.OUT a_1859_712# 0.0964f
C4 a_1859_1312# OUT 0.069f
C5 mux_2x1_1.I0 OUT 5.19e-19
C6 S0 I3 0.0665f
C7 mux_2x1_1.nand2_1.IN2 mux_2x1_1.I1 0.11f
C8 mux_2x1_1.I0 mux_2x1_1.nand2_2.IN2 0.0646f
C9 mux_2x1_1.I0 I0 0.0148f
C10 VDD a_n956_1312# 3.14e-19
C11 mux_2x1_2.nand2_2.OUT I0 0.202f
C12 I2 mux_2x1_1.I1 1.36e-19
C13 mux_2x1_0.nand2_2.IN2 I0 0.0036f
C14 S0 mux_2x1_1.I1 0.0109f
C15 mux_2x1_1.I0 mux_2x1_2.nand2_2.IN2 0.0048f
C16 mux_2x1_2.nand2_2.OUT mux_2x1_2.nand2_2.IN2 0.12f
C17 mux_2x1_1.I0 a_170_1312# 0.00211f
C18 OUT S1 0.00946f
C19 mux_2x1_2.nand2_1.IN2 a_n956_1312# 0.069f
C20 a_733_712# mux_2x1_1.I0 8.2e-19
C21 VDD OUT 0.234f
C22 mux_2x1_1.nand2_1.IN2 a_1859_1312# 0.00372f
C23 mux_2x1_1.nand2_2.IN2 S1 0.136f
C24 a_733_712# mux_2x1_0.nand2_2.IN2 0.00372f
C25 mux_2x1_1.nand2_1.IN2 mux_2x1_1.I0 0.00155f
C26 VDD mux_2x1_1.nand2_2.IN2 0.402f
C27 VDD I0 0.254f
C28 mux_2x1_1.nand2_1.IN2 a_1296_1312# 0.069f
C29 I2 mux_2x1_1.I0 0.0101f
C30 mux_2x1_1.nand2_2.IN2 a_1859_712# 0.00372f
C31 I1 S0 0.0576f
C32 I2 mux_2x1_0.nand2_2.IN2 0.0473f
C33 mux_2x1_1.I0 S0 0.198f
C34 mux_2x1_1.nand2_2.IN2 mux_2x1_0.nand2_2.OUT 0.0113f
C35 mux_2x1_2.nand2_2.IN2 VDD 0.401f
C36 mux_2x1_0.nand2_1.IN2 a_170_1312# 0.069f
C37 mux_2x1_2.nand2_2.OUT S0 0.0521f
C38 S0 mux_2x1_0.nand2_2.IN2 0.136f
C39 VDD a_170_1312# 3.14e-19
C40 a_n393_712# I0 0.00293f
C41 mux_2x1_1.I0 I3 0.0454f
C42 a_733_712# S1 2.15e-19
C43 mux_2x1_2.nand2_2.OUT I3 0.0174f
C44 OUT mux_2x1_1.nand2_2.OUT 0.303f
C45 a_733_712# VDD 0.00444f
C46 mux_2x1_1.nand2_1.IN2 S1 0.341f
C47 mux_2x1_2.nand2_2.IN2 a_n393_712# 0.00372f
C48 mux_2x1_2.nand2_2.IN2 mux_2x1_2.nand2_1.IN2 0.00212f
C49 mux_2x1_1.nand2_1.IN2 VDD 0.461f
C50 I2 S1 0.00408f
C51 mux_2x1_1.nand2_2.IN2 mux_2x1_1.nand2_2.OUT 0.12f
C52 mux_2x1_1.I0 mux_2x1_1.I1 0.00147f
C53 a_733_712# mux_2x1_0.nand2_2.OUT 0.0964f
C54 I2 VDD 0.255f
C55 S0 S1 0.00205f
C56 a_1296_1312# mux_2x1_1.I1 0.00372f
C57 mux_2x1_0.nand2_1.IN2 S0 0.378f
C58 mux_2x1_1.nand2_1.IN2 mux_2x1_0.nand2_2.OUT 0.0106f
C59 S0 VDD 1.56f
C60 I2 mux_2x1_0.nand2_2.OUT 0.202f
C61 mux_2x1_0.nand2_1.IN2 I3 0.0959f
C62 VDD I3 0.153f
C63 S0 mux_2x1_0.nand2_2.OUT 0.00113f
C64 S0 a_n393_1312# 9.5e-19
C65 S0 a_n393_712# 6.89e-19
C66 mux_2x1_2.nand2_1.IN2 S0 0.368f
C67 mux_2x1_1.I1 S1 0.0593f
C68 mux_2x1_1.nand2_1.IN2 mux_2x1_1.nand2_2.OUT 0.053f
C69 mux_2x1_1.I0 a_1859_1312# 2.44e-19
C70 mux_2x1_0.nand2_1.IN2 mux_2x1_1.I1 0.109f
C71 a_733_1312# mux_2x1_1.I1 0.069f
C72 VDD mux_2x1_1.I1 0.423f
C73 mux_2x1_2.nand2_2.OUT mux_2x1_1.I0 0.63f
C74 mux_2x1_1.I0 a_1296_1312# 1.04e-19
C75 mux_2x1_1.I0 mux_2x1_0.nand2_2.IN2 0.019f
C76 mux_2x1_2.nand2_2.OUT mux_2x1_0.nand2_2.IN2 0.0113f
C77 mux_2x1_1.I1 mux_2x1_0.nand2_2.OUT 0.328f
C78 mux_2x1_1.I0 S1 0.0157f
C79 VDD a_1859_1312# 0.00444f
C80 mux_2x1_1.I0 mux_2x1_0.nand2_1.IN2 0.0169f
C81 a_1296_1312# S1 0.0144f
C82 I1 VDD 0.146f
C83 mux_2x1_1.I0 a_733_1312# 2.44e-19
C84 S1 mux_2x1_0.nand2_2.IN2 3.65e-19
C85 mux_2x1_1.I0 VDD 1.29f
C86 mux_2x1_2.nand2_2.OUT mux_2x1_0.nand2_1.IN2 0.0102f
C87 mux_2x1_0.nand2_1.IN2 mux_2x1_0.nand2_2.IN2 0.00212f
C88 mux_2x1_2.nand2_2.OUT VDD 0.662f
C89 VDD a_1296_1312# 3.14e-19
C90 VDD mux_2x1_0.nand2_2.IN2 0.402f
C91 mux_2x1_1.I0 a_1859_712# 0.00375f
C92 S0 a_n956_1312# 0.0144f
C93 mux_2x1_2.nand2_2.IN2 I0 0.0473f
C94 mux_2x1_1.I0 mux_2x1_0.nand2_2.OUT 0.0242f
C95 a_1296_1312# mux_2x1_0.nand2_2.OUT 9.43e-19
C96 I1 mux_2x1_2.nand2_1.IN2 0.0959f
C97 mux_2x1_0.nand2_2.IN2 mux_2x1_0.nand2_2.OUT 0.12f
C98 mux_2x1_1.I0 a_n393_1312# 0.069f
C99 mux_2x1_1.I0 mux_2x1_2.nand2_1.IN2 0.109f
C100 mux_2x1_1.I0 a_n393_712# 1.5e-19
C101 mux_2x1_1.nand2_1.IN2 OUT 0.109f
C102 mux_2x1_2.nand2_2.OUT a_n393_1312# 0.00949f
C103 mux_2x1_2.nand2_2.OUT mux_2x1_2.nand2_1.IN2 0.053f
C104 mux_2x1_2.nand2_2.OUT a_n393_712# 0.0964f
C105 mux_2x1_0.nand2_1.IN2 S1 4.51e-21
C106 mux_2x1_1.nand2_1.IN2 mux_2x1_1.nand2_2.IN2 0.00212f
C107 VDD S1 0.594f
C108 a_1859_1312# mux_2x1_1.nand2_2.OUT 0.00949f
C109 mux_2x1_0.nand2_1.IN2 a_733_1312# 0.00372f
C110 S0 OUT 6.5e-20
C111 mux_2x1_0.nand2_1.IN2 VDD 0.46f
C112 mux_2x1_1.I0 mux_2x1_1.nand2_2.OUT 0.25f
C113 VDD a_733_1312# 0.00444f
C114 I2 mux_2x1_1.nand2_2.IN2 0.0036f
C115 S1 a_1859_712# 2.62e-19
C116 S0 I0 0.00438f
C117 S1 mux_2x1_0.nand2_2.OUT 0.108f
C118 VDD a_1859_712# 0.00444f
C119 mux_2x1_0.nand2_1.IN2 mux_2x1_0.nand2_2.OUT 0.053f
C120 a_733_1312# mux_2x1_0.nand2_2.OUT 0.00949f
C121 VDD mux_2x1_0.nand2_2.OUT 0.666f
C122 VDD a_n393_1312# 0.00444f
C123 mux_2x1_2.nand2_2.IN2 S0 0.137f
C124 mux_2x1_2.nand2_1.IN2 VDD 0.456f
C125 VDD a_n393_712# 0.00444f
C126 S0 a_170_1312# 0.0151f
C127 a_733_712# I2 0.00293f
C128 mux_2x1_1.nand2_2.OUT S1 4.46e-19
C129 I1 a_n956_1312# 0.00347f
C130 I3 a_170_1312# 0.00347f
C131 a_733_712# S0 2.62e-19
C132 a_1859_712# VSS 0.0676f
C133 mux_2x1_1.nand2_2.IN2 VSS 0.422f
C134 a_733_712# VSS 0.0676f
C135 I2 VSS 0.232f
C136 mux_2x1_0.nand2_2.IN2 VSS 0.422f
C137 a_n393_712# VSS 0.0676f
C138 I0 VSS 0.232f
C139 mux_2x1_2.nand2_2.IN2 VSS 0.437f
C140 a_1859_1312# VSS 0.0676f
C141 a_1296_1312# VSS 0.0676f
C142 a_733_1312# VSS 0.0676f
C143 a_170_1312# VSS 0.0676f
C144 a_n393_1312# VSS 0.0676f
C145 a_n956_1312# VSS 0.0678f
C146 OUT VSS 0.14f
C147 mux_2x1_1.I0 VSS 1.1f
C148 mux_2x1_1.nand2_2.OUT VSS 0.651f
C149 mux_2x1_1.nand2_1.IN2 VSS 0.412f
C150 S1 VSS 0.702f
C151 mux_2x1_1.I1 VSS 0.416f
C152 mux_2x1_0.nand2_2.OUT VSS 0.489f
C153 mux_2x1_0.nand2_1.IN2 VSS 0.412f
C154 I3 VSS 0.257f
C155 mux_2x1_2.nand2_2.OUT VSS 0.437f
C156 mux_2x1_2.nand2_1.IN2 VSS 0.435f
C157 S0 VSS 1.75f
C158 I1 VSS 0.292f
C159 VDD VSS 12.3f
.ends

