* NGSPICE file created from PFD_T2_flat.ext - technology: gf180mcuC

.subckt PFD_ver_2_pex UP VDD VSS FIN FDIV DOWN
X0 Buffer_V_2_1.IN INV_mag_0.IN.t17 VDD.t43 VDD.t42 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X1 Buffer_V_2_0.IN INV_mag_0.OUT VSS.t35 VSS.t34 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X2 Buffer_V_2_0.IN INV_mag_1.IN.t17 VDD.t81 VDD.t80 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X3 VDD INV_mag_0.IN.t18 Buffer_V_2_1.IN VDD.t39 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X4 UP a_2895_3200# VSS.t42 VSS.t16 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X5 Buffer_V_2_1.IN INV_mag_1.OUT VSS.t64 VSS.t62 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X6 VSS INV_mag_1.IN.t18 a_1176_1116# VSS.t19 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X7 INV_mag_1.IN a_306_350.t4 VDD.t82 VDD.t67 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X8 INV_mag_0.IN a_305_3341.t4 VDD.t110 VDD.t21 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X9 VDD FIN.t0 a_305_3341.t0 VDD.t0 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X10 VDD INV_mag_1.IN.t19 Buffer_V_2_0.IN VDD.t49 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X11 VSS INV_mag_0.IN.t19 a_1175_2256# VSS.t10 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X12 a_218_2267# INV_mag_1.OUT VSS.t63 VSS.t62 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X13 DOWN a_2896_302# VSS.t4 VSS.t3 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X14 VDD Buffer_V_2_1.IN a_2895_3200# VDD.t46 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X15 INV_mag_0.IN FIN.t1 a_219_2510# VSS.t32 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X16 VDD INV_mag_0.IN.t20 INV_mag_0.OUT VDD.t36 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X17 a_2896_302# Buffer_V_2_0.IN VDD.t66 VDD.t65 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X18 a_219_1360# INV_mag_1.OUT VSS.t60 VSS.t34 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X19 VDD a_306_350.t5 INV_mag_1.IN.t5 VDD.t71 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X20 VSS Buffer_V_2_1.IN a_2895_3200# VSS.t16 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X21 VSS INV_mag_1.OUT Buffer_V_2_1.IN VSS.t58 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X22 Buffer_V_2_0.IN INV_mag_1.IN.t20 a_1176_1116# VSS.t19 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X23 VDD Buffer_V_2_0.IN a_2896_302# VDD.t62 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X24 INV_mag_0.OUT INV_mag_0.IN.t21 VSS.t13 VSS.t12 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.5u
X25 INV_mag_1.IN a_306_350.t6 VDD.t5 VDD.t4 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X26 VDD INV_mag_0.IN.t22 Buffer_V_2_1.IN VDD.t31 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X27 VSS INV_mag_1.IN.t21 a_1176_1116# VSS.t20 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X28 a_220_1117# FDIV.t0 INV_mag_1.IN.t3 VSS.t5 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X29 INV_mag_0.IN a_305_3341.t5 VDD.t111 VDD.t42 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X30 INV_mag_0.IN a_305_3341.t6 VDD.t113 VDD.t112 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X31 Buffer_V_2_0.IN INV_mag_1.IN.t22 VDD.t68 VDD.t67 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X32 VDD a_306_350.t7 INV_mag_1.IN.t1 VDD.t6 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X33 VDD INV_mag_1.IN.t23 INV_mag_1.OUT VDD.t36 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X34 DOWN a_2896_302# VDD.t19 VDD.t18 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X35 VDD a_305_3341.t7 INV_mag_0.IN.t5 VDD.t0 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X36 VDD a_305_3341.t8 INV_mag_0.IN.t6 VDD.t39 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X37 VSS a_305_3341.t9 a_219_2510# VSS.t36 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X38 a_1175_2256# INV_mag_0.IN.t23 VSS.t11 VSS.t6 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X39 a_1776_787# INV_mag_0.IN.t24 VDD.t34 VDD.t33 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X40 VDD a_306_350.t8 INV_mag_1.IN.t2 VDD.t9 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X41 VDD a_305_3341.t10 INV_mag_0.IN.t7 VDD.t93 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X42 INV_mag_0.OUT INV_mag_0.IN.t25 VDD.t30 VDD.t29 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X43 VDD INV_mag_1.IN.t24 Buffer_V_2_0.IN VDD.t71 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X44 Buffer_V_2_0.IN INV_mag_1.IN.t25 a_1176_1116# VSS.t20 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X45 INV_mag_1.IN INV_mag_1.IN.t15 a_1776_787# VDD.t79 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X46 INV_mag_1.IN a_306_350.t9 VDD.t101 VDD.t100 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X47 INV_mag_1.IN a_306_350.t10 VDD.t103 VDD.t102 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X48 VDD a_2895_3200# UP.t2 VDD.t76 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X49 INV_mag_0.IN INV_mag_0.IN.t3 a_1775_2840# VDD.t28 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X50 VDD a_2896_302# DOWN.t1 VDD.t15 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X51 Buffer_V_2_1.IN INV_mag_0.IN.t27 a_1175_2256# VSS.t7 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X52 Buffer_V_2_0.IN INV_mag_1.IN.t27 VDD.t55 VDD.t4 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X53 VDD INV_mag_0.IN.t28 a_1776_787# VDD.t25 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X54 a_1176_1116# INV_mag_1.IN.t28 VSS.t24 VSS.t23 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X55 INV_mag_1.IN FDIV.t1 a_220_1117# VSS.t48 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X56 a_220_1117# a_306_350.t11 VSS.t50 VSS.t49 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X57 VSS INV_mag_0.OUT Buffer_V_2_0.IN VSS.t29 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X58 VDD a_305_3341.t11 INV_mag_0.IN.t8 VDD.t31 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X59 a_1776_787# INV_mag_1.IN.t13 INV_mag_1.IN.t14 VDD.t3 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X60 Buffer_V_2_1.IN INV_mag_0.IN.t29 VDD.t24 VDD.t23 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X61 INV_mag_1.OUT INV_mag_1.IN.t29 VDD.t52 VDD.t29 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X62 INV_mag_1.IN a_306_350.t12 VDD.t89 VDD.t88 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X63 INV_mag_0.IN a_305_3341.t12 VDD.t98 VDD.t56 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X64 a_2895_3200# Buffer_V_2_1.IN VDD.t45 VDD.t44 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X65 VSS INV_mag_1.OUT a_219_1360# VSS.t29 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X66 a_1176_1116# INV_mag_1.IN.t30 Buffer_V_2_0.IN VSS.t23 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X67 VDD a_306_350.t13 INV_mag_1.IN.t9 VDD.t90 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X68 a_1775_2840# INV_mag_1.IN.t31 VDD.t54 VDD.t53 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X69 Buffer_V_2_1.IN INV_mag_0.IN.t30 a_1175_2256# VSS.t10 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X70 VSS a_306_350.t14 a_220_1117# VSS.t45 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X71 INV_mag_1.IN a_306_350.t15 VDD.t85 VDD.t80 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X72 VDD a_305_3341.t13 INV_mag_0.IN.t10 VDD.t104 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X73 Buffer_V_2_1.IN INV_mag_0.IN.t31 VDD.t22 VDD.t21 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X74 VSS INV_mag_1.OUT Buffer_V_2_1.IN VSS.t51 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X75 INV_mag_1.OUT INV_mag_1.IN.t32 VSS.t2 VSS.t1 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.5u
X76 INV_mag_0.IN a_305_3341.t14 VDD.t107 VDD.t23 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X77 INV_mag_0.IN a_305_3341.t15 VDD.t109 VDD.t108 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X78 VDD INV_mag_1.IN.t33 a_1775_2840# VDD.t12 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X79 a_219_2510# a_305_3341.t16 VSS.t66 VSS.t65 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X80 VSS INV_mag_1.OUT a_218_2267# VSS.t51 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X81 VDD a_306_350.t16 INV_mag_1.IN.t7 VDD.t49 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X82 a_219_2510# FIN.t3 INV_mag_0.IN.t0 VSS.t0 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X83 a_218_2267# INV_mag_0.OUT a_305_3341.t2 VSS.t28 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X84 VSS INV_mag_0.IN.t32 a_1175_2256# VSS.t7 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X85 VDD FDIV.t3 a_306_350.t3 VDD.t90 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X86 a_1775_2840# INV_mag_0.IN.t1 INV_mag_0.IN.t2 VDD.t20 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X87 VSS INV_mag_0.OUT Buffer_V_2_0.IN VSS.t25 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X88 UP a_2895_3200# VDD.t75 VDD.t74 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X89 a_1175_2256# INV_mag_0.IN.t33 Buffer_V_2_1.IN VSS.t6 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X90 a_219_1360# INV_mag_0.OUT a_306_350.t0 VSS.t0 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X91 VSS Buffer_V_2_0.IN a_2896_302# VSS.t39 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
R0 INV_mag_0.IN.n24 INV_mag_0.IN.t3 219.017
R1 INV_mag_0.IN.n3 INV_mag_0.IN.t20 116.993
R2 INV_mag_0.IN.n27 INV_mag_0.IN.t29 33.8279
R3 INV_mag_0.IN.n28 INV_mag_0.IN.n27 30.2144
R4 INV_mag_0.IN.t17 INV_mag_0.IN.n1 25.0458
R5 INV_mag_0.IN.n30 INV_mag_0.IN.n29 16.5048
R6 INV_mag_0.IN.n31 INV_mag_0.IN.n30 16.5048
R7 INV_mag_0.IN.n1 INV_mag_0.IN.t27 15.3305
R8 INV_mag_0.IN.n5 INV_mag_0.IN.t28 15.2644
R9 INV_mag_0.IN.n1 INV_mag_0.IN.n28 12.8616
R10 INV_mag_0.IN.n5 INV_mag_0.IN.t24 12.7717
R11 INV_mag_0.IN.n6 INV_mag_0.IN.t17 12.0785
R12 INV_mag_0.IN.n4 INV_mag_0.IN.n3 11.3197
R13 INV_mag_0.IN.n24 INV_mag_0.IN.t1 10.8543
R14 INV_mag_0.IN.n3 INV_mag_0.IN.t21 10.2935
R15 INV_mag_0.IN.n29 INV_mag_0.IN.t30 9.4175
R16 INV_mag_0.IN.n30 INV_mag_0.IN.t33 9.4175
R17 INV_mag_0.IN.t27 INV_mag_0.IN.n31 9.4175
R18 INV_mag_0.IN.n29 INV_mag_0.IN.t19 9.1985
R19 INV_mag_0.IN.n30 INV_mag_0.IN.t23 9.1985
R20 INV_mag_0.IN.n31 INV_mag_0.IN.t32 9.1985
R21 INV_mag_0.IN.n32 INV_mag_0.IN.n5 8.99637
R22 INV_mag_0.IN.n4 INV_mag_0.IN.t25 8.74171
R23 INV_mag_0.IN.n1 INV_mag_0.IN.t22 8.05323
R24 INV_mag_0.IN.n15 INV_mag_0.IN.n14 6.76657
R25 INV_mag_0.IN.n2 INV_mag_0.IN.n23 6.46389
R26 INV_mag_0.IN.n20 INV_mag_0.IN.n8 5.77603
R27 INV_mag_0.IN.n15 INV_mag_0.IN.n12 5.58741
R28 INV_mag_0.IN INV_mag_0.IN.n32 5.21028
R29 INV_mag_0.IN.n2 INV_mag_0.IN.n24 4.7386
R30 INV_mag_0.IN INV_mag_0.IN.n4 4.69432
R31 INV_mag_0.IN.n27 INV_mag_0.IN.t18 3.6505
R32 INV_mag_0.IN.n28 INV_mag_0.IN.t31 3.6505
R33 INV_mag_0.IN.n22 INV_mag_0.IN.t10 3.6405
R34 INV_mag_0.IN.n22 INV_mag_0.IN.n21 3.6405
R35 INV_mag_0.IN.n10 INV_mag_0.IN.t8 3.6405
R36 INV_mag_0.IN.n10 INV_mag_0.IN.n9 3.6405
R37 INV_mag_0.IN.n12 INV_mag_0.IN.t5 3.6405
R38 INV_mag_0.IN.n12 INV_mag_0.IN.n11 3.6405
R39 INV_mag_0.IN.n17 INV_mag_0.IN.t6 3.6405
R40 INV_mag_0.IN.n17 INV_mag_0.IN.n16 3.6405
R41 INV_mag_0.IN.n8 INV_mag_0.IN.t7 3.6405
R42 INV_mag_0.IN.n8 INV_mag_0.IN.n7 3.6405
R43 INV_mag_0.IN.n26 INV_mag_0.IN.t2 3.6405
R44 INV_mag_0.IN.n26 INV_mag_0.IN.n25 3.6405
R45 INV_mag_0.IN.n14 INV_mag_0.IN.t0 3.2765
R46 INV_mag_0.IN.n14 INV_mag_0.IN.n13 3.2765
R47 INV_mag_0.IN.n20 INV_mag_0.IN.n19 3.15378
R48 INV_mag_0.IN.n2 INV_mag_0.IN.n26 2.94651
R49 INV_mag_0.IN.n18 INV_mag_0.IN.n17 2.92863
R50 INV_mag_0.IN.n19 INV_mag_0.IN.n10 2.6005
R51 INV_mag_0.IN.n0 INV_mag_0.IN.n22 2.6005
R52 INV_mag_0.IN.n0 INV_mag_0.IN.n20 2.57308
R53 INV_mag_0.IN.n18 INV_mag_0.IN.n15 2.26925
R54 INV_mag_0.IN.n19 INV_mag_0.IN.n18 1.00114
R55 INV_mag_0.IN.n32 INV_mag_0.IN.n6 3.21412
R56 INV_mag_0.IN.n0 INV_mag_0.IN.n2 1.67584
R57 INV_mag_0.IN.n6 INV_mag_0.IN.n0 0.431204
R58 VDD.t65 VDD.t3 432.243
R59 VDD.t44 VDD.t20 339.613
R60 VDD.t18 VDD.t15 316.279
R61 VDD.t62 VDD.t65 316.279
R62 VDD.t74 VDD.t76 282.159
R63 VDD.t46 VDD.t44 282.159
R64 VDD.t104 VDD.t42 188.018
R65 VDD.t42 VDD.t31 188.018
R66 VDD.t31 VDD.t21 188.018
R67 VDD.t21 VDD.t39 188.018
R68 VDD.t39 VDD.t23 188.018
R69 VDD.t23 VDD.t0 188.018
R70 VDD.t0 VDD.t56 188.018
R71 VDD.n56 VDD.t62 184.496
R72 VDD.t4 VDD.t9 180.213
R73 VDD.t71 VDD.t4 180.213
R74 VDD.t67 VDD.t49 180.213
R75 VDD.t49 VDD.t80 180.213
R76 VDD.t80 VDD.t90 180.213
R77 VDD.t90 VDD.t88 180.213
R78 VDD.n13 VDD.t46 164.593
R79 VDD.n64 VDD.t67 161.661
R80 VDD.n56 VDD.t18 131.784
R81 VDD.n49 VDD.t36 120.213
R82 VDD.t20 VDD.t108 118.191
R83 VDD.t28 VDD.t93 118.191
R84 VDD.t53 VDD.t112 118.191
R85 VDD.n13 VDD.t74 117.567
R86 VDD.t6 VDD.t79 113.275
R87 VDD.t100 VDD.t33 113.275
R88 VDD.t12 VDD.t104 108.948
R89 VDD.t9 VDD.t25 104.418
R90 VDD.n49 VDD.t29 96.809
R91 VDD.t108 VDD.t28 70.1759
R92 VDD.t93 VDD.t53 70.1759
R93 VDD.t112 VDD.t12 70.1759
R94 VDD.t79 VDD.t102 67.2571
R95 VDD.t33 VDD.t6 67.2571
R96 VDD.t25 VDD.t100 67.2571
R97 VDD.n64 VDD.t71 18.5517
R98 VDD.n38 VDD.t57 6.94485
R99 VDD.n79 VDD.t99 6.94485
R100 VDD.n44 VDD.t45 6.68267
R101 VDD.n52 VDD.n51 6.61305
R102 VDD.n47 VDD.n12 6.58706
R103 VDD.n50 VDD.t30 6.54616
R104 VDD.n50 VDD.t52 6.54616
R105 VDD.n59 VDD.t66 6.52811
R106 VDD.n55 VDD.n11 6.52199
R107 VDD.n53 VDD.n48 6.51831
R108 VDD.n46 VDD.n13 6.3005
R109 VDD.n57 VDD.n56 6.3005
R110 VDD.n38 VDD.t98 6.2405
R111 VDD.n79 VDD.t89 6.2405
R112 VDD.n54 VDD.n47 5.1934
R113 VDD.n8 VDD.n7 3.99669
R114 VDD.n20 VDD.n19 3.99665
R115 VDD.n7 VDD.t34 3.80383
R116 VDD.n19 VDD.t54 3.80304
R117 VDD.n28 VDD.t107 3.6405
R118 VDD.n28 VDD.n27 3.6405
R119 VDD.n30 VDD.t24 3.6405
R120 VDD.n30 VDD.n29 3.6405
R121 VDD.n32 VDD.t22 3.6405
R122 VDD.n32 VDD.n31 3.6405
R123 VDD.n34 VDD.t43 3.6405
R124 VDD.n34 VDD.n33 3.6405
R125 VDD.n26 VDD.t110 3.6405
R126 VDD.n26 VDD.n25 3.6405
R127 VDD.n24 VDD.t111 3.6405
R128 VDD.n24 VDD.n23 3.6405
R129 VDD.n22 VDD.t113 3.6405
R130 VDD.n22 VDD.n21 3.6405
R131 VDD.n17 VDD.t109 3.6405
R132 VDD.n17 VDD.n16 3.6405
R133 VDD.n15 VDD.t75 3.6405
R134 VDD.n15 VDD.n14 3.6405
R135 VDD.n10 VDD.t19 3.6405
R136 VDD.n10 VDD.n9 3.6405
R137 VDD.n5 VDD.t103 3.6405
R138 VDD.n5 VDD.n4 3.6405
R139 VDD.n3 VDD.t101 3.6405
R140 VDD.n3 VDD.n2 3.6405
R141 VDD.n1 VDD.t5 3.6405
R142 VDD.n1 VDD.n0 3.6405
R143 VDD.n67 VDD.t82 3.6405
R144 VDD.n67 VDD.n66 3.6405
R145 VDD.n77 VDD.t85 3.6405
R146 VDD.n77 VDD.n76 3.6405
R147 VDD.n69 VDD.t81 3.6405
R148 VDD.n69 VDD.n68 3.6405
R149 VDD.n73 VDD.t55 3.6405
R150 VDD.n73 VDD.n72 3.6405
R151 VDD.n71 VDD.t68 3.6405
R152 VDD.n71 VDD.n70 3.6405
R153 VDD.n35 VDD.n34 3.54622
R154 VDD.n74 VDD.n73 3.54622
R155 VDD.n7 VDD.n6 3.20353
R156 VDD.n19 VDD.n18 3.20342
R157 VDD VDD.n49 3.15269
R158 VDD VDD.n65 3.1505
R159 VDD.n65 VDD.n64 3.1505
R160 VDD.n40 VDD.n26 3.13854
R161 VDD.n41 VDD.n24 3.13854
R162 VDD.n42 VDD.n22 3.13854
R163 VDD.n61 VDD.n3 3.13659
R164 VDD.n62 VDD.n1 3.13659
R165 VDD.n81 VDD.n67 3.13659
R166 VDD.n45 VDD.n15 3.04267
R167 VDD.n58 VDD.n10 2.88811
R168 VDD.n36 VDD.n30 2.78441
R169 VDD.n35 VDD.n32 2.78441
R170 VDD.n75 VDD.n69 2.78441
R171 VDD.n74 VDD.n71 2.78441
R172 VDD.n37 VDD.n28 2.6005
R173 VDD.n78 VDD.n77 2.6005
R174 VDD.n20 VDD.n17 1.64018
R175 VDD.n8 VDD.n5 1.64018
R176 VDD.n55 VDD.n54 0.800311
R177 VDD.n36 VDD.n35 0.798761
R178 VDD.n75 VDD.n74 0.798761
R179 VDD.n39 VDD.n38 0.674543
R180 VDD.n80 VDD.n79 0.652059
R181 VDD.n39 VDD.n37 0.538543
R182 VDD.n80 VDD.n78 0.536587
R183 VDD.n43 VDD.n20 0.502171
R184 VDD.n60 VDD.n8 0.500214
R185 VDD.n37 VDD.n36 0.430935
R186 VDD.n78 VDD.n75 0.430935
R187 VDD.n54 VDD.n53 0.153071
R188 VDD.n44 VDD.n43 0.139165
R189 VDD.n43 VDD.n42 0.1365
R190 VDD.n42 VDD.n41 0.1365
R191 VDD.n41 VDD.n40 0.1365
R192 VDD.n40 VDD.n39 0.1365
R193 VDD.n60 VDD.n59 0.127292
R194 VDD.n59 VDD.n58 0.115972
R195 VDD.n61 VDD.n60 0.115972
R196 VDD.n62 VDD.n61 0.115972
R197 VDD.n81 VDD.n80 0.115972
R198 VDD VDD.n55 0.110028
R199 VDD.n45 VDD.n44 0.101936
R200 VDD.n47 VDD 0.0967155
R201 VDD VDD.n81 0.0811604
R202 VDD VDD.n50 0.0798636
R203 VDD.n52 VDD 0.0778182
R204 VDD.n53 VDD.n52 0.0363784
R205 VDD VDD.n62 0.0353113
R206 VDD.n65 VDD.n63 0.00534988
R207 VDD.n58 VDD.n57 0.00531132
R208 VDD.n46 VDD.n45 0.00497514
R209 VDD.n57 VDD 0.00134906
R210 VDD VDD.n46 0.00124586
R211 VSS.t12 VSS.t3 9017.57
R212 VSS.n41 VSS.n25 5518.87
R213 VSS.t29 VSS.n41 898.405
R214 VSS.n40 VSS.t39 803.232
R215 VSS.n42 VSS.t49 650.385
R216 VSS.n26 VSS.n25 493.043
R217 VSS.n33 VSS.t39 490.178
R218 VSS.t23 VSS.t10 390.616
R219 VSS.t19 VSS.t6 390.616
R220 VSS.t65 VSS.t45 390.616
R221 VSS.t36 VSS.t5 390.616
R222 VSS.t20 VSS.t58 390.072
R223 VSS.t34 VSS.t51 389.693
R224 VSS.t25 VSS.t62 389.693
R225 VSS.t28 VSS.t48 388.692
R226 VSS.n32 VSS.n26 364.678
R227 VSS.n40 VSS.n32 323.834
R228 VSS.t3 VSS.n39 321.293
R229 VSS.n40 VSS.t12 242.145
R230 VSS.n25 VSS.t16 128.367
R231 VSS.n41 VSS.n40 100.385
R232 VSS.n39 VSS.t1 24.7153
R233 VSS.n42 VSS.t7 9.62158
R234 VSS.n21 VSS.n5 6.8902
R235 VSS.n22 VSS.n4 6.87063
R236 VSS.n37 VSS.t2 6.71903
R237 VSS.n30 VSS.t13 6.71644
R238 VSS.n9 VSS.t63 6.62607
R239 VSS.n17 VSS.t60 6.62607
R240 VSS.n10 VSS.n6 6.6202
R241 VSS.n18 VSS.n14 6.6202
R242 VSS.n12 VSS.n11 6.4265
R243 VSS.n19 VSS.n13 6.4265
R244 VSS VSS.n43 5.2005
R245 VSS VSS.n43 5.2005
R246 VSS.n33 VSS.t1 4.11964
R247 VSS.n48 VSS.n45 4.11115
R248 VSS.n48 VSS.n47 4.0918
R249 VSS.n23 VSS.n3 3.60687
R250 VSS.n24 VSS.n1 3.5873
R251 VSS.n30 VSS.n29 3.40289
R252 VSS.n37 VSS.n36 3.40289
R253 VSS.n9 VSS.n8 3.3442
R254 VSS.n17 VSS.n16 3.3442
R255 VSS.n29 VSS.t42 3.2765
R256 VSS.n29 VSS.n28 3.2765
R257 VSS.n36 VSS.t4 3.2765
R258 VSS.n36 VSS.n35 3.2765
R259 VSS.n8 VSS.t64 3.2765
R260 VSS.n8 VSS.n7 3.2765
R261 VSS.n1 VSS.t11 3.2765
R262 VSS.n1 VSS.n0 3.2765
R263 VSS.n47 VSS.t66 3.2765
R264 VSS.n47 VSS.n46 3.2765
R265 VSS.n45 VSS.t50 3.2765
R266 VSS.n45 VSS.n44 3.2765
R267 VSS.n3 VSS.t24 3.2765
R268 VSS.n3 VSS.n2 3.2765
R269 VSS.n16 VSS.t35 3.2765
R270 VSS.n16 VSS.n15 3.2765
R271 VSS VSS.n34 2.6005
R272 VSS.n34 VSS.n33 2.6005
R273 VSS.n38 VSS 2.6005
R274 VSS.n39 VSS.n38 2.6005
R275 VSS VSS.n27 2.6005
R276 VSS.n27 VSS.n26 2.6005
R277 VSS.n31 VSS 2.6005
R278 VSS.n32 VSS.n31 2.6005
R279 VSS.n43 VSS.n42 2.6005
R280 VSS.t10 VSS.t20 1.92472
R281 VSS.t6 VSS.t23 1.92472
R282 VSS.t7 VSS.t19 1.92472
R283 VSS.t49 VSS.t65 1.92472
R284 VSS.t45 VSS.t36 1.92472
R285 VSS.t5 VSS.t0 1.92472
R286 VSS.t0 VSS.t28 1.92472
R287 VSS.t48 VSS.t32 1.92472
R288 VSS.t32 VSS.t33 1.92472
R289 VSS.t51 VSS.t29 1.92017
R290 VSS.t62 VSS.t34 1.92017
R291 VSS.t58 VSS.t25 1.92017
R292 VSS.n10 VSS.n9 0.781777
R293 VSS.n18 VSS.n17 0.781777
R294 VSS.n20 VSS.n19 0.478105
R295 VSS.n20 VSS.n12 0.458326
R296 VSS.n38 VSS.n34 0.241879
R297 VSS.n12 VSS.n10 0.200065
R298 VSS.n19 VSS.n18 0.200065
R299 VSS.n31 VSS.n27 0.188841
R300 VSS.n21 VSS.n20 0.131118
R301 VSS VSS.n48 0.0945618
R302 VSS.n23 VSS.n22 0.0877209
R303 VSS VSS.n24 0.0231603
R304 VSS VSS.n37 0.00664458
R305 VSS VSS.n30 0.00652231
R306 VSS.n22 VSS.n21 0.000713777
R307 VSS.n24 VSS.n23 0.000713777
R308 INV_mag_1.IN.n26 INV_mag_1.IN.t15 226.316
R309 INV_mag_1.IN.n6 INV_mag_1.IN.t23 116.993
R310 INV_mag_1.IN.n31 INV_mag_1.IN.t17 33.8279
R311 INV_mag_1.IN.n32 INV_mag_1.IN.n31 30.2144
R312 INV_mag_1.IN.t27 INV_mag_1.IN.n2 25.0458
R313 INV_mag_1.IN.n29 INV_mag_1.IN.n28 16.5048
R314 INV_mag_1.IN.n30 INV_mag_1.IN.n29 16.5048
R315 INV_mag_1.IN.n2 INV_mag_1.IN.t20 15.3305
R316 INV_mag_1.IN.n4 INV_mag_1.IN.t33 15.1914
R317 INV_mag_1.IN.n2 INV_mag_1.IN.n32 12.8616
R318 INV_mag_1.IN.n4 INV_mag_1.IN.t31 12.6987
R319 INV_mag_1.IN.n5 INV_mag_1.IN.t27 12.1515
R320 INV_mag_1.IN.n7 INV_mag_1.IN.n6 11.3159
R321 INV_mag_1.IN.n26 INV_mag_1.IN.t13 10.9468
R322 INV_mag_1.IN.n6 INV_mag_1.IN.t32 10.2935
R323 INV_mag_1.IN.n0 INV_mag_1.IN.n4 10.261
R324 INV_mag_1.IN.n28 INV_mag_1.IN.t25 9.4175
R325 INV_mag_1.IN.n29 INV_mag_1.IN.t30 9.4175
R326 INV_mag_1.IN.t20 INV_mag_1.IN.n30 9.4175
R327 INV_mag_1.IN.n28 INV_mag_1.IN.t21 9.1985
R328 INV_mag_1.IN.n29 INV_mag_1.IN.t28 9.1985
R329 INV_mag_1.IN.n30 INV_mag_1.IN.t18 9.1985
R330 INV_mag_1.IN.n7 INV_mag_1.IN.t29 8.74974
R331 INV_mag_1.IN.n2 INV_mag_1.IN.t24 8.05323
R332 INV_mag_1.IN.n16 INV_mag_1.IN.n15 6.76657
R333 INV_mag_1.IN.n3 INV_mag_1.IN.n27 6.46231
R334 INV_mag_1.IN.n16 INV_mag_1.IN.n13 5.58741
R335 INV_mag_1.IN.n23 INV_mag_1.IN.n11 5.17308
R336 INV_mag_1.IN.n3 INV_mag_1.IN.n26 4.73858
R337 INV_mag_1.IN.n31 INV_mag_1.IN.t19 3.6505
R338 INV_mag_1.IN.n32 INV_mag_1.IN.t22 3.6505
R339 INV_mag_1.IN.n9 INV_mag_1.IN.t1 3.6405
R340 INV_mag_1.IN.n9 INV_mag_1.IN.n8 3.6405
R341 INV_mag_1.IN.n11 INV_mag_1.IN.t2 3.6405
R342 INV_mag_1.IN.n11 INV_mag_1.IN.n10 3.6405
R343 INV_mag_1.IN.n21 INV_mag_1.IN.t5 3.6405
R344 INV_mag_1.IN.n21 INV_mag_1.IN.n20 3.6405
R345 INV_mag_1.IN.n13 INV_mag_1.IN.t9 3.6405
R346 INV_mag_1.IN.n13 INV_mag_1.IN.n12 3.6405
R347 INV_mag_1.IN.n18 INV_mag_1.IN.t7 3.6405
R348 INV_mag_1.IN.n18 INV_mag_1.IN.n17 3.6405
R349 INV_mag_1.IN.n25 INV_mag_1.IN.t14 3.6405
R350 INV_mag_1.IN.n25 INV_mag_1.IN.n24 3.6405
R351 INV_mag_1.IN.n15 INV_mag_1.IN.t3 3.2765
R352 INV_mag_1.IN.n15 INV_mag_1.IN.n14 3.2765
R353 INV_mag_1.IN.n1 INV_mag_1.IN.n23 3.17603
R354 INV_mag_1.IN.n23 INV_mag_1.IN.n22 3.15378
R355 INV_mag_1.IN.n3 INV_mag_1.IN.n25 2.94791
R356 INV_mag_1.IN.n19 INV_mag_1.IN.n18 2.92863
R357 INV_mag_1.IN.n22 INV_mag_1.IN.n21 2.6005
R358 INV_mag_1.IN.n1 INV_mag_1.IN.n9 2.6005
R359 INV_mag_1.IN.n19 INV_mag_1.IN.n16 2.26925
R360 INV_mag_1.IN INV_mag_1.IN.n0 6.76224
R361 INV_mag_1.IN INV_mag_1.IN.n7 4.69745
R362 INV_mag_1.IN.n0 INV_mag_1.IN.n5 2.6584
R363 INV_mag_1.IN.n1 INV_mag_1.IN.n3 1.0806
R364 INV_mag_1.IN.n5 INV_mag_1.IN.n1 1.06506
R365 INV_mag_1.IN.n22 INV_mag_1.IN.n19 1.00114
R366 UP.n3 UP.n2 6.76498
R367 UP.n1 UP.t2 3.6405
R368 UP.n1 UP.n0 3.6405
R369 UP.n3 UP.n1 2.78441
R370 UP UP.n3 0.610296
R371 a_306_350.n0 a_306_350.t10 33.8126
R372 a_306_350.n1 a_306_350.n0 30.3299
R373 a_306_350.n2 a_306_350.n1 30.3299
R374 a_306_350.n3 a_306_350.n2 30.3299
R375 a_306_350.n4 a_306_350.n3 30.3299
R376 a_306_350.n5 a_306_350.n4 30.3299
R377 a_306_350.n6 a_306_350.n5 30.3299
R378 a_306_350.n7 a_306_350.n6 30.3299
R379 a_306_350.n8 a_306_350.n7 30.3299
R380 a_306_350.n13 a_306_350.t14 26.2202
R381 a_306_350.n9 a_306_350.t12 12.8368
R382 a_306_350.n9 a_306_350.n8 12.0257
R383 a_306_350.n14 a_306_350.n13 8.40022
R384 a_306_350.n12 a_306_350.n9 5.21433
R385 a_306_350.n0 a_306_350.t7 3.6505
R386 a_306_350.n1 a_306_350.t9 3.6505
R387 a_306_350.n2 a_306_350.t8 3.6505
R388 a_306_350.n3 a_306_350.t6 3.6505
R389 a_306_350.n4 a_306_350.t5 3.6505
R390 a_306_350.n5 a_306_350.t4 3.6505
R391 a_306_350.n6 a_306_350.t16 3.6505
R392 a_306_350.n7 a_306_350.t15 3.6505
R393 a_306_350.n8 a_306_350.t13 3.6505
R394 a_306_350.n13 a_306_350.t11 3.6505
R395 a_306_350.n11 a_306_350.t3 3.6405
R396 a_306_350.n11 a_306_350.n10 3.6405
R397 a_306_350.n14 a_306_350.n12 3.38916
R398 a_306_350.n15 a_306_350.t0 3.38754
R399 a_306_350.n16 a_306_350.n15 2.9777
R400 a_306_350.n15 a_306_350.n14 2.4743
R401 a_306_350.n12 a_306_350.n11 1.25598
R402 a_305_3341.n2 a_305_3341.t15 33.8126
R403 a_305_3341.n3 a_305_3341.n2 30.3299
R404 a_305_3341.n4 a_305_3341.n3 30.3299
R405 a_305_3341.n5 a_305_3341.n4 30.3299
R406 a_305_3341.n6 a_305_3341.n5 30.3299
R407 a_305_3341.n7 a_305_3341.n6 30.3299
R408 a_305_3341.n8 a_305_3341.n7 30.3299
R409 a_305_3341.n9 a_305_3341.n8 30.3299
R410 a_305_3341.n10 a_305_3341.n9 30.3299
R411 a_305_3341.n13 a_305_3341.t9 26.2932
R412 a_305_3341.n11 a_305_3341.t12 12.8368
R413 a_305_3341.n11 a_305_3341.n10 12.0257
R414 a_305_3341.n14 a_305_3341.n13 8.47283
R415 a_305_3341.n12 a_305_3341.n11 5.21433
R416 a_305_3341.n2 a_305_3341.t10 3.6505
R417 a_305_3341.n3 a_305_3341.t6 3.6505
R418 a_305_3341.n4 a_305_3341.t13 3.6505
R419 a_305_3341.n5 a_305_3341.t5 3.6505
R420 a_305_3341.n6 a_305_3341.t11 3.6505
R421 a_305_3341.n7 a_305_3341.t4 3.6505
R422 a_305_3341.n8 a_305_3341.t8 3.6505
R423 a_305_3341.n9 a_305_3341.t14 3.6505
R424 a_305_3341.n10 a_305_3341.t7 3.6505
R425 a_305_3341.n13 a_305_3341.t16 3.6505
R426 a_305_3341.n1 a_305_3341.t0 3.6405
R427 a_305_3341.n1 a_305_3341.n0 3.6405
R428 a_305_3341.n14 a_305_3341.n12 3.50583
R429 a_305_3341.n15 a_305_3341.t2 3.38777
R430 a_305_3341.n16 a_305_3341.n15 2.97653
R431 a_305_3341.n15 a_305_3341.n14 2.47455
R432 a_305_3341.n12 a_305_3341.n1 1.25598
R433 FIN.n0 FIN.t0 12.4835
R434 FIN.n2 FIN.t2 11.5345
R435 FIN.n0 FIN.t3 11.4615
R436 FIN.n1 FIN.t1 11.4615
R437 FIN.n1 FIN.n0 10.6935
R438 FIN FIN.n2 5.27048
R439 FIN.n2 FIN.n1 0.9495
R440 DOWN.n3 DOWN.n0 6.76498
R441 DOWN.n2 DOWN.t1 3.6405
R442 DOWN.n2 DOWN.n1 3.6405
R443 DOWN.n3 DOWN.n2 2.78441
R444 DOWN DOWN.n3 0.610296
R445 FDIV.n1 FDIV.n0 13.9524
R446 FDIV.n0 FDIV.t3 12.4105
R447 FDIV.n0 FDIV.t0 11.5345
R448 FDIV FDIV.n1 8.49358
R449 FDIV.n1 FDIV.t2 8.1035
R450 FDIV.n1 FDIV.t1 7.6655
C0 VDD UP 0.293f
C1 VDD a_219_1360# 0.048f
C2 INV_mag_1.IN a_1776_787# 0.354f
C3 VDD INV_mag_0.IN 4.71f
C4 INV_mag_1.IN Buffer_V_2_0.IN 0.595f
C5 VDD a_2895_3200# 0.498f
C6 FDIV a_219_2510# 3e-20
C7 INV_mag_0.OUT a_219_1360# 0.304f
C8 INV_mag_0.IN a_218_2267# 0.251f
C9 INV_mag_0.IN INV_mag_0.OUT 0.321f
C10 VDD INV_mag_1.IN 4.96f
C11 a_2895_3200# INV_mag_0.OUT 5.66e-19
C12 a_1176_1116# INV_mag_1.OUT 1.35e-20
C13 INV_mag_1.IN a_218_2267# 0.0588f
C14 INV_mag_1.IN INV_mag_0.OUT 0.219f
C15 Buffer_V_2_0.IN DOWN 0.00536f
C16 INV_mag_0.IN a_1775_2840# 0.342f
C17 VDD a_1175_2256# 0.0011f
C18 VDD DOWN 0.316f
C19 a_2895_3200# a_1775_2840# 0.00805f
C20 a_218_2267# a_1175_2256# 0.0428f
C21 a_220_1117# FDIV 0.0859f
C22 INV_mag_1.IN a_1775_2840# 0.0617f
C23 INV_mag_0.IN a_219_2510# 0.22f
C24 a_219_1360# INV_mag_1.OUT 0.037f
C25 INV_mag_0.OUT a_1175_2256# 7.19e-20
C26 UP INV_mag_1.OUT 0.00335f
C27 INV_mag_0.OUT DOWN 7.95e-19
C28 Buffer_V_2_1.IN UP 0.0051f
C29 INV_mag_0.IN INV_mag_1.OUT 0.409f
C30 VDD FIN 0.359f
C31 Buffer_V_2_1.IN INV_mag_0.IN 0.428f
C32 a_1176_1116# a_220_1117# 0.0514f
C33 a_2895_3200# INV_mag_1.OUT 0.00986f
C34 Buffer_V_2_1.IN a_2895_3200# 0.172f
C35 INV_mag_1.IN a_219_2510# 0.00927f
C36 Buffer_V_2_0.IN a_1776_787# 0.603f
C37 INV_mag_1.IN a_2896_302# 0.0341f
C38 a_218_2267# FIN 0.0424f
C39 INV_mag_1.IN INV_mag_1.OUT 0.229f
C40 INV_mag_0.OUT FIN 0.0514f
C41 Buffer_V_2_1.IN INV_mag_1.IN 0.0388f
C42 VDD a_1776_787# 0.272f
C43 VDD Buffer_V_2_0.IN 1.3f
C44 a_219_1360# FDIV 0.0426f
C45 INV_mag_0.IN FDIV 3.6e-22
C46 a_220_1117# a_219_1360# 0.145f
C47 a_1776_787# INV_mag_0.OUT 0.371f
C48 a_219_2510# a_1175_2256# 0.0514f
C49 a_2896_302# DOWN 0.13f
C50 INV_mag_0.IN a_220_1117# 1.57e-19
C51 a_1176_1116# a_219_1360# 0.0428f
C52 Buffer_V_2_0.IN INV_mag_0.OUT 0.187f
C53 INV_mag_1.OUT a_1175_2256# 0.00331f
C54 DOWN INV_mag_1.OUT 4.18e-19
C55 Buffer_V_2_1.IN a_1175_2256# 0.262f
C56 INV_mag_0.IN a_1176_1116# 0.00872f
C57 VDD a_218_2267# 0.0499f
C58 INV_mag_1.IN FDIV 0.142f
C59 VDD INV_mag_0.OUT 0.678f
C60 INV_mag_1.IN a_220_1117# 0.231f
C61 FIN a_219_2510# 0.0772f
C62 INV_mag_0.OUT a_218_2267# 0.305f
C63 INV_mag_1.IN a_1176_1116# 0.155f
C64 Buffer_V_2_1.IN FIN 0.00602f
C65 VDD a_1775_2840# 0.275f
C66 INV_mag_0.IN UP 4.32e-20
C67 INV_mag_0.IN a_219_1360# 0.0939f
C68 a_1776_787# INV_mag_1.OUT 4.79e-19
C69 a_2895_3200# UP 0.13f
C70 Buffer_V_2_0.IN a_2896_302# 0.182f
C71 a_218_2267# a_1775_2840# 0.00339f
C72 Buffer_V_2_0.IN INV_mag_1.OUT 0.0183f
C73 a_2895_3200# INV_mag_0.IN 0.0258f
C74 INV_mag_0.OUT a_1775_2840# 0.00268f
C75 INV_mag_1.IN a_219_1360# 0.196f
C76 UP INV_mag_1.IN 8.12e-19
C77 VDD a_219_2510# 0.0314f
C78 VDD a_2896_302# 0.507f
C79 INV_mag_0.IN INV_mag_1.IN 1.33f
C80 VDD INV_mag_1.OUT 0.805f
C81 VDD Buffer_V_2_1.IN 1.18f
C82 a_218_2267# a_219_2510# 0.145f
C83 a_2895_3200# INV_mag_1.IN 0.00286f
C84 a_220_1117# FIN 2.24e-20
C85 a_218_2267# INV_mag_1.OUT 0.0502f
C86 INV_mag_0.OUT a_219_2510# 0.00145f
C87 INV_mag_0.OUT a_2896_302# 0.00304f
C88 Buffer_V_2_1.IN a_218_2267# 0.0325f
C89 INV_mag_0.OUT INV_mag_1.OUT 0.482f
C90 Buffer_V_2_1.IN INV_mag_0.OUT 0.00202f
C91 Buffer_V_2_0.IN FDIV 0.00647f
C92 INV_mag_0.IN a_1175_2256# 0.145f
C93 a_220_1117# Buffer_V_2_0.IN 0.0369f
C94 VDD FDIV 0.372f
C95 a_1176_1116# Buffer_V_2_0.IN 0.262f
C96 a_1775_2840# INV_mag_1.OUT 0.0143f
C97 VDD a_220_1117# 0.0315f
C98 INV_mag_1.IN a_1175_2256# 0.017f
C99 Buffer_V_2_1.IN a_1775_2840# 0.619f
C100 a_218_2267# FDIV 5.53e-20
C101 a_219_1360# FIN 3.78e-20
C102 INV_mag_1.IN DOWN 0.00201f
C103 VDD a_1176_1116# 0.0011f
C104 INV_mag_0.IN FIN 0.134f
C105 INV_mag_0.OUT FDIV 0.0514f
C106 a_220_1117# INV_mag_0.OUT 0.00219f
C107 INV_mag_1.OUT a_219_2510# 7.65e-19
C108 a_2896_302# INV_mag_1.OUT 6.07e-19
C109 Buffer_V_2_1.IN a_219_2510# 0.0368f
C110 a_1176_1116# INV_mag_0.OUT 0.0019f
C111 a_1776_787# a_219_1360# 0.00315f
C112 INV_mag_1.IN FIN 0.00539f
C113 Buffer_V_2_1.IN INV_mag_1.OUT 0.135f
C114 Buffer_V_2_0.IN a_219_1360# 0.038f
C115 INV_mag_0.IN a_1776_787# 0.0719f
C116 INV_mag_0.IN Buffer_V_2_0.IN 0.0412f
C117 FDIV VSS 0.581f
C118 FIN VSS 0.536f
C119 DOWN VSS 0.171f
C120 a_2896_302# VSS 0.517f
C121 a_1776_787# VSS 0.161f
C122 Buffer_V_2_0.IN VSS 1.13f
C123 a_220_1117# VSS 0.155f
C124 a_1176_1116# VSS 0.324f
C125 a_219_1360# VSS 0.707f
C126 a_218_2267# VSS 0.709f
C127 INV_mag_0.OUT VSS 3.57f
C128 a_1175_2256# VSS 0.324f
C129 a_219_2510# VSS 0.157f
C130 INV_mag_1.OUT VSS 3.13f
C131 a_1775_2840# VSS 0.157f
C132 INV_mag_1.IN VSS 3.55f
C133 UP VSS 0.171f
C134 INV_mag_0.IN VSS 3.07f
C135 a_2895_3200# VSS 0.512f
C136 Buffer_V_2_1.IN VSS 1.15f
C137 VDD VSS 27f
C138 a_305_3341.t0 VSS 0.0172f
C139 a_305_3341.n0 VSS 0.0172f
C140 a_305_3341.n1 VSS 0.0347f
C141 a_305_3341.t7 VSS 0.0205f
C142 a_305_3341.t14 VSS 0.0205f
C143 a_305_3341.t8 VSS 0.0205f
C144 a_305_3341.t4 VSS 0.0205f
C145 a_305_3341.t11 VSS 0.0205f
C146 a_305_3341.t5 VSS 0.0205f
C147 a_305_3341.t13 VSS 0.0205f
C148 a_305_3341.t6 VSS 0.0205f
C149 a_305_3341.t10 VSS 0.0205f
C150 a_305_3341.t15 VSS 0.0907f
C151 a_305_3341.n2 VSS 0.105f
C152 a_305_3341.n3 VSS 0.0937f
C153 a_305_3341.n4 VSS 0.0937f
C154 a_305_3341.n5 VSS 0.0937f
C155 a_305_3341.n6 VSS 0.0937f
C156 a_305_3341.n7 VSS 0.0937f
C157 a_305_3341.n8 VSS 0.0937f
C158 a_305_3341.n9 VSS 0.0937f
C159 a_305_3341.n10 VSS 0.0815f
C160 a_305_3341.t12 VSS 0.0681f
C161 a_305_3341.n11 VSS 0.101f
C162 a_305_3341.n12 VSS 0.4f
C163 a_305_3341.t16 VSS 0.0205f
C164 a_305_3341.t9 VSS 0.0995f
C165 a_305_3341.n13 VSS 0.166f
C166 a_305_3341.n14 VSS 0.667f
C167 a_305_3341.t2 VSS 0.0182f
C168 a_305_3341.n15 VSS 0.0552f
C169 a_305_3341.n16 VSS 0.0163f
C170 a_306_350.t13 VSS 0.0205f
C171 a_306_350.t15 VSS 0.0205f
C172 a_306_350.t16 VSS 0.0205f
C173 a_306_350.t4 VSS 0.0205f
C174 a_306_350.t5 VSS 0.0205f
C175 a_306_350.t6 VSS 0.0205f
C176 a_306_350.t8 VSS 0.0205f
C177 a_306_350.t9 VSS 0.0205f
C178 a_306_350.t7 VSS 0.0205f
C179 a_306_350.t10 VSS 0.0907f
C180 a_306_350.n0 VSS 0.105f
C181 a_306_350.n1 VSS 0.0937f
C182 a_306_350.n2 VSS 0.0937f
C183 a_306_350.n3 VSS 0.0937f
C184 a_306_350.n4 VSS 0.0937f
C185 a_306_350.n5 VSS 0.0937f
C186 a_306_350.n6 VSS 0.0937f
C187 a_306_350.n7 VSS 0.0937f
C188 a_306_350.n8 VSS 0.0815f
C189 a_306_350.t12 VSS 0.0681f
C190 a_306_350.n9 VSS 0.101f
C191 a_306_350.t3 VSS 0.0172f
C192 a_306_350.n10 VSS 0.0172f
C193 a_306_350.n11 VSS 0.0347f
C194 a_306_350.n12 VSS 0.389f
C195 a_306_350.t11 VSS 0.0205f
C196 a_306_350.t14 VSS 0.0996f
C197 a_306_350.n13 VSS 0.166f
C198 a_306_350.n14 VSS 0.679f
C199 a_306_350.t0 VSS 0.0182f
C200 a_306_350.n15 VSS 0.0552f
C201 a_306_350.n16 VSS 0.0163f
C202 INV_mag_1.IN.n0 VSS 1.41f
C203 INV_mag_1.IN.n1 VSS 0.168f
C204 INV_mag_1.IN.n2 VSS 0.11f
C205 INV_mag_1.IN.n3 VSS 0.162f
C206 INV_mag_1.IN.n4 VSS 0.329f
C207 INV_mag_1.IN.n5 VSS 0.129f
C208 INV_mag_1.IN.t32 VSS 0.0309f
C209 INV_mag_1.IN.t23 VSS 0.0685f
C210 INV_mag_1.IN.n6 VSS 0.0554f
C211 INV_mag_1.IN.t29 VSS 0.0269f
C212 INV_mag_1.IN.n7 VSS 0.0465f
C213 INV_mag_1.IN.t31 VSS 0.0376f
C214 INV_mag_1.IN.t33 VSS 0.0413f
C215 INV_mag_1.IN.t1 VSS 0.0105f
C216 INV_mag_1.IN.n8 VSS 0.0105f
C217 INV_mag_1.IN.n9 VSS 0.021f
C218 INV_mag_1.IN.t2 VSS 0.0105f
C219 INV_mag_1.IN.n10 VSS 0.0105f
C220 INV_mag_1.IN.n11 VSS 0.0491f
C221 INV_mag_1.IN.t9 VSS 0.0105f
C222 INV_mag_1.IN.n12 VSS 0.0105f
C223 INV_mag_1.IN.n13 VSS 0.0554f
C224 INV_mag_1.IN.t3 VSS 0.0105f
C225 INV_mag_1.IN.n14 VSS 0.0105f
C226 INV_mag_1.IN.n15 VSS 0.0638f
C227 INV_mag_1.IN.n16 VSS 0.32f
C228 INV_mag_1.IN.t7 VSS 0.0105f
C229 INV_mag_1.IN.n17 VSS 0.0105f
C230 INV_mag_1.IN.n18 VSS 0.0226f
C231 INV_mag_1.IN.n19 VSS 0.109f
C232 INV_mag_1.IN.t5 VSS 0.0105f
C233 INV_mag_1.IN.n20 VSS 0.0105f
C234 INV_mag_1.IN.n21 VSS 0.021f
C235 INV_mag_1.IN.n22 VSS 0.124f
C236 INV_mag_1.IN.n23 VSS 0.249f
C237 INV_mag_1.IN.t14 VSS 0.0105f
C238 INV_mag_1.IN.n24 VSS 0.0105f
C239 INV_mag_1.IN.n25 VSS 0.0254f
C240 INV_mag_1.IN.t15 VSS 0.067f
C241 INV_mag_1.IN.t13 VSS 0.0321f
C242 INV_mag_1.IN.n26 VSS 0.0397f
C243 INV_mag_1.IN.n27 VSS 0.0221f
C244 INV_mag_1.IN.t21 VSS 0.0279f
C245 INV_mag_1.IN.t25 VSS 0.0285f
C246 INV_mag_1.IN.n28 VSS 0.0612f
C247 INV_mag_1.IN.t28 VSS 0.0279f
C248 INV_mag_1.IN.t30 VSS 0.0285f
C249 INV_mag_1.IN.n29 VSS 0.0708f
C250 INV_mag_1.IN.t18 VSS 0.0279f
C251 INV_mag_1.IN.n30 VSS 0.0612f
C252 INV_mag_1.IN.t20 VSS 0.0685f
C253 INV_mag_1.IN.t24 VSS 0.0247f
C254 INV_mag_1.IN.t22 VSS 0.0125f
C255 INV_mag_1.IN.t19 VSS 0.0125f
C256 INV_mag_1.IN.t17 VSS 0.0555f
C257 INV_mag_1.IN.n31 VSS 0.0645f
C258 INV_mag_1.IN.n32 VSS 0.0491f
C259 INV_mag_1.IN.t27 VSS 0.0873f
C260 VDD.t5 VSS 0.00328f
C261 VDD.n0 VSS 0.00328f
C262 VDD.n1 VSS 0.0084f
C263 VDD.t101 VSS 0.00328f
C264 VDD.n2 VSS 0.00328f
C265 VDD.n3 VSS 0.0084f
C266 VDD.t103 VSS 0.00328f
C267 VDD.n4 VSS 0.00328f
C268 VDD.n5 VSS 0.00657f
C269 VDD.n6 VSS 0.00303f
C270 VDD.t34 VSS 0.0035f
C271 VDD.n7 VSS 0.0305f
C272 VDD.n8 VSS 0.0569f
C273 VDD.t66 VSS 0.00706f
C274 VDD.t19 VSS 0.00328f
C275 VDD.n9 VSS 0.00328f
C276 VDD.n10 VSS 0.00727f
C277 VDD.n11 VSS 0.00704f
C278 VDD.n12 VSS 0.00721f
C279 VDD.t76 VSS 0.296f
C280 VDD.t74 VSS 0.132f
C281 VDD.t56 VSS 0.447f
C282 VDD.t0 VSS 0.28f
C283 VDD.t23 VSS 0.28f
C284 VDD.t39 VSS 0.28f
C285 VDD.t21 VSS 0.28f
C286 VDD.t31 VSS 0.28f
C287 VDD.t42 VSS 0.28f
C288 VDD.t104 VSS 0.232f
C289 VDD.t12 VSS 0.134f
C290 VDD.t112 VSS 0.14f
C291 VDD.t53 VSS 0.14f
C292 VDD.t93 VSS 0.14f
C293 VDD.t28 VSS 0.14f
C294 VDD.t108 VSS 0.14f
C295 VDD.t20 VSS 0.318f
C296 VDD.t44 VSS 0.257f
C297 VDD.t46 VSS 0.147f
C298 VDD.n13 VSS 0.137f
C299 VDD.t75 VSS 0.00328f
C300 VDD.n14 VSS 0.00328f
C301 VDD.n15 VSS 0.00789f
C302 VDD.t45 VSS 0.00745f
C303 VDD.t109 VSS 0.00328f
C304 VDD.n16 VSS 0.00328f
C305 VDD.n17 VSS 0.00657f
C306 VDD.n18 VSS 0.00303f
C307 VDD.t54 VSS 0.0035f
C308 VDD.n19 VSS 0.0305f
C309 VDD.n20 VSS 0.0569f
C310 VDD.t113 VSS 0.00328f
C311 VDD.n21 VSS 0.00328f
C312 VDD.n22 VSS 0.00841f
C313 VDD.t111 VSS 0.00328f
C314 VDD.n23 VSS 0.00328f
C315 VDD.n24 VSS 0.00841f
C316 VDD.t110 VSS 0.00328f
C317 VDD.n25 VSS 0.00328f
C318 VDD.n26 VSS 0.00841f
C319 VDD.t107 VSS 0.00328f
C320 VDD.n27 VSS 0.00328f
C321 VDD.n28 VSS 0.00657f
C322 VDD.t24 VSS 0.00328f
C323 VDD.n29 VSS 0.00328f
C324 VDD.n30 VSS 0.00693f
C325 VDD.t22 VSS 0.00328f
C326 VDD.n31 VSS 0.00328f
C327 VDD.n32 VSS 0.00693f
C328 VDD.t43 VSS 0.00328f
C329 VDD.n33 VSS 0.00328f
C330 VDD.n34 VSS 0.0107f
C331 VDD.n35 VSS 0.0458f
C332 VDD.n36 VSS 0.0275f
C333 VDD.n37 VSS 0.0144f
C334 VDD.t98 VSS 0.00655f
C335 VDD.t57 VSS 0.00835f
C336 VDD.n38 VSS 0.063f
C337 VDD.n39 VSS 0.242f
C338 VDD.n40 VSS 0.156f
C339 VDD.n41 VSS 0.156f
C340 VDD.n42 VSS 0.156f
C341 VDD.n43 VSS 0.151f
C342 VDD.n44 VSS 0.203f
C343 VDD.n45 VSS 0.109f
C344 VDD.n46 VSS 0.0488f
C345 VDD.n47 VSS 0.199f
C346 VDD.n48 VSS 0.0072f
C347 VDD.t36 VSS 0.333f
C348 VDD.t29 VSS 0.32f
C349 VDD.n49 VSS 0.168f
C350 VDD.t30 VSS 0.00718f
C351 VDD.t52 VSS 0.00718f
C352 VDD.n50 VSS 0.0985f
C353 VDD.n51 VSS 0.00749f
C354 VDD.n52 VSS 0.0713f
C355 VDD.n53 VSS 0.088f
C356 VDD.n54 VSS 0.784f
C357 VDD.n55 VSS 0.392f
C358 VDD.t15 VSS 0.266f
C359 VDD.t18 VSS 0.118f
C360 VDD.t3 VSS 0.241f
C361 VDD.t65 VSS 0.194f
C362 VDD.t62 VSS 0.132f
C363 VDD.n56 VSS 0.127f
C364 VDD.n57 VSS 0.048f
C365 VDD.n58 VSS 0.096f
C366 VDD.n59 VSS 0.187f
C367 VDD.n60 VSS 0.179f
C368 VDD.n61 VSS 0.181f
C369 VDD.n62 VSS 0.123f
C370 VDD.n63 VSS 0.145f
C371 VDD.t102 VSS 0.146f
C372 VDD.t79 VSS 0.146f
C373 VDD.t6 VSS 0.146f
C374 VDD.t33 VSS 0.146f
C375 VDD.t100 VSS 0.146f
C376 VDD.t25 VSS 0.14f
C377 VDD.t9 VSS 0.243f
C378 VDD.t4 VSS 0.292f
C379 VDD.t71 VSS 0.161f
C380 VDD.t88 VSS 0.466f
C381 VDD.t90 VSS 0.292f
C382 VDD.t80 VSS 0.292f
C383 VDD.t49 VSS 0.292f
C384 VDD.t67 VSS 0.277f
C385 VDD.n64 VSS 0.146f
C386 VDD.n65 VSS 0.157f
C387 VDD.t82 VSS 0.00328f
C388 VDD.n66 VSS 0.00328f
C389 VDD.n67 VSS 0.0084f
C390 VDD.t81 VSS 0.00328f
C391 VDD.n68 VSS 0.00328f
C392 VDD.n69 VSS 0.00693f
C393 VDD.t68 VSS 0.00328f
C394 VDD.n70 VSS 0.00328f
C395 VDD.n71 VSS 0.00693f
C396 VDD.t55 VSS 0.00328f
C397 VDD.n72 VSS 0.00328f
C398 VDD.n73 VSS 0.0107f
C399 VDD.n74 VSS 0.0458f
C400 VDD.n75 VSS 0.0275f
C401 VDD.t85 VSS 0.00328f
C402 VDD.n76 VSS 0.00328f
C403 VDD.n77 VSS 0.00657f
C404 VDD.n78 VSS 0.0143f
C405 VDD.t99 VSS 0.00835f
C406 VDD.t89 VSS 0.00655f
C407 VDD.n79 VSS 0.0637f
C408 VDD.n80 VSS 0.286f
C409 VDD.n81 VSS 0.156f
C410 INV_mag_0.IN.n0 VSS 0.166f
C411 INV_mag_0.IN.n1 VSS 0.115f
C412 INV_mag_0.IN.n2 VSS 0.21f
C413 INV_mag_0.IN.t21 VSS 0.0324f
C414 INV_mag_0.IN.t20 VSS 0.0717f
C415 INV_mag_0.IN.n3 VSS 0.058f
C416 INV_mag_0.IN.t25 VSS 0.0282f
C417 INV_mag_0.IN.n4 VSS 0.0487f
C418 INV_mag_0.IN.t24 VSS 0.0395f
C419 INV_mag_0.IN.t28 VSS 0.0432f
C420 INV_mag_0.IN.n5 VSS 0.168f
C421 INV_mag_0.IN.n6 VSS 0.128f
C422 INV_mag_0.IN.t7 VSS 0.011f
C423 INV_mag_0.IN.n7 VSS 0.011f
C424 INV_mag_0.IN.n8 VSS 0.0625f
C425 INV_mag_0.IN.t8 VSS 0.011f
C426 INV_mag_0.IN.n9 VSS 0.011f
C427 INV_mag_0.IN.n10 VSS 0.022f
C428 INV_mag_0.IN.t5 VSS 0.011f
C429 INV_mag_0.IN.n11 VSS 0.011f
C430 INV_mag_0.IN.n12 VSS 0.058f
C431 INV_mag_0.IN.t0 VSS 0.011f
C432 INV_mag_0.IN.n13 VSS 0.011f
C433 INV_mag_0.IN.n14 VSS 0.0668f
C434 INV_mag_0.IN.n15 VSS 0.335f
C435 INV_mag_0.IN.t6 VSS 0.011f
C436 INV_mag_0.IN.n16 VSS 0.011f
C437 INV_mag_0.IN.n17 VSS 0.0237f
C438 INV_mag_0.IN.n18 VSS 0.114f
C439 INV_mag_0.IN.n19 VSS 0.13f
C440 INV_mag_0.IN.n20 VSS 0.265f
C441 INV_mag_0.IN.t10 VSS 0.011f
C442 INV_mag_0.IN.n21 VSS 0.011f
C443 INV_mag_0.IN.n22 VSS 0.022f
C444 INV_mag_0.IN.n23 VSS 0.0232f
C445 INV_mag_0.IN.t3 VSS 0.0701f
C446 INV_mag_0.IN.t1 VSS 0.0334f
C447 INV_mag_0.IN.n24 VSS 0.0418f
C448 INV_mag_0.IN.t2 VSS 0.011f
C449 INV_mag_0.IN.n25 VSS 0.011f
C450 INV_mag_0.IN.n26 VSS 0.0266f
C451 INV_mag_0.IN.t22 VSS 0.0258f
C452 INV_mag_0.IN.t31 VSS 0.0131f
C453 INV_mag_0.IN.t18 VSS 0.0131f
C454 INV_mag_0.IN.t29 VSS 0.0582f
C455 INV_mag_0.IN.n27 VSS 0.0675f
C456 INV_mag_0.IN.n28 VSS 0.0515f
C457 INV_mag_0.IN.t30 VSS 0.0298f
C458 INV_mag_0.IN.t19 VSS 0.0292f
C459 INV_mag_0.IN.n29 VSS 0.064f
C460 INV_mag_0.IN.t33 VSS 0.0298f
C461 INV_mag_0.IN.t23 VSS 0.0292f
C462 INV_mag_0.IN.n30 VSS 0.0742f
C463 INV_mag_0.IN.t32 VSS 0.0292f
C464 INV_mag_0.IN.n31 VSS 0.064f
C465 INV_mag_0.IN.t27 VSS 0.0717f
C466 INV_mag_0.IN.t17 VSS 0.0914f
C467 INV_mag_0.IN.n32 VSS 1.19f
.ends

