* NGSPICE file created from LF_mag.ext - technology: gf180mcuC

.subckt mim_2p0fF_WS3THJ m4_n4490_n4370# m4_n4370_n4250#
X0 m4_n4370_n4250# m4_n4490_n4370# cap_mim_2f0_m4m5_noshield c_width=42.5u c_length=42.5u
.ends

.subckt cap3p_layout Pp Nn
Xmim_2p0fF_WS3THJ_0 Nn Pp mim_2p0fF_WS3THJ
.ends

.subckt ppolyf_u_TPG873 a_1000_n1102# a_280_1000# a_n440_1000# a_n920_n1102# a_n440_n1102#
+ a_520_n1102# a_40_1000# a_n200_1000# a_n1160_1000# a_n200_n1102# a_n1160_n1102#
+ w_n1344_n1286# a_1000_1000# a_760_1000# a_n680_n1102# a_n920_1000# a_760_n1102#
+ a_520_1000# a_280_n1102# a_n680_1000# a_40_n1102#
X0 a_n680_1000# a_n680_n1102# w_n1344_n1286# ppolyf_u r_width=0.8u r_length=10u
X1 a_n920_1000# a_n920_n1102# w_n1344_n1286# ppolyf_u r_width=0.8u r_length=10u
X2 a_280_1000# a_280_n1102# w_n1344_n1286# ppolyf_u r_width=0.8u r_length=10u
X3 a_520_1000# a_520_n1102# w_n1344_n1286# ppolyf_u r_width=0.8u r_length=10u
X4 a_40_1000# a_40_n1102# w_n1344_n1286# ppolyf_u r_width=0.8u r_length=10u
X5 a_n1160_1000# a_n1160_n1102# w_n1344_n1286# ppolyf_u r_width=0.8u r_length=10u
X6 a_760_1000# a_760_n1102# w_n1344_n1286# ppolyf_u r_width=0.8u r_length=10u
X7 a_1000_1000# a_1000_n1102# w_n1344_n1286# ppolyf_u r_width=0.8u r_length=10u
X8 a_n200_1000# a_n200_n1102# w_n1344_n1286# ppolyf_u r_width=0.8u r_length=10u
X9 a_n440_1000# a_n440_n1102# w_n1344_n1286# ppolyf_u r_width=0.8u r_length=10u
.ends

.subckt res_48k_mag A B VDD
Xppolyf_u_TPG873_0 m1_n2577_205# m1_n3297_2306# m1_n3777_2306# m1_n4497_204# m1_n4017_204#
+ m1_n3057_204# m1_n3297_2306# m1_n3777_2306# A m1_n3537_204# m1_n4497_204# VDD B
+ m1_n2817_2306# m1_n4017_204# m1_n4257_2306# m1_n2577_205# m1_n2817_2306# m1_n3057_204#
+ m1_n4257_2306# m1_n3537_204# ppolyf_u_TPG873
.ends

.subckt mim_2p0fF_Q67PCK m4_5681_n21380# m4_11295_n21380# m4_n16775_n21380# m4_n22389_n21380#
+ m4_n11041_n21260# m4_17029_n21260# m4_5801_n21260# m4_11415_n21260# m4_67_n21380#
+ m4_n16655_n21260# m4_187_n21260# m4_n5547_n21380# m4_n22269_n21260# m4_16909_n21380#
+ m4_n11161_n21380# m4_n5427_n21260#
X0 m4_5801_n21260# m4_5681_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X1 m4_187_n21260# m4_67_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X2 m4_187_n21260# m4_67_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X3 m4_n11041_n21260# m4_n11161_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X4 m4_17029_n21260# m4_16909_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X5 m4_17029_n21260# m4_16909_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X6 m4_n5427_n21260# m4_n5547_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X7 m4_17029_n21260# m4_16909_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X8 m4_n22269_n21260# m4_n22389_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X9 m4_n16655_n21260# m4_n16775_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X10 m4_11415_n21260# m4_11295_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X11 m4_n22269_n21260# m4_n22389_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X12 m4_11415_n21260# m4_11295_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X13 m4_n16655_n21260# m4_n16775_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X14 m4_n11041_n21260# m4_n11161_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X15 m4_5801_n21260# m4_5681_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X16 m4_17029_n21260# m4_16909_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X17 m4_5801_n21260# m4_5681_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X18 m4_n22269_n21260# m4_n22389_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X19 m4_n16655_n21260# m4_n16775_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X20 m4_5801_n21260# m4_5681_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X21 m4_n5427_n21260# m4_n5547_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X22 m4_n5427_n21260# m4_n5547_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X23 m4_n11041_n21260# m4_n11161_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X24 m4_n11041_n21260# m4_n11161_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X25 m4_187_n21260# m4_67_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X26 m4_n5427_n21260# m4_n5547_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X27 m4_n16655_n21260# m4_n16775_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X28 m4_5801_n21260# m4_5681_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X29 m4_n22269_n21260# m4_n22389_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X30 m4_11415_n21260# m4_11295_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X31 m4_n5427_n21260# m4_n5547_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X32 m4_n22269_n21260# m4_n22389_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X33 m4_n5427_n21260# m4_n5547_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X34 m4_n16655_n21260# m4_n16775_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X35 m4_11415_n21260# m4_11295_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X36 m4_n22269_n21260# m4_n22389_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X37 m4_n11041_n21260# m4_n11161_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X38 m4_187_n21260# m4_67_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X39 m4_17029_n21260# m4_16909_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X40 m4_n11041_n21260# m4_n11161_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X41 m4_187_n21260# m4_67_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X42 m4_187_n21260# m4_67_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X43 m4_5801_n21260# m4_5681_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X44 m4_n22269_n21260# m4_n22389_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X45 m4_17029_n21260# m4_16909_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X46 m4_n16655_n21260# m4_n16775_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X47 m4_17029_n21260# m4_16909_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X48 m4_n11041_n21260# m4_n11161_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X49 m4_17029_n21260# m4_16909_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X50 m4_n11041_n21260# m4_n11161_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X51 m4_5801_n21260# m4_5681_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X52 m4_5801_n21260# m4_5681_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X53 m4_11415_n21260# m4_11295_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X54 m4_n16655_n21260# m4_n16775_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X55 m4_n16655_n21260# m4_n16775_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X56 m4_11415_n21260# m4_11295_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X57 m4_n5427_n21260# m4_n5547_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X58 m4_n5427_n21260# m4_n5547_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X59 m4_11415_n21260# m4_11295_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X60 m4_187_n21260# m4_67_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X61 m4_187_n21260# m4_67_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X62 m4_n22269_n21260# m4_n22389_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X63 m4_11415_n21260# m4_11295_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
.ends

.subckt cap80p_mag P N
Xmim_2p0fF_Q67PCK_0 N N N N P P P P N P P N P N N P mim_2p0fF_Q67PCK
.ends

.subckt LF_mag VCNTL VSS VDD
Xcap3p_layout_0 VCNTL VSS cap3p_layout
Xres_48k_mag_0 VCNTL cap80p_mag_0/P VDD res_48k_mag
Xcap80p_mag_0 cap80p_mag_0/P VSS cap80p_mag
.ends

