magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2750 -2045 2750 2045
<< psubdiff >>
rect -750 23 750 45
rect -750 -23 -728 23
rect 728 -23 750 23
rect -750 -45 750 -23
<< psubdiffcont >>
rect -728 -23 728 23
<< metal1 >>
rect -739 23 739 34
rect -739 -23 -728 23
rect 728 -23 739 23
rect -739 -34 739 -23
<< end >>
