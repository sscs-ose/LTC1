magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1461 1019 1461
<< metal1 >>
rect -19 455 19 461
rect -19 -455 -13 455
rect 13 -455 19 455
rect -19 -461 19 -455
<< via1 >>
rect -13 -455 13 455
<< metal2 >>
rect -19 455 19 461
rect -19 -455 -13 455
rect 13 -455 19 455
rect -19 -461 19 -455
<< end >>
