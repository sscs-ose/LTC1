** sch_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_MUX/TB_TOP_MUX.sch
**.subckt TB_TOP_MUX
V1 VSS GND 0
.save i(v1)
V2 VDD1 VSS 3.3
.save i(v2)
V3 VCTRL2 VSS 3.3
.save i(v3)
V4 VCTRL_IN VSS 1
.save i(v4)
V5 DIV_OUT1 VSS pulse(0 3.3 200n 100p 100p 500n 1000n)
.save i(v5)
V6 F_IN VSS pulse(0 3.3 0 100p 100p 500n 1000n)
.save i(v6)
I1 ITAIL VSS 20u
I4 VDD ITAIL1 20u
V8 S1 VSS 0
.save i(v8)
V9 S2 VSS 0
.save i(v9)
V10 S3 VSS 0
.save i(v10)
V11 S4 VSS 0
.save i(v11)
V12 S6 VSS 0
.save i(v12)
V7 PRE_SCALAR VSS pulse(0 3.3 0 100p 100p 0.5u 1u)
.save i(v7)
V13 DN_INPUT VSS pulse(0 3.3 10n 100p 100p 500n 1000n)
.save i(v13)
V14 UP_INPUT VSS pulse(0 3.3 0 100p 100p 500n 1000n)
.save i(v14)
V15 VDD VSS PWL(0 0 0.1US 0 0.101US 3.3)
.save i(v15)
x2 UP_INPUT VDD DN_INPUT VSS PRE_SCALAR UP F_IN DN ITAIL DIV_OUT S1 ITAIL1 VCTRL_IN S6 VCTRL2 S2 OUT
+ S3 S4 OUTB LF_OFFCHIP S5 pex_PLL_TOP_MUX_2
C1 LF_OFFCHIP VSS 11.27p m=1
R1 LF_OFFCHIP net1 74k m=1
C2 net1 VSS 239p m=1
V16 S5 VSS 0
.save i(v16)
x6 VDD1 net2 VDD net3 VDD net4 VSS VSS net5 net6 VSS VSS net7 VDD net8 net9 OUTB VSS DIV_OUT net10
+ 7b_divider_pex
**** begin user architecture code


.include pex_7b_divider_magic.spice
.include pex_PLL_TOP_MUX_2.spice
.include Tappered-Buffer_1_pex.spice
.control
save out  outb  x2.up1  x2.dn1  x2.vco_dff_c_0.vctrl.t35  div_out  f_in  pre_scalar

tran 300n 50u

write TB_TOP_MUX.raw
.endc



.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice res_typical
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice cap_mim
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice moscap_typical
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice mimcap_typical

**** end user architecture code
**.ends
.GLOBAL GND
.end
