magic
tech gf180mcuC
magscale 1 10
timestamp 1698512721
<< nwell >>
rect 61 2680 2865 2894
rect 1120 2594 1326 2595
rect 1440 2594 1486 2595
rect 2125 2538 2126 2640
rect 2080 2537 2126 2538
rect 1440 1438 1486 1541
rect 260 1398 664 1399
rect 61 1087 664 1398
rect 61 573 260 1087
<< pwell >>
rect 1280 120 1646 144
<< pdiff >>
rect 2125 2538 2126 2544
rect 2080 2537 2126 2538
rect 1440 1528 1486 1541
<< psubdiff >>
rect 111 -73 2815 -60
rect 111 -119 124 -73
rect 170 -119 218 -73
rect 264 -119 312 -73
rect 358 -119 406 -73
rect 452 -119 500 -73
rect 546 -119 594 -73
rect 640 -119 688 -73
rect 734 -119 782 -73
rect 828 -119 876 -73
rect 922 -119 970 -73
rect 1016 -119 1064 -73
rect 1110 -119 1158 -73
rect 1204 -119 1252 -73
rect 1298 -119 1346 -73
rect 1392 -119 1440 -73
rect 1486 -119 1534 -73
rect 1580 -119 1628 -73
rect 1674 -119 1722 -73
rect 1768 -119 1816 -73
rect 1862 -119 1910 -73
rect 1956 -119 2004 -73
rect 2050 -119 2098 -73
rect 2144 -119 2192 -73
rect 2238 -119 2286 -73
rect 2332 -119 2380 -73
rect 2426 -119 2474 -73
rect 2520 -119 2568 -73
rect 2614 -119 2662 -73
rect 2708 -119 2756 -73
rect 2802 -119 2815 -73
rect 111 -132 2815 -119
<< nsubdiff >>
rect 111 2857 2815 2870
rect 111 2811 124 2857
rect 170 2811 218 2857
rect 264 2811 312 2857
rect 358 2811 406 2857
rect 452 2811 500 2857
rect 546 2811 594 2857
rect 640 2811 688 2857
rect 734 2811 782 2857
rect 828 2811 876 2857
rect 922 2811 970 2857
rect 1016 2811 1064 2857
rect 1110 2811 1158 2857
rect 1204 2811 1252 2857
rect 1298 2811 1346 2857
rect 1392 2811 1440 2857
rect 1486 2811 1534 2857
rect 1580 2811 1628 2857
rect 1674 2811 1722 2857
rect 1768 2811 1816 2857
rect 1862 2811 1910 2857
rect 1956 2811 2004 2857
rect 2050 2811 2098 2857
rect 2144 2811 2192 2857
rect 2238 2811 2286 2857
rect 2332 2811 2380 2857
rect 2426 2811 2474 2857
rect 2520 2811 2568 2857
rect 2614 2811 2662 2857
rect 2708 2811 2756 2857
rect 2802 2811 2815 2857
rect 111 2798 2815 2811
<< psubdiffcont >>
rect 124 -119 170 -73
rect 218 -119 264 -73
rect 312 -119 358 -73
rect 406 -119 452 -73
rect 500 -119 546 -73
rect 594 -119 640 -73
rect 688 -119 734 -73
rect 782 -119 828 -73
rect 876 -119 922 -73
rect 970 -119 1016 -73
rect 1064 -119 1110 -73
rect 1158 -119 1204 -73
rect 1252 -119 1298 -73
rect 1346 -119 1392 -73
rect 1440 -119 1486 -73
rect 1534 -119 1580 -73
rect 1628 -119 1674 -73
rect 1722 -119 1768 -73
rect 1816 -119 1862 -73
rect 1910 -119 1956 -73
rect 2004 -119 2050 -73
rect 2098 -119 2144 -73
rect 2192 -119 2238 -73
rect 2286 -119 2332 -73
rect 2380 -119 2426 -73
rect 2474 -119 2520 -73
rect 2568 -119 2614 -73
rect 2662 -119 2708 -73
rect 2756 -119 2802 -73
<< nsubdiffcont >>
rect 124 2811 170 2857
rect 218 2811 264 2857
rect 312 2811 358 2857
rect 406 2811 452 2857
rect 500 2811 546 2857
rect 594 2811 640 2857
rect 688 2811 734 2857
rect 782 2811 828 2857
rect 876 2811 922 2857
rect 970 2811 1016 2857
rect 1064 2811 1110 2857
rect 1158 2811 1204 2857
rect 1252 2811 1298 2857
rect 1346 2811 1392 2857
rect 1440 2811 1486 2857
rect 1534 2811 1580 2857
rect 1628 2811 1674 2857
rect 1722 2811 1768 2857
rect 1816 2811 1862 2857
rect 1910 2811 1956 2857
rect 2004 2811 2050 2857
rect 2098 2811 2144 2857
rect 2192 2811 2238 2857
rect 2286 2811 2332 2857
rect 2380 2811 2426 2857
rect 2474 2811 2520 2857
rect 2568 2811 2614 2857
rect 2662 2811 2708 2857
rect 2756 2811 2802 2857
<< polysilicon >>
rect 235 2570 2691 2626
rect 235 1768 291 2296
rect 395 1768 451 2296
rect 555 1768 611 2296
rect 715 1768 771 2296
rect 875 1768 931 2296
rect 1035 1768 1091 2296
rect 1195 1768 1251 2296
rect 1355 1768 1411 2296
rect 1515 1768 1571 2296
rect 1675 1768 1731 2296
rect 1835 1768 1891 2296
rect 1995 1768 2051 2296
rect 2155 1768 2211 2296
rect 2315 1768 2371 2296
rect 2475 1768 2531 2296
rect 2635 1768 2691 2296
rect 235 1346 291 1534
rect 227 1333 299 1346
rect 227 1287 240 1333
rect 286 1287 299 1333
rect 227 1274 299 1287
rect 163 537 235 545
rect 163 532 741 537
rect 163 486 176 532
rect 222 486 741 532
rect 163 481 741 486
rect 163 473 235 481
rect 685 168 741 481
rect 875 432 931 960
rect 1035 432 1091 960
rect 1195 432 1251 960
rect 1355 432 1411 960
rect 1515 432 1571 960
rect 1675 432 1731 960
rect 1835 432 1891 960
rect 1995 432 2051 960
rect 685 112 2051 168
<< polycontact >>
rect 240 1287 286 1333
rect 176 486 222 532
<< metal1 >>
rect 61 2857 2865 2890
rect 61 2811 124 2857
rect 170 2811 218 2857
rect 264 2811 312 2857
rect 358 2811 406 2857
rect 452 2811 500 2857
rect 546 2811 594 2857
rect 640 2811 688 2857
rect 734 2811 782 2857
rect 828 2811 876 2857
rect 922 2811 970 2857
rect 1016 2811 1064 2857
rect 1110 2811 1158 2857
rect 1204 2811 1252 2857
rect 1298 2811 1346 2857
rect 1392 2811 1440 2857
rect 1486 2811 1534 2857
rect 1580 2811 1628 2857
rect 1674 2811 1722 2857
rect 1768 2811 1816 2857
rect 1862 2811 1910 2857
rect 1956 2811 2004 2857
rect 2050 2811 2098 2857
rect 2144 2811 2192 2857
rect 2238 2811 2286 2857
rect 2332 2811 2380 2857
rect 2426 2811 2474 2857
rect 2520 2811 2568 2857
rect 2614 2811 2662 2857
rect 2708 2811 2756 2857
rect 2802 2811 2865 2857
rect 61 2778 2865 2811
rect 160 2686 1166 2732
rect 160 2537 206 2686
rect 1120 2640 1166 2686
rect 1440 2686 2446 2732
rect 1440 2640 1486 2686
rect 2400 2640 2446 2686
rect 320 2594 1006 2640
rect 320 2537 366 2594
rect 640 2537 686 2594
rect 960 2537 1006 2594
rect 1120 2594 1486 2640
rect 1120 2537 1166 2594
rect 1440 2537 1486 2594
rect 1600 2594 2286 2640
rect 1600 2537 1646 2594
rect 1920 2537 1966 2594
rect 2240 2537 2286 2594
rect 2400 2594 2766 2640
rect 2400 2537 2446 2594
rect 1920 2519 1966 2520
rect 2720 2500 2766 2594
rect 160 1747 206 2326
rect 320 1747 366 2326
rect 480 1747 526 2326
rect 640 1747 686 2326
rect 160 1484 206 1558
rect 480 1484 526 1558
rect 160 1438 526 1484
rect 229 1333 297 1344
rect 229 1287 240 1333
rect 286 1287 297 1333
rect 229 1276 297 1287
rect 480 1300 526 1438
rect 640 1392 686 1582
rect 800 1484 846 2330
rect 960 1541 1006 2330
rect 1120 1484 1166 2330
rect 800 1438 1166 1484
rect 1280 1392 1326 2330
rect 1440 1484 1486 2330
rect 1600 1541 1646 2330
rect 1760 1484 1806 2330
rect 1440 1438 1806 1484
rect 1920 1392 1966 2330
rect 2080 1484 2126 2330
rect 2240 1747 2286 2326
rect 2400 1484 2446 2330
rect 2560 1747 2606 2326
rect 2720 1765 2766 2330
rect 2080 1438 2447 1484
rect 2560 1392 2606 1541
rect 640 1346 2717 1392
rect 240 1221 286 1276
rect 480 1254 1166 1300
rect 168 1175 286 1221
rect 168 659 214 1175
rect 260 994 664 1106
rect 168 613 405 659
rect 165 534 233 543
rect 45 532 233 534
rect 45 488 176 532
rect 165 486 176 488
rect 222 486 233 532
rect 165 475 233 486
rect 312 139 612 251
rect 406 -40 518 139
rect 800 52 846 1254
rect 960 144 1006 1197
rect 1120 403 1166 1254
rect 1280 144 1326 1346
rect 1440 1254 1806 1300
rect 1440 403 1486 1254
rect 1600 403 1646 1197
rect 1760 403 1806 1254
rect 1920 403 1966 1346
rect 2080 1239 2305 1285
rect 2080 403 2126 1239
rect 1600 144 1646 201
rect 960 98 1646 144
rect 1760 144 1806 201
rect 2080 144 2126 238
rect 1760 98 2126 144
rect 1760 52 1806 98
rect 800 6 1806 52
rect 61 -73 2865 -40
rect 61 -119 124 -73
rect 170 -119 218 -73
rect 264 -119 312 -73
rect 358 -119 406 -73
rect 452 -119 500 -73
rect 546 -119 594 -73
rect 640 -119 688 -73
rect 734 -119 782 -73
rect 828 -119 876 -73
rect 922 -119 970 -73
rect 1016 -119 1064 -73
rect 1110 -119 1158 -73
rect 1204 -119 1252 -73
rect 1298 -119 1346 -73
rect 1392 -119 1440 -73
rect 1486 -119 1534 -73
rect 1580 -119 1628 -73
rect 1674 -119 1722 -73
rect 1768 -119 1816 -73
rect 1862 -119 1910 -73
rect 1956 -119 2004 -73
rect 2050 -119 2098 -73
rect 2144 -119 2192 -73
rect 2238 -119 2286 -73
rect 2332 -119 2380 -73
rect 2426 -119 2474 -73
rect 2520 -119 2568 -73
rect 2614 -119 2662 -73
rect 2708 -119 2756 -73
rect 2802 -119 2865 -73
rect 61 -152 2865 -119
use Inverter_Layout  Inverter_Layout_0 ~/GF180Projects/Tapeout/Magic/Logic_Gates/Inverter
timestamp 1698512688
transform -1 0 602 0 1 263
box -62 -124 342 856
use nfet_03v3_DNGK9V  nfet_03v3_DNGK9V_0
timestamp 1698512460
transform 1 0 1463 0 1 699
box -700 -579 700 579
use pmos_3p3_QKQ23Q  pmos_3p3_QKQ23Q_0
timestamp 1691402935
transform 1 0 1463 0 1 2039
box -1402 -641 1402 641
<< labels >>
flabel metal1 2211 1262 2211 1262 0 FreeSans 320 0 0 0 VIN
port 5 nsew
flabel metal1 2628 1369 2628 1369 0 FreeSans 320 0 0 0 VOUT
port 7 nsew
flabel metal1 509 1050 509 1050 0 FreeSans 320 0 0 0 VDD
port 8 nsew
flabel metal1 462 194 462 194 0 FreeSans 320 0 0 0 VSS
port 9 nsew
flabel metal1 111 511 111 511 0 FreeSans 320 0 0 0 CLK
port 2 nsew
<< end >>
