magic
tech gf180mcuC
magscale 1 10
timestamp 1695275716
<< metal1 >>
rect 19130 45942 48057 46220
rect 19130 45607 48060 45942
rect 45035 44323 45911 44483
rect 45037 44084 45911 44323
rect 47682 44119 48060 45607
rect 45037 39647 45436 44084
rect 45740 44049 45900 44084
rect 47900 44049 48060 44119
rect 45556 41371 48244 41551
rect 45037 39597 46938 39647
rect 45037 39276 46305 39597
rect 46886 39276 46938 39597
rect 45037 39187 46938 39276
rect 45931 29867 46616 29872
rect 45820 602 46616 29867
rect 26584 45 46616 602
<< metal4 >>
rect 33253 33603 33465 33670
rect 33298 33560 33365 33603
rect 38867 33598 39079 33665
rect 44481 33600 44693 33667
rect 38932 33560 38999 33598
rect 44547 33560 44614 33600
<< metal5 >>
rect 38867 33627 39079 33634
use cap3p_layout  cap3p_layout_0
timestamp 1694760847
transform -1 0 54857 0 -1 38823
box -120 -826 8884 9253
use cap80p_mag  cap80p_mag_0
timestamp 1695275716
transform 1 0 39213 0 1 39107
box -39298 -39064 5480 6870
use res_48k_mag  res_48k_mag_0
timestamp 1693460400
transform 1 0 50236 0 1 41531
box -4680 -160 -1992 2678
<< labels >>
flabel metal1 45105 40745 45105 40745 0 FreeSans 1600 0 0 0 VCNTL
port 0 nsew
flabel metal1 39651 288 39651 288 0 FreeSans 1600 0 0 0 VSS
port 1 nsew
flabel metal1 46961 41452 46961 41452 0 FreeSans 1600 0 0 0 VDD
port 2 nsew
<< end >>
