magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2201 -9695 2201 9695
<< psubdiff >>
rect -201 7637 201 7695
rect -201 -7637 -179 7637
rect -133 -7637 -75 7637
rect -29 -7637 29 7637
rect 75 -7637 133 7637
rect 179 -7637 201 7637
rect -201 -7695 201 -7637
<< psubdiffcont >>
rect -179 -7637 -133 7637
rect -75 -7637 -29 7637
rect 29 -7637 75 7637
rect 133 -7637 179 7637
<< metal1 >>
rect -190 7637 190 7684
rect -190 -7637 -179 7637
rect -133 -7637 -75 7637
rect -29 -7637 29 7637
rect 75 -7637 133 7637
rect 179 -7637 190 7637
rect -190 -7684 190 -7637
<< end >>
