magic
tech gf180mcuC
magscale 1 10
timestamp 1690007892
<< nwell >>
rect 0 391 404 813
rect 536 391 1360 813
rect 0 372 204 391
<< pwell >>
rect 58 148 346 346
rect 536 148 824 342
rect 1072 148 1360 342
<< nmos >>
rect 174 222 230 272
rect 652 223 708 267
rect 1188 223 1244 267
<< pmos >>
rect 174 521 230 621
rect 714 528 770 572
rect 1126 528 1182 572
<< ndiff >>
rect 82 272 154 283
rect 250 272 322 283
rect 82 270 174 272
rect 82 224 95 270
rect 141 224 174 270
rect 82 222 174 224
rect 230 270 322 272
rect 230 224 263 270
rect 309 224 322 270
rect 560 268 632 281
rect 230 222 322 224
rect 82 211 154 222
rect 250 211 322 222
rect 560 222 573 268
rect 619 267 632 268
rect 728 268 800 281
rect 728 267 741 268
rect 619 223 652 267
rect 708 223 741 267
rect 619 222 632 223
rect 560 209 632 222
rect 728 222 741 223
rect 787 222 800 268
rect 728 209 800 222
rect 1096 268 1168 281
rect 1096 222 1109 268
rect 1155 267 1168 268
rect 1264 268 1336 281
rect 1264 267 1277 268
rect 1155 223 1188 267
rect 1244 223 1277 267
rect 1155 222 1168 223
rect 1096 209 1168 222
rect 1264 222 1277 223
rect 1323 222 1336 268
rect 1264 209 1336 222
<< pdiff >>
rect 86 608 174 621
rect 86 534 99 608
rect 145 534 174 608
rect 86 521 174 534
rect 230 608 318 621
rect 230 534 259 608
rect 305 534 318 608
rect 230 521 318 534
rect 622 573 694 586
rect 622 527 635 573
rect 681 572 694 573
rect 790 573 862 586
rect 790 572 803 573
rect 681 528 714 572
rect 770 528 803 572
rect 681 527 694 528
rect 622 514 694 527
rect 790 527 803 528
rect 849 527 862 573
rect 790 514 862 527
rect 1034 573 1106 586
rect 1034 527 1047 573
rect 1093 572 1106 573
rect 1202 573 1274 586
rect 1202 572 1215 573
rect 1093 528 1126 572
rect 1182 528 1215 572
rect 1093 527 1106 528
rect 1034 514 1106 527
rect 1202 527 1215 528
rect 1261 527 1274 573
rect 1202 514 1274 527
<< ndiffc >>
rect 95 224 141 270
rect 263 224 309 270
rect 573 222 619 268
rect 741 222 787 268
rect 1109 222 1155 268
rect 1277 222 1323 268
<< pdiffc >>
rect 99 534 145 608
rect 259 534 305 608
rect 635 527 681 573
rect 803 527 849 573
rect 1047 527 1093 573
rect 1215 527 1261 573
<< psubdiff >>
rect 26 78 374 91
rect 26 29 45 78
rect 354 29 374 78
rect 26 14 374 29
rect 558 80 1329 95
rect 558 34 577 80
rect 1306 34 1329 80
rect 558 19 1329 34
<< nsubdiff >>
rect 40 769 332 786
rect 40 718 60 769
rect 310 718 332 769
rect 40 701 332 718
rect 564 774 1327 789
rect 564 728 593 774
rect 1305 728 1327 774
rect 564 715 1327 728
<< psubdiffcont >>
rect 45 29 354 78
rect 577 34 1306 80
<< nsubdiffcont >>
rect 60 718 310 769
rect 593 728 1305 774
<< polysilicon >>
rect 174 621 230 665
rect 1412 664 1501 678
rect 1412 658 1425 664
rect 714 572 770 616
rect 1126 606 1425 658
rect 174 459 230 521
rect 714 473 770 528
rect 1126 572 1182 606
rect 1412 604 1425 606
rect 1488 604 1501 664
rect 1412 591 1501 604
rect 1126 484 1182 528
rect 115 445 230 459
rect 115 386 129 445
rect 192 386 230 445
rect 703 460 792 473
rect 703 400 716 460
rect 779 400 792 460
rect 703 386 792 400
rect 115 372 230 386
rect 174 272 230 372
rect 413 301 502 315
rect 413 241 426 301
rect 489 241 502 301
rect 413 228 502 241
rect 174 178 230 222
rect 451 179 496 228
rect 652 267 708 311
rect 652 179 708 223
rect 1188 267 1244 311
rect 451 132 708 179
rect 1188 188 1244 223
rect 1414 206 1503 220
rect 1414 188 1427 206
rect 1188 146 1427 188
rect 1490 146 1503 206
rect 1188 142 1503 146
rect 1414 133 1503 142
<< polycontact >>
rect 1425 604 1488 664
rect 129 386 192 445
rect 716 400 779 460
rect 426 241 489 301
rect 1427 146 1490 206
<< metal1 >>
rect 0 774 1360 813
rect 0 769 593 774
rect 0 718 60 769
rect 310 728 593 769
rect 1305 728 1360 774
rect 310 718 1360 728
rect 0 700 1360 718
rect 76 608 146 700
rect 76 534 99 608
rect 145 534 146 608
rect 76 519 146 534
rect 258 608 322 621
rect 258 534 259 608
rect 305 534 322 608
rect 440 614 527 632
rect 440 549 453 614
rect 518 576 527 614
rect 518 573 692 576
rect 518 549 635 573
rect 440 547 635 549
rect 0 445 204 453
rect 0 415 129 445
rect -23 398 129 415
rect -23 340 2 398
rect 60 386 129 398
rect 192 386 204 445
rect 60 372 204 386
rect 258 418 322 534
rect 446 527 635 547
rect 681 527 692 573
rect 446 525 692 527
rect 790 573 861 700
rect 790 527 803 573
rect 849 527 861 573
rect 790 525 861 527
rect 1035 573 1106 700
rect 1412 664 1501 678
rect 1412 604 1425 664
rect 1488 604 1501 664
rect 1412 591 1501 604
rect 1035 527 1047 573
rect 1093 527 1106 573
rect 1035 525 1106 527
rect 1204 573 1335 574
rect 1204 527 1215 573
rect 1261 527 1335 573
rect 1204 525 1335 527
rect 446 505 631 525
rect 60 340 74 372
rect -23 337 74 340
rect 258 371 459 418
rect 73 270 154 275
rect 258 270 322 371
rect 412 315 459 371
rect 412 301 502 315
rect 412 287 426 301
rect 73 224 95 270
rect 141 224 154 270
rect 252 224 263 270
rect 309 224 322 270
rect 413 241 426 287
rect 489 241 502 301
rect 413 228 502 241
rect 560 268 631 505
rect 703 460 792 473
rect 703 400 716 460
rect 779 400 792 460
rect 703 386 792 400
rect 1266 456 1335 525
rect 1266 397 1275 456
rect 1327 397 1335 456
rect 1266 268 1335 397
rect 73 113 154 224
rect 258 223 322 224
rect 560 222 573 268
rect 619 222 631 268
rect 560 221 631 222
rect 729 222 741 268
rect 787 222 801 268
rect 729 113 801 222
rect 1097 222 1109 268
rect 1155 222 1167 268
rect 1097 113 1167 222
rect 1266 222 1277 268
rect 1323 222 1335 268
rect 1266 221 1335 222
rect 1414 206 1503 220
rect 1414 146 1427 206
rect 1490 146 1503 206
rect 1414 133 1503 146
rect 0 80 1360 113
rect 0 78 577 80
rect 0 29 45 78
rect 354 34 577 78
rect 1306 34 1360 80
rect 354 29 1360 34
rect 0 0 1360 29
<< via1 >>
rect 453 549 518 614
rect 2 340 60 398
rect 1425 604 1488 664
rect 716 400 779 460
rect 1275 397 1327 456
rect 1427 146 1490 206
<< metal2 >>
rect 1412 672 1501 678
rect 453 664 1501 672
rect 453 632 1425 664
rect 440 614 1425 632
rect 440 549 453 614
rect 518 607 1425 614
rect 518 549 530 607
rect 1412 604 1425 607
rect 1488 604 1501 664
rect 1412 591 1501 604
rect 440 547 530 549
rect 703 460 792 473
rect -23 398 74 415
rect -23 340 2 398
rect 60 340 74 398
rect 703 400 716 460
rect 779 456 1339 460
rect 779 400 1275 456
rect 703 397 1275 400
rect 1327 397 1339 456
rect 703 393 1339 397
rect 703 386 792 393
rect -23 337 74 340
rect 2 202 60 337
rect 1414 206 1503 220
rect 1414 202 1427 206
rect 2 146 1427 202
rect 1490 146 1503 206
rect 2 144 1503 146
rect 1372 138 1503 144
rect 1414 133 1503 138
<< labels >>
flabel nsubdiffcont 185 744 185 744 0 FreeSans 640 0 0 0 Inverter_0.VDD
flabel psubdiffcont 199 52 199 52 0 FreeSans 640 0 0 0 Inverter_0.VSS
flabel metal1 390 386 390 386 0 FreeSans 640 0 0 0 Inverter_0.OUT
flabel via1 1451 633 1451 633 0 FreeSans 640 0 0 0 OUT
port 1 nsew
flabel via1 1301 419 1301 419 0 FreeSans 640 0 0 0 OUT_B
port 2 nsew
flabel nsubdiffcont 942 749 942 749 0 FreeSans 640 0 0 0 VDD
port 3 nsew
flabel psubdiffcont 938 56 938 56 0 FreeSans 640 0 0 0 VSS
port 4 nsew
flabel via1 29 371 29 371 0 FreeSans 640 0 0 0 VIN
port 5 nsew
<< end >>
