magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -2394 -2180 2394 2180
<< nwell >>
rect -394 -180 394 180
<< pmos >>
rect -220 -50 -52 50
rect 52 -50 220 50
<< pdiff >>
rect -308 23 -220 50
rect -308 -23 -295 23
rect -249 -23 -220 23
rect -308 -50 -220 -23
rect -52 23 52 50
rect -52 -23 -23 23
rect 23 -23 52 23
rect -52 -50 52 -23
rect 220 23 308 50
rect 220 -23 249 23
rect 295 -23 308 23
rect 220 -50 308 -23
<< pdiffc >>
rect -295 -23 -249 23
rect -23 -23 23 23
rect 249 -23 295 23
<< polysilicon >>
rect -220 50 -52 94
rect 52 50 220 94
rect -220 -94 -52 -50
rect 52 -94 220 -50
<< metal1 >>
rect -295 23 -249 48
rect -295 -48 -249 -23
rect -23 23 23 48
rect -23 -48 23 -23
rect 249 23 295 48
rect 249 -48 295 -23
<< end >>
