magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1071 -1149 1071 1149
<< metal1 >>
rect -71 143 71 149
rect -71 -143 -65 143
rect 65 -143 71 143
rect -71 -149 71 -143
<< via1 >>
rect -65 -143 65 143
<< metal2 >>
rect -71 143 71 149
rect -71 -143 -65 143
rect 65 -143 71 143
rect -71 -149 71 -143
<< end >>
