magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1877 -1349 1877 1349
<< metal3 >>
rect -877 344 877 349
rect -877 316 -872 344
rect -844 316 -806 344
rect -778 316 -740 344
rect -712 316 -674 344
rect -646 316 -608 344
rect -580 316 -542 344
rect -514 316 -476 344
rect -448 316 -410 344
rect -382 316 -344 344
rect -316 316 -278 344
rect -250 316 -212 344
rect -184 316 -146 344
rect -118 316 -80 344
rect -52 316 -14 344
rect 14 316 52 344
rect 80 316 118 344
rect 146 316 184 344
rect 212 316 250 344
rect 278 316 316 344
rect 344 316 382 344
rect 410 316 448 344
rect 476 316 514 344
rect 542 316 580 344
rect 608 316 646 344
rect 674 316 712 344
rect 740 316 778 344
rect 806 316 844 344
rect 872 316 877 344
rect -877 278 877 316
rect -877 250 -872 278
rect -844 250 -806 278
rect -778 250 -740 278
rect -712 250 -674 278
rect -646 250 -608 278
rect -580 250 -542 278
rect -514 250 -476 278
rect -448 250 -410 278
rect -382 250 -344 278
rect -316 250 -278 278
rect -250 250 -212 278
rect -184 250 -146 278
rect -118 250 -80 278
rect -52 250 -14 278
rect 14 250 52 278
rect 80 250 118 278
rect 146 250 184 278
rect 212 250 250 278
rect 278 250 316 278
rect 344 250 382 278
rect 410 250 448 278
rect 476 250 514 278
rect 542 250 580 278
rect 608 250 646 278
rect 674 250 712 278
rect 740 250 778 278
rect 806 250 844 278
rect 872 250 877 278
rect -877 212 877 250
rect -877 184 -872 212
rect -844 184 -806 212
rect -778 184 -740 212
rect -712 184 -674 212
rect -646 184 -608 212
rect -580 184 -542 212
rect -514 184 -476 212
rect -448 184 -410 212
rect -382 184 -344 212
rect -316 184 -278 212
rect -250 184 -212 212
rect -184 184 -146 212
rect -118 184 -80 212
rect -52 184 -14 212
rect 14 184 52 212
rect 80 184 118 212
rect 146 184 184 212
rect 212 184 250 212
rect 278 184 316 212
rect 344 184 382 212
rect 410 184 448 212
rect 476 184 514 212
rect 542 184 580 212
rect 608 184 646 212
rect 674 184 712 212
rect 740 184 778 212
rect 806 184 844 212
rect 872 184 877 212
rect -877 146 877 184
rect -877 118 -872 146
rect -844 118 -806 146
rect -778 118 -740 146
rect -712 118 -674 146
rect -646 118 -608 146
rect -580 118 -542 146
rect -514 118 -476 146
rect -448 118 -410 146
rect -382 118 -344 146
rect -316 118 -278 146
rect -250 118 -212 146
rect -184 118 -146 146
rect -118 118 -80 146
rect -52 118 -14 146
rect 14 118 52 146
rect 80 118 118 146
rect 146 118 184 146
rect 212 118 250 146
rect 278 118 316 146
rect 344 118 382 146
rect 410 118 448 146
rect 476 118 514 146
rect 542 118 580 146
rect 608 118 646 146
rect 674 118 712 146
rect 740 118 778 146
rect 806 118 844 146
rect 872 118 877 146
rect -877 80 877 118
rect -877 52 -872 80
rect -844 52 -806 80
rect -778 52 -740 80
rect -712 52 -674 80
rect -646 52 -608 80
rect -580 52 -542 80
rect -514 52 -476 80
rect -448 52 -410 80
rect -382 52 -344 80
rect -316 52 -278 80
rect -250 52 -212 80
rect -184 52 -146 80
rect -118 52 -80 80
rect -52 52 -14 80
rect 14 52 52 80
rect 80 52 118 80
rect 146 52 184 80
rect 212 52 250 80
rect 278 52 316 80
rect 344 52 382 80
rect 410 52 448 80
rect 476 52 514 80
rect 542 52 580 80
rect 608 52 646 80
rect 674 52 712 80
rect 740 52 778 80
rect 806 52 844 80
rect 872 52 877 80
rect -877 14 877 52
rect -877 -14 -872 14
rect -844 -14 -806 14
rect -778 -14 -740 14
rect -712 -14 -674 14
rect -646 -14 -608 14
rect -580 -14 -542 14
rect -514 -14 -476 14
rect -448 -14 -410 14
rect -382 -14 -344 14
rect -316 -14 -278 14
rect -250 -14 -212 14
rect -184 -14 -146 14
rect -118 -14 -80 14
rect -52 -14 -14 14
rect 14 -14 52 14
rect 80 -14 118 14
rect 146 -14 184 14
rect 212 -14 250 14
rect 278 -14 316 14
rect 344 -14 382 14
rect 410 -14 448 14
rect 476 -14 514 14
rect 542 -14 580 14
rect 608 -14 646 14
rect 674 -14 712 14
rect 740 -14 778 14
rect 806 -14 844 14
rect 872 -14 877 14
rect -877 -52 877 -14
rect -877 -80 -872 -52
rect -844 -80 -806 -52
rect -778 -80 -740 -52
rect -712 -80 -674 -52
rect -646 -80 -608 -52
rect -580 -80 -542 -52
rect -514 -80 -476 -52
rect -448 -80 -410 -52
rect -382 -80 -344 -52
rect -316 -80 -278 -52
rect -250 -80 -212 -52
rect -184 -80 -146 -52
rect -118 -80 -80 -52
rect -52 -80 -14 -52
rect 14 -80 52 -52
rect 80 -80 118 -52
rect 146 -80 184 -52
rect 212 -80 250 -52
rect 278 -80 316 -52
rect 344 -80 382 -52
rect 410 -80 448 -52
rect 476 -80 514 -52
rect 542 -80 580 -52
rect 608 -80 646 -52
rect 674 -80 712 -52
rect 740 -80 778 -52
rect 806 -80 844 -52
rect 872 -80 877 -52
rect -877 -118 877 -80
rect -877 -146 -872 -118
rect -844 -146 -806 -118
rect -778 -146 -740 -118
rect -712 -146 -674 -118
rect -646 -146 -608 -118
rect -580 -146 -542 -118
rect -514 -146 -476 -118
rect -448 -146 -410 -118
rect -382 -146 -344 -118
rect -316 -146 -278 -118
rect -250 -146 -212 -118
rect -184 -146 -146 -118
rect -118 -146 -80 -118
rect -52 -146 -14 -118
rect 14 -146 52 -118
rect 80 -146 118 -118
rect 146 -146 184 -118
rect 212 -146 250 -118
rect 278 -146 316 -118
rect 344 -146 382 -118
rect 410 -146 448 -118
rect 476 -146 514 -118
rect 542 -146 580 -118
rect 608 -146 646 -118
rect 674 -146 712 -118
rect 740 -146 778 -118
rect 806 -146 844 -118
rect 872 -146 877 -118
rect -877 -184 877 -146
rect -877 -212 -872 -184
rect -844 -212 -806 -184
rect -778 -212 -740 -184
rect -712 -212 -674 -184
rect -646 -212 -608 -184
rect -580 -212 -542 -184
rect -514 -212 -476 -184
rect -448 -212 -410 -184
rect -382 -212 -344 -184
rect -316 -212 -278 -184
rect -250 -212 -212 -184
rect -184 -212 -146 -184
rect -118 -212 -80 -184
rect -52 -212 -14 -184
rect 14 -212 52 -184
rect 80 -212 118 -184
rect 146 -212 184 -184
rect 212 -212 250 -184
rect 278 -212 316 -184
rect 344 -212 382 -184
rect 410 -212 448 -184
rect 476 -212 514 -184
rect 542 -212 580 -184
rect 608 -212 646 -184
rect 674 -212 712 -184
rect 740 -212 778 -184
rect 806 -212 844 -184
rect 872 -212 877 -184
rect -877 -250 877 -212
rect -877 -278 -872 -250
rect -844 -278 -806 -250
rect -778 -278 -740 -250
rect -712 -278 -674 -250
rect -646 -278 -608 -250
rect -580 -278 -542 -250
rect -514 -278 -476 -250
rect -448 -278 -410 -250
rect -382 -278 -344 -250
rect -316 -278 -278 -250
rect -250 -278 -212 -250
rect -184 -278 -146 -250
rect -118 -278 -80 -250
rect -52 -278 -14 -250
rect 14 -278 52 -250
rect 80 -278 118 -250
rect 146 -278 184 -250
rect 212 -278 250 -250
rect 278 -278 316 -250
rect 344 -278 382 -250
rect 410 -278 448 -250
rect 476 -278 514 -250
rect 542 -278 580 -250
rect 608 -278 646 -250
rect 674 -278 712 -250
rect 740 -278 778 -250
rect 806 -278 844 -250
rect 872 -278 877 -250
rect -877 -316 877 -278
rect -877 -344 -872 -316
rect -844 -344 -806 -316
rect -778 -344 -740 -316
rect -712 -344 -674 -316
rect -646 -344 -608 -316
rect -580 -344 -542 -316
rect -514 -344 -476 -316
rect -448 -344 -410 -316
rect -382 -344 -344 -316
rect -316 -344 -278 -316
rect -250 -344 -212 -316
rect -184 -344 -146 -316
rect -118 -344 -80 -316
rect -52 -344 -14 -316
rect 14 -344 52 -316
rect 80 -344 118 -316
rect 146 -344 184 -316
rect 212 -344 250 -316
rect 278 -344 316 -316
rect 344 -344 382 -316
rect 410 -344 448 -316
rect 476 -344 514 -316
rect 542 -344 580 -316
rect 608 -344 646 -316
rect 674 -344 712 -316
rect 740 -344 778 -316
rect 806 -344 844 -316
rect 872 -344 877 -316
rect -877 -349 877 -344
<< via3 >>
rect -872 316 -844 344
rect -806 316 -778 344
rect -740 316 -712 344
rect -674 316 -646 344
rect -608 316 -580 344
rect -542 316 -514 344
rect -476 316 -448 344
rect -410 316 -382 344
rect -344 316 -316 344
rect -278 316 -250 344
rect -212 316 -184 344
rect -146 316 -118 344
rect -80 316 -52 344
rect -14 316 14 344
rect 52 316 80 344
rect 118 316 146 344
rect 184 316 212 344
rect 250 316 278 344
rect 316 316 344 344
rect 382 316 410 344
rect 448 316 476 344
rect 514 316 542 344
rect 580 316 608 344
rect 646 316 674 344
rect 712 316 740 344
rect 778 316 806 344
rect 844 316 872 344
rect -872 250 -844 278
rect -806 250 -778 278
rect -740 250 -712 278
rect -674 250 -646 278
rect -608 250 -580 278
rect -542 250 -514 278
rect -476 250 -448 278
rect -410 250 -382 278
rect -344 250 -316 278
rect -278 250 -250 278
rect -212 250 -184 278
rect -146 250 -118 278
rect -80 250 -52 278
rect -14 250 14 278
rect 52 250 80 278
rect 118 250 146 278
rect 184 250 212 278
rect 250 250 278 278
rect 316 250 344 278
rect 382 250 410 278
rect 448 250 476 278
rect 514 250 542 278
rect 580 250 608 278
rect 646 250 674 278
rect 712 250 740 278
rect 778 250 806 278
rect 844 250 872 278
rect -872 184 -844 212
rect -806 184 -778 212
rect -740 184 -712 212
rect -674 184 -646 212
rect -608 184 -580 212
rect -542 184 -514 212
rect -476 184 -448 212
rect -410 184 -382 212
rect -344 184 -316 212
rect -278 184 -250 212
rect -212 184 -184 212
rect -146 184 -118 212
rect -80 184 -52 212
rect -14 184 14 212
rect 52 184 80 212
rect 118 184 146 212
rect 184 184 212 212
rect 250 184 278 212
rect 316 184 344 212
rect 382 184 410 212
rect 448 184 476 212
rect 514 184 542 212
rect 580 184 608 212
rect 646 184 674 212
rect 712 184 740 212
rect 778 184 806 212
rect 844 184 872 212
rect -872 118 -844 146
rect -806 118 -778 146
rect -740 118 -712 146
rect -674 118 -646 146
rect -608 118 -580 146
rect -542 118 -514 146
rect -476 118 -448 146
rect -410 118 -382 146
rect -344 118 -316 146
rect -278 118 -250 146
rect -212 118 -184 146
rect -146 118 -118 146
rect -80 118 -52 146
rect -14 118 14 146
rect 52 118 80 146
rect 118 118 146 146
rect 184 118 212 146
rect 250 118 278 146
rect 316 118 344 146
rect 382 118 410 146
rect 448 118 476 146
rect 514 118 542 146
rect 580 118 608 146
rect 646 118 674 146
rect 712 118 740 146
rect 778 118 806 146
rect 844 118 872 146
rect -872 52 -844 80
rect -806 52 -778 80
rect -740 52 -712 80
rect -674 52 -646 80
rect -608 52 -580 80
rect -542 52 -514 80
rect -476 52 -448 80
rect -410 52 -382 80
rect -344 52 -316 80
rect -278 52 -250 80
rect -212 52 -184 80
rect -146 52 -118 80
rect -80 52 -52 80
rect -14 52 14 80
rect 52 52 80 80
rect 118 52 146 80
rect 184 52 212 80
rect 250 52 278 80
rect 316 52 344 80
rect 382 52 410 80
rect 448 52 476 80
rect 514 52 542 80
rect 580 52 608 80
rect 646 52 674 80
rect 712 52 740 80
rect 778 52 806 80
rect 844 52 872 80
rect -872 -14 -844 14
rect -806 -14 -778 14
rect -740 -14 -712 14
rect -674 -14 -646 14
rect -608 -14 -580 14
rect -542 -14 -514 14
rect -476 -14 -448 14
rect -410 -14 -382 14
rect -344 -14 -316 14
rect -278 -14 -250 14
rect -212 -14 -184 14
rect -146 -14 -118 14
rect -80 -14 -52 14
rect -14 -14 14 14
rect 52 -14 80 14
rect 118 -14 146 14
rect 184 -14 212 14
rect 250 -14 278 14
rect 316 -14 344 14
rect 382 -14 410 14
rect 448 -14 476 14
rect 514 -14 542 14
rect 580 -14 608 14
rect 646 -14 674 14
rect 712 -14 740 14
rect 778 -14 806 14
rect 844 -14 872 14
rect -872 -80 -844 -52
rect -806 -80 -778 -52
rect -740 -80 -712 -52
rect -674 -80 -646 -52
rect -608 -80 -580 -52
rect -542 -80 -514 -52
rect -476 -80 -448 -52
rect -410 -80 -382 -52
rect -344 -80 -316 -52
rect -278 -80 -250 -52
rect -212 -80 -184 -52
rect -146 -80 -118 -52
rect -80 -80 -52 -52
rect -14 -80 14 -52
rect 52 -80 80 -52
rect 118 -80 146 -52
rect 184 -80 212 -52
rect 250 -80 278 -52
rect 316 -80 344 -52
rect 382 -80 410 -52
rect 448 -80 476 -52
rect 514 -80 542 -52
rect 580 -80 608 -52
rect 646 -80 674 -52
rect 712 -80 740 -52
rect 778 -80 806 -52
rect 844 -80 872 -52
rect -872 -146 -844 -118
rect -806 -146 -778 -118
rect -740 -146 -712 -118
rect -674 -146 -646 -118
rect -608 -146 -580 -118
rect -542 -146 -514 -118
rect -476 -146 -448 -118
rect -410 -146 -382 -118
rect -344 -146 -316 -118
rect -278 -146 -250 -118
rect -212 -146 -184 -118
rect -146 -146 -118 -118
rect -80 -146 -52 -118
rect -14 -146 14 -118
rect 52 -146 80 -118
rect 118 -146 146 -118
rect 184 -146 212 -118
rect 250 -146 278 -118
rect 316 -146 344 -118
rect 382 -146 410 -118
rect 448 -146 476 -118
rect 514 -146 542 -118
rect 580 -146 608 -118
rect 646 -146 674 -118
rect 712 -146 740 -118
rect 778 -146 806 -118
rect 844 -146 872 -118
rect -872 -212 -844 -184
rect -806 -212 -778 -184
rect -740 -212 -712 -184
rect -674 -212 -646 -184
rect -608 -212 -580 -184
rect -542 -212 -514 -184
rect -476 -212 -448 -184
rect -410 -212 -382 -184
rect -344 -212 -316 -184
rect -278 -212 -250 -184
rect -212 -212 -184 -184
rect -146 -212 -118 -184
rect -80 -212 -52 -184
rect -14 -212 14 -184
rect 52 -212 80 -184
rect 118 -212 146 -184
rect 184 -212 212 -184
rect 250 -212 278 -184
rect 316 -212 344 -184
rect 382 -212 410 -184
rect 448 -212 476 -184
rect 514 -212 542 -184
rect 580 -212 608 -184
rect 646 -212 674 -184
rect 712 -212 740 -184
rect 778 -212 806 -184
rect 844 -212 872 -184
rect -872 -278 -844 -250
rect -806 -278 -778 -250
rect -740 -278 -712 -250
rect -674 -278 -646 -250
rect -608 -278 -580 -250
rect -542 -278 -514 -250
rect -476 -278 -448 -250
rect -410 -278 -382 -250
rect -344 -278 -316 -250
rect -278 -278 -250 -250
rect -212 -278 -184 -250
rect -146 -278 -118 -250
rect -80 -278 -52 -250
rect -14 -278 14 -250
rect 52 -278 80 -250
rect 118 -278 146 -250
rect 184 -278 212 -250
rect 250 -278 278 -250
rect 316 -278 344 -250
rect 382 -278 410 -250
rect 448 -278 476 -250
rect 514 -278 542 -250
rect 580 -278 608 -250
rect 646 -278 674 -250
rect 712 -278 740 -250
rect 778 -278 806 -250
rect 844 -278 872 -250
rect -872 -344 -844 -316
rect -806 -344 -778 -316
rect -740 -344 -712 -316
rect -674 -344 -646 -316
rect -608 -344 -580 -316
rect -542 -344 -514 -316
rect -476 -344 -448 -316
rect -410 -344 -382 -316
rect -344 -344 -316 -316
rect -278 -344 -250 -316
rect -212 -344 -184 -316
rect -146 -344 -118 -316
rect -80 -344 -52 -316
rect -14 -344 14 -316
rect 52 -344 80 -316
rect 118 -344 146 -316
rect 184 -344 212 -316
rect 250 -344 278 -316
rect 316 -344 344 -316
rect 382 -344 410 -316
rect 448 -344 476 -316
rect 514 -344 542 -316
rect 580 -344 608 -316
rect 646 -344 674 -316
rect 712 -344 740 -316
rect 778 -344 806 -316
rect 844 -344 872 -316
<< metal4 >>
rect -877 344 877 349
rect -877 316 -872 344
rect -844 316 -806 344
rect -778 316 -740 344
rect -712 316 -674 344
rect -646 316 -608 344
rect -580 316 -542 344
rect -514 316 -476 344
rect -448 316 -410 344
rect -382 316 -344 344
rect -316 316 -278 344
rect -250 316 -212 344
rect -184 316 -146 344
rect -118 316 -80 344
rect -52 316 -14 344
rect 14 316 52 344
rect 80 316 118 344
rect 146 316 184 344
rect 212 316 250 344
rect 278 316 316 344
rect 344 316 382 344
rect 410 316 448 344
rect 476 316 514 344
rect 542 316 580 344
rect 608 316 646 344
rect 674 316 712 344
rect 740 316 778 344
rect 806 316 844 344
rect 872 316 877 344
rect -877 278 877 316
rect -877 250 -872 278
rect -844 250 -806 278
rect -778 250 -740 278
rect -712 250 -674 278
rect -646 250 -608 278
rect -580 250 -542 278
rect -514 250 -476 278
rect -448 250 -410 278
rect -382 250 -344 278
rect -316 250 -278 278
rect -250 250 -212 278
rect -184 250 -146 278
rect -118 250 -80 278
rect -52 250 -14 278
rect 14 250 52 278
rect 80 250 118 278
rect 146 250 184 278
rect 212 250 250 278
rect 278 250 316 278
rect 344 250 382 278
rect 410 250 448 278
rect 476 250 514 278
rect 542 250 580 278
rect 608 250 646 278
rect 674 250 712 278
rect 740 250 778 278
rect 806 250 844 278
rect 872 250 877 278
rect -877 212 877 250
rect -877 184 -872 212
rect -844 184 -806 212
rect -778 184 -740 212
rect -712 184 -674 212
rect -646 184 -608 212
rect -580 184 -542 212
rect -514 184 -476 212
rect -448 184 -410 212
rect -382 184 -344 212
rect -316 184 -278 212
rect -250 184 -212 212
rect -184 184 -146 212
rect -118 184 -80 212
rect -52 184 -14 212
rect 14 184 52 212
rect 80 184 118 212
rect 146 184 184 212
rect 212 184 250 212
rect 278 184 316 212
rect 344 184 382 212
rect 410 184 448 212
rect 476 184 514 212
rect 542 184 580 212
rect 608 184 646 212
rect 674 184 712 212
rect 740 184 778 212
rect 806 184 844 212
rect 872 184 877 212
rect -877 146 877 184
rect -877 118 -872 146
rect -844 118 -806 146
rect -778 118 -740 146
rect -712 118 -674 146
rect -646 118 -608 146
rect -580 118 -542 146
rect -514 118 -476 146
rect -448 118 -410 146
rect -382 118 -344 146
rect -316 118 -278 146
rect -250 118 -212 146
rect -184 118 -146 146
rect -118 118 -80 146
rect -52 118 -14 146
rect 14 118 52 146
rect 80 118 118 146
rect 146 118 184 146
rect 212 118 250 146
rect 278 118 316 146
rect 344 118 382 146
rect 410 118 448 146
rect 476 118 514 146
rect 542 118 580 146
rect 608 118 646 146
rect 674 118 712 146
rect 740 118 778 146
rect 806 118 844 146
rect 872 118 877 146
rect -877 80 877 118
rect -877 52 -872 80
rect -844 52 -806 80
rect -778 52 -740 80
rect -712 52 -674 80
rect -646 52 -608 80
rect -580 52 -542 80
rect -514 52 -476 80
rect -448 52 -410 80
rect -382 52 -344 80
rect -316 52 -278 80
rect -250 52 -212 80
rect -184 52 -146 80
rect -118 52 -80 80
rect -52 52 -14 80
rect 14 52 52 80
rect 80 52 118 80
rect 146 52 184 80
rect 212 52 250 80
rect 278 52 316 80
rect 344 52 382 80
rect 410 52 448 80
rect 476 52 514 80
rect 542 52 580 80
rect 608 52 646 80
rect 674 52 712 80
rect 740 52 778 80
rect 806 52 844 80
rect 872 52 877 80
rect -877 14 877 52
rect -877 -14 -872 14
rect -844 -14 -806 14
rect -778 -14 -740 14
rect -712 -14 -674 14
rect -646 -14 -608 14
rect -580 -14 -542 14
rect -514 -14 -476 14
rect -448 -14 -410 14
rect -382 -14 -344 14
rect -316 -14 -278 14
rect -250 -14 -212 14
rect -184 -14 -146 14
rect -118 -14 -80 14
rect -52 -14 -14 14
rect 14 -14 52 14
rect 80 -14 118 14
rect 146 -14 184 14
rect 212 -14 250 14
rect 278 -14 316 14
rect 344 -14 382 14
rect 410 -14 448 14
rect 476 -14 514 14
rect 542 -14 580 14
rect 608 -14 646 14
rect 674 -14 712 14
rect 740 -14 778 14
rect 806 -14 844 14
rect 872 -14 877 14
rect -877 -52 877 -14
rect -877 -80 -872 -52
rect -844 -80 -806 -52
rect -778 -80 -740 -52
rect -712 -80 -674 -52
rect -646 -80 -608 -52
rect -580 -80 -542 -52
rect -514 -80 -476 -52
rect -448 -80 -410 -52
rect -382 -80 -344 -52
rect -316 -80 -278 -52
rect -250 -80 -212 -52
rect -184 -80 -146 -52
rect -118 -80 -80 -52
rect -52 -80 -14 -52
rect 14 -80 52 -52
rect 80 -80 118 -52
rect 146 -80 184 -52
rect 212 -80 250 -52
rect 278 -80 316 -52
rect 344 -80 382 -52
rect 410 -80 448 -52
rect 476 -80 514 -52
rect 542 -80 580 -52
rect 608 -80 646 -52
rect 674 -80 712 -52
rect 740 -80 778 -52
rect 806 -80 844 -52
rect 872 -80 877 -52
rect -877 -118 877 -80
rect -877 -146 -872 -118
rect -844 -146 -806 -118
rect -778 -146 -740 -118
rect -712 -146 -674 -118
rect -646 -146 -608 -118
rect -580 -146 -542 -118
rect -514 -146 -476 -118
rect -448 -146 -410 -118
rect -382 -146 -344 -118
rect -316 -146 -278 -118
rect -250 -146 -212 -118
rect -184 -146 -146 -118
rect -118 -146 -80 -118
rect -52 -146 -14 -118
rect 14 -146 52 -118
rect 80 -146 118 -118
rect 146 -146 184 -118
rect 212 -146 250 -118
rect 278 -146 316 -118
rect 344 -146 382 -118
rect 410 -146 448 -118
rect 476 -146 514 -118
rect 542 -146 580 -118
rect 608 -146 646 -118
rect 674 -146 712 -118
rect 740 -146 778 -118
rect 806 -146 844 -118
rect 872 -146 877 -118
rect -877 -184 877 -146
rect -877 -212 -872 -184
rect -844 -212 -806 -184
rect -778 -212 -740 -184
rect -712 -212 -674 -184
rect -646 -212 -608 -184
rect -580 -212 -542 -184
rect -514 -212 -476 -184
rect -448 -212 -410 -184
rect -382 -212 -344 -184
rect -316 -212 -278 -184
rect -250 -212 -212 -184
rect -184 -212 -146 -184
rect -118 -212 -80 -184
rect -52 -212 -14 -184
rect 14 -212 52 -184
rect 80 -212 118 -184
rect 146 -212 184 -184
rect 212 -212 250 -184
rect 278 -212 316 -184
rect 344 -212 382 -184
rect 410 -212 448 -184
rect 476 -212 514 -184
rect 542 -212 580 -184
rect 608 -212 646 -184
rect 674 -212 712 -184
rect 740 -212 778 -184
rect 806 -212 844 -184
rect 872 -212 877 -184
rect -877 -250 877 -212
rect -877 -278 -872 -250
rect -844 -278 -806 -250
rect -778 -278 -740 -250
rect -712 -278 -674 -250
rect -646 -278 -608 -250
rect -580 -278 -542 -250
rect -514 -278 -476 -250
rect -448 -278 -410 -250
rect -382 -278 -344 -250
rect -316 -278 -278 -250
rect -250 -278 -212 -250
rect -184 -278 -146 -250
rect -118 -278 -80 -250
rect -52 -278 -14 -250
rect 14 -278 52 -250
rect 80 -278 118 -250
rect 146 -278 184 -250
rect 212 -278 250 -250
rect 278 -278 316 -250
rect 344 -278 382 -250
rect 410 -278 448 -250
rect 476 -278 514 -250
rect 542 -278 580 -250
rect 608 -278 646 -250
rect 674 -278 712 -250
rect 740 -278 778 -250
rect 806 -278 844 -250
rect 872 -278 877 -250
rect -877 -316 877 -278
rect -877 -344 -872 -316
rect -844 -344 -806 -316
rect -778 -344 -740 -316
rect -712 -344 -674 -316
rect -646 -344 -608 -316
rect -580 -344 -542 -316
rect -514 -344 -476 -316
rect -448 -344 -410 -316
rect -382 -344 -344 -316
rect -316 -344 -278 -316
rect -250 -344 -212 -316
rect -184 -344 -146 -316
rect -118 -344 -80 -316
rect -52 -344 -14 -316
rect 14 -344 52 -316
rect 80 -344 118 -316
rect 146 -344 184 -316
rect 212 -344 250 -316
rect 278 -344 316 -316
rect 344 -344 382 -316
rect 410 -344 448 -316
rect 476 -344 514 -316
rect 542 -344 580 -316
rect 608 -344 646 -316
rect 674 -344 712 -316
rect 740 -344 778 -316
rect 806 -344 844 -316
rect 872 -344 877 -316
rect -877 -349 877 -344
<< end >>
