magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1775 1019 1775
<< metal1 >>
rect -19 769 19 775
rect -19 743 -13 769
rect 13 743 19 769
rect -19 715 19 743
rect -19 689 -13 715
rect 13 689 19 715
rect -19 661 19 689
rect -19 635 -13 661
rect 13 635 19 661
rect -19 607 19 635
rect -19 581 -13 607
rect 13 581 19 607
rect -19 553 19 581
rect -19 527 -13 553
rect 13 527 19 553
rect -19 499 19 527
rect -19 473 -13 499
rect 13 473 19 499
rect -19 445 19 473
rect -19 419 -13 445
rect 13 419 19 445
rect -19 391 19 419
rect -19 365 -13 391
rect 13 365 19 391
rect -19 337 19 365
rect -19 311 -13 337
rect 13 311 19 337
rect -19 283 19 311
rect -19 257 -13 283
rect 13 257 19 283
rect -19 229 19 257
rect -19 203 -13 229
rect 13 203 19 229
rect -19 175 19 203
rect -19 149 -13 175
rect 13 149 19 175
rect -19 121 19 149
rect -19 95 -13 121
rect 13 95 19 121
rect -19 67 19 95
rect -19 41 -13 67
rect 13 41 19 67
rect -19 13 19 41
rect -19 -13 -13 13
rect 13 -13 19 13
rect -19 -41 19 -13
rect -19 -67 -13 -41
rect 13 -67 19 -41
rect -19 -95 19 -67
rect -19 -121 -13 -95
rect 13 -121 19 -95
rect -19 -149 19 -121
rect -19 -175 -13 -149
rect 13 -175 19 -149
rect -19 -203 19 -175
rect -19 -229 -13 -203
rect 13 -229 19 -203
rect -19 -257 19 -229
rect -19 -283 -13 -257
rect 13 -283 19 -257
rect -19 -311 19 -283
rect -19 -337 -13 -311
rect 13 -337 19 -311
rect -19 -365 19 -337
rect -19 -391 -13 -365
rect 13 -391 19 -365
rect -19 -419 19 -391
rect -19 -445 -13 -419
rect 13 -445 19 -419
rect -19 -473 19 -445
rect -19 -499 -13 -473
rect 13 -499 19 -473
rect -19 -527 19 -499
rect -19 -553 -13 -527
rect 13 -553 19 -527
rect -19 -581 19 -553
rect -19 -607 -13 -581
rect 13 -607 19 -581
rect -19 -635 19 -607
rect -19 -661 -13 -635
rect 13 -661 19 -635
rect -19 -689 19 -661
rect -19 -715 -13 -689
rect 13 -715 19 -689
rect -19 -743 19 -715
rect -19 -769 -13 -743
rect 13 -769 19 -743
rect -19 -775 19 -769
<< via1 >>
rect -13 743 13 769
rect -13 689 13 715
rect -13 635 13 661
rect -13 581 13 607
rect -13 527 13 553
rect -13 473 13 499
rect -13 419 13 445
rect -13 365 13 391
rect -13 311 13 337
rect -13 257 13 283
rect -13 203 13 229
rect -13 149 13 175
rect -13 95 13 121
rect -13 41 13 67
rect -13 -13 13 13
rect -13 -67 13 -41
rect -13 -121 13 -95
rect -13 -175 13 -149
rect -13 -229 13 -203
rect -13 -283 13 -257
rect -13 -337 13 -311
rect -13 -391 13 -365
rect -13 -445 13 -419
rect -13 -499 13 -473
rect -13 -553 13 -527
rect -13 -607 13 -581
rect -13 -661 13 -635
rect -13 -715 13 -689
rect -13 -769 13 -743
<< metal2 >>
rect -19 769 19 775
rect -19 743 -13 769
rect 13 743 19 769
rect -19 715 19 743
rect -19 689 -13 715
rect 13 689 19 715
rect -19 661 19 689
rect -19 635 -13 661
rect 13 635 19 661
rect -19 607 19 635
rect -19 581 -13 607
rect 13 581 19 607
rect -19 553 19 581
rect -19 527 -13 553
rect 13 527 19 553
rect -19 499 19 527
rect -19 473 -13 499
rect 13 473 19 499
rect -19 445 19 473
rect -19 419 -13 445
rect 13 419 19 445
rect -19 391 19 419
rect -19 365 -13 391
rect 13 365 19 391
rect -19 337 19 365
rect -19 311 -13 337
rect 13 311 19 337
rect -19 283 19 311
rect -19 257 -13 283
rect 13 257 19 283
rect -19 229 19 257
rect -19 203 -13 229
rect 13 203 19 229
rect -19 175 19 203
rect -19 149 -13 175
rect 13 149 19 175
rect -19 121 19 149
rect -19 95 -13 121
rect 13 95 19 121
rect -19 67 19 95
rect -19 41 -13 67
rect 13 41 19 67
rect -19 13 19 41
rect -19 -13 -13 13
rect 13 -13 19 13
rect -19 -41 19 -13
rect -19 -67 -13 -41
rect 13 -67 19 -41
rect -19 -95 19 -67
rect -19 -121 -13 -95
rect 13 -121 19 -95
rect -19 -149 19 -121
rect -19 -175 -13 -149
rect 13 -175 19 -149
rect -19 -203 19 -175
rect -19 -229 -13 -203
rect 13 -229 19 -203
rect -19 -257 19 -229
rect -19 -283 -13 -257
rect 13 -283 19 -257
rect -19 -311 19 -283
rect -19 -337 -13 -311
rect 13 -337 19 -311
rect -19 -365 19 -337
rect -19 -391 -13 -365
rect 13 -391 19 -365
rect -19 -419 19 -391
rect -19 -445 -13 -419
rect 13 -445 19 -419
rect -19 -473 19 -445
rect -19 -499 -13 -473
rect 13 -499 19 -473
rect -19 -527 19 -499
rect -19 -553 -13 -527
rect 13 -553 19 -527
rect -19 -581 19 -553
rect -19 -607 -13 -581
rect 13 -607 19 -581
rect -19 -635 19 -607
rect -19 -661 -13 -635
rect 13 -661 19 -635
rect -19 -689 19 -661
rect -19 -715 -13 -689
rect 13 -715 19 -689
rect -19 -743 19 -715
rect -19 -769 -13 -743
rect 13 -769 19 -743
rect -19 -775 19 -769
<< end >>
