magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1127 -1046 1127 1046
<< metal1 >>
rect -127 40 127 46
rect -127 14 -121 40
rect -95 14 -67 40
rect -41 14 -13 40
rect 13 14 41 40
rect 67 14 95 40
rect 121 14 127 40
rect -127 -14 127 14
rect -127 -40 -121 -14
rect -95 -40 -67 -14
rect -41 -40 -13 -14
rect 13 -40 41 -14
rect 67 -40 95 -14
rect 121 -40 127 -14
rect -127 -46 127 -40
<< via1 >>
rect -121 14 -95 40
rect -67 14 -41 40
rect -13 14 13 40
rect 41 14 67 40
rect 95 14 121 40
rect -121 -40 -95 -14
rect -67 -40 -41 -14
rect -13 -40 13 -14
rect 41 -40 67 -14
rect 95 -40 121 -14
<< metal2 >>
rect -127 40 127 46
rect -127 14 -121 40
rect -95 14 -67 40
rect -41 14 -13 40
rect 13 14 41 40
rect 67 14 95 40
rect 121 14 127 40
rect -127 -14 127 14
rect -127 -40 -121 -14
rect -95 -40 -67 -14
rect -41 -40 -13 -14
rect 13 -40 41 -14
rect 67 -40 95 -14
rect 121 -40 127 -14
rect -127 -46 127 -40
<< end >>
