* NGSPICE file created from resis_magic_flat.ext - technology: gf180mcuC

.subckt pex_resis_magic r1 r2 VDD
X0 VDD.t1 VDD.t2 VDD.t0 ppolyf_u r_width=0.8u r_length=6.46u
X1 r1.t3 r2.t3 VDD.t9 ppolyf_u r_width=0.8u r_length=6.46u
X2 r1.t1 r2.t1 VDD.t7 ppolyf_u r_width=0.8u r_length=6.46u
X3 r1.t0 r2.t0 VDD.t3 ppolyf_u r_width=0.8u r_length=6.46u
X4 VDD.t5 VDD.t6 VDD.t4 ppolyf_u r_width=0.8u r_length=6.46u
X5 r1.t2 r2.t2 VDD.t8 ppolyf_u r_width=0.8u r_length=6.46u
R0 VDD.t3 VDD.t7 128.618
R1 VDD.t9 VDD.t8 128.618
R2 VDD.n0 VDD.t4 112.475
R3 VDD.n7 VDD.t0 112.475
R4 VDD.n3 VDD.t3 64.3092
R5 VDD.n3 VDD.t9 64.3092
R6 VDD.n6 VDD.t1 7.05738
R7 VDD.n2 VDD.t5 7.05738
R8 VDD.n8 VDD.t6 7.05738
R9 VDD.n11 VDD.t2 7.05738
R10 VDD.n12 VDD.n7 3.1505
R11 VDD.n10 VDD.n9 3.1505
R12 VDD.n1 VDD.n0 3.1505
R13 VDD.n5 VDD.n4 3.1505
R14 VDD.n4 VDD.n3 3.1505
R15 VDD.n2 VDD.n1 1.93858
R16 VDD.n12 VDD.n11 1.92634
R17 VDD VDD.n12 1.918
R18 VDD.n6 VDD.n5 1.04752
R19 VDD.n11 VDD.n10 1.04582
R20 VDD.n5 VDD.n2 1.0396
R21 VDD.n10 VDD.n8 1.03824
R22 VDD VDD.n6 0.00745455
R23 r1.n0 r1.t1 7.34172
R24 r1.n9 r1.t2 7.33651
R25 r1.n12 r1.n11 4.5005
R26 r1.n4 r1.n3 4.5005
R27 r1.n10 r1.n8 3.85802
R28 r1.n2 r1.n1 3.84744
R29 r1.n8 r1.t3 2.75071
R30 r1.n1 r1.t0 2.72624
R31 r1.n17 r1.n13 2.24952
R32 r1 r1.n18 0.180045
R33 r1.n7 r1.n6 0.0810714
R34 r1.n4 r1.n2 0.0426491
R35 r1.n12 r1.n10 0.0356429
R36 r1.n10 r1.n9 0.0339658
R37 r1.n2 r1.n0 0.0291957
R38 r1.n13 r1.n7 0.0227857
R39 r1.n6 r1.n5 0.0193571
R40 r1.n16 r1.n15 0.00777273
R41 r1.n5 r1.n4 0.00735714
R42 r1.n17 r1.n16 0.00440715
R43 r1.n18 r1.n17 0.00395261
R44 r1.n13 r1.n12 0.00392857
R45 r1.n15 r1.n14 0.000954545
R46 r2.n10 r2.t2 7.34824
R47 r2.n1 r2.t1 7.32998
R48 r2.n13 r2.n12 4.5005
R49 r2.n11 r2.n9 3.8901
R50 r2.n5 r2.n4 2.87542
R51 r2.n9 r2.t3 2.82343
R52 r2.n3 r2.t0 2.82343
R53 r2.n15 r2.n14 2.24986
R54 r2.n7 r2.n6 2.24862
R55 r2.n4 r2.n3 0.815925
R56 r2 r2.n16 0.202318
R57 r2.n13 r2.n11 0.0469348
R58 r2.n2 r2.n1 0.0336304
R59 r2.n6 r2.n2 0.0278913
R60 r2.n11 r2.n10 0.0226739
R61 r2.n14 r2.n8 0.0138043
R62 r2.n14 r2.n13 0.0114565
R63 r2.n6 r2.n5 0.00971699
R64 r2.n15 r2.n7 0.00853925
R65 r2.n7 r2.n0 0.00576767
R66 r2.n16 r2.n15 0.00327158
C0 r2 r1 0.0346f
C1 r1 VDD 1.19f
C2 r2 VDD 1.18f
C3 r2 VSUBS 0.548f
C4 r1 VSUBS 0.527f
C5 VDD VSUBS 11.9f
.ends

