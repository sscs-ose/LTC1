magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1517 -1022 989 1022
<< metal4 >>
rect -514 14 -14 19
rect -514 -14 -509 14
rect -481 -14 -443 14
rect -415 -14 -377 14
rect -349 -14 -311 14
rect -283 -14 -245 14
rect -217 -14 -179 14
rect -151 -14 -113 14
rect -85 -14 -47 14
rect -19 -14 -14 14
rect -514 -19 -14 -14
<< via4 >>
rect -509 -14 -481 14
rect -443 -14 -415 14
rect -377 -14 -349 14
rect -311 -14 -283 14
rect -245 -14 -217 14
rect -179 -14 -151 14
rect -113 -14 -85 14
rect -47 -14 -19 14
<< metal5 >>
rect -517 14 -11 22
rect -517 -14 -509 14
rect -481 -14 -443 14
rect -415 -14 -377 14
rect -349 -14 -311 14
rect -283 -14 -245 14
rect -217 -14 -179 14
rect -151 -14 -113 14
rect -85 -14 -47 14
rect -19 -14 -11 14
rect -517 -22 -11 -14
<< end >>
