magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1712 -1019 986 1019
<< metal3 >>
rect -712 14 -14 19
rect -712 -14 -707 14
rect -679 -14 -641 14
rect -613 -14 -575 14
rect -547 -14 -509 14
rect -481 -14 -443 14
rect -415 -14 -377 14
rect -349 -14 -311 14
rect -283 -14 -245 14
rect -217 -14 -179 14
rect -151 -14 -113 14
rect -85 -14 -47 14
rect -19 -14 -14 14
rect -712 -19 -14 -14
<< via3 >>
rect -707 -14 -679 14
rect -641 -14 -613 14
rect -575 -14 -547 14
rect -509 -14 -481 14
rect -443 -14 -415 14
rect -377 -14 -349 14
rect -311 -14 -283 14
rect -245 -14 -217 14
rect -179 -14 -151 14
rect -113 -14 -85 14
rect -47 -14 -19 14
<< metal4 >>
rect -712 14 -14 19
rect -712 -14 -707 14
rect -679 -14 -641 14
rect -613 -14 -575 14
rect -547 -14 -509 14
rect -481 -14 -443 14
rect -415 -14 -377 14
rect -349 -14 -311 14
rect -283 -14 -245 14
rect -217 -14 -179 14
rect -151 -14 -113 14
rect -85 -14 -47 14
rect -19 -14 -14 14
rect -712 -19 -14 -14
<< end >>
