magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1050 -1143 1050 1143
<< metal1 >>
rect -50 137 50 143
rect -50 111 -44 137
rect -18 111 18 137
rect 44 111 50 137
rect -50 75 50 111
rect -50 49 -44 75
rect -18 49 18 75
rect 44 49 50 75
rect -50 13 50 49
rect -50 -13 -44 13
rect -18 -13 18 13
rect 44 -13 50 13
rect -50 -49 50 -13
rect -50 -75 -44 -49
rect -18 -75 18 -49
rect 44 -75 50 -49
rect -50 -111 50 -75
rect -50 -137 -44 -111
rect -18 -137 18 -111
rect 44 -137 50 -111
rect -50 -143 50 -137
<< via1 >>
rect -44 111 -18 137
rect 18 111 44 137
rect -44 49 -18 75
rect 18 49 44 75
rect -44 -13 -18 13
rect 18 -13 44 13
rect -44 -75 -18 -49
rect 18 -75 44 -49
rect -44 -137 -18 -111
rect 18 -137 44 -111
<< metal2 >>
rect -50 137 50 143
rect -50 111 -44 137
rect -18 111 18 137
rect 44 111 50 137
rect -50 75 50 111
rect -50 49 -44 75
rect -18 49 18 75
rect 44 49 50 75
rect -50 13 50 49
rect -50 -13 -44 13
rect -18 -13 18 13
rect 44 -13 50 13
rect -50 -49 50 -13
rect -50 -75 -44 -49
rect -18 -75 18 -49
rect 44 -75 50 -49
rect -50 -111 50 -75
rect -50 -137 -44 -111
rect -18 -137 18 -111
rect 44 -137 50 -111
rect -50 -143 50 -137
<< end >>
