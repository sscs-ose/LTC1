magic
tech gf180mcuC
magscale 1 10
timestamp 1692335619
<< nwell >>
rect -762 -1016 762 1016
<< pmos >>
rect -588 386 -532 886
rect -428 386 -372 886
rect -268 386 -212 886
rect -108 386 -52 886
rect 52 386 108 886
rect 212 386 268 886
rect 372 386 428 886
rect 532 386 588 886
rect -588 -250 -532 250
rect -428 -250 -372 250
rect -268 -250 -212 250
rect -108 -250 -52 250
rect 52 -250 108 250
rect 212 -250 268 250
rect 372 -250 428 250
rect 532 -250 588 250
rect -588 -886 -532 -386
rect -428 -886 -372 -386
rect -268 -886 -212 -386
rect -108 -886 -52 -386
rect 52 -886 108 -386
rect 212 -886 268 -386
rect 372 -886 428 -386
rect 532 -886 588 -386
<< pdiff >>
rect -676 873 -588 886
rect -676 399 -663 873
rect -617 399 -588 873
rect -676 386 -588 399
rect -532 873 -428 886
rect -532 399 -503 873
rect -457 399 -428 873
rect -532 386 -428 399
rect -372 873 -268 886
rect -372 399 -343 873
rect -297 399 -268 873
rect -372 386 -268 399
rect -212 873 -108 886
rect -212 399 -183 873
rect -137 399 -108 873
rect -212 386 -108 399
rect -52 873 52 886
rect -52 399 -23 873
rect 23 399 52 873
rect -52 386 52 399
rect 108 873 212 886
rect 108 399 137 873
rect 183 399 212 873
rect 108 386 212 399
rect 268 873 372 886
rect 268 399 297 873
rect 343 399 372 873
rect 268 386 372 399
rect 428 873 532 886
rect 428 399 457 873
rect 503 399 532 873
rect 428 386 532 399
rect 588 873 676 886
rect 588 399 617 873
rect 663 399 676 873
rect 588 386 676 399
rect -676 237 -588 250
rect -676 -237 -663 237
rect -617 -237 -588 237
rect -676 -250 -588 -237
rect -532 237 -428 250
rect -532 -237 -503 237
rect -457 -237 -428 237
rect -532 -250 -428 -237
rect -372 237 -268 250
rect -372 -237 -343 237
rect -297 -237 -268 237
rect -372 -250 -268 -237
rect -212 237 -108 250
rect -212 -237 -183 237
rect -137 -237 -108 237
rect -212 -250 -108 -237
rect -52 237 52 250
rect -52 -237 -23 237
rect 23 -237 52 237
rect -52 -250 52 -237
rect 108 237 212 250
rect 108 -237 137 237
rect 183 -237 212 237
rect 108 -250 212 -237
rect 268 237 372 250
rect 268 -237 297 237
rect 343 -237 372 237
rect 268 -250 372 -237
rect 428 237 532 250
rect 428 -237 457 237
rect 503 -237 532 237
rect 428 -250 532 -237
rect 588 237 676 250
rect 588 -237 617 237
rect 663 -237 676 237
rect 588 -250 676 -237
rect -676 -399 -588 -386
rect -676 -873 -663 -399
rect -617 -873 -588 -399
rect -676 -886 -588 -873
rect -532 -399 -428 -386
rect -532 -873 -503 -399
rect -457 -873 -428 -399
rect -532 -886 -428 -873
rect -372 -399 -268 -386
rect -372 -873 -343 -399
rect -297 -873 -268 -399
rect -372 -886 -268 -873
rect -212 -399 -108 -386
rect -212 -873 -183 -399
rect -137 -873 -108 -399
rect -212 -886 -108 -873
rect -52 -399 52 -386
rect -52 -873 -23 -399
rect 23 -873 52 -399
rect -52 -886 52 -873
rect 108 -399 212 -386
rect 108 -873 137 -399
rect 183 -873 212 -399
rect 108 -886 212 -873
rect 268 -399 372 -386
rect 268 -873 297 -399
rect 343 -873 372 -399
rect 268 -886 372 -873
rect 428 -399 532 -386
rect 428 -873 457 -399
rect 503 -873 532 -399
rect 428 -886 532 -873
rect 588 -399 676 -386
rect 588 -873 617 -399
rect 663 -873 676 -399
rect 588 -886 676 -873
<< pdiffc >>
rect -663 399 -617 873
rect -503 399 -457 873
rect -343 399 -297 873
rect -183 399 -137 873
rect -23 399 23 873
rect 137 399 183 873
rect 297 399 343 873
rect 457 399 503 873
rect 617 399 663 873
rect -663 -237 -617 237
rect -503 -237 -457 237
rect -343 -237 -297 237
rect -183 -237 -137 237
rect -23 -237 23 237
rect 137 -237 183 237
rect 297 -237 343 237
rect 457 -237 503 237
rect 617 -237 663 237
rect -663 -873 -617 -399
rect -503 -873 -457 -399
rect -343 -873 -297 -399
rect -183 -873 -137 -399
rect -23 -873 23 -399
rect 137 -873 183 -399
rect 297 -873 343 -399
rect 457 -873 503 -399
rect 617 -873 663 -399
<< polysilicon >>
rect -588 886 -532 930
rect -428 886 -372 930
rect -268 886 -212 930
rect -108 886 -52 930
rect 52 886 108 930
rect 212 886 268 930
rect 372 886 428 930
rect 532 886 588 930
rect -588 342 -532 386
rect -428 342 -372 386
rect -268 342 -212 386
rect -108 342 -52 386
rect 52 342 108 386
rect 212 342 268 386
rect 372 342 428 386
rect 532 342 588 386
rect -588 250 -532 294
rect -428 250 -372 294
rect -268 250 -212 294
rect -108 250 -52 294
rect 52 250 108 294
rect 212 250 268 294
rect 372 250 428 294
rect 532 250 588 294
rect -588 -294 -532 -250
rect -428 -294 -372 -250
rect -268 -294 -212 -250
rect -108 -294 -52 -250
rect 52 -294 108 -250
rect 212 -294 268 -250
rect 372 -294 428 -250
rect 532 -294 588 -250
rect -588 -386 -532 -342
rect -428 -386 -372 -342
rect -268 -386 -212 -342
rect -108 -386 -52 -342
rect 52 -386 108 -342
rect 212 -386 268 -342
rect 372 -386 428 -342
rect 532 -386 588 -342
rect -588 -930 -532 -886
rect -428 -930 -372 -886
rect -268 -930 -212 -886
rect -108 -930 -52 -886
rect 52 -930 108 -886
rect 212 -930 268 -886
rect 372 -930 428 -886
rect 532 -930 588 -886
<< metal1 >>
rect -663 873 -617 884
rect -663 388 -617 399
rect -503 873 -457 884
rect -503 388 -457 399
rect -343 873 -297 884
rect -343 388 -297 399
rect -183 873 -137 884
rect -183 388 -137 399
rect -23 873 23 884
rect -23 388 23 399
rect 137 873 183 884
rect 137 388 183 399
rect 297 873 343 884
rect 297 388 343 399
rect 457 873 503 884
rect 457 388 503 399
rect 617 873 663 884
rect 617 388 663 399
rect -663 237 -617 248
rect -663 -248 -617 -237
rect -503 237 -457 248
rect -503 -248 -457 -237
rect -343 237 -297 248
rect -343 -248 -297 -237
rect -183 237 -137 248
rect -183 -248 -137 -237
rect -23 237 23 248
rect -23 -248 23 -237
rect 137 237 183 248
rect 137 -248 183 -237
rect 297 237 343 248
rect 297 -248 343 -237
rect 457 237 503 248
rect 457 -248 503 -237
rect 617 237 663 248
rect 617 -248 663 -237
rect -663 -399 -617 -388
rect -663 -884 -617 -873
rect -503 -399 -457 -388
rect -503 -884 -457 -873
rect -343 -399 -297 -388
rect -343 -884 -297 -873
rect -183 -399 -137 -388
rect -183 -884 -137 -873
rect -23 -399 23 -388
rect -23 -884 23 -873
rect 137 -399 183 -388
rect 137 -884 183 -873
rect 297 -399 343 -388
rect 297 -884 343 -873
rect 457 -399 503 -388
rect 457 -884 503 -873
rect 617 -399 663 -388
rect 617 -884 663 -873
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 2.5 l 0.280 m 3 nf 8 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
