magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -5194 -2045 5194 2045
<< psubdiff >>
rect -3194 23 3194 45
rect -3194 -23 -3172 23
rect 3172 -23 3194 23
rect -3194 -45 3194 -23
<< psubdiffcont >>
rect -3172 -23 3172 23
<< metal1 >>
rect -3183 23 3183 34
rect -3183 -23 -3172 23
rect 3172 -23 3183 23
rect -3183 -34 3183 -23
<< end >>
