magic
tech gf180mcuC
magscale 1 10
timestamp 1692798605
<< metal1 >>
rect 2590 6714 2668 6726
rect 2590 6706 2602 6714
rect 2101 6660 2602 6706
rect 2656 6660 2668 6714
rect 2101 6652 2668 6660
rect 2590 6648 2668 6652
rect -393 6560 -315 6572
rect -393 6506 -381 6560
rect -327 6556 -315 6560
rect -327 6510 295 6556
rect -327 6506 -315 6510
rect -393 6494 -315 6506
rect -129 6292 -51 6304
rect -129 6238 -117 6292
rect -63 6288 -51 6292
rect -63 6242 324 6288
rect -63 6238 -51 6242
rect -129 6226 -51 6238
rect 2223 6134 2713 6180
rect -647 5893 -569 5905
rect -647 5839 -635 5893
rect -581 5891 -569 5893
rect -581 5845 292 5891
rect -581 5839 -569 5845
rect -647 5827 -569 5839
rect 2450 5750 2528 5762
rect 2450 5748 2462 5750
rect 2041 5697 2462 5748
rect 2450 5696 2462 5697
rect 2516 5696 2528 5750
rect 2450 5684 2528 5696
rect -520 5602 -442 5614
rect -520 5548 -508 5602
rect -454 5598 -442 5602
rect -454 5552 333 5598
rect -454 5548 -442 5552
rect -520 5536 -442 5548
rect 2231 5263 2713 5309
rect -129 5205 -51 5217
rect -129 5151 -117 5205
rect -63 5201 -51 5205
rect -63 5155 291 5201
rect -63 5151 -51 5155
rect -129 5139 -51 5151
rect -393 4937 -315 4949
rect -393 4883 -381 4937
rect -327 4933 -315 4937
rect -327 4887 294 4933
rect -327 4883 -315 4887
rect -393 4871 -315 4883
rect 2590 4792 2668 4804
rect 2590 4791 2602 4792
rect 2153 4738 2602 4791
rect 2656 4738 2668 4792
rect 2590 4726 2668 4738
rect -266 4646 -188 4658
rect -266 4592 -254 4646
rect -200 4642 -188 4646
rect -200 4596 309 4642
rect -200 4592 -188 4596
rect -266 4580 -188 4592
rect -129 4378 -51 4390
rect -129 4324 -117 4378
rect -63 4374 -51 4378
rect -63 4328 290 4374
rect -63 4324 -51 4328
rect -129 4312 -51 4324
rect 2220 4220 2713 4266
rect -647 3981 -569 3993
rect -647 3927 -635 3981
rect -581 3977 -569 3981
rect -581 3931 301 3977
rect -581 3927 -569 3931
rect -647 3915 -569 3927
rect 2450 3834 2528 3846
rect 2450 3832 2462 3834
rect 2016 3782 2462 3832
rect 2450 3780 2462 3782
rect 2516 3780 2528 3834
rect 2450 3768 2528 3780
rect -520 3688 -442 3700
rect -520 3634 -508 3688
rect -454 3684 -442 3688
rect -454 3638 303 3684
rect -454 3634 -442 3638
rect -520 3622 -442 3634
rect 2224 3349 2713 3395
rect -129 3291 -51 3303
rect -129 3237 -117 3291
rect -63 3287 -51 3291
rect -63 3241 322 3287
rect -63 3237 -51 3241
rect -129 3225 -51 3237
rect -266 3023 -188 3035
rect -266 2969 -254 3023
rect -200 3019 -188 3023
rect -200 2973 288 3019
rect -200 2969 -188 2973
rect -266 2957 -188 2969
rect 2590 2878 2668 2890
rect 2590 2876 2602 2878
rect 2156 2826 2602 2876
rect 2590 2824 2602 2826
rect 2656 2824 2668 2878
rect 2590 2812 2668 2824
rect -393 2732 -315 2744
rect -393 2678 -381 2732
rect -327 2728 -315 2732
rect -327 2682 288 2728
rect -327 2678 -315 2682
rect -393 2666 -315 2678
rect -4 2464 74 2476
rect -4 2410 8 2464
rect 62 2460 74 2464
rect 62 2414 288 2460
rect 62 2410 74 2414
rect -4 2398 74 2410
rect 2231 2306 2713 2352
rect -647 2067 -569 2079
rect -647 2013 -635 2067
rect -581 2063 -569 2067
rect -581 2017 305 2063
rect -581 2013 -569 2017
rect -647 2001 -569 2013
rect 2450 1921 2528 1933
rect 2450 1918 2462 1921
rect 1225 1759 1273 1876
rect 2055 1869 2462 1918
rect 2450 1867 2462 1869
rect 2516 1867 2528 1921
rect 2450 1855 2528 1867
rect 974 1711 1273 1759
rect 1225 1569 1273 1711
rect -520 1391 -442 1403
rect -520 1337 -508 1391
rect -454 1387 -442 1391
rect -454 1341 157 1387
rect -454 1337 -442 1341
rect -520 1325 -442 1337
rect 1111 1174 1190 1220
rect 1111 1041 1157 1174
rect 1032 995 1157 1041
rect 2272 969 2713 1016
rect -266 808 -188 820
rect -266 754 -254 808
rect -200 804 -188 808
rect -200 758 146 804
rect 1120 780 1198 792
rect -200 754 -188 758
rect -266 742 -188 754
rect 1120 726 1132 780
rect 1186 726 1198 780
rect 1205 730 1229 776
rect 1120 714 1198 726
rect 947 588 1351 636
rect -4 525 74 537
rect -4 471 8 525
rect 62 506 74 525
rect 1120 525 1198 537
rect 1120 506 1132 525
rect 62 471 1132 506
rect 1186 471 1198 525
rect -4 459 1198 471
rect -520 432 -442 444
rect -520 378 -508 432
rect -454 413 -442 432
rect -454 378 1675 413
rect -520 373 1675 378
rect -520 366 1609 373
rect -255 307 -177 319
rect -255 253 -243 307
rect -189 303 -177 307
rect 822 308 900 320
rect 822 303 834 308
rect -189 256 834 303
rect -189 253 -177 256
rect -255 241 -177 253
rect 822 254 834 256
rect 888 254 900 308
rect 1597 319 1609 366
rect 1663 319 1675 373
rect 1597 307 1675 319
rect 822 242 900 254
rect 648 138 1119 186
rect 1374 143 1845 191
rect 1870 156 1941 623
rect 2590 198 2668 210
rect 2590 194 2602 198
rect 2200 148 2602 194
rect 2590 144 2602 148
rect 2656 144 2668 198
rect 2590 132 2668 144
rect -4 75 74 87
rect -4 21 8 75
rect 62 70 74 75
rect 62 24 181 70
rect 866 66 944 78
rect 62 21 74 24
rect -4 9 74 21
rect 866 12 878 66
rect 932 12 944 66
rect 866 0 944 12
rect 1596 70 1674 72
rect 1596 16 1608 70
rect 1662 66 1674 70
rect 1662 20 1683 66
rect 1662 16 1674 20
rect 1596 7 1674 16
rect 790 -195 868 -183
rect 790 -199 802 -195
rect 731 -245 802 -199
rect 790 -249 802 -245
rect 856 -249 868 -195
rect 1547 -199 1625 -187
rect 1547 -203 1559 -199
rect 1528 -249 1559 -203
rect 790 -261 868 -249
rect 1547 -253 1559 -249
rect 1613 -253 1625 -199
rect 2297 -199 2375 -187
rect 2297 -203 2309 -199
rect 2285 -249 2309 -203
rect 1547 -265 1625 -253
rect 2297 -253 2309 -249
rect 2363 -253 2375 -199
rect 2297 -265 2375 -253
rect 686 -557 942 -549
rect 685 -589 942 -557
rect 685 -596 941 -589
rect 685 -597 724 -596
rect 932 -597 941 -596
rect 1443 -598 1713 -550
rect 2450 -562 2528 -550
rect 2450 -566 2462 -562
rect 2150 -612 2462 -566
rect 2450 -616 2462 -612
rect 2516 -616 2528 -562
rect 2450 -628 2528 -616
rect -129 -654 -51 -642
rect -129 -708 -117 -654
rect -63 -673 -51 -654
rect 790 -654 868 -642
rect 790 -673 802 -654
rect -63 -708 802 -673
rect 856 -708 868 -654
rect -129 -720 868 -708
rect -392 -748 -314 -736
rect -392 -802 -380 -748
rect -326 -767 -314 -748
rect 1547 -748 1625 -736
rect 1547 -767 1559 -748
rect -326 -802 1559 -767
rect 1613 -802 1625 -748
rect -392 -814 1625 -802
rect -647 -844 -569 -832
rect -647 -898 -635 -844
rect -581 -863 -569 -844
rect 2296 -844 2374 -832
rect 2296 -863 2308 -844
rect -581 -898 2308 -863
rect 2362 -898 2374 -844
rect -647 -910 2374 -898
<< via1 >>
rect 2602 6660 2656 6714
rect -381 6506 -327 6560
rect -117 6238 -63 6292
rect -635 5839 -581 5893
rect 2462 5696 2516 5750
rect -508 5548 -454 5602
rect -117 5151 -63 5205
rect -381 4883 -327 4937
rect 2602 4738 2656 4792
rect -254 4592 -200 4646
rect -117 4324 -63 4378
rect -635 3927 -581 3981
rect 2462 3780 2516 3834
rect -508 3634 -454 3688
rect -117 3237 -63 3291
rect -254 2969 -200 3023
rect 2602 2824 2656 2878
rect -381 2678 -327 2732
rect 8 2410 62 2464
rect -635 2013 -581 2067
rect 2462 1867 2516 1921
rect -508 1337 -454 1391
rect -254 754 -200 808
rect 1132 726 1186 780
rect 8 471 62 525
rect 1132 471 1186 525
rect -508 378 -454 432
rect -243 253 -189 307
rect 834 254 888 308
rect 1609 319 1663 373
rect 2602 144 2656 198
rect 8 21 62 75
rect 878 12 932 66
rect 1608 16 1662 70
rect 802 -249 856 -195
rect 1559 -253 1613 -199
rect 2309 -253 2363 -199
rect 2462 -616 2516 -562
rect -117 -708 -63 -654
rect 802 -708 856 -654
rect -380 -802 -326 -748
rect 1559 -802 1613 -748
rect -635 -898 -581 -844
rect 2308 -898 2362 -844
<< metal2 >>
rect -636 5905 -580 6754
rect -647 5893 -569 5905
rect -647 5839 -635 5893
rect -581 5839 -569 5893
rect -647 5827 -569 5839
rect -636 3993 -580 5827
rect -509 5614 -453 6754
rect -382 6572 -326 6754
rect -393 6560 -315 6572
rect -393 6506 -381 6560
rect -327 6506 -315 6560
rect -393 6494 -315 6506
rect -520 5602 -442 5614
rect -520 5548 -508 5602
rect -454 5548 -442 5602
rect -520 5536 -442 5548
rect -647 3981 -569 3993
rect -647 3927 -635 3981
rect -581 3927 -569 3981
rect -647 3915 -569 3927
rect -636 2079 -580 3915
rect -509 3700 -453 5536
rect -382 4949 -326 6494
rect -393 4937 -315 4949
rect -393 4883 -381 4937
rect -327 4883 -315 4937
rect -393 4871 -315 4883
rect -520 3688 -442 3700
rect -520 3634 -508 3688
rect -454 3634 -442 3688
rect -520 3622 -442 3634
rect -647 2067 -569 2079
rect -647 2013 -635 2067
rect -581 2013 -569 2067
rect -647 2001 -569 2013
rect -636 -832 -580 2001
rect -509 1403 -453 3622
rect -382 2744 -326 4871
rect -255 4658 -199 6754
rect -118 6304 -62 6754
rect -129 6292 -51 6304
rect -129 6238 -117 6292
rect -63 6238 -51 6292
rect -129 6226 -51 6238
rect -118 5217 -62 6226
rect -129 5205 -51 5217
rect -129 5151 -117 5205
rect -63 5151 -51 5205
rect -129 5139 -51 5151
rect -266 4646 -188 4658
rect -266 4592 -254 4646
rect -200 4592 -188 4646
rect -266 4580 -188 4592
rect -255 3035 -199 4580
rect -118 4390 -62 5139
rect -129 4378 -51 4390
rect -129 4324 -117 4378
rect -63 4324 -51 4378
rect -129 4312 -51 4324
rect -118 3303 -62 4312
rect -129 3291 -51 3303
rect -129 3237 -117 3291
rect -63 3237 -51 3291
rect -129 3225 -51 3237
rect -266 3023 -188 3035
rect -266 2969 -254 3023
rect -200 2969 -188 3023
rect -266 2957 -188 2969
rect -393 2732 -315 2744
rect -393 2678 -381 2732
rect -327 2678 -315 2732
rect -393 2666 -315 2678
rect -520 1391 -442 1403
rect -520 1337 -508 1391
rect -454 1337 -442 1391
rect -520 1325 -442 1337
rect -509 444 -453 1325
rect -520 432 -442 444
rect -520 378 -508 432
rect -454 378 -442 432
rect -520 366 -442 378
rect -647 -844 -569 -832
rect -647 -898 -635 -844
rect -581 -898 -569 -844
rect -647 -910 -569 -898
rect -636 -950 -580 -910
rect -509 -950 -453 366
rect -382 -736 -326 2666
rect -255 820 -199 2957
rect -266 808 -188 820
rect -266 754 -254 808
rect -200 754 -188 808
rect -266 742 -188 754
rect -255 319 -199 742
rect -255 307 -177 319
rect -255 253 -243 307
rect -189 253 -177 307
rect -255 241 -177 253
rect -392 -748 -314 -736
rect -392 -802 -380 -748
rect -326 -802 -314 -748
rect -392 -814 -314 -802
rect -382 -950 -326 -814
rect -255 -950 -199 241
rect -118 -642 -62 3225
rect 7 2476 63 6754
rect 2454 5762 2524 6752
rect 2594 6726 2664 6752
rect 2590 6714 2668 6726
rect 2590 6660 2602 6714
rect 2656 6660 2668 6714
rect 2590 6648 2668 6660
rect 2450 5750 2528 5762
rect 2450 5696 2462 5750
rect 2516 5696 2528 5750
rect 2450 5684 2528 5696
rect 2454 3846 2524 5684
rect 2594 4804 2664 6648
rect 2590 4792 2668 4804
rect 2590 4738 2602 4792
rect 2656 4738 2668 4792
rect 2590 4726 2668 4738
rect 2450 3834 2528 3846
rect 2450 3780 2462 3834
rect 2516 3780 2528 3834
rect 2450 3768 2528 3780
rect -4 2464 74 2476
rect -4 2410 8 2464
rect 62 2410 74 2464
rect -4 2398 74 2410
rect 7 537 63 2398
rect 2454 1933 2524 3768
rect 2594 2890 2664 4726
rect 2590 2878 2668 2890
rect 2590 2824 2602 2878
rect 2656 2824 2668 2878
rect 2590 2812 2668 2824
rect 2450 1921 2528 1933
rect 2450 1867 2462 1921
rect 2516 1867 2528 1921
rect 2450 1855 2528 1867
rect 1120 780 1198 792
rect 1120 726 1132 780
rect 1186 726 1198 780
rect 1120 714 1198 726
rect 1131 537 1187 714
rect -4 525 74 537
rect -4 471 8 525
rect 62 471 74 525
rect -4 459 74 471
rect 1120 525 1198 537
rect 1120 471 1132 525
rect 1186 471 1198 525
rect 1120 459 1198 471
rect 7 87 63 459
rect 1597 373 1675 385
rect 822 308 934 320
rect 822 254 834 308
rect 888 254 934 308
rect 1597 319 1609 373
rect 1663 319 1675 373
rect 1597 307 1675 319
rect 822 242 934 254
rect -4 75 74 87
rect 878 78 934 242
rect -4 21 8 75
rect 62 21 74 75
rect -4 9 74 21
rect 866 66 944 78
rect 1608 72 1664 307
rect 866 12 878 66
rect 932 12 944 66
rect -129 -654 -51 -642
rect -129 -708 -117 -654
rect -63 -708 -51 -654
rect -129 -720 -51 -708
rect -118 -950 -62 -720
rect 7 -950 63 9
rect 866 0 944 12
rect 1596 70 1674 72
rect 1596 16 1608 70
rect 1662 16 1674 70
rect 1596 7 1674 16
rect 790 -195 868 -183
rect 790 -249 802 -195
rect 856 -249 868 -195
rect 790 -261 868 -249
rect 1547 -199 1625 -187
rect 1547 -253 1559 -199
rect 1613 -253 1625 -199
rect 801 -642 857 -261
rect 1547 -265 1625 -253
rect 2297 -199 2375 -187
rect 2297 -253 2309 -199
rect 2363 -253 2375 -199
rect 2297 -265 2375 -253
rect 790 -654 868 -642
rect 790 -708 802 -654
rect 856 -708 868 -654
rect 790 -720 868 -708
rect 1558 -736 1614 -265
rect 1547 -748 1625 -736
rect 1547 -802 1559 -748
rect 1613 -802 1625 -748
rect 1547 -814 1625 -802
rect 2308 -832 2364 -265
rect 2454 -550 2524 1855
rect 2594 210 2664 2812
rect 2590 198 2668 210
rect 2590 144 2602 198
rect 2656 144 2668 198
rect 2590 132 2668 144
rect 2450 -562 2528 -550
rect 2450 -616 2462 -562
rect 2516 -616 2528 -562
rect 2450 -628 2528 -616
rect 2296 -844 2374 -832
rect 2296 -898 2308 -844
rect 2362 -898 2374 -844
rect 2296 -910 2374 -898
rect 2454 -950 2524 -628
rect 2594 -950 2664 132
use AND  AND_1
timestamp 1692688043
transform 1 0 1157 0 -1 1488
box -4 -102 1174 945
use AND_3_magic  AND_3_magic_0
timestamp 1692688043
transform 1 0 353 0 -1 5220
box -111 -552 1925 531
use AND_3_magic  AND_3_magic_1
timestamp 1692688043
transform 1 0 353 0 1 6223
box -111 -552 1925 531
use AND_3_magic  AND_3_magic_2
timestamp 1692688043
transform 1 0 353 0 -1 3306
box -111 -552 1925 531
use AND_3_magic  AND_3_magic_3
timestamp 1692688043
transform 1 0 353 0 1 4309
box -111 -552 1925 531
use AND_3_magic  AND_3_magic_5
timestamp 1692688043
transform 1 0 353 0 1 2395
box -111 -552 1925 531
use INVERTER_magic  INVERTER_magic_0
timestamp 1692688043
transform 1 0 160 0 1 -238
box -34 -387 617 468
use INVERTER_magic  INVERTER_magic_1
timestamp 1692688043
transform 1 0 1671 0 1 -242
box -34 -387 617 468
use INVERTER_magic  INVERTER_magic_2
timestamp 1692688043
transform 1 0 916 0 1 -242
box -34 -387 617 468
use OR_magic  OR_magic_1
timestamp 1692688043
transform 1 0 166 0 -1 1027
box -66 -768 912 484
<< labels >>
flabel metal2 33 6712 33 6712 0 FreeSans 480 0 0 0 A
port 1 nsew
flabel metal2 -229 6711 -229 6711 0 FreeSans 480 0 0 0 B
port 3 nsew
flabel metal2 -486 6714 -486 6714 0 FreeSans 480 0 0 0 C
port 5 nsew
flabel metal2 2634 6737 2634 6737 0 FreeSans 480 0 0 0 VDD
port 7 nsew
flabel metal2 2491 6582 2491 6582 0 FreeSans 480 0 0 0 VSS
port 11 nsew
flabel metal1 2689 6159 2689 6159 0 FreeSans 400 0 0 0 S1
port 13 nsew
flabel metal1 2689 5287 2689 5287 0 FreeSans 400 0 0 0 S2
port 15 nsew
flabel metal1 2690 4244 2690 4244 0 FreeSans 400 0 0 0 S3
port 17 nsew
flabel metal1 2690 3374 2690 3374 0 FreeSans 400 0 0 0 S4
port 19 nsew
flabel metal1 2689 2330 2689 2330 0 FreeSans 400 0 0 0 S5
port 21 nsew
flabel metal1 2688 993 2688 993 0 FreeSans 400 0 0 0 S6
port 23 nsew
<< end >>
