magic
tech gf180mcuC
magscale 1 10
timestamp 1691396512
<< pwell >>
rect -540 -840 540 840
<< nmos >>
rect -428 572 -372 772
rect -268 572 -212 772
rect -108 572 -52 772
rect 52 572 108 772
rect 212 572 268 772
rect 372 572 428 772
rect -428 236 -372 436
rect -268 236 -212 436
rect -108 236 -52 436
rect 52 236 108 436
rect 212 236 268 436
rect 372 236 428 436
rect -428 -100 -372 100
rect -268 -100 -212 100
rect -108 -100 -52 100
rect 52 -100 108 100
rect 212 -100 268 100
rect 372 -100 428 100
rect -428 -436 -372 -236
rect -268 -436 -212 -236
rect -108 -436 -52 -236
rect 52 -436 108 -236
rect 212 -436 268 -236
rect 372 -436 428 -236
rect -428 -772 -372 -572
rect -268 -772 -212 -572
rect -108 -772 -52 -572
rect 52 -772 108 -572
rect 212 -772 268 -572
rect 372 -772 428 -572
<< ndiff >>
rect -516 759 -428 772
rect -516 585 -503 759
rect -457 585 -428 759
rect -516 572 -428 585
rect -372 759 -268 772
rect -372 585 -343 759
rect -297 585 -268 759
rect -372 572 -268 585
rect -212 759 -108 772
rect -212 585 -183 759
rect -137 585 -108 759
rect -212 572 -108 585
rect -52 759 52 772
rect -52 585 -23 759
rect 23 585 52 759
rect -52 572 52 585
rect 108 759 212 772
rect 108 585 137 759
rect 183 585 212 759
rect 108 572 212 585
rect 268 759 372 772
rect 268 585 297 759
rect 343 585 372 759
rect 268 572 372 585
rect 428 759 516 772
rect 428 585 457 759
rect 503 585 516 759
rect 428 572 516 585
rect -516 423 -428 436
rect -516 249 -503 423
rect -457 249 -428 423
rect -516 236 -428 249
rect -372 423 -268 436
rect -372 249 -343 423
rect -297 249 -268 423
rect -372 236 -268 249
rect -212 423 -108 436
rect -212 249 -183 423
rect -137 249 -108 423
rect -212 236 -108 249
rect -52 423 52 436
rect -52 249 -23 423
rect 23 249 52 423
rect -52 236 52 249
rect 108 423 212 436
rect 108 249 137 423
rect 183 249 212 423
rect 108 236 212 249
rect 268 423 372 436
rect 268 249 297 423
rect 343 249 372 423
rect 268 236 372 249
rect 428 423 516 436
rect 428 249 457 423
rect 503 249 516 423
rect 428 236 516 249
rect -516 87 -428 100
rect -516 -87 -503 87
rect -457 -87 -428 87
rect -516 -100 -428 -87
rect -372 87 -268 100
rect -372 -87 -343 87
rect -297 -87 -268 87
rect -372 -100 -268 -87
rect -212 87 -108 100
rect -212 -87 -183 87
rect -137 -87 -108 87
rect -212 -100 -108 -87
rect -52 87 52 100
rect -52 -87 -23 87
rect 23 -87 52 87
rect -52 -100 52 -87
rect 108 87 212 100
rect 108 -87 137 87
rect 183 -87 212 87
rect 108 -100 212 -87
rect 268 87 372 100
rect 268 -87 297 87
rect 343 -87 372 87
rect 268 -100 372 -87
rect 428 87 516 100
rect 428 -87 457 87
rect 503 -87 516 87
rect 428 -100 516 -87
rect -516 -249 -428 -236
rect -516 -423 -503 -249
rect -457 -423 -428 -249
rect -516 -436 -428 -423
rect -372 -249 -268 -236
rect -372 -423 -343 -249
rect -297 -423 -268 -249
rect -372 -436 -268 -423
rect -212 -249 -108 -236
rect -212 -423 -183 -249
rect -137 -423 -108 -249
rect -212 -436 -108 -423
rect -52 -249 52 -236
rect -52 -423 -23 -249
rect 23 -423 52 -249
rect -52 -436 52 -423
rect 108 -249 212 -236
rect 108 -423 137 -249
rect 183 -423 212 -249
rect 108 -436 212 -423
rect 268 -249 372 -236
rect 268 -423 297 -249
rect 343 -423 372 -249
rect 268 -436 372 -423
rect 428 -249 516 -236
rect 428 -423 457 -249
rect 503 -423 516 -249
rect 428 -436 516 -423
rect -516 -585 -428 -572
rect -516 -759 -503 -585
rect -457 -759 -428 -585
rect -516 -772 -428 -759
rect -372 -585 -268 -572
rect -372 -759 -343 -585
rect -297 -759 -268 -585
rect -372 -772 -268 -759
rect -212 -585 -108 -572
rect -212 -759 -183 -585
rect -137 -759 -108 -585
rect -212 -772 -108 -759
rect -52 -585 52 -572
rect -52 -759 -23 -585
rect 23 -759 52 -585
rect -52 -772 52 -759
rect 108 -585 212 -572
rect 108 -759 137 -585
rect 183 -759 212 -585
rect 108 -772 212 -759
rect 268 -585 372 -572
rect 268 -759 297 -585
rect 343 -759 372 -585
rect 268 -772 372 -759
rect 428 -585 516 -572
rect 428 -759 457 -585
rect 503 -759 516 -585
rect 428 -772 516 -759
<< ndiffc >>
rect -503 585 -457 759
rect -343 585 -297 759
rect -183 585 -137 759
rect -23 585 23 759
rect 137 585 183 759
rect 297 585 343 759
rect 457 585 503 759
rect -503 249 -457 423
rect -343 249 -297 423
rect -183 249 -137 423
rect -23 249 23 423
rect 137 249 183 423
rect 297 249 343 423
rect 457 249 503 423
rect -503 -87 -457 87
rect -343 -87 -297 87
rect -183 -87 -137 87
rect -23 -87 23 87
rect 137 -87 183 87
rect 297 -87 343 87
rect 457 -87 503 87
rect -503 -423 -457 -249
rect -343 -423 -297 -249
rect -183 -423 -137 -249
rect -23 -423 23 -249
rect 137 -423 183 -249
rect 297 -423 343 -249
rect 457 -423 503 -249
rect -503 -759 -457 -585
rect -343 -759 -297 -585
rect -183 -759 -137 -585
rect -23 -759 23 -585
rect 137 -759 183 -585
rect 297 -759 343 -585
rect 457 -759 503 -585
<< polysilicon >>
rect -428 772 -372 816
rect -268 772 -212 816
rect -108 772 -52 816
rect 52 772 108 816
rect 212 772 268 816
rect 372 772 428 816
rect -428 528 -372 572
rect -268 528 -212 572
rect -108 528 -52 572
rect 52 528 108 572
rect 212 528 268 572
rect 372 528 428 572
rect -428 436 -372 480
rect -268 436 -212 480
rect -108 436 -52 480
rect 52 436 108 480
rect 212 436 268 480
rect 372 436 428 480
rect -428 192 -372 236
rect -268 192 -212 236
rect -108 192 -52 236
rect 52 192 108 236
rect 212 192 268 236
rect 372 192 428 236
rect -428 100 -372 144
rect -268 100 -212 144
rect -108 100 -52 144
rect 52 100 108 144
rect 212 100 268 144
rect 372 100 428 144
rect -428 -144 -372 -100
rect -268 -144 -212 -100
rect -108 -144 -52 -100
rect 52 -144 108 -100
rect 212 -144 268 -100
rect 372 -144 428 -100
rect -428 -236 -372 -192
rect -268 -236 -212 -192
rect -108 -236 -52 -192
rect 52 -236 108 -192
rect 212 -236 268 -192
rect 372 -236 428 -192
rect -428 -480 -372 -436
rect -268 -480 -212 -436
rect -108 -480 -52 -436
rect 52 -480 108 -436
rect 212 -480 268 -436
rect 372 -480 428 -436
rect -428 -572 -372 -528
rect -268 -572 -212 -528
rect -108 -572 -52 -528
rect 52 -572 108 -528
rect 212 -572 268 -528
rect 372 -572 428 -528
rect -428 -816 -372 -772
rect -268 -816 -212 -772
rect -108 -816 -52 -772
rect 52 -816 108 -772
rect 212 -816 268 -772
rect 372 -816 428 -772
<< metal1 >>
rect -503 759 -457 770
rect -503 574 -457 585
rect -343 759 -297 770
rect -343 574 -297 585
rect -183 759 -137 770
rect -183 574 -137 585
rect -23 759 23 770
rect -23 574 23 585
rect 137 759 183 770
rect 137 574 183 585
rect 297 759 343 770
rect 297 574 343 585
rect 457 759 503 770
rect 457 574 503 585
rect -503 423 -457 434
rect -503 238 -457 249
rect -343 423 -297 434
rect -343 238 -297 249
rect -183 423 -137 434
rect -183 238 -137 249
rect -23 423 23 434
rect -23 238 23 249
rect 137 423 183 434
rect 137 238 183 249
rect 297 423 343 434
rect 297 238 343 249
rect 457 423 503 434
rect 457 238 503 249
rect -503 87 -457 98
rect -503 -98 -457 -87
rect -343 87 -297 98
rect -343 -98 -297 -87
rect -183 87 -137 98
rect -183 -98 -137 -87
rect -23 87 23 98
rect -23 -98 23 -87
rect 137 87 183 98
rect 137 -98 183 -87
rect 297 87 343 98
rect 297 -98 343 -87
rect 457 87 503 98
rect 457 -98 503 -87
rect -503 -249 -457 -238
rect -503 -434 -457 -423
rect -343 -249 -297 -238
rect -343 -434 -297 -423
rect -183 -249 -137 -238
rect -183 -434 -137 -423
rect -23 -249 23 -238
rect -23 -434 23 -423
rect 137 -249 183 -238
rect 137 -434 183 -423
rect 297 -249 343 -238
rect 297 -434 343 -423
rect 457 -249 503 -238
rect 457 -434 503 -423
rect -503 -585 -457 -574
rect -503 -770 -457 -759
rect -343 -585 -297 -574
rect -343 -770 -297 -759
rect -183 -585 -137 -574
rect -183 -770 -137 -759
rect -23 -585 23 -574
rect -23 -770 23 -759
rect 137 -585 183 -574
rect 137 -770 183 -759
rect 297 -585 343 -574
rect 297 -770 343 -759
rect 457 -585 503 -574
rect 457 -770 503 -759
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 1 l 0.280 m 5 nf 6 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
