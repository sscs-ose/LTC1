magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1424 -1019 1424 1019
<< metal1 >>
rect -424 13 424 19
rect -424 -13 -418 13
rect -392 -13 -364 13
rect -338 -13 -310 13
rect -284 -13 -256 13
rect -230 -13 -202 13
rect -176 -13 -148 13
rect -122 -13 -94 13
rect -68 -13 -40 13
rect -14 -13 14 13
rect 40 -13 68 13
rect 94 -13 122 13
rect 148 -13 176 13
rect 202 -13 230 13
rect 256 -13 284 13
rect 310 -13 338 13
rect 364 -13 392 13
rect 418 -13 424 13
rect -424 -19 424 -13
<< via1 >>
rect -418 -13 -392 13
rect -364 -13 -338 13
rect -310 -13 -284 13
rect -256 -13 -230 13
rect -202 -13 -176 13
rect -148 -13 -122 13
rect -94 -13 -68 13
rect -40 -13 -14 13
rect 14 -13 40 13
rect 68 -13 94 13
rect 122 -13 148 13
rect 176 -13 202 13
rect 230 -13 256 13
rect 284 -13 310 13
rect 338 -13 364 13
rect 392 -13 418 13
<< metal2 >>
rect -424 13 424 19
rect -424 -13 -418 13
rect -392 -13 -364 13
rect -338 -13 -310 13
rect -284 -13 -256 13
rect -230 -13 -202 13
rect -176 -13 -148 13
rect -122 -13 -94 13
rect -68 -13 -40 13
rect -14 -13 14 13
rect 40 -13 68 13
rect 94 -13 122 13
rect 148 -13 176 13
rect 202 -13 230 13
rect 256 -13 284 13
rect 310 -13 338 13
rect 364 -13 392 13
rect 418 -13 424 13
rect -424 -19 424 -13
<< end >>
