magic
tech gf180mcuC
magscale 1 10
timestamp 1699859038
<< nwell >>
rect -1124 -1136 1124 1136
<< nsubdiff >>
rect -1100 1040 1100 1112
rect -1100 996 -1028 1040
rect -1100 -996 -1087 996
rect -1041 -996 -1028 996
rect 1028 996 1100 1040
rect -1100 -1040 -1028 -996
rect 1028 -996 1041 996
rect 1087 -996 1100 996
rect 1028 -1040 1100 -996
rect -1100 -1112 1100 -1040
<< nsubdiffcont >>
rect -1087 -996 -1041 996
rect 1041 -996 1087 996
<< polysilicon >>
rect -940 939 -740 952
rect -940 893 -927 939
rect -753 893 -740 939
rect -940 850 -740 893
rect -940 -893 -740 -850
rect -940 -939 -927 -893
rect -753 -939 -740 -893
rect -940 -952 -740 -939
rect -660 939 -460 952
rect -660 893 -647 939
rect -473 893 -460 939
rect -660 850 -460 893
rect -660 -893 -460 -850
rect -660 -939 -647 -893
rect -473 -939 -460 -893
rect -660 -952 -460 -939
rect -380 939 -180 952
rect -380 893 -367 939
rect -193 893 -180 939
rect -380 850 -180 893
rect -380 -893 -180 -850
rect -380 -939 -367 -893
rect -193 -939 -180 -893
rect -380 -952 -180 -939
rect -100 939 100 952
rect -100 893 -87 939
rect 87 893 100 939
rect -100 850 100 893
rect -100 -893 100 -850
rect -100 -939 -87 -893
rect 87 -939 100 -893
rect -100 -952 100 -939
rect 180 939 380 952
rect 180 893 193 939
rect 367 893 380 939
rect 180 850 380 893
rect 180 -893 380 -850
rect 180 -939 193 -893
rect 367 -939 380 -893
rect 180 -952 380 -939
rect 460 939 660 952
rect 460 893 473 939
rect 647 893 660 939
rect 460 850 660 893
rect 460 -893 660 -850
rect 460 -939 473 -893
rect 647 -939 660 -893
rect 460 -952 660 -939
rect 740 939 940 952
rect 740 893 753 939
rect 927 893 940 939
rect 740 850 940 893
rect 740 -893 940 -850
rect 740 -939 753 -893
rect 927 -939 940 -893
rect 740 -952 940 -939
<< polycontact >>
rect -927 893 -753 939
rect -927 -939 -753 -893
rect -647 893 -473 939
rect -647 -939 -473 -893
rect -367 893 -193 939
rect -367 -939 -193 -893
rect -87 893 87 939
rect -87 -939 87 -893
rect 193 893 367 939
rect 193 -939 367 -893
rect 473 893 647 939
rect 473 -939 647 -893
rect 753 893 927 939
rect 753 -939 927 -893
<< ppolyres >>
rect -940 -850 -740 850
rect -660 -850 -460 850
rect -380 -850 -180 850
rect -100 -850 100 850
rect 180 -850 380 850
rect 460 -850 660 850
rect 740 -850 940 850
<< metal1 >>
rect -1087 1053 1087 1099
rect -1087 996 -1041 1053
rect 1041 996 1087 1053
rect -938 893 -927 939
rect -753 893 -742 939
rect -658 893 -647 939
rect -473 893 -462 939
rect -378 893 -367 939
rect -193 893 -182 939
rect -98 893 -87 939
rect 87 893 98 939
rect 182 893 193 939
rect 367 893 378 939
rect 462 893 473 939
rect 647 893 658 939
rect 742 893 753 939
rect 927 893 938 939
rect -938 -939 -927 -893
rect -753 -939 -742 -893
rect -658 -939 -647 -893
rect -473 -939 -462 -893
rect -378 -939 -367 -893
rect -193 -939 -182 -893
rect -98 -939 -87 -893
rect 87 -939 98 -893
rect 182 -939 193 -893
rect 367 -939 378 -893
rect 462 -939 473 -893
rect 647 -939 658 -893
rect 742 -939 753 -893
rect 927 -939 938 -893
rect -1087 -1053 -1041 -996
rect 1041 -1053 1087 -996
rect -1087 -1099 1087 -1053
<< properties >>
string FIXED_BBOX -1064 -1076 1064 1076
string gencell ppolyf_u
string library gf180mcu
string parameters w 1.0 l 8.5 m 1 nx 7 wmin 0.80 lmin 1.00 rho 315 val 2.879k dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 1 grc 1 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 1
<< end >>
