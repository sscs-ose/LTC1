magic
tech gf180mcuC
magscale 1 10
timestamp 1691316535
<< error_p >>
rect -538 -23 -527 23
rect 470 -23 481 23
<< pwell >>
rect -564 -97 564 97
<< nmos >>
rect -448 -22 448 22
<< ndiff >>
rect -540 23 -468 36
rect -540 -23 -527 23
rect -481 22 -468 23
rect 468 23 540 36
rect 468 22 481 23
rect -481 -22 -448 22
rect 448 -22 481 22
rect -481 -23 -468 -22
rect -540 -36 -468 -23
rect 468 -23 481 -22
rect 527 -23 540 23
rect 468 -36 540 -23
<< ndiffc >>
rect -527 -23 -481 23
rect 481 -23 527 23
<< polysilicon >>
rect -448 22 448 66
rect -448 -66 448 -22
<< metal1 >>
rect -538 -23 -527 23
rect -481 -23 -470 23
rect 470 -23 481 23
rect 527 -23 538 23
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 0.220 l 4.48 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
