magic
tech gf180mcuC
magscale 1 10
timestamp 1699205295
<< nwell >>
rect -277 1001 3734 1163
rect -277 -1865 -77 1001
rect 3571 -1865 3734 1001
rect -277 -2247 3734 -1865
rect -277 -5113 -77 -2247
rect 3571 -5113 3734 -2247
rect -277 -5275 3734 -5113
<< nsubdiff >>
rect -227 1096 3684 1113
rect -227 1050 -210 1096
rect -164 1050 -112 1096
rect -66 1050 -14 1096
rect 32 1050 84 1096
rect 130 1050 182 1096
rect 228 1050 280 1096
rect 326 1050 378 1096
rect 424 1050 476 1096
rect 522 1050 574 1096
rect 620 1050 672 1096
rect 718 1050 770 1096
rect 816 1050 868 1096
rect 914 1050 966 1096
rect 1012 1050 1064 1096
rect 1110 1050 1162 1096
rect 1208 1050 1260 1096
rect 1306 1050 1358 1096
rect 1404 1050 1456 1096
rect 1502 1050 1554 1096
rect 1600 1050 1652 1096
rect 1698 1050 1750 1096
rect 1796 1050 1848 1096
rect 1894 1050 1946 1096
rect 1992 1050 2044 1096
rect 2090 1050 2142 1096
rect 2188 1050 2240 1096
rect 2286 1050 2338 1096
rect 2384 1050 2436 1096
rect 2482 1050 2534 1096
rect 2580 1050 2632 1096
rect 2678 1050 2730 1096
rect 2776 1050 2828 1096
rect 2874 1050 2926 1096
rect 2972 1050 3024 1096
rect 3070 1050 3122 1096
rect 3168 1050 3220 1096
rect 3266 1050 3318 1096
rect 3364 1050 3416 1096
rect 3462 1050 3514 1096
rect 3560 1050 3621 1096
rect 3667 1050 3684 1096
rect -227 1033 3684 1050
rect -227 988 -147 1033
rect -227 942 -210 988
rect -164 942 -147 988
rect -227 890 -147 942
rect -227 844 -210 890
rect -164 844 -147 890
rect -227 792 -147 844
rect -227 746 -210 792
rect -164 746 -147 792
rect -227 694 -147 746
rect -227 648 -210 694
rect -164 648 -147 694
rect -227 596 -147 648
rect -227 550 -210 596
rect -164 550 -147 596
rect -227 498 -147 550
rect -227 452 -210 498
rect -164 452 -147 498
rect -227 400 -147 452
rect -227 354 -210 400
rect -164 354 -147 400
rect -227 302 -147 354
rect -227 256 -210 302
rect -164 256 -147 302
rect -227 204 -147 256
rect -227 158 -210 204
rect -164 158 -147 204
rect -227 106 -147 158
rect -227 60 -210 106
rect -164 60 -147 106
rect -227 8 -147 60
rect -227 -38 -210 8
rect -164 -38 -147 8
rect -227 -90 -147 -38
rect -227 -136 -210 -90
rect -164 -136 -147 -90
rect -227 -188 -147 -136
rect -227 -234 -210 -188
rect -164 -234 -147 -188
rect -227 -286 -147 -234
rect -227 -332 -210 -286
rect -164 -332 -147 -286
rect -227 -384 -147 -332
rect -227 -430 -210 -384
rect -164 -430 -147 -384
rect -227 -482 -147 -430
rect -227 -528 -210 -482
rect -164 -528 -147 -482
rect -227 -580 -147 -528
rect -227 -626 -210 -580
rect -164 -626 -147 -580
rect -227 -678 -147 -626
rect -227 -724 -210 -678
rect -164 -724 -147 -678
rect -227 -776 -147 -724
rect -227 -822 -210 -776
rect -164 -822 -147 -776
rect -227 -874 -147 -822
rect -227 -920 -210 -874
rect -164 -920 -147 -874
rect -227 -972 -147 -920
rect -227 -1018 -210 -972
rect -164 -1018 -147 -972
rect -227 -1070 -147 -1018
rect -227 -1116 -210 -1070
rect -164 -1116 -147 -1070
rect -227 -1168 -147 -1116
rect -227 -1214 -210 -1168
rect -164 -1214 -147 -1168
rect -227 -1266 -147 -1214
rect -227 -1312 -210 -1266
rect -164 -1312 -147 -1266
rect -227 -1364 -147 -1312
rect -227 -1410 -210 -1364
rect -164 -1410 -147 -1364
rect -227 -1462 -147 -1410
rect -227 -1508 -210 -1462
rect -164 -1508 -147 -1462
rect -227 -1560 -147 -1508
rect -227 -1606 -210 -1560
rect -164 -1606 -147 -1560
rect -227 -1658 -147 -1606
rect -227 -1704 -210 -1658
rect -164 -1704 -147 -1658
rect -227 -1756 -147 -1704
rect -227 -1802 -210 -1756
rect -164 -1802 -147 -1756
rect -227 -1854 -147 -1802
rect -227 -1900 -210 -1854
rect -164 -1900 -147 -1854
rect -227 -1935 -147 -1900
rect 3604 988 3684 1033
rect 3604 942 3621 988
rect 3667 942 3684 988
rect 3604 890 3684 942
rect 3604 844 3621 890
rect 3667 844 3684 890
rect 3604 792 3684 844
rect 3604 746 3621 792
rect 3667 746 3684 792
rect 3604 694 3684 746
rect 3604 648 3621 694
rect 3667 648 3684 694
rect 3604 596 3684 648
rect 3604 550 3621 596
rect 3667 550 3684 596
rect 3604 498 3684 550
rect 3604 452 3621 498
rect 3667 452 3684 498
rect 3604 400 3684 452
rect 3604 354 3621 400
rect 3667 354 3684 400
rect 3604 302 3684 354
rect 3604 256 3621 302
rect 3667 256 3684 302
rect 3604 204 3684 256
rect 3604 158 3621 204
rect 3667 158 3684 204
rect 3604 106 3684 158
rect 3604 60 3621 106
rect 3667 60 3684 106
rect 3604 8 3684 60
rect 3604 -38 3621 8
rect 3667 -38 3684 8
rect 3604 -90 3684 -38
rect 3604 -136 3621 -90
rect 3667 -136 3684 -90
rect 3604 -188 3684 -136
rect 3604 -234 3621 -188
rect 3667 -234 3684 -188
rect 3604 -286 3684 -234
rect 3604 -332 3621 -286
rect 3667 -332 3684 -286
rect 3604 -384 3684 -332
rect 3604 -430 3621 -384
rect 3667 -430 3684 -384
rect 3604 -482 3684 -430
rect 3604 -528 3621 -482
rect 3667 -528 3684 -482
rect 3604 -580 3684 -528
rect 3604 -626 3621 -580
rect 3667 -626 3684 -580
rect 3604 -678 3684 -626
rect 3604 -724 3621 -678
rect 3667 -724 3684 -678
rect 3604 -776 3684 -724
rect 3604 -822 3621 -776
rect 3667 -822 3684 -776
rect 3604 -874 3684 -822
rect 3604 -920 3621 -874
rect 3667 -920 3684 -874
rect 3604 -972 3684 -920
rect 3604 -1018 3621 -972
rect 3667 -1018 3684 -972
rect 3604 -1070 3684 -1018
rect 3604 -1116 3621 -1070
rect 3667 -1116 3684 -1070
rect 3604 -1168 3684 -1116
rect 3604 -1214 3621 -1168
rect 3667 -1214 3684 -1168
rect 3604 -1266 3684 -1214
rect 3604 -1312 3621 -1266
rect 3667 -1312 3684 -1266
rect 3604 -1364 3684 -1312
rect 3604 -1410 3621 -1364
rect 3667 -1410 3684 -1364
rect 3604 -1462 3684 -1410
rect 3604 -1508 3621 -1462
rect 3667 -1508 3684 -1462
rect 3604 -1560 3684 -1508
rect 3604 -1606 3621 -1560
rect 3667 -1606 3684 -1560
rect 3604 -1658 3684 -1606
rect 3604 -1704 3621 -1658
rect 3667 -1704 3684 -1658
rect 3604 -1756 3684 -1704
rect 3604 -1802 3621 -1756
rect 3667 -1802 3684 -1756
rect 3604 -1854 3684 -1802
rect 3604 -1900 3621 -1854
rect 3667 -1900 3684 -1854
rect 3604 -1935 3684 -1900
rect -227 -1952 3684 -1935
rect -227 -1998 -210 -1952
rect -164 -1998 -112 -1952
rect -66 -1998 -14 -1952
rect 32 -1998 84 -1952
rect 130 -1998 182 -1952
rect 228 -1998 280 -1952
rect 326 -1998 378 -1952
rect 424 -1998 476 -1952
rect 522 -1998 574 -1952
rect 620 -1998 672 -1952
rect 718 -1998 770 -1952
rect 816 -1998 868 -1952
rect 914 -1998 966 -1952
rect 1012 -1998 1064 -1952
rect 1110 -1998 1162 -1952
rect 1208 -1998 1260 -1952
rect 1306 -1998 1358 -1952
rect 1404 -1998 1456 -1952
rect 1502 -1998 1554 -1952
rect 1600 -1998 1652 -1952
rect 1698 -1998 1750 -1952
rect 1796 -1998 1848 -1952
rect 1894 -1998 1946 -1952
rect 1992 -1998 2044 -1952
rect 2090 -1998 2142 -1952
rect 2188 -1998 2240 -1952
rect 2286 -1998 2338 -1952
rect 2384 -1998 2436 -1952
rect 2482 -1998 2534 -1952
rect 2580 -1998 2632 -1952
rect 2678 -1998 2730 -1952
rect 2776 -1998 2828 -1952
rect 2874 -1998 2926 -1952
rect 2972 -1998 3024 -1952
rect 3070 -1998 3122 -1952
rect 3168 -1998 3220 -1952
rect 3266 -1998 3318 -1952
rect 3364 -1998 3416 -1952
rect 3462 -1998 3514 -1952
rect 3560 -1998 3621 -1952
rect 3667 -1998 3684 -1952
rect -227 -2015 3684 -1998
rect -227 -2114 3684 -2097
rect -227 -2160 -210 -2114
rect -164 -2160 -112 -2114
rect -66 -2160 -14 -2114
rect 32 -2160 84 -2114
rect 130 -2160 182 -2114
rect 228 -2160 280 -2114
rect 326 -2160 378 -2114
rect 424 -2160 476 -2114
rect 522 -2160 574 -2114
rect 620 -2160 672 -2114
rect 718 -2160 770 -2114
rect 816 -2160 868 -2114
rect 914 -2160 966 -2114
rect 1012 -2160 1064 -2114
rect 1110 -2160 1162 -2114
rect 1208 -2160 1260 -2114
rect 1306 -2160 1358 -2114
rect 1404 -2160 1456 -2114
rect 1502 -2160 1554 -2114
rect 1600 -2160 1652 -2114
rect 1698 -2160 1750 -2114
rect 1796 -2160 1848 -2114
rect 1894 -2160 1946 -2114
rect 1992 -2160 2044 -2114
rect 2090 -2160 2142 -2114
rect 2188 -2160 2240 -2114
rect 2286 -2160 2338 -2114
rect 2384 -2160 2436 -2114
rect 2482 -2160 2534 -2114
rect 2580 -2160 2632 -2114
rect 2678 -2160 2730 -2114
rect 2776 -2160 2828 -2114
rect 2874 -2160 2926 -2114
rect 2972 -2160 3024 -2114
rect 3070 -2160 3122 -2114
rect 3168 -2160 3220 -2114
rect 3266 -2160 3318 -2114
rect 3364 -2160 3416 -2114
rect 3462 -2160 3514 -2114
rect 3560 -2160 3621 -2114
rect 3667 -2160 3684 -2114
rect -227 -2177 3684 -2160
rect -227 -2212 -147 -2177
rect -227 -2258 -210 -2212
rect -164 -2258 -147 -2212
rect -227 -2310 -147 -2258
rect -227 -2356 -210 -2310
rect -164 -2356 -147 -2310
rect -227 -2408 -147 -2356
rect -227 -2454 -210 -2408
rect -164 -2454 -147 -2408
rect -227 -2506 -147 -2454
rect -227 -2552 -210 -2506
rect -164 -2552 -147 -2506
rect -227 -2604 -147 -2552
rect -227 -2650 -210 -2604
rect -164 -2650 -147 -2604
rect -227 -2702 -147 -2650
rect -227 -2748 -210 -2702
rect -164 -2748 -147 -2702
rect -227 -2800 -147 -2748
rect -227 -2846 -210 -2800
rect -164 -2846 -147 -2800
rect -227 -2898 -147 -2846
rect -227 -2944 -210 -2898
rect -164 -2944 -147 -2898
rect -227 -2996 -147 -2944
rect -227 -3042 -210 -2996
rect -164 -3042 -147 -2996
rect -227 -3094 -147 -3042
rect -227 -3140 -210 -3094
rect -164 -3140 -147 -3094
rect -227 -3192 -147 -3140
rect -227 -3238 -210 -3192
rect -164 -3238 -147 -3192
rect -227 -3290 -147 -3238
rect -227 -3336 -210 -3290
rect -164 -3336 -147 -3290
rect -227 -3388 -147 -3336
rect -227 -3434 -210 -3388
rect -164 -3434 -147 -3388
rect -227 -3486 -147 -3434
rect -227 -3532 -210 -3486
rect -164 -3532 -147 -3486
rect -227 -3584 -147 -3532
rect -227 -3630 -210 -3584
rect -164 -3630 -147 -3584
rect -227 -3682 -147 -3630
rect -227 -3728 -210 -3682
rect -164 -3728 -147 -3682
rect -227 -3780 -147 -3728
rect -227 -3826 -210 -3780
rect -164 -3826 -147 -3780
rect -227 -3878 -147 -3826
rect -227 -3924 -210 -3878
rect -164 -3924 -147 -3878
rect -227 -3976 -147 -3924
rect -227 -4022 -210 -3976
rect -164 -4022 -147 -3976
rect -227 -4074 -147 -4022
rect -227 -4120 -210 -4074
rect -164 -4120 -147 -4074
rect -227 -4172 -147 -4120
rect -227 -4218 -210 -4172
rect -164 -4218 -147 -4172
rect -227 -4270 -147 -4218
rect -227 -4316 -210 -4270
rect -164 -4316 -147 -4270
rect -227 -4368 -147 -4316
rect -227 -4414 -210 -4368
rect -164 -4414 -147 -4368
rect -227 -4466 -147 -4414
rect -227 -4512 -210 -4466
rect -164 -4512 -147 -4466
rect -227 -4564 -147 -4512
rect -227 -4610 -210 -4564
rect -164 -4610 -147 -4564
rect -227 -4662 -147 -4610
rect -227 -4708 -210 -4662
rect -164 -4708 -147 -4662
rect -227 -4760 -147 -4708
rect -227 -4806 -210 -4760
rect -164 -4806 -147 -4760
rect -227 -4858 -147 -4806
rect -227 -4904 -210 -4858
rect -164 -4904 -147 -4858
rect -227 -4956 -147 -4904
rect -227 -5002 -210 -4956
rect -164 -5002 -147 -4956
rect -227 -5054 -147 -5002
rect -227 -5100 -210 -5054
rect -164 -5100 -147 -5054
rect -227 -5145 -147 -5100
rect 3604 -2212 3684 -2177
rect 3604 -2258 3621 -2212
rect 3667 -2258 3684 -2212
rect 3604 -2310 3684 -2258
rect 3604 -2356 3621 -2310
rect 3667 -2356 3684 -2310
rect 3604 -2408 3684 -2356
rect 3604 -2454 3621 -2408
rect 3667 -2454 3684 -2408
rect 3604 -2506 3684 -2454
rect 3604 -2552 3621 -2506
rect 3667 -2552 3684 -2506
rect 3604 -2604 3684 -2552
rect 3604 -2650 3621 -2604
rect 3667 -2650 3684 -2604
rect 3604 -2702 3684 -2650
rect 3604 -2748 3621 -2702
rect 3667 -2748 3684 -2702
rect 3604 -2800 3684 -2748
rect 3604 -2846 3621 -2800
rect 3667 -2846 3684 -2800
rect 3604 -2898 3684 -2846
rect 3604 -2944 3621 -2898
rect 3667 -2944 3684 -2898
rect 3604 -2996 3684 -2944
rect 3604 -3042 3621 -2996
rect 3667 -3042 3684 -2996
rect 3604 -3094 3684 -3042
rect 3604 -3140 3621 -3094
rect 3667 -3140 3684 -3094
rect 3604 -3192 3684 -3140
rect 3604 -3238 3621 -3192
rect 3667 -3238 3684 -3192
rect 3604 -3290 3684 -3238
rect 3604 -3336 3621 -3290
rect 3667 -3336 3684 -3290
rect 3604 -3388 3684 -3336
rect 3604 -3434 3621 -3388
rect 3667 -3434 3684 -3388
rect 3604 -3486 3684 -3434
rect 3604 -3532 3621 -3486
rect 3667 -3532 3684 -3486
rect 3604 -3584 3684 -3532
rect 3604 -3630 3621 -3584
rect 3667 -3630 3684 -3584
rect 3604 -3682 3684 -3630
rect 3604 -3728 3621 -3682
rect 3667 -3728 3684 -3682
rect 3604 -3780 3684 -3728
rect 3604 -3826 3621 -3780
rect 3667 -3826 3684 -3780
rect 3604 -3878 3684 -3826
rect 3604 -3924 3621 -3878
rect 3667 -3924 3684 -3878
rect 3604 -3976 3684 -3924
rect 3604 -4022 3621 -3976
rect 3667 -4022 3684 -3976
rect 3604 -4074 3684 -4022
rect 3604 -4120 3621 -4074
rect 3667 -4120 3684 -4074
rect 3604 -4172 3684 -4120
rect 3604 -4218 3621 -4172
rect 3667 -4218 3684 -4172
rect 3604 -4270 3684 -4218
rect 3604 -4316 3621 -4270
rect 3667 -4316 3684 -4270
rect 3604 -4368 3684 -4316
rect 3604 -4414 3621 -4368
rect 3667 -4414 3684 -4368
rect 3604 -4466 3684 -4414
rect 3604 -4512 3621 -4466
rect 3667 -4512 3684 -4466
rect 3604 -4564 3684 -4512
rect 3604 -4610 3621 -4564
rect 3667 -4610 3684 -4564
rect 3604 -4662 3684 -4610
rect 3604 -4708 3621 -4662
rect 3667 -4708 3684 -4662
rect 3604 -4760 3684 -4708
rect 3604 -4806 3621 -4760
rect 3667 -4806 3684 -4760
rect 3604 -4858 3684 -4806
rect 3604 -4904 3621 -4858
rect 3667 -4904 3684 -4858
rect 3604 -4956 3684 -4904
rect 3604 -5002 3621 -4956
rect 3667 -5002 3684 -4956
rect 3604 -5054 3684 -5002
rect 3604 -5100 3621 -5054
rect 3667 -5100 3684 -5054
rect 3604 -5145 3684 -5100
rect -227 -5162 3684 -5145
rect -227 -5208 -210 -5162
rect -164 -5208 -112 -5162
rect -66 -5208 -14 -5162
rect 32 -5208 84 -5162
rect 130 -5208 182 -5162
rect 228 -5208 280 -5162
rect 326 -5208 378 -5162
rect 424 -5208 476 -5162
rect 522 -5208 574 -5162
rect 620 -5208 672 -5162
rect 718 -5208 770 -5162
rect 816 -5208 868 -5162
rect 914 -5208 966 -5162
rect 1012 -5208 1064 -5162
rect 1110 -5208 1162 -5162
rect 1208 -5208 1260 -5162
rect 1306 -5208 1358 -5162
rect 1404 -5208 1456 -5162
rect 1502 -5208 1554 -5162
rect 1600 -5208 1652 -5162
rect 1698 -5208 1750 -5162
rect 1796 -5208 1848 -5162
rect 1894 -5208 1946 -5162
rect 1992 -5208 2044 -5162
rect 2090 -5208 2142 -5162
rect 2188 -5208 2240 -5162
rect 2286 -5208 2338 -5162
rect 2384 -5208 2436 -5162
rect 2482 -5208 2534 -5162
rect 2580 -5208 2632 -5162
rect 2678 -5208 2730 -5162
rect 2776 -5208 2828 -5162
rect 2874 -5208 2926 -5162
rect 2972 -5208 3024 -5162
rect 3070 -5208 3122 -5162
rect 3168 -5208 3220 -5162
rect 3266 -5208 3318 -5162
rect 3364 -5208 3416 -5162
rect 3462 -5208 3514 -5162
rect 3560 -5208 3621 -5162
rect 3667 -5208 3684 -5162
rect -227 -5225 3684 -5208
<< nsubdiffcont >>
rect -210 1050 -164 1096
rect -112 1050 -66 1096
rect -14 1050 32 1096
rect 84 1050 130 1096
rect 182 1050 228 1096
rect 280 1050 326 1096
rect 378 1050 424 1096
rect 476 1050 522 1096
rect 574 1050 620 1096
rect 672 1050 718 1096
rect 770 1050 816 1096
rect 868 1050 914 1096
rect 966 1050 1012 1096
rect 1064 1050 1110 1096
rect 1162 1050 1208 1096
rect 1260 1050 1306 1096
rect 1358 1050 1404 1096
rect 1456 1050 1502 1096
rect 1554 1050 1600 1096
rect 1652 1050 1698 1096
rect 1750 1050 1796 1096
rect 1848 1050 1894 1096
rect 1946 1050 1992 1096
rect 2044 1050 2090 1096
rect 2142 1050 2188 1096
rect 2240 1050 2286 1096
rect 2338 1050 2384 1096
rect 2436 1050 2482 1096
rect 2534 1050 2580 1096
rect 2632 1050 2678 1096
rect 2730 1050 2776 1096
rect 2828 1050 2874 1096
rect 2926 1050 2972 1096
rect 3024 1050 3070 1096
rect 3122 1050 3168 1096
rect 3220 1050 3266 1096
rect 3318 1050 3364 1096
rect 3416 1050 3462 1096
rect 3514 1050 3560 1096
rect 3621 1050 3667 1096
rect -210 942 -164 988
rect -210 844 -164 890
rect -210 746 -164 792
rect -210 648 -164 694
rect -210 550 -164 596
rect -210 452 -164 498
rect -210 354 -164 400
rect -210 256 -164 302
rect -210 158 -164 204
rect -210 60 -164 106
rect -210 -38 -164 8
rect -210 -136 -164 -90
rect -210 -234 -164 -188
rect -210 -332 -164 -286
rect -210 -430 -164 -384
rect -210 -528 -164 -482
rect -210 -626 -164 -580
rect -210 -724 -164 -678
rect -210 -822 -164 -776
rect -210 -920 -164 -874
rect -210 -1018 -164 -972
rect -210 -1116 -164 -1070
rect -210 -1214 -164 -1168
rect -210 -1312 -164 -1266
rect -210 -1410 -164 -1364
rect -210 -1508 -164 -1462
rect -210 -1606 -164 -1560
rect -210 -1704 -164 -1658
rect -210 -1802 -164 -1756
rect -210 -1900 -164 -1854
rect 3621 942 3667 988
rect 3621 844 3667 890
rect 3621 746 3667 792
rect 3621 648 3667 694
rect 3621 550 3667 596
rect 3621 452 3667 498
rect 3621 354 3667 400
rect 3621 256 3667 302
rect 3621 158 3667 204
rect 3621 60 3667 106
rect 3621 -38 3667 8
rect 3621 -136 3667 -90
rect 3621 -234 3667 -188
rect 3621 -332 3667 -286
rect 3621 -430 3667 -384
rect 3621 -528 3667 -482
rect 3621 -626 3667 -580
rect 3621 -724 3667 -678
rect 3621 -822 3667 -776
rect 3621 -920 3667 -874
rect 3621 -1018 3667 -972
rect 3621 -1116 3667 -1070
rect 3621 -1214 3667 -1168
rect 3621 -1312 3667 -1266
rect 3621 -1410 3667 -1364
rect 3621 -1508 3667 -1462
rect 3621 -1606 3667 -1560
rect 3621 -1704 3667 -1658
rect 3621 -1802 3667 -1756
rect 3621 -1900 3667 -1854
rect -210 -1998 -164 -1952
rect -112 -1998 -66 -1952
rect -14 -1998 32 -1952
rect 84 -1998 130 -1952
rect 182 -1998 228 -1952
rect 280 -1998 326 -1952
rect 378 -1998 424 -1952
rect 476 -1998 522 -1952
rect 574 -1998 620 -1952
rect 672 -1998 718 -1952
rect 770 -1998 816 -1952
rect 868 -1998 914 -1952
rect 966 -1998 1012 -1952
rect 1064 -1998 1110 -1952
rect 1162 -1998 1208 -1952
rect 1260 -1998 1306 -1952
rect 1358 -1998 1404 -1952
rect 1456 -1998 1502 -1952
rect 1554 -1998 1600 -1952
rect 1652 -1998 1698 -1952
rect 1750 -1998 1796 -1952
rect 1848 -1998 1894 -1952
rect 1946 -1998 1992 -1952
rect 2044 -1998 2090 -1952
rect 2142 -1998 2188 -1952
rect 2240 -1998 2286 -1952
rect 2338 -1998 2384 -1952
rect 2436 -1998 2482 -1952
rect 2534 -1998 2580 -1952
rect 2632 -1998 2678 -1952
rect 2730 -1998 2776 -1952
rect 2828 -1998 2874 -1952
rect 2926 -1998 2972 -1952
rect 3024 -1998 3070 -1952
rect 3122 -1998 3168 -1952
rect 3220 -1998 3266 -1952
rect 3318 -1998 3364 -1952
rect 3416 -1998 3462 -1952
rect 3514 -1998 3560 -1952
rect 3621 -1998 3667 -1952
rect -210 -2160 -164 -2114
rect -112 -2160 -66 -2114
rect -14 -2160 32 -2114
rect 84 -2160 130 -2114
rect 182 -2160 228 -2114
rect 280 -2160 326 -2114
rect 378 -2160 424 -2114
rect 476 -2160 522 -2114
rect 574 -2160 620 -2114
rect 672 -2160 718 -2114
rect 770 -2160 816 -2114
rect 868 -2160 914 -2114
rect 966 -2160 1012 -2114
rect 1064 -2160 1110 -2114
rect 1162 -2160 1208 -2114
rect 1260 -2160 1306 -2114
rect 1358 -2160 1404 -2114
rect 1456 -2160 1502 -2114
rect 1554 -2160 1600 -2114
rect 1652 -2160 1698 -2114
rect 1750 -2160 1796 -2114
rect 1848 -2160 1894 -2114
rect 1946 -2160 1992 -2114
rect 2044 -2160 2090 -2114
rect 2142 -2160 2188 -2114
rect 2240 -2160 2286 -2114
rect 2338 -2160 2384 -2114
rect 2436 -2160 2482 -2114
rect 2534 -2160 2580 -2114
rect 2632 -2160 2678 -2114
rect 2730 -2160 2776 -2114
rect 2828 -2160 2874 -2114
rect 2926 -2160 2972 -2114
rect 3024 -2160 3070 -2114
rect 3122 -2160 3168 -2114
rect 3220 -2160 3266 -2114
rect 3318 -2160 3364 -2114
rect 3416 -2160 3462 -2114
rect 3514 -2160 3560 -2114
rect 3621 -2160 3667 -2114
rect -210 -2258 -164 -2212
rect -210 -2356 -164 -2310
rect -210 -2454 -164 -2408
rect -210 -2552 -164 -2506
rect -210 -2650 -164 -2604
rect -210 -2748 -164 -2702
rect -210 -2846 -164 -2800
rect -210 -2944 -164 -2898
rect -210 -3042 -164 -2996
rect -210 -3140 -164 -3094
rect -210 -3238 -164 -3192
rect -210 -3336 -164 -3290
rect -210 -3434 -164 -3388
rect -210 -3532 -164 -3486
rect -210 -3630 -164 -3584
rect -210 -3728 -164 -3682
rect -210 -3826 -164 -3780
rect -210 -3924 -164 -3878
rect -210 -4022 -164 -3976
rect -210 -4120 -164 -4074
rect -210 -4218 -164 -4172
rect -210 -4316 -164 -4270
rect -210 -4414 -164 -4368
rect -210 -4512 -164 -4466
rect -210 -4610 -164 -4564
rect -210 -4708 -164 -4662
rect -210 -4806 -164 -4760
rect -210 -4904 -164 -4858
rect -210 -5002 -164 -4956
rect -210 -5100 -164 -5054
rect 3621 -2258 3667 -2212
rect 3621 -2356 3667 -2310
rect 3621 -2454 3667 -2408
rect 3621 -2552 3667 -2506
rect 3621 -2650 3667 -2604
rect 3621 -2748 3667 -2702
rect 3621 -2846 3667 -2800
rect 3621 -2944 3667 -2898
rect 3621 -3042 3667 -2996
rect 3621 -3140 3667 -3094
rect 3621 -3238 3667 -3192
rect 3621 -3336 3667 -3290
rect 3621 -3434 3667 -3388
rect 3621 -3532 3667 -3486
rect 3621 -3630 3667 -3584
rect 3621 -3728 3667 -3682
rect 3621 -3826 3667 -3780
rect 3621 -3924 3667 -3878
rect 3621 -4022 3667 -3976
rect 3621 -4120 3667 -4074
rect 3621 -4218 3667 -4172
rect 3621 -4316 3667 -4270
rect 3621 -4414 3667 -4368
rect 3621 -4512 3667 -4466
rect 3621 -4610 3667 -4564
rect 3621 -4708 3667 -4662
rect 3621 -4806 3667 -4760
rect 3621 -4904 3667 -4858
rect 3621 -5002 3667 -4956
rect 3621 -5100 3667 -5054
rect -210 -5208 -164 -5162
rect -112 -5208 -66 -5162
rect -14 -5208 32 -5162
rect 84 -5208 130 -5162
rect 182 -5208 228 -5162
rect 280 -5208 326 -5162
rect 378 -5208 424 -5162
rect 476 -5208 522 -5162
rect 574 -5208 620 -5162
rect 672 -5208 718 -5162
rect 770 -5208 816 -5162
rect 868 -5208 914 -5162
rect 966 -5208 1012 -5162
rect 1064 -5208 1110 -5162
rect 1162 -5208 1208 -5162
rect 1260 -5208 1306 -5162
rect 1358 -5208 1404 -5162
rect 1456 -5208 1502 -5162
rect 1554 -5208 1600 -5162
rect 1652 -5208 1698 -5162
rect 1750 -5208 1796 -5162
rect 1848 -5208 1894 -5162
rect 1946 -5208 1992 -5162
rect 2044 -5208 2090 -5162
rect 2142 -5208 2188 -5162
rect 2240 -5208 2286 -5162
rect 2338 -5208 2384 -5162
rect 2436 -5208 2482 -5162
rect 2534 -5208 2580 -5162
rect 2632 -5208 2678 -5162
rect 2730 -5208 2776 -5162
rect 2828 -5208 2874 -5162
rect 2926 -5208 2972 -5162
rect 3024 -5208 3070 -5162
rect 3122 -5208 3168 -5162
rect 3220 -5208 3266 -5162
rect 3318 -5208 3364 -5162
rect 3416 -5208 3462 -5162
rect 3514 -5208 3560 -5162
rect 3621 -5208 3667 -5162
<< metal1 >>
rect -227 1096 3684 1113
rect -227 1050 -210 1096
rect -164 1050 -112 1096
rect -66 1050 -14 1096
rect 32 1050 84 1096
rect 130 1050 182 1096
rect 228 1050 280 1096
rect 326 1050 378 1096
rect 424 1050 476 1096
rect 522 1050 574 1096
rect 620 1050 672 1096
rect 718 1050 770 1096
rect 816 1050 868 1096
rect 914 1050 966 1096
rect 1012 1050 1064 1096
rect 1110 1050 1162 1096
rect 1208 1050 1260 1096
rect 1306 1050 1358 1096
rect 1404 1050 1456 1096
rect 1502 1050 1554 1096
rect 1600 1050 1652 1096
rect 1698 1050 1750 1096
rect 1796 1050 1848 1096
rect 1894 1050 1946 1096
rect 1992 1050 2044 1096
rect 2090 1050 2142 1096
rect 2188 1050 2240 1096
rect 2286 1050 2338 1096
rect 2384 1050 2436 1096
rect 2482 1050 2534 1096
rect 2580 1050 2632 1096
rect 2678 1050 2730 1096
rect 2776 1050 2828 1096
rect 2874 1050 2926 1096
rect 2972 1050 3024 1096
rect 3070 1050 3122 1096
rect 3168 1050 3220 1096
rect 3266 1050 3318 1096
rect 3364 1050 3416 1096
rect 3462 1050 3514 1096
rect 3560 1050 3621 1096
rect 3667 1050 3684 1096
rect -227 1033 3684 1050
rect -227 988 -147 1033
rect -227 942 -210 988
rect -164 942 -147 988
rect -227 890 -147 942
rect 3604 988 3684 1033
rect 3604 942 3621 988
rect 3667 942 3684 988
rect -227 844 -210 890
rect -164 844 -147 890
rect -227 811 -147 844
rect 1047 850 1607 918
rect -227 792 305 811
rect -227 746 -210 792
rect -164 746 305 792
rect -227 743 305 746
rect 387 793 587 804
rect -227 694 -147 743
rect 387 737 404 793
rect 460 737 514 793
rect 570 737 587 793
rect 387 731 587 737
rect 667 793 867 804
rect 667 737 684 793
rect 740 737 794 793
rect 850 737 867 793
rect 1047 758 1134 850
rect 667 731 867 737
rect -227 648 -210 694
rect -164 648 -147 694
rect -227 596 -147 648
rect 1326 712 1413 804
rect 1520 758 1607 850
rect 2167 850 2727 918
rect 2167 804 2254 850
rect 2640 804 2727 850
rect 3604 890 3684 942
rect 3604 844 3621 890
rect 3667 844 3684 890
rect 3604 811 3684 844
rect 1789 758 1886 804
rect 2167 758 2265 804
rect 1799 712 1886 758
rect 1326 644 1886 712
rect 2446 712 2533 804
rect 2629 758 2727 804
rect 2909 758 3006 804
rect 2919 712 3006 758
rect 3190 792 3684 811
rect 3190 746 3621 792
rect 3667 746 3684 792
rect 3190 743 3684 746
rect 2446 644 3006 712
rect 3604 694 3684 743
rect 3604 648 3621 694
rect 3667 648 3684 694
rect -227 550 -210 596
rect -164 550 -147 596
rect -227 498 -147 550
rect -227 452 -210 498
rect -164 452 -147 498
rect -227 400 -147 452
rect -227 354 -210 400
rect -164 354 -147 400
rect -227 302 -147 354
rect 3604 596 3684 648
rect 3604 550 3621 596
rect 3667 550 3684 596
rect 3604 498 3684 550
rect 3604 452 3621 498
rect 3667 452 3684 498
rect 3604 400 3684 452
rect 3604 354 3621 400
rect 3667 354 3684 400
rect -227 256 -210 302
rect -164 256 -147 302
rect -227 235 -147 256
rect 767 258 1327 326
rect -227 204 306 235
rect 767 212 854 258
rect 1240 212 1327 258
rect 1887 258 2447 326
rect 1887 212 1974 258
rect 2360 212 2447 258
rect 3604 302 3684 354
rect 3604 256 3621 302
rect 3667 256 3684 302
rect -227 158 -210 204
rect -164 167 306 204
rect -164 158 -147 167
rect -227 106 -147 158
rect -227 60 -210 106
rect -164 60 -147 106
rect -227 8 -147 60
rect 486 120 573 212
rect 767 166 865 212
rect 959 120 1046 212
rect 1229 166 1327 212
rect 486 52 1046 120
rect 1607 120 1694 212
rect 1887 166 1985 212
rect 2080 120 2167 212
rect 2349 166 2447 212
rect 2907 228 3107 239
rect 1607 52 2167 120
rect 2704 119 2791 211
rect 2907 172 2924 228
rect 2980 172 3034 228
rect 3090 172 3107 228
rect 3604 224 3684 256
rect 2907 166 3107 172
rect 3187 204 3684 224
rect 3187 158 3621 204
rect 3667 158 3684 204
rect 3187 156 3684 158
rect 2704 51 2988 119
rect -227 -38 -210 8
rect -164 -38 -147 8
rect -227 -90 -147 -38
rect -227 -136 -210 -90
rect -164 -113 -147 -90
rect 767 -67 1327 1
rect 767 -113 854 -67
rect 1240 -113 1327 -67
rect 1887 -67 2447 1
rect 1887 -113 1974 -67
rect 2360 -113 2447 -67
rect 2920 -113 2988 51
rect 3604 106 3684 156
rect 3604 60 3621 106
rect 3667 60 3684 106
rect 3604 8 3684 60
rect 3604 -38 3621 8
rect 3667 -38 3684 8
rect 3604 -90 3684 -38
rect 3604 -107 3621 -90
rect -164 -136 305 -113
rect -227 -181 305 -136
rect 387 -124 587 -113
rect 387 -180 404 -124
rect 460 -180 514 -124
rect 570 -180 587 -124
rect 767 -159 865 -113
rect -227 -188 -147 -181
rect 387 -186 587 -180
rect -227 -234 -210 -188
rect -164 -234 -147 -188
rect -227 -286 -147 -234
rect 976 -257 1055 -114
rect 1229 -159 1327 -113
rect 1607 -159 1705 -113
rect 1887 -159 1985 -113
rect 2067 -124 2267 -113
rect -227 -332 -210 -286
rect -164 -332 -147 -286
rect -227 -384 -147 -332
rect -227 -430 -210 -384
rect -164 -430 -147 -384
rect -227 -482 -147 -430
rect -227 -528 -210 -482
rect -164 -528 -147 -482
rect -227 -580 -147 -528
rect -227 -626 -210 -580
rect -164 -626 -147 -580
rect -227 -678 -147 -626
rect 707 -336 1055 -257
rect 1607 -232 1694 -159
rect 2067 -180 2084 -124
rect 2140 -180 2194 -124
rect 2250 -180 2267 -124
rect 2349 -159 2447 -113
rect 2067 -186 2267 -180
rect 2685 -232 2753 -117
rect 2907 -124 3107 -113
rect 2907 -180 2924 -124
rect 2980 -180 3034 -124
rect 3090 -180 3107 -124
rect 3188 -136 3621 -107
rect 3667 -136 3684 -90
rect 3188 -175 3684 -136
rect 2907 -186 3107 -180
rect 1607 -300 2753 -232
rect 3604 -188 3684 -175
rect 3604 -234 3621 -188
rect 3667 -234 3684 -188
rect 3604 -286 3684 -234
rect 3604 -332 3621 -286
rect 3667 -332 3684 -286
rect 707 -678 786 -336
rect 3604 -384 3684 -332
rect 3604 -430 3621 -384
rect 3667 -430 3684 -384
rect 1047 -544 2193 -476
rect -227 -724 -210 -678
rect -164 -683 -147 -678
rect -164 -724 305 -683
rect 667 -689 867 -678
rect -227 -751 305 -724
rect -227 -776 -147 -751
rect -227 -822 -210 -776
rect -164 -822 -147 -776
rect -227 -874 -147 -822
rect 488 -797 575 -705
rect 667 -745 684 -689
rect 740 -745 794 -689
rect 850 -745 867 -689
rect 667 -751 867 -745
rect 1047 -705 1134 -544
rect 1327 -659 1887 -591
rect 1327 -705 1414 -659
rect 1800 -705 1887 -659
rect 1047 -751 1145 -705
rect 1327 -751 1425 -705
rect 1547 -797 1634 -705
rect 1789 -751 1887 -705
rect 2125 -747 2193 -544
rect 3604 -482 3684 -430
rect 3604 -528 3621 -482
rect 3667 -528 3684 -482
rect 3604 -580 3684 -528
rect 3604 -626 3621 -580
rect 3667 -626 3684 -580
rect 3604 -678 3684 -626
rect 2627 -689 2827 -678
rect 2447 -751 2545 -705
rect 2627 -745 2644 -689
rect 2700 -745 2754 -689
rect 2810 -745 2827 -689
rect 3604 -692 3621 -678
rect 2627 -751 2827 -745
rect 2909 -751 3007 -705
rect 488 -865 1634 -797
rect 2447 -797 2534 -751
rect 2920 -797 3007 -751
rect 3187 -724 3621 -692
rect 3667 -724 3684 -678
rect 3187 -760 3684 -724
rect 2447 -865 3007 -797
rect 3604 -776 3684 -760
rect 3604 -822 3621 -776
rect 3667 -822 3684 -776
rect -227 -920 -210 -874
rect -164 -920 -147 -874
rect -227 -972 -147 -920
rect -227 -1018 -210 -972
rect -164 -1018 -147 -972
rect 3604 -874 3684 -822
rect 3604 -920 3621 -874
rect 3667 -920 3684 -874
rect 3604 -972 3684 -920
rect -227 -1028 -147 -1018
rect -227 -1070 305 -1028
rect 665 -1029 1148 -1016
rect -227 -1116 -210 -1070
rect -164 -1096 305 -1070
rect 387 -1041 587 -1030
rect -164 -1116 -147 -1096
rect 387 -1097 404 -1041
rect 460 -1097 514 -1041
rect 570 -1097 587 -1041
rect 387 -1103 587 -1097
rect 665 -1087 1149 -1029
rect 1225 -1030 1705 -1028
rect 1783 -1030 2264 -1016
rect 3604 -1018 3621 -972
rect 3667 -1018 3684 -972
rect 2343 -1030 2824 -1020
rect 3604 -1023 3684 -1018
rect -227 -1168 -147 -1116
rect -227 -1214 -210 -1168
rect -164 -1214 -147 -1168
rect 665 -1170 1148 -1087
rect 1225 -1159 1709 -1030
rect 1226 -1184 1709 -1159
rect 1783 -1088 2269 -1030
rect 2343 -1088 2829 -1030
rect 2907 -1041 3107 -1030
rect 2907 -1065 2924 -1041
rect 1783 -1186 2264 -1088
rect 2343 -1190 2824 -1088
rect 2903 -1097 2924 -1065
rect 2980 -1097 3034 -1041
rect 3090 -1097 3107 -1041
rect 3187 -1070 3684 -1023
rect 3187 -1091 3621 -1070
rect 2903 -1103 3107 -1097
rect -227 -1266 -147 -1214
rect -227 -1312 -210 -1266
rect -164 -1312 -147 -1266
rect -227 -1364 -147 -1312
rect -227 -1410 -210 -1364
rect -164 -1410 -147 -1364
rect -227 -1462 -147 -1410
rect -227 -1508 -210 -1462
rect -164 -1508 -147 -1462
rect -227 -1560 -147 -1508
rect -227 -1606 -210 -1560
rect -164 -1606 -147 -1560
rect -227 -1612 -147 -1606
rect -227 -1658 307 -1612
rect -227 -1704 -210 -1658
rect -164 -1680 307 -1658
rect -164 -1704 -147 -1680
rect 387 -1682 870 -1528
rect 945 -1610 1428 -1527
rect 1506 -1610 1986 -1546
rect 2064 -1610 2545 -1509
rect 2674 -1516 2820 -1190
rect 2903 -1516 3092 -1103
rect 3604 -1116 3621 -1091
rect 3667 -1116 3684 -1070
rect 3604 -1168 3684 -1116
rect 3604 -1214 3621 -1168
rect 3667 -1214 3684 -1168
rect 3604 -1266 3684 -1214
rect 3604 -1312 3621 -1266
rect 3667 -1312 3684 -1266
rect 3604 -1364 3684 -1312
rect 3604 -1410 3621 -1364
rect 3667 -1410 3684 -1364
rect 3604 -1462 3684 -1410
rect 3604 -1508 3621 -1462
rect 3667 -1508 3684 -1462
rect 945 -1668 1429 -1610
rect 1506 -1668 1989 -1610
rect 2064 -1668 2549 -1610
rect 945 -1681 1428 -1668
rect 1506 -1677 1986 -1668
rect 2064 -1679 2545 -1668
rect 2628 -1686 3109 -1516
rect 3604 -1560 3684 -1508
rect 3604 -1606 3621 -1560
rect 3667 -1606 3684 -1560
rect 3604 -1612 3684 -1606
rect 3187 -1658 3684 -1612
rect 3187 -1680 3621 -1658
rect -227 -1756 -147 -1704
rect -227 -1802 -210 -1756
rect -164 -1802 -147 -1756
rect -227 -1854 -147 -1802
rect -227 -1900 -210 -1854
rect -164 -1900 -147 -1854
rect -227 -1935 -147 -1900
rect 3604 -1704 3621 -1680
rect 3667 -1704 3684 -1658
rect 3604 -1756 3684 -1704
rect 3604 -1802 3621 -1756
rect 3667 -1802 3684 -1756
rect 3604 -1854 3684 -1802
rect 3604 -1900 3621 -1854
rect 3667 -1900 3684 -1854
rect 3604 -1935 3684 -1900
rect -227 -1952 3684 -1935
rect -227 -1998 -210 -1952
rect -164 -1998 -112 -1952
rect -66 -1998 -14 -1952
rect 32 -1998 84 -1952
rect 130 -1998 182 -1952
rect 228 -1998 280 -1952
rect 326 -1998 378 -1952
rect 424 -1998 476 -1952
rect 522 -1998 574 -1952
rect 620 -1998 672 -1952
rect 718 -1998 770 -1952
rect 816 -1998 868 -1952
rect 914 -1998 966 -1952
rect 1012 -1998 1064 -1952
rect 1110 -1998 1162 -1952
rect 1208 -1998 1260 -1952
rect 1306 -1998 1358 -1952
rect 1404 -1998 1456 -1952
rect 1502 -1998 1554 -1952
rect 1600 -1998 1652 -1952
rect 1698 -1998 1750 -1952
rect 1796 -1998 1848 -1952
rect 1894 -1998 1946 -1952
rect 1992 -1998 2044 -1952
rect 2090 -1998 2142 -1952
rect 2188 -1998 2240 -1952
rect 2286 -1998 2338 -1952
rect 2384 -1998 2436 -1952
rect 2482 -1998 2534 -1952
rect 2580 -1998 2632 -1952
rect 2678 -1998 2730 -1952
rect 2776 -1998 2828 -1952
rect 2874 -1998 2926 -1952
rect 2972 -1998 3024 -1952
rect 3070 -1998 3122 -1952
rect 3168 -1998 3220 -1952
rect 3266 -1998 3318 -1952
rect 3364 -1998 3416 -1952
rect 3462 -1998 3514 -1952
rect 3560 -1998 3621 -1952
rect 3667 -1998 3684 -1952
rect -227 -2015 3684 -1998
rect -119 -2097 3584 -2015
rect -227 -2114 3684 -2097
rect -227 -2160 -210 -2114
rect -164 -2160 -112 -2114
rect -66 -2160 -14 -2114
rect 32 -2160 84 -2114
rect 130 -2160 182 -2114
rect 228 -2160 280 -2114
rect 326 -2160 378 -2114
rect 424 -2160 476 -2114
rect 522 -2160 574 -2114
rect 620 -2160 672 -2114
rect 718 -2160 770 -2114
rect 816 -2160 868 -2114
rect 914 -2160 966 -2114
rect 1012 -2160 1064 -2114
rect 1110 -2160 1162 -2114
rect 1208 -2160 1260 -2114
rect 1306 -2160 1358 -2114
rect 1404 -2160 1456 -2114
rect 1502 -2160 1554 -2114
rect 1600 -2160 1652 -2114
rect 1698 -2160 1750 -2114
rect 1796 -2160 1848 -2114
rect 1894 -2160 1946 -2114
rect 1992 -2160 2044 -2114
rect 2090 -2160 2142 -2114
rect 2188 -2160 2240 -2114
rect 2286 -2160 2338 -2114
rect 2384 -2160 2436 -2114
rect 2482 -2160 2534 -2114
rect 2580 -2160 2632 -2114
rect 2678 -2160 2730 -2114
rect 2776 -2160 2828 -2114
rect 2874 -2160 2926 -2114
rect 2972 -2160 3024 -2114
rect 3070 -2160 3122 -2114
rect 3168 -2160 3220 -2114
rect 3266 -2160 3318 -2114
rect 3364 -2160 3416 -2114
rect 3462 -2160 3514 -2114
rect 3560 -2160 3621 -2114
rect 3667 -2160 3684 -2114
rect -227 -2177 3684 -2160
rect -227 -2212 -147 -2177
rect -227 -2258 -210 -2212
rect -164 -2258 -147 -2212
rect -227 -2310 -147 -2258
rect -227 -2356 -210 -2310
rect -164 -2356 -147 -2310
rect -227 -2408 -147 -2356
rect -227 -2454 -210 -2408
rect -164 -2432 -147 -2408
rect 3604 -2212 3684 -2177
rect 3604 -2258 3621 -2212
rect 3667 -2258 3684 -2212
rect 3604 -2310 3684 -2258
rect 3604 -2356 3621 -2310
rect 3667 -2356 3684 -2310
rect 3604 -2408 3684 -2356
rect -164 -2454 307 -2432
rect -227 -2500 307 -2454
rect -227 -2506 -147 -2500
rect -227 -2552 -210 -2506
rect -164 -2552 -147 -2506
rect -227 -2604 -147 -2552
rect 384 -2588 867 -2434
rect 946 -2582 1429 -2428
rect 1506 -2582 1989 -2428
rect 2066 -2585 2549 -2431
rect 2627 -2583 3110 -2429
rect 3604 -2432 3621 -2408
rect 3187 -2454 3621 -2432
rect 3667 -2454 3684 -2408
rect 3187 -2500 3684 -2454
rect 3604 -2506 3684 -2500
rect 3604 -2552 3621 -2506
rect 3667 -2552 3684 -2506
rect -227 -2650 -210 -2604
rect -164 -2650 -147 -2604
rect -227 -2702 -147 -2650
rect -227 -2748 -210 -2702
rect -164 -2748 -147 -2702
rect -227 -2800 -147 -2748
rect -227 -2846 -210 -2800
rect -164 -2846 -147 -2800
rect -227 -2898 -147 -2846
rect -227 -2944 -210 -2898
rect -164 -2944 -147 -2898
rect -227 -2996 -147 -2944
rect -227 -3042 -210 -2996
rect -164 -3016 -147 -2996
rect 387 -3015 587 -3009
rect -164 -3042 305 -3016
rect -227 -3084 305 -3042
rect 387 -3071 404 -3015
rect 460 -3071 514 -3015
rect 570 -3071 587 -3015
rect 387 -3082 587 -3071
rect -227 -3094 -147 -3084
rect 667 -3094 1150 -2940
rect 1227 -3094 1710 -2940
rect 2647 -2943 2807 -2583
rect -227 -3140 -210 -3094
rect -164 -3140 -147 -3094
rect 1789 -3097 2272 -2943
rect 2346 -3097 2829 -2943
rect 2925 -3009 3085 -2583
rect 3604 -2604 3684 -2552
rect 3604 -2650 3621 -2604
rect 3667 -2650 3684 -2604
rect 3604 -2702 3684 -2650
rect 3604 -2748 3621 -2702
rect 3667 -2748 3684 -2702
rect 3604 -2800 3684 -2748
rect 3604 -2846 3621 -2800
rect 3667 -2846 3684 -2800
rect 3604 -2898 3684 -2846
rect 3604 -2944 3621 -2898
rect 3667 -2944 3684 -2898
rect 3604 -2996 3684 -2944
rect 2907 -3015 3107 -3009
rect 2907 -3071 2924 -3015
rect 2980 -3071 3034 -3015
rect 3090 -3071 3107 -3015
rect 3604 -3021 3621 -2996
rect 2907 -3082 3107 -3071
rect 3187 -3042 3621 -3021
rect 3667 -3042 3684 -2996
rect 3187 -3089 3684 -3042
rect 3604 -3094 3684 -3089
rect -227 -3192 -147 -3140
rect -227 -3238 -210 -3192
rect -164 -3238 -147 -3192
rect -227 -3290 -147 -3238
rect 3604 -3140 3621 -3094
rect 3667 -3140 3684 -3094
rect 3604 -3192 3684 -3140
rect 3604 -3238 3621 -3192
rect 3667 -3238 3684 -3192
rect -227 -3336 -210 -3290
rect -164 -3336 -147 -3290
rect -227 -3361 -147 -3336
rect 488 -3315 1634 -3247
rect -227 -3388 305 -3361
rect -227 -3434 -210 -3388
rect -164 -3429 305 -3388
rect 488 -3407 575 -3315
rect 667 -3367 867 -3361
rect 667 -3423 684 -3367
rect 740 -3423 794 -3367
rect 850 -3423 867 -3367
rect -164 -3434 -147 -3429
rect 667 -3434 867 -3423
rect 1047 -3407 1145 -3361
rect 1327 -3407 1425 -3361
rect 1547 -3407 1634 -3315
rect 2447 -3315 3007 -3247
rect 2447 -3361 2534 -3315
rect 2920 -3361 3007 -3315
rect 3604 -3290 3684 -3238
rect 3604 -3336 3621 -3290
rect 3667 -3336 3684 -3290
rect 3604 -3352 3684 -3336
rect 1789 -3407 1887 -3361
rect -227 -3486 -147 -3434
rect -227 -3532 -210 -3486
rect -164 -3532 -147 -3486
rect -227 -3584 -147 -3532
rect -227 -3630 -210 -3584
rect -164 -3630 -147 -3584
rect -227 -3682 -147 -3630
rect -227 -3728 -210 -3682
rect -164 -3728 -147 -3682
rect -227 -3780 -147 -3728
rect -227 -3826 -210 -3780
rect -164 -3826 -147 -3780
rect -227 -3878 -147 -3826
rect 707 -3776 786 -3434
rect 1047 -3568 1134 -3407
rect 1327 -3453 1414 -3407
rect 1800 -3453 1887 -3407
rect 1327 -3521 1887 -3453
rect 2125 -3568 2193 -3365
rect 2447 -3407 2545 -3361
rect 2627 -3367 2827 -3361
rect 2627 -3423 2644 -3367
rect 2700 -3423 2754 -3367
rect 2810 -3423 2827 -3367
rect 2909 -3407 3007 -3361
rect 3187 -3388 3684 -3352
rect 3187 -3420 3621 -3388
rect 2627 -3434 2827 -3423
rect 3604 -3434 3621 -3420
rect 3667 -3434 3684 -3388
rect 1047 -3636 2193 -3568
rect 3604 -3486 3684 -3434
rect 3604 -3532 3621 -3486
rect 3667 -3532 3684 -3486
rect 3604 -3584 3684 -3532
rect 3604 -3630 3621 -3584
rect 3667 -3630 3684 -3584
rect 3604 -3682 3684 -3630
rect 3604 -3728 3621 -3682
rect 3667 -3728 3684 -3682
rect 707 -3855 1055 -3776
rect 3604 -3780 3684 -3728
rect -227 -3924 -210 -3878
rect -164 -3924 -147 -3878
rect -227 -3931 -147 -3924
rect -227 -3976 305 -3931
rect -227 -4022 -210 -3976
rect -164 -3999 305 -3976
rect 387 -3932 587 -3926
rect 387 -3988 404 -3932
rect 460 -3988 514 -3932
rect 570 -3988 587 -3932
rect 387 -3999 587 -3988
rect 767 -3999 865 -3953
rect 976 -3998 1055 -3855
rect 1607 -3880 2753 -3812
rect 1607 -3953 1694 -3880
rect 2067 -3932 2267 -3926
rect 1229 -3999 1327 -3953
rect 1607 -3999 1705 -3953
rect 1887 -3999 1985 -3953
rect 2067 -3988 2084 -3932
rect 2140 -3988 2194 -3932
rect 2250 -3988 2267 -3932
rect 2067 -3999 2267 -3988
rect 2349 -3999 2447 -3953
rect 2685 -3995 2753 -3880
rect 3604 -3826 3621 -3780
rect 3667 -3826 3684 -3780
rect 3604 -3878 3684 -3826
rect 3604 -3924 3621 -3878
rect 3667 -3924 3684 -3878
rect 2907 -3932 3107 -3926
rect 2907 -3988 2924 -3932
rect 2980 -3988 3034 -3932
rect 3090 -3988 3107 -3932
rect 3604 -3937 3684 -3924
rect 2907 -3999 3107 -3988
rect 3188 -3976 3684 -3937
rect -164 -4022 -147 -3999
rect -227 -4074 -147 -4022
rect -227 -4120 -210 -4074
rect -164 -4120 -147 -4074
rect 767 -4045 854 -3999
rect 1240 -4045 1327 -3999
rect 767 -4113 1327 -4045
rect 1887 -4045 1974 -3999
rect 2360 -4045 2447 -3999
rect 1887 -4113 2447 -4045
rect -227 -4172 -147 -4120
rect 2920 -4163 2988 -3999
rect 3188 -4005 3621 -3976
rect -227 -4218 -210 -4172
rect -164 -4218 -147 -4172
rect -227 -4270 -147 -4218
rect -227 -4316 -210 -4270
rect -164 -4279 -147 -4270
rect 486 -4232 1046 -4164
rect -164 -4316 306 -4279
rect -227 -4347 306 -4316
rect 486 -4324 573 -4232
rect 767 -4324 865 -4278
rect 959 -4324 1046 -4232
rect 1607 -4232 2167 -4164
rect 1229 -4324 1327 -4278
rect 1607 -4324 1694 -4232
rect 1887 -4324 1985 -4278
rect 2080 -4324 2167 -4232
rect 2704 -4231 2988 -4163
rect 3604 -4022 3621 -4005
rect 3667 -4022 3684 -3976
rect 3604 -4074 3684 -4022
rect 3604 -4120 3621 -4074
rect 3667 -4120 3684 -4074
rect 3604 -4172 3684 -4120
rect 3604 -4218 3621 -4172
rect 3667 -4218 3684 -4172
rect 2349 -4324 2447 -4278
rect 2704 -4323 2791 -4231
rect 3604 -4268 3684 -4218
rect 3187 -4270 3684 -4268
rect 2907 -4284 3107 -4278
rect -227 -4368 -147 -4347
rect -227 -4414 -210 -4368
rect -164 -4414 -147 -4368
rect -227 -4466 -147 -4414
rect 767 -4370 854 -4324
rect 1240 -4370 1327 -4324
rect 767 -4438 1327 -4370
rect 1887 -4370 1974 -4324
rect 2360 -4370 2447 -4324
rect 2907 -4340 2924 -4284
rect 2980 -4340 3034 -4284
rect 3090 -4340 3107 -4284
rect 3187 -4316 3621 -4270
rect 3667 -4316 3684 -4270
rect 3187 -4336 3684 -4316
rect 2907 -4351 3107 -4340
rect 1887 -4438 2447 -4370
rect 3604 -4368 3684 -4336
rect 3604 -4414 3621 -4368
rect 3667 -4414 3684 -4368
rect -227 -4512 -210 -4466
rect -164 -4512 -147 -4466
rect -227 -4564 -147 -4512
rect -227 -4610 -210 -4564
rect -164 -4610 -147 -4564
rect -227 -4662 -147 -4610
rect -227 -4708 -210 -4662
rect -164 -4708 -147 -4662
rect -227 -4760 -147 -4708
rect 3604 -4466 3684 -4414
rect 3604 -4512 3621 -4466
rect 3667 -4512 3684 -4466
rect 3604 -4564 3684 -4512
rect 3604 -4610 3621 -4564
rect 3667 -4610 3684 -4564
rect 3604 -4662 3684 -4610
rect 3604 -4708 3621 -4662
rect 3667 -4708 3684 -4662
rect -227 -4806 -210 -4760
rect -164 -4806 -147 -4760
rect -227 -4855 -147 -4806
rect 1326 -4824 1886 -4756
rect 387 -4849 587 -4843
rect -227 -4858 305 -4855
rect -227 -4904 -210 -4858
rect -164 -4904 305 -4858
rect -227 -4923 305 -4904
rect 387 -4905 404 -4849
rect 460 -4905 514 -4849
rect 570 -4905 587 -4849
rect 387 -4916 587 -4905
rect 667 -4849 867 -4843
rect 667 -4905 684 -4849
rect 740 -4905 794 -4849
rect 850 -4905 867 -4849
rect 667 -4916 867 -4905
rect -227 -4956 -147 -4923
rect -227 -5002 -210 -4956
rect -164 -5002 -147 -4956
rect -227 -5054 -147 -5002
rect 1047 -4962 1134 -4870
rect 1326 -4916 1413 -4824
rect 1799 -4870 1886 -4824
rect 2446 -4824 3006 -4756
rect 1520 -4962 1607 -4870
rect 1789 -4916 1886 -4870
rect 2167 -4916 2265 -4870
rect 2446 -4916 2533 -4824
rect 2919 -4870 3006 -4824
rect 3604 -4760 3684 -4708
rect 3604 -4806 3621 -4760
rect 3667 -4806 3684 -4760
rect 3604 -4855 3684 -4806
rect 2629 -4916 2727 -4870
rect 2909 -4916 3006 -4870
rect 3190 -4858 3684 -4855
rect 3190 -4904 3621 -4858
rect 3667 -4904 3684 -4858
rect 1047 -5030 1607 -4962
rect 2167 -4962 2254 -4916
rect 2640 -4962 2727 -4916
rect 3190 -4923 3684 -4904
rect 2167 -5030 2727 -4962
rect 3604 -4956 3684 -4923
rect 3604 -5002 3621 -4956
rect 3667 -5002 3684 -4956
rect -227 -5100 -210 -5054
rect -164 -5100 -147 -5054
rect -227 -5145 -147 -5100
rect 3604 -5054 3684 -5002
rect 3604 -5100 3621 -5054
rect 3667 -5100 3684 -5054
rect 3604 -5145 3684 -5100
rect -227 -5162 3684 -5145
rect -227 -5208 -210 -5162
rect -164 -5208 -112 -5162
rect -66 -5208 -14 -5162
rect 32 -5208 84 -5162
rect 130 -5208 182 -5162
rect 228 -5208 280 -5162
rect 326 -5208 378 -5162
rect 424 -5208 476 -5162
rect 522 -5208 574 -5162
rect 620 -5208 672 -5162
rect 718 -5208 770 -5162
rect 816 -5208 868 -5162
rect 914 -5208 966 -5162
rect 1012 -5208 1064 -5162
rect 1110 -5208 1162 -5162
rect 1208 -5208 1260 -5162
rect 1306 -5208 1358 -5162
rect 1404 -5208 1456 -5162
rect 1502 -5208 1554 -5162
rect 1600 -5208 1652 -5162
rect 1698 -5208 1750 -5162
rect 1796 -5208 1848 -5162
rect 1894 -5208 1946 -5162
rect 1992 -5208 2044 -5162
rect 2090 -5208 2142 -5162
rect 2188 -5208 2240 -5162
rect 2286 -5208 2338 -5162
rect 2384 -5208 2436 -5162
rect 2482 -5208 2534 -5162
rect 2580 -5208 2632 -5162
rect 2678 -5208 2730 -5162
rect 2776 -5208 2828 -5162
rect 2874 -5208 2926 -5162
rect 2972 -5208 3024 -5162
rect 3070 -5208 3122 -5162
rect 3168 -5208 3220 -5162
rect 3266 -5208 3318 -5162
rect 3364 -5208 3416 -5162
rect 3462 -5208 3514 -5162
rect 3560 -5208 3621 -5162
rect 3667 -5208 3684 -5162
rect -227 -5225 3684 -5208
<< via1 >>
rect 404 737 460 793
rect 514 737 570 793
rect 684 737 740 793
rect 794 737 850 793
rect 2924 172 2980 228
rect 3034 172 3090 228
rect 404 -180 460 -124
rect 514 -180 570 -124
rect 2084 -180 2140 -124
rect 2194 -180 2250 -124
rect 2924 -180 2980 -124
rect 3034 -180 3090 -124
rect 684 -745 740 -689
rect 794 -745 850 -689
rect 2644 -745 2700 -689
rect 2754 -745 2810 -689
rect 404 -1097 460 -1041
rect 514 -1097 570 -1041
rect 2924 -1097 2980 -1041
rect 3034 -1097 3090 -1041
rect 404 -3071 460 -3015
rect 514 -3071 570 -3015
rect 2924 -3071 2980 -3015
rect 3034 -3071 3090 -3015
rect 684 -3423 740 -3367
rect 794 -3423 850 -3367
rect 2644 -3423 2700 -3367
rect 2754 -3423 2810 -3367
rect 404 -3988 460 -3932
rect 514 -3988 570 -3932
rect 2084 -3988 2140 -3932
rect 2194 -3988 2250 -3932
rect 2924 -3988 2980 -3932
rect 3034 -3988 3090 -3932
rect 2924 -4340 2980 -4284
rect 3034 -4340 3090 -4284
rect 404 -4905 460 -4849
rect 514 -4905 570 -4849
rect 684 -4905 740 -4849
rect 794 -4905 850 -4849
<< metal2 >>
rect -680 3503 -468 3515
rect -680 3447 -665 3503
rect -609 3447 -555 3503
rect -499 3493 -468 3503
rect -499 3447 562 3493
rect -680 3393 562 3447
rect -680 3337 -665 3393
rect -609 3337 -555 3393
rect -499 3337 562 3393
rect -680 3336 562 3337
rect -680 3303 -468 3336
rect 405 804 562 3336
rect 3867 1127 4079 1150
rect 3867 1071 3889 1127
rect 3945 1071 3999 1127
rect 4055 1071 4079 1127
rect 3867 1017 4079 1071
rect 3867 961 3889 1017
rect 3945 961 3999 1017
rect 4055 961 4079 1017
rect 3867 938 4079 961
rect 387 793 587 804
rect 387 737 404 793
rect 460 737 514 793
rect 570 737 587 793
rect 387 731 587 737
rect 667 793 867 804
rect 667 737 684 793
rect 740 737 794 793
rect 850 737 867 793
rect 667 731 867 737
rect -661 159 -449 169
rect -661 103 -648 159
rect -592 103 -538 159
rect -482 103 -449 159
rect -661 94 -449 103
rect 697 94 808 731
rect 2907 228 3107 239
rect 2907 172 2924 228
rect 2980 172 3034 228
rect 3090 172 3107 228
rect 2907 166 3107 172
rect 2968 106 3068 166
rect -661 54 808 94
rect -661 -2 -648 54
rect -592 -2 -538 54
rect -482 -2 808 54
rect -661 -51 808 -2
rect -661 -107 -648 -51
rect -592 -107 -538 -51
rect -482 -59 808 -51
rect 2145 6 3068 106
rect -482 -107 -449 -59
rect -661 -122 -449 -107
rect 387 -124 587 -59
rect 2145 -113 2245 6
rect 387 -180 404 -124
rect 460 -180 514 -124
rect 570 -180 587 -124
rect 387 -186 587 -180
rect 2067 -124 2267 -113
rect 2067 -180 2084 -124
rect 2140 -180 2194 -124
rect 2250 -180 2267 -124
rect 2067 -186 2267 -180
rect 2907 -124 3107 -113
rect 2907 -180 2924 -124
rect 2980 -180 3034 -124
rect 3090 -180 3107 -124
rect 2907 -186 3107 -180
rect -447 -449 2827 -352
rect -449 -580 2827 -449
rect 667 -689 867 -678
rect 667 -745 684 -689
rect 740 -745 794 -689
rect 850 -745 867 -689
rect -1020 -803 -810 -798
rect 667 -803 867 -745
rect 2625 -689 2827 -580
rect 2625 -745 2644 -689
rect 2700 -745 2754 -689
rect 2810 -745 2827 -689
rect 2625 -749 2827 -745
rect 2627 -751 2827 -749
rect -1020 -810 867 -803
rect -1020 -866 -998 -810
rect -942 -866 -888 -810
rect -832 -866 867 -810
rect -1020 -920 867 -866
rect -1020 -976 -998 -920
rect -942 -976 -888 -920
rect -832 -974 867 -920
rect -832 -975 824 -974
rect -832 -976 -810 -975
rect -1020 -1030 -810 -976
rect -1020 -1086 -998 -1030
rect -942 -1086 -888 -1030
rect -832 -1086 -810 -1030
rect -1020 -1140 -810 -1086
rect 387 -1041 587 -975
rect 387 -1097 404 -1041
rect 460 -1097 514 -1041
rect 570 -1097 587 -1041
rect 387 -1103 587 -1097
rect 2907 -1041 3107 -1030
rect 2907 -1097 2924 -1041
rect 2980 -1097 3034 -1041
rect 3090 -1097 3107 -1041
rect 2907 -1103 3107 -1097
rect -1020 -1196 -998 -1140
rect -942 -1196 -888 -1140
rect -832 -1196 -810 -1140
rect -1020 -1224 -810 -1196
rect 2929 -1263 3086 -1103
rect 3892 -1263 4049 938
rect 2929 -1420 4049 -1263
rect -3329 -1477 -2914 -1456
rect -3329 -1482 -763 -1477
rect -3329 -1538 -3312 -1482
rect -3256 -1538 -3202 -1482
rect -3146 -1538 -3092 -1482
rect -3036 -1538 -2982 -1482
rect -2926 -1538 -763 -1482
rect -3329 -1592 -763 -1538
rect -3329 -1648 -3312 -1592
rect -3256 -1648 -3202 -1592
rect -3146 -1648 -3092 -1592
rect -3036 -1648 -2982 -1592
rect -2926 -1648 -763 -1592
rect -3329 -1649 -763 -1648
rect -3329 -1681 -2914 -1649
rect -935 -3137 -763 -1649
rect 2929 -2849 4049 -2692
rect 2929 -3009 3086 -2849
rect 387 -3015 587 -3009
rect 387 -3071 404 -3015
rect 460 -3071 514 -3015
rect 570 -3071 587 -3015
rect 387 -3078 587 -3071
rect 386 -3137 587 -3078
rect 2907 -3015 3107 -3009
rect 2907 -3071 2924 -3015
rect 2980 -3071 3034 -3015
rect 3090 -3071 3107 -3015
rect 2907 -3082 3107 -3071
rect -935 -3309 867 -3137
rect 667 -3367 867 -3309
rect 667 -3423 684 -3367
rect 740 -3423 794 -3367
rect 850 -3423 867 -3367
rect 667 -3434 867 -3423
rect 2627 -3367 2827 -3361
rect 2627 -3423 2644 -3367
rect 2700 -3423 2754 -3367
rect 2810 -3423 2827 -3367
rect 2627 -3532 2827 -3423
rect -370 -3644 2827 -3532
rect -371 -3774 2827 -3644
rect -371 -3775 2781 -3774
rect 387 -3932 587 -3926
rect 387 -3988 404 -3932
rect 460 -3988 514 -3932
rect 570 -3988 587 -3932
rect 387 -3999 587 -3988
rect 2067 -3932 2267 -3926
rect 2067 -3988 2084 -3932
rect 2140 -3988 2194 -3932
rect 2250 -3988 2267 -3932
rect 2067 -3999 2267 -3988
rect 2907 -3932 3107 -3926
rect 2907 -3988 2924 -3932
rect 2980 -3988 3034 -3932
rect 3090 -3988 3107 -3932
rect 2907 -3999 3107 -3988
rect -666 -4020 -370 -4002
rect 387 -4020 504 -3999
rect -722 -4076 -653 -4020
rect -597 -4076 -548 -4020
rect -492 -4076 -443 -4020
rect -387 -4076 504 -4020
rect -722 -4077 504 -4076
rect -722 -4130 808 -4077
rect -722 -4186 -653 -4130
rect -597 -4186 -548 -4130
rect -492 -4186 -443 -4130
rect -387 -4186 808 -4130
rect -722 -4188 808 -4186
rect -722 -4190 385 -4188
rect -666 -4214 -370 -4190
rect 697 -4843 808 -4188
rect 2145 -4118 2245 -3999
rect 2145 -4218 3068 -4118
rect 2968 -4278 3068 -4218
rect 2907 -4284 3107 -4278
rect 2907 -4340 2924 -4284
rect 2980 -4340 3034 -4284
rect 3090 -4340 3107 -4284
rect 2907 -4351 3107 -4340
rect 387 -4849 587 -4843
rect 387 -4905 404 -4849
rect 460 -4905 514 -4849
rect 570 -4905 587 -4849
rect 387 -4916 587 -4905
rect 667 -4849 867 -4843
rect 667 -4905 684 -4849
rect 740 -4905 794 -4849
rect 850 -4905 867 -4849
rect 667 -4916 867 -4905
rect -680 -7448 -468 -7415
rect 405 -7448 562 -4916
rect 3892 -5100 4049 -2849
rect 3867 -5123 4079 -5100
rect 3867 -5179 3889 -5123
rect 3945 -5179 3999 -5123
rect 4055 -5179 4079 -5123
rect 3867 -5233 4079 -5179
rect 3867 -5289 3889 -5233
rect 3945 -5289 3999 -5233
rect 4055 -5289 4079 -5233
rect 3867 -5312 4079 -5289
rect -680 -7449 562 -7448
rect -680 -7505 -665 -7449
rect -609 -7505 -555 -7449
rect -499 -7505 562 -7449
rect -680 -7559 562 -7505
rect -680 -7615 -665 -7559
rect -609 -7615 -555 -7559
rect -499 -7605 562 -7559
rect -499 -7615 -468 -7605
rect -680 -7627 -468 -7615
<< via2 >>
rect -665 3447 -609 3503
rect -555 3447 -499 3503
rect -665 3337 -609 3393
rect -555 3337 -499 3393
rect 3889 1071 3945 1127
rect 3999 1071 4055 1127
rect 3889 961 3945 1017
rect 3999 961 4055 1017
rect -648 103 -592 159
rect -538 103 -482 159
rect -648 -2 -592 54
rect -538 -2 -482 54
rect -648 -107 -592 -51
rect -538 -107 -482 -51
rect -998 -866 -942 -810
rect -888 -866 -832 -810
rect -998 -976 -942 -920
rect -888 -976 -832 -920
rect -998 -1086 -942 -1030
rect -888 -1086 -832 -1030
rect -998 -1196 -942 -1140
rect -888 -1196 -832 -1140
rect -3312 -1538 -3256 -1482
rect -3202 -1538 -3146 -1482
rect -3092 -1538 -3036 -1482
rect -2982 -1538 -2926 -1482
rect -3312 -1648 -3256 -1592
rect -3202 -1648 -3146 -1592
rect -3092 -1648 -3036 -1592
rect -2982 -1648 -2926 -1592
rect -653 -4076 -597 -4020
rect -548 -4076 -492 -4020
rect -443 -4076 -387 -4020
rect -653 -4186 -597 -4130
rect -548 -4186 -492 -4130
rect -443 -4186 -387 -4130
rect 3889 -5179 3945 -5123
rect 3999 -5179 4055 -5123
rect 3889 -5289 3945 -5233
rect 3999 -5289 4055 -5233
rect -665 -7505 -609 -7449
rect -555 -7505 -499 -7449
rect -665 -7615 -609 -7559
rect -555 -7615 -499 -7559
<< metal3 >>
rect -680 3503 -468 3515
rect -680 3447 -665 3503
rect -609 3447 -555 3503
rect -499 3447 -468 3503
rect -680 3393 -468 3447
rect -680 3337 -665 3393
rect -609 3337 -555 3393
rect -499 3337 -468 3393
rect -680 3303 -468 3337
rect -2949 2707 -2861 2795
rect 3867 1127 4079 1150
rect 3867 1071 3889 1127
rect 3945 1071 3999 1127
rect 4055 1071 4079 1127
rect 3867 1017 4079 1071
rect 3867 961 3889 1017
rect 3945 961 3999 1017
rect 4055 961 4079 1017
rect 3867 938 4079 961
rect -661 159 -449 169
rect -661 103 -648 159
rect -592 103 -538 159
rect -482 103 -449 159
rect -661 54 -449 103
rect -661 -2 -648 54
rect -592 -2 -538 54
rect -482 -2 -449 54
rect -661 -51 -449 -2
rect -661 -107 -648 -51
rect -592 -107 -538 -51
rect -482 -107 -449 -51
rect -661 -122 -449 -107
rect -1020 -810 -810 -798
rect -1020 -866 -998 -810
rect -942 -866 -888 -810
rect -832 -866 -810 -810
rect -1020 -920 -810 -866
rect -1020 -976 -998 -920
rect -942 -976 -888 -920
rect -832 -976 -810 -920
rect -1020 -1030 -810 -976
rect -1020 -1086 -998 -1030
rect -942 -1086 -888 -1030
rect -832 -1086 -810 -1030
rect -1020 -1140 -810 -1086
rect -1020 -1196 -998 -1140
rect -942 -1196 -888 -1140
rect -832 -1196 -810 -1140
rect -1020 -1224 -810 -1196
rect -3329 -1482 -2914 -1456
rect -3329 -1538 -3312 -1482
rect -3256 -1538 -3202 -1482
rect -3146 -1538 -3092 -1482
rect -3036 -1538 -2982 -1482
rect -2926 -1538 -2914 -1482
rect -3329 -1592 -2914 -1538
rect -3329 -1648 -3312 -1592
rect -3256 -1648 -3202 -1592
rect -3146 -1648 -3092 -1592
rect -3036 -1648 -2982 -1592
rect -2926 -1648 -2914 -1592
rect -3329 -1681 -2914 -1648
rect -666 -4020 -370 -4002
rect -666 -4076 -653 -4020
rect -597 -4076 -548 -4020
rect -492 -4076 -443 -4020
rect -387 -4076 -370 -4020
rect -666 -4130 -370 -4076
rect -666 -4186 -653 -4130
rect -597 -4186 -548 -4130
rect -492 -4186 -443 -4130
rect -387 -4186 -370 -4130
rect -666 -4214 -370 -4186
rect 3867 -5123 4079 -5100
rect 3867 -5179 3889 -5123
rect 3945 -5179 3999 -5123
rect 4055 -5179 4079 -5123
rect 3867 -5233 4079 -5179
rect 3867 -5289 3889 -5233
rect 3945 -5289 3999 -5233
rect 4055 -5289 4079 -5233
rect 3867 -5312 4079 -5289
rect -680 -7449 -468 -7415
rect -680 -7505 -665 -7449
rect -609 -7505 -555 -7449
rect -499 -7505 -468 -7449
rect -680 -7559 -468 -7505
rect -680 -7615 -665 -7559
rect -609 -7615 -555 -7559
rect -499 -7615 -468 -7559
rect -680 -7627 -468 -7615
<< via3 >>
rect -665 3447 -609 3503
rect -555 3447 -499 3503
rect -665 3337 -609 3393
rect -555 3337 -499 3393
rect 3889 1071 3945 1127
rect 3999 1071 4055 1127
rect 3889 961 3945 1017
rect 3999 961 4055 1017
rect -648 103 -592 159
rect -538 103 -482 159
rect -648 -2 -592 54
rect -538 -2 -482 54
rect -648 -107 -592 -51
rect -538 -107 -482 -51
rect -998 -866 -942 -810
rect -888 -866 -832 -810
rect -998 -976 -942 -920
rect -888 -976 -832 -920
rect -998 -1086 -942 -1030
rect -888 -1086 -832 -1030
rect -998 -1196 -942 -1140
rect -888 -1196 -832 -1140
rect -3312 -1538 -3256 -1482
rect -3202 -1538 -3146 -1482
rect -3092 -1538 -3036 -1482
rect -2982 -1538 -2926 -1482
rect -3312 -1648 -3256 -1592
rect -3202 -1648 -3146 -1592
rect -3092 -1648 -3036 -1592
rect -2982 -1648 -2926 -1592
rect -653 -4076 -597 -4020
rect -548 -4076 -492 -4020
rect -443 -4076 -387 -4020
rect -653 -4186 -597 -4130
rect -548 -4186 -492 -4130
rect -443 -4186 -387 -4130
rect 3889 -5179 3945 -5123
rect 3999 -5179 4055 -5123
rect 3889 -5289 3945 -5233
rect 3999 -5289 4055 -5233
rect -665 -7505 -609 -7449
rect -555 -7505 -499 -7449
rect -665 -7615 -609 -7559
rect -555 -7615 -499 -7559
<< metal4 >>
rect -680 3503 -468 3515
rect -680 3447 -665 3503
rect -609 3447 -555 3503
rect -499 3447 -468 3503
rect -680 3393 -468 3447
rect -680 3337 -665 3393
rect -609 3337 -555 3393
rect -499 3337 -468 3393
rect -680 3303 -468 3337
rect 3867 1127 4079 1150
rect 3867 1071 3889 1127
rect 3945 1071 3999 1127
rect 4055 1071 4079 1127
rect 3867 1017 4079 1071
rect 3867 961 3889 1017
rect 3945 961 3999 1017
rect 4055 961 4079 1017
rect 3867 938 4079 961
rect -661 159 -449 169
rect -661 103 -648 159
rect -592 103 -538 159
rect -482 103 -449 159
rect -661 54 -449 103
rect -661 -2 -648 54
rect -592 -2 -538 54
rect -482 -2 -449 54
rect -661 -51 -449 -2
rect -661 -107 -648 -51
rect -592 -107 -538 -51
rect -482 -107 -449 -51
rect -661 -122 -449 -107
rect -1020 -810 -810 -798
rect -1020 -866 -998 -810
rect -942 -866 -888 -810
rect -832 -866 -810 -810
rect -1020 -920 -810 -866
rect -1020 -976 -998 -920
rect -942 -976 -888 -920
rect -832 -976 -810 -920
rect -1020 -1030 -810 -976
rect -1020 -1086 -998 -1030
rect -942 -1086 -888 -1030
rect -832 -1086 -810 -1030
rect -5409 -2439 -5197 -1100
rect -1020 -1140 -810 -1086
rect -1020 -1196 -998 -1140
rect -942 -1196 -888 -1140
rect -832 -1196 -810 -1140
rect -1020 -1224 -810 -1196
rect -3329 -1482 -2914 -1456
rect -3329 -1538 -3312 -1482
rect -3256 -1538 -3202 -1482
rect -3146 -1538 -3092 -1482
rect -3036 -1538 -2982 -1482
rect -2926 -1538 -2914 -1482
rect -3329 -1592 -2914 -1538
rect -3329 -1648 -3312 -1592
rect -3256 -1648 -3202 -1592
rect -3146 -1648 -3092 -1592
rect -3036 -1648 -2982 -1592
rect -2926 -1648 -2914 -1592
rect -3329 -1681 -2914 -1648
rect -666 -4020 -370 -4002
rect -666 -4076 -653 -4020
rect -597 -4076 -548 -4020
rect -492 -4076 -443 -4020
rect -387 -4076 -370 -4020
rect -666 -4130 -370 -4076
rect -666 -4186 -653 -4130
rect -597 -4186 -548 -4130
rect -492 -4186 -443 -4130
rect -387 -4186 -370 -4130
rect -666 -4214 -370 -4186
rect 3867 -5123 4079 -5100
rect 3867 -5179 3889 -5123
rect 3945 -5179 3999 -5123
rect 4055 -5179 4079 -5123
rect 3867 -5233 4079 -5179
rect 3867 -5289 3889 -5233
rect 3945 -5289 3999 -5233
rect 4055 -5289 4079 -5233
rect 3867 -5312 4079 -5289
rect -680 -7449 -468 -7415
rect -680 -7505 -665 -7449
rect -609 -7505 -555 -7449
rect -499 -7505 -468 -7449
rect -680 -7559 -468 -7505
rect -680 -7615 -665 -7559
rect -609 -7615 -555 -7559
rect -499 -7615 -468 -7559
rect -680 -7627 -468 -7615
<< via4 >>
rect -665 3447 -609 3503
rect -555 3447 -499 3503
rect -665 3337 -609 3393
rect -555 3337 -499 3393
rect 3889 1071 3945 1127
rect 3999 1071 4055 1127
rect 3889 961 3945 1017
rect 3999 961 4055 1017
rect -648 103 -592 159
rect -538 103 -482 159
rect -648 -2 -592 54
rect -538 -2 -482 54
rect -648 -107 -592 -51
rect -538 -107 -482 -51
rect -998 -866 -942 -810
rect -888 -866 -832 -810
rect -998 -976 -942 -920
rect -888 -976 -832 -920
rect -998 -1086 -942 -1030
rect -888 -1086 -832 -1030
rect -998 -1196 -942 -1140
rect -888 -1196 -832 -1140
rect -3312 -1538 -3256 -1482
rect -3202 -1538 -3146 -1482
rect -3092 -1538 -3036 -1482
rect -2982 -1538 -2926 -1482
rect -3312 -1648 -3256 -1592
rect -3202 -1648 -3146 -1592
rect -3092 -1648 -3036 -1592
rect -2982 -1648 -2926 -1592
rect -653 -4076 -597 -4020
rect -548 -4076 -492 -4020
rect -443 -4076 -387 -4020
rect -653 -4186 -597 -4130
rect -548 -4186 -492 -4130
rect -443 -4186 -387 -4130
rect 3889 -5179 3945 -5123
rect 3999 -5179 4055 -5123
rect 3889 -5289 3945 -5233
rect 3999 -5289 4055 -5233
rect -665 -7505 -609 -7449
rect -555 -7505 -499 -7449
rect -665 -7615 -609 -7559
rect -555 -7615 -499 -7559
<< metal5 >>
rect -680 3503 -74 3515
rect -680 3447 -665 3503
rect -609 3447 -555 3503
rect -499 3447 -74 3503
rect -680 3393 -74 3447
rect -680 3337 -665 3393
rect -609 3337 -555 3393
rect -499 3337 -74 3393
rect -680 3303 -74 3337
rect 3892 1150 4049 1517
rect 3867 1127 4079 1150
rect 3867 1071 3889 1127
rect 3945 1071 3999 1127
rect 4055 1071 4079 1127
rect 3867 1017 4079 1071
rect 3867 961 3889 1017
rect 3945 961 3999 1017
rect 4055 961 4079 1017
rect 3867 938 4079 961
rect -661 159 -449 169
rect -661 103 -648 159
rect -592 103 -538 159
rect -482 103 -449 159
rect -661 54 -449 103
rect -661 -2 -648 54
rect -592 -2 -538 54
rect -482 -2 -449 54
rect -661 -51 -449 -2
rect -661 -107 -648 -51
rect -592 -107 -538 -51
rect -482 -107 -449 -51
rect -1276 -796 -1260 -547
rect -1276 -798 -881 -796
rect -1276 -810 -810 -798
rect -1276 -853 -998 -810
rect -1311 -866 -998 -853
rect -942 -866 -888 -810
rect -832 -866 -810 -810
rect -1311 -920 -810 -866
rect -1311 -976 -998 -920
rect -942 -976 -888 -920
rect -832 -976 -810 -920
rect -1311 -1030 -810 -976
rect -7265 -1841 -7053 -1059
rect -1311 -1086 -998 -1030
rect -942 -1086 -888 -1030
rect -832 -1086 -810 -1030
rect -1311 -1140 -810 -1086
rect -1311 -1152 -998 -1140
rect -3328 -1456 -3116 -1184
rect -1020 -1196 -998 -1152
rect -942 -1196 -888 -1140
rect -832 -1196 -810 -1140
rect -1020 -1224 -810 -1196
rect -3329 -1482 -2914 -1456
rect -3329 -1538 -3312 -1482
rect -3256 -1538 -3202 -1482
rect -3146 -1538 -3092 -1482
rect -3036 -1538 -2982 -1482
rect -2926 -1538 -2914 -1482
rect -3329 -1592 -2914 -1538
rect -3329 -1648 -3312 -1592
rect -3256 -1648 -3202 -1592
rect -3146 -1648 -3092 -1592
rect -3036 -1648 -2982 -1592
rect -2926 -1648 -2914 -1592
rect -3329 -1681 -2914 -1648
rect -661 -1841 -449 -107
rect -7268 -2053 -449 -1841
rect -7265 -2529 -7053 -2053
rect -3079 -2387 -2867 -2053
rect -3099 -2468 -2887 -2435
rect -1024 -4020 -370 -4002
rect -1024 -4076 -653 -4020
rect -597 -4076 -548 -4020
rect -492 -4076 -443 -4020
rect -387 -4076 -370 -4020
rect -1024 -4130 -370 -4076
rect -1024 -4186 -653 -4130
rect -597 -4186 -548 -4130
rect -492 -4186 -443 -4130
rect -387 -4186 -370 -4130
rect -1024 -4214 -370 -4186
rect 3867 -5123 4079 -5100
rect 3867 -5179 3889 -5123
rect 3945 -5179 3999 -5123
rect 4055 -5179 4079 -5123
rect 3867 -5233 4079 -5179
rect 3867 -5289 3889 -5233
rect 3945 -5289 3999 -5233
rect 4055 -5289 4079 -5233
rect 3867 -5312 4079 -5289
rect 3897 -5635 4054 -5312
rect -680 -7449 -74 -7415
rect -680 -7505 -665 -7449
rect -609 -7505 -555 -7449
rect -499 -7505 -74 -7449
rect -680 -7559 -74 -7505
rect -680 -7615 -665 -7559
rect -609 -7615 -555 -7559
rect -499 -7615 -74 -7559
rect -680 -7627 -74 -7615
rect -5380 -8976 -5253 -8848
rect -5411 -9070 -5199 -8976
rect -1225 -9070 -1013 -8975
rect -5411 -9282 -1013 -9070
use cap_mim_2p0fF_NEQE26  cap_mim_2p0fF_NEQE26_0
timestamp 1699205295
transform 0 1 3114 1 0 -7401
box -1840 -3400 1840 3400
use cap_mim_2p0fF_NEQE26  cap_mim_2p0fF_NEQE26_1
timestamp 1699205295
transform 1 0 -2853 0 1 -5575
box -1840 -3400 1840 3400
use cap_mim_2p0fF_NEQE26  cap_mim_2p0fF_NEQE26_2
timestamp 1699205295
transform 0 1 3114 -1 0 3289
box -1840 -3400 1840 3400
use cap_mim_2p0fF_NEQE26  cap_mim_2p0fF_NEQE26_3
timestamp 1699205295
transform 1 0 -7039 0 1 2207
box -1840 -3400 1840 3400
use cap_mim_2p0fF_NEQE26  cap_mim_2p0fF_NEQE26_4
timestamp 1699205295
transform 1 0 -7039 0 -1 -5717
box -1840 -3400 1840 3400
use cap_mim_2p0fF_NEQE26  cap_mim_2p0fF_NEQE26_5
timestamp 1699205295
transform 1 0 -3102 0 -1 2216
box -1840 -3400 1840 3400
use ppolyf_u_6V6NLJ  ppolyf_u_6V6NLJ_0
timestamp 1699203423
transform 1 0 1747 0 -1 -2763
box -1824 -516 1824 516
use ppolyf_u_6V6NLJ  ppolyf_u_6V6NLJ_1
timestamp 1699203423
transform 1 0 1747 0 -1 -4597
box -1824 -516 1824 516
use ppolyf_u_6V6NLJ  ppolyf_u_6V6NLJ_2
timestamp 1699203423
transform 1 0 1747 0 -1 -3680
box -1824 -516 1824 516
use ppolyf_u_6V6NLJ  ppolyf_u_6V6NLJ_3
timestamp 1699203423
transform 1 0 1747 0 1 -1349
box -1824 -516 1824 516
use ppolyf_u_6V6NLJ  ppolyf_u_6V6NLJ_4
timestamp 1699203423
transform 1 0 1747 0 1 485
box -1824 -516 1824 516
use ppolyf_u_6V6NLJ  ppolyf_u_6V6NLJ_5
timestamp 1699203423
transform 1 0 1747 0 1 -432
box -1824 -516 1824 516
<< labels >>
flabel metal2 -119 -4152 -119 -4152 0 FreeSans 800 0 0 0 R3_R7
port 3 nsew
flabel metal2 -111 -3198 -111 -3198 0 FreeSans 800 0 0 0 R7_R8_R10_C
port 1 nsew
flabel space -397 -3623 -397 -3623 0 FreeSans 1600 0 0 0 INN_N
port 5 nsew
flabel metal2 -386 -512 -386 -512 0 FreeSans 1600 0 0 0 INN_P
port 7 nsew
flabel metal1 1718 1077 1718 1077 0 FreeSans 1600 0 0 0 VDD
port 8 nsew
flabel metal2 3949 -1295 3949 -1295 0 FreeSans 1600 0 0 0 OP_AMP_IN_P
port 9 nsew
flabel metal2 3928 -2832 3928 -2832 0 FreeSans 1600 0 0 0 OP_AMP_IN_N
port 10 nsew
<< end >>
