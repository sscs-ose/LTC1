magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1045 1019 1045
<< metal1 >>
rect -19 39 19 45
rect -19 -39 -13 39
rect 13 -39 19 39
rect -19 -45 19 -39
<< via1 >>
rect -13 -39 13 39
<< metal2 >>
rect -19 39 19 45
rect -19 -39 -13 39
rect 13 -39 19 39
rect -19 -45 19 -39
<< end >>
