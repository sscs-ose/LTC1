magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -6189 -2222 4082 6087
<< nwell >>
rect -817 1943 -712 1945
rect -511 1943 -452 1961
rect -3723 1885 -2663 1906
rect -817 1905 243 1943
<< psubdiff >>
rect -4178 4057 2072 4075
rect -4178 4011 -4125 4057
rect -4079 4011 -3975 4057
rect -3929 4011 -3825 4057
rect -3779 4011 -3675 4057
rect -3629 4011 -3525 4057
rect -3479 4011 -3375 4057
rect -3329 4011 -3225 4057
rect -3179 4011 -3075 4057
rect -3029 4011 -2925 4057
rect -2879 4011 -2775 4057
rect -2729 4011 -2625 4057
rect -2579 4011 -2475 4057
rect -2429 4011 -2325 4057
rect -2279 4011 -2175 4057
rect -2129 4011 -2025 4057
rect -1979 4011 -1875 4057
rect -1829 4011 -1725 4057
rect -1679 4011 -1575 4057
rect -1529 4011 -1425 4057
rect -1379 4011 -1275 4057
rect -1229 4011 -1125 4057
rect -1079 4011 -975 4057
rect -929 4011 -825 4057
rect -779 4011 -675 4057
rect -629 4011 -525 4057
rect -479 4011 -375 4057
rect -329 4011 -225 4057
rect -179 4011 -75 4057
rect -29 4011 75 4057
rect 121 4011 225 4057
rect 271 4011 375 4057
rect 421 4011 525 4057
rect 571 4011 675 4057
rect 721 4011 825 4057
rect 871 4011 975 4057
rect 1021 4011 1125 4057
rect 1171 4011 1275 4057
rect 1321 4011 1425 4057
rect 1471 4011 1575 4057
rect 1621 4011 1725 4057
rect 1771 4011 1875 4057
rect 1921 4030 2072 4057
rect 1921 4011 2004 4030
rect -4178 3985 2004 4011
rect -4178 3950 -4088 3985
rect -4178 3904 -4158 3950
rect -4112 3904 -4088 3950
rect -4178 3800 -4088 3904
rect -4178 3754 -4158 3800
rect -4112 3754 -4088 3800
rect -4178 3650 -4088 3754
rect -4178 3604 -4158 3650
rect -4112 3604 -4088 3650
rect -4178 3500 -4088 3604
rect -4178 3454 -4158 3500
rect -4112 3454 -4088 3500
rect -4178 3350 -4088 3454
rect -4178 3304 -4158 3350
rect -4112 3304 -4088 3350
rect -4178 3200 -4088 3304
rect -4178 3154 -4158 3200
rect -4112 3154 -4088 3200
rect -4178 3050 -4088 3154
rect -4178 3004 -4158 3050
rect -4112 3004 -4088 3050
rect -4178 2900 -4088 3004
rect -4178 2854 -4158 2900
rect -4112 2854 -4088 2900
rect -4178 2750 -4088 2854
rect -4178 2704 -4158 2750
rect -4112 2704 -4088 2750
rect -4178 2600 -4088 2704
rect -4178 2554 -4158 2600
rect -4112 2554 -4088 2600
rect -4178 2450 -4088 2554
rect -4178 2404 -4158 2450
rect -4112 2404 -4088 2450
rect -4178 2300 -4088 2404
rect -4178 2254 -4158 2300
rect -4112 2254 -4088 2300
rect -4178 2150 -4088 2254
rect -4178 2104 -4158 2150
rect -4112 2104 -4088 2150
rect -4178 2000 -4088 2104
rect -4178 1954 -4158 2000
rect -4112 1954 -4088 2000
rect -4178 1850 -4088 1954
rect -4178 1804 -4158 1850
rect -4112 1804 -4088 1850
rect -4178 1700 -4088 1804
rect -4178 1654 -4158 1700
rect -4112 1654 -4088 1700
rect -4178 1550 -4088 1654
rect -4178 1504 -4158 1550
rect -4112 1504 -4088 1550
rect -4178 1400 -4088 1504
rect -4178 1354 -4158 1400
rect -4112 1354 -4088 1400
rect -4178 1250 -4088 1354
rect -4178 1204 -4158 1250
rect -4112 1204 -4088 1250
rect -4178 1100 -4088 1204
rect -4178 1054 -4158 1100
rect -4112 1054 -4088 1100
rect -4178 950 -4088 1054
rect -4178 904 -4158 950
rect -4112 904 -4088 950
rect -4178 800 -4088 904
rect -4178 754 -4158 800
rect -4112 754 -4088 800
rect -4178 650 -4088 754
rect -4178 604 -4158 650
rect -4112 604 -4088 650
rect -4178 500 -4088 604
rect -4178 454 -4158 500
rect -4112 454 -4088 500
rect -4178 350 -4088 454
rect -4178 304 -4158 350
rect -4112 304 -4088 350
rect -4178 200 -4088 304
rect -4178 154 -4158 200
rect -4112 154 -4088 200
rect -4178 50 -4088 154
rect -4178 4 -4158 50
rect -4112 4 -4088 50
rect -4178 -115 -4088 4
rect 1982 3984 2004 3985
rect 2050 3984 2072 4030
rect 1982 3880 2072 3984
rect 1982 3834 2004 3880
rect 2050 3834 2072 3880
rect 1982 3730 2072 3834
rect 1982 3684 2004 3730
rect 2050 3684 2072 3730
rect 1982 3580 2072 3684
rect 1982 3534 2004 3580
rect 2050 3534 2072 3580
rect 1982 3430 2072 3534
rect 1982 3384 2004 3430
rect 2050 3384 2072 3430
rect 1982 3280 2072 3384
rect 1982 3234 2004 3280
rect 2050 3234 2072 3280
rect 1982 3130 2072 3234
rect 1982 3084 2004 3130
rect 2050 3084 2072 3130
rect 1982 2980 2072 3084
rect 1982 2934 2004 2980
rect 2050 2934 2072 2980
rect 1982 2830 2072 2934
rect 1982 2784 2004 2830
rect 2050 2784 2072 2830
rect 1982 2680 2072 2784
rect 1982 2634 2004 2680
rect 2050 2634 2072 2680
rect 1982 2530 2072 2634
rect 1982 2484 2004 2530
rect 2050 2484 2072 2530
rect 1982 2380 2072 2484
rect 1982 2334 2004 2380
rect 2050 2334 2072 2380
rect 1982 2230 2072 2334
rect 1982 2184 2004 2230
rect 2050 2184 2072 2230
rect 1982 2080 2072 2184
rect 1982 2034 2004 2080
rect 2050 2034 2072 2080
rect 1982 1930 2072 2034
rect 1982 1884 2004 1930
rect 2050 1884 2072 1930
rect 1982 1780 2072 1884
rect 1982 1734 2004 1780
rect 2050 1734 2072 1780
rect 1982 1630 2072 1734
rect 1982 1584 2004 1630
rect 2050 1584 2072 1630
rect 1982 1480 2072 1584
rect 1982 1434 2004 1480
rect 2050 1434 2072 1480
rect 1982 1330 2072 1434
rect 1982 1284 2004 1330
rect 2050 1284 2072 1330
rect 1982 1180 2072 1284
rect 1982 1134 2004 1180
rect 2050 1134 2072 1180
rect 1982 1030 2072 1134
rect 1982 984 2004 1030
rect 2050 984 2072 1030
rect 1982 880 2072 984
rect 1982 834 2004 880
rect 2050 834 2072 880
rect 1982 730 2072 834
rect 1982 684 2004 730
rect 2050 684 2072 730
rect 1982 580 2072 684
rect 1982 534 2004 580
rect 2050 534 2072 580
rect 1982 430 2072 534
rect 1982 384 2004 430
rect 2050 384 2072 430
rect 1982 280 2072 384
rect 1982 234 2004 280
rect 2050 234 2072 280
rect 1982 130 2072 234
rect 1982 84 2004 130
rect 2050 84 2072 130
rect 1982 -20 2072 84
rect 1982 -66 2004 -20
rect 2050 -66 2072 -20
rect 1982 -115 2072 -66
rect -4178 -136 2072 -115
rect -4178 -182 -4058 -136
rect -4012 -182 -3908 -136
rect -3862 -182 -3758 -136
rect -3712 -182 -3608 -136
rect -3562 -182 -3458 -136
rect -3412 -182 -3308 -136
rect -3262 -182 -3158 -136
rect -3112 -182 -3008 -136
rect -2962 -182 -2858 -136
rect -2812 -182 -2708 -136
rect -2662 -182 -2558 -136
rect -2512 -182 -2408 -136
rect -2362 -182 -2258 -136
rect -2212 -182 -2108 -136
rect -2062 -182 -1958 -136
rect -1912 -182 -1808 -136
rect -1762 -182 -1658 -136
rect -1612 -182 -1508 -136
rect -1462 -182 -1358 -136
rect -1312 -182 -1208 -136
rect -1162 -182 -1058 -136
rect -1012 -182 -908 -136
rect -862 -182 -758 -136
rect -712 -182 -608 -136
rect -562 -182 -458 -136
rect -412 -182 -308 -136
rect -262 -182 -158 -136
rect -112 -182 -8 -136
rect 38 -182 142 -136
rect 188 -182 292 -136
rect 338 -182 442 -136
rect 488 -182 592 -136
rect 638 -182 742 -136
rect 788 -182 892 -136
rect 938 -182 1042 -136
rect 1088 -182 1192 -136
rect 1238 -182 1342 -136
rect 1388 -182 1492 -136
rect 1538 -182 1642 -136
rect 1688 -182 1792 -136
rect 1838 -182 1942 -136
rect 1988 -182 2072 -136
rect -4178 -205 2072 -182
<< psubdiffcont >>
rect -4125 4011 -4079 4057
rect -3975 4011 -3929 4057
rect -3825 4011 -3779 4057
rect -3675 4011 -3629 4057
rect -3525 4011 -3479 4057
rect -3375 4011 -3329 4057
rect -3225 4011 -3179 4057
rect -3075 4011 -3029 4057
rect -2925 4011 -2879 4057
rect -2775 4011 -2729 4057
rect -2625 4011 -2579 4057
rect -2475 4011 -2429 4057
rect -2325 4011 -2279 4057
rect -2175 4011 -2129 4057
rect -2025 4011 -1979 4057
rect -1875 4011 -1829 4057
rect -1725 4011 -1679 4057
rect -1575 4011 -1529 4057
rect -1425 4011 -1379 4057
rect -1275 4011 -1229 4057
rect -1125 4011 -1079 4057
rect -975 4011 -929 4057
rect -825 4011 -779 4057
rect -675 4011 -629 4057
rect -525 4011 -479 4057
rect -375 4011 -329 4057
rect -225 4011 -179 4057
rect -75 4011 -29 4057
rect 75 4011 121 4057
rect 225 4011 271 4057
rect 375 4011 421 4057
rect 525 4011 571 4057
rect 675 4011 721 4057
rect 825 4011 871 4057
rect 975 4011 1021 4057
rect 1125 4011 1171 4057
rect 1275 4011 1321 4057
rect 1425 4011 1471 4057
rect 1575 4011 1621 4057
rect 1725 4011 1771 4057
rect 1875 4011 1921 4057
rect -4158 3904 -4112 3950
rect -4158 3754 -4112 3800
rect -4158 3604 -4112 3650
rect -4158 3454 -4112 3500
rect -4158 3304 -4112 3350
rect -4158 3154 -4112 3200
rect -4158 3004 -4112 3050
rect -4158 2854 -4112 2900
rect -4158 2704 -4112 2750
rect -4158 2554 -4112 2600
rect -4158 2404 -4112 2450
rect -4158 2254 -4112 2300
rect -4158 2104 -4112 2150
rect -4158 1954 -4112 2000
rect -4158 1804 -4112 1850
rect -4158 1654 -4112 1700
rect -4158 1504 -4112 1550
rect -4158 1354 -4112 1400
rect -4158 1204 -4112 1250
rect -4158 1054 -4112 1100
rect -4158 904 -4112 950
rect -4158 754 -4112 800
rect -4158 604 -4112 650
rect -4158 454 -4112 500
rect -4158 304 -4112 350
rect -4158 154 -4112 200
rect -4158 4 -4112 50
rect 2004 3984 2050 4030
rect 2004 3834 2050 3880
rect 2004 3684 2050 3730
rect 2004 3534 2050 3580
rect 2004 3384 2050 3430
rect 2004 3234 2050 3280
rect 2004 3084 2050 3130
rect 2004 2934 2050 2980
rect 2004 2784 2050 2830
rect 2004 2634 2050 2680
rect 2004 2484 2050 2530
rect 2004 2334 2050 2380
rect 2004 2184 2050 2230
rect 2004 2034 2050 2080
rect 2004 1884 2050 1930
rect 2004 1734 2050 1780
rect 2004 1584 2050 1630
rect 2004 1434 2050 1480
rect 2004 1284 2050 1330
rect 2004 1134 2050 1180
rect 2004 984 2050 1030
rect 2004 834 2050 880
rect 2004 684 2050 730
rect 2004 534 2050 580
rect 2004 384 2050 430
rect 2004 234 2050 280
rect 2004 84 2050 130
rect 2004 -66 2050 -20
rect -4058 -182 -4012 -136
rect -3908 -182 -3862 -136
rect -3758 -182 -3712 -136
rect -3608 -182 -3562 -136
rect -3458 -182 -3412 -136
rect -3308 -182 -3262 -136
rect -3158 -182 -3112 -136
rect -3008 -182 -2962 -136
rect -2858 -182 -2812 -136
rect -2708 -182 -2662 -136
rect -2558 -182 -2512 -136
rect -2408 -182 -2362 -136
rect -2258 -182 -2212 -136
rect -2108 -182 -2062 -136
rect -1958 -182 -1912 -136
rect -1808 -182 -1762 -136
rect -1658 -182 -1612 -136
rect -1508 -182 -1462 -136
rect -1358 -182 -1312 -136
rect -1208 -182 -1162 -136
rect -1058 -182 -1012 -136
rect -908 -182 -862 -136
rect -758 -182 -712 -136
rect -608 -182 -562 -136
rect -458 -182 -412 -136
rect -308 -182 -262 -136
rect -158 -182 -112 -136
rect -8 -182 38 -136
rect 142 -182 188 -136
rect 292 -182 338 -136
rect 442 -182 488 -136
rect 592 -182 638 -136
rect 742 -182 788 -136
rect 892 -182 938 -136
rect 1042 -182 1088 -136
rect 1192 -182 1238 -136
rect 1342 -182 1388 -136
rect 1492 -182 1538 -136
rect 1642 -182 1688 -136
rect 1792 -182 1838 -136
rect 1942 -182 1988 -136
<< metal1 >>
rect -4189 4057 2082 4087
rect -4189 4011 -4125 4057
rect -4079 4011 -3975 4057
rect -3929 4011 -3825 4057
rect -3779 4011 -3675 4057
rect -3629 4011 -3525 4057
rect -3479 4011 -3375 4057
rect -3329 4011 -3225 4057
rect -3179 4011 -3075 4057
rect -3029 4011 -2925 4057
rect -2879 4011 -2775 4057
rect -2729 4011 -2625 4057
rect -2579 4011 -2475 4057
rect -2429 4011 -2325 4057
rect -2279 4011 -2175 4057
rect -2129 4011 -2025 4057
rect -1979 4011 -1875 4057
rect -1829 4011 -1725 4057
rect -1679 4011 -1575 4057
rect -1529 4011 -1425 4057
rect -1379 4011 -1275 4057
rect -1229 4011 -1125 4057
rect -1079 4011 -975 4057
rect -929 4011 -825 4057
rect -779 4011 -675 4057
rect -629 4011 -525 4057
rect -479 4011 -375 4057
rect -329 4011 -225 4057
rect -179 4011 -75 4057
rect -29 4011 75 4057
rect 121 4011 225 4057
rect 271 4011 375 4057
rect 421 4011 525 4057
rect 571 4011 675 4057
rect 721 4011 825 4057
rect 871 4011 975 4057
rect 1021 4011 1125 4057
rect 1171 4011 1275 4057
rect 1321 4011 1425 4057
rect 1471 4011 1575 4057
rect 1621 4011 1725 4057
rect 1771 4011 1875 4057
rect 1921 4030 2082 4057
rect 1921 4011 2004 4030
rect -4189 3984 2004 4011
rect 2050 3984 2082 4030
rect -4189 3964 2082 3984
rect -4189 3950 -4066 3964
rect -4189 3904 -4158 3950
rect -4112 3904 -4066 3950
rect -4189 3800 -4066 3904
rect -1211 3884 -1137 3916
rect -4189 3754 -4158 3800
rect -4112 3754 -4066 3800
rect -1227 3863 -1119 3884
rect -1227 3811 -1200 3863
rect -1148 3811 -1119 3863
rect -1227 3790 -1119 3811
rect 1959 3880 2082 3964
rect 1959 3834 2004 3880
rect 2050 3834 2082 3880
rect -4189 3650 -4066 3754
rect 1959 3730 2082 3834
rect -4189 3604 -4158 3650
rect -4112 3604 -4066 3650
rect -2895 3671 -2836 3673
rect -2895 3619 -2892 3671
rect -2840 3619 -2836 3671
rect -2895 3617 -2836 3619
rect -2780 3609 -2240 3668
rect -2057 3653 -1571 3670
rect -2057 3651 -1659 3653
rect -2057 3647 -1848 3651
rect -4189 3500 -4066 3604
rect -2057 3595 -2043 3647
rect -1991 3599 -1848 3647
rect -1796 3601 -1659 3651
rect -1607 3601 -1571 3653
rect -1299 3642 -759 3701
rect 93 3648 633 3707
rect 1959 3684 2004 3730
rect 2050 3684 2082 3730
rect 679 3672 777 3677
rect 1049 3674 1147 3679
rect 673 3660 987 3672
rect -1796 3599 -1571 3601
rect -1991 3595 -1571 3599
rect -2057 3573 -1571 3595
rect 673 3608 694 3660
rect 746 3653 987 3660
rect 746 3608 877 3653
rect 673 3601 877 3608
rect 929 3601 987 3653
rect 673 3582 987 3601
rect 1049 3664 1095 3674
rect 1049 3662 1120 3664
rect 1049 3610 1064 3662
rect 1116 3628 1120 3662
rect 1141 3628 1147 3674
rect 1116 3610 1147 3628
rect 1049 3594 1147 3610
rect 1249 3674 1347 3679
rect 1249 3664 1295 3674
rect 1249 3662 1320 3664
rect 1249 3610 1264 3662
rect 1316 3628 1320 3662
rect 1341 3628 1347 3674
rect 1316 3610 1347 3628
rect 1249 3594 1347 3610
rect 1959 3580 2082 3684
rect -4189 3454 -4158 3500
rect -4112 3454 -4066 3500
rect -4189 3350 -4066 3454
rect -4189 3304 -4158 3350
rect -4112 3304 -4066 3350
rect 1959 3534 2004 3580
rect 2050 3534 2082 3580
rect 1959 3430 2082 3534
rect 1959 3384 2004 3430
rect 2050 3384 2082 3430
rect -1224 3325 -1116 3335
rect 489 3333 574 3346
rect -4189 3200 -4066 3304
rect -1323 3315 -827 3325
rect -4189 3154 -4158 3200
rect -4112 3154 -4066 3200
rect -3721 3187 -3618 3233
rect -2652 3224 -2233 3270
rect -1323 3263 -1200 3315
rect -1148 3263 -827 3315
rect -1323 3253 -827 3263
rect 489 3323 709 3333
rect 489 3271 511 3323
rect 563 3271 709 3323
rect 1959 3280 2082 3384
rect 489 3261 709 3271
rect 489 3259 574 3261
rect -1224 3241 -1116 3253
rect 1588 3232 1858 3278
rect 1959 3234 2004 3280
rect 2050 3234 2082 3280
rect -4189 3050 -4066 3154
rect -4189 3004 -4158 3050
rect -4112 3004 -4066 3050
rect -4189 2900 -4066 3004
rect -4189 2854 -4158 2900
rect -4112 2854 -4066 2900
rect -4189 2750 -4066 2854
rect 1959 3130 2082 3234
rect 1959 3084 2004 3130
rect 2050 3084 2082 3130
rect 1959 2980 2082 3084
rect 1959 2934 2004 2980
rect 2050 2934 2082 2980
rect 1959 2830 2082 2934
rect 1959 2784 2004 2830
rect 2050 2784 2082 2830
rect -4189 2704 -4158 2750
rect -4112 2704 -4066 2750
rect -1144 2726 -1068 2748
rect -4189 2600 -4066 2704
rect -4189 2554 -4158 2600
rect -4112 2554 -4066 2600
rect -4189 2450 -4066 2554
rect -4189 2404 -4158 2450
rect -4112 2404 -4066 2450
rect -4189 2300 -4066 2404
rect -4189 2254 -4158 2300
rect -4112 2254 -4066 2300
rect -4189 2150 -4066 2254
rect -4189 2104 -4158 2150
rect -4112 2104 -4066 2150
rect -4189 2000 -4066 2104
rect -4189 1954 -4158 2000
rect -4112 1954 -4066 2000
rect -4189 1850 -4066 1954
rect -4189 1804 -4158 1850
rect -4112 1804 -4066 1850
rect -4189 1700 -4066 1804
rect -4189 1654 -4158 1700
rect -4112 1654 -4066 1700
rect -4189 1550 -4066 1654
rect -4189 1504 -4158 1550
rect -4112 1504 -4066 1550
rect -4189 1400 -4066 1504
rect -4189 1354 -4158 1400
rect -4112 1354 -4066 1400
rect -4189 1250 -4066 1354
rect -4189 1204 -4158 1250
rect -4112 1204 -4066 1250
rect -4189 1100 -4066 1204
rect -4189 1054 -4158 1100
rect -4112 1054 -4066 1100
rect -3945 1877 -3848 2722
rect -1144 2674 -1130 2726
rect -1078 2674 -1068 2726
rect -2363 2645 -2096 2674
rect -1144 2658 -1068 2674
rect -738 2727 -652 2744
rect -738 2675 -720 2727
rect -668 2675 -652 2727
rect -738 2659 -652 2675
rect -2363 2641 -2185 2645
rect -2363 2589 -2337 2641
rect -2285 2593 -2185 2641
rect -2133 2593 -2096 2645
rect -2285 2589 -2096 2593
rect -2363 2559 -2096 2589
rect -1754 2629 -1389 2656
rect -1754 2577 -1737 2629
rect -1685 2623 -1458 2629
rect -1685 2577 -1597 2623
rect -1754 2571 -1597 2577
rect -1545 2577 -1458 2623
rect -1406 2577 -1389 2629
rect -1545 2571 -1389 2577
rect -1754 2549 -1389 2571
rect -2666 2389 -2358 2444
rect -3767 2244 -3603 2261
rect -3767 2192 -3723 2244
rect -3671 2192 -3603 2244
rect -3767 2113 -3603 2192
rect -2413 2176 -2358 2389
rect -2413 2162 -2314 2176
rect -3767 2086 -3583 2113
rect -2413 2110 -2377 2162
rect -2325 2110 -2314 2162
rect -2413 2108 -2314 2110
rect -2380 2097 -2314 2108
rect -3767 2034 -3733 2086
rect -3681 2034 -3583 2086
rect -3767 2011 -3583 2034
rect -2509 2014 -2424 2029
rect -3767 2010 -3603 2011
rect -2509 1962 -2493 2014
rect -2441 1962 -2424 2014
rect -2509 1958 -2424 1962
rect -3723 1885 -2663 1906
rect -3945 1825 -3923 1877
rect -3871 1825 -3848 1877
rect -3945 1167 -3848 1825
rect -2495 1407 -2440 1958
rect -1134 1932 -1071 2658
rect -667 1964 -283 1982
rect -667 1961 -364 1964
rect -667 1957 -506 1961
rect -2327 1877 -2250 1909
rect -1293 1887 -1071 1932
rect -817 1943 -712 1945
rect -667 1943 -634 1957
rect -817 1905 -634 1943
rect -582 1909 -506 1957
rect -454 1912 -364 1961
rect -312 1943 -283 1964
rect -312 1912 243 1943
rect -454 1909 243 1912
rect -582 1905 243 1909
rect 324 1911 421 2761
rect 1959 2680 2082 2784
rect 1959 2634 2004 2680
rect 2050 2634 2082 2680
rect 494 2518 663 2532
rect 1959 2530 2082 2634
rect 494 2516 687 2518
rect 494 2464 631 2516
rect 683 2464 687 2516
rect 494 2462 687 2464
rect 1959 2484 2004 2530
rect 2050 2484 2082 2530
rect 494 2395 663 2462
rect 494 2343 525 2395
rect 577 2343 663 2395
rect 494 2320 663 2343
rect 1959 2380 2082 2484
rect 1959 2334 2004 2380
rect 2050 2334 2082 2380
rect 494 2275 735 2320
rect 494 2223 523 2275
rect 575 2223 735 2275
rect 494 2193 735 2223
rect 1959 2230 2082 2334
rect 1959 2184 2004 2230
rect 2050 2184 2082 2230
rect 1959 2080 2082 2184
rect 1959 2034 2004 2080
rect 2050 2034 2082 2080
rect 1753 1954 1854 1968
rect 1753 1940 1775 1954
rect -667 1888 -283 1905
rect -1293 1886 -1087 1887
rect -2327 1825 -2317 1877
rect -2265 1825 -2250 1877
rect -2327 1807 -2250 1825
rect -2153 1499 -1730 1521
rect -2153 1491 -1818 1499
rect -2153 1439 -2136 1491
rect -2084 1489 -1818 1491
rect -2084 1439 -1976 1489
rect -2153 1437 -1976 1439
rect -1924 1447 -1818 1489
rect -1766 1447 -1730 1499
rect -1924 1437 -1730 1447
rect -2153 1421 -1730 1437
rect -2666 1352 -2440 1407
rect -3945 1070 -3753 1167
rect -4189 950 -4066 1054
rect -1133 1033 -1087 1886
rect 324 1839 688 1911
rect 1600 1902 1775 1940
rect 1827 1902 1854 1954
rect 1600 1894 1854 1902
rect 1743 1879 1854 1894
rect 1959 1930 2082 2034
rect 1959 1884 2004 1930
rect 2050 1884 2082 1930
rect -908 1430 -833 1449
rect -908 1378 -901 1430
rect -849 1378 -833 1430
rect -908 1359 -833 1378
rect 324 1188 421 1839
rect 902 1524 1288 1532
rect 902 1507 1291 1524
rect 902 1502 1208 1507
rect 902 1487 1045 1502
rect 902 1435 921 1487
rect 973 1450 1045 1487
rect 1097 1455 1208 1502
rect 1260 1455 1291 1507
rect 1097 1450 1291 1455
rect 973 1439 1291 1450
rect 973 1435 1288 1439
rect 902 1425 1288 1435
rect 273 1091 421 1188
rect 1743 1067 1815 1879
rect -4189 904 -4158 950
rect -4112 904 -4066 950
rect -4189 800 -4066 904
rect -4189 754 -4158 800
rect -4112 754 -4066 800
rect -4189 650 -4066 754
rect -4189 604 -4158 650
rect -4112 604 -4066 650
rect -2465 958 -2263 1004
rect -1283 987 -1087 1033
rect 563 1007 615 1018
rect 361 961 615 1007
rect 1570 995 1815 1067
rect 1959 1780 2082 1884
rect 1959 1734 2004 1780
rect 2050 1734 2082 1780
rect 1959 1630 2082 1734
rect 1959 1584 2004 1630
rect 2050 1584 2082 1630
rect 1959 1480 2082 1584
rect 1959 1434 2004 1480
rect 2050 1434 2082 1480
rect 1959 1330 2082 1434
rect 1959 1284 2004 1330
rect 2050 1284 2082 1330
rect 1959 1180 2082 1284
rect 1959 1134 2004 1180
rect 2050 1134 2082 1180
rect 1959 1030 2082 1134
rect -4189 500 -4066 604
rect -4189 454 -4158 500
rect -4112 454 -4066 500
rect -4189 350 -4066 454
rect -4189 304 -4158 350
rect -4112 304 -4066 350
rect -4189 200 -4066 304
rect -4189 154 -4158 200
rect -4112 154 -4066 200
rect -4189 50 -4066 154
rect -4189 4 -4158 50
rect -4112 4 -4066 50
rect -4189 -99 -4066 4
rect -3722 559 -3618 605
rect -3722 35 -3676 559
rect -3198 170 -2820 183
rect -3198 162 -2888 170
rect -3198 110 -3180 162
rect -3128 159 -2888 162
rect -3128 110 -3045 159
rect -3198 107 -3045 110
rect -2993 118 -2888 159
rect -2836 118 -2820 170
rect -2993 107 -2820 118
rect -3198 89 -2820 107
rect -2465 35 -2419 958
rect 361 626 407 961
rect 563 957 615 961
rect 1959 984 2004 1030
rect 2050 984 2082 1030
rect 138 580 407 626
rect 1959 880 2082 984
rect 1959 834 2004 880
rect 2050 834 2082 880
rect 1959 730 2082 834
rect 1959 684 2004 730
rect 2050 684 2082 730
rect 1959 580 2082 684
rect 1959 534 2004 580
rect 2050 534 2082 580
rect -1581 407 -1170 430
rect -1581 404 -1263 407
rect -1581 352 -1559 404
rect -1507 399 -1263 404
rect -1507 352 -1438 399
rect -1581 347 -1438 352
rect -1386 355 -1263 399
rect -1211 355 -1170 407
rect -1386 347 -1170 355
rect -1581 328 -1170 347
rect 370 406 756 432
rect 370 405 553 406
rect 370 353 406 405
rect 458 354 553 405
rect 605 400 756 406
rect 605 354 681 400
rect 458 353 681 354
rect 370 348 681 353
rect 733 348 756 400
rect 370 325 756 348
rect 1959 430 2082 534
rect 1959 384 2004 430
rect 2050 384 2082 430
rect 1959 280 2082 384
rect 1959 234 2004 280
rect 2050 234 2082 280
rect -679 206 -141 213
rect -679 204 -139 206
rect -679 152 -671 204
rect -619 189 -139 204
rect -619 167 -222 189
rect -619 152 -484 167
rect -679 115 -484 152
rect -432 137 -222 167
rect -170 137 -139 189
rect -432 121 -139 137
rect 1959 130 2082 234
rect -432 115 -141 121
rect -679 113 -141 115
rect -499 99 -401 113
rect -3722 -11 -2419 35
rect 1959 84 2004 130
rect 2050 84 2082 130
rect 1959 -20 2082 84
rect 1959 -66 2004 -20
rect 2050 -66 2082 -20
rect 1959 -99 2082 -66
rect -4189 -136 2082 -99
rect -4189 -182 -4058 -136
rect -4012 -182 -3908 -136
rect -3862 -182 -3758 -136
rect -3712 -182 -3608 -136
rect -3562 -182 -3458 -136
rect -3412 -182 -3308 -136
rect -3262 -182 -3158 -136
rect -3112 -182 -3008 -136
rect -2962 -182 -2858 -136
rect -2812 -182 -2708 -136
rect -2662 -182 -2558 -136
rect -2512 -182 -2408 -136
rect -2362 -182 -2258 -136
rect -2212 -182 -2108 -136
rect -2062 -182 -1958 -136
rect -1912 -182 -1808 -136
rect -1762 -182 -1658 -136
rect -1612 -182 -1508 -136
rect -1462 -182 -1358 -136
rect -1312 -182 -1208 -136
rect -1162 -182 -1058 -136
rect -1012 -182 -908 -136
rect -862 -182 -758 -136
rect -712 -182 -608 -136
rect -562 -182 -458 -136
rect -412 -182 -308 -136
rect -262 -182 -158 -136
rect -112 -182 -8 -136
rect 38 -182 142 -136
rect 188 -182 292 -136
rect 338 -182 442 -136
rect 488 -182 592 -136
rect 638 -182 742 -136
rect 788 -182 892 -136
rect 938 -182 1042 -136
rect 1088 -182 1192 -136
rect 1238 -182 1342 -136
rect 1388 -182 1492 -136
rect 1538 -182 1642 -136
rect 1688 -182 1792 -136
rect 1838 -182 1942 -136
rect 1988 -182 2082 -136
rect -4189 -221 2082 -182
rect -3706 -222 2082 -221
<< via1 >>
rect -1200 3811 -1148 3863
rect -2892 3619 -2840 3671
rect -2043 3595 -1991 3647
rect -1848 3599 -1796 3651
rect -1659 3601 -1607 3653
rect 694 3608 746 3660
rect 877 3601 929 3653
rect 1064 3610 1116 3662
rect 1264 3610 1316 3662
rect -1200 3263 -1148 3315
rect 511 3271 563 3323
rect -1130 2674 -1078 2726
rect -720 2675 -668 2727
rect -2337 2589 -2285 2641
rect -2185 2593 -2133 2645
rect -1737 2577 -1685 2629
rect -1597 2571 -1545 2623
rect -1458 2577 -1406 2629
rect -3723 2192 -3671 2244
rect -2377 2110 -2325 2162
rect -3733 2034 -3681 2086
rect -2493 1962 -2441 2014
rect -3923 1825 -3871 1877
rect -634 1905 -582 1957
rect -506 1909 -454 1961
rect -364 1912 -312 1964
rect 631 2464 683 2516
rect 525 2343 577 2395
rect 523 2223 575 2275
rect -2317 1825 -2265 1877
rect -2136 1439 -2084 1491
rect -1976 1437 -1924 1489
rect -1818 1447 -1766 1499
rect 1775 1902 1827 1954
rect -901 1378 -849 1430
rect 921 1435 973 1487
rect 1045 1450 1097 1502
rect 1208 1455 1260 1507
rect -3180 110 -3128 162
rect -3045 107 -2993 159
rect -2888 118 -2836 170
rect -1559 352 -1507 404
rect -1438 347 -1386 399
rect -1263 355 -1211 407
rect 406 353 458 405
rect 553 354 605 406
rect 681 348 733 400
rect -671 152 -619 204
rect -484 115 -432 167
rect -222 137 -170 189
<< metal2 >>
rect -1227 3863 -1119 3884
rect -1227 3811 -1200 3863
rect -1148 3811 -1119 3863
rect -1227 3801 -1119 3811
rect -2495 3790 -1119 3801
rect -2495 3745 -1138 3790
rect -2907 3673 -2822 3685
rect -2907 3617 -2894 3673
rect -2838 3617 -2822 3673
rect -2907 3603 -2822 3617
rect -3767 2246 -3603 2261
rect -3767 2190 -3725 2246
rect -3669 2190 -3603 2246
rect -3767 2088 -3603 2190
rect -3767 2032 -3735 2088
rect -3679 2032 -3603 2088
rect -3767 2010 -3603 2032
rect -2495 2029 -2439 3745
rect -2057 3661 -1571 3670
rect -2058 3655 -1571 3661
rect -2058 3653 -1661 3655
rect -2058 3649 -1850 3653
rect -2058 3593 -2045 3649
rect -1989 3597 -1850 3649
rect -1794 3599 -1661 3653
rect -1605 3599 -1571 3655
rect -1794 3597 -1571 3599
rect -1989 3593 -1571 3597
rect -2058 3579 -1571 3593
rect -2057 3573 -1571 3579
rect -1210 3335 -1138 3745
rect 679 3672 764 3674
rect 673 3662 987 3672
rect 673 3606 692 3662
rect 748 3655 987 3662
rect 748 3606 875 3655
rect 673 3599 875 3606
rect 931 3599 987 3655
rect 673 3582 987 3599
rect 1049 3664 1134 3676
rect 1049 3608 1062 3664
rect 1118 3608 1134 3664
rect 1049 3594 1134 3608
rect 1249 3664 1334 3676
rect 1249 3608 1262 3664
rect 1318 3608 1334 3664
rect 1249 3594 1334 3608
rect -1224 3315 -1116 3335
rect -1224 3263 -1200 3315
rect -1148 3263 -1116 3315
rect -1224 3241 -1116 3263
rect 489 3323 574 3346
rect 489 3271 511 3323
rect 563 3271 574 3323
rect 489 3259 574 3271
rect -1144 2732 -1068 2748
rect -738 2732 -652 2744
rect -1144 2727 -652 2732
rect -1144 2726 -720 2727
rect -1144 2674 -1130 2726
rect -1078 2675 -720 2726
rect -668 2675 -652 2727
rect -1078 2674 -652 2675
rect -2363 2647 -2096 2674
rect -1144 2669 -652 2674
rect -1144 2658 -1068 2669
rect -738 2659 -652 2669
rect 501 2658 573 3259
rect -2363 2643 -2187 2647
rect -2363 2587 -2339 2643
rect -2283 2591 -2187 2643
rect -2131 2591 -2096 2647
rect -2283 2587 -2096 2591
rect -2363 2559 -2096 2587
rect -1754 2643 -1389 2656
rect -1754 2631 -1388 2643
rect -1754 2575 -1739 2631
rect -1683 2625 -1460 2631
rect -1683 2575 -1599 2625
rect -1754 2569 -1599 2575
rect -1543 2575 -1460 2625
rect -1404 2575 -1388 2631
rect 501 2589 1837 2658
rect 879 2586 1837 2589
rect -1543 2569 -1388 2575
rect -1754 2561 -1388 2569
rect -1754 2549 -1389 2561
rect 494 2530 663 2532
rect 494 2518 701 2530
rect 494 2462 629 2518
rect 685 2462 701 2518
rect 494 2448 701 2462
rect 494 2397 663 2448
rect 494 2341 523 2397
rect 579 2341 663 2397
rect 494 2277 663 2341
rect 494 2221 521 2277
rect 577 2221 663 2277
rect 494 2193 663 2221
rect -2380 2167 -2314 2176
rect -2380 2162 -939 2167
rect -2380 2110 -2377 2162
rect -2325 2110 -939 2162
rect -2380 2102 -939 2110
rect -2380 2097 -2314 2102
rect -2509 2014 -2424 2029
rect -2509 1962 -2493 2014
rect -2441 1962 -2424 2014
rect -2509 1958 -2424 1962
rect -3941 1880 -3865 1892
rect -2327 1880 -2250 1909
rect -3941 1877 -2250 1880
rect -3941 1825 -3923 1877
rect -3871 1825 -2317 1877
rect -2265 1825 -2250 1877
rect -3941 1822 -2250 1825
rect -3941 1811 -3865 1822
rect -2327 1807 -2250 1822
rect -2153 1501 -1730 1521
rect -2153 1493 -1820 1501
rect -2153 1437 -2138 1493
rect -2082 1491 -1820 1493
rect -2082 1437 -1978 1491
rect -1922 1445 -1820 1491
rect -1764 1445 -1730 1501
rect -2153 1435 -1978 1437
rect -1922 1435 -1730 1445
rect -2153 1421 -1730 1435
rect -1004 1449 -939 2102
rect -667 1966 -283 1982
rect 1765 1968 1837 2586
rect -667 1963 -366 1966
rect -667 1959 -508 1963
rect -667 1903 -636 1959
rect -580 1907 -508 1959
rect -452 1910 -366 1963
rect -310 1910 -283 1966
rect -452 1907 -283 1910
rect -580 1903 -283 1907
rect -667 1888 -283 1903
rect 1753 1954 1854 1968
rect 1753 1902 1775 1954
rect 1827 1902 1854 1954
rect 1753 1879 1854 1902
rect 902 1509 1288 1532
rect 902 1504 1206 1509
rect 902 1489 1043 1504
rect -1004 1430 -833 1449
rect -1004 1378 -901 1430
rect -849 1378 -833 1430
rect 902 1433 919 1489
rect 975 1448 1043 1489
rect 1099 1453 1206 1504
rect 1262 1453 1288 1509
rect 1099 1448 1288 1453
rect 975 1433 1288 1448
rect 902 1425 1288 1433
rect 906 1419 991 1425
rect -1004 1372 -833 1378
rect -912 1359 -833 1372
rect -1581 409 -1170 430
rect -1581 406 -1265 409
rect -1581 350 -1561 406
rect -1505 401 -1265 406
rect -1505 350 -1440 401
rect -1581 345 -1440 350
rect -1384 353 -1265 401
rect -1209 353 -1170 409
rect -1384 345 -1170 353
rect -1581 328 -1170 345
rect 370 408 756 432
rect 370 407 551 408
rect 370 351 404 407
rect 460 352 551 407
rect 607 402 756 408
rect 607 352 679 402
rect 460 351 679 352
rect 370 346 679 351
rect 735 346 756 402
rect 370 325 756 346
rect -686 211 -601 218
rect -686 206 -150 211
rect -2903 183 -2818 184
rect -3187 176 -2803 183
rect -3195 172 -2803 176
rect -3195 164 -2890 172
rect -3195 108 -3182 164
rect -3126 161 -2890 164
rect -3126 108 -3047 161
rect -3195 105 -3047 108
rect -2991 116 -2890 161
rect -2834 116 -2803 172
rect -686 150 -673 206
rect -617 191 -150 206
rect -617 169 -224 191
rect -617 150 -486 169
rect -686 136 -486 150
rect -2991 105 -2803 116
rect -679 113 -486 136
rect -430 135 -224 169
rect -168 135 -150 191
rect -430 113 -150 135
rect -3195 94 -2803 105
rect -499 99 -414 113
rect -3187 74 -2803 94
<< via2 >>
rect -2894 3671 -2838 3673
rect -2894 3619 -2892 3671
rect -2892 3619 -2840 3671
rect -2840 3619 -2838 3671
rect -2894 3617 -2838 3619
rect -3725 2244 -3669 2246
rect -3725 2192 -3723 2244
rect -3723 2192 -3671 2244
rect -3671 2192 -3669 2244
rect -3725 2190 -3669 2192
rect -3735 2086 -3679 2088
rect -3735 2034 -3733 2086
rect -3733 2034 -3681 2086
rect -3681 2034 -3679 2086
rect -3735 2032 -3679 2034
rect -1661 3653 -1605 3655
rect -1850 3651 -1794 3653
rect -2045 3647 -1989 3649
rect -2045 3595 -2043 3647
rect -2043 3595 -1991 3647
rect -1991 3595 -1989 3647
rect -1850 3599 -1848 3651
rect -1848 3599 -1796 3651
rect -1796 3599 -1794 3651
rect -1661 3601 -1659 3653
rect -1659 3601 -1607 3653
rect -1607 3601 -1605 3653
rect -1661 3599 -1605 3601
rect -1850 3597 -1794 3599
rect -2045 3593 -1989 3595
rect 692 3660 748 3662
rect 692 3608 694 3660
rect 694 3608 746 3660
rect 746 3608 748 3660
rect 692 3606 748 3608
rect 875 3653 931 3655
rect 875 3601 877 3653
rect 877 3601 929 3653
rect 929 3601 931 3653
rect 875 3599 931 3601
rect 1062 3662 1118 3664
rect 1062 3610 1064 3662
rect 1064 3610 1116 3662
rect 1116 3610 1118 3662
rect 1062 3608 1118 3610
rect 1262 3662 1318 3664
rect 1262 3610 1264 3662
rect 1264 3610 1316 3662
rect 1316 3610 1318 3662
rect 1262 3608 1318 3610
rect -2187 2645 -2131 2647
rect -2339 2641 -2283 2643
rect -2339 2589 -2337 2641
rect -2337 2589 -2285 2641
rect -2285 2589 -2283 2641
rect -2187 2593 -2185 2645
rect -2185 2593 -2133 2645
rect -2133 2593 -2131 2645
rect -2187 2591 -2131 2593
rect -2339 2587 -2283 2589
rect -1739 2629 -1683 2631
rect -1739 2577 -1737 2629
rect -1737 2577 -1685 2629
rect -1685 2577 -1683 2629
rect -1460 2629 -1404 2631
rect -1739 2575 -1683 2577
rect -1599 2623 -1543 2625
rect -1599 2571 -1597 2623
rect -1597 2571 -1545 2623
rect -1545 2571 -1543 2623
rect -1460 2577 -1458 2629
rect -1458 2577 -1406 2629
rect -1406 2577 -1404 2629
rect -1460 2575 -1404 2577
rect -1599 2569 -1543 2571
rect 629 2516 685 2518
rect 629 2464 631 2516
rect 631 2464 683 2516
rect 683 2464 685 2516
rect 629 2462 685 2464
rect 523 2395 579 2397
rect 523 2343 525 2395
rect 525 2343 577 2395
rect 577 2343 579 2395
rect 523 2341 579 2343
rect 521 2275 577 2277
rect 521 2223 523 2275
rect 523 2223 575 2275
rect 575 2223 577 2275
rect 521 2221 577 2223
rect -1820 1499 -1764 1501
rect -2138 1491 -2082 1493
rect -2138 1439 -2136 1491
rect -2136 1439 -2084 1491
rect -2084 1439 -2082 1491
rect -2138 1437 -2082 1439
rect -1978 1489 -1922 1491
rect -1978 1437 -1976 1489
rect -1976 1437 -1924 1489
rect -1924 1437 -1922 1489
rect -1820 1447 -1818 1499
rect -1818 1447 -1766 1499
rect -1766 1447 -1764 1499
rect -1820 1445 -1764 1447
rect -1978 1435 -1922 1437
rect -366 1964 -310 1966
rect -508 1961 -452 1963
rect -636 1957 -580 1959
rect -636 1905 -634 1957
rect -634 1905 -582 1957
rect -582 1905 -580 1957
rect -508 1909 -506 1961
rect -506 1909 -454 1961
rect -454 1909 -452 1961
rect -366 1912 -364 1964
rect -364 1912 -312 1964
rect -312 1912 -310 1964
rect -366 1910 -310 1912
rect -508 1907 -452 1909
rect -636 1903 -580 1905
rect 1206 1507 1262 1509
rect 1043 1502 1099 1504
rect 919 1487 975 1489
rect 919 1435 921 1487
rect 921 1435 973 1487
rect 973 1435 975 1487
rect 1043 1450 1045 1502
rect 1045 1450 1097 1502
rect 1097 1450 1099 1502
rect 1206 1455 1208 1507
rect 1208 1455 1260 1507
rect 1260 1455 1262 1507
rect 1206 1453 1262 1455
rect 1043 1448 1099 1450
rect 919 1433 975 1435
rect -1265 407 -1209 409
rect -1561 404 -1505 406
rect -1561 352 -1559 404
rect -1559 352 -1507 404
rect -1507 352 -1505 404
rect -1561 350 -1505 352
rect -1440 399 -1384 401
rect -1440 347 -1438 399
rect -1438 347 -1386 399
rect -1386 347 -1384 399
rect -1265 355 -1263 407
rect -1263 355 -1211 407
rect -1211 355 -1209 407
rect -1265 353 -1209 355
rect -1440 345 -1384 347
rect 404 405 460 407
rect 404 353 406 405
rect 406 353 458 405
rect 458 353 460 405
rect 404 351 460 353
rect 551 406 607 408
rect 551 354 553 406
rect 553 354 605 406
rect 605 354 607 406
rect 551 352 607 354
rect 679 400 735 402
rect 679 348 681 400
rect 681 348 733 400
rect 733 348 735 400
rect 679 346 735 348
rect -2890 170 -2834 172
rect -3182 162 -3126 164
rect -3182 110 -3180 162
rect -3180 110 -3128 162
rect -3128 110 -3126 162
rect -3182 108 -3126 110
rect -3047 159 -2991 161
rect -3047 107 -3045 159
rect -3045 107 -2993 159
rect -2993 107 -2991 159
rect -2890 118 -2888 170
rect -2888 118 -2836 170
rect -2836 118 -2834 170
rect -2890 116 -2834 118
rect -673 204 -617 206
rect -673 152 -671 204
rect -671 152 -619 204
rect -619 152 -617 204
rect -224 189 -168 191
rect -673 150 -617 152
rect -486 167 -430 169
rect -3047 105 -2991 107
rect -486 115 -484 167
rect -484 115 -432 167
rect -432 115 -430 167
rect -224 137 -222 189
rect -222 137 -170 189
rect -170 137 -168 189
rect -224 135 -168 137
rect -486 113 -430 115
<< metal3 >>
rect -2907 3673 -2822 3685
rect 1049 3674 1134 3676
rect 1249 3674 1334 3676
rect -2907 3617 -2894 3673
rect -2838 3617 -2822 3673
rect 679 3672 764 3674
rect -2057 3661 -1571 3670
rect -2907 3603 -2822 3617
rect -2058 3655 -1571 3661
rect -2058 3653 -1661 3655
rect -2058 3649 -1850 3653
rect -2058 3593 -2045 3649
rect -1989 3597 -1850 3649
rect -1794 3599 -1661 3653
rect -1605 3599 -1571 3655
rect -1794 3597 -1571 3599
rect -1989 3593 -1571 3597
rect -2058 3574 -1571 3593
rect 673 3662 987 3672
rect 673 3606 692 3662
rect 748 3655 987 3662
rect 748 3606 875 3655
rect 673 3599 875 3606
rect 931 3599 987 3655
rect 673 3582 987 3599
rect 1049 3664 1147 3674
rect 1049 3608 1062 3664
rect 1118 3608 1147 3664
rect 1049 3594 1147 3608
rect 1249 3664 1347 3674
rect 1249 3608 1262 3664
rect 1318 3608 1347 3664
rect 1249 3594 1347 3608
rect -2057 3573 -1571 3574
rect -2363 2662 -2096 2674
rect -3525 2647 -2096 2662
rect -3525 2643 -2187 2647
rect -3525 2587 -2339 2643
rect -2283 2591 -2187 2643
rect -2131 2591 -2096 2647
rect -2283 2587 -2096 2591
rect -3525 2562 -2096 2587
rect -3767 2246 -3603 2261
rect -3767 2190 -3725 2246
rect -3669 2190 -3603 2246
rect -3767 2105 -3603 2190
rect -3525 2105 -3425 2562
rect -2363 2559 -2096 2562
rect -3767 2088 -3425 2105
rect -3767 2032 -3735 2088
rect -3679 2032 -3425 2088
rect -3767 2010 -3425 2032
rect -3659 2005 -3425 2010
rect -2010 1521 -1905 3573
rect -1754 2643 -1389 2656
rect -1754 2631 -1388 2643
rect -1754 2575 -1739 2631
rect -1683 2625 -1460 2631
rect -1683 2575 -1599 2625
rect -1754 2569 -1599 2575
rect -1543 2575 -1460 2625
rect -1404 2575 -1388 2631
rect -1543 2569 -1388 2575
rect -1754 2561 -1388 2569
rect -1754 2549 -1389 2561
rect -1484 1992 -1391 2549
rect 609 2532 702 2538
rect 494 2518 702 2532
rect 494 2462 629 2518
rect 685 2462 702 2518
rect 494 2397 702 2462
rect 494 2341 523 2397
rect 579 2341 702 2397
rect 494 2277 702 2341
rect 494 2221 521 2277
rect 577 2221 702 2277
rect 494 2193 702 2221
rect 609 1992 702 2193
rect -1484 1966 702 1992
rect -1484 1963 -366 1966
rect -1484 1959 -508 1963
rect -1484 1903 -636 1959
rect -580 1907 -508 1959
rect -452 1910 -366 1963
rect -310 1910 702 1966
rect -452 1907 702 1910
rect -580 1903 702 1907
rect -1484 1899 702 1903
rect -2153 1501 -1730 1521
rect -2153 1493 -1820 1501
rect -2153 1437 -2138 1493
rect -2082 1491 -1820 1493
rect -2082 1437 -1978 1491
rect -2153 1435 -1978 1437
rect -1922 1445 -1820 1491
rect -1764 1445 -1730 1501
rect -1922 1435 -1730 1445
rect -2153 1421 -1730 1435
rect -2903 183 -2818 184
rect -3187 178 -2803 183
rect -2010 178 -1905 1421
rect -1484 430 -1391 1899
rect -667 1888 -283 1899
rect 609 432 702 1899
rect 879 1532 984 3582
rect 879 1519 1288 1532
rect 879 1509 1291 1519
rect 879 1504 1206 1509
rect 879 1489 1043 1504
rect 879 1433 919 1489
rect 975 1448 1043 1489
rect 1099 1453 1206 1504
rect 1262 1453 1291 1509
rect 1099 1448 1291 1453
rect 975 1439 1291 1448
rect 975 1433 1288 1439
rect 879 1425 1288 1433
rect 879 1419 991 1425
rect -1581 409 -1170 430
rect -1581 406 -1265 409
rect -1581 350 -1561 406
rect -1505 401 -1265 406
rect -1505 350 -1440 401
rect -1581 345 -1440 350
rect -1384 353 -1265 401
rect -1209 353 -1170 409
rect -1384 345 -1170 353
rect -1581 328 -1170 345
rect 370 408 756 432
rect 370 407 551 408
rect 370 351 404 407
rect 460 352 551 407
rect 607 402 756 408
rect 607 352 679 402
rect 460 351 679 352
rect 370 346 679 351
rect 735 346 756 402
rect 370 325 756 346
rect -686 211 -601 218
rect -686 206 -150 211
rect -686 178 -673 206
rect -3187 176 -673 178
rect -3195 172 -673 176
rect -3195 164 -2890 172
rect -3195 108 -3182 164
rect -3126 161 -2890 164
rect -3126 108 -3047 161
rect -3195 105 -3047 108
rect -2991 116 -2890 161
rect -2834 150 -673 172
rect -617 201 -150 206
rect -617 191 -139 201
rect -617 169 -224 191
rect -617 150 -486 169
rect -2834 116 -486 150
rect -2991 113 -486 116
rect -430 135 -224 169
rect -168 178 -139 191
rect 879 178 984 1419
rect -168 135 984 178
rect -430 113 984 135
rect -2991 105 984 113
rect -3195 94 984 105
rect -3187 74 984 94
rect -2937 73 984 74
use INV_2  INV_2_0
timestamp 1713185578
transform -1 0 -1216 0 -1 3226
box 21 -485 1081 648
use INV_2  INV_2_1
timestamp 1713185578
transform 1 0 -2318 0 1 1930
box 21 -485 1081 648
use INV_2  INV_2_2
timestamp 1713185578
transform 1 0 575 0 -1 3234
box 21 -485 1081 648
use INV_2  INV_2_3
timestamp 1713185578
transform 1 0 575 0 1 1938
box 21 -485 1081 648
use INV_2  INV_2_4
timestamp 1713185578
transform -1 0 1677 0 -1 968
box 21 -485 1081 648
use INV_2  INV_2_5
timestamp 1713185578
transform -1 0 -1216 0 -1 960
box 21 -485 1081 648
use Tr_Gate  Tr_Gate_0
timestamp 1713185578
transform 1 0 -817 0 1 1343
box -53 -1233 1187 569
use Tr_Gate  Tr_Gate_1
timestamp 1713185578
transform 1 0 -817 0 -1 2509
box -53 -1233 1187 569
use Tr_Gate  Tr_Gate_2
timestamp 1713185578
transform -1 0 -2663 0 -1 2470
box -53 -1233 1187 569
use Tr_Gate  Tr_Gate_3
timestamp 1713185578
transform -1 0 -2663 0 1 1322
box -53 -1233 1187 569
<< labels >>
flabel metal1 s -3700 3207 -3699 3208 0 FreeSans 1250 0 0 0 D
port 1 nsew
flabel metal1 s -1178 3898 -1178 3898 0 FreeSans 1250 0 0 0 CLK
port 2 nsew
flabel metal1 s 1813 1916 1813 1916 0 FreeSans 1250 0 0 0 Q
port 3 nsew
flabel metal1 s 1835 3254 1835 3254 0 FreeSans 1250 0 0 0 Q-
port 4 nsew
flabel metal1 s 324 3679 324 3679 0 FreeSans 1250 0 0 0 VSS
port 5 nsew
flabel metal1 s -3762 2064 -3762 2064 0 FreeSans 1250 0 0 0 VDD
port 6 nsew
<< end >>
