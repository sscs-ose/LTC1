magic
tech gf180mcuC
magscale 1 10
timestamp 1692705520
<< error_p >>
rect -140 -23 -129 23
rect 72 -23 83 23
<< pwell >>
rect -166 -101 166 101
<< nmos >>
rect -50 -30 50 30
<< ndiff >>
rect -142 30 -70 36
rect 70 30 142 36
rect -142 23 -50 30
rect -142 -23 -129 23
rect -83 -23 -50 23
rect -142 -30 -50 -23
rect 50 23 142 30
rect 50 -23 83 23
rect 129 -23 142 23
rect 50 -30 142 -23
rect -142 -36 -70 -30
rect 70 -36 142 -30
<< ndiffc >>
rect -129 -23 -83 23
rect 83 -23 129 23
<< polysilicon >>
rect -50 30 50 74
rect -50 -74 50 -30
<< metal1 >>
rect -140 -23 -129 23
rect -83 -23 -72 23
rect 72 -23 83 23
rect 129 -23 140 23
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 0.3 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
