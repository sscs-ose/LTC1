magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2345 -2095 2345 2095
<< psubdiff >>
rect -345 70 345 95
rect -345 -70 -305 70
rect 305 -70 345 70
rect -345 -95 345 -70
<< psubdiffcont >>
rect -305 -70 305 70
<< metal1 >>
rect -334 70 334 84
rect -334 -70 -305 70
rect 305 -70 334 70
rect -334 -84 334 -70
<< end >>
