magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -3173 -2045 3173 2045
<< psubdiff >>
rect -1173 23 1173 45
rect -1173 -23 -1151 23
rect 1151 -23 1173 23
rect -1173 -45 1173 -23
<< psubdiffcont >>
rect -1151 -23 1151 23
<< metal1 >>
rect -1162 23 1162 34
rect -1162 -23 -1151 23
rect 1151 -23 1162 23
rect -1162 -34 1162 -23
<< end >>
