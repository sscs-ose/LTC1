magic
tech gf180mcuC
magscale 1 10
timestamp 1692688043
<< nwell >>
rect 0 321 1924 531
<< psubdiff >>
rect 31 -478 1884 -464
rect 31 -525 44 -478
rect 96 -525 154 -478
rect 206 -525 264 -478
rect 316 -525 374 -478
rect 426 -525 484 -478
rect 536 -525 594 -478
rect 646 -525 704 -478
rect 756 -525 814 -478
rect 866 -525 924 -478
rect 976 -525 1034 -478
rect 1086 -525 1144 -478
rect 1196 -525 1254 -478
rect 1306 -525 1364 -478
rect 1416 -525 1474 -478
rect 1526 -525 1584 -478
rect 1636 -525 1694 -478
rect 1746 -525 1804 -478
rect 1856 -525 1884 -478
rect 31 -538 1884 -525
<< nsubdiff >>
rect 30 481 1887 494
rect 30 430 44 481
rect 95 430 154 481
rect 205 430 264 481
rect 315 430 374 481
rect 425 430 484 481
rect 535 430 594 481
rect 645 430 704 481
rect 755 430 814 481
rect 865 430 924 481
rect 975 430 1034 481
rect 1085 430 1144 481
rect 1195 430 1254 481
rect 1305 430 1364 481
rect 1415 430 1474 481
rect 1525 430 1584 481
rect 1635 430 1694 481
rect 1745 430 1804 481
rect 1855 430 1887 481
rect 30 416 1887 430
<< psubdiffcont >>
rect 44 -525 96 -478
rect 154 -525 206 -478
rect 264 -525 316 -478
rect 374 -525 426 -478
rect 484 -525 536 -478
rect 594 -525 646 -478
rect 704 -525 756 -478
rect 814 -525 866 -478
rect 924 -525 976 -478
rect 1034 -525 1086 -478
rect 1144 -525 1196 -478
rect 1254 -525 1306 -478
rect 1364 -525 1416 -478
rect 1474 -525 1526 -478
rect 1584 -525 1636 -478
rect 1694 -525 1746 -478
rect 1804 -525 1856 -478
<< nsubdiffcont >>
rect 44 430 95 481
rect 154 430 205 481
rect 264 430 315 481
rect 374 430 425 481
rect 484 430 535 481
rect 594 430 645 481
rect 704 430 755 481
rect 814 430 865 481
rect 924 430 975 481
rect 1034 430 1085 481
rect 1144 430 1195 481
rect 1254 430 1305 481
rect 1364 430 1415 481
rect 1474 430 1525 481
rect 1584 430 1635 481
rect 1694 430 1745 481
rect 1804 430 1855 481
<< polysilicon >>
rect -32 338 40 346
rect -32 333 570 338
rect -32 287 -19 333
rect 27 287 570 333
rect -32 282 570 287
rect -32 274 40 282
rect 514 230 570 282
rect 842 303 914 316
rect 842 257 855 303
rect 901 257 914 303
rect 1346 303 1418 316
rect 842 244 914 257
rect 850 230 906 244
rect 1018 230 1242 266
rect 1346 257 1359 303
rect 1405 257 1418 303
rect 1346 244 1418 257
rect 1354 230 1410 244
rect 178 92 234 93
rect 682 92 738 112
rect 1522 92 1578 94
rect 178 78 402 92
rect 120 65 402 78
rect 120 19 133 65
rect 179 55 402 65
rect 514 56 738 92
rect 179 19 234 55
rect 120 6 234 19
rect 178 -69 234 6
rect 178 -105 570 -69
rect 682 -79 738 56
rect 178 -114 234 -105
rect 682 -115 1074 -79
rect 1186 -150 1242 92
rect 1522 62 1746 92
rect 1469 56 1746 62
rect 1469 49 1578 56
rect 1469 3 1482 49
rect 1528 3 1578 49
rect 1469 -10 1578 3
rect 1690 -150 1746 56
rect 1186 -266 1578 -230
rect 1186 -332 1242 -266
rect 1170 -345 1242 -332
rect 1170 -391 1183 -345
rect 1229 -391 1242 -345
rect 1170 -404 1242 -391
<< polycontact >>
rect -19 287 27 333
rect 855 257 901 303
rect 1359 257 1405 303
rect 133 19 179 65
rect 1482 3 1528 49
rect 1183 -391 1229 -345
<< metal1 >>
rect 18 481 1899 506
rect 18 430 44 481
rect 95 430 154 481
rect 205 430 264 481
rect 315 430 374 481
rect 425 430 484 481
rect 535 430 594 481
rect 645 430 704 481
rect 755 430 814 481
rect 865 430 924 481
rect 975 430 1034 481
rect 1085 430 1144 481
rect 1195 430 1254 481
rect 1305 430 1364 481
rect 1415 430 1474 481
rect 1525 430 1584 481
rect 1635 430 1694 481
rect 1745 430 1804 481
rect 1855 430 1899 481
rect 18 404 1899 430
rect -32 333 40 346
rect -111 287 -19 333
rect 27 287 40 333
rect -32 274 40 287
rect 99 184 145 404
rect 435 184 481 404
rect 855 316 901 404
rect 1359 316 1405 404
rect 842 303 914 316
rect 1346 303 1418 316
rect 771 257 855 303
rect 901 257 985 303
rect 771 244 985 257
rect 771 184 817 244
rect 939 184 985 244
rect 1275 257 1359 303
rect 1405 257 1489 303
rect 1275 244 1489 257
rect 1275 184 1321 244
rect 1443 184 1489 244
rect 1779 184 1825 404
rect 267 92 313 138
rect 603 92 649 138
rect 1107 92 1153 138
rect 120 65 192 78
rect -111 19 133 65
rect 179 19 192 65
rect 267 49 1313 92
rect 1611 90 1657 138
rect 1469 49 1539 62
rect 267 46 1482 49
rect 120 6 192 19
rect 395 -56 441 46
rect 1267 3 1482 46
rect 1528 3 1539 49
rect 1611 44 1825 90
rect 1469 -10 1539 3
rect 1779 -43 1825 44
rect 99 -102 481 -56
rect 99 -148 145 -102
rect 435 -148 481 -102
rect 603 -102 985 -56
rect 603 -148 649 -102
rect 939 -148 985 -102
rect 1107 -102 1489 -56
rect 1107 -148 1153 -102
rect 1443 -148 1489 -102
rect 1779 -89 1925 -43
rect 267 -240 313 -194
rect 603 -240 649 -194
rect 267 -286 649 -240
rect 771 -240 817 -194
rect 1107 -240 1153 -194
rect 771 -286 1153 -240
rect 1275 -240 1321 -194
rect 1611 -240 1657 -194
rect 1779 -196 1825 -89
rect 1275 -286 1657 -240
rect -111 -345 1242 -332
rect -111 -378 1183 -345
rect 1170 -391 1183 -378
rect 1229 -391 1242 -345
rect 1170 -404 1242 -391
rect 1611 -450 1657 -286
rect 17 -478 1898 -450
rect 17 -525 44 -478
rect 96 -525 154 -478
rect 206 -525 264 -478
rect 316 -525 374 -478
rect 426 -525 484 -478
rect 536 -525 594 -478
rect 646 -525 704 -478
rect 756 -525 814 -478
rect 866 -525 924 -478
rect 976 -525 1034 -478
rect 1086 -525 1144 -478
rect 1196 -525 1254 -478
rect 1306 -525 1364 -478
rect 1416 -525 1474 -478
rect 1526 -525 1584 -478
rect 1636 -525 1694 -478
rect 1746 -525 1804 -478
rect 1856 -525 1898 -478
rect 17 -552 1898 -525
use nmos_3p3_F9QVWA  nmos_3p3_F9QVWA_0
timestamp 1692519410
transform 1 0 878 0 1 -171
box -312 -99 312 99
use nmos_3p3_F9QVWA  nmos_3p3_F9QVWA_1
timestamp 1692519410
transform 1 0 374 0 1 -171
box -312 -99 312 99
use nmos_3p3_F9QVWA  nmos_3p3_F9QVWA_2
timestamp 1692519410
transform 1 0 1382 0 1 -171
box -312 -99 312 99
use nmos_3p3_H9QVWA  nmos_3p3_H9QVWA_0
timestamp 1692686659
transform 1 0 1718 0 1 -171
box -144 -99 144 99
use pmos_3p3_M8RCNG  pmos_3p3_M8RCNG_0
timestamp 1692567440
transform 1 0 1382 0 1 161
box -206 -161 206 161
use pmos_3p3_M8RCNG  pmos_3p3_M8RCNG_1
timestamp 1692567440
transform 1 0 878 0 1 161
box -206 -161 206 161
use pmos_3p3_MGRCNG  pmos_3p3_MGRCNG_0
timestamp 1692619765
transform 1 0 290 0 1 161
box -290 -161 290 161
use pmos_3p3_MGRCNG  pmos_3p3_MGRCNG_1
timestamp 1692619765
transform 1 0 1634 0 1 161
box -290 -161 290 161
use pmos_3p3_MGRCNG  pmos_3p3_MGRCNG_2
timestamp 1692619765
transform -1 0 626 0 1 161
box -290 -161 290 161
use pmos_3p3_MGRCNG  pmos_3p3_MGRCNG_4
timestamp 1692619765
transform 1 0 1130 0 1 161
box -290 -161 290 161
<< labels >>
flabel metal1 -94 311 -94 311 0 FreeSans 480 0 0 0 B
port 0 nsew
flabel metal1 1841 -70 1841 -70 0 FreeSans 480 0 0 0 OUT
port 6 nsew
flabel nsubdiffcont 951 457 951 457 0 FreeSans 480 0 0 0 VDD
port 7 nsew
flabel metal1 -92 -356 -92 -356 0 FreeSans 480 0 0 0 C
port 4 nsew
flabel psubdiffcont 949 -498 949 -498 0 FreeSans 480 0 0 0 VSS
port 9 nsew
flabel metal1 -91 45 -91 45 0 FreeSans 480 0 0 0 A
port 10 nsew
<< end >>
