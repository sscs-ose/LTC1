* NGSPICE file created from folded_single_check8_flat.ext - technology: gf180mcuC

.subckt folded_single_check8_flat VDD VSS VINP VINN OUT IBIAS
X0 VSS a_n2814_n10181.t20 a_n3063_n8710.t15 VSS.t43 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1 OUT.t25 OUT.t24 OUT.t25 VSS.t10 nfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X2 VSS a_n2814_n10181.t21 a_n3063_n9510.t22 VSS.t18 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X3 a_n453_n1964.t7 a_n453_n1964.t6 a_n453_n1964.t7 VDD.t17 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.56u
X4 VSS a_n89_n10306.t0 a_n89_n10306.t1 VSS.t3 nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.56u
X5 VDD IBIAS.t3 a_n2983_n1659.t30 VDD.t48 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X6 a_n453_n3002.t19 a_n453_n3002.t18 a_n453_n3002.t19 VDD.t17 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.56u
X7 VSS a_n2814_n10181.t22 a_n3063_n9510.t21 VSS.t33 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X8 OUT.t23 OUT.t22 OUT.t23 VSS.t10 nfet_03v3 ad=0 pd=0 as=0.78p ps=3.52u w=3u l=0.28u
X9 VDD IBIAS.t7 a_n453_n3002.t11 VDD.t23 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X10 a_n2983_n1659.t15 a_n2983_n1659.t14 a_n2983_n1659.t15 VDD.t31 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.56u
X11 VDD IBIAS.t8 a_n2983_n1659.t26 VDD.t26 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X12 VDD IBIAS.t9 a_n2983_n1659.t25 VDD.t26 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X13 a_n2983_n1659.t13 a_n2983_n1659.t12 a_n2983_n1659.t13 VDD.t31 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.56u
X14 a_n3063_n8710.t31 a_n3063_n8710.t30 a_n3063_n8710.t31 VSS.t6 nfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X15 a_n2983_n1659.t11 a_n2983_n1659.t10 a_n2983_n1659.t11 VDD.t31 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.56u
X16 a_n453_n3002.t17 a_n453_n3002.t16 a_n453_n3002.t17 VDD.t17 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.56u
X17 OUT a_n168_n4318.t6 a_n453_n1964.t18 VDD.t39 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X18 VDD IBIAS.t10 a_n453_n1964.t17 VDD.t23 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X19 a_n2814_n10181.t17 a_n2814_n10181.t16 a_n2814_n10181.t17 VSS.t0 nfet_03v3 ad=0 pd=0 as=1.32p ps=6.88u w=3u l=0.28u
X20 VDD IBIAS.t11 a_n2983_n1659.t24 VDD.t26 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X21 a_n3063_n8710.t29 a_n3063_n8710.t28 a_n3063_n8710.t29 VSS.t6 nfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X22 OUT.t21 OUT.t20 OUT.t21 VSS.t0 nfet_03v3 ad=0 pd=0 as=1.32p ps=6.88u w=3u l=0.28u
X23 OUT a_n89_n10306.t7 a_n3063_n8710.t1 VSS.t1 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X24 VSS a_n2814_n10181.t29 a_n3063_n8710.t14 VSS.t22 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X25 VSS a_n2814_n10181.t30 a_n3063_n8710.t13 VSS.t22 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X26 a_n3063_n9510.t31 a_n3063_n9510.t30 a_n3063_n9510.t31 VSS.t9 nfet_03v3 ad=0 pd=0 as=1.32p ps=6.88u w=3u l=0.28u
X27 a_n453_n1964.t5 a_n453_n1964.t4 a_n453_n1964.t5 VDD.t17 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.56u
X28 VSS a_n2814_n10181.t32 a_n3063_n8710.t12 VSS.t18 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X29 OUT a_n168_n4318.t8 a_n453_n1964.t19 VDD.t39 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X30 VSS a_n2814_n10181.t33 a_n3063_n8710.t11 VSS.t43 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X31 a_n3063_n9510.t29 a_n3063_n9510.t28 a_n3063_n9510.t29 VSS.t9 nfet_03v3 ad=0 pd=0 as=1.32p ps=6.88u w=3u l=0.28u
X32 VDD IBIAS.t17 a_n453_n1964.t14 VDD.t33 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X33 VSS a_n2814_n10181.t34 a_n3063_n9510.t16 VSS.t43 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X34 VSS a_n2814_n10181.t36 a_n3063_n8710.t10 VSS.t18 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X35 a_n2814_n10181.t15 a_n2814_n10181.t14 a_n2814_n10181.t15 VSS.t10 nfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X36 OUT a_n89_n10306.t11 a_n3063_n8710.t5 VSS.t8 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X37 VSS a_n2814_n10181.t37 a_n3063_n9510.t15 VSS.t43 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X38 a_n2983_n1659.t9 a_n2983_n1659.t8 a_n2983_n1659.t9 VDD.t31 pfet_03v3 ad=0 pd=0 as=0.78p ps=3.52u w=3u l=0.56u
X39 OUT.t19 OUT.t18 OUT.t19 VDD.t8 pfet_03v3 ad=0 pd=0 as=1.32p ps=6.88u w=3u l=0.28u
X40 VSS a_n2814_n10181.t38 a_n3063_n8710.t9 VSS.t33 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X41 VDD IBIAS.t24 a_n453_n1964.t12 VDD.t33 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X42 a_n2983_n1659.t7 a_n2983_n1659.t6 a_n2983_n1659.t7 VDD.t64 pfet_03v3 ad=0 pd=0 as=1.32p ps=6.88u w=3u l=0.56u
X43 VSS a_n2814_n10181.t39 a_n3063_n9510.t14 VSS.t33 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X44 VDD IBIAS.t26 a_n453_n3002.t7 VDD.t33 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X45 a_n453_n1964.t3 a_n453_n1964.t2 a_n453_n1964.t3 VDD.t30 pfet_03v3 ad=0 pd=0 as=1.32p ps=6.88u w=3u l=0.56u
X46 VSS a_3734_n7493.t3 a_n168_n4318.t2 VSS.t3 nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.56u
X47 OUT a_n89_n10306.t12 a_n3063_n8710.t4 VSS.t8 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X48 VSS a_n2814_n10181.t43 a_n3063_n8710.t8 VSS.t33 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X49 a_n453_n3002.t15 a_n453_n3002.t14 a_n453_n3002.t15 VDD.t30 pfet_03v3 ad=0 pd=0 as=1.32p ps=6.88u w=3u l=0.56u
X50 a_n3063_n9510.t27 a_n3063_n9510.t26 a_n3063_n9510.t27 VSS.t6 nfet_03v3 ad=0 pd=0 as=0.78p ps=3.52u w=3u l=0.28u
X51 VDD IBIAS.t28 a_n2983_n1659.t19 VDD.t48 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X52 VDD IBIAS.t29 a_n453_n1964.t10 VDD.t23 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X53 a_n2814_n10181.t13 a_n2814_n10181.t12 a_n2814_n10181.t13 VSS.t0 nfet_03v3 ad=0 pd=0 as=1.32p ps=6.88u w=3u l=0.28u
X54 a_n2983_n1659.t5 a_n2983_n1659.t4 a_n2983_n1659.t5 VDD.t64 pfet_03v3 ad=0 pd=0 as=1.32p ps=6.88u w=3u l=0.56u
X55 VDD IBIAS.t30 a_n453_n3002.t5 VDD.t23 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X56 a_n3063_n9510.t25 a_n3063_n9510.t24 a_n3063_n9510.t25 VSS.t6 nfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X57 OUT.t17 OUT.t16 OUT.t17 VDD.t8 pfet_03v3 ad=0 pd=0 as=1.32p ps=6.88u w=3u l=0.28u
X58 OUT.t15 OUT.t14 OUT.t15 VDD.t3 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X59 a_n2983_n1659.t3 a_n2983_n1659.t2 a_n2983_n1659.t3 VDD.t64 pfet_03v3 ad=0 pd=0 as=1.32p ps=6.88u w=3u l=0.56u
X60 VDD IBIAS.t31 a_n453_n3002.t4 VDD.t33 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X61 OUT a_n89_n10306.t14 a_n3063_n8710.t7 VSS.t1 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X62 VDD IBIAS.t32 a_n2983_n1659.t18 VDD.t26 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X63 VDD IBIAS.t33 a_n2983_n1659.t17 VDD.t48 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X64 VDD IBIAS.t34 a_n2983_n1659.t16 VDD.t48 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X65 a_n453_n1964.t1 a_n453_n1964.t0 a_n453_n1964.t1 VDD.t30 pfet_03v3 ad=0 pd=0 as=1.32p ps=6.88u w=3u l=0.56u
X66 VSS a_n2814_n10181.t47 a_n3063_n9510.t11 VSS.t22 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X67 a_n3063_n8710.t27 a_n3063_n8710.t26 a_n3063_n8710.t27 VSS.t9 nfet_03v3 ad=0 pd=0 as=1.32p ps=6.88u w=3u l=0.28u
X68 OUT.t13 OUT.t12 OUT.t13 VDD.t3 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X69 a_n2983_n1659.t1 a_n2983_n1659.t0 a_n2983_n1659.t1 VDD.t64 pfet_03v3 ad=0 pd=0 as=1.32p ps=6.88u w=3u l=0.56u
X70 VDD IBIAS.t0 IBIAS.t1 VDD.t65 pfet_03v3 ad=1.76p pd=8.88u as=1.76p ps=8.88u w=4u l=0.56u
X71 OUT.t11 OUT.t10 OUT.t11 VSS.t0 nfet_03v3 ad=0 pd=0 as=1.32p ps=6.88u w=3u l=0.28u
X72 a_n453_n3002.t13 a_n453_n3002.t12 a_n453_n3002.t13 VDD.t30 pfet_03v3 ad=0 pd=0 as=1.32p ps=6.88u w=3u l=0.56u
X73 VSS a_3734_n7493.t1 a_3734_n7493.t2 VSS.t11 nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.56u
X74 VSS a_n2814_n10181.t49 a_n3063_n9510.t9 VSS.t22 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X75 VSS a_n2814_n10181.t50 a_n3063_n9510.t8 VSS.t18 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X76 a_n2814_n10181.t11 a_n2814_n10181.t10 a_n2814_n10181.t11 VSS.t10 nfet_03v3 ad=0 pd=0 as=0.78p ps=3.52u w=3u l=0.28u
X77 a_n3063_n8710.t25 a_n3063_n8710.t24 a_n3063_n8710.t25 VSS.t9 nfet_03v3 ad=0 pd=0 as=1.32p ps=6.88u w=3u l=0.28u
R0 a_n2777_n5169.n0 a_n2777_n5169.t1 1.21383
R1 a_n2617_n5169.t0 a_n2617_n5169.n0 1.21383
R2 VDD.t62 VDD.t83 409.736
R3 VDD.t79 VDD.t65 363.524
R4 VDD.n195 VDD.t62 255.7
R5 VDD.n195 VDD.t79 153.421
R6 VDD.n254 VDD.t3 19.3637
R7 VDD.n1068 VDD.t26 12.698
R8 VDD.n266 VDD.t22 11.6184
R9 VDD.n622 VDD.t9 11.4588
R10 VDD.n1049 VDD.t64 11.005
R11 VDD.n640 VDD.t14 10.4172
R12 VDD.n287 VDD.t8 9.89723
R13 VDD.n902 VDD.t23 9.61159
R14 VDD.n864 VDD.t17 9.16456
R15 VDD.n257 VDD.t39 9.03664
R16 VDD.n607 VDD.t11 8.85467
R17 VDD.n604 VDD.t10 8.33383
R18 VDD.n873 VDD.t4 7.15294
R19 VDD.n643 VDD.t1 6.77133
R20 VDD.n911 VDD.t30 6.70591
R21 VDD.n194 VDD.t84 6.50617
R22 VDD.n196 VDD.n195 6.3005
R23 VDD.n1078 VDD.t20 5.92601
R24 VDD.n619 VDD.t12 5.72967
R25 VDD.n1062 VDD.t18 4.79734
R26 VDD.n194 VDD.t63 4.41333
R27 VDD.n198 VDD.n193 4.41137
R28 VDD.n197 VDD.t80 4.41137
R29 VDD.n628 VDD.t16 4.16717
R30 VDD.n707 VDD.n706 3.54072
R31 VDD.n707 VDD.n705 3.54072
R32 VDD.n201 VDD.n200 3.48503
R33 VDD.n201 VDD.n199 3.48503
R34 VDD.n383 VDD.n381 3.48503
R35 VDD.n359 VDD.n357 3.48503
R36 VDD.n359 VDD.n358 3.48503
R37 VDD.n886 VDD.t6 3.3532
R38 VDD.n835 VDD.n834 3.1505
R39 VDD.n14 VDD.n13 3.1505
R40 VDD.n12 VDD.n11 3.1505
R41 VDD.n10 VDD.n9 3.1505
R42 VDD.n8 VDD.n7 3.1505
R43 VDD.n752 VDD.n751 3.1505
R44 VDD.n754 VDD.n753 3.1505
R45 VDD.n756 VDD.n755 3.1505
R46 VDD.n758 VDD.n757 3.1505
R47 VDD.n760 VDD.n759 3.1505
R48 VDD.n762 VDD.n761 3.1505
R49 VDD.n764 VDD.n763 3.1505
R50 VDD.n766 VDD.n765 3.1505
R51 VDD.n768 VDD.n767 3.1505
R52 VDD.n770 VDD.n769 3.1505
R53 VDD.n772 VDD.n771 3.1505
R54 VDD.n774 VDD.n773 3.1505
R55 VDD.n776 VDD.n775 3.1505
R56 VDD.n778 VDD.n777 3.1505
R57 VDD.n780 VDD.n779 3.1505
R58 VDD.n782 VDD.n781 3.1505
R59 VDD.n784 VDD.n783 3.1505
R60 VDD.n786 VDD.n785 3.1505
R61 VDD.n788 VDD.n787 3.1505
R62 VDD.n790 VDD.n789 3.1505
R63 VDD.n792 VDD.n791 3.1505
R64 VDD.n794 VDD.n793 3.1505
R65 VDD.n796 VDD.n795 3.1505
R66 VDD.n798 VDD.n797 3.1505
R67 VDD.n800 VDD.n799 3.1505
R68 VDD.n803 VDD.n802 3.1505
R69 VDD.n805 VDD.n804 3.1505
R70 VDD.n808 VDD.n807 3.1505
R71 VDD.n810 VDD.n809 3.1505
R72 VDD.n813 VDD.n812 3.1505
R73 VDD.n815 VDD.n814 3.1505
R74 VDD.n818 VDD.n817 3.1505
R75 VDD.n820 VDD.n819 3.1505
R76 VDD.n823 VDD.n822 3.1505
R77 VDD.n825 VDD.n824 3.1505
R78 VDD.n828 VDD.n827 3.1505
R79 VDD.n830 VDD.n829 3.1505
R80 VDD.n833 VDD.n832 3.1505
R81 VDD.n16 VDD.n15 3.1505
R82 VDD.n854 VDD.n853 3.1505
R83 VDD.n857 VDD.n856 3.1505
R84 VDD.n856 VDD.n855 3.1505
R85 VDD.n860 VDD.n859 3.1505
R86 VDD.n859 VDD.n858 3.1505
R87 VDD.n863 VDD.n862 3.1505
R88 VDD.n862 VDD.n861 3.1505
R89 VDD.n866 VDD.n865 3.1505
R90 VDD.n865 VDD.n864 3.1505
R91 VDD.n869 VDD.n868 3.1505
R92 VDD.n868 VDD.n867 3.1505
R93 VDD.n872 VDD.n871 3.1505
R94 VDD.n871 VDD.n870 3.1505
R95 VDD.n875 VDD.n874 3.1505
R96 VDD.n874 VDD.n873 3.1505
R97 VDD.n879 VDD.n878 3.1505
R98 VDD.n878 VDD.n877 3.1505
R99 VDD.n882 VDD.n881 3.1505
R100 VDD.n881 VDD.n880 3.1505
R101 VDD.n885 VDD.n884 3.1505
R102 VDD.n884 VDD.n883 3.1505
R103 VDD.n888 VDD.n887 3.1505
R104 VDD.n887 VDD.n886 3.1505
R105 VDD.n891 VDD.n890 3.1505
R106 VDD.n890 VDD.n889 3.1505
R107 VDD.n904 VDD.n903 3.1505
R108 VDD.n903 VDD.n902 3.1505
R109 VDD.n907 VDD.n906 3.1505
R110 VDD.n906 VDD.n905 3.1505
R111 VDD.n910 VDD.n909 3.1505
R112 VDD.n909 VDD.n908 3.1505
R113 VDD.n913 VDD.n912 3.1505
R114 VDD.n912 VDD.n911 3.1505
R115 VDD.n916 VDD.n915 3.1505
R116 VDD.n915 VDD.n914 3.1505
R117 VDD.n919 VDD.n918 3.1505
R118 VDD.n918 VDD.n917 3.1505
R119 VDD.n922 VDD.n921 3.1505
R120 VDD.n921 VDD.n920 3.1505
R121 VDD.n924 VDD.n923 3.1505
R122 VDD.n58 VDD.n57 3.1505
R123 VDD.n20 VDD.n19 3.1505
R124 VDD.n22 VDD.n21 3.1505
R125 VDD.n24 VDD.n23 3.1505
R126 VDD.n26 VDD.n25 3.1505
R127 VDD.n28 VDD.n27 3.1505
R128 VDD.n30 VDD.n29 3.1505
R129 VDD.n32 VDD.n31 3.1505
R130 VDD.n35 VDD.n34 3.1505
R131 VDD.n37 VDD.n36 3.1505
R132 VDD.n39 VDD.n38 3.1505
R133 VDD.n41 VDD.n40 3.1505
R134 VDD.n43 VDD.n42 3.1505
R135 VDD.n46 VDD.n45 3.1505
R136 VDD.n48 VDD.n47 3.1505
R137 VDD.n50 VDD.n49 3.1505
R138 VDD.n52 VDD.n51 3.1505
R139 VDD.n54 VDD.n53 3.1505
R140 VDD.n56 VDD.n55 3.1505
R141 VDD.n18 VDD.n17 3.1505
R142 VDD.n741 VDD.n740 3.1505
R143 VDD.n724 VDD.n723 3.1505
R144 VDD.n724 VDD.n722 3.1505
R145 VDD.n693 VDD.n692 3.1505
R146 VDD.n681 VDD.n425 3.1505
R147 VDD.n410 VDD.n409 3.1505
R148 VDD.n412 VDD.n411 3.1505
R149 VDD.n414 VDD.n413 3.1505
R150 VDD.n416 VDD.n415 3.1505
R151 VDD.n418 VDD.n417 3.1505
R152 VDD.n420 VDD.n419 3.1505
R153 VDD.n422 VDD.n421 3.1505
R154 VDD.n424 VDD.n423 3.1505
R155 VDD.n683 VDD.n682 3.1505
R156 VDD.n685 VDD.n684 3.1505
R157 VDD.n687 VDD.n686 3.1505
R158 VDD.n689 VDD.n688 3.1505
R159 VDD.n691 VDD.n690 3.1505
R160 VDD.n695 VDD.n694 3.1505
R161 VDD.n697 VDD.n696 3.1505
R162 VDD.n699 VDD.n698 3.1505
R163 VDD.n702 VDD.n701 3.1505
R164 VDD.n704 VDD.n703 3.1505
R165 VDD.n710 VDD.n709 3.1505
R166 VDD.n712 VDD.n711 3.1505
R167 VDD.n715 VDD.n714 3.1505
R168 VDD.n717 VDD.n716 3.1505
R169 VDD.n720 VDD.n719 3.1505
R170 VDD.n726 VDD.n725 3.1505
R171 VDD.n729 VDD.n728 3.1505
R172 VDD.n731 VDD.n730 3.1505
R173 VDD.n734 VDD.n733 3.1505
R174 VDD.n736 VDD.n735 3.1505
R175 VDD.n739 VDD.n738 3.1505
R176 VDD.n940 VDD.n939 3.1505
R177 VDD.n408 VDD.n0 3.1505
R178 VDD.n60 VDD.n59 3.1505
R179 VDD.n399 VDD.n398 3.1505
R180 VDD.n401 VDD.n400 3.1505
R181 VDD.n403 VDD.n402 3.1505
R182 VDD.n405 VDD.n404 3.1505
R183 VDD.n407 VDD.n406 3.1505
R184 VDD.n244 VDD.n243 3.1505
R185 VDD.n250 VDD.n249 3.1505
R186 VDD.n249 VDD.n248 3.1505
R187 VDD.n253 VDD.n252 3.1505
R188 VDD.n252 VDD.n251 3.1505
R189 VDD.n256 VDD.n255 3.1505
R190 VDD.n255 VDD.n254 3.1505
R191 VDD.n259 VDD.n258 3.1505
R192 VDD.n258 VDD.n257 3.1505
R193 VDD.n262 VDD.n261 3.1505
R194 VDD.n261 VDD.n260 3.1505
R195 VDD.n265 VDD.n264 3.1505
R196 VDD.n264 VDD.n263 3.1505
R197 VDD.n268 VDD.n267 3.1505
R198 VDD.n267 VDD.n266 3.1505
R199 VDD.n271 VDD.n270 3.1505
R200 VDD.n270 VDD.n269 3.1505
R201 VDD.n274 VDD.n273 3.1505
R202 VDD.n273 VDD.n272 3.1505
R203 VDD.n277 VDD.n276 3.1505
R204 VDD.n276 VDD.n275 3.1505
R205 VDD.n280 VDD.n279 3.1505
R206 VDD.n279 VDD.n278 3.1505
R207 VDD.n283 VDD.n282 3.1505
R208 VDD.n282 VDD.n281 3.1505
R209 VDD.n286 VDD.n285 3.1505
R210 VDD.n285 VDD.n284 3.1505
R211 VDD.n289 VDD.n288 3.1505
R212 VDD.n288 VDD.n287 3.1505
R213 VDD.n292 VDD.n291 3.1505
R214 VDD.n291 VDD.n290 3.1505
R215 VDD.n295 VDD.n294 3.1505
R216 VDD.n294 VDD.n293 3.1505
R217 VDD.n297 VDD.n296 3.1505
R218 VDD.n247 VDD.n246 3.1505
R219 VDD.n246 VDD.n245 3.1505
R220 VDD.n242 VDD.n241 3.1505
R221 VDD.n236 VDD.n235 3.1505
R222 VDD.n234 VDD.n233 3.1505
R223 VDD.n231 VDD.n230 3.1505
R224 VDD.n229 VDD.n228 3.1505
R225 VDD.n226 VDD.n225 3.1505
R226 VDD.n224 VDD.n223 3.1505
R227 VDD.n221 VDD.n220 3.1505
R228 VDD.n219 VDD.n218 3.1505
R229 VDD.n216 VDD.n215 3.1505
R230 VDD.n214 VDD.n213 3.1505
R231 VDD.n211 VDD.n210 3.1505
R232 VDD.n209 VDD.n208 3.1505
R233 VDD.n206 VDD.n205 3.1505
R234 VDD.n204 VDD.n203 3.1505
R235 VDD.n192 VDD.n191 3.1505
R236 VDD.n190 VDD.n189 3.1505
R237 VDD.n188 VDD.n187 3.1505
R238 VDD.n302 VDD.n301 3.1505
R239 VDD.n305 VDD.n304 3.1505
R240 VDD.n343 VDD.n342 3.1505
R241 VDD.n307 VDD.n306 3.1505
R242 VDD.n309 VDD.n308 3.1505
R243 VDD.n311 VDD.n310 3.1505
R244 VDD.n313 VDD.n312 3.1505
R245 VDD.n315 VDD.n314 3.1505
R246 VDD.n317 VDD.n316 3.1505
R247 VDD.n319 VDD.n318 3.1505
R248 VDD.n321 VDD.n320 3.1505
R249 VDD.n323 VDD.n322 3.1505
R250 VDD.n325 VDD.n324 3.1505
R251 VDD.n327 VDD.n326 3.1505
R252 VDD.n329 VDD.n328 3.1505
R253 VDD.n331 VDD.n330 3.1505
R254 VDD.n333 VDD.n332 3.1505
R255 VDD.n335 VDD.n334 3.1505
R256 VDD.n337 VDD.n336 3.1505
R257 VDD.n339 VDD.n338 3.1505
R258 VDD.n341 VDD.n340 3.1505
R259 VDD.n393 VDD.n392 3.1505
R260 VDD.n391 VDD.n390 3.1505
R261 VDD.n388 VDD.n387 3.1505
R262 VDD.n386 VDD.n385 3.1505
R263 VDD.n377 VDD.n376 3.1505
R264 VDD.n374 VDD.n373 3.1505
R265 VDD.n372 VDD.n371 3.1505
R266 VDD.n369 VDD.n368 3.1505
R267 VDD.n367 VDD.n366 3.1505
R268 VDD.n364 VDD.n363 3.1505
R269 VDD.n362 VDD.n361 3.1505
R270 VDD.n356 VDD.n355 3.1505
R271 VDD.n354 VDD.n353 3.1505
R272 VDD.n352 VDD.n351 3.1505
R273 VDD.n350 VDD.n349 3.1505
R274 VDD.n346 VDD.n345 3.1505
R275 VDD.n300 VDD.n299 3.1505
R276 VDD.n348 VDD.n347 3.1505
R277 VDD.n90 VDD.n89 3.1505
R278 VDD.n590 VDD.n589 3.1505
R279 VDD.n588 VDD.n587 3.1505
R280 VDD.n585 VDD.n584 3.1505
R281 VDD.n583 VDD.n582 3.1505
R282 VDD.n580 VDD.n579 3.1505
R283 VDD.n578 VDD.n577 3.1505
R284 VDD.n575 VDD.n574 3.1505
R285 VDD.n573 VDD.n572 3.1505
R286 VDD.n570 VDD.n569 3.1505
R287 VDD.n568 VDD.n567 3.1505
R288 VDD.n565 VDD.n564 3.1505
R289 VDD.n563 VDD.n562 3.1505
R290 VDD.n560 VDD.n559 3.1505
R291 VDD.n558 VDD.n557 3.1505
R292 VDD.n555 VDD.n554 3.1505
R293 VDD.n553 VDD.n552 3.1505
R294 VDD.n551 VDD.n550 3.1505
R295 VDD.n549 VDD.n548 3.1505
R296 VDD.n547 VDD.n546 3.1505
R297 VDD.n545 VDD.n544 3.1505
R298 VDD.n543 VDD.n542 3.1505
R299 VDD.n541 VDD.n540 3.1505
R300 VDD.n539 VDD.n538 3.1505
R301 VDD.n537 VDD.n536 3.1505
R302 VDD.n535 VDD.n534 3.1505
R303 VDD.n533 VDD.n532 3.1505
R304 VDD.n531 VDD.n530 3.1505
R305 VDD.n529 VDD.n528 3.1505
R306 VDD.n527 VDD.n526 3.1505
R307 VDD.n525 VDD.n524 3.1505
R308 VDD.n523 VDD.n522 3.1505
R309 VDD.n521 VDD.n520 3.1505
R310 VDD.n519 VDD.n518 3.1505
R311 VDD.n517 VDD.n516 3.1505
R312 VDD.n515 VDD.n514 3.1505
R313 VDD.n513 VDD.n512 3.1505
R314 VDD.n511 VDD.n510 3.1505
R315 VDD.n132 VDD.n131 3.1505
R316 VDD.n130 VDD.n129 3.1505
R317 VDD.n128 VDD.n127 3.1505
R318 VDD.n126 VDD.n125 3.1505
R319 VDD.n124 VDD.n123 3.1505
R320 VDD.n122 VDD.n121 3.1505
R321 VDD.n120 VDD.n119 3.1505
R322 VDD.n118 VDD.n117 3.1505
R323 VDD.n116 VDD.n115 3.1505
R324 VDD.n114 VDD.n113 3.1505
R325 VDD.n112 VDD.n111 3.1505
R326 VDD.n110 VDD.n109 3.1505
R327 VDD.n108 VDD.n107 3.1505
R328 VDD.n106 VDD.n105 3.1505
R329 VDD.n104 VDD.n103 3.1505
R330 VDD.n102 VDD.n101 3.1505
R331 VDD.n100 VDD.n99 3.1505
R332 VDD.n98 VDD.n97 3.1505
R333 VDD.n96 VDD.n95 3.1505
R334 VDD.n94 VDD.n93 3.1505
R335 VDD.n92 VDD.n91 3.1505
R336 VDD.n134 VDD.n133 3.1505
R337 VDD.n668 VDD.n667 3.1505
R338 VDD.n655 VDD.n654 3.1505
R339 VDD.n650 VDD.n649 3.1505
R340 VDD.n653 VDD.n652 3.1505
R341 VDD.n648 VDD.n647 3.1505
R342 VDD.n62 VDD.n61 3.1505
R343 VDD.n82 VDD.n81 3.1505
R344 VDD.n64 VDD.n63 3.1505
R345 VDD.n67 VDD.n66 3.1505
R346 VDD.n69 VDD.n68 3.1505
R347 VDD.n72 VDD.n71 3.1505
R348 VDD.n74 VDD.n73 3.1505
R349 VDD.n77 VDD.n76 3.1505
R350 VDD.n79 VDD.n78 3.1505
R351 VDD.n85 VDD.n84 3.1505
R352 VDD.n88 VDD.n87 3.1505
R353 VDD.n185 VDD.n184 3.1505
R354 VDD.n177 VDD.n176 3.1505
R355 VDD.n180 VDD.n179 3.1505
R356 VDD.n182 VDD.n181 3.1505
R357 VDD.n175 VDD.n174 3.1505
R358 VDD.n172 VDD.n171 3.1505
R359 VDD.n156 VDD.n155 3.1505
R360 VDD.n158 VDD.n157 3.1505
R361 VDD.n160 VDD.n159 3.1505
R362 VDD.n162 VDD.n161 3.1505
R363 VDD.n164 VDD.n163 3.1505
R364 VDD.n166 VDD.n165 3.1505
R365 VDD.n169 VDD.n168 3.1505
R366 VDD.n154 VDD.n153 3.1505
R367 VDD.n152 VDD.n151 3.1505
R368 VDD.n145 VDD.n144 3.1505
R369 VDD.n147 VDD.n146 3.1505
R370 VDD.n149 VDD.n148 3.1505
R371 VDD.n143 VDD.n142 3.1505
R372 VDD.n141 VDD.n140 3.1505
R373 VDD.n138 VDD.n137 3.1505
R374 VDD.n136 VDD.n135 3.1505
R375 VDD.n591 VDD.n509 3.1505
R376 VDD.n645 VDD.n644 3.1505
R377 VDD.n644 VDD.n643 3.1505
R378 VDD.n642 VDD.n641 3.1505
R379 VDD.n641 VDD.n640 3.1505
R380 VDD.n639 VDD.n638 3.1505
R381 VDD.n638 VDD.n637 3.1505
R382 VDD.n636 VDD.n635 3.1505
R383 VDD.n635 VDD.n634 3.1505
R384 VDD.n633 VDD.n632 3.1505
R385 VDD.n632 VDD.n631 3.1505
R386 VDD.n630 VDD.n629 3.1505
R387 VDD.n629 VDD.n628 3.1505
R388 VDD.n627 VDD.n626 3.1505
R389 VDD.n626 VDD.n625 3.1505
R390 VDD.n624 VDD.n623 3.1505
R391 VDD.n623 VDD.n622 3.1505
R392 VDD.n621 VDD.n620 3.1505
R393 VDD.n620 VDD.n619 3.1505
R394 VDD.n618 VDD.n617 3.1505
R395 VDD.n617 VDD.n616 3.1505
R396 VDD.n615 VDD.n614 3.1505
R397 VDD.n614 VDD.n613 3.1505
R398 VDD.n612 VDD.n611 3.1505
R399 VDD.n611 VDD.n610 3.1505
R400 VDD.n609 VDD.n608 3.1505
R401 VDD.n608 VDD.n607 3.1505
R402 VDD.n606 VDD.n605 3.1505
R403 VDD.n605 VDD.n604 3.1505
R404 VDD.n603 VDD.n602 3.1505
R405 VDD.n602 VDD.n601 3.1505
R406 VDD.n600 VDD.n599 3.1505
R407 VDD.n599 VDD.n598 3.1505
R408 VDD.n597 VDD.n596 3.1505
R409 VDD.n596 VDD.n595 3.1505
R410 VDD.n594 VDD.n593 3.1505
R411 VDD.n593 VDD.n592 3.1505
R412 VDD.n670 VDD.n669 3.1505
R413 VDD.n673 VDD.n672 3.1505
R414 VDD.n672 VDD.n671 3.1505
R415 VDD.n676 VDD.n675 3.1505
R416 VDD.n675 VDD.n674 3.1505
R417 VDD.n448 VDD.n447 3.1505
R418 VDD.n1021 VDD.n1020 3.1505
R419 VDD.n1018 VDD.n1017 3.1505
R420 VDD.n1015 VDD.n1014 3.1505
R421 VDD.n1013 VDD.n1012 3.1505
R422 VDD.n1010 VDD.n1009 3.1505
R423 VDD.n1008 VDD.n1007 3.1505
R424 VDD.n1005 VDD.n1004 3.1505
R425 VDD.n1003 VDD.n1002 3.1505
R426 VDD.n1000 VDD.n999 3.1505
R427 VDD.n998 VDD.n997 3.1505
R428 VDD.n995 VDD.n994 3.1505
R429 VDD.n993 VDD.n992 3.1505
R430 VDD.n990 VDD.n989 3.1505
R431 VDD.n988 VDD.n987 3.1505
R432 VDD.n985 VDD.n984 3.1505
R433 VDD.n983 VDD.n982 3.1505
R434 VDD.n981 VDD.n980 3.1505
R435 VDD.n979 VDD.n978 3.1505
R436 VDD.n977 VDD.n976 3.1505
R437 VDD.n975 VDD.n974 3.1505
R438 VDD.n973 VDD.n972 3.1505
R439 VDD.n971 VDD.n970 3.1505
R440 VDD.n969 VDD.n968 3.1505
R441 VDD.n967 VDD.n966 3.1505
R442 VDD.n965 VDD.n964 3.1505
R443 VDD.n963 VDD.n962 3.1505
R444 VDD.n432 VDD.n431 3.1505
R445 VDD.n434 VDD.n433 3.1505
R446 VDD.n436 VDD.n435 3.1505
R447 VDD.n438 VDD.n437 3.1505
R448 VDD.n440 VDD.n439 3.1505
R449 VDD.n443 VDD.n442 3.1505
R450 VDD.n445 VDD.n444 3.1505
R451 VDD.n1023 VDD.n1022 3.1505
R452 VDD.n491 VDD.n490 3.1505
R453 VDD.n489 VDD.n488 3.1505
R454 VDD.n487 VDD.n486 3.1505
R455 VDD.n485 VDD.n484 3.1505
R456 VDD.n483 VDD.n482 3.1505
R457 VDD.n481 VDD.n480 3.1505
R458 VDD.n475 VDD.n474 3.1505
R459 VDD.n473 VDD.n472 3.1505
R460 VDD.n471 VDD.n470 3.1505
R461 VDD.n469 VDD.n468 3.1505
R462 VDD.n466 VDD.n465 3.1505
R463 VDD.n464 VDD.n463 3.1505
R464 VDD.n462 VDD.n461 3.1505
R465 VDD.n460 VDD.n459 3.1505
R466 VDD.n458 VDD.n457 3.1505
R467 VDD.n456 VDD.n455 3.1505
R468 VDD.n454 VDD.n453 3.1505
R469 VDD.n452 VDD.n451 3.1505
R470 VDD.n450 VDD.n449 3.1505
R471 VDD.n1094 VDD.n1093 3.1505
R472 VDD.n1039 VDD.n1038 3.1505
R473 VDD.n1038 VDD.n1037 3.1505
R474 VDD.n1042 VDD.n1041 3.1505
R475 VDD.n1041 VDD.n1040 3.1505
R476 VDD.n1045 VDD.n1044 3.1505
R477 VDD.n1044 VDD.n1043 3.1505
R478 VDD.n1048 VDD.n1047 3.1505
R479 VDD.n1047 VDD.n1046 3.1505
R480 VDD.n1051 VDD.n1050 3.1505
R481 VDD.n1050 VDD.n1049 3.1505
R482 VDD.n1054 VDD.n1053 3.1505
R483 VDD.n1053 VDD.n1052 3.1505
R484 VDD.n1057 VDD.n1056 3.1505
R485 VDD.n1056 VDD.n1055 3.1505
R486 VDD.n1060 VDD.n1059 3.1505
R487 VDD.n1059 VDD.n1058 3.1505
R488 VDD.n1064 VDD.n1063 3.1505
R489 VDD.n1063 VDD.n1062 3.1505
R490 VDD.n1067 VDD.n1066 3.1505
R491 VDD.n1066 VDD.n1065 3.1505
R492 VDD.n1070 VDD.n1069 3.1505
R493 VDD.n1069 VDD.n1068 3.1505
R494 VDD.n1073 VDD.n1072 3.1505
R495 VDD.n1072 VDD.n1071 3.1505
R496 VDD.n1077 VDD.n1076 3.1505
R497 VDD.n1076 VDD.n1075 3.1505
R498 VDD.n1080 VDD.n1079 3.1505
R499 VDD.n1079 VDD.n1078 3.1505
R500 VDD.n1083 VDD.n1082 3.1505
R501 VDD.n1082 VDD.n1081 3.1505
R502 VDD.n1086 VDD.n1085 3.1505
R503 VDD.n1085 VDD.n1084 3.1505
R504 VDD.n1089 VDD.n1088 3.1505
R505 VDD.n1088 VDD.n1087 3.1505
R506 VDD.n1092 VDD.n1091 3.1505
R507 VDD.n1091 VDD.n1090 3.1505
R508 VDD.n1095 VDD.n1094 3.1505
R509 VDD.n1098 VDD.n1097 3.1505
R510 VDD.n1097 VDD.n1096 3.1505
R511 VDD.n1100 VDD.n1099 3.1505
R512 VDD.n1036 VDD.n1035 3.1505
R513 VDD.n427 VDD.n426 3.1505
R514 VDD.n1126 VDD.n1125 3.1505
R515 VDD.n1123 VDD.n1122 3.1505
R516 VDD.n1121 VDD.n1120 3.1505
R517 VDD.n1119 VDD.n1118 3.1505
R518 VDD.n1128 VDD.n1127 3.1505
R519 VDD.n1131 VDD.n1130 3.1505
R520 VDD.n1135 VDD.n1134 3.1505
R521 VDD.n1146 VDD.n1145 3.1505
R522 VDD.n1143 VDD.n1142 3.1505
R523 VDD.n1140 VDD.n1139 3.1505
R524 VDD.n1138 VDD.n1137 3.1505
R525 VDD.n1148 VDD.n1147 3.1505
R526 VDD.n1152 VDD.n1151 3.1505
R527 VDD.n1166 VDD.n1165 3.1505
R528 VDD.n1163 VDD.n1162 3.1505
R529 VDD.n1160 VDD.n1159 3.1505
R530 VDD.n1158 VDD.n1157 3.1505
R531 VDD.n1155 VDD.n1154 3.1505
R532 VDD.n1168 VDD.n1167 3.1505
R533 VDD.n1172 VDD.n1171 3.1505
R534 VDD.n1192 VDD.n1191 3.1505
R535 VDD.n1189 VDD.n1188 3.1505
R536 VDD.n1182 VDD.n1181 3.1505
R537 VDD.n1180 VDD.n1179 3.1505
R538 VDD.n1177 VDD.n1176 3.1505
R539 VDD.n1175 VDD.n1174 3.1505
R540 VDD.n1194 VDD.n1193 3.1505
R541 VDD.n1198 VDD.n1197 3.1505
R542 VDD.n1117 VDD.n1116 3.1505
R543 VDD.n1114 VDD.n1113 3.1505
R544 VDD.n1111 VDD.n1110 3.1505
R545 VDD.n1108 VDD.n1107 3.1505
R546 VDD.n1105 VDD.n1104 3.1505
R547 VDD.n1103 VDD.n1102 3.1505
R548 VDD.n679 VDD.n678 3.1505
R549 VDD.n943 VDD.n942 3.1505
R550 VDD.n634 VDD.t13 3.1255
R551 VDD.n1055 VDD.t48 3.10434
R552 VDD.n430 VDD.n429 2.6005
R553 VDD.n959 VDD.n958 2.6005
R554 VDD.n960 VDD.n956 2.6005
R555 VDD.n961 VDD.n954 2.6005
R556 VDD.n6 VDD.n5 2.6005
R557 VDD.n748 VDD.n747 2.6005
R558 VDD.n749 VDD.n745 2.6005
R559 VDD.n750 VDD.n743 2.6005
R560 VDD.n3 VDD.n2 2.6005
R561 VDD.n898 VDD.n897 2.6005
R562 VDD.n899 VDD.n895 2.6005
R563 VDD.n900 VDD.n893 2.6005
R564 VDD.n478 VDD.n477 2.6005
R565 VDD.n950 VDD.n949 2.6005
R566 VDD.n951 VDD.n947 2.6005
R567 VDD.n952 VDD.n945 2.6005
R568 VDD.n1107 VDD.n1106 2.40832
R569 VDD.n1110 VDD.n1109 2.40832
R570 VDD.n1113 VDD.n1112 2.40832
R571 VDD.n1116 VDD.n1115 2.40832
R572 VDD.n1197 VDD.n1195 2.40832
R573 VDD.n1197 VDD.n1196 2.40832
R574 VDD.n1171 VDD.n1170 2.40832
R575 VDD.n1151 VDD.n1150 2.40832
R576 VDD.n1134 VDD.n1133 2.40832
R577 VDD.n1130 VDD.n1129 2.40832
R578 VDD.n1154 VDD.n1153 2.40832
R579 VDD.n281 VDD.t0 2.15196
R580 VDD.n749 VDD.n748 2.03528
R581 VDD.n899 VDD.n898 2.03528
R582 VDD.n750 VDD.n749 2.03137
R583 VDD.n900 VDD.n899 2.03137
R584 VDD.n1084 VDD.t31 1.97567
R585 VDD.n241 VDD.n240 1.7598
R586 VDD.n299 VDD.n298 1.75914
R587 VDD.n942 VDD.n941 1.75914
R588 VDD.n667 VDD.n666 1.74343
R589 VDD.n1017 VDD.n1016 1.74343
R590 VDD.n1012 VDD.n1011 1.74343
R591 VDD.n1007 VDD.n1006 1.74343
R592 VDD.n1002 VDD.n1001 1.74343
R593 VDD.n997 VDD.n996 1.74343
R594 VDD.n992 VDD.n991 1.74343
R595 VDD.n987 VDD.n986 1.74343
R596 VDD.n1142 VDD.n1141 1.74343
R597 VDD.n1162 VDD.n1161 1.74343
R598 VDD.n1188 VDD.n1187 1.74343
R599 VDD.n1179 VDD.n1178 1.74343
R600 VDD.n832 VDD.n831 1.74276
R601 VDD.n827 VDD.n826 1.74276
R602 VDD.n822 VDD.n821 1.74276
R603 VDD.n817 VDD.n816 1.74276
R604 VDD.n812 VDD.n811 1.74276
R605 VDD.n807 VDD.n806 1.74276
R606 VDD.n802 VDD.n801 1.74276
R607 VDD.n722 VDD.n721 1.74276
R608 VDD.n701 VDD.n700 1.74276
R609 VDD.n714 VDD.n713 1.74276
R610 VDD.n719 VDD.n718 1.74276
R611 VDD.n728 VDD.n727 1.74276
R612 VDD.n733 VDD.n732 1.74276
R613 VDD.n738 VDD.n737 1.74276
R614 VDD.n304 VDD.n303 1.74276
R615 VDD.n233 VDD.n232 1.74276
R616 VDD.n228 VDD.n227 1.74276
R617 VDD.n223 VDD.n222 1.74276
R618 VDD.n218 VDD.n217 1.74276
R619 VDD.n213 VDD.n212 1.74276
R620 VDD.n208 VDD.n207 1.74276
R621 VDD.n383 VDD.n382 1.74276
R622 VDD.n390 VDD.n389 1.74276
R623 VDD.n376 VDD.n375 1.74276
R624 VDD.n371 VDD.n370 1.74276
R625 VDD.n366 VDD.n365 1.74276
R626 VDD.n587 VDD.n586 1.74276
R627 VDD.n582 VDD.n581 1.74276
R628 VDD.n577 VDD.n576 1.74276
R629 VDD.n572 VDD.n571 1.74276
R630 VDD.n567 VDD.n566 1.74276
R631 VDD.n562 VDD.n561 1.74276
R632 VDD.n557 VDD.n556 1.74276
R633 VDD.n87 VDD.n86 1.74276
R634 VDD.n652 VDD.n651 1.74276
R635 VDD.n647 VDD.n646 1.74276
R636 VDD.n81 VDD.n80 1.74276
R637 VDD.n66 VDD.n65 1.74276
R638 VDD.n71 VDD.n70 1.74276
R639 VDD.n76 VDD.n75 1.74276
R640 VDD.n184 VDD.n183 1.74276
R641 VDD.n179 VDD.n178 1.74276
R642 VDD.n174 VDD.n173 1.74276
R643 VDD.n168 VDD.n167 1.74276
R644 VDD.n494 VDD.n492 1.74276
R645 VDD.n494 VDD.n493 1.74276
R646 VDD.n613 VDD.t15 1.563
R647 VDD.n1102 VDD.n1101 1.42472
R648 VDD.n1137 VDD.n1136 1.42472
R649 VDD.n1174 VDD.n1173 1.42472
R650 VDD.n1191 VDD.n1190 1.42456
R651 VDD.n1165 VDD.n1164 1.42456
R652 VDD.n1157 VDD.n1156 1.42456
R653 VDD.n1145 VDD.n1144 1.42456
R654 VDD.n1125 VDD.n1124 1.42456
R655 VDD.n1020 VDD.n1019 1.42456
R656 VDD.n442 VDD.n441 1.42456
R657 VDD.n447 VDD.n446 1.42456
R658 VDD.n1034 VDD.n1033 1.40117
R659 VDD.n853 VDD.n852 1.36443
R660 VDD.n939 VDD.n938 1.36443
R661 VDD.n345 VDD.n344 1.351
R662 VDD.n509 VDD.n508 1.351
R663 VDD.n880 VDD.t33 1.34158
R664 VDD.n961 VDD.n960 1.27435
R665 VDD.n960 VDD.n959 1.27435
R666 VDD.n952 VDD.n951 1.27435
R667 VDD.n951 VDD.n950 1.27435
R668 VDD.n202 VDD.n198 1.21458
R669 VDD.n33 VDD.n6 1.1255
R670 VDD.n44 VDD.n3 1.1255
R671 VDD.n1035 VDD.n1034 1.0512
R672 VDD.n598 VDD.t2 1.04217
R673 VDD.n876 VDD.n750 1.03159
R674 VDD.n901 VDD.n900 1.03159
R675 VDD.n467 VDD.n430 0.968
R676 VDD.n479 VDD.n478 0.968
R677 VDD.n508 VDD.n507 0.901
R678 VDD.n1061 VDD.n961 0.9005
R679 VDD.n1074 VDD.n952 0.9005
R680 VDD.n852 VDD.n851 0.894284
R681 VDD.n851 VDD.n836 0.894284
R682 VDD.n938 VDD.n937 0.894284
R683 VDD.n937 VDD.n925 0.894284
R684 VDD.n666 VDD.n665 0.705355
R685 VDD.n1033 VDD.n1032 0.705355
R686 VDD.n1033 VDD.n1031 0.705355
R687 VDD.n1033 VDD.n1030 0.705355
R688 VDD.n1033 VDD.n1029 0.705355
R689 VDD.n1033 VDD.n1028 0.705355
R690 VDD.n1033 VDD.n1027 0.705355
R691 VDD.n1033 VDD.n1026 0.705355
R692 VDD.n1033 VDD.n1025 0.705355
R693 VDD.n1186 VDD.n1185 0.705355
R694 VDD.n1186 VDD.n1184 0.705355
R695 VDD.n1187 VDD.n1186 0.705355
R696 VDD.n851 VDD.n850 0.705118
R697 VDD.n851 VDD.n849 0.705118
R698 VDD.n851 VDD.n846 0.705118
R699 VDD.n851 VDD.n842 0.705118
R700 VDD.n851 VDD.n838 0.705118
R701 VDD.n851 VDD.n837 0.705118
R702 VDD.n937 VDD.n931 0.705118
R703 VDD.n937 VDD.n935 0.705118
R704 VDD.n937 VDD.n936 0.705118
R705 VDD.n937 VDD.n927 0.705118
R706 VDD.n202 VDD.n201 0.705118
R707 VDD.n239 VDD.n238 0.705118
R708 VDD.n360 VDD.n359 0.705118
R709 VDD.n384 VDD.n383 0.705118
R710 VDD.n381 VDD.n380 0.705118
R711 VDD.n380 VDD.n379 0.705118
R712 VDD.n380 VDD.n378 0.705118
R713 VDD.n507 VDD.n506 0.705118
R714 VDD.n507 VDD.n505 0.705118
R715 VDD.n507 VDD.n504 0.705118
R716 VDD.n507 VDD.n503 0.705118
R717 VDD.n507 VDD.n502 0.705118
R718 VDD.n507 VDD.n501 0.705118
R719 VDD.n507 VDD.n500 0.705118
R720 VDD.n507 VDD.n499 0.705118
R721 VDD.n507 VDD.n498 0.705118
R722 VDD.n507 VDD.n497 0.705118
R723 VDD.n507 VDD.n496 0.705118
R724 VDD.n665 VDD.n663 0.705118
R725 VDD.n665 VDD.n664 0.705118
R726 VDD.n665 VDD.n662 0.705118
R727 VDD.n665 VDD.n660 0.705118
R728 VDD.n665 VDD.n661 0.705118
R729 VDD.n665 VDD.n659 0.705118
R730 VDD.n665 VDD.n658 0.705118
R731 VDD.n677 VDD.n494 0.705118
R732 VDD.n240 VDD.n239 0.697168
R733 VDD.n851 VDD.n848 0.69693
R734 VDD.n851 VDD.n844 0.69693
R735 VDD.n851 VDD.n840 0.69693
R736 VDD.n937 VDD.n929 0.69693
R737 VDD.n937 VDD.n933 0.69693
R738 VDD.n851 VDD.n847 0.677271
R739 VDD.n851 VDD.n845 0.677271
R740 VDD.n851 VDD.n843 0.677271
R741 VDD.n851 VDD.n841 0.677271
R742 VDD.n851 VDD.n839 0.677271
R743 VDD.n708 VDD.n707 0.677271
R744 VDD.n937 VDD.n930 0.677271
R745 VDD.n937 VDD.n932 0.677271
R746 VDD.n937 VDD.n934 0.677271
R747 VDD.n937 VDD.n928 0.677271
R748 VDD.n937 VDD.n926 0.677271
R749 VDD.n945 VDD.t51 0.607167
R750 VDD.n945 VDD.n944 0.607167
R751 VDD.n947 VDD.t21 0.607167
R752 VDD.n947 VDD.n946 0.607167
R753 VDD.n949 VDD.t40 0.607167
R754 VDD.n949 VDD.n948 0.607167
R755 VDD.n477 VDD.t68 0.607167
R756 VDD.n477 VDD.n476 0.607167
R757 VDD.n954 VDD.t19 0.607167
R758 VDD.n954 VDD.n953 0.607167
R759 VDD.n956 VDD.t81 0.607167
R760 VDD.n956 VDD.n955 0.607167
R761 VDD.n958 VDD.t82 0.607167
R762 VDD.n958 VDD.n957 0.607167
R763 VDD.n429 VDD.t38 0.607167
R764 VDD.n429 VDD.n428 0.607167
R765 VDD.n893 VDD.t56 0.607167
R766 VDD.n893 VDD.n892 0.607167
R767 VDD.n895 VDD.t7 0.607167
R768 VDD.n895 VDD.n894 0.607167
R769 VDD.n897 VDD.t32 0.607167
R770 VDD.n897 VDD.n896 0.607167
R771 VDD.n2 VDD.t47 0.607167
R772 VDD.n2 VDD.n1 0.607167
R773 VDD.n743 VDD.t59 0.607167
R774 VDD.n743 VDD.n742 0.607167
R775 VDD.n745 VDD.t5 0.607167
R776 VDD.n745 VDD.n744 0.607167
R777 VDD.n747 VDD.t41 0.607167
R778 VDD.n747 VDD.n746 0.607167
R779 VDD.n5 VDD.t46 0.607167
R780 VDD.n5 VDD.n4 0.607167
R781 VDD.n396 VDD.n395 0.530311
R782 VDD.n239 VDD.n237 0.430793
R783 VDD.n272 VDD.t29 0.430793
R784 VDD.n677 VDD.n676 0.356659
R785 VDD.n681 VDD.n680 0.34342
R786 VDD.n1186 VDD.n1183 0.282667
R787 VDD.n1033 VDD.n1024 0.282667
R788 VDD.n665 VDD.n657 0.260917
R789 VDD.n507 VDD.n495 0.260917
R790 VDD.n395 VDD.n394 0.260092
R791 VDD VDD.n943 0.222544
R792 VDD.n198 VDD.n197 0.129466
R793 VDD.n197 VDD.n196 0.123603
R794 VDD VDD.n1199 0.121376
R795 VDD.n196 VDD.n194 0.106362
R796 VDD.n396 VDD.n83 0.0963273
R797 VDD.n418 VDD.n416 0.0932551
R798 VDD.n689 VDD.n687 0.0932551
R799 VDD.n699 VDD.n697 0.0932551
R800 VDD.n717 VDD.n715 0.0932551
R801 VDD.n736 VDD.n734 0.0932551
R802 VDD.n835 VDD.n833 0.0932551
R803 VDD.n825 VDD.n823 0.0932551
R804 VDD.n815 VDD.n813 0.0932551
R805 VDD.n805 VDD.n803 0.0932551
R806 VDD.n796 VDD.n794 0.0932551
R807 VDD.n786 VDD.n784 0.0932551
R808 VDD.n778 VDD.n776 0.0932551
R809 VDD.n770 VDD.n768 0.0932551
R810 VDD.n762 VDD.n760 0.0932551
R811 VDD.n754 VDD.n752 0.0932551
R812 VDD.n863 VDD.n860 0.0932551
R813 VDD.n875 VDD.n872 0.0932551
R814 VDD.n888 VDD.n885 0.0932551
R815 VDD.n910 VDD.n907 0.0932551
R816 VDD.n922 VDD.n919 0.0932551
R817 VDD.n24 VDD.n22 0.0932551
R818 VDD.n32 VDD.n30 0.0932551
R819 VDD.n41 VDD.n39 0.0932551
R820 VDD.n50 VDD.n48 0.0932551
R821 VDD.n58 VDD.n56 0.0932551
R822 VDD.n403 VDD.n401 0.0932551
R823 VDD.n395 VDD.n186 0.0911122
R824 VDD.n397 VDD.n396 0.0905
R825 VDD.n414 VDD.n412 0.0886633
R826 VDD.n685 VDD.n683 0.0886633
R827 VDD.n712 VDD.n710 0.0886633
R828 VDD.n731 VDD.n729 0.0886633
R829 VDD.n820 VDD.n818 0.0886633
R830 VDD.n800 VDD.n798 0.0886633
R831 VDD.n790 VDD.n788 0.0886633
R832 VDD.n774 VDD.n772 0.0886633
R833 VDD.n758 VDD.n756 0.0886633
R834 VDD.n12 VDD.n10 0.0886633
R835 VDD.n882 VDD.n879 0.0886633
R836 VDD.n916 VDD.n913 0.0886633
R837 VDD.n37 VDD.n35 0.0886633
R838 VDD.n54 VDD.n52 0.0886633
R839 VDD.n300 VDD.n297 0.0886633
R840 VDD.n242 VDD.n236 0.0886633
R841 VDD.n594 VDD.n591 0.0877449
R842 VDD.n343 VDD.n341 0.0877449
R843 VDD.n1039 VDD.n1036 0.0877449
R844 VDD.n645 VDD.n642 0.0868265
R845 VDD.n642 VDD.n639 0.0868265
R846 VDD.n639 VDD.n636 0.0868265
R847 VDD.n636 VDD.n633 0.0868265
R848 VDD.n633 VDD.n630 0.0868265
R849 VDD.n630 VDD.n627 0.0868265
R850 VDD.n627 VDD.n624 0.0868265
R851 VDD.n624 VDD.n621 0.0868265
R852 VDD.n621 VDD.n618 0.0868265
R853 VDD.n618 VDD.n615 0.0868265
R854 VDD.n615 VDD.n612 0.0868265
R855 VDD.n612 VDD.n609 0.0868265
R856 VDD.n609 VDD.n606 0.0868265
R857 VDD.n606 VDD.n603 0.0868265
R858 VDD.n603 VDD.n600 0.0868265
R859 VDD.n600 VDD.n597 0.0868265
R860 VDD.n597 VDD.n594 0.0868265
R861 VDD.n424 VDD.n422 0.0868265
R862 VDD.n422 VDD.n420 0.0868265
R863 VDD.n420 VDD.n418 0.0868265
R864 VDD.n416 VDD.n414 0.0868265
R865 VDD.n412 VDD.n410 0.0868265
R866 VDD.n691 VDD.n689 0.0868265
R867 VDD.n687 VDD.n685 0.0868265
R868 VDD.n704 VDD.n702 0.0868265
R869 VDD.n702 VDD.n699 0.0868265
R870 VDD.n697 VDD.n695 0.0868265
R871 VDD.n720 VDD.n717 0.0868265
R872 VDD.n715 VDD.n712 0.0868265
R873 VDD.n741 VDD.n739 0.0868265
R874 VDD.n739 VDD.n736 0.0868265
R875 VDD.n734 VDD.n731 0.0868265
R876 VDD.n729 VDD.n726 0.0868265
R877 VDD.n833 VDD.n830 0.0868265
R878 VDD.n830 VDD.n828 0.0868265
R879 VDD.n828 VDD.n825 0.0868265
R880 VDD.n823 VDD.n820 0.0868265
R881 VDD.n818 VDD.n815 0.0868265
R882 VDD.n813 VDD.n810 0.0868265
R883 VDD.n810 VDD.n808 0.0868265
R884 VDD.n808 VDD.n805 0.0868265
R885 VDD.n803 VDD.n800 0.0868265
R886 VDD.n798 VDD.n796 0.0868265
R887 VDD.n794 VDD.n792 0.0868265
R888 VDD.n792 VDD.n790 0.0868265
R889 VDD.n788 VDD.n786 0.0868265
R890 VDD.n784 VDD.n782 0.0868265
R891 VDD.n782 VDD.n780 0.0868265
R892 VDD.n780 VDD.n778 0.0868265
R893 VDD.n776 VDD.n774 0.0868265
R894 VDD.n772 VDD.n770 0.0868265
R895 VDD.n768 VDD.n766 0.0868265
R896 VDD.n766 VDD.n764 0.0868265
R897 VDD.n764 VDD.n762 0.0868265
R898 VDD.n760 VDD.n758 0.0868265
R899 VDD.n756 VDD.n754 0.0868265
R900 VDD.n10 VDD.n8 0.0868265
R901 VDD.n14 VDD.n12 0.0868265
R902 VDD.n16 VDD.n14 0.0868265
R903 VDD.n857 VDD.n854 0.0868265
R904 VDD.n860 VDD.n857 0.0868265
R905 VDD.n866 VDD.n863 0.0868265
R906 VDD.n869 VDD.n866 0.0868265
R907 VDD.n872 VDD.n869 0.0868265
R908 VDD.n885 VDD.n882 0.0868265
R909 VDD.n891 VDD.n888 0.0868265
R910 VDD.n907 VDD.n904 0.0868265
R911 VDD.n913 VDD.n910 0.0868265
R912 VDD.n919 VDD.n916 0.0868265
R913 VDD.n924 VDD.n922 0.0868265
R914 VDD.n20 VDD.n18 0.0868265
R915 VDD.n22 VDD.n20 0.0868265
R916 VDD.n26 VDD.n24 0.0868265
R917 VDD.n28 VDD.n26 0.0868265
R918 VDD.n30 VDD.n28 0.0868265
R919 VDD.n39 VDD.n37 0.0868265
R920 VDD.n43 VDD.n41 0.0868265
R921 VDD.n48 VDD.n46 0.0868265
R922 VDD.n52 VDD.n50 0.0868265
R923 VDD.n56 VDD.n54 0.0868265
R924 VDD.n407 VDD.n405 0.0868265
R925 VDD.n405 VDD.n403 0.0868265
R926 VDD.n401 VDD.n399 0.0868265
R927 VDD.n356 VDD.n354 0.0868265
R928 VDD.n354 VDD.n352 0.0868265
R929 VDD.n352 VDD.n350 0.0868265
R930 VDD.n377 VDD.n374 0.0868265
R931 VDD.n374 VDD.n372 0.0868265
R932 VDD.n372 VDD.n369 0.0868265
R933 VDD.n369 VDD.n367 0.0868265
R934 VDD.n367 VDD.n364 0.0868265
R935 VDD.n364 VDD.n362 0.0868265
R936 VDD.n393 VDD.n391 0.0868265
R937 VDD.n391 VDD.n388 0.0868265
R938 VDD.n388 VDD.n386 0.0868265
R939 VDD.n309 VDD.n307 0.0868265
R940 VDD.n311 VDD.n309 0.0868265
R941 VDD.n313 VDD.n311 0.0868265
R942 VDD.n315 VDD.n313 0.0868265
R943 VDD.n317 VDD.n315 0.0868265
R944 VDD.n319 VDD.n317 0.0868265
R945 VDD.n321 VDD.n319 0.0868265
R946 VDD.n323 VDD.n321 0.0868265
R947 VDD.n325 VDD.n323 0.0868265
R948 VDD.n327 VDD.n325 0.0868265
R949 VDD.n329 VDD.n327 0.0868265
R950 VDD.n331 VDD.n329 0.0868265
R951 VDD.n333 VDD.n331 0.0868265
R952 VDD.n335 VDD.n333 0.0868265
R953 VDD.n337 VDD.n335 0.0868265
R954 VDD.n339 VDD.n337 0.0868265
R955 VDD.n341 VDD.n339 0.0868265
R956 VDD.n192 VDD.n190 0.0868265
R957 VDD.n190 VDD.n188 0.0868265
R958 VDD.n305 VDD.n302 0.0868265
R959 VDD.n236 VDD.n234 0.0868265
R960 VDD.n234 VDD.n231 0.0868265
R961 VDD.n231 VDD.n229 0.0868265
R962 VDD.n229 VDD.n226 0.0868265
R963 VDD.n226 VDD.n224 0.0868265
R964 VDD.n224 VDD.n221 0.0868265
R965 VDD.n221 VDD.n219 0.0868265
R966 VDD.n219 VDD.n216 0.0868265
R967 VDD.n216 VDD.n214 0.0868265
R968 VDD.n214 VDD.n211 0.0868265
R969 VDD.n211 VDD.n209 0.0868265
R970 VDD.n209 VDD.n206 0.0868265
R971 VDD.n206 VDD.n204 0.0868265
R972 VDD.n247 VDD.n244 0.0868265
R973 VDD.n250 VDD.n247 0.0868265
R974 VDD.n253 VDD.n250 0.0868265
R975 VDD.n256 VDD.n253 0.0868265
R976 VDD.n259 VDD.n256 0.0868265
R977 VDD.n262 VDD.n259 0.0868265
R978 VDD.n265 VDD.n262 0.0868265
R979 VDD.n268 VDD.n265 0.0868265
R980 VDD.n271 VDD.n268 0.0868265
R981 VDD.n274 VDD.n271 0.0868265
R982 VDD.n277 VDD.n274 0.0868265
R983 VDD.n280 VDD.n277 0.0868265
R984 VDD.n283 VDD.n280 0.0868265
R985 VDD.n286 VDD.n283 0.0868265
R986 VDD.n289 VDD.n286 0.0868265
R987 VDD.n292 VDD.n289 0.0868265
R988 VDD.n295 VDD.n292 0.0868265
R989 VDD.n670 VDD.n668 0.0868265
R990 VDD.n655 VDD.n653 0.0868265
R991 VDD.n653 VDD.n650 0.0868265
R992 VDD.n650 VDD.n648 0.0868265
R993 VDD.n82 VDD.n79 0.0868265
R994 VDD.n79 VDD.n77 0.0868265
R995 VDD.n77 VDD.n74 0.0868265
R996 VDD.n74 VDD.n72 0.0868265
R997 VDD.n72 VDD.n69 0.0868265
R998 VDD.n69 VDD.n67 0.0868265
R999 VDD.n67 VDD.n64 0.0868265
R1000 VDD.n88 VDD.n85 0.0868265
R1001 VDD.n185 VDD.n182 0.0868265
R1002 VDD.n182 VDD.n180 0.0868265
R1003 VDD.n180 VDD.n177 0.0868265
R1004 VDD.n177 VDD.n175 0.0868265
R1005 VDD.n175 VDD.n172 0.0868265
R1006 VDD.n169 VDD.n166 0.0868265
R1007 VDD.n166 VDD.n164 0.0868265
R1008 VDD.n164 VDD.n162 0.0868265
R1009 VDD.n162 VDD.n160 0.0868265
R1010 VDD.n160 VDD.n158 0.0868265
R1011 VDD.n158 VDD.n156 0.0868265
R1012 VDD.n156 VDD.n154 0.0868265
R1013 VDD.n154 VDD.n152 0.0868265
R1014 VDD.n149 VDD.n147 0.0868265
R1015 VDD.n147 VDD.n145 0.0868265
R1016 VDD.n145 VDD.n143 0.0868265
R1017 VDD.n143 VDD.n141 0.0868265
R1018 VDD.n138 VDD.n136 0.0868265
R1019 VDD.n134 VDD.n132 0.0868265
R1020 VDD.n132 VDD.n130 0.0868265
R1021 VDD.n130 VDD.n128 0.0868265
R1022 VDD.n128 VDD.n126 0.0868265
R1023 VDD.n126 VDD.n124 0.0868265
R1024 VDD.n124 VDD.n122 0.0868265
R1025 VDD.n122 VDD.n120 0.0868265
R1026 VDD.n120 VDD.n118 0.0868265
R1027 VDD.n118 VDD.n116 0.0868265
R1028 VDD.n116 VDD.n114 0.0868265
R1029 VDD.n114 VDD.n112 0.0868265
R1030 VDD.n112 VDD.n110 0.0868265
R1031 VDD.n110 VDD.n108 0.0868265
R1032 VDD.n108 VDD.n106 0.0868265
R1033 VDD.n106 VDD.n104 0.0868265
R1034 VDD.n104 VDD.n102 0.0868265
R1035 VDD.n102 VDD.n100 0.0868265
R1036 VDD.n100 VDD.n98 0.0868265
R1037 VDD.n98 VDD.n96 0.0868265
R1038 VDD.n96 VDD.n94 0.0868265
R1039 VDD.n94 VDD.n92 0.0868265
R1040 VDD.n590 VDD.n588 0.0868265
R1041 VDD.n588 VDD.n585 0.0868265
R1042 VDD.n585 VDD.n583 0.0868265
R1043 VDD.n583 VDD.n580 0.0868265
R1044 VDD.n580 VDD.n578 0.0868265
R1045 VDD.n578 VDD.n575 0.0868265
R1046 VDD.n575 VDD.n573 0.0868265
R1047 VDD.n573 VDD.n570 0.0868265
R1048 VDD.n570 VDD.n568 0.0868265
R1049 VDD.n568 VDD.n565 0.0868265
R1050 VDD.n565 VDD.n563 0.0868265
R1051 VDD.n563 VDD.n560 0.0868265
R1052 VDD.n560 VDD.n558 0.0868265
R1053 VDD.n558 VDD.n555 0.0868265
R1054 VDD.n555 VDD.n553 0.0868265
R1055 VDD.n553 VDD.n551 0.0868265
R1056 VDD.n551 VDD.n549 0.0868265
R1057 VDD.n549 VDD.n547 0.0868265
R1058 VDD.n547 VDD.n545 0.0868265
R1059 VDD.n545 VDD.n543 0.0868265
R1060 VDD.n543 VDD.n541 0.0868265
R1061 VDD.n541 VDD.n539 0.0868265
R1062 VDD.n539 VDD.n537 0.0868265
R1063 VDD.n537 VDD.n535 0.0868265
R1064 VDD.n535 VDD.n533 0.0868265
R1065 VDD.n533 VDD.n531 0.0868265
R1066 VDD.n531 VDD.n529 0.0868265
R1067 VDD.n529 VDD.n527 0.0868265
R1068 VDD.n527 VDD.n525 0.0868265
R1069 VDD.n525 VDD.n523 0.0868265
R1070 VDD.n523 VDD.n521 0.0868265
R1071 VDD.n521 VDD.n519 0.0868265
R1072 VDD.n519 VDD.n517 0.0868265
R1073 VDD.n517 VDD.n515 0.0868265
R1074 VDD.n515 VDD.n513 0.0868265
R1075 VDD.n513 VDD.n511 0.0868265
R1076 VDD.n1023 VDD.n1021 0.0868265
R1077 VDD.n1021 VDD.n1018 0.0868265
R1078 VDD.n1018 VDD.n1015 0.0868265
R1079 VDD.n1015 VDD.n1013 0.0868265
R1080 VDD.n1013 VDD.n1010 0.0868265
R1081 VDD.n1010 VDD.n1008 0.0868265
R1082 VDD.n1008 VDD.n1005 0.0868265
R1083 VDD.n1005 VDD.n1003 0.0868265
R1084 VDD.n1003 VDD.n1000 0.0868265
R1085 VDD.n1000 VDD.n998 0.0868265
R1086 VDD.n998 VDD.n995 0.0868265
R1087 VDD.n995 VDD.n993 0.0868265
R1088 VDD.n993 VDD.n990 0.0868265
R1089 VDD.n990 VDD.n988 0.0868265
R1090 VDD.n988 VDD.n985 0.0868265
R1091 VDD.n985 VDD.n983 0.0868265
R1092 VDD.n983 VDD.n981 0.0868265
R1093 VDD.n981 VDD.n979 0.0868265
R1094 VDD.n979 VDD.n977 0.0868265
R1095 VDD.n977 VDD.n975 0.0868265
R1096 VDD.n975 VDD.n973 0.0868265
R1097 VDD.n973 VDD.n971 0.0868265
R1098 VDD.n971 VDD.n969 0.0868265
R1099 VDD.n969 VDD.n967 0.0868265
R1100 VDD.n967 VDD.n965 0.0868265
R1101 VDD.n965 VDD.n963 0.0868265
R1102 VDD.n434 VDD.n432 0.0868265
R1103 VDD.n436 VDD.n434 0.0868265
R1104 VDD.n438 VDD.n436 0.0868265
R1105 VDD.n440 VDD.n438 0.0868265
R1106 VDD.n443 VDD.n440 0.0868265
R1107 VDD.n445 VDD.n443 0.0868265
R1108 VDD.n448 VDD.n445 0.0868265
R1109 VDD.n491 VDD.n489 0.0868265
R1110 VDD.n489 VDD.n487 0.0868265
R1111 VDD.n487 VDD.n485 0.0868265
R1112 VDD.n485 VDD.n483 0.0868265
R1113 VDD.n483 VDD.n481 0.0868265
R1114 VDD.n475 VDD.n473 0.0868265
R1115 VDD.n473 VDD.n471 0.0868265
R1116 VDD.n471 VDD.n469 0.0868265
R1117 VDD.n466 VDD.n464 0.0868265
R1118 VDD.n464 VDD.n462 0.0868265
R1119 VDD.n462 VDD.n460 0.0868265
R1120 VDD.n460 VDD.n458 0.0868265
R1121 VDD.n458 VDD.n456 0.0868265
R1122 VDD.n456 VDD.n454 0.0868265
R1123 VDD.n454 VDD.n452 0.0868265
R1124 VDD.n452 VDD.n450 0.0868265
R1125 VDD.n1100 VDD.n1098 0.0868265
R1126 VDD.n1098 VDD.n1095 0.0868265
R1127 VDD.n1095 VDD.n1092 0.0868265
R1128 VDD.n1092 VDD.n1089 0.0868265
R1129 VDD.n1089 VDD.n1086 0.0868265
R1130 VDD.n1086 VDD.n1083 0.0868265
R1131 VDD.n1083 VDD.n1080 0.0868265
R1132 VDD.n1080 VDD.n1077 0.0868265
R1133 VDD.n1073 VDD.n1070 0.0868265
R1134 VDD.n1070 VDD.n1067 0.0868265
R1135 VDD.n1067 VDD.n1064 0.0868265
R1136 VDD.n1060 VDD.n1057 0.0868265
R1137 VDD.n1057 VDD.n1054 0.0868265
R1138 VDD.n1054 VDD.n1051 0.0868265
R1139 VDD.n1051 VDD.n1048 0.0868265
R1140 VDD.n1048 VDD.n1045 0.0868265
R1141 VDD.n1045 VDD.n1042 0.0868265
R1142 VDD.n1042 VDD.n1039 0.0868265
R1143 VDD.n1105 VDD.n1103 0.0868265
R1144 VDD.n1108 VDD.n1105 0.0868265
R1145 VDD.n1111 VDD.n1108 0.0868265
R1146 VDD.n1114 VDD.n1111 0.0868265
R1147 VDD.n1117 VDD.n1114 0.0868265
R1148 VDD.n1198 VDD.n1194 0.0868265
R1149 VDD.n1194 VDD.n1192 0.0868265
R1150 VDD.n1192 VDD.n1189 0.0868265
R1151 VDD.n1189 VDD.n1182 0.0868265
R1152 VDD.n1182 VDD.n1180 0.0868265
R1153 VDD.n1180 VDD.n1177 0.0868265
R1154 VDD.n1177 VDD.n1175 0.0868265
R1155 VDD.n1175 VDD.n1172 0.0868265
R1156 VDD.n1168 VDD.n1166 0.0868265
R1157 VDD.n1166 VDD.n1163 0.0868265
R1158 VDD.n1163 VDD.n1160 0.0868265
R1159 VDD.n1160 VDD.n1158 0.0868265
R1160 VDD.n1158 VDD.n1155 0.0868265
R1161 VDD.n1155 VDD.n1152 0.0868265
R1162 VDD.n1148 VDD.n1146 0.0868265
R1163 VDD.n1146 VDD.n1143 0.0868265
R1164 VDD.n1143 VDD.n1140 0.0868265
R1165 VDD.n1140 VDD.n1138 0.0868265
R1166 VDD.n1138 VDD.n1135 0.0868265
R1167 VDD.n1131 VDD.n1128 0.0868265
R1168 VDD.n1128 VDD.n1126 0.0868265
R1169 VDD.n1126 VDD.n1123 0.0868265
R1170 VDD.n1123 VDD.n1121 0.0868265
R1171 VDD.n1121 VDD.n1119 0.0868265
R1172 VDD.n1135 VDD.n1132 0.0849898
R1173 VDD.n469 VDD.n467 0.0840714
R1174 VDD.n1064 VDD.n1061 0.0840714
R1175 VDD.n394 VDD.n393 0.0822347
R1176 VDD.n170 VDD.n169 0.0794796
R1177 VDD.n680 VDD.n679 0.0785612
R1178 VDD.n141 VDD.n139 0.0776429
R1179 VDD.n384 VDD.n377 0.0758061
R1180 VDD.n150 VDD.n149 0.0758061
R1181 VDD.n708 VDD.n704 0.0748878
R1182 VDD.n656 VDD.n655 0.0748878
R1183 VDD.n724 VDD.n720 0.073051
R1184 VDD.n360 VDD.n356 0.0721327
R1185 VDD.n83 VDD.n62 0.0721327
R1186 VDD.n202 VDD.n192 0.0712143
R1187 VDD.n1199 VDD.n1117 0.0712143
R1188 VDD.n876 VDD.n875 0.0702959
R1189 VDD.n33 VDD.n32 0.0702959
R1190 VDD.n1169 VDD.n1168 0.0702959
R1191 VDD.n186 VDD.n88 0.0684592
R1192 VDD.n726 VDD.n724 0.0675408
R1193 VDD.n204 VDD.n202 0.0675408
R1194 VDD.n710 VDD.n708 0.0657041
R1195 VDD.n397 VDD.n60 0.0620306
R1196 VDD.n904 VDD.n901 0.0601939
R1197 VDD.n46 VDD.n44 0.0601939
R1198 VDD.n1149 VDD.n1148 0.0574388
R1199 VDD.n479 VDD.n475 0.0546837
R1200 VDD.n1074 VDD.n1073 0.0546837
R1201 VDD.n362 VDD.n360 0.0528469
R1202 VDD.n408 VDD.n407 0.0500918
R1203 VDD.n386 VDD.n384 0.0491735
R1204 VDD.n943 VDD.n940 0.0455
R1205 VDD.n244 VDD.n242 0.0455
R1206 VDD.n673 VDD.n670 0.0436633
R1207 VDD.n940 VDD.n924 0.0436633
R1208 VDD.n854 VDD.n835 0.0436633
R1209 VDD.n18 VDD.n16 0.0436633
R1210 VDD.n297 VDD.n295 0.0436633
R1211 VDD.n307 VDD.n305 0.0436633
R1212 VDD.n1103 VDD.n1100 0.0436633
R1213 VDD.n346 VDD.n343 0.0427449
R1214 VDD.n591 VDD.n590 0.0427449
R1215 VDD.n1036 VDD.n1023 0.0427449
R1216 VDD.n136 VDD.n134 0.0427449
R1217 VDD.n92 VDD.n90 0.0427449
R1218 VDD.n450 VDD.n448 0.0427449
R1219 VDD.n60 VDD.n58 0.0418265
R1220 VDD.n677 VDD.n491 0.0390714
R1221 VDD.n681 VDD.n424 0.0326429
R1222 VDD.n350 VDD.n348 0.0326429
R1223 VDD.n481 VDD.n479 0.0326429
R1224 VDD.n1077 VDD.n1074 0.0326429
R1225 VDD.n1152 VDD.n1149 0.0298878
R1226 VDD.n693 VDD.n691 0.028051
R1227 VDD.n901 VDD.n891 0.0271327
R1228 VDD.n44 VDD.n43 0.0271327
R1229 VDD.n399 VDD.n397 0.0271327
R1230 VDD.n679 VDD.n677 0.0262143
R1231 VDD.n683 VDD.n681 0.0216225
R1232 VDD.n695 VDD.n693 0.0216225
R1233 VDD.n186 VDD.n185 0.0188673
R1234 VDD.n879 VDD.n876 0.0170306
R1235 VDD.n35 VDD.n33 0.0170306
R1236 VDD.n1172 VDD.n1169 0.0170306
R1237 VDD.n1199 VDD.n1198 0.0161122
R1238 VDD.n83 VDD.n82 0.0151939
R1239 VDD.n676 VDD.n645 0.0142755
R1240 VDD.n668 VDD.n656 0.0124388
R1241 VDD.n152 VDD.n150 0.0115204
R1242 VDD.n139 VDD.n138 0.00968367
R1243 VDD.n676 VDD.n673 0.00876531
R1244 VDD.n680 VDD.n427 0.00876531
R1245 VDD.n172 VDD.n170 0.00784694
R1246 VDD.n394 VDD.n300 0.00692857
R1247 VDD.n348 VDD.n346 0.0060102
R1248 VDD.n943 VDD.n741 0.00417347
R1249 VDD.n467 VDD.n466 0.0032551
R1250 VDD.n1061 VDD.n1060 0.0032551
R1251 VDD.n410 VDD.n408 0.00233673
R1252 VDD.n1132 VDD.n1131 0.00233673
R1253 a_n2814_n10181.n0 a_n2814_n10181.t12 52.4934
R1254 a_n2814_n10181.n6 a_n2814_n10181.t14 52.1689
R1255 a_n2814_n10181.n57 a_n2814_n10181.t16 51.5691
R1256 a_n2814_n10181.n2 a_n2814_n10181.t10 50.3958
R1257 a_n2814_n10181.n19 a_n2814_n10181.t46 45.8862
R1258 a_n2814_n10181.n20 a_n2814_n10181.t37 45.8862
R1259 a_n2814_n10181.n21 a_n2814_n10181.t28 45.8862
R1260 a_n2814_n10181.n22 a_n2814_n10181.t43 45.8862
R1261 a_n2814_n10181.n26 a_n2814_n10181.t35 45.8862
R1262 a_n2814_n10181.n25 a_n2814_n10181.t49 45.8862
R1263 a_n2814_n10181.n24 a_n2814_n10181.t45 45.8862
R1264 a_n2814_n10181.n23 a_n2814_n10181.t36 45.8862
R1265 a_n2814_n10181.n19 a_n2814_n10181.t27 45.6255
R1266 a_n2814_n10181.n20 a_n2814_n10181.t20 45.6255
R1267 a_n2814_n10181.n21 a_n2814_n10181.t41 45.6255
R1268 a_n2814_n10181.n22 a_n2814_n10181.t22 45.6255
R1269 a_n2814_n10181.n26 a_n2814_n10181.t48 45.6255
R1270 a_n2814_n10181.n25 a_n2814_n10181.t29 45.6255
R1271 a_n2814_n10181.n24 a_n2814_n10181.t25 45.6255
R1272 a_n2814_n10181.n33 a_n2814_n10181.t44 45.6255
R1273 a_n2814_n10181.n28 a_n2814_n10181.t23 45.6255
R1274 a_n2814_n10181.n37 a_n2814_n10181.t42 45.6255
R1275 a_n2814_n10181.n29 a_n2814_n10181.t33 45.6255
R1276 a_n2814_n10181.n38 a_n2814_n10181.t34 45.6255
R1277 a_n2814_n10181.n30 a_n2814_n10181.t26 45.6255
R1278 a_n2814_n10181.n39 a_n2814_n10181.t24 45.6255
R1279 a_n2814_n10181.n31 a_n2814_n10181.t39 45.6255
R1280 a_n2814_n10181.n40 a_n2814_n10181.t38 45.6255
R1281 a_n2814_n10181.n35 a_n2814_n10181.t51 45.6255
R1282 a_n2814_n10181.n44 a_n2814_n10181.t31 45.6255
R1283 a_n2814_n10181.n34 a_n2814_n10181.t30 45.6255
R1284 a_n2814_n10181.n43 a_n2814_n10181.t47 45.6255
R1285 a_n2814_n10181.n32 a_n2814_n10181.t21 45.6255
R1286 a_n2814_n10181.n41 a_n2814_n10181.t32 45.6255
R1287 a_n2814_n10181.n42 a_n2814_n10181.t40 45.6255
R1288 a_n2814_n10181.n23 a_n2814_n10181.t50 45.6255
R1289 a_n2814_n10181.n29 a_n2814_n10181.n28 11.9189
R1290 a_n2814_n10181.n30 a_n2814_n10181.n29 11.9189
R1291 a_n2814_n10181.n31 a_n2814_n10181.n30 11.9189
R1292 a_n2814_n10181.n35 a_n2814_n10181.n34 11.9189
R1293 a_n2814_n10181.n34 a_n2814_n10181.n33 11.9189
R1294 a_n2814_n10181.n33 a_n2814_n10181.n32 11.9189
R1295 a_n2814_n10181.n38 a_n2814_n10181.n37 11.9189
R1296 a_n2814_n10181.n39 a_n2814_n10181.n38 11.9189
R1297 a_n2814_n10181.n40 a_n2814_n10181.n39 11.9189
R1298 a_n2814_n10181.n44 a_n2814_n10181.n43 11.9189
R1299 a_n2814_n10181.n43 a_n2814_n10181.n42 11.9189
R1300 a_n2814_n10181.n42 a_n2814_n10181.n41 11.9189
R1301 a_n2814_n10181.n20 a_n2814_n10181.n19 11.9189
R1302 a_n2814_n10181.n21 a_n2814_n10181.n20 11.9189
R1303 a_n2814_n10181.n22 a_n2814_n10181.n21 11.9189
R1304 a_n2814_n10181.n26 a_n2814_n10181.n25 11.9189
R1305 a_n2814_n10181.n25 a_n2814_n10181.n24 11.9189
R1306 a_n2814_n10181.n24 a_n2814_n10181.n23 11.9189
R1307 a_n2814_n10181.n52 a_n2814_n10181.n51 7.2292
R1308 a_n2814_n10181.n46 a_n2814_n10181.n36 6.65848
R1309 a_n2814_n10181.n36 a_n2814_n10181.n31 6.10866
R1310 a_n2814_n10181.n45 a_n2814_n10181.n40 6.03417
R1311 a_n2814_n10181.n27 a_n2814_n10181.n22 6.03417
R1312 a_n2814_n10181.n48 a_n2814_n10181.n47 5.89239
R1313 a_n2814_n10181.n45 a_n2814_n10181.n44 5.88519
R1314 a_n2814_n10181.n27 a_n2814_n10181.n26 5.88519
R1315 a_n2814_n10181.n46 a_n2814_n10181.n45 5.88439
R1316 a_n2814_n10181.n47 a_n2814_n10181.n27 5.88428
R1317 a_n2814_n10181.n36 a_n2814_n10181.n35 5.8107
R1318 a_n2814_n10181.n15 a_n2814_n10181.t9 4.61117
R1319 a_n2814_n10181.n14 a_n2814_n10181.n12 4.61117
R1320 a_n2814_n10181.n49 a_n2814_n10181.n16 4.61089
R1321 a_n2814_n10181.n48 a_n2814_n10181.n18 4.2863
R1322 a_n2814_n10181.n15 a_n2814_n10181.t7 3.20717
R1323 a_n2814_n10181.n14 a_n2814_n10181.n13 3.20717
R1324 a_n2814_n10181.n7 a_n2814_n10181.n5 3.1505
R1325 a_n2814_n10181.n59 a_n2814_n10181.n58 3.1505
R1326 a_n2814_n10181.n10 a_n2814_n10181.n9 2.60819
R1327 a_n2814_n10181.n56 a_n2814_n10181.n55 2.60725
R1328 a_n2814_n10181.n53 a_n2814_n10181.n52 2.50614
R1329 a_n2814_n10181.n53 a_n2814_n10181.n11 2.30722
R1330 a_n2814_n10181.n49 a_n2814_n10181.n48 2.2505
R1331 a_n2814_n10181.n52 a_n2814_n10181.n49 1.62755
R1332 a_n2814_n10181.n58 a_n2814_n10181.n56 1.45274
R1333 a_n2814_n10181.n10 a_n2814_n10181.n7 1.44462
R1334 a_n2814_n10181.n54 a_n2814_n10181.n53 1.1178
R1335 a_n2814_n10181.n16 a_n2814_n10181.n15 0.9533
R1336 a_n2814_n10181.n16 a_n2814_n10181.n14 0.9527
R1337 a_n2814_n10181.n7 a_n2814_n10181.n6 0.863826
R1338 a_n2814_n10181.n58 a_n2814_n10181.n57 0.851587
R1339 a_n2814_n10181.n1 a_n2814_n10181.n0 0.800639
R1340 a_n2814_n10181.n47 a_n2814_n10181.n46 0.775661
R1341 a_n2814_n10181.n3 a_n2814_n10181.n2 0.768411
R1342 a_n2814_n10181.n59 a_n2814_n10181.t1 0.5465
R1343 a_n2814_n10181.t17 a_n2814_n10181.n59 0.5465
R1344 a_n2814_n10181.n18 a_n2814_n10181.t2 0.5465
R1345 a_n2814_n10181.n18 a_n2814_n10181.n17 0.5465
R1346 a_n2814_n10181.n51 a_n2814_n10181.t19 0.5465
R1347 a_n2814_n10181.n51 a_n2814_n10181.n50 0.5465
R1348 a_n2814_n10181.n9 a_n2814_n10181.t11 0.5465
R1349 a_n2814_n10181.n9 a_n2814_n10181.n8 0.5465
R1350 a_n2814_n10181.n5 a_n2814_n10181.t15 0.5465
R1351 a_n2814_n10181.n5 a_n2814_n10181.n4 0.5465
R1352 a_n2814_n10181.n55 a_n2814_n10181.t8 0.5465
R1353 a_n2814_n10181.n55 a_n2814_n10181.t13 0.5465
R1354 a_n2814_n10181.n11 a_n2814_n10181.n3 0.41197
R1355 a_n2814_n10181.n54 a_n2814_n10181.n1 0.405068
R1356 a_n2814_n10181.n56 a_n2814_n10181.n54 0.0331417
R1357 a_n2814_n10181.n11 a_n2814_n10181.n10 0.0315339
R1358 a_n3063_n8710.n54 a_n3063_n8710.t26 55.0215
R1359 a_n3063_n8710.n5 a_n3063_n8710.t30 55.0195
R1360 a_n3063_n8710.n32 a_n3063_n8710.t28 55.0161
R1361 a_n3063_n8710.n34 a_n3063_n8710.t24 55.0146
R1362 a_n3063_n8710.n14 a_n3063_n8710.t4 5.39224
R1363 a_n3063_n8710.n10 a_n3063_n8710.n9 5.38071
R1364 a_n3063_n8710.n11 a_n3063_n8710.n10 5.11785
R1365 a_n3063_n8710.n15 a_n3063_n8710.n14 5.06689
R1366 a_n3063_n8710.n10 a_n3063_n8710.t5 4.77202
R1367 a_n3063_n8710.n16 a_n3063_n8710.t1 4.77006
R1368 a_n3063_n8710.n14 a_n3063_n8710.n13 4.76049
R1369 a_n3063_n8710.n12 a_n3063_n8710.n7 4.44941
R1370 a_n3063_n8710.n18 a_n3063_n8710.n17 4.09252
R1371 a_n3063_n8710.n22 a_n3063_n8710.n21 3.4449
R1372 a_n3063_n8710.n0 a_n3063_n8710.n46 3.47423
R1373 a_n3063_n8710.n17 a_n3063_n8710.n12 2.6551
R1374 a_n3063_n8710.n39 a_n3063_n8710.n38 2.62158
R1375 a_n3063_n8710.n33 a_n3063_n8710.n31 2.62158
R1376 a_n3063_n8710.n36 a_n3063_n8710.n35 2.62146
R1377 a_n3063_n8710.n6 a_n3063_n8710.n4 2.6208
R1378 a_n3063_n8710.n51 a_n3063_n8710.n2 2.62078
R1379 a_n3063_n8710.n53 a_n3063_n8710.n52 2.62065
R1380 a_n3063_n8710.n17 a_n3063_n8710.n16 2.2505
R1381 a_n3063_n8710.n41 a_n3063_n8710.n40 2.2505
R1382 a_n3063_n8710.n50 a_n3063_n8710.n49 2.2505
R1383 a_n3063_n8710.n26 a_n3063_n8710.n25 2.2449
R1384 a_n3063_n8710.t27 a_n3063_n8710.n54 2.02927
R1385 a_n3063_n8710.n11 a_n3063_n8710.n8 1.89811
R1386 a_n3063_n8710.n15 a_n3063_n8710.t7 1.88742
R1387 a_n3063_n8710.n48 a_n3063_n8710.n0 1.50488
R1388 a_n3063_n8710.n0 a_n3063_n8710.n44 1.50096
R1389 a_n3063_n8710.n44 a_n3063_n8710.n43 1.49517
R1390 a_n3063_n8710.n25 a_n3063_n8710.n24 1.4938
R1391 a_n3063_n8710.n6 a_n3063_n8710.n5 1.34058
R1392 a_n3063_n8710.n33 a_n3063_n8710.n32 1.33904
R1393 a_n3063_n8710.n36 a_n3063_n8710.n34 1.33895
R1394 a_n3063_n8710.n12 a_n3063_n8710.n11 1.16362
R1395 a_n3063_n8710.n49 a_n3063_n8710.n48 1.15831
R1396 a_n3063_n8710.n29 a_n3063_n8710.n27 1.1218
R1397 a_n3063_n8710.n16 a_n3063_n8710.n15 0.881391
R1398 a_n3063_n8710.n39 a_n3063_n8710.n36 0.875886
R1399 a_n3063_n8710.n52 a_n3063_n8710.n51 0.875886
R1400 a_n3063_n8710.n49 a_n3063_n8710.n41 0.836663
R1401 a_n3063_n8710.n53 a_n3063_n8710.t12 0.5465
R1402 a_n3063_n8710.t27 a_n3063_n8710.n53 0.5465
R1403 a_n3063_n8710.n2 a_n3063_n8710.t9 0.5465
R1404 a_n3063_n8710.n2 a_n3063_n8710.n1 0.5465
R1405 a_n3063_n8710.n43 a_n3063_n8710.t11 0.5465
R1406 a_n3063_n8710.n43 a_n3063_n8710.n42 0.5465
R1407 a_n3063_n8710.n46 a_n3063_n8710.t13 0.5465
R1408 a_n3063_n8710.n46 a_n3063_n8710.n45 0.5465
R1409 a_n3063_n8710.n38 a_n3063_n8710.t8 0.5465
R1410 a_n3063_n8710.n38 a_n3063_n8710.n37 0.5465
R1411 a_n3063_n8710.n35 a_n3063_n8710.t10 0.5465
R1412 a_n3063_n8710.n35 a_n3063_n8710.t25 0.5465
R1413 a_n3063_n8710.n31 a_n3063_n8710.t29 0.5465
R1414 a_n3063_n8710.n31 a_n3063_n8710.n30 0.5465
R1415 a_n3063_n8710.n24 a_n3063_n8710.t15 0.5465
R1416 a_n3063_n8710.n24 a_n3063_n8710.n23 0.5465
R1417 a_n3063_n8710.n21 a_n3063_n8710.t14 0.5465
R1418 a_n3063_n8710.n21 a_n3063_n8710.n20 0.5465
R1419 a_n3063_n8710.n4 a_n3063_n8710.t31 0.5465
R1420 a_n3063_n8710.n4 a_n3063_n8710.n3 0.5465
R1421 a_n3063_n8710.n41 a_n3063_n8710.n29 0.499525
R1422 a_n3063_n8710.n40 a_n3063_n8710.n33 0.421979
R1423 a_n3063_n8710.n50 a_n3063_n8710.n6 0.421979
R1424 a_n3063_n8710.n40 a_n3063_n8710.n39 0.416316
R1425 a_n3063_n8710.n51 a_n3063_n8710.n50 0.416316
R1426 a_n3063_n8710.n26 a_n3063_n8710.n22 0.0180864
R1427 a_n3063_n8710.n19 a_n3063_n8710.n18 0.0171082
R1428 a_n3063_n8710.n27 a_n3063_n8710.n19 0.0141734
R1429 a_n3063_n8710.n27 a_n3063_n8710.n26 0.0131951
R1430 a_n3063_n8710.n48 a_n3063_n8710.n47 0.0114473
R1431 a_n3063_n8710.n29 a_n3063_n8710.n28 0.00965828
R1432 VSS.n197 VSS.t11 615.511
R1433 VSS.n472 VSS.t33 35.8214
R1434 VSS.n251 VSS.t10 32.0901
R1435 VSS.n459 VSS.t30 29.8512
R1436 VSS.n489 VSS.t28 28.3587
R1437 VSS.n267 VSS.t7 25.3736
R1438 VSS.n446 VSS.t9 23.8811
R1439 VSS.n282 VSS.t2 18.6572
R1440 VSS.n485 VSS.t43 17.9109
R1441 VSS.n462 VSS.t22 16.4184
R1442 VSS.t8 VSS.n257 15.6721
R1443 VSS.n469 VSS.t16 10.4483
R1444 VSS.n479 VSS.t37 8.95572
R1445 VSS.n288 VSS.t0 8.20945
R1446 VSS.n258 VSS.t8 5.22438
R1447 VSS.n198 VSS.n197 5.2005
R1448 VSS.n196 VSS.n195 4.86554
R1449 VSS.n199 VSS.n193 4.70124
R1450 VSS.n196 VSS.n194 4.69928
R1451 VSS.n89 VSS.n87 3.30147
R1452 VSS.n101 VSS.n99 3.30147
R1453 VSS.n101 VSS.n100 3.30091
R1454 VSS.n89 VSS.n88 3.30091
R1455 VSS.n340 VSS.n333 3.1505
R1456 VSS.n339 VSS.n335 3.1505
R1457 VSS.n338 VSS.n337 3.1505
R1458 VSS.n525 VSS.n524 3.1505
R1459 VSS.n349 VSS.n342 3.1505
R1460 VSS.n348 VSS.n344 3.1505
R1461 VSS.n347 VSS.n346 3.1505
R1462 VSS.n528 VSS.n527 3.1505
R1463 VSS.n358 VSS.n351 3.1505
R1464 VSS.n357 VSS.n353 3.1505
R1465 VSS.n356 VSS.n355 3.1505
R1466 VSS.n531 VSS.n530 3.1505
R1467 VSS.n331 VSS.n324 3.1505
R1468 VSS.n330 VSS.n326 3.1505
R1469 VSS.n329 VSS.n328 3.1505
R1470 VSS.n579 VSS.n578 3.1505
R1471 VSS.n452 VSS.t18 2.98557
R1472 VSS.n591 VSS.n522 2.60143
R1473 VSS.n504 VSS.n322 2.60143
R1474 VSS.n243 VSS.n242 2.6005
R1475 VSS.n192 VSS.n191 2.6005
R1476 VSS.n15 VSS.n14 2.6005
R1477 VSS.n13 VSS.n12 2.6005
R1478 VSS.n11 VSS.n10 2.6005
R1479 VSS.n9 VSS.n8 2.6005
R1480 VSS.n7 VSS.n6 2.6005
R1481 VSS.n5 VSS.n4 2.6005
R1482 VSS.n3 VSS.n2 2.6005
R1483 VSS.n1 VSS.n0 2.6005
R1484 VSS.n162 VSS.n161 2.6005
R1485 VSS.n164 VSS.n163 2.6005
R1486 VSS.n166 VSS.n165 2.6005
R1487 VSS.n168 VSS.n167 2.6005
R1488 VSS.n170 VSS.n169 2.6005
R1489 VSS.n172 VSS.n171 2.6005
R1490 VSS.n174 VSS.n173 2.6005
R1491 VSS.n176 VSS.n175 2.6005
R1492 VSS.n178 VSS.n177 2.6005
R1493 VSS.n180 VSS.n179 2.6005
R1494 VSS.n182 VSS.n181 2.6005
R1495 VSS.n184 VSS.n183 2.6005
R1496 VSS.n186 VSS.n185 2.6005
R1497 VSS.n188 VSS.n187 2.6005
R1498 VSS.n190 VSS.n189 2.6005
R1499 VSS.n201 VSS.n200 2.6005
R1500 VSS.n203 VSS.n202 2.6005
R1501 VSS.n205 VSS.n204 2.6005
R1502 VSS.n207 VSS.n206 2.6005
R1503 VSS.n209 VSS.n208 2.6005
R1504 VSS.n211 VSS.n210 2.6005
R1505 VSS.n214 VSS.n213 2.6005
R1506 VSS.n217 VSS.n216 2.6005
R1507 VSS.n220 VSS.n219 2.6005
R1508 VSS.n223 VSS.n222 2.6005
R1509 VSS.n226 VSS.n225 2.6005
R1510 VSS.n229 VSS.n228 2.6005
R1511 VSS.n232 VSS.n231 2.6005
R1512 VSS.n235 VSS.n234 2.6005
R1513 VSS.n238 VSS.n237 2.6005
R1514 VSS.n241 VSS.n240 2.6005
R1515 VSS.n651 VSS.n650 2.6005
R1516 VSS.n638 VSS.n637 2.6005
R1517 VSS.n541 VSS.n540 2.6005
R1518 VSS.n422 VSS.n421 2.6005
R1519 VSS.n420 VSS.n419 2.6005
R1520 VSS.n417 VSS.n416 2.6005
R1521 VSS.n415 VSS.n414 2.6005
R1522 VSS.n412 VSS.n411 2.6005
R1523 VSS.n410 VSS.n409 2.6005
R1524 VSS.n407 VSS.n406 2.6005
R1525 VSS.n405 VSS.n404 2.6005
R1526 VSS.n402 VSS.n401 2.6005
R1527 VSS.n400 VSS.n399 2.6005
R1528 VSS.n398 VSS.n397 2.6005
R1529 VSS.n396 VSS.n395 2.6005
R1530 VSS.n394 VSS.n393 2.6005
R1531 VSS.n392 VSS.n391 2.6005
R1532 VSS.n390 VSS.n389 2.6005
R1533 VSS.n388 VSS.n387 2.6005
R1534 VSS.n386 VSS.n385 2.6005
R1535 VSS.n384 VSS.n383 2.6005
R1536 VSS.n382 VSS.n381 2.6005
R1537 VSS.n380 VSS.n379 2.6005
R1538 VSS.n378 VSS.n377 2.6005
R1539 VSS.n376 VSS.n375 2.6005
R1540 VSS.n374 VSS.n373 2.6005
R1541 VSS.n372 VSS.n371 2.6005
R1542 VSS.n370 VSS.n369 2.6005
R1543 VSS.n368 VSS.n367 2.6005
R1544 VSS.n366 VSS.n365 2.6005
R1545 VSS.n364 VSS.n363 2.6005
R1546 VSS.n362 VSS.n361 2.6005
R1547 VSS.n360 VSS.n359 2.6005
R1548 VSS.n533 VSS.n532 2.6005
R1549 VSS.n535 VSS.n534 2.6005
R1550 VSS.n537 VSS.n536 2.6005
R1551 VSS.n539 VSS.n538 2.6005
R1552 VSS.n644 VSS.n643 2.6005
R1553 VSS.n646 VSS.n645 2.6005
R1554 VSS.n649 VSS.n648 2.6005
R1555 VSS.n641 VSS.n640 2.6005
R1556 VSS.n629 VSS.n628 2.6005
R1557 VSS.n631 VSS.n630 2.6005
R1558 VSS.n633 VSS.n632 2.6005
R1559 VSS.n636 VSS.n635 2.6005
R1560 VSS.n626 VSS.n625 2.6005
R1561 VSS.n623 VSS.n622 2.6005
R1562 VSS.n616 VSS.n615 2.6005
R1563 VSS.n618 VSS.n617 2.6005
R1564 VSS.n621 VSS.n620 2.6005
R1565 VSS.n614 VSS.n613 2.6005
R1566 VSS.n611 VSS.n610 2.6005
R1567 VSS.n605 VSS.n604 2.6005
R1568 VSS.n607 VSS.n606 2.6005
R1569 VSS.n609 VSS.n608 2.6005
R1570 VSS.n603 VSS.n602 2.6005
R1571 VSS.n600 VSS.n599 2.6005
R1572 VSS.n596 VSS.n595 2.6005
R1573 VSS.n598 VSS.n597 2.6005
R1574 VSS.n594 VSS.n593 2.6005
R1575 VSS.n244 VSS.n160 2.6005
R1576 VSS.n247 VSS.n246 2.6005
R1577 VSS.n246 VSS.n245 2.6005
R1578 VSS.n250 VSS.n249 2.6005
R1579 VSS.n249 VSS.n248 2.6005
R1580 VSS.n253 VSS.n252 2.6005
R1581 VSS.n252 VSS.n251 2.6005
R1582 VSS.n256 VSS.n255 2.6005
R1583 VSS.n255 VSS.n254 2.6005
R1584 VSS.n260 VSS.n259 2.6005
R1585 VSS.n259 VSS.n258 2.6005
R1586 VSS.n263 VSS.n262 2.6005
R1587 VSS.n262 VSS.n261 2.6005
R1588 VSS.n266 VSS.n265 2.6005
R1589 VSS.n265 VSS.n264 2.6005
R1590 VSS.n269 VSS.n268 2.6005
R1591 VSS.n268 VSS.n267 2.6005
R1592 VSS.n272 VSS.n271 2.6005
R1593 VSS.n271 VSS.n270 2.6005
R1594 VSS.n275 VSS.n274 2.6005
R1595 VSS.n274 VSS.n273 2.6005
R1596 VSS.n278 VSS.n277 2.6005
R1597 VSS.n277 VSS.n276 2.6005
R1598 VSS.n281 VSS.n280 2.6005
R1599 VSS.n280 VSS.n279 2.6005
R1600 VSS.n284 VSS.n283 2.6005
R1601 VSS.n283 VSS.n282 2.6005
R1602 VSS.n287 VSS.n286 2.6005
R1603 VSS.n286 VSS.n285 2.6005
R1604 VSS.n290 VSS.n289 2.6005
R1605 VSS.n289 VSS.n288 2.6005
R1606 VSS.n293 VSS.n292 2.6005
R1607 VSS.n292 VSS.n291 2.6005
R1608 VSS.n296 VSS.n295 2.6005
R1609 VSS.n295 VSS.n294 2.6005
R1610 VSS.n298 VSS.n297 2.6005
R1611 VSS.n53 VSS.n52 2.6005
R1612 VSS.n19 VSS.n18 2.6005
R1613 VSS.n21 VSS.n20 2.6005
R1614 VSS.n23 VSS.n22 2.6005
R1615 VSS.n25 VSS.n24 2.6005
R1616 VSS.n27 VSS.n26 2.6005
R1617 VSS.n29 VSS.n28 2.6005
R1618 VSS.n31 VSS.n30 2.6005
R1619 VSS.n33 VSS.n32 2.6005
R1620 VSS.n35 VSS.n34 2.6005
R1621 VSS.n37 VSS.n36 2.6005
R1622 VSS.n39 VSS.n38 2.6005
R1623 VSS.n41 VSS.n40 2.6005
R1624 VSS.n43 VSS.n42 2.6005
R1625 VSS.n45 VSS.n44 2.6005
R1626 VSS.n47 VSS.n46 2.6005
R1627 VSS.n49 VSS.n48 2.6005
R1628 VSS.n51 VSS.n50 2.6005
R1629 VSS.n17 VSS.n16 2.6005
R1630 VSS.n63 VSS.n62 2.6005
R1631 VSS.n73 VSS.n72 2.6005
R1632 VSS.n82 VSS.n81 2.6005
R1633 VSS.n92 VSS.n91 2.6005
R1634 VSS.n104 VSS.n103 2.6005
R1635 VSS.n115 VSS.n114 2.6005
R1636 VSS.n303 VSS.n302 2.6005
R1637 VSS.n306 VSS.n305 2.6005
R1638 VSS.n308 VSS.n307 2.6005
R1639 VSS.n128 VSS.n127 2.6005
R1640 VSS.n125 VSS.n124 2.6005
R1641 VSS.n123 VSS.n122 2.6005
R1642 VSS.n120 VSS.n119 2.6005
R1643 VSS.n118 VSS.n117 2.6005
R1644 VSS.n113 VSS.n111 2.6005
R1645 VSS.n113 VSS.n112 2.6005
R1646 VSS.n109 VSS.n108 2.6005
R1647 VSS.n106 VSS.n105 2.6005
R1648 VSS.n98 VSS.n97 2.6005
R1649 VSS.n96 VSS.n95 2.6005
R1650 VSS.n94 VSS.n93 2.6005
R1651 VSS.n86 VSS.n85 2.6005
R1652 VSS.n84 VSS.n83 2.6005
R1653 VSS.n80 VSS.n78 2.6005
R1654 VSS.n80 VSS.n79 2.6005
R1655 VSS.n77 VSS.n76 2.6005
R1656 VSS.n75 VSS.n74 2.6005
R1657 VSS.n71 VSS.n70 2.6005
R1658 VSS.n69 VSS.n68 2.6005
R1659 VSS.n67 VSS.n66 2.6005
R1660 VSS.n65 VSS.n64 2.6005
R1661 VSS.n59 VSS.n58 2.6005
R1662 VSS.n57 VSS.n56 2.6005
R1663 VSS.n55 VSS.n54 2.6005
R1664 VSS.n301 VSS.n300 2.6005
R1665 VSS.n61 VSS.n60 2.6005
R1666 VSS.n590 VSS.n589 2.6005
R1667 VSS.n588 VSS.n587 2.6005
R1668 VSS.n586 VSS.n585 2.6005
R1669 VSS.n584 VSS.n583 2.6005
R1670 VSS.n582 VSS.n581 2.6005
R1671 VSS.n576 VSS.n575 2.6005
R1672 VSS.n574 VSS.n573 2.6005
R1673 VSS.n572 VSS.n571 2.6005
R1674 VSS.n569 VSS.n568 2.6005
R1675 VSS.n567 VSS.n566 2.6005
R1676 VSS.n565 VSS.n564 2.6005
R1677 VSS.n562 VSS.n561 2.6005
R1678 VSS.n560 VSS.n559 2.6005
R1679 VSS.n558 VSS.n557 2.6005
R1680 VSS.n556 VSS.n555 2.6005
R1681 VSS.n553 VSS.n552 2.6005
R1682 VSS.n551 VSS.n550 2.6005
R1683 VSS.n549 VSS.n548 2.6005
R1684 VSS.n547 VSS.n546 2.6005
R1685 VSS.n545 VSS.n544 2.6005
R1686 VSS.n543 VSS.n542 2.6005
R1687 VSS.n503 VSS.n502 2.6005
R1688 VSS.n502 VSS.n501 2.6005
R1689 VSS.n500 VSS.n499 2.6005
R1690 VSS.n499 VSS.n498 2.6005
R1691 VSS.n497 VSS.n496 2.6005
R1692 VSS.n496 VSS.n495 2.6005
R1693 VSS.n494 VSS.n493 2.6005
R1694 VSS.n493 VSS.n492 2.6005
R1695 VSS.n491 VSS.n490 2.6005
R1696 VSS.n490 VSS.n489 2.6005
R1697 VSS.n487 VSS.n486 2.6005
R1698 VSS.n486 VSS.n485 2.6005
R1699 VSS.n484 VSS.n483 2.6005
R1700 VSS.n483 VSS.n482 2.6005
R1701 VSS.n481 VSS.n480 2.6005
R1702 VSS.n480 VSS.n479 2.6005
R1703 VSS.n477 VSS.n476 2.6005
R1704 VSS.n476 VSS.n475 2.6005
R1705 VSS.n474 VSS.n473 2.6005
R1706 VSS.n473 VSS.n472 2.6005
R1707 VSS.n471 VSS.n470 2.6005
R1708 VSS.n470 VSS.n469 2.6005
R1709 VSS.n467 VSS.n466 2.6005
R1710 VSS.n466 VSS.n465 2.6005
R1711 VSS.n464 VSS.n463 2.6005
R1712 VSS.n463 VSS.n462 2.6005
R1713 VSS.n461 VSS.n460 2.6005
R1714 VSS.n460 VSS.n459 2.6005
R1715 VSS.n458 VSS.n457 2.6005
R1716 VSS.n457 VSS.n456 2.6005
R1717 VSS.n454 VSS.n453 2.6005
R1718 VSS.n453 VSS.n452 2.6005
R1719 VSS.n451 VSS.n450 2.6005
R1720 VSS.n450 VSS.n449 2.6005
R1721 VSS.n448 VSS.n447 2.6005
R1722 VSS.n447 VSS.n446 2.6005
R1723 VSS.n445 VSS.n444 2.6005
R1724 VSS.n444 VSS.n443 2.6005
R1725 VSS.n442 VSS.n441 2.6005
R1726 VSS.n441 VSS.n440 2.6005
R1727 VSS.n439 VSS.n438 2.6005
R1728 VSS.n519 VSS.n518 2.6005
R1729 VSS.n657 VSS.n656 2.6005
R1730 VSS.n660 VSS.n659 2.6005
R1731 VSS.n662 VSS.n661 2.6005
R1732 VSS.n665 VSS.n664 2.6005
R1733 VSS.n667 VSS.n666 2.6005
R1734 VSS.n655 VSS.n654 2.6005
R1735 VSS.n321 VSS.n320 2.6005
R1736 VSS.n671 VSS.n670 2.6005
R1737 VSS.n237 VSS.n236 2.41715
R1738 VSS.n234 VSS.n233 2.41715
R1739 VSS.n231 VSS.n230 2.41715
R1740 VSS.n228 VSS.n227 2.41715
R1741 VSS.n225 VSS.n224 2.41715
R1742 VSS.n222 VSS.n221 2.41715
R1743 VSS.n219 VSS.n218 2.41715
R1744 VSS.n216 VSS.n215 2.41715
R1745 VSS.n213 VSS.n212 2.41715
R1746 VSS.n201 VSS.n199 1.73826
R1747 VSS.n419 VSS.n418 1.65132
R1748 VSS.n414 VSS.n413 1.65132
R1749 VSS.n409 VSS.n408 1.65132
R1750 VSS.n404 VSS.n403 1.65132
R1751 VSS.n654 VSS.n653 1.65076
R1752 VSS.n127 VSS.n126 1.65065
R1753 VSS.n122 VSS.n121 1.65065
R1754 VSS.n117 VSS.n116 1.65065
R1755 VSS.n111 VSS.n110 1.65065
R1756 VSS.n108 VSS.n107 1.65065
R1757 VSS.n305 VSS.n304 1.65065
R1758 VSS.n659 VSS.n658 1.65065
R1759 VSS.n664 VSS.n663 1.65065
R1760 VSS.n320 VSS.n319 1.65065
R1761 VSS.n670 VSS.n669 1.65065
R1762 VSS.n273 VSS.t1 1.49304
R1763 VSS.n495 VSS.t6 1.49304
R1764 VSS.n340 VSS.n339 1.4405
R1765 VSS.n349 VSS.n348 1.4405
R1766 VSS.n358 VSS.n357 1.4405
R1767 VSS.n331 VSS.n330 1.4405
R1768 VSS.n339 VSS.n338 1.4369
R1769 VSS.n348 VSS.n347 1.4369
R1770 VSS.n357 VSS.n356 1.4369
R1771 VSS.n330 VSS.n329 1.4369
R1772 VSS.n240 VSS.n239 1.39588
R1773 VSS.n648 VSS.n647 1.39588
R1774 VSS.n635 VSS.n634 1.39588
R1775 VSS.n620 VSS.n619 1.39588
R1776 VSS.n643 VSS.n642 1.39574
R1777 VSS.n628 VSS.n627 1.39574
R1778 VSS.n158 VSS.n130 1.39293
R1779 VSS.n158 VSS.n131 1.39293
R1780 VSS.n158 VSS.n132 1.39293
R1781 VSS.n158 VSS.n133 1.39293
R1782 VSS.n158 VSS.n134 1.39293
R1783 VSS.n158 VSS.n135 1.39293
R1784 VSS.n158 VSS.n136 1.39293
R1785 VSS.n158 VSS.n137 1.39293
R1786 VSS.n158 VSS.n138 1.39293
R1787 VSS.n158 VSS.n139 1.39293
R1788 VSS.n158 VSS.n140 1.39293
R1789 VSS.n158 VSS.n141 1.39293
R1790 VSS.n158 VSS.n142 1.39293
R1791 VSS.n158 VSS.n143 1.39293
R1792 VSS.n158 VSS.n144 1.39293
R1793 VSS.n158 VSS.n145 1.39293
R1794 VSS.n158 VSS.n146 1.39293
R1795 VSS.n158 VSS.n147 1.39293
R1796 VSS.n158 VSS.n148 1.39293
R1797 VSS.n158 VSS.n149 1.39293
R1798 VSS.n158 VSS.n150 1.39293
R1799 VSS.n158 VSS.n151 1.39293
R1800 VSS.n158 VSS.n152 1.39293
R1801 VSS.n158 VSS.n153 1.39293
R1802 VSS.n158 VSS.n154 1.39293
R1803 VSS.n158 VSS.n155 1.39293
R1804 VSS.n158 VSS.n156 1.39293
R1805 VSS.n158 VSS.n157 1.39293
R1806 VSS.n516 VSS.n514 1.39293
R1807 VSS.n160 VSS.n159 1.34121
R1808 VSS.n438 VSS.n437 1.3407
R1809 VSS.n518 VSS.n517 1.3407
R1810 VSS.n300 VSS.n299 1.34055
R1811 VSS.t11 VSS.t3 1.25921
R1812 VSS.n478 VSS.n340 0.9455
R1813 VSS.n468 VSS.n349 0.9455
R1814 VSS.n455 VSS.n358 0.9455
R1815 VSS.n488 VSS.n331 0.9455
R1816 VSS.n570 VSS.n525 0.9131
R1817 VSS.n563 VSS.n528 0.9131
R1818 VSS.n554 VSS.n531 0.9131
R1819 VSS.n580 VSS.n579 0.9131
R1820 VSS.n516 VSS.n510 0.804703
R1821 VSS.n158 VSS.n129 0.804503
R1822 VSS.n516 VSS.n512 0.804503
R1823 VSS.n516 VSS.n509 0.804503
R1824 VSS.n159 VSS.n158 0.631461
R1825 VSS.n516 VSS.n505 0.631461
R1826 VSS.n437 VSS.n436 0.631461
R1827 VSS.n517 VSS.n516 0.631461
R1828 VSS.n578 VSS.t65 0.5465
R1829 VSS.n578 VSS.n577 0.5465
R1830 VSS.n328 VSS.t36 0.5465
R1831 VSS.n328 VSS.n327 0.5465
R1832 VSS.n326 VSS.t29 0.5465
R1833 VSS.n326 VSS.n325 0.5465
R1834 VSS.n324 VSS.t61 0.5465
R1835 VSS.n324 VSS.n323 0.5465
R1836 VSS.n524 VSS.t62 0.5465
R1837 VSS.n524 VSS.n523 0.5465
R1838 VSS.n337 VSS.t64 0.5465
R1839 VSS.n337 VSS.n336 0.5465
R1840 VSS.n335 VSS.t60 0.5465
R1841 VSS.n335 VSS.n334 0.5465
R1842 VSS.n333 VSS.t38 0.5465
R1843 VSS.n333 VSS.n332 0.5465
R1844 VSS.n527 VSS.t17 0.5465
R1845 VSS.n527 VSS.n526 0.5465
R1846 VSS.n346 VSS.t55 0.5465
R1847 VSS.n346 VSS.n345 0.5465
R1848 VSS.n344 VSS.t48 0.5465
R1849 VSS.n344 VSS.n343 0.5465
R1850 VSS.n342 VSS.t25 0.5465
R1851 VSS.n342 VSS.n341 0.5465
R1852 VSS.n530 VSS.t32 0.5465
R1853 VSS.n530 VSS.n529 0.5465
R1854 VSS.n355 VSS.t39 0.5465
R1855 VSS.n355 VSS.n354 0.5465
R1856 VSS.n353 VSS.t31 0.5465
R1857 VSS.n353 VSS.n352 0.5465
R1858 VSS.n351 VSS.t63 0.5465
R1859 VSS.n351 VSS.n350 0.5465
R1860 VSS.n436 VSS.n435 0.476417
R1861 VSS.n436 VSS.n434 0.476417
R1862 VSS.n436 VSS.n433 0.476417
R1863 VSS.n436 VSS.n432 0.476417
R1864 VSS.n436 VSS.n431 0.476417
R1865 VSS.n436 VSS.n430 0.476417
R1866 VSS.n436 VSS.n429 0.476417
R1867 VSS.n436 VSS.n428 0.476417
R1868 VSS.n436 VSS.n427 0.476417
R1869 VSS.n436 VSS.n426 0.476417
R1870 VSS.n436 VSS.n425 0.476417
R1871 VSS.n436 VSS.n424 0.476417
R1872 VSS.n436 VSS.n423 0.476417
R1873 VSS.n516 VSS.n515 0.476417
R1874 VSS.n516 VSS.n513 0.476417
R1875 VSS.n516 VSS.n511 0.476417
R1876 VSS.n516 VSS.n508 0.476417
R1877 VSS.n516 VSS.n507 0.476417
R1878 VSS.n102 VSS.n101 0.476417
R1879 VSS.n90 VSS.n89 0.476417
R1880 VSS.n521 VSS.n520 0.476417
R1881 VSS.n516 VSS.n506 0.476417
R1882 VSS.n318 VSS.n317 0.476176
R1883 VSS.n318 VSS.n315 0.476176
R1884 VSS.n318 VSS.n314 0.476176
R1885 VSS.n318 VSS.n313 0.476176
R1886 VSS.n318 VSS.n312 0.476176
R1887 VSS.n318 VSS.n311 0.476176
R1888 VSS.n318 VSS.n310 0.476176
R1889 VSS.n318 VSS.n309 0.476176
R1890 VSS.n319 VSS.n318 0.476176
R1891 VSS.n318 VSS.n316 0.476176
R1892 VSS VSS.n321 0.263861
R1893 VSS VSS.n671 0.24468
R1894 VSS.n199 VSS.n198 0.119223
R1895 VSS.n128 VSS.n125 0.0914278
R1896 VSS.n125 VSS.n123 0.0914278
R1897 VSS.n123 VSS.n120 0.0914278
R1898 VSS.n120 VSS.n118 0.0914278
R1899 VSS.n118 VSS.n115 0.0914278
R1900 VSS.n113 VSS.n109 0.0914278
R1901 VSS.n109 VSS.n106 0.0914278
R1902 VSS.n106 VSS.n104 0.0914278
R1903 VSS.n98 VSS.n96 0.0914278
R1904 VSS.n96 VSS.n94 0.0914278
R1905 VSS.n94 VSS.n92 0.0914278
R1906 VSS.n86 VSS.n84 0.0914278
R1907 VSS.n84 VSS.n82 0.0914278
R1908 VSS.n77 VSS.n75 0.0914278
R1909 VSS.n75 VSS.n73 0.0914278
R1910 VSS.n69 VSS.n67 0.0914278
R1911 VSS.n67 VSS.n65 0.0914278
R1912 VSS.n65 VSS.n63 0.0914278
R1913 VSS.n303 VSS.n301 0.0914278
R1914 VSS.n306 VSS.n303 0.0914278
R1915 VSS.n308 VSS.n306 0.0914278
R1916 VSS.n422 VSS.n420 0.0914278
R1917 VSS.n420 VSS.n417 0.0914278
R1918 VSS.n417 VSS.n415 0.0914278
R1919 VSS.n415 VSS.n412 0.0914278
R1920 VSS.n412 VSS.n410 0.0914278
R1921 VSS.n410 VSS.n407 0.0914278
R1922 VSS.n407 VSS.n405 0.0914278
R1923 VSS.n405 VSS.n402 0.0914278
R1924 VSS.n402 VSS.n400 0.0914278
R1925 VSS.n400 VSS.n398 0.0914278
R1926 VSS.n398 VSS.n396 0.0914278
R1927 VSS.n396 VSS.n394 0.0914278
R1928 VSS.n394 VSS.n392 0.0914278
R1929 VSS.n392 VSS.n390 0.0914278
R1930 VSS.n390 VSS.n388 0.0914278
R1931 VSS.n388 VSS.n386 0.0914278
R1932 VSS.n386 VSS.n384 0.0914278
R1933 VSS.n384 VSS.n382 0.0914278
R1934 VSS.n382 VSS.n380 0.0914278
R1935 VSS.n380 VSS.n378 0.0914278
R1936 VSS.n378 VSS.n376 0.0914278
R1937 VSS.n376 VSS.n374 0.0914278
R1938 VSS.n374 VSS.n372 0.0914278
R1939 VSS.n372 VSS.n370 0.0914278
R1940 VSS.n370 VSS.n368 0.0914278
R1941 VSS.n368 VSS.n366 0.0914278
R1942 VSS.n366 VSS.n364 0.0914278
R1943 VSS.n364 VSS.n362 0.0914278
R1944 VSS.n362 VSS.n360 0.0914278
R1945 VSS.n535 VSS.n533 0.0914278
R1946 VSS.n537 VSS.n535 0.0914278
R1947 VSS.n539 VSS.n537 0.0914278
R1948 VSS.n541 VSS.n539 0.0914278
R1949 VSS.n598 VSS.n596 0.0914278
R1950 VSS.n596 VSS.n594 0.0914278
R1951 VSS.n609 VSS.n607 0.0914278
R1952 VSS.n607 VSS.n605 0.0914278
R1953 VSS.n605 VSS.n603 0.0914278
R1954 VSS.n621 VSS.n618 0.0914278
R1955 VSS.n618 VSS.n616 0.0914278
R1956 VSS.n616 VSS.n614 0.0914278
R1957 VSS.n649 VSS.n646 0.0914278
R1958 VSS.n646 VSS.n644 0.0914278
R1959 VSS.n644 VSS.n641 0.0914278
R1960 VSS.n636 VSS.n633 0.0914278
R1961 VSS.n633 VSS.n631 0.0914278
R1962 VSS.n631 VSS.n629 0.0914278
R1963 VSS.n629 VSS.n626 0.0914278
R1964 VSS.n192 VSS.n190 0.0914278
R1965 VSS.n190 VSS.n188 0.0914278
R1966 VSS.n188 VSS.n186 0.0914278
R1967 VSS.n186 VSS.n184 0.0914278
R1968 VSS.n184 VSS.n182 0.0914278
R1969 VSS.n182 VSS.n180 0.0914278
R1970 VSS.n180 VSS.n178 0.0914278
R1971 VSS.n178 VSS.n176 0.0914278
R1972 VSS.n176 VSS.n174 0.0914278
R1973 VSS.n174 VSS.n172 0.0914278
R1974 VSS.n172 VSS.n170 0.0914278
R1975 VSS.n170 VSS.n168 0.0914278
R1976 VSS.n168 VSS.n166 0.0914278
R1977 VSS.n166 VSS.n164 0.0914278
R1978 VSS.n164 VSS.n162 0.0914278
R1979 VSS.n3 VSS.n1 0.0914278
R1980 VSS.n5 VSS.n3 0.0914278
R1981 VSS.n7 VSS.n5 0.0914278
R1982 VSS.n9 VSS.n7 0.0914278
R1983 VSS.n11 VSS.n9 0.0914278
R1984 VSS.n13 VSS.n11 0.0914278
R1985 VSS.n15 VSS.n13 0.0914278
R1986 VSS.n247 VSS.n244 0.0914278
R1987 VSS.n250 VSS.n247 0.0914278
R1988 VSS.n253 VSS.n250 0.0914278
R1989 VSS.n256 VSS.n253 0.0914278
R1990 VSS.n260 VSS.n256 0.0914278
R1991 VSS.n263 VSS.n260 0.0914278
R1992 VSS.n266 VSS.n263 0.0914278
R1993 VSS.n269 VSS.n266 0.0914278
R1994 VSS.n272 VSS.n269 0.0914278
R1995 VSS.n275 VSS.n272 0.0914278
R1996 VSS.n278 VSS.n275 0.0914278
R1997 VSS.n281 VSS.n278 0.0914278
R1998 VSS.n284 VSS.n281 0.0914278
R1999 VSS.n287 VSS.n284 0.0914278
R2000 VSS.n290 VSS.n287 0.0914278
R2001 VSS.n293 VSS.n290 0.0914278
R2002 VSS.n296 VSS.n293 0.0914278
R2003 VSS.n298 VSS.n296 0.0914278
R2004 VSS.n243 VSS.n241 0.0914278
R2005 VSS.n241 VSS.n238 0.0914278
R2006 VSS.n238 VSS.n235 0.0914278
R2007 VSS.n235 VSS.n232 0.0914278
R2008 VSS.n232 VSS.n229 0.0914278
R2009 VSS.n229 VSS.n226 0.0914278
R2010 VSS.n226 VSS.n223 0.0914278
R2011 VSS.n223 VSS.n220 0.0914278
R2012 VSS.n220 VSS.n217 0.0914278
R2013 VSS.n217 VSS.n214 0.0914278
R2014 VSS.n214 VSS.n211 0.0914278
R2015 VSS.n211 VSS.n209 0.0914278
R2016 VSS.n209 VSS.n207 0.0914278
R2017 VSS.n207 VSS.n205 0.0914278
R2018 VSS.n205 VSS.n203 0.0914278
R2019 VSS.n59 VSS.n57 0.0914278
R2020 VSS.n57 VSS.n55 0.0914278
R2021 VSS.n19 VSS.n17 0.0914278
R2022 VSS.n21 VSS.n19 0.0914278
R2023 VSS.n23 VSS.n21 0.0914278
R2024 VSS.n25 VSS.n23 0.0914278
R2025 VSS.n27 VSS.n25 0.0914278
R2026 VSS.n29 VSS.n27 0.0914278
R2027 VSS.n31 VSS.n29 0.0914278
R2028 VSS.n33 VSS.n31 0.0914278
R2029 VSS.n35 VSS.n33 0.0914278
R2030 VSS.n37 VSS.n35 0.0914278
R2031 VSS.n39 VSS.n37 0.0914278
R2032 VSS.n41 VSS.n39 0.0914278
R2033 VSS.n43 VSS.n41 0.0914278
R2034 VSS.n45 VSS.n43 0.0914278
R2035 VSS.n47 VSS.n45 0.0914278
R2036 VSS.n49 VSS.n47 0.0914278
R2037 VSS.n51 VSS.n49 0.0914278
R2038 VSS.n53 VSS.n51 0.0914278
R2039 VSS.n590 VSS.n588 0.0914278
R2040 VSS.n588 VSS.n586 0.0914278
R2041 VSS.n586 VSS.n584 0.0914278
R2042 VSS.n584 VSS.n582 0.0914278
R2043 VSS.n576 VSS.n574 0.0914278
R2044 VSS.n574 VSS.n572 0.0914278
R2045 VSS.n569 VSS.n567 0.0914278
R2046 VSS.n567 VSS.n565 0.0914278
R2047 VSS.n562 VSS.n560 0.0914278
R2048 VSS.n560 VSS.n558 0.0914278
R2049 VSS.n558 VSS.n556 0.0914278
R2050 VSS.n553 VSS.n551 0.0914278
R2051 VSS.n551 VSS.n549 0.0914278
R2052 VSS.n549 VSS.n547 0.0914278
R2053 VSS.n547 VSS.n545 0.0914278
R2054 VSS.n545 VSS.n543 0.0914278
R2055 VSS.n503 VSS.n500 0.0914278
R2056 VSS.n500 VSS.n497 0.0914278
R2057 VSS.n497 VSS.n494 0.0914278
R2058 VSS.n494 VSS.n491 0.0914278
R2059 VSS.n487 VSS.n484 0.0914278
R2060 VSS.n484 VSS.n481 0.0914278
R2061 VSS.n477 VSS.n474 0.0914278
R2062 VSS.n474 VSS.n471 0.0914278
R2063 VSS.n467 VSS.n464 0.0914278
R2064 VSS.n464 VSS.n461 0.0914278
R2065 VSS.n461 VSS.n458 0.0914278
R2066 VSS.n454 VSS.n451 0.0914278
R2067 VSS.n451 VSS.n448 0.0914278
R2068 VSS.n448 VSS.n445 0.0914278
R2069 VSS.n445 VSS.n442 0.0914278
R2070 VSS.n442 VSS.n439 0.0914278
R2071 VSS.n667 VSS.n665 0.0914278
R2072 VSS.n665 VSS.n662 0.0914278
R2073 VSS.n662 VSS.n660 0.0914278
R2074 VSS.n660 VSS.n657 0.0914278
R2075 VSS.n657 VSS.n655 0.0914278
R2076 VSS.n591 VSS.n590 0.0905
R2077 VSS.n504 VSS.n503 0.0905
R2078 VSS.n92 VSS.n90 0.0895722
R2079 VSS.n565 VSS.n563 0.0877165
R2080 VSS.n471 VSS.n468 0.0877165
R2081 VSS.n594 VSS.n592 0.0858608
R2082 VSS.n82 VSS.n80 0.0830773
R2083 VSS.n104 VSS.n102 0.0821495
R2084 VSS.n102 VSS.n98 0.0784381
R2085 VSS.n80 VSS.n77 0.0775103
R2086 VSS.n90 VSS.n86 0.0710155
R2087 VSS.n554 VSS.n553 0.0710155
R2088 VSS.n455 VSS.n454 0.0710155
R2089 VSS.n115 VSS.n113 0.0691598
R2090 VSS.n73 VSS.n71 0.068232
R2091 VSS.n572 VSS.n570 0.0635928
R2092 VSS.n481 VSS.n478 0.0635928
R2093 VSS.n626 VSS.n624 0.0561701
R2094 VSS.n203 VSS.n201 0.0533866
R2095 VSS.n580 VSS.n576 0.0524588
R2096 VSS.n488 VSS.n487 0.0524588
R2097 VSS.n198 VSS.n196 0.0518191
R2098 VSS.n321 VSS.n308 0.0515309
R2099 VSS.n668 VSS.n667 0.0515309
R2100 VSS.n614 VSS.n612 0.0496753
R2101 VSS.n641 VSS.n639 0.0487474
R2102 VSS.n301 VSS.n298 0.0459639
R2103 VSS.n439 VSS.n422 0.0459639
R2104 VSS.n543 VSS.n541 0.0459639
R2105 VSS.n17 VSS.n15 0.0459639
R2106 VSS.n244 VSS.n243 0.0459639
R2107 VSS.n55 VSS.n53 0.0459639
R2108 VSS.n519 VSS.n504 0.0459639
R2109 VSS.n61 VSS.n59 0.0413247
R2110 VSS.n582 VSS.n580 0.0394691
R2111 VSS.n491 VSS.n488 0.0394691
R2112 VSS.n655 VSS.n652 0.0357577
R2113 VSS.n601 VSS.n598 0.0348299
R2114 VSS.n603 VSS.n601 0.0348299
R2115 VSS.n652 VSS.n649 0.0339021
R2116 VSS.n201 VSS.n192 0.0339021
R2117 VSS.n592 VSS.n591 0.0292629
R2118 VSS.n63 VSS.n61 0.0283351
R2119 VSS.n570 VSS.n569 0.0283351
R2120 VSS.n478 VSS.n477 0.0283351
R2121 VSS.n639 VSS.n636 0.0209124
R2122 VSS.n556 VSS.n554 0.0209124
R2123 VSS.n458 VSS.n455 0.0209124
R2124 VSS.n612 VSS.n609 0.0199845
R2125 VSS.n321 VSS.n128 0.0181289
R2126 VSS.n668 VSS.n519 0.0181289
R2127 VSS.n624 VSS.n621 0.0134897
R2128 VSS.n563 VSS.n562 0.00421134
R2129 VSS.n468 VSS.n467 0.00421134
R2130 VSS.n71 VSS.n69 0.00142783
R2131 VSS.n601 VSS.n600 0.0012377
R2132 VSS.n612 VSS.n611 0.0012377
R2133 VSS.n624 VSS.n623 0.0012377
R2134 VSS.n639 VSS.n638 0.0012377
R2135 VSS.n652 VSS.n651 0.0012377
R2136 VSS.n592 VSS.n521 0.0012377
R2137 VSS.n671 VSS.n668 0.0012377
R2138 OUT.n24 OUT.t24 55.2511
R2139 OUT.n14 OUT.t10 53.6484
R2140 OUT.n26 OUT.t20 52.4934
R2141 OUT.n12 OUT.t22 51.4031
R2142 OUT.n33 OUT.t16 50.0561
R2143 OUT.n3 OUT.t12 49.577
R2144 OUT.n3 OUT.t14 48.7525
R2145 OUT.n33 OUT.t18 48.2735
R2146 OUT.n30 OUT.n18 5.49154
R2147 OUT.n29 OUT.n20 5.48524
R2148 OUT.n29 OUT.n28 4.52226
R2149 OUT.n39 OUT.n31 4.38577
R2150 OUT.n35 OUT.n33 4.0005
R2151 OUT.n4 OUT.n3 4.0005
R2152 OUT.n25 OUT.n23 3.86659
R2153 OUT.n13 OUT.n11 3.83724
R2154 OUT.n31 OUT.n16 3.3987
R2155 OUT.n5 OUT.n1 3.2449
R2156 OUT.n36 OUT.n32 3.2377
R2157 OUT.n38 OUT.n37 2.6005
R2158 OUT.n8 OUT.n7 2.6005
R2159 OUT.n15 OUT.n13 2.32876
R2160 OUT.n27 OUT.n25 2.31115
R2161 OUT.n16 OUT.n9 1.48952
R2162 OUT.n28 OUT.n21 1.44997
R2163 OUT OUT.n8 1.2011
R2164 OUT.n31 OUT.n30 1.19168
R2165 OUT.n30 OUT.n29 1.18495
R2166 OUT.n39 OUT.n38 1.12137
R2167 OUT OUT.n39 1.01517
R2168 OUT.n38 OUT.n36 0.6611
R2169 OUT.n8 OUT.n5 0.6539
R2170 OUT.n37 OUT.t0 0.607167
R2171 OUT.n37 OUT.t17 0.607167
R2172 OUT.n32 OUT.t2 0.607167
R2173 OUT.n32 OUT.t19 0.607167
R2174 OUT.n7 OUT.t13 0.607167
R2175 OUT.n7 OUT.n6 0.607167
R2176 OUT.n1 OUT.t15 0.607167
R2177 OUT.n1 OUT.n0 0.607167
R2178 OUT.n11 OUT.t23 0.5465
R2179 OUT.n11 OUT.n10 0.5465
R2180 OUT.n9 OUT.t4 0.5465
R2181 OUT.n9 OUT.t11 0.5465
R2182 OUT.n18 OUT.t1 0.5465
R2183 OUT.n18 OUT.n17 0.5465
R2184 OUT.n20 OUT.t9 0.5465
R2185 OUT.n20 OUT.n19 0.5465
R2186 OUT.n21 OUT.t5 0.5465
R2187 OUT.n21 OUT.t21 0.5465
R2188 OUT.n23 OUT.t25 0.5465
R2189 OUT.n23 OUT.n22 0.5465
R2190 OUT.n28 OUT.n27 0.389832
R2191 OUT.n16 OUT.n15 0.28107
R2192 OUT.n25 OUT.n24 0.277411
R2193 OUT.n27 OUT.n26 0.160935
R2194 OUT.n15 OUT.n14 0.158978
R2195 OUT.n13 OUT.n12 0.157022
R2196 OUT.n5 OUT.n4 0.124059
R2197 OUT.n36 OUT.n35 0.122534
R2198 OUT.n35 OUT.n34 0.122534
R2199 OUT.n4 OUT.n2 0.121008
R2200 IBIAS.n1 IBIAS.t35 35.4861
R2201 IBIAS.n0 IBIAS.t18 31.1559
R2202 IBIAS.n11 IBIAS.t13 29.7219
R2203 IBIAS.n12 IBIAS.t26 29.7219
R2204 IBIAS.n13 IBIAS.t14 29.7219
R2205 IBIAS.n14 IBIAS.t29 29.7219
R2206 IBIAS.n17 IBIAS.t22 29.5264
R2207 IBIAS.n18 IBIAS.t31 29.5264
R2208 IBIAS.n2 IBIAS.t0 28.8746
R2209 IBIAS.n19 IBIAS.t7 28.6139
R2210 IBIAS.n17 IBIAS.t15 28.6139
R2211 IBIAS.n18 IBIAS.t24 28.6139
R2212 IBIAS.n20 IBIAS.t16 28.6139
R2213 IBIAS.n13 IBIAS.t23 28.5487
R2214 IBIAS.n14 IBIAS.t10 28.5487
R2215 IBIAS.n9 IBIAS.t30 27.4407
R2216 IBIAS.n6 IBIAS.t27 27.4407
R2217 IBIAS.n7 IBIAS.t17 27.4407
R2218 IBIAS.n8 IBIAS.t25 27.4407
R2219 IBIAS.n29 IBIAS.t4 24.0514
R2220 IBIAS.n30 IBIAS.t11 24.0514
R2221 IBIAS.n43 IBIAS.t28 24.0514
R2222 IBIAS.n23 IBIAS.t2 23.921
R2223 IBIAS.n26 IBIAS.t21 23.921
R2224 IBIAS.n29 IBIAS.t20 23.921
R2225 IBIAS.n27 IBIAS.t9 23.921
R2226 IBIAS.n30 IBIAS.t8 23.921
R2227 IBIAS.n44 IBIAS.t5 23.921
R2228 IBIAS.n43 IBIAS.t33 23.921
R2229 IBIAS.n36 IBIAS.t34 23.921
R2230 IBIAS.n39 IBIAS.t3 23.921
R2231 IBIAS.n37 IBIAS.t6 23.921
R2232 IBIAS.n25 IBIAS.t32 23.7907
R2233 IBIAS.n45 IBIAS.t19 23.7907
R2234 IBIAS.n41 IBIAS.t12 23.7907
R2235 IBIAS.n49 IBIAS.n5 10.8465
R2236 IBIAS.n18 IBIAS.n17 10.8005
R2237 IBIAS.n20 IBIAS.n19 10.8005
R2238 IBIAS.n7 IBIAS.n6 10.8005
R2239 IBIAS.n8 IBIAS.n7 10.8005
R2240 IBIAS.n12 IBIAS.n11 10.8005
R2241 IBIAS.n13 IBIAS.n12 10.8005
R2242 IBIAS.n10 IBIAS.n9 10.7505
R2243 IBIAS.n15 IBIAS.n14 10.7505
R2244 IBIAS.n37 IBIAS.n36 10.4005
R2245 IBIAS.n30 IBIAS.n29 10.4005
R2246 IBIAS.n27 IBIAS.n26 10.4005
R2247 IBIAS.n24 IBIAS.n23 10.4005
R2248 IBIAS.n44 IBIAS.n43 10.4005
R2249 IBIAS.n40 IBIAS.n39 10.4005
R2250 IBIAS.n21 IBIAS.n18 9.3005
R2251 IBIAS.n34 IBIAS.n32 7.82535
R2252 IBIAS.n34 IBIAS.n33 7.65154
R2253 IBIAS.n48 IBIAS.n22 7.45984
R2254 IBIAS.n16 IBIAS.n10 5.86108
R2255 IBIAS.n42 IBIAS.n41 5.27954
R2256 IBIAS.n28 IBIAS.n25 5.27781
R2257 IBIAS.n35 IBIAS.n34 4.0005
R2258 IBIAS.n28 IBIAS.n27 4.0005
R2259 IBIAS.n31 IBIAS.n30 4.0005
R2260 IBIAS.n42 IBIAS.n38 4.0005
R2261 IBIAS.n46 IBIAS.n45 4.0005
R2262 IBIAS.n16 IBIAS.n15 4.0005
R2263 IBIAS.n22 IBIAS.n21 4.0005
R2264 IBIAS.n4 IBIAS.n3 4.0005
R2265 IBIAS.n5 IBIAS.t1 3.97702
R2266 IBIAS.n48 IBIAS.n47 3.87374
R2267 IBIAS.n1 IBIAS.n0 3.23007
R2268 IBIAS IBIAS.n49 2.41755
R2269 IBIAS.n22 IBIAS.n16 1.75796
R2270 IBIAS.n49 IBIAS.n48 1.71832
R2271 IBIAS.n21 IBIAS.n20 1.5005
R2272 IBIAS.n35 IBIAS.n31 1.37101
R2273 IBIAS.n46 IBIAS.n42 1.27954
R2274 IBIAS.n31 IBIAS.n28 1.27435
R2275 IBIAS.n47 IBIAS.n46 1.26642
R2276 IBIAS.n4 IBIAS.n1 0.87189
R2277 IBIAS.n3 IBIAS.n2 0.8035
R2278 IBIAS.n45 IBIAS.n44 0.261214
R2279 IBIAS.n25 IBIAS.n24 0.130857
R2280 IBIAS.n41 IBIAS.n40 0.130857
R2281 IBIAS.n5 IBIAS.n4 0.0878546
R2282 IBIAS.n38 IBIAS.n37 0.0656786
R2283 IBIAS.n47 IBIAS.n35 0.0593781
R2284 IBIAS.n10 IBIAS.n8 0.0505
R2285 IBIAS.n15 IBIAS.n13 0.0505
R2286 a_n2983_n1659.n27 a_n2983_n1659.t0 23.9862
R2287 a_n2983_n1659.n42 a_n2983_n1659.t6 23.9862
R2288 a_n2983_n1659.n42 a_n2983_n1659.t2 23.9862
R2289 a_n2983_n1659.n32 a_n2983_n1659.t4 23.9862
R2290 a_n2983_n1659.n53 a_n2983_n1659.t14 23.9862
R2291 a_n2983_n1659.n53 a_n2983_n1659.t12 23.9862
R2292 a_n2983_n1659.n4 a_n2983_n1659.t10 23.9862
R2293 a_n2983_n1659.n0 a_n2983_n1659.t8 23.9862
R2294 a_n2983_n1659.n48 a_n2983_n1659.n47 6.23075
R2295 a_n2983_n1659.n47 a_n2983_n1659.n46 6.22569
R2296 a_n2983_n1659.n47 a_n2983_n1659.n25 5.8995
R2297 a_n2983_n1659.n28 a_n2983_n1659.n27 4.0005
R2298 a_n2983_n1659.n33 a_n2983_n1659.n32 4.0005
R2299 a_n2983_n1659.n43 a_n2983_n1659.n42 4.0005
R2300 a_n2983_n1659.n1 a_n2983_n1659.n0 4.0005
R2301 a_n2983_n1659.n5 a_n2983_n1659.n4 4.0005
R2302 a_n2983_n1659.n54 a_n2983_n1659.n53 4.0005
R2303 a_n2983_n1659.n19 a_n2983_n1659.n16 3.87435
R2304 a_n2983_n1659.t15 a_n2983_n1659.n8 3.79909
R2305 a_n2983_n1659.n57 a_n2983_n1659.n55 3.19242
R2306 a_n2983_n1659.n29 a_n2983_n1659.n26 3.19069
R2307 a_n2983_n1659.n31 a_n2983_n1659.n30 2.6005
R2308 a_n2983_n1659.n36 a_n2983_n1659.n35 2.6005
R2309 a_n2983_n1659.n46 a_n2983_n1659.n45 2.6005
R2310 a_n2983_n1659.n25 a_n2983_n1659.n24 2.6005
R2311 a_n2983_n1659.n22 a_n2983_n1659.n21 2.6005
R2312 a_n2983_n1659.n19 a_n2983_n1659.n18 2.6005
R2313 a_n2983_n1659.n48 a_n2983_n1659.n14 2.6005
R2314 a_n2983_n1659.n52 a_n2983_n1659.n10 2.6005
R2315 a_n2983_n1659.n50 a_n2983_n1659.n12 2.6005
R2316 a_n2983_n1659.n22 a_n2983_n1659.n19 1.27435
R2317 a_n2983_n1659.n25 a_n2983_n1659.n22 1.27435
R2318 a_n2983_n1659.n12 a_n2983_n1659.t11 0.607167
R2319 a_n2983_n1659.n12 a_n2983_n1659.n11 0.607167
R2320 a_n2983_n1659.n14 a_n2983_n1659.t9 0.607167
R2321 a_n2983_n1659.n14 a_n2983_n1659.n13 0.607167
R2322 a_n2983_n1659.n45 a_n2983_n1659.t30 0.607167
R2323 a_n2983_n1659.n45 a_n2983_n1659.t7 0.607167
R2324 a_n2983_n1659.n35 a_n2983_n1659.t16 0.607167
R2325 a_n2983_n1659.n35 a_n2983_n1659.t3 0.607167
R2326 a_n2983_n1659.n30 a_n2983_n1659.t17 0.607167
R2327 a_n2983_n1659.n30 a_n2983_n1659.t5 0.607167
R2328 a_n2983_n1659.n26 a_n2983_n1659.t19 0.607167
R2329 a_n2983_n1659.n26 a_n2983_n1659.t1 0.607167
R2330 a_n2983_n1659.n16 a_n2983_n1659.t24 0.607167
R2331 a_n2983_n1659.n16 a_n2983_n1659.n15 0.607167
R2332 a_n2983_n1659.n18 a_n2983_n1659.t26 0.607167
R2333 a_n2983_n1659.n18 a_n2983_n1659.n17 0.607167
R2334 a_n2983_n1659.n21 a_n2983_n1659.t25 0.607167
R2335 a_n2983_n1659.n21 a_n2983_n1659.n20 0.607167
R2336 a_n2983_n1659.n24 a_n2983_n1659.t18 0.607167
R2337 a_n2983_n1659.n24 a_n2983_n1659.n23 0.607167
R2338 a_n2983_n1659.n10 a_n2983_n1659.t13 0.607167
R2339 a_n2983_n1659.n10 a_n2983_n1659.n9 0.607167
R2340 a_n2983_n1659.t15 a_n2983_n1659.n57 0.607167
R2341 a_n2983_n1659.n57 a_n2983_n1659.n56 0.607167
R2342 a_n2983_n1659.n38 a_n2983_n1659.n37 0.590692
R2343 a_n2983_n1659.n39 a_n2983_n1659.n38 0.590692
R2344 a_n2983_n1659.n31 a_n2983_n1659.n29 0.590692
R2345 a_n2983_n1659.n34 a_n2983_n1659.n31 0.590692
R2346 a_n2983_n1659.n36 a_n2983_n1659.n34 0.590692
R2347 a_n2983_n1659.n44 a_n2983_n1659.n36 0.590692
R2348 a_n2983_n1659.n40 a_n2983_n1659.n39 0.590692
R2349 a_n2983_n1659.n41 a_n2983_n1659.n40 0.590692
R2350 a_n2983_n1659.n46 a_n2983_n1659.n44 0.590692
R2351 a_n2983_n1659.n49 a_n2983_n1659.n48 0.590692
R2352 a_n2983_n1659.n6 a_n2983_n1659.n3 0.590692
R2353 a_n2983_n1659.n3 a_n2983_n1659.n2 0.590692
R2354 a_n2983_n1659.n52 a_n2983_n1659.n51 0.590692
R2355 a_n2983_n1659.n51 a_n2983_n1659.n50 0.590692
R2356 a_n2983_n1659.n50 a_n2983_n1659.n49 0.590692
R2357 a_n2983_n1659.n7 a_n2983_n1659.n6 0.590692
R2358 a_n2983_n1659.n55 a_n2983_n1659.n52 0.588962
R2359 a_n2983_n1659.n8 a_n2983_n1659.n7 0.588962
R2360 a_n2983_n1659.n29 a_n2983_n1659.n28 0.183833
R2361 a_n2983_n1659.n34 a_n2983_n1659.n33 0.183833
R2362 a_n2983_n1659.n44 a_n2983_n1659.n43 0.182167
R2363 a_n2983_n1659.n55 a_n2983_n1659.n54 0.1805
R2364 a_n2983_n1659.n43 a_n2983_n1659.n41 0.178833
R2365 a_n2983_n1659.n2 a_n2983_n1659.n1 0.178833
R2366 a_n2983_n1659.n6 a_n2983_n1659.n5 0.178833
R2367 a_n3081_n3465.t1 a_n3081_n3465.t0 58.9303
R2368 a_n2937_n3465.n0 a_n2937_n3465.t1 1.21383
R2369 a_n3063_n9510.n2 a_n3063_n9510.t28 55.0195
R2370 a_n3063_n9510.n7 a_n3063_n9510.t26 55.0195
R2371 a_n3063_n9510.n14 a_n3063_n9510.t24 55.0161
R2372 a_n3063_n9510.n17 a_n3063_n9510.t30 55.0112
R2373 a_n3063_n9510.n30 a_n3063_n9510.t0 5.58454
R2374 a_n3063_n9510.n32 a_n3063_n9510.t4 5.58454
R2375 a_n3063_n9510.n25 a_n3063_n9510.n24 5.58454
R2376 a_n3063_n9510.n27 a_n3063_n9510.n26 5.58454
R2377 a_n3063_n9510.n30 a_n3063_n9510.n29 3.6965
R2378 a_n3063_n9510.n32 a_n3063_n9510.n31 3.6965
R2379 a_n3063_n9510.n25 a_n3063_n9510.t3 3.6965
R2380 a_n3063_n9510.n27 a_n3063_n9510.t5 3.6965
R2381 a_n3063_n9510.n0 a_n3063_n9510.n45 3.48152
R2382 a_n3063_n9510.n21 a_n3063_n9510.n20 3.38017
R2383 a_n3063_n9510.n34 a_n3063_n9510.n28 3.09912
R2384 a_n3063_n9510.n35 a_n3063_n9510.n34 3.04779
R2385 a_n3063_n9510.n51 a_n3063_n9510.n50 2.74437
R2386 a_n3063_n9510.n15 a_n3063_n9510.n13 2.62186
R2387 a_n3063_n9510.n16 a_n3063_n9510.n11 2.62184
R2388 a_n3063_n9510.n19 a_n3063_n9510.n18 2.62171
R2389 a_n3063_n9510.n8 a_n3063_n9510.n6 2.62053
R2390 a_n3063_n9510.n9 a_n3063_n9510.n4 2.62053
R2391 a_n3063_n9510.n53 a_n3063_n9510.n52 2.61995
R2392 a_n3063_n9510.n35 a_n3063_n9510.n23 2.60908
R2393 a_n3063_n9510.n1 a_n3063_n9510.n38 2.25075
R2394 a_n3063_n9510.n0 a_n3063_n9510.n48 2.25074
R2395 a_n3063_n9510.n34 a_n3063_n9510.n33 2.2505
R2396 a_n3063_n9510.n40 a_n3063_n9510.n39 2.24582
R2397 a_n3063_n9510.n50 a_n3063_n9510.n0 2.24292
R2398 a_n3063_n9510.t29 a_n3063_n9510.n2 2.02965
R2399 a_n3063_n9510.n48 a_n3063_n9510.n47 1.49462
R2400 a_n3063_n9510.n38 a_n3063_n9510.n37 1.4938
R2401 a_n3063_n9510.n8 a_n3063_n9510.n7 1.34068
R2402 a_n3063_n9510.n19 a_n3063_n9510.n17 1.33871
R2403 a_n3063_n9510.n15 a_n3063_n9510.n14 1.33839
R2404 a_n3063_n9510.n33 a_n3063_n9510.n30 1.06058
R2405 a_n3063_n9510.n28 a_n3063_n9510.n25 1.06058
R2406 a_n3063_n9510.n16 a_n3063_n9510.n15 0.876314
R2407 a_n3063_n9510.n9 a_n3063_n9510.n8 0.876314
R2408 a_n3063_n9510.n1 a_n3063_n9510.n35 0.869485
R2409 a_n3063_n9510.n42 a_n3063_n9510.n41 0.774919
R2410 a_n3063_n9510.n33 a_n3063_n9510.n32 0.768847
R2411 a_n3063_n9510.n28 a_n3063_n9510.n27 0.768847
R2412 a_n3063_n9510.n47 a_n3063_n9510.t11 0.5465
R2413 a_n3063_n9510.n47 a_n3063_n9510.n46 0.5465
R2414 a_n3063_n9510.n45 a_n3063_n9510.t16 0.5465
R2415 a_n3063_n9510.n45 a_n3063_n9510.n44 0.5465
R2416 a_n3063_n9510.n37 a_n3063_n9510.t9 0.5465
R2417 a_n3063_n9510.n37 a_n3063_n9510.n36 0.5465
R2418 a_n3063_n9510.n23 a_n3063_n9510.t15 0.5465
R2419 a_n3063_n9510.n23 a_n3063_n9510.n22 0.5465
R2420 a_n3063_n9510.n18 a_n3063_n9510.t8 0.5465
R2421 a_n3063_n9510.n18 a_n3063_n9510.t31 0.5465
R2422 a_n3063_n9510.n11 a_n3063_n9510.t21 0.5465
R2423 a_n3063_n9510.n11 a_n3063_n9510.n10 0.5465
R2424 a_n3063_n9510.n13 a_n3063_n9510.t25 0.5465
R2425 a_n3063_n9510.n13 a_n3063_n9510.n12 0.5465
R2426 a_n3063_n9510.n4 a_n3063_n9510.t14 0.5465
R2427 a_n3063_n9510.n4 a_n3063_n9510.n3 0.5465
R2428 a_n3063_n9510.n6 a_n3063_n9510.t27 0.5465
R2429 a_n3063_n9510.n6 a_n3063_n9510.n5 0.5465
R2430 a_n3063_n9510.t22 a_n3063_n9510.n53 0.5465
R2431 a_n3063_n9510.n53 a_n3063_n9510.t29 0.5465
R2432 a_n3063_n9510.n51 a_n3063_n9510.n9 0.422148
R2433 a_n3063_n9510.n20 a_n3063_n9510.n16 0.422093
R2434 a_n3063_n9510.n52 a_n3063_n9510.n51 0.419432
R2435 a_n3063_n9510.n20 a_n3063_n9510.n19 0.418828
R2436 a_n3063_n9510.n40 a_n3063_n9510.n21 0.0329419
R2437 a_n3063_n9510.n41 a_n3063_n9510.n40 0.0329419
R2438 a_n3063_n9510.n43 a_n3063_n9510.n42 0.0318953
R2439 a_n3063_n9510.n0 a_n3063_n9510.n49 0.0290293
R2440 a_n3063_n9510.n50 a_n3063_n9510.n43 0.0182092
R2441 a_n3063_n9510.n39 a_n3063_n9510.n1 0.0153123
R2442 a_n3086_n6147.t1 a_n3086_n6147.t0 59.8509
R2443 a_n2937_n6021.t0 a_n2937_n6021.n0 1.21383
R2444 a_n2457_n4317.t0 a_n2457_n4317.n0 1.21383
R2445 a_n2297_n4317.n0 a_n2297_n4317.t1 1.21383
R2446 a_n453_n1964.n16 a_n453_n1964.t2 34.0237
R2447 a_n453_n1964.n0 a_n453_n1964.t6 34.0237
R2448 a_n453_n1964.n16 a_n453_n1964.t0 33.763
R2449 a_n453_n1964.n0 a_n453_n1964.t4 33.763
R2450 a_n453_n1964.n13 a_n453_n1964.n4 13.4076
R2451 a_n453_n1964.n13 a_n453_n1964.n12 8.57505
R2452 a_n453_n1964.n12 a_n453_n1964.n6 6.43511
R2453 a_n453_n1964.n21 a_n453_n1964.n20 6.30469
R2454 a_n453_n1964.n25 a_n453_n1964.n21 5.43808
R2455 a_n453_n1964.n10 a_n453_n1964.n9 4.61117
R2456 a_n453_n1964.n7 a_n453_n1964.t19 4.61117
R2457 a_n453_n1964.t7 a_n453_n1964.n2 4.17956
R2458 a_n453_n1964.n18 a_n453_n1964.n16 4.0005
R2459 a_n453_n1964.n1 a_n453_n1964.n0 4.0005
R2460 a_n453_n1964.n19 a_n453_n1964.n15 3.56311
R2461 a_n453_n1964.n24 a_n453_n1964.n23 3.56311
R2462 a_n453_n1964.n10 a_n453_n1964.n8 3.20717
R2463 a_n453_n1964.n7 a_n453_n1964.t18 3.20717
R2464 a_n453_n1964.n21 a_n453_n1964.n13 3.20621
R2465 a_n453_n1964.n12 a_n453_n1964.n11 2.89327
R2466 a_n453_n1964.n20 a_n453_n1964.n14 2.6005
R2467 a_n453_n1964.n27 a_n453_n1964.n25 2.6005
R2468 a_n453_n1964.n11 a_n453_n1964.n7 1.70296
R2469 a_n453_n1964.n11 a_n453_n1964.n10 1.09816
R2470 a_n453_n1964.n20 a_n453_n1964.n19 0.972891
R2471 a_n453_n1964.n25 a_n453_n1964.n24 0.972891
R2472 a_n453_n1964.n14 a_n453_n1964.t10 0.607167
R2473 a_n453_n1964.n14 a_n453_n1964.t3 0.607167
R2474 a_n453_n1964.n15 a_n453_n1964.t17 0.607167
R2475 a_n453_n1964.n15 a_n453_n1964.t1 0.607167
R2476 a_n453_n1964.n4 a_n453_n1964.t14 0.607167
R2477 a_n453_n1964.n4 a_n453_n1964.n3 0.607167
R2478 a_n453_n1964.n6 a_n453_n1964.t12 0.607167
R2479 a_n453_n1964.n6 a_n453_n1964.n5 0.607167
R2480 a_n453_n1964.n23 a_n453_n1964.t5 0.607167
R2481 a_n453_n1964.n23 a_n453_n1964.n22 0.607167
R2482 a_n453_n1964.t7 a_n453_n1964.n27 0.607167
R2483 a_n453_n1964.n27 a_n453_n1964.n26 0.607167
R2484 a_n453_n1964.n18 a_n453_n1964.n17 0.194618
R2485 a_n453_n1964.n19 a_n453_n1964.n18 0.187559
R2486 a_n453_n1964.n2 a_n453_n1964.n1 0.184029
R2487 a_n89_n10306.n8 a_n89_n10306.t10 56.0541
R2488 a_n89_n10306.n8 a_n89_n10306.t3 55.5326
R2489 a_n89_n10306.n9 a_n89_n10306.t11 47.3201
R2490 a_n89_n10306.n10 a_n89_n10306.t4 47.3201
R2491 a_n89_n10306.n12 a_n89_n10306.t13 47.3201
R2492 a_n89_n10306.n11 a_n89_n10306.t17 47.3201
R2493 a_n89_n10306.n10 a_n89_n10306.t15 47.3201
R2494 a_n89_n10306.n12 a_n89_n10306.t7 47.3201
R2495 a_n89_n10306.n3 a_n89_n10306.t18 47.3201
R2496 a_n89_n10306.n0 a_n89_n10306.t12 47.3201
R2497 a_n89_n10306.n1 a_n89_n10306.t5 47.3201
R2498 a_n89_n10306.n1 a_n89_n10306.t9 47.3201
R2499 a_n89_n10306.n2 a_n89_n10306.t6 47.3201
R2500 a_n89_n10306.n2 a_n89_n10306.t8 47.3201
R2501 a_n89_n10306.n3 a_n89_n10306.t14 47.3201
R2502 a_n89_n10306.n11 a_n89_n10306.t16 47.3201
R2503 a_n89_n10306.n16 a_n89_n10306.t0 26.8782
R2504 a_n89_n10306.n1 a_n89_n10306.n0 18.8981
R2505 a_n89_n10306.n3 a_n89_n10306.n2 18.8981
R2506 a_n89_n10306.n8 a_n89_n10306.n7 18.8981
R2507 a_n89_n10306.n6 a_n89_n10306.n5 18.8981
R2508 a_n89_n10306.n10 a_n89_n10306.n9 18.8981
R2509 a_n89_n10306.n12 a_n89_n10306.n11 18.8981
R2510 a_n89_n10306.n14 a_n89_n10306.n8 17.4226
R2511 a_n89_n10306.n7 a_n89_n10306.n6 9.41985
R2512 a_n89_n10306.n14 a_n89_n10306.n13 7.65668
R2513 a_n89_n10306.n15 a_n89_n10306.n4 6.6153
R2514 a_n89_n10306.n17 a_n89_n10306.n15 6.60167
R2515 a_n89_n10306.n18 a_n89_n10306.n17 6.4841
R2516 a_n89_n10306.n13 a_n89_n10306.n10 5.12227
R2517 a_n89_n10306.n4 a_n89_n10306.n3 4.82792
R2518 a_n89_n10306.n4 a_n89_n10306.n1 4.59244
R2519 a_n89_n10306.n16 a_n89_n10306.t1 4.47258
R2520 a_n89_n10306.n13 a_n89_n10306.n12 4.29808
R2521 a_n89_n10306.n15 a_n89_n10306.n14 1.0215
R2522 a_n89_n10306.n17 a_n89_n10306.n16 0.324731
R2523 a_n2937_n4317.n0 a_n2937_n4317.t1 1.21383
R2524 a_n2777_n4317.n0 a_n2777_n4317.t1 1.21383
R2525 a_n168_n4318.n2 a_n168_n4318.t6 70.1735
R2526 a_n168_n4318.n8 a_n168_n4318.t5 45.8988
R2527 a_n168_n4318.n4 a_n168_n4318.t8 44.8434
R2528 a_n168_n4318.n5 a_n168_n4318.t10 44.8434
R2529 a_n168_n4318.n2 a_n168_n4318.t9 44.8434
R2530 a_n168_n4318.n6 a_n168_n4318.t3 44.8434
R2531 a_n168_n4318.n3 a_n168_n4318.t11 44.8434
R2532 a_n168_n4318.n7 a_n168_n4318.t7 44.8434
R2533 a_n168_n4318.t5 a_n168_n4318.n7 44.8434
R2534 a_n168_n4318.n9 a_n168_n4318.n8 33.6473
R2535 a_n168_n4318.n8 a_n168_n4318.n3 24.2752
R2536 a_n168_n4318.n5 a_n168_n4318.n4 22.8527
R2537 a_n168_n4318.n7 a_n168_n4318.n6 22.8527
R2538 a_n168_n4318.n1 a_n168_n4318.t0 19.6434
R2539 a_n168_n4318.n3 a_n168_n4318.n2 14.0728
R2540 a_n168_n4318.n6 a_n168_n4318.n5 12.6962
R2541 a_n168_n4318.t2 a_n168_n4318.n9 6.33333
R2542 a_n168_n4318.n1 a_n168_n4318.n0 4.95
R2543 a_n168_n4318.n9 a_n168_n4318.n1 0.541581
R2544 a_n453_n3002.n25 a_n453_n3002.t14 33.7219
R2545 a_n453_n3002.n16 a_n453_n3002.t16 33.5264
R2546 a_n453_n3002.n2 a_n453_n3002.t18 30.5282
R2547 a_n453_n3002.n5 a_n453_n3002.t12 30.3978
R2548 a_n453_n3002.n13 a_n453_n3002.n12 7.77975
R2549 a_n453_n3002.n7 a_n453_n3002.n6 5.8123
R2550 a_n453_n3002.n26 a_n453_n3002.n24 5.73119
R2551 a_n453_n3002.n7 a_n453_n3002.n3 5.04829
R2552 a_n453_n3002.n24 a_n453_n3002.n13 4.82813
R2553 a_n453_n3002.n13 a_n453_n3002.n7 4.79057
R2554 a_n453_n3002.n23 a_n453_n3002.n22 4.49732
R2555 a_n453_n3002.n22 a_n453_n3002.n21 4.0045
R2556 a_n453_n3002.n12 a_n453_n3002.n9 3.56623
R2557 a_n453_n3002.n12 a_n453_n3002.n11 3.548
R2558 a_n453_n3002.n27 a_n453_n3002.n26 3.40873
R2559 a_n453_n3002.n17 a_n453_n3002.n15 3.40267
R2560 a_n453_n3002.n3 a_n453_n3002.n1 3.3205
R2561 a_n453_n3002.n6 a_n453_n3002.n4 3.31659
R2562 a_n453_n3002.n23 a_n453_n3002.n17 2.80473
R2563 a_n453_n3002.n22 a_n453_n3002.n19 2.6005
R2564 a_n453_n3002.n24 a_n453_n3002.n23 2.2505
R2565 a_n453_n3002.n15 a_n453_n3002.t17 0.607167
R2566 a_n453_n3002.n15 a_n453_n3002.n14 0.607167
R2567 a_n453_n3002.n21 a_n453_n3002.t1 0.607167
R2568 a_n453_n3002.n21 a_n453_n3002.n20 0.607167
R2569 a_n453_n3002.n19 a_n453_n3002.t2 0.607167
R2570 a_n453_n3002.n19 a_n453_n3002.n18 0.607167
R2571 a_n453_n3002.n9 a_n453_n3002.t7 0.607167
R2572 a_n453_n3002.n9 a_n453_n3002.n8 0.607167
R2573 a_n453_n3002.n11 a_n453_n3002.t4 0.607167
R2574 a_n453_n3002.n11 a_n453_n3002.n10 0.607167
R2575 a_n453_n3002.n4 a_n453_n3002.t5 0.607167
R2576 a_n453_n3002.n4 a_n453_n3002.t13 0.607167
R2577 a_n453_n3002.n1 a_n453_n3002.t19 0.607167
R2578 a_n453_n3002.n1 a_n453_n3002.n0 0.607167
R2579 a_n453_n3002.n27 a_n453_n3002.t11 0.607167
R2580 a_n453_n3002.t15 a_n453_n3002.n27 0.607167
R2581 a_n453_n3002.n6 a_n453_n3002.n5 0.1265
R2582 a_n453_n3002.n3 a_n453_n3002.n2 0.121232
R2583 a_n453_n3002.n26 a_n453_n3002.n25 0.109786
R2584 a_n453_n3002.n17 a_n453_n3002.n16 0.109337
R2585 a_n1977_n4317.t0 a_n1977_n4317.n0 1.21383
R2586 a_n1817_n4317.t0 a_n1817_n4317.n0 1.21383
R2587 a_n1817_n3465.t0 a_n1817_n3465.n0 1.21383
R2588 a_n1657_n3465.t0 a_n1657_n3465.n0 1.21383
R2589 a_n1817_n6021.n0 a_n1817_n6021.t1 1.21383
R2590 a_n1657_n6021.n0 a_n1657_n6021.t1 1.21383
R2591 a_n3083_n5296.t1 a_n3083_n5296.t0 59.7744
R2592 a_n2937_n5169.t0 a_n2937_n5169.n0 1.21383
R2593 a_n2137_n4317.n0 a_n2137_n4317.t1 1.21383
R2594 a_n2617_n4317.t0 a_n2617_n4317.n0 1.21383
R2595 a_n2137_n6021.t0 a_n2137_n6021.n0 1.21383
R2596 a_n1977_n6021.n0 a_n1977_n6021.t1 1.21383
R2597 a_n2137_n3465.n0 a_n2137_n3465.t1 1.21383
R2598 a_n1977_n3465.n0 a_n1977_n3465.t1 1.21383
R2599 a_n2617_n6021.t0 a_n2617_n6021.n0 1.21383
R2600 a_n2457_n6021.n0 a_n2457_n6021.t1 1.21383
R2601 a_n2617_n3465.t0 a_n2617_n3465.n0 1.21383
R2602 a_n2457_n3465.t0 a_n2457_n3465.n0 1.21383
R2603 a_n1553_n3596.n0 a_n1553_n3596.t0 59.4423
R2604 a_n1553_n6152.n0 a_n1553_n6152.t0 59.4488
R2605 a_n1817_n5169.t0 a_n1817_n5169.n0 1.21383
R2606 a_n1657_n5169.t0 a_n1657_n5169.n0 1.21383
R2607 a_n3086_n4453.t1 a_n3086_n4453.t0 59.0853
R2608 a_n2137_n5169.n0 a_n2137_n5169.t1 1.21383
R2609 a_n1977_n5169.n0 a_n1977_n5169.t1 1.21383
R2610 a_n2297_n3465.t0 a_n2297_n3465.n0 1.21383
R2611 a_n2297_n6021.t0 a_n2297_n6021.n0 1.21383
R2612 a_n2457_n5169.t0 a_n2457_n5169.n0 1.21383
R2613 a_n2777_n3465.n0 a_n2777_n3465.t1 1.21383
R2614 a_n2777_n6021.t0 a_n2777_n6021.n0 1.21383
R2615 a_n1553_n5305.n0 a_n1553_n5305.t0 59.0914
R2616 a_n1657_n4317.n0 a_n1657_n4317.t1 1.21383
R2617 a_3734_n7493.n0 a_3734_n7493.t3 48.7904
R2618 a_3734_n7493.n0 a_3734_n7493.t1 15.8389
R2619 a_3734_n7493.n1 a_3734_n7493.n0 10.7971
R2620 a_3734_n7493.n2 a_3734_n7493.n1 6.99401
R2621 a_3734_n7493.n1 a_3734_n7493.t2 4.51305
R2622 a_n2297_n5169.n0 a_n2297_n5169.t1 1.21383
R2623 a_n1553_n4448.n0 a_n1553_n4448.t0 59.4488
R2624 VINP VINP.n0 2.26502
R2625 VINN VINN.n0 2.26502
C0 VDD a_n2849_n6153# 1.21f
C1 VDD OUT 2.23f
C2 a_n2845_n5323# VINN 0.0367f
C3 m1_n3664_n2831# VINN 2.76e-20
C4 a_n2845_n5323# a_n2688_n4484# 0.192f
C5 m1_n3668_n2597# VINN 0.0295f
C6 a_n2845_n3640# VDD 1.1f
C7 OUT a_n2849_n6153# 4.07e-22
C8 IBIAS VINN 0.017f
C9 VDD VINP 0.216f
C10 a_n2849_n2813# VDD 1.38f
C11 VINP a_n2849_n6153# 0.0225f
C12 VINN a_n2688_n4484# 0.0579f
C13 a_n2845_n3640# VINP 0.0635f
C14 a_n2849_n2813# a_n2845_n3640# 0.213f
C15 a_n2849_n2813# VINP 0.0315f
C16 a_n2845_n5323# VDD 1.09f
C17 m1_n3664_n2831# VDD 0.0221f
C18 m1_n3668_n2597# VDD 0.00962f
C19 VDD IBIAS 17.6f
C20 a_n2845_n5323# a_n2849_n6153# 0.213f
C21 a_n2845_n5323# OUT 1.33e-20
C22 VDD VINN 0.474f
C23 IBIAS OUT 0.00148f
C24 a_n2845_n5323# a_n2845_n3640# 0.0177f
C25 VDD a_n2688_n4484# 0.869f
C26 a_n2845_n5323# VINP 0.0602f
C27 m1_n3664_n2831# VINP 0.0266f
C28 a_n2849_n2813# m1_n3664_n2831# 1.24e-19
C29 a_n2845_n3640# IBIAS 0.00116f
C30 VINN a_n2849_n6153# 0.0472f
C31 OUT VINN 0.006f
C32 a_n2849_n6153# a_n2688_n4484# 2.58e-22
C33 OUT a_n2688_n4484# 1.75e-20
C34 a_n2849_n2813# IBIAS 0.00118f
C35 a_n2845_n3640# VINN 0.0471f
C36 a_n2845_n3640# a_n2688_n4484# 0.192f
C37 VINN VINP 0.297f
C38 VINP a_n2688_n4484# 0.0181f
C39 a_n2849_n2813# VINN 0.0734f
C40 a_n2849_n2813# a_n2688_n4484# 5.88e-22
C41 m1_n3668_n2597# m1_n3664_n2831# 0.0478f
.ends

