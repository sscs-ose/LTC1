magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -3726 -2128 3726 2128
<< nwell >>
rect -1726 -128 1726 128
<< nsubdiff >>
rect -1643 23 1643 45
rect -1643 -23 -1621 23
rect 1621 -23 1643 23
rect -1643 -45 1643 -23
<< nsubdiffcont >>
rect -1621 -23 1621 23
<< metal1 >>
rect -1632 23 1632 34
rect -1632 -23 -1621 23
rect 1621 -23 1632 23
rect -1632 -34 1632 -23
<< end >>
