magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1100 -1073 1100 1073
<< metal1 >>
rect -100 67 100 73
rect -100 41 -94 67
rect -68 41 -40 67
rect -14 41 14 67
rect 40 41 68 67
rect 94 41 100 67
rect -100 13 100 41
rect -100 -13 -94 13
rect -68 -13 -40 13
rect -14 -13 14 13
rect 40 -13 68 13
rect 94 -13 100 13
rect -100 -41 100 -13
rect -100 -67 -94 -41
rect -68 -67 -40 -41
rect -14 -67 14 -41
rect 40 -67 68 -41
rect 94 -67 100 -41
rect -100 -73 100 -67
<< via1 >>
rect -94 41 -68 67
rect -40 41 -14 67
rect 14 41 40 67
rect 68 41 94 67
rect -94 -13 -68 13
rect -40 -13 -14 13
rect 14 -13 40 13
rect 68 -13 94 13
rect -94 -67 -68 -41
rect -40 -67 -14 -41
rect 14 -67 40 -41
rect 68 -67 94 -41
<< metal2 >>
rect -100 67 100 73
rect -100 41 -94 67
rect -68 41 -40 67
rect -14 41 14 67
rect 40 41 68 67
rect 94 41 100 67
rect -100 13 100 41
rect -100 -13 -94 13
rect -68 -13 -40 13
rect -14 -13 14 13
rect 40 -13 68 13
rect 94 -13 100 13
rect -100 -41 100 -13
rect -100 -67 -94 -41
rect -68 -67 -40 -41
rect -14 -67 14 -41
rect 40 -67 68 -41
rect 94 -67 100 -41
rect -100 -73 100 -67
<< end >>
